// Benchmark "top" written by ABC on Wed May 27 23:35:13 2020

module rf_multiplier ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , a16 ,
    a17 , a18 , a19 , a20 , a21 , a22 , a23 , a24 ,
    a25 , a26 , a27 , a28 , a29 , a30 , a31 , a32 ,
    a33 , a34 , a35 , a36 , a37 , a38 , a39 , a40 ,
    a41 , a42 , a43 , a44 , a45 , a46 , a47 , a48 ,
    a49 , a50 , a51 , a52 , a53 , a54 , a55 , a56 ,
    a57 , a58 , a59 , a60 , a61 , a62 , a63 , b0 ,
    b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 , b9 ,
    b10 , b11 , b12 , b13 , b14 , b15 , b16 , b17 ,
    b18 , b19 , b20 , b21 , b22 , b23 , b24 , b25 ,
    b26 , b27 , b28 , b29 , b30 , b31 , b32 , b33 ,
    b34 , b35 , b36 , b37 , b38 , b39 , b40 , b41 ,
    b42 , b43 , b44 , b45 , b46 , b47 , b48 , b49 ,
    b50 , b51 , b52 , b53 , b54 , b55 , b56 , b57 ,
    b58 , b59 , b60 , b61 , b62 , b63 ,
    f0 , f1 , f2 , f3 , f4 , f5 , f6 , f7 , f8 ,
    f9 , f10 , f11 , f12 , f13 , f14 , f15 , f16 ,
    f17 , f18 , f19 , f20 , f21 , f22 , f23 , f24 ,
    f25 , f26 , f27 , f28 , f29 , f30 , f31 , f32 ,
    f33 , f34 , f35 , f36 , f37 , f38 , f39 , f40 ,
    f41 , f42 , f43 , f44 , f45 , f46 , f47 , f48 ,
    f49 , f50 , f51 , f52 , f53 , f54 , f55 , f56 ,
    f57 , f58 , f59 , f60 , f61 , f62 , f63 , f64 ,
    f65 , f66 , f67 , f68 , f69 , f70 , f71 , f72 ,
    f73 , f74 , f75 , f76 , f77 , f78 , f79 , f80 ,
    f81 , f82 , f83 , f84 , f85 , f86 , f87 , f88 ,
    f89 , f90 , f91 , f92 , f93 , f94 , f95 , f96 ,
    f97 , f98 , f99 , f100 , f101 , f102 , f103 ,
    f104 , f105 , f106 , f107 , f108 , f109 , f110 ,
    f111 , f112 , f113 , f114 , f115 , f116 , f117 ,
    f118 , f119 , f120 , f121 , f122 , f123 , f124 ,
    f125 , f126 , f127   );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    a16 , a17 , a18 , a19 , a20 , a21 , a22 , a23 ,
    a24 , a25 , a26 , a27 , a28 , a29 , a30 , a31 ,
    a32 , a33 , a34 , a35 , a36 , a37 , a38 , a39 ,
    a40 , a41 , a42 , a43 , a44 , a45 , a46 , a47 ,
    a48 , a49 , a50 , a51 , a52 , a53 , a54 , a55 ,
    a56 , a57 , a58 , a59 , a60 , a61 , a62 , a63 ,
    b0 , b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 ,
    b9 , b10 , b11 , b12 , b13 , b14 , b15 , b16 ,
    b17 , b18 , b19 , b20 , b21 , b22 , b23 , b24 ,
    b25 , b26 , b27 , b28 , b29 , b30 , b31 , b32 ,
    b33 , b34 , b35 , b36 , b37 , b38 , b39 , b40 ,
    b41 , b42 , b43 , b44 , b45 , b46 , b47 , b48 ,
    b49 , b50 , b51 , b52 , b53 , b54 , b55 , b56 ,
    b57 , b58 , b59 , b60 , b61 , b62 , b63 ;
  output f0 , f1 , f2 , f3 , f4 , f5 , f6 , f7 ,
    f8 , f9 , f10 , f11 , f12 , f13 , f14 , f15 ,
    f16 , f17 , f18 , f19 , f20 , f21 , f22 , f23 ,
    f24 , f25 , f26 , f27 , f28 , f29 , f30 , f31 ,
    f32 , f33 , f34 , f35 , f36 , f37 , f38 , f39 ,
    f40 , f41 , f42 , f43 , f44 , f45 , f46 , f47 ,
    f48 , f49 , f50 , f51 , f52 , f53 , f54 , f55 ,
    f56 , f57 , f58 , f59 , f60 , f61 , f62 , f63 ,
    f64 , f65 , f66 , f67 , f68 , f69 , f70 , f71 ,
    f72 , f73 , f74 , f75 , f76 , f77 , f78 , f79 ,
    f80 , f81 , f82 , f83 , f84 , f85 , f86 , f87 ,
    f88 , f89 , f90 , f91 , f92 , f93 , f94 , f95 ,
    f96 , f97 , f98 , f99 , f100 , f101 , f102 ,
    f103 , f104 , f105 , f106 , f107 , f108 , f109 ,
    f110 , f111 , f112 , f113 , f114 , f115 , f116 ,
    f117 , f118 , f119 , f120 , f121 , f122 , f123 ,
    f124 , f125 , f126 , f127 ;
  wire n256, n257, n258, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n636, n637,
    n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
    n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
    n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
    n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
    n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
    n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
    n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
    n3570, n3571, n3572, n3573, n3574, n3575, n3577, n3578, n3579, n3580,
    n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
    n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
    n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
    n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
    n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
    n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
    n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
    n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
    n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
    n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
    n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
    n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
    n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
    n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
    n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
    n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4349, n4350, n4351, n4352, n4353, n4354,
    n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
    n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
    n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
    n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
    n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
    n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
    n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
    n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
    n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
    n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
    n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
    n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
    n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
    n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
    n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
    n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
    n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
    n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
    n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
    n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
    n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
    n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
    n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
    n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
    n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
    n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
    n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
    n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
    n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
    n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
    n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
    n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
    n5640, n5641, n5642, n5643, n5644, n5645, n5647, n5648, n5649, n5650,
    n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
    n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
    n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
    n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
    n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
    n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
    n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
    n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
    n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
    n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
    n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
    n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
    n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
    n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5871,
    n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
    n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
    n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
    n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
    n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
    n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
    n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
    n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
    n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
    n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
    n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
    n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
    n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
    n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
    n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
    n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
    n6112, n6113, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
    n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
    n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
    n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
    n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
    n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
    n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
    n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
    n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
    n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
    n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
    n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
    n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
    n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
    n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
    n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
    n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
    n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
    n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
    n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
    n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
    n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
    n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
    n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
    n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
    n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
    n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
    n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
    n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
    n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
    n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
    n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
    n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
    n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
    n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
    n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
    n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
    n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
    n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
    n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
    n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
    n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
    n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
    n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
    n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
    n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
    n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
    n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
    n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
    n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
    n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
    n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
    n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
    n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
    n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
    n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
    n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
    n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
    n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
    n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
    n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
    n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
    n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
    n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
    n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
    n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
    n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
    n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
    n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
    n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
    n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
    n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
    n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
    n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
    n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
    n7668, n7669, n7670, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
    n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
    n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
    n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
    n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
    n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
    n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
    n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
    n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7949,
    n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
    n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
    n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
    n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
    n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
    n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
    n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
    n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
    n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
    n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
    n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
    n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
    n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
    n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
    n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
    n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
    n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
    n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
    n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
    n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
    n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
    n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
    n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
    n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
    n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8506, n8507, n8508, n8509, n8510, n8511,
    n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
    n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
    n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
    n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
    n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
    n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
    n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
    n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
    n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
    n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
    n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
    n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
    n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
    n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
    n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
    n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
    n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
    n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
    n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
    n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
    n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
    n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
    n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
    n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
    n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
    n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
    n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
    n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
    n8792, n8793, n8794, n8795, n8796, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
    n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
    n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
    n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
    n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
    n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
    n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
    n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
    n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
    n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
    n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
    n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
    n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
    n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
    n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
    n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
    n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
    n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
    n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
    n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
    n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
    n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
    n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
    n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
    n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
    n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
    n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
    n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
    n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
    n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
    n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
    n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
    n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
    n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
    n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
    n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
    n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
    n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
    n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
    n9394, n9395, n9396, n9397, n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
    n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
    n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
    n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
    n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
    n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
    n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
    n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
    n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
    n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
    n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
    n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
    n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
    n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
    n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
    n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
    n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
    n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
    n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
    n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
    n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9711, n9712, n9713, n9714, n9715,
    n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
    n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
    n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
    n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
    n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
    n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
    n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
    n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
    n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
    n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
    n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
    n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
    n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
    n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
    n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
    n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
    n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
    n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
    n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
    n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
    n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
    n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
    n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
    n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
    n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
    n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
    n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
    n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
    n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
    n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
    n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
    n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
    n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
    n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
    n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
    n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
    n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
    n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
    n10321, n10322, n10323, n10324, n10325, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
    n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
    n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
    n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
    n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
    n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
    n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
    n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
    n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
    n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
    n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
    n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
    n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
    n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
    n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
    n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
    n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
    n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
    n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10655,
    n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
    n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
    n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
    n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
    n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
    n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
    n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
    n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
    n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
    n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
    n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
    n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
    n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
    n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
    n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
    n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
    n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
    n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
    n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
    n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
    n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
    n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
    n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
    n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
    n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
    n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
    n11107, n11108, n11109, n11110, n11111, n11112, n11116, n11117, n11118,
    n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
    n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
    n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
    n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
    n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
    n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
    n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
    n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
    n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
    n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
    n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
    n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
    n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
    n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
    n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
    n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
    n11281, n11282, n11283, n11284, n11285, n11286, n11288, n11289, n11290,
    n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
    n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
    n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
    n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
    n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
    n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
    n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
    n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
    n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
    n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
    n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
    n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
    n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
    n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
    n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
    n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
    n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
    n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
    n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
    n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
    n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
    n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
    n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
    n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
    n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
    n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
    n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
    n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
    n11597, n11598, n11599, n11600, n11601, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
    n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
    n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
    n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
    n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
    n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
    n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
    n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
    n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
    n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
    n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
    n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
    n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
    n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
    n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
    n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
    n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
    n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
    n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
    n11904, n11905, n11906, n11907, n11908, n11910, n11911, n11912, n11913,
    n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
    n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
    n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
    n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
    n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
    n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
    n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
    n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
    n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
    n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
    n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
    n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
    n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
    n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
    n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
    n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
    n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
    n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
    n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
    n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
    n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
    n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
    n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
    n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
    n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
    n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
    n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
    n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
    n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
    n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
    n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
    n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
    n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
    n12211, n12212, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
    n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
    n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
    n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
    n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
    n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
    n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
    n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
    n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
    n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
    n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
    n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
    n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
    n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
    n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
    n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
    n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
    n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
    n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
    n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
    n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
    n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
    n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
    n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
    n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
    n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
    n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
    n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
    n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
    n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
    n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12526, n12527,
    n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
    n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
    n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
    n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
    n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12831, n12832, n12833, n12834,
    n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
    n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
    n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
    n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
    n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
    n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
    n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
    n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
    n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
    n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
    n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
    n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
    n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
    n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
    n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
    n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
    n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
    n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
    n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
    n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
    n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
    n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
    n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
    n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
    n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
    n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
    n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
    n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
    n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
    n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
    n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
    n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
    n13123, n13124, n13125, n13126, n13127, n13128, n13130, n13131, n13132,
    n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
    n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
    n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
    n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
    n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
    n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
    n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
    n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
    n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
    n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
    n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
    n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
    n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
    n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
    n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
    n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
    n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
    n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
    n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
    n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
    n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
    n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
    n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
    n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
    n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
    n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
    n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
    n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
    n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
    n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
    n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
    n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
    n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
    n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
    n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
    n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
    n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
    n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
    n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
    n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
    n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
    n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
    n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
    n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
    n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
    n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
    n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
    n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
    n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
    n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
    n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
    n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
    n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
    n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13719,
    n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
    n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
    n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
    n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
    n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
    n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
    n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
    n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
    n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
    n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
    n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
    n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
    n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
    n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
    n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
    n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
    n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
    n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
    n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
    n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
    n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
    n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
    n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
    n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
    n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
    n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
    n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
    n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
    n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
    n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
    n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13998, n13999,
    n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
    n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
    n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
    n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
    n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
    n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
    n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
    n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
    n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
    n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
    n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
    n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
    n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
    n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
    n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
    n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
    n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
    n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
    n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
    n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
    n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
    n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
    n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
    n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
    n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
    n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
    n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
    n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
    n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
    n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
    n14270, n14271, n14272, n14273, n14275, n14276, n14277, n14278, n14279,
    n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
    n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
    n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
    n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
    n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
    n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
    n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
    n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
    n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
    n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
    n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
    n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
    n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
    n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
    n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
    n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
    n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
    n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
    n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
    n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
    n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
    n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14546, n14547, n14548, n14549, n14550,
    n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
    n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
    n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
    n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
    n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
    n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
    n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
    n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
    n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
    n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
    n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
    n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
    n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
    n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
    n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
    n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
    n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
    n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
    n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
    n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
    n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
    n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
    n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
    n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
    n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
    n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
    n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
    n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
    n14803, n14804, n14805, n14806, n14807, n14809, n14810, n14811, n14812,
    n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
    n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
    n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
    n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
    n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
    n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
    n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
    n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
    n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
    n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
    n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
    n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
    n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
    n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
    n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
    n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
    n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
    n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
    n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
    n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
    n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
    n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
    n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
    n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
    n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
    n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
    n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
    n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
    n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
    n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
    n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
    n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
    n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
    n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
    n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
    n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
    n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
    n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
    n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
    n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
    n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
    n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15332, n15333, n15334, n15335, n15336,
    n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
    n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
    n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
    n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
    n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
    n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
    n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
    n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
    n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
    n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
    n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
    n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
    n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
    n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
    n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
    n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
    n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
    n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
    n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
    n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
    n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
    n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
    n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
    n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
    n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
    n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
    n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
    n15580, n15581, n15582, n15583, n15584, n15586, n15587, n15588, n15589,
    n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
    n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
    n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
    n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
    n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
    n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
    n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
    n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
    n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
    n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
    n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
    n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
    n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
    n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
    n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
    n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
    n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
    n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
    n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
    n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
    n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
    n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
    n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
    n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
    n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
    n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
    n15833, n15834, n15835, n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
    n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
    n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
    n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
    n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
    n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
    n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
    n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
    n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
    n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
    n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
    n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
    n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
    n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
    n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
    n16068, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
    n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
    n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
    n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
    n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
    n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
    n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
    n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
    n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
    n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
    n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
    n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
    n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
    n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
    n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
    n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
    n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
    n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
    n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
    n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
    n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
    n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
    n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
    n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
    n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
    n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
    n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16311, n16312,
    n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
    n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
    n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
    n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
    n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
    n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
    n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
    n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
    n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
    n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
    n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
    n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
    n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
    n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
    n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
    n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
    n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
    n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
    n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
    n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
    n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
    n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
    n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
    n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
    n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
    n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
    n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
    n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
    n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
    n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
    n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
    n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
    n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
    n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
    n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
    n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
    n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
    n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
    n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
    n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
    n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
    n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
    n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
    n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
    n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
    n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
    n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
    n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
    n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
    n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
    n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
    n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
    n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
    n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
    n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
    n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
    n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
    n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
    n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
    n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
    n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
    n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
    n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16998, n16999,
    n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
    n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
    n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
    n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
    n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
    n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
    n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
    n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
    n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
    n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
    n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
    n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
    n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
    n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
    n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
    n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
    n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
    n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
    n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
    n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
    n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
    n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
    n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
    n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
    n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17224, n17225,
    n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
    n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
    n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
    n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
    n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
    n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
    n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
    n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
    n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
    n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
    n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
    n17424, n17425, n17426, n17427, n17428, n17430, n17431, n17432, n17433,
    n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
    n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
    n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
    n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
    n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
    n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
    n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
    n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
    n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
    n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
    n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
    n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
    n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
    n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
    n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
    n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
    n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
    n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
    n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
    n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
    n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
    n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
    n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17640, n17641,
    n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
    n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
    n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
    n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
    n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
    n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
    n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
    n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
    n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
    n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
    n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
    n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
    n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
    n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
    n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
    n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
    n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
    n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
    n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
    n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
    n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
    n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
    n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
    n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
    n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
    n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
    n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
    n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
    n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
    n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
    n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
    n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
    n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
    n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
    n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
    n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
    n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
    n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
    n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
    n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
    n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
    n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
    n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
    n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
    n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
    n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
    n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
    n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
    n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
    n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
    n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
    n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
    n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
    n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
    n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
    n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
    n18229, n18230, n18231, n18232, n18233, n18234, n18236, n18237, n18238,
    n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
    n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
    n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
    n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
    n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
    n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
    n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
    n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
    n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
    n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
    n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
    n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
    n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
    n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
    n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
    n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
    n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
    n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18427, n18428,
    n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
    n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
    n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
    n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
    n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
    n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
    n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
    n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
    n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
    n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
    n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
    n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
    n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
    n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
    n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
    n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
    n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
    n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
    n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18599, n18600,
    n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
    n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
    n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
    n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
    n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
    n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
    n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
    n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
    n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
    n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
    n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
    n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
    n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
    n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
    n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
    n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
    n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
    n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
    n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
    n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18780, n18781,
    n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
    n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
    n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
    n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
    n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
    n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
    n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
    n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
    n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
    n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
    n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
    n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
    n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
    n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
    n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
    n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
    n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
    n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
    n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
    n18953, n18954, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
    n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
    n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
    n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
    n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
    n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
    n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
    n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
    n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
    n19116, n19117, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
    n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
    n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
    n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
    n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
    n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
    n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
    n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
    n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
    n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
    n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
    n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
    n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
    n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
    n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
    n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
    n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
    n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
    n19279, n19280, n19281, n19282, n19284, n19285, n19286, n19287, n19288,
    n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
    n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
    n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
    n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
    n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
    n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
    n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
    n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
    n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
    n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
    n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
    n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
    n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
    n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
    n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
    n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
    n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
    n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
    n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
    n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
    n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
    n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
    n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
    n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19596,
    n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
    n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
    n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
    n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
    n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
    n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
    n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
    n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
    n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
    n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
    n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
    n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
    n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
    n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
    n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
    n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
    n19741, n19742, n19743, n19745, n19746, n19747, n19748, n19749, n19750,
    n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
    n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
    n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
    n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
    n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
    n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
    n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
    n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
    n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
    n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
    n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
    n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
    n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
    n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
    n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
    n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
    n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976,
    n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
    n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
    n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
    n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
    n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
    n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
    n20031, n20032, n20034, n20035, n20036, n20037, n20038, n20039, n20040,
    n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
    n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
    n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
    n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
    n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
    n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
    n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
    n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
    n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
    n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
    n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
    n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
    n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
    n20158, n20159, n20160, n20161, n20162, n20164, n20165, n20166, n20167,
    n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176,
    n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
    n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
    n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
    n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
    n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
    n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
    n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
    n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248,
    n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
    n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
    n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
    n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
    n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
    n20294, n20295, n20296, n20298, n20299, n20300, n20301, n20302, n20303,
    n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
    n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
    n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
    n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
    n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384,
    n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
    n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
    n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
    n20412, n20413, n20414, n20415, n20416, n20418, n20419, n20420, n20421,
    n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
    n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
    n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
    n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
    n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
    n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
    n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
    n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
    n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
    n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
    n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520,
    n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
    n20530, n20531, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
    n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
    n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
    n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584,
    n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
    n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
    n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
    n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
    n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
    n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
    n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
    n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
    n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
    n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
    n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
    n20748, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
    n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
    n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
    n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784,
    n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
    n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
    n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
    n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
    n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
    n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
    n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20847, n20848,
    n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
    n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
    n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
    n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
    n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
    n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
    n20939, n20940, n20941, n20942, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
    n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
    n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
    n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
    n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21030,
    n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
    n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048,
    n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
    n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
    n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
    n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
    n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
    n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
    n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21112,
    n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
    n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
    n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
    n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
    n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
    n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
    n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175,
    n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184,
    n21185, n21186, n21187, n21188, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
    n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
    n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239,
    n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
    n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
    n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
    n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
    n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303,
    n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312,
    n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
    n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
    n21331, n21332, n21333, n21334, n21335, n21337, n21338, n21339, n21340,
    n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
    n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
    n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367,
    n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376,
    n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
    n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
    n21395, n21396, n21397, n21398, n21399, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
    n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
    n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
    n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21464, n21465, n21466, n21467, n21468,
    n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
    n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486,
    n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
    n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504,
    n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
    n21514, n21515, n21516, n21518, n21519, n21520, n21521, n21522, n21523,
    n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
    n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
    n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
    n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
    n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21568, n21569,
    n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
    n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
    n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
    n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
    n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21615,
    n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624,
    n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
    n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
    n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
    n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
    n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670,
    n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
    n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21688, n21689,
    n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
    n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
    n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21717,
    n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
    n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
    n21736, n21737, n21738, n21739, n21741, n21742, n21743, n21744, n21745,
    n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
    n21755, n21756, n21757, n21758, n21760, n21761, n21762, n21763, n21764,
    n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773,
    n21774, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
    n21784, n21785;
  jnot g00000(.din(a0 ), .dout(n256));
  jnot g00001(.din(b0 ), .dout(n257));
  jor  g00002(.dina(n257), .dinb(n256), .dout(n258));
  jnot g00003(.din(n258), .dout(f0 ));
  jnot g00004(.din(a2 ), .dout(n260));
  jor  g00005(.dina(n258), .dinb(n260), .dout(n261));
  jnot g00006(.din(a1 ), .dout(n262));
  jxor g00007(.dina(a2 ), .dinb(n262), .dout(n263));
  jor  g00008(.dina(n263), .dinb(n256), .dout(n264));
  jxor g00009(.dina(b1 ), .dinb(n257), .dout(n265));
  jor  g00010(.dina(n265), .dinb(n264), .dout(n266));
  jnot g00011(.din(b1 ), .dout(n267));
  jxor g00012(.dina(a2 ), .dinb(a1 ), .dout(n268));
  jor  g00013(.dina(n268), .dinb(n256), .dout(n269));
  jor  g00014(.dina(n269), .dinb(n267), .dout(n270));
  jor  g00015(.dina(n262), .dinb(a0 ), .dout(n271));
  jor  g00016(.dina(n271), .dinb(n257), .dout(n272));
  jand g00017(.dina(n272), .dinb(n270), .dout(n273));
  jand g00018(.dina(n273), .dinb(n266), .dout(n274));
  jxor g00019(.dina(n274), .dinb(n261), .dout(f1 ));
  jand g00020(.dina(n258), .dinb(a2 ), .dout(n276));
  jand g00021(.dina(n276), .dinb(n274), .dout(n277));
  jor  g00022(.dina(n277), .dinb(n260), .dout(n278));
  jnot g00023(.din(b2 ), .dout(n279));
  jor  g00024(.dina(n269), .dinb(n279), .dout(n280));
  jor  g00025(.dina(n271), .dinb(n267), .dout(n281));
  jand g00026(.dina(n281), .dinb(n280), .dout(n282));
  jor  g00027(.dina(a1 ), .dinb(a0 ), .dout(n283));
  jor  g00028(.dina(n283), .dinb(n263), .dout(n284));
  jor  g00029(.dina(n284), .dinb(n257), .dout(n285));
  jand g00030(.dina(b1 ), .dinb(n257), .dout(n286));
  jxor g00031(.dina(n286), .dinb(n279), .dout(n287));
  jor  g00032(.dina(n287), .dinb(n264), .dout(n288));
  jand g00033(.dina(n288), .dinb(n285), .dout(n289));
  jand g00034(.dina(n289), .dinb(n282), .dout(n290));
  jxor g00035(.dina(n290), .dinb(n278), .dout(f2 ));
  jxor g00036(.dina(b3 ), .dinb(b2 ), .dout(n292));
  jnot g00037(.din(n292), .dout(n293));
  jor  g00038(.dina(b2 ), .dinb(b0 ), .dout(n294));
  jand g00039(.dina(n294), .dinb(b1 ), .dout(n295));
  jxor g00040(.dina(n295), .dinb(n293), .dout(n296));
  jor  g00041(.dina(n296), .dinb(n264), .dout(n297));
  jor  g00042(.dina(n284), .dinb(n267), .dout(n298));
  jnot g00043(.din(b3 ), .dout(n299));
  jor  g00044(.dina(n269), .dinb(n299), .dout(n300));
  jor  g00045(.dina(n271), .dinb(n279), .dout(n301));
  jand g00046(.dina(n301), .dinb(n300), .dout(n302));
  jand g00047(.dina(n302), .dinb(n298), .dout(n303));
  jand g00048(.dina(n303), .dinb(n297), .dout(n304));
  jxor g00049(.dina(n304), .dinb(n260), .dout(n305));
  jxor g00050(.dina(a3 ), .dinb(a2 ), .dout(n306));
  jand g00051(.dina(n306), .dinb(b0 ), .dout(n307));
  jxor g00052(.dina(n307), .dinb(n305), .dout(n308));
  jand g00053(.dina(n290), .dinb(n277), .dout(n309));
  jxor g00054(.dina(n309), .dinb(n308), .dout(f3 ));
  jand g00055(.dina(n307), .dinb(n305), .dout(n311));
  jand g00056(.dina(n309), .dinb(n308), .dout(n312));
  jor  g00057(.dina(n312), .dinb(n311), .dout(n313));
  jand g00058(.dina(b3 ), .dinb(b2 ), .dout(n314));
  jand g00059(.dina(n295), .dinb(n292), .dout(n315));
  jor  g00060(.dina(n315), .dinb(n314), .dout(n316));
  jxor g00061(.dina(b4 ), .dinb(b3 ), .dout(n317));
  jnot g00062(.din(n317), .dout(n318));
  jxor g00063(.dina(n318), .dinb(n316), .dout(n319));
  jor  g00064(.dina(n319), .dinb(n264), .dout(n320));
  jor  g00065(.dina(n284), .dinb(n279), .dout(n321));
  jnot g00066(.din(b4 ), .dout(n322));
  jor  g00067(.dina(n269), .dinb(n322), .dout(n323));
  jor  g00068(.dina(n271), .dinb(n299), .dout(n324));
  jand g00069(.dina(n324), .dinb(n323), .dout(n325));
  jand g00070(.dina(n325), .dinb(n321), .dout(n326));
  jand g00071(.dina(n326), .dinb(n320), .dout(n327));
  jxor g00072(.dina(n327), .dinb(n260), .dout(n328));
  jand g00073(.dina(n307), .dinb(a5 ), .dout(n329));
  jnot g00074(.din(n306), .dout(n330));
  jxor g00075(.dina(a5 ), .dinb(a4 ), .dout(n331));
  jor  g00076(.dina(n331), .dinb(n330), .dout(n332));
  jor  g00077(.dina(n332), .dinb(n267), .dout(n333));
  jnot g00078(.din(n333), .dout(n334));
  jxor g00079(.dina(a4 ), .dinb(a3 ), .dout(n335));
  jand g00080(.dina(n335), .dinb(n330), .dout(n336));
  jand g00081(.dina(n336), .dinb(b0 ), .dout(n337));
  jnot g00082(.din(n265), .dout(n338));
  jand g00083(.dina(n331), .dinb(n306), .dout(n339));
  jand g00084(.dina(n339), .dinb(n338), .dout(n340));
  jor  g00085(.dina(n340), .dinb(n337), .dout(n341));
  jor  g00086(.dina(n341), .dinb(n334), .dout(n342));
  jxor g00087(.dina(n342), .dinb(n329), .dout(n343));
  jxor g00088(.dina(n343), .dinb(n328), .dout(n344));
  jxor g00089(.dina(n344), .dinb(n313), .dout(f4 ));
  jand g00090(.dina(n343), .dinb(n328), .dout(n346));
  jand g00091(.dina(n344), .dinb(n313), .dout(n347));
  jor  g00092(.dina(n347), .dinb(n346), .dout(n348));
  jand g00093(.dina(b4 ), .dinb(b3 ), .dout(n349));
  jand g00094(.dina(n317), .dinb(n316), .dout(n350));
  jor  g00095(.dina(n350), .dinb(n349), .dout(n351));
  jxor g00096(.dina(b5 ), .dinb(b4 ), .dout(n352));
  jnot g00097(.din(n352), .dout(n353));
  jxor g00098(.dina(n353), .dinb(n351), .dout(n354));
  jor  g00099(.dina(n354), .dinb(n264), .dout(n355));
  jor  g00100(.dina(n284), .dinb(n299), .dout(n356));
  jnot g00101(.din(b5 ), .dout(n357));
  jor  g00102(.dina(n269), .dinb(n357), .dout(n358));
  jor  g00103(.dina(n271), .dinb(n322), .dout(n359));
  jand g00104(.dina(n359), .dinb(n358), .dout(n360));
  jand g00105(.dina(n360), .dinb(n356), .dout(n361));
  jand g00106(.dina(n361), .dinb(n355), .dout(n362));
  jxor g00107(.dina(n362), .dinb(n260), .dout(n363));
  jnot g00108(.din(a5 ), .dout(n364));
  jor  g00109(.dina(n307), .dinb(n364), .dout(n365));
  jor  g00110(.dina(n365), .dinb(n342), .dout(n366));
  jnot g00111(.din(n366), .dout(n367));
  jor  g00112(.dina(n367), .dinb(n364), .dout(n368));
  jnot g00113(.din(n331), .dout(n369));
  jor  g00114(.dina(n335), .dinb(n369), .dout(n370));
  jor  g00115(.dina(n370), .dinb(n306), .dout(n371));
  jor  g00116(.dina(n371), .dinb(n257), .dout(n372));
  jor  g00117(.dina(n332), .dinb(n279), .dout(n373));
  jand g00118(.dina(n336), .dinb(b1 ), .dout(n374));
  jnot g00119(.din(n287), .dout(n375));
  jand g00120(.dina(n339), .dinb(n375), .dout(n376));
  jor  g00121(.dina(n376), .dinb(n374), .dout(n377));
  jnot g00122(.din(n377), .dout(n378));
  jand g00123(.dina(n378), .dinb(n373), .dout(n379));
  jand g00124(.dina(n379), .dinb(n372), .dout(n380));
  jxor g00125(.dina(n380), .dinb(n368), .dout(n381));
  jxor g00126(.dina(n381), .dinb(n363), .dout(n382));
  jxor g00127(.dina(n382), .dinb(n348), .dout(f5 ));
  jand g00128(.dina(n381), .dinb(n363), .dout(n384));
  jand g00129(.dina(n382), .dinb(n348), .dout(n385));
  jor  g00130(.dina(n385), .dinb(n384), .dout(n386));
  jand g00131(.dina(b5 ), .dinb(b4 ), .dout(n387));
  jand g00132(.dina(n352), .dinb(n351), .dout(n388));
  jor  g00133(.dina(n388), .dinb(n387), .dout(n389));
  jxor g00134(.dina(b6 ), .dinb(b5 ), .dout(n390));
  jnot g00135(.din(n390), .dout(n391));
  jxor g00136(.dina(n391), .dinb(n389), .dout(n392));
  jor  g00137(.dina(n392), .dinb(n264), .dout(n393));
  jor  g00138(.dina(n284), .dinb(n322), .dout(n394));
  jnot g00139(.din(b6 ), .dout(n395));
  jor  g00140(.dina(n269), .dinb(n395), .dout(n396));
  jor  g00141(.dina(n271), .dinb(n357), .dout(n397));
  jand g00142(.dina(n397), .dinb(n396), .dout(n398));
  jand g00143(.dina(n398), .dinb(n394), .dout(n399));
  jand g00144(.dina(n399), .dinb(n393), .dout(n400));
  jxor g00145(.dina(n400), .dinb(n260), .dout(n401));
  jnot g00146(.din(n339), .dout(n402));
  jor  g00147(.dina(n402), .dinb(n296), .dout(n403));
  jor  g00148(.dina(n371), .dinb(n267), .dout(n404));
  jnot g00149(.din(n336), .dout(n405));
  jor  g00150(.dina(n405), .dinb(n279), .dout(n406));
  jor  g00151(.dina(n332), .dinb(n299), .dout(n407));
  jand g00152(.dina(n407), .dinb(n406), .dout(n408));
  jand g00153(.dina(n408), .dinb(n404), .dout(n409));
  jand g00154(.dina(n409), .dinb(n403), .dout(n410));
  jxor g00155(.dina(n410), .dinb(a5 ), .dout(n411));
  jnot g00156(.din(n411), .dout(n412));
  jxor g00157(.dina(a6 ), .dinb(a5 ), .dout(n413));
  jand g00158(.dina(n413), .dinb(b0 ), .dout(n414));
  jand g00159(.dina(n380), .dinb(n367), .dout(n415));
  jxor g00160(.dina(n415), .dinb(n414), .dout(n416));
  jxor g00161(.dina(n416), .dinb(n412), .dout(n417));
  jxor g00162(.dina(n417), .dinb(n401), .dout(n418));
  jxor g00163(.dina(n418), .dinb(n386), .dout(f6 ));
  jand g00164(.dina(n417), .dinb(n401), .dout(n420));
  jand g00165(.dina(n418), .dinb(n386), .dout(n421));
  jor  g00166(.dina(n421), .dinb(n420), .dout(n422));
  jand g00167(.dina(b6 ), .dinb(b5 ), .dout(n423));
  jand g00168(.dina(n390), .dinb(n389), .dout(n424));
  jor  g00169(.dina(n424), .dinb(n423), .dout(n425));
  jxor g00170(.dina(b7 ), .dinb(b6 ), .dout(n426));
  jnot g00171(.din(n426), .dout(n427));
  jxor g00172(.dina(n427), .dinb(n425), .dout(n428));
  jor  g00173(.dina(n428), .dinb(n264), .dout(n429));
  jor  g00174(.dina(n284), .dinb(n357), .dout(n430));
  jnot g00175(.din(b7 ), .dout(n431));
  jor  g00176(.dina(n269), .dinb(n431), .dout(n432));
  jor  g00177(.dina(n271), .dinb(n395), .dout(n433));
  jand g00178(.dina(n433), .dinb(n432), .dout(n434));
  jand g00179(.dina(n434), .dinb(n430), .dout(n435));
  jand g00180(.dina(n435), .dinb(n429), .dout(n436));
  jxor g00181(.dina(n436), .dinb(n260), .dout(n437));
  jand g00182(.dina(n415), .dinb(n414), .dout(n438));
  jand g00183(.dina(n416), .dinb(n412), .dout(n439));
  jor  g00184(.dina(n439), .dinb(n438), .dout(n440));
  jor  g00185(.dina(n402), .dinb(n319), .dout(n441));
  jor  g00186(.dina(n371), .dinb(n279), .dout(n442));
  jor  g00187(.dina(n405), .dinb(n299), .dout(n443));
  jor  g00188(.dina(n332), .dinb(n322), .dout(n444));
  jand g00189(.dina(n444), .dinb(n443), .dout(n445));
  jand g00190(.dina(n445), .dinb(n442), .dout(n446));
  jand g00191(.dina(n446), .dinb(n441), .dout(n447));
  jxor g00192(.dina(n447), .dinb(a5 ), .dout(n448));
  jand g00193(.dina(n414), .dinb(a8 ), .dout(n449));
  jxor g00194(.dina(a8 ), .dinb(a7 ), .dout(n450));
  jnot g00195(.din(n450), .dout(n451));
  jand g00196(.dina(n451), .dinb(n413), .dout(n452));
  jand g00197(.dina(n452), .dinb(b1 ), .dout(n453));
  jnot g00198(.din(n413), .dout(n454));
  jxor g00199(.dina(a7 ), .dinb(a6 ), .dout(n455));
  jand g00200(.dina(n455), .dinb(n454), .dout(n456));
  jand g00201(.dina(n456), .dinb(b0 ), .dout(n457));
  jand g00202(.dina(n450), .dinb(n413), .dout(n458));
  jand g00203(.dina(n458), .dinb(n338), .dout(n459));
  jor  g00204(.dina(n459), .dinb(n457), .dout(n460));
  jor  g00205(.dina(n460), .dinb(n453), .dout(n461));
  jxor g00206(.dina(n461), .dinb(n449), .dout(n462));
  jxor g00207(.dina(n462), .dinb(n448), .dout(n463));
  jnot g00208(.din(n463), .dout(n464));
  jxor g00209(.dina(n464), .dinb(n440), .dout(n465));
  jxor g00210(.dina(n465), .dinb(n437), .dout(n466));
  jxor g00211(.dina(n466), .dinb(n422), .dout(f7 ));
  jand g00212(.dina(n465), .dinb(n437), .dout(n468));
  jand g00213(.dina(n466), .dinb(n422), .dout(n469));
  jor  g00214(.dina(n469), .dinb(n468), .dout(n470));
  jnot g00215(.din(n448), .dout(n471));
  jand g00216(.dina(n462), .dinb(n471), .dout(n472));
  jand g00217(.dina(n464), .dinb(n440), .dout(n473));
  jor  g00218(.dina(n473), .dinb(n472), .dout(n474));
  jor  g00219(.dina(n354), .dinb(n402), .dout(n475));
  jor  g00220(.dina(n371), .dinb(n299), .dout(n476));
  jor  g00221(.dina(n405), .dinb(n322), .dout(n477));
  jor  g00222(.dina(n332), .dinb(n357), .dout(n478));
  jand g00223(.dina(n478), .dinb(n477), .dout(n479));
  jand g00224(.dina(n479), .dinb(n476), .dout(n480));
  jand g00225(.dina(n480), .dinb(n475), .dout(n481));
  jxor g00226(.dina(n481), .dinb(a5 ), .dout(n482));
  jnot g00227(.din(a8 ), .dout(n483));
  jnot g00228(.din(n461), .dout(n484));
  jnot g00229(.din(n414), .dout(n485));
  jand g00230(.dina(n485), .dinb(a8 ), .dout(n486));
  jand g00231(.dina(n486), .dinb(n484), .dout(n487));
  jor  g00232(.dina(n487), .dinb(n483), .dout(n488));
  jor  g00233(.dina(n455), .dinb(n451), .dout(n489));
  jor  g00234(.dina(n489), .dinb(n413), .dout(n490));
  jnot g00235(.din(n490), .dout(n491));
  jand g00236(.dina(n491), .dinb(b0 ), .dout(n492));
  jand g00237(.dina(n452), .dinb(b2 ), .dout(n493));
  jand g00238(.dina(n456), .dinb(b1 ), .dout(n494));
  jand g00239(.dina(n458), .dinb(n375), .dout(n495));
  jor  g00240(.dina(n495), .dinb(n494), .dout(n496));
  jor  g00241(.dina(n496), .dinb(n493), .dout(n497));
  jor  g00242(.dina(n497), .dinb(n492), .dout(n498));
  jnot g00243(.din(n498), .dout(n499));
  jxor g00244(.dina(n499), .dinb(n488), .dout(n500));
  jxor g00245(.dina(n500), .dinb(n482), .dout(n501));
  jnot g00246(.din(n501), .dout(n502));
  jxor g00247(.dina(n502), .dinb(n474), .dout(n503));
  jand g00248(.dina(b7 ), .dinb(b6 ), .dout(n504));
  jand g00249(.dina(n426), .dinb(n425), .dout(n505));
  jor  g00250(.dina(n505), .dinb(n504), .dout(n506));
  jxor g00251(.dina(b8 ), .dinb(b7 ), .dout(n507));
  jnot g00252(.din(n507), .dout(n508));
  jxor g00253(.dina(n508), .dinb(n506), .dout(n509));
  jor  g00254(.dina(n509), .dinb(n264), .dout(n510));
  jor  g00255(.dina(n284), .dinb(n395), .dout(n511));
  jnot g00256(.din(b8 ), .dout(n512));
  jor  g00257(.dina(n269), .dinb(n512), .dout(n513));
  jor  g00258(.dina(n271), .dinb(n431), .dout(n514));
  jand g00259(.dina(n514), .dinb(n513), .dout(n515));
  jand g00260(.dina(n515), .dinb(n511), .dout(n516));
  jand g00261(.dina(n516), .dinb(n510), .dout(n517));
  jxor g00262(.dina(n517), .dinb(n260), .dout(n518));
  jxor g00263(.dina(n518), .dinb(n503), .dout(n519));
  jxor g00264(.dina(n519), .dinb(n470), .dout(f8 ));
  jand g00265(.dina(n518), .dinb(n503), .dout(n521));
  jand g00266(.dina(n519), .dinb(n470), .dout(n522));
  jor  g00267(.dina(n522), .dinb(n521), .dout(n523));
  jnot g00268(.din(n482), .dout(n524));
  jand g00269(.dina(n500), .dinb(n524), .dout(n525));
  jand g00270(.dina(n502), .dinb(n474), .dout(n526));
  jor  g00271(.dina(n526), .dinb(n525), .dout(n527));
  jnot g00272(.din(n458), .dout(n528));
  jor  g00273(.dina(n528), .dinb(n296), .dout(n529));
  jor  g00274(.dina(n490), .dinb(n267), .dout(n530));
  jnot g00275(.din(n456), .dout(n531));
  jor  g00276(.dina(n531), .dinb(n279), .dout(n532));
  jnot g00277(.din(n452), .dout(n533));
  jor  g00278(.dina(n533), .dinb(n299), .dout(n534));
  jand g00279(.dina(n534), .dinb(n532), .dout(n535));
  jand g00280(.dina(n535), .dinb(n530), .dout(n536));
  jand g00281(.dina(n536), .dinb(n529), .dout(n537));
  jxor g00282(.dina(n537), .dinb(a8 ), .dout(n538));
  jnot g00283(.din(n538), .dout(n539));
  jxor g00284(.dina(a9 ), .dinb(a8 ), .dout(n540));
  jand g00285(.dina(n540), .dinb(b0 ), .dout(n541));
  jand g00286(.dina(n499), .dinb(n487), .dout(n542));
  jxor g00287(.dina(n542), .dinb(n541), .dout(n543));
  jxor g00288(.dina(n543), .dinb(n539), .dout(n544));
  jnot g00289(.din(n544), .dout(n545));
  jor  g00290(.dina(n392), .dinb(n402), .dout(n546));
  jor  g00291(.dina(n371), .dinb(n322), .dout(n547));
  jor  g00292(.dina(n405), .dinb(n357), .dout(n548));
  jor  g00293(.dina(n332), .dinb(n395), .dout(n549));
  jand g00294(.dina(n549), .dinb(n548), .dout(n550));
  jand g00295(.dina(n550), .dinb(n547), .dout(n551));
  jand g00296(.dina(n551), .dinb(n546), .dout(n552));
  jxor g00297(.dina(n552), .dinb(a5 ), .dout(n553));
  jxor g00298(.dina(n553), .dinb(n545), .dout(n554));
  jxor g00299(.dina(n554), .dinb(n527), .dout(n555));
  jand g00300(.dina(b8 ), .dinb(b7 ), .dout(n556));
  jand g00301(.dina(n507), .dinb(n506), .dout(n557));
  jor  g00302(.dina(n557), .dinb(n556), .dout(n558));
  jxor g00303(.dina(b9 ), .dinb(b8 ), .dout(n559));
  jnot g00304(.din(n559), .dout(n560));
  jxor g00305(.dina(n560), .dinb(n558), .dout(n561));
  jor  g00306(.dina(n561), .dinb(n264), .dout(n562));
  jor  g00307(.dina(n284), .dinb(n431), .dout(n563));
  jnot g00308(.din(b9 ), .dout(n564));
  jor  g00309(.dina(n269), .dinb(n564), .dout(n565));
  jor  g00310(.dina(n271), .dinb(n512), .dout(n566));
  jand g00311(.dina(n566), .dinb(n565), .dout(n567));
  jand g00312(.dina(n567), .dinb(n563), .dout(n568));
  jand g00313(.dina(n568), .dinb(n562), .dout(n569));
  jxor g00314(.dina(n569), .dinb(n260), .dout(n570));
  jxor g00315(.dina(n570), .dinb(n555), .dout(n571));
  jxor g00316(.dina(n571), .dinb(n523), .dout(f9 ));
  jand g00317(.dina(n570), .dinb(n555), .dout(n573));
  jand g00318(.dina(n571), .dinb(n523), .dout(n574));
  jor  g00319(.dina(n574), .dinb(n573), .dout(n575));
  jor  g00320(.dina(n553), .dinb(n545), .dout(n576));
  jnot g00321(.din(n576), .dout(n577));
  jand g00322(.dina(n554), .dinb(n527), .dout(n578));
  jor  g00323(.dina(n578), .dinb(n577), .dout(n579));
  jand g00324(.dina(n542), .dinb(n541), .dout(n580));
  jand g00325(.dina(n543), .dinb(n539), .dout(n581));
  jor  g00326(.dina(n581), .dinb(n580), .dout(n582));
  jor  g00327(.dina(n528), .dinb(n319), .dout(n583));
  jor  g00328(.dina(n490), .dinb(n279), .dout(n584));
  jor  g00329(.dina(n531), .dinb(n299), .dout(n585));
  jor  g00330(.dina(n533), .dinb(n322), .dout(n586));
  jand g00331(.dina(n586), .dinb(n585), .dout(n587));
  jand g00332(.dina(n587), .dinb(n584), .dout(n588));
  jand g00333(.dina(n588), .dinb(n583), .dout(n589));
  jxor g00334(.dina(n589), .dinb(a8 ), .dout(n590));
  jnot g00335(.din(n590), .dout(n591));
  jand g00336(.dina(n541), .dinb(a11 ), .dout(n592));
  jxor g00337(.dina(a11 ), .dinb(a10 ), .dout(n593));
  jnot g00338(.din(n593), .dout(n594));
  jand g00339(.dina(n594), .dinb(n540), .dout(n595));
  jand g00340(.dina(n595), .dinb(b1 ), .dout(n596));
  jnot g00341(.din(n540), .dout(n597));
  jxor g00342(.dina(a10 ), .dinb(a9 ), .dout(n598));
  jand g00343(.dina(n598), .dinb(n597), .dout(n599));
  jand g00344(.dina(n599), .dinb(b0 ), .dout(n600));
  jand g00345(.dina(n593), .dinb(n540), .dout(n601));
  jand g00346(.dina(n601), .dinb(n338), .dout(n602));
  jor  g00347(.dina(n602), .dinb(n600), .dout(n603));
  jor  g00348(.dina(n603), .dinb(n596), .dout(n604));
  jxor g00349(.dina(n604), .dinb(n592), .dout(n605));
  jxor g00350(.dina(n605), .dinb(n591), .dout(n606));
  jxor g00351(.dina(n606), .dinb(n582), .dout(n607));
  jnot g00352(.din(n607), .dout(n608));
  jor  g00353(.dina(n428), .dinb(n402), .dout(n609));
  jor  g00354(.dina(n371), .dinb(n357), .dout(n610));
  jor  g00355(.dina(n405), .dinb(n395), .dout(n611));
  jor  g00356(.dina(n332), .dinb(n431), .dout(n612));
  jand g00357(.dina(n612), .dinb(n611), .dout(n613));
  jand g00358(.dina(n613), .dinb(n610), .dout(n614));
  jand g00359(.dina(n614), .dinb(n609), .dout(n615));
  jxor g00360(.dina(n615), .dinb(a5 ), .dout(n616));
  jxor g00361(.dina(n616), .dinb(n608), .dout(n617));
  jxor g00362(.dina(n617), .dinb(n579), .dout(n618));
  jand g00363(.dina(b9 ), .dinb(b8 ), .dout(n619));
  jand g00364(.dina(n559), .dinb(n558), .dout(n620));
  jor  g00365(.dina(n620), .dinb(n619), .dout(n621));
  jxor g00366(.dina(b10 ), .dinb(b9 ), .dout(n622));
  jnot g00367(.din(n622), .dout(n623));
  jxor g00368(.dina(n623), .dinb(n621), .dout(n624));
  jor  g00369(.dina(n624), .dinb(n264), .dout(n625));
  jor  g00370(.dina(n284), .dinb(n512), .dout(n626));
  jnot g00371(.din(b10 ), .dout(n627));
  jor  g00372(.dina(n269), .dinb(n627), .dout(n628));
  jor  g00373(.dina(n271), .dinb(n564), .dout(n629));
  jand g00374(.dina(n629), .dinb(n628), .dout(n630));
  jand g00375(.dina(n630), .dinb(n626), .dout(n631));
  jand g00376(.dina(n631), .dinb(n625), .dout(n632));
  jxor g00377(.dina(n632), .dinb(n260), .dout(n633));
  jxor g00378(.dina(n633), .dinb(n618), .dout(n634));
  jxor g00379(.dina(n634), .dinb(n575), .dout(f10 ));
  jand g00380(.dina(n633), .dinb(n618), .dout(n636));
  jand g00381(.dina(n634), .dinb(n575), .dout(n637));
  jor  g00382(.dina(n637), .dinb(n636), .dout(n638));
  jand g00383(.dina(b10 ), .dinb(b9 ), .dout(n639));
  jand g00384(.dina(n622), .dinb(n621), .dout(n640));
  jor  g00385(.dina(n640), .dinb(n639), .dout(n641));
  jxor g00386(.dina(b11 ), .dinb(b10 ), .dout(n642));
  jnot g00387(.din(n642), .dout(n643));
  jxor g00388(.dina(n643), .dinb(n641), .dout(n644));
  jor  g00389(.dina(n644), .dinb(n264), .dout(n645));
  jor  g00390(.dina(n284), .dinb(n564), .dout(n646));
  jnot g00391(.din(b11 ), .dout(n647));
  jor  g00392(.dina(n269), .dinb(n647), .dout(n648));
  jor  g00393(.dina(n271), .dinb(n627), .dout(n649));
  jand g00394(.dina(n649), .dinb(n648), .dout(n650));
  jand g00395(.dina(n650), .dinb(n646), .dout(n651));
  jand g00396(.dina(n651), .dinb(n645), .dout(n652));
  jxor g00397(.dina(n652), .dinb(n260), .dout(n653));
  jor  g00398(.dina(n616), .dinb(n608), .dout(n654));
  jnot g00399(.din(n654), .dout(n655));
  jand g00400(.dina(n617), .dinb(n579), .dout(n656));
  jor  g00401(.dina(n656), .dinb(n655), .dout(n657));
  jor  g00402(.dina(n509), .dinb(n402), .dout(n658));
  jor  g00403(.dina(n371), .dinb(n395), .dout(n659));
  jor  g00404(.dina(n405), .dinb(n431), .dout(n660));
  jor  g00405(.dina(n332), .dinb(n512), .dout(n661));
  jand g00406(.dina(n661), .dinb(n660), .dout(n662));
  jand g00407(.dina(n662), .dinb(n659), .dout(n663));
  jand g00408(.dina(n663), .dinb(n658), .dout(n664));
  jxor g00409(.dina(n664), .dinb(a5 ), .dout(n665));
  jand g00410(.dina(n605), .dinb(n591), .dout(n666));
  jand g00411(.dina(n606), .dinb(n582), .dout(n667));
  jor  g00412(.dina(n667), .dinb(n666), .dout(n668));
  jor  g00413(.dina(n528), .dinb(n354), .dout(n669));
  jor  g00414(.dina(n490), .dinb(n299), .dout(n670));
  jor  g00415(.dina(n531), .dinb(n322), .dout(n671));
  jor  g00416(.dina(n533), .dinb(n357), .dout(n672));
  jand g00417(.dina(n672), .dinb(n671), .dout(n673));
  jand g00418(.dina(n673), .dinb(n670), .dout(n674));
  jand g00419(.dina(n674), .dinb(n669), .dout(n675));
  jxor g00420(.dina(n675), .dinb(a8 ), .dout(n676));
  jnot g00421(.din(n676), .dout(n677));
  jnot g00422(.din(a11 ), .dout(n678));
  jor  g00423(.dina(n541), .dinb(n678), .dout(n679));
  jor  g00424(.dina(n679), .dinb(n604), .dout(n680));
  jand g00425(.dina(n680), .dinb(a11 ), .dout(n681));
  jor  g00426(.dina(n598), .dinb(n594), .dout(n682));
  jor  g00427(.dina(n682), .dinb(n540), .dout(n683));
  jnot g00428(.din(n683), .dout(n684));
  jand g00429(.dina(n684), .dinb(b0 ), .dout(n685));
  jand g00430(.dina(n595), .dinb(b2 ), .dout(n686));
  jand g00431(.dina(n599), .dinb(b1 ), .dout(n687));
  jand g00432(.dina(n601), .dinb(n375), .dout(n688));
  jor  g00433(.dina(n688), .dinb(n687), .dout(n689));
  jor  g00434(.dina(n689), .dinb(n686), .dout(n690));
  jor  g00435(.dina(n690), .dinb(n685), .dout(n691));
  jxor g00436(.dina(n691), .dinb(n681), .dout(n692));
  jxor g00437(.dina(n692), .dinb(n677), .dout(n693));
  jxor g00438(.dina(n693), .dinb(n668), .dout(n694));
  jxor g00439(.dina(n694), .dinb(n665), .dout(n695));
  jnot g00440(.din(n695), .dout(n696));
  jxor g00441(.dina(n696), .dinb(n657), .dout(n697));
  jxor g00442(.dina(n697), .dinb(n653), .dout(n698));
  jxor g00443(.dina(n698), .dinb(n638), .dout(f11 ));
  jand g00444(.dina(n697), .dinb(n653), .dout(n700));
  jand g00445(.dina(n698), .dinb(n638), .dout(n701));
  jor  g00446(.dina(n701), .dinb(n700), .dout(n702));
  jand g00447(.dina(n692), .dinb(n677), .dout(n703));
  jand g00448(.dina(n693), .dinb(n668), .dout(n704));
  jor  g00449(.dina(n704), .dinb(n703), .dout(n705));
  jnot g00450(.din(n601), .dout(n706));
  jor  g00451(.dina(n706), .dinb(n296), .dout(n707));
  jor  g00452(.dina(n683), .dinb(n267), .dout(n708));
  jnot g00453(.din(n599), .dout(n709));
  jor  g00454(.dina(n709), .dinb(n279), .dout(n710));
  jnot g00455(.din(n595), .dout(n711));
  jor  g00456(.dina(n711), .dinb(n299), .dout(n712));
  jand g00457(.dina(n712), .dinb(n710), .dout(n713));
  jand g00458(.dina(n713), .dinb(n708), .dout(n714));
  jand g00459(.dina(n714), .dinb(n707), .dout(n715));
  jxor g00460(.dina(n715), .dinb(a11 ), .dout(n716));
  jnot g00461(.din(n716), .dout(n717));
  jxor g00462(.dina(a12 ), .dinb(a11 ), .dout(n718));
  jand g00463(.dina(n718), .dinb(b0 ), .dout(n719));
  jnot g00464(.din(n719), .dout(n720));
  jor  g00465(.dina(n691), .dinb(n680), .dout(n721));
  jxor g00466(.dina(n721), .dinb(n720), .dout(n722));
  jxor g00467(.dina(n722), .dinb(n717), .dout(n723));
  jnot g00468(.din(n723), .dout(n724));
  jor  g00469(.dina(n528), .dinb(n392), .dout(n725));
  jor  g00470(.dina(n490), .dinb(n322), .dout(n726));
  jor  g00471(.dina(n531), .dinb(n357), .dout(n727));
  jor  g00472(.dina(n533), .dinb(n395), .dout(n728));
  jand g00473(.dina(n728), .dinb(n727), .dout(n729));
  jand g00474(.dina(n729), .dinb(n726), .dout(n730));
  jand g00475(.dina(n730), .dinb(n725), .dout(n731));
  jxor g00476(.dina(n731), .dinb(a8 ), .dout(n732));
  jxor g00477(.dina(n732), .dinb(n724), .dout(n733));
  jxor g00478(.dina(n733), .dinb(n705), .dout(n734));
  jnot g00479(.din(n734), .dout(n735));
  jor  g00480(.dina(n561), .dinb(n402), .dout(n736));
  jor  g00481(.dina(n371), .dinb(n431), .dout(n737));
  jor  g00482(.dina(n405), .dinb(n512), .dout(n738));
  jor  g00483(.dina(n332), .dinb(n564), .dout(n739));
  jand g00484(.dina(n739), .dinb(n738), .dout(n740));
  jand g00485(.dina(n740), .dinb(n737), .dout(n741));
  jand g00486(.dina(n741), .dinb(n736), .dout(n742));
  jxor g00487(.dina(n742), .dinb(a5 ), .dout(n743));
  jxor g00488(.dina(n743), .dinb(n735), .dout(n744));
  jnot g00489(.din(n665), .dout(n745));
  jand g00490(.dina(n694), .dinb(n745), .dout(n746));
  jand g00491(.dina(n696), .dinb(n657), .dout(n747));
  jor  g00492(.dina(n747), .dinb(n746), .dout(n748));
  jxor g00493(.dina(n748), .dinb(n744), .dout(n749));
  jand g00494(.dina(b11 ), .dinb(b10 ), .dout(n750));
  jand g00495(.dina(n642), .dinb(n641), .dout(n751));
  jor  g00496(.dina(n751), .dinb(n750), .dout(n752));
  jxor g00497(.dina(b12 ), .dinb(b11 ), .dout(n753));
  jnot g00498(.din(n753), .dout(n754));
  jxor g00499(.dina(n754), .dinb(n752), .dout(n755));
  jor  g00500(.dina(n755), .dinb(n264), .dout(n756));
  jor  g00501(.dina(n284), .dinb(n627), .dout(n757));
  jnot g00502(.din(b12 ), .dout(n758));
  jor  g00503(.dina(n269), .dinb(n758), .dout(n759));
  jor  g00504(.dina(n271), .dinb(n647), .dout(n760));
  jand g00505(.dina(n760), .dinb(n759), .dout(n761));
  jand g00506(.dina(n761), .dinb(n757), .dout(n762));
  jand g00507(.dina(n762), .dinb(n756), .dout(n763));
  jxor g00508(.dina(n763), .dinb(n260), .dout(n764));
  jxor g00509(.dina(n764), .dinb(n749), .dout(n765));
  jxor g00510(.dina(n765), .dinb(n702), .dout(f12 ));
  jand g00511(.dina(n764), .dinb(n749), .dout(n767));
  jand g00512(.dina(n765), .dinb(n702), .dout(n768));
  jor  g00513(.dina(n768), .dinb(n767), .dout(n769));
  jand g00514(.dina(b12 ), .dinb(b11 ), .dout(n770));
  jand g00515(.dina(n753), .dinb(n752), .dout(n771));
  jor  g00516(.dina(n771), .dinb(n770), .dout(n772));
  jxor g00517(.dina(b13 ), .dinb(b12 ), .dout(n773));
  jnot g00518(.din(n773), .dout(n774));
  jxor g00519(.dina(n774), .dinb(n772), .dout(n775));
  jor  g00520(.dina(n775), .dinb(n264), .dout(n776));
  jor  g00521(.dina(n284), .dinb(n647), .dout(n777));
  jnot g00522(.din(b13 ), .dout(n778));
  jor  g00523(.dina(n269), .dinb(n778), .dout(n779));
  jor  g00524(.dina(n271), .dinb(n758), .dout(n780));
  jand g00525(.dina(n780), .dinb(n779), .dout(n781));
  jand g00526(.dina(n781), .dinb(n777), .dout(n782));
  jand g00527(.dina(n782), .dinb(n776), .dout(n783));
  jxor g00528(.dina(n783), .dinb(n260), .dout(n784));
  jor  g00529(.dina(n743), .dinb(n735), .dout(n785));
  jnot g00530(.din(n785), .dout(n786));
  jand g00531(.dina(n748), .dinb(n744), .dout(n787));
  jor  g00532(.dina(n787), .dinb(n786), .dout(n788));
  jor  g00533(.dina(n732), .dinb(n724), .dout(n789));
  jand g00534(.dina(n733), .dinb(n705), .dout(n790));
  jnot g00535(.din(n790), .dout(n791));
  jand g00536(.dina(n791), .dinb(n789), .dout(n792));
  jnot g00537(.din(n721), .dout(n793));
  jand g00538(.dina(n793), .dinb(n719), .dout(n794));
  jand g00539(.dina(n722), .dinb(n717), .dout(n795));
  jor  g00540(.dina(n795), .dinb(n794), .dout(n796));
  jor  g00541(.dina(n706), .dinb(n319), .dout(n797));
  jor  g00542(.dina(n683), .dinb(n279), .dout(n798));
  jor  g00543(.dina(n709), .dinb(n299), .dout(n799));
  jor  g00544(.dina(n711), .dinb(n322), .dout(n800));
  jand g00545(.dina(n800), .dinb(n799), .dout(n801));
  jand g00546(.dina(n801), .dinb(n798), .dout(n802));
  jand g00547(.dina(n802), .dinb(n797), .dout(n803));
  jxor g00548(.dina(n803), .dinb(a11 ), .dout(n804));
  jnot g00549(.din(n804), .dout(n805));
  jand g00550(.dina(n719), .dinb(a14 ), .dout(n806));
  jxor g00551(.dina(a14 ), .dinb(a13 ), .dout(n807));
  jnot g00552(.din(n807), .dout(n808));
  jand g00553(.dina(n808), .dinb(n718), .dout(n809));
  jand g00554(.dina(n809), .dinb(b1 ), .dout(n810));
  jnot g00555(.din(n718), .dout(n811));
  jxor g00556(.dina(a13 ), .dinb(a12 ), .dout(n812));
  jand g00557(.dina(n812), .dinb(n811), .dout(n813));
  jand g00558(.dina(n813), .dinb(b0 ), .dout(n814));
  jand g00559(.dina(n807), .dinb(n718), .dout(n815));
  jand g00560(.dina(n815), .dinb(n338), .dout(n816));
  jor  g00561(.dina(n816), .dinb(n814), .dout(n817));
  jor  g00562(.dina(n817), .dinb(n810), .dout(n818));
  jxor g00563(.dina(n818), .dinb(n806), .dout(n819));
  jxor g00564(.dina(n819), .dinb(n805), .dout(n820));
  jxor g00565(.dina(n820), .dinb(n796), .dout(n821));
  jnot g00566(.din(n821), .dout(n822));
  jor  g00567(.dina(n528), .dinb(n428), .dout(n823));
  jor  g00568(.dina(n490), .dinb(n357), .dout(n824));
  jor  g00569(.dina(n531), .dinb(n395), .dout(n825));
  jor  g00570(.dina(n533), .dinb(n431), .dout(n826));
  jand g00571(.dina(n826), .dinb(n825), .dout(n827));
  jand g00572(.dina(n827), .dinb(n824), .dout(n828));
  jand g00573(.dina(n828), .dinb(n823), .dout(n829));
  jxor g00574(.dina(n829), .dinb(a8 ), .dout(n830));
  jxor g00575(.dina(n830), .dinb(n822), .dout(n831));
  jnot g00576(.din(n831), .dout(n832));
  jxor g00577(.dina(n832), .dinb(n792), .dout(n833));
  jor  g00578(.dina(n624), .dinb(n402), .dout(n834));
  jor  g00579(.dina(n371), .dinb(n512), .dout(n835));
  jor  g00580(.dina(n405), .dinb(n564), .dout(n836));
  jor  g00581(.dina(n332), .dinb(n627), .dout(n837));
  jand g00582(.dina(n837), .dinb(n836), .dout(n838));
  jand g00583(.dina(n838), .dinb(n835), .dout(n839));
  jand g00584(.dina(n839), .dinb(n834), .dout(n840));
  jxor g00585(.dina(n840), .dinb(a5 ), .dout(n841));
  jxor g00586(.dina(n841), .dinb(n833), .dout(n842));
  jnot g00587(.din(n842), .dout(n843));
  jxor g00588(.dina(n843), .dinb(n788), .dout(n844));
  jxor g00589(.dina(n844), .dinb(n784), .dout(n845));
  jxor g00590(.dina(n845), .dinb(n769), .dout(f13 ));
  jand g00591(.dina(n844), .dinb(n784), .dout(n847));
  jand g00592(.dina(n845), .dinb(n769), .dout(n848));
  jor  g00593(.dina(n848), .dinb(n847), .dout(n849));
  jand g00594(.dina(b13 ), .dinb(b12 ), .dout(n850));
  jand g00595(.dina(n773), .dinb(n772), .dout(n851));
  jor  g00596(.dina(n851), .dinb(n850), .dout(n852));
  jxor g00597(.dina(b14 ), .dinb(b13 ), .dout(n853));
  jnot g00598(.din(n853), .dout(n854));
  jxor g00599(.dina(n854), .dinb(n852), .dout(n855));
  jor  g00600(.dina(n855), .dinb(n264), .dout(n856));
  jor  g00601(.dina(n284), .dinb(n758), .dout(n857));
  jnot g00602(.din(b14 ), .dout(n858));
  jor  g00603(.dina(n269), .dinb(n858), .dout(n859));
  jor  g00604(.dina(n271), .dinb(n778), .dout(n860));
  jand g00605(.dina(n860), .dinb(n859), .dout(n861));
  jand g00606(.dina(n861), .dinb(n857), .dout(n862));
  jand g00607(.dina(n862), .dinb(n856), .dout(n863));
  jxor g00608(.dina(n863), .dinb(n260), .dout(n864));
  jnot g00609(.din(n833), .dout(n865));
  jor  g00610(.dina(n841), .dinb(n865), .dout(n866));
  jnot g00611(.din(n866), .dout(n867));
  jand g00612(.dina(n843), .dinb(n788), .dout(n868));
  jor  g00613(.dina(n868), .dinb(n867), .dout(n869));
  jor  g00614(.dina(n644), .dinb(n402), .dout(n870));
  jor  g00615(.dina(n371), .dinb(n564), .dout(n871));
  jor  g00616(.dina(n405), .dinb(n627), .dout(n872));
  jor  g00617(.dina(n332), .dinb(n647), .dout(n873));
  jand g00618(.dina(n873), .dinb(n872), .dout(n874));
  jand g00619(.dina(n874), .dinb(n871), .dout(n875));
  jand g00620(.dina(n875), .dinb(n870), .dout(n876));
  jxor g00621(.dina(n876), .dinb(a5 ), .dout(n877));
  jor  g00622(.dina(n830), .dinb(n822), .dout(n878));
  jor  g00623(.dina(n832), .dinb(n792), .dout(n879));
  jand g00624(.dina(n879), .dinb(n878), .dout(n880));
  jor  g00625(.dina(n509), .dinb(n528), .dout(n881));
  jor  g00626(.dina(n490), .dinb(n395), .dout(n882));
  jor  g00627(.dina(n531), .dinb(n431), .dout(n883));
  jor  g00628(.dina(n533), .dinb(n512), .dout(n884));
  jand g00629(.dina(n884), .dinb(n883), .dout(n885));
  jand g00630(.dina(n885), .dinb(n882), .dout(n886));
  jand g00631(.dina(n886), .dinb(n881), .dout(n887));
  jxor g00632(.dina(n887), .dinb(a8 ), .dout(n888));
  jnot g00633(.din(n888), .dout(n889));
  jand g00634(.dina(n819), .dinb(n805), .dout(n890));
  jand g00635(.dina(n820), .dinb(n796), .dout(n891));
  jor  g00636(.dina(n891), .dinb(n890), .dout(n892));
  jor  g00637(.dina(n706), .dinb(n354), .dout(n893));
  jor  g00638(.dina(n683), .dinb(n299), .dout(n894));
  jor  g00639(.dina(n709), .dinb(n322), .dout(n895));
  jor  g00640(.dina(n711), .dinb(n357), .dout(n896));
  jand g00641(.dina(n896), .dinb(n895), .dout(n897));
  jand g00642(.dina(n897), .dinb(n894), .dout(n898));
  jand g00643(.dina(n898), .dinb(n893), .dout(n899));
  jxor g00644(.dina(n899), .dinb(a11 ), .dout(n900));
  jnot g00645(.din(n900), .dout(n901));
  jnot g00646(.din(n818), .dout(n902));
  jand g00647(.dina(n720), .dinb(a14 ), .dout(n903));
  jand g00648(.dina(n903), .dinb(n902), .dout(n904));
  jnot g00649(.din(n904), .dout(n905));
  jand g00650(.dina(n905), .dinb(a14 ), .dout(n906));
  jor  g00651(.dina(n812), .dinb(n808), .dout(n907));
  jor  g00652(.dina(n907), .dinb(n718), .dout(n908));
  jnot g00653(.din(n908), .dout(n909));
  jand g00654(.dina(n909), .dinb(b0 ), .dout(n910));
  jand g00655(.dina(n809), .dinb(b2 ), .dout(n911));
  jand g00656(.dina(n813), .dinb(b1 ), .dout(n912));
  jand g00657(.dina(n815), .dinb(n375), .dout(n913));
  jor  g00658(.dina(n913), .dinb(n912), .dout(n914));
  jor  g00659(.dina(n914), .dinb(n911), .dout(n915));
  jor  g00660(.dina(n915), .dinb(n910), .dout(n916));
  jxor g00661(.dina(n916), .dinb(n906), .dout(n917));
  jxor g00662(.dina(n917), .dinb(n901), .dout(n918));
  jxor g00663(.dina(n918), .dinb(n892), .dout(n919));
  jxor g00664(.dina(n919), .dinb(n889), .dout(n920));
  jnot g00665(.din(n920), .dout(n921));
  jxor g00666(.dina(n921), .dinb(n880), .dout(n922));
  jxor g00667(.dina(n922), .dinb(n877), .dout(n923));
  jnot g00668(.din(n923), .dout(n924));
  jxor g00669(.dina(n924), .dinb(n869), .dout(n925));
  jxor g00670(.dina(n925), .dinb(n864), .dout(n926));
  jxor g00671(.dina(n926), .dinb(n849), .dout(f14 ));
  jand g00672(.dina(n925), .dinb(n864), .dout(n928));
  jand g00673(.dina(n926), .dinb(n849), .dout(n929));
  jor  g00674(.dina(n929), .dinb(n928), .dout(n930));
  jand g00675(.dina(b14 ), .dinb(b13 ), .dout(n931));
  jand g00676(.dina(n853), .dinb(n852), .dout(n932));
  jor  g00677(.dina(n932), .dinb(n931), .dout(n933));
  jxor g00678(.dina(b15 ), .dinb(b14 ), .dout(n934));
  jnot g00679(.din(n934), .dout(n935));
  jxor g00680(.dina(n935), .dinb(n933), .dout(n936));
  jor  g00681(.dina(n936), .dinb(n264), .dout(n937));
  jor  g00682(.dina(n284), .dinb(n778), .dout(n938));
  jnot g00683(.din(b15 ), .dout(n939));
  jor  g00684(.dina(n269), .dinb(n939), .dout(n940));
  jor  g00685(.dina(n271), .dinb(n858), .dout(n941));
  jand g00686(.dina(n941), .dinb(n940), .dout(n942));
  jand g00687(.dina(n942), .dinb(n938), .dout(n943));
  jand g00688(.dina(n943), .dinb(n937), .dout(n944));
  jxor g00689(.dina(n944), .dinb(n260), .dout(n945));
  jnot g00690(.din(n877), .dout(n946));
  jand g00691(.dina(n922), .dinb(n946), .dout(n947));
  jand g00692(.dina(n924), .dinb(n869), .dout(n948));
  jor  g00693(.dina(n948), .dinb(n947), .dout(n949));
  jor  g00694(.dina(n755), .dinb(n402), .dout(n950));
  jor  g00695(.dina(n371), .dinb(n627), .dout(n951));
  jor  g00696(.dina(n405), .dinb(n647), .dout(n952));
  jor  g00697(.dina(n332), .dinb(n758), .dout(n953));
  jand g00698(.dina(n953), .dinb(n952), .dout(n954));
  jand g00699(.dina(n954), .dinb(n951), .dout(n955));
  jand g00700(.dina(n955), .dinb(n950), .dout(n956));
  jxor g00701(.dina(n956), .dinb(a5 ), .dout(n957));
  jand g00702(.dina(n919), .dinb(n889), .dout(n958));
  jnot g00703(.din(n958), .dout(n959));
  jor  g00704(.dina(n921), .dinb(n880), .dout(n960));
  jand g00705(.dina(n960), .dinb(n959), .dout(n961));
  jor  g00706(.dina(n561), .dinb(n528), .dout(n962));
  jor  g00707(.dina(n490), .dinb(n431), .dout(n963));
  jor  g00708(.dina(n531), .dinb(n512), .dout(n964));
  jor  g00709(.dina(n533), .dinb(n564), .dout(n965));
  jand g00710(.dina(n965), .dinb(n964), .dout(n966));
  jand g00711(.dina(n966), .dinb(n963), .dout(n967));
  jand g00712(.dina(n967), .dinb(n962), .dout(n968));
  jxor g00713(.dina(n968), .dinb(a8 ), .dout(n969));
  jnot g00714(.din(n969), .dout(n970));
  jand g00715(.dina(n917), .dinb(n901), .dout(n971));
  jand g00716(.dina(n918), .dinb(n892), .dout(n972));
  jor  g00717(.dina(n972), .dinb(n971), .dout(n973));
  jnot g00718(.din(n815), .dout(n974));
  jor  g00719(.dina(n974), .dinb(n296), .dout(n975));
  jor  g00720(.dina(n908), .dinb(n267), .dout(n976));
  jnot g00721(.din(n813), .dout(n977));
  jor  g00722(.dina(n977), .dinb(n279), .dout(n978));
  jnot g00723(.din(n809), .dout(n979));
  jor  g00724(.dina(n979), .dinb(n299), .dout(n980));
  jand g00725(.dina(n980), .dinb(n978), .dout(n981));
  jand g00726(.dina(n981), .dinb(n976), .dout(n982));
  jand g00727(.dina(n982), .dinb(n975), .dout(n983));
  jxor g00728(.dina(n983), .dinb(a14 ), .dout(n984));
  jnot g00729(.din(n984), .dout(n985));
  jxor g00730(.dina(a15 ), .dinb(a14 ), .dout(n986));
  jand g00731(.dina(n986), .dinb(b0 ), .dout(n987));
  jnot g00732(.din(n987), .dout(n988));
  jor  g00733(.dina(n916), .dinb(n905), .dout(n989));
  jxor g00734(.dina(n989), .dinb(n988), .dout(n990));
  jxor g00735(.dina(n990), .dinb(n985), .dout(n991));
  jnot g00736(.din(n991), .dout(n992));
  jor  g00737(.dina(n706), .dinb(n392), .dout(n993));
  jor  g00738(.dina(n683), .dinb(n322), .dout(n994));
  jor  g00739(.dina(n709), .dinb(n357), .dout(n995));
  jor  g00740(.dina(n711), .dinb(n395), .dout(n996));
  jand g00741(.dina(n996), .dinb(n995), .dout(n997));
  jand g00742(.dina(n997), .dinb(n994), .dout(n998));
  jand g00743(.dina(n998), .dinb(n993), .dout(n999));
  jxor g00744(.dina(n999), .dinb(a11 ), .dout(n1000));
  jxor g00745(.dina(n1000), .dinb(n992), .dout(n1001));
  jxor g00746(.dina(n1001), .dinb(n973), .dout(n1002));
  jxor g00747(.dina(n1002), .dinb(n970), .dout(n1003));
  jnot g00748(.din(n1003), .dout(n1004));
  jxor g00749(.dina(n1004), .dinb(n961), .dout(n1005));
  jxor g00750(.dina(n1005), .dinb(n957), .dout(n1006));
  jnot g00751(.din(n1006), .dout(n1007));
  jxor g00752(.dina(n1007), .dinb(n949), .dout(n1008));
  jxor g00753(.dina(n1008), .dinb(n945), .dout(n1009));
  jxor g00754(.dina(n1009), .dinb(n930), .dout(f15 ));
  jand g00755(.dina(n1008), .dinb(n945), .dout(n1011));
  jand g00756(.dina(n1009), .dinb(n930), .dout(n1012));
  jor  g00757(.dina(n1012), .dinb(n1011), .dout(n1013));
  jand g00758(.dina(b15 ), .dinb(b14 ), .dout(n1014));
  jand g00759(.dina(n934), .dinb(n933), .dout(n1015));
  jor  g00760(.dina(n1015), .dinb(n1014), .dout(n1016));
  jxor g00761(.dina(b16 ), .dinb(b15 ), .dout(n1017));
  jnot g00762(.din(n1017), .dout(n1018));
  jxor g00763(.dina(n1018), .dinb(n1016), .dout(n1019));
  jor  g00764(.dina(n1019), .dinb(n264), .dout(n1020));
  jor  g00765(.dina(n284), .dinb(n858), .dout(n1021));
  jnot g00766(.din(b16 ), .dout(n1022));
  jor  g00767(.dina(n269), .dinb(n1022), .dout(n1023));
  jor  g00768(.dina(n271), .dinb(n939), .dout(n1024));
  jand g00769(.dina(n1024), .dinb(n1023), .dout(n1025));
  jand g00770(.dina(n1025), .dinb(n1021), .dout(n1026));
  jand g00771(.dina(n1026), .dinb(n1020), .dout(n1027));
  jxor g00772(.dina(n1027), .dinb(n260), .dout(n1028));
  jnot g00773(.din(n957), .dout(n1029));
  jand g00774(.dina(n1005), .dinb(n1029), .dout(n1030));
  jand g00775(.dina(n1007), .dinb(n949), .dout(n1031));
  jor  g00776(.dina(n1031), .dinb(n1030), .dout(n1032));
  jor  g00777(.dina(n775), .dinb(n402), .dout(n1033));
  jor  g00778(.dina(n371), .dinb(n647), .dout(n1034));
  jor  g00779(.dina(n405), .dinb(n758), .dout(n1035));
  jor  g00780(.dina(n332), .dinb(n778), .dout(n1036));
  jand g00781(.dina(n1036), .dinb(n1035), .dout(n1037));
  jand g00782(.dina(n1037), .dinb(n1034), .dout(n1038));
  jand g00783(.dina(n1038), .dinb(n1033), .dout(n1039));
  jxor g00784(.dina(n1039), .dinb(a5 ), .dout(n1040));
  jand g00785(.dina(n1002), .dinb(n970), .dout(n1041));
  jnot g00786(.din(n1041), .dout(n1042));
  jor  g00787(.dina(n1004), .dinb(n961), .dout(n1043));
  jand g00788(.dina(n1043), .dinb(n1042), .dout(n1044));
  jor  g00789(.dina(n624), .dinb(n528), .dout(n1045));
  jor  g00790(.dina(n490), .dinb(n512), .dout(n1046));
  jor  g00791(.dina(n531), .dinb(n564), .dout(n1047));
  jor  g00792(.dina(n533), .dinb(n627), .dout(n1048));
  jand g00793(.dina(n1048), .dinb(n1047), .dout(n1049));
  jand g00794(.dina(n1049), .dinb(n1046), .dout(n1050));
  jand g00795(.dina(n1050), .dinb(n1045), .dout(n1051));
  jxor g00796(.dina(n1051), .dinb(a8 ), .dout(n1052));
  jnot g00797(.din(n1052), .dout(n1053));
  jor  g00798(.dina(n1000), .dinb(n992), .dout(n1054));
  jand g00799(.dina(n1001), .dinb(n973), .dout(n1055));
  jnot g00800(.din(n1055), .dout(n1056));
  jand g00801(.dina(n1056), .dinb(n1054), .dout(n1057));
  jnot g00802(.din(n1057), .dout(n1058));
  jor  g00803(.dina(n706), .dinb(n428), .dout(n1059));
  jor  g00804(.dina(n683), .dinb(n357), .dout(n1060));
  jor  g00805(.dina(n709), .dinb(n395), .dout(n1061));
  jor  g00806(.dina(n711), .dinb(n431), .dout(n1062));
  jand g00807(.dina(n1062), .dinb(n1061), .dout(n1063));
  jand g00808(.dina(n1063), .dinb(n1060), .dout(n1064));
  jand g00809(.dina(n1064), .dinb(n1059), .dout(n1065));
  jxor g00810(.dina(n1065), .dinb(a11 ), .dout(n1066));
  jnot g00811(.din(n1066), .dout(n1067));
  jnot g00812(.din(n989), .dout(n1068));
  jand g00813(.dina(n1068), .dinb(n987), .dout(n1069));
  jand g00814(.dina(n990), .dinb(n985), .dout(n1070));
  jor  g00815(.dina(n1070), .dinb(n1069), .dout(n1071));
  jor  g00816(.dina(n974), .dinb(n319), .dout(n1072));
  jor  g00817(.dina(n908), .dinb(n279), .dout(n1073));
  jor  g00818(.dina(n977), .dinb(n299), .dout(n1074));
  jor  g00819(.dina(n979), .dinb(n322), .dout(n1075));
  jand g00820(.dina(n1075), .dinb(n1074), .dout(n1076));
  jand g00821(.dina(n1076), .dinb(n1073), .dout(n1077));
  jand g00822(.dina(n1077), .dinb(n1072), .dout(n1078));
  jxor g00823(.dina(n1078), .dinb(a14 ), .dout(n1079));
  jnot g00824(.din(n1079), .dout(n1080));
  jand g00825(.dina(n987), .dinb(a17 ), .dout(n1081));
  jxor g00826(.dina(a17 ), .dinb(a16 ), .dout(n1082));
  jnot g00827(.din(n1082), .dout(n1083));
  jand g00828(.dina(n1083), .dinb(n986), .dout(n1084));
  jand g00829(.dina(n1084), .dinb(b1 ), .dout(n1085));
  jnot g00830(.din(n986), .dout(n1086));
  jxor g00831(.dina(a16 ), .dinb(a15 ), .dout(n1087));
  jand g00832(.dina(n1087), .dinb(n1086), .dout(n1088));
  jand g00833(.dina(n1088), .dinb(b0 ), .dout(n1089));
  jand g00834(.dina(n1082), .dinb(n986), .dout(n1090));
  jand g00835(.dina(n1090), .dinb(n338), .dout(n1091));
  jor  g00836(.dina(n1091), .dinb(n1089), .dout(n1092));
  jor  g00837(.dina(n1092), .dinb(n1085), .dout(n1093));
  jxor g00838(.dina(n1093), .dinb(n1081), .dout(n1094));
  jxor g00839(.dina(n1094), .dinb(n1080), .dout(n1095));
  jxor g00840(.dina(n1095), .dinb(n1071), .dout(n1096));
  jxor g00841(.dina(n1096), .dinb(n1067), .dout(n1097));
  jxor g00842(.dina(n1097), .dinb(n1058), .dout(n1098));
  jxor g00843(.dina(n1098), .dinb(n1053), .dout(n1099));
  jnot g00844(.din(n1099), .dout(n1100));
  jxor g00845(.dina(n1100), .dinb(n1044), .dout(n1101));
  jxor g00846(.dina(n1101), .dinb(n1040), .dout(n1102));
  jnot g00847(.din(n1102), .dout(n1103));
  jxor g00848(.dina(n1103), .dinb(n1032), .dout(n1104));
  jxor g00849(.dina(n1104), .dinb(n1028), .dout(n1105));
  jxor g00850(.dina(n1105), .dinb(n1013), .dout(f16 ));
  jand g00851(.dina(n1104), .dinb(n1028), .dout(n1107));
  jand g00852(.dina(n1105), .dinb(n1013), .dout(n1108));
  jor  g00853(.dina(n1108), .dinb(n1107), .dout(n1109));
  jnot g00854(.din(n1040), .dout(n1110));
  jand g00855(.dina(n1101), .dinb(n1110), .dout(n1111));
  jand g00856(.dina(n1103), .dinb(n1032), .dout(n1112));
  jor  g00857(.dina(n1112), .dinb(n1111), .dout(n1113));
  jor  g00858(.dina(n855), .dinb(n402), .dout(n1114));
  jor  g00859(.dina(n371), .dinb(n758), .dout(n1115));
  jor  g00860(.dina(n405), .dinb(n778), .dout(n1116));
  jor  g00861(.dina(n332), .dinb(n858), .dout(n1117));
  jand g00862(.dina(n1117), .dinb(n1116), .dout(n1118));
  jand g00863(.dina(n1118), .dinb(n1115), .dout(n1119));
  jand g00864(.dina(n1119), .dinb(n1114), .dout(n1120));
  jxor g00865(.dina(n1120), .dinb(a5 ), .dout(n1121));
  jand g00866(.dina(n1098), .dinb(n1053), .dout(n1122));
  jnot g00867(.din(n1122), .dout(n1123));
  jor  g00868(.dina(n1100), .dinb(n1044), .dout(n1124));
  jand g00869(.dina(n1124), .dinb(n1123), .dout(n1125));
  jor  g00870(.dina(n644), .dinb(n528), .dout(n1126));
  jor  g00871(.dina(n490), .dinb(n564), .dout(n1127));
  jor  g00872(.dina(n531), .dinb(n627), .dout(n1128));
  jor  g00873(.dina(n533), .dinb(n647), .dout(n1129));
  jand g00874(.dina(n1129), .dinb(n1128), .dout(n1130));
  jand g00875(.dina(n1130), .dinb(n1127), .dout(n1131));
  jand g00876(.dina(n1131), .dinb(n1126), .dout(n1132));
  jxor g00877(.dina(n1132), .dinb(a8 ), .dout(n1133));
  jnot g00878(.din(n1133), .dout(n1134));
  jand g00879(.dina(n1096), .dinb(n1067), .dout(n1135));
  jand g00880(.dina(n1097), .dinb(n1058), .dout(n1136));
  jor  g00881(.dina(n1136), .dinb(n1135), .dout(n1137));
  jor  g00882(.dina(n706), .dinb(n509), .dout(n1138));
  jor  g00883(.dina(n683), .dinb(n395), .dout(n1139));
  jor  g00884(.dina(n709), .dinb(n431), .dout(n1140));
  jor  g00885(.dina(n711), .dinb(n512), .dout(n1141));
  jand g00886(.dina(n1141), .dinb(n1140), .dout(n1142));
  jand g00887(.dina(n1142), .dinb(n1139), .dout(n1143));
  jand g00888(.dina(n1143), .dinb(n1138), .dout(n1144));
  jxor g00889(.dina(n1144), .dinb(a11 ), .dout(n1145));
  jnot g00890(.din(n1145), .dout(n1146));
  jand g00891(.dina(n1094), .dinb(n1080), .dout(n1147));
  jand g00892(.dina(n1095), .dinb(n1071), .dout(n1148));
  jor  g00893(.dina(n1148), .dinb(n1147), .dout(n1149));
  jor  g00894(.dina(n974), .dinb(n354), .dout(n1150));
  jor  g00895(.dina(n908), .dinb(n299), .dout(n1151));
  jor  g00896(.dina(n977), .dinb(n322), .dout(n1152));
  jor  g00897(.dina(n979), .dinb(n357), .dout(n1153));
  jand g00898(.dina(n1153), .dinb(n1152), .dout(n1154));
  jand g00899(.dina(n1154), .dinb(n1151), .dout(n1155));
  jand g00900(.dina(n1155), .dinb(n1150), .dout(n1156));
  jxor g00901(.dina(n1156), .dinb(a14 ), .dout(n1157));
  jnot g00902(.din(n1157), .dout(n1158));
  jnot g00903(.din(n1093), .dout(n1159));
  jand g00904(.dina(n988), .dinb(a17 ), .dout(n1160));
  jand g00905(.dina(n1160), .dinb(n1159), .dout(n1161));
  jnot g00906(.din(n1161), .dout(n1162));
  jand g00907(.dina(n1162), .dinb(a17 ), .dout(n1163));
  jor  g00908(.dina(n1087), .dinb(n1083), .dout(n1164));
  jor  g00909(.dina(n1164), .dinb(n986), .dout(n1165));
  jnot g00910(.din(n1165), .dout(n1166));
  jand g00911(.dina(n1166), .dinb(b0 ), .dout(n1167));
  jand g00912(.dina(n1084), .dinb(b2 ), .dout(n1168));
  jand g00913(.dina(n1088), .dinb(b1 ), .dout(n1169));
  jand g00914(.dina(n1090), .dinb(n375), .dout(n1170));
  jor  g00915(.dina(n1170), .dinb(n1169), .dout(n1171));
  jor  g00916(.dina(n1171), .dinb(n1168), .dout(n1172));
  jor  g00917(.dina(n1172), .dinb(n1167), .dout(n1173));
  jxor g00918(.dina(n1173), .dinb(n1163), .dout(n1174));
  jxor g00919(.dina(n1174), .dinb(n1158), .dout(n1175));
  jxor g00920(.dina(n1175), .dinb(n1149), .dout(n1176));
  jxor g00921(.dina(n1176), .dinb(n1146), .dout(n1177));
  jxor g00922(.dina(n1177), .dinb(n1137), .dout(n1178));
  jxor g00923(.dina(n1178), .dinb(n1134), .dout(n1179));
  jnot g00924(.din(n1179), .dout(n1180));
  jxor g00925(.dina(n1180), .dinb(n1125), .dout(n1181));
  jxor g00926(.dina(n1181), .dinb(n1121), .dout(n1182));
  jnot g00927(.din(n1182), .dout(n1183));
  jxor g00928(.dina(n1183), .dinb(n1113), .dout(n1184));
  jand g00929(.dina(b16 ), .dinb(b15 ), .dout(n1185));
  jand g00930(.dina(n1017), .dinb(n1016), .dout(n1186));
  jor  g00931(.dina(n1186), .dinb(n1185), .dout(n1187));
  jxor g00932(.dina(b17 ), .dinb(b16 ), .dout(n1188));
  jnot g00933(.din(n1188), .dout(n1189));
  jxor g00934(.dina(n1189), .dinb(n1187), .dout(n1190));
  jor  g00935(.dina(n1190), .dinb(n264), .dout(n1191));
  jor  g00936(.dina(n284), .dinb(n939), .dout(n1192));
  jnot g00937(.din(b17 ), .dout(n1193));
  jor  g00938(.dina(n269), .dinb(n1193), .dout(n1194));
  jor  g00939(.dina(n271), .dinb(n1022), .dout(n1195));
  jand g00940(.dina(n1195), .dinb(n1194), .dout(n1196));
  jand g00941(.dina(n1196), .dinb(n1192), .dout(n1197));
  jand g00942(.dina(n1197), .dinb(n1191), .dout(n1198));
  jxor g00943(.dina(n1198), .dinb(n260), .dout(n1199));
  jxor g00944(.dina(n1199), .dinb(n1184), .dout(n1200));
  jxor g00945(.dina(n1200), .dinb(n1109), .dout(f17 ));
  jand g00946(.dina(n1199), .dinb(n1184), .dout(n1202));
  jand g00947(.dina(n1200), .dinb(n1109), .dout(n1203));
  jor  g00948(.dina(n1203), .dinb(n1202), .dout(n1204));
  jnot g00949(.din(n1121), .dout(n1205));
  jand g00950(.dina(n1181), .dinb(n1205), .dout(n1206));
  jand g00951(.dina(n1183), .dinb(n1113), .dout(n1207));
  jor  g00952(.dina(n1207), .dinb(n1206), .dout(n1208));
  jor  g00953(.dina(n936), .dinb(n402), .dout(n1209));
  jor  g00954(.dina(n371), .dinb(n778), .dout(n1210));
  jor  g00955(.dina(n405), .dinb(n858), .dout(n1211));
  jor  g00956(.dina(n332), .dinb(n939), .dout(n1212));
  jand g00957(.dina(n1212), .dinb(n1211), .dout(n1213));
  jand g00958(.dina(n1213), .dinb(n1210), .dout(n1214));
  jand g00959(.dina(n1214), .dinb(n1209), .dout(n1215));
  jxor g00960(.dina(n1215), .dinb(a5 ), .dout(n1216));
  jand g00961(.dina(n1178), .dinb(n1134), .dout(n1217));
  jnot g00962(.din(n1217), .dout(n1218));
  jor  g00963(.dina(n1180), .dinb(n1125), .dout(n1219));
  jand g00964(.dina(n1219), .dinb(n1218), .dout(n1220));
  jor  g00965(.dina(n755), .dinb(n528), .dout(n1221));
  jor  g00966(.dina(n490), .dinb(n627), .dout(n1222));
  jor  g00967(.dina(n531), .dinb(n647), .dout(n1223));
  jor  g00968(.dina(n533), .dinb(n758), .dout(n1224));
  jand g00969(.dina(n1224), .dinb(n1223), .dout(n1225));
  jand g00970(.dina(n1225), .dinb(n1222), .dout(n1226));
  jand g00971(.dina(n1226), .dinb(n1221), .dout(n1227));
  jxor g00972(.dina(n1227), .dinb(a8 ), .dout(n1228));
  jnot g00973(.din(n1228), .dout(n1229));
  jand g00974(.dina(n1176), .dinb(n1146), .dout(n1230));
  jand g00975(.dina(n1177), .dinb(n1137), .dout(n1231));
  jor  g00976(.dina(n1231), .dinb(n1230), .dout(n1232));
  jor  g00977(.dina(n706), .dinb(n561), .dout(n1233));
  jor  g00978(.dina(n683), .dinb(n431), .dout(n1234));
  jor  g00979(.dina(n709), .dinb(n512), .dout(n1235));
  jor  g00980(.dina(n711), .dinb(n564), .dout(n1236));
  jand g00981(.dina(n1236), .dinb(n1235), .dout(n1237));
  jand g00982(.dina(n1237), .dinb(n1234), .dout(n1238));
  jand g00983(.dina(n1238), .dinb(n1233), .dout(n1239));
  jxor g00984(.dina(n1239), .dinb(a11 ), .dout(n1240));
  jnot g00985(.din(n1240), .dout(n1241));
  jand g00986(.dina(n1174), .dinb(n1158), .dout(n1242));
  jand g00987(.dina(n1175), .dinb(n1149), .dout(n1243));
  jor  g00988(.dina(n1243), .dinb(n1242), .dout(n1244));
  jnot g00989(.din(n1090), .dout(n1245));
  jor  g00990(.dina(n1245), .dinb(n296), .dout(n1246));
  jor  g00991(.dina(n1165), .dinb(n267), .dout(n1247));
  jnot g00992(.din(n1088), .dout(n1248));
  jor  g00993(.dina(n1248), .dinb(n279), .dout(n1249));
  jnot g00994(.din(n1084), .dout(n1250));
  jor  g00995(.dina(n1250), .dinb(n299), .dout(n1251));
  jand g00996(.dina(n1251), .dinb(n1249), .dout(n1252));
  jand g00997(.dina(n1252), .dinb(n1247), .dout(n1253));
  jand g00998(.dina(n1253), .dinb(n1246), .dout(n1254));
  jxor g00999(.dina(n1254), .dinb(a17 ), .dout(n1255));
  jnot g01000(.din(n1255), .dout(n1256));
  jxor g01001(.dina(a18 ), .dinb(a17 ), .dout(n1257));
  jand g01002(.dina(n1257), .dinb(b0 ), .dout(n1258));
  jnot g01003(.din(n1258), .dout(n1259));
  jor  g01004(.dina(n1173), .dinb(n1162), .dout(n1260));
  jxor g01005(.dina(n1260), .dinb(n1259), .dout(n1261));
  jxor g01006(.dina(n1261), .dinb(n1256), .dout(n1262));
  jnot g01007(.din(n1262), .dout(n1263));
  jor  g01008(.dina(n974), .dinb(n392), .dout(n1264));
  jor  g01009(.dina(n908), .dinb(n322), .dout(n1265));
  jor  g01010(.dina(n977), .dinb(n357), .dout(n1266));
  jor  g01011(.dina(n979), .dinb(n395), .dout(n1267));
  jand g01012(.dina(n1267), .dinb(n1266), .dout(n1268));
  jand g01013(.dina(n1268), .dinb(n1265), .dout(n1269));
  jand g01014(.dina(n1269), .dinb(n1264), .dout(n1270));
  jxor g01015(.dina(n1270), .dinb(a14 ), .dout(n1271));
  jxor g01016(.dina(n1271), .dinb(n1263), .dout(n1272));
  jxor g01017(.dina(n1272), .dinb(n1244), .dout(n1273));
  jxor g01018(.dina(n1273), .dinb(n1241), .dout(n1274));
  jxor g01019(.dina(n1274), .dinb(n1232), .dout(n1275));
  jxor g01020(.dina(n1275), .dinb(n1229), .dout(n1276));
  jnot g01021(.din(n1276), .dout(n1277));
  jxor g01022(.dina(n1277), .dinb(n1220), .dout(n1278));
  jxor g01023(.dina(n1278), .dinb(n1216), .dout(n1279));
  jnot g01024(.din(n1279), .dout(n1280));
  jxor g01025(.dina(n1280), .dinb(n1208), .dout(n1281));
  jand g01026(.dina(b17 ), .dinb(b16 ), .dout(n1282));
  jand g01027(.dina(n1188), .dinb(n1187), .dout(n1283));
  jor  g01028(.dina(n1283), .dinb(n1282), .dout(n1284));
  jxor g01029(.dina(b18 ), .dinb(b17 ), .dout(n1285));
  jnot g01030(.din(n1285), .dout(n1286));
  jxor g01031(.dina(n1286), .dinb(n1284), .dout(n1287));
  jor  g01032(.dina(n1287), .dinb(n264), .dout(n1288));
  jor  g01033(.dina(n284), .dinb(n1022), .dout(n1289));
  jnot g01034(.din(b18 ), .dout(n1290));
  jor  g01035(.dina(n269), .dinb(n1290), .dout(n1291));
  jor  g01036(.dina(n271), .dinb(n1193), .dout(n1292));
  jand g01037(.dina(n1292), .dinb(n1291), .dout(n1293));
  jand g01038(.dina(n1293), .dinb(n1289), .dout(n1294));
  jand g01039(.dina(n1294), .dinb(n1288), .dout(n1295));
  jxor g01040(.dina(n1295), .dinb(n260), .dout(n1296));
  jxor g01041(.dina(n1296), .dinb(n1281), .dout(n1297));
  jxor g01042(.dina(n1297), .dinb(n1204), .dout(f18 ));
  jand g01043(.dina(n1296), .dinb(n1281), .dout(n1299));
  jand g01044(.dina(n1297), .dinb(n1204), .dout(n1300));
  jor  g01045(.dina(n1300), .dinb(n1299), .dout(n1301));
  jnot g01046(.din(n1216), .dout(n1302));
  jand g01047(.dina(n1278), .dinb(n1302), .dout(n1303));
  jand g01048(.dina(n1280), .dinb(n1208), .dout(n1304));
  jor  g01049(.dina(n1304), .dinb(n1303), .dout(n1305));
  jand g01050(.dina(n1273), .dinb(n1241), .dout(n1306));
  jand g01051(.dina(n1274), .dinb(n1232), .dout(n1307));
  jor  g01052(.dina(n1307), .dinb(n1306), .dout(n1308));
  jor  g01053(.dina(n1271), .dinb(n1263), .dout(n1309));
  jand g01054(.dina(n1272), .dinb(n1244), .dout(n1310));
  jnot g01055(.din(n1310), .dout(n1311));
  jand g01056(.dina(n1311), .dinb(n1309), .dout(n1312));
  jnot g01057(.din(n1312), .dout(n1313));
  jor  g01058(.dina(n974), .dinb(n428), .dout(n1314));
  jor  g01059(.dina(n908), .dinb(n357), .dout(n1315));
  jor  g01060(.dina(n977), .dinb(n395), .dout(n1316));
  jor  g01061(.dina(n979), .dinb(n431), .dout(n1317));
  jand g01062(.dina(n1317), .dinb(n1316), .dout(n1318));
  jand g01063(.dina(n1318), .dinb(n1315), .dout(n1319));
  jand g01064(.dina(n1319), .dinb(n1314), .dout(n1320));
  jxor g01065(.dina(n1320), .dinb(a14 ), .dout(n1321));
  jnot g01066(.din(n1321), .dout(n1322));
  jnot g01067(.din(n1260), .dout(n1323));
  jand g01068(.dina(n1323), .dinb(n1258), .dout(n1324));
  jand g01069(.dina(n1261), .dinb(n1256), .dout(n1325));
  jor  g01070(.dina(n1325), .dinb(n1324), .dout(n1326));
  jor  g01071(.dina(n1245), .dinb(n319), .dout(n1327));
  jor  g01072(.dina(n1165), .dinb(n279), .dout(n1328));
  jor  g01073(.dina(n1248), .dinb(n299), .dout(n1329));
  jor  g01074(.dina(n1250), .dinb(n322), .dout(n1330));
  jand g01075(.dina(n1330), .dinb(n1329), .dout(n1331));
  jand g01076(.dina(n1331), .dinb(n1328), .dout(n1332));
  jand g01077(.dina(n1332), .dinb(n1327), .dout(n1333));
  jxor g01078(.dina(n1333), .dinb(a17 ), .dout(n1334));
  jnot g01079(.din(n1334), .dout(n1335));
  jand g01080(.dina(n1258), .dinb(a20 ), .dout(n1336));
  jxor g01081(.dina(a20 ), .dinb(a19 ), .dout(n1337));
  jnot g01082(.din(n1337), .dout(n1338));
  jand g01083(.dina(n1338), .dinb(n1257), .dout(n1339));
  jand g01084(.dina(n1339), .dinb(b1 ), .dout(n1340));
  jnot g01085(.din(n1257), .dout(n1341));
  jxor g01086(.dina(a19 ), .dinb(a18 ), .dout(n1342));
  jand g01087(.dina(n1342), .dinb(n1341), .dout(n1343));
  jand g01088(.dina(n1343), .dinb(b0 ), .dout(n1344));
  jand g01089(.dina(n1337), .dinb(n1257), .dout(n1345));
  jand g01090(.dina(n1345), .dinb(n338), .dout(n1346));
  jor  g01091(.dina(n1346), .dinb(n1344), .dout(n1347));
  jor  g01092(.dina(n1347), .dinb(n1340), .dout(n1348));
  jxor g01093(.dina(n1348), .dinb(n1336), .dout(n1349));
  jxor g01094(.dina(n1349), .dinb(n1335), .dout(n1350));
  jxor g01095(.dina(n1350), .dinb(n1326), .dout(n1351));
  jxor g01096(.dina(n1351), .dinb(n1322), .dout(n1352));
  jxor g01097(.dina(n1352), .dinb(n1313), .dout(n1353));
  jnot g01098(.din(n1353), .dout(n1354));
  jor  g01099(.dina(n624), .dinb(n706), .dout(n1355));
  jor  g01100(.dina(n683), .dinb(n512), .dout(n1356));
  jor  g01101(.dina(n709), .dinb(n564), .dout(n1357));
  jor  g01102(.dina(n711), .dinb(n627), .dout(n1358));
  jand g01103(.dina(n1358), .dinb(n1357), .dout(n1359));
  jand g01104(.dina(n1359), .dinb(n1356), .dout(n1360));
  jand g01105(.dina(n1360), .dinb(n1355), .dout(n1361));
  jxor g01106(.dina(n1361), .dinb(a11 ), .dout(n1362));
  jxor g01107(.dina(n1362), .dinb(n1354), .dout(n1363));
  jxor g01108(.dina(n1363), .dinb(n1308), .dout(n1364));
  jnot g01109(.din(n1364), .dout(n1365));
  jor  g01110(.dina(n775), .dinb(n528), .dout(n1366));
  jor  g01111(.dina(n490), .dinb(n647), .dout(n1367));
  jor  g01112(.dina(n531), .dinb(n758), .dout(n1368));
  jor  g01113(.dina(n533), .dinb(n778), .dout(n1369));
  jand g01114(.dina(n1369), .dinb(n1368), .dout(n1370));
  jand g01115(.dina(n1370), .dinb(n1367), .dout(n1371));
  jand g01116(.dina(n1371), .dinb(n1366), .dout(n1372));
  jxor g01117(.dina(n1372), .dinb(a8 ), .dout(n1373));
  jxor g01118(.dina(n1373), .dinb(n1365), .dout(n1374));
  jnot g01119(.din(n1374), .dout(n1375));
  jand g01120(.dina(n1275), .dinb(n1229), .dout(n1376));
  jnot g01121(.din(n1376), .dout(n1377));
  jor  g01122(.dina(n1277), .dinb(n1220), .dout(n1378));
  jand g01123(.dina(n1378), .dinb(n1377), .dout(n1379));
  jxor g01124(.dina(n1379), .dinb(n1375), .dout(n1380));
  jor  g01125(.dina(n1019), .dinb(n402), .dout(n1381));
  jor  g01126(.dina(n371), .dinb(n858), .dout(n1382));
  jor  g01127(.dina(n405), .dinb(n939), .dout(n1383));
  jor  g01128(.dina(n332), .dinb(n1022), .dout(n1384));
  jand g01129(.dina(n1384), .dinb(n1383), .dout(n1385));
  jand g01130(.dina(n1385), .dinb(n1382), .dout(n1386));
  jand g01131(.dina(n1386), .dinb(n1381), .dout(n1387));
  jxor g01132(.dina(n1387), .dinb(a5 ), .dout(n1388));
  jxor g01133(.dina(n1388), .dinb(n1380), .dout(n1389));
  jnot g01134(.din(n1389), .dout(n1390));
  jxor g01135(.dina(n1390), .dinb(n1305), .dout(n1391));
  jand g01136(.dina(b18 ), .dinb(b17 ), .dout(n1392));
  jand g01137(.dina(n1285), .dinb(n1284), .dout(n1393));
  jor  g01138(.dina(n1393), .dinb(n1392), .dout(n1394));
  jxor g01139(.dina(b19 ), .dinb(b18 ), .dout(n1395));
  jnot g01140(.din(n1395), .dout(n1396));
  jxor g01141(.dina(n1396), .dinb(n1394), .dout(n1397));
  jor  g01142(.dina(n1397), .dinb(n264), .dout(n1398));
  jor  g01143(.dina(n284), .dinb(n1193), .dout(n1399));
  jnot g01144(.din(b19 ), .dout(n1400));
  jor  g01145(.dina(n269), .dinb(n1400), .dout(n1401));
  jor  g01146(.dina(n271), .dinb(n1290), .dout(n1402));
  jand g01147(.dina(n1402), .dinb(n1401), .dout(n1403));
  jand g01148(.dina(n1403), .dinb(n1399), .dout(n1404));
  jand g01149(.dina(n1404), .dinb(n1398), .dout(n1405));
  jxor g01150(.dina(n1405), .dinb(n260), .dout(n1406));
  jxor g01151(.dina(n1406), .dinb(n1391), .dout(n1407));
  jxor g01152(.dina(n1407), .dinb(n1301), .dout(f19 ));
  jand g01153(.dina(n1406), .dinb(n1391), .dout(n1409));
  jand g01154(.dina(n1407), .dinb(n1301), .dout(n1410));
  jor  g01155(.dina(n1410), .dinb(n1409), .dout(n1411));
  jand g01156(.dina(b19 ), .dinb(b18 ), .dout(n1412));
  jand g01157(.dina(n1395), .dinb(n1394), .dout(n1413));
  jor  g01158(.dina(n1413), .dinb(n1412), .dout(n1414));
  jxor g01159(.dina(b20 ), .dinb(b19 ), .dout(n1415));
  jnot g01160(.din(n1415), .dout(n1416));
  jxor g01161(.dina(n1416), .dinb(n1414), .dout(n1417));
  jor  g01162(.dina(n1417), .dinb(n264), .dout(n1418));
  jor  g01163(.dina(n284), .dinb(n1290), .dout(n1419));
  jnot g01164(.din(b20 ), .dout(n1420));
  jor  g01165(.dina(n269), .dinb(n1420), .dout(n1421));
  jor  g01166(.dina(n271), .dinb(n1400), .dout(n1422));
  jand g01167(.dina(n1422), .dinb(n1421), .dout(n1423));
  jand g01168(.dina(n1423), .dinb(n1419), .dout(n1424));
  jand g01169(.dina(n1424), .dinb(n1418), .dout(n1425));
  jxor g01170(.dina(n1425), .dinb(n260), .dout(n1426));
  jnot g01171(.din(n1380), .dout(n1427));
  jor  g01172(.dina(n1388), .dinb(n1427), .dout(n1428));
  jnot g01173(.din(n1428), .dout(n1429));
  jand g01174(.dina(n1390), .dinb(n1305), .dout(n1430));
  jor  g01175(.dina(n1430), .dinb(n1429), .dout(n1431));
  jor  g01176(.dina(n1190), .dinb(n402), .dout(n1432));
  jor  g01177(.dina(n371), .dinb(n939), .dout(n1433));
  jor  g01178(.dina(n405), .dinb(n1022), .dout(n1434));
  jor  g01179(.dina(n332), .dinb(n1193), .dout(n1435));
  jand g01180(.dina(n1435), .dinb(n1434), .dout(n1436));
  jand g01181(.dina(n1436), .dinb(n1433), .dout(n1437));
  jand g01182(.dina(n1437), .dinb(n1432), .dout(n1438));
  jxor g01183(.dina(n1438), .dinb(a5 ), .dout(n1439));
  jnot g01184(.din(n1439), .dout(n1440));
  jor  g01185(.dina(n1373), .dinb(n1365), .dout(n1441));
  jor  g01186(.dina(n1379), .dinb(n1375), .dout(n1442));
  jand g01187(.dina(n1442), .dinb(n1441), .dout(n1443));
  jnot g01188(.din(n1443), .dout(n1444));
  jor  g01189(.dina(n1362), .dinb(n1354), .dout(n1445));
  jand g01190(.dina(n1363), .dinb(n1308), .dout(n1446));
  jnot g01191(.din(n1446), .dout(n1447));
  jand g01192(.dina(n1447), .dinb(n1445), .dout(n1448));
  jnot g01193(.din(n1448), .dout(n1449));
  jor  g01194(.dina(n644), .dinb(n706), .dout(n1450));
  jor  g01195(.dina(n683), .dinb(n564), .dout(n1451));
  jor  g01196(.dina(n709), .dinb(n627), .dout(n1452));
  jor  g01197(.dina(n711), .dinb(n647), .dout(n1453));
  jand g01198(.dina(n1453), .dinb(n1452), .dout(n1454));
  jand g01199(.dina(n1454), .dinb(n1451), .dout(n1455));
  jand g01200(.dina(n1455), .dinb(n1450), .dout(n1456));
  jxor g01201(.dina(n1456), .dinb(a11 ), .dout(n1457));
  jnot g01202(.din(n1457), .dout(n1458));
  jand g01203(.dina(n1351), .dinb(n1322), .dout(n1459));
  jand g01204(.dina(n1352), .dinb(n1313), .dout(n1460));
  jor  g01205(.dina(n1460), .dinb(n1459), .dout(n1461));
  jor  g01206(.dina(n974), .dinb(n509), .dout(n1462));
  jor  g01207(.dina(n908), .dinb(n395), .dout(n1463));
  jor  g01208(.dina(n977), .dinb(n431), .dout(n1464));
  jor  g01209(.dina(n979), .dinb(n512), .dout(n1465));
  jand g01210(.dina(n1465), .dinb(n1464), .dout(n1466));
  jand g01211(.dina(n1466), .dinb(n1463), .dout(n1467));
  jand g01212(.dina(n1467), .dinb(n1462), .dout(n1468));
  jxor g01213(.dina(n1468), .dinb(a14 ), .dout(n1469));
  jnot g01214(.din(n1469), .dout(n1470));
  jand g01215(.dina(n1349), .dinb(n1335), .dout(n1471));
  jand g01216(.dina(n1350), .dinb(n1326), .dout(n1472));
  jor  g01217(.dina(n1472), .dinb(n1471), .dout(n1473));
  jor  g01218(.dina(n1245), .dinb(n354), .dout(n1474));
  jor  g01219(.dina(n1165), .dinb(n299), .dout(n1475));
  jor  g01220(.dina(n1248), .dinb(n322), .dout(n1476));
  jor  g01221(.dina(n1250), .dinb(n357), .dout(n1477));
  jand g01222(.dina(n1477), .dinb(n1476), .dout(n1478));
  jand g01223(.dina(n1478), .dinb(n1475), .dout(n1479));
  jand g01224(.dina(n1479), .dinb(n1474), .dout(n1480));
  jxor g01225(.dina(n1480), .dinb(a17 ), .dout(n1481));
  jnot g01226(.din(n1481), .dout(n1482));
  jnot g01227(.din(n1348), .dout(n1483));
  jand g01228(.dina(n1259), .dinb(a20 ), .dout(n1484));
  jand g01229(.dina(n1484), .dinb(n1483), .dout(n1485));
  jnot g01230(.din(n1485), .dout(n1486));
  jand g01231(.dina(n1486), .dinb(a20 ), .dout(n1487));
  jor  g01232(.dina(n1342), .dinb(n1338), .dout(n1488));
  jor  g01233(.dina(n1488), .dinb(n1257), .dout(n1489));
  jnot g01234(.din(n1489), .dout(n1490));
  jand g01235(.dina(n1490), .dinb(b0 ), .dout(n1491));
  jand g01236(.dina(n1339), .dinb(b2 ), .dout(n1492));
  jand g01237(.dina(n1343), .dinb(b1 ), .dout(n1493));
  jand g01238(.dina(n1345), .dinb(n375), .dout(n1494));
  jor  g01239(.dina(n1494), .dinb(n1493), .dout(n1495));
  jor  g01240(.dina(n1495), .dinb(n1492), .dout(n1496));
  jor  g01241(.dina(n1496), .dinb(n1491), .dout(n1497));
  jxor g01242(.dina(n1497), .dinb(n1487), .dout(n1498));
  jxor g01243(.dina(n1498), .dinb(n1482), .dout(n1499));
  jxor g01244(.dina(n1499), .dinb(n1473), .dout(n1500));
  jxor g01245(.dina(n1500), .dinb(n1470), .dout(n1501));
  jxor g01246(.dina(n1501), .dinb(n1461), .dout(n1502));
  jxor g01247(.dina(n1502), .dinb(n1458), .dout(n1503));
  jxor g01248(.dina(n1503), .dinb(n1449), .dout(n1504));
  jnot g01249(.din(n1504), .dout(n1505));
  jor  g01250(.dina(n855), .dinb(n528), .dout(n1506));
  jor  g01251(.dina(n490), .dinb(n758), .dout(n1507));
  jor  g01252(.dina(n531), .dinb(n778), .dout(n1508));
  jor  g01253(.dina(n533), .dinb(n858), .dout(n1509));
  jand g01254(.dina(n1509), .dinb(n1508), .dout(n1510));
  jand g01255(.dina(n1510), .dinb(n1507), .dout(n1511));
  jand g01256(.dina(n1511), .dinb(n1506), .dout(n1512));
  jxor g01257(.dina(n1512), .dinb(a8 ), .dout(n1513));
  jxor g01258(.dina(n1513), .dinb(n1505), .dout(n1514));
  jxor g01259(.dina(n1514), .dinb(n1444), .dout(n1515));
  jxor g01260(.dina(n1515), .dinb(n1440), .dout(n1516));
  jxor g01261(.dina(n1516), .dinb(n1431), .dout(n1517));
  jxor g01262(.dina(n1517), .dinb(n1426), .dout(n1518));
  jxor g01263(.dina(n1518), .dinb(n1411), .dout(f20 ));
  jand g01264(.dina(n1517), .dinb(n1426), .dout(n1520));
  jand g01265(.dina(n1518), .dinb(n1411), .dout(n1521));
  jor  g01266(.dina(n1521), .dinb(n1520), .dout(n1522));
  jand g01267(.dina(n1515), .dinb(n1440), .dout(n1523));
  jand g01268(.dina(n1516), .dinb(n1431), .dout(n1524));
  jor  g01269(.dina(n1524), .dinb(n1523), .dout(n1525));
  jor  g01270(.dina(n1513), .dinb(n1505), .dout(n1526));
  jnot g01271(.din(n1526), .dout(n1527));
  jand g01272(.dina(n1514), .dinb(n1444), .dout(n1528));
  jor  g01273(.dina(n1528), .dinb(n1527), .dout(n1529));
  jor  g01274(.dina(n936), .dinb(n528), .dout(n1530));
  jor  g01275(.dina(n490), .dinb(n778), .dout(n1531));
  jor  g01276(.dina(n531), .dinb(n858), .dout(n1532));
  jor  g01277(.dina(n533), .dinb(n939), .dout(n1533));
  jand g01278(.dina(n1533), .dinb(n1532), .dout(n1534));
  jand g01279(.dina(n1534), .dinb(n1531), .dout(n1535));
  jand g01280(.dina(n1535), .dinb(n1530), .dout(n1536));
  jxor g01281(.dina(n1536), .dinb(a8 ), .dout(n1537));
  jnot g01282(.din(n1537), .dout(n1538));
  jand g01283(.dina(n1502), .dinb(n1458), .dout(n1539));
  jand g01284(.dina(n1503), .dinb(n1449), .dout(n1540));
  jor  g01285(.dina(n1540), .dinb(n1539), .dout(n1541));
  jor  g01286(.dina(n755), .dinb(n706), .dout(n1542));
  jor  g01287(.dina(n683), .dinb(n627), .dout(n1543));
  jor  g01288(.dina(n709), .dinb(n647), .dout(n1544));
  jor  g01289(.dina(n711), .dinb(n758), .dout(n1545));
  jand g01290(.dina(n1545), .dinb(n1544), .dout(n1546));
  jand g01291(.dina(n1546), .dinb(n1543), .dout(n1547));
  jand g01292(.dina(n1547), .dinb(n1542), .dout(n1548));
  jxor g01293(.dina(n1548), .dinb(a11 ), .dout(n1549));
  jnot g01294(.din(n1549), .dout(n1550));
  jand g01295(.dina(n1500), .dinb(n1470), .dout(n1551));
  jand g01296(.dina(n1501), .dinb(n1461), .dout(n1552));
  jor  g01297(.dina(n1552), .dinb(n1551), .dout(n1553));
  jor  g01298(.dina(n974), .dinb(n561), .dout(n1554));
  jor  g01299(.dina(n908), .dinb(n431), .dout(n1555));
  jor  g01300(.dina(n977), .dinb(n512), .dout(n1556));
  jor  g01301(.dina(n979), .dinb(n564), .dout(n1557));
  jand g01302(.dina(n1557), .dinb(n1556), .dout(n1558));
  jand g01303(.dina(n1558), .dinb(n1555), .dout(n1559));
  jand g01304(.dina(n1559), .dinb(n1554), .dout(n1560));
  jxor g01305(.dina(n1560), .dinb(a14 ), .dout(n1561));
  jnot g01306(.din(n1561), .dout(n1562));
  jand g01307(.dina(n1498), .dinb(n1482), .dout(n1563));
  jand g01308(.dina(n1499), .dinb(n1473), .dout(n1564));
  jor  g01309(.dina(n1564), .dinb(n1563), .dout(n1565));
  jnot g01310(.din(n1345), .dout(n1566));
  jor  g01311(.dina(n1566), .dinb(n296), .dout(n1567));
  jor  g01312(.dina(n1489), .dinb(n267), .dout(n1568));
  jnot g01313(.din(n1343), .dout(n1569));
  jor  g01314(.dina(n1569), .dinb(n279), .dout(n1570));
  jnot g01315(.din(n1339), .dout(n1571));
  jor  g01316(.dina(n1571), .dinb(n299), .dout(n1572));
  jand g01317(.dina(n1572), .dinb(n1570), .dout(n1573));
  jand g01318(.dina(n1573), .dinb(n1568), .dout(n1574));
  jand g01319(.dina(n1574), .dinb(n1567), .dout(n1575));
  jxor g01320(.dina(n1575), .dinb(a20 ), .dout(n1576));
  jnot g01321(.din(n1576), .dout(n1577));
  jxor g01322(.dina(a21 ), .dinb(a20 ), .dout(n1578));
  jand g01323(.dina(n1578), .dinb(b0 ), .dout(n1579));
  jnot g01324(.din(n1579), .dout(n1580));
  jor  g01325(.dina(n1497), .dinb(n1486), .dout(n1581));
  jxor g01326(.dina(n1581), .dinb(n1580), .dout(n1582));
  jxor g01327(.dina(n1582), .dinb(n1577), .dout(n1583));
  jnot g01328(.din(n1583), .dout(n1584));
  jor  g01329(.dina(n1245), .dinb(n392), .dout(n1585));
  jor  g01330(.dina(n1165), .dinb(n322), .dout(n1586));
  jor  g01331(.dina(n1248), .dinb(n357), .dout(n1587));
  jor  g01332(.dina(n1250), .dinb(n395), .dout(n1588));
  jand g01333(.dina(n1588), .dinb(n1587), .dout(n1589));
  jand g01334(.dina(n1589), .dinb(n1586), .dout(n1590));
  jand g01335(.dina(n1590), .dinb(n1585), .dout(n1591));
  jxor g01336(.dina(n1591), .dinb(a17 ), .dout(n1592));
  jxor g01337(.dina(n1592), .dinb(n1584), .dout(n1593));
  jxor g01338(.dina(n1593), .dinb(n1565), .dout(n1594));
  jxor g01339(.dina(n1594), .dinb(n1562), .dout(n1595));
  jxor g01340(.dina(n1595), .dinb(n1553), .dout(n1596));
  jxor g01341(.dina(n1596), .dinb(n1550), .dout(n1597));
  jxor g01342(.dina(n1597), .dinb(n1541), .dout(n1598));
  jxor g01343(.dina(n1598), .dinb(n1538), .dout(n1599));
  jnot g01344(.din(n1599), .dout(n1600));
  jxor g01345(.dina(n1600), .dinb(n1529), .dout(n1601));
  jor  g01346(.dina(n1287), .dinb(n402), .dout(n1602));
  jor  g01347(.dina(n371), .dinb(n1022), .dout(n1603));
  jor  g01348(.dina(n405), .dinb(n1193), .dout(n1604));
  jor  g01349(.dina(n332), .dinb(n1290), .dout(n1605));
  jand g01350(.dina(n1605), .dinb(n1604), .dout(n1606));
  jand g01351(.dina(n1606), .dinb(n1603), .dout(n1607));
  jand g01352(.dina(n1607), .dinb(n1602), .dout(n1608));
  jxor g01353(.dina(n1608), .dinb(a5 ), .dout(n1609));
  jxor g01354(.dina(n1609), .dinb(n1601), .dout(n1610));
  jxor g01355(.dina(n1610), .dinb(n1525), .dout(n1611));
  jand g01356(.dina(b20 ), .dinb(b19 ), .dout(n1612));
  jand g01357(.dina(n1415), .dinb(n1414), .dout(n1613));
  jor  g01358(.dina(n1613), .dinb(n1612), .dout(n1614));
  jxor g01359(.dina(b21 ), .dinb(b20 ), .dout(n1615));
  jnot g01360(.din(n1615), .dout(n1616));
  jxor g01361(.dina(n1616), .dinb(n1614), .dout(n1617));
  jor  g01362(.dina(n1617), .dinb(n264), .dout(n1618));
  jor  g01363(.dina(n284), .dinb(n1400), .dout(n1619));
  jnot g01364(.din(b21 ), .dout(n1620));
  jor  g01365(.dina(n269), .dinb(n1620), .dout(n1621));
  jor  g01366(.dina(n271), .dinb(n1420), .dout(n1622));
  jand g01367(.dina(n1622), .dinb(n1621), .dout(n1623));
  jand g01368(.dina(n1623), .dinb(n1619), .dout(n1624));
  jand g01369(.dina(n1624), .dinb(n1618), .dout(n1625));
  jxor g01370(.dina(n1625), .dinb(n260), .dout(n1626));
  jxor g01371(.dina(n1626), .dinb(n1611), .dout(n1627));
  jxor g01372(.dina(n1627), .dinb(n1522), .dout(f21 ));
  jand g01373(.dina(n1626), .dinb(n1611), .dout(n1629));
  jand g01374(.dina(n1627), .dinb(n1522), .dout(n1630));
  jor  g01375(.dina(n1630), .dinb(n1629), .dout(n1631));
  jor  g01376(.dina(n1609), .dinb(n1601), .dout(n1632));
  jnot g01377(.din(n1632), .dout(n1633));
  jand g01378(.dina(n1610), .dinb(n1525), .dout(n1634));
  jor  g01379(.dina(n1634), .dinb(n1633), .dout(n1635));
  jand g01380(.dina(n1598), .dinb(n1538), .dout(n1636));
  jand g01381(.dina(n1599), .dinb(n1529), .dout(n1637));
  jor  g01382(.dina(n1637), .dinb(n1636), .dout(n1638));
  jor  g01383(.dina(n1019), .dinb(n528), .dout(n1639));
  jor  g01384(.dina(n490), .dinb(n858), .dout(n1640));
  jor  g01385(.dina(n531), .dinb(n939), .dout(n1641));
  jor  g01386(.dina(n533), .dinb(n1022), .dout(n1642));
  jand g01387(.dina(n1642), .dinb(n1641), .dout(n1643));
  jand g01388(.dina(n1643), .dinb(n1640), .dout(n1644));
  jand g01389(.dina(n1644), .dinb(n1639), .dout(n1645));
  jxor g01390(.dina(n1645), .dinb(a8 ), .dout(n1646));
  jnot g01391(.din(n1646), .dout(n1647));
  jand g01392(.dina(n1596), .dinb(n1550), .dout(n1648));
  jand g01393(.dina(n1597), .dinb(n1541), .dout(n1649));
  jor  g01394(.dina(n1649), .dinb(n1648), .dout(n1650));
  jand g01395(.dina(n1594), .dinb(n1562), .dout(n1651));
  jand g01396(.dina(n1595), .dinb(n1553), .dout(n1652));
  jor  g01397(.dina(n1652), .dinb(n1651), .dout(n1653));
  jor  g01398(.dina(n1592), .dinb(n1584), .dout(n1654));
  jand g01399(.dina(n1593), .dinb(n1565), .dout(n1655));
  jnot g01400(.din(n1655), .dout(n1656));
  jand g01401(.dina(n1656), .dinb(n1654), .dout(n1657));
  jnot g01402(.din(n1657), .dout(n1658));
  jor  g01403(.dina(n1245), .dinb(n428), .dout(n1659));
  jor  g01404(.dina(n1165), .dinb(n357), .dout(n1660));
  jor  g01405(.dina(n1248), .dinb(n395), .dout(n1661));
  jor  g01406(.dina(n1250), .dinb(n431), .dout(n1662));
  jand g01407(.dina(n1662), .dinb(n1661), .dout(n1663));
  jand g01408(.dina(n1663), .dinb(n1660), .dout(n1664));
  jand g01409(.dina(n1664), .dinb(n1659), .dout(n1665));
  jxor g01410(.dina(n1665), .dinb(a17 ), .dout(n1666));
  jnot g01411(.din(n1666), .dout(n1667));
  jnot g01412(.din(n1581), .dout(n1668));
  jand g01413(.dina(n1668), .dinb(n1579), .dout(n1669));
  jand g01414(.dina(n1582), .dinb(n1577), .dout(n1670));
  jor  g01415(.dina(n1670), .dinb(n1669), .dout(n1671));
  jor  g01416(.dina(n1566), .dinb(n319), .dout(n1672));
  jor  g01417(.dina(n1489), .dinb(n279), .dout(n1673));
  jor  g01418(.dina(n1569), .dinb(n299), .dout(n1674));
  jor  g01419(.dina(n1571), .dinb(n322), .dout(n1675));
  jand g01420(.dina(n1675), .dinb(n1674), .dout(n1676));
  jand g01421(.dina(n1676), .dinb(n1673), .dout(n1677));
  jand g01422(.dina(n1677), .dinb(n1672), .dout(n1678));
  jxor g01423(.dina(n1678), .dinb(a20 ), .dout(n1679));
  jnot g01424(.din(n1679), .dout(n1680));
  jand g01425(.dina(n1579), .dinb(a23 ), .dout(n1681));
  jxor g01426(.dina(a23 ), .dinb(a22 ), .dout(n1682));
  jnot g01427(.din(n1682), .dout(n1683));
  jand g01428(.dina(n1683), .dinb(n1578), .dout(n1684));
  jand g01429(.dina(n1684), .dinb(b1 ), .dout(n1685));
  jnot g01430(.din(n1578), .dout(n1686));
  jxor g01431(.dina(a22 ), .dinb(a21 ), .dout(n1687));
  jand g01432(.dina(n1687), .dinb(n1686), .dout(n1688));
  jand g01433(.dina(n1688), .dinb(b0 ), .dout(n1689));
  jand g01434(.dina(n1682), .dinb(n1578), .dout(n1690));
  jand g01435(.dina(n1690), .dinb(n338), .dout(n1691));
  jor  g01436(.dina(n1691), .dinb(n1689), .dout(n1692));
  jor  g01437(.dina(n1692), .dinb(n1685), .dout(n1693));
  jxor g01438(.dina(n1693), .dinb(n1681), .dout(n1694));
  jxor g01439(.dina(n1694), .dinb(n1680), .dout(n1695));
  jxor g01440(.dina(n1695), .dinb(n1671), .dout(n1696));
  jxor g01441(.dina(n1696), .dinb(n1667), .dout(n1697));
  jxor g01442(.dina(n1697), .dinb(n1658), .dout(n1698));
  jnot g01443(.din(n1698), .dout(n1699));
  jor  g01444(.dina(n974), .dinb(n624), .dout(n1700));
  jor  g01445(.dina(n908), .dinb(n512), .dout(n1701));
  jor  g01446(.dina(n977), .dinb(n564), .dout(n1702));
  jor  g01447(.dina(n979), .dinb(n627), .dout(n1703));
  jand g01448(.dina(n1703), .dinb(n1702), .dout(n1704));
  jand g01449(.dina(n1704), .dinb(n1701), .dout(n1705));
  jand g01450(.dina(n1705), .dinb(n1700), .dout(n1706));
  jxor g01451(.dina(n1706), .dinb(a14 ), .dout(n1707));
  jxor g01452(.dina(n1707), .dinb(n1699), .dout(n1708));
  jxor g01453(.dina(n1708), .dinb(n1653), .dout(n1709));
  jnot g01454(.din(n1709), .dout(n1710));
  jor  g01455(.dina(n775), .dinb(n706), .dout(n1711));
  jor  g01456(.dina(n683), .dinb(n647), .dout(n1712));
  jor  g01457(.dina(n709), .dinb(n758), .dout(n1713));
  jor  g01458(.dina(n711), .dinb(n778), .dout(n1714));
  jand g01459(.dina(n1714), .dinb(n1713), .dout(n1715));
  jand g01460(.dina(n1715), .dinb(n1712), .dout(n1716));
  jand g01461(.dina(n1716), .dinb(n1711), .dout(n1717));
  jxor g01462(.dina(n1717), .dinb(a11 ), .dout(n1718));
  jxor g01463(.dina(n1718), .dinb(n1710), .dout(n1719));
  jxor g01464(.dina(n1719), .dinb(n1650), .dout(n1720));
  jxor g01465(.dina(n1720), .dinb(n1647), .dout(n1721));
  jnot g01466(.din(n1721), .dout(n1722));
  jxor g01467(.dina(n1722), .dinb(n1638), .dout(n1723));
  jor  g01468(.dina(n1397), .dinb(n402), .dout(n1724));
  jor  g01469(.dina(n371), .dinb(n1193), .dout(n1725));
  jor  g01470(.dina(n405), .dinb(n1290), .dout(n1726));
  jor  g01471(.dina(n332), .dinb(n1400), .dout(n1727));
  jand g01472(.dina(n1727), .dinb(n1726), .dout(n1728));
  jand g01473(.dina(n1728), .dinb(n1725), .dout(n1729));
  jand g01474(.dina(n1729), .dinb(n1724), .dout(n1730));
  jxor g01475(.dina(n1730), .dinb(a5 ), .dout(n1731));
  jxor g01476(.dina(n1731), .dinb(n1723), .dout(n1732));
  jxor g01477(.dina(n1732), .dinb(n1635), .dout(n1733));
  jand g01478(.dina(b21 ), .dinb(b20 ), .dout(n1734));
  jand g01479(.dina(n1615), .dinb(n1614), .dout(n1735));
  jor  g01480(.dina(n1735), .dinb(n1734), .dout(n1736));
  jxor g01481(.dina(b22 ), .dinb(b21 ), .dout(n1737));
  jnot g01482(.din(n1737), .dout(n1738));
  jxor g01483(.dina(n1738), .dinb(n1736), .dout(n1739));
  jor  g01484(.dina(n1739), .dinb(n264), .dout(n1740));
  jor  g01485(.dina(n284), .dinb(n1420), .dout(n1741));
  jnot g01486(.din(b22 ), .dout(n1742));
  jor  g01487(.dina(n269), .dinb(n1742), .dout(n1743));
  jor  g01488(.dina(n271), .dinb(n1620), .dout(n1744));
  jand g01489(.dina(n1744), .dinb(n1743), .dout(n1745));
  jand g01490(.dina(n1745), .dinb(n1741), .dout(n1746));
  jand g01491(.dina(n1746), .dinb(n1740), .dout(n1747));
  jxor g01492(.dina(n1747), .dinb(n260), .dout(n1748));
  jxor g01493(.dina(n1748), .dinb(n1733), .dout(n1749));
  jxor g01494(.dina(n1749), .dinb(n1631), .dout(f22 ));
  jand g01495(.dina(n1748), .dinb(n1733), .dout(n1751));
  jand g01496(.dina(n1749), .dinb(n1631), .dout(n1752));
  jor  g01497(.dina(n1752), .dinb(n1751), .dout(n1753));
  jor  g01498(.dina(n1731), .dinb(n1723), .dout(n1754));
  jnot g01499(.din(n1754), .dout(n1755));
  jand g01500(.dina(n1732), .dinb(n1635), .dout(n1756));
  jor  g01501(.dina(n1756), .dinb(n1755), .dout(n1757));
  jor  g01502(.dina(n1417), .dinb(n402), .dout(n1758));
  jor  g01503(.dina(n371), .dinb(n1290), .dout(n1759));
  jor  g01504(.dina(n405), .dinb(n1400), .dout(n1760));
  jor  g01505(.dina(n332), .dinb(n1420), .dout(n1761));
  jand g01506(.dina(n1761), .dinb(n1760), .dout(n1762));
  jand g01507(.dina(n1762), .dinb(n1759), .dout(n1763));
  jand g01508(.dina(n1763), .dinb(n1758), .dout(n1764));
  jxor g01509(.dina(n1764), .dinb(a5 ), .dout(n1765));
  jnot g01510(.din(n1765), .dout(n1766));
  jand g01511(.dina(n1720), .dinb(n1647), .dout(n1767));
  jand g01512(.dina(n1721), .dinb(n1638), .dout(n1768));
  jor  g01513(.dina(n1768), .dinb(n1767), .dout(n1769));
  jor  g01514(.dina(n1190), .dinb(n528), .dout(n1770));
  jor  g01515(.dina(n490), .dinb(n939), .dout(n1771));
  jor  g01516(.dina(n531), .dinb(n1022), .dout(n1772));
  jor  g01517(.dina(n533), .dinb(n1193), .dout(n1773));
  jand g01518(.dina(n1773), .dinb(n1772), .dout(n1774));
  jand g01519(.dina(n1774), .dinb(n1771), .dout(n1775));
  jand g01520(.dina(n1775), .dinb(n1770), .dout(n1776));
  jxor g01521(.dina(n1776), .dinb(a8 ), .dout(n1777));
  jnot g01522(.din(n1777), .dout(n1778));
  jor  g01523(.dina(n1718), .dinb(n1710), .dout(n1779));
  jand g01524(.dina(n1719), .dinb(n1650), .dout(n1780));
  jnot g01525(.din(n1780), .dout(n1781));
  jand g01526(.dina(n1781), .dinb(n1779), .dout(n1782));
  jor  g01527(.dina(n1707), .dinb(n1699), .dout(n1783));
  jand g01528(.dina(n1708), .dinb(n1653), .dout(n1784));
  jnot g01529(.din(n1784), .dout(n1785));
  jand g01530(.dina(n1785), .dinb(n1783), .dout(n1786));
  jnot g01531(.din(n1786), .dout(n1787));
  jor  g01532(.dina(n974), .dinb(n644), .dout(n1788));
  jor  g01533(.dina(n908), .dinb(n564), .dout(n1789));
  jor  g01534(.dina(n977), .dinb(n627), .dout(n1790));
  jor  g01535(.dina(n979), .dinb(n647), .dout(n1791));
  jand g01536(.dina(n1791), .dinb(n1790), .dout(n1792));
  jand g01537(.dina(n1792), .dinb(n1789), .dout(n1793));
  jand g01538(.dina(n1793), .dinb(n1788), .dout(n1794));
  jxor g01539(.dina(n1794), .dinb(a14 ), .dout(n1795));
  jnot g01540(.din(n1795), .dout(n1796));
  jand g01541(.dina(n1696), .dinb(n1667), .dout(n1797));
  jand g01542(.dina(n1697), .dinb(n1658), .dout(n1798));
  jor  g01543(.dina(n1798), .dinb(n1797), .dout(n1799));
  jor  g01544(.dina(n1245), .dinb(n509), .dout(n1800));
  jor  g01545(.dina(n1165), .dinb(n395), .dout(n1801));
  jor  g01546(.dina(n1248), .dinb(n431), .dout(n1802));
  jor  g01547(.dina(n1250), .dinb(n512), .dout(n1803));
  jand g01548(.dina(n1803), .dinb(n1802), .dout(n1804));
  jand g01549(.dina(n1804), .dinb(n1801), .dout(n1805));
  jand g01550(.dina(n1805), .dinb(n1800), .dout(n1806));
  jxor g01551(.dina(n1806), .dinb(a17 ), .dout(n1807));
  jnot g01552(.din(n1807), .dout(n1808));
  jand g01553(.dina(n1694), .dinb(n1680), .dout(n1809));
  jand g01554(.dina(n1695), .dinb(n1671), .dout(n1810));
  jor  g01555(.dina(n1810), .dinb(n1809), .dout(n1811));
  jor  g01556(.dina(n1566), .dinb(n354), .dout(n1812));
  jor  g01557(.dina(n1489), .dinb(n299), .dout(n1813));
  jor  g01558(.dina(n1569), .dinb(n322), .dout(n1814));
  jor  g01559(.dina(n1571), .dinb(n357), .dout(n1815));
  jand g01560(.dina(n1815), .dinb(n1814), .dout(n1816));
  jand g01561(.dina(n1816), .dinb(n1813), .dout(n1817));
  jand g01562(.dina(n1817), .dinb(n1812), .dout(n1818));
  jxor g01563(.dina(n1818), .dinb(a20 ), .dout(n1819));
  jnot g01564(.din(n1819), .dout(n1820));
  jnot g01565(.din(n1693), .dout(n1821));
  jand g01566(.dina(n1580), .dinb(a23 ), .dout(n1822));
  jand g01567(.dina(n1822), .dinb(n1821), .dout(n1823));
  jnot g01568(.din(n1823), .dout(n1824));
  jand g01569(.dina(n1824), .dinb(a23 ), .dout(n1825));
  jor  g01570(.dina(n1687), .dinb(n1683), .dout(n1826));
  jor  g01571(.dina(n1826), .dinb(n1578), .dout(n1827));
  jnot g01572(.din(n1827), .dout(n1828));
  jand g01573(.dina(n1828), .dinb(b0 ), .dout(n1829));
  jand g01574(.dina(n1684), .dinb(b2 ), .dout(n1830));
  jand g01575(.dina(n1688), .dinb(b1 ), .dout(n1831));
  jand g01576(.dina(n1690), .dinb(n375), .dout(n1832));
  jor  g01577(.dina(n1832), .dinb(n1831), .dout(n1833));
  jor  g01578(.dina(n1833), .dinb(n1830), .dout(n1834));
  jor  g01579(.dina(n1834), .dinb(n1829), .dout(n1835));
  jxor g01580(.dina(n1835), .dinb(n1825), .dout(n1836));
  jxor g01581(.dina(n1836), .dinb(n1820), .dout(n1837));
  jxor g01582(.dina(n1837), .dinb(n1811), .dout(n1838));
  jxor g01583(.dina(n1838), .dinb(n1808), .dout(n1839));
  jxor g01584(.dina(n1839), .dinb(n1799), .dout(n1840));
  jxor g01585(.dina(n1840), .dinb(n1796), .dout(n1841));
  jxor g01586(.dina(n1841), .dinb(n1787), .dout(n1842));
  jnot g01587(.din(n1842), .dout(n1843));
  jor  g01588(.dina(n855), .dinb(n706), .dout(n1844));
  jor  g01589(.dina(n683), .dinb(n758), .dout(n1845));
  jor  g01590(.dina(n709), .dinb(n778), .dout(n1846));
  jor  g01591(.dina(n711), .dinb(n858), .dout(n1847));
  jand g01592(.dina(n1847), .dinb(n1846), .dout(n1848));
  jand g01593(.dina(n1848), .dinb(n1845), .dout(n1849));
  jand g01594(.dina(n1849), .dinb(n1844), .dout(n1850));
  jxor g01595(.dina(n1850), .dinb(a11 ), .dout(n1851));
  jxor g01596(.dina(n1851), .dinb(n1843), .dout(n1852));
  jnot g01597(.din(n1852), .dout(n1853));
  jxor g01598(.dina(n1853), .dinb(n1782), .dout(n1854));
  jxor g01599(.dina(n1854), .dinb(n1778), .dout(n1855));
  jxor g01600(.dina(n1855), .dinb(n1769), .dout(n1856));
  jxor g01601(.dina(n1856), .dinb(n1766), .dout(n1857));
  jxor g01602(.dina(n1857), .dinb(n1757), .dout(n1858));
  jand g01603(.dina(b22 ), .dinb(b21 ), .dout(n1859));
  jand g01604(.dina(n1737), .dinb(n1736), .dout(n1860));
  jor  g01605(.dina(n1860), .dinb(n1859), .dout(n1861));
  jxor g01606(.dina(b23 ), .dinb(b22 ), .dout(n1862));
  jnot g01607(.din(n1862), .dout(n1863));
  jxor g01608(.dina(n1863), .dinb(n1861), .dout(n1864));
  jor  g01609(.dina(n1864), .dinb(n264), .dout(n1865));
  jor  g01610(.dina(n284), .dinb(n1620), .dout(n1866));
  jnot g01611(.din(b23 ), .dout(n1867));
  jor  g01612(.dina(n269), .dinb(n1867), .dout(n1868));
  jor  g01613(.dina(n271), .dinb(n1742), .dout(n1869));
  jand g01614(.dina(n1869), .dinb(n1868), .dout(n1870));
  jand g01615(.dina(n1870), .dinb(n1866), .dout(n1871));
  jand g01616(.dina(n1871), .dinb(n1865), .dout(n1872));
  jxor g01617(.dina(n1872), .dinb(n260), .dout(n1873));
  jxor g01618(.dina(n1873), .dinb(n1858), .dout(n1874));
  jxor g01619(.dina(n1874), .dinb(n1753), .dout(f23 ));
  jand g01620(.dina(n1873), .dinb(n1858), .dout(n1876));
  jand g01621(.dina(n1874), .dinb(n1753), .dout(n1877));
  jor  g01622(.dina(n1877), .dinb(n1876), .dout(n1878));
  jand g01623(.dina(b23 ), .dinb(b22 ), .dout(n1879));
  jand g01624(.dina(n1862), .dinb(n1861), .dout(n1880));
  jor  g01625(.dina(n1880), .dinb(n1879), .dout(n1881));
  jxor g01626(.dina(b24 ), .dinb(b23 ), .dout(n1882));
  jnot g01627(.din(n1882), .dout(n1883));
  jxor g01628(.dina(n1883), .dinb(n1881), .dout(n1884));
  jor  g01629(.dina(n1884), .dinb(n264), .dout(n1885));
  jor  g01630(.dina(n284), .dinb(n1742), .dout(n1886));
  jnot g01631(.din(b24 ), .dout(n1887));
  jor  g01632(.dina(n269), .dinb(n1887), .dout(n1888));
  jor  g01633(.dina(n271), .dinb(n1867), .dout(n1889));
  jand g01634(.dina(n1889), .dinb(n1888), .dout(n1890));
  jand g01635(.dina(n1890), .dinb(n1886), .dout(n1891));
  jand g01636(.dina(n1891), .dinb(n1885), .dout(n1892));
  jxor g01637(.dina(n1892), .dinb(n260), .dout(n1893));
  jand g01638(.dina(n1856), .dinb(n1766), .dout(n1894));
  jand g01639(.dina(n1857), .dinb(n1757), .dout(n1895));
  jor  g01640(.dina(n1895), .dinb(n1894), .dout(n1896));
  jor  g01641(.dina(n1617), .dinb(n402), .dout(n1897));
  jor  g01642(.dina(n371), .dinb(n1400), .dout(n1898));
  jor  g01643(.dina(n405), .dinb(n1420), .dout(n1899));
  jor  g01644(.dina(n332), .dinb(n1620), .dout(n1900));
  jand g01645(.dina(n1900), .dinb(n1899), .dout(n1901));
  jand g01646(.dina(n1901), .dinb(n1898), .dout(n1902));
  jand g01647(.dina(n1902), .dinb(n1897), .dout(n1903));
  jxor g01648(.dina(n1903), .dinb(a5 ), .dout(n1904));
  jnot g01649(.din(n1904), .dout(n1905));
  jand g01650(.dina(n1854), .dinb(n1778), .dout(n1906));
  jand g01651(.dina(n1855), .dinb(n1769), .dout(n1907));
  jor  g01652(.dina(n1907), .dinb(n1906), .dout(n1908));
  jor  g01653(.dina(n1851), .dinb(n1843), .dout(n1909));
  jor  g01654(.dina(n1853), .dinb(n1782), .dout(n1910));
  jand g01655(.dina(n1910), .dinb(n1909), .dout(n1911));
  jand g01656(.dina(n1840), .dinb(n1796), .dout(n1912));
  jand g01657(.dina(n1841), .dinb(n1787), .dout(n1913));
  jor  g01658(.dina(n1913), .dinb(n1912), .dout(n1914));
  jor  g01659(.dina(n974), .dinb(n755), .dout(n1915));
  jor  g01660(.dina(n908), .dinb(n627), .dout(n1916));
  jor  g01661(.dina(n977), .dinb(n647), .dout(n1917));
  jor  g01662(.dina(n979), .dinb(n758), .dout(n1918));
  jand g01663(.dina(n1918), .dinb(n1917), .dout(n1919));
  jand g01664(.dina(n1919), .dinb(n1916), .dout(n1920));
  jand g01665(.dina(n1920), .dinb(n1915), .dout(n1921));
  jxor g01666(.dina(n1921), .dinb(a14 ), .dout(n1922));
  jnot g01667(.din(n1922), .dout(n1923));
  jand g01668(.dina(n1838), .dinb(n1808), .dout(n1924));
  jand g01669(.dina(n1839), .dinb(n1799), .dout(n1925));
  jor  g01670(.dina(n1925), .dinb(n1924), .dout(n1926));
  jor  g01671(.dina(n1245), .dinb(n561), .dout(n1927));
  jor  g01672(.dina(n1165), .dinb(n431), .dout(n1928));
  jor  g01673(.dina(n1248), .dinb(n512), .dout(n1929));
  jor  g01674(.dina(n1250), .dinb(n564), .dout(n1930));
  jand g01675(.dina(n1930), .dinb(n1929), .dout(n1931));
  jand g01676(.dina(n1931), .dinb(n1928), .dout(n1932));
  jand g01677(.dina(n1932), .dinb(n1927), .dout(n1933));
  jxor g01678(.dina(n1933), .dinb(a17 ), .dout(n1934));
  jnot g01679(.din(n1934), .dout(n1935));
  jand g01680(.dina(n1836), .dinb(n1820), .dout(n1936));
  jand g01681(.dina(n1837), .dinb(n1811), .dout(n1937));
  jor  g01682(.dina(n1937), .dinb(n1936), .dout(n1938));
  jnot g01683(.din(n1690), .dout(n1939));
  jor  g01684(.dina(n1939), .dinb(n296), .dout(n1940));
  jor  g01685(.dina(n1827), .dinb(n267), .dout(n1941));
  jnot g01686(.din(n1688), .dout(n1942));
  jor  g01687(.dina(n1942), .dinb(n279), .dout(n1943));
  jnot g01688(.din(n1684), .dout(n1944));
  jor  g01689(.dina(n1944), .dinb(n299), .dout(n1945));
  jand g01690(.dina(n1945), .dinb(n1943), .dout(n1946));
  jand g01691(.dina(n1946), .dinb(n1941), .dout(n1947));
  jand g01692(.dina(n1947), .dinb(n1940), .dout(n1948));
  jxor g01693(.dina(n1948), .dinb(a23 ), .dout(n1949));
  jnot g01694(.din(n1949), .dout(n1950));
  jxor g01695(.dina(a24 ), .dinb(a23 ), .dout(n1951));
  jand g01696(.dina(n1951), .dinb(b0 ), .dout(n1952));
  jnot g01697(.din(n1952), .dout(n1953));
  jor  g01698(.dina(n1835), .dinb(n1824), .dout(n1954));
  jxor g01699(.dina(n1954), .dinb(n1953), .dout(n1955));
  jxor g01700(.dina(n1955), .dinb(n1950), .dout(n1956));
  jnot g01701(.din(n1956), .dout(n1957));
  jor  g01702(.dina(n1566), .dinb(n392), .dout(n1958));
  jor  g01703(.dina(n1489), .dinb(n322), .dout(n1959));
  jor  g01704(.dina(n1569), .dinb(n357), .dout(n1960));
  jor  g01705(.dina(n1571), .dinb(n395), .dout(n1961));
  jand g01706(.dina(n1961), .dinb(n1960), .dout(n1962));
  jand g01707(.dina(n1962), .dinb(n1959), .dout(n1963));
  jand g01708(.dina(n1963), .dinb(n1958), .dout(n1964));
  jxor g01709(.dina(n1964), .dinb(a20 ), .dout(n1965));
  jxor g01710(.dina(n1965), .dinb(n1957), .dout(n1966));
  jxor g01711(.dina(n1966), .dinb(n1938), .dout(n1967));
  jxor g01712(.dina(n1967), .dinb(n1935), .dout(n1968));
  jxor g01713(.dina(n1968), .dinb(n1926), .dout(n1969));
  jxor g01714(.dina(n1969), .dinb(n1923), .dout(n1970));
  jxor g01715(.dina(n1970), .dinb(n1914), .dout(n1971));
  jnot g01716(.din(n1971), .dout(n1972));
  jor  g01717(.dina(n936), .dinb(n706), .dout(n1973));
  jor  g01718(.dina(n683), .dinb(n778), .dout(n1974));
  jor  g01719(.dina(n709), .dinb(n858), .dout(n1975));
  jor  g01720(.dina(n711), .dinb(n939), .dout(n1976));
  jand g01721(.dina(n1976), .dinb(n1975), .dout(n1977));
  jand g01722(.dina(n1977), .dinb(n1974), .dout(n1978));
  jand g01723(.dina(n1978), .dinb(n1973), .dout(n1979));
  jxor g01724(.dina(n1979), .dinb(a11 ), .dout(n1980));
  jxor g01725(.dina(n1980), .dinb(n1972), .dout(n1981));
  jnot g01726(.din(n1981), .dout(n1982));
  jxor g01727(.dina(n1982), .dinb(n1911), .dout(n1983));
  jor  g01728(.dina(n1287), .dinb(n528), .dout(n1984));
  jor  g01729(.dina(n490), .dinb(n1022), .dout(n1985));
  jor  g01730(.dina(n531), .dinb(n1193), .dout(n1986));
  jor  g01731(.dina(n533), .dinb(n1290), .dout(n1987));
  jand g01732(.dina(n1987), .dinb(n1986), .dout(n1988));
  jand g01733(.dina(n1988), .dinb(n1985), .dout(n1989));
  jand g01734(.dina(n1989), .dinb(n1984), .dout(n1990));
  jxor g01735(.dina(n1990), .dinb(a8 ), .dout(n1991));
  jxor g01736(.dina(n1991), .dinb(n1983), .dout(n1992));
  jnot g01737(.din(n1992), .dout(n1993));
  jxor g01738(.dina(n1993), .dinb(n1908), .dout(n1994));
  jxor g01739(.dina(n1994), .dinb(n1905), .dout(n1995));
  jxor g01740(.dina(n1995), .dinb(n1896), .dout(n1996));
  jxor g01741(.dina(n1996), .dinb(n1893), .dout(n1997));
  jxor g01742(.dina(n1997), .dinb(n1878), .dout(f24 ));
  jand g01743(.dina(n1996), .dinb(n1893), .dout(n1999));
  jand g01744(.dina(n1997), .dinb(n1878), .dout(n2000));
  jor  g01745(.dina(n2000), .dinb(n1999), .dout(n2001));
  jand g01746(.dina(b24 ), .dinb(b23 ), .dout(n2002));
  jand g01747(.dina(n1882), .dinb(n1881), .dout(n2003));
  jor  g01748(.dina(n2003), .dinb(n2002), .dout(n2004));
  jxor g01749(.dina(b25 ), .dinb(b24 ), .dout(n2005));
  jnot g01750(.din(n2005), .dout(n2006));
  jxor g01751(.dina(n2006), .dinb(n2004), .dout(n2007));
  jor  g01752(.dina(n2007), .dinb(n264), .dout(n2008));
  jor  g01753(.dina(n284), .dinb(n1867), .dout(n2009));
  jnot g01754(.din(b25 ), .dout(n2010));
  jor  g01755(.dina(n269), .dinb(n2010), .dout(n2011));
  jor  g01756(.dina(n271), .dinb(n1887), .dout(n2012));
  jand g01757(.dina(n2012), .dinb(n2011), .dout(n2013));
  jand g01758(.dina(n2013), .dinb(n2009), .dout(n2014));
  jand g01759(.dina(n2014), .dinb(n2008), .dout(n2015));
  jxor g01760(.dina(n2015), .dinb(n260), .dout(n2016));
  jand g01761(.dina(n1994), .dinb(n1905), .dout(n2017));
  jand g01762(.dina(n1995), .dinb(n1896), .dout(n2018));
  jor  g01763(.dina(n2018), .dinb(n2017), .dout(n2019));
  jor  g01764(.dina(n1739), .dinb(n402), .dout(n2020));
  jor  g01765(.dina(n371), .dinb(n1420), .dout(n2021));
  jor  g01766(.dina(n405), .dinb(n1620), .dout(n2022));
  jor  g01767(.dina(n332), .dinb(n1742), .dout(n2023));
  jand g01768(.dina(n2023), .dinb(n2022), .dout(n2024));
  jand g01769(.dina(n2024), .dinb(n2021), .dout(n2025));
  jand g01770(.dina(n2025), .dinb(n2020), .dout(n2026));
  jxor g01771(.dina(n2026), .dinb(a5 ), .dout(n2027));
  jnot g01772(.din(n2027), .dout(n2028));
  jnot g01773(.din(n1983), .dout(n2029));
  jor  g01774(.dina(n1991), .dinb(n2029), .dout(n2030));
  jnot g01775(.din(n2030), .dout(n2031));
  jand g01776(.dina(n1993), .dinb(n1908), .dout(n2032));
  jor  g01777(.dina(n2032), .dinb(n2031), .dout(n2033));
  jor  g01778(.dina(n1980), .dinb(n1972), .dout(n2034));
  jor  g01779(.dina(n1982), .dinb(n1911), .dout(n2035));
  jand g01780(.dina(n2035), .dinb(n2034), .dout(n2036));
  jand g01781(.dina(n1967), .dinb(n1935), .dout(n2037));
  jand g01782(.dina(n1968), .dinb(n1926), .dout(n2038));
  jor  g01783(.dina(n2038), .dinb(n2037), .dout(n2039));
  jor  g01784(.dina(n1965), .dinb(n1957), .dout(n2040));
  jand g01785(.dina(n1966), .dinb(n1938), .dout(n2041));
  jnot g01786(.din(n2041), .dout(n2042));
  jand g01787(.dina(n2042), .dinb(n2040), .dout(n2043));
  jnot g01788(.din(n2043), .dout(n2044));
  jor  g01789(.dina(n1566), .dinb(n428), .dout(n2045));
  jor  g01790(.dina(n1489), .dinb(n357), .dout(n2046));
  jor  g01791(.dina(n1569), .dinb(n395), .dout(n2047));
  jor  g01792(.dina(n1571), .dinb(n431), .dout(n2048));
  jand g01793(.dina(n2048), .dinb(n2047), .dout(n2049));
  jand g01794(.dina(n2049), .dinb(n2046), .dout(n2050));
  jand g01795(.dina(n2050), .dinb(n2045), .dout(n2051));
  jxor g01796(.dina(n2051), .dinb(a20 ), .dout(n2052));
  jnot g01797(.din(n2052), .dout(n2053));
  jnot g01798(.din(n1954), .dout(n2054));
  jand g01799(.dina(n2054), .dinb(n1952), .dout(n2055));
  jand g01800(.dina(n1955), .dinb(n1950), .dout(n2056));
  jor  g01801(.dina(n2056), .dinb(n2055), .dout(n2057));
  jor  g01802(.dina(n1939), .dinb(n319), .dout(n2058));
  jor  g01803(.dina(n1827), .dinb(n279), .dout(n2059));
  jor  g01804(.dina(n1942), .dinb(n299), .dout(n2060));
  jor  g01805(.dina(n1944), .dinb(n322), .dout(n2061));
  jand g01806(.dina(n2061), .dinb(n2060), .dout(n2062));
  jand g01807(.dina(n2062), .dinb(n2059), .dout(n2063));
  jand g01808(.dina(n2063), .dinb(n2058), .dout(n2064));
  jxor g01809(.dina(n2064), .dinb(a23 ), .dout(n2065));
  jnot g01810(.din(n2065), .dout(n2066));
  jand g01811(.dina(n1952), .dinb(a26 ), .dout(n2067));
  jxor g01812(.dina(a26 ), .dinb(a25 ), .dout(n2068));
  jnot g01813(.din(n2068), .dout(n2069));
  jand g01814(.dina(n2069), .dinb(n1951), .dout(n2070));
  jand g01815(.dina(n2070), .dinb(b1 ), .dout(n2071));
  jnot g01816(.din(n1951), .dout(n2072));
  jxor g01817(.dina(a25 ), .dinb(a24 ), .dout(n2073));
  jand g01818(.dina(n2073), .dinb(n2072), .dout(n2074));
  jand g01819(.dina(n2074), .dinb(b0 ), .dout(n2075));
  jand g01820(.dina(n2068), .dinb(n1951), .dout(n2076));
  jand g01821(.dina(n2076), .dinb(n338), .dout(n2077));
  jor  g01822(.dina(n2077), .dinb(n2075), .dout(n2078));
  jor  g01823(.dina(n2078), .dinb(n2071), .dout(n2079));
  jxor g01824(.dina(n2079), .dinb(n2067), .dout(n2080));
  jxor g01825(.dina(n2080), .dinb(n2066), .dout(n2081));
  jxor g01826(.dina(n2081), .dinb(n2057), .dout(n2082));
  jxor g01827(.dina(n2082), .dinb(n2053), .dout(n2083));
  jxor g01828(.dina(n2083), .dinb(n2044), .dout(n2084));
  jnot g01829(.din(n2084), .dout(n2085));
  jor  g01830(.dina(n1245), .dinb(n624), .dout(n2086));
  jor  g01831(.dina(n1165), .dinb(n512), .dout(n2087));
  jor  g01832(.dina(n1248), .dinb(n564), .dout(n2088));
  jor  g01833(.dina(n1250), .dinb(n627), .dout(n2089));
  jand g01834(.dina(n2089), .dinb(n2088), .dout(n2090));
  jand g01835(.dina(n2090), .dinb(n2087), .dout(n2091));
  jand g01836(.dina(n2091), .dinb(n2086), .dout(n2092));
  jxor g01837(.dina(n2092), .dinb(a17 ), .dout(n2093));
  jxor g01838(.dina(n2093), .dinb(n2085), .dout(n2094));
  jxor g01839(.dina(n2094), .dinb(n2039), .dout(n2095));
  jnot g01840(.din(n2095), .dout(n2096));
  jor  g01841(.dina(n974), .dinb(n775), .dout(n2097));
  jor  g01842(.dina(n908), .dinb(n647), .dout(n2098));
  jor  g01843(.dina(n977), .dinb(n758), .dout(n2099));
  jor  g01844(.dina(n979), .dinb(n778), .dout(n2100));
  jand g01845(.dina(n2100), .dinb(n2099), .dout(n2101));
  jand g01846(.dina(n2101), .dinb(n2098), .dout(n2102));
  jand g01847(.dina(n2102), .dinb(n2097), .dout(n2103));
  jxor g01848(.dina(n2103), .dinb(a14 ), .dout(n2104));
  jxor g01849(.dina(n2104), .dinb(n2096), .dout(n2105));
  jand g01850(.dina(n1969), .dinb(n1923), .dout(n2106));
  jand g01851(.dina(n1970), .dinb(n1914), .dout(n2107));
  jor  g01852(.dina(n2107), .dinb(n2106), .dout(n2108));
  jxor g01853(.dina(n2108), .dinb(n2105), .dout(n2109));
  jnot g01854(.din(n2109), .dout(n2110));
  jor  g01855(.dina(n1019), .dinb(n706), .dout(n2111));
  jor  g01856(.dina(n683), .dinb(n858), .dout(n2112));
  jor  g01857(.dina(n709), .dinb(n939), .dout(n2113));
  jor  g01858(.dina(n711), .dinb(n1022), .dout(n2114));
  jand g01859(.dina(n2114), .dinb(n2113), .dout(n2115));
  jand g01860(.dina(n2115), .dinb(n2112), .dout(n2116));
  jand g01861(.dina(n2116), .dinb(n2111), .dout(n2117));
  jxor g01862(.dina(n2117), .dinb(a11 ), .dout(n2118));
  jxor g01863(.dina(n2118), .dinb(n2110), .dout(n2119));
  jnot g01864(.din(n2119), .dout(n2120));
  jxor g01865(.dina(n2120), .dinb(n2036), .dout(n2121));
  jor  g01866(.dina(n1397), .dinb(n528), .dout(n2122));
  jor  g01867(.dina(n490), .dinb(n1193), .dout(n2123));
  jor  g01868(.dina(n531), .dinb(n1290), .dout(n2124));
  jor  g01869(.dina(n533), .dinb(n1400), .dout(n2125));
  jand g01870(.dina(n2125), .dinb(n2124), .dout(n2126));
  jand g01871(.dina(n2126), .dinb(n2123), .dout(n2127));
  jand g01872(.dina(n2127), .dinb(n2122), .dout(n2128));
  jxor g01873(.dina(n2128), .dinb(a8 ), .dout(n2129));
  jxor g01874(.dina(n2129), .dinb(n2121), .dout(n2130));
  jnot g01875(.din(n2130), .dout(n2131));
  jxor g01876(.dina(n2131), .dinb(n2033), .dout(n2132));
  jxor g01877(.dina(n2132), .dinb(n2028), .dout(n2133));
  jxor g01878(.dina(n2133), .dinb(n2019), .dout(n2134));
  jxor g01879(.dina(n2134), .dinb(n2016), .dout(n2135));
  jxor g01880(.dina(n2135), .dinb(n2001), .dout(f25 ));
  jand g01881(.dina(n2134), .dinb(n2016), .dout(n2137));
  jand g01882(.dina(n2135), .dinb(n2001), .dout(n2138));
  jor  g01883(.dina(n2138), .dinb(n2137), .dout(n2139));
  jand g01884(.dina(b25 ), .dinb(b24 ), .dout(n2140));
  jand g01885(.dina(n2005), .dinb(n2004), .dout(n2141));
  jor  g01886(.dina(n2141), .dinb(n2140), .dout(n2142));
  jxor g01887(.dina(b26 ), .dinb(b25 ), .dout(n2143));
  jnot g01888(.din(n2143), .dout(n2144));
  jxor g01889(.dina(n2144), .dinb(n2142), .dout(n2145));
  jor  g01890(.dina(n2145), .dinb(n264), .dout(n2146));
  jor  g01891(.dina(n284), .dinb(n1887), .dout(n2147));
  jnot g01892(.din(b26 ), .dout(n2148));
  jor  g01893(.dina(n269), .dinb(n2148), .dout(n2149));
  jor  g01894(.dina(n271), .dinb(n2010), .dout(n2150));
  jand g01895(.dina(n2150), .dinb(n2149), .dout(n2151));
  jand g01896(.dina(n2151), .dinb(n2147), .dout(n2152));
  jand g01897(.dina(n2152), .dinb(n2146), .dout(n2153));
  jxor g01898(.dina(n2153), .dinb(n260), .dout(n2154));
  jand g01899(.dina(n2132), .dinb(n2028), .dout(n2155));
  jand g01900(.dina(n2133), .dinb(n2019), .dout(n2156));
  jor  g01901(.dina(n2156), .dinb(n2155), .dout(n2157));
  jnot g01902(.din(n2121), .dout(n2158));
  jor  g01903(.dina(n2129), .dinb(n2158), .dout(n2159));
  jnot g01904(.din(n2159), .dout(n2160));
  jand g01905(.dina(n2131), .dinb(n2033), .dout(n2161));
  jor  g01906(.dina(n2161), .dinb(n2160), .dout(n2162));
  jor  g01907(.dina(n2118), .dinb(n2110), .dout(n2163));
  jor  g01908(.dina(n2120), .dinb(n2036), .dout(n2164));
  jand g01909(.dina(n2164), .dinb(n2163), .dout(n2165));
  jor  g01910(.dina(n1190), .dinb(n706), .dout(n2166));
  jor  g01911(.dina(n683), .dinb(n939), .dout(n2167));
  jor  g01912(.dina(n709), .dinb(n1022), .dout(n2168));
  jor  g01913(.dina(n711), .dinb(n1193), .dout(n2169));
  jand g01914(.dina(n2169), .dinb(n2168), .dout(n2170));
  jand g01915(.dina(n2170), .dinb(n2167), .dout(n2171));
  jand g01916(.dina(n2171), .dinb(n2166), .dout(n2172));
  jxor g01917(.dina(n2172), .dinb(a11 ), .dout(n2173));
  jnot g01918(.din(n2173), .dout(n2174));
  jor  g01919(.dina(n2104), .dinb(n2096), .dout(n2175));
  jand g01920(.dina(n2108), .dinb(n2105), .dout(n2176));
  jnot g01921(.din(n2176), .dout(n2177));
  jand g01922(.dina(n2177), .dinb(n2175), .dout(n2178));
  jnot g01923(.din(n2178), .dout(n2179));
  jor  g01924(.dina(n2093), .dinb(n2085), .dout(n2180));
  jand g01925(.dina(n2094), .dinb(n2039), .dout(n2181));
  jnot g01926(.din(n2181), .dout(n2182));
  jand g01927(.dina(n2182), .dinb(n2180), .dout(n2183));
  jnot g01928(.din(n2183), .dout(n2184));
  jor  g01929(.dina(n1245), .dinb(n644), .dout(n2185));
  jor  g01930(.dina(n1165), .dinb(n564), .dout(n2186));
  jor  g01931(.dina(n1248), .dinb(n627), .dout(n2187));
  jor  g01932(.dina(n1250), .dinb(n647), .dout(n2188));
  jand g01933(.dina(n2188), .dinb(n2187), .dout(n2189));
  jand g01934(.dina(n2189), .dinb(n2186), .dout(n2190));
  jand g01935(.dina(n2190), .dinb(n2185), .dout(n2191));
  jxor g01936(.dina(n2191), .dinb(a17 ), .dout(n2192));
  jnot g01937(.din(n2192), .dout(n2193));
  jand g01938(.dina(n2082), .dinb(n2053), .dout(n2194));
  jand g01939(.dina(n2083), .dinb(n2044), .dout(n2195));
  jor  g01940(.dina(n2195), .dinb(n2194), .dout(n2196));
  jor  g01941(.dina(n1566), .dinb(n509), .dout(n2197));
  jor  g01942(.dina(n1489), .dinb(n395), .dout(n2198));
  jor  g01943(.dina(n1569), .dinb(n431), .dout(n2199));
  jor  g01944(.dina(n1571), .dinb(n512), .dout(n2200));
  jand g01945(.dina(n2200), .dinb(n2199), .dout(n2201));
  jand g01946(.dina(n2201), .dinb(n2198), .dout(n2202));
  jand g01947(.dina(n2202), .dinb(n2197), .dout(n2203));
  jxor g01948(.dina(n2203), .dinb(a20 ), .dout(n2204));
  jnot g01949(.din(n2204), .dout(n2205));
  jand g01950(.dina(n2080), .dinb(n2066), .dout(n2206));
  jand g01951(.dina(n2081), .dinb(n2057), .dout(n2207));
  jor  g01952(.dina(n2207), .dinb(n2206), .dout(n2208));
  jor  g01953(.dina(n1939), .dinb(n354), .dout(n2209));
  jor  g01954(.dina(n1827), .dinb(n299), .dout(n2210));
  jor  g01955(.dina(n1942), .dinb(n322), .dout(n2211));
  jor  g01956(.dina(n1944), .dinb(n357), .dout(n2212));
  jand g01957(.dina(n2212), .dinb(n2211), .dout(n2213));
  jand g01958(.dina(n2213), .dinb(n2210), .dout(n2214));
  jand g01959(.dina(n2214), .dinb(n2209), .dout(n2215));
  jxor g01960(.dina(n2215), .dinb(a23 ), .dout(n2216));
  jnot g01961(.din(n2216), .dout(n2217));
  jnot g01962(.din(n2079), .dout(n2218));
  jand g01963(.dina(n1953), .dinb(a26 ), .dout(n2219));
  jand g01964(.dina(n2219), .dinb(n2218), .dout(n2220));
  jnot g01965(.din(n2220), .dout(n2221));
  jand g01966(.dina(n2221), .dinb(a26 ), .dout(n2222));
  jor  g01967(.dina(n2073), .dinb(n2069), .dout(n2223));
  jor  g01968(.dina(n2223), .dinb(n1951), .dout(n2224));
  jnot g01969(.din(n2224), .dout(n2225));
  jand g01970(.dina(n2225), .dinb(b0 ), .dout(n2226));
  jand g01971(.dina(n2070), .dinb(b2 ), .dout(n2227));
  jand g01972(.dina(n2074), .dinb(b1 ), .dout(n2228));
  jand g01973(.dina(n2076), .dinb(n375), .dout(n2229));
  jor  g01974(.dina(n2229), .dinb(n2228), .dout(n2230));
  jor  g01975(.dina(n2230), .dinb(n2227), .dout(n2231));
  jor  g01976(.dina(n2231), .dinb(n2226), .dout(n2232));
  jxor g01977(.dina(n2232), .dinb(n2222), .dout(n2233));
  jxor g01978(.dina(n2233), .dinb(n2217), .dout(n2234));
  jxor g01979(.dina(n2234), .dinb(n2208), .dout(n2235));
  jxor g01980(.dina(n2235), .dinb(n2205), .dout(n2236));
  jxor g01981(.dina(n2236), .dinb(n2196), .dout(n2237));
  jxor g01982(.dina(n2237), .dinb(n2193), .dout(n2238));
  jxor g01983(.dina(n2238), .dinb(n2184), .dout(n2239));
  jnot g01984(.din(n2239), .dout(n2240));
  jor  g01985(.dina(n855), .dinb(n974), .dout(n2241));
  jor  g01986(.dina(n908), .dinb(n758), .dout(n2242));
  jor  g01987(.dina(n977), .dinb(n778), .dout(n2243));
  jor  g01988(.dina(n979), .dinb(n858), .dout(n2244));
  jand g01989(.dina(n2244), .dinb(n2243), .dout(n2245));
  jand g01990(.dina(n2245), .dinb(n2242), .dout(n2246));
  jand g01991(.dina(n2246), .dinb(n2241), .dout(n2247));
  jxor g01992(.dina(n2247), .dinb(a14 ), .dout(n2248));
  jxor g01993(.dina(n2248), .dinb(n2240), .dout(n2249));
  jxor g01994(.dina(n2249), .dinb(n2179), .dout(n2250));
  jxor g01995(.dina(n2250), .dinb(n2174), .dout(n2251));
  jnot g01996(.din(n2251), .dout(n2252));
  jxor g01997(.dina(n2252), .dinb(n2165), .dout(n2253));
  jor  g01998(.dina(n1417), .dinb(n528), .dout(n2254));
  jor  g01999(.dina(n490), .dinb(n1290), .dout(n2255));
  jor  g02000(.dina(n531), .dinb(n1400), .dout(n2256));
  jor  g02001(.dina(n533), .dinb(n1420), .dout(n2257));
  jand g02002(.dina(n2257), .dinb(n2256), .dout(n2258));
  jand g02003(.dina(n2258), .dinb(n2255), .dout(n2259));
  jand g02004(.dina(n2259), .dinb(n2254), .dout(n2260));
  jxor g02005(.dina(n2260), .dinb(a8 ), .dout(n2261));
  jxor g02006(.dina(n2261), .dinb(n2253), .dout(n2262));
  jxor g02007(.dina(n2262), .dinb(n2162), .dout(n2263));
  jor  g02008(.dina(n1864), .dinb(n402), .dout(n2264));
  jor  g02009(.dina(n371), .dinb(n1620), .dout(n2265));
  jor  g02010(.dina(n405), .dinb(n1742), .dout(n2266));
  jor  g02011(.dina(n332), .dinb(n1867), .dout(n2267));
  jand g02012(.dina(n2267), .dinb(n2266), .dout(n2268));
  jand g02013(.dina(n2268), .dinb(n2265), .dout(n2269));
  jand g02014(.dina(n2269), .dinb(n2264), .dout(n2270));
  jxor g02015(.dina(n2270), .dinb(a5 ), .dout(n2271));
  jxor g02016(.dina(n2271), .dinb(n2263), .dout(n2272));
  jxor g02017(.dina(n2272), .dinb(n2157), .dout(n2273));
  jxor g02018(.dina(n2273), .dinb(n2154), .dout(n2274));
  jxor g02019(.dina(n2274), .dinb(n2139), .dout(f26 ));
  jand g02020(.dina(n2273), .dinb(n2154), .dout(n2276));
  jand g02021(.dina(n2274), .dinb(n2139), .dout(n2277));
  jor  g02022(.dina(n2277), .dinb(n2276), .dout(n2278));
  jor  g02023(.dina(n2271), .dinb(n2263), .dout(n2279));
  jnot g02024(.din(n2279), .dout(n2280));
  jand g02025(.dina(n2272), .dinb(n2157), .dout(n2281));
  jor  g02026(.dina(n2281), .dinb(n2280), .dout(n2282));
  jand g02027(.dina(n2250), .dinb(n2174), .dout(n2283));
  jnot g02028(.din(n2283), .dout(n2284));
  jor  g02029(.dina(n2252), .dinb(n2165), .dout(n2285));
  jand g02030(.dina(n2285), .dinb(n2284), .dout(n2286));
  jor  g02031(.dina(n2248), .dinb(n2240), .dout(n2287));
  jand g02032(.dina(n2249), .dinb(n2179), .dout(n2288));
  jnot g02033(.din(n2288), .dout(n2289));
  jand g02034(.dina(n2289), .dinb(n2287), .dout(n2290));
  jnot g02035(.din(n2290), .dout(n2291));
  jand g02036(.dina(n2237), .dinb(n2193), .dout(n2292));
  jand g02037(.dina(n2238), .dinb(n2184), .dout(n2293));
  jor  g02038(.dina(n2293), .dinb(n2292), .dout(n2294));
  jor  g02039(.dina(n1245), .dinb(n755), .dout(n2295));
  jor  g02040(.dina(n1165), .dinb(n627), .dout(n2296));
  jor  g02041(.dina(n1248), .dinb(n647), .dout(n2297));
  jor  g02042(.dina(n1250), .dinb(n758), .dout(n2298));
  jand g02043(.dina(n2298), .dinb(n2297), .dout(n2299));
  jand g02044(.dina(n2299), .dinb(n2296), .dout(n2300));
  jand g02045(.dina(n2300), .dinb(n2295), .dout(n2301));
  jxor g02046(.dina(n2301), .dinb(a17 ), .dout(n2302));
  jnot g02047(.din(n2302), .dout(n2303));
  jand g02048(.dina(n2235), .dinb(n2205), .dout(n2304));
  jand g02049(.dina(n2236), .dinb(n2196), .dout(n2305));
  jor  g02050(.dina(n2305), .dinb(n2304), .dout(n2306));
  jor  g02051(.dina(n1566), .dinb(n561), .dout(n2307));
  jor  g02052(.dina(n1489), .dinb(n431), .dout(n2308));
  jor  g02053(.dina(n1569), .dinb(n512), .dout(n2309));
  jor  g02054(.dina(n1571), .dinb(n564), .dout(n2310));
  jand g02055(.dina(n2310), .dinb(n2309), .dout(n2311));
  jand g02056(.dina(n2311), .dinb(n2308), .dout(n2312));
  jand g02057(.dina(n2312), .dinb(n2307), .dout(n2313));
  jxor g02058(.dina(n2313), .dinb(a20 ), .dout(n2314));
  jnot g02059(.din(n2314), .dout(n2315));
  jand g02060(.dina(n2233), .dinb(n2217), .dout(n2316));
  jand g02061(.dina(n2234), .dinb(n2208), .dout(n2317));
  jor  g02062(.dina(n2317), .dinb(n2316), .dout(n2318));
  jnot g02063(.din(n2076), .dout(n2319));
  jor  g02064(.dina(n2319), .dinb(n296), .dout(n2320));
  jor  g02065(.dina(n2224), .dinb(n267), .dout(n2321));
  jnot g02066(.din(n2074), .dout(n2322));
  jor  g02067(.dina(n2322), .dinb(n279), .dout(n2323));
  jnot g02068(.din(n2070), .dout(n2324));
  jor  g02069(.dina(n2324), .dinb(n299), .dout(n2325));
  jand g02070(.dina(n2325), .dinb(n2323), .dout(n2326));
  jand g02071(.dina(n2326), .dinb(n2321), .dout(n2327));
  jand g02072(.dina(n2327), .dinb(n2320), .dout(n2328));
  jxor g02073(.dina(n2328), .dinb(a26 ), .dout(n2329));
  jnot g02074(.din(n2329), .dout(n2330));
  jxor g02075(.dina(a27 ), .dinb(a26 ), .dout(n2331));
  jand g02076(.dina(n2331), .dinb(b0 ), .dout(n2332));
  jnot g02077(.din(n2332), .dout(n2333));
  jor  g02078(.dina(n2232), .dinb(n2221), .dout(n2334));
  jxor g02079(.dina(n2334), .dinb(n2333), .dout(n2335));
  jxor g02080(.dina(n2335), .dinb(n2330), .dout(n2336));
  jnot g02081(.din(n2336), .dout(n2337));
  jor  g02082(.dina(n1939), .dinb(n392), .dout(n2338));
  jor  g02083(.dina(n1827), .dinb(n322), .dout(n2339));
  jor  g02084(.dina(n1942), .dinb(n357), .dout(n2340));
  jor  g02085(.dina(n1944), .dinb(n395), .dout(n2341));
  jand g02086(.dina(n2341), .dinb(n2340), .dout(n2342));
  jand g02087(.dina(n2342), .dinb(n2339), .dout(n2343));
  jand g02088(.dina(n2343), .dinb(n2338), .dout(n2344));
  jxor g02089(.dina(n2344), .dinb(a23 ), .dout(n2345));
  jxor g02090(.dina(n2345), .dinb(n2337), .dout(n2346));
  jxor g02091(.dina(n2346), .dinb(n2318), .dout(n2347));
  jxor g02092(.dina(n2347), .dinb(n2315), .dout(n2348));
  jxor g02093(.dina(n2348), .dinb(n2306), .dout(n2349));
  jxor g02094(.dina(n2349), .dinb(n2303), .dout(n2350));
  jxor g02095(.dina(n2350), .dinb(n2294), .dout(n2351));
  jnot g02096(.din(n2351), .dout(n2352));
  jor  g02097(.dina(n936), .dinb(n974), .dout(n2353));
  jor  g02098(.dina(n908), .dinb(n778), .dout(n2354));
  jor  g02099(.dina(n977), .dinb(n858), .dout(n2355));
  jor  g02100(.dina(n979), .dinb(n939), .dout(n2356));
  jand g02101(.dina(n2356), .dinb(n2355), .dout(n2357));
  jand g02102(.dina(n2357), .dinb(n2354), .dout(n2358));
  jand g02103(.dina(n2358), .dinb(n2353), .dout(n2359));
  jxor g02104(.dina(n2359), .dinb(a14 ), .dout(n2360));
  jxor g02105(.dina(n2360), .dinb(n2352), .dout(n2361));
  jxor g02106(.dina(n2361), .dinb(n2291), .dout(n2362));
  jor  g02107(.dina(n1287), .dinb(n706), .dout(n2363));
  jor  g02108(.dina(n683), .dinb(n1022), .dout(n2364));
  jor  g02109(.dina(n709), .dinb(n1193), .dout(n2365));
  jor  g02110(.dina(n711), .dinb(n1290), .dout(n2366));
  jand g02111(.dina(n2366), .dinb(n2365), .dout(n2367));
  jand g02112(.dina(n2367), .dinb(n2364), .dout(n2368));
  jand g02113(.dina(n2368), .dinb(n2363), .dout(n2369));
  jxor g02114(.dina(n2369), .dinb(a11 ), .dout(n2370));
  jxor g02115(.dina(n2370), .dinb(n2362), .dout(n2371));
  jxor g02116(.dina(n2371), .dinb(n2286), .dout(n2372));
  jor  g02117(.dina(n1617), .dinb(n528), .dout(n2373));
  jor  g02118(.dina(n490), .dinb(n1400), .dout(n2374));
  jor  g02119(.dina(n531), .dinb(n1420), .dout(n2375));
  jor  g02120(.dina(n533), .dinb(n1620), .dout(n2376));
  jand g02121(.dina(n2376), .dinb(n2375), .dout(n2377));
  jand g02122(.dina(n2377), .dinb(n2374), .dout(n2378));
  jand g02123(.dina(n2378), .dinb(n2373), .dout(n2379));
  jxor g02124(.dina(n2379), .dinb(a8 ), .dout(n2380));
  jxor g02125(.dina(n2380), .dinb(n2372), .dout(n2381));
  jnot g02126(.din(n2253), .dout(n2382));
  jor  g02127(.dina(n2261), .dinb(n2382), .dout(n2383));
  jnot g02128(.din(n2383), .dout(n2384));
  jnot g02129(.din(n2262), .dout(n2385));
  jand g02130(.dina(n2385), .dinb(n2162), .dout(n2386));
  jor  g02131(.dina(n2386), .dinb(n2384), .dout(n2387));
  jxor g02132(.dina(n2387), .dinb(n2381), .dout(n2388));
  jor  g02133(.dina(n1884), .dinb(n402), .dout(n2389));
  jor  g02134(.dina(n371), .dinb(n1742), .dout(n2390));
  jor  g02135(.dina(n405), .dinb(n1867), .dout(n2391));
  jor  g02136(.dina(n332), .dinb(n1887), .dout(n2392));
  jand g02137(.dina(n2392), .dinb(n2391), .dout(n2393));
  jand g02138(.dina(n2393), .dinb(n2390), .dout(n2394));
  jand g02139(.dina(n2394), .dinb(n2389), .dout(n2395));
  jxor g02140(.dina(n2395), .dinb(a5 ), .dout(n2396));
  jxor g02141(.dina(n2396), .dinb(n2388), .dout(n2397));
  jxor g02142(.dina(n2397), .dinb(n2282), .dout(n2398));
  jand g02143(.dina(b26 ), .dinb(b25 ), .dout(n2399));
  jand g02144(.dina(n2143), .dinb(n2142), .dout(n2400));
  jor  g02145(.dina(n2400), .dinb(n2399), .dout(n2401));
  jxor g02146(.dina(b27 ), .dinb(b26 ), .dout(n2402));
  jnot g02147(.din(n2402), .dout(n2403));
  jxor g02148(.dina(n2403), .dinb(n2401), .dout(n2404));
  jor  g02149(.dina(n2404), .dinb(n264), .dout(n2405));
  jor  g02150(.dina(n284), .dinb(n2010), .dout(n2406));
  jnot g02151(.din(b27 ), .dout(n2407));
  jor  g02152(.dina(n269), .dinb(n2407), .dout(n2408));
  jor  g02153(.dina(n271), .dinb(n2148), .dout(n2409));
  jand g02154(.dina(n2409), .dinb(n2408), .dout(n2410));
  jand g02155(.dina(n2410), .dinb(n2406), .dout(n2411));
  jand g02156(.dina(n2411), .dinb(n2405), .dout(n2412));
  jxor g02157(.dina(n2412), .dinb(n260), .dout(n2413));
  jxor g02158(.dina(n2413), .dinb(n2398), .dout(n2414));
  jxor g02159(.dina(n2414), .dinb(n2278), .dout(f27 ));
  jand g02160(.dina(n2413), .dinb(n2398), .dout(n2416));
  jand g02161(.dina(n2414), .dinb(n2278), .dout(n2417));
  jor  g02162(.dina(n2417), .dinb(n2416), .dout(n2418));
  jor  g02163(.dina(n2396), .dinb(n2388), .dout(n2419));
  jnot g02164(.din(n2419), .dout(n2420));
  jand g02165(.dina(n2397), .dinb(n2282), .dout(n2421));
  jor  g02166(.dina(n2421), .dinb(n2420), .dout(n2422));
  jnot g02167(.din(n2362), .dout(n2423));
  jor  g02168(.dina(n2370), .dinb(n2423), .dout(n2424));
  jor  g02169(.dina(n2371), .dinb(n2286), .dout(n2425));
  jand g02170(.dina(n2425), .dinb(n2424), .dout(n2426));
  jor  g02171(.dina(n2360), .dinb(n2352), .dout(n2427));
  jnot g02172(.din(n2427), .dout(n2428));
  jand g02173(.dina(n2361), .dinb(n2291), .dout(n2429));
  jor  g02174(.dina(n2429), .dinb(n2428), .dout(n2430));
  jor  g02175(.dina(n1019), .dinb(n974), .dout(n2431));
  jor  g02176(.dina(n908), .dinb(n858), .dout(n2432));
  jor  g02177(.dina(n977), .dinb(n939), .dout(n2433));
  jor  g02178(.dina(n979), .dinb(n1022), .dout(n2434));
  jand g02179(.dina(n2434), .dinb(n2433), .dout(n2435));
  jand g02180(.dina(n2435), .dinb(n2432), .dout(n2436));
  jand g02181(.dina(n2436), .dinb(n2431), .dout(n2437));
  jxor g02182(.dina(n2437), .dinb(a14 ), .dout(n2438));
  jnot g02183(.din(n2438), .dout(n2439));
  jand g02184(.dina(n2349), .dinb(n2303), .dout(n2440));
  jand g02185(.dina(n2350), .dinb(n2294), .dout(n2441));
  jor  g02186(.dina(n2441), .dinb(n2440), .dout(n2442));
  jand g02187(.dina(n2347), .dinb(n2315), .dout(n2443));
  jand g02188(.dina(n2348), .dinb(n2306), .dout(n2444));
  jor  g02189(.dina(n2444), .dinb(n2443), .dout(n2445));
  jor  g02190(.dina(n2345), .dinb(n2337), .dout(n2446));
  jand g02191(.dina(n2346), .dinb(n2318), .dout(n2447));
  jnot g02192(.din(n2447), .dout(n2448));
  jand g02193(.dina(n2448), .dinb(n2446), .dout(n2449));
  jnot g02194(.din(n2449), .dout(n2450));
  jor  g02195(.dina(n1939), .dinb(n428), .dout(n2451));
  jor  g02196(.dina(n1827), .dinb(n357), .dout(n2452));
  jor  g02197(.dina(n1942), .dinb(n395), .dout(n2453));
  jor  g02198(.dina(n1944), .dinb(n431), .dout(n2454));
  jand g02199(.dina(n2454), .dinb(n2453), .dout(n2455));
  jand g02200(.dina(n2455), .dinb(n2452), .dout(n2456));
  jand g02201(.dina(n2456), .dinb(n2451), .dout(n2457));
  jxor g02202(.dina(n2457), .dinb(a23 ), .dout(n2458));
  jnot g02203(.din(n2458), .dout(n2459));
  jnot g02204(.din(n2334), .dout(n2460));
  jand g02205(.dina(n2460), .dinb(n2332), .dout(n2461));
  jand g02206(.dina(n2335), .dinb(n2330), .dout(n2462));
  jor  g02207(.dina(n2462), .dinb(n2461), .dout(n2463));
  jor  g02208(.dina(n2319), .dinb(n319), .dout(n2464));
  jor  g02209(.dina(n2224), .dinb(n279), .dout(n2465));
  jor  g02210(.dina(n2322), .dinb(n299), .dout(n2466));
  jor  g02211(.dina(n2324), .dinb(n322), .dout(n2467));
  jand g02212(.dina(n2467), .dinb(n2466), .dout(n2468));
  jand g02213(.dina(n2468), .dinb(n2465), .dout(n2469));
  jand g02214(.dina(n2469), .dinb(n2464), .dout(n2470));
  jxor g02215(.dina(n2470), .dinb(a26 ), .dout(n2471));
  jnot g02216(.din(n2471), .dout(n2472));
  jand g02217(.dina(n2332), .dinb(a29 ), .dout(n2473));
  jxor g02218(.dina(a29 ), .dinb(a28 ), .dout(n2474));
  jnot g02219(.din(n2474), .dout(n2475));
  jand g02220(.dina(n2475), .dinb(n2331), .dout(n2476));
  jand g02221(.dina(n2476), .dinb(b1 ), .dout(n2477));
  jnot g02222(.din(n2331), .dout(n2478));
  jxor g02223(.dina(a28 ), .dinb(a27 ), .dout(n2479));
  jand g02224(.dina(n2479), .dinb(n2478), .dout(n2480));
  jand g02225(.dina(n2480), .dinb(b0 ), .dout(n2481));
  jand g02226(.dina(n2474), .dinb(n2331), .dout(n2482));
  jand g02227(.dina(n2482), .dinb(n338), .dout(n2483));
  jor  g02228(.dina(n2483), .dinb(n2481), .dout(n2484));
  jor  g02229(.dina(n2484), .dinb(n2477), .dout(n2485));
  jxor g02230(.dina(n2485), .dinb(n2473), .dout(n2486));
  jxor g02231(.dina(n2486), .dinb(n2472), .dout(n2487));
  jxor g02232(.dina(n2487), .dinb(n2463), .dout(n2488));
  jxor g02233(.dina(n2488), .dinb(n2459), .dout(n2489));
  jxor g02234(.dina(n2489), .dinb(n2450), .dout(n2490));
  jnot g02235(.din(n2490), .dout(n2491));
  jor  g02236(.dina(n1566), .dinb(n624), .dout(n2492));
  jor  g02237(.dina(n1489), .dinb(n512), .dout(n2493));
  jor  g02238(.dina(n1569), .dinb(n564), .dout(n2494));
  jor  g02239(.dina(n1571), .dinb(n627), .dout(n2495));
  jand g02240(.dina(n2495), .dinb(n2494), .dout(n2496));
  jand g02241(.dina(n2496), .dinb(n2493), .dout(n2497));
  jand g02242(.dina(n2497), .dinb(n2492), .dout(n2498));
  jxor g02243(.dina(n2498), .dinb(a20 ), .dout(n2499));
  jxor g02244(.dina(n2499), .dinb(n2491), .dout(n2500));
  jxor g02245(.dina(n2500), .dinb(n2445), .dout(n2501));
  jnot g02246(.din(n2501), .dout(n2502));
  jor  g02247(.dina(n1245), .dinb(n775), .dout(n2503));
  jor  g02248(.dina(n1165), .dinb(n647), .dout(n2504));
  jor  g02249(.dina(n1248), .dinb(n758), .dout(n2505));
  jor  g02250(.dina(n1250), .dinb(n778), .dout(n2506));
  jand g02251(.dina(n2506), .dinb(n2505), .dout(n2507));
  jand g02252(.dina(n2507), .dinb(n2504), .dout(n2508));
  jand g02253(.dina(n2508), .dinb(n2503), .dout(n2509));
  jxor g02254(.dina(n2509), .dinb(a17 ), .dout(n2510));
  jxor g02255(.dina(n2510), .dinb(n2502), .dout(n2511));
  jxor g02256(.dina(n2511), .dinb(n2442), .dout(n2512));
  jxor g02257(.dina(n2512), .dinb(n2439), .dout(n2513));
  jxor g02258(.dina(n2513), .dinb(n2430), .dout(n2514));
  jor  g02259(.dina(n1397), .dinb(n706), .dout(n2515));
  jor  g02260(.dina(n683), .dinb(n1193), .dout(n2516));
  jor  g02261(.dina(n709), .dinb(n1290), .dout(n2517));
  jor  g02262(.dina(n711), .dinb(n1400), .dout(n2518));
  jand g02263(.dina(n2518), .dinb(n2517), .dout(n2519));
  jand g02264(.dina(n2519), .dinb(n2516), .dout(n2520));
  jand g02265(.dina(n2520), .dinb(n2515), .dout(n2521));
  jxor g02266(.dina(n2521), .dinb(a11 ), .dout(n2522));
  jxor g02267(.dina(n2522), .dinb(n2514), .dout(n2523));
  jxor g02268(.dina(n2523), .dinb(n2426), .dout(n2524));
  jor  g02269(.dina(n1739), .dinb(n528), .dout(n2525));
  jor  g02270(.dina(n490), .dinb(n1420), .dout(n2526));
  jor  g02271(.dina(n531), .dinb(n1620), .dout(n2527));
  jor  g02272(.dina(n533), .dinb(n1742), .dout(n2528));
  jand g02273(.dina(n2528), .dinb(n2527), .dout(n2529));
  jand g02274(.dina(n2529), .dinb(n2526), .dout(n2530));
  jand g02275(.dina(n2530), .dinb(n2525), .dout(n2531));
  jxor g02276(.dina(n2531), .dinb(a8 ), .dout(n2532));
  jxor g02277(.dina(n2532), .dinb(n2524), .dout(n2533));
  jnot g02278(.din(n2372), .dout(n2534));
  jor  g02279(.dina(n2380), .dinb(n2534), .dout(n2535));
  jnot g02280(.din(n2535), .dout(n2536));
  jnot g02281(.din(n2381), .dout(n2537));
  jand g02282(.dina(n2387), .dinb(n2537), .dout(n2538));
  jor  g02283(.dina(n2538), .dinb(n2536), .dout(n2539));
  jxor g02284(.dina(n2539), .dinb(n2533), .dout(n2540));
  jor  g02285(.dina(n2007), .dinb(n402), .dout(n2541));
  jor  g02286(.dina(n371), .dinb(n1867), .dout(n2542));
  jor  g02287(.dina(n405), .dinb(n1887), .dout(n2543));
  jor  g02288(.dina(n332), .dinb(n2010), .dout(n2544));
  jand g02289(.dina(n2544), .dinb(n2543), .dout(n2545));
  jand g02290(.dina(n2545), .dinb(n2542), .dout(n2546));
  jand g02291(.dina(n2546), .dinb(n2541), .dout(n2547));
  jxor g02292(.dina(n2547), .dinb(a5 ), .dout(n2548));
  jxor g02293(.dina(n2548), .dinb(n2540), .dout(n2549));
  jxor g02294(.dina(n2549), .dinb(n2422), .dout(n2550));
  jand g02295(.dina(b27 ), .dinb(b26 ), .dout(n2551));
  jand g02296(.dina(n2402), .dinb(n2401), .dout(n2552));
  jor  g02297(.dina(n2552), .dinb(n2551), .dout(n2553));
  jxor g02298(.dina(b28 ), .dinb(b27 ), .dout(n2554));
  jnot g02299(.din(n2554), .dout(n2555));
  jxor g02300(.dina(n2555), .dinb(n2553), .dout(n2556));
  jor  g02301(.dina(n2556), .dinb(n264), .dout(n2557));
  jor  g02302(.dina(n284), .dinb(n2148), .dout(n2558));
  jnot g02303(.din(b28 ), .dout(n2559));
  jor  g02304(.dina(n269), .dinb(n2559), .dout(n2560));
  jor  g02305(.dina(n271), .dinb(n2407), .dout(n2561));
  jand g02306(.dina(n2561), .dinb(n2560), .dout(n2562));
  jand g02307(.dina(n2562), .dinb(n2558), .dout(n2563));
  jand g02308(.dina(n2563), .dinb(n2557), .dout(n2564));
  jxor g02309(.dina(n2564), .dinb(n260), .dout(n2565));
  jxor g02310(.dina(n2565), .dinb(n2550), .dout(n2566));
  jxor g02311(.dina(n2566), .dinb(n2418), .dout(f28 ));
  jand g02312(.dina(n2565), .dinb(n2550), .dout(n2568));
  jand g02313(.dina(n2566), .dinb(n2418), .dout(n2569));
  jor  g02314(.dina(n2569), .dinb(n2568), .dout(n2570));
  jand g02315(.dina(b28 ), .dinb(b27 ), .dout(n2571));
  jand g02316(.dina(n2554), .dinb(n2553), .dout(n2572));
  jor  g02317(.dina(n2572), .dinb(n2571), .dout(n2573));
  jxor g02318(.dina(b29 ), .dinb(b28 ), .dout(n2574));
  jnot g02319(.din(n2574), .dout(n2575));
  jxor g02320(.dina(n2575), .dinb(n2573), .dout(n2576));
  jor  g02321(.dina(n2576), .dinb(n264), .dout(n2577));
  jor  g02322(.dina(n284), .dinb(n2407), .dout(n2578));
  jnot g02323(.din(b29 ), .dout(n2579));
  jor  g02324(.dina(n269), .dinb(n2579), .dout(n2580));
  jor  g02325(.dina(n271), .dinb(n2559), .dout(n2581));
  jand g02326(.dina(n2581), .dinb(n2580), .dout(n2582));
  jand g02327(.dina(n2582), .dinb(n2578), .dout(n2583));
  jand g02328(.dina(n2583), .dinb(n2577), .dout(n2584));
  jxor g02329(.dina(n2584), .dinb(n260), .dout(n2585));
  jor  g02330(.dina(n2548), .dinb(n2540), .dout(n2586));
  jnot g02331(.din(n2586), .dout(n2587));
  jand g02332(.dina(n2549), .dinb(n2422), .dout(n2588));
  jor  g02333(.dina(n2588), .dinb(n2587), .dout(n2589));
  jor  g02334(.dina(n2145), .dinb(n402), .dout(n2590));
  jor  g02335(.dina(n371), .dinb(n1887), .dout(n2591));
  jor  g02336(.dina(n405), .dinb(n2010), .dout(n2592));
  jor  g02337(.dina(n332), .dinb(n2148), .dout(n2593));
  jand g02338(.dina(n2593), .dinb(n2592), .dout(n2594));
  jand g02339(.dina(n2594), .dinb(n2591), .dout(n2595));
  jand g02340(.dina(n2595), .dinb(n2590), .dout(n2596));
  jxor g02341(.dina(n2596), .dinb(a5 ), .dout(n2597));
  jnot g02342(.din(n2597), .dout(n2598));
  jnot g02343(.din(n2524), .dout(n2599));
  jor  g02344(.dina(n2532), .dinb(n2599), .dout(n2600));
  jnot g02345(.din(n2600), .dout(n2601));
  jnot g02346(.din(n2533), .dout(n2602));
  jand g02347(.dina(n2539), .dinb(n2602), .dout(n2603));
  jor  g02348(.dina(n2603), .dinb(n2601), .dout(n2604));
  jnot g02349(.din(n2514), .dout(n2605));
  jor  g02350(.dina(n2522), .dinb(n2605), .dout(n2606));
  jor  g02351(.dina(n2523), .dinb(n2426), .dout(n2607));
  jand g02352(.dina(n2607), .dinb(n2606), .dout(n2608));
  jand g02353(.dina(n2512), .dinb(n2439), .dout(n2609));
  jand g02354(.dina(n2513), .dinb(n2430), .dout(n2610));
  jor  g02355(.dina(n2610), .dinb(n2609), .dout(n2611));
  jor  g02356(.dina(n2510), .dinb(n2502), .dout(n2612));
  jand g02357(.dina(n2511), .dinb(n2442), .dout(n2613));
  jnot g02358(.din(n2613), .dout(n2614));
  jand g02359(.dina(n2614), .dinb(n2612), .dout(n2615));
  jnot g02360(.din(n2615), .dout(n2616));
  jor  g02361(.dina(n2499), .dinb(n2491), .dout(n2617));
  jand g02362(.dina(n2500), .dinb(n2445), .dout(n2618));
  jnot g02363(.din(n2618), .dout(n2619));
  jand g02364(.dina(n2619), .dinb(n2617), .dout(n2620));
  jnot g02365(.din(n2620), .dout(n2621));
  jor  g02366(.dina(n1566), .dinb(n644), .dout(n2622));
  jor  g02367(.dina(n1489), .dinb(n564), .dout(n2623));
  jor  g02368(.dina(n1569), .dinb(n627), .dout(n2624));
  jor  g02369(.dina(n1571), .dinb(n647), .dout(n2625));
  jand g02370(.dina(n2625), .dinb(n2624), .dout(n2626));
  jand g02371(.dina(n2626), .dinb(n2623), .dout(n2627));
  jand g02372(.dina(n2627), .dinb(n2622), .dout(n2628));
  jxor g02373(.dina(n2628), .dinb(a20 ), .dout(n2629));
  jnot g02374(.din(n2629), .dout(n2630));
  jand g02375(.dina(n2488), .dinb(n2459), .dout(n2631));
  jand g02376(.dina(n2489), .dinb(n2450), .dout(n2632));
  jor  g02377(.dina(n2632), .dinb(n2631), .dout(n2633));
  jor  g02378(.dina(n1939), .dinb(n509), .dout(n2634));
  jor  g02379(.dina(n1827), .dinb(n395), .dout(n2635));
  jor  g02380(.dina(n1942), .dinb(n431), .dout(n2636));
  jor  g02381(.dina(n1944), .dinb(n512), .dout(n2637));
  jand g02382(.dina(n2637), .dinb(n2636), .dout(n2638));
  jand g02383(.dina(n2638), .dinb(n2635), .dout(n2639));
  jand g02384(.dina(n2639), .dinb(n2634), .dout(n2640));
  jxor g02385(.dina(n2640), .dinb(a23 ), .dout(n2641));
  jnot g02386(.din(n2641), .dout(n2642));
  jand g02387(.dina(n2486), .dinb(n2472), .dout(n2643));
  jand g02388(.dina(n2487), .dinb(n2463), .dout(n2644));
  jor  g02389(.dina(n2644), .dinb(n2643), .dout(n2645));
  jor  g02390(.dina(n2319), .dinb(n354), .dout(n2646));
  jor  g02391(.dina(n2224), .dinb(n299), .dout(n2647));
  jor  g02392(.dina(n2322), .dinb(n322), .dout(n2648));
  jor  g02393(.dina(n2324), .dinb(n357), .dout(n2649));
  jand g02394(.dina(n2649), .dinb(n2648), .dout(n2650));
  jand g02395(.dina(n2650), .dinb(n2647), .dout(n2651));
  jand g02396(.dina(n2651), .dinb(n2646), .dout(n2652));
  jxor g02397(.dina(n2652), .dinb(a26 ), .dout(n2653));
  jnot g02398(.din(n2653), .dout(n2654));
  jnot g02399(.din(n2485), .dout(n2655));
  jand g02400(.dina(n2333), .dinb(a29 ), .dout(n2656));
  jand g02401(.dina(n2656), .dinb(n2655), .dout(n2657));
  jnot g02402(.din(n2657), .dout(n2658));
  jand g02403(.dina(n2658), .dinb(a29 ), .dout(n2659));
  jor  g02404(.dina(n2479), .dinb(n2475), .dout(n2660));
  jor  g02405(.dina(n2660), .dinb(n2331), .dout(n2661));
  jnot g02406(.din(n2661), .dout(n2662));
  jand g02407(.dina(n2662), .dinb(b0 ), .dout(n2663));
  jand g02408(.dina(n2476), .dinb(b2 ), .dout(n2664));
  jand g02409(.dina(n2480), .dinb(b1 ), .dout(n2665));
  jand g02410(.dina(n2482), .dinb(n375), .dout(n2666));
  jor  g02411(.dina(n2666), .dinb(n2665), .dout(n2667));
  jor  g02412(.dina(n2667), .dinb(n2664), .dout(n2668));
  jor  g02413(.dina(n2668), .dinb(n2663), .dout(n2669));
  jxor g02414(.dina(n2669), .dinb(n2659), .dout(n2670));
  jxor g02415(.dina(n2670), .dinb(n2654), .dout(n2671));
  jxor g02416(.dina(n2671), .dinb(n2645), .dout(n2672));
  jxor g02417(.dina(n2672), .dinb(n2642), .dout(n2673));
  jxor g02418(.dina(n2673), .dinb(n2633), .dout(n2674));
  jxor g02419(.dina(n2674), .dinb(n2630), .dout(n2675));
  jxor g02420(.dina(n2675), .dinb(n2621), .dout(n2676));
  jnot g02421(.din(n2676), .dout(n2677));
  jor  g02422(.dina(n1245), .dinb(n855), .dout(n2678));
  jor  g02423(.dina(n1165), .dinb(n758), .dout(n2679));
  jor  g02424(.dina(n1248), .dinb(n778), .dout(n2680));
  jor  g02425(.dina(n1250), .dinb(n858), .dout(n2681));
  jand g02426(.dina(n2681), .dinb(n2680), .dout(n2682));
  jand g02427(.dina(n2682), .dinb(n2679), .dout(n2683));
  jand g02428(.dina(n2683), .dinb(n2678), .dout(n2684));
  jxor g02429(.dina(n2684), .dinb(a17 ), .dout(n2685));
  jxor g02430(.dina(n2685), .dinb(n2677), .dout(n2686));
  jxor g02431(.dina(n2686), .dinb(n2616), .dout(n2687));
  jnot g02432(.din(n2687), .dout(n2688));
  jor  g02433(.dina(n1190), .dinb(n974), .dout(n2689));
  jor  g02434(.dina(n908), .dinb(n939), .dout(n2690));
  jor  g02435(.dina(n977), .dinb(n1022), .dout(n2691));
  jor  g02436(.dina(n979), .dinb(n1193), .dout(n2692));
  jand g02437(.dina(n2692), .dinb(n2691), .dout(n2693));
  jand g02438(.dina(n2693), .dinb(n2690), .dout(n2694));
  jand g02439(.dina(n2694), .dinb(n2689), .dout(n2695));
  jxor g02440(.dina(n2695), .dinb(a14 ), .dout(n2696));
  jxor g02441(.dina(n2696), .dinb(n2688), .dout(n2697));
  jxor g02442(.dina(n2697), .dinb(n2611), .dout(n2698));
  jor  g02443(.dina(n1417), .dinb(n706), .dout(n2699));
  jor  g02444(.dina(n683), .dinb(n1290), .dout(n2700));
  jor  g02445(.dina(n709), .dinb(n1400), .dout(n2701));
  jor  g02446(.dina(n711), .dinb(n1420), .dout(n2702));
  jand g02447(.dina(n2702), .dinb(n2701), .dout(n2703));
  jand g02448(.dina(n2703), .dinb(n2700), .dout(n2704));
  jand g02449(.dina(n2704), .dinb(n2699), .dout(n2705));
  jxor g02450(.dina(n2705), .dinb(a11 ), .dout(n2706));
  jxor g02451(.dina(n2706), .dinb(n2698), .dout(n2707));
  jxor g02452(.dina(n2707), .dinb(n2608), .dout(n2708));
  jor  g02453(.dina(n1864), .dinb(n528), .dout(n2709));
  jor  g02454(.dina(n490), .dinb(n1620), .dout(n2710));
  jor  g02455(.dina(n531), .dinb(n1742), .dout(n2711));
  jor  g02456(.dina(n533), .dinb(n1867), .dout(n2712));
  jand g02457(.dina(n2712), .dinb(n2711), .dout(n2713));
  jand g02458(.dina(n2713), .dinb(n2710), .dout(n2714));
  jand g02459(.dina(n2714), .dinb(n2709), .dout(n2715));
  jxor g02460(.dina(n2715), .dinb(a8 ), .dout(n2716));
  jxor g02461(.dina(n2716), .dinb(n2708), .dout(n2717));
  jnot g02462(.din(n2717), .dout(n2718));
  jxor g02463(.dina(n2718), .dinb(n2604), .dout(n2719));
  jxor g02464(.dina(n2719), .dinb(n2598), .dout(n2720));
  jxor g02465(.dina(n2720), .dinb(n2589), .dout(n2721));
  jxor g02466(.dina(n2721), .dinb(n2585), .dout(n2722));
  jxor g02467(.dina(n2722), .dinb(n2570), .dout(f29 ));
  jand g02468(.dina(n2721), .dinb(n2585), .dout(n2724));
  jand g02469(.dina(n2722), .dinb(n2570), .dout(n2725));
  jor  g02470(.dina(n2725), .dinb(n2724), .dout(n2726));
  jand g02471(.dina(n2719), .dinb(n2598), .dout(n2727));
  jand g02472(.dina(n2720), .dinb(n2589), .dout(n2728));
  jor  g02473(.dina(n2728), .dinb(n2727), .dout(n2729));
  jnot g02474(.din(n2708), .dout(n2730));
  jor  g02475(.dina(n2716), .dinb(n2730), .dout(n2731));
  jnot g02476(.din(n2731), .dout(n2732));
  jand g02477(.dina(n2718), .dinb(n2604), .dout(n2733));
  jor  g02478(.dina(n2733), .dinb(n2732), .dout(n2734));
  jor  g02479(.dina(n1884), .dinb(n528), .dout(n2735));
  jor  g02480(.dina(n490), .dinb(n1742), .dout(n2736));
  jor  g02481(.dina(n531), .dinb(n1867), .dout(n2737));
  jor  g02482(.dina(n533), .dinb(n1887), .dout(n2738));
  jand g02483(.dina(n2738), .dinb(n2737), .dout(n2739));
  jand g02484(.dina(n2739), .dinb(n2736), .dout(n2740));
  jand g02485(.dina(n2740), .dinb(n2735), .dout(n2741));
  jxor g02486(.dina(n2741), .dinb(a8 ), .dout(n2742));
  jnot g02487(.din(n2742), .dout(n2743));
  jnot g02488(.din(n2698), .dout(n2744));
  jor  g02489(.dina(n2706), .dinb(n2744), .dout(n2745));
  jor  g02490(.dina(n2707), .dinb(n2608), .dout(n2746));
  jand g02491(.dina(n2746), .dinb(n2745), .dout(n2747));
  jor  g02492(.dina(n2696), .dinb(n2688), .dout(n2748));
  jnot g02493(.din(n2748), .dout(n2749));
  jand g02494(.dina(n2697), .dinb(n2611), .dout(n2750));
  jor  g02495(.dina(n2750), .dinb(n2749), .dout(n2751));
  jor  g02496(.dina(n2685), .dinb(n2677), .dout(n2752));
  jand g02497(.dina(n2686), .dinb(n2616), .dout(n2753));
  jnot g02498(.din(n2753), .dout(n2754));
  jand g02499(.dina(n2754), .dinb(n2752), .dout(n2755));
  jnot g02500(.din(n2755), .dout(n2756));
  jand g02501(.dina(n2674), .dinb(n2630), .dout(n2757));
  jand g02502(.dina(n2675), .dinb(n2621), .dout(n2758));
  jor  g02503(.dina(n2758), .dinb(n2757), .dout(n2759));
  jor  g02504(.dina(n1566), .dinb(n755), .dout(n2760));
  jor  g02505(.dina(n1489), .dinb(n627), .dout(n2761));
  jor  g02506(.dina(n1569), .dinb(n647), .dout(n2762));
  jor  g02507(.dina(n1571), .dinb(n758), .dout(n2763));
  jand g02508(.dina(n2763), .dinb(n2762), .dout(n2764));
  jand g02509(.dina(n2764), .dinb(n2761), .dout(n2765));
  jand g02510(.dina(n2765), .dinb(n2760), .dout(n2766));
  jxor g02511(.dina(n2766), .dinb(a20 ), .dout(n2767));
  jnot g02512(.din(n2767), .dout(n2768));
  jand g02513(.dina(n2672), .dinb(n2642), .dout(n2769));
  jand g02514(.dina(n2673), .dinb(n2633), .dout(n2770));
  jor  g02515(.dina(n2770), .dinb(n2769), .dout(n2771));
  jor  g02516(.dina(n1939), .dinb(n561), .dout(n2772));
  jor  g02517(.dina(n1827), .dinb(n431), .dout(n2773));
  jor  g02518(.dina(n1942), .dinb(n512), .dout(n2774));
  jor  g02519(.dina(n1944), .dinb(n564), .dout(n2775));
  jand g02520(.dina(n2775), .dinb(n2774), .dout(n2776));
  jand g02521(.dina(n2776), .dinb(n2773), .dout(n2777));
  jand g02522(.dina(n2777), .dinb(n2772), .dout(n2778));
  jxor g02523(.dina(n2778), .dinb(a23 ), .dout(n2779));
  jnot g02524(.din(n2779), .dout(n2780));
  jand g02525(.dina(n2670), .dinb(n2654), .dout(n2781));
  jand g02526(.dina(n2671), .dinb(n2645), .dout(n2782));
  jor  g02527(.dina(n2782), .dinb(n2781), .dout(n2783));
  jnot g02528(.din(n2482), .dout(n2784));
  jor  g02529(.dina(n2784), .dinb(n296), .dout(n2785));
  jor  g02530(.dina(n2661), .dinb(n267), .dout(n2786));
  jnot g02531(.din(n2480), .dout(n2787));
  jor  g02532(.dina(n2787), .dinb(n279), .dout(n2788));
  jnot g02533(.din(n2476), .dout(n2789));
  jor  g02534(.dina(n2789), .dinb(n299), .dout(n2790));
  jand g02535(.dina(n2790), .dinb(n2788), .dout(n2791));
  jand g02536(.dina(n2791), .dinb(n2786), .dout(n2792));
  jand g02537(.dina(n2792), .dinb(n2785), .dout(n2793));
  jxor g02538(.dina(n2793), .dinb(a29 ), .dout(n2794));
  jnot g02539(.din(n2794), .dout(n2795));
  jxor g02540(.dina(a30 ), .dinb(a29 ), .dout(n2796));
  jand g02541(.dina(n2796), .dinb(b0 ), .dout(n2797));
  jnot g02542(.din(n2797), .dout(n2798));
  jor  g02543(.dina(n2669), .dinb(n2658), .dout(n2799));
  jxor g02544(.dina(n2799), .dinb(n2798), .dout(n2800));
  jxor g02545(.dina(n2800), .dinb(n2795), .dout(n2801));
  jnot g02546(.din(n2801), .dout(n2802));
  jor  g02547(.dina(n2319), .dinb(n392), .dout(n2803));
  jor  g02548(.dina(n2224), .dinb(n322), .dout(n2804));
  jor  g02549(.dina(n2322), .dinb(n357), .dout(n2805));
  jor  g02550(.dina(n2324), .dinb(n395), .dout(n2806));
  jand g02551(.dina(n2806), .dinb(n2805), .dout(n2807));
  jand g02552(.dina(n2807), .dinb(n2804), .dout(n2808));
  jand g02553(.dina(n2808), .dinb(n2803), .dout(n2809));
  jxor g02554(.dina(n2809), .dinb(a26 ), .dout(n2810));
  jxor g02555(.dina(n2810), .dinb(n2802), .dout(n2811));
  jxor g02556(.dina(n2811), .dinb(n2783), .dout(n2812));
  jxor g02557(.dina(n2812), .dinb(n2780), .dout(n2813));
  jxor g02558(.dina(n2813), .dinb(n2771), .dout(n2814));
  jxor g02559(.dina(n2814), .dinb(n2768), .dout(n2815));
  jxor g02560(.dina(n2815), .dinb(n2759), .dout(n2816));
  jnot g02561(.din(n2816), .dout(n2817));
  jor  g02562(.dina(n1245), .dinb(n936), .dout(n2818));
  jor  g02563(.dina(n1165), .dinb(n778), .dout(n2819));
  jor  g02564(.dina(n1248), .dinb(n858), .dout(n2820));
  jor  g02565(.dina(n1250), .dinb(n939), .dout(n2821));
  jand g02566(.dina(n2821), .dinb(n2820), .dout(n2822));
  jand g02567(.dina(n2822), .dinb(n2819), .dout(n2823));
  jand g02568(.dina(n2823), .dinb(n2818), .dout(n2824));
  jxor g02569(.dina(n2824), .dinb(a17 ), .dout(n2825));
  jxor g02570(.dina(n2825), .dinb(n2817), .dout(n2826));
  jxor g02571(.dina(n2826), .dinb(n2756), .dout(n2827));
  jnot g02572(.din(n2827), .dout(n2828));
  jor  g02573(.dina(n1287), .dinb(n974), .dout(n2829));
  jor  g02574(.dina(n908), .dinb(n1022), .dout(n2830));
  jor  g02575(.dina(n977), .dinb(n1193), .dout(n2831));
  jor  g02576(.dina(n979), .dinb(n1290), .dout(n2832));
  jand g02577(.dina(n2832), .dinb(n2831), .dout(n2833));
  jand g02578(.dina(n2833), .dinb(n2830), .dout(n2834));
  jand g02579(.dina(n2834), .dinb(n2829), .dout(n2835));
  jxor g02580(.dina(n2835), .dinb(a14 ), .dout(n2836));
  jxor g02581(.dina(n2836), .dinb(n2828), .dout(n2837));
  jxor g02582(.dina(n2837), .dinb(n2751), .dout(n2838));
  jor  g02583(.dina(n1617), .dinb(n706), .dout(n2839));
  jor  g02584(.dina(n683), .dinb(n1400), .dout(n2840));
  jor  g02585(.dina(n709), .dinb(n1420), .dout(n2841));
  jor  g02586(.dina(n711), .dinb(n1620), .dout(n2842));
  jand g02587(.dina(n2842), .dinb(n2841), .dout(n2843));
  jand g02588(.dina(n2843), .dinb(n2840), .dout(n2844));
  jand g02589(.dina(n2844), .dinb(n2839), .dout(n2845));
  jxor g02590(.dina(n2845), .dinb(a11 ), .dout(n2846));
  jxor g02591(.dina(n2846), .dinb(n2838), .dout(n2847));
  jxor g02592(.dina(n2847), .dinb(n2747), .dout(n2848));
  jxor g02593(.dina(n2848), .dinb(n2743), .dout(n2849));
  jnot g02594(.din(n2849), .dout(n2850));
  jxor g02595(.dina(n2850), .dinb(n2734), .dout(n2851));
  jor  g02596(.dina(n2404), .dinb(n402), .dout(n2852));
  jor  g02597(.dina(n371), .dinb(n2010), .dout(n2853));
  jor  g02598(.dina(n405), .dinb(n2148), .dout(n2854));
  jor  g02599(.dina(n332), .dinb(n2407), .dout(n2855));
  jand g02600(.dina(n2855), .dinb(n2854), .dout(n2856));
  jand g02601(.dina(n2856), .dinb(n2853), .dout(n2857));
  jand g02602(.dina(n2857), .dinb(n2852), .dout(n2858));
  jxor g02603(.dina(n2858), .dinb(a5 ), .dout(n2859));
  jxor g02604(.dina(n2859), .dinb(n2851), .dout(n2860));
  jxor g02605(.dina(n2860), .dinb(n2729), .dout(n2861));
  jand g02606(.dina(b29 ), .dinb(b28 ), .dout(n2862));
  jand g02607(.dina(n2574), .dinb(n2573), .dout(n2863));
  jor  g02608(.dina(n2863), .dinb(n2862), .dout(n2864));
  jxor g02609(.dina(b30 ), .dinb(b29 ), .dout(n2865));
  jnot g02610(.din(n2865), .dout(n2866));
  jxor g02611(.dina(n2866), .dinb(n2864), .dout(n2867));
  jor  g02612(.dina(n2867), .dinb(n264), .dout(n2868));
  jor  g02613(.dina(n284), .dinb(n2559), .dout(n2869));
  jnot g02614(.din(b30 ), .dout(n2870));
  jor  g02615(.dina(n269), .dinb(n2870), .dout(n2871));
  jor  g02616(.dina(n271), .dinb(n2579), .dout(n2872));
  jand g02617(.dina(n2872), .dinb(n2871), .dout(n2873));
  jand g02618(.dina(n2873), .dinb(n2869), .dout(n2874));
  jand g02619(.dina(n2874), .dinb(n2868), .dout(n2875));
  jxor g02620(.dina(n2875), .dinb(n260), .dout(n2876));
  jxor g02621(.dina(n2876), .dinb(n2861), .dout(n2877));
  jxor g02622(.dina(n2877), .dinb(n2726), .dout(f30 ));
  jand g02623(.dina(n2876), .dinb(n2861), .dout(n2879));
  jand g02624(.dina(n2877), .dinb(n2726), .dout(n2880));
  jor  g02625(.dina(n2880), .dinb(n2879), .dout(n2881));
  jor  g02626(.dina(n2859), .dinb(n2851), .dout(n2882));
  jnot g02627(.din(n2882), .dout(n2883));
  jand g02628(.dina(n2860), .dinb(n2729), .dout(n2884));
  jor  g02629(.dina(n2884), .dinb(n2883), .dout(n2885));
  jand g02630(.dina(n2848), .dinb(n2743), .dout(n2886));
  jand g02631(.dina(n2849), .dinb(n2734), .dout(n2887));
  jor  g02632(.dina(n2887), .dinb(n2886), .dout(n2888));
  jnot g02633(.din(n2838), .dout(n2889));
  jor  g02634(.dina(n2846), .dinb(n2889), .dout(n2890));
  jor  g02635(.dina(n2847), .dinb(n2747), .dout(n2891));
  jand g02636(.dina(n2891), .dinb(n2890), .dout(n2892));
  jor  g02637(.dina(n2836), .dinb(n2828), .dout(n2893));
  jnot g02638(.din(n2893), .dout(n2894));
  jand g02639(.dina(n2837), .dinb(n2751), .dout(n2895));
  jor  g02640(.dina(n2895), .dinb(n2894), .dout(n2896));
  jor  g02641(.dina(n2825), .dinb(n2817), .dout(n2897));
  jand g02642(.dina(n2826), .dinb(n2756), .dout(n2898));
  jnot g02643(.din(n2898), .dout(n2899));
  jand g02644(.dina(n2899), .dinb(n2897), .dout(n2900));
  jnot g02645(.din(n2900), .dout(n2901));
  jand g02646(.dina(n2812), .dinb(n2780), .dout(n2902));
  jand g02647(.dina(n2813), .dinb(n2771), .dout(n2903));
  jor  g02648(.dina(n2903), .dinb(n2902), .dout(n2904));
  jor  g02649(.dina(n2810), .dinb(n2802), .dout(n2905));
  jand g02650(.dina(n2811), .dinb(n2783), .dout(n2906));
  jnot g02651(.din(n2906), .dout(n2907));
  jand g02652(.dina(n2907), .dinb(n2905), .dout(n2908));
  jnot g02653(.din(n2908), .dout(n2909));
  jor  g02654(.dina(n2319), .dinb(n428), .dout(n2910));
  jor  g02655(.dina(n2224), .dinb(n357), .dout(n2911));
  jor  g02656(.dina(n2322), .dinb(n395), .dout(n2912));
  jor  g02657(.dina(n2324), .dinb(n431), .dout(n2913));
  jand g02658(.dina(n2913), .dinb(n2912), .dout(n2914));
  jand g02659(.dina(n2914), .dinb(n2911), .dout(n2915));
  jand g02660(.dina(n2915), .dinb(n2910), .dout(n2916));
  jxor g02661(.dina(n2916), .dinb(a26 ), .dout(n2917));
  jnot g02662(.din(n2917), .dout(n2918));
  jnot g02663(.din(n2799), .dout(n2919));
  jand g02664(.dina(n2919), .dinb(n2797), .dout(n2920));
  jand g02665(.dina(n2800), .dinb(n2795), .dout(n2921));
  jor  g02666(.dina(n2921), .dinb(n2920), .dout(n2922));
  jor  g02667(.dina(n2784), .dinb(n319), .dout(n2923));
  jor  g02668(.dina(n2661), .dinb(n279), .dout(n2924));
  jor  g02669(.dina(n2787), .dinb(n299), .dout(n2925));
  jor  g02670(.dina(n2789), .dinb(n322), .dout(n2926));
  jand g02671(.dina(n2926), .dinb(n2925), .dout(n2927));
  jand g02672(.dina(n2927), .dinb(n2924), .dout(n2928));
  jand g02673(.dina(n2928), .dinb(n2923), .dout(n2929));
  jxor g02674(.dina(n2929), .dinb(a29 ), .dout(n2930));
  jnot g02675(.din(n2930), .dout(n2931));
  jand g02676(.dina(n2797), .dinb(a32 ), .dout(n2932));
  jxor g02677(.dina(a32 ), .dinb(a31 ), .dout(n2933));
  jnot g02678(.din(n2933), .dout(n2934));
  jand g02679(.dina(n2934), .dinb(n2796), .dout(n2935));
  jand g02680(.dina(n2935), .dinb(b1 ), .dout(n2936));
  jnot g02681(.din(n2796), .dout(n2937));
  jxor g02682(.dina(a31 ), .dinb(a30 ), .dout(n2938));
  jand g02683(.dina(n2938), .dinb(n2937), .dout(n2939));
  jand g02684(.dina(n2939), .dinb(b0 ), .dout(n2940));
  jand g02685(.dina(n2933), .dinb(n2796), .dout(n2941));
  jand g02686(.dina(n2941), .dinb(n338), .dout(n2942));
  jor  g02687(.dina(n2942), .dinb(n2940), .dout(n2943));
  jor  g02688(.dina(n2943), .dinb(n2936), .dout(n2944));
  jxor g02689(.dina(n2944), .dinb(n2932), .dout(n2945));
  jxor g02690(.dina(n2945), .dinb(n2931), .dout(n2946));
  jxor g02691(.dina(n2946), .dinb(n2922), .dout(n2947));
  jxor g02692(.dina(n2947), .dinb(n2918), .dout(n2948));
  jxor g02693(.dina(n2948), .dinb(n2909), .dout(n2949));
  jnot g02694(.din(n2949), .dout(n2950));
  jor  g02695(.dina(n1939), .dinb(n624), .dout(n2951));
  jor  g02696(.dina(n1827), .dinb(n512), .dout(n2952));
  jor  g02697(.dina(n1942), .dinb(n564), .dout(n2953));
  jor  g02698(.dina(n1944), .dinb(n627), .dout(n2954));
  jand g02699(.dina(n2954), .dinb(n2953), .dout(n2955));
  jand g02700(.dina(n2955), .dinb(n2952), .dout(n2956));
  jand g02701(.dina(n2956), .dinb(n2951), .dout(n2957));
  jxor g02702(.dina(n2957), .dinb(a23 ), .dout(n2958));
  jxor g02703(.dina(n2958), .dinb(n2950), .dout(n2959));
  jxor g02704(.dina(n2959), .dinb(n2904), .dout(n2960));
  jnot g02705(.din(n2960), .dout(n2961));
  jor  g02706(.dina(n1566), .dinb(n775), .dout(n2962));
  jor  g02707(.dina(n1489), .dinb(n647), .dout(n2963));
  jor  g02708(.dina(n1569), .dinb(n758), .dout(n2964));
  jor  g02709(.dina(n1571), .dinb(n778), .dout(n2965));
  jand g02710(.dina(n2965), .dinb(n2964), .dout(n2966));
  jand g02711(.dina(n2966), .dinb(n2963), .dout(n2967));
  jand g02712(.dina(n2967), .dinb(n2962), .dout(n2968));
  jxor g02713(.dina(n2968), .dinb(a20 ), .dout(n2969));
  jxor g02714(.dina(n2969), .dinb(n2961), .dout(n2970));
  jand g02715(.dina(n2814), .dinb(n2768), .dout(n2971));
  jand g02716(.dina(n2815), .dinb(n2759), .dout(n2972));
  jor  g02717(.dina(n2972), .dinb(n2971), .dout(n2973));
  jxor g02718(.dina(n2973), .dinb(n2970), .dout(n2974));
  jnot g02719(.din(n2974), .dout(n2975));
  jor  g02720(.dina(n1245), .dinb(n1019), .dout(n2976));
  jor  g02721(.dina(n1165), .dinb(n858), .dout(n2977));
  jor  g02722(.dina(n1248), .dinb(n939), .dout(n2978));
  jor  g02723(.dina(n1250), .dinb(n1022), .dout(n2979));
  jand g02724(.dina(n2979), .dinb(n2978), .dout(n2980));
  jand g02725(.dina(n2980), .dinb(n2977), .dout(n2981));
  jand g02726(.dina(n2981), .dinb(n2976), .dout(n2982));
  jxor g02727(.dina(n2982), .dinb(a17 ), .dout(n2983));
  jxor g02728(.dina(n2983), .dinb(n2975), .dout(n2984));
  jxor g02729(.dina(n2984), .dinb(n2901), .dout(n2985));
  jnot g02730(.din(n2985), .dout(n2986));
  jor  g02731(.dina(n1397), .dinb(n974), .dout(n2987));
  jor  g02732(.dina(n908), .dinb(n1193), .dout(n2988));
  jor  g02733(.dina(n977), .dinb(n1290), .dout(n2989));
  jor  g02734(.dina(n979), .dinb(n1400), .dout(n2990));
  jand g02735(.dina(n2990), .dinb(n2989), .dout(n2991));
  jand g02736(.dina(n2991), .dinb(n2988), .dout(n2992));
  jand g02737(.dina(n2992), .dinb(n2987), .dout(n2993));
  jxor g02738(.dina(n2993), .dinb(a14 ), .dout(n2994));
  jxor g02739(.dina(n2994), .dinb(n2986), .dout(n2995));
  jxor g02740(.dina(n2995), .dinb(n2896), .dout(n2996));
  jor  g02741(.dina(n1739), .dinb(n706), .dout(n2997));
  jor  g02742(.dina(n683), .dinb(n1420), .dout(n2998));
  jor  g02743(.dina(n709), .dinb(n1620), .dout(n2999));
  jor  g02744(.dina(n711), .dinb(n1742), .dout(n3000));
  jand g02745(.dina(n3000), .dinb(n2999), .dout(n3001));
  jand g02746(.dina(n3001), .dinb(n2998), .dout(n3002));
  jand g02747(.dina(n3002), .dinb(n2997), .dout(n3003));
  jxor g02748(.dina(n3003), .dinb(a11 ), .dout(n3004));
  jxor g02749(.dina(n3004), .dinb(n2996), .dout(n3005));
  jxor g02750(.dina(n3005), .dinb(n2892), .dout(n3006));
  jor  g02751(.dina(n2007), .dinb(n528), .dout(n3007));
  jor  g02752(.dina(n490), .dinb(n1867), .dout(n3008));
  jor  g02753(.dina(n531), .dinb(n1887), .dout(n3009));
  jor  g02754(.dina(n533), .dinb(n2010), .dout(n3010));
  jand g02755(.dina(n3010), .dinb(n3009), .dout(n3011));
  jand g02756(.dina(n3011), .dinb(n3008), .dout(n3012));
  jand g02757(.dina(n3012), .dinb(n3007), .dout(n3013));
  jxor g02758(.dina(n3013), .dinb(a8 ), .dout(n3014));
  jxor g02759(.dina(n3014), .dinb(n3006), .dout(n3015));
  jxor g02760(.dina(n3015), .dinb(n2888), .dout(n3016));
  jor  g02761(.dina(n2556), .dinb(n402), .dout(n3017));
  jor  g02762(.dina(n371), .dinb(n2148), .dout(n3018));
  jor  g02763(.dina(n405), .dinb(n2407), .dout(n3019));
  jor  g02764(.dina(n332), .dinb(n2559), .dout(n3020));
  jand g02765(.dina(n3020), .dinb(n3019), .dout(n3021));
  jand g02766(.dina(n3021), .dinb(n3018), .dout(n3022));
  jand g02767(.dina(n3022), .dinb(n3017), .dout(n3023));
  jxor g02768(.dina(n3023), .dinb(a5 ), .dout(n3024));
  jxor g02769(.dina(n3024), .dinb(n3016), .dout(n3025));
  jxor g02770(.dina(n3025), .dinb(n2885), .dout(n3026));
  jand g02771(.dina(b30 ), .dinb(b29 ), .dout(n3027));
  jand g02772(.dina(n2865), .dinb(n2864), .dout(n3028));
  jor  g02773(.dina(n3028), .dinb(n3027), .dout(n3029));
  jxor g02774(.dina(b31 ), .dinb(b30 ), .dout(n3030));
  jnot g02775(.din(n3030), .dout(n3031));
  jxor g02776(.dina(n3031), .dinb(n3029), .dout(n3032));
  jor  g02777(.dina(n3032), .dinb(n264), .dout(n3033));
  jor  g02778(.dina(n284), .dinb(n2579), .dout(n3034));
  jnot g02779(.din(b31 ), .dout(n3035));
  jor  g02780(.dina(n269), .dinb(n3035), .dout(n3036));
  jor  g02781(.dina(n271), .dinb(n2870), .dout(n3037));
  jand g02782(.dina(n3037), .dinb(n3036), .dout(n3038));
  jand g02783(.dina(n3038), .dinb(n3034), .dout(n3039));
  jand g02784(.dina(n3039), .dinb(n3033), .dout(n3040));
  jxor g02785(.dina(n3040), .dinb(n260), .dout(n3041));
  jxor g02786(.dina(n3041), .dinb(n3026), .dout(n3042));
  jxor g02787(.dina(n3042), .dinb(n2881), .dout(f31 ));
  jand g02788(.dina(n3041), .dinb(n3026), .dout(n3044));
  jand g02789(.dina(n3042), .dinb(n2881), .dout(n3045));
  jor  g02790(.dina(n3045), .dinb(n3044), .dout(n3046));
  jand g02791(.dina(b31 ), .dinb(b30 ), .dout(n3047));
  jand g02792(.dina(n3030), .dinb(n3029), .dout(n3048));
  jor  g02793(.dina(n3048), .dinb(n3047), .dout(n3049));
  jxor g02794(.dina(b32 ), .dinb(b31 ), .dout(n3050));
  jnot g02795(.din(n3050), .dout(n3051));
  jxor g02796(.dina(n3051), .dinb(n3049), .dout(n3052));
  jor  g02797(.dina(n3052), .dinb(n264), .dout(n3053));
  jor  g02798(.dina(n284), .dinb(n2870), .dout(n3054));
  jnot g02799(.din(b32 ), .dout(n3055));
  jor  g02800(.dina(n269), .dinb(n3055), .dout(n3056));
  jor  g02801(.dina(n271), .dinb(n3035), .dout(n3057));
  jand g02802(.dina(n3057), .dinb(n3056), .dout(n3058));
  jand g02803(.dina(n3058), .dinb(n3054), .dout(n3059));
  jand g02804(.dina(n3059), .dinb(n3053), .dout(n3060));
  jxor g02805(.dina(n3060), .dinb(n260), .dout(n3061));
  jor  g02806(.dina(n3024), .dinb(n3016), .dout(n3062));
  jnot g02807(.din(n3062), .dout(n3063));
  jand g02808(.dina(n3025), .dinb(n2885), .dout(n3064));
  jor  g02809(.dina(n3064), .dinb(n3063), .dout(n3065));
  jnot g02810(.din(n3006), .dout(n3066));
  jor  g02811(.dina(n3014), .dinb(n3066), .dout(n3067));
  jnot g02812(.din(n3067), .dout(n3068));
  jnot g02813(.din(n3015), .dout(n3069));
  jand g02814(.dina(n3069), .dinb(n2888), .dout(n3070));
  jor  g02815(.dina(n3070), .dinb(n3068), .dout(n3071));
  jnot g02816(.din(n3071), .dout(n3072));
  jnot g02817(.din(n2996), .dout(n3073));
  jor  g02818(.dina(n3004), .dinb(n3073), .dout(n3074));
  jor  g02819(.dina(n3005), .dinb(n2892), .dout(n3075));
  jand g02820(.dina(n3075), .dinb(n3074), .dout(n3076));
  jnot g02821(.din(n3076), .dout(n3077));
  jor  g02822(.dina(n1864), .dinb(n706), .dout(n3078));
  jor  g02823(.dina(n683), .dinb(n1620), .dout(n3079));
  jor  g02824(.dina(n709), .dinb(n1742), .dout(n3080));
  jor  g02825(.dina(n711), .dinb(n1867), .dout(n3081));
  jand g02826(.dina(n3081), .dinb(n3080), .dout(n3082));
  jand g02827(.dina(n3082), .dinb(n3079), .dout(n3083));
  jand g02828(.dina(n3083), .dinb(n3078), .dout(n3084));
  jxor g02829(.dina(n3084), .dinb(a11 ), .dout(n3085));
  jnot g02830(.din(n3085), .dout(n3086));
  jor  g02831(.dina(n2994), .dinb(n2986), .dout(n3087));
  jnot g02832(.din(n3087), .dout(n3088));
  jand g02833(.dina(n2995), .dinb(n2896), .dout(n3089));
  jor  g02834(.dina(n3089), .dinb(n3088), .dout(n3090));
  jor  g02835(.dina(n2983), .dinb(n2975), .dout(n3091));
  jand g02836(.dina(n2984), .dinb(n2901), .dout(n3092));
  jnot g02837(.din(n3092), .dout(n3093));
  jand g02838(.dina(n3093), .dinb(n3091), .dout(n3094));
  jnot g02839(.din(n3094), .dout(n3095));
  jor  g02840(.dina(n2969), .dinb(n2961), .dout(n3096));
  jand g02841(.dina(n2973), .dinb(n2970), .dout(n3097));
  jnot g02842(.din(n3097), .dout(n3098));
  jand g02843(.dina(n3098), .dinb(n3096), .dout(n3099));
  jnot g02844(.din(n3099), .dout(n3100));
  jor  g02845(.dina(n1566), .dinb(n855), .dout(n3101));
  jor  g02846(.dina(n1489), .dinb(n758), .dout(n3102));
  jor  g02847(.dina(n1569), .dinb(n778), .dout(n3103));
  jor  g02848(.dina(n1571), .dinb(n858), .dout(n3104));
  jand g02849(.dina(n3104), .dinb(n3103), .dout(n3105));
  jand g02850(.dina(n3105), .dinb(n3102), .dout(n3106));
  jand g02851(.dina(n3106), .dinb(n3101), .dout(n3107));
  jxor g02852(.dina(n3107), .dinb(a20 ), .dout(n3108));
  jnot g02853(.din(n3108), .dout(n3109));
  jor  g02854(.dina(n2958), .dinb(n2950), .dout(n3110));
  jand g02855(.dina(n2959), .dinb(n2904), .dout(n3111));
  jnot g02856(.din(n3111), .dout(n3112));
  jand g02857(.dina(n3112), .dinb(n3110), .dout(n3113));
  jnot g02858(.din(n3113), .dout(n3114));
  jand g02859(.dina(n2947), .dinb(n2918), .dout(n3115));
  jand g02860(.dina(n2948), .dinb(n2909), .dout(n3116));
  jor  g02861(.dina(n3116), .dinb(n3115), .dout(n3117));
  jand g02862(.dina(n2945), .dinb(n2931), .dout(n3118));
  jand g02863(.dina(n2946), .dinb(n2922), .dout(n3119));
  jor  g02864(.dina(n3119), .dinb(n3118), .dout(n3120));
  jor  g02865(.dina(n2784), .dinb(n354), .dout(n3121));
  jor  g02866(.dina(n2661), .dinb(n299), .dout(n3122));
  jor  g02867(.dina(n2787), .dinb(n322), .dout(n3123));
  jor  g02868(.dina(n2789), .dinb(n357), .dout(n3124));
  jand g02869(.dina(n3124), .dinb(n3123), .dout(n3125));
  jand g02870(.dina(n3125), .dinb(n3122), .dout(n3126));
  jand g02871(.dina(n3126), .dinb(n3121), .dout(n3127));
  jxor g02872(.dina(n3127), .dinb(a29 ), .dout(n3128));
  jnot g02873(.din(n3128), .dout(n3129));
  jnot g02874(.din(n2944), .dout(n3130));
  jand g02875(.dina(n2798), .dinb(a32 ), .dout(n3131));
  jand g02876(.dina(n3131), .dinb(n3130), .dout(n3132));
  jnot g02877(.din(n3132), .dout(n3133));
  jand g02878(.dina(n3133), .dinb(a32 ), .dout(n3134));
  jor  g02879(.dina(n2938), .dinb(n2934), .dout(n3135));
  jor  g02880(.dina(n3135), .dinb(n2796), .dout(n3136));
  jnot g02881(.din(n3136), .dout(n3137));
  jand g02882(.dina(n3137), .dinb(b0 ), .dout(n3138));
  jand g02883(.dina(n2935), .dinb(b2 ), .dout(n3139));
  jand g02884(.dina(n2939), .dinb(b1 ), .dout(n3140));
  jand g02885(.dina(n2941), .dinb(n375), .dout(n3141));
  jor  g02886(.dina(n3141), .dinb(n3140), .dout(n3142));
  jor  g02887(.dina(n3142), .dinb(n3139), .dout(n3143));
  jor  g02888(.dina(n3143), .dinb(n3138), .dout(n3144));
  jxor g02889(.dina(n3144), .dinb(n3134), .dout(n3145));
  jxor g02890(.dina(n3145), .dinb(n3129), .dout(n3146));
  jxor g02891(.dina(n3146), .dinb(n3120), .dout(n3147));
  jnot g02892(.din(n3147), .dout(n3148));
  jor  g02893(.dina(n2319), .dinb(n509), .dout(n3149));
  jor  g02894(.dina(n2224), .dinb(n395), .dout(n3150));
  jor  g02895(.dina(n2322), .dinb(n431), .dout(n3151));
  jor  g02896(.dina(n2324), .dinb(n512), .dout(n3152));
  jand g02897(.dina(n3152), .dinb(n3151), .dout(n3153));
  jand g02898(.dina(n3153), .dinb(n3150), .dout(n3154));
  jand g02899(.dina(n3154), .dinb(n3149), .dout(n3155));
  jxor g02900(.dina(n3155), .dinb(a26 ), .dout(n3156));
  jxor g02901(.dina(n3156), .dinb(n3148), .dout(n3157));
  jxor g02902(.dina(n3157), .dinb(n3117), .dout(n3158));
  jnot g02903(.din(n3158), .dout(n3159));
  jor  g02904(.dina(n1939), .dinb(n644), .dout(n3160));
  jor  g02905(.dina(n1827), .dinb(n564), .dout(n3161));
  jor  g02906(.dina(n1942), .dinb(n627), .dout(n3162));
  jor  g02907(.dina(n1944), .dinb(n647), .dout(n3163));
  jand g02908(.dina(n3163), .dinb(n3162), .dout(n3164));
  jand g02909(.dina(n3164), .dinb(n3161), .dout(n3165));
  jand g02910(.dina(n3165), .dinb(n3160), .dout(n3166));
  jxor g02911(.dina(n3166), .dinb(a23 ), .dout(n3167));
  jxor g02912(.dina(n3167), .dinb(n3159), .dout(n3168));
  jxor g02913(.dina(n3168), .dinb(n3114), .dout(n3169));
  jxor g02914(.dina(n3169), .dinb(n3109), .dout(n3170));
  jxor g02915(.dina(n3170), .dinb(n3100), .dout(n3171));
  jnot g02916(.din(n3171), .dout(n3172));
  jor  g02917(.dina(n1190), .dinb(n1245), .dout(n3173));
  jor  g02918(.dina(n1165), .dinb(n939), .dout(n3174));
  jor  g02919(.dina(n1248), .dinb(n1022), .dout(n3175));
  jor  g02920(.dina(n1250), .dinb(n1193), .dout(n3176));
  jand g02921(.dina(n3176), .dinb(n3175), .dout(n3177));
  jand g02922(.dina(n3177), .dinb(n3174), .dout(n3178));
  jand g02923(.dina(n3178), .dinb(n3173), .dout(n3179));
  jxor g02924(.dina(n3179), .dinb(a17 ), .dout(n3180));
  jxor g02925(.dina(n3180), .dinb(n3172), .dout(n3181));
  jxor g02926(.dina(n3181), .dinb(n3095), .dout(n3182));
  jor  g02927(.dina(n1417), .dinb(n974), .dout(n3183));
  jor  g02928(.dina(n908), .dinb(n1290), .dout(n3184));
  jor  g02929(.dina(n977), .dinb(n1400), .dout(n3185));
  jor  g02930(.dina(n979), .dinb(n1420), .dout(n3186));
  jand g02931(.dina(n3186), .dinb(n3185), .dout(n3187));
  jand g02932(.dina(n3187), .dinb(n3184), .dout(n3188));
  jand g02933(.dina(n3188), .dinb(n3183), .dout(n3189));
  jxor g02934(.dina(n3189), .dinb(a14 ), .dout(n3190));
  jxor g02935(.dina(n3190), .dinb(n3182), .dout(n3191));
  jnot g02936(.din(n3191), .dout(n3192));
  jxor g02937(.dina(n3192), .dinb(n3090), .dout(n3193));
  jxor g02938(.dina(n3193), .dinb(n3086), .dout(n3194));
  jxor g02939(.dina(n3194), .dinb(n3077), .dout(n3195));
  jnot g02940(.din(n3195), .dout(n3196));
  jor  g02941(.dina(n2145), .dinb(n528), .dout(n3197));
  jor  g02942(.dina(n490), .dinb(n1887), .dout(n3198));
  jor  g02943(.dina(n531), .dinb(n2010), .dout(n3199));
  jor  g02944(.dina(n533), .dinb(n2148), .dout(n3200));
  jand g02945(.dina(n3200), .dinb(n3199), .dout(n3201));
  jand g02946(.dina(n3201), .dinb(n3198), .dout(n3202));
  jand g02947(.dina(n3202), .dinb(n3197), .dout(n3203));
  jxor g02948(.dina(n3203), .dinb(a8 ), .dout(n3204));
  jxor g02949(.dina(n3204), .dinb(n3196), .dout(n3205));
  jxor g02950(.dina(n3205), .dinb(n3072), .dout(n3206));
  jor  g02951(.dina(n2576), .dinb(n402), .dout(n3207));
  jor  g02952(.dina(n371), .dinb(n2407), .dout(n3208));
  jor  g02953(.dina(n405), .dinb(n2559), .dout(n3209));
  jor  g02954(.dina(n332), .dinb(n2579), .dout(n3210));
  jand g02955(.dina(n3210), .dinb(n3209), .dout(n3211));
  jand g02956(.dina(n3211), .dinb(n3208), .dout(n3212));
  jand g02957(.dina(n3212), .dinb(n3207), .dout(n3213));
  jxor g02958(.dina(n3213), .dinb(a5 ), .dout(n3214));
  jxor g02959(.dina(n3214), .dinb(n3206), .dout(n3215));
  jxor g02960(.dina(n3215), .dinb(n3065), .dout(n3216));
  jxor g02961(.dina(n3216), .dinb(n3061), .dout(n3217));
  jxor g02962(.dina(n3217), .dinb(n3046), .dout(f32 ));
  jand g02963(.dina(n3216), .dinb(n3061), .dout(n3219));
  jand g02964(.dina(n3217), .dinb(n3046), .dout(n3220));
  jor  g02965(.dina(n3220), .dinb(n3219), .dout(n3221));
  jand g02966(.dina(b32 ), .dinb(b31 ), .dout(n3222));
  jand g02967(.dina(n3050), .dinb(n3049), .dout(n3223));
  jor  g02968(.dina(n3223), .dinb(n3222), .dout(n3224));
  jxor g02969(.dina(b33 ), .dinb(b32 ), .dout(n3225));
  jnot g02970(.din(n3225), .dout(n3226));
  jxor g02971(.dina(n3226), .dinb(n3224), .dout(n3227));
  jor  g02972(.dina(n3227), .dinb(n264), .dout(n3228));
  jor  g02973(.dina(n284), .dinb(n3035), .dout(n3229));
  jnot g02974(.din(b33 ), .dout(n3230));
  jor  g02975(.dina(n269), .dinb(n3230), .dout(n3231));
  jor  g02976(.dina(n271), .dinb(n3055), .dout(n3232));
  jand g02977(.dina(n3232), .dinb(n3231), .dout(n3233));
  jand g02978(.dina(n3233), .dinb(n3229), .dout(n3234));
  jand g02979(.dina(n3234), .dinb(n3228), .dout(n3235));
  jxor g02980(.dina(n3235), .dinb(n260), .dout(n3236));
  jor  g02981(.dina(n3214), .dinb(n3206), .dout(n3237));
  jnot g02982(.din(n3237), .dout(n3238));
  jand g02983(.dina(n3215), .dinb(n3065), .dout(n3239));
  jor  g02984(.dina(n3239), .dinb(n3238), .dout(n3240));
  jor  g02985(.dina(n3204), .dinb(n3196), .dout(n3241));
  jnot g02986(.din(n3241), .dout(n3242));
  jand g02987(.dina(n3205), .dinb(n3071), .dout(n3243));
  jor  g02988(.dina(n3243), .dinb(n3242), .dout(n3244));
  jnot g02989(.din(n3244), .dout(n3245));
  jand g02990(.dina(n3193), .dinb(n3086), .dout(n3246));
  jand g02991(.dina(n3194), .dinb(n3077), .dout(n3247));
  jor  g02992(.dina(n3247), .dinb(n3246), .dout(n3248));
  jor  g02993(.dina(n1884), .dinb(n706), .dout(n3249));
  jor  g02994(.dina(n683), .dinb(n1742), .dout(n3250));
  jor  g02995(.dina(n709), .dinb(n1867), .dout(n3251));
  jor  g02996(.dina(n711), .dinb(n1887), .dout(n3252));
  jand g02997(.dina(n3252), .dinb(n3251), .dout(n3253));
  jand g02998(.dina(n3253), .dinb(n3250), .dout(n3254));
  jand g02999(.dina(n3254), .dinb(n3249), .dout(n3255));
  jxor g03000(.dina(n3255), .dinb(a11 ), .dout(n3256));
  jnot g03001(.din(n3256), .dout(n3257));
  jnot g03002(.din(n3182), .dout(n3258));
  jor  g03003(.dina(n3190), .dinb(n3258), .dout(n3259));
  jnot g03004(.din(n3259), .dout(n3260));
  jand g03005(.dina(n3192), .dinb(n3090), .dout(n3261));
  jor  g03006(.dina(n3261), .dinb(n3260), .dout(n3262));
  jor  g03007(.dina(n3180), .dinb(n3172), .dout(n3263));
  jnot g03008(.din(n3263), .dout(n3264));
  jand g03009(.dina(n3181), .dinb(n3095), .dout(n3265));
  jor  g03010(.dina(n3265), .dinb(n3264), .dout(n3266));
  jor  g03011(.dina(n1287), .dinb(n1245), .dout(n3267));
  jor  g03012(.dina(n1165), .dinb(n1022), .dout(n3268));
  jor  g03013(.dina(n1248), .dinb(n1193), .dout(n3269));
  jor  g03014(.dina(n1250), .dinb(n1290), .dout(n3270));
  jand g03015(.dina(n3270), .dinb(n3269), .dout(n3271));
  jand g03016(.dina(n3271), .dinb(n3268), .dout(n3272));
  jand g03017(.dina(n3272), .dinb(n3267), .dout(n3273));
  jxor g03018(.dina(n3273), .dinb(a17 ), .dout(n3274));
  jnot g03019(.din(n3274), .dout(n3275));
  jand g03020(.dina(n3169), .dinb(n3109), .dout(n3276));
  jand g03021(.dina(n3170), .dinb(n3100), .dout(n3277));
  jor  g03022(.dina(n3277), .dinb(n3276), .dout(n3278));
  jor  g03023(.dina(n3167), .dinb(n3159), .dout(n3279));
  jand g03024(.dina(n3168), .dinb(n3114), .dout(n3280));
  jnot g03025(.din(n3280), .dout(n3281));
  jand g03026(.dina(n3281), .dinb(n3279), .dout(n3282));
  jnot g03027(.din(n3282), .dout(n3283));
  jor  g03028(.dina(n3156), .dinb(n3148), .dout(n3284));
  jand g03029(.dina(n3157), .dinb(n3117), .dout(n3285));
  jnot g03030(.din(n3285), .dout(n3286));
  jand g03031(.dina(n3286), .dinb(n3284), .dout(n3287));
  jnot g03032(.din(n3287), .dout(n3288));
  jor  g03033(.dina(n2319), .dinb(n561), .dout(n3289));
  jor  g03034(.dina(n2224), .dinb(n431), .dout(n3290));
  jor  g03035(.dina(n2322), .dinb(n512), .dout(n3291));
  jor  g03036(.dina(n2324), .dinb(n564), .dout(n3292));
  jand g03037(.dina(n3292), .dinb(n3291), .dout(n3293));
  jand g03038(.dina(n3293), .dinb(n3290), .dout(n3294));
  jand g03039(.dina(n3294), .dinb(n3289), .dout(n3295));
  jxor g03040(.dina(n3295), .dinb(a26 ), .dout(n3296));
  jnot g03041(.din(n3296), .dout(n3297));
  jand g03042(.dina(n3145), .dinb(n3129), .dout(n3298));
  jand g03043(.dina(n3146), .dinb(n3120), .dout(n3299));
  jor  g03044(.dina(n3299), .dinb(n3298), .dout(n3300));
  jnot g03045(.din(n2941), .dout(n3301));
  jor  g03046(.dina(n3301), .dinb(n296), .dout(n3302));
  jor  g03047(.dina(n3136), .dinb(n267), .dout(n3303));
  jnot g03048(.din(n2939), .dout(n3304));
  jor  g03049(.dina(n3304), .dinb(n279), .dout(n3305));
  jnot g03050(.din(n2935), .dout(n3306));
  jor  g03051(.dina(n3306), .dinb(n299), .dout(n3307));
  jand g03052(.dina(n3307), .dinb(n3305), .dout(n3308));
  jand g03053(.dina(n3308), .dinb(n3303), .dout(n3309));
  jand g03054(.dina(n3309), .dinb(n3302), .dout(n3310));
  jxor g03055(.dina(n3310), .dinb(a32 ), .dout(n3311));
  jnot g03056(.din(n3311), .dout(n3312));
  jxor g03057(.dina(a33 ), .dinb(a32 ), .dout(n3313));
  jand g03058(.dina(n3313), .dinb(b0 ), .dout(n3314));
  jnot g03059(.din(n3314), .dout(n3315));
  jor  g03060(.dina(n3144), .dinb(n3133), .dout(n3316));
  jxor g03061(.dina(n3316), .dinb(n3315), .dout(n3317));
  jxor g03062(.dina(n3317), .dinb(n3312), .dout(n3318));
  jnot g03063(.din(n3318), .dout(n3319));
  jor  g03064(.dina(n2784), .dinb(n392), .dout(n3320));
  jor  g03065(.dina(n2661), .dinb(n322), .dout(n3321));
  jor  g03066(.dina(n2787), .dinb(n357), .dout(n3322));
  jor  g03067(.dina(n2789), .dinb(n395), .dout(n3323));
  jand g03068(.dina(n3323), .dinb(n3322), .dout(n3324));
  jand g03069(.dina(n3324), .dinb(n3321), .dout(n3325));
  jand g03070(.dina(n3325), .dinb(n3320), .dout(n3326));
  jxor g03071(.dina(n3326), .dinb(a29 ), .dout(n3327));
  jxor g03072(.dina(n3327), .dinb(n3319), .dout(n3328));
  jxor g03073(.dina(n3328), .dinb(n3300), .dout(n3329));
  jxor g03074(.dina(n3329), .dinb(n3297), .dout(n3330));
  jxor g03075(.dina(n3330), .dinb(n3288), .dout(n3331));
  jnot g03076(.din(n3331), .dout(n3332));
  jor  g03077(.dina(n1939), .dinb(n755), .dout(n3333));
  jor  g03078(.dina(n1827), .dinb(n627), .dout(n3334));
  jor  g03079(.dina(n1942), .dinb(n647), .dout(n3335));
  jor  g03080(.dina(n1944), .dinb(n758), .dout(n3336));
  jand g03081(.dina(n3336), .dinb(n3335), .dout(n3337));
  jand g03082(.dina(n3337), .dinb(n3334), .dout(n3338));
  jand g03083(.dina(n3338), .dinb(n3333), .dout(n3339));
  jxor g03084(.dina(n3339), .dinb(a23 ), .dout(n3340));
  jxor g03085(.dina(n3340), .dinb(n3332), .dout(n3341));
  jxor g03086(.dina(n3341), .dinb(n3283), .dout(n3342));
  jnot g03087(.din(n3342), .dout(n3343));
  jor  g03088(.dina(n1566), .dinb(n936), .dout(n3344));
  jor  g03089(.dina(n1489), .dinb(n778), .dout(n3345));
  jor  g03090(.dina(n1569), .dinb(n858), .dout(n3346));
  jor  g03091(.dina(n1571), .dinb(n939), .dout(n3347));
  jand g03092(.dina(n3347), .dinb(n3346), .dout(n3348));
  jand g03093(.dina(n3348), .dinb(n3345), .dout(n3349));
  jand g03094(.dina(n3349), .dinb(n3344), .dout(n3350));
  jxor g03095(.dina(n3350), .dinb(a20 ), .dout(n3351));
  jxor g03096(.dina(n3351), .dinb(n3343), .dout(n3352));
  jxor g03097(.dina(n3352), .dinb(n3278), .dout(n3353));
  jxor g03098(.dina(n3353), .dinb(n3275), .dout(n3354));
  jxor g03099(.dina(n3354), .dinb(n3266), .dout(n3355));
  jor  g03100(.dina(n1617), .dinb(n974), .dout(n3356));
  jor  g03101(.dina(n908), .dinb(n1400), .dout(n3357));
  jor  g03102(.dina(n977), .dinb(n1420), .dout(n3358));
  jor  g03103(.dina(n979), .dinb(n1620), .dout(n3359));
  jand g03104(.dina(n3359), .dinb(n3358), .dout(n3360));
  jand g03105(.dina(n3360), .dinb(n3357), .dout(n3361));
  jand g03106(.dina(n3361), .dinb(n3356), .dout(n3362));
  jxor g03107(.dina(n3362), .dinb(a14 ), .dout(n3363));
  jxor g03108(.dina(n3363), .dinb(n3355), .dout(n3364));
  jnot g03109(.din(n3364), .dout(n3365));
  jxor g03110(.dina(n3365), .dinb(n3262), .dout(n3366));
  jxor g03111(.dina(n3366), .dinb(n3257), .dout(n3367));
  jxor g03112(.dina(n3367), .dinb(n3248), .dout(n3368));
  jnot g03113(.din(n3368), .dout(n3369));
  jor  g03114(.dina(n2404), .dinb(n528), .dout(n3370));
  jor  g03115(.dina(n490), .dinb(n2010), .dout(n3371));
  jor  g03116(.dina(n531), .dinb(n2148), .dout(n3372));
  jor  g03117(.dina(n533), .dinb(n2407), .dout(n3373));
  jand g03118(.dina(n3373), .dinb(n3372), .dout(n3374));
  jand g03119(.dina(n3374), .dinb(n3371), .dout(n3375));
  jand g03120(.dina(n3375), .dinb(n3370), .dout(n3376));
  jxor g03121(.dina(n3376), .dinb(a8 ), .dout(n3377));
  jxor g03122(.dina(n3377), .dinb(n3369), .dout(n3378));
  jxor g03123(.dina(n3378), .dinb(n3245), .dout(n3379));
  jor  g03124(.dina(n2867), .dinb(n402), .dout(n3380));
  jor  g03125(.dina(n371), .dinb(n2559), .dout(n3381));
  jor  g03126(.dina(n405), .dinb(n2579), .dout(n3382));
  jor  g03127(.dina(n332), .dinb(n2870), .dout(n3383));
  jand g03128(.dina(n3383), .dinb(n3382), .dout(n3384));
  jand g03129(.dina(n3384), .dinb(n3381), .dout(n3385));
  jand g03130(.dina(n3385), .dinb(n3380), .dout(n3386));
  jxor g03131(.dina(n3386), .dinb(a5 ), .dout(n3387));
  jxor g03132(.dina(n3387), .dinb(n3379), .dout(n3388));
  jxor g03133(.dina(n3388), .dinb(n3240), .dout(n3389));
  jxor g03134(.dina(n3389), .dinb(n3236), .dout(n3390));
  jxor g03135(.dina(n3390), .dinb(n3221), .dout(f33 ));
  jand g03136(.dina(n3389), .dinb(n3236), .dout(n3392));
  jand g03137(.dina(n3390), .dinb(n3221), .dout(n3393));
  jor  g03138(.dina(n3393), .dinb(n3392), .dout(n3394));
  jand g03139(.dina(b33 ), .dinb(b32 ), .dout(n3395));
  jand g03140(.dina(n3225), .dinb(n3224), .dout(n3396));
  jor  g03141(.dina(n3396), .dinb(n3395), .dout(n3397));
  jxor g03142(.dina(b34 ), .dinb(b33 ), .dout(n3398));
  jnot g03143(.din(n3398), .dout(n3399));
  jxor g03144(.dina(n3399), .dinb(n3397), .dout(n3400));
  jor  g03145(.dina(n3400), .dinb(n264), .dout(n3401));
  jor  g03146(.dina(n284), .dinb(n3055), .dout(n3402));
  jnot g03147(.din(b34 ), .dout(n3403));
  jor  g03148(.dina(n269), .dinb(n3403), .dout(n3404));
  jor  g03149(.dina(n271), .dinb(n3230), .dout(n3405));
  jand g03150(.dina(n3405), .dinb(n3404), .dout(n3406));
  jand g03151(.dina(n3406), .dinb(n3402), .dout(n3407));
  jand g03152(.dina(n3407), .dinb(n3401), .dout(n3408));
  jxor g03153(.dina(n3408), .dinb(n260), .dout(n3409));
  jor  g03154(.dina(n3387), .dinb(n3379), .dout(n3410));
  jnot g03155(.din(n3410), .dout(n3411));
  jand g03156(.dina(n3388), .dinb(n3240), .dout(n3412));
  jor  g03157(.dina(n3412), .dinb(n3411), .dout(n3413));
  jor  g03158(.dina(n3377), .dinb(n3369), .dout(n3414));
  jnot g03159(.din(n3414), .dout(n3415));
  jand g03160(.dina(n3378), .dinb(n3244), .dout(n3416));
  jor  g03161(.dina(n3416), .dinb(n3415), .dout(n3417));
  jnot g03162(.din(n3417), .dout(n3418));
  jand g03163(.dina(n3366), .dinb(n3257), .dout(n3419));
  jand g03164(.dina(n3367), .dinb(n3248), .dout(n3420));
  jor  g03165(.dina(n3420), .dinb(n3419), .dout(n3421));
  jnot g03166(.din(n3421), .dout(n3422));
  jnot g03167(.din(n3355), .dout(n3423));
  jor  g03168(.dina(n3363), .dinb(n3423), .dout(n3424));
  jnot g03169(.din(n3424), .dout(n3425));
  jand g03170(.dina(n3365), .dinb(n3262), .dout(n3426));
  jor  g03171(.dina(n3426), .dinb(n3425), .dout(n3427));
  jand g03172(.dina(n3353), .dinb(n3275), .dout(n3428));
  jand g03173(.dina(n3354), .dinb(n3266), .dout(n3429));
  jor  g03174(.dina(n3429), .dinb(n3428), .dout(n3430));
  jor  g03175(.dina(n3351), .dinb(n3343), .dout(n3431));
  jand g03176(.dina(n3352), .dinb(n3278), .dout(n3432));
  jnot g03177(.din(n3432), .dout(n3433));
  jand g03178(.dina(n3433), .dinb(n3431), .dout(n3434));
  jnot g03179(.din(n3434), .dout(n3435));
  jor  g03180(.dina(n3340), .dinb(n3332), .dout(n3436));
  jand g03181(.dina(n3341), .dinb(n3283), .dout(n3437));
  jnot g03182(.din(n3437), .dout(n3438));
  jand g03183(.dina(n3438), .dinb(n3436), .dout(n3439));
  jnot g03184(.din(n3439), .dout(n3440));
  jand g03185(.dina(n3329), .dinb(n3297), .dout(n3441));
  jand g03186(.dina(n3330), .dinb(n3288), .dout(n3442));
  jor  g03187(.dina(n3442), .dinb(n3441), .dout(n3443));
  jor  g03188(.dina(n3327), .dinb(n3319), .dout(n3444));
  jand g03189(.dina(n3328), .dinb(n3300), .dout(n3445));
  jnot g03190(.din(n3445), .dout(n3446));
  jand g03191(.dina(n3446), .dinb(n3444), .dout(n3447));
  jnot g03192(.din(n3447), .dout(n3448));
  jor  g03193(.dina(n2784), .dinb(n428), .dout(n3449));
  jor  g03194(.dina(n2661), .dinb(n357), .dout(n3450));
  jor  g03195(.dina(n2787), .dinb(n395), .dout(n3451));
  jor  g03196(.dina(n2789), .dinb(n431), .dout(n3452));
  jand g03197(.dina(n3452), .dinb(n3451), .dout(n3453));
  jand g03198(.dina(n3453), .dinb(n3450), .dout(n3454));
  jand g03199(.dina(n3454), .dinb(n3449), .dout(n3455));
  jxor g03200(.dina(n3455), .dinb(a29 ), .dout(n3456));
  jnot g03201(.din(n3456), .dout(n3457));
  jnot g03202(.din(n3316), .dout(n3458));
  jand g03203(.dina(n3458), .dinb(n3314), .dout(n3459));
  jand g03204(.dina(n3317), .dinb(n3312), .dout(n3460));
  jor  g03205(.dina(n3460), .dinb(n3459), .dout(n3461));
  jor  g03206(.dina(n3301), .dinb(n319), .dout(n3462));
  jor  g03207(.dina(n3136), .dinb(n279), .dout(n3463));
  jor  g03208(.dina(n3304), .dinb(n299), .dout(n3464));
  jor  g03209(.dina(n3306), .dinb(n322), .dout(n3465));
  jand g03210(.dina(n3465), .dinb(n3464), .dout(n3466));
  jand g03211(.dina(n3466), .dinb(n3463), .dout(n3467));
  jand g03212(.dina(n3467), .dinb(n3462), .dout(n3468));
  jxor g03213(.dina(n3468), .dinb(a32 ), .dout(n3469));
  jnot g03214(.din(n3469), .dout(n3470));
  jand g03215(.dina(n3314), .dinb(a35 ), .dout(n3471));
  jxor g03216(.dina(a35 ), .dinb(a34 ), .dout(n3472));
  jnot g03217(.din(n3472), .dout(n3473));
  jand g03218(.dina(n3473), .dinb(n3313), .dout(n3474));
  jand g03219(.dina(n3474), .dinb(b1 ), .dout(n3475));
  jnot g03220(.din(n3313), .dout(n3476));
  jxor g03221(.dina(a34 ), .dinb(a33 ), .dout(n3477));
  jand g03222(.dina(n3477), .dinb(n3476), .dout(n3478));
  jand g03223(.dina(n3478), .dinb(b0 ), .dout(n3479));
  jand g03224(.dina(n3472), .dinb(n3313), .dout(n3480));
  jand g03225(.dina(n3480), .dinb(n338), .dout(n3481));
  jor  g03226(.dina(n3481), .dinb(n3479), .dout(n3482));
  jor  g03227(.dina(n3482), .dinb(n3475), .dout(n3483));
  jxor g03228(.dina(n3483), .dinb(n3471), .dout(n3484));
  jxor g03229(.dina(n3484), .dinb(n3470), .dout(n3485));
  jxor g03230(.dina(n3485), .dinb(n3461), .dout(n3486));
  jxor g03231(.dina(n3486), .dinb(n3457), .dout(n3487));
  jxor g03232(.dina(n3487), .dinb(n3448), .dout(n3488));
  jnot g03233(.din(n3488), .dout(n3489));
  jor  g03234(.dina(n2319), .dinb(n624), .dout(n3490));
  jor  g03235(.dina(n2224), .dinb(n512), .dout(n3491));
  jor  g03236(.dina(n2322), .dinb(n564), .dout(n3492));
  jor  g03237(.dina(n2324), .dinb(n627), .dout(n3493));
  jand g03238(.dina(n3493), .dinb(n3492), .dout(n3494));
  jand g03239(.dina(n3494), .dinb(n3491), .dout(n3495));
  jand g03240(.dina(n3495), .dinb(n3490), .dout(n3496));
  jxor g03241(.dina(n3496), .dinb(a26 ), .dout(n3497));
  jxor g03242(.dina(n3497), .dinb(n3489), .dout(n3498));
  jxor g03243(.dina(n3498), .dinb(n3443), .dout(n3499));
  jnot g03244(.din(n3499), .dout(n3500));
  jor  g03245(.dina(n1939), .dinb(n775), .dout(n3501));
  jor  g03246(.dina(n1827), .dinb(n647), .dout(n3502));
  jor  g03247(.dina(n1942), .dinb(n758), .dout(n3503));
  jor  g03248(.dina(n1944), .dinb(n778), .dout(n3504));
  jand g03249(.dina(n3504), .dinb(n3503), .dout(n3505));
  jand g03250(.dina(n3505), .dinb(n3502), .dout(n3506));
  jand g03251(.dina(n3506), .dinb(n3501), .dout(n3507));
  jxor g03252(.dina(n3507), .dinb(a23 ), .dout(n3508));
  jxor g03253(.dina(n3508), .dinb(n3500), .dout(n3509));
  jxor g03254(.dina(n3509), .dinb(n3440), .dout(n3510));
  jnot g03255(.din(n3510), .dout(n3511));
  jor  g03256(.dina(n1566), .dinb(n1019), .dout(n3512));
  jor  g03257(.dina(n1489), .dinb(n858), .dout(n3513));
  jor  g03258(.dina(n1569), .dinb(n939), .dout(n3514));
  jor  g03259(.dina(n1571), .dinb(n1022), .dout(n3515));
  jand g03260(.dina(n3515), .dinb(n3514), .dout(n3516));
  jand g03261(.dina(n3516), .dinb(n3513), .dout(n3517));
  jand g03262(.dina(n3517), .dinb(n3512), .dout(n3518));
  jxor g03263(.dina(n3518), .dinb(a20 ), .dout(n3519));
  jxor g03264(.dina(n3519), .dinb(n3511), .dout(n3520));
  jxor g03265(.dina(n3520), .dinb(n3435), .dout(n3521));
  jnot g03266(.din(n3521), .dout(n3522));
  jor  g03267(.dina(n1397), .dinb(n1245), .dout(n3523));
  jor  g03268(.dina(n1165), .dinb(n1193), .dout(n3524));
  jor  g03269(.dina(n1248), .dinb(n1290), .dout(n3525));
  jor  g03270(.dina(n1250), .dinb(n1400), .dout(n3526));
  jand g03271(.dina(n3526), .dinb(n3525), .dout(n3527));
  jand g03272(.dina(n3527), .dinb(n3524), .dout(n3528));
  jand g03273(.dina(n3528), .dinb(n3523), .dout(n3529));
  jxor g03274(.dina(n3529), .dinb(a17 ), .dout(n3530));
  jxor g03275(.dina(n3530), .dinb(n3522), .dout(n3531));
  jxor g03276(.dina(n3531), .dinb(n3430), .dout(n3532));
  jor  g03277(.dina(n1739), .dinb(n974), .dout(n3533));
  jor  g03278(.dina(n908), .dinb(n1420), .dout(n3534));
  jor  g03279(.dina(n977), .dinb(n1620), .dout(n3535));
  jor  g03280(.dina(n979), .dinb(n1742), .dout(n3536));
  jand g03281(.dina(n3536), .dinb(n3535), .dout(n3537));
  jand g03282(.dina(n3537), .dinb(n3534), .dout(n3538));
  jand g03283(.dina(n3538), .dinb(n3533), .dout(n3539));
  jxor g03284(.dina(n3539), .dinb(a14 ), .dout(n3540));
  jxor g03285(.dina(n3540), .dinb(n3532), .dout(n3541));
  jnot g03286(.din(n3541), .dout(n3542));
  jxor g03287(.dina(n3542), .dinb(n3427), .dout(n3543));
  jor  g03288(.dina(n2007), .dinb(n706), .dout(n3544));
  jor  g03289(.dina(n683), .dinb(n1867), .dout(n3545));
  jor  g03290(.dina(n709), .dinb(n1887), .dout(n3546));
  jor  g03291(.dina(n711), .dinb(n2010), .dout(n3547));
  jand g03292(.dina(n3547), .dinb(n3546), .dout(n3548));
  jand g03293(.dina(n3548), .dinb(n3545), .dout(n3549));
  jand g03294(.dina(n3549), .dinb(n3544), .dout(n3550));
  jxor g03295(.dina(n3550), .dinb(a11 ), .dout(n3551));
  jxor g03296(.dina(n3551), .dinb(n3543), .dout(n3552));
  jxor g03297(.dina(n3552), .dinb(n3422), .dout(n3553));
  jnot g03298(.din(n3553), .dout(n3554));
  jor  g03299(.dina(n2556), .dinb(n528), .dout(n3555));
  jor  g03300(.dina(n490), .dinb(n2148), .dout(n3556));
  jor  g03301(.dina(n531), .dinb(n2407), .dout(n3557));
  jor  g03302(.dina(n533), .dinb(n2559), .dout(n3558));
  jand g03303(.dina(n3558), .dinb(n3557), .dout(n3559));
  jand g03304(.dina(n3559), .dinb(n3556), .dout(n3560));
  jand g03305(.dina(n3560), .dinb(n3555), .dout(n3561));
  jxor g03306(.dina(n3561), .dinb(a8 ), .dout(n3562));
  jxor g03307(.dina(n3562), .dinb(n3554), .dout(n3563));
  jxor g03308(.dina(n3563), .dinb(n3418), .dout(n3564));
  jor  g03309(.dina(n3032), .dinb(n402), .dout(n3565));
  jor  g03310(.dina(n371), .dinb(n2579), .dout(n3566));
  jor  g03311(.dina(n405), .dinb(n2870), .dout(n3567));
  jor  g03312(.dina(n332), .dinb(n3035), .dout(n3568));
  jand g03313(.dina(n3568), .dinb(n3567), .dout(n3569));
  jand g03314(.dina(n3569), .dinb(n3566), .dout(n3570));
  jand g03315(.dina(n3570), .dinb(n3565), .dout(n3571));
  jxor g03316(.dina(n3571), .dinb(a5 ), .dout(n3572));
  jxor g03317(.dina(n3572), .dinb(n3564), .dout(n3573));
  jxor g03318(.dina(n3573), .dinb(n3413), .dout(n3574));
  jxor g03319(.dina(n3574), .dinb(n3409), .dout(n3575));
  jxor g03320(.dina(n3575), .dinb(n3394), .dout(f34 ));
  jand g03321(.dina(n3574), .dinb(n3409), .dout(n3577));
  jand g03322(.dina(n3575), .dinb(n3394), .dout(n3578));
  jor  g03323(.dina(n3578), .dinb(n3577), .dout(n3579));
  jand g03324(.dina(b34 ), .dinb(b33 ), .dout(n3580));
  jand g03325(.dina(n3398), .dinb(n3397), .dout(n3581));
  jor  g03326(.dina(n3581), .dinb(n3580), .dout(n3582));
  jxor g03327(.dina(b35 ), .dinb(b34 ), .dout(n3583));
  jnot g03328(.din(n3583), .dout(n3584));
  jxor g03329(.dina(n3584), .dinb(n3582), .dout(n3585));
  jor  g03330(.dina(n3585), .dinb(n264), .dout(n3586));
  jor  g03331(.dina(n284), .dinb(n3230), .dout(n3587));
  jnot g03332(.din(b35 ), .dout(n3588));
  jor  g03333(.dina(n269), .dinb(n3588), .dout(n3589));
  jor  g03334(.dina(n271), .dinb(n3403), .dout(n3590));
  jand g03335(.dina(n3590), .dinb(n3589), .dout(n3591));
  jand g03336(.dina(n3591), .dinb(n3587), .dout(n3592));
  jand g03337(.dina(n3592), .dinb(n3586), .dout(n3593));
  jxor g03338(.dina(n3593), .dinb(n260), .dout(n3594));
  jor  g03339(.dina(n3572), .dinb(n3564), .dout(n3595));
  jnot g03340(.din(n3595), .dout(n3596));
  jand g03341(.dina(n3573), .dinb(n3413), .dout(n3597));
  jor  g03342(.dina(n3597), .dinb(n3596), .dout(n3598));
  jor  g03343(.dina(n3562), .dinb(n3554), .dout(n3599));
  jnot g03344(.din(n3599), .dout(n3600));
  jand g03345(.dina(n3563), .dinb(n3417), .dout(n3601));
  jor  g03346(.dina(n3601), .dinb(n3600), .dout(n3602));
  jnot g03347(.din(n3602), .dout(n3603));
  jnot g03348(.din(n3543), .dout(n3604));
  jor  g03349(.dina(n3551), .dinb(n3604), .dout(n3605));
  jor  g03350(.dina(n3552), .dinb(n3422), .dout(n3606));
  jand g03351(.dina(n3606), .dinb(n3605), .dout(n3607));
  jor  g03352(.dina(n2145), .dinb(n706), .dout(n3608));
  jor  g03353(.dina(n683), .dinb(n1887), .dout(n3609));
  jor  g03354(.dina(n709), .dinb(n2010), .dout(n3610));
  jor  g03355(.dina(n711), .dinb(n2148), .dout(n3611));
  jand g03356(.dina(n3611), .dinb(n3610), .dout(n3612));
  jand g03357(.dina(n3612), .dinb(n3609), .dout(n3613));
  jand g03358(.dina(n3613), .dinb(n3608), .dout(n3614));
  jxor g03359(.dina(n3614), .dinb(a11 ), .dout(n3615));
  jnot g03360(.din(n3615), .dout(n3616));
  jnot g03361(.din(n3532), .dout(n3617));
  jor  g03362(.dina(n3540), .dinb(n3617), .dout(n3618));
  jnot g03363(.din(n3618), .dout(n3619));
  jand g03364(.dina(n3542), .dinb(n3427), .dout(n3620));
  jor  g03365(.dina(n3620), .dinb(n3619), .dout(n3621));
  jor  g03366(.dina(n1864), .dinb(n974), .dout(n3622));
  jor  g03367(.dina(n908), .dinb(n1620), .dout(n3623));
  jor  g03368(.dina(n977), .dinb(n1742), .dout(n3624));
  jor  g03369(.dina(n979), .dinb(n1867), .dout(n3625));
  jand g03370(.dina(n3625), .dinb(n3624), .dout(n3626));
  jand g03371(.dina(n3626), .dinb(n3623), .dout(n3627));
  jand g03372(.dina(n3627), .dinb(n3622), .dout(n3628));
  jxor g03373(.dina(n3628), .dinb(a14 ), .dout(n3629));
  jnot g03374(.din(n3629), .dout(n3630));
  jor  g03375(.dina(n3530), .dinb(n3522), .dout(n3631));
  jnot g03376(.din(n3631), .dout(n3632));
  jand g03377(.dina(n3531), .dinb(n3430), .dout(n3633));
  jor  g03378(.dina(n3633), .dinb(n3632), .dout(n3634));
  jor  g03379(.dina(n3519), .dinb(n3511), .dout(n3635));
  jand g03380(.dina(n3520), .dinb(n3435), .dout(n3636));
  jnot g03381(.din(n3636), .dout(n3637));
  jand g03382(.dina(n3637), .dinb(n3635), .dout(n3638));
  jnot g03383(.din(n3638), .dout(n3639));
  jor  g03384(.dina(n3508), .dinb(n3500), .dout(n3640));
  jand g03385(.dina(n3509), .dinb(n3440), .dout(n3641));
  jnot g03386(.din(n3641), .dout(n3642));
  jand g03387(.dina(n3642), .dinb(n3640), .dout(n3643));
  jnot g03388(.din(n3643), .dout(n3644));
  jor  g03389(.dina(n1939), .dinb(n855), .dout(n3645));
  jor  g03390(.dina(n1827), .dinb(n758), .dout(n3646));
  jor  g03391(.dina(n1942), .dinb(n778), .dout(n3647));
  jor  g03392(.dina(n1944), .dinb(n858), .dout(n3648));
  jand g03393(.dina(n3648), .dinb(n3647), .dout(n3649));
  jand g03394(.dina(n3649), .dinb(n3646), .dout(n3650));
  jand g03395(.dina(n3650), .dinb(n3645), .dout(n3651));
  jxor g03396(.dina(n3651), .dinb(a23 ), .dout(n3652));
  jnot g03397(.din(n3652), .dout(n3653));
  jor  g03398(.dina(n3497), .dinb(n3489), .dout(n3654));
  jand g03399(.dina(n3498), .dinb(n3443), .dout(n3655));
  jnot g03400(.din(n3655), .dout(n3656));
  jand g03401(.dina(n3656), .dinb(n3654), .dout(n3657));
  jnot g03402(.din(n3657), .dout(n3658));
  jor  g03403(.dina(n2319), .dinb(n644), .dout(n3659));
  jor  g03404(.dina(n2224), .dinb(n564), .dout(n3660));
  jor  g03405(.dina(n2322), .dinb(n627), .dout(n3661));
  jor  g03406(.dina(n2324), .dinb(n647), .dout(n3662));
  jand g03407(.dina(n3662), .dinb(n3661), .dout(n3663));
  jand g03408(.dina(n3663), .dinb(n3660), .dout(n3664));
  jand g03409(.dina(n3664), .dinb(n3659), .dout(n3665));
  jxor g03410(.dina(n3665), .dinb(a26 ), .dout(n3666));
  jnot g03411(.din(n3666), .dout(n3667));
  jand g03412(.dina(n3486), .dinb(n3457), .dout(n3668));
  jand g03413(.dina(n3487), .dinb(n3448), .dout(n3669));
  jor  g03414(.dina(n3669), .dinb(n3668), .dout(n3670));
  jand g03415(.dina(n3484), .dinb(n3470), .dout(n3671));
  jand g03416(.dina(n3485), .dinb(n3461), .dout(n3672));
  jor  g03417(.dina(n3672), .dinb(n3671), .dout(n3673));
  jor  g03418(.dina(n3301), .dinb(n354), .dout(n3674));
  jor  g03419(.dina(n3136), .dinb(n299), .dout(n3675));
  jor  g03420(.dina(n3304), .dinb(n322), .dout(n3676));
  jor  g03421(.dina(n3306), .dinb(n357), .dout(n3677));
  jand g03422(.dina(n3677), .dinb(n3676), .dout(n3678));
  jand g03423(.dina(n3678), .dinb(n3675), .dout(n3679));
  jand g03424(.dina(n3679), .dinb(n3674), .dout(n3680));
  jxor g03425(.dina(n3680), .dinb(a32 ), .dout(n3681));
  jnot g03426(.din(n3681), .dout(n3682));
  jnot g03427(.din(n3483), .dout(n3683));
  jand g03428(.dina(n3315), .dinb(a35 ), .dout(n3684));
  jand g03429(.dina(n3684), .dinb(n3683), .dout(n3685));
  jnot g03430(.din(n3685), .dout(n3686));
  jand g03431(.dina(n3686), .dinb(a35 ), .dout(n3687));
  jor  g03432(.dina(n3477), .dinb(n3473), .dout(n3688));
  jor  g03433(.dina(n3688), .dinb(n3313), .dout(n3689));
  jnot g03434(.din(n3689), .dout(n3690));
  jand g03435(.dina(n3690), .dinb(b0 ), .dout(n3691));
  jand g03436(.dina(n3474), .dinb(b2 ), .dout(n3692));
  jand g03437(.dina(n3478), .dinb(b1 ), .dout(n3693));
  jand g03438(.dina(n3480), .dinb(n375), .dout(n3694));
  jor  g03439(.dina(n3694), .dinb(n3693), .dout(n3695));
  jor  g03440(.dina(n3695), .dinb(n3692), .dout(n3696));
  jor  g03441(.dina(n3696), .dinb(n3691), .dout(n3697));
  jxor g03442(.dina(n3697), .dinb(n3687), .dout(n3698));
  jxor g03443(.dina(n3698), .dinb(n3682), .dout(n3699));
  jxor g03444(.dina(n3699), .dinb(n3673), .dout(n3700));
  jnot g03445(.din(n3700), .dout(n3701));
  jor  g03446(.dina(n2784), .dinb(n509), .dout(n3702));
  jor  g03447(.dina(n2661), .dinb(n395), .dout(n3703));
  jor  g03448(.dina(n2787), .dinb(n431), .dout(n3704));
  jor  g03449(.dina(n2789), .dinb(n512), .dout(n3705));
  jand g03450(.dina(n3705), .dinb(n3704), .dout(n3706));
  jand g03451(.dina(n3706), .dinb(n3703), .dout(n3707));
  jand g03452(.dina(n3707), .dinb(n3702), .dout(n3708));
  jxor g03453(.dina(n3708), .dinb(a29 ), .dout(n3709));
  jxor g03454(.dina(n3709), .dinb(n3701), .dout(n3710));
  jxor g03455(.dina(n3710), .dinb(n3670), .dout(n3711));
  jxor g03456(.dina(n3711), .dinb(n3667), .dout(n3712));
  jxor g03457(.dina(n3712), .dinb(n3658), .dout(n3713));
  jxor g03458(.dina(n3713), .dinb(n3653), .dout(n3714));
  jxor g03459(.dina(n3714), .dinb(n3644), .dout(n3715));
  jnot g03460(.din(n3715), .dout(n3716));
  jor  g03461(.dina(n1566), .dinb(n1190), .dout(n3717));
  jor  g03462(.dina(n1489), .dinb(n939), .dout(n3718));
  jor  g03463(.dina(n1569), .dinb(n1022), .dout(n3719));
  jor  g03464(.dina(n1571), .dinb(n1193), .dout(n3720));
  jand g03465(.dina(n3720), .dinb(n3719), .dout(n3721));
  jand g03466(.dina(n3721), .dinb(n3718), .dout(n3722));
  jand g03467(.dina(n3722), .dinb(n3717), .dout(n3723));
  jxor g03468(.dina(n3723), .dinb(a20 ), .dout(n3724));
  jxor g03469(.dina(n3724), .dinb(n3716), .dout(n3725));
  jxor g03470(.dina(n3725), .dinb(n3639), .dout(n3726));
  jnot g03471(.din(n3726), .dout(n3727));
  jor  g03472(.dina(n1417), .dinb(n1245), .dout(n3728));
  jor  g03473(.dina(n1165), .dinb(n1290), .dout(n3729));
  jor  g03474(.dina(n1248), .dinb(n1400), .dout(n3730));
  jor  g03475(.dina(n1250), .dinb(n1420), .dout(n3731));
  jand g03476(.dina(n3731), .dinb(n3730), .dout(n3732));
  jand g03477(.dina(n3732), .dinb(n3729), .dout(n3733));
  jand g03478(.dina(n3733), .dinb(n3728), .dout(n3734));
  jxor g03479(.dina(n3734), .dinb(a17 ), .dout(n3735));
  jxor g03480(.dina(n3735), .dinb(n3727), .dout(n3736));
  jxor g03481(.dina(n3736), .dinb(n3634), .dout(n3737));
  jxor g03482(.dina(n3737), .dinb(n3630), .dout(n3738));
  jxor g03483(.dina(n3738), .dinb(n3621), .dout(n3739));
  jxor g03484(.dina(n3739), .dinb(n3616), .dout(n3740));
  jnot g03485(.din(n3740), .dout(n3741));
  jxor g03486(.dina(n3741), .dinb(n3607), .dout(n3742));
  jnot g03487(.din(n3742), .dout(n3743));
  jor  g03488(.dina(n2576), .dinb(n528), .dout(n3744));
  jor  g03489(.dina(n490), .dinb(n2407), .dout(n3745));
  jor  g03490(.dina(n531), .dinb(n2559), .dout(n3746));
  jor  g03491(.dina(n533), .dinb(n2579), .dout(n3747));
  jand g03492(.dina(n3747), .dinb(n3746), .dout(n3748));
  jand g03493(.dina(n3748), .dinb(n3745), .dout(n3749));
  jand g03494(.dina(n3749), .dinb(n3744), .dout(n3750));
  jxor g03495(.dina(n3750), .dinb(a8 ), .dout(n3751));
  jxor g03496(.dina(n3751), .dinb(n3743), .dout(n3752));
  jxor g03497(.dina(n3752), .dinb(n3603), .dout(n3753));
  jor  g03498(.dina(n3052), .dinb(n402), .dout(n3754));
  jor  g03499(.dina(n371), .dinb(n2870), .dout(n3755));
  jor  g03500(.dina(n405), .dinb(n3035), .dout(n3756));
  jor  g03501(.dina(n332), .dinb(n3055), .dout(n3757));
  jand g03502(.dina(n3757), .dinb(n3756), .dout(n3758));
  jand g03503(.dina(n3758), .dinb(n3755), .dout(n3759));
  jand g03504(.dina(n3759), .dinb(n3754), .dout(n3760));
  jxor g03505(.dina(n3760), .dinb(a5 ), .dout(n3761));
  jxor g03506(.dina(n3761), .dinb(n3753), .dout(n3762));
  jxor g03507(.dina(n3762), .dinb(n3598), .dout(n3763));
  jxor g03508(.dina(n3763), .dinb(n3594), .dout(n3764));
  jxor g03509(.dina(n3764), .dinb(n3579), .dout(f35 ));
  jand g03510(.dina(n3763), .dinb(n3594), .dout(n3766));
  jand g03511(.dina(n3764), .dinb(n3579), .dout(n3767));
  jor  g03512(.dina(n3767), .dinb(n3766), .dout(n3768));
  jor  g03513(.dina(n3761), .dinb(n3753), .dout(n3769));
  jnot g03514(.din(n3769), .dout(n3770));
  jand g03515(.dina(n3762), .dinb(n3598), .dout(n3771));
  jor  g03516(.dina(n3771), .dinb(n3770), .dout(n3772));
  jor  g03517(.dina(n3227), .dinb(n402), .dout(n3773));
  jor  g03518(.dina(n371), .dinb(n3035), .dout(n3774));
  jor  g03519(.dina(n405), .dinb(n3055), .dout(n3775));
  jor  g03520(.dina(n332), .dinb(n3230), .dout(n3776));
  jand g03521(.dina(n3776), .dinb(n3775), .dout(n3777));
  jand g03522(.dina(n3777), .dinb(n3774), .dout(n3778));
  jand g03523(.dina(n3778), .dinb(n3773), .dout(n3779));
  jxor g03524(.dina(n3779), .dinb(a5 ), .dout(n3780));
  jnot g03525(.din(n3780), .dout(n3781));
  jor  g03526(.dina(n3751), .dinb(n3743), .dout(n3782));
  jnot g03527(.din(n3782), .dout(n3783));
  jand g03528(.dina(n3752), .dinb(n3602), .dout(n3784));
  jor  g03529(.dina(n3784), .dinb(n3783), .dout(n3785));
  jor  g03530(.dina(n2867), .dinb(n528), .dout(n3786));
  jor  g03531(.dina(n490), .dinb(n2559), .dout(n3787));
  jor  g03532(.dina(n531), .dinb(n2579), .dout(n3788));
  jor  g03533(.dina(n533), .dinb(n2870), .dout(n3789));
  jand g03534(.dina(n3789), .dinb(n3788), .dout(n3790));
  jand g03535(.dina(n3790), .dinb(n3787), .dout(n3791));
  jand g03536(.dina(n3791), .dinb(n3786), .dout(n3792));
  jxor g03537(.dina(n3792), .dinb(a8 ), .dout(n3793));
  jnot g03538(.din(n3793), .dout(n3794));
  jand g03539(.dina(n3739), .dinb(n3616), .dout(n3795));
  jnot g03540(.din(n3795), .dout(n3796));
  jor  g03541(.dina(n3741), .dinb(n3607), .dout(n3797));
  jand g03542(.dina(n3797), .dinb(n3796), .dout(n3798));
  jand g03543(.dina(n3737), .dinb(n3630), .dout(n3799));
  jand g03544(.dina(n3738), .dinb(n3621), .dout(n3800));
  jor  g03545(.dina(n3800), .dinb(n3799), .dout(n3801));
  jor  g03546(.dina(n1884), .dinb(n974), .dout(n3802));
  jor  g03547(.dina(n908), .dinb(n1742), .dout(n3803));
  jor  g03548(.dina(n977), .dinb(n1867), .dout(n3804));
  jor  g03549(.dina(n979), .dinb(n1887), .dout(n3805));
  jand g03550(.dina(n3805), .dinb(n3804), .dout(n3806));
  jand g03551(.dina(n3806), .dinb(n3803), .dout(n3807));
  jand g03552(.dina(n3807), .dinb(n3802), .dout(n3808));
  jxor g03553(.dina(n3808), .dinb(a14 ), .dout(n3809));
  jnot g03554(.din(n3809), .dout(n3810));
  jor  g03555(.dina(n3735), .dinb(n3727), .dout(n3811));
  jnot g03556(.din(n3811), .dout(n3812));
  jand g03557(.dina(n3736), .dinb(n3634), .dout(n3813));
  jor  g03558(.dina(n3813), .dinb(n3812), .dout(n3814));
  jor  g03559(.dina(n3724), .dinb(n3716), .dout(n3815));
  jand g03560(.dina(n3725), .dinb(n3639), .dout(n3816));
  jnot g03561(.din(n3816), .dout(n3817));
  jand g03562(.dina(n3817), .dinb(n3815), .dout(n3818));
  jnot g03563(.din(n3818), .dout(n3819));
  jor  g03564(.dina(n1566), .dinb(n1287), .dout(n3820));
  jor  g03565(.dina(n1489), .dinb(n1022), .dout(n3821));
  jor  g03566(.dina(n1569), .dinb(n1193), .dout(n3822));
  jor  g03567(.dina(n1571), .dinb(n1290), .dout(n3823));
  jand g03568(.dina(n3823), .dinb(n3822), .dout(n3824));
  jand g03569(.dina(n3824), .dinb(n3821), .dout(n3825));
  jand g03570(.dina(n3825), .dinb(n3820), .dout(n3826));
  jxor g03571(.dina(n3826), .dinb(a20 ), .dout(n3827));
  jnot g03572(.din(n3827), .dout(n3828));
  jand g03573(.dina(n3713), .dinb(n3653), .dout(n3829));
  jand g03574(.dina(n3714), .dinb(n3644), .dout(n3830));
  jor  g03575(.dina(n3830), .dinb(n3829), .dout(n3831));
  jor  g03576(.dina(n3709), .dinb(n3701), .dout(n3832));
  jand g03577(.dina(n3710), .dinb(n3670), .dout(n3833));
  jnot g03578(.din(n3833), .dout(n3834));
  jand g03579(.dina(n3834), .dinb(n3832), .dout(n3835));
  jnot g03580(.din(n3835), .dout(n3836));
  jor  g03581(.dina(n2784), .dinb(n561), .dout(n3837));
  jor  g03582(.dina(n2661), .dinb(n431), .dout(n3838));
  jor  g03583(.dina(n2787), .dinb(n512), .dout(n3839));
  jor  g03584(.dina(n2789), .dinb(n564), .dout(n3840));
  jand g03585(.dina(n3840), .dinb(n3839), .dout(n3841));
  jand g03586(.dina(n3841), .dinb(n3838), .dout(n3842));
  jand g03587(.dina(n3842), .dinb(n3837), .dout(n3843));
  jxor g03588(.dina(n3843), .dinb(a29 ), .dout(n3844));
  jnot g03589(.din(n3844), .dout(n3845));
  jand g03590(.dina(n3698), .dinb(n3682), .dout(n3846));
  jand g03591(.dina(n3699), .dinb(n3673), .dout(n3847));
  jor  g03592(.dina(n3847), .dinb(n3846), .dout(n3848));
  jnot g03593(.din(n3480), .dout(n3849));
  jor  g03594(.dina(n3849), .dinb(n296), .dout(n3850));
  jor  g03595(.dina(n3689), .dinb(n267), .dout(n3851));
  jnot g03596(.din(n3478), .dout(n3852));
  jor  g03597(.dina(n3852), .dinb(n279), .dout(n3853));
  jnot g03598(.din(n3474), .dout(n3854));
  jor  g03599(.dina(n3854), .dinb(n299), .dout(n3855));
  jand g03600(.dina(n3855), .dinb(n3853), .dout(n3856));
  jand g03601(.dina(n3856), .dinb(n3851), .dout(n3857));
  jand g03602(.dina(n3857), .dinb(n3850), .dout(n3858));
  jxor g03603(.dina(n3858), .dinb(a35 ), .dout(n3859));
  jnot g03604(.din(n3859), .dout(n3860));
  jxor g03605(.dina(a36 ), .dinb(a35 ), .dout(n3861));
  jand g03606(.dina(n3861), .dinb(b0 ), .dout(n3862));
  jnot g03607(.din(n3862), .dout(n3863));
  jor  g03608(.dina(n3697), .dinb(n3686), .dout(n3864));
  jxor g03609(.dina(n3864), .dinb(n3863), .dout(n3865));
  jxor g03610(.dina(n3865), .dinb(n3860), .dout(n3866));
  jnot g03611(.din(n3866), .dout(n3867));
  jor  g03612(.dina(n3301), .dinb(n392), .dout(n3868));
  jor  g03613(.dina(n3136), .dinb(n322), .dout(n3869));
  jor  g03614(.dina(n3304), .dinb(n357), .dout(n3870));
  jor  g03615(.dina(n3306), .dinb(n395), .dout(n3871));
  jand g03616(.dina(n3871), .dinb(n3870), .dout(n3872));
  jand g03617(.dina(n3872), .dinb(n3869), .dout(n3873));
  jand g03618(.dina(n3873), .dinb(n3868), .dout(n3874));
  jxor g03619(.dina(n3874), .dinb(a32 ), .dout(n3875));
  jxor g03620(.dina(n3875), .dinb(n3867), .dout(n3876));
  jxor g03621(.dina(n3876), .dinb(n3848), .dout(n3877));
  jxor g03622(.dina(n3877), .dinb(n3845), .dout(n3878));
  jxor g03623(.dina(n3878), .dinb(n3836), .dout(n3879));
  jnot g03624(.din(n3879), .dout(n3880));
  jor  g03625(.dina(n2319), .dinb(n755), .dout(n3881));
  jor  g03626(.dina(n2224), .dinb(n627), .dout(n3882));
  jor  g03627(.dina(n2322), .dinb(n647), .dout(n3883));
  jor  g03628(.dina(n2324), .dinb(n758), .dout(n3884));
  jand g03629(.dina(n3884), .dinb(n3883), .dout(n3885));
  jand g03630(.dina(n3885), .dinb(n3882), .dout(n3886));
  jand g03631(.dina(n3886), .dinb(n3881), .dout(n3887));
  jxor g03632(.dina(n3887), .dinb(a26 ), .dout(n3888));
  jxor g03633(.dina(n3888), .dinb(n3880), .dout(n3889));
  jand g03634(.dina(n3711), .dinb(n3667), .dout(n3890));
  jand g03635(.dina(n3712), .dinb(n3658), .dout(n3891));
  jor  g03636(.dina(n3891), .dinb(n3890), .dout(n3892));
  jxor g03637(.dina(n3892), .dinb(n3889), .dout(n3893));
  jnot g03638(.din(n3893), .dout(n3894));
  jor  g03639(.dina(n1939), .dinb(n936), .dout(n3895));
  jor  g03640(.dina(n1827), .dinb(n778), .dout(n3896));
  jor  g03641(.dina(n1942), .dinb(n858), .dout(n3897));
  jor  g03642(.dina(n1944), .dinb(n939), .dout(n3898));
  jand g03643(.dina(n3898), .dinb(n3897), .dout(n3899));
  jand g03644(.dina(n3899), .dinb(n3896), .dout(n3900));
  jand g03645(.dina(n3900), .dinb(n3895), .dout(n3901));
  jxor g03646(.dina(n3901), .dinb(a23 ), .dout(n3902));
  jxor g03647(.dina(n3902), .dinb(n3894), .dout(n3903));
  jxor g03648(.dina(n3903), .dinb(n3831), .dout(n3904));
  jxor g03649(.dina(n3904), .dinb(n3828), .dout(n3905));
  jxor g03650(.dina(n3905), .dinb(n3819), .dout(n3906));
  jnot g03651(.din(n3906), .dout(n3907));
  jor  g03652(.dina(n1617), .dinb(n1245), .dout(n3908));
  jor  g03653(.dina(n1165), .dinb(n1400), .dout(n3909));
  jor  g03654(.dina(n1248), .dinb(n1420), .dout(n3910));
  jor  g03655(.dina(n1250), .dinb(n1620), .dout(n3911));
  jand g03656(.dina(n3911), .dinb(n3910), .dout(n3912));
  jand g03657(.dina(n3912), .dinb(n3909), .dout(n3913));
  jand g03658(.dina(n3913), .dinb(n3908), .dout(n3914));
  jxor g03659(.dina(n3914), .dinb(a17 ), .dout(n3915));
  jxor g03660(.dina(n3915), .dinb(n3907), .dout(n3916));
  jxor g03661(.dina(n3916), .dinb(n3814), .dout(n3917));
  jxor g03662(.dina(n3917), .dinb(n3810), .dout(n3918));
  jxor g03663(.dina(n3918), .dinb(n3801), .dout(n3919));
  jor  g03664(.dina(n2404), .dinb(n706), .dout(n3920));
  jor  g03665(.dina(n683), .dinb(n2010), .dout(n3921));
  jor  g03666(.dina(n709), .dinb(n2148), .dout(n3922));
  jor  g03667(.dina(n711), .dinb(n2407), .dout(n3923));
  jand g03668(.dina(n3923), .dinb(n3922), .dout(n3924));
  jand g03669(.dina(n3924), .dinb(n3921), .dout(n3925));
  jand g03670(.dina(n3925), .dinb(n3920), .dout(n3926));
  jxor g03671(.dina(n3926), .dinb(a11 ), .dout(n3927));
  jxor g03672(.dina(n3927), .dinb(n3919), .dout(n3928));
  jxor g03673(.dina(n3928), .dinb(n3798), .dout(n3929));
  jxor g03674(.dina(n3929), .dinb(n3794), .dout(n3930));
  jxor g03675(.dina(n3930), .dinb(n3785), .dout(n3931));
  jxor g03676(.dina(n3931), .dinb(n3781), .dout(n3932));
  jxor g03677(.dina(n3932), .dinb(n3772), .dout(n3933));
  jand g03678(.dina(b35 ), .dinb(b34 ), .dout(n3934));
  jand g03679(.dina(n3583), .dinb(n3582), .dout(n3935));
  jor  g03680(.dina(n3935), .dinb(n3934), .dout(n3936));
  jxor g03681(.dina(b36 ), .dinb(b35 ), .dout(n3937));
  jnot g03682(.din(n3937), .dout(n3938));
  jxor g03683(.dina(n3938), .dinb(n3936), .dout(n3939));
  jor  g03684(.dina(n3939), .dinb(n264), .dout(n3940));
  jor  g03685(.dina(n284), .dinb(n3403), .dout(n3941));
  jnot g03686(.din(b36 ), .dout(n3942));
  jor  g03687(.dina(n269), .dinb(n3942), .dout(n3943));
  jor  g03688(.dina(n271), .dinb(n3588), .dout(n3944));
  jand g03689(.dina(n3944), .dinb(n3943), .dout(n3945));
  jand g03690(.dina(n3945), .dinb(n3941), .dout(n3946));
  jand g03691(.dina(n3946), .dinb(n3940), .dout(n3947));
  jxor g03692(.dina(n3947), .dinb(n260), .dout(n3948));
  jxor g03693(.dina(n3948), .dinb(n3933), .dout(n3949));
  jxor g03694(.dina(n3949), .dinb(n3768), .dout(f36 ));
  jand g03695(.dina(n3948), .dinb(n3933), .dout(n3951));
  jand g03696(.dina(n3949), .dinb(n3768), .dout(n3952));
  jor  g03697(.dina(n3952), .dinb(n3951), .dout(n3953));
  jand g03698(.dina(n3931), .dinb(n3781), .dout(n3954));
  jand g03699(.dina(n3932), .dinb(n3772), .dout(n3955));
  jor  g03700(.dina(n3955), .dinb(n3954), .dout(n3956));
  jand g03701(.dina(n3929), .dinb(n3794), .dout(n3957));
  jand g03702(.dina(n3930), .dinb(n3785), .dout(n3958));
  jor  g03703(.dina(n3958), .dinb(n3957), .dout(n3959));
  jor  g03704(.dina(n3032), .dinb(n528), .dout(n3960));
  jor  g03705(.dina(n490), .dinb(n2579), .dout(n3961));
  jor  g03706(.dina(n531), .dinb(n2870), .dout(n3962));
  jor  g03707(.dina(n533), .dinb(n3035), .dout(n3963));
  jand g03708(.dina(n3963), .dinb(n3962), .dout(n3964));
  jand g03709(.dina(n3964), .dinb(n3961), .dout(n3965));
  jand g03710(.dina(n3965), .dinb(n3960), .dout(n3966));
  jxor g03711(.dina(n3966), .dinb(a8 ), .dout(n3967));
  jnot g03712(.din(n3967), .dout(n3968));
  jnot g03713(.din(n3919), .dout(n3969));
  jor  g03714(.dina(n3927), .dinb(n3969), .dout(n3970));
  jor  g03715(.dina(n3928), .dinb(n3798), .dout(n3971));
  jand g03716(.dina(n3971), .dinb(n3970), .dout(n3972));
  jor  g03717(.dina(n2556), .dinb(n706), .dout(n3973));
  jor  g03718(.dina(n683), .dinb(n2148), .dout(n3974));
  jor  g03719(.dina(n709), .dinb(n2407), .dout(n3975));
  jor  g03720(.dina(n711), .dinb(n2559), .dout(n3976));
  jand g03721(.dina(n3976), .dinb(n3975), .dout(n3977));
  jand g03722(.dina(n3977), .dinb(n3974), .dout(n3978));
  jand g03723(.dina(n3978), .dinb(n3973), .dout(n3979));
  jxor g03724(.dina(n3979), .dinb(a11 ), .dout(n3980));
  jnot g03725(.din(n3980), .dout(n3981));
  jand g03726(.dina(n3917), .dinb(n3810), .dout(n3982));
  jand g03727(.dina(n3918), .dinb(n3801), .dout(n3983));
  jor  g03728(.dina(n3983), .dinb(n3982), .dout(n3984));
  jor  g03729(.dina(n3915), .dinb(n3907), .dout(n3985));
  jnot g03730(.din(n3985), .dout(n3986));
  jand g03731(.dina(n3916), .dinb(n3814), .dout(n3987));
  jor  g03732(.dina(n3987), .dinb(n3986), .dout(n3988));
  jand g03733(.dina(n3904), .dinb(n3828), .dout(n3989));
  jand g03734(.dina(n3905), .dinb(n3819), .dout(n3990));
  jor  g03735(.dina(n3990), .dinb(n3989), .dout(n3991));
  jor  g03736(.dina(n3902), .dinb(n3894), .dout(n3992));
  jand g03737(.dina(n3903), .dinb(n3831), .dout(n3993));
  jnot g03738(.din(n3993), .dout(n3994));
  jand g03739(.dina(n3994), .dinb(n3992), .dout(n3995));
  jnot g03740(.din(n3995), .dout(n3996));
  jor  g03741(.dina(n3888), .dinb(n3880), .dout(n3997));
  jand g03742(.dina(n3892), .dinb(n3889), .dout(n3998));
  jnot g03743(.din(n3998), .dout(n3999));
  jand g03744(.dina(n3999), .dinb(n3997), .dout(n4000));
  jnot g03745(.din(n4000), .dout(n4001));
  jor  g03746(.dina(n2319), .dinb(n775), .dout(n4002));
  jor  g03747(.dina(n2224), .dinb(n647), .dout(n4003));
  jor  g03748(.dina(n2322), .dinb(n758), .dout(n4004));
  jor  g03749(.dina(n2324), .dinb(n778), .dout(n4005));
  jand g03750(.dina(n4005), .dinb(n4004), .dout(n4006));
  jand g03751(.dina(n4006), .dinb(n4003), .dout(n4007));
  jand g03752(.dina(n4007), .dinb(n4002), .dout(n4008));
  jxor g03753(.dina(n4008), .dinb(a26 ), .dout(n4009));
  jnot g03754(.din(n4009), .dout(n4010));
  jand g03755(.dina(n3877), .dinb(n3845), .dout(n4011));
  jand g03756(.dina(n3878), .dinb(n3836), .dout(n4012));
  jor  g03757(.dina(n4012), .dinb(n4011), .dout(n4013));
  jor  g03758(.dina(n2784), .dinb(n624), .dout(n4014));
  jor  g03759(.dina(n2661), .dinb(n512), .dout(n4015));
  jor  g03760(.dina(n2787), .dinb(n564), .dout(n4016));
  jor  g03761(.dina(n2789), .dinb(n627), .dout(n4017));
  jand g03762(.dina(n4017), .dinb(n4016), .dout(n4018));
  jand g03763(.dina(n4018), .dinb(n4015), .dout(n4019));
  jand g03764(.dina(n4019), .dinb(n4014), .dout(n4020));
  jxor g03765(.dina(n4020), .dinb(a29 ), .dout(n4021));
  jnot g03766(.din(n4021), .dout(n4022));
  jor  g03767(.dina(n3875), .dinb(n3867), .dout(n4023));
  jand g03768(.dina(n3876), .dinb(n3848), .dout(n4024));
  jnot g03769(.din(n4024), .dout(n4025));
  jand g03770(.dina(n4025), .dinb(n4023), .dout(n4026));
  jnot g03771(.din(n4026), .dout(n4027));
  jor  g03772(.dina(n3301), .dinb(n428), .dout(n4028));
  jor  g03773(.dina(n3136), .dinb(n357), .dout(n4029));
  jor  g03774(.dina(n3304), .dinb(n395), .dout(n4030));
  jor  g03775(.dina(n3306), .dinb(n431), .dout(n4031));
  jand g03776(.dina(n4031), .dinb(n4030), .dout(n4032));
  jand g03777(.dina(n4032), .dinb(n4029), .dout(n4033));
  jand g03778(.dina(n4033), .dinb(n4028), .dout(n4034));
  jxor g03779(.dina(n4034), .dinb(a32 ), .dout(n4035));
  jnot g03780(.din(n4035), .dout(n4036));
  jnot g03781(.din(n3864), .dout(n4037));
  jand g03782(.dina(n4037), .dinb(n3862), .dout(n4038));
  jand g03783(.dina(n3865), .dinb(n3860), .dout(n4039));
  jor  g03784(.dina(n4039), .dinb(n4038), .dout(n4040));
  jor  g03785(.dina(n3849), .dinb(n319), .dout(n4041));
  jor  g03786(.dina(n3689), .dinb(n279), .dout(n4042));
  jor  g03787(.dina(n3852), .dinb(n299), .dout(n4043));
  jor  g03788(.dina(n3854), .dinb(n322), .dout(n4044));
  jand g03789(.dina(n4044), .dinb(n4043), .dout(n4045));
  jand g03790(.dina(n4045), .dinb(n4042), .dout(n4046));
  jand g03791(.dina(n4046), .dinb(n4041), .dout(n4047));
  jxor g03792(.dina(n4047), .dinb(a35 ), .dout(n4048));
  jnot g03793(.din(n4048), .dout(n4049));
  jand g03794(.dina(n3862), .dinb(a38 ), .dout(n4050));
  jxor g03795(.dina(a38 ), .dinb(a37 ), .dout(n4051));
  jnot g03796(.din(n4051), .dout(n4052));
  jand g03797(.dina(n4052), .dinb(n3861), .dout(n4053));
  jand g03798(.dina(n4053), .dinb(b1 ), .dout(n4054));
  jnot g03799(.din(n3861), .dout(n4055));
  jxor g03800(.dina(a37 ), .dinb(a36 ), .dout(n4056));
  jand g03801(.dina(n4056), .dinb(n4055), .dout(n4057));
  jand g03802(.dina(n4057), .dinb(b0 ), .dout(n4058));
  jand g03803(.dina(n4051), .dinb(n3861), .dout(n4059));
  jand g03804(.dina(n4059), .dinb(n338), .dout(n4060));
  jor  g03805(.dina(n4060), .dinb(n4058), .dout(n4061));
  jor  g03806(.dina(n4061), .dinb(n4054), .dout(n4062));
  jxor g03807(.dina(n4062), .dinb(n4050), .dout(n4063));
  jxor g03808(.dina(n4063), .dinb(n4049), .dout(n4064));
  jxor g03809(.dina(n4064), .dinb(n4040), .dout(n4065));
  jxor g03810(.dina(n4065), .dinb(n4036), .dout(n4066));
  jxor g03811(.dina(n4066), .dinb(n4027), .dout(n4067));
  jxor g03812(.dina(n4067), .dinb(n4022), .dout(n4068));
  jxor g03813(.dina(n4068), .dinb(n4013), .dout(n4069));
  jxor g03814(.dina(n4069), .dinb(n4010), .dout(n4070));
  jxor g03815(.dina(n4070), .dinb(n4001), .dout(n4071));
  jnot g03816(.din(n4071), .dout(n4072));
  jor  g03817(.dina(n1939), .dinb(n1019), .dout(n4073));
  jor  g03818(.dina(n1827), .dinb(n858), .dout(n4074));
  jor  g03819(.dina(n1942), .dinb(n939), .dout(n4075));
  jor  g03820(.dina(n1944), .dinb(n1022), .dout(n4076));
  jand g03821(.dina(n4076), .dinb(n4075), .dout(n4077));
  jand g03822(.dina(n4077), .dinb(n4074), .dout(n4078));
  jand g03823(.dina(n4078), .dinb(n4073), .dout(n4079));
  jxor g03824(.dina(n4079), .dinb(a23 ), .dout(n4080));
  jxor g03825(.dina(n4080), .dinb(n4072), .dout(n4081));
  jxor g03826(.dina(n4081), .dinb(n3996), .dout(n4082));
  jnot g03827(.din(n4082), .dout(n4083));
  jor  g03828(.dina(n1397), .dinb(n1566), .dout(n4084));
  jor  g03829(.dina(n1489), .dinb(n1193), .dout(n4085));
  jor  g03830(.dina(n1569), .dinb(n1290), .dout(n4086));
  jor  g03831(.dina(n1571), .dinb(n1400), .dout(n4087));
  jand g03832(.dina(n4087), .dinb(n4086), .dout(n4088));
  jand g03833(.dina(n4088), .dinb(n4085), .dout(n4089));
  jand g03834(.dina(n4089), .dinb(n4084), .dout(n4090));
  jxor g03835(.dina(n4090), .dinb(a20 ), .dout(n4091));
  jxor g03836(.dina(n4091), .dinb(n4083), .dout(n4092));
  jxor g03837(.dina(n4092), .dinb(n3991), .dout(n4093));
  jnot g03838(.din(n4093), .dout(n4094));
  jor  g03839(.dina(n1739), .dinb(n1245), .dout(n4095));
  jor  g03840(.dina(n1165), .dinb(n1420), .dout(n4096));
  jor  g03841(.dina(n1248), .dinb(n1620), .dout(n4097));
  jor  g03842(.dina(n1250), .dinb(n1742), .dout(n4098));
  jand g03843(.dina(n4098), .dinb(n4097), .dout(n4099));
  jand g03844(.dina(n4099), .dinb(n4096), .dout(n4100));
  jand g03845(.dina(n4100), .dinb(n4095), .dout(n4101));
  jxor g03846(.dina(n4101), .dinb(a17 ), .dout(n4102));
  jxor g03847(.dina(n4102), .dinb(n4094), .dout(n4103));
  jxor g03848(.dina(n4103), .dinb(n3988), .dout(n4104));
  jor  g03849(.dina(n2007), .dinb(n974), .dout(n4105));
  jor  g03850(.dina(n908), .dinb(n1867), .dout(n4106));
  jor  g03851(.dina(n977), .dinb(n1887), .dout(n4107));
  jor  g03852(.dina(n979), .dinb(n2010), .dout(n4108));
  jand g03853(.dina(n4108), .dinb(n4107), .dout(n4109));
  jand g03854(.dina(n4109), .dinb(n4106), .dout(n4110));
  jand g03855(.dina(n4110), .dinb(n4105), .dout(n4111));
  jxor g03856(.dina(n4111), .dinb(a14 ), .dout(n4112));
  jxor g03857(.dina(n4112), .dinb(n4104), .dout(n4113));
  jnot g03858(.din(n4113), .dout(n4114));
  jxor g03859(.dina(n4114), .dinb(n3984), .dout(n4115));
  jxor g03860(.dina(n4115), .dinb(n3981), .dout(n4116));
  jnot g03861(.din(n4116), .dout(n4117));
  jxor g03862(.dina(n4117), .dinb(n3972), .dout(n4118));
  jxor g03863(.dina(n4118), .dinb(n3968), .dout(n4119));
  jnot g03864(.din(n4119), .dout(n4120));
  jxor g03865(.dina(n4120), .dinb(n3959), .dout(n4121));
  jor  g03866(.dina(n3400), .dinb(n402), .dout(n4122));
  jor  g03867(.dina(n371), .dinb(n3055), .dout(n4123));
  jor  g03868(.dina(n405), .dinb(n3230), .dout(n4124));
  jor  g03869(.dina(n332), .dinb(n3403), .dout(n4125));
  jand g03870(.dina(n4125), .dinb(n4124), .dout(n4126));
  jand g03871(.dina(n4126), .dinb(n4123), .dout(n4127));
  jand g03872(.dina(n4127), .dinb(n4122), .dout(n4128));
  jxor g03873(.dina(n4128), .dinb(a5 ), .dout(n4129));
  jxor g03874(.dina(n4129), .dinb(n4121), .dout(n4130));
  jxor g03875(.dina(n4130), .dinb(n3956), .dout(n4131));
  jand g03876(.dina(b36 ), .dinb(b35 ), .dout(n4132));
  jand g03877(.dina(n3937), .dinb(n3936), .dout(n4133));
  jor  g03878(.dina(n4133), .dinb(n4132), .dout(n4134));
  jxor g03879(.dina(b37 ), .dinb(b36 ), .dout(n4135));
  jnot g03880(.din(n4135), .dout(n4136));
  jxor g03881(.dina(n4136), .dinb(n4134), .dout(n4137));
  jor  g03882(.dina(n4137), .dinb(n264), .dout(n4138));
  jor  g03883(.dina(n284), .dinb(n3588), .dout(n4139));
  jnot g03884(.din(b37 ), .dout(n4140));
  jor  g03885(.dina(n269), .dinb(n4140), .dout(n4141));
  jor  g03886(.dina(n271), .dinb(n3942), .dout(n4142));
  jand g03887(.dina(n4142), .dinb(n4141), .dout(n4143));
  jand g03888(.dina(n4143), .dinb(n4139), .dout(n4144));
  jand g03889(.dina(n4144), .dinb(n4138), .dout(n4145));
  jxor g03890(.dina(n4145), .dinb(n260), .dout(n4146));
  jxor g03891(.dina(n4146), .dinb(n4131), .dout(n4147));
  jxor g03892(.dina(n4147), .dinb(n3953), .dout(f37 ));
  jand g03893(.dina(n4146), .dinb(n4131), .dout(n4149));
  jand g03894(.dina(n4147), .dinb(n3953), .dout(n4150));
  jor  g03895(.dina(n4150), .dinb(n4149), .dout(n4151));
  jor  g03896(.dina(n4129), .dinb(n4121), .dout(n4152));
  jnot g03897(.din(n4152), .dout(n4153));
  jand g03898(.dina(n4130), .dinb(n3956), .dout(n4154));
  jor  g03899(.dina(n4154), .dinb(n4153), .dout(n4155));
  jor  g03900(.dina(n3585), .dinb(n402), .dout(n4156));
  jor  g03901(.dina(n371), .dinb(n3230), .dout(n4157));
  jor  g03902(.dina(n405), .dinb(n3403), .dout(n4158));
  jor  g03903(.dina(n332), .dinb(n3588), .dout(n4159));
  jand g03904(.dina(n4159), .dinb(n4158), .dout(n4160));
  jand g03905(.dina(n4160), .dinb(n4157), .dout(n4161));
  jand g03906(.dina(n4161), .dinb(n4156), .dout(n4162));
  jxor g03907(.dina(n4162), .dinb(a5 ), .dout(n4163));
  jnot g03908(.din(n4163), .dout(n4164));
  jand g03909(.dina(n4118), .dinb(n3968), .dout(n4165));
  jand g03910(.dina(n4119), .dinb(n3959), .dout(n4166));
  jor  g03911(.dina(n4166), .dinb(n4165), .dout(n4167));
  jor  g03912(.dina(n3052), .dinb(n528), .dout(n4168));
  jor  g03913(.dina(n490), .dinb(n2870), .dout(n4169));
  jor  g03914(.dina(n531), .dinb(n3035), .dout(n4170));
  jor  g03915(.dina(n533), .dinb(n3055), .dout(n4171));
  jand g03916(.dina(n4171), .dinb(n4170), .dout(n4172));
  jand g03917(.dina(n4172), .dinb(n4169), .dout(n4173));
  jand g03918(.dina(n4173), .dinb(n4168), .dout(n4174));
  jxor g03919(.dina(n4174), .dinb(a8 ), .dout(n4175));
  jnot g03920(.din(n4175), .dout(n4176));
  jand g03921(.dina(n4115), .dinb(n3981), .dout(n4177));
  jnot g03922(.din(n4177), .dout(n4178));
  jor  g03923(.dina(n4117), .dinb(n3972), .dout(n4179));
  jand g03924(.dina(n4179), .dinb(n4178), .dout(n4180));
  jor  g03925(.dina(n2576), .dinb(n706), .dout(n4181));
  jor  g03926(.dina(n683), .dinb(n2407), .dout(n4182));
  jor  g03927(.dina(n709), .dinb(n2559), .dout(n4183));
  jor  g03928(.dina(n711), .dinb(n2579), .dout(n4184));
  jand g03929(.dina(n4184), .dinb(n4183), .dout(n4185));
  jand g03930(.dina(n4185), .dinb(n4182), .dout(n4186));
  jand g03931(.dina(n4186), .dinb(n4181), .dout(n4187));
  jxor g03932(.dina(n4187), .dinb(a11 ), .dout(n4188));
  jnot g03933(.din(n4188), .dout(n4189));
  jnot g03934(.din(n4104), .dout(n4190));
  jor  g03935(.dina(n4112), .dinb(n4190), .dout(n4191));
  jnot g03936(.din(n4191), .dout(n4192));
  jand g03937(.dina(n4114), .dinb(n3984), .dout(n4193));
  jor  g03938(.dina(n4193), .dinb(n4192), .dout(n4194));
  jor  g03939(.dina(n2145), .dinb(n974), .dout(n4195));
  jor  g03940(.dina(n908), .dinb(n1887), .dout(n4196));
  jor  g03941(.dina(n977), .dinb(n2010), .dout(n4197));
  jor  g03942(.dina(n979), .dinb(n2148), .dout(n4198));
  jand g03943(.dina(n4198), .dinb(n4197), .dout(n4199));
  jand g03944(.dina(n4199), .dinb(n4196), .dout(n4200));
  jand g03945(.dina(n4200), .dinb(n4195), .dout(n4201));
  jxor g03946(.dina(n4201), .dinb(a14 ), .dout(n4202));
  jnot g03947(.din(n4202), .dout(n4203));
  jor  g03948(.dina(n4102), .dinb(n4094), .dout(n4204));
  jnot g03949(.din(n4204), .dout(n4205));
  jand g03950(.dina(n4103), .dinb(n3988), .dout(n4206));
  jor  g03951(.dina(n4206), .dinb(n4205), .dout(n4207));
  jor  g03952(.dina(n4091), .dinb(n4083), .dout(n4208));
  jand g03953(.dina(n4092), .dinb(n3991), .dout(n4209));
  jnot g03954(.din(n4209), .dout(n4210));
  jand g03955(.dina(n4210), .dinb(n4208), .dout(n4211));
  jnot g03956(.din(n4211), .dout(n4212));
  jor  g03957(.dina(n4080), .dinb(n4072), .dout(n4213));
  jand g03958(.dina(n4081), .dinb(n3996), .dout(n4214));
  jnot g03959(.din(n4214), .dout(n4215));
  jand g03960(.dina(n4215), .dinb(n4213), .dout(n4216));
  jnot g03961(.din(n4216), .dout(n4217));
  jand g03962(.dina(n4069), .dinb(n4010), .dout(n4218));
  jand g03963(.dina(n4070), .dinb(n4001), .dout(n4219));
  jor  g03964(.dina(n4219), .dinb(n4218), .dout(n4220));
  jor  g03965(.dina(n2319), .dinb(n855), .dout(n4221));
  jor  g03966(.dina(n2224), .dinb(n758), .dout(n4222));
  jor  g03967(.dina(n2322), .dinb(n778), .dout(n4223));
  jor  g03968(.dina(n2324), .dinb(n858), .dout(n4224));
  jand g03969(.dina(n4224), .dinb(n4223), .dout(n4225));
  jand g03970(.dina(n4225), .dinb(n4222), .dout(n4226));
  jand g03971(.dina(n4226), .dinb(n4221), .dout(n4227));
  jxor g03972(.dina(n4227), .dinb(a26 ), .dout(n4228));
  jnot g03973(.din(n4228), .dout(n4229));
  jand g03974(.dina(n4067), .dinb(n4022), .dout(n4230));
  jand g03975(.dina(n4068), .dinb(n4013), .dout(n4231));
  jor  g03976(.dina(n4231), .dinb(n4230), .dout(n4232));
  jor  g03977(.dina(n2784), .dinb(n644), .dout(n4233));
  jor  g03978(.dina(n2661), .dinb(n564), .dout(n4234));
  jor  g03979(.dina(n2787), .dinb(n627), .dout(n4235));
  jor  g03980(.dina(n2789), .dinb(n647), .dout(n4236));
  jand g03981(.dina(n4236), .dinb(n4235), .dout(n4237));
  jand g03982(.dina(n4237), .dinb(n4234), .dout(n4238));
  jand g03983(.dina(n4238), .dinb(n4233), .dout(n4239));
  jxor g03984(.dina(n4239), .dinb(a29 ), .dout(n4240));
  jnot g03985(.din(n4240), .dout(n4241));
  jand g03986(.dina(n4065), .dinb(n4036), .dout(n4242));
  jand g03987(.dina(n4066), .dinb(n4027), .dout(n4243));
  jor  g03988(.dina(n4243), .dinb(n4242), .dout(n4244));
  jor  g03989(.dina(n3301), .dinb(n509), .dout(n4245));
  jor  g03990(.dina(n3136), .dinb(n395), .dout(n4246));
  jor  g03991(.dina(n3304), .dinb(n431), .dout(n4247));
  jor  g03992(.dina(n3306), .dinb(n512), .dout(n4248));
  jand g03993(.dina(n4248), .dinb(n4247), .dout(n4249));
  jand g03994(.dina(n4249), .dinb(n4246), .dout(n4250));
  jand g03995(.dina(n4250), .dinb(n4245), .dout(n4251));
  jxor g03996(.dina(n4251), .dinb(a32 ), .dout(n4252));
  jnot g03997(.din(n4252), .dout(n4253));
  jand g03998(.dina(n4063), .dinb(n4049), .dout(n4254));
  jand g03999(.dina(n4064), .dinb(n4040), .dout(n4255));
  jor  g04000(.dina(n4255), .dinb(n4254), .dout(n4256));
  jor  g04001(.dina(n3849), .dinb(n354), .dout(n4257));
  jor  g04002(.dina(n3689), .dinb(n299), .dout(n4258));
  jor  g04003(.dina(n3852), .dinb(n322), .dout(n4259));
  jor  g04004(.dina(n3854), .dinb(n357), .dout(n4260));
  jand g04005(.dina(n4260), .dinb(n4259), .dout(n4261));
  jand g04006(.dina(n4261), .dinb(n4258), .dout(n4262));
  jand g04007(.dina(n4262), .dinb(n4257), .dout(n4263));
  jxor g04008(.dina(n4263), .dinb(a35 ), .dout(n4264));
  jnot g04009(.din(n4264), .dout(n4265));
  jnot g04010(.din(n4062), .dout(n4266));
  jand g04011(.dina(n3863), .dinb(a38 ), .dout(n4267));
  jand g04012(.dina(n4267), .dinb(n4266), .dout(n4268));
  jnot g04013(.din(n4268), .dout(n4269));
  jand g04014(.dina(n4269), .dinb(a38 ), .dout(n4270));
  jor  g04015(.dina(n4056), .dinb(n4052), .dout(n4271));
  jor  g04016(.dina(n4271), .dinb(n3861), .dout(n4272));
  jnot g04017(.din(n4272), .dout(n4273));
  jand g04018(.dina(n4273), .dinb(b0 ), .dout(n4274));
  jand g04019(.dina(n4053), .dinb(b2 ), .dout(n4275));
  jand g04020(.dina(n4057), .dinb(b1 ), .dout(n4276));
  jand g04021(.dina(n4059), .dinb(n375), .dout(n4277));
  jor  g04022(.dina(n4277), .dinb(n4276), .dout(n4278));
  jor  g04023(.dina(n4278), .dinb(n4275), .dout(n4279));
  jor  g04024(.dina(n4279), .dinb(n4274), .dout(n4280));
  jxor g04025(.dina(n4280), .dinb(n4270), .dout(n4281));
  jxor g04026(.dina(n4281), .dinb(n4265), .dout(n4282));
  jxor g04027(.dina(n4282), .dinb(n4256), .dout(n4283));
  jxor g04028(.dina(n4283), .dinb(n4253), .dout(n4284));
  jxor g04029(.dina(n4284), .dinb(n4244), .dout(n4285));
  jxor g04030(.dina(n4285), .dinb(n4241), .dout(n4286));
  jxor g04031(.dina(n4286), .dinb(n4232), .dout(n4287));
  jxor g04032(.dina(n4287), .dinb(n4229), .dout(n4288));
  jxor g04033(.dina(n4288), .dinb(n4220), .dout(n4289));
  jnot g04034(.din(n4289), .dout(n4290));
  jor  g04035(.dina(n1939), .dinb(n1190), .dout(n4291));
  jor  g04036(.dina(n1827), .dinb(n939), .dout(n4292));
  jor  g04037(.dina(n1942), .dinb(n1022), .dout(n4293));
  jor  g04038(.dina(n1944), .dinb(n1193), .dout(n4294));
  jand g04039(.dina(n4294), .dinb(n4293), .dout(n4295));
  jand g04040(.dina(n4295), .dinb(n4292), .dout(n4296));
  jand g04041(.dina(n4296), .dinb(n4291), .dout(n4297));
  jxor g04042(.dina(n4297), .dinb(a23 ), .dout(n4298));
  jxor g04043(.dina(n4298), .dinb(n4290), .dout(n4299));
  jxor g04044(.dina(n4299), .dinb(n4217), .dout(n4300));
  jnot g04045(.din(n4300), .dout(n4301));
  jor  g04046(.dina(n1417), .dinb(n1566), .dout(n4302));
  jor  g04047(.dina(n1489), .dinb(n1290), .dout(n4303));
  jor  g04048(.dina(n1569), .dinb(n1400), .dout(n4304));
  jor  g04049(.dina(n1571), .dinb(n1420), .dout(n4305));
  jand g04050(.dina(n4305), .dinb(n4304), .dout(n4306));
  jand g04051(.dina(n4306), .dinb(n4303), .dout(n4307));
  jand g04052(.dina(n4307), .dinb(n4302), .dout(n4308));
  jxor g04053(.dina(n4308), .dinb(a20 ), .dout(n4309));
  jxor g04054(.dina(n4309), .dinb(n4301), .dout(n4310));
  jxor g04055(.dina(n4310), .dinb(n4212), .dout(n4311));
  jnot g04056(.din(n4311), .dout(n4312));
  jor  g04057(.dina(n1864), .dinb(n1245), .dout(n4313));
  jor  g04058(.dina(n1165), .dinb(n1620), .dout(n4314));
  jor  g04059(.dina(n1248), .dinb(n1742), .dout(n4315));
  jor  g04060(.dina(n1250), .dinb(n1867), .dout(n4316));
  jand g04061(.dina(n4316), .dinb(n4315), .dout(n4317));
  jand g04062(.dina(n4317), .dinb(n4314), .dout(n4318));
  jand g04063(.dina(n4318), .dinb(n4313), .dout(n4319));
  jxor g04064(.dina(n4319), .dinb(a17 ), .dout(n4320));
  jxor g04065(.dina(n4320), .dinb(n4312), .dout(n4321));
  jxor g04066(.dina(n4321), .dinb(n4207), .dout(n4322));
  jxor g04067(.dina(n4322), .dinb(n4203), .dout(n4323));
  jxor g04068(.dina(n4323), .dinb(n4194), .dout(n4324));
  jxor g04069(.dina(n4324), .dinb(n4189), .dout(n4325));
  jnot g04070(.din(n4325), .dout(n4326));
  jxor g04071(.dina(n4326), .dinb(n4180), .dout(n4327));
  jxor g04072(.dina(n4327), .dinb(n4176), .dout(n4328));
  jxor g04073(.dina(n4328), .dinb(n4167), .dout(n4329));
  jxor g04074(.dina(n4329), .dinb(n4164), .dout(n4330));
  jxor g04075(.dina(n4330), .dinb(n4155), .dout(n4331));
  jand g04076(.dina(b37 ), .dinb(b36 ), .dout(n4332));
  jand g04077(.dina(n4135), .dinb(n4134), .dout(n4333));
  jor  g04078(.dina(n4333), .dinb(n4332), .dout(n4334));
  jxor g04079(.dina(b38 ), .dinb(b37 ), .dout(n4335));
  jnot g04080(.din(n4335), .dout(n4336));
  jxor g04081(.dina(n4336), .dinb(n4334), .dout(n4337));
  jor  g04082(.dina(n4337), .dinb(n264), .dout(n4338));
  jor  g04083(.dina(n284), .dinb(n3942), .dout(n4339));
  jnot g04084(.din(b38 ), .dout(n4340));
  jor  g04085(.dina(n269), .dinb(n4340), .dout(n4341));
  jor  g04086(.dina(n271), .dinb(n4140), .dout(n4342));
  jand g04087(.dina(n4342), .dinb(n4341), .dout(n4343));
  jand g04088(.dina(n4343), .dinb(n4339), .dout(n4344));
  jand g04089(.dina(n4344), .dinb(n4338), .dout(n4345));
  jxor g04090(.dina(n4345), .dinb(n260), .dout(n4346));
  jxor g04091(.dina(n4346), .dinb(n4331), .dout(n4347));
  jxor g04092(.dina(n4347), .dinb(n4151), .dout(f38 ));
  jand g04093(.dina(n4346), .dinb(n4331), .dout(n4349));
  jand g04094(.dina(n4347), .dinb(n4151), .dout(n4350));
  jor  g04095(.dina(n4350), .dinb(n4349), .dout(n4351));
  jand g04096(.dina(n4329), .dinb(n4164), .dout(n4352));
  jand g04097(.dina(n4330), .dinb(n4155), .dout(n4353));
  jor  g04098(.dina(n4353), .dinb(n4352), .dout(n4354));
  jor  g04099(.dina(n3939), .dinb(n402), .dout(n4355));
  jor  g04100(.dina(n371), .dinb(n3403), .dout(n4356));
  jor  g04101(.dina(n405), .dinb(n3588), .dout(n4357));
  jor  g04102(.dina(n332), .dinb(n3942), .dout(n4358));
  jand g04103(.dina(n4358), .dinb(n4357), .dout(n4359));
  jand g04104(.dina(n4359), .dinb(n4356), .dout(n4360));
  jand g04105(.dina(n4360), .dinb(n4355), .dout(n4361));
  jxor g04106(.dina(n4361), .dinb(a5 ), .dout(n4362));
  jnot g04107(.din(n4362), .dout(n4363));
  jand g04108(.dina(n4327), .dinb(n4176), .dout(n4364));
  jand g04109(.dina(n4328), .dinb(n4167), .dout(n4365));
  jor  g04110(.dina(n4365), .dinb(n4364), .dout(n4366));
  jand g04111(.dina(n4324), .dinb(n4189), .dout(n4367));
  jnot g04112(.din(n4367), .dout(n4368));
  jor  g04113(.dina(n4326), .dinb(n4180), .dout(n4369));
  jand g04114(.dina(n4369), .dinb(n4368), .dout(n4370));
  jor  g04115(.dina(n2867), .dinb(n706), .dout(n4371));
  jor  g04116(.dina(n683), .dinb(n2559), .dout(n4372));
  jor  g04117(.dina(n709), .dinb(n2579), .dout(n4373));
  jor  g04118(.dina(n711), .dinb(n2870), .dout(n4374));
  jand g04119(.dina(n4374), .dinb(n4373), .dout(n4375));
  jand g04120(.dina(n4375), .dinb(n4372), .dout(n4376));
  jand g04121(.dina(n4376), .dinb(n4371), .dout(n4377));
  jxor g04122(.dina(n4377), .dinb(a11 ), .dout(n4378));
  jnot g04123(.din(n4378), .dout(n4379));
  jand g04124(.dina(n4322), .dinb(n4203), .dout(n4380));
  jand g04125(.dina(n4323), .dinb(n4194), .dout(n4381));
  jor  g04126(.dina(n4381), .dinb(n4380), .dout(n4382));
  jor  g04127(.dina(n4320), .dinb(n4312), .dout(n4383));
  jnot g04128(.din(n4383), .dout(n4384));
  jand g04129(.dina(n4321), .dinb(n4207), .dout(n4385));
  jor  g04130(.dina(n4385), .dinb(n4384), .dout(n4386));
  jor  g04131(.dina(n4309), .dinb(n4301), .dout(n4387));
  jand g04132(.dina(n4310), .dinb(n4212), .dout(n4388));
  jnot g04133(.din(n4388), .dout(n4389));
  jand g04134(.dina(n4389), .dinb(n4387), .dout(n4390));
  jnot g04135(.din(n4390), .dout(n4391));
  jor  g04136(.dina(n4298), .dinb(n4290), .dout(n4392));
  jand g04137(.dina(n4299), .dinb(n4217), .dout(n4393));
  jnot g04138(.din(n4393), .dout(n4394));
  jand g04139(.dina(n4394), .dinb(n4392), .dout(n4395));
  jnot g04140(.din(n4395), .dout(n4396));
  jor  g04141(.dina(n1939), .dinb(n1287), .dout(n4397));
  jor  g04142(.dina(n1827), .dinb(n1022), .dout(n4398));
  jor  g04143(.dina(n1942), .dinb(n1193), .dout(n4399));
  jor  g04144(.dina(n1944), .dinb(n1290), .dout(n4400));
  jand g04145(.dina(n4400), .dinb(n4399), .dout(n4401));
  jand g04146(.dina(n4401), .dinb(n4398), .dout(n4402));
  jand g04147(.dina(n4402), .dinb(n4397), .dout(n4403));
  jxor g04148(.dina(n4403), .dinb(a23 ), .dout(n4404));
  jnot g04149(.din(n4404), .dout(n4405));
  jand g04150(.dina(n4287), .dinb(n4229), .dout(n4406));
  jand g04151(.dina(n4288), .dinb(n4220), .dout(n4407));
  jor  g04152(.dina(n4407), .dinb(n4406), .dout(n4408));
  jand g04153(.dina(n4283), .dinb(n4253), .dout(n4409));
  jand g04154(.dina(n4284), .dinb(n4244), .dout(n4410));
  jor  g04155(.dina(n4410), .dinb(n4409), .dout(n4411));
  jand g04156(.dina(n4281), .dinb(n4265), .dout(n4412));
  jand g04157(.dina(n4282), .dinb(n4256), .dout(n4413));
  jor  g04158(.dina(n4413), .dinb(n4412), .dout(n4414));
  jnot g04159(.din(n4059), .dout(n4415));
  jor  g04160(.dina(n4415), .dinb(n296), .dout(n4416));
  jor  g04161(.dina(n4272), .dinb(n267), .dout(n4417));
  jnot g04162(.din(n4057), .dout(n4418));
  jor  g04163(.dina(n4418), .dinb(n279), .dout(n4419));
  jnot g04164(.din(n4053), .dout(n4420));
  jor  g04165(.dina(n4420), .dinb(n299), .dout(n4421));
  jand g04166(.dina(n4421), .dinb(n4419), .dout(n4422));
  jand g04167(.dina(n4422), .dinb(n4417), .dout(n4423));
  jand g04168(.dina(n4423), .dinb(n4416), .dout(n4424));
  jxor g04169(.dina(n4424), .dinb(a38 ), .dout(n4425));
  jnot g04170(.din(n4425), .dout(n4426));
  jxor g04171(.dina(a39 ), .dinb(a38 ), .dout(n4427));
  jand g04172(.dina(n4427), .dinb(b0 ), .dout(n4428));
  jnot g04173(.din(n4428), .dout(n4429));
  jor  g04174(.dina(n4280), .dinb(n4269), .dout(n4430));
  jxor g04175(.dina(n4430), .dinb(n4429), .dout(n4431));
  jxor g04176(.dina(n4431), .dinb(n4426), .dout(n4432));
  jnot g04177(.din(n4432), .dout(n4433));
  jor  g04178(.dina(n3849), .dinb(n392), .dout(n4434));
  jor  g04179(.dina(n3689), .dinb(n322), .dout(n4435));
  jor  g04180(.dina(n3852), .dinb(n357), .dout(n4436));
  jor  g04181(.dina(n3854), .dinb(n395), .dout(n4437));
  jand g04182(.dina(n4437), .dinb(n4436), .dout(n4438));
  jand g04183(.dina(n4438), .dinb(n4435), .dout(n4439));
  jand g04184(.dina(n4439), .dinb(n4434), .dout(n4440));
  jxor g04185(.dina(n4440), .dinb(a35 ), .dout(n4441));
  jxor g04186(.dina(n4441), .dinb(n4433), .dout(n4442));
  jxor g04187(.dina(n4442), .dinb(n4414), .dout(n4443));
  jnot g04188(.din(n4443), .dout(n4444));
  jor  g04189(.dina(n3301), .dinb(n561), .dout(n4445));
  jor  g04190(.dina(n3136), .dinb(n431), .dout(n4446));
  jor  g04191(.dina(n3304), .dinb(n512), .dout(n4447));
  jor  g04192(.dina(n3306), .dinb(n564), .dout(n4448));
  jand g04193(.dina(n4448), .dinb(n4447), .dout(n4449));
  jand g04194(.dina(n4449), .dinb(n4446), .dout(n4450));
  jand g04195(.dina(n4450), .dinb(n4445), .dout(n4451));
  jxor g04196(.dina(n4451), .dinb(a32 ), .dout(n4452));
  jxor g04197(.dina(n4452), .dinb(n4444), .dout(n4453));
  jxor g04198(.dina(n4453), .dinb(n4411), .dout(n4454));
  jnot g04199(.din(n4454), .dout(n4455));
  jor  g04200(.dina(n2784), .dinb(n755), .dout(n4456));
  jor  g04201(.dina(n2661), .dinb(n627), .dout(n4457));
  jor  g04202(.dina(n2787), .dinb(n647), .dout(n4458));
  jor  g04203(.dina(n2789), .dinb(n758), .dout(n4459));
  jand g04204(.dina(n4459), .dinb(n4458), .dout(n4460));
  jand g04205(.dina(n4460), .dinb(n4457), .dout(n4461));
  jand g04206(.dina(n4461), .dinb(n4456), .dout(n4462));
  jxor g04207(.dina(n4462), .dinb(a29 ), .dout(n4463));
  jxor g04208(.dina(n4463), .dinb(n4455), .dout(n4464));
  jand g04209(.dina(n4285), .dinb(n4241), .dout(n4465));
  jand g04210(.dina(n4286), .dinb(n4232), .dout(n4466));
  jor  g04211(.dina(n4466), .dinb(n4465), .dout(n4467));
  jxor g04212(.dina(n4467), .dinb(n4464), .dout(n4468));
  jnot g04213(.din(n4468), .dout(n4469));
  jor  g04214(.dina(n2319), .dinb(n936), .dout(n4470));
  jor  g04215(.dina(n2224), .dinb(n778), .dout(n4471));
  jor  g04216(.dina(n2322), .dinb(n858), .dout(n4472));
  jor  g04217(.dina(n2324), .dinb(n939), .dout(n4473));
  jand g04218(.dina(n4473), .dinb(n4472), .dout(n4474));
  jand g04219(.dina(n4474), .dinb(n4471), .dout(n4475));
  jand g04220(.dina(n4475), .dinb(n4470), .dout(n4476));
  jxor g04221(.dina(n4476), .dinb(a26 ), .dout(n4477));
  jxor g04222(.dina(n4477), .dinb(n4469), .dout(n4478));
  jxor g04223(.dina(n4478), .dinb(n4408), .dout(n4479));
  jxor g04224(.dina(n4479), .dinb(n4405), .dout(n4480));
  jxor g04225(.dina(n4480), .dinb(n4396), .dout(n4481));
  jnot g04226(.din(n4481), .dout(n4482));
  jor  g04227(.dina(n1617), .dinb(n1566), .dout(n4483));
  jor  g04228(.dina(n1489), .dinb(n1400), .dout(n4484));
  jor  g04229(.dina(n1569), .dinb(n1420), .dout(n4485));
  jor  g04230(.dina(n1571), .dinb(n1620), .dout(n4486));
  jand g04231(.dina(n4486), .dinb(n4485), .dout(n4487));
  jand g04232(.dina(n4487), .dinb(n4484), .dout(n4488));
  jand g04233(.dina(n4488), .dinb(n4483), .dout(n4489));
  jxor g04234(.dina(n4489), .dinb(a20 ), .dout(n4490));
  jxor g04235(.dina(n4490), .dinb(n4482), .dout(n4491));
  jxor g04236(.dina(n4491), .dinb(n4391), .dout(n4492));
  jor  g04237(.dina(n1884), .dinb(n1245), .dout(n4493));
  jor  g04238(.dina(n1165), .dinb(n1742), .dout(n4494));
  jor  g04239(.dina(n1248), .dinb(n1867), .dout(n4495));
  jor  g04240(.dina(n1250), .dinb(n1887), .dout(n4496));
  jand g04241(.dina(n4496), .dinb(n4495), .dout(n4497));
  jand g04242(.dina(n4497), .dinb(n4494), .dout(n4498));
  jand g04243(.dina(n4498), .dinb(n4493), .dout(n4499));
  jxor g04244(.dina(n4499), .dinb(a17 ), .dout(n4500));
  jxor g04245(.dina(n4500), .dinb(n4492), .dout(n4501));
  jxor g04246(.dina(n4501), .dinb(n4386), .dout(n4502));
  jor  g04247(.dina(n2404), .dinb(n974), .dout(n4503));
  jor  g04248(.dina(n908), .dinb(n2010), .dout(n4504));
  jor  g04249(.dina(n977), .dinb(n2148), .dout(n4505));
  jor  g04250(.dina(n979), .dinb(n2407), .dout(n4506));
  jand g04251(.dina(n4506), .dinb(n4505), .dout(n4507));
  jand g04252(.dina(n4507), .dinb(n4504), .dout(n4508));
  jand g04253(.dina(n4508), .dinb(n4503), .dout(n4509));
  jxor g04254(.dina(n4509), .dinb(a14 ), .dout(n4510));
  jxor g04255(.dina(n4510), .dinb(n4502), .dout(n4511));
  jxor g04256(.dina(n4511), .dinb(n4382), .dout(n4512));
  jxor g04257(.dina(n4512), .dinb(n4379), .dout(n4513));
  jnot g04258(.din(n4513), .dout(n4514));
  jxor g04259(.dina(n4514), .dinb(n4370), .dout(n4515));
  jnot g04260(.din(n4515), .dout(n4516));
  jor  g04261(.dina(n3227), .dinb(n528), .dout(n4517));
  jor  g04262(.dina(n490), .dinb(n3035), .dout(n4518));
  jor  g04263(.dina(n531), .dinb(n3055), .dout(n4519));
  jor  g04264(.dina(n533), .dinb(n3230), .dout(n4520));
  jand g04265(.dina(n4520), .dinb(n4519), .dout(n4521));
  jand g04266(.dina(n4521), .dinb(n4518), .dout(n4522));
  jand g04267(.dina(n4522), .dinb(n4517), .dout(n4523));
  jxor g04268(.dina(n4523), .dinb(a8 ), .dout(n4524));
  jxor g04269(.dina(n4524), .dinb(n4516), .dout(n4525));
  jxor g04270(.dina(n4525), .dinb(n4366), .dout(n4526));
  jxor g04271(.dina(n4526), .dinb(n4363), .dout(n4527));
  jxor g04272(.dina(n4527), .dinb(n4354), .dout(n4528));
  jand g04273(.dina(b38 ), .dinb(b37 ), .dout(n4529));
  jand g04274(.dina(n4335), .dinb(n4334), .dout(n4530));
  jor  g04275(.dina(n4530), .dinb(n4529), .dout(n4531));
  jxor g04276(.dina(b39 ), .dinb(b38 ), .dout(n4532));
  jnot g04277(.din(n4532), .dout(n4533));
  jxor g04278(.dina(n4533), .dinb(n4531), .dout(n4534));
  jor  g04279(.dina(n4534), .dinb(n264), .dout(n4535));
  jor  g04280(.dina(n284), .dinb(n4140), .dout(n4536));
  jnot g04281(.din(b39 ), .dout(n4537));
  jor  g04282(.dina(n269), .dinb(n4537), .dout(n4538));
  jor  g04283(.dina(n271), .dinb(n4340), .dout(n4539));
  jand g04284(.dina(n4539), .dinb(n4538), .dout(n4540));
  jand g04285(.dina(n4540), .dinb(n4536), .dout(n4541));
  jand g04286(.dina(n4541), .dinb(n4535), .dout(n4542));
  jxor g04287(.dina(n4542), .dinb(n260), .dout(n4543));
  jxor g04288(.dina(n4543), .dinb(n4528), .dout(n4544));
  jxor g04289(.dina(n4544), .dinb(n4351), .dout(f39 ));
  jand g04290(.dina(n4543), .dinb(n4528), .dout(n4546));
  jand g04291(.dina(n4544), .dinb(n4351), .dout(n4547));
  jor  g04292(.dina(n4547), .dinb(n4546), .dout(n4548));
  jand g04293(.dina(b39 ), .dinb(b38 ), .dout(n4549));
  jand g04294(.dina(n4532), .dinb(n4531), .dout(n4550));
  jor  g04295(.dina(n4550), .dinb(n4549), .dout(n4551));
  jxor g04296(.dina(b40 ), .dinb(b39 ), .dout(n4552));
  jnot g04297(.din(n4552), .dout(n4553));
  jxor g04298(.dina(n4553), .dinb(n4551), .dout(n4554));
  jor  g04299(.dina(n4554), .dinb(n264), .dout(n4555));
  jor  g04300(.dina(n284), .dinb(n4340), .dout(n4556));
  jnot g04301(.din(b40 ), .dout(n4557));
  jor  g04302(.dina(n269), .dinb(n4557), .dout(n4558));
  jor  g04303(.dina(n271), .dinb(n4537), .dout(n4559));
  jand g04304(.dina(n4559), .dinb(n4558), .dout(n4560));
  jand g04305(.dina(n4560), .dinb(n4556), .dout(n4561));
  jand g04306(.dina(n4561), .dinb(n4555), .dout(n4562));
  jxor g04307(.dina(n4562), .dinb(n260), .dout(n4563));
  jand g04308(.dina(n4526), .dinb(n4363), .dout(n4564));
  jand g04309(.dina(n4527), .dinb(n4354), .dout(n4565));
  jor  g04310(.dina(n4565), .dinb(n4564), .dout(n4566));
  jor  g04311(.dina(n4524), .dinb(n4516), .dout(n4567));
  jnot g04312(.din(n4567), .dout(n4568));
  jand g04313(.dina(n4525), .dinb(n4366), .dout(n4569));
  jor  g04314(.dina(n4569), .dinb(n4568), .dout(n4570));
  jor  g04315(.dina(n3400), .dinb(n528), .dout(n4571));
  jor  g04316(.dina(n490), .dinb(n3055), .dout(n4572));
  jor  g04317(.dina(n531), .dinb(n3230), .dout(n4573));
  jor  g04318(.dina(n533), .dinb(n3403), .dout(n4574));
  jand g04319(.dina(n4574), .dinb(n4573), .dout(n4575));
  jand g04320(.dina(n4575), .dinb(n4572), .dout(n4576));
  jand g04321(.dina(n4576), .dinb(n4571), .dout(n4577));
  jxor g04322(.dina(n4577), .dinb(a8 ), .dout(n4578));
  jnot g04323(.din(n4578), .dout(n4579));
  jand g04324(.dina(n4512), .dinb(n4379), .dout(n4580));
  jnot g04325(.din(n4580), .dout(n4581));
  jor  g04326(.dina(n4514), .dinb(n4370), .dout(n4582));
  jand g04327(.dina(n4582), .dinb(n4581), .dout(n4583));
  jor  g04328(.dina(n3032), .dinb(n706), .dout(n4584));
  jor  g04329(.dina(n683), .dinb(n2579), .dout(n4585));
  jor  g04330(.dina(n709), .dinb(n2870), .dout(n4586));
  jor  g04331(.dina(n711), .dinb(n3035), .dout(n4587));
  jand g04332(.dina(n4587), .dinb(n4586), .dout(n4588));
  jand g04333(.dina(n4588), .dinb(n4585), .dout(n4589));
  jand g04334(.dina(n4589), .dinb(n4584), .dout(n4590));
  jxor g04335(.dina(n4590), .dinb(a11 ), .dout(n4591));
  jnot g04336(.din(n4591), .dout(n4592));
  jor  g04337(.dina(n4510), .dinb(n4502), .dout(n4593));
  jnot g04338(.din(n4593), .dout(n4594));
  jand g04339(.dina(n4511), .dinb(n4382), .dout(n4595));
  jor  g04340(.dina(n4595), .dinb(n4594), .dout(n4596));
  jor  g04341(.dina(n2556), .dinb(n974), .dout(n4597));
  jor  g04342(.dina(n908), .dinb(n2148), .dout(n4598));
  jor  g04343(.dina(n977), .dinb(n2407), .dout(n4599));
  jor  g04344(.dina(n979), .dinb(n2559), .dout(n4600));
  jand g04345(.dina(n4600), .dinb(n4599), .dout(n4601));
  jand g04346(.dina(n4601), .dinb(n4598), .dout(n4602));
  jand g04347(.dina(n4602), .dinb(n4597), .dout(n4603));
  jxor g04348(.dina(n4603), .dinb(a14 ), .dout(n4604));
  jnot g04349(.din(n4604), .dout(n4605));
  jnot g04350(.din(n4492), .dout(n4606));
  jor  g04351(.dina(n4500), .dinb(n4606), .dout(n4607));
  jnot g04352(.din(n4607), .dout(n4608));
  jnot g04353(.din(n4501), .dout(n4609));
  jand g04354(.dina(n4609), .dinb(n4386), .dout(n4610));
  jor  g04355(.dina(n4610), .dinb(n4608), .dout(n4611));
  jor  g04356(.dina(n4490), .dinb(n4482), .dout(n4612));
  jnot g04357(.din(n4612), .dout(n4613));
  jand g04358(.dina(n4491), .dinb(n4391), .dout(n4614));
  jor  g04359(.dina(n4614), .dinb(n4613), .dout(n4615));
  jand g04360(.dina(n4479), .dinb(n4405), .dout(n4616));
  jand g04361(.dina(n4480), .dinb(n4396), .dout(n4617));
  jor  g04362(.dina(n4617), .dinb(n4616), .dout(n4618));
  jor  g04363(.dina(n4477), .dinb(n4469), .dout(n4619));
  jand g04364(.dina(n4478), .dinb(n4408), .dout(n4620));
  jnot g04365(.din(n4620), .dout(n4621));
  jand g04366(.dina(n4621), .dinb(n4619), .dout(n4622));
  jnot g04367(.din(n4622), .dout(n4623));
  jor  g04368(.dina(n4463), .dinb(n4455), .dout(n4624));
  jand g04369(.dina(n4467), .dinb(n4464), .dout(n4625));
  jnot g04370(.din(n4625), .dout(n4626));
  jand g04371(.dina(n4626), .dinb(n4624), .dout(n4627));
  jnot g04372(.din(n4627), .dout(n4628));
  jor  g04373(.dina(n2784), .dinb(n775), .dout(n4629));
  jor  g04374(.dina(n2661), .dinb(n647), .dout(n4630));
  jor  g04375(.dina(n2787), .dinb(n758), .dout(n4631));
  jor  g04376(.dina(n2789), .dinb(n778), .dout(n4632));
  jand g04377(.dina(n4632), .dinb(n4631), .dout(n4633));
  jand g04378(.dina(n4633), .dinb(n4630), .dout(n4634));
  jand g04379(.dina(n4634), .dinb(n4629), .dout(n4635));
  jxor g04380(.dina(n4635), .dinb(a29 ), .dout(n4636));
  jnot g04381(.din(n4636), .dout(n4637));
  jor  g04382(.dina(n4452), .dinb(n4444), .dout(n4638));
  jand g04383(.dina(n4453), .dinb(n4411), .dout(n4639));
  jnot g04384(.din(n4639), .dout(n4640));
  jand g04385(.dina(n4640), .dinb(n4638), .dout(n4641));
  jnot g04386(.din(n4641), .dout(n4642));
  jor  g04387(.dina(n4441), .dinb(n4433), .dout(n4643));
  jand g04388(.dina(n4442), .dinb(n4414), .dout(n4644));
  jnot g04389(.din(n4644), .dout(n4645));
  jand g04390(.dina(n4645), .dinb(n4643), .dout(n4646));
  jnot g04391(.din(n4646), .dout(n4647));
  jnot g04392(.din(n4430), .dout(n4648));
  jand g04393(.dina(n4648), .dinb(n4428), .dout(n4649));
  jand g04394(.dina(n4431), .dinb(n4426), .dout(n4650));
  jor  g04395(.dina(n4650), .dinb(n4649), .dout(n4651));
  jor  g04396(.dina(n4415), .dinb(n319), .dout(n4652));
  jor  g04397(.dina(n4272), .dinb(n279), .dout(n4653));
  jor  g04398(.dina(n4418), .dinb(n299), .dout(n4654));
  jor  g04399(.dina(n4420), .dinb(n322), .dout(n4655));
  jand g04400(.dina(n4655), .dinb(n4654), .dout(n4656));
  jand g04401(.dina(n4656), .dinb(n4653), .dout(n4657));
  jand g04402(.dina(n4657), .dinb(n4652), .dout(n4658));
  jxor g04403(.dina(n4658), .dinb(a38 ), .dout(n4659));
  jnot g04404(.din(n4659), .dout(n4660));
  jand g04405(.dina(n4428), .dinb(a41 ), .dout(n4661));
  jxor g04406(.dina(a41 ), .dinb(a40 ), .dout(n4662));
  jnot g04407(.din(n4662), .dout(n4663));
  jand g04408(.dina(n4663), .dinb(n4427), .dout(n4664));
  jand g04409(.dina(n4664), .dinb(b1 ), .dout(n4665));
  jnot g04410(.din(n4427), .dout(n4666));
  jxor g04411(.dina(a40 ), .dinb(a39 ), .dout(n4667));
  jand g04412(.dina(n4667), .dinb(n4666), .dout(n4668));
  jand g04413(.dina(n4668), .dinb(b0 ), .dout(n4669));
  jand g04414(.dina(n4662), .dinb(n4427), .dout(n4670));
  jand g04415(.dina(n4670), .dinb(n338), .dout(n4671));
  jor  g04416(.dina(n4671), .dinb(n4669), .dout(n4672));
  jor  g04417(.dina(n4672), .dinb(n4665), .dout(n4673));
  jxor g04418(.dina(n4673), .dinb(n4661), .dout(n4674));
  jxor g04419(.dina(n4674), .dinb(n4660), .dout(n4675));
  jxor g04420(.dina(n4675), .dinb(n4651), .dout(n4676));
  jnot g04421(.din(n4676), .dout(n4677));
  jor  g04422(.dina(n3849), .dinb(n428), .dout(n4678));
  jor  g04423(.dina(n3689), .dinb(n357), .dout(n4679));
  jor  g04424(.dina(n3852), .dinb(n395), .dout(n4680));
  jor  g04425(.dina(n3854), .dinb(n431), .dout(n4681));
  jand g04426(.dina(n4681), .dinb(n4680), .dout(n4682));
  jand g04427(.dina(n4682), .dinb(n4679), .dout(n4683));
  jand g04428(.dina(n4683), .dinb(n4678), .dout(n4684));
  jxor g04429(.dina(n4684), .dinb(a35 ), .dout(n4685));
  jxor g04430(.dina(n4685), .dinb(n4677), .dout(n4686));
  jxor g04431(.dina(n4686), .dinb(n4647), .dout(n4687));
  jnot g04432(.din(n4687), .dout(n4688));
  jor  g04433(.dina(n3301), .dinb(n624), .dout(n4689));
  jor  g04434(.dina(n3136), .dinb(n512), .dout(n4690));
  jor  g04435(.dina(n3304), .dinb(n564), .dout(n4691));
  jor  g04436(.dina(n3306), .dinb(n627), .dout(n4692));
  jand g04437(.dina(n4692), .dinb(n4691), .dout(n4693));
  jand g04438(.dina(n4693), .dinb(n4690), .dout(n4694));
  jand g04439(.dina(n4694), .dinb(n4689), .dout(n4695));
  jxor g04440(.dina(n4695), .dinb(a32 ), .dout(n4696));
  jxor g04441(.dina(n4696), .dinb(n4688), .dout(n4697));
  jxor g04442(.dina(n4697), .dinb(n4642), .dout(n4698));
  jxor g04443(.dina(n4698), .dinb(n4637), .dout(n4699));
  jxor g04444(.dina(n4699), .dinb(n4628), .dout(n4700));
  jnot g04445(.din(n4700), .dout(n4701));
  jor  g04446(.dina(n2319), .dinb(n1019), .dout(n4702));
  jor  g04447(.dina(n2224), .dinb(n858), .dout(n4703));
  jor  g04448(.dina(n2322), .dinb(n939), .dout(n4704));
  jor  g04449(.dina(n2324), .dinb(n1022), .dout(n4705));
  jand g04450(.dina(n4705), .dinb(n4704), .dout(n4706));
  jand g04451(.dina(n4706), .dinb(n4703), .dout(n4707));
  jand g04452(.dina(n4707), .dinb(n4702), .dout(n4708));
  jxor g04453(.dina(n4708), .dinb(a26 ), .dout(n4709));
  jxor g04454(.dina(n4709), .dinb(n4701), .dout(n4710));
  jxor g04455(.dina(n4710), .dinb(n4623), .dout(n4711));
  jnot g04456(.din(n4711), .dout(n4712));
  jor  g04457(.dina(n1939), .dinb(n1397), .dout(n4713));
  jor  g04458(.dina(n1827), .dinb(n1193), .dout(n4714));
  jor  g04459(.dina(n1942), .dinb(n1290), .dout(n4715));
  jor  g04460(.dina(n1944), .dinb(n1400), .dout(n4716));
  jand g04461(.dina(n4716), .dinb(n4715), .dout(n4717));
  jand g04462(.dina(n4717), .dinb(n4714), .dout(n4718));
  jand g04463(.dina(n4718), .dinb(n4713), .dout(n4719));
  jxor g04464(.dina(n4719), .dinb(a23 ), .dout(n4720));
  jxor g04465(.dina(n4720), .dinb(n4712), .dout(n4721));
  jxor g04466(.dina(n4721), .dinb(n4618), .dout(n4722));
  jnot g04467(.din(n4722), .dout(n4723));
  jor  g04468(.dina(n1739), .dinb(n1566), .dout(n4724));
  jor  g04469(.dina(n1489), .dinb(n1420), .dout(n4725));
  jor  g04470(.dina(n1569), .dinb(n1620), .dout(n4726));
  jor  g04471(.dina(n1571), .dinb(n1742), .dout(n4727));
  jand g04472(.dina(n4727), .dinb(n4726), .dout(n4728));
  jand g04473(.dina(n4728), .dinb(n4725), .dout(n4729));
  jand g04474(.dina(n4729), .dinb(n4724), .dout(n4730));
  jxor g04475(.dina(n4730), .dinb(a20 ), .dout(n4731));
  jxor g04476(.dina(n4731), .dinb(n4723), .dout(n4732));
  jxor g04477(.dina(n4732), .dinb(n4615), .dout(n4733));
  jor  g04478(.dina(n2007), .dinb(n1245), .dout(n4734));
  jor  g04479(.dina(n1165), .dinb(n1867), .dout(n4735));
  jor  g04480(.dina(n1248), .dinb(n1887), .dout(n4736));
  jor  g04481(.dina(n1250), .dinb(n2010), .dout(n4737));
  jand g04482(.dina(n4737), .dinb(n4736), .dout(n4738));
  jand g04483(.dina(n4738), .dinb(n4735), .dout(n4739));
  jand g04484(.dina(n4739), .dinb(n4734), .dout(n4740));
  jxor g04485(.dina(n4740), .dinb(a17 ), .dout(n4741));
  jxor g04486(.dina(n4741), .dinb(n4733), .dout(n4742));
  jnot g04487(.din(n4742), .dout(n4743));
  jxor g04488(.dina(n4743), .dinb(n4611), .dout(n4744));
  jxor g04489(.dina(n4744), .dinb(n4605), .dout(n4745));
  jxor g04490(.dina(n4745), .dinb(n4596), .dout(n4746));
  jxor g04491(.dina(n4746), .dinb(n4592), .dout(n4747));
  jnot g04492(.din(n4747), .dout(n4748));
  jxor g04493(.dina(n4748), .dinb(n4583), .dout(n4749));
  jxor g04494(.dina(n4749), .dinb(n4579), .dout(n4750));
  jnot g04495(.din(n4750), .dout(n4751));
  jxor g04496(.dina(n4751), .dinb(n4570), .dout(n4752));
  jor  g04497(.dina(n4137), .dinb(n402), .dout(n4753));
  jor  g04498(.dina(n371), .dinb(n3588), .dout(n4754));
  jor  g04499(.dina(n405), .dinb(n3942), .dout(n4755));
  jor  g04500(.dina(n332), .dinb(n4140), .dout(n4756));
  jand g04501(.dina(n4756), .dinb(n4755), .dout(n4757));
  jand g04502(.dina(n4757), .dinb(n4754), .dout(n4758));
  jand g04503(.dina(n4758), .dinb(n4753), .dout(n4759));
  jxor g04504(.dina(n4759), .dinb(a5 ), .dout(n4760));
  jxor g04505(.dina(n4760), .dinb(n4752), .dout(n4761));
  jxor g04506(.dina(n4761), .dinb(n4566), .dout(n4762));
  jxor g04507(.dina(n4762), .dinb(n4563), .dout(n4763));
  jxor g04508(.dina(n4763), .dinb(n4548), .dout(f40 ));
  jand g04509(.dina(n4762), .dinb(n4563), .dout(n4765));
  jand g04510(.dina(n4763), .dinb(n4548), .dout(n4766));
  jor  g04511(.dina(n4766), .dinb(n4765), .dout(n4767));
  jor  g04512(.dina(n4760), .dinb(n4752), .dout(n4768));
  jnot g04513(.din(n4768), .dout(n4769));
  jand g04514(.dina(n4761), .dinb(n4566), .dout(n4770));
  jor  g04515(.dina(n4770), .dinb(n4769), .dout(n4771));
  jor  g04516(.dina(n4337), .dinb(n402), .dout(n4772));
  jor  g04517(.dina(n371), .dinb(n3942), .dout(n4773));
  jor  g04518(.dina(n405), .dinb(n4140), .dout(n4774));
  jor  g04519(.dina(n332), .dinb(n4340), .dout(n4775));
  jand g04520(.dina(n4775), .dinb(n4774), .dout(n4776));
  jand g04521(.dina(n4776), .dinb(n4773), .dout(n4777));
  jand g04522(.dina(n4777), .dinb(n4772), .dout(n4778));
  jxor g04523(.dina(n4778), .dinb(a5 ), .dout(n4779));
  jnot g04524(.din(n4779), .dout(n4780));
  jand g04525(.dina(n4749), .dinb(n4579), .dout(n4781));
  jand g04526(.dina(n4750), .dinb(n4570), .dout(n4782));
  jor  g04527(.dina(n4782), .dinb(n4781), .dout(n4783));
  jand g04528(.dina(n4746), .dinb(n4592), .dout(n4784));
  jnot g04529(.din(n4784), .dout(n4785));
  jor  g04530(.dina(n4748), .dinb(n4583), .dout(n4786));
  jand g04531(.dina(n4786), .dinb(n4785), .dout(n4787));
  jor  g04532(.dina(n3052), .dinb(n706), .dout(n4788));
  jor  g04533(.dina(n683), .dinb(n2870), .dout(n4789));
  jor  g04534(.dina(n709), .dinb(n3035), .dout(n4790));
  jor  g04535(.dina(n711), .dinb(n3055), .dout(n4791));
  jand g04536(.dina(n4791), .dinb(n4790), .dout(n4792));
  jand g04537(.dina(n4792), .dinb(n4789), .dout(n4793));
  jand g04538(.dina(n4793), .dinb(n4788), .dout(n4794));
  jxor g04539(.dina(n4794), .dinb(a11 ), .dout(n4795));
  jnot g04540(.din(n4795), .dout(n4796));
  jand g04541(.dina(n4744), .dinb(n4605), .dout(n4797));
  jand g04542(.dina(n4745), .dinb(n4596), .dout(n4798));
  jor  g04543(.dina(n4798), .dinb(n4797), .dout(n4799));
  jor  g04544(.dina(n2576), .dinb(n974), .dout(n4800));
  jor  g04545(.dina(n908), .dinb(n2407), .dout(n4801));
  jor  g04546(.dina(n977), .dinb(n2559), .dout(n4802));
  jor  g04547(.dina(n979), .dinb(n2579), .dout(n4803));
  jand g04548(.dina(n4803), .dinb(n4802), .dout(n4804));
  jand g04549(.dina(n4804), .dinb(n4801), .dout(n4805));
  jand g04550(.dina(n4805), .dinb(n4800), .dout(n4806));
  jxor g04551(.dina(n4806), .dinb(a14 ), .dout(n4807));
  jnot g04552(.din(n4807), .dout(n4808));
  jnot g04553(.din(n4733), .dout(n4809));
  jor  g04554(.dina(n4741), .dinb(n4809), .dout(n4810));
  jnot g04555(.din(n4810), .dout(n4811));
  jand g04556(.dina(n4743), .dinb(n4611), .dout(n4812));
  jor  g04557(.dina(n4812), .dinb(n4811), .dout(n4813));
  jor  g04558(.dina(n2145), .dinb(n1245), .dout(n4814));
  jor  g04559(.dina(n1165), .dinb(n1887), .dout(n4815));
  jor  g04560(.dina(n1248), .dinb(n2010), .dout(n4816));
  jor  g04561(.dina(n1250), .dinb(n2148), .dout(n4817));
  jand g04562(.dina(n4817), .dinb(n4816), .dout(n4818));
  jand g04563(.dina(n4818), .dinb(n4815), .dout(n4819));
  jand g04564(.dina(n4819), .dinb(n4814), .dout(n4820));
  jxor g04565(.dina(n4820), .dinb(a17 ), .dout(n4821));
  jnot g04566(.din(n4821), .dout(n4822));
  jor  g04567(.dina(n4731), .dinb(n4723), .dout(n4823));
  jnot g04568(.din(n4823), .dout(n4824));
  jand g04569(.dina(n4732), .dinb(n4615), .dout(n4825));
  jor  g04570(.dina(n4825), .dinb(n4824), .dout(n4826));
  jor  g04571(.dina(n4720), .dinb(n4712), .dout(n4827));
  jand g04572(.dina(n4721), .dinb(n4618), .dout(n4828));
  jnot g04573(.din(n4828), .dout(n4829));
  jand g04574(.dina(n4829), .dinb(n4827), .dout(n4830));
  jnot g04575(.din(n4830), .dout(n4831));
  jor  g04576(.dina(n4709), .dinb(n4701), .dout(n4832));
  jand g04577(.dina(n4710), .dinb(n4623), .dout(n4833));
  jnot g04578(.din(n4833), .dout(n4834));
  jand g04579(.dina(n4834), .dinb(n4832), .dout(n4835));
  jnot g04580(.din(n4835), .dout(n4836));
  jor  g04581(.dina(n2319), .dinb(n1190), .dout(n4837));
  jor  g04582(.dina(n2224), .dinb(n939), .dout(n4838));
  jor  g04583(.dina(n2322), .dinb(n1022), .dout(n4839));
  jor  g04584(.dina(n2324), .dinb(n1193), .dout(n4840));
  jand g04585(.dina(n4840), .dinb(n4839), .dout(n4841));
  jand g04586(.dina(n4841), .dinb(n4838), .dout(n4842));
  jand g04587(.dina(n4842), .dinb(n4837), .dout(n4843));
  jxor g04588(.dina(n4843), .dinb(a26 ), .dout(n4844));
  jnot g04589(.din(n4844), .dout(n4845));
  jand g04590(.dina(n4698), .dinb(n4637), .dout(n4846));
  jand g04591(.dina(n4699), .dinb(n4628), .dout(n4847));
  jor  g04592(.dina(n4847), .dinb(n4846), .dout(n4848));
  jor  g04593(.dina(n2784), .dinb(n855), .dout(n4849));
  jor  g04594(.dina(n2661), .dinb(n758), .dout(n4850));
  jor  g04595(.dina(n2787), .dinb(n778), .dout(n4851));
  jor  g04596(.dina(n2789), .dinb(n858), .dout(n4852));
  jand g04597(.dina(n4852), .dinb(n4851), .dout(n4853));
  jand g04598(.dina(n4853), .dinb(n4850), .dout(n4854));
  jand g04599(.dina(n4854), .dinb(n4849), .dout(n4855));
  jxor g04600(.dina(n4855), .dinb(a29 ), .dout(n4856));
  jnot g04601(.din(n4856), .dout(n4857));
  jor  g04602(.dina(n4696), .dinb(n4688), .dout(n4858));
  jand g04603(.dina(n4697), .dinb(n4642), .dout(n4859));
  jnot g04604(.din(n4859), .dout(n4860));
  jand g04605(.dina(n4860), .dinb(n4858), .dout(n4861));
  jnot g04606(.din(n4861), .dout(n4862));
  jor  g04607(.dina(n3301), .dinb(n644), .dout(n4863));
  jor  g04608(.dina(n3136), .dinb(n564), .dout(n4864));
  jor  g04609(.dina(n3304), .dinb(n627), .dout(n4865));
  jor  g04610(.dina(n3306), .dinb(n647), .dout(n4866));
  jand g04611(.dina(n4866), .dinb(n4865), .dout(n4867));
  jand g04612(.dina(n4867), .dinb(n4864), .dout(n4868));
  jand g04613(.dina(n4868), .dinb(n4863), .dout(n4869));
  jxor g04614(.dina(n4869), .dinb(a32 ), .dout(n4870));
  jnot g04615(.din(n4870), .dout(n4871));
  jor  g04616(.dina(n4685), .dinb(n4677), .dout(n4872));
  jand g04617(.dina(n4686), .dinb(n4647), .dout(n4873));
  jnot g04618(.din(n4873), .dout(n4874));
  jand g04619(.dina(n4874), .dinb(n4872), .dout(n4875));
  jnot g04620(.din(n4875), .dout(n4876));
  jor  g04621(.dina(n3849), .dinb(n509), .dout(n4877));
  jor  g04622(.dina(n3689), .dinb(n395), .dout(n4878));
  jor  g04623(.dina(n3852), .dinb(n431), .dout(n4879));
  jor  g04624(.dina(n3854), .dinb(n512), .dout(n4880));
  jand g04625(.dina(n4880), .dinb(n4879), .dout(n4881));
  jand g04626(.dina(n4881), .dinb(n4878), .dout(n4882));
  jand g04627(.dina(n4882), .dinb(n4877), .dout(n4883));
  jxor g04628(.dina(n4883), .dinb(a35 ), .dout(n4884));
  jnot g04629(.din(n4884), .dout(n4885));
  jand g04630(.dina(n4674), .dinb(n4660), .dout(n4886));
  jand g04631(.dina(n4675), .dinb(n4651), .dout(n4887));
  jor  g04632(.dina(n4887), .dinb(n4886), .dout(n4888));
  jor  g04633(.dina(n4415), .dinb(n354), .dout(n4889));
  jor  g04634(.dina(n4272), .dinb(n299), .dout(n4890));
  jor  g04635(.dina(n4418), .dinb(n322), .dout(n4891));
  jor  g04636(.dina(n4420), .dinb(n357), .dout(n4892));
  jand g04637(.dina(n4892), .dinb(n4891), .dout(n4893));
  jand g04638(.dina(n4893), .dinb(n4890), .dout(n4894));
  jand g04639(.dina(n4894), .dinb(n4889), .dout(n4895));
  jxor g04640(.dina(n4895), .dinb(a38 ), .dout(n4896));
  jnot g04641(.din(n4896), .dout(n4897));
  jnot g04642(.din(n4673), .dout(n4898));
  jand g04643(.dina(n4429), .dinb(a41 ), .dout(n4899));
  jand g04644(.dina(n4899), .dinb(n4898), .dout(n4900));
  jnot g04645(.din(n4900), .dout(n4901));
  jand g04646(.dina(n4901), .dinb(a41 ), .dout(n4902));
  jor  g04647(.dina(n4667), .dinb(n4663), .dout(n4903));
  jor  g04648(.dina(n4903), .dinb(n4427), .dout(n4904));
  jnot g04649(.din(n4904), .dout(n4905));
  jand g04650(.dina(n4905), .dinb(b0 ), .dout(n4906));
  jand g04651(.dina(n4664), .dinb(b2 ), .dout(n4907));
  jand g04652(.dina(n4668), .dinb(b1 ), .dout(n4908));
  jand g04653(.dina(n4670), .dinb(n375), .dout(n4909));
  jor  g04654(.dina(n4909), .dinb(n4908), .dout(n4910));
  jor  g04655(.dina(n4910), .dinb(n4907), .dout(n4911));
  jor  g04656(.dina(n4911), .dinb(n4906), .dout(n4912));
  jxor g04657(.dina(n4912), .dinb(n4902), .dout(n4913));
  jxor g04658(.dina(n4913), .dinb(n4897), .dout(n4914));
  jxor g04659(.dina(n4914), .dinb(n4888), .dout(n4915));
  jxor g04660(.dina(n4915), .dinb(n4885), .dout(n4916));
  jxor g04661(.dina(n4916), .dinb(n4876), .dout(n4917));
  jxor g04662(.dina(n4917), .dinb(n4871), .dout(n4918));
  jxor g04663(.dina(n4918), .dinb(n4862), .dout(n4919));
  jxor g04664(.dina(n4919), .dinb(n4857), .dout(n4920));
  jxor g04665(.dina(n4920), .dinb(n4848), .dout(n4921));
  jxor g04666(.dina(n4921), .dinb(n4845), .dout(n4922));
  jxor g04667(.dina(n4922), .dinb(n4836), .dout(n4923));
  jnot g04668(.din(n4923), .dout(n4924));
  jor  g04669(.dina(n1939), .dinb(n1417), .dout(n4925));
  jor  g04670(.dina(n1827), .dinb(n1290), .dout(n4926));
  jor  g04671(.dina(n1942), .dinb(n1400), .dout(n4927));
  jor  g04672(.dina(n1944), .dinb(n1420), .dout(n4928));
  jand g04673(.dina(n4928), .dinb(n4927), .dout(n4929));
  jand g04674(.dina(n4929), .dinb(n4926), .dout(n4930));
  jand g04675(.dina(n4930), .dinb(n4925), .dout(n4931));
  jxor g04676(.dina(n4931), .dinb(a23 ), .dout(n4932));
  jxor g04677(.dina(n4932), .dinb(n4924), .dout(n4933));
  jxor g04678(.dina(n4933), .dinb(n4831), .dout(n4934));
  jnot g04679(.din(n4934), .dout(n4935));
  jor  g04680(.dina(n1864), .dinb(n1566), .dout(n4936));
  jor  g04681(.dina(n1489), .dinb(n1620), .dout(n4937));
  jor  g04682(.dina(n1569), .dinb(n1742), .dout(n4938));
  jor  g04683(.dina(n1571), .dinb(n1867), .dout(n4939));
  jand g04684(.dina(n4939), .dinb(n4938), .dout(n4940));
  jand g04685(.dina(n4940), .dinb(n4937), .dout(n4941));
  jand g04686(.dina(n4941), .dinb(n4936), .dout(n4942));
  jxor g04687(.dina(n4942), .dinb(a20 ), .dout(n4943));
  jxor g04688(.dina(n4943), .dinb(n4935), .dout(n4944));
  jxor g04689(.dina(n4944), .dinb(n4826), .dout(n4945));
  jxor g04690(.dina(n4945), .dinb(n4822), .dout(n4946));
  jxor g04691(.dina(n4946), .dinb(n4813), .dout(n4947));
  jxor g04692(.dina(n4947), .dinb(n4808), .dout(n4948));
  jxor g04693(.dina(n4948), .dinb(n4799), .dout(n4949));
  jxor g04694(.dina(n4949), .dinb(n4796), .dout(n4950));
  jnot g04695(.din(n4950), .dout(n4951));
  jxor g04696(.dina(n4951), .dinb(n4787), .dout(n4952));
  jnot g04697(.din(n4952), .dout(n4953));
  jor  g04698(.dina(n3585), .dinb(n528), .dout(n4954));
  jor  g04699(.dina(n490), .dinb(n3230), .dout(n4955));
  jor  g04700(.dina(n531), .dinb(n3403), .dout(n4956));
  jor  g04701(.dina(n533), .dinb(n3588), .dout(n4957));
  jand g04702(.dina(n4957), .dinb(n4956), .dout(n4958));
  jand g04703(.dina(n4958), .dinb(n4955), .dout(n4959));
  jand g04704(.dina(n4959), .dinb(n4954), .dout(n4960));
  jxor g04705(.dina(n4960), .dinb(a8 ), .dout(n4961));
  jxor g04706(.dina(n4961), .dinb(n4953), .dout(n4962));
  jxor g04707(.dina(n4962), .dinb(n4783), .dout(n4963));
  jxor g04708(.dina(n4963), .dinb(n4780), .dout(n4964));
  jxor g04709(.dina(n4964), .dinb(n4771), .dout(n4965));
  jand g04710(.dina(b40 ), .dinb(b39 ), .dout(n4966));
  jand g04711(.dina(n4552), .dinb(n4551), .dout(n4967));
  jor  g04712(.dina(n4967), .dinb(n4966), .dout(n4968));
  jxor g04713(.dina(b41 ), .dinb(b40 ), .dout(n4969));
  jnot g04714(.din(n4969), .dout(n4970));
  jxor g04715(.dina(n4970), .dinb(n4968), .dout(n4971));
  jor  g04716(.dina(n4971), .dinb(n264), .dout(n4972));
  jor  g04717(.dina(n284), .dinb(n4537), .dout(n4973));
  jnot g04718(.din(b41 ), .dout(n4974));
  jor  g04719(.dina(n269), .dinb(n4974), .dout(n4975));
  jor  g04720(.dina(n271), .dinb(n4557), .dout(n4976));
  jand g04721(.dina(n4976), .dinb(n4975), .dout(n4977));
  jand g04722(.dina(n4977), .dinb(n4973), .dout(n4978));
  jand g04723(.dina(n4978), .dinb(n4972), .dout(n4979));
  jxor g04724(.dina(n4979), .dinb(n260), .dout(n4980));
  jxor g04725(.dina(n4980), .dinb(n4965), .dout(n4981));
  jxor g04726(.dina(n4981), .dinb(n4767), .dout(f41 ));
  jand g04727(.dina(n4980), .dinb(n4965), .dout(n4983));
  jand g04728(.dina(n4981), .dinb(n4767), .dout(n4984));
  jor  g04729(.dina(n4984), .dinb(n4983), .dout(n4985));
  jand g04730(.dina(b41 ), .dinb(b40 ), .dout(n4986));
  jand g04731(.dina(n4969), .dinb(n4968), .dout(n4987));
  jor  g04732(.dina(n4987), .dinb(n4986), .dout(n4988));
  jxor g04733(.dina(b42 ), .dinb(b41 ), .dout(n4989));
  jnot g04734(.din(n4989), .dout(n4990));
  jxor g04735(.dina(n4990), .dinb(n4988), .dout(n4991));
  jor  g04736(.dina(n4991), .dinb(n264), .dout(n4992));
  jor  g04737(.dina(n284), .dinb(n4557), .dout(n4993));
  jnot g04738(.din(b42 ), .dout(n4994));
  jor  g04739(.dina(n269), .dinb(n4994), .dout(n4995));
  jor  g04740(.dina(n271), .dinb(n4974), .dout(n4996));
  jand g04741(.dina(n4996), .dinb(n4995), .dout(n4997));
  jand g04742(.dina(n4997), .dinb(n4993), .dout(n4998));
  jand g04743(.dina(n4998), .dinb(n4992), .dout(n4999));
  jxor g04744(.dina(n4999), .dinb(n260), .dout(n5000));
  jand g04745(.dina(n4963), .dinb(n4780), .dout(n5001));
  jand g04746(.dina(n4964), .dinb(n4771), .dout(n5002));
  jor  g04747(.dina(n5002), .dinb(n5001), .dout(n5003));
  jor  g04748(.dina(n4534), .dinb(n402), .dout(n5004));
  jor  g04749(.dina(n371), .dinb(n4140), .dout(n5005));
  jor  g04750(.dina(n405), .dinb(n4340), .dout(n5006));
  jor  g04751(.dina(n332), .dinb(n4537), .dout(n5007));
  jand g04752(.dina(n5007), .dinb(n5006), .dout(n5008));
  jand g04753(.dina(n5008), .dinb(n5005), .dout(n5009));
  jand g04754(.dina(n5009), .dinb(n5004), .dout(n5010));
  jxor g04755(.dina(n5010), .dinb(a5 ), .dout(n5011));
  jnot g04756(.din(n5011), .dout(n5012));
  jor  g04757(.dina(n4961), .dinb(n4953), .dout(n5013));
  jnot g04758(.din(n5013), .dout(n5014));
  jand g04759(.dina(n4962), .dinb(n4783), .dout(n5015));
  jor  g04760(.dina(n5015), .dinb(n5014), .dout(n5016));
  jor  g04761(.dina(n3939), .dinb(n528), .dout(n5017));
  jor  g04762(.dina(n490), .dinb(n3403), .dout(n5018));
  jor  g04763(.dina(n531), .dinb(n3588), .dout(n5019));
  jor  g04764(.dina(n533), .dinb(n3942), .dout(n5020));
  jand g04765(.dina(n5020), .dinb(n5019), .dout(n5021));
  jand g04766(.dina(n5021), .dinb(n5018), .dout(n5022));
  jand g04767(.dina(n5022), .dinb(n5017), .dout(n5023));
  jxor g04768(.dina(n5023), .dinb(a8 ), .dout(n5024));
  jnot g04769(.din(n5024), .dout(n5025));
  jand g04770(.dina(n4949), .dinb(n4796), .dout(n5026));
  jnot g04771(.din(n5026), .dout(n5027));
  jor  g04772(.dina(n4951), .dinb(n4787), .dout(n5028));
  jand g04773(.dina(n5028), .dinb(n5027), .dout(n5029));
  jand g04774(.dina(n4947), .dinb(n4808), .dout(n5030));
  jand g04775(.dina(n4948), .dinb(n4799), .dout(n5031));
  jor  g04776(.dina(n5031), .dinb(n5030), .dout(n5032));
  jor  g04777(.dina(n2867), .dinb(n974), .dout(n5033));
  jor  g04778(.dina(n908), .dinb(n2559), .dout(n5034));
  jor  g04779(.dina(n977), .dinb(n2579), .dout(n5035));
  jor  g04780(.dina(n979), .dinb(n2870), .dout(n5036));
  jand g04781(.dina(n5036), .dinb(n5035), .dout(n5037));
  jand g04782(.dina(n5037), .dinb(n5034), .dout(n5038));
  jand g04783(.dina(n5038), .dinb(n5033), .dout(n5039));
  jxor g04784(.dina(n5039), .dinb(a14 ), .dout(n5040));
  jnot g04785(.din(n5040), .dout(n5041));
  jand g04786(.dina(n4945), .dinb(n4822), .dout(n5042));
  jand g04787(.dina(n4946), .dinb(n4813), .dout(n5043));
  jor  g04788(.dina(n5043), .dinb(n5042), .dout(n5044));
  jor  g04789(.dina(n4943), .dinb(n4935), .dout(n5045));
  jnot g04790(.din(n5045), .dout(n5046));
  jand g04791(.dina(n4944), .dinb(n4826), .dout(n5047));
  jor  g04792(.dina(n5047), .dinb(n5046), .dout(n5048));
  jor  g04793(.dina(n4932), .dinb(n4924), .dout(n5049));
  jand g04794(.dina(n4933), .dinb(n4831), .dout(n5050));
  jnot g04795(.din(n5050), .dout(n5051));
  jand g04796(.dina(n5051), .dinb(n5049), .dout(n5052));
  jnot g04797(.din(n5052), .dout(n5053));
  jand g04798(.dina(n4921), .dinb(n4845), .dout(n5054));
  jand g04799(.dina(n4922), .dinb(n4836), .dout(n5055));
  jor  g04800(.dina(n5055), .dinb(n5054), .dout(n5056));
  jor  g04801(.dina(n2319), .dinb(n1287), .dout(n5057));
  jor  g04802(.dina(n2224), .dinb(n1022), .dout(n5058));
  jor  g04803(.dina(n2322), .dinb(n1193), .dout(n5059));
  jor  g04804(.dina(n2324), .dinb(n1290), .dout(n5060));
  jand g04805(.dina(n5060), .dinb(n5059), .dout(n5061));
  jand g04806(.dina(n5061), .dinb(n5058), .dout(n5062));
  jand g04807(.dina(n5062), .dinb(n5057), .dout(n5063));
  jxor g04808(.dina(n5063), .dinb(a26 ), .dout(n5064));
  jnot g04809(.din(n5064), .dout(n5065));
  jand g04810(.dina(n4919), .dinb(n4857), .dout(n5066));
  jand g04811(.dina(n4920), .dinb(n4848), .dout(n5067));
  jor  g04812(.dina(n5067), .dinb(n5066), .dout(n5068));
  jor  g04813(.dina(n2784), .dinb(n936), .dout(n5069));
  jor  g04814(.dina(n2661), .dinb(n778), .dout(n5070));
  jor  g04815(.dina(n2787), .dinb(n858), .dout(n5071));
  jor  g04816(.dina(n2789), .dinb(n939), .dout(n5072));
  jand g04817(.dina(n5072), .dinb(n5071), .dout(n5073));
  jand g04818(.dina(n5073), .dinb(n5070), .dout(n5074));
  jand g04819(.dina(n5074), .dinb(n5069), .dout(n5075));
  jxor g04820(.dina(n5075), .dinb(a29 ), .dout(n5076));
  jnot g04821(.din(n5076), .dout(n5077));
  jand g04822(.dina(n4917), .dinb(n4871), .dout(n5078));
  jand g04823(.dina(n4918), .dinb(n4862), .dout(n5079));
  jor  g04824(.dina(n5079), .dinb(n5078), .dout(n5080));
  jor  g04825(.dina(n3301), .dinb(n755), .dout(n5081));
  jor  g04826(.dina(n3136), .dinb(n627), .dout(n5082));
  jor  g04827(.dina(n3304), .dinb(n647), .dout(n5083));
  jor  g04828(.dina(n3306), .dinb(n758), .dout(n5084));
  jand g04829(.dina(n5084), .dinb(n5083), .dout(n5085));
  jand g04830(.dina(n5085), .dinb(n5082), .dout(n5086));
  jand g04831(.dina(n5086), .dinb(n5081), .dout(n5087));
  jxor g04832(.dina(n5087), .dinb(a32 ), .dout(n5088));
  jnot g04833(.din(n5088), .dout(n5089));
  jand g04834(.dina(n4915), .dinb(n4885), .dout(n5090));
  jand g04835(.dina(n4916), .dinb(n4876), .dout(n5091));
  jor  g04836(.dina(n5091), .dinb(n5090), .dout(n5092));
  jand g04837(.dina(n4913), .dinb(n4897), .dout(n5093));
  jand g04838(.dina(n4914), .dinb(n4888), .dout(n5094));
  jor  g04839(.dina(n5094), .dinb(n5093), .dout(n5095));
  jnot g04840(.din(n4670), .dout(n5096));
  jor  g04841(.dina(n5096), .dinb(n296), .dout(n5097));
  jor  g04842(.dina(n4904), .dinb(n267), .dout(n5098));
  jnot g04843(.din(n4668), .dout(n5099));
  jor  g04844(.dina(n5099), .dinb(n279), .dout(n5100));
  jnot g04845(.din(n4664), .dout(n5101));
  jor  g04846(.dina(n5101), .dinb(n299), .dout(n5102));
  jand g04847(.dina(n5102), .dinb(n5100), .dout(n5103));
  jand g04848(.dina(n5103), .dinb(n5098), .dout(n5104));
  jand g04849(.dina(n5104), .dinb(n5097), .dout(n5105));
  jxor g04850(.dina(n5105), .dinb(a41 ), .dout(n5106));
  jnot g04851(.din(n5106), .dout(n5107));
  jxor g04852(.dina(a42 ), .dinb(a41 ), .dout(n5108));
  jand g04853(.dina(n5108), .dinb(b0 ), .dout(n5109));
  jnot g04854(.din(n5109), .dout(n5110));
  jor  g04855(.dina(n4912), .dinb(n4901), .dout(n5111));
  jxor g04856(.dina(n5111), .dinb(n5110), .dout(n5112));
  jxor g04857(.dina(n5112), .dinb(n5107), .dout(n5113));
  jnot g04858(.din(n5113), .dout(n5114));
  jor  g04859(.dina(n4415), .dinb(n392), .dout(n5115));
  jor  g04860(.dina(n4272), .dinb(n322), .dout(n5116));
  jor  g04861(.dina(n4418), .dinb(n357), .dout(n5117));
  jor  g04862(.dina(n4420), .dinb(n395), .dout(n5118));
  jand g04863(.dina(n5118), .dinb(n5117), .dout(n5119));
  jand g04864(.dina(n5119), .dinb(n5116), .dout(n5120));
  jand g04865(.dina(n5120), .dinb(n5115), .dout(n5121));
  jxor g04866(.dina(n5121), .dinb(a38 ), .dout(n5122));
  jxor g04867(.dina(n5122), .dinb(n5114), .dout(n5123));
  jxor g04868(.dina(n5123), .dinb(n5095), .dout(n5124));
  jnot g04869(.din(n5124), .dout(n5125));
  jor  g04870(.dina(n3849), .dinb(n561), .dout(n5126));
  jor  g04871(.dina(n3689), .dinb(n431), .dout(n5127));
  jor  g04872(.dina(n3852), .dinb(n512), .dout(n5128));
  jor  g04873(.dina(n3854), .dinb(n564), .dout(n5129));
  jand g04874(.dina(n5129), .dinb(n5128), .dout(n5130));
  jand g04875(.dina(n5130), .dinb(n5127), .dout(n5131));
  jand g04876(.dina(n5131), .dinb(n5126), .dout(n5132));
  jxor g04877(.dina(n5132), .dinb(a35 ), .dout(n5133));
  jxor g04878(.dina(n5133), .dinb(n5125), .dout(n5134));
  jxor g04879(.dina(n5134), .dinb(n5092), .dout(n5135));
  jxor g04880(.dina(n5135), .dinb(n5089), .dout(n5136));
  jxor g04881(.dina(n5136), .dinb(n5080), .dout(n5137));
  jxor g04882(.dina(n5137), .dinb(n5077), .dout(n5138));
  jxor g04883(.dina(n5138), .dinb(n5068), .dout(n5139));
  jxor g04884(.dina(n5139), .dinb(n5065), .dout(n5140));
  jxor g04885(.dina(n5140), .dinb(n5056), .dout(n5141));
  jnot g04886(.din(n5141), .dout(n5142));
  jor  g04887(.dina(n1939), .dinb(n1617), .dout(n5143));
  jor  g04888(.dina(n1827), .dinb(n1400), .dout(n5144));
  jor  g04889(.dina(n1942), .dinb(n1420), .dout(n5145));
  jor  g04890(.dina(n1944), .dinb(n1620), .dout(n5146));
  jand g04891(.dina(n5146), .dinb(n5145), .dout(n5147));
  jand g04892(.dina(n5147), .dinb(n5144), .dout(n5148));
  jand g04893(.dina(n5148), .dinb(n5143), .dout(n5149));
  jxor g04894(.dina(n5149), .dinb(a23 ), .dout(n5150));
  jxor g04895(.dina(n5150), .dinb(n5142), .dout(n5151));
  jxor g04896(.dina(n5151), .dinb(n5053), .dout(n5152));
  jor  g04897(.dina(n1884), .dinb(n1566), .dout(n5153));
  jor  g04898(.dina(n1489), .dinb(n1742), .dout(n5154));
  jor  g04899(.dina(n1569), .dinb(n1867), .dout(n5155));
  jor  g04900(.dina(n1571), .dinb(n1887), .dout(n5156));
  jand g04901(.dina(n5156), .dinb(n5155), .dout(n5157));
  jand g04902(.dina(n5157), .dinb(n5154), .dout(n5158));
  jand g04903(.dina(n5158), .dinb(n5153), .dout(n5159));
  jxor g04904(.dina(n5159), .dinb(a20 ), .dout(n5160));
  jxor g04905(.dina(n5160), .dinb(n5152), .dout(n5161));
  jxor g04906(.dina(n5161), .dinb(n5048), .dout(n5162));
  jor  g04907(.dina(n2404), .dinb(n1245), .dout(n5163));
  jor  g04908(.dina(n1165), .dinb(n2010), .dout(n5164));
  jor  g04909(.dina(n1248), .dinb(n2148), .dout(n5165));
  jor  g04910(.dina(n1250), .dinb(n2407), .dout(n5166));
  jand g04911(.dina(n5166), .dinb(n5165), .dout(n5167));
  jand g04912(.dina(n5167), .dinb(n5164), .dout(n5168));
  jand g04913(.dina(n5168), .dinb(n5163), .dout(n5169));
  jxor g04914(.dina(n5169), .dinb(a17 ), .dout(n5170));
  jxor g04915(.dina(n5170), .dinb(n5162), .dout(n5171));
  jxor g04916(.dina(n5171), .dinb(n5044), .dout(n5172));
  jxor g04917(.dina(n5172), .dinb(n5041), .dout(n5173));
  jxor g04918(.dina(n5173), .dinb(n5032), .dout(n5174));
  jor  g04919(.dina(n3227), .dinb(n706), .dout(n5175));
  jor  g04920(.dina(n683), .dinb(n3035), .dout(n5176));
  jor  g04921(.dina(n709), .dinb(n3055), .dout(n5177));
  jor  g04922(.dina(n711), .dinb(n3230), .dout(n5178));
  jand g04923(.dina(n5178), .dinb(n5177), .dout(n5179));
  jand g04924(.dina(n5179), .dinb(n5176), .dout(n5180));
  jand g04925(.dina(n5180), .dinb(n5175), .dout(n5181));
  jxor g04926(.dina(n5181), .dinb(a11 ), .dout(n5182));
  jxor g04927(.dina(n5182), .dinb(n5174), .dout(n5183));
  jxor g04928(.dina(n5183), .dinb(n5029), .dout(n5184));
  jxor g04929(.dina(n5184), .dinb(n5025), .dout(n5185));
  jxor g04930(.dina(n5185), .dinb(n5016), .dout(n5186));
  jxor g04931(.dina(n5186), .dinb(n5012), .dout(n5187));
  jxor g04932(.dina(n5187), .dinb(n5003), .dout(n5188));
  jxor g04933(.dina(n5188), .dinb(n5000), .dout(n5189));
  jxor g04934(.dina(n5189), .dinb(n4985), .dout(f42 ));
  jand g04935(.dina(n5188), .dinb(n5000), .dout(n5191));
  jand g04936(.dina(n5189), .dinb(n4985), .dout(n5192));
  jor  g04937(.dina(n5192), .dinb(n5191), .dout(n5193));
  jand g04938(.dina(n5186), .dinb(n5012), .dout(n5194));
  jand g04939(.dina(n5187), .dinb(n5003), .dout(n5195));
  jor  g04940(.dina(n5195), .dinb(n5194), .dout(n5196));
  jor  g04941(.dina(n4554), .dinb(n402), .dout(n5197));
  jor  g04942(.dina(n371), .dinb(n4340), .dout(n5198));
  jor  g04943(.dina(n405), .dinb(n4537), .dout(n5199));
  jor  g04944(.dina(n332), .dinb(n4557), .dout(n5200));
  jand g04945(.dina(n5200), .dinb(n5199), .dout(n5201));
  jand g04946(.dina(n5201), .dinb(n5198), .dout(n5202));
  jand g04947(.dina(n5202), .dinb(n5197), .dout(n5203));
  jxor g04948(.dina(n5203), .dinb(a5 ), .dout(n5204));
  jnot g04949(.din(n5204), .dout(n5205));
  jand g04950(.dina(n5184), .dinb(n5025), .dout(n5206));
  jand g04951(.dina(n5185), .dinb(n5016), .dout(n5207));
  jor  g04952(.dina(n5207), .dinb(n5206), .dout(n5208));
  jnot g04953(.din(n5174), .dout(n5209));
  jor  g04954(.dina(n5182), .dinb(n5209), .dout(n5210));
  jor  g04955(.dina(n5183), .dinb(n5029), .dout(n5211));
  jand g04956(.dina(n5211), .dinb(n5210), .dout(n5212));
  jand g04957(.dina(n5172), .dinb(n5041), .dout(n5213));
  jand g04958(.dina(n5173), .dinb(n5032), .dout(n5214));
  jor  g04959(.dina(n5214), .dinb(n5213), .dout(n5215));
  jor  g04960(.dina(n3032), .dinb(n974), .dout(n5216));
  jor  g04961(.dina(n908), .dinb(n2579), .dout(n5217));
  jor  g04962(.dina(n977), .dinb(n2870), .dout(n5218));
  jor  g04963(.dina(n979), .dinb(n3035), .dout(n5219));
  jand g04964(.dina(n5219), .dinb(n5218), .dout(n5220));
  jand g04965(.dina(n5220), .dinb(n5217), .dout(n5221));
  jand g04966(.dina(n5221), .dinb(n5216), .dout(n5222));
  jxor g04967(.dina(n5222), .dinb(a14 ), .dout(n5223));
  jnot g04968(.din(n5223), .dout(n5224));
  jor  g04969(.dina(n5170), .dinb(n5162), .dout(n5225));
  jnot g04970(.din(n5225), .dout(n5226));
  jand g04971(.dina(n5171), .dinb(n5044), .dout(n5227));
  jor  g04972(.dina(n5227), .dinb(n5226), .dout(n5228));
  jor  g04973(.dina(n2556), .dinb(n1245), .dout(n5229));
  jor  g04974(.dina(n1165), .dinb(n2148), .dout(n5230));
  jor  g04975(.dina(n1248), .dinb(n2407), .dout(n5231));
  jor  g04976(.dina(n1250), .dinb(n2559), .dout(n5232));
  jand g04977(.dina(n5232), .dinb(n5231), .dout(n5233));
  jand g04978(.dina(n5233), .dinb(n5230), .dout(n5234));
  jand g04979(.dina(n5234), .dinb(n5229), .dout(n5235));
  jxor g04980(.dina(n5235), .dinb(a17 ), .dout(n5236));
  jnot g04981(.din(n5236), .dout(n5237));
  jnot g04982(.din(n5152), .dout(n5238));
  jor  g04983(.dina(n5160), .dinb(n5238), .dout(n5239));
  jnot g04984(.din(n5239), .dout(n5240));
  jnot g04985(.din(n5161), .dout(n5241));
  jand g04986(.dina(n5241), .dinb(n5048), .dout(n5242));
  jor  g04987(.dina(n5242), .dinb(n5240), .dout(n5243));
  jor  g04988(.dina(n5150), .dinb(n5142), .dout(n5244));
  jnot g04989(.din(n5244), .dout(n5245));
  jand g04990(.dina(n5151), .dinb(n5053), .dout(n5246));
  jor  g04991(.dina(n5246), .dinb(n5245), .dout(n5247));
  jand g04992(.dina(n5139), .dinb(n5065), .dout(n5248));
  jand g04993(.dina(n5140), .dinb(n5056), .dout(n5249));
  jor  g04994(.dina(n5249), .dinb(n5248), .dout(n5250));
  jand g04995(.dina(n5137), .dinb(n5077), .dout(n5251));
  jand g04996(.dina(n5138), .dinb(n5068), .dout(n5252));
  jor  g04997(.dina(n5252), .dinb(n5251), .dout(n5253));
  jand g04998(.dina(n5135), .dinb(n5089), .dout(n5254));
  jand g04999(.dina(n5136), .dinb(n5080), .dout(n5255));
  jor  g05000(.dina(n5255), .dinb(n5254), .dout(n5256));
  jor  g05001(.dina(n3301), .dinb(n775), .dout(n5257));
  jor  g05002(.dina(n3136), .dinb(n647), .dout(n5258));
  jor  g05003(.dina(n3304), .dinb(n758), .dout(n5259));
  jor  g05004(.dina(n3306), .dinb(n778), .dout(n5260));
  jand g05005(.dina(n5260), .dinb(n5259), .dout(n5261));
  jand g05006(.dina(n5261), .dinb(n5258), .dout(n5262));
  jand g05007(.dina(n5262), .dinb(n5257), .dout(n5263));
  jxor g05008(.dina(n5263), .dinb(a32 ), .dout(n5264));
  jnot g05009(.din(n5264), .dout(n5265));
  jor  g05010(.dina(n5133), .dinb(n5125), .dout(n5266));
  jand g05011(.dina(n5134), .dinb(n5092), .dout(n5267));
  jnot g05012(.din(n5267), .dout(n5268));
  jand g05013(.dina(n5268), .dinb(n5266), .dout(n5269));
  jnot g05014(.din(n5269), .dout(n5270));
  jor  g05015(.dina(n5122), .dinb(n5114), .dout(n5271));
  jand g05016(.dina(n5123), .dinb(n5095), .dout(n5272));
  jnot g05017(.din(n5272), .dout(n5273));
  jand g05018(.dina(n5273), .dinb(n5271), .dout(n5274));
  jnot g05019(.din(n5274), .dout(n5275));
  jnot g05020(.din(n5111), .dout(n5276));
  jand g05021(.dina(n5276), .dinb(n5109), .dout(n5277));
  jand g05022(.dina(n5112), .dinb(n5107), .dout(n5278));
  jor  g05023(.dina(n5278), .dinb(n5277), .dout(n5279));
  jor  g05024(.dina(n5096), .dinb(n319), .dout(n5280));
  jor  g05025(.dina(n4904), .dinb(n279), .dout(n5281));
  jor  g05026(.dina(n5099), .dinb(n299), .dout(n5282));
  jor  g05027(.dina(n5101), .dinb(n322), .dout(n5283));
  jand g05028(.dina(n5283), .dinb(n5282), .dout(n5284));
  jand g05029(.dina(n5284), .dinb(n5281), .dout(n5285));
  jand g05030(.dina(n5285), .dinb(n5280), .dout(n5286));
  jxor g05031(.dina(n5286), .dinb(a41 ), .dout(n5287));
  jnot g05032(.din(n5287), .dout(n5288));
  jand g05033(.dina(n5109), .dinb(a44 ), .dout(n5289));
  jxor g05034(.dina(a44 ), .dinb(a43 ), .dout(n5290));
  jnot g05035(.din(n5290), .dout(n5291));
  jand g05036(.dina(n5291), .dinb(n5108), .dout(n5292));
  jand g05037(.dina(n5292), .dinb(b1 ), .dout(n5293));
  jnot g05038(.din(n5108), .dout(n5294));
  jxor g05039(.dina(a43 ), .dinb(a42 ), .dout(n5295));
  jand g05040(.dina(n5295), .dinb(n5294), .dout(n5296));
  jand g05041(.dina(n5296), .dinb(b0 ), .dout(n5297));
  jand g05042(.dina(n5290), .dinb(n5108), .dout(n5298));
  jand g05043(.dina(n5298), .dinb(n338), .dout(n5299));
  jor  g05044(.dina(n5299), .dinb(n5297), .dout(n5300));
  jor  g05045(.dina(n5300), .dinb(n5293), .dout(n5301));
  jxor g05046(.dina(n5301), .dinb(n5289), .dout(n5302));
  jxor g05047(.dina(n5302), .dinb(n5288), .dout(n5303));
  jxor g05048(.dina(n5303), .dinb(n5279), .dout(n5304));
  jnot g05049(.din(n5304), .dout(n5305));
  jor  g05050(.dina(n4415), .dinb(n428), .dout(n5306));
  jor  g05051(.dina(n4272), .dinb(n357), .dout(n5307));
  jor  g05052(.dina(n4418), .dinb(n395), .dout(n5308));
  jor  g05053(.dina(n4420), .dinb(n431), .dout(n5309));
  jand g05054(.dina(n5309), .dinb(n5308), .dout(n5310));
  jand g05055(.dina(n5310), .dinb(n5307), .dout(n5311));
  jand g05056(.dina(n5311), .dinb(n5306), .dout(n5312));
  jxor g05057(.dina(n5312), .dinb(a38 ), .dout(n5313));
  jxor g05058(.dina(n5313), .dinb(n5305), .dout(n5314));
  jxor g05059(.dina(n5314), .dinb(n5275), .dout(n5315));
  jnot g05060(.din(n5315), .dout(n5316));
  jor  g05061(.dina(n3849), .dinb(n624), .dout(n5317));
  jor  g05062(.dina(n3689), .dinb(n512), .dout(n5318));
  jor  g05063(.dina(n3852), .dinb(n564), .dout(n5319));
  jor  g05064(.dina(n3854), .dinb(n627), .dout(n5320));
  jand g05065(.dina(n5320), .dinb(n5319), .dout(n5321));
  jand g05066(.dina(n5321), .dinb(n5318), .dout(n5322));
  jand g05067(.dina(n5322), .dinb(n5317), .dout(n5323));
  jxor g05068(.dina(n5323), .dinb(a35 ), .dout(n5324));
  jxor g05069(.dina(n5324), .dinb(n5316), .dout(n5325));
  jxor g05070(.dina(n5325), .dinb(n5270), .dout(n5326));
  jxor g05071(.dina(n5326), .dinb(n5265), .dout(n5327));
  jxor g05072(.dina(n5327), .dinb(n5256), .dout(n5328));
  jnot g05073(.din(n5328), .dout(n5329));
  jor  g05074(.dina(n2784), .dinb(n1019), .dout(n5330));
  jor  g05075(.dina(n2661), .dinb(n858), .dout(n5331));
  jor  g05076(.dina(n2787), .dinb(n939), .dout(n5332));
  jor  g05077(.dina(n2789), .dinb(n1022), .dout(n5333));
  jand g05078(.dina(n5333), .dinb(n5332), .dout(n5334));
  jand g05079(.dina(n5334), .dinb(n5331), .dout(n5335));
  jand g05080(.dina(n5335), .dinb(n5330), .dout(n5336));
  jxor g05081(.dina(n5336), .dinb(a29 ), .dout(n5337));
  jxor g05082(.dina(n5337), .dinb(n5329), .dout(n5338));
  jxor g05083(.dina(n5338), .dinb(n5253), .dout(n5339));
  jnot g05084(.din(n5339), .dout(n5340));
  jor  g05085(.dina(n2319), .dinb(n1397), .dout(n5341));
  jor  g05086(.dina(n2224), .dinb(n1193), .dout(n5342));
  jor  g05087(.dina(n2322), .dinb(n1290), .dout(n5343));
  jor  g05088(.dina(n2324), .dinb(n1400), .dout(n5344));
  jand g05089(.dina(n5344), .dinb(n5343), .dout(n5345));
  jand g05090(.dina(n5345), .dinb(n5342), .dout(n5346));
  jand g05091(.dina(n5346), .dinb(n5341), .dout(n5347));
  jxor g05092(.dina(n5347), .dinb(a26 ), .dout(n5348));
  jxor g05093(.dina(n5348), .dinb(n5340), .dout(n5349));
  jxor g05094(.dina(n5349), .dinb(n5250), .dout(n5350));
  jnot g05095(.din(n5350), .dout(n5351));
  jor  g05096(.dina(n1739), .dinb(n1939), .dout(n5352));
  jor  g05097(.dina(n1827), .dinb(n1420), .dout(n5353));
  jor  g05098(.dina(n1942), .dinb(n1620), .dout(n5354));
  jor  g05099(.dina(n1944), .dinb(n1742), .dout(n5355));
  jand g05100(.dina(n5355), .dinb(n5354), .dout(n5356));
  jand g05101(.dina(n5356), .dinb(n5353), .dout(n5357));
  jand g05102(.dina(n5357), .dinb(n5352), .dout(n5358));
  jxor g05103(.dina(n5358), .dinb(a23 ), .dout(n5359));
  jxor g05104(.dina(n5359), .dinb(n5351), .dout(n5360));
  jxor g05105(.dina(n5360), .dinb(n5247), .dout(n5361));
  jor  g05106(.dina(n2007), .dinb(n1566), .dout(n5362));
  jor  g05107(.dina(n1489), .dinb(n1867), .dout(n5363));
  jor  g05108(.dina(n1569), .dinb(n1887), .dout(n5364));
  jor  g05109(.dina(n1571), .dinb(n2010), .dout(n5365));
  jand g05110(.dina(n5365), .dinb(n5364), .dout(n5366));
  jand g05111(.dina(n5366), .dinb(n5363), .dout(n5367));
  jand g05112(.dina(n5367), .dinb(n5362), .dout(n5368));
  jxor g05113(.dina(n5368), .dinb(a20 ), .dout(n5369));
  jxor g05114(.dina(n5369), .dinb(n5361), .dout(n5370));
  jnot g05115(.din(n5370), .dout(n5371));
  jxor g05116(.dina(n5371), .dinb(n5243), .dout(n5372));
  jxor g05117(.dina(n5372), .dinb(n5237), .dout(n5373));
  jxor g05118(.dina(n5373), .dinb(n5228), .dout(n5374));
  jxor g05119(.dina(n5374), .dinb(n5224), .dout(n5375));
  jxor g05120(.dina(n5375), .dinb(n5215), .dout(n5376));
  jor  g05121(.dina(n3400), .dinb(n706), .dout(n5377));
  jor  g05122(.dina(n683), .dinb(n3055), .dout(n5378));
  jor  g05123(.dina(n709), .dinb(n3230), .dout(n5379));
  jor  g05124(.dina(n711), .dinb(n3403), .dout(n5380));
  jand g05125(.dina(n5380), .dinb(n5379), .dout(n5381));
  jand g05126(.dina(n5381), .dinb(n5378), .dout(n5382));
  jand g05127(.dina(n5382), .dinb(n5377), .dout(n5383));
  jxor g05128(.dina(n5383), .dinb(a11 ), .dout(n5384));
  jxor g05129(.dina(n5384), .dinb(n5376), .dout(n5385));
  jxor g05130(.dina(n5385), .dinb(n5212), .dout(n5386));
  jnot g05131(.din(n5386), .dout(n5387));
  jor  g05132(.dina(n4137), .dinb(n528), .dout(n5388));
  jor  g05133(.dina(n490), .dinb(n3588), .dout(n5389));
  jor  g05134(.dina(n531), .dinb(n3942), .dout(n5390));
  jor  g05135(.dina(n533), .dinb(n4140), .dout(n5391));
  jand g05136(.dina(n5391), .dinb(n5390), .dout(n5392));
  jand g05137(.dina(n5392), .dinb(n5389), .dout(n5393));
  jand g05138(.dina(n5393), .dinb(n5388), .dout(n5394));
  jxor g05139(.dina(n5394), .dinb(a8 ), .dout(n5395));
  jxor g05140(.dina(n5395), .dinb(n5387), .dout(n5396));
  jxor g05141(.dina(n5396), .dinb(n5208), .dout(n5397));
  jxor g05142(.dina(n5397), .dinb(n5205), .dout(n5398));
  jxor g05143(.dina(n5398), .dinb(n5196), .dout(n5399));
  jand g05144(.dina(b42 ), .dinb(b41 ), .dout(n5400));
  jand g05145(.dina(n4989), .dinb(n4988), .dout(n5401));
  jor  g05146(.dina(n5401), .dinb(n5400), .dout(n5402));
  jxor g05147(.dina(b43 ), .dinb(b42 ), .dout(n5403));
  jnot g05148(.din(n5403), .dout(n5404));
  jxor g05149(.dina(n5404), .dinb(n5402), .dout(n5405));
  jor  g05150(.dina(n5405), .dinb(n264), .dout(n5406));
  jor  g05151(.dina(n284), .dinb(n4974), .dout(n5407));
  jnot g05152(.din(b43 ), .dout(n5408));
  jor  g05153(.dina(n269), .dinb(n5408), .dout(n5409));
  jor  g05154(.dina(n271), .dinb(n4994), .dout(n5410));
  jand g05155(.dina(n5410), .dinb(n5409), .dout(n5411));
  jand g05156(.dina(n5411), .dinb(n5407), .dout(n5412));
  jand g05157(.dina(n5412), .dinb(n5406), .dout(n5413));
  jxor g05158(.dina(n5413), .dinb(n260), .dout(n5414));
  jxor g05159(.dina(n5414), .dinb(n5399), .dout(n5415));
  jxor g05160(.dina(n5415), .dinb(n5193), .dout(f43 ));
  jand g05161(.dina(n5414), .dinb(n5399), .dout(n5417));
  jand g05162(.dina(n5415), .dinb(n5193), .dout(n5418));
  jor  g05163(.dina(n5418), .dinb(n5417), .dout(n5419));
  jand g05164(.dina(b43 ), .dinb(b42 ), .dout(n5420));
  jand g05165(.dina(n5403), .dinb(n5402), .dout(n5421));
  jor  g05166(.dina(n5421), .dinb(n5420), .dout(n5422));
  jxor g05167(.dina(b44 ), .dinb(b43 ), .dout(n5423));
  jnot g05168(.din(n5423), .dout(n5424));
  jxor g05169(.dina(n5424), .dinb(n5422), .dout(n5425));
  jor  g05170(.dina(n5425), .dinb(n264), .dout(n5426));
  jor  g05171(.dina(n284), .dinb(n4994), .dout(n5427));
  jnot g05172(.din(b44 ), .dout(n5428));
  jor  g05173(.dina(n269), .dinb(n5428), .dout(n5429));
  jor  g05174(.dina(n271), .dinb(n5408), .dout(n5430));
  jand g05175(.dina(n5430), .dinb(n5429), .dout(n5431));
  jand g05176(.dina(n5431), .dinb(n5427), .dout(n5432));
  jand g05177(.dina(n5432), .dinb(n5426), .dout(n5433));
  jxor g05178(.dina(n5433), .dinb(n260), .dout(n5434));
  jand g05179(.dina(n5397), .dinb(n5205), .dout(n5435));
  jand g05180(.dina(n5398), .dinb(n5196), .dout(n5436));
  jor  g05181(.dina(n5436), .dinb(n5435), .dout(n5437));
  jor  g05182(.dina(n4971), .dinb(n402), .dout(n5438));
  jor  g05183(.dina(n371), .dinb(n4537), .dout(n5439));
  jor  g05184(.dina(n405), .dinb(n4557), .dout(n5440));
  jor  g05185(.dina(n332), .dinb(n4974), .dout(n5441));
  jand g05186(.dina(n5441), .dinb(n5440), .dout(n5442));
  jand g05187(.dina(n5442), .dinb(n5439), .dout(n5443));
  jand g05188(.dina(n5443), .dinb(n5438), .dout(n5444));
  jxor g05189(.dina(n5444), .dinb(a5 ), .dout(n5445));
  jnot g05190(.din(n5445), .dout(n5446));
  jor  g05191(.dina(n5395), .dinb(n5387), .dout(n5447));
  jnot g05192(.din(n5447), .dout(n5448));
  jand g05193(.dina(n5396), .dinb(n5208), .dout(n5449));
  jor  g05194(.dina(n5449), .dinb(n5448), .dout(n5450));
  jnot g05195(.din(n5376), .dout(n5451));
  jor  g05196(.dina(n5384), .dinb(n5451), .dout(n5452));
  jor  g05197(.dina(n5385), .dinb(n5212), .dout(n5453));
  jand g05198(.dina(n5453), .dinb(n5452), .dout(n5454));
  jand g05199(.dina(n5374), .dinb(n5224), .dout(n5455));
  jand g05200(.dina(n5375), .dinb(n5215), .dout(n5456));
  jor  g05201(.dina(n5456), .dinb(n5455), .dout(n5457));
  jor  g05202(.dina(n3052), .dinb(n974), .dout(n5458));
  jor  g05203(.dina(n908), .dinb(n2870), .dout(n5459));
  jor  g05204(.dina(n977), .dinb(n3035), .dout(n5460));
  jor  g05205(.dina(n979), .dinb(n3055), .dout(n5461));
  jand g05206(.dina(n5461), .dinb(n5460), .dout(n5462));
  jand g05207(.dina(n5462), .dinb(n5459), .dout(n5463));
  jand g05208(.dina(n5463), .dinb(n5458), .dout(n5464));
  jxor g05209(.dina(n5464), .dinb(a14 ), .dout(n5465));
  jnot g05210(.din(n5465), .dout(n5466));
  jand g05211(.dina(n5372), .dinb(n5237), .dout(n5467));
  jand g05212(.dina(n5373), .dinb(n5228), .dout(n5468));
  jor  g05213(.dina(n5468), .dinb(n5467), .dout(n5469));
  jor  g05214(.dina(n2576), .dinb(n1245), .dout(n5470));
  jor  g05215(.dina(n1165), .dinb(n2407), .dout(n5471));
  jor  g05216(.dina(n1248), .dinb(n2559), .dout(n5472));
  jor  g05217(.dina(n1250), .dinb(n2579), .dout(n5473));
  jand g05218(.dina(n5473), .dinb(n5472), .dout(n5474));
  jand g05219(.dina(n5474), .dinb(n5471), .dout(n5475));
  jand g05220(.dina(n5475), .dinb(n5470), .dout(n5476));
  jxor g05221(.dina(n5476), .dinb(a17 ), .dout(n5477));
  jnot g05222(.din(n5477), .dout(n5478));
  jnot g05223(.din(n5361), .dout(n5479));
  jor  g05224(.dina(n5369), .dinb(n5479), .dout(n5480));
  jnot g05225(.din(n5480), .dout(n5481));
  jand g05226(.dina(n5371), .dinb(n5243), .dout(n5482));
  jor  g05227(.dina(n5482), .dinb(n5481), .dout(n5483));
  jor  g05228(.dina(n2145), .dinb(n1566), .dout(n5484));
  jor  g05229(.dina(n1489), .dinb(n1887), .dout(n5485));
  jor  g05230(.dina(n1569), .dinb(n2010), .dout(n5486));
  jor  g05231(.dina(n1571), .dinb(n2148), .dout(n5487));
  jand g05232(.dina(n5487), .dinb(n5486), .dout(n5488));
  jand g05233(.dina(n5488), .dinb(n5485), .dout(n5489));
  jand g05234(.dina(n5489), .dinb(n5484), .dout(n5490));
  jxor g05235(.dina(n5490), .dinb(a20 ), .dout(n5491));
  jnot g05236(.din(n5491), .dout(n5492));
  jor  g05237(.dina(n5359), .dinb(n5351), .dout(n5493));
  jnot g05238(.din(n5493), .dout(n5494));
  jand g05239(.dina(n5360), .dinb(n5247), .dout(n5495));
  jor  g05240(.dina(n5495), .dinb(n5494), .dout(n5496));
  jor  g05241(.dina(n5348), .dinb(n5340), .dout(n5497));
  jand g05242(.dina(n5349), .dinb(n5250), .dout(n5498));
  jnot g05243(.din(n5498), .dout(n5499));
  jand g05244(.dina(n5499), .dinb(n5497), .dout(n5500));
  jnot g05245(.din(n5500), .dout(n5501));
  jor  g05246(.dina(n5337), .dinb(n5329), .dout(n5502));
  jand g05247(.dina(n5338), .dinb(n5253), .dout(n5503));
  jnot g05248(.din(n5503), .dout(n5504));
  jand g05249(.dina(n5504), .dinb(n5502), .dout(n5505));
  jnot g05250(.din(n5505), .dout(n5506));
  jor  g05251(.dina(n2784), .dinb(n1190), .dout(n5507));
  jor  g05252(.dina(n2661), .dinb(n939), .dout(n5508));
  jor  g05253(.dina(n2787), .dinb(n1022), .dout(n5509));
  jor  g05254(.dina(n2789), .dinb(n1193), .dout(n5510));
  jand g05255(.dina(n5510), .dinb(n5509), .dout(n5511));
  jand g05256(.dina(n5511), .dinb(n5508), .dout(n5512));
  jand g05257(.dina(n5512), .dinb(n5507), .dout(n5513));
  jxor g05258(.dina(n5513), .dinb(a29 ), .dout(n5514));
  jnot g05259(.din(n5514), .dout(n5515));
  jand g05260(.dina(n5326), .dinb(n5265), .dout(n5516));
  jand g05261(.dina(n5327), .dinb(n5256), .dout(n5517));
  jor  g05262(.dina(n5517), .dinb(n5516), .dout(n5518));
  jor  g05263(.dina(n3301), .dinb(n855), .dout(n5519));
  jor  g05264(.dina(n3136), .dinb(n758), .dout(n5520));
  jor  g05265(.dina(n3304), .dinb(n778), .dout(n5521));
  jor  g05266(.dina(n3306), .dinb(n858), .dout(n5522));
  jand g05267(.dina(n5522), .dinb(n5521), .dout(n5523));
  jand g05268(.dina(n5523), .dinb(n5520), .dout(n5524));
  jand g05269(.dina(n5524), .dinb(n5519), .dout(n5525));
  jxor g05270(.dina(n5525), .dinb(a32 ), .dout(n5526));
  jnot g05271(.din(n5526), .dout(n5527));
  jor  g05272(.dina(n5324), .dinb(n5316), .dout(n5528));
  jand g05273(.dina(n5325), .dinb(n5270), .dout(n5529));
  jnot g05274(.din(n5529), .dout(n5530));
  jand g05275(.dina(n5530), .dinb(n5528), .dout(n5531));
  jnot g05276(.din(n5531), .dout(n5532));
  jor  g05277(.dina(n3849), .dinb(n644), .dout(n5533));
  jor  g05278(.dina(n3689), .dinb(n564), .dout(n5534));
  jor  g05279(.dina(n3852), .dinb(n627), .dout(n5535));
  jor  g05280(.dina(n3854), .dinb(n647), .dout(n5536));
  jand g05281(.dina(n5536), .dinb(n5535), .dout(n5537));
  jand g05282(.dina(n5537), .dinb(n5534), .dout(n5538));
  jand g05283(.dina(n5538), .dinb(n5533), .dout(n5539));
  jxor g05284(.dina(n5539), .dinb(a35 ), .dout(n5540));
  jnot g05285(.din(n5540), .dout(n5541));
  jor  g05286(.dina(n5313), .dinb(n5305), .dout(n5542));
  jand g05287(.dina(n5314), .dinb(n5275), .dout(n5543));
  jnot g05288(.din(n5543), .dout(n5544));
  jand g05289(.dina(n5544), .dinb(n5542), .dout(n5545));
  jnot g05290(.din(n5545), .dout(n5546));
  jor  g05291(.dina(n4415), .dinb(n509), .dout(n5547));
  jor  g05292(.dina(n4272), .dinb(n395), .dout(n5548));
  jor  g05293(.dina(n4418), .dinb(n431), .dout(n5549));
  jor  g05294(.dina(n4420), .dinb(n512), .dout(n5550));
  jand g05295(.dina(n5550), .dinb(n5549), .dout(n5551));
  jand g05296(.dina(n5551), .dinb(n5548), .dout(n5552));
  jand g05297(.dina(n5552), .dinb(n5547), .dout(n5553));
  jxor g05298(.dina(n5553), .dinb(a38 ), .dout(n5554));
  jnot g05299(.din(n5554), .dout(n5555));
  jand g05300(.dina(n5302), .dinb(n5288), .dout(n5556));
  jand g05301(.dina(n5303), .dinb(n5279), .dout(n5557));
  jor  g05302(.dina(n5557), .dinb(n5556), .dout(n5558));
  jor  g05303(.dina(n5096), .dinb(n354), .dout(n5559));
  jor  g05304(.dina(n4904), .dinb(n299), .dout(n5560));
  jor  g05305(.dina(n5099), .dinb(n322), .dout(n5561));
  jor  g05306(.dina(n5101), .dinb(n357), .dout(n5562));
  jand g05307(.dina(n5562), .dinb(n5561), .dout(n5563));
  jand g05308(.dina(n5563), .dinb(n5560), .dout(n5564));
  jand g05309(.dina(n5564), .dinb(n5559), .dout(n5565));
  jxor g05310(.dina(n5565), .dinb(a41 ), .dout(n5566));
  jnot g05311(.din(n5566), .dout(n5567));
  jnot g05312(.din(n5301), .dout(n5568));
  jand g05313(.dina(n5110), .dinb(a44 ), .dout(n5569));
  jand g05314(.dina(n5569), .dinb(n5568), .dout(n5570));
  jnot g05315(.din(n5570), .dout(n5571));
  jand g05316(.dina(n5571), .dinb(a44 ), .dout(n5572));
  jor  g05317(.dina(n5295), .dinb(n5291), .dout(n5573));
  jor  g05318(.dina(n5573), .dinb(n5108), .dout(n5574));
  jnot g05319(.din(n5574), .dout(n5575));
  jand g05320(.dina(n5575), .dinb(b0 ), .dout(n5576));
  jand g05321(.dina(n5292), .dinb(b2 ), .dout(n5577));
  jand g05322(.dina(n5296), .dinb(b1 ), .dout(n5578));
  jand g05323(.dina(n5298), .dinb(n375), .dout(n5579));
  jor  g05324(.dina(n5579), .dinb(n5578), .dout(n5580));
  jor  g05325(.dina(n5580), .dinb(n5577), .dout(n5581));
  jor  g05326(.dina(n5581), .dinb(n5576), .dout(n5582));
  jxor g05327(.dina(n5582), .dinb(n5572), .dout(n5583));
  jxor g05328(.dina(n5583), .dinb(n5567), .dout(n5584));
  jxor g05329(.dina(n5584), .dinb(n5558), .dout(n5585));
  jxor g05330(.dina(n5585), .dinb(n5555), .dout(n5586));
  jxor g05331(.dina(n5586), .dinb(n5546), .dout(n5587));
  jxor g05332(.dina(n5587), .dinb(n5541), .dout(n5588));
  jxor g05333(.dina(n5588), .dinb(n5532), .dout(n5589));
  jxor g05334(.dina(n5589), .dinb(n5527), .dout(n5590));
  jxor g05335(.dina(n5590), .dinb(n5518), .dout(n5591));
  jxor g05336(.dina(n5591), .dinb(n5515), .dout(n5592));
  jxor g05337(.dina(n5592), .dinb(n5506), .dout(n5593));
  jnot g05338(.din(n5593), .dout(n5594));
  jor  g05339(.dina(n2319), .dinb(n1417), .dout(n5595));
  jor  g05340(.dina(n2224), .dinb(n1290), .dout(n5596));
  jor  g05341(.dina(n2322), .dinb(n1400), .dout(n5597));
  jor  g05342(.dina(n2324), .dinb(n1420), .dout(n5598));
  jand g05343(.dina(n5598), .dinb(n5597), .dout(n5599));
  jand g05344(.dina(n5599), .dinb(n5596), .dout(n5600));
  jand g05345(.dina(n5600), .dinb(n5595), .dout(n5601));
  jxor g05346(.dina(n5601), .dinb(a26 ), .dout(n5602));
  jxor g05347(.dina(n5602), .dinb(n5594), .dout(n5603));
  jxor g05348(.dina(n5603), .dinb(n5501), .dout(n5604));
  jnot g05349(.din(n5604), .dout(n5605));
  jor  g05350(.dina(n1864), .dinb(n1939), .dout(n5606));
  jor  g05351(.dina(n1827), .dinb(n1620), .dout(n5607));
  jor  g05352(.dina(n1942), .dinb(n1742), .dout(n5608));
  jor  g05353(.dina(n1944), .dinb(n1867), .dout(n5609));
  jand g05354(.dina(n5609), .dinb(n5608), .dout(n5610));
  jand g05355(.dina(n5610), .dinb(n5607), .dout(n5611));
  jand g05356(.dina(n5611), .dinb(n5606), .dout(n5612));
  jxor g05357(.dina(n5612), .dinb(a23 ), .dout(n5613));
  jxor g05358(.dina(n5613), .dinb(n5605), .dout(n5614));
  jxor g05359(.dina(n5614), .dinb(n5496), .dout(n5615));
  jxor g05360(.dina(n5615), .dinb(n5492), .dout(n5616));
  jxor g05361(.dina(n5616), .dinb(n5483), .dout(n5617));
  jxor g05362(.dina(n5617), .dinb(n5478), .dout(n5618));
  jxor g05363(.dina(n5618), .dinb(n5469), .dout(n5619));
  jxor g05364(.dina(n5619), .dinb(n5466), .dout(n5620));
  jxor g05365(.dina(n5620), .dinb(n5457), .dout(n5621));
  jor  g05366(.dina(n3585), .dinb(n706), .dout(n5622));
  jor  g05367(.dina(n683), .dinb(n3230), .dout(n5623));
  jor  g05368(.dina(n709), .dinb(n3403), .dout(n5624));
  jor  g05369(.dina(n711), .dinb(n3588), .dout(n5625));
  jand g05370(.dina(n5625), .dinb(n5624), .dout(n5626));
  jand g05371(.dina(n5626), .dinb(n5623), .dout(n5627));
  jand g05372(.dina(n5627), .dinb(n5622), .dout(n5628));
  jxor g05373(.dina(n5628), .dinb(a11 ), .dout(n5629));
  jxor g05374(.dina(n5629), .dinb(n5621), .dout(n5630));
  jxor g05375(.dina(n5630), .dinb(n5454), .dout(n5631));
  jnot g05376(.din(n5631), .dout(n5632));
  jor  g05377(.dina(n4337), .dinb(n528), .dout(n5633));
  jor  g05378(.dina(n490), .dinb(n3942), .dout(n5634));
  jor  g05379(.dina(n531), .dinb(n4140), .dout(n5635));
  jor  g05380(.dina(n533), .dinb(n4340), .dout(n5636));
  jand g05381(.dina(n5636), .dinb(n5635), .dout(n5637));
  jand g05382(.dina(n5637), .dinb(n5634), .dout(n5638));
  jand g05383(.dina(n5638), .dinb(n5633), .dout(n5639));
  jxor g05384(.dina(n5639), .dinb(a8 ), .dout(n5640));
  jxor g05385(.dina(n5640), .dinb(n5632), .dout(n5641));
  jxor g05386(.dina(n5641), .dinb(n5450), .dout(n5642));
  jxor g05387(.dina(n5642), .dinb(n5446), .dout(n5643));
  jxor g05388(.dina(n5643), .dinb(n5437), .dout(n5644));
  jxor g05389(.dina(n5644), .dinb(n5434), .dout(n5645));
  jxor g05390(.dina(n5645), .dinb(n5419), .dout(f44 ));
  jand g05391(.dina(n5644), .dinb(n5434), .dout(n5647));
  jand g05392(.dina(n5645), .dinb(n5419), .dout(n5648));
  jor  g05393(.dina(n5648), .dinb(n5647), .dout(n5649));
  jand g05394(.dina(n5642), .dinb(n5446), .dout(n5650));
  jand g05395(.dina(n5643), .dinb(n5437), .dout(n5651));
  jor  g05396(.dina(n5651), .dinb(n5650), .dout(n5652));
  jor  g05397(.dina(n5640), .dinb(n5632), .dout(n5653));
  jnot g05398(.din(n5653), .dout(n5654));
  jand g05399(.dina(n5641), .dinb(n5450), .dout(n5655));
  jor  g05400(.dina(n5655), .dinb(n5654), .dout(n5656));
  jnot g05401(.din(n5656), .dout(n5657));
  jnot g05402(.din(n5621), .dout(n5658));
  jor  g05403(.dina(n5629), .dinb(n5658), .dout(n5659));
  jor  g05404(.dina(n5630), .dinb(n5454), .dout(n5660));
  jand g05405(.dina(n5660), .dinb(n5659), .dout(n5661));
  jor  g05406(.dina(n3939), .dinb(n706), .dout(n5662));
  jor  g05407(.dina(n683), .dinb(n3403), .dout(n5663));
  jor  g05408(.dina(n709), .dinb(n3588), .dout(n5664));
  jor  g05409(.dina(n711), .dinb(n3942), .dout(n5665));
  jand g05410(.dina(n5665), .dinb(n5664), .dout(n5666));
  jand g05411(.dina(n5666), .dinb(n5663), .dout(n5667));
  jand g05412(.dina(n5667), .dinb(n5662), .dout(n5668));
  jxor g05413(.dina(n5668), .dinb(a11 ), .dout(n5669));
  jand g05414(.dina(n5619), .dinb(n5466), .dout(n5670));
  jand g05415(.dina(n5620), .dinb(n5457), .dout(n5671));
  jor  g05416(.dina(n5671), .dinb(n5670), .dout(n5672));
  jand g05417(.dina(n5617), .dinb(n5478), .dout(n5673));
  jand g05418(.dina(n5618), .dinb(n5469), .dout(n5674));
  jor  g05419(.dina(n5674), .dinb(n5673), .dout(n5675));
  jor  g05420(.dina(n2867), .dinb(n1245), .dout(n5676));
  jor  g05421(.dina(n1165), .dinb(n2559), .dout(n5677));
  jor  g05422(.dina(n1248), .dinb(n2579), .dout(n5678));
  jor  g05423(.dina(n1250), .dinb(n2870), .dout(n5679));
  jand g05424(.dina(n5679), .dinb(n5678), .dout(n5680));
  jand g05425(.dina(n5680), .dinb(n5677), .dout(n5681));
  jand g05426(.dina(n5681), .dinb(n5676), .dout(n5682));
  jxor g05427(.dina(n5682), .dinb(a17 ), .dout(n5683));
  jnot g05428(.din(n5683), .dout(n5684));
  jand g05429(.dina(n5615), .dinb(n5492), .dout(n5685));
  jand g05430(.dina(n5616), .dinb(n5483), .dout(n5686));
  jor  g05431(.dina(n5686), .dinb(n5685), .dout(n5687));
  jor  g05432(.dina(n5613), .dinb(n5605), .dout(n5688));
  jnot g05433(.din(n5688), .dout(n5689));
  jand g05434(.dina(n5614), .dinb(n5496), .dout(n5690));
  jor  g05435(.dina(n5690), .dinb(n5689), .dout(n5691));
  jor  g05436(.dina(n5602), .dinb(n5594), .dout(n5692));
  jand g05437(.dina(n5603), .dinb(n5501), .dout(n5693));
  jnot g05438(.din(n5693), .dout(n5694));
  jand g05439(.dina(n5694), .dinb(n5692), .dout(n5695));
  jnot g05440(.din(n5695), .dout(n5696));
  jand g05441(.dina(n5591), .dinb(n5515), .dout(n5697));
  jand g05442(.dina(n5592), .dinb(n5506), .dout(n5698));
  jor  g05443(.dina(n5698), .dinb(n5697), .dout(n5699));
  jor  g05444(.dina(n2784), .dinb(n1287), .dout(n5700));
  jor  g05445(.dina(n2661), .dinb(n1022), .dout(n5701));
  jor  g05446(.dina(n2787), .dinb(n1193), .dout(n5702));
  jor  g05447(.dina(n2789), .dinb(n1290), .dout(n5703));
  jand g05448(.dina(n5703), .dinb(n5702), .dout(n5704));
  jand g05449(.dina(n5704), .dinb(n5701), .dout(n5705));
  jand g05450(.dina(n5705), .dinb(n5700), .dout(n5706));
  jxor g05451(.dina(n5706), .dinb(a29 ), .dout(n5707));
  jnot g05452(.din(n5707), .dout(n5708));
  jand g05453(.dina(n5589), .dinb(n5527), .dout(n5709));
  jand g05454(.dina(n5590), .dinb(n5518), .dout(n5710));
  jor  g05455(.dina(n5710), .dinb(n5709), .dout(n5711));
  jor  g05456(.dina(n3301), .dinb(n936), .dout(n5712));
  jor  g05457(.dina(n3136), .dinb(n778), .dout(n5713));
  jor  g05458(.dina(n3304), .dinb(n858), .dout(n5714));
  jor  g05459(.dina(n3306), .dinb(n939), .dout(n5715));
  jand g05460(.dina(n5715), .dinb(n5714), .dout(n5716));
  jand g05461(.dina(n5716), .dinb(n5713), .dout(n5717));
  jand g05462(.dina(n5717), .dinb(n5712), .dout(n5718));
  jxor g05463(.dina(n5718), .dinb(a32 ), .dout(n5719));
  jnot g05464(.din(n5719), .dout(n5720));
  jand g05465(.dina(n5587), .dinb(n5541), .dout(n5721));
  jand g05466(.dina(n5588), .dinb(n5532), .dout(n5722));
  jor  g05467(.dina(n5722), .dinb(n5721), .dout(n5723));
  jor  g05468(.dina(n3849), .dinb(n755), .dout(n5724));
  jor  g05469(.dina(n3689), .dinb(n627), .dout(n5725));
  jor  g05470(.dina(n3852), .dinb(n647), .dout(n5726));
  jor  g05471(.dina(n3854), .dinb(n758), .dout(n5727));
  jand g05472(.dina(n5727), .dinb(n5726), .dout(n5728));
  jand g05473(.dina(n5728), .dinb(n5725), .dout(n5729));
  jand g05474(.dina(n5729), .dinb(n5724), .dout(n5730));
  jxor g05475(.dina(n5730), .dinb(a35 ), .dout(n5731));
  jnot g05476(.din(n5731), .dout(n5732));
  jand g05477(.dina(n5585), .dinb(n5555), .dout(n5733));
  jand g05478(.dina(n5586), .dinb(n5546), .dout(n5734));
  jor  g05479(.dina(n5734), .dinb(n5733), .dout(n5735));
  jand g05480(.dina(n5583), .dinb(n5567), .dout(n5736));
  jand g05481(.dina(n5584), .dinb(n5558), .dout(n5737));
  jor  g05482(.dina(n5737), .dinb(n5736), .dout(n5738));
  jnot g05483(.din(n5298), .dout(n5739));
  jor  g05484(.dina(n5739), .dinb(n296), .dout(n5740));
  jor  g05485(.dina(n5574), .dinb(n267), .dout(n5741));
  jnot g05486(.din(n5296), .dout(n5742));
  jor  g05487(.dina(n5742), .dinb(n279), .dout(n5743));
  jnot g05488(.din(n5292), .dout(n5744));
  jor  g05489(.dina(n5744), .dinb(n299), .dout(n5745));
  jand g05490(.dina(n5745), .dinb(n5743), .dout(n5746));
  jand g05491(.dina(n5746), .dinb(n5741), .dout(n5747));
  jand g05492(.dina(n5747), .dinb(n5740), .dout(n5748));
  jxor g05493(.dina(n5748), .dinb(a44 ), .dout(n5749));
  jnot g05494(.din(n5749), .dout(n5750));
  jxor g05495(.dina(a45 ), .dinb(a44 ), .dout(n5751));
  jand g05496(.dina(n5751), .dinb(b0 ), .dout(n5752));
  jnot g05497(.din(n5752), .dout(n5753));
  jor  g05498(.dina(n5582), .dinb(n5571), .dout(n5754));
  jxor g05499(.dina(n5754), .dinb(n5753), .dout(n5755));
  jxor g05500(.dina(n5755), .dinb(n5750), .dout(n5756));
  jnot g05501(.din(n5756), .dout(n5757));
  jor  g05502(.dina(n5096), .dinb(n392), .dout(n5758));
  jor  g05503(.dina(n4904), .dinb(n322), .dout(n5759));
  jor  g05504(.dina(n5099), .dinb(n357), .dout(n5760));
  jor  g05505(.dina(n5101), .dinb(n395), .dout(n5761));
  jand g05506(.dina(n5761), .dinb(n5760), .dout(n5762));
  jand g05507(.dina(n5762), .dinb(n5759), .dout(n5763));
  jand g05508(.dina(n5763), .dinb(n5758), .dout(n5764));
  jxor g05509(.dina(n5764), .dinb(a41 ), .dout(n5765));
  jxor g05510(.dina(n5765), .dinb(n5757), .dout(n5766));
  jxor g05511(.dina(n5766), .dinb(n5738), .dout(n5767));
  jnot g05512(.din(n5767), .dout(n5768));
  jor  g05513(.dina(n4415), .dinb(n561), .dout(n5769));
  jor  g05514(.dina(n4272), .dinb(n431), .dout(n5770));
  jor  g05515(.dina(n4418), .dinb(n512), .dout(n5771));
  jor  g05516(.dina(n4420), .dinb(n564), .dout(n5772));
  jand g05517(.dina(n5772), .dinb(n5771), .dout(n5773));
  jand g05518(.dina(n5773), .dinb(n5770), .dout(n5774));
  jand g05519(.dina(n5774), .dinb(n5769), .dout(n5775));
  jxor g05520(.dina(n5775), .dinb(a38 ), .dout(n5776));
  jxor g05521(.dina(n5776), .dinb(n5768), .dout(n5777));
  jxor g05522(.dina(n5777), .dinb(n5735), .dout(n5778));
  jxor g05523(.dina(n5778), .dinb(n5732), .dout(n5779));
  jxor g05524(.dina(n5779), .dinb(n5723), .dout(n5780));
  jxor g05525(.dina(n5780), .dinb(n5720), .dout(n5781));
  jxor g05526(.dina(n5781), .dinb(n5711), .dout(n5782));
  jxor g05527(.dina(n5782), .dinb(n5708), .dout(n5783));
  jxor g05528(.dina(n5783), .dinb(n5699), .dout(n5784));
  jnot g05529(.din(n5784), .dout(n5785));
  jor  g05530(.dina(n2319), .dinb(n1617), .dout(n5786));
  jor  g05531(.dina(n2224), .dinb(n1400), .dout(n5787));
  jor  g05532(.dina(n2322), .dinb(n1420), .dout(n5788));
  jor  g05533(.dina(n2324), .dinb(n1620), .dout(n5789));
  jand g05534(.dina(n5789), .dinb(n5788), .dout(n5790));
  jand g05535(.dina(n5790), .dinb(n5787), .dout(n5791));
  jand g05536(.dina(n5791), .dinb(n5786), .dout(n5792));
  jxor g05537(.dina(n5792), .dinb(a26 ), .dout(n5793));
  jxor g05538(.dina(n5793), .dinb(n5785), .dout(n5794));
  jxor g05539(.dina(n5794), .dinb(n5696), .dout(n5795));
  jnot g05540(.din(n5795), .dout(n5796));
  jor  g05541(.dina(n1884), .dinb(n1939), .dout(n5797));
  jor  g05542(.dina(n1827), .dinb(n1742), .dout(n5798));
  jor  g05543(.dina(n1942), .dinb(n1867), .dout(n5799));
  jor  g05544(.dina(n1944), .dinb(n1887), .dout(n5800));
  jand g05545(.dina(n5800), .dinb(n5799), .dout(n5801));
  jand g05546(.dina(n5801), .dinb(n5798), .dout(n5802));
  jand g05547(.dina(n5802), .dinb(n5797), .dout(n5803));
  jxor g05548(.dina(n5803), .dinb(a23 ), .dout(n5804));
  jxor g05549(.dina(n5804), .dinb(n5796), .dout(n5805));
  jxor g05550(.dina(n5805), .dinb(n5691), .dout(n5806));
  jor  g05551(.dina(n2404), .dinb(n1566), .dout(n5807));
  jor  g05552(.dina(n1489), .dinb(n2010), .dout(n5808));
  jor  g05553(.dina(n1569), .dinb(n2148), .dout(n5809));
  jor  g05554(.dina(n1571), .dinb(n2407), .dout(n5810));
  jand g05555(.dina(n5810), .dinb(n5809), .dout(n5811));
  jand g05556(.dina(n5811), .dinb(n5808), .dout(n5812));
  jand g05557(.dina(n5812), .dinb(n5807), .dout(n5813));
  jxor g05558(.dina(n5813), .dinb(a20 ), .dout(n5814));
  jxor g05559(.dina(n5814), .dinb(n5806), .dout(n5815));
  jnot g05560(.din(n5815), .dout(n5816));
  jxor g05561(.dina(n5816), .dinb(n5687), .dout(n5817));
  jxor g05562(.dina(n5817), .dinb(n5684), .dout(n5818));
  jxor g05563(.dina(n5818), .dinb(n5675), .dout(n5819));
  jnot g05564(.din(n5819), .dout(n5820));
  jor  g05565(.dina(n3227), .dinb(n974), .dout(n5821));
  jor  g05566(.dina(n908), .dinb(n3035), .dout(n5822));
  jor  g05567(.dina(n977), .dinb(n3055), .dout(n5823));
  jor  g05568(.dina(n979), .dinb(n3230), .dout(n5824));
  jand g05569(.dina(n5824), .dinb(n5823), .dout(n5825));
  jand g05570(.dina(n5825), .dinb(n5822), .dout(n5826));
  jand g05571(.dina(n5826), .dinb(n5821), .dout(n5827));
  jxor g05572(.dina(n5827), .dinb(a14 ), .dout(n5828));
  jxor g05573(.dina(n5828), .dinb(n5820), .dout(n5829));
  jxor g05574(.dina(n5829), .dinb(n5672), .dout(n5830));
  jxor g05575(.dina(n5830), .dinb(n5669), .dout(n5831));
  jxor g05576(.dina(n5831), .dinb(n5661), .dout(n5832));
  jnot g05577(.din(n5832), .dout(n5833));
  jor  g05578(.dina(n4534), .dinb(n528), .dout(n5834));
  jor  g05579(.dina(n490), .dinb(n4140), .dout(n5835));
  jor  g05580(.dina(n531), .dinb(n4340), .dout(n5836));
  jor  g05581(.dina(n533), .dinb(n4537), .dout(n5837));
  jand g05582(.dina(n5837), .dinb(n5836), .dout(n5838));
  jand g05583(.dina(n5838), .dinb(n5835), .dout(n5839));
  jand g05584(.dina(n5839), .dinb(n5834), .dout(n5840));
  jxor g05585(.dina(n5840), .dinb(a8 ), .dout(n5841));
  jxor g05586(.dina(n5841), .dinb(n5833), .dout(n5842));
  jxor g05587(.dina(n5842), .dinb(n5657), .dout(n5843));
  jor  g05588(.dina(n4991), .dinb(n402), .dout(n5844));
  jor  g05589(.dina(n371), .dinb(n4557), .dout(n5845));
  jor  g05590(.dina(n405), .dinb(n4974), .dout(n5846));
  jor  g05591(.dina(n332), .dinb(n4994), .dout(n5847));
  jand g05592(.dina(n5847), .dinb(n5846), .dout(n5848));
  jand g05593(.dina(n5848), .dinb(n5845), .dout(n5849));
  jand g05594(.dina(n5849), .dinb(n5844), .dout(n5850));
  jxor g05595(.dina(n5850), .dinb(a5 ), .dout(n5851));
  jxor g05596(.dina(n5851), .dinb(n5843), .dout(n5852));
  jxor g05597(.dina(n5852), .dinb(n5652), .dout(n5853));
  jand g05598(.dina(b44 ), .dinb(b43 ), .dout(n5854));
  jand g05599(.dina(n5423), .dinb(n5422), .dout(n5855));
  jor  g05600(.dina(n5855), .dinb(n5854), .dout(n5856));
  jxor g05601(.dina(b45 ), .dinb(b44 ), .dout(n5857));
  jnot g05602(.din(n5857), .dout(n5858));
  jxor g05603(.dina(n5858), .dinb(n5856), .dout(n5859));
  jor  g05604(.dina(n5859), .dinb(n264), .dout(n5860));
  jor  g05605(.dina(n284), .dinb(n5408), .dout(n5861));
  jnot g05606(.din(b45 ), .dout(n5862));
  jor  g05607(.dina(n269), .dinb(n5862), .dout(n5863));
  jor  g05608(.dina(n271), .dinb(n5428), .dout(n5864));
  jand g05609(.dina(n5864), .dinb(n5863), .dout(n5865));
  jand g05610(.dina(n5865), .dinb(n5861), .dout(n5866));
  jand g05611(.dina(n5866), .dinb(n5860), .dout(n5867));
  jxor g05612(.dina(n5867), .dinb(n260), .dout(n5868));
  jxor g05613(.dina(n5868), .dinb(n5853), .dout(n5869));
  jxor g05614(.dina(n5869), .dinb(n5649), .dout(f45 ));
  jand g05615(.dina(n5868), .dinb(n5853), .dout(n5871));
  jand g05616(.dina(n5869), .dinb(n5649), .dout(n5872));
  jor  g05617(.dina(n5872), .dinb(n5871), .dout(n5873));
  jor  g05618(.dina(n5851), .dinb(n5843), .dout(n5874));
  jnot g05619(.din(n5874), .dout(n5875));
  jand g05620(.dina(n5852), .dinb(n5652), .dout(n5876));
  jor  g05621(.dina(n5876), .dinb(n5875), .dout(n5877));
  jor  g05622(.dina(n5841), .dinb(n5833), .dout(n5878));
  jnot g05623(.din(n5878), .dout(n5879));
  jand g05624(.dina(n5842), .dinb(n5656), .dout(n5880));
  jor  g05625(.dina(n5880), .dinb(n5879), .dout(n5881));
  jnot g05626(.din(n5881), .dout(n5882));
  jnot g05627(.din(n5669), .dout(n5883));
  jand g05628(.dina(n5830), .dinb(n5883), .dout(n5884));
  jnot g05629(.din(n5884), .dout(n5885));
  jor  g05630(.dina(n5831), .dinb(n5661), .dout(n5886));
  jand g05631(.dina(n5886), .dinb(n5885), .dout(n5887));
  jor  g05632(.dina(n5828), .dinb(n5820), .dout(n5888));
  jnot g05633(.din(n5888), .dout(n5889));
  jand g05634(.dina(n5829), .dinb(n5672), .dout(n5890));
  jor  g05635(.dina(n5890), .dinb(n5889), .dout(n5891));
  jand g05636(.dina(n5817), .dinb(n5684), .dout(n5892));
  jand g05637(.dina(n5818), .dinb(n5675), .dout(n5893));
  jor  g05638(.dina(n5893), .dinb(n5892), .dout(n5894));
  jor  g05639(.dina(n3032), .dinb(n1245), .dout(n5895));
  jor  g05640(.dina(n1165), .dinb(n2579), .dout(n5896));
  jor  g05641(.dina(n1248), .dinb(n2870), .dout(n5897));
  jor  g05642(.dina(n1250), .dinb(n3035), .dout(n5898));
  jand g05643(.dina(n5898), .dinb(n5897), .dout(n5899));
  jand g05644(.dina(n5899), .dinb(n5896), .dout(n5900));
  jand g05645(.dina(n5900), .dinb(n5895), .dout(n5901));
  jxor g05646(.dina(n5901), .dinb(a17 ), .dout(n5902));
  jnot g05647(.din(n5902), .dout(n5903));
  jnot g05648(.din(n5806), .dout(n5904));
  jor  g05649(.dina(n5814), .dinb(n5904), .dout(n5905));
  jnot g05650(.din(n5905), .dout(n5906));
  jand g05651(.dina(n5816), .dinb(n5687), .dout(n5907));
  jor  g05652(.dina(n5907), .dinb(n5906), .dout(n5908));
  jor  g05653(.dina(n2556), .dinb(n1566), .dout(n5909));
  jor  g05654(.dina(n1489), .dinb(n2148), .dout(n5910));
  jor  g05655(.dina(n1569), .dinb(n2407), .dout(n5911));
  jor  g05656(.dina(n1571), .dinb(n2559), .dout(n5912));
  jand g05657(.dina(n5912), .dinb(n5911), .dout(n5913));
  jand g05658(.dina(n5913), .dinb(n5910), .dout(n5914));
  jand g05659(.dina(n5914), .dinb(n5909), .dout(n5915));
  jxor g05660(.dina(n5915), .dinb(a20 ), .dout(n5916));
  jnot g05661(.din(n5916), .dout(n5917));
  jor  g05662(.dina(n5804), .dinb(n5796), .dout(n5918));
  jnot g05663(.din(n5918), .dout(n5919));
  jand g05664(.dina(n5805), .dinb(n5691), .dout(n5920));
  jor  g05665(.dina(n5920), .dinb(n5919), .dout(n5921));
  jor  g05666(.dina(n5793), .dinb(n5785), .dout(n5922));
  jand g05667(.dina(n5794), .dinb(n5696), .dout(n5923));
  jnot g05668(.din(n5923), .dout(n5924));
  jand g05669(.dina(n5924), .dinb(n5922), .dout(n5925));
  jnot g05670(.din(n5925), .dout(n5926));
  jand g05671(.dina(n5782), .dinb(n5708), .dout(n5927));
  jand g05672(.dina(n5783), .dinb(n5699), .dout(n5928));
  jor  g05673(.dina(n5928), .dinb(n5927), .dout(n5929));
  jand g05674(.dina(n5780), .dinb(n5720), .dout(n5930));
  jand g05675(.dina(n5781), .dinb(n5711), .dout(n5931));
  jor  g05676(.dina(n5931), .dinb(n5930), .dout(n5932));
  jand g05677(.dina(n5778), .dinb(n5732), .dout(n5933));
  jand g05678(.dina(n5779), .dinb(n5723), .dout(n5934));
  jor  g05679(.dina(n5934), .dinb(n5933), .dout(n5935));
  jor  g05680(.dina(n3849), .dinb(n775), .dout(n5936));
  jor  g05681(.dina(n3689), .dinb(n647), .dout(n5937));
  jor  g05682(.dina(n3852), .dinb(n758), .dout(n5938));
  jor  g05683(.dina(n3854), .dinb(n778), .dout(n5939));
  jand g05684(.dina(n5939), .dinb(n5938), .dout(n5940));
  jand g05685(.dina(n5940), .dinb(n5937), .dout(n5941));
  jand g05686(.dina(n5941), .dinb(n5936), .dout(n5942));
  jxor g05687(.dina(n5942), .dinb(a35 ), .dout(n5943));
  jnot g05688(.din(n5943), .dout(n5944));
  jor  g05689(.dina(n5776), .dinb(n5768), .dout(n5945));
  jand g05690(.dina(n5777), .dinb(n5735), .dout(n5946));
  jnot g05691(.din(n5946), .dout(n5947));
  jand g05692(.dina(n5947), .dinb(n5945), .dout(n5948));
  jnot g05693(.din(n5948), .dout(n5949));
  jor  g05694(.dina(n5765), .dinb(n5757), .dout(n5950));
  jand g05695(.dina(n5766), .dinb(n5738), .dout(n5951));
  jnot g05696(.din(n5951), .dout(n5952));
  jand g05697(.dina(n5952), .dinb(n5950), .dout(n5953));
  jnot g05698(.din(n5953), .dout(n5954));
  jnot g05699(.din(n5754), .dout(n5955));
  jand g05700(.dina(n5955), .dinb(n5752), .dout(n5956));
  jand g05701(.dina(n5755), .dinb(n5750), .dout(n5957));
  jor  g05702(.dina(n5957), .dinb(n5956), .dout(n5958));
  jor  g05703(.dina(n5739), .dinb(n319), .dout(n5959));
  jor  g05704(.dina(n5574), .dinb(n279), .dout(n5960));
  jor  g05705(.dina(n5742), .dinb(n299), .dout(n5961));
  jor  g05706(.dina(n5744), .dinb(n322), .dout(n5962));
  jand g05707(.dina(n5962), .dinb(n5961), .dout(n5963));
  jand g05708(.dina(n5963), .dinb(n5960), .dout(n5964));
  jand g05709(.dina(n5964), .dinb(n5959), .dout(n5965));
  jxor g05710(.dina(n5965), .dinb(a44 ), .dout(n5966));
  jnot g05711(.din(n5966), .dout(n5967));
  jand g05712(.dina(n5752), .dinb(a47 ), .dout(n5968));
  jxor g05713(.dina(a47 ), .dinb(a46 ), .dout(n5969));
  jnot g05714(.din(n5969), .dout(n5970));
  jand g05715(.dina(n5970), .dinb(n5751), .dout(n5971));
  jand g05716(.dina(n5971), .dinb(b1 ), .dout(n5972));
  jnot g05717(.din(n5751), .dout(n5973));
  jxor g05718(.dina(a46 ), .dinb(a45 ), .dout(n5974));
  jand g05719(.dina(n5974), .dinb(n5973), .dout(n5975));
  jand g05720(.dina(n5975), .dinb(b0 ), .dout(n5976));
  jand g05721(.dina(n5969), .dinb(n5751), .dout(n5977));
  jand g05722(.dina(n5977), .dinb(n338), .dout(n5978));
  jor  g05723(.dina(n5978), .dinb(n5976), .dout(n5979));
  jor  g05724(.dina(n5979), .dinb(n5972), .dout(n5980));
  jxor g05725(.dina(n5980), .dinb(n5968), .dout(n5981));
  jxor g05726(.dina(n5981), .dinb(n5967), .dout(n5982));
  jxor g05727(.dina(n5982), .dinb(n5958), .dout(n5983));
  jnot g05728(.din(n5983), .dout(n5984));
  jor  g05729(.dina(n5096), .dinb(n428), .dout(n5985));
  jor  g05730(.dina(n4904), .dinb(n357), .dout(n5986));
  jor  g05731(.dina(n5099), .dinb(n395), .dout(n5987));
  jor  g05732(.dina(n5101), .dinb(n431), .dout(n5988));
  jand g05733(.dina(n5988), .dinb(n5987), .dout(n5989));
  jand g05734(.dina(n5989), .dinb(n5986), .dout(n5990));
  jand g05735(.dina(n5990), .dinb(n5985), .dout(n5991));
  jxor g05736(.dina(n5991), .dinb(a41 ), .dout(n5992));
  jxor g05737(.dina(n5992), .dinb(n5984), .dout(n5993));
  jxor g05738(.dina(n5993), .dinb(n5954), .dout(n5994));
  jnot g05739(.din(n5994), .dout(n5995));
  jor  g05740(.dina(n4415), .dinb(n624), .dout(n5996));
  jor  g05741(.dina(n4272), .dinb(n512), .dout(n5997));
  jor  g05742(.dina(n4418), .dinb(n564), .dout(n5998));
  jor  g05743(.dina(n4420), .dinb(n627), .dout(n5999));
  jand g05744(.dina(n5999), .dinb(n5998), .dout(n6000));
  jand g05745(.dina(n6000), .dinb(n5997), .dout(n6001));
  jand g05746(.dina(n6001), .dinb(n5996), .dout(n6002));
  jxor g05747(.dina(n6002), .dinb(a38 ), .dout(n6003));
  jxor g05748(.dina(n6003), .dinb(n5995), .dout(n6004));
  jxor g05749(.dina(n6004), .dinb(n5949), .dout(n6005));
  jxor g05750(.dina(n6005), .dinb(n5944), .dout(n6006));
  jxor g05751(.dina(n6006), .dinb(n5935), .dout(n6007));
  jnot g05752(.din(n6007), .dout(n6008));
  jor  g05753(.dina(n3301), .dinb(n1019), .dout(n6009));
  jor  g05754(.dina(n3136), .dinb(n858), .dout(n6010));
  jor  g05755(.dina(n3304), .dinb(n939), .dout(n6011));
  jor  g05756(.dina(n3306), .dinb(n1022), .dout(n6012));
  jand g05757(.dina(n6012), .dinb(n6011), .dout(n6013));
  jand g05758(.dina(n6013), .dinb(n6010), .dout(n6014));
  jand g05759(.dina(n6014), .dinb(n6009), .dout(n6015));
  jxor g05760(.dina(n6015), .dinb(a32 ), .dout(n6016));
  jxor g05761(.dina(n6016), .dinb(n6008), .dout(n6017));
  jxor g05762(.dina(n6017), .dinb(n5932), .dout(n6018));
  jnot g05763(.din(n6018), .dout(n6019));
  jor  g05764(.dina(n2784), .dinb(n1397), .dout(n6020));
  jor  g05765(.dina(n2661), .dinb(n1193), .dout(n6021));
  jor  g05766(.dina(n2787), .dinb(n1290), .dout(n6022));
  jor  g05767(.dina(n2789), .dinb(n1400), .dout(n6023));
  jand g05768(.dina(n6023), .dinb(n6022), .dout(n6024));
  jand g05769(.dina(n6024), .dinb(n6021), .dout(n6025));
  jand g05770(.dina(n6025), .dinb(n6020), .dout(n6026));
  jxor g05771(.dina(n6026), .dinb(a29 ), .dout(n6027));
  jxor g05772(.dina(n6027), .dinb(n6019), .dout(n6028));
  jxor g05773(.dina(n6028), .dinb(n5929), .dout(n6029));
  jnot g05774(.din(n6029), .dout(n6030));
  jor  g05775(.dina(n2319), .dinb(n1739), .dout(n6031));
  jor  g05776(.dina(n2224), .dinb(n1420), .dout(n6032));
  jor  g05777(.dina(n2322), .dinb(n1620), .dout(n6033));
  jor  g05778(.dina(n2324), .dinb(n1742), .dout(n6034));
  jand g05779(.dina(n6034), .dinb(n6033), .dout(n6035));
  jand g05780(.dina(n6035), .dinb(n6032), .dout(n6036));
  jand g05781(.dina(n6036), .dinb(n6031), .dout(n6037));
  jxor g05782(.dina(n6037), .dinb(a26 ), .dout(n6038));
  jxor g05783(.dina(n6038), .dinb(n6030), .dout(n6039));
  jxor g05784(.dina(n6039), .dinb(n5926), .dout(n6040));
  jnot g05785(.din(n6040), .dout(n6041));
  jor  g05786(.dina(n2007), .dinb(n1939), .dout(n6042));
  jor  g05787(.dina(n1827), .dinb(n1867), .dout(n6043));
  jor  g05788(.dina(n1942), .dinb(n1887), .dout(n6044));
  jor  g05789(.dina(n1944), .dinb(n2010), .dout(n6045));
  jand g05790(.dina(n6045), .dinb(n6044), .dout(n6046));
  jand g05791(.dina(n6046), .dinb(n6043), .dout(n6047));
  jand g05792(.dina(n6047), .dinb(n6042), .dout(n6048));
  jxor g05793(.dina(n6048), .dinb(a23 ), .dout(n6049));
  jxor g05794(.dina(n6049), .dinb(n6041), .dout(n6050));
  jxor g05795(.dina(n6050), .dinb(n5921), .dout(n6051));
  jxor g05796(.dina(n6051), .dinb(n5917), .dout(n6052));
  jxor g05797(.dina(n6052), .dinb(n5908), .dout(n6053));
  jxor g05798(.dina(n6053), .dinb(n5903), .dout(n6054));
  jxor g05799(.dina(n6054), .dinb(n5894), .dout(n6055));
  jnot g05800(.din(n6055), .dout(n6056));
  jor  g05801(.dina(n3400), .dinb(n974), .dout(n6057));
  jor  g05802(.dina(n908), .dinb(n3055), .dout(n6058));
  jor  g05803(.dina(n977), .dinb(n3230), .dout(n6059));
  jor  g05804(.dina(n979), .dinb(n3403), .dout(n6060));
  jand g05805(.dina(n6060), .dinb(n6059), .dout(n6061));
  jand g05806(.dina(n6061), .dinb(n6058), .dout(n6062));
  jand g05807(.dina(n6062), .dinb(n6057), .dout(n6063));
  jxor g05808(.dina(n6063), .dinb(a14 ), .dout(n6064));
  jxor g05809(.dina(n6064), .dinb(n6056), .dout(n6065));
  jxor g05810(.dina(n6065), .dinb(n5891), .dout(n6066));
  jor  g05811(.dina(n4137), .dinb(n706), .dout(n6067));
  jor  g05812(.dina(n683), .dinb(n3588), .dout(n6068));
  jor  g05813(.dina(n709), .dinb(n3942), .dout(n6069));
  jor  g05814(.dina(n711), .dinb(n4140), .dout(n6070));
  jand g05815(.dina(n6070), .dinb(n6069), .dout(n6071));
  jand g05816(.dina(n6071), .dinb(n6068), .dout(n6072));
  jand g05817(.dina(n6072), .dinb(n6067), .dout(n6073));
  jxor g05818(.dina(n6073), .dinb(a11 ), .dout(n6074));
  jxor g05819(.dina(n6074), .dinb(n6066), .dout(n6075));
  jxor g05820(.dina(n6075), .dinb(n5887), .dout(n6076));
  jnot g05821(.din(n6076), .dout(n6077));
  jor  g05822(.dina(n4554), .dinb(n528), .dout(n6078));
  jor  g05823(.dina(n490), .dinb(n4340), .dout(n6079));
  jor  g05824(.dina(n531), .dinb(n4537), .dout(n6080));
  jor  g05825(.dina(n533), .dinb(n4557), .dout(n6081));
  jand g05826(.dina(n6081), .dinb(n6080), .dout(n6082));
  jand g05827(.dina(n6082), .dinb(n6079), .dout(n6083));
  jand g05828(.dina(n6083), .dinb(n6078), .dout(n6084));
  jxor g05829(.dina(n6084), .dinb(a8 ), .dout(n6085));
  jxor g05830(.dina(n6085), .dinb(n6077), .dout(n6086));
  jxor g05831(.dina(n6086), .dinb(n5882), .dout(n6087));
  jor  g05832(.dina(n5405), .dinb(n402), .dout(n6088));
  jor  g05833(.dina(n371), .dinb(n4974), .dout(n6089));
  jor  g05834(.dina(n405), .dinb(n4994), .dout(n6090));
  jor  g05835(.dina(n332), .dinb(n5408), .dout(n6091));
  jand g05836(.dina(n6091), .dinb(n6090), .dout(n6092));
  jand g05837(.dina(n6092), .dinb(n6089), .dout(n6093));
  jand g05838(.dina(n6093), .dinb(n6088), .dout(n6094));
  jxor g05839(.dina(n6094), .dinb(a5 ), .dout(n6095));
  jxor g05840(.dina(n6095), .dinb(n6087), .dout(n6096));
  jxor g05841(.dina(n6096), .dinb(n5877), .dout(n6097));
  jand g05842(.dina(b45 ), .dinb(b44 ), .dout(n6098));
  jand g05843(.dina(n5857), .dinb(n5856), .dout(n6099));
  jor  g05844(.dina(n6099), .dinb(n6098), .dout(n6100));
  jxor g05845(.dina(b46 ), .dinb(b45 ), .dout(n6101));
  jnot g05846(.din(n6101), .dout(n6102));
  jxor g05847(.dina(n6102), .dinb(n6100), .dout(n6103));
  jor  g05848(.dina(n6103), .dinb(n264), .dout(n6104));
  jor  g05849(.dina(n284), .dinb(n5428), .dout(n6105));
  jnot g05850(.din(b46 ), .dout(n6106));
  jor  g05851(.dina(n269), .dinb(n6106), .dout(n6107));
  jor  g05852(.dina(n271), .dinb(n5862), .dout(n6108));
  jand g05853(.dina(n6108), .dinb(n6107), .dout(n6109));
  jand g05854(.dina(n6109), .dinb(n6105), .dout(n6110));
  jand g05855(.dina(n6110), .dinb(n6104), .dout(n6111));
  jxor g05856(.dina(n6111), .dinb(n260), .dout(n6112));
  jxor g05857(.dina(n6112), .dinb(n6097), .dout(n6113));
  jxor g05858(.dina(n6113), .dinb(n5873), .dout(f46 ));
  jand g05859(.dina(n6112), .dinb(n6097), .dout(n6115));
  jand g05860(.dina(n6113), .dinb(n5873), .dout(n6116));
  jor  g05861(.dina(n6116), .dinb(n6115), .dout(n6117));
  jor  g05862(.dina(n6095), .dinb(n6087), .dout(n6118));
  jnot g05863(.din(n6118), .dout(n6119));
  jand g05864(.dina(n6096), .dinb(n5877), .dout(n6120));
  jor  g05865(.dina(n6120), .dinb(n6119), .dout(n6121));
  jor  g05866(.dina(n5425), .dinb(n402), .dout(n6122));
  jor  g05867(.dina(n371), .dinb(n4994), .dout(n6123));
  jor  g05868(.dina(n405), .dinb(n5408), .dout(n6124));
  jor  g05869(.dina(n332), .dinb(n5428), .dout(n6125));
  jand g05870(.dina(n6125), .dinb(n6124), .dout(n6126));
  jand g05871(.dina(n6126), .dinb(n6123), .dout(n6127));
  jand g05872(.dina(n6127), .dinb(n6122), .dout(n6128));
  jxor g05873(.dina(n6128), .dinb(a5 ), .dout(n6129));
  jnot g05874(.din(n6129), .dout(n6130));
  jor  g05875(.dina(n6085), .dinb(n6077), .dout(n6131));
  jnot g05876(.din(n6131), .dout(n6132));
  jand g05877(.dina(n6086), .dinb(n5881), .dout(n6133));
  jor  g05878(.dina(n6133), .dinb(n6132), .dout(n6134));
  jnot g05879(.din(n6066), .dout(n6135));
  jor  g05880(.dina(n6074), .dinb(n6135), .dout(n6136));
  jor  g05881(.dina(n6075), .dinb(n5887), .dout(n6137));
  jand g05882(.dina(n6137), .dinb(n6136), .dout(n6138));
  jor  g05883(.dina(n6064), .dinb(n6056), .dout(n6139));
  jnot g05884(.din(n6139), .dout(n6140));
  jand g05885(.dina(n6065), .dinb(n5891), .dout(n6141));
  jor  g05886(.dina(n6141), .dinb(n6140), .dout(n6142));
  jand g05887(.dina(n6053), .dinb(n5903), .dout(n6143));
  jand g05888(.dina(n6054), .dinb(n5894), .dout(n6144));
  jor  g05889(.dina(n6144), .dinb(n6143), .dout(n6145));
  jor  g05890(.dina(n3052), .dinb(n1245), .dout(n6146));
  jor  g05891(.dina(n1165), .dinb(n2870), .dout(n6147));
  jor  g05892(.dina(n1248), .dinb(n3035), .dout(n6148));
  jor  g05893(.dina(n1250), .dinb(n3055), .dout(n6149));
  jand g05894(.dina(n6149), .dinb(n6148), .dout(n6150));
  jand g05895(.dina(n6150), .dinb(n6147), .dout(n6151));
  jand g05896(.dina(n6151), .dinb(n6146), .dout(n6152));
  jxor g05897(.dina(n6152), .dinb(a17 ), .dout(n6153));
  jnot g05898(.din(n6153), .dout(n6154));
  jand g05899(.dina(n6051), .dinb(n5917), .dout(n6155));
  jand g05900(.dina(n6052), .dinb(n5908), .dout(n6156));
  jor  g05901(.dina(n6156), .dinb(n6155), .dout(n6157));
  jor  g05902(.dina(n2576), .dinb(n1566), .dout(n6158));
  jor  g05903(.dina(n1489), .dinb(n2407), .dout(n6159));
  jor  g05904(.dina(n1569), .dinb(n2559), .dout(n6160));
  jor  g05905(.dina(n1571), .dinb(n2579), .dout(n6161));
  jand g05906(.dina(n6161), .dinb(n6160), .dout(n6162));
  jand g05907(.dina(n6162), .dinb(n6159), .dout(n6163));
  jand g05908(.dina(n6163), .dinb(n6158), .dout(n6164));
  jxor g05909(.dina(n6164), .dinb(a20 ), .dout(n6165));
  jnot g05910(.din(n6165), .dout(n6166));
  jor  g05911(.dina(n6049), .dinb(n6041), .dout(n6167));
  jnot g05912(.din(n6167), .dout(n6168));
  jand g05913(.dina(n6050), .dinb(n5921), .dout(n6169));
  jor  g05914(.dina(n6169), .dinb(n6168), .dout(n6170));
  jor  g05915(.dina(n2145), .dinb(n1939), .dout(n6171));
  jor  g05916(.dina(n1827), .dinb(n1887), .dout(n6172));
  jor  g05917(.dina(n1942), .dinb(n2010), .dout(n6173));
  jor  g05918(.dina(n1944), .dinb(n2148), .dout(n6174));
  jand g05919(.dina(n6174), .dinb(n6173), .dout(n6175));
  jand g05920(.dina(n6175), .dinb(n6172), .dout(n6176));
  jand g05921(.dina(n6176), .dinb(n6171), .dout(n6177));
  jxor g05922(.dina(n6177), .dinb(a23 ), .dout(n6178));
  jnot g05923(.din(n6178), .dout(n6179));
  jor  g05924(.dina(n6038), .dinb(n6030), .dout(n6180));
  jand g05925(.dina(n6039), .dinb(n5926), .dout(n6181));
  jnot g05926(.din(n6181), .dout(n6182));
  jand g05927(.dina(n6182), .dinb(n6180), .dout(n6183));
  jnot g05928(.din(n6183), .dout(n6184));
  jor  g05929(.dina(n6027), .dinb(n6019), .dout(n6185));
  jand g05930(.dina(n6028), .dinb(n5929), .dout(n6186));
  jnot g05931(.din(n6186), .dout(n6187));
  jand g05932(.dina(n6187), .dinb(n6185), .dout(n6188));
  jnot g05933(.din(n6188), .dout(n6189));
  jor  g05934(.dina(n2784), .dinb(n1417), .dout(n6190));
  jor  g05935(.dina(n2661), .dinb(n1290), .dout(n6191));
  jor  g05936(.dina(n2787), .dinb(n1400), .dout(n6192));
  jor  g05937(.dina(n2789), .dinb(n1420), .dout(n6193));
  jand g05938(.dina(n6193), .dinb(n6192), .dout(n6194));
  jand g05939(.dina(n6194), .dinb(n6191), .dout(n6195));
  jand g05940(.dina(n6195), .dinb(n6190), .dout(n6196));
  jxor g05941(.dina(n6196), .dinb(a29 ), .dout(n6197));
  jnot g05942(.din(n6197), .dout(n6198));
  jor  g05943(.dina(n6016), .dinb(n6008), .dout(n6199));
  jand g05944(.dina(n6017), .dinb(n5932), .dout(n6200));
  jnot g05945(.din(n6200), .dout(n6201));
  jand g05946(.dina(n6201), .dinb(n6199), .dout(n6202));
  jnot g05947(.din(n6202), .dout(n6203));
  jor  g05948(.dina(n3301), .dinb(n1190), .dout(n6204));
  jor  g05949(.dina(n3136), .dinb(n939), .dout(n6205));
  jor  g05950(.dina(n3304), .dinb(n1022), .dout(n6206));
  jor  g05951(.dina(n3306), .dinb(n1193), .dout(n6207));
  jand g05952(.dina(n6207), .dinb(n6206), .dout(n6208));
  jand g05953(.dina(n6208), .dinb(n6205), .dout(n6209));
  jand g05954(.dina(n6209), .dinb(n6204), .dout(n6210));
  jxor g05955(.dina(n6210), .dinb(a32 ), .dout(n6211));
  jnot g05956(.din(n6211), .dout(n6212));
  jand g05957(.dina(n6005), .dinb(n5944), .dout(n6213));
  jand g05958(.dina(n6006), .dinb(n5935), .dout(n6214));
  jor  g05959(.dina(n6214), .dinb(n6213), .dout(n6215));
  jor  g05960(.dina(n6003), .dinb(n5995), .dout(n6216));
  jand g05961(.dina(n6004), .dinb(n5949), .dout(n6217));
  jnot g05962(.din(n6217), .dout(n6218));
  jand g05963(.dina(n6218), .dinb(n6216), .dout(n6219));
  jnot g05964(.din(n6219), .dout(n6220));
  jor  g05965(.dina(n4415), .dinb(n644), .dout(n6221));
  jor  g05966(.dina(n4272), .dinb(n564), .dout(n6222));
  jor  g05967(.dina(n4418), .dinb(n627), .dout(n6223));
  jor  g05968(.dina(n4420), .dinb(n647), .dout(n6224));
  jand g05969(.dina(n6224), .dinb(n6223), .dout(n6225));
  jand g05970(.dina(n6225), .dinb(n6222), .dout(n6226));
  jand g05971(.dina(n6226), .dinb(n6221), .dout(n6227));
  jxor g05972(.dina(n6227), .dinb(a38 ), .dout(n6228));
  jnot g05973(.din(n6228), .dout(n6229));
  jor  g05974(.dina(n5992), .dinb(n5984), .dout(n6230));
  jand g05975(.dina(n5993), .dinb(n5954), .dout(n6231));
  jnot g05976(.din(n6231), .dout(n6232));
  jand g05977(.dina(n6232), .dinb(n6230), .dout(n6233));
  jnot g05978(.din(n6233), .dout(n6234));
  jor  g05979(.dina(n5096), .dinb(n509), .dout(n6235));
  jor  g05980(.dina(n4904), .dinb(n395), .dout(n6236));
  jor  g05981(.dina(n5099), .dinb(n431), .dout(n6237));
  jor  g05982(.dina(n5101), .dinb(n512), .dout(n6238));
  jand g05983(.dina(n6238), .dinb(n6237), .dout(n6239));
  jand g05984(.dina(n6239), .dinb(n6236), .dout(n6240));
  jand g05985(.dina(n6240), .dinb(n6235), .dout(n6241));
  jxor g05986(.dina(n6241), .dinb(a41 ), .dout(n6242));
  jnot g05987(.din(n6242), .dout(n6243));
  jand g05988(.dina(n5981), .dinb(n5967), .dout(n6244));
  jand g05989(.dina(n5982), .dinb(n5958), .dout(n6245));
  jor  g05990(.dina(n6245), .dinb(n6244), .dout(n6246));
  jor  g05991(.dina(n5739), .dinb(n354), .dout(n6247));
  jor  g05992(.dina(n5574), .dinb(n299), .dout(n6248));
  jor  g05993(.dina(n5742), .dinb(n322), .dout(n6249));
  jor  g05994(.dina(n5744), .dinb(n357), .dout(n6250));
  jand g05995(.dina(n6250), .dinb(n6249), .dout(n6251));
  jand g05996(.dina(n6251), .dinb(n6248), .dout(n6252));
  jand g05997(.dina(n6252), .dinb(n6247), .dout(n6253));
  jxor g05998(.dina(n6253), .dinb(a44 ), .dout(n6254));
  jnot g05999(.din(n6254), .dout(n6255));
  jnot g06000(.din(n5980), .dout(n6256));
  jand g06001(.dina(n5753), .dinb(a47 ), .dout(n6257));
  jand g06002(.dina(n6257), .dinb(n6256), .dout(n6258));
  jnot g06003(.din(n6258), .dout(n6259));
  jand g06004(.dina(n6259), .dinb(a47 ), .dout(n6260));
  jor  g06005(.dina(n5974), .dinb(n5970), .dout(n6261));
  jor  g06006(.dina(n6261), .dinb(n5751), .dout(n6262));
  jnot g06007(.din(n6262), .dout(n6263));
  jand g06008(.dina(n6263), .dinb(b0 ), .dout(n6264));
  jand g06009(.dina(n5971), .dinb(b2 ), .dout(n6265));
  jand g06010(.dina(n5975), .dinb(b1 ), .dout(n6266));
  jand g06011(.dina(n5977), .dinb(n375), .dout(n6267));
  jor  g06012(.dina(n6267), .dinb(n6266), .dout(n6268));
  jor  g06013(.dina(n6268), .dinb(n6265), .dout(n6269));
  jor  g06014(.dina(n6269), .dinb(n6264), .dout(n6270));
  jxor g06015(.dina(n6270), .dinb(n6260), .dout(n6271));
  jxor g06016(.dina(n6271), .dinb(n6255), .dout(n6272));
  jxor g06017(.dina(n6272), .dinb(n6246), .dout(n6273));
  jxor g06018(.dina(n6273), .dinb(n6243), .dout(n6274));
  jxor g06019(.dina(n6274), .dinb(n6234), .dout(n6275));
  jxor g06020(.dina(n6275), .dinb(n6229), .dout(n6276));
  jxor g06021(.dina(n6276), .dinb(n6220), .dout(n6277));
  jnot g06022(.din(n6277), .dout(n6278));
  jor  g06023(.dina(n3849), .dinb(n855), .dout(n6279));
  jor  g06024(.dina(n3689), .dinb(n758), .dout(n6280));
  jor  g06025(.dina(n3852), .dinb(n778), .dout(n6281));
  jor  g06026(.dina(n3854), .dinb(n858), .dout(n6282));
  jand g06027(.dina(n6282), .dinb(n6281), .dout(n6283));
  jand g06028(.dina(n6283), .dinb(n6280), .dout(n6284));
  jand g06029(.dina(n6284), .dinb(n6279), .dout(n6285));
  jxor g06030(.dina(n6285), .dinb(a35 ), .dout(n6286));
  jxor g06031(.dina(n6286), .dinb(n6278), .dout(n6287));
  jxor g06032(.dina(n6287), .dinb(n6215), .dout(n6288));
  jxor g06033(.dina(n6288), .dinb(n6212), .dout(n6289));
  jxor g06034(.dina(n6289), .dinb(n6203), .dout(n6290));
  jxor g06035(.dina(n6290), .dinb(n6198), .dout(n6291));
  jxor g06036(.dina(n6291), .dinb(n6189), .dout(n6292));
  jnot g06037(.din(n6292), .dout(n6293));
  jor  g06038(.dina(n2319), .dinb(n1864), .dout(n6294));
  jor  g06039(.dina(n2224), .dinb(n1620), .dout(n6295));
  jor  g06040(.dina(n2322), .dinb(n1742), .dout(n6296));
  jor  g06041(.dina(n2324), .dinb(n1867), .dout(n6297));
  jand g06042(.dina(n6297), .dinb(n6296), .dout(n6298));
  jand g06043(.dina(n6298), .dinb(n6295), .dout(n6299));
  jand g06044(.dina(n6299), .dinb(n6294), .dout(n6300));
  jxor g06045(.dina(n6300), .dinb(a26 ), .dout(n6301));
  jxor g06046(.dina(n6301), .dinb(n6293), .dout(n6302));
  jxor g06047(.dina(n6302), .dinb(n6184), .dout(n6303));
  jxor g06048(.dina(n6303), .dinb(n6179), .dout(n6304));
  jxor g06049(.dina(n6304), .dinb(n6170), .dout(n6305));
  jxor g06050(.dina(n6305), .dinb(n6166), .dout(n6306));
  jxor g06051(.dina(n6306), .dinb(n6157), .dout(n6307));
  jxor g06052(.dina(n6307), .dinb(n6154), .dout(n6308));
  jxor g06053(.dina(n6308), .dinb(n6145), .dout(n6309));
  jnot g06054(.din(n6309), .dout(n6310));
  jor  g06055(.dina(n3585), .dinb(n974), .dout(n6311));
  jor  g06056(.dina(n908), .dinb(n3230), .dout(n6312));
  jor  g06057(.dina(n977), .dinb(n3403), .dout(n6313));
  jor  g06058(.dina(n979), .dinb(n3588), .dout(n6314));
  jand g06059(.dina(n6314), .dinb(n6313), .dout(n6315));
  jand g06060(.dina(n6315), .dinb(n6312), .dout(n6316));
  jand g06061(.dina(n6316), .dinb(n6311), .dout(n6317));
  jxor g06062(.dina(n6317), .dinb(a14 ), .dout(n6318));
  jxor g06063(.dina(n6318), .dinb(n6310), .dout(n6319));
  jxor g06064(.dina(n6319), .dinb(n6142), .dout(n6320));
  jor  g06065(.dina(n4337), .dinb(n706), .dout(n6321));
  jor  g06066(.dina(n683), .dinb(n3942), .dout(n6322));
  jor  g06067(.dina(n709), .dinb(n4140), .dout(n6323));
  jor  g06068(.dina(n711), .dinb(n4340), .dout(n6324));
  jand g06069(.dina(n6324), .dinb(n6323), .dout(n6325));
  jand g06070(.dina(n6325), .dinb(n6322), .dout(n6326));
  jand g06071(.dina(n6326), .dinb(n6321), .dout(n6327));
  jxor g06072(.dina(n6327), .dinb(a11 ), .dout(n6328));
  jxor g06073(.dina(n6328), .dinb(n6320), .dout(n6329));
  jxor g06074(.dina(n6329), .dinb(n6138), .dout(n6330));
  jnot g06075(.din(n6330), .dout(n6331));
  jor  g06076(.dina(n4971), .dinb(n528), .dout(n6332));
  jor  g06077(.dina(n490), .dinb(n4537), .dout(n6333));
  jor  g06078(.dina(n531), .dinb(n4557), .dout(n6334));
  jor  g06079(.dina(n533), .dinb(n4974), .dout(n6335));
  jand g06080(.dina(n6335), .dinb(n6334), .dout(n6336));
  jand g06081(.dina(n6336), .dinb(n6333), .dout(n6337));
  jand g06082(.dina(n6337), .dinb(n6332), .dout(n6338));
  jxor g06083(.dina(n6338), .dinb(a8 ), .dout(n6339));
  jxor g06084(.dina(n6339), .dinb(n6331), .dout(n6340));
  jxor g06085(.dina(n6340), .dinb(n6134), .dout(n6341));
  jxor g06086(.dina(n6341), .dinb(n6130), .dout(n6342));
  jxor g06087(.dina(n6342), .dinb(n6121), .dout(n6343));
  jand g06088(.dina(b46 ), .dinb(b45 ), .dout(n6344));
  jand g06089(.dina(n6101), .dinb(n6100), .dout(n6345));
  jor  g06090(.dina(n6345), .dinb(n6344), .dout(n6346));
  jxor g06091(.dina(b47 ), .dinb(b46 ), .dout(n6347));
  jnot g06092(.din(n6347), .dout(n6348));
  jxor g06093(.dina(n6348), .dinb(n6346), .dout(n6349));
  jor  g06094(.dina(n6349), .dinb(n264), .dout(n6350));
  jor  g06095(.dina(n284), .dinb(n5862), .dout(n6351));
  jnot g06096(.din(b47 ), .dout(n6352));
  jor  g06097(.dina(n269), .dinb(n6352), .dout(n6353));
  jor  g06098(.dina(n271), .dinb(n6106), .dout(n6354));
  jand g06099(.dina(n6354), .dinb(n6353), .dout(n6355));
  jand g06100(.dina(n6355), .dinb(n6351), .dout(n6356));
  jand g06101(.dina(n6356), .dinb(n6350), .dout(n6357));
  jxor g06102(.dina(n6357), .dinb(n260), .dout(n6358));
  jxor g06103(.dina(n6358), .dinb(n6343), .dout(n6359));
  jxor g06104(.dina(n6359), .dinb(n6117), .dout(f47 ));
  jand g06105(.dina(n6358), .dinb(n6343), .dout(n6361));
  jand g06106(.dina(n6359), .dinb(n6117), .dout(n6362));
  jor  g06107(.dina(n6362), .dinb(n6361), .dout(n6363));
  jand g06108(.dina(b47 ), .dinb(b46 ), .dout(n6364));
  jand g06109(.dina(n6347), .dinb(n6346), .dout(n6365));
  jor  g06110(.dina(n6365), .dinb(n6364), .dout(n6366));
  jxor g06111(.dina(b48 ), .dinb(b47 ), .dout(n6367));
  jnot g06112(.din(n6367), .dout(n6368));
  jxor g06113(.dina(n6368), .dinb(n6366), .dout(n6369));
  jor  g06114(.dina(n6369), .dinb(n264), .dout(n6370));
  jor  g06115(.dina(n284), .dinb(n6106), .dout(n6371));
  jnot g06116(.din(b48 ), .dout(n6372));
  jor  g06117(.dina(n269), .dinb(n6372), .dout(n6373));
  jor  g06118(.dina(n271), .dinb(n6352), .dout(n6374));
  jand g06119(.dina(n6374), .dinb(n6373), .dout(n6375));
  jand g06120(.dina(n6375), .dinb(n6371), .dout(n6376));
  jand g06121(.dina(n6376), .dinb(n6370), .dout(n6377));
  jxor g06122(.dina(n6377), .dinb(n260), .dout(n6378));
  jand g06123(.dina(n6341), .dinb(n6130), .dout(n6379));
  jand g06124(.dina(n6342), .dinb(n6121), .dout(n6380));
  jor  g06125(.dina(n6380), .dinb(n6379), .dout(n6381));
  jor  g06126(.dina(n5859), .dinb(n402), .dout(n6382));
  jor  g06127(.dina(n371), .dinb(n5408), .dout(n6383));
  jor  g06128(.dina(n405), .dinb(n5428), .dout(n6384));
  jor  g06129(.dina(n332), .dinb(n5862), .dout(n6385));
  jand g06130(.dina(n6385), .dinb(n6384), .dout(n6386));
  jand g06131(.dina(n6386), .dinb(n6383), .dout(n6387));
  jand g06132(.dina(n6387), .dinb(n6382), .dout(n6388));
  jxor g06133(.dina(n6388), .dinb(a5 ), .dout(n6389));
  jnot g06134(.din(n6389), .dout(n6390));
  jor  g06135(.dina(n6339), .dinb(n6331), .dout(n6391));
  jnot g06136(.din(n6391), .dout(n6392));
  jand g06137(.dina(n6340), .dinb(n6134), .dout(n6393));
  jor  g06138(.dina(n6393), .dinb(n6392), .dout(n6394));
  jnot g06139(.din(n6320), .dout(n6395));
  jor  g06140(.dina(n6328), .dinb(n6395), .dout(n6396));
  jor  g06141(.dina(n6329), .dinb(n6138), .dout(n6397));
  jand g06142(.dina(n6397), .dinb(n6396), .dout(n6398));
  jor  g06143(.dina(n6318), .dinb(n6310), .dout(n6399));
  jnot g06144(.din(n6399), .dout(n6400));
  jand g06145(.dina(n6319), .dinb(n6142), .dout(n6401));
  jor  g06146(.dina(n6401), .dinb(n6400), .dout(n6402));
  jor  g06147(.dina(n3939), .dinb(n974), .dout(n6403));
  jor  g06148(.dina(n908), .dinb(n3403), .dout(n6404));
  jor  g06149(.dina(n977), .dinb(n3588), .dout(n6405));
  jor  g06150(.dina(n979), .dinb(n3942), .dout(n6406));
  jand g06151(.dina(n6406), .dinb(n6405), .dout(n6407));
  jand g06152(.dina(n6407), .dinb(n6404), .dout(n6408));
  jand g06153(.dina(n6408), .dinb(n6403), .dout(n6409));
  jxor g06154(.dina(n6409), .dinb(a14 ), .dout(n6410));
  jnot g06155(.din(n6410), .dout(n6411));
  jand g06156(.dina(n6307), .dinb(n6154), .dout(n6412));
  jand g06157(.dina(n6308), .dinb(n6145), .dout(n6413));
  jor  g06158(.dina(n6413), .dinb(n6412), .dout(n6414));
  jand g06159(.dina(n6305), .dinb(n6166), .dout(n6415));
  jnot g06160(.din(n6415), .dout(n6416));
  jnot g06161(.din(n6155), .dout(n6417));
  jnot g06162(.din(n5685), .dout(n6418));
  jnot g06163(.din(n5048), .dout(n6419));
  jor  g06164(.dina(n5161), .dinb(n6419), .dout(n6420));
  jand g06165(.dina(n6420), .dinb(n5239), .dout(n6421));
  jor  g06166(.dina(n5370), .dinb(n6421), .dout(n6422));
  jand g06167(.dina(n6422), .dinb(n5480), .dout(n6423));
  jnot g06168(.din(n5616), .dout(n6424));
  jor  g06169(.dina(n6424), .dinb(n6423), .dout(n6425));
  jand g06170(.dina(n6425), .dinb(n6418), .dout(n6426));
  jor  g06171(.dina(n5815), .dinb(n6426), .dout(n6427));
  jand g06172(.dina(n6427), .dinb(n5905), .dout(n6428));
  jnot g06173(.din(n6052), .dout(n6429));
  jor  g06174(.dina(n6429), .dinb(n6428), .dout(n6430));
  jand g06175(.dina(n6430), .dinb(n6417), .dout(n6431));
  jnot g06176(.din(n6306), .dout(n6432));
  jor  g06177(.dina(n6432), .dinb(n6431), .dout(n6433));
  jand g06178(.dina(n6433), .dinb(n6416), .dout(n6434));
  jor  g06179(.dina(n2867), .dinb(n1566), .dout(n6435));
  jor  g06180(.dina(n1489), .dinb(n2559), .dout(n6436));
  jor  g06181(.dina(n1569), .dinb(n2579), .dout(n6437));
  jor  g06182(.dina(n1571), .dinb(n2870), .dout(n6438));
  jand g06183(.dina(n6438), .dinb(n6437), .dout(n6439));
  jand g06184(.dina(n6439), .dinb(n6436), .dout(n6440));
  jand g06185(.dina(n6440), .dinb(n6435), .dout(n6441));
  jxor g06186(.dina(n6441), .dinb(a20 ), .dout(n6442));
  jnot g06187(.din(n6442), .dout(n6443));
  jand g06188(.dina(n6303), .dinb(n6179), .dout(n6444));
  jand g06189(.dina(n6304), .dinb(n6170), .dout(n6445));
  jor  g06190(.dina(n6445), .dinb(n6444), .dout(n6446));
  jor  g06191(.dina(n6301), .dinb(n6293), .dout(n6447));
  jand g06192(.dina(n6302), .dinb(n6184), .dout(n6448));
  jnot g06193(.din(n6448), .dout(n6449));
  jand g06194(.dina(n6449), .dinb(n6447), .dout(n6450));
  jnot g06195(.din(n6450), .dout(n6451));
  jand g06196(.dina(n6290), .dinb(n6198), .dout(n6452));
  jand g06197(.dina(n6291), .dinb(n6189), .dout(n6453));
  jor  g06198(.dina(n6453), .dinb(n6452), .dout(n6454));
  jand g06199(.dina(n6288), .dinb(n6212), .dout(n6455));
  jand g06200(.dina(n6289), .dinb(n6203), .dout(n6456));
  jor  g06201(.dina(n6456), .dinb(n6455), .dout(n6457));
  jor  g06202(.dina(n6286), .dinb(n6278), .dout(n6458));
  jand g06203(.dina(n6287), .dinb(n6215), .dout(n6459));
  jnot g06204(.din(n6459), .dout(n6460));
  jand g06205(.dina(n6460), .dinb(n6458), .dout(n6461));
  jnot g06206(.din(n6461), .dout(n6462));
  jor  g06207(.dina(n3849), .dinb(n936), .dout(n6463));
  jor  g06208(.dina(n3689), .dinb(n778), .dout(n6464));
  jor  g06209(.dina(n3852), .dinb(n858), .dout(n6465));
  jor  g06210(.dina(n3854), .dinb(n939), .dout(n6466));
  jand g06211(.dina(n6466), .dinb(n6465), .dout(n6467));
  jand g06212(.dina(n6467), .dinb(n6464), .dout(n6468));
  jand g06213(.dina(n6468), .dinb(n6463), .dout(n6469));
  jxor g06214(.dina(n6469), .dinb(a35 ), .dout(n6470));
  jnot g06215(.din(n6470), .dout(n6471));
  jand g06216(.dina(n6275), .dinb(n6229), .dout(n6472));
  jand g06217(.dina(n6276), .dinb(n6220), .dout(n6473));
  jor  g06218(.dina(n6473), .dinb(n6472), .dout(n6474));
  jor  g06219(.dina(n4415), .dinb(n755), .dout(n6475));
  jor  g06220(.dina(n4272), .dinb(n627), .dout(n6476));
  jor  g06221(.dina(n4418), .dinb(n647), .dout(n6477));
  jor  g06222(.dina(n4420), .dinb(n758), .dout(n6478));
  jand g06223(.dina(n6478), .dinb(n6477), .dout(n6479));
  jand g06224(.dina(n6479), .dinb(n6476), .dout(n6480));
  jand g06225(.dina(n6480), .dinb(n6475), .dout(n6481));
  jxor g06226(.dina(n6481), .dinb(a38 ), .dout(n6482));
  jnot g06227(.din(n6482), .dout(n6483));
  jand g06228(.dina(n6273), .dinb(n6243), .dout(n6484));
  jand g06229(.dina(n6274), .dinb(n6234), .dout(n6485));
  jor  g06230(.dina(n6485), .dinb(n6484), .dout(n6486));
  jand g06231(.dina(n6271), .dinb(n6255), .dout(n6487));
  jand g06232(.dina(n6272), .dinb(n6246), .dout(n6488));
  jor  g06233(.dina(n6488), .dinb(n6487), .dout(n6489));
  jnot g06234(.din(n5977), .dout(n6490));
  jor  g06235(.dina(n6490), .dinb(n296), .dout(n6491));
  jor  g06236(.dina(n6262), .dinb(n267), .dout(n6492));
  jnot g06237(.din(n5975), .dout(n6493));
  jor  g06238(.dina(n6493), .dinb(n279), .dout(n6494));
  jnot g06239(.din(n5971), .dout(n6495));
  jor  g06240(.dina(n6495), .dinb(n299), .dout(n6496));
  jand g06241(.dina(n6496), .dinb(n6494), .dout(n6497));
  jand g06242(.dina(n6497), .dinb(n6492), .dout(n6498));
  jand g06243(.dina(n6498), .dinb(n6491), .dout(n6499));
  jxor g06244(.dina(n6499), .dinb(a47 ), .dout(n6500));
  jnot g06245(.din(n6500), .dout(n6501));
  jxor g06246(.dina(a48 ), .dinb(a47 ), .dout(n6502));
  jand g06247(.dina(n6502), .dinb(b0 ), .dout(n6503));
  jnot g06248(.din(n6503), .dout(n6504));
  jor  g06249(.dina(n6270), .dinb(n6259), .dout(n6505));
  jxor g06250(.dina(n6505), .dinb(n6504), .dout(n6506));
  jxor g06251(.dina(n6506), .dinb(n6501), .dout(n6507));
  jnot g06252(.din(n6507), .dout(n6508));
  jor  g06253(.dina(n5739), .dinb(n392), .dout(n6509));
  jor  g06254(.dina(n5574), .dinb(n322), .dout(n6510));
  jor  g06255(.dina(n5742), .dinb(n357), .dout(n6511));
  jor  g06256(.dina(n5744), .dinb(n395), .dout(n6512));
  jand g06257(.dina(n6512), .dinb(n6511), .dout(n6513));
  jand g06258(.dina(n6513), .dinb(n6510), .dout(n6514));
  jand g06259(.dina(n6514), .dinb(n6509), .dout(n6515));
  jxor g06260(.dina(n6515), .dinb(a44 ), .dout(n6516));
  jxor g06261(.dina(n6516), .dinb(n6508), .dout(n6517));
  jxor g06262(.dina(n6517), .dinb(n6489), .dout(n6518));
  jnot g06263(.din(n6518), .dout(n6519));
  jor  g06264(.dina(n5096), .dinb(n561), .dout(n6520));
  jor  g06265(.dina(n4904), .dinb(n431), .dout(n6521));
  jor  g06266(.dina(n5099), .dinb(n512), .dout(n6522));
  jor  g06267(.dina(n5101), .dinb(n564), .dout(n6523));
  jand g06268(.dina(n6523), .dinb(n6522), .dout(n6524));
  jand g06269(.dina(n6524), .dinb(n6521), .dout(n6525));
  jand g06270(.dina(n6525), .dinb(n6520), .dout(n6526));
  jxor g06271(.dina(n6526), .dinb(a41 ), .dout(n6527));
  jxor g06272(.dina(n6527), .dinb(n6519), .dout(n6528));
  jxor g06273(.dina(n6528), .dinb(n6486), .dout(n6529));
  jxor g06274(.dina(n6529), .dinb(n6483), .dout(n6530));
  jxor g06275(.dina(n6530), .dinb(n6474), .dout(n6531));
  jxor g06276(.dina(n6531), .dinb(n6471), .dout(n6532));
  jxor g06277(.dina(n6532), .dinb(n6462), .dout(n6533));
  jnot g06278(.din(n6533), .dout(n6534));
  jor  g06279(.dina(n3301), .dinb(n1287), .dout(n6535));
  jor  g06280(.dina(n3136), .dinb(n1022), .dout(n6536));
  jor  g06281(.dina(n3304), .dinb(n1193), .dout(n6537));
  jor  g06282(.dina(n3306), .dinb(n1290), .dout(n6538));
  jand g06283(.dina(n6538), .dinb(n6537), .dout(n6539));
  jand g06284(.dina(n6539), .dinb(n6536), .dout(n6540));
  jand g06285(.dina(n6540), .dinb(n6535), .dout(n6541));
  jxor g06286(.dina(n6541), .dinb(a32 ), .dout(n6542));
  jxor g06287(.dina(n6542), .dinb(n6534), .dout(n6543));
  jxor g06288(.dina(n6543), .dinb(n6457), .dout(n6544));
  jnot g06289(.din(n6544), .dout(n6545));
  jor  g06290(.dina(n2784), .dinb(n1617), .dout(n6546));
  jor  g06291(.dina(n2661), .dinb(n1400), .dout(n6547));
  jor  g06292(.dina(n2787), .dinb(n1420), .dout(n6548));
  jor  g06293(.dina(n2789), .dinb(n1620), .dout(n6549));
  jand g06294(.dina(n6549), .dinb(n6548), .dout(n6550));
  jand g06295(.dina(n6550), .dinb(n6547), .dout(n6551));
  jand g06296(.dina(n6551), .dinb(n6546), .dout(n6552));
  jxor g06297(.dina(n6552), .dinb(a29 ), .dout(n6553));
  jxor g06298(.dina(n6553), .dinb(n6545), .dout(n6554));
  jxor g06299(.dina(n6554), .dinb(n6454), .dout(n6555));
  jnot g06300(.din(n6555), .dout(n6556));
  jor  g06301(.dina(n2319), .dinb(n1884), .dout(n6557));
  jor  g06302(.dina(n2224), .dinb(n1742), .dout(n6558));
  jor  g06303(.dina(n2322), .dinb(n1867), .dout(n6559));
  jor  g06304(.dina(n2324), .dinb(n1887), .dout(n6560));
  jand g06305(.dina(n6560), .dinb(n6559), .dout(n6561));
  jand g06306(.dina(n6561), .dinb(n6558), .dout(n6562));
  jand g06307(.dina(n6562), .dinb(n6557), .dout(n6563));
  jxor g06308(.dina(n6563), .dinb(a26 ), .dout(n6564));
  jxor g06309(.dina(n6564), .dinb(n6556), .dout(n6565));
  jxor g06310(.dina(n6565), .dinb(n6451), .dout(n6566));
  jnot g06311(.din(n6566), .dout(n6567));
  jor  g06312(.dina(n2404), .dinb(n1939), .dout(n6568));
  jor  g06313(.dina(n1827), .dinb(n2010), .dout(n6569));
  jor  g06314(.dina(n1942), .dinb(n2148), .dout(n6570));
  jor  g06315(.dina(n1944), .dinb(n2407), .dout(n6571));
  jand g06316(.dina(n6571), .dinb(n6570), .dout(n6572));
  jand g06317(.dina(n6572), .dinb(n6569), .dout(n6573));
  jand g06318(.dina(n6573), .dinb(n6568), .dout(n6574));
  jxor g06319(.dina(n6574), .dinb(a23 ), .dout(n6575));
  jxor g06320(.dina(n6575), .dinb(n6567), .dout(n6576));
  jxor g06321(.dina(n6576), .dinb(n6446), .dout(n6577));
  jxor g06322(.dina(n6577), .dinb(n6443), .dout(n6578));
  jxor g06323(.dina(n6578), .dinb(n6434), .dout(n6579));
  jor  g06324(.dina(n3227), .dinb(n1245), .dout(n6580));
  jor  g06325(.dina(n1165), .dinb(n3035), .dout(n6581));
  jor  g06326(.dina(n1248), .dinb(n3055), .dout(n6582));
  jor  g06327(.dina(n1250), .dinb(n3230), .dout(n6583));
  jand g06328(.dina(n6583), .dinb(n6582), .dout(n6584));
  jand g06329(.dina(n6584), .dinb(n6581), .dout(n6585));
  jand g06330(.dina(n6585), .dinb(n6580), .dout(n6586));
  jxor g06331(.dina(n6586), .dinb(a17 ), .dout(n6587));
  jxor g06332(.dina(n6587), .dinb(n6579), .dout(n6588));
  jxor g06333(.dina(n6588), .dinb(n6414), .dout(n6589));
  jxor g06334(.dina(n6589), .dinb(n6411), .dout(n6590));
  jxor g06335(.dina(n6590), .dinb(n6402), .dout(n6591));
  jor  g06336(.dina(n4534), .dinb(n706), .dout(n6592));
  jor  g06337(.dina(n683), .dinb(n4140), .dout(n6593));
  jor  g06338(.dina(n709), .dinb(n4340), .dout(n6594));
  jor  g06339(.dina(n711), .dinb(n4537), .dout(n6595));
  jand g06340(.dina(n6595), .dinb(n6594), .dout(n6596));
  jand g06341(.dina(n6596), .dinb(n6593), .dout(n6597));
  jand g06342(.dina(n6597), .dinb(n6592), .dout(n6598));
  jxor g06343(.dina(n6598), .dinb(a11 ), .dout(n6599));
  jxor g06344(.dina(n6599), .dinb(n6591), .dout(n6600));
  jxor g06345(.dina(n6600), .dinb(n6398), .dout(n6601));
  jnot g06346(.din(n6601), .dout(n6602));
  jor  g06347(.dina(n4991), .dinb(n528), .dout(n6603));
  jor  g06348(.dina(n490), .dinb(n4557), .dout(n6604));
  jor  g06349(.dina(n531), .dinb(n4974), .dout(n6605));
  jor  g06350(.dina(n533), .dinb(n4994), .dout(n6606));
  jand g06351(.dina(n6606), .dinb(n6605), .dout(n6607));
  jand g06352(.dina(n6607), .dinb(n6604), .dout(n6608));
  jand g06353(.dina(n6608), .dinb(n6603), .dout(n6609));
  jxor g06354(.dina(n6609), .dinb(a8 ), .dout(n6610));
  jxor g06355(.dina(n6610), .dinb(n6602), .dout(n6611));
  jxor g06356(.dina(n6611), .dinb(n6394), .dout(n6612));
  jxor g06357(.dina(n6612), .dinb(n6390), .dout(n6613));
  jxor g06358(.dina(n6613), .dinb(n6381), .dout(n6614));
  jxor g06359(.dina(n6614), .dinb(n6378), .dout(n6615));
  jxor g06360(.dina(n6615), .dinb(n6363), .dout(f48 ));
  jand g06361(.dina(n6614), .dinb(n6378), .dout(n6617));
  jand g06362(.dina(n6615), .dinb(n6363), .dout(n6618));
  jor  g06363(.dina(n6618), .dinb(n6617), .dout(n6619));
  jand g06364(.dina(n6612), .dinb(n6390), .dout(n6620));
  jand g06365(.dina(n6613), .dinb(n6381), .dout(n6621));
  jor  g06366(.dina(n6621), .dinb(n6620), .dout(n6622));
  jor  g06367(.dina(n6610), .dinb(n6602), .dout(n6623));
  jnot g06368(.din(n6623), .dout(n6624));
  jand g06369(.dina(n6611), .dinb(n6394), .dout(n6625));
  jor  g06370(.dina(n6625), .dinb(n6624), .dout(n6626));
  jnot g06371(.din(n6626), .dout(n6627));
  jnot g06372(.din(n6591), .dout(n6628));
  jor  g06373(.dina(n6599), .dinb(n6628), .dout(n6629));
  jor  g06374(.dina(n6600), .dinb(n6398), .dout(n6630));
  jand g06375(.dina(n6630), .dinb(n6629), .dout(n6631));
  jand g06376(.dina(n6589), .dinb(n6411), .dout(n6632));
  jand g06377(.dina(n6590), .dinb(n6402), .dout(n6633));
  jor  g06378(.dina(n6633), .dinb(n6632), .dout(n6634));
  jor  g06379(.dina(n6587), .dinb(n6579), .dout(n6635));
  jnot g06380(.din(n6635), .dout(n6636));
  jand g06381(.dina(n6588), .dinb(n6414), .dout(n6637));
  jor  g06382(.dina(n6637), .dinb(n6636), .dout(n6638));
  jand g06383(.dina(n6577), .dinb(n6443), .dout(n6639));
  jnot g06384(.din(n6639), .dout(n6640));
  jnot g06385(.din(n6578), .dout(n6641));
  jor  g06386(.dina(n6641), .dinb(n6434), .dout(n6642));
  jand g06387(.dina(n6642), .dinb(n6640), .dout(n6643));
  jor  g06388(.dina(n3032), .dinb(n1566), .dout(n6644));
  jor  g06389(.dina(n1489), .dinb(n2579), .dout(n6645));
  jor  g06390(.dina(n1569), .dinb(n2870), .dout(n6646));
  jor  g06391(.dina(n1571), .dinb(n3035), .dout(n6647));
  jand g06392(.dina(n6647), .dinb(n6646), .dout(n6648));
  jand g06393(.dina(n6648), .dinb(n6645), .dout(n6649));
  jand g06394(.dina(n6649), .dinb(n6644), .dout(n6650));
  jxor g06395(.dina(n6650), .dinb(a20 ), .dout(n6651));
  jnot g06396(.din(n6651), .dout(n6652));
  jor  g06397(.dina(n6575), .dinb(n6567), .dout(n6653));
  jnot g06398(.din(n6653), .dout(n6654));
  jand g06399(.dina(n6576), .dinb(n6446), .dout(n6655));
  jor  g06400(.dina(n6655), .dinb(n6654), .dout(n6656));
  jor  g06401(.dina(n2556), .dinb(n1939), .dout(n6657));
  jor  g06402(.dina(n1827), .dinb(n2148), .dout(n6658));
  jor  g06403(.dina(n1942), .dinb(n2407), .dout(n6659));
  jor  g06404(.dina(n1944), .dinb(n2559), .dout(n6660));
  jand g06405(.dina(n6660), .dinb(n6659), .dout(n6661));
  jand g06406(.dina(n6661), .dinb(n6658), .dout(n6662));
  jand g06407(.dina(n6662), .dinb(n6657), .dout(n6663));
  jxor g06408(.dina(n6663), .dinb(a23 ), .dout(n6664));
  jnot g06409(.din(n6664), .dout(n6665));
  jor  g06410(.dina(n6564), .dinb(n6556), .dout(n6666));
  jand g06411(.dina(n6565), .dinb(n6451), .dout(n6667));
  jnot g06412(.din(n6667), .dout(n6668));
  jand g06413(.dina(n6668), .dinb(n6666), .dout(n6669));
  jnot g06414(.din(n6669), .dout(n6670));
  jor  g06415(.dina(n6553), .dinb(n6545), .dout(n6671));
  jand g06416(.dina(n6554), .dinb(n6454), .dout(n6672));
  jnot g06417(.din(n6672), .dout(n6673));
  jand g06418(.dina(n6673), .dinb(n6671), .dout(n6674));
  jnot g06419(.din(n6674), .dout(n6675));
  jor  g06420(.dina(n6542), .dinb(n6534), .dout(n6676));
  jand g06421(.dina(n6543), .dinb(n6457), .dout(n6677));
  jnot g06422(.din(n6677), .dout(n6678));
  jand g06423(.dina(n6678), .dinb(n6676), .dout(n6679));
  jnot g06424(.din(n6679), .dout(n6680));
  jand g06425(.dina(n6531), .dinb(n6471), .dout(n6681));
  jand g06426(.dina(n6532), .dinb(n6462), .dout(n6682));
  jor  g06427(.dina(n6682), .dinb(n6681), .dout(n6683));
  jand g06428(.dina(n6529), .dinb(n6483), .dout(n6684));
  jand g06429(.dina(n6530), .dinb(n6474), .dout(n6685));
  jor  g06430(.dina(n6685), .dinb(n6684), .dout(n6686));
  jor  g06431(.dina(n4415), .dinb(n775), .dout(n6687));
  jor  g06432(.dina(n4272), .dinb(n647), .dout(n6688));
  jor  g06433(.dina(n4418), .dinb(n758), .dout(n6689));
  jor  g06434(.dina(n4420), .dinb(n778), .dout(n6690));
  jand g06435(.dina(n6690), .dinb(n6689), .dout(n6691));
  jand g06436(.dina(n6691), .dinb(n6688), .dout(n6692));
  jand g06437(.dina(n6692), .dinb(n6687), .dout(n6693));
  jxor g06438(.dina(n6693), .dinb(a38 ), .dout(n6694));
  jnot g06439(.din(n6694), .dout(n6695));
  jor  g06440(.dina(n6527), .dinb(n6519), .dout(n6696));
  jand g06441(.dina(n6528), .dinb(n6486), .dout(n6697));
  jnot g06442(.din(n6697), .dout(n6698));
  jand g06443(.dina(n6698), .dinb(n6696), .dout(n6699));
  jnot g06444(.din(n6699), .dout(n6700));
  jor  g06445(.dina(n6516), .dinb(n6508), .dout(n6701));
  jand g06446(.dina(n6517), .dinb(n6489), .dout(n6702));
  jnot g06447(.din(n6702), .dout(n6703));
  jand g06448(.dina(n6703), .dinb(n6701), .dout(n6704));
  jnot g06449(.din(n6704), .dout(n6705));
  jnot g06450(.din(n6505), .dout(n6706));
  jand g06451(.dina(n6706), .dinb(n6503), .dout(n6707));
  jand g06452(.dina(n6506), .dinb(n6501), .dout(n6708));
  jor  g06453(.dina(n6708), .dinb(n6707), .dout(n6709));
  jor  g06454(.dina(n6490), .dinb(n319), .dout(n6710));
  jor  g06455(.dina(n6262), .dinb(n279), .dout(n6711));
  jor  g06456(.dina(n6493), .dinb(n299), .dout(n6712));
  jor  g06457(.dina(n6495), .dinb(n322), .dout(n6713));
  jand g06458(.dina(n6713), .dinb(n6712), .dout(n6714));
  jand g06459(.dina(n6714), .dinb(n6711), .dout(n6715));
  jand g06460(.dina(n6715), .dinb(n6710), .dout(n6716));
  jxor g06461(.dina(n6716), .dinb(a47 ), .dout(n6717));
  jnot g06462(.din(n6717), .dout(n6718));
  jand g06463(.dina(n6503), .dinb(a50 ), .dout(n6719));
  jxor g06464(.dina(a50 ), .dinb(a49 ), .dout(n6720));
  jnot g06465(.din(n6720), .dout(n6721));
  jand g06466(.dina(n6721), .dinb(n6502), .dout(n6722));
  jand g06467(.dina(n6722), .dinb(b1 ), .dout(n6723));
  jnot g06468(.din(n6502), .dout(n6724));
  jxor g06469(.dina(a49 ), .dinb(a48 ), .dout(n6725));
  jand g06470(.dina(n6725), .dinb(n6724), .dout(n6726));
  jand g06471(.dina(n6726), .dinb(b0 ), .dout(n6727));
  jand g06472(.dina(n6720), .dinb(n6502), .dout(n6728));
  jand g06473(.dina(n6728), .dinb(n338), .dout(n6729));
  jor  g06474(.dina(n6729), .dinb(n6727), .dout(n6730));
  jor  g06475(.dina(n6730), .dinb(n6723), .dout(n6731));
  jxor g06476(.dina(n6731), .dinb(n6719), .dout(n6732));
  jxor g06477(.dina(n6732), .dinb(n6718), .dout(n6733));
  jxor g06478(.dina(n6733), .dinb(n6709), .dout(n6734));
  jnot g06479(.din(n6734), .dout(n6735));
  jor  g06480(.dina(n5739), .dinb(n428), .dout(n6736));
  jor  g06481(.dina(n5574), .dinb(n357), .dout(n6737));
  jor  g06482(.dina(n5742), .dinb(n395), .dout(n6738));
  jor  g06483(.dina(n5744), .dinb(n431), .dout(n6739));
  jand g06484(.dina(n6739), .dinb(n6738), .dout(n6740));
  jand g06485(.dina(n6740), .dinb(n6737), .dout(n6741));
  jand g06486(.dina(n6741), .dinb(n6736), .dout(n6742));
  jxor g06487(.dina(n6742), .dinb(a44 ), .dout(n6743));
  jxor g06488(.dina(n6743), .dinb(n6735), .dout(n6744));
  jxor g06489(.dina(n6744), .dinb(n6705), .dout(n6745));
  jnot g06490(.din(n6745), .dout(n6746));
  jor  g06491(.dina(n5096), .dinb(n624), .dout(n6747));
  jor  g06492(.dina(n4904), .dinb(n512), .dout(n6748));
  jor  g06493(.dina(n5099), .dinb(n564), .dout(n6749));
  jor  g06494(.dina(n5101), .dinb(n627), .dout(n6750));
  jand g06495(.dina(n6750), .dinb(n6749), .dout(n6751));
  jand g06496(.dina(n6751), .dinb(n6748), .dout(n6752));
  jand g06497(.dina(n6752), .dinb(n6747), .dout(n6753));
  jxor g06498(.dina(n6753), .dinb(a41 ), .dout(n6754));
  jxor g06499(.dina(n6754), .dinb(n6746), .dout(n6755));
  jxor g06500(.dina(n6755), .dinb(n6700), .dout(n6756));
  jxor g06501(.dina(n6756), .dinb(n6695), .dout(n6757));
  jxor g06502(.dina(n6757), .dinb(n6686), .dout(n6758));
  jnot g06503(.din(n6758), .dout(n6759));
  jor  g06504(.dina(n3849), .dinb(n1019), .dout(n6760));
  jor  g06505(.dina(n3689), .dinb(n858), .dout(n6761));
  jor  g06506(.dina(n3852), .dinb(n939), .dout(n6762));
  jor  g06507(.dina(n3854), .dinb(n1022), .dout(n6763));
  jand g06508(.dina(n6763), .dinb(n6762), .dout(n6764));
  jand g06509(.dina(n6764), .dinb(n6761), .dout(n6765));
  jand g06510(.dina(n6765), .dinb(n6760), .dout(n6766));
  jxor g06511(.dina(n6766), .dinb(a35 ), .dout(n6767));
  jxor g06512(.dina(n6767), .dinb(n6759), .dout(n6768));
  jxor g06513(.dina(n6768), .dinb(n6683), .dout(n6769));
  jnot g06514(.din(n6769), .dout(n6770));
  jor  g06515(.dina(n3301), .dinb(n1397), .dout(n6771));
  jor  g06516(.dina(n3136), .dinb(n1193), .dout(n6772));
  jor  g06517(.dina(n3304), .dinb(n1290), .dout(n6773));
  jor  g06518(.dina(n3306), .dinb(n1400), .dout(n6774));
  jand g06519(.dina(n6774), .dinb(n6773), .dout(n6775));
  jand g06520(.dina(n6775), .dinb(n6772), .dout(n6776));
  jand g06521(.dina(n6776), .dinb(n6771), .dout(n6777));
  jxor g06522(.dina(n6777), .dinb(a32 ), .dout(n6778));
  jxor g06523(.dina(n6778), .dinb(n6770), .dout(n6779));
  jxor g06524(.dina(n6779), .dinb(n6680), .dout(n6780));
  jnot g06525(.din(n6780), .dout(n6781));
  jor  g06526(.dina(n2784), .dinb(n1739), .dout(n6782));
  jor  g06527(.dina(n2661), .dinb(n1420), .dout(n6783));
  jor  g06528(.dina(n2787), .dinb(n1620), .dout(n6784));
  jor  g06529(.dina(n2789), .dinb(n1742), .dout(n6785));
  jand g06530(.dina(n6785), .dinb(n6784), .dout(n6786));
  jand g06531(.dina(n6786), .dinb(n6783), .dout(n6787));
  jand g06532(.dina(n6787), .dinb(n6782), .dout(n6788));
  jxor g06533(.dina(n6788), .dinb(a29 ), .dout(n6789));
  jxor g06534(.dina(n6789), .dinb(n6781), .dout(n6790));
  jxor g06535(.dina(n6790), .dinb(n6675), .dout(n6791));
  jnot g06536(.din(n6791), .dout(n6792));
  jor  g06537(.dina(n2319), .dinb(n2007), .dout(n6793));
  jor  g06538(.dina(n2224), .dinb(n1867), .dout(n6794));
  jor  g06539(.dina(n2322), .dinb(n1887), .dout(n6795));
  jor  g06540(.dina(n2324), .dinb(n2010), .dout(n6796));
  jand g06541(.dina(n6796), .dinb(n6795), .dout(n6797));
  jand g06542(.dina(n6797), .dinb(n6794), .dout(n6798));
  jand g06543(.dina(n6798), .dinb(n6793), .dout(n6799));
  jxor g06544(.dina(n6799), .dinb(a26 ), .dout(n6800));
  jxor g06545(.dina(n6800), .dinb(n6792), .dout(n6801));
  jxor g06546(.dina(n6801), .dinb(n6670), .dout(n6802));
  jxor g06547(.dina(n6802), .dinb(n6665), .dout(n6803));
  jxor g06548(.dina(n6803), .dinb(n6656), .dout(n6804));
  jxor g06549(.dina(n6804), .dinb(n6652), .dout(n6805));
  jxor g06550(.dina(n6805), .dinb(n6643), .dout(n6806));
  jor  g06551(.dina(n3400), .dinb(n1245), .dout(n6807));
  jor  g06552(.dina(n1165), .dinb(n3055), .dout(n6808));
  jor  g06553(.dina(n1248), .dinb(n3230), .dout(n6809));
  jor  g06554(.dina(n1250), .dinb(n3403), .dout(n6810));
  jand g06555(.dina(n6810), .dinb(n6809), .dout(n6811));
  jand g06556(.dina(n6811), .dinb(n6808), .dout(n6812));
  jand g06557(.dina(n6812), .dinb(n6807), .dout(n6813));
  jxor g06558(.dina(n6813), .dinb(a17 ), .dout(n6814));
  jxor g06559(.dina(n6814), .dinb(n6806), .dout(n6815));
  jxor g06560(.dina(n6815), .dinb(n6638), .dout(n6816));
  jnot g06561(.din(n6816), .dout(n6817));
  jor  g06562(.dina(n4137), .dinb(n974), .dout(n6818));
  jor  g06563(.dina(n908), .dinb(n3588), .dout(n6819));
  jor  g06564(.dina(n977), .dinb(n3942), .dout(n6820));
  jor  g06565(.dina(n979), .dinb(n4140), .dout(n6821));
  jand g06566(.dina(n6821), .dinb(n6820), .dout(n6822));
  jand g06567(.dina(n6822), .dinb(n6819), .dout(n6823));
  jand g06568(.dina(n6823), .dinb(n6818), .dout(n6824));
  jxor g06569(.dina(n6824), .dinb(a14 ), .dout(n6825));
  jxor g06570(.dina(n6825), .dinb(n6817), .dout(n6826));
  jxor g06571(.dina(n6826), .dinb(n6634), .dout(n6827));
  jor  g06572(.dina(n4554), .dinb(n706), .dout(n6828));
  jor  g06573(.dina(n683), .dinb(n4340), .dout(n6829));
  jor  g06574(.dina(n709), .dinb(n4537), .dout(n6830));
  jor  g06575(.dina(n711), .dinb(n4557), .dout(n6831));
  jand g06576(.dina(n6831), .dinb(n6830), .dout(n6832));
  jand g06577(.dina(n6832), .dinb(n6829), .dout(n6833));
  jand g06578(.dina(n6833), .dinb(n6828), .dout(n6834));
  jxor g06579(.dina(n6834), .dinb(a11 ), .dout(n6835));
  jxor g06580(.dina(n6835), .dinb(n6827), .dout(n6836));
  jxor g06581(.dina(n6836), .dinb(n6631), .dout(n6837));
  jnot g06582(.din(n6837), .dout(n6838));
  jor  g06583(.dina(n5405), .dinb(n528), .dout(n6839));
  jor  g06584(.dina(n490), .dinb(n4974), .dout(n6840));
  jor  g06585(.dina(n531), .dinb(n4994), .dout(n6841));
  jor  g06586(.dina(n533), .dinb(n5408), .dout(n6842));
  jand g06587(.dina(n6842), .dinb(n6841), .dout(n6843));
  jand g06588(.dina(n6843), .dinb(n6840), .dout(n6844));
  jand g06589(.dina(n6844), .dinb(n6839), .dout(n6845));
  jxor g06590(.dina(n6845), .dinb(a8 ), .dout(n6846));
  jxor g06591(.dina(n6846), .dinb(n6838), .dout(n6847));
  jxor g06592(.dina(n6847), .dinb(n6627), .dout(n6848));
  jor  g06593(.dina(n6103), .dinb(n402), .dout(n6849));
  jor  g06594(.dina(n371), .dinb(n5428), .dout(n6850));
  jor  g06595(.dina(n405), .dinb(n5862), .dout(n6851));
  jor  g06596(.dina(n332), .dinb(n6106), .dout(n6852));
  jand g06597(.dina(n6852), .dinb(n6851), .dout(n6853));
  jand g06598(.dina(n6853), .dinb(n6850), .dout(n6854));
  jand g06599(.dina(n6854), .dinb(n6849), .dout(n6855));
  jxor g06600(.dina(n6855), .dinb(a5 ), .dout(n6856));
  jxor g06601(.dina(n6856), .dinb(n6848), .dout(n6857));
  jxor g06602(.dina(n6857), .dinb(n6622), .dout(n6858));
  jand g06603(.dina(b48 ), .dinb(b47 ), .dout(n6859));
  jand g06604(.dina(n6367), .dinb(n6366), .dout(n6860));
  jor  g06605(.dina(n6860), .dinb(n6859), .dout(n6861));
  jxor g06606(.dina(b49 ), .dinb(b48 ), .dout(n6862));
  jnot g06607(.din(n6862), .dout(n6863));
  jxor g06608(.dina(n6863), .dinb(n6861), .dout(n6864));
  jor  g06609(.dina(n6864), .dinb(n264), .dout(n6865));
  jor  g06610(.dina(n284), .dinb(n6352), .dout(n6866));
  jnot g06611(.din(b49 ), .dout(n6867));
  jor  g06612(.dina(n269), .dinb(n6867), .dout(n6868));
  jor  g06613(.dina(n271), .dinb(n6372), .dout(n6869));
  jand g06614(.dina(n6869), .dinb(n6868), .dout(n6870));
  jand g06615(.dina(n6870), .dinb(n6866), .dout(n6871));
  jand g06616(.dina(n6871), .dinb(n6865), .dout(n6872));
  jxor g06617(.dina(n6872), .dinb(n260), .dout(n6873));
  jxor g06618(.dina(n6873), .dinb(n6858), .dout(n6874));
  jxor g06619(.dina(n6874), .dinb(n6619), .dout(f49 ));
  jand g06620(.dina(n6873), .dinb(n6858), .dout(n6876));
  jand g06621(.dina(n6874), .dinb(n6619), .dout(n6877));
  jor  g06622(.dina(n6877), .dinb(n6876), .dout(n6878));
  jor  g06623(.dina(n6856), .dinb(n6848), .dout(n6879));
  jnot g06624(.din(n6879), .dout(n6880));
  jand g06625(.dina(n6857), .dinb(n6622), .dout(n6881));
  jor  g06626(.dina(n6881), .dinb(n6880), .dout(n6882));
  jor  g06627(.dina(n6846), .dinb(n6838), .dout(n6883));
  jnot g06628(.din(n6883), .dout(n6884));
  jand g06629(.dina(n6847), .dinb(n6626), .dout(n6885));
  jor  g06630(.dina(n6885), .dinb(n6884), .dout(n6886));
  jnot g06631(.din(n6886), .dout(n6887));
  jnot g06632(.din(n6827), .dout(n6888));
  jor  g06633(.dina(n6835), .dinb(n6888), .dout(n6889));
  jor  g06634(.dina(n6836), .dinb(n6631), .dout(n6890));
  jand g06635(.dina(n6890), .dinb(n6889), .dout(n6891));
  jor  g06636(.dina(n6825), .dinb(n6817), .dout(n6892));
  jnot g06637(.din(n6892), .dout(n6893));
  jand g06638(.dina(n6826), .dinb(n6634), .dout(n6894));
  jor  g06639(.dina(n6894), .dinb(n6893), .dout(n6895));
  jor  g06640(.dina(n6814), .dinb(n6806), .dout(n6896));
  jnot g06641(.din(n6896), .dout(n6897));
  jand g06642(.dina(n6815), .dinb(n6638), .dout(n6898));
  jor  g06643(.dina(n6898), .dinb(n6897), .dout(n6899));
  jand g06644(.dina(n6804), .dinb(n6652), .dout(n6900));
  jnot g06645(.din(n6900), .dout(n6901));
  jnot g06646(.din(n6805), .dout(n6902));
  jor  g06647(.dina(n6902), .dinb(n6643), .dout(n6903));
  jand g06648(.dina(n6903), .dinb(n6901), .dout(n6904));
  jor  g06649(.dina(n3052), .dinb(n1566), .dout(n6905));
  jor  g06650(.dina(n1489), .dinb(n2870), .dout(n6906));
  jor  g06651(.dina(n1569), .dinb(n3035), .dout(n6907));
  jor  g06652(.dina(n1571), .dinb(n3055), .dout(n6908));
  jand g06653(.dina(n6908), .dinb(n6907), .dout(n6909));
  jand g06654(.dina(n6909), .dinb(n6906), .dout(n6910));
  jand g06655(.dina(n6910), .dinb(n6905), .dout(n6911));
  jxor g06656(.dina(n6911), .dinb(a20 ), .dout(n6912));
  jnot g06657(.din(n6912), .dout(n6913));
  jand g06658(.dina(n6802), .dinb(n6665), .dout(n6914));
  jand g06659(.dina(n6803), .dinb(n6656), .dout(n6915));
  jor  g06660(.dina(n6915), .dinb(n6914), .dout(n6916));
  jor  g06661(.dina(n2576), .dinb(n1939), .dout(n6917));
  jor  g06662(.dina(n1827), .dinb(n2407), .dout(n6918));
  jor  g06663(.dina(n1942), .dinb(n2559), .dout(n6919));
  jor  g06664(.dina(n1944), .dinb(n2579), .dout(n6920));
  jand g06665(.dina(n6920), .dinb(n6919), .dout(n6921));
  jand g06666(.dina(n6921), .dinb(n6918), .dout(n6922));
  jand g06667(.dina(n6922), .dinb(n6917), .dout(n6923));
  jxor g06668(.dina(n6923), .dinb(a23 ), .dout(n6924));
  jnot g06669(.din(n6924), .dout(n6925));
  jor  g06670(.dina(n6800), .dinb(n6792), .dout(n6926));
  jnot g06671(.din(n6926), .dout(n6927));
  jand g06672(.dina(n6801), .dinb(n6670), .dout(n6928));
  jor  g06673(.dina(n6928), .dinb(n6927), .dout(n6929));
  jor  g06674(.dina(n2145), .dinb(n2319), .dout(n6930));
  jor  g06675(.dina(n2224), .dinb(n1887), .dout(n6931));
  jor  g06676(.dina(n2322), .dinb(n2010), .dout(n6932));
  jor  g06677(.dina(n2324), .dinb(n2148), .dout(n6933));
  jand g06678(.dina(n6933), .dinb(n6932), .dout(n6934));
  jand g06679(.dina(n6934), .dinb(n6931), .dout(n6935));
  jand g06680(.dina(n6935), .dinb(n6930), .dout(n6936));
  jxor g06681(.dina(n6936), .dinb(a26 ), .dout(n6937));
  jnot g06682(.din(n6937), .dout(n6938));
  jor  g06683(.dina(n6789), .dinb(n6781), .dout(n6939));
  jand g06684(.dina(n6790), .dinb(n6675), .dout(n6940));
  jnot g06685(.din(n6940), .dout(n6941));
  jand g06686(.dina(n6941), .dinb(n6939), .dout(n6942));
  jnot g06687(.din(n6942), .dout(n6943));
  jor  g06688(.dina(n6778), .dinb(n6770), .dout(n6944));
  jand g06689(.dina(n6779), .dinb(n6680), .dout(n6945));
  jnot g06690(.din(n6945), .dout(n6946));
  jand g06691(.dina(n6946), .dinb(n6944), .dout(n6947));
  jnot g06692(.din(n6947), .dout(n6948));
  jor  g06693(.dina(n3301), .dinb(n1417), .dout(n6949));
  jor  g06694(.dina(n3136), .dinb(n1290), .dout(n6950));
  jor  g06695(.dina(n3304), .dinb(n1400), .dout(n6951));
  jor  g06696(.dina(n3306), .dinb(n1420), .dout(n6952));
  jand g06697(.dina(n6952), .dinb(n6951), .dout(n6953));
  jand g06698(.dina(n6953), .dinb(n6950), .dout(n6954));
  jand g06699(.dina(n6954), .dinb(n6949), .dout(n6955));
  jxor g06700(.dina(n6955), .dinb(a32 ), .dout(n6956));
  jnot g06701(.din(n6956), .dout(n6957));
  jor  g06702(.dina(n6767), .dinb(n6759), .dout(n6958));
  jand g06703(.dina(n6768), .dinb(n6683), .dout(n6959));
  jnot g06704(.din(n6959), .dout(n6960));
  jand g06705(.dina(n6960), .dinb(n6958), .dout(n6961));
  jnot g06706(.din(n6961), .dout(n6962));
  jor  g06707(.dina(n3849), .dinb(n1190), .dout(n6963));
  jor  g06708(.dina(n3689), .dinb(n939), .dout(n6964));
  jor  g06709(.dina(n3852), .dinb(n1022), .dout(n6965));
  jor  g06710(.dina(n3854), .dinb(n1193), .dout(n6966));
  jand g06711(.dina(n6966), .dinb(n6965), .dout(n6967));
  jand g06712(.dina(n6967), .dinb(n6964), .dout(n6968));
  jand g06713(.dina(n6968), .dinb(n6963), .dout(n6969));
  jxor g06714(.dina(n6969), .dinb(a35 ), .dout(n6970));
  jnot g06715(.din(n6970), .dout(n6971));
  jand g06716(.dina(n6756), .dinb(n6695), .dout(n6972));
  jand g06717(.dina(n6757), .dinb(n6686), .dout(n6973));
  jor  g06718(.dina(n6973), .dinb(n6972), .dout(n6974));
  jor  g06719(.dina(n6754), .dinb(n6746), .dout(n6975));
  jand g06720(.dina(n6755), .dinb(n6700), .dout(n6976));
  jnot g06721(.din(n6976), .dout(n6977));
  jand g06722(.dina(n6977), .dinb(n6975), .dout(n6978));
  jnot g06723(.din(n6978), .dout(n6979));
  jor  g06724(.dina(n5096), .dinb(n644), .dout(n6980));
  jor  g06725(.dina(n4904), .dinb(n564), .dout(n6981));
  jor  g06726(.dina(n5099), .dinb(n627), .dout(n6982));
  jor  g06727(.dina(n5101), .dinb(n647), .dout(n6983));
  jand g06728(.dina(n6983), .dinb(n6982), .dout(n6984));
  jand g06729(.dina(n6984), .dinb(n6981), .dout(n6985));
  jand g06730(.dina(n6985), .dinb(n6980), .dout(n6986));
  jxor g06731(.dina(n6986), .dinb(a41 ), .dout(n6987));
  jnot g06732(.din(n6987), .dout(n6988));
  jor  g06733(.dina(n6743), .dinb(n6735), .dout(n6989));
  jand g06734(.dina(n6744), .dinb(n6705), .dout(n6990));
  jnot g06735(.din(n6990), .dout(n6991));
  jand g06736(.dina(n6991), .dinb(n6989), .dout(n6992));
  jnot g06737(.din(n6992), .dout(n6993));
  jor  g06738(.dina(n5739), .dinb(n509), .dout(n6994));
  jor  g06739(.dina(n5574), .dinb(n395), .dout(n6995));
  jor  g06740(.dina(n5742), .dinb(n431), .dout(n6996));
  jor  g06741(.dina(n5744), .dinb(n512), .dout(n6997));
  jand g06742(.dina(n6997), .dinb(n6996), .dout(n6998));
  jand g06743(.dina(n6998), .dinb(n6995), .dout(n6999));
  jand g06744(.dina(n6999), .dinb(n6994), .dout(n7000));
  jxor g06745(.dina(n7000), .dinb(a44 ), .dout(n7001));
  jnot g06746(.din(n7001), .dout(n7002));
  jand g06747(.dina(n6732), .dinb(n6718), .dout(n7003));
  jand g06748(.dina(n6733), .dinb(n6709), .dout(n7004));
  jor  g06749(.dina(n7004), .dinb(n7003), .dout(n7005));
  jor  g06750(.dina(n6490), .dinb(n354), .dout(n7006));
  jor  g06751(.dina(n6262), .dinb(n299), .dout(n7007));
  jor  g06752(.dina(n6493), .dinb(n322), .dout(n7008));
  jor  g06753(.dina(n6495), .dinb(n357), .dout(n7009));
  jand g06754(.dina(n7009), .dinb(n7008), .dout(n7010));
  jand g06755(.dina(n7010), .dinb(n7007), .dout(n7011));
  jand g06756(.dina(n7011), .dinb(n7006), .dout(n7012));
  jxor g06757(.dina(n7012), .dinb(a47 ), .dout(n7013));
  jnot g06758(.din(n7013), .dout(n7014));
  jnot g06759(.din(n6731), .dout(n7015));
  jand g06760(.dina(n6504), .dinb(a50 ), .dout(n7016));
  jand g06761(.dina(n7016), .dinb(n7015), .dout(n7017));
  jnot g06762(.din(n7017), .dout(n7018));
  jand g06763(.dina(n7018), .dinb(a50 ), .dout(n7019));
  jor  g06764(.dina(n6725), .dinb(n6721), .dout(n7020));
  jor  g06765(.dina(n7020), .dinb(n6502), .dout(n7021));
  jnot g06766(.din(n7021), .dout(n7022));
  jand g06767(.dina(n7022), .dinb(b0 ), .dout(n7023));
  jand g06768(.dina(n6722), .dinb(b2 ), .dout(n7024));
  jand g06769(.dina(n6726), .dinb(b1 ), .dout(n7025));
  jand g06770(.dina(n6728), .dinb(n375), .dout(n7026));
  jor  g06771(.dina(n7026), .dinb(n7025), .dout(n7027));
  jor  g06772(.dina(n7027), .dinb(n7024), .dout(n7028));
  jor  g06773(.dina(n7028), .dinb(n7023), .dout(n7029));
  jxor g06774(.dina(n7029), .dinb(n7019), .dout(n7030));
  jxor g06775(.dina(n7030), .dinb(n7014), .dout(n7031));
  jxor g06776(.dina(n7031), .dinb(n7005), .dout(n7032));
  jxor g06777(.dina(n7032), .dinb(n7002), .dout(n7033));
  jxor g06778(.dina(n7033), .dinb(n6993), .dout(n7034));
  jxor g06779(.dina(n7034), .dinb(n6988), .dout(n7035));
  jxor g06780(.dina(n7035), .dinb(n6979), .dout(n7036));
  jnot g06781(.din(n7036), .dout(n7037));
  jor  g06782(.dina(n4415), .dinb(n855), .dout(n7038));
  jor  g06783(.dina(n4272), .dinb(n758), .dout(n7039));
  jor  g06784(.dina(n4418), .dinb(n778), .dout(n7040));
  jor  g06785(.dina(n4420), .dinb(n858), .dout(n7041));
  jand g06786(.dina(n7041), .dinb(n7040), .dout(n7042));
  jand g06787(.dina(n7042), .dinb(n7039), .dout(n7043));
  jand g06788(.dina(n7043), .dinb(n7038), .dout(n7044));
  jxor g06789(.dina(n7044), .dinb(a38 ), .dout(n7045));
  jxor g06790(.dina(n7045), .dinb(n7037), .dout(n7046));
  jxor g06791(.dina(n7046), .dinb(n6974), .dout(n7047));
  jxor g06792(.dina(n7047), .dinb(n6971), .dout(n7048));
  jxor g06793(.dina(n7048), .dinb(n6962), .dout(n7049));
  jxor g06794(.dina(n7049), .dinb(n6957), .dout(n7050));
  jxor g06795(.dina(n7050), .dinb(n6948), .dout(n7051));
  jnot g06796(.din(n7051), .dout(n7052));
  jor  g06797(.dina(n2784), .dinb(n1864), .dout(n7053));
  jor  g06798(.dina(n2661), .dinb(n1620), .dout(n7054));
  jor  g06799(.dina(n2787), .dinb(n1742), .dout(n7055));
  jor  g06800(.dina(n2789), .dinb(n1867), .dout(n7056));
  jand g06801(.dina(n7056), .dinb(n7055), .dout(n7057));
  jand g06802(.dina(n7057), .dinb(n7054), .dout(n7058));
  jand g06803(.dina(n7058), .dinb(n7053), .dout(n7059));
  jxor g06804(.dina(n7059), .dinb(a29 ), .dout(n7060));
  jxor g06805(.dina(n7060), .dinb(n7052), .dout(n7061));
  jxor g06806(.dina(n7061), .dinb(n6943), .dout(n7062));
  jxor g06807(.dina(n7062), .dinb(n6938), .dout(n7063));
  jxor g06808(.dina(n7063), .dinb(n6929), .dout(n7064));
  jxor g06809(.dina(n7064), .dinb(n6925), .dout(n7065));
  jxor g06810(.dina(n7065), .dinb(n6916), .dout(n7066));
  jxor g06811(.dina(n7066), .dinb(n6913), .dout(n7067));
  jxor g06812(.dina(n7067), .dinb(n6904), .dout(n7068));
  jor  g06813(.dina(n3585), .dinb(n1245), .dout(n7069));
  jor  g06814(.dina(n1165), .dinb(n3230), .dout(n7070));
  jor  g06815(.dina(n1248), .dinb(n3403), .dout(n7071));
  jor  g06816(.dina(n1250), .dinb(n3588), .dout(n7072));
  jand g06817(.dina(n7072), .dinb(n7071), .dout(n7073));
  jand g06818(.dina(n7073), .dinb(n7070), .dout(n7074));
  jand g06819(.dina(n7074), .dinb(n7069), .dout(n7075));
  jxor g06820(.dina(n7075), .dinb(a17 ), .dout(n7076));
  jxor g06821(.dina(n7076), .dinb(n7068), .dout(n7077));
  jxor g06822(.dina(n7077), .dinb(n6899), .dout(n7078));
  jnot g06823(.din(n7078), .dout(n7079));
  jor  g06824(.dina(n4337), .dinb(n974), .dout(n7080));
  jor  g06825(.dina(n908), .dinb(n3942), .dout(n7081));
  jor  g06826(.dina(n977), .dinb(n4140), .dout(n7082));
  jor  g06827(.dina(n979), .dinb(n4340), .dout(n7083));
  jand g06828(.dina(n7083), .dinb(n7082), .dout(n7084));
  jand g06829(.dina(n7084), .dinb(n7081), .dout(n7085));
  jand g06830(.dina(n7085), .dinb(n7080), .dout(n7086));
  jxor g06831(.dina(n7086), .dinb(a14 ), .dout(n7087));
  jxor g06832(.dina(n7087), .dinb(n7079), .dout(n7088));
  jxor g06833(.dina(n7088), .dinb(n6895), .dout(n7089));
  jor  g06834(.dina(n4971), .dinb(n706), .dout(n7090));
  jor  g06835(.dina(n683), .dinb(n4537), .dout(n7091));
  jor  g06836(.dina(n709), .dinb(n4557), .dout(n7092));
  jor  g06837(.dina(n711), .dinb(n4974), .dout(n7093));
  jand g06838(.dina(n7093), .dinb(n7092), .dout(n7094));
  jand g06839(.dina(n7094), .dinb(n7091), .dout(n7095));
  jand g06840(.dina(n7095), .dinb(n7090), .dout(n7096));
  jxor g06841(.dina(n7096), .dinb(a11 ), .dout(n7097));
  jxor g06842(.dina(n7097), .dinb(n7089), .dout(n7098));
  jxor g06843(.dina(n7098), .dinb(n6891), .dout(n7099));
  jnot g06844(.din(n7099), .dout(n7100));
  jor  g06845(.dina(n5425), .dinb(n528), .dout(n7101));
  jor  g06846(.dina(n490), .dinb(n4994), .dout(n7102));
  jor  g06847(.dina(n531), .dinb(n5408), .dout(n7103));
  jor  g06848(.dina(n533), .dinb(n5428), .dout(n7104));
  jand g06849(.dina(n7104), .dinb(n7103), .dout(n7105));
  jand g06850(.dina(n7105), .dinb(n7102), .dout(n7106));
  jand g06851(.dina(n7106), .dinb(n7101), .dout(n7107));
  jxor g06852(.dina(n7107), .dinb(a8 ), .dout(n7108));
  jxor g06853(.dina(n7108), .dinb(n7100), .dout(n7109));
  jxor g06854(.dina(n7109), .dinb(n6887), .dout(n7110));
  jor  g06855(.dina(n6349), .dinb(n402), .dout(n7111));
  jor  g06856(.dina(n371), .dinb(n5862), .dout(n7112));
  jor  g06857(.dina(n405), .dinb(n6106), .dout(n7113));
  jor  g06858(.dina(n332), .dinb(n6352), .dout(n7114));
  jand g06859(.dina(n7114), .dinb(n7113), .dout(n7115));
  jand g06860(.dina(n7115), .dinb(n7112), .dout(n7116));
  jand g06861(.dina(n7116), .dinb(n7111), .dout(n7117));
  jxor g06862(.dina(n7117), .dinb(a5 ), .dout(n7118));
  jxor g06863(.dina(n7118), .dinb(n7110), .dout(n7119));
  jxor g06864(.dina(n7119), .dinb(n6882), .dout(n7120));
  jand g06865(.dina(b49 ), .dinb(b48 ), .dout(n7121));
  jand g06866(.dina(n6862), .dinb(n6861), .dout(n7122));
  jor  g06867(.dina(n7122), .dinb(n7121), .dout(n7123));
  jxor g06868(.dina(b50 ), .dinb(b49 ), .dout(n7124));
  jnot g06869(.din(n7124), .dout(n7125));
  jxor g06870(.dina(n7125), .dinb(n7123), .dout(n7126));
  jor  g06871(.dina(n7126), .dinb(n264), .dout(n7127));
  jor  g06872(.dina(n284), .dinb(n6372), .dout(n7128));
  jnot g06873(.din(b50 ), .dout(n7129));
  jor  g06874(.dina(n269), .dinb(n7129), .dout(n7130));
  jor  g06875(.dina(n271), .dinb(n6867), .dout(n7131));
  jand g06876(.dina(n7131), .dinb(n7130), .dout(n7132));
  jand g06877(.dina(n7132), .dinb(n7128), .dout(n7133));
  jand g06878(.dina(n7133), .dinb(n7127), .dout(n7134));
  jxor g06879(.dina(n7134), .dinb(n260), .dout(n7135));
  jxor g06880(.dina(n7135), .dinb(n7120), .dout(n7136));
  jxor g06881(.dina(n7136), .dinb(n6878), .dout(f50 ));
  jand g06882(.dina(n7135), .dinb(n7120), .dout(n7138));
  jand g06883(.dina(n7136), .dinb(n6878), .dout(n7139));
  jor  g06884(.dina(n7139), .dinb(n7138), .dout(n7140));
  jand g06885(.dina(b50 ), .dinb(b49 ), .dout(n7141));
  jand g06886(.dina(n7124), .dinb(n7123), .dout(n7142));
  jor  g06887(.dina(n7142), .dinb(n7141), .dout(n7143));
  jxor g06888(.dina(b51 ), .dinb(b50 ), .dout(n7144));
  jnot g06889(.din(n7144), .dout(n7145));
  jxor g06890(.dina(n7145), .dinb(n7143), .dout(n7146));
  jor  g06891(.dina(n7146), .dinb(n264), .dout(n7147));
  jor  g06892(.dina(n284), .dinb(n6867), .dout(n7148));
  jnot g06893(.din(b51 ), .dout(n7149));
  jor  g06894(.dina(n269), .dinb(n7149), .dout(n7150));
  jor  g06895(.dina(n271), .dinb(n7129), .dout(n7151));
  jand g06896(.dina(n7151), .dinb(n7150), .dout(n7152));
  jand g06897(.dina(n7152), .dinb(n7148), .dout(n7153));
  jand g06898(.dina(n7153), .dinb(n7147), .dout(n7154));
  jxor g06899(.dina(n7154), .dinb(n260), .dout(n7155));
  jor  g06900(.dina(n7118), .dinb(n7110), .dout(n7156));
  jnot g06901(.din(n7156), .dout(n7157));
  jand g06902(.dina(n7119), .dinb(n6882), .dout(n7158));
  jor  g06903(.dina(n7158), .dinb(n7157), .dout(n7159));
  jor  g06904(.dina(n6369), .dinb(n402), .dout(n7160));
  jor  g06905(.dina(n371), .dinb(n6106), .dout(n7161));
  jor  g06906(.dina(n405), .dinb(n6352), .dout(n7162));
  jor  g06907(.dina(n332), .dinb(n6372), .dout(n7163));
  jand g06908(.dina(n7163), .dinb(n7162), .dout(n7164));
  jand g06909(.dina(n7164), .dinb(n7161), .dout(n7165));
  jand g06910(.dina(n7165), .dinb(n7160), .dout(n7166));
  jxor g06911(.dina(n7166), .dinb(a5 ), .dout(n7167));
  jnot g06912(.din(n7167), .dout(n7168));
  jor  g06913(.dina(n7108), .dinb(n7100), .dout(n7169));
  jnot g06914(.din(n7169), .dout(n7170));
  jand g06915(.dina(n7109), .dinb(n6886), .dout(n7171));
  jor  g06916(.dina(n7171), .dinb(n7170), .dout(n7172));
  jor  g06917(.dina(n7087), .dinb(n7079), .dout(n7173));
  jnot g06918(.din(n7173), .dout(n7174));
  jand g06919(.dina(n7088), .dinb(n6895), .dout(n7175));
  jor  g06920(.dina(n7175), .dinb(n7174), .dout(n7176));
  jor  g06921(.dina(n7076), .dinb(n7068), .dout(n7177));
  jnot g06922(.din(n7177), .dout(n7178));
  jand g06923(.dina(n7077), .dinb(n6899), .dout(n7179));
  jor  g06924(.dina(n7179), .dinb(n7178), .dout(n7180));
  jor  g06925(.dina(n3939), .dinb(n1245), .dout(n7181));
  jor  g06926(.dina(n1165), .dinb(n3403), .dout(n7182));
  jor  g06927(.dina(n1248), .dinb(n3588), .dout(n7183));
  jor  g06928(.dina(n1250), .dinb(n3942), .dout(n7184));
  jand g06929(.dina(n7184), .dinb(n7183), .dout(n7185));
  jand g06930(.dina(n7185), .dinb(n7182), .dout(n7186));
  jand g06931(.dina(n7186), .dinb(n7181), .dout(n7187));
  jxor g06932(.dina(n7187), .dinb(a17 ), .dout(n7188));
  jnot g06933(.din(n7188), .dout(n7189));
  jand g06934(.dina(n7066), .dinb(n6913), .dout(n7190));
  jand g06935(.dina(n6306), .dinb(n6157), .dout(n7191));
  jor  g06936(.dina(n7191), .dinb(n6415), .dout(n7192));
  jand g06937(.dina(n6578), .dinb(n7192), .dout(n7193));
  jor  g06938(.dina(n7193), .dinb(n6639), .dout(n7194));
  jand g06939(.dina(n6805), .dinb(n7194), .dout(n7195));
  jor  g06940(.dina(n7195), .dinb(n6900), .dout(n7196));
  jand g06941(.dina(n7067), .dinb(n7196), .dout(n7197));
  jor  g06942(.dina(n7197), .dinb(n7190), .dout(n7198));
  jand g06943(.dina(n7064), .dinb(n6925), .dout(n7199));
  jand g06944(.dina(n7065), .dinb(n6916), .dout(n7200));
  jor  g06945(.dina(n7200), .dinb(n7199), .dout(n7201));
  jor  g06946(.dina(n2867), .dinb(n1939), .dout(n7202));
  jor  g06947(.dina(n1827), .dinb(n2559), .dout(n7203));
  jor  g06948(.dina(n1942), .dinb(n2579), .dout(n7204));
  jor  g06949(.dina(n1944), .dinb(n2870), .dout(n7205));
  jand g06950(.dina(n7205), .dinb(n7204), .dout(n7206));
  jand g06951(.dina(n7206), .dinb(n7203), .dout(n7207));
  jand g06952(.dina(n7207), .dinb(n7202), .dout(n7208));
  jxor g06953(.dina(n7208), .dinb(a23 ), .dout(n7209));
  jnot g06954(.din(n7209), .dout(n7210));
  jand g06955(.dina(n7062), .dinb(n6938), .dout(n7211));
  jand g06956(.dina(n7063), .dinb(n6929), .dout(n7212));
  jor  g06957(.dina(n7212), .dinb(n7211), .dout(n7213));
  jor  g06958(.dina(n7060), .dinb(n7052), .dout(n7214));
  jand g06959(.dina(n7061), .dinb(n6943), .dout(n7215));
  jnot g06960(.din(n7215), .dout(n7216));
  jand g06961(.dina(n7216), .dinb(n7214), .dout(n7217));
  jnot g06962(.din(n7217), .dout(n7218));
  jand g06963(.dina(n7049), .dinb(n6957), .dout(n7219));
  jand g06964(.dina(n7050), .dinb(n6948), .dout(n7220));
  jor  g06965(.dina(n7220), .dinb(n7219), .dout(n7221));
  jand g06966(.dina(n7047), .dinb(n6971), .dout(n7222));
  jand g06967(.dina(n7048), .dinb(n6962), .dout(n7223));
  jor  g06968(.dina(n7223), .dinb(n7222), .dout(n7224));
  jor  g06969(.dina(n3849), .dinb(n1287), .dout(n7225));
  jor  g06970(.dina(n3689), .dinb(n1022), .dout(n7226));
  jor  g06971(.dina(n3852), .dinb(n1193), .dout(n7227));
  jor  g06972(.dina(n3854), .dinb(n1290), .dout(n7228));
  jand g06973(.dina(n7228), .dinb(n7227), .dout(n7229));
  jand g06974(.dina(n7229), .dinb(n7226), .dout(n7230));
  jand g06975(.dina(n7230), .dinb(n7225), .dout(n7231));
  jxor g06976(.dina(n7231), .dinb(a35 ), .dout(n7232));
  jnot g06977(.din(n7232), .dout(n7233));
  jor  g06978(.dina(n7045), .dinb(n7037), .dout(n7234));
  jand g06979(.dina(n7046), .dinb(n6974), .dout(n7235));
  jnot g06980(.din(n7235), .dout(n7236));
  jand g06981(.dina(n7236), .dinb(n7234), .dout(n7237));
  jnot g06982(.din(n7237), .dout(n7238));
  jor  g06983(.dina(n4415), .dinb(n936), .dout(n7239));
  jor  g06984(.dina(n4272), .dinb(n778), .dout(n7240));
  jor  g06985(.dina(n4418), .dinb(n858), .dout(n7241));
  jor  g06986(.dina(n4420), .dinb(n939), .dout(n7242));
  jand g06987(.dina(n7242), .dinb(n7241), .dout(n7243));
  jand g06988(.dina(n7243), .dinb(n7240), .dout(n7244));
  jand g06989(.dina(n7244), .dinb(n7239), .dout(n7245));
  jxor g06990(.dina(n7245), .dinb(a38 ), .dout(n7246));
  jnot g06991(.din(n7246), .dout(n7247));
  jand g06992(.dina(n7034), .dinb(n6988), .dout(n7248));
  jand g06993(.dina(n7035), .dinb(n6979), .dout(n7249));
  jor  g06994(.dina(n7249), .dinb(n7248), .dout(n7250));
  jor  g06995(.dina(n5096), .dinb(n755), .dout(n7251));
  jor  g06996(.dina(n4904), .dinb(n627), .dout(n7252));
  jor  g06997(.dina(n5099), .dinb(n647), .dout(n7253));
  jor  g06998(.dina(n5101), .dinb(n758), .dout(n7254));
  jand g06999(.dina(n7254), .dinb(n7253), .dout(n7255));
  jand g07000(.dina(n7255), .dinb(n7252), .dout(n7256));
  jand g07001(.dina(n7256), .dinb(n7251), .dout(n7257));
  jxor g07002(.dina(n7257), .dinb(a41 ), .dout(n7258));
  jnot g07003(.din(n7258), .dout(n7259));
  jand g07004(.dina(n7032), .dinb(n7002), .dout(n7260));
  jand g07005(.dina(n7033), .dinb(n6993), .dout(n7261));
  jor  g07006(.dina(n7261), .dinb(n7260), .dout(n7262));
  jand g07007(.dina(n7030), .dinb(n7014), .dout(n7263));
  jand g07008(.dina(n7031), .dinb(n7005), .dout(n7264));
  jor  g07009(.dina(n7264), .dinb(n7263), .dout(n7265));
  jnot g07010(.din(n6728), .dout(n7266));
  jor  g07011(.dina(n7266), .dinb(n296), .dout(n7267));
  jor  g07012(.dina(n7021), .dinb(n267), .dout(n7268));
  jnot g07013(.din(n6726), .dout(n7269));
  jor  g07014(.dina(n7269), .dinb(n279), .dout(n7270));
  jnot g07015(.din(n6722), .dout(n7271));
  jor  g07016(.dina(n7271), .dinb(n299), .dout(n7272));
  jand g07017(.dina(n7272), .dinb(n7270), .dout(n7273));
  jand g07018(.dina(n7273), .dinb(n7268), .dout(n7274));
  jand g07019(.dina(n7274), .dinb(n7267), .dout(n7275));
  jxor g07020(.dina(n7275), .dinb(a50 ), .dout(n7276));
  jnot g07021(.din(n7276), .dout(n7277));
  jxor g07022(.dina(a51 ), .dinb(a50 ), .dout(n7278));
  jand g07023(.dina(n7278), .dinb(b0 ), .dout(n7279));
  jnot g07024(.din(n7279), .dout(n7280));
  jor  g07025(.dina(n7029), .dinb(n7018), .dout(n7281));
  jxor g07026(.dina(n7281), .dinb(n7280), .dout(n7282));
  jxor g07027(.dina(n7282), .dinb(n7277), .dout(n7283));
  jnot g07028(.din(n7283), .dout(n7284));
  jor  g07029(.dina(n6490), .dinb(n392), .dout(n7285));
  jor  g07030(.dina(n6262), .dinb(n322), .dout(n7286));
  jor  g07031(.dina(n6493), .dinb(n357), .dout(n7287));
  jor  g07032(.dina(n6495), .dinb(n395), .dout(n7288));
  jand g07033(.dina(n7288), .dinb(n7287), .dout(n7289));
  jand g07034(.dina(n7289), .dinb(n7286), .dout(n7290));
  jand g07035(.dina(n7290), .dinb(n7285), .dout(n7291));
  jxor g07036(.dina(n7291), .dinb(a47 ), .dout(n7292));
  jxor g07037(.dina(n7292), .dinb(n7284), .dout(n7293));
  jxor g07038(.dina(n7293), .dinb(n7265), .dout(n7294));
  jnot g07039(.din(n7294), .dout(n7295));
  jor  g07040(.dina(n5739), .dinb(n561), .dout(n7296));
  jor  g07041(.dina(n5574), .dinb(n431), .dout(n7297));
  jor  g07042(.dina(n5742), .dinb(n512), .dout(n7298));
  jor  g07043(.dina(n5744), .dinb(n564), .dout(n7299));
  jand g07044(.dina(n7299), .dinb(n7298), .dout(n7300));
  jand g07045(.dina(n7300), .dinb(n7297), .dout(n7301));
  jand g07046(.dina(n7301), .dinb(n7296), .dout(n7302));
  jxor g07047(.dina(n7302), .dinb(a44 ), .dout(n7303));
  jxor g07048(.dina(n7303), .dinb(n7295), .dout(n7304));
  jxor g07049(.dina(n7304), .dinb(n7262), .dout(n7305));
  jxor g07050(.dina(n7305), .dinb(n7259), .dout(n7306));
  jxor g07051(.dina(n7306), .dinb(n7250), .dout(n7307));
  jxor g07052(.dina(n7307), .dinb(n7247), .dout(n7308));
  jxor g07053(.dina(n7308), .dinb(n7238), .dout(n7309));
  jxor g07054(.dina(n7309), .dinb(n7233), .dout(n7310));
  jxor g07055(.dina(n7310), .dinb(n7224), .dout(n7311));
  jnot g07056(.din(n7311), .dout(n7312));
  jor  g07057(.dina(n3301), .dinb(n1617), .dout(n7313));
  jor  g07058(.dina(n3136), .dinb(n1400), .dout(n7314));
  jor  g07059(.dina(n3304), .dinb(n1420), .dout(n7315));
  jor  g07060(.dina(n3306), .dinb(n1620), .dout(n7316));
  jand g07061(.dina(n7316), .dinb(n7315), .dout(n7317));
  jand g07062(.dina(n7317), .dinb(n7314), .dout(n7318));
  jand g07063(.dina(n7318), .dinb(n7313), .dout(n7319));
  jxor g07064(.dina(n7319), .dinb(a32 ), .dout(n7320));
  jxor g07065(.dina(n7320), .dinb(n7312), .dout(n7321));
  jxor g07066(.dina(n7321), .dinb(n7221), .dout(n7322));
  jnot g07067(.din(n7322), .dout(n7323));
  jor  g07068(.dina(n2784), .dinb(n1884), .dout(n7324));
  jor  g07069(.dina(n2661), .dinb(n1742), .dout(n7325));
  jor  g07070(.dina(n2787), .dinb(n1867), .dout(n7326));
  jor  g07071(.dina(n2789), .dinb(n1887), .dout(n7327));
  jand g07072(.dina(n7327), .dinb(n7326), .dout(n7328));
  jand g07073(.dina(n7328), .dinb(n7325), .dout(n7329));
  jand g07074(.dina(n7329), .dinb(n7324), .dout(n7330));
  jxor g07075(.dina(n7330), .dinb(a29 ), .dout(n7331));
  jxor g07076(.dina(n7331), .dinb(n7323), .dout(n7332));
  jxor g07077(.dina(n7332), .dinb(n7218), .dout(n7333));
  jnot g07078(.din(n7333), .dout(n7334));
  jor  g07079(.dina(n2404), .dinb(n2319), .dout(n7335));
  jor  g07080(.dina(n2224), .dinb(n2010), .dout(n7336));
  jor  g07081(.dina(n2322), .dinb(n2148), .dout(n7337));
  jor  g07082(.dina(n2324), .dinb(n2407), .dout(n7338));
  jand g07083(.dina(n7338), .dinb(n7337), .dout(n7339));
  jand g07084(.dina(n7339), .dinb(n7336), .dout(n7340));
  jand g07085(.dina(n7340), .dinb(n7335), .dout(n7341));
  jxor g07086(.dina(n7341), .dinb(a26 ), .dout(n7342));
  jxor g07087(.dina(n7342), .dinb(n7334), .dout(n7343));
  jxor g07088(.dina(n7343), .dinb(n7213), .dout(n7344));
  jxor g07089(.dina(n7344), .dinb(n7210), .dout(n7345));
  jxor g07090(.dina(n7345), .dinb(n7201), .dout(n7346));
  jor  g07091(.dina(n3227), .dinb(n1566), .dout(n7347));
  jor  g07092(.dina(n1489), .dinb(n3035), .dout(n7348));
  jor  g07093(.dina(n1569), .dinb(n3055), .dout(n7349));
  jor  g07094(.dina(n1571), .dinb(n3230), .dout(n7350));
  jand g07095(.dina(n7350), .dinb(n7349), .dout(n7351));
  jand g07096(.dina(n7351), .dinb(n7348), .dout(n7352));
  jand g07097(.dina(n7352), .dinb(n7347), .dout(n7353));
  jxor g07098(.dina(n7353), .dinb(a20 ), .dout(n7354));
  jxor g07099(.dina(n7354), .dinb(n7346), .dout(n7355));
  jnot g07100(.din(n7355), .dout(n7356));
  jxor g07101(.dina(n7356), .dinb(n7198), .dout(n7357));
  jxor g07102(.dina(n7357), .dinb(n7189), .dout(n7358));
  jxor g07103(.dina(n7358), .dinb(n7180), .dout(n7359));
  jnot g07104(.din(n7359), .dout(n7360));
  jor  g07105(.dina(n4534), .dinb(n974), .dout(n7361));
  jor  g07106(.dina(n908), .dinb(n4140), .dout(n7362));
  jor  g07107(.dina(n977), .dinb(n4340), .dout(n7363));
  jor  g07108(.dina(n979), .dinb(n4537), .dout(n7364));
  jand g07109(.dina(n7364), .dinb(n7363), .dout(n7365));
  jand g07110(.dina(n7365), .dinb(n7362), .dout(n7366));
  jand g07111(.dina(n7366), .dinb(n7361), .dout(n7367));
  jxor g07112(.dina(n7367), .dinb(a14 ), .dout(n7368));
  jxor g07113(.dina(n7368), .dinb(n7360), .dout(n7369));
  jxor g07114(.dina(n7369), .dinb(n7176), .dout(n7370));
  jor  g07115(.dina(n4991), .dinb(n706), .dout(n7371));
  jor  g07116(.dina(n683), .dinb(n4557), .dout(n7372));
  jor  g07117(.dina(n709), .dinb(n4974), .dout(n7373));
  jor  g07118(.dina(n711), .dinb(n4994), .dout(n7374));
  jand g07119(.dina(n7374), .dinb(n7373), .dout(n7375));
  jand g07120(.dina(n7375), .dinb(n7372), .dout(n7376));
  jand g07121(.dina(n7376), .dinb(n7371), .dout(n7377));
  jxor g07122(.dina(n7377), .dinb(a11 ), .dout(n7378));
  jxor g07123(.dina(n7378), .dinb(n7370), .dout(n7379));
  jnot g07124(.din(n7089), .dout(n7380));
  jor  g07125(.dina(n7097), .dinb(n7380), .dout(n7381));
  jor  g07126(.dina(n7098), .dinb(n6891), .dout(n7382));
  jand g07127(.dina(n7382), .dinb(n7381), .dout(n7383));
  jxor g07128(.dina(n7383), .dinb(n7379), .dout(n7384));
  jnot g07129(.din(n7384), .dout(n7385));
  jor  g07130(.dina(n5859), .dinb(n528), .dout(n7386));
  jor  g07131(.dina(n490), .dinb(n5408), .dout(n7387));
  jor  g07132(.dina(n531), .dinb(n5428), .dout(n7388));
  jor  g07133(.dina(n533), .dinb(n5862), .dout(n7389));
  jand g07134(.dina(n7389), .dinb(n7388), .dout(n7390));
  jand g07135(.dina(n7390), .dinb(n7387), .dout(n7391));
  jand g07136(.dina(n7391), .dinb(n7386), .dout(n7392));
  jxor g07137(.dina(n7392), .dinb(a8 ), .dout(n7393));
  jxor g07138(.dina(n7393), .dinb(n7385), .dout(n7394));
  jxor g07139(.dina(n7394), .dinb(n7172), .dout(n7395));
  jxor g07140(.dina(n7395), .dinb(n7168), .dout(n7396));
  jxor g07141(.dina(n7396), .dinb(n7159), .dout(n7397));
  jxor g07142(.dina(n7397), .dinb(n7155), .dout(n7398));
  jxor g07143(.dina(n7398), .dinb(n7140), .dout(f51 ));
  jand g07144(.dina(n7397), .dinb(n7155), .dout(n7400));
  jand g07145(.dina(n7398), .dinb(n7140), .dout(n7401));
  jor  g07146(.dina(n7401), .dinb(n7400), .dout(n7402));
  jand g07147(.dina(b51 ), .dinb(b50 ), .dout(n7403));
  jand g07148(.dina(n7144), .dinb(n7143), .dout(n7404));
  jor  g07149(.dina(n7404), .dinb(n7403), .dout(n7405));
  jxor g07150(.dina(b52 ), .dinb(b51 ), .dout(n7406));
  jnot g07151(.din(n7406), .dout(n7407));
  jxor g07152(.dina(n7407), .dinb(n7405), .dout(n7408));
  jor  g07153(.dina(n7408), .dinb(n264), .dout(n7409));
  jor  g07154(.dina(n284), .dinb(n7129), .dout(n7410));
  jnot g07155(.din(b52 ), .dout(n7411));
  jor  g07156(.dina(n269), .dinb(n7411), .dout(n7412));
  jor  g07157(.dina(n271), .dinb(n7149), .dout(n7413));
  jand g07158(.dina(n7413), .dinb(n7412), .dout(n7414));
  jand g07159(.dina(n7414), .dinb(n7410), .dout(n7415));
  jand g07160(.dina(n7415), .dinb(n7409), .dout(n7416));
  jxor g07161(.dina(n7416), .dinb(n260), .dout(n7417));
  jand g07162(.dina(n7395), .dinb(n7168), .dout(n7418));
  jand g07163(.dina(n7396), .dinb(n7159), .dout(n7419));
  jor  g07164(.dina(n7419), .dinb(n7418), .dout(n7420));
  jor  g07165(.dina(n7393), .dinb(n7385), .dout(n7421));
  jnot g07166(.din(n7421), .dout(n7422));
  jand g07167(.dina(n7394), .dinb(n7172), .dout(n7423));
  jor  g07168(.dina(n7423), .dinb(n7422), .dout(n7424));
  jnot g07169(.din(n7424), .dout(n7425));
  jnot g07170(.din(n7370), .dout(n7426));
  jor  g07171(.dina(n7378), .dinb(n7426), .dout(n7427));
  jor  g07172(.dina(n7383), .dinb(n7379), .dout(n7428));
  jand g07173(.dina(n7428), .dinb(n7427), .dout(n7429));
  jor  g07174(.dina(n7368), .dinb(n7360), .dout(n7430));
  jnot g07175(.din(n7430), .dout(n7431));
  jand g07176(.dina(n7369), .dinb(n7176), .dout(n7432));
  jor  g07177(.dina(n7432), .dinb(n7431), .dout(n7433));
  jand g07178(.dina(n7357), .dinb(n7189), .dout(n7434));
  jand g07179(.dina(n7358), .dinb(n7180), .dout(n7435));
  jor  g07180(.dina(n7435), .dinb(n7434), .dout(n7436));
  jnot g07181(.din(n7346), .dout(n7437));
  jor  g07182(.dina(n7354), .dinb(n7437), .dout(n7438));
  jnot g07183(.din(n7190), .dout(n7439));
  jnot g07184(.din(n7067), .dout(n7440));
  jor  g07185(.dina(n7440), .dinb(n6904), .dout(n7441));
  jand g07186(.dina(n7441), .dinb(n7439), .dout(n7442));
  jor  g07187(.dina(n7355), .dinb(n7442), .dout(n7443));
  jand g07188(.dina(n7443), .dinb(n7438), .dout(n7444));
  jand g07189(.dina(n7344), .dinb(n7210), .dout(n7445));
  jand g07190(.dina(n7345), .dinb(n7201), .dout(n7446));
  jor  g07191(.dina(n7446), .dinb(n7445), .dout(n7447));
  jor  g07192(.dina(n7342), .dinb(n7334), .dout(n7448));
  jnot g07193(.din(n7448), .dout(n7449));
  jand g07194(.dina(n7343), .dinb(n7213), .dout(n7450));
  jor  g07195(.dina(n7450), .dinb(n7449), .dout(n7451));
  jor  g07196(.dina(n2556), .dinb(n2319), .dout(n7452));
  jor  g07197(.dina(n2224), .dinb(n2148), .dout(n7453));
  jor  g07198(.dina(n2322), .dinb(n2407), .dout(n7454));
  jor  g07199(.dina(n2324), .dinb(n2559), .dout(n7455));
  jand g07200(.dina(n7455), .dinb(n7454), .dout(n7456));
  jand g07201(.dina(n7456), .dinb(n7453), .dout(n7457));
  jand g07202(.dina(n7457), .dinb(n7452), .dout(n7458));
  jxor g07203(.dina(n7458), .dinb(a26 ), .dout(n7459));
  jnot g07204(.din(n7459), .dout(n7460));
  jor  g07205(.dina(n7331), .dinb(n7323), .dout(n7461));
  jand g07206(.dina(n7332), .dinb(n7218), .dout(n7462));
  jnot g07207(.din(n7462), .dout(n7463));
  jand g07208(.dina(n7463), .dinb(n7461), .dout(n7464));
  jnot g07209(.din(n7464), .dout(n7465));
  jor  g07210(.dina(n7320), .dinb(n7312), .dout(n7466));
  jand g07211(.dina(n7321), .dinb(n7221), .dout(n7467));
  jnot g07212(.din(n7467), .dout(n7468));
  jand g07213(.dina(n7468), .dinb(n7466), .dout(n7469));
  jnot g07214(.din(n7469), .dout(n7470));
  jand g07215(.dina(n7309), .dinb(n7233), .dout(n7471));
  jand g07216(.dina(n7310), .dinb(n7224), .dout(n7472));
  jor  g07217(.dina(n7472), .dinb(n7471), .dout(n7473));
  jand g07218(.dina(n7307), .dinb(n7247), .dout(n7474));
  jand g07219(.dina(n7308), .dinb(n7238), .dout(n7475));
  jor  g07220(.dina(n7475), .dinb(n7474), .dout(n7476));
  jand g07221(.dina(n7305), .dinb(n7259), .dout(n7477));
  jand g07222(.dina(n7306), .dinb(n7250), .dout(n7478));
  jor  g07223(.dina(n7478), .dinb(n7477), .dout(n7479));
  jor  g07224(.dina(n5096), .dinb(n775), .dout(n7480));
  jor  g07225(.dina(n4904), .dinb(n647), .dout(n7481));
  jor  g07226(.dina(n5099), .dinb(n758), .dout(n7482));
  jor  g07227(.dina(n5101), .dinb(n778), .dout(n7483));
  jand g07228(.dina(n7483), .dinb(n7482), .dout(n7484));
  jand g07229(.dina(n7484), .dinb(n7481), .dout(n7485));
  jand g07230(.dina(n7485), .dinb(n7480), .dout(n7486));
  jxor g07231(.dina(n7486), .dinb(a41 ), .dout(n7487));
  jnot g07232(.din(n7487), .dout(n7488));
  jor  g07233(.dina(n7303), .dinb(n7295), .dout(n7489));
  jand g07234(.dina(n7304), .dinb(n7262), .dout(n7490));
  jnot g07235(.din(n7490), .dout(n7491));
  jand g07236(.dina(n7491), .dinb(n7489), .dout(n7492));
  jnot g07237(.din(n7492), .dout(n7493));
  jor  g07238(.dina(n7292), .dinb(n7284), .dout(n7494));
  jand g07239(.dina(n7293), .dinb(n7265), .dout(n7495));
  jnot g07240(.din(n7495), .dout(n7496));
  jand g07241(.dina(n7496), .dinb(n7494), .dout(n7497));
  jnot g07242(.din(n7497), .dout(n7498));
  jnot g07243(.din(n7281), .dout(n7499));
  jand g07244(.dina(n7499), .dinb(n7279), .dout(n7500));
  jand g07245(.dina(n7282), .dinb(n7277), .dout(n7501));
  jor  g07246(.dina(n7501), .dinb(n7500), .dout(n7502));
  jor  g07247(.dina(n7266), .dinb(n319), .dout(n7503));
  jor  g07248(.dina(n7021), .dinb(n279), .dout(n7504));
  jor  g07249(.dina(n7269), .dinb(n299), .dout(n7505));
  jor  g07250(.dina(n7271), .dinb(n322), .dout(n7506));
  jand g07251(.dina(n7506), .dinb(n7505), .dout(n7507));
  jand g07252(.dina(n7507), .dinb(n7504), .dout(n7508));
  jand g07253(.dina(n7508), .dinb(n7503), .dout(n7509));
  jxor g07254(.dina(n7509), .dinb(a50 ), .dout(n7510));
  jnot g07255(.din(n7510), .dout(n7511));
  jand g07256(.dina(n7279), .dinb(a53 ), .dout(n7512));
  jxor g07257(.dina(a53 ), .dinb(a52 ), .dout(n7513));
  jnot g07258(.din(n7513), .dout(n7514));
  jand g07259(.dina(n7514), .dinb(n7278), .dout(n7515));
  jand g07260(.dina(n7515), .dinb(b1 ), .dout(n7516));
  jnot g07261(.din(n7278), .dout(n7517));
  jxor g07262(.dina(a52 ), .dinb(a51 ), .dout(n7518));
  jand g07263(.dina(n7518), .dinb(n7517), .dout(n7519));
  jand g07264(.dina(n7519), .dinb(b0 ), .dout(n7520));
  jand g07265(.dina(n7513), .dinb(n7278), .dout(n7521));
  jand g07266(.dina(n7521), .dinb(n338), .dout(n7522));
  jor  g07267(.dina(n7522), .dinb(n7520), .dout(n7523));
  jor  g07268(.dina(n7523), .dinb(n7516), .dout(n7524));
  jxor g07269(.dina(n7524), .dinb(n7512), .dout(n7525));
  jxor g07270(.dina(n7525), .dinb(n7511), .dout(n7526));
  jxor g07271(.dina(n7526), .dinb(n7502), .dout(n7527));
  jnot g07272(.din(n7527), .dout(n7528));
  jor  g07273(.dina(n6490), .dinb(n428), .dout(n7529));
  jor  g07274(.dina(n6262), .dinb(n357), .dout(n7530));
  jor  g07275(.dina(n6493), .dinb(n395), .dout(n7531));
  jor  g07276(.dina(n6495), .dinb(n431), .dout(n7532));
  jand g07277(.dina(n7532), .dinb(n7531), .dout(n7533));
  jand g07278(.dina(n7533), .dinb(n7530), .dout(n7534));
  jand g07279(.dina(n7534), .dinb(n7529), .dout(n7535));
  jxor g07280(.dina(n7535), .dinb(a47 ), .dout(n7536));
  jxor g07281(.dina(n7536), .dinb(n7528), .dout(n7537));
  jxor g07282(.dina(n7537), .dinb(n7498), .dout(n7538));
  jnot g07283(.din(n7538), .dout(n7539));
  jor  g07284(.dina(n5739), .dinb(n624), .dout(n7540));
  jor  g07285(.dina(n5574), .dinb(n512), .dout(n7541));
  jor  g07286(.dina(n5742), .dinb(n564), .dout(n7542));
  jor  g07287(.dina(n5744), .dinb(n627), .dout(n7543));
  jand g07288(.dina(n7543), .dinb(n7542), .dout(n7544));
  jand g07289(.dina(n7544), .dinb(n7541), .dout(n7545));
  jand g07290(.dina(n7545), .dinb(n7540), .dout(n7546));
  jxor g07291(.dina(n7546), .dinb(a44 ), .dout(n7547));
  jxor g07292(.dina(n7547), .dinb(n7539), .dout(n7548));
  jxor g07293(.dina(n7548), .dinb(n7493), .dout(n7549));
  jxor g07294(.dina(n7549), .dinb(n7488), .dout(n7550));
  jxor g07295(.dina(n7550), .dinb(n7479), .dout(n7551));
  jnot g07296(.din(n7551), .dout(n7552));
  jor  g07297(.dina(n4415), .dinb(n1019), .dout(n7553));
  jor  g07298(.dina(n4272), .dinb(n858), .dout(n7554));
  jor  g07299(.dina(n4418), .dinb(n939), .dout(n7555));
  jor  g07300(.dina(n4420), .dinb(n1022), .dout(n7556));
  jand g07301(.dina(n7556), .dinb(n7555), .dout(n7557));
  jand g07302(.dina(n7557), .dinb(n7554), .dout(n7558));
  jand g07303(.dina(n7558), .dinb(n7553), .dout(n7559));
  jxor g07304(.dina(n7559), .dinb(a38 ), .dout(n7560));
  jxor g07305(.dina(n7560), .dinb(n7552), .dout(n7561));
  jxor g07306(.dina(n7561), .dinb(n7476), .dout(n7562));
  jnot g07307(.din(n7562), .dout(n7563));
  jor  g07308(.dina(n3849), .dinb(n1397), .dout(n7564));
  jor  g07309(.dina(n3689), .dinb(n1193), .dout(n7565));
  jor  g07310(.dina(n3852), .dinb(n1290), .dout(n7566));
  jor  g07311(.dina(n3854), .dinb(n1400), .dout(n7567));
  jand g07312(.dina(n7567), .dinb(n7566), .dout(n7568));
  jand g07313(.dina(n7568), .dinb(n7565), .dout(n7569));
  jand g07314(.dina(n7569), .dinb(n7564), .dout(n7570));
  jxor g07315(.dina(n7570), .dinb(a35 ), .dout(n7571));
  jxor g07316(.dina(n7571), .dinb(n7563), .dout(n7572));
  jxor g07317(.dina(n7572), .dinb(n7473), .dout(n7573));
  jnot g07318(.din(n7573), .dout(n7574));
  jor  g07319(.dina(n3301), .dinb(n1739), .dout(n7575));
  jor  g07320(.dina(n3136), .dinb(n1420), .dout(n7576));
  jor  g07321(.dina(n3304), .dinb(n1620), .dout(n7577));
  jor  g07322(.dina(n3306), .dinb(n1742), .dout(n7578));
  jand g07323(.dina(n7578), .dinb(n7577), .dout(n7579));
  jand g07324(.dina(n7579), .dinb(n7576), .dout(n7580));
  jand g07325(.dina(n7580), .dinb(n7575), .dout(n7581));
  jxor g07326(.dina(n7581), .dinb(a32 ), .dout(n7582));
  jxor g07327(.dina(n7582), .dinb(n7574), .dout(n7583));
  jxor g07328(.dina(n7583), .dinb(n7470), .dout(n7584));
  jnot g07329(.din(n7584), .dout(n7585));
  jor  g07330(.dina(n2784), .dinb(n2007), .dout(n7586));
  jor  g07331(.dina(n2661), .dinb(n1867), .dout(n7587));
  jor  g07332(.dina(n2787), .dinb(n1887), .dout(n7588));
  jor  g07333(.dina(n2789), .dinb(n2010), .dout(n7589));
  jand g07334(.dina(n7589), .dinb(n7588), .dout(n7590));
  jand g07335(.dina(n7590), .dinb(n7587), .dout(n7591));
  jand g07336(.dina(n7591), .dinb(n7586), .dout(n7592));
  jxor g07337(.dina(n7592), .dinb(a29 ), .dout(n7593));
  jxor g07338(.dina(n7593), .dinb(n7585), .dout(n7594));
  jxor g07339(.dina(n7594), .dinb(n7465), .dout(n7595));
  jxor g07340(.dina(n7595), .dinb(n7460), .dout(n7596));
  jxor g07341(.dina(n7596), .dinb(n7451), .dout(n7597));
  jor  g07342(.dina(n3032), .dinb(n1939), .dout(n7598));
  jor  g07343(.dina(n1827), .dinb(n2579), .dout(n7599));
  jor  g07344(.dina(n1942), .dinb(n2870), .dout(n7600));
  jor  g07345(.dina(n1944), .dinb(n3035), .dout(n7601));
  jand g07346(.dina(n7601), .dinb(n7600), .dout(n7602));
  jand g07347(.dina(n7602), .dinb(n7599), .dout(n7603));
  jand g07348(.dina(n7603), .dinb(n7598), .dout(n7604));
  jxor g07349(.dina(n7604), .dinb(a23 ), .dout(n7605));
  jxor g07350(.dina(n7605), .dinb(n7597), .dout(n7606));
  jxor g07351(.dina(n7606), .dinb(n7447), .dout(n7607));
  jor  g07352(.dina(n3400), .dinb(n1566), .dout(n7608));
  jor  g07353(.dina(n1489), .dinb(n3055), .dout(n7609));
  jor  g07354(.dina(n1569), .dinb(n3230), .dout(n7610));
  jor  g07355(.dina(n1571), .dinb(n3403), .dout(n7611));
  jand g07356(.dina(n7611), .dinb(n7610), .dout(n7612));
  jand g07357(.dina(n7612), .dinb(n7609), .dout(n7613));
  jand g07358(.dina(n7613), .dinb(n7608), .dout(n7614));
  jxor g07359(.dina(n7614), .dinb(a20 ), .dout(n7615));
  jxor g07360(.dina(n7615), .dinb(n7607), .dout(n7616));
  jxor g07361(.dina(n7616), .dinb(n7444), .dout(n7617));
  jor  g07362(.dina(n4137), .dinb(n1245), .dout(n7618));
  jor  g07363(.dina(n1165), .dinb(n3588), .dout(n7619));
  jor  g07364(.dina(n1248), .dinb(n3942), .dout(n7620));
  jor  g07365(.dina(n1250), .dinb(n4140), .dout(n7621));
  jand g07366(.dina(n7621), .dinb(n7620), .dout(n7622));
  jand g07367(.dina(n7622), .dinb(n7619), .dout(n7623));
  jand g07368(.dina(n7623), .dinb(n7618), .dout(n7624));
  jxor g07369(.dina(n7624), .dinb(a17 ), .dout(n7625));
  jxor g07370(.dina(n7625), .dinb(n7617), .dout(n7626));
  jxor g07371(.dina(n7626), .dinb(n7436), .dout(n7627));
  jnot g07372(.din(n7627), .dout(n7628));
  jor  g07373(.dina(n4554), .dinb(n974), .dout(n7629));
  jor  g07374(.dina(n908), .dinb(n4340), .dout(n7630));
  jor  g07375(.dina(n977), .dinb(n4537), .dout(n7631));
  jor  g07376(.dina(n979), .dinb(n4557), .dout(n7632));
  jand g07377(.dina(n7632), .dinb(n7631), .dout(n7633));
  jand g07378(.dina(n7633), .dinb(n7630), .dout(n7634));
  jand g07379(.dina(n7634), .dinb(n7629), .dout(n7635));
  jxor g07380(.dina(n7635), .dinb(a14 ), .dout(n7636));
  jxor g07381(.dina(n7636), .dinb(n7628), .dout(n7637));
  jxor g07382(.dina(n7637), .dinb(n7433), .dout(n7638));
  jor  g07383(.dina(n5405), .dinb(n706), .dout(n7639));
  jor  g07384(.dina(n683), .dinb(n4974), .dout(n7640));
  jor  g07385(.dina(n709), .dinb(n4994), .dout(n7641));
  jor  g07386(.dina(n711), .dinb(n5408), .dout(n7642));
  jand g07387(.dina(n7642), .dinb(n7641), .dout(n7643));
  jand g07388(.dina(n7643), .dinb(n7640), .dout(n7644));
  jand g07389(.dina(n7644), .dinb(n7639), .dout(n7645));
  jxor g07390(.dina(n7645), .dinb(a11 ), .dout(n7646));
  jxor g07391(.dina(n7646), .dinb(n7638), .dout(n7647));
  jxor g07392(.dina(n7647), .dinb(n7429), .dout(n7648));
  jnot g07393(.din(n7648), .dout(n7649));
  jor  g07394(.dina(n6103), .dinb(n528), .dout(n7650));
  jor  g07395(.dina(n490), .dinb(n5428), .dout(n7651));
  jor  g07396(.dina(n531), .dinb(n5862), .dout(n7652));
  jor  g07397(.dina(n533), .dinb(n6106), .dout(n7653));
  jand g07398(.dina(n7653), .dinb(n7652), .dout(n7654));
  jand g07399(.dina(n7654), .dinb(n7651), .dout(n7655));
  jand g07400(.dina(n7655), .dinb(n7650), .dout(n7656));
  jxor g07401(.dina(n7656), .dinb(a8 ), .dout(n7657));
  jxor g07402(.dina(n7657), .dinb(n7649), .dout(n7658));
  jxor g07403(.dina(n7658), .dinb(n7425), .dout(n7659));
  jor  g07404(.dina(n6864), .dinb(n402), .dout(n7660));
  jor  g07405(.dina(n371), .dinb(n6352), .dout(n7661));
  jor  g07406(.dina(n405), .dinb(n6372), .dout(n7662));
  jor  g07407(.dina(n332), .dinb(n6867), .dout(n7663));
  jand g07408(.dina(n7663), .dinb(n7662), .dout(n7664));
  jand g07409(.dina(n7664), .dinb(n7661), .dout(n7665));
  jand g07410(.dina(n7665), .dinb(n7660), .dout(n7666));
  jxor g07411(.dina(n7666), .dinb(a5 ), .dout(n7667));
  jxor g07412(.dina(n7667), .dinb(n7659), .dout(n7668));
  jxor g07413(.dina(n7668), .dinb(n7420), .dout(n7669));
  jxor g07414(.dina(n7669), .dinb(n7417), .dout(n7670));
  jxor g07415(.dina(n7670), .dinb(n7402), .dout(f52 ));
  jand g07416(.dina(n7669), .dinb(n7417), .dout(n7672));
  jand g07417(.dina(n7670), .dinb(n7402), .dout(n7673));
  jor  g07418(.dina(n7673), .dinb(n7672), .dout(n7674));
  jand g07419(.dina(b52 ), .dinb(b51 ), .dout(n7675));
  jand g07420(.dina(n7406), .dinb(n7405), .dout(n7676));
  jor  g07421(.dina(n7676), .dinb(n7675), .dout(n7677));
  jxor g07422(.dina(b53 ), .dinb(b52 ), .dout(n7678));
  jnot g07423(.din(n7678), .dout(n7679));
  jxor g07424(.dina(n7679), .dinb(n7677), .dout(n7680));
  jor  g07425(.dina(n7680), .dinb(n264), .dout(n7681));
  jor  g07426(.dina(n284), .dinb(n7149), .dout(n7682));
  jnot g07427(.din(b53 ), .dout(n7683));
  jor  g07428(.dina(n269), .dinb(n7683), .dout(n7684));
  jor  g07429(.dina(n271), .dinb(n7411), .dout(n7685));
  jand g07430(.dina(n7685), .dinb(n7684), .dout(n7686));
  jand g07431(.dina(n7686), .dinb(n7682), .dout(n7687));
  jand g07432(.dina(n7687), .dinb(n7681), .dout(n7688));
  jxor g07433(.dina(n7688), .dinb(n260), .dout(n7689));
  jor  g07434(.dina(n7667), .dinb(n7659), .dout(n7690));
  jnot g07435(.din(n7690), .dout(n7691));
  jand g07436(.dina(n7668), .dinb(n7420), .dout(n7692));
  jor  g07437(.dina(n7692), .dinb(n7691), .dout(n7693));
  jor  g07438(.dina(n7657), .dinb(n7649), .dout(n7694));
  jnot g07439(.din(n7694), .dout(n7695));
  jand g07440(.dina(n7658), .dinb(n7424), .dout(n7696));
  jor  g07441(.dina(n7696), .dinb(n7695), .dout(n7697));
  jnot g07442(.din(n7697), .dout(n7698));
  jnot g07443(.din(n7638), .dout(n7699));
  jor  g07444(.dina(n7646), .dinb(n7699), .dout(n7700));
  jor  g07445(.dina(n7647), .dinb(n7429), .dout(n7701));
  jand g07446(.dina(n7701), .dinb(n7700), .dout(n7702));
  jor  g07447(.dina(n7636), .dinb(n7628), .dout(n7703));
  jnot g07448(.din(n7703), .dout(n7704));
  jand g07449(.dina(n7637), .dinb(n7433), .dout(n7705));
  jor  g07450(.dina(n7705), .dinb(n7704), .dout(n7706));
  jor  g07451(.dina(n7625), .dinb(n7617), .dout(n7707));
  jnot g07452(.din(n7707), .dout(n7708));
  jand g07453(.dina(n7626), .dinb(n7436), .dout(n7709));
  jor  g07454(.dina(n7709), .dinb(n7708), .dout(n7710));
  jor  g07455(.dina(n7615), .dinb(n7607), .dout(n7711));
  jnot g07456(.din(n7616), .dout(n7712));
  jor  g07457(.dina(n7712), .dinb(n7444), .dout(n7713));
  jand g07458(.dina(n7713), .dinb(n7711), .dout(n7714));
  jnot g07459(.din(n7597), .dout(n7715));
  jor  g07460(.dina(n7605), .dinb(n7715), .dout(n7716));
  jnot g07461(.din(n7447), .dout(n7717));
  jor  g07462(.dina(n7606), .dinb(n7717), .dout(n7718));
  jand g07463(.dina(n7718), .dinb(n7716), .dout(n7719));
  jor  g07464(.dina(n3052), .dinb(n1939), .dout(n7720));
  jor  g07465(.dina(n1827), .dinb(n2870), .dout(n7721));
  jor  g07466(.dina(n1942), .dinb(n3035), .dout(n7722));
  jor  g07467(.dina(n1944), .dinb(n3055), .dout(n7723));
  jand g07468(.dina(n7723), .dinb(n7722), .dout(n7724));
  jand g07469(.dina(n7724), .dinb(n7721), .dout(n7725));
  jand g07470(.dina(n7725), .dinb(n7720), .dout(n7726));
  jxor g07471(.dina(n7726), .dinb(a23 ), .dout(n7727));
  jnot g07472(.din(n7727), .dout(n7728));
  jand g07473(.dina(n7595), .dinb(n7460), .dout(n7729));
  jand g07474(.dina(n7596), .dinb(n7451), .dout(n7730));
  jor  g07475(.dina(n7730), .dinb(n7729), .dout(n7731));
  jor  g07476(.dina(n2576), .dinb(n2319), .dout(n7732));
  jor  g07477(.dina(n2224), .dinb(n2407), .dout(n7733));
  jor  g07478(.dina(n2322), .dinb(n2559), .dout(n7734));
  jor  g07479(.dina(n2324), .dinb(n2579), .dout(n7735));
  jand g07480(.dina(n7735), .dinb(n7734), .dout(n7736));
  jand g07481(.dina(n7736), .dinb(n7733), .dout(n7737));
  jand g07482(.dina(n7737), .dinb(n7732), .dout(n7738));
  jxor g07483(.dina(n7738), .dinb(a26 ), .dout(n7739));
  jnot g07484(.din(n7739), .dout(n7740));
  jor  g07485(.dina(n7593), .dinb(n7585), .dout(n7741));
  jand g07486(.dina(n7594), .dinb(n7465), .dout(n7742));
  jnot g07487(.din(n7742), .dout(n7743));
  jand g07488(.dina(n7743), .dinb(n7741), .dout(n7744));
  jnot g07489(.din(n7744), .dout(n7745));
  jor  g07490(.dina(n2784), .dinb(n2145), .dout(n7746));
  jor  g07491(.dina(n2661), .dinb(n1887), .dout(n7747));
  jor  g07492(.dina(n2787), .dinb(n2010), .dout(n7748));
  jor  g07493(.dina(n2789), .dinb(n2148), .dout(n7749));
  jand g07494(.dina(n7749), .dinb(n7748), .dout(n7750));
  jand g07495(.dina(n7750), .dinb(n7747), .dout(n7751));
  jand g07496(.dina(n7751), .dinb(n7746), .dout(n7752));
  jxor g07497(.dina(n7752), .dinb(a29 ), .dout(n7753));
  jnot g07498(.din(n7753), .dout(n7754));
  jor  g07499(.dina(n7582), .dinb(n7574), .dout(n7755));
  jand g07500(.dina(n7583), .dinb(n7470), .dout(n7756));
  jnot g07501(.din(n7756), .dout(n7757));
  jand g07502(.dina(n7757), .dinb(n7755), .dout(n7758));
  jnot g07503(.din(n7758), .dout(n7759));
  jor  g07504(.dina(n3301), .dinb(n1864), .dout(n7760));
  jor  g07505(.dina(n3136), .dinb(n1620), .dout(n7761));
  jor  g07506(.dina(n3304), .dinb(n1742), .dout(n7762));
  jor  g07507(.dina(n3306), .dinb(n1867), .dout(n7763));
  jand g07508(.dina(n7763), .dinb(n7762), .dout(n7764));
  jand g07509(.dina(n7764), .dinb(n7761), .dout(n7765));
  jand g07510(.dina(n7765), .dinb(n7760), .dout(n7766));
  jxor g07511(.dina(n7766), .dinb(a32 ), .dout(n7767));
  jnot g07512(.din(n7767), .dout(n7768));
  jor  g07513(.dina(n7571), .dinb(n7563), .dout(n7769));
  jand g07514(.dina(n7572), .dinb(n7473), .dout(n7770));
  jnot g07515(.din(n7770), .dout(n7771));
  jand g07516(.dina(n7771), .dinb(n7769), .dout(n7772));
  jnot g07517(.din(n7772), .dout(n7773));
  jor  g07518(.dina(n3849), .dinb(n1417), .dout(n7774));
  jor  g07519(.dina(n3689), .dinb(n1290), .dout(n7775));
  jor  g07520(.dina(n3852), .dinb(n1400), .dout(n7776));
  jor  g07521(.dina(n3854), .dinb(n1420), .dout(n7777));
  jand g07522(.dina(n7777), .dinb(n7776), .dout(n7778));
  jand g07523(.dina(n7778), .dinb(n7775), .dout(n7779));
  jand g07524(.dina(n7779), .dinb(n7774), .dout(n7780));
  jxor g07525(.dina(n7780), .dinb(a35 ), .dout(n7781));
  jnot g07526(.din(n7781), .dout(n7782));
  jor  g07527(.dina(n7560), .dinb(n7552), .dout(n7783));
  jand g07528(.dina(n7561), .dinb(n7476), .dout(n7784));
  jnot g07529(.din(n7784), .dout(n7785));
  jand g07530(.dina(n7785), .dinb(n7783), .dout(n7786));
  jnot g07531(.din(n7786), .dout(n7787));
  jor  g07532(.dina(n4415), .dinb(n1190), .dout(n7788));
  jor  g07533(.dina(n4272), .dinb(n939), .dout(n7789));
  jor  g07534(.dina(n4418), .dinb(n1022), .dout(n7790));
  jor  g07535(.dina(n4420), .dinb(n1193), .dout(n7791));
  jand g07536(.dina(n7791), .dinb(n7790), .dout(n7792));
  jand g07537(.dina(n7792), .dinb(n7789), .dout(n7793));
  jand g07538(.dina(n7793), .dinb(n7788), .dout(n7794));
  jxor g07539(.dina(n7794), .dinb(a38 ), .dout(n7795));
  jnot g07540(.din(n7795), .dout(n7796));
  jand g07541(.dina(n7549), .dinb(n7488), .dout(n7797));
  jand g07542(.dina(n7550), .dinb(n7479), .dout(n7798));
  jor  g07543(.dina(n7798), .dinb(n7797), .dout(n7799));
  jor  g07544(.dina(n7547), .dinb(n7539), .dout(n7800));
  jand g07545(.dina(n7548), .dinb(n7493), .dout(n7801));
  jnot g07546(.din(n7801), .dout(n7802));
  jand g07547(.dina(n7802), .dinb(n7800), .dout(n7803));
  jnot g07548(.din(n7803), .dout(n7804));
  jor  g07549(.dina(n5739), .dinb(n644), .dout(n7805));
  jor  g07550(.dina(n5574), .dinb(n564), .dout(n7806));
  jor  g07551(.dina(n5742), .dinb(n627), .dout(n7807));
  jor  g07552(.dina(n5744), .dinb(n647), .dout(n7808));
  jand g07553(.dina(n7808), .dinb(n7807), .dout(n7809));
  jand g07554(.dina(n7809), .dinb(n7806), .dout(n7810));
  jand g07555(.dina(n7810), .dinb(n7805), .dout(n7811));
  jxor g07556(.dina(n7811), .dinb(a44 ), .dout(n7812));
  jnot g07557(.din(n7812), .dout(n7813));
  jor  g07558(.dina(n7536), .dinb(n7528), .dout(n7814));
  jand g07559(.dina(n7537), .dinb(n7498), .dout(n7815));
  jnot g07560(.din(n7815), .dout(n7816));
  jand g07561(.dina(n7816), .dinb(n7814), .dout(n7817));
  jnot g07562(.din(n7817), .dout(n7818));
  jor  g07563(.dina(n6490), .dinb(n509), .dout(n7819));
  jor  g07564(.dina(n6262), .dinb(n395), .dout(n7820));
  jor  g07565(.dina(n6493), .dinb(n431), .dout(n7821));
  jor  g07566(.dina(n6495), .dinb(n512), .dout(n7822));
  jand g07567(.dina(n7822), .dinb(n7821), .dout(n7823));
  jand g07568(.dina(n7823), .dinb(n7820), .dout(n7824));
  jand g07569(.dina(n7824), .dinb(n7819), .dout(n7825));
  jxor g07570(.dina(n7825), .dinb(a47 ), .dout(n7826));
  jnot g07571(.din(n7826), .dout(n7827));
  jand g07572(.dina(n7525), .dinb(n7511), .dout(n7828));
  jand g07573(.dina(n7526), .dinb(n7502), .dout(n7829));
  jor  g07574(.dina(n7829), .dinb(n7828), .dout(n7830));
  jor  g07575(.dina(n7266), .dinb(n354), .dout(n7831));
  jor  g07576(.dina(n7021), .dinb(n299), .dout(n7832));
  jor  g07577(.dina(n7269), .dinb(n322), .dout(n7833));
  jor  g07578(.dina(n7271), .dinb(n357), .dout(n7834));
  jand g07579(.dina(n7834), .dinb(n7833), .dout(n7835));
  jand g07580(.dina(n7835), .dinb(n7832), .dout(n7836));
  jand g07581(.dina(n7836), .dinb(n7831), .dout(n7837));
  jxor g07582(.dina(n7837), .dinb(a50 ), .dout(n7838));
  jnot g07583(.din(n7838), .dout(n7839));
  jnot g07584(.din(n7524), .dout(n7840));
  jand g07585(.dina(n7280), .dinb(a53 ), .dout(n7841));
  jand g07586(.dina(n7841), .dinb(n7840), .dout(n7842));
  jnot g07587(.din(n7842), .dout(n7843));
  jand g07588(.dina(n7843), .dinb(a53 ), .dout(n7844));
  jor  g07589(.dina(n7518), .dinb(n7514), .dout(n7845));
  jor  g07590(.dina(n7845), .dinb(n7278), .dout(n7846));
  jnot g07591(.din(n7846), .dout(n7847));
  jand g07592(.dina(n7847), .dinb(b0 ), .dout(n7848));
  jand g07593(.dina(n7515), .dinb(b2 ), .dout(n7849));
  jand g07594(.dina(n7519), .dinb(b1 ), .dout(n7850));
  jand g07595(.dina(n7521), .dinb(n375), .dout(n7851));
  jor  g07596(.dina(n7851), .dinb(n7850), .dout(n7852));
  jor  g07597(.dina(n7852), .dinb(n7849), .dout(n7853));
  jor  g07598(.dina(n7853), .dinb(n7848), .dout(n7854));
  jxor g07599(.dina(n7854), .dinb(n7844), .dout(n7855));
  jxor g07600(.dina(n7855), .dinb(n7839), .dout(n7856));
  jxor g07601(.dina(n7856), .dinb(n7830), .dout(n7857));
  jxor g07602(.dina(n7857), .dinb(n7827), .dout(n7858));
  jxor g07603(.dina(n7858), .dinb(n7818), .dout(n7859));
  jxor g07604(.dina(n7859), .dinb(n7813), .dout(n7860));
  jxor g07605(.dina(n7860), .dinb(n7804), .dout(n7861));
  jnot g07606(.din(n7861), .dout(n7862));
  jor  g07607(.dina(n5096), .dinb(n855), .dout(n7863));
  jor  g07608(.dina(n4904), .dinb(n758), .dout(n7864));
  jor  g07609(.dina(n5099), .dinb(n778), .dout(n7865));
  jor  g07610(.dina(n5101), .dinb(n858), .dout(n7866));
  jand g07611(.dina(n7866), .dinb(n7865), .dout(n7867));
  jand g07612(.dina(n7867), .dinb(n7864), .dout(n7868));
  jand g07613(.dina(n7868), .dinb(n7863), .dout(n7869));
  jxor g07614(.dina(n7869), .dinb(a41 ), .dout(n7870));
  jxor g07615(.dina(n7870), .dinb(n7862), .dout(n7871));
  jxor g07616(.dina(n7871), .dinb(n7799), .dout(n7872));
  jxor g07617(.dina(n7872), .dinb(n7796), .dout(n7873));
  jxor g07618(.dina(n7873), .dinb(n7787), .dout(n7874));
  jxor g07619(.dina(n7874), .dinb(n7782), .dout(n7875));
  jxor g07620(.dina(n7875), .dinb(n7773), .dout(n7876));
  jxor g07621(.dina(n7876), .dinb(n7768), .dout(n7877));
  jxor g07622(.dina(n7877), .dinb(n7759), .dout(n7878));
  jxor g07623(.dina(n7878), .dinb(n7754), .dout(n7879));
  jxor g07624(.dina(n7879), .dinb(n7745), .dout(n7880));
  jxor g07625(.dina(n7880), .dinb(n7740), .dout(n7881));
  jxor g07626(.dina(n7881), .dinb(n7731), .dout(n7882));
  jxor g07627(.dina(n7882), .dinb(n7728), .dout(n7883));
  jxor g07628(.dina(n7883), .dinb(n7719), .dout(n7884));
  jor  g07629(.dina(n3585), .dinb(n1566), .dout(n7885));
  jor  g07630(.dina(n1489), .dinb(n3230), .dout(n7886));
  jor  g07631(.dina(n1569), .dinb(n3403), .dout(n7887));
  jor  g07632(.dina(n1571), .dinb(n3588), .dout(n7888));
  jand g07633(.dina(n7888), .dinb(n7887), .dout(n7889));
  jand g07634(.dina(n7889), .dinb(n7886), .dout(n7890));
  jand g07635(.dina(n7890), .dinb(n7885), .dout(n7891));
  jxor g07636(.dina(n7891), .dinb(a20 ), .dout(n7892));
  jxor g07637(.dina(n7892), .dinb(n7884), .dout(n7893));
  jxor g07638(.dina(n7893), .dinb(n7714), .dout(n7894));
  jor  g07639(.dina(n4337), .dinb(n1245), .dout(n7895));
  jor  g07640(.dina(n1165), .dinb(n3942), .dout(n7896));
  jor  g07641(.dina(n1248), .dinb(n4140), .dout(n7897));
  jor  g07642(.dina(n1250), .dinb(n4340), .dout(n7898));
  jand g07643(.dina(n7898), .dinb(n7897), .dout(n7899));
  jand g07644(.dina(n7899), .dinb(n7896), .dout(n7900));
  jand g07645(.dina(n7900), .dinb(n7895), .dout(n7901));
  jxor g07646(.dina(n7901), .dinb(a17 ), .dout(n7902));
  jxor g07647(.dina(n7902), .dinb(n7894), .dout(n7903));
  jxor g07648(.dina(n7903), .dinb(n7710), .dout(n7904));
  jnot g07649(.din(n7904), .dout(n7905));
  jor  g07650(.dina(n4971), .dinb(n974), .dout(n7906));
  jor  g07651(.dina(n908), .dinb(n4537), .dout(n7907));
  jor  g07652(.dina(n977), .dinb(n4557), .dout(n7908));
  jor  g07653(.dina(n979), .dinb(n4974), .dout(n7909));
  jand g07654(.dina(n7909), .dinb(n7908), .dout(n7910));
  jand g07655(.dina(n7910), .dinb(n7907), .dout(n7911));
  jand g07656(.dina(n7911), .dinb(n7906), .dout(n7912));
  jxor g07657(.dina(n7912), .dinb(a14 ), .dout(n7913));
  jxor g07658(.dina(n7913), .dinb(n7905), .dout(n7914));
  jxor g07659(.dina(n7914), .dinb(n7706), .dout(n7915));
  jor  g07660(.dina(n5425), .dinb(n706), .dout(n7916));
  jor  g07661(.dina(n683), .dinb(n4994), .dout(n7917));
  jor  g07662(.dina(n709), .dinb(n5408), .dout(n7918));
  jor  g07663(.dina(n711), .dinb(n5428), .dout(n7919));
  jand g07664(.dina(n7919), .dinb(n7918), .dout(n7920));
  jand g07665(.dina(n7920), .dinb(n7917), .dout(n7921));
  jand g07666(.dina(n7921), .dinb(n7916), .dout(n7922));
  jxor g07667(.dina(n7922), .dinb(a11 ), .dout(n7923));
  jxor g07668(.dina(n7923), .dinb(n7915), .dout(n7924));
  jxor g07669(.dina(n7924), .dinb(n7702), .dout(n7925));
  jnot g07670(.din(n7925), .dout(n7926));
  jor  g07671(.dina(n6349), .dinb(n528), .dout(n7927));
  jor  g07672(.dina(n490), .dinb(n5862), .dout(n7928));
  jor  g07673(.dina(n531), .dinb(n6106), .dout(n7929));
  jor  g07674(.dina(n533), .dinb(n6352), .dout(n7930));
  jand g07675(.dina(n7930), .dinb(n7929), .dout(n7931));
  jand g07676(.dina(n7931), .dinb(n7928), .dout(n7932));
  jand g07677(.dina(n7932), .dinb(n7927), .dout(n7933));
  jxor g07678(.dina(n7933), .dinb(a8 ), .dout(n7934));
  jxor g07679(.dina(n7934), .dinb(n7926), .dout(n7935));
  jxor g07680(.dina(n7935), .dinb(n7698), .dout(n7936));
  jor  g07681(.dina(n7126), .dinb(n402), .dout(n7937));
  jor  g07682(.dina(n371), .dinb(n6372), .dout(n7938));
  jor  g07683(.dina(n405), .dinb(n6867), .dout(n7939));
  jor  g07684(.dina(n332), .dinb(n7129), .dout(n7940));
  jand g07685(.dina(n7940), .dinb(n7939), .dout(n7941));
  jand g07686(.dina(n7941), .dinb(n7938), .dout(n7942));
  jand g07687(.dina(n7942), .dinb(n7937), .dout(n7943));
  jxor g07688(.dina(n7943), .dinb(a5 ), .dout(n7944));
  jxor g07689(.dina(n7944), .dinb(n7936), .dout(n7945));
  jxor g07690(.dina(n7945), .dinb(n7693), .dout(n7946));
  jxor g07691(.dina(n7946), .dinb(n7689), .dout(n7947));
  jxor g07692(.dina(n7947), .dinb(n7674), .dout(f53 ));
  jand g07693(.dina(n7946), .dinb(n7689), .dout(n7949));
  jand g07694(.dina(n7947), .dinb(n7674), .dout(n7950));
  jor  g07695(.dina(n7950), .dinb(n7949), .dout(n7951));
  jand g07696(.dina(b53 ), .dinb(b52 ), .dout(n7952));
  jand g07697(.dina(n7678), .dinb(n7677), .dout(n7953));
  jor  g07698(.dina(n7953), .dinb(n7952), .dout(n7954));
  jxor g07699(.dina(b54 ), .dinb(b53 ), .dout(n7955));
  jnot g07700(.din(n7955), .dout(n7956));
  jxor g07701(.dina(n7956), .dinb(n7954), .dout(n7957));
  jor  g07702(.dina(n7957), .dinb(n264), .dout(n7958));
  jor  g07703(.dina(n284), .dinb(n7411), .dout(n7959));
  jnot g07704(.din(b54 ), .dout(n7960));
  jor  g07705(.dina(n269), .dinb(n7960), .dout(n7961));
  jor  g07706(.dina(n271), .dinb(n7683), .dout(n7962));
  jand g07707(.dina(n7962), .dinb(n7961), .dout(n7963));
  jand g07708(.dina(n7963), .dinb(n7959), .dout(n7964));
  jand g07709(.dina(n7964), .dinb(n7958), .dout(n7965));
  jxor g07710(.dina(n7965), .dinb(n260), .dout(n7966));
  jor  g07711(.dina(n7944), .dinb(n7936), .dout(n7967));
  jnot g07712(.din(n7967), .dout(n7968));
  jand g07713(.dina(n7945), .dinb(n7693), .dout(n7969));
  jor  g07714(.dina(n7969), .dinb(n7968), .dout(n7970));
  jor  g07715(.dina(n7934), .dinb(n7926), .dout(n7971));
  jnot g07716(.din(n7971), .dout(n7972));
  jand g07717(.dina(n7935), .dinb(n7697), .dout(n7973));
  jor  g07718(.dina(n7973), .dinb(n7972), .dout(n7974));
  jor  g07719(.dina(n6369), .dinb(n528), .dout(n7975));
  jor  g07720(.dina(n490), .dinb(n6106), .dout(n7976));
  jor  g07721(.dina(n531), .dinb(n6352), .dout(n7977));
  jor  g07722(.dina(n533), .dinb(n6372), .dout(n7978));
  jand g07723(.dina(n7978), .dinb(n7977), .dout(n7979));
  jand g07724(.dina(n7979), .dinb(n7976), .dout(n7980));
  jand g07725(.dina(n7980), .dinb(n7975), .dout(n7981));
  jxor g07726(.dina(n7981), .dinb(a8 ), .dout(n7982));
  jnot g07727(.din(n7915), .dout(n7983));
  jor  g07728(.dina(n7923), .dinb(n7983), .dout(n7984));
  jor  g07729(.dina(n7924), .dinb(n7702), .dout(n7985));
  jand g07730(.dina(n7985), .dinb(n7984), .dout(n7986));
  jor  g07731(.dina(n5859), .dinb(n706), .dout(n7987));
  jor  g07732(.dina(n683), .dinb(n5408), .dout(n7988));
  jor  g07733(.dina(n709), .dinb(n5428), .dout(n7989));
  jor  g07734(.dina(n711), .dinb(n5862), .dout(n7990));
  jand g07735(.dina(n7990), .dinb(n7989), .dout(n7991));
  jand g07736(.dina(n7991), .dinb(n7988), .dout(n7992));
  jand g07737(.dina(n7992), .dinb(n7987), .dout(n7993));
  jxor g07738(.dina(n7993), .dinb(a11 ), .dout(n7994));
  jor  g07739(.dina(n7913), .dinb(n7905), .dout(n7995));
  jnot g07740(.din(n7995), .dout(n7996));
  jand g07741(.dina(n7914), .dinb(n7706), .dout(n7997));
  jor  g07742(.dina(n7997), .dinb(n7996), .dout(n7998));
  jor  g07743(.dina(n7902), .dinb(n7894), .dout(n7999));
  jnot g07744(.din(n7999), .dout(n8000));
  jand g07745(.dina(n7903), .dinb(n7710), .dout(n8001));
  jor  g07746(.dina(n8001), .dinb(n8000), .dout(n8002));
  jor  g07747(.dina(n7892), .dinb(n7884), .dout(n8003));
  jnot g07748(.din(n7716), .dout(n8004));
  jnot g07749(.din(n7606), .dout(n8005));
  jand g07750(.dina(n8005), .dinb(n7447), .dout(n8006));
  jor  g07751(.dina(n8006), .dinb(n8004), .dout(n8007));
  jxor g07752(.dina(n7883), .dinb(n8007), .dout(n8008));
  jxor g07753(.dina(n7892), .dinb(n8008), .dout(n8009));
  jor  g07754(.dina(n8009), .dinb(n7714), .dout(n8010));
  jand g07755(.dina(n8010), .dinb(n8003), .dout(n8011));
  jor  g07756(.dina(n3939), .dinb(n1566), .dout(n8012));
  jor  g07757(.dina(n1489), .dinb(n3403), .dout(n8013));
  jor  g07758(.dina(n1569), .dinb(n3588), .dout(n8014));
  jor  g07759(.dina(n1571), .dinb(n3942), .dout(n8015));
  jand g07760(.dina(n8015), .dinb(n8014), .dout(n8016));
  jand g07761(.dina(n8016), .dinb(n8013), .dout(n8017));
  jand g07762(.dina(n8017), .dinb(n8012), .dout(n8018));
  jxor g07763(.dina(n8018), .dinb(a20 ), .dout(n8019));
  jnot g07764(.din(n8019), .dout(n8020));
  jand g07765(.dina(n7882), .dinb(n7728), .dout(n8021));
  jand g07766(.dina(n7883), .dinb(n8007), .dout(n8022));
  jor  g07767(.dina(n8022), .dinb(n8021), .dout(n8023));
  jand g07768(.dina(n7880), .dinb(n7740), .dout(n8024));
  jand g07769(.dina(n7881), .dinb(n7731), .dout(n8025));
  jor  g07770(.dina(n8025), .dinb(n8024), .dout(n8026));
  jor  g07771(.dina(n2867), .dinb(n2319), .dout(n8027));
  jor  g07772(.dina(n2224), .dinb(n2559), .dout(n8028));
  jor  g07773(.dina(n2322), .dinb(n2579), .dout(n8029));
  jor  g07774(.dina(n2324), .dinb(n2870), .dout(n8030));
  jand g07775(.dina(n8030), .dinb(n8029), .dout(n8031));
  jand g07776(.dina(n8031), .dinb(n8028), .dout(n8032));
  jand g07777(.dina(n8032), .dinb(n8027), .dout(n8033));
  jxor g07778(.dina(n8033), .dinb(a26 ), .dout(n8034));
  jnot g07779(.din(n8034), .dout(n8035));
  jand g07780(.dina(n7878), .dinb(n7754), .dout(n8036));
  jand g07781(.dina(n7879), .dinb(n7745), .dout(n8037));
  jor  g07782(.dina(n8037), .dinb(n8036), .dout(n8038));
  jor  g07783(.dina(n2784), .dinb(n2404), .dout(n8039));
  jor  g07784(.dina(n2661), .dinb(n2010), .dout(n8040));
  jor  g07785(.dina(n2787), .dinb(n2148), .dout(n8041));
  jor  g07786(.dina(n2789), .dinb(n2407), .dout(n8042));
  jand g07787(.dina(n8042), .dinb(n8041), .dout(n8043));
  jand g07788(.dina(n8043), .dinb(n8040), .dout(n8044));
  jand g07789(.dina(n8044), .dinb(n8039), .dout(n8045));
  jxor g07790(.dina(n8045), .dinb(a29 ), .dout(n8046));
  jnot g07791(.din(n8046), .dout(n8047));
  jand g07792(.dina(n7876), .dinb(n7768), .dout(n8048));
  jand g07793(.dina(n7877), .dinb(n7759), .dout(n8049));
  jor  g07794(.dina(n8049), .dinb(n8048), .dout(n8050));
  jor  g07795(.dina(n3301), .dinb(n1884), .dout(n8051));
  jor  g07796(.dina(n3136), .dinb(n1742), .dout(n8052));
  jor  g07797(.dina(n3304), .dinb(n1867), .dout(n8053));
  jor  g07798(.dina(n3306), .dinb(n1887), .dout(n8054));
  jand g07799(.dina(n8054), .dinb(n8053), .dout(n8055));
  jand g07800(.dina(n8055), .dinb(n8052), .dout(n8056));
  jand g07801(.dina(n8056), .dinb(n8051), .dout(n8057));
  jxor g07802(.dina(n8057), .dinb(a32 ), .dout(n8058));
  jnot g07803(.din(n8058), .dout(n8059));
  jand g07804(.dina(n7874), .dinb(n7782), .dout(n8060));
  jand g07805(.dina(n7875), .dinb(n7773), .dout(n8061));
  jor  g07806(.dina(n8061), .dinb(n8060), .dout(n8062));
  jor  g07807(.dina(n3849), .dinb(n1617), .dout(n8063));
  jor  g07808(.dina(n3689), .dinb(n1400), .dout(n8064));
  jor  g07809(.dina(n3852), .dinb(n1420), .dout(n8065));
  jor  g07810(.dina(n3854), .dinb(n1620), .dout(n8066));
  jand g07811(.dina(n8066), .dinb(n8065), .dout(n8067));
  jand g07812(.dina(n8067), .dinb(n8064), .dout(n8068));
  jand g07813(.dina(n8068), .dinb(n8063), .dout(n8069));
  jxor g07814(.dina(n8069), .dinb(a35 ), .dout(n8070));
  jnot g07815(.din(n8070), .dout(n8071));
  jand g07816(.dina(n7872), .dinb(n7796), .dout(n8072));
  jand g07817(.dina(n7873), .dinb(n7787), .dout(n8073));
  jor  g07818(.dina(n8073), .dinb(n8072), .dout(n8074));
  jor  g07819(.dina(n4415), .dinb(n1287), .dout(n8075));
  jor  g07820(.dina(n4272), .dinb(n1022), .dout(n8076));
  jor  g07821(.dina(n4418), .dinb(n1193), .dout(n8077));
  jor  g07822(.dina(n4420), .dinb(n1290), .dout(n8078));
  jand g07823(.dina(n8078), .dinb(n8077), .dout(n8079));
  jand g07824(.dina(n8079), .dinb(n8076), .dout(n8080));
  jand g07825(.dina(n8080), .dinb(n8075), .dout(n8081));
  jxor g07826(.dina(n8081), .dinb(a38 ), .dout(n8082));
  jnot g07827(.din(n8082), .dout(n8083));
  jor  g07828(.dina(n7870), .dinb(n7862), .dout(n8084));
  jand g07829(.dina(n7871), .dinb(n7799), .dout(n8085));
  jnot g07830(.din(n8085), .dout(n8086));
  jand g07831(.dina(n8086), .dinb(n8084), .dout(n8087));
  jnot g07832(.din(n8087), .dout(n8088));
  jor  g07833(.dina(n5096), .dinb(n936), .dout(n8089));
  jor  g07834(.dina(n4904), .dinb(n778), .dout(n8090));
  jor  g07835(.dina(n5099), .dinb(n858), .dout(n8091));
  jor  g07836(.dina(n5101), .dinb(n939), .dout(n8092));
  jand g07837(.dina(n8092), .dinb(n8091), .dout(n8093));
  jand g07838(.dina(n8093), .dinb(n8090), .dout(n8094));
  jand g07839(.dina(n8094), .dinb(n8089), .dout(n8095));
  jxor g07840(.dina(n8095), .dinb(a41 ), .dout(n8096));
  jnot g07841(.din(n8096), .dout(n8097));
  jand g07842(.dina(n7859), .dinb(n7813), .dout(n8098));
  jand g07843(.dina(n7860), .dinb(n7804), .dout(n8099));
  jor  g07844(.dina(n8099), .dinb(n8098), .dout(n8100));
  jor  g07845(.dina(n5739), .dinb(n755), .dout(n8101));
  jor  g07846(.dina(n5574), .dinb(n627), .dout(n8102));
  jor  g07847(.dina(n5742), .dinb(n647), .dout(n8103));
  jor  g07848(.dina(n5744), .dinb(n758), .dout(n8104));
  jand g07849(.dina(n8104), .dinb(n8103), .dout(n8105));
  jand g07850(.dina(n8105), .dinb(n8102), .dout(n8106));
  jand g07851(.dina(n8106), .dinb(n8101), .dout(n8107));
  jxor g07852(.dina(n8107), .dinb(a44 ), .dout(n8108));
  jnot g07853(.din(n8108), .dout(n8109));
  jand g07854(.dina(n7857), .dinb(n7827), .dout(n8110));
  jand g07855(.dina(n7858), .dinb(n7818), .dout(n8111));
  jor  g07856(.dina(n8111), .dinb(n8110), .dout(n8112));
  jor  g07857(.dina(n6490), .dinb(n561), .dout(n8113));
  jor  g07858(.dina(n6262), .dinb(n431), .dout(n8114));
  jor  g07859(.dina(n6493), .dinb(n512), .dout(n8115));
  jor  g07860(.dina(n6495), .dinb(n564), .dout(n8116));
  jand g07861(.dina(n8116), .dinb(n8115), .dout(n8117));
  jand g07862(.dina(n8117), .dinb(n8114), .dout(n8118));
  jand g07863(.dina(n8118), .dinb(n8113), .dout(n8119));
  jxor g07864(.dina(n8119), .dinb(a47 ), .dout(n8120));
  jnot g07865(.din(n8120), .dout(n8121));
  jand g07866(.dina(n7855), .dinb(n7839), .dout(n8122));
  jand g07867(.dina(n7856), .dinb(n7830), .dout(n8123));
  jor  g07868(.dina(n8123), .dinb(n8122), .dout(n8124));
  jnot g07869(.din(n7521), .dout(n8125));
  jor  g07870(.dina(n8125), .dinb(n296), .dout(n8126));
  jor  g07871(.dina(n7846), .dinb(n267), .dout(n8127));
  jnot g07872(.din(n7519), .dout(n8128));
  jor  g07873(.dina(n8128), .dinb(n279), .dout(n8129));
  jnot g07874(.din(n7515), .dout(n8130));
  jor  g07875(.dina(n8130), .dinb(n299), .dout(n8131));
  jand g07876(.dina(n8131), .dinb(n8129), .dout(n8132));
  jand g07877(.dina(n8132), .dinb(n8127), .dout(n8133));
  jand g07878(.dina(n8133), .dinb(n8126), .dout(n8134));
  jxor g07879(.dina(n8134), .dinb(a53 ), .dout(n8135));
  jnot g07880(.din(n8135), .dout(n8136));
  jxor g07881(.dina(a54 ), .dinb(a53 ), .dout(n8137));
  jand g07882(.dina(n8137), .dinb(b0 ), .dout(n8138));
  jnot g07883(.din(n8138), .dout(n8139));
  jor  g07884(.dina(n7854), .dinb(n7843), .dout(n8140));
  jxor g07885(.dina(n8140), .dinb(n8139), .dout(n8141));
  jxor g07886(.dina(n8141), .dinb(n8136), .dout(n8142));
  jnot g07887(.din(n8142), .dout(n8143));
  jor  g07888(.dina(n7266), .dinb(n392), .dout(n8144));
  jor  g07889(.dina(n7021), .dinb(n322), .dout(n8145));
  jor  g07890(.dina(n7269), .dinb(n357), .dout(n8146));
  jor  g07891(.dina(n7271), .dinb(n395), .dout(n8147));
  jand g07892(.dina(n8147), .dinb(n8146), .dout(n8148));
  jand g07893(.dina(n8148), .dinb(n8145), .dout(n8149));
  jand g07894(.dina(n8149), .dinb(n8144), .dout(n8150));
  jxor g07895(.dina(n8150), .dinb(a50 ), .dout(n8151));
  jxor g07896(.dina(n8151), .dinb(n8143), .dout(n8152));
  jxor g07897(.dina(n8152), .dinb(n8124), .dout(n8153));
  jxor g07898(.dina(n8153), .dinb(n8121), .dout(n8154));
  jxor g07899(.dina(n8154), .dinb(n8112), .dout(n8155));
  jxor g07900(.dina(n8155), .dinb(n8109), .dout(n8156));
  jxor g07901(.dina(n8156), .dinb(n8100), .dout(n8157));
  jxor g07902(.dina(n8157), .dinb(n8097), .dout(n8158));
  jxor g07903(.dina(n8158), .dinb(n8088), .dout(n8159));
  jxor g07904(.dina(n8159), .dinb(n8083), .dout(n8160));
  jxor g07905(.dina(n8160), .dinb(n8074), .dout(n8161));
  jxor g07906(.dina(n8161), .dinb(n8071), .dout(n8162));
  jxor g07907(.dina(n8162), .dinb(n8062), .dout(n8163));
  jxor g07908(.dina(n8163), .dinb(n8059), .dout(n8164));
  jxor g07909(.dina(n8164), .dinb(n8050), .dout(n8165));
  jxor g07910(.dina(n8165), .dinb(n8047), .dout(n8166));
  jxor g07911(.dina(n8166), .dinb(n8038), .dout(n8167));
  jxor g07912(.dina(n8167), .dinb(n8035), .dout(n8168));
  jxor g07913(.dina(n8168), .dinb(n8026), .dout(n8169));
  jor  g07914(.dina(n3227), .dinb(n1939), .dout(n8170));
  jor  g07915(.dina(n1827), .dinb(n3035), .dout(n8171));
  jor  g07916(.dina(n1942), .dinb(n3055), .dout(n8172));
  jor  g07917(.dina(n1944), .dinb(n3230), .dout(n8173));
  jand g07918(.dina(n8173), .dinb(n8172), .dout(n8174));
  jand g07919(.dina(n8174), .dinb(n8171), .dout(n8175));
  jand g07920(.dina(n8175), .dinb(n8170), .dout(n8176));
  jxor g07921(.dina(n8176), .dinb(a23 ), .dout(n8177));
  jxor g07922(.dina(n8177), .dinb(n8169), .dout(n8178));
  jnot g07923(.din(n8178), .dout(n8179));
  jxor g07924(.dina(n8179), .dinb(n8023), .dout(n8180));
  jxor g07925(.dina(n8180), .dinb(n8020), .dout(n8181));
  jxor g07926(.dina(n8181), .dinb(n8011), .dout(n8182));
  jor  g07927(.dina(n4534), .dinb(n1245), .dout(n8183));
  jor  g07928(.dina(n1165), .dinb(n4140), .dout(n8184));
  jor  g07929(.dina(n1248), .dinb(n4340), .dout(n8185));
  jor  g07930(.dina(n1250), .dinb(n4537), .dout(n8186));
  jand g07931(.dina(n8186), .dinb(n8185), .dout(n8187));
  jand g07932(.dina(n8187), .dinb(n8184), .dout(n8188));
  jand g07933(.dina(n8188), .dinb(n8183), .dout(n8189));
  jxor g07934(.dina(n8189), .dinb(a17 ), .dout(n8190));
  jxor g07935(.dina(n8190), .dinb(n8182), .dout(n8191));
  jxor g07936(.dina(n8191), .dinb(n8002), .dout(n8192));
  jnot g07937(.din(n8192), .dout(n8193));
  jor  g07938(.dina(n4991), .dinb(n974), .dout(n8194));
  jor  g07939(.dina(n908), .dinb(n4557), .dout(n8195));
  jor  g07940(.dina(n977), .dinb(n4974), .dout(n8196));
  jor  g07941(.dina(n979), .dinb(n4994), .dout(n8197));
  jand g07942(.dina(n8197), .dinb(n8196), .dout(n8198));
  jand g07943(.dina(n8198), .dinb(n8195), .dout(n8199));
  jand g07944(.dina(n8199), .dinb(n8194), .dout(n8200));
  jxor g07945(.dina(n8200), .dinb(a14 ), .dout(n8201));
  jxor g07946(.dina(n8201), .dinb(n8193), .dout(n8202));
  jxor g07947(.dina(n8202), .dinb(n7998), .dout(n8203));
  jxor g07948(.dina(n8203), .dinb(n7994), .dout(n8204));
  jxor g07949(.dina(n8204), .dinb(n7986), .dout(n8205));
  jxor g07950(.dina(n8205), .dinb(n7982), .dout(n8206));
  jxor g07951(.dina(n8206), .dinb(n7974), .dout(n8207));
  jor  g07952(.dina(n7146), .dinb(n402), .dout(n8208));
  jor  g07953(.dina(n371), .dinb(n6867), .dout(n8209));
  jor  g07954(.dina(n405), .dinb(n7129), .dout(n8210));
  jor  g07955(.dina(n332), .dinb(n7149), .dout(n8211));
  jand g07956(.dina(n8211), .dinb(n8210), .dout(n8212));
  jand g07957(.dina(n8212), .dinb(n8209), .dout(n8213));
  jand g07958(.dina(n8213), .dinb(n8208), .dout(n8214));
  jxor g07959(.dina(n8214), .dinb(a5 ), .dout(n8215));
  jxor g07960(.dina(n8215), .dinb(n8207), .dout(n8216));
  jxor g07961(.dina(n8216), .dinb(n7970), .dout(n8217));
  jxor g07962(.dina(n8217), .dinb(n7966), .dout(n8218));
  jxor g07963(.dina(n8218), .dinb(n7951), .dout(f54 ));
  jand g07964(.dina(n8217), .dinb(n7966), .dout(n8220));
  jand g07965(.dina(n8218), .dinb(n7951), .dout(n8221));
  jor  g07966(.dina(n8221), .dinb(n8220), .dout(n8222));
  jand g07967(.dina(b54 ), .dinb(b53 ), .dout(n8223));
  jand g07968(.dina(n7955), .dinb(n7954), .dout(n8224));
  jor  g07969(.dina(n8224), .dinb(n8223), .dout(n8225));
  jxor g07970(.dina(b55 ), .dinb(b54 ), .dout(n8226));
  jnot g07971(.din(n8226), .dout(n8227));
  jxor g07972(.dina(n8227), .dinb(n8225), .dout(n8228));
  jor  g07973(.dina(n8228), .dinb(n264), .dout(n8229));
  jor  g07974(.dina(n284), .dinb(n7683), .dout(n8230));
  jnot g07975(.din(b55 ), .dout(n8231));
  jor  g07976(.dina(n269), .dinb(n8231), .dout(n8232));
  jor  g07977(.dina(n271), .dinb(n7960), .dout(n8233));
  jand g07978(.dina(n8233), .dinb(n8232), .dout(n8234));
  jand g07979(.dina(n8234), .dinb(n8230), .dout(n8235));
  jand g07980(.dina(n8235), .dinb(n8229), .dout(n8236));
  jxor g07981(.dina(n8236), .dinb(n260), .dout(n8237));
  jor  g07982(.dina(n8215), .dinb(n8207), .dout(n8238));
  jnot g07983(.din(n8238), .dout(n8239));
  jand g07984(.dina(n8216), .dinb(n7970), .dout(n8240));
  jor  g07985(.dina(n8240), .dinb(n8239), .dout(n8241));
  jnot g07986(.din(n7982), .dout(n8242));
  jand g07987(.dina(n8205), .dinb(n8242), .dout(n8243));
  jxor g07988(.dina(n8205), .dinb(n8242), .dout(n8244));
  jand g07989(.dina(n8244), .dinb(n7974), .dout(n8245));
  jor  g07990(.dina(n8245), .dinb(n8243), .dout(n8246));
  jor  g07991(.dina(n6864), .dinb(n528), .dout(n8247));
  jor  g07992(.dina(n490), .dinb(n6352), .dout(n8248));
  jor  g07993(.dina(n531), .dinb(n6372), .dout(n8249));
  jor  g07994(.dina(n533), .dinb(n6867), .dout(n8250));
  jand g07995(.dina(n8250), .dinb(n8249), .dout(n8251));
  jand g07996(.dina(n8251), .dinb(n8248), .dout(n8252));
  jand g07997(.dina(n8252), .dinb(n8247), .dout(n8253));
  jxor g07998(.dina(n8253), .dinb(a8 ), .dout(n8254));
  jnot g07999(.din(n8254), .dout(n8255));
  jnot g08000(.din(n7994), .dout(n8256));
  jand g08001(.dina(n8203), .dinb(n8256), .dout(n8257));
  jnot g08002(.din(n8257), .dout(n8258));
  jor  g08003(.dina(n8204), .dinb(n7986), .dout(n8259));
  jand g08004(.dina(n8259), .dinb(n8258), .dout(n8260));
  jor  g08005(.dina(n6103), .dinb(n706), .dout(n8261));
  jor  g08006(.dina(n683), .dinb(n5428), .dout(n8262));
  jor  g08007(.dina(n709), .dinb(n5862), .dout(n8263));
  jor  g08008(.dina(n711), .dinb(n6106), .dout(n8264));
  jand g08009(.dina(n8264), .dinb(n8263), .dout(n8265));
  jand g08010(.dina(n8265), .dinb(n8262), .dout(n8266));
  jand g08011(.dina(n8266), .dinb(n8261), .dout(n8267));
  jxor g08012(.dina(n8267), .dinb(a11 ), .dout(n8268));
  jor  g08013(.dina(n8201), .dinb(n8193), .dout(n8269));
  jnot g08014(.din(n8269), .dout(n8270));
  jand g08015(.dina(n8202), .dinb(n7998), .dout(n8271));
  jor  g08016(.dina(n8271), .dinb(n8270), .dout(n8272));
  jor  g08017(.dina(n8190), .dinb(n8182), .dout(n8273));
  jnot g08018(.din(n8273), .dout(n8274));
  jand g08019(.dina(n8191), .dinb(n8002), .dout(n8275));
  jor  g08020(.dina(n8275), .dinb(n8274), .dout(n8276));
  jand g08021(.dina(n8180), .dinb(n8020), .dout(n8277));
  jnot g08022(.din(n8277), .dout(n8278));
  jxor g08023(.dina(n8180), .dinb(n8019), .dout(n8279));
  jor  g08024(.dina(n8279), .dinb(n8011), .dout(n8280));
  jand g08025(.dina(n8280), .dinb(n8278), .dout(n8281));
  jnot g08026(.din(n8169), .dout(n8282));
  jor  g08027(.dina(n8177), .dinb(n8282), .dout(n8283));
  jnot g08028(.din(n8021), .dout(n8284));
  jnot g08029(.din(n7883), .dout(n8285));
  jor  g08030(.dina(n8285), .dinb(n7719), .dout(n8286));
  jand g08031(.dina(n8286), .dinb(n8284), .dout(n8287));
  jor  g08032(.dina(n8178), .dinb(n8287), .dout(n8288));
  jand g08033(.dina(n8288), .dinb(n8283), .dout(n8289));
  jand g08034(.dina(n8167), .dinb(n8035), .dout(n8290));
  jand g08035(.dina(n8168), .dinb(n8026), .dout(n8291));
  jor  g08036(.dina(n8291), .dinb(n8290), .dout(n8292));
  jand g08037(.dina(n8165), .dinb(n8047), .dout(n8293));
  jand g08038(.dina(n8166), .dinb(n8038), .dout(n8294));
  jor  g08039(.dina(n8294), .dinb(n8293), .dout(n8295));
  jand g08040(.dina(n8163), .dinb(n8059), .dout(n8296));
  jand g08041(.dina(n8164), .dinb(n8050), .dout(n8297));
  jor  g08042(.dina(n8297), .dinb(n8296), .dout(n8298));
  jand g08043(.dina(n8161), .dinb(n8071), .dout(n8299));
  jand g08044(.dina(n8162), .dinb(n8062), .dout(n8300));
  jor  g08045(.dina(n8300), .dinb(n8299), .dout(n8301));
  jand g08046(.dina(n8159), .dinb(n8083), .dout(n8302));
  jand g08047(.dina(n8160), .dinb(n8074), .dout(n8303));
  jor  g08048(.dina(n8303), .dinb(n8302), .dout(n8304));
  jand g08049(.dina(n8157), .dinb(n8097), .dout(n8305));
  jand g08050(.dina(n8158), .dinb(n8088), .dout(n8306));
  jor  g08051(.dina(n8306), .dinb(n8305), .dout(n8307));
  jand g08052(.dina(n8155), .dinb(n8109), .dout(n8308));
  jand g08053(.dina(n8156), .dinb(n8100), .dout(n8309));
  jor  g08054(.dina(n8309), .dinb(n8308), .dout(n8310));
  jor  g08055(.dina(n5739), .dinb(n775), .dout(n8311));
  jor  g08056(.dina(n5574), .dinb(n647), .dout(n8312));
  jor  g08057(.dina(n5742), .dinb(n758), .dout(n8313));
  jor  g08058(.dina(n5744), .dinb(n778), .dout(n8314));
  jand g08059(.dina(n8314), .dinb(n8313), .dout(n8315));
  jand g08060(.dina(n8315), .dinb(n8312), .dout(n8316));
  jand g08061(.dina(n8316), .dinb(n8311), .dout(n8317));
  jxor g08062(.dina(n8317), .dinb(a44 ), .dout(n8318));
  jnot g08063(.din(n8318), .dout(n8319));
  jand g08064(.dina(n8153), .dinb(n8121), .dout(n8320));
  jand g08065(.dina(n8154), .dinb(n8112), .dout(n8321));
  jor  g08066(.dina(n8321), .dinb(n8320), .dout(n8322));
  jor  g08067(.dina(n6490), .dinb(n624), .dout(n8323));
  jor  g08068(.dina(n6262), .dinb(n512), .dout(n8324));
  jor  g08069(.dina(n6493), .dinb(n564), .dout(n8325));
  jor  g08070(.dina(n6495), .dinb(n627), .dout(n8326));
  jand g08071(.dina(n8326), .dinb(n8325), .dout(n8327));
  jand g08072(.dina(n8327), .dinb(n8324), .dout(n8328));
  jand g08073(.dina(n8328), .dinb(n8323), .dout(n8329));
  jxor g08074(.dina(n8329), .dinb(a47 ), .dout(n8330));
  jnot g08075(.din(n8330), .dout(n8331));
  jor  g08076(.dina(n8151), .dinb(n8143), .dout(n8332));
  jand g08077(.dina(n8152), .dinb(n8124), .dout(n8333));
  jnot g08078(.din(n8333), .dout(n8334));
  jand g08079(.dina(n8334), .dinb(n8332), .dout(n8335));
  jnot g08080(.din(n8335), .dout(n8336));
  jor  g08081(.dina(n7266), .dinb(n428), .dout(n8337));
  jor  g08082(.dina(n7021), .dinb(n357), .dout(n8338));
  jor  g08083(.dina(n7269), .dinb(n395), .dout(n8339));
  jor  g08084(.dina(n7271), .dinb(n431), .dout(n8340));
  jand g08085(.dina(n8340), .dinb(n8339), .dout(n8341));
  jand g08086(.dina(n8341), .dinb(n8338), .dout(n8342));
  jand g08087(.dina(n8342), .dinb(n8337), .dout(n8343));
  jxor g08088(.dina(n8343), .dinb(a50 ), .dout(n8344));
  jnot g08089(.din(n8344), .dout(n8345));
  jnot g08090(.din(n8140), .dout(n8346));
  jand g08091(.dina(n8346), .dinb(n8138), .dout(n8347));
  jand g08092(.dina(n8141), .dinb(n8136), .dout(n8348));
  jor  g08093(.dina(n8348), .dinb(n8347), .dout(n8349));
  jor  g08094(.dina(n8125), .dinb(n319), .dout(n8350));
  jor  g08095(.dina(n7846), .dinb(n279), .dout(n8351));
  jor  g08096(.dina(n8128), .dinb(n299), .dout(n8352));
  jor  g08097(.dina(n8130), .dinb(n322), .dout(n8353));
  jand g08098(.dina(n8353), .dinb(n8352), .dout(n8354));
  jand g08099(.dina(n8354), .dinb(n8351), .dout(n8355));
  jand g08100(.dina(n8355), .dinb(n8350), .dout(n8356));
  jxor g08101(.dina(n8356), .dinb(a53 ), .dout(n8357));
  jnot g08102(.din(n8357), .dout(n8358));
  jand g08103(.dina(n8138), .dinb(a56 ), .dout(n8359));
  jxor g08104(.dina(a56 ), .dinb(a55 ), .dout(n8360));
  jnot g08105(.din(n8360), .dout(n8361));
  jand g08106(.dina(n8361), .dinb(n8137), .dout(n8362));
  jand g08107(.dina(n8362), .dinb(b1 ), .dout(n8363));
  jnot g08108(.din(n8137), .dout(n8364));
  jxor g08109(.dina(a55 ), .dinb(a54 ), .dout(n8365));
  jand g08110(.dina(n8365), .dinb(n8364), .dout(n8366));
  jand g08111(.dina(n8366), .dinb(b0 ), .dout(n8367));
  jand g08112(.dina(n8360), .dinb(n8137), .dout(n8368));
  jand g08113(.dina(n8368), .dinb(n338), .dout(n8369));
  jor  g08114(.dina(n8369), .dinb(n8367), .dout(n8370));
  jor  g08115(.dina(n8370), .dinb(n8363), .dout(n8371));
  jxor g08116(.dina(n8371), .dinb(n8359), .dout(n8372));
  jxor g08117(.dina(n8372), .dinb(n8358), .dout(n8373));
  jxor g08118(.dina(n8373), .dinb(n8349), .dout(n8374));
  jxor g08119(.dina(n8374), .dinb(n8345), .dout(n8375));
  jxor g08120(.dina(n8375), .dinb(n8336), .dout(n8376));
  jxor g08121(.dina(n8376), .dinb(n8331), .dout(n8377));
  jxor g08122(.dina(n8377), .dinb(n8322), .dout(n8378));
  jxor g08123(.dina(n8378), .dinb(n8319), .dout(n8379));
  jxor g08124(.dina(n8379), .dinb(n8310), .dout(n8380));
  jnot g08125(.din(n8380), .dout(n8381));
  jor  g08126(.dina(n5096), .dinb(n1019), .dout(n8382));
  jor  g08127(.dina(n4904), .dinb(n858), .dout(n8383));
  jor  g08128(.dina(n5099), .dinb(n939), .dout(n8384));
  jor  g08129(.dina(n5101), .dinb(n1022), .dout(n8385));
  jand g08130(.dina(n8385), .dinb(n8384), .dout(n8386));
  jand g08131(.dina(n8386), .dinb(n8383), .dout(n8387));
  jand g08132(.dina(n8387), .dinb(n8382), .dout(n8388));
  jxor g08133(.dina(n8388), .dinb(a41 ), .dout(n8389));
  jxor g08134(.dina(n8389), .dinb(n8381), .dout(n8390));
  jxor g08135(.dina(n8390), .dinb(n8307), .dout(n8391));
  jnot g08136(.din(n8391), .dout(n8392));
  jor  g08137(.dina(n4415), .dinb(n1397), .dout(n8393));
  jor  g08138(.dina(n4272), .dinb(n1193), .dout(n8394));
  jor  g08139(.dina(n4418), .dinb(n1290), .dout(n8395));
  jor  g08140(.dina(n4420), .dinb(n1400), .dout(n8396));
  jand g08141(.dina(n8396), .dinb(n8395), .dout(n8397));
  jand g08142(.dina(n8397), .dinb(n8394), .dout(n8398));
  jand g08143(.dina(n8398), .dinb(n8393), .dout(n8399));
  jxor g08144(.dina(n8399), .dinb(a38 ), .dout(n8400));
  jxor g08145(.dina(n8400), .dinb(n8392), .dout(n8401));
  jxor g08146(.dina(n8401), .dinb(n8304), .dout(n8402));
  jnot g08147(.din(n8402), .dout(n8403));
  jor  g08148(.dina(n3849), .dinb(n1739), .dout(n8404));
  jor  g08149(.dina(n3689), .dinb(n1420), .dout(n8405));
  jor  g08150(.dina(n3852), .dinb(n1620), .dout(n8406));
  jor  g08151(.dina(n3854), .dinb(n1742), .dout(n8407));
  jand g08152(.dina(n8407), .dinb(n8406), .dout(n8408));
  jand g08153(.dina(n8408), .dinb(n8405), .dout(n8409));
  jand g08154(.dina(n8409), .dinb(n8404), .dout(n8410));
  jxor g08155(.dina(n8410), .dinb(a35 ), .dout(n8411));
  jxor g08156(.dina(n8411), .dinb(n8403), .dout(n8412));
  jxor g08157(.dina(n8412), .dinb(n8301), .dout(n8413));
  jnot g08158(.din(n8413), .dout(n8414));
  jor  g08159(.dina(n3301), .dinb(n2007), .dout(n8415));
  jor  g08160(.dina(n3136), .dinb(n1867), .dout(n8416));
  jor  g08161(.dina(n3304), .dinb(n1887), .dout(n8417));
  jor  g08162(.dina(n3306), .dinb(n2010), .dout(n8418));
  jand g08163(.dina(n8418), .dinb(n8417), .dout(n8419));
  jand g08164(.dina(n8419), .dinb(n8416), .dout(n8420));
  jand g08165(.dina(n8420), .dinb(n8415), .dout(n8421));
  jxor g08166(.dina(n8421), .dinb(a32 ), .dout(n8422));
  jxor g08167(.dina(n8422), .dinb(n8414), .dout(n8423));
  jxor g08168(.dina(n8423), .dinb(n8298), .dout(n8424));
  jnot g08169(.din(n8424), .dout(n8425));
  jor  g08170(.dina(n2556), .dinb(n2784), .dout(n8426));
  jor  g08171(.dina(n2661), .dinb(n2148), .dout(n8427));
  jor  g08172(.dina(n2787), .dinb(n2407), .dout(n8428));
  jor  g08173(.dina(n2789), .dinb(n2559), .dout(n8429));
  jand g08174(.dina(n8429), .dinb(n8428), .dout(n8430));
  jand g08175(.dina(n8430), .dinb(n8427), .dout(n8431));
  jand g08176(.dina(n8431), .dinb(n8426), .dout(n8432));
  jxor g08177(.dina(n8432), .dinb(a29 ), .dout(n8433));
  jxor g08178(.dina(n8433), .dinb(n8425), .dout(n8434));
  jxor g08179(.dina(n8434), .dinb(n8295), .dout(n8435));
  jnot g08180(.din(n8435), .dout(n8436));
  jor  g08181(.dina(n3032), .dinb(n2319), .dout(n8437));
  jor  g08182(.dina(n2224), .dinb(n2579), .dout(n8438));
  jor  g08183(.dina(n2322), .dinb(n2870), .dout(n8439));
  jor  g08184(.dina(n2324), .dinb(n3035), .dout(n8440));
  jand g08185(.dina(n8440), .dinb(n8439), .dout(n8441));
  jand g08186(.dina(n8441), .dinb(n8438), .dout(n8442));
  jand g08187(.dina(n8442), .dinb(n8437), .dout(n8443));
  jxor g08188(.dina(n8443), .dinb(a26 ), .dout(n8444));
  jxor g08189(.dina(n8444), .dinb(n8436), .dout(n8445));
  jxor g08190(.dina(n8445), .dinb(n8292), .dout(n8446));
  jor  g08191(.dina(n3400), .dinb(n1939), .dout(n8447));
  jor  g08192(.dina(n1827), .dinb(n3055), .dout(n8448));
  jor  g08193(.dina(n1942), .dinb(n3230), .dout(n8449));
  jor  g08194(.dina(n1944), .dinb(n3403), .dout(n8450));
  jand g08195(.dina(n8450), .dinb(n8449), .dout(n8451));
  jand g08196(.dina(n8451), .dinb(n8448), .dout(n8452));
  jand g08197(.dina(n8452), .dinb(n8447), .dout(n8453));
  jxor g08198(.dina(n8453), .dinb(a23 ), .dout(n8454));
  jxor g08199(.dina(n8454), .dinb(n8446), .dout(n8455));
  jnot g08200(.din(n8455), .dout(n8456));
  jxor g08201(.dina(n8456), .dinb(n8289), .dout(n8457));
  jor  g08202(.dina(n4137), .dinb(n1566), .dout(n8458));
  jor  g08203(.dina(n1489), .dinb(n3588), .dout(n8459));
  jor  g08204(.dina(n1569), .dinb(n3942), .dout(n8460));
  jor  g08205(.dina(n1571), .dinb(n4140), .dout(n8461));
  jand g08206(.dina(n8461), .dinb(n8460), .dout(n8462));
  jand g08207(.dina(n8462), .dinb(n8459), .dout(n8463));
  jand g08208(.dina(n8463), .dinb(n8458), .dout(n8464));
  jxor g08209(.dina(n8464), .dinb(a20 ), .dout(n8465));
  jxor g08210(.dina(n8465), .dinb(n8457), .dout(n8466));
  jxor g08211(.dina(n8466), .dinb(n8281), .dout(n8467));
  jor  g08212(.dina(n4554), .dinb(n1245), .dout(n8468));
  jor  g08213(.dina(n1165), .dinb(n4340), .dout(n8469));
  jor  g08214(.dina(n1248), .dinb(n4537), .dout(n8470));
  jor  g08215(.dina(n1250), .dinb(n4557), .dout(n8471));
  jand g08216(.dina(n8471), .dinb(n8470), .dout(n8472));
  jand g08217(.dina(n8472), .dinb(n8469), .dout(n8473));
  jand g08218(.dina(n8473), .dinb(n8468), .dout(n8474));
  jxor g08219(.dina(n8474), .dinb(a17 ), .dout(n8475));
  jxor g08220(.dina(n8475), .dinb(n8467), .dout(n8476));
  jxor g08221(.dina(n8476), .dinb(n8276), .dout(n8477));
  jnot g08222(.din(n8477), .dout(n8478));
  jor  g08223(.dina(n5405), .dinb(n974), .dout(n8479));
  jor  g08224(.dina(n908), .dinb(n4974), .dout(n8480));
  jor  g08225(.dina(n977), .dinb(n4994), .dout(n8481));
  jor  g08226(.dina(n979), .dinb(n5408), .dout(n8482));
  jand g08227(.dina(n8482), .dinb(n8481), .dout(n8483));
  jand g08228(.dina(n8483), .dinb(n8480), .dout(n8484));
  jand g08229(.dina(n8484), .dinb(n8479), .dout(n8485));
  jxor g08230(.dina(n8485), .dinb(a14 ), .dout(n8486));
  jxor g08231(.dina(n8486), .dinb(n8478), .dout(n8487));
  jxor g08232(.dina(n8487), .dinb(n8272), .dout(n8488));
  jxor g08233(.dina(n8488), .dinb(n8268), .dout(n8489));
  jxor g08234(.dina(n8489), .dinb(n8260), .dout(n8490));
  jxor g08235(.dina(n8490), .dinb(n8255), .dout(n8491));
  jxor g08236(.dina(n8491), .dinb(n8246), .dout(n8492));
  jor  g08237(.dina(n7408), .dinb(n402), .dout(n8493));
  jor  g08238(.dina(n371), .dinb(n7129), .dout(n8494));
  jor  g08239(.dina(n405), .dinb(n7149), .dout(n8495));
  jor  g08240(.dina(n332), .dinb(n7411), .dout(n8496));
  jand g08241(.dina(n8496), .dinb(n8495), .dout(n8497));
  jand g08242(.dina(n8497), .dinb(n8494), .dout(n8498));
  jand g08243(.dina(n8498), .dinb(n8493), .dout(n8499));
  jxor g08244(.dina(n8499), .dinb(a5 ), .dout(n8500));
  jnot g08245(.din(n8500), .dout(n8501));
  jxor g08246(.dina(n8501), .dinb(n8492), .dout(n8502));
  jxor g08247(.dina(n8502), .dinb(n8241), .dout(n8503));
  jxor g08248(.dina(n8503), .dinb(n8237), .dout(n8504));
  jxor g08249(.dina(n8504), .dinb(n8222), .dout(f55 ));
  jand g08250(.dina(n8503), .dinb(n8237), .dout(n8506));
  jand g08251(.dina(n8504), .dinb(n8222), .dout(n8507));
  jor  g08252(.dina(n8507), .dinb(n8506), .dout(n8508));
  jand g08253(.dina(n8501), .dinb(n8492), .dout(n8509));
  jand g08254(.dina(n8502), .dinb(n8241), .dout(n8510));
  jor  g08255(.dina(n8510), .dinb(n8509), .dout(n8511));
  jor  g08256(.dina(n7680), .dinb(n402), .dout(n8512));
  jor  g08257(.dina(n371), .dinb(n7149), .dout(n8513));
  jor  g08258(.dina(n405), .dinb(n7411), .dout(n8514));
  jor  g08259(.dina(n332), .dinb(n7683), .dout(n8515));
  jand g08260(.dina(n8515), .dinb(n8514), .dout(n8516));
  jand g08261(.dina(n8516), .dinb(n8513), .dout(n8517));
  jand g08262(.dina(n8517), .dinb(n8512), .dout(n8518));
  jxor g08263(.dina(n8518), .dinb(a5 ), .dout(n8519));
  jnot g08264(.din(n8519), .dout(n8520));
  jand g08265(.dina(n8490), .dinb(n8255), .dout(n8521));
  jand g08266(.dina(n8491), .dinb(n8246), .dout(n8522));
  jor  g08267(.dina(n8522), .dinb(n8521), .dout(n8523));
  jor  g08268(.dina(n7126), .dinb(n528), .dout(n8524));
  jor  g08269(.dina(n490), .dinb(n6372), .dout(n8525));
  jor  g08270(.dina(n531), .dinb(n6867), .dout(n8526));
  jor  g08271(.dina(n533), .dinb(n7129), .dout(n8527));
  jand g08272(.dina(n8527), .dinb(n8526), .dout(n8528));
  jand g08273(.dina(n8528), .dinb(n8525), .dout(n8529));
  jand g08274(.dina(n8529), .dinb(n8524), .dout(n8530));
  jxor g08275(.dina(n8530), .dinb(a8 ), .dout(n8531));
  jnot g08276(.din(n8531), .dout(n8532));
  jnot g08277(.din(n8268), .dout(n8533));
  jand g08278(.dina(n8488), .dinb(n8533), .dout(n8534));
  jnot g08279(.din(n8534), .dout(n8535));
  jor  g08280(.dina(n8489), .dinb(n8260), .dout(n8536));
  jand g08281(.dina(n8536), .dinb(n8535), .dout(n8537));
  jor  g08282(.dina(n8486), .dinb(n8478), .dout(n8538));
  jnot g08283(.din(n8538), .dout(n8539));
  jand g08284(.dina(n8487), .dinb(n8272), .dout(n8540));
  jor  g08285(.dina(n8540), .dinb(n8539), .dout(n8541));
  jor  g08286(.dina(n8475), .dinb(n8467), .dout(n8542));
  jnot g08287(.din(n8542), .dout(n8543));
  jand g08288(.dina(n8476), .dinb(n8276), .dout(n8544));
  jor  g08289(.dina(n8544), .dinb(n8543), .dout(n8545));
  jor  g08290(.dina(n8465), .dinb(n8457), .dout(n8546));
  jnot g08291(.din(n8283), .dout(n8547));
  jand g08292(.dina(n8179), .dinb(n8023), .dout(n8548));
  jor  g08293(.dina(n8548), .dinb(n8547), .dout(n8549));
  jxor g08294(.dina(n8456), .dinb(n8549), .dout(n8550));
  jxor g08295(.dina(n8465), .dinb(n8550), .dout(n8551));
  jor  g08296(.dina(n8551), .dinb(n8281), .dout(n8552));
  jand g08297(.dina(n8552), .dinb(n8546), .dout(n8553));
  jnot g08298(.din(n8446), .dout(n8554));
  jor  g08299(.dina(n8454), .dinb(n8554), .dout(n8555));
  jor  g08300(.dina(n8455), .dinb(n8289), .dout(n8556));
  jand g08301(.dina(n8556), .dinb(n8555), .dout(n8557));
  jor  g08302(.dina(n8444), .dinb(n8436), .dout(n8558));
  jnot g08303(.din(n8558), .dout(n8559));
  jand g08304(.dina(n8445), .dinb(n8292), .dout(n8560));
  jor  g08305(.dina(n8560), .dinb(n8559), .dout(n8561));
  jor  g08306(.dina(n3052), .dinb(n2319), .dout(n8562));
  jor  g08307(.dina(n2224), .dinb(n2870), .dout(n8563));
  jor  g08308(.dina(n2322), .dinb(n3035), .dout(n8564));
  jor  g08309(.dina(n2324), .dinb(n3055), .dout(n8565));
  jand g08310(.dina(n8565), .dinb(n8564), .dout(n8566));
  jand g08311(.dina(n8566), .dinb(n8563), .dout(n8567));
  jand g08312(.dina(n8567), .dinb(n8562), .dout(n8568));
  jxor g08313(.dina(n8568), .dinb(a26 ), .dout(n8569));
  jnot g08314(.din(n8569), .dout(n8570));
  jor  g08315(.dina(n8433), .dinb(n8425), .dout(n8571));
  jand g08316(.dina(n8434), .dinb(n8295), .dout(n8572));
  jnot g08317(.din(n8572), .dout(n8573));
  jand g08318(.dina(n8573), .dinb(n8571), .dout(n8574));
  jnot g08319(.din(n8574), .dout(n8575));
  jor  g08320(.dina(n2576), .dinb(n2784), .dout(n8576));
  jor  g08321(.dina(n2661), .dinb(n2407), .dout(n8577));
  jor  g08322(.dina(n2787), .dinb(n2559), .dout(n8578));
  jor  g08323(.dina(n2789), .dinb(n2579), .dout(n8579));
  jand g08324(.dina(n8579), .dinb(n8578), .dout(n8580));
  jand g08325(.dina(n8580), .dinb(n8577), .dout(n8581));
  jand g08326(.dina(n8581), .dinb(n8576), .dout(n8582));
  jxor g08327(.dina(n8582), .dinb(a29 ), .dout(n8583));
  jnot g08328(.din(n8583), .dout(n8584));
  jor  g08329(.dina(n8422), .dinb(n8414), .dout(n8585));
  jand g08330(.dina(n8423), .dinb(n8298), .dout(n8586));
  jnot g08331(.din(n8586), .dout(n8587));
  jand g08332(.dina(n8587), .dinb(n8585), .dout(n8588));
  jnot g08333(.din(n8588), .dout(n8589));
  jor  g08334(.dina(n8411), .dinb(n8403), .dout(n8590));
  jand g08335(.dina(n8412), .dinb(n8301), .dout(n8591));
  jnot g08336(.din(n8591), .dout(n8592));
  jand g08337(.dina(n8592), .dinb(n8590), .dout(n8593));
  jnot g08338(.din(n8593), .dout(n8594));
  jor  g08339(.dina(n3849), .dinb(n1864), .dout(n8595));
  jor  g08340(.dina(n3689), .dinb(n1620), .dout(n8596));
  jor  g08341(.dina(n3852), .dinb(n1742), .dout(n8597));
  jor  g08342(.dina(n3854), .dinb(n1867), .dout(n8598));
  jand g08343(.dina(n8598), .dinb(n8597), .dout(n8599));
  jand g08344(.dina(n8599), .dinb(n8596), .dout(n8600));
  jand g08345(.dina(n8600), .dinb(n8595), .dout(n8601));
  jxor g08346(.dina(n8601), .dinb(a35 ), .dout(n8602));
  jnot g08347(.din(n8602), .dout(n8603));
  jor  g08348(.dina(n8400), .dinb(n8392), .dout(n8604));
  jand g08349(.dina(n8401), .dinb(n8304), .dout(n8605));
  jnot g08350(.din(n8605), .dout(n8606));
  jand g08351(.dina(n8606), .dinb(n8604), .dout(n8607));
  jnot g08352(.din(n8607), .dout(n8608));
  jor  g08353(.dina(n4415), .dinb(n1417), .dout(n8609));
  jor  g08354(.dina(n4272), .dinb(n1290), .dout(n8610));
  jor  g08355(.dina(n4418), .dinb(n1400), .dout(n8611));
  jor  g08356(.dina(n4420), .dinb(n1420), .dout(n8612));
  jand g08357(.dina(n8612), .dinb(n8611), .dout(n8613));
  jand g08358(.dina(n8613), .dinb(n8610), .dout(n8614));
  jand g08359(.dina(n8614), .dinb(n8609), .dout(n8615));
  jxor g08360(.dina(n8615), .dinb(a38 ), .dout(n8616));
  jnot g08361(.din(n8616), .dout(n8617));
  jor  g08362(.dina(n8389), .dinb(n8381), .dout(n8618));
  jand g08363(.dina(n8390), .dinb(n8307), .dout(n8619));
  jnot g08364(.din(n8619), .dout(n8620));
  jand g08365(.dina(n8620), .dinb(n8618), .dout(n8621));
  jnot g08366(.din(n8621), .dout(n8622));
  jor  g08367(.dina(n5096), .dinb(n1190), .dout(n8623));
  jor  g08368(.dina(n4904), .dinb(n939), .dout(n8624));
  jor  g08369(.dina(n5099), .dinb(n1022), .dout(n8625));
  jor  g08370(.dina(n5101), .dinb(n1193), .dout(n8626));
  jand g08371(.dina(n8626), .dinb(n8625), .dout(n8627));
  jand g08372(.dina(n8627), .dinb(n8624), .dout(n8628));
  jand g08373(.dina(n8628), .dinb(n8623), .dout(n8629));
  jxor g08374(.dina(n8629), .dinb(a41 ), .dout(n8630));
  jnot g08375(.din(n8630), .dout(n8631));
  jand g08376(.dina(n8378), .dinb(n8319), .dout(n8632));
  jand g08377(.dina(n8379), .dinb(n8310), .dout(n8633));
  jor  g08378(.dina(n8633), .dinb(n8632), .dout(n8634));
  jand g08379(.dina(n8376), .dinb(n8331), .dout(n8635));
  jand g08380(.dina(n8377), .dinb(n8322), .dout(n8636));
  jor  g08381(.dina(n8636), .dinb(n8635), .dout(n8637));
  jor  g08382(.dina(n6490), .dinb(n644), .dout(n8638));
  jor  g08383(.dina(n6262), .dinb(n564), .dout(n8639));
  jor  g08384(.dina(n6493), .dinb(n627), .dout(n8640));
  jor  g08385(.dina(n6495), .dinb(n647), .dout(n8641));
  jand g08386(.dina(n8641), .dinb(n8640), .dout(n8642));
  jand g08387(.dina(n8642), .dinb(n8639), .dout(n8643));
  jand g08388(.dina(n8643), .dinb(n8638), .dout(n8644));
  jxor g08389(.dina(n8644), .dinb(a47 ), .dout(n8645));
  jnot g08390(.din(n8645), .dout(n8646));
  jand g08391(.dina(n8374), .dinb(n8345), .dout(n8647));
  jand g08392(.dina(n8375), .dinb(n8336), .dout(n8648));
  jor  g08393(.dina(n8648), .dinb(n8647), .dout(n8649));
  jor  g08394(.dina(n7266), .dinb(n509), .dout(n8650));
  jor  g08395(.dina(n7021), .dinb(n395), .dout(n8651));
  jor  g08396(.dina(n7269), .dinb(n431), .dout(n8652));
  jor  g08397(.dina(n7271), .dinb(n512), .dout(n8653));
  jand g08398(.dina(n8653), .dinb(n8652), .dout(n8654));
  jand g08399(.dina(n8654), .dinb(n8651), .dout(n8655));
  jand g08400(.dina(n8655), .dinb(n8650), .dout(n8656));
  jxor g08401(.dina(n8656), .dinb(a50 ), .dout(n8657));
  jnot g08402(.din(n8657), .dout(n8658));
  jand g08403(.dina(n8372), .dinb(n8358), .dout(n8659));
  jand g08404(.dina(n8373), .dinb(n8349), .dout(n8660));
  jor  g08405(.dina(n8660), .dinb(n8659), .dout(n8661));
  jor  g08406(.dina(n8125), .dinb(n354), .dout(n8662));
  jor  g08407(.dina(n7846), .dinb(n299), .dout(n8663));
  jor  g08408(.dina(n8128), .dinb(n322), .dout(n8664));
  jor  g08409(.dina(n8130), .dinb(n357), .dout(n8665));
  jand g08410(.dina(n8665), .dinb(n8664), .dout(n8666));
  jand g08411(.dina(n8666), .dinb(n8663), .dout(n8667));
  jand g08412(.dina(n8667), .dinb(n8662), .dout(n8668));
  jxor g08413(.dina(n8668), .dinb(a53 ), .dout(n8669));
  jnot g08414(.din(n8669), .dout(n8670));
  jnot g08415(.din(n8371), .dout(n8671));
  jand g08416(.dina(n8139), .dinb(a56 ), .dout(n8672));
  jand g08417(.dina(n8672), .dinb(n8671), .dout(n8673));
  jnot g08418(.din(n8673), .dout(n8674));
  jand g08419(.dina(n8674), .dinb(a56 ), .dout(n8675));
  jor  g08420(.dina(n8365), .dinb(n8361), .dout(n8676));
  jor  g08421(.dina(n8676), .dinb(n8137), .dout(n8677));
  jnot g08422(.din(n8677), .dout(n8678));
  jand g08423(.dina(n8678), .dinb(b0 ), .dout(n8679));
  jand g08424(.dina(n8362), .dinb(b2 ), .dout(n8680));
  jand g08425(.dina(n8366), .dinb(b1 ), .dout(n8681));
  jand g08426(.dina(n8368), .dinb(n375), .dout(n8682));
  jor  g08427(.dina(n8682), .dinb(n8681), .dout(n8683));
  jor  g08428(.dina(n8683), .dinb(n8680), .dout(n8684));
  jor  g08429(.dina(n8684), .dinb(n8679), .dout(n8685));
  jxor g08430(.dina(n8685), .dinb(n8675), .dout(n8686));
  jxor g08431(.dina(n8686), .dinb(n8670), .dout(n8687));
  jxor g08432(.dina(n8687), .dinb(n8661), .dout(n8688));
  jxor g08433(.dina(n8688), .dinb(n8658), .dout(n8689));
  jxor g08434(.dina(n8689), .dinb(n8649), .dout(n8690));
  jxor g08435(.dina(n8690), .dinb(n8646), .dout(n8691));
  jxor g08436(.dina(n8691), .dinb(n8637), .dout(n8692));
  jnot g08437(.din(n8692), .dout(n8693));
  jor  g08438(.dina(n5739), .dinb(n855), .dout(n8694));
  jor  g08439(.dina(n5574), .dinb(n758), .dout(n8695));
  jor  g08440(.dina(n5742), .dinb(n778), .dout(n8696));
  jor  g08441(.dina(n5744), .dinb(n858), .dout(n8697));
  jand g08442(.dina(n8697), .dinb(n8696), .dout(n8698));
  jand g08443(.dina(n8698), .dinb(n8695), .dout(n8699));
  jand g08444(.dina(n8699), .dinb(n8694), .dout(n8700));
  jxor g08445(.dina(n8700), .dinb(a44 ), .dout(n8701));
  jxor g08446(.dina(n8701), .dinb(n8693), .dout(n8702));
  jxor g08447(.dina(n8702), .dinb(n8634), .dout(n8703));
  jxor g08448(.dina(n8703), .dinb(n8631), .dout(n8704));
  jxor g08449(.dina(n8704), .dinb(n8622), .dout(n8705));
  jxor g08450(.dina(n8705), .dinb(n8617), .dout(n8706));
  jxor g08451(.dina(n8706), .dinb(n8608), .dout(n8707));
  jxor g08452(.dina(n8707), .dinb(n8603), .dout(n8708));
  jxor g08453(.dina(n8708), .dinb(n8594), .dout(n8709));
  jnot g08454(.din(n8709), .dout(n8710));
  jor  g08455(.dina(n3301), .dinb(n2145), .dout(n8711));
  jor  g08456(.dina(n3136), .dinb(n1887), .dout(n8712));
  jor  g08457(.dina(n3304), .dinb(n2010), .dout(n8713));
  jor  g08458(.dina(n3306), .dinb(n2148), .dout(n8714));
  jand g08459(.dina(n8714), .dinb(n8713), .dout(n8715));
  jand g08460(.dina(n8715), .dinb(n8712), .dout(n8716));
  jand g08461(.dina(n8716), .dinb(n8711), .dout(n8717));
  jxor g08462(.dina(n8717), .dinb(a32 ), .dout(n8718));
  jxor g08463(.dina(n8718), .dinb(n8710), .dout(n8719));
  jxor g08464(.dina(n8719), .dinb(n8589), .dout(n8720));
  jxor g08465(.dina(n8720), .dinb(n8584), .dout(n8721));
  jxor g08466(.dina(n8721), .dinb(n8575), .dout(n8722));
  jxor g08467(.dina(n8722), .dinb(n8570), .dout(n8723));
  jxor g08468(.dina(n8723), .dinb(n8561), .dout(n8724));
  jor  g08469(.dina(n3585), .dinb(n1939), .dout(n8725));
  jor  g08470(.dina(n1827), .dinb(n3230), .dout(n8726));
  jor  g08471(.dina(n1942), .dinb(n3403), .dout(n8727));
  jor  g08472(.dina(n1944), .dinb(n3588), .dout(n8728));
  jand g08473(.dina(n8728), .dinb(n8727), .dout(n8729));
  jand g08474(.dina(n8729), .dinb(n8726), .dout(n8730));
  jand g08475(.dina(n8730), .dinb(n8725), .dout(n8731));
  jxor g08476(.dina(n8731), .dinb(a23 ), .dout(n8732));
  jxor g08477(.dina(n8732), .dinb(n8724), .dout(n8733));
  jnot g08478(.din(n8733), .dout(n8734));
  jxor g08479(.dina(n8734), .dinb(n8557), .dout(n8735));
  jor  g08480(.dina(n4337), .dinb(n1566), .dout(n8736));
  jor  g08481(.dina(n1489), .dinb(n3942), .dout(n8737));
  jor  g08482(.dina(n1569), .dinb(n4140), .dout(n8738));
  jor  g08483(.dina(n1571), .dinb(n4340), .dout(n8739));
  jand g08484(.dina(n8739), .dinb(n8738), .dout(n8740));
  jand g08485(.dina(n8740), .dinb(n8737), .dout(n8741));
  jand g08486(.dina(n8741), .dinb(n8736), .dout(n8742));
  jxor g08487(.dina(n8742), .dinb(a20 ), .dout(n8743));
  jxor g08488(.dina(n8743), .dinb(n8735), .dout(n8744));
  jxor g08489(.dina(n8744), .dinb(n8553), .dout(n8745));
  jor  g08490(.dina(n4971), .dinb(n1245), .dout(n8746));
  jor  g08491(.dina(n1165), .dinb(n4537), .dout(n8747));
  jor  g08492(.dina(n1248), .dinb(n4557), .dout(n8748));
  jor  g08493(.dina(n1250), .dinb(n4974), .dout(n8749));
  jand g08494(.dina(n8749), .dinb(n8748), .dout(n8750));
  jand g08495(.dina(n8750), .dinb(n8747), .dout(n8751));
  jand g08496(.dina(n8751), .dinb(n8746), .dout(n8752));
  jxor g08497(.dina(n8752), .dinb(a17 ), .dout(n8753));
  jxor g08498(.dina(n8753), .dinb(n8745), .dout(n8754));
  jxor g08499(.dina(n8754), .dinb(n8545), .dout(n8755));
  jnot g08500(.din(n8755), .dout(n8756));
  jor  g08501(.dina(n5425), .dinb(n974), .dout(n8757));
  jor  g08502(.dina(n908), .dinb(n4994), .dout(n8758));
  jor  g08503(.dina(n977), .dinb(n5408), .dout(n8759));
  jor  g08504(.dina(n979), .dinb(n5428), .dout(n8760));
  jand g08505(.dina(n8760), .dinb(n8759), .dout(n8761));
  jand g08506(.dina(n8761), .dinb(n8758), .dout(n8762));
  jand g08507(.dina(n8762), .dinb(n8757), .dout(n8763));
  jxor g08508(.dina(n8763), .dinb(a14 ), .dout(n8764));
  jxor g08509(.dina(n8764), .dinb(n8756), .dout(n8765));
  jxor g08510(.dina(n8765), .dinb(n8541), .dout(n8766));
  jor  g08511(.dina(n6349), .dinb(n706), .dout(n8767));
  jor  g08512(.dina(n683), .dinb(n5862), .dout(n8768));
  jor  g08513(.dina(n709), .dinb(n6106), .dout(n8769));
  jor  g08514(.dina(n711), .dinb(n6352), .dout(n8770));
  jand g08515(.dina(n8770), .dinb(n8769), .dout(n8771));
  jand g08516(.dina(n8771), .dinb(n8768), .dout(n8772));
  jand g08517(.dina(n8772), .dinb(n8767), .dout(n8773));
  jxor g08518(.dina(n8773), .dinb(a11 ), .dout(n8774));
  jxor g08519(.dina(n8774), .dinb(n8766), .dout(n8775));
  jxor g08520(.dina(n8775), .dinb(n8537), .dout(n8776));
  jxor g08521(.dina(n8776), .dinb(n8532), .dout(n8777));
  jxor g08522(.dina(n8777), .dinb(n8523), .dout(n8778));
  jxor g08523(.dina(n8778), .dinb(n8520), .dout(n8779));
  jxor g08524(.dina(n8779), .dinb(n8511), .dout(n8780));
  jand g08525(.dina(b55 ), .dinb(b54 ), .dout(n8781));
  jand g08526(.dina(n8226), .dinb(n8225), .dout(n8782));
  jor  g08527(.dina(n8782), .dinb(n8781), .dout(n8783));
  jxor g08528(.dina(b56 ), .dinb(b55 ), .dout(n8784));
  jnot g08529(.din(n8784), .dout(n8785));
  jxor g08530(.dina(n8785), .dinb(n8783), .dout(n8786));
  jor  g08531(.dina(n8786), .dinb(n264), .dout(n8787));
  jor  g08532(.dina(n284), .dinb(n7960), .dout(n8788));
  jnot g08533(.din(b56 ), .dout(n8789));
  jor  g08534(.dina(n269), .dinb(n8789), .dout(n8790));
  jor  g08535(.dina(n271), .dinb(n8231), .dout(n8791));
  jand g08536(.dina(n8791), .dinb(n8790), .dout(n8792));
  jand g08537(.dina(n8792), .dinb(n8788), .dout(n8793));
  jand g08538(.dina(n8793), .dinb(n8787), .dout(n8794));
  jxor g08539(.dina(n8794), .dinb(n260), .dout(n8795));
  jxor g08540(.dina(n8795), .dinb(n8780), .dout(n8796));
  jxor g08541(.dina(n8796), .dinb(n8508), .dout(f56 ));
  jand g08542(.dina(n8795), .dinb(n8780), .dout(n8798));
  jand g08543(.dina(n8796), .dinb(n8508), .dout(n8799));
  jor  g08544(.dina(n8799), .dinb(n8798), .dout(n8800));
  jand g08545(.dina(b56 ), .dinb(b55 ), .dout(n8801));
  jand g08546(.dina(n8784), .dinb(n8783), .dout(n8802));
  jor  g08547(.dina(n8802), .dinb(n8801), .dout(n8803));
  jxor g08548(.dina(b57 ), .dinb(b56 ), .dout(n8804));
  jnot g08549(.din(n8804), .dout(n8805));
  jxor g08550(.dina(n8805), .dinb(n8803), .dout(n8806));
  jor  g08551(.dina(n8806), .dinb(n264), .dout(n8807));
  jor  g08552(.dina(n284), .dinb(n8231), .dout(n8808));
  jnot g08553(.din(b57 ), .dout(n8809));
  jor  g08554(.dina(n269), .dinb(n8809), .dout(n8810));
  jor  g08555(.dina(n271), .dinb(n8789), .dout(n8811));
  jand g08556(.dina(n8811), .dinb(n8810), .dout(n8812));
  jand g08557(.dina(n8812), .dinb(n8808), .dout(n8813));
  jand g08558(.dina(n8813), .dinb(n8807), .dout(n8814));
  jxor g08559(.dina(n8814), .dinb(n260), .dout(n8815));
  jand g08560(.dina(n8778), .dinb(n8520), .dout(n8816));
  jand g08561(.dina(n8779), .dinb(n8511), .dout(n8817));
  jor  g08562(.dina(n8817), .dinb(n8816), .dout(n8818));
  jor  g08563(.dina(n7957), .dinb(n402), .dout(n8819));
  jor  g08564(.dina(n371), .dinb(n7411), .dout(n8820));
  jor  g08565(.dina(n405), .dinb(n7683), .dout(n8821));
  jor  g08566(.dina(n332), .dinb(n7960), .dout(n8822));
  jand g08567(.dina(n8822), .dinb(n8821), .dout(n8823));
  jand g08568(.dina(n8823), .dinb(n8820), .dout(n8824));
  jand g08569(.dina(n8824), .dinb(n8819), .dout(n8825));
  jxor g08570(.dina(n8825), .dinb(a5 ), .dout(n8826));
  jnot g08571(.din(n8826), .dout(n8827));
  jand g08572(.dina(n8776), .dinb(n8532), .dout(n8828));
  jand g08573(.dina(n8777), .dinb(n8523), .dout(n8829));
  jor  g08574(.dina(n8829), .dinb(n8828), .dout(n8830));
  jor  g08575(.dina(n7146), .dinb(n528), .dout(n8831));
  jor  g08576(.dina(n490), .dinb(n6867), .dout(n8832));
  jor  g08577(.dina(n531), .dinb(n7129), .dout(n8833));
  jor  g08578(.dina(n533), .dinb(n7149), .dout(n8834));
  jand g08579(.dina(n8834), .dinb(n8833), .dout(n8835));
  jand g08580(.dina(n8835), .dinb(n8832), .dout(n8836));
  jand g08581(.dina(n8836), .dinb(n8831), .dout(n8837));
  jxor g08582(.dina(n8837), .dinb(a8 ), .dout(n8838));
  jnot g08583(.din(n8838), .dout(n8839));
  jnot g08584(.din(n8766), .dout(n8840));
  jor  g08585(.dina(n8774), .dinb(n8840), .dout(n8841));
  jor  g08586(.dina(n8775), .dinb(n8537), .dout(n8842));
  jand g08587(.dina(n8842), .dinb(n8841), .dout(n8843));
  jor  g08588(.dina(n6369), .dinb(n706), .dout(n8844));
  jor  g08589(.dina(n683), .dinb(n6106), .dout(n8845));
  jor  g08590(.dina(n709), .dinb(n6352), .dout(n8846));
  jor  g08591(.dina(n711), .dinb(n6372), .dout(n8847));
  jand g08592(.dina(n8847), .dinb(n8846), .dout(n8848));
  jand g08593(.dina(n8848), .dinb(n8845), .dout(n8849));
  jand g08594(.dina(n8849), .dinb(n8844), .dout(n8850));
  jxor g08595(.dina(n8850), .dinb(a11 ), .dout(n8851));
  jor  g08596(.dina(n8764), .dinb(n8756), .dout(n8852));
  jnot g08597(.din(n8852), .dout(n8853));
  jand g08598(.dina(n8765), .dinb(n8541), .dout(n8854));
  jor  g08599(.dina(n8854), .dinb(n8853), .dout(n8855));
  jor  g08600(.dina(n5859), .dinb(n974), .dout(n8856));
  jor  g08601(.dina(n908), .dinb(n5408), .dout(n8857));
  jor  g08602(.dina(n977), .dinb(n5428), .dout(n8858));
  jor  g08603(.dina(n979), .dinb(n5862), .dout(n8859));
  jand g08604(.dina(n8859), .dinb(n8858), .dout(n8860));
  jand g08605(.dina(n8860), .dinb(n8857), .dout(n8861));
  jand g08606(.dina(n8861), .dinb(n8856), .dout(n8862));
  jxor g08607(.dina(n8862), .dinb(a14 ), .dout(n8863));
  jnot g08608(.din(n8863), .dout(n8864));
  jor  g08609(.dina(n8753), .dinb(n8745), .dout(n8865));
  jnot g08610(.din(n8865), .dout(n8866));
  jand g08611(.dina(n8754), .dinb(n8545), .dout(n8867));
  jor  g08612(.dina(n8867), .dinb(n8866), .dout(n8868));
  jor  g08613(.dina(n8743), .dinb(n8735), .dout(n8869));
  jnot g08614(.din(n8555), .dout(n8870));
  jand g08615(.dina(n8456), .dinb(n8549), .dout(n8871));
  jor  g08616(.dina(n8871), .dinb(n8870), .dout(n8872));
  jxor g08617(.dina(n8734), .dinb(n8872), .dout(n8873));
  jxor g08618(.dina(n8743), .dinb(n8873), .dout(n8874));
  jor  g08619(.dina(n8874), .dinb(n8553), .dout(n8875));
  jand g08620(.dina(n8875), .dinb(n8869), .dout(n8876));
  jnot g08621(.din(n8724), .dout(n8877));
  jor  g08622(.dina(n8732), .dinb(n8877), .dout(n8878));
  jor  g08623(.dina(n8733), .dinb(n8557), .dout(n8879));
  jand g08624(.dina(n8879), .dinb(n8878), .dout(n8880));
  jor  g08625(.dina(n3939), .dinb(n1939), .dout(n8881));
  jor  g08626(.dina(n1827), .dinb(n3403), .dout(n8882));
  jor  g08627(.dina(n1942), .dinb(n3588), .dout(n8883));
  jor  g08628(.dina(n1944), .dinb(n3942), .dout(n8884));
  jand g08629(.dina(n8884), .dinb(n8883), .dout(n8885));
  jand g08630(.dina(n8885), .dinb(n8882), .dout(n8886));
  jand g08631(.dina(n8886), .dinb(n8881), .dout(n8887));
  jxor g08632(.dina(n8887), .dinb(a23 ), .dout(n8888));
  jnot g08633(.din(n8888), .dout(n8889));
  jand g08634(.dina(n8722), .dinb(n8570), .dout(n8890));
  jand g08635(.dina(n8723), .dinb(n8561), .dout(n8891));
  jor  g08636(.dina(n8891), .dinb(n8890), .dout(n8892));
  jand g08637(.dina(n8720), .dinb(n8584), .dout(n8893));
  jand g08638(.dina(n8721), .dinb(n8575), .dout(n8894));
  jor  g08639(.dina(n8894), .dinb(n8893), .dout(n8895));
  jor  g08640(.dina(n2867), .dinb(n2784), .dout(n8896));
  jor  g08641(.dina(n2661), .dinb(n2559), .dout(n8897));
  jor  g08642(.dina(n2787), .dinb(n2579), .dout(n8898));
  jor  g08643(.dina(n2789), .dinb(n2870), .dout(n8899));
  jand g08644(.dina(n8899), .dinb(n8898), .dout(n8900));
  jand g08645(.dina(n8900), .dinb(n8897), .dout(n8901));
  jand g08646(.dina(n8901), .dinb(n8896), .dout(n8902));
  jxor g08647(.dina(n8902), .dinb(a29 ), .dout(n8903));
  jnot g08648(.din(n8903), .dout(n8904));
  jor  g08649(.dina(n8718), .dinb(n8710), .dout(n8905));
  jand g08650(.dina(n8719), .dinb(n8589), .dout(n8906));
  jnot g08651(.din(n8906), .dout(n8907));
  jand g08652(.dina(n8907), .dinb(n8905), .dout(n8908));
  jnot g08653(.din(n8908), .dout(n8909));
  jand g08654(.dina(n8707), .dinb(n8603), .dout(n8910));
  jand g08655(.dina(n8708), .dinb(n8594), .dout(n8911));
  jor  g08656(.dina(n8911), .dinb(n8910), .dout(n8912));
  jand g08657(.dina(n8705), .dinb(n8617), .dout(n8913));
  jand g08658(.dina(n8706), .dinb(n8608), .dout(n8914));
  jor  g08659(.dina(n8914), .dinb(n8913), .dout(n8915));
  jor  g08660(.dina(n4415), .dinb(n1617), .dout(n8916));
  jor  g08661(.dina(n4272), .dinb(n1400), .dout(n8917));
  jor  g08662(.dina(n4418), .dinb(n1420), .dout(n8918));
  jor  g08663(.dina(n4420), .dinb(n1620), .dout(n8919));
  jand g08664(.dina(n8919), .dinb(n8918), .dout(n8920));
  jand g08665(.dina(n8920), .dinb(n8917), .dout(n8921));
  jand g08666(.dina(n8921), .dinb(n8916), .dout(n8922));
  jxor g08667(.dina(n8922), .dinb(a38 ), .dout(n8923));
  jnot g08668(.din(n8923), .dout(n8924));
  jand g08669(.dina(n8703), .dinb(n8631), .dout(n8925));
  jand g08670(.dina(n8704), .dinb(n8622), .dout(n8926));
  jor  g08671(.dina(n8926), .dinb(n8925), .dout(n8927));
  jor  g08672(.dina(n5096), .dinb(n1287), .dout(n8928));
  jor  g08673(.dina(n4904), .dinb(n1022), .dout(n8929));
  jor  g08674(.dina(n5099), .dinb(n1193), .dout(n8930));
  jor  g08675(.dina(n5101), .dinb(n1290), .dout(n8931));
  jand g08676(.dina(n8931), .dinb(n8930), .dout(n8932));
  jand g08677(.dina(n8932), .dinb(n8929), .dout(n8933));
  jand g08678(.dina(n8933), .dinb(n8928), .dout(n8934));
  jxor g08679(.dina(n8934), .dinb(a41 ), .dout(n8935));
  jnot g08680(.din(n8935), .dout(n8936));
  jor  g08681(.dina(n8701), .dinb(n8693), .dout(n8937));
  jand g08682(.dina(n8702), .dinb(n8634), .dout(n8938));
  jnot g08683(.din(n8938), .dout(n8939));
  jand g08684(.dina(n8939), .dinb(n8937), .dout(n8940));
  jnot g08685(.din(n8940), .dout(n8941));
  jor  g08686(.dina(n5739), .dinb(n936), .dout(n8942));
  jor  g08687(.dina(n5574), .dinb(n778), .dout(n8943));
  jor  g08688(.dina(n5742), .dinb(n858), .dout(n8944));
  jor  g08689(.dina(n5744), .dinb(n939), .dout(n8945));
  jand g08690(.dina(n8945), .dinb(n8944), .dout(n8946));
  jand g08691(.dina(n8946), .dinb(n8943), .dout(n8947));
  jand g08692(.dina(n8947), .dinb(n8942), .dout(n8948));
  jxor g08693(.dina(n8948), .dinb(a44 ), .dout(n8949));
  jnot g08694(.din(n8949), .dout(n8950));
  jand g08695(.dina(n8690), .dinb(n8646), .dout(n8951));
  jand g08696(.dina(n8691), .dinb(n8637), .dout(n8952));
  jor  g08697(.dina(n8952), .dinb(n8951), .dout(n8953));
  jor  g08698(.dina(n6490), .dinb(n755), .dout(n8954));
  jor  g08699(.dina(n6262), .dinb(n627), .dout(n8955));
  jor  g08700(.dina(n6493), .dinb(n647), .dout(n8956));
  jor  g08701(.dina(n6495), .dinb(n758), .dout(n8957));
  jand g08702(.dina(n8957), .dinb(n8956), .dout(n8958));
  jand g08703(.dina(n8958), .dinb(n8955), .dout(n8959));
  jand g08704(.dina(n8959), .dinb(n8954), .dout(n8960));
  jxor g08705(.dina(n8960), .dinb(a47 ), .dout(n8961));
  jnot g08706(.din(n8961), .dout(n8962));
  jand g08707(.dina(n8688), .dinb(n8658), .dout(n8963));
  jand g08708(.dina(n8689), .dinb(n8649), .dout(n8964));
  jor  g08709(.dina(n8964), .dinb(n8963), .dout(n8965));
  jor  g08710(.dina(n7266), .dinb(n561), .dout(n8966));
  jor  g08711(.dina(n7021), .dinb(n431), .dout(n8967));
  jor  g08712(.dina(n7269), .dinb(n512), .dout(n8968));
  jor  g08713(.dina(n7271), .dinb(n564), .dout(n8969));
  jand g08714(.dina(n8969), .dinb(n8968), .dout(n8970));
  jand g08715(.dina(n8970), .dinb(n8967), .dout(n8971));
  jand g08716(.dina(n8971), .dinb(n8966), .dout(n8972));
  jxor g08717(.dina(n8972), .dinb(a50 ), .dout(n8973));
  jnot g08718(.din(n8973), .dout(n8974));
  jand g08719(.dina(n8686), .dinb(n8670), .dout(n8975));
  jand g08720(.dina(n8687), .dinb(n8661), .dout(n8976));
  jor  g08721(.dina(n8976), .dinb(n8975), .dout(n8977));
  jnot g08722(.din(n8368), .dout(n8978));
  jor  g08723(.dina(n8978), .dinb(n296), .dout(n8979));
  jor  g08724(.dina(n8677), .dinb(n267), .dout(n8980));
  jnot g08725(.din(n8366), .dout(n8981));
  jor  g08726(.dina(n8981), .dinb(n279), .dout(n8982));
  jnot g08727(.din(n8362), .dout(n8983));
  jor  g08728(.dina(n8983), .dinb(n299), .dout(n8984));
  jand g08729(.dina(n8984), .dinb(n8982), .dout(n8985));
  jand g08730(.dina(n8985), .dinb(n8980), .dout(n8986));
  jand g08731(.dina(n8986), .dinb(n8979), .dout(n8987));
  jxor g08732(.dina(n8987), .dinb(a56 ), .dout(n8988));
  jnot g08733(.din(n8988), .dout(n8989));
  jxor g08734(.dina(a57 ), .dinb(a56 ), .dout(n8990));
  jand g08735(.dina(n8990), .dinb(b0 ), .dout(n8991));
  jnot g08736(.din(n8991), .dout(n8992));
  jor  g08737(.dina(n8685), .dinb(n8674), .dout(n8993));
  jxor g08738(.dina(n8993), .dinb(n8992), .dout(n8994));
  jxor g08739(.dina(n8994), .dinb(n8989), .dout(n8995));
  jnot g08740(.din(n8995), .dout(n8996));
  jor  g08741(.dina(n8125), .dinb(n392), .dout(n8997));
  jor  g08742(.dina(n7846), .dinb(n322), .dout(n8998));
  jor  g08743(.dina(n8128), .dinb(n357), .dout(n8999));
  jor  g08744(.dina(n8130), .dinb(n395), .dout(n9000));
  jand g08745(.dina(n9000), .dinb(n8999), .dout(n9001));
  jand g08746(.dina(n9001), .dinb(n8998), .dout(n9002));
  jand g08747(.dina(n9002), .dinb(n8997), .dout(n9003));
  jxor g08748(.dina(n9003), .dinb(a53 ), .dout(n9004));
  jxor g08749(.dina(n9004), .dinb(n8996), .dout(n9005));
  jxor g08750(.dina(n9005), .dinb(n8977), .dout(n9006));
  jxor g08751(.dina(n9006), .dinb(n8974), .dout(n9007));
  jxor g08752(.dina(n9007), .dinb(n8965), .dout(n9008));
  jxor g08753(.dina(n9008), .dinb(n8962), .dout(n9009));
  jxor g08754(.dina(n9009), .dinb(n8953), .dout(n9010));
  jxor g08755(.dina(n9010), .dinb(n8950), .dout(n9011));
  jxor g08756(.dina(n9011), .dinb(n8941), .dout(n9012));
  jxor g08757(.dina(n9012), .dinb(n8936), .dout(n9013));
  jxor g08758(.dina(n9013), .dinb(n8927), .dout(n9014));
  jxor g08759(.dina(n9014), .dinb(n8924), .dout(n9015));
  jxor g08760(.dina(n9015), .dinb(n8915), .dout(n9016));
  jnot g08761(.din(n9016), .dout(n9017));
  jor  g08762(.dina(n3849), .dinb(n1884), .dout(n9018));
  jor  g08763(.dina(n3689), .dinb(n1742), .dout(n9019));
  jor  g08764(.dina(n3852), .dinb(n1867), .dout(n9020));
  jor  g08765(.dina(n3854), .dinb(n1887), .dout(n9021));
  jand g08766(.dina(n9021), .dinb(n9020), .dout(n9022));
  jand g08767(.dina(n9022), .dinb(n9019), .dout(n9023));
  jand g08768(.dina(n9023), .dinb(n9018), .dout(n9024));
  jxor g08769(.dina(n9024), .dinb(a35 ), .dout(n9025));
  jxor g08770(.dina(n9025), .dinb(n9017), .dout(n9026));
  jxor g08771(.dina(n9026), .dinb(n8912), .dout(n9027));
  jnot g08772(.din(n9027), .dout(n9028));
  jor  g08773(.dina(n3301), .dinb(n2404), .dout(n9029));
  jor  g08774(.dina(n3136), .dinb(n2010), .dout(n9030));
  jor  g08775(.dina(n3304), .dinb(n2148), .dout(n9031));
  jor  g08776(.dina(n3306), .dinb(n2407), .dout(n9032));
  jand g08777(.dina(n9032), .dinb(n9031), .dout(n9033));
  jand g08778(.dina(n9033), .dinb(n9030), .dout(n9034));
  jand g08779(.dina(n9034), .dinb(n9029), .dout(n9035));
  jxor g08780(.dina(n9035), .dinb(a32 ), .dout(n9036));
  jxor g08781(.dina(n9036), .dinb(n9028), .dout(n9037));
  jxor g08782(.dina(n9037), .dinb(n8909), .dout(n9038));
  jxor g08783(.dina(n9038), .dinb(n8904), .dout(n9039));
  jxor g08784(.dina(n9039), .dinb(n8895), .dout(n9040));
  jnot g08785(.din(n9040), .dout(n9041));
  jor  g08786(.dina(n3227), .dinb(n2319), .dout(n9042));
  jor  g08787(.dina(n2224), .dinb(n3035), .dout(n9043));
  jor  g08788(.dina(n2322), .dinb(n3055), .dout(n9044));
  jor  g08789(.dina(n2324), .dinb(n3230), .dout(n9045));
  jand g08790(.dina(n9045), .dinb(n9044), .dout(n9046));
  jand g08791(.dina(n9046), .dinb(n9043), .dout(n9047));
  jand g08792(.dina(n9047), .dinb(n9042), .dout(n9048));
  jxor g08793(.dina(n9048), .dinb(a26 ), .dout(n9049));
  jxor g08794(.dina(n9049), .dinb(n9041), .dout(n9050));
  jxor g08795(.dina(n9050), .dinb(n8892), .dout(n9051));
  jxor g08796(.dina(n9051), .dinb(n8889), .dout(n9052));
  jxor g08797(.dina(n9052), .dinb(n8880), .dout(n9053));
  jor  g08798(.dina(n4534), .dinb(n1566), .dout(n9054));
  jor  g08799(.dina(n1489), .dinb(n4140), .dout(n9055));
  jor  g08800(.dina(n1569), .dinb(n4340), .dout(n9056));
  jor  g08801(.dina(n1571), .dinb(n4537), .dout(n9057));
  jand g08802(.dina(n9057), .dinb(n9056), .dout(n9058));
  jand g08803(.dina(n9058), .dinb(n9055), .dout(n9059));
  jand g08804(.dina(n9059), .dinb(n9054), .dout(n9060));
  jxor g08805(.dina(n9060), .dinb(a20 ), .dout(n9061));
  jxor g08806(.dina(n9061), .dinb(n9053), .dout(n9062));
  jxor g08807(.dina(n9062), .dinb(n8876), .dout(n9063));
  jor  g08808(.dina(n4991), .dinb(n1245), .dout(n9064));
  jor  g08809(.dina(n1165), .dinb(n4557), .dout(n9065));
  jor  g08810(.dina(n1248), .dinb(n4974), .dout(n9066));
  jor  g08811(.dina(n1250), .dinb(n4994), .dout(n9067));
  jand g08812(.dina(n9067), .dinb(n9066), .dout(n9068));
  jand g08813(.dina(n9068), .dinb(n9065), .dout(n9069));
  jand g08814(.dina(n9069), .dinb(n9064), .dout(n9070));
  jxor g08815(.dina(n9070), .dinb(a17 ), .dout(n9071));
  jxor g08816(.dina(n9071), .dinb(n9063), .dout(n9072));
  jxor g08817(.dina(n9072), .dinb(n8868), .dout(n9073));
  jxor g08818(.dina(n9073), .dinb(n8864), .dout(n9074));
  jxor g08819(.dina(n9074), .dinb(n8855), .dout(n9075));
  jxor g08820(.dina(n9075), .dinb(n8851), .dout(n9076));
  jxor g08821(.dina(n9076), .dinb(n8843), .dout(n9077));
  jxor g08822(.dina(n9077), .dinb(n8839), .dout(n9078));
  jxor g08823(.dina(n9078), .dinb(n8830), .dout(n9079));
  jxor g08824(.dina(n9079), .dinb(n8827), .dout(n9080));
  jxor g08825(.dina(n9080), .dinb(n8818), .dout(n9081));
  jxor g08826(.dina(n9081), .dinb(n8815), .dout(n9082));
  jxor g08827(.dina(n9082), .dinb(n8800), .dout(f57 ));
  jand g08828(.dina(n9081), .dinb(n8815), .dout(n9084));
  jand g08829(.dina(n9082), .dinb(n8800), .dout(n9085));
  jor  g08830(.dina(n9085), .dinb(n9084), .dout(n9086));
  jand g08831(.dina(n9079), .dinb(n8827), .dout(n9087));
  jand g08832(.dina(n9080), .dinb(n8818), .dout(n9088));
  jor  g08833(.dina(n9088), .dinb(n9087), .dout(n9089));
  jor  g08834(.dina(n8228), .dinb(n402), .dout(n9090));
  jor  g08835(.dina(n371), .dinb(n7683), .dout(n9091));
  jor  g08836(.dina(n405), .dinb(n7960), .dout(n9092));
  jor  g08837(.dina(n332), .dinb(n8231), .dout(n9093));
  jand g08838(.dina(n9093), .dinb(n9092), .dout(n9094));
  jand g08839(.dina(n9094), .dinb(n9091), .dout(n9095));
  jand g08840(.dina(n9095), .dinb(n9090), .dout(n9096));
  jxor g08841(.dina(n9096), .dinb(a5 ), .dout(n9097));
  jnot g08842(.din(n9097), .dout(n9098));
  jand g08843(.dina(n9077), .dinb(n8839), .dout(n9099));
  jand g08844(.dina(n9078), .dinb(n8830), .dout(n9100));
  jor  g08845(.dina(n9100), .dinb(n9099), .dout(n9101));
  jor  g08846(.dina(n7408), .dinb(n528), .dout(n9102));
  jor  g08847(.dina(n490), .dinb(n7129), .dout(n9103));
  jor  g08848(.dina(n531), .dinb(n7149), .dout(n9104));
  jor  g08849(.dina(n533), .dinb(n7411), .dout(n9105));
  jand g08850(.dina(n9105), .dinb(n9104), .dout(n9106));
  jand g08851(.dina(n9106), .dinb(n9103), .dout(n9107));
  jand g08852(.dina(n9107), .dinb(n9102), .dout(n9108));
  jxor g08853(.dina(n9108), .dinb(a8 ), .dout(n9109));
  jnot g08854(.din(n9109), .dout(n9110));
  jnot g08855(.din(n8851), .dout(n9111));
  jand g08856(.dina(n9075), .dinb(n9111), .dout(n9112));
  jnot g08857(.din(n9112), .dout(n9113));
  jor  g08858(.dina(n9076), .dinb(n8843), .dout(n9114));
  jand g08859(.dina(n9114), .dinb(n9113), .dout(n9115));
  jor  g08860(.dina(n6864), .dinb(n706), .dout(n9116));
  jor  g08861(.dina(n683), .dinb(n6352), .dout(n9117));
  jor  g08862(.dina(n709), .dinb(n6372), .dout(n9118));
  jor  g08863(.dina(n711), .dinb(n6867), .dout(n9119));
  jand g08864(.dina(n9119), .dinb(n9118), .dout(n9120));
  jand g08865(.dina(n9120), .dinb(n9117), .dout(n9121));
  jand g08866(.dina(n9121), .dinb(n9116), .dout(n9122));
  jxor g08867(.dina(n9122), .dinb(a11 ), .dout(n9123));
  jand g08868(.dina(n9073), .dinb(n8864), .dout(n9124));
  jand g08869(.dina(n9074), .dinb(n8855), .dout(n9125));
  jor  g08870(.dina(n9125), .dinb(n9124), .dout(n9126));
  jor  g08871(.dina(n6103), .dinb(n974), .dout(n9127));
  jor  g08872(.dina(n908), .dinb(n5428), .dout(n9128));
  jor  g08873(.dina(n977), .dinb(n5862), .dout(n9129));
  jor  g08874(.dina(n979), .dinb(n6106), .dout(n9130));
  jand g08875(.dina(n9130), .dinb(n9129), .dout(n9131));
  jand g08876(.dina(n9131), .dinb(n9128), .dout(n9132));
  jand g08877(.dina(n9132), .dinb(n9127), .dout(n9133));
  jxor g08878(.dina(n9133), .dinb(a14 ), .dout(n9134));
  jnot g08879(.din(n9134), .dout(n9135));
  jor  g08880(.dina(n9071), .dinb(n9063), .dout(n9136));
  jnot g08881(.din(n9136), .dout(n9137));
  jand g08882(.dina(n9072), .dinb(n8868), .dout(n9138));
  jor  g08883(.dina(n9138), .dinb(n9137), .dout(n9139));
  jor  g08884(.dina(n9061), .dinb(n9053), .dout(n9140));
  jnot g08885(.din(n9140), .dout(n9141));
  jnot g08886(.din(n8869), .dout(n9142));
  jnot g08887(.din(n8546), .dout(n9143));
  jnot g08888(.din(n8003), .dout(n9144));
  jnot g08889(.din(n7711), .dout(n9145));
  jnot g08890(.din(n7438), .dout(n9146));
  jand g08891(.dina(n7356), .dinb(n7198), .dout(n9147));
  jor  g08892(.dina(n9147), .dinb(n9146), .dout(n9148));
  jand g08893(.dina(n7616), .dinb(n9148), .dout(n9149));
  jor  g08894(.dina(n9149), .dinb(n9145), .dout(n9150));
  jand g08895(.dina(n7893), .dinb(n9150), .dout(n9151));
  jor  g08896(.dina(n9151), .dinb(n9144), .dout(n9152));
  jand g08897(.dina(n8181), .dinb(n9152), .dout(n9153));
  jor  g08898(.dina(n9153), .dinb(n8277), .dout(n9154));
  jand g08899(.dina(n8466), .dinb(n9154), .dout(n9155));
  jor  g08900(.dina(n9155), .dinb(n9143), .dout(n9156));
  jand g08901(.dina(n8744), .dinb(n9156), .dout(n9157));
  jor  g08902(.dina(n9157), .dinb(n9142), .dout(n9158));
  jand g08903(.dina(n9062), .dinb(n9158), .dout(n9159));
  jor  g08904(.dina(n9159), .dinb(n9141), .dout(n9160));
  jand g08905(.dina(n9051), .dinb(n8889), .dout(n9161));
  jnot g08906(.din(n8878), .dout(n9162));
  jand g08907(.dina(n8734), .dinb(n8872), .dout(n9163));
  jor  g08908(.dina(n9163), .dinb(n9162), .dout(n9164));
  jand g08909(.dina(n9052), .dinb(n9164), .dout(n9165));
  jor  g08910(.dina(n9165), .dinb(n9161), .dout(n9166));
  jor  g08911(.dina(n9049), .dinb(n9041), .dout(n9167));
  jnot g08912(.din(n9167), .dout(n9168));
  jand g08913(.dina(n9050), .dinb(n8892), .dout(n9169));
  jor  g08914(.dina(n9169), .dinb(n9168), .dout(n9170));
  jand g08915(.dina(n9038), .dinb(n8904), .dout(n9171));
  jand g08916(.dina(n9039), .dinb(n8895), .dout(n9172));
  jor  g08917(.dina(n9172), .dinb(n9171), .dout(n9173));
  jor  g08918(.dina(n3032), .dinb(n2784), .dout(n9174));
  jor  g08919(.dina(n2661), .dinb(n2579), .dout(n9175));
  jor  g08920(.dina(n2787), .dinb(n2870), .dout(n9176));
  jor  g08921(.dina(n2789), .dinb(n3035), .dout(n9177));
  jand g08922(.dina(n9177), .dinb(n9176), .dout(n9178));
  jand g08923(.dina(n9178), .dinb(n9175), .dout(n9179));
  jand g08924(.dina(n9179), .dinb(n9174), .dout(n9180));
  jxor g08925(.dina(n9180), .dinb(a29 ), .dout(n9181));
  jnot g08926(.din(n9181), .dout(n9182));
  jor  g08927(.dina(n9036), .dinb(n9028), .dout(n9183));
  jand g08928(.dina(n9037), .dinb(n8909), .dout(n9184));
  jnot g08929(.din(n9184), .dout(n9185));
  jand g08930(.dina(n9185), .dinb(n9183), .dout(n9186));
  jnot g08931(.din(n9186), .dout(n9187));
  jor  g08932(.dina(n9025), .dinb(n9017), .dout(n9188));
  jand g08933(.dina(n9026), .dinb(n8912), .dout(n9189));
  jnot g08934(.din(n9189), .dout(n9190));
  jand g08935(.dina(n9190), .dinb(n9188), .dout(n9191));
  jnot g08936(.din(n9191), .dout(n9192));
  jand g08937(.dina(n9014), .dinb(n8924), .dout(n9193));
  jand g08938(.dina(n9015), .dinb(n8915), .dout(n9194));
  jor  g08939(.dina(n9194), .dinb(n9193), .dout(n9195));
  jand g08940(.dina(n9012), .dinb(n8936), .dout(n9196));
  jand g08941(.dina(n9013), .dinb(n8927), .dout(n9197));
  jor  g08942(.dina(n9197), .dinb(n9196), .dout(n9198));
  jand g08943(.dina(n9010), .dinb(n8950), .dout(n9199));
  jand g08944(.dina(n9011), .dinb(n8941), .dout(n9200));
  jor  g08945(.dina(n9200), .dinb(n9199), .dout(n9201));
  jand g08946(.dina(n9008), .dinb(n8962), .dout(n9202));
  jand g08947(.dina(n9009), .dinb(n8953), .dout(n9203));
  jor  g08948(.dina(n9203), .dinb(n9202), .dout(n9204));
  jand g08949(.dina(n9006), .dinb(n8974), .dout(n9205));
  jand g08950(.dina(n9007), .dinb(n8965), .dout(n9206));
  jor  g08951(.dina(n9206), .dinb(n9205), .dout(n9207));
  jor  g08952(.dina(n9004), .dinb(n8996), .dout(n9208));
  jand g08953(.dina(n9005), .dinb(n8977), .dout(n9209));
  jnot g08954(.din(n9209), .dout(n9210));
  jand g08955(.dina(n9210), .dinb(n9208), .dout(n9211));
  jnot g08956(.din(n9211), .dout(n9212));
  jor  g08957(.dina(n8125), .dinb(n428), .dout(n9213));
  jor  g08958(.dina(n7846), .dinb(n357), .dout(n9214));
  jor  g08959(.dina(n8128), .dinb(n395), .dout(n9215));
  jor  g08960(.dina(n8130), .dinb(n431), .dout(n9216));
  jand g08961(.dina(n9216), .dinb(n9215), .dout(n9217));
  jand g08962(.dina(n9217), .dinb(n9214), .dout(n9218));
  jand g08963(.dina(n9218), .dinb(n9213), .dout(n9219));
  jxor g08964(.dina(n9219), .dinb(a53 ), .dout(n9220));
  jnot g08965(.din(n9220), .dout(n9221));
  jnot g08966(.din(n8993), .dout(n9222));
  jand g08967(.dina(n9222), .dinb(n8991), .dout(n9223));
  jand g08968(.dina(n8994), .dinb(n8989), .dout(n9224));
  jor  g08969(.dina(n9224), .dinb(n9223), .dout(n9225));
  jor  g08970(.dina(n8978), .dinb(n319), .dout(n9226));
  jor  g08971(.dina(n8677), .dinb(n279), .dout(n9227));
  jor  g08972(.dina(n8981), .dinb(n299), .dout(n9228));
  jor  g08973(.dina(n8983), .dinb(n322), .dout(n9229));
  jand g08974(.dina(n9229), .dinb(n9228), .dout(n9230));
  jand g08975(.dina(n9230), .dinb(n9227), .dout(n9231));
  jand g08976(.dina(n9231), .dinb(n9226), .dout(n9232));
  jxor g08977(.dina(n9232), .dinb(a56 ), .dout(n9233));
  jnot g08978(.din(n9233), .dout(n9234));
  jand g08979(.dina(n8991), .dinb(a59 ), .dout(n9235));
  jxor g08980(.dina(a59 ), .dinb(a58 ), .dout(n9236));
  jnot g08981(.din(n9236), .dout(n9237));
  jand g08982(.dina(n9237), .dinb(n8990), .dout(n9238));
  jand g08983(.dina(n9238), .dinb(b1 ), .dout(n9239));
  jnot g08984(.din(n8990), .dout(n9240));
  jxor g08985(.dina(a58 ), .dinb(a57 ), .dout(n9241));
  jand g08986(.dina(n9241), .dinb(n9240), .dout(n9242));
  jand g08987(.dina(n9242), .dinb(b0 ), .dout(n9243));
  jand g08988(.dina(n9236), .dinb(n8990), .dout(n9244));
  jand g08989(.dina(n9244), .dinb(n338), .dout(n9245));
  jor  g08990(.dina(n9245), .dinb(n9243), .dout(n9246));
  jor  g08991(.dina(n9246), .dinb(n9239), .dout(n9247));
  jxor g08992(.dina(n9247), .dinb(n9235), .dout(n9248));
  jxor g08993(.dina(n9248), .dinb(n9234), .dout(n9249));
  jxor g08994(.dina(n9249), .dinb(n9225), .dout(n9250));
  jxor g08995(.dina(n9250), .dinb(n9221), .dout(n9251));
  jxor g08996(.dina(n9251), .dinb(n9212), .dout(n9252));
  jnot g08997(.din(n9252), .dout(n9253));
  jor  g08998(.dina(n7266), .dinb(n624), .dout(n9254));
  jor  g08999(.dina(n7021), .dinb(n512), .dout(n9255));
  jor  g09000(.dina(n7269), .dinb(n564), .dout(n9256));
  jor  g09001(.dina(n7271), .dinb(n627), .dout(n9257));
  jand g09002(.dina(n9257), .dinb(n9256), .dout(n9258));
  jand g09003(.dina(n9258), .dinb(n9255), .dout(n9259));
  jand g09004(.dina(n9259), .dinb(n9254), .dout(n9260));
  jxor g09005(.dina(n9260), .dinb(a50 ), .dout(n9261));
  jxor g09006(.dina(n9261), .dinb(n9253), .dout(n9262));
  jxor g09007(.dina(n9262), .dinb(n9207), .dout(n9263));
  jnot g09008(.din(n9263), .dout(n9264));
  jor  g09009(.dina(n6490), .dinb(n775), .dout(n9265));
  jor  g09010(.dina(n6262), .dinb(n647), .dout(n9266));
  jor  g09011(.dina(n6493), .dinb(n758), .dout(n9267));
  jor  g09012(.dina(n6495), .dinb(n778), .dout(n9268));
  jand g09013(.dina(n9268), .dinb(n9267), .dout(n9269));
  jand g09014(.dina(n9269), .dinb(n9266), .dout(n9270));
  jand g09015(.dina(n9270), .dinb(n9265), .dout(n9271));
  jxor g09016(.dina(n9271), .dinb(a47 ), .dout(n9272));
  jxor g09017(.dina(n9272), .dinb(n9264), .dout(n9273));
  jxor g09018(.dina(n9273), .dinb(n9204), .dout(n9274));
  jnot g09019(.din(n9274), .dout(n9275));
  jor  g09020(.dina(n5739), .dinb(n1019), .dout(n9276));
  jor  g09021(.dina(n5574), .dinb(n858), .dout(n9277));
  jor  g09022(.dina(n5742), .dinb(n939), .dout(n9278));
  jor  g09023(.dina(n5744), .dinb(n1022), .dout(n9279));
  jand g09024(.dina(n9279), .dinb(n9278), .dout(n9280));
  jand g09025(.dina(n9280), .dinb(n9277), .dout(n9281));
  jand g09026(.dina(n9281), .dinb(n9276), .dout(n9282));
  jxor g09027(.dina(n9282), .dinb(a44 ), .dout(n9283));
  jxor g09028(.dina(n9283), .dinb(n9275), .dout(n9284));
  jxor g09029(.dina(n9284), .dinb(n9201), .dout(n9285));
  jnot g09030(.din(n9285), .dout(n9286));
  jor  g09031(.dina(n5096), .dinb(n1397), .dout(n9287));
  jor  g09032(.dina(n4904), .dinb(n1193), .dout(n9288));
  jor  g09033(.dina(n5099), .dinb(n1290), .dout(n9289));
  jor  g09034(.dina(n5101), .dinb(n1400), .dout(n9290));
  jand g09035(.dina(n9290), .dinb(n9289), .dout(n9291));
  jand g09036(.dina(n9291), .dinb(n9288), .dout(n9292));
  jand g09037(.dina(n9292), .dinb(n9287), .dout(n9293));
  jxor g09038(.dina(n9293), .dinb(a41 ), .dout(n9294));
  jxor g09039(.dina(n9294), .dinb(n9286), .dout(n9295));
  jxor g09040(.dina(n9295), .dinb(n9198), .dout(n9296));
  jnot g09041(.din(n9296), .dout(n9297));
  jor  g09042(.dina(n4415), .dinb(n1739), .dout(n9298));
  jor  g09043(.dina(n4272), .dinb(n1420), .dout(n9299));
  jor  g09044(.dina(n4418), .dinb(n1620), .dout(n9300));
  jor  g09045(.dina(n4420), .dinb(n1742), .dout(n9301));
  jand g09046(.dina(n9301), .dinb(n9300), .dout(n9302));
  jand g09047(.dina(n9302), .dinb(n9299), .dout(n9303));
  jand g09048(.dina(n9303), .dinb(n9298), .dout(n9304));
  jxor g09049(.dina(n9304), .dinb(a38 ), .dout(n9305));
  jxor g09050(.dina(n9305), .dinb(n9297), .dout(n9306));
  jxor g09051(.dina(n9306), .dinb(n9195), .dout(n9307));
  jnot g09052(.din(n9307), .dout(n9308));
  jor  g09053(.dina(n3849), .dinb(n2007), .dout(n9309));
  jor  g09054(.dina(n3689), .dinb(n1867), .dout(n9310));
  jor  g09055(.dina(n3852), .dinb(n1887), .dout(n9311));
  jor  g09056(.dina(n3854), .dinb(n2010), .dout(n9312));
  jand g09057(.dina(n9312), .dinb(n9311), .dout(n9313));
  jand g09058(.dina(n9313), .dinb(n9310), .dout(n9314));
  jand g09059(.dina(n9314), .dinb(n9309), .dout(n9315));
  jxor g09060(.dina(n9315), .dinb(a35 ), .dout(n9316));
  jxor g09061(.dina(n9316), .dinb(n9308), .dout(n9317));
  jxor g09062(.dina(n9317), .dinb(n9192), .dout(n9318));
  jnot g09063(.din(n9318), .dout(n9319));
  jor  g09064(.dina(n3301), .dinb(n2556), .dout(n9320));
  jor  g09065(.dina(n3136), .dinb(n2148), .dout(n9321));
  jor  g09066(.dina(n3304), .dinb(n2407), .dout(n9322));
  jor  g09067(.dina(n3306), .dinb(n2559), .dout(n9323));
  jand g09068(.dina(n9323), .dinb(n9322), .dout(n9324));
  jand g09069(.dina(n9324), .dinb(n9321), .dout(n9325));
  jand g09070(.dina(n9325), .dinb(n9320), .dout(n9326));
  jxor g09071(.dina(n9326), .dinb(a32 ), .dout(n9327));
  jxor g09072(.dina(n9327), .dinb(n9319), .dout(n9328));
  jxor g09073(.dina(n9328), .dinb(n9187), .dout(n9329));
  jxor g09074(.dina(n9329), .dinb(n9182), .dout(n9330));
  jxor g09075(.dina(n9330), .dinb(n9173), .dout(n9331));
  jnot g09076(.din(n9331), .dout(n9332));
  jor  g09077(.dina(n3400), .dinb(n2319), .dout(n9333));
  jor  g09078(.dina(n2224), .dinb(n3055), .dout(n9334));
  jor  g09079(.dina(n2322), .dinb(n3230), .dout(n9335));
  jor  g09080(.dina(n2324), .dinb(n3403), .dout(n9336));
  jand g09081(.dina(n9336), .dinb(n9335), .dout(n9337));
  jand g09082(.dina(n9337), .dinb(n9334), .dout(n9338));
  jand g09083(.dina(n9338), .dinb(n9333), .dout(n9339));
  jxor g09084(.dina(n9339), .dinb(a26 ), .dout(n9340));
  jxor g09085(.dina(n9340), .dinb(n9332), .dout(n9341));
  jxor g09086(.dina(n9341), .dinb(n9170), .dout(n9342));
  jor  g09087(.dina(n4137), .dinb(n1939), .dout(n9343));
  jor  g09088(.dina(n1827), .dinb(n3588), .dout(n9344));
  jor  g09089(.dina(n1942), .dinb(n3942), .dout(n9345));
  jor  g09090(.dina(n1944), .dinb(n4140), .dout(n9346));
  jand g09091(.dina(n9346), .dinb(n9345), .dout(n9347));
  jand g09092(.dina(n9347), .dinb(n9344), .dout(n9348));
  jand g09093(.dina(n9348), .dinb(n9343), .dout(n9349));
  jxor g09094(.dina(n9349), .dinb(a23 ), .dout(n9350));
  jxor g09095(.dina(n9350), .dinb(n9342), .dout(n9351));
  jnot g09096(.din(n9351), .dout(n9352));
  jxor g09097(.dina(n9352), .dinb(n9166), .dout(n9353));
  jor  g09098(.dina(n4554), .dinb(n1566), .dout(n9354));
  jor  g09099(.dina(n1489), .dinb(n4340), .dout(n9355));
  jor  g09100(.dina(n1569), .dinb(n4537), .dout(n9356));
  jor  g09101(.dina(n1571), .dinb(n4557), .dout(n9357));
  jand g09102(.dina(n9357), .dinb(n9356), .dout(n9358));
  jand g09103(.dina(n9358), .dinb(n9355), .dout(n9359));
  jand g09104(.dina(n9359), .dinb(n9354), .dout(n9360));
  jxor g09105(.dina(n9360), .dinb(a20 ), .dout(n9361));
  jxor g09106(.dina(n9361), .dinb(n9353), .dout(n9362));
  jxor g09107(.dina(n9362), .dinb(n9160), .dout(n9363));
  jor  g09108(.dina(n5405), .dinb(n1245), .dout(n9364));
  jor  g09109(.dina(n1165), .dinb(n4974), .dout(n9365));
  jor  g09110(.dina(n1248), .dinb(n4994), .dout(n9366));
  jor  g09111(.dina(n1250), .dinb(n5408), .dout(n9367));
  jand g09112(.dina(n9367), .dinb(n9366), .dout(n9368));
  jand g09113(.dina(n9368), .dinb(n9365), .dout(n9369));
  jand g09114(.dina(n9369), .dinb(n9364), .dout(n9370));
  jxor g09115(.dina(n9370), .dinb(a17 ), .dout(n9371));
  jxor g09116(.dina(n9371), .dinb(n9363), .dout(n9372));
  jxor g09117(.dina(n9372), .dinb(n9139), .dout(n9373));
  jxor g09118(.dina(n9373), .dinb(n9135), .dout(n9374));
  jxor g09119(.dina(n9374), .dinb(n9126), .dout(n9375));
  jxor g09120(.dina(n9375), .dinb(n9123), .dout(n9376));
  jxor g09121(.dina(n9376), .dinb(n9115), .dout(n9377));
  jxor g09122(.dina(n9377), .dinb(n9110), .dout(n9378));
  jxor g09123(.dina(n9378), .dinb(n9101), .dout(n9379));
  jxor g09124(.dina(n9379), .dinb(n9098), .dout(n9380));
  jxor g09125(.dina(n9380), .dinb(n9089), .dout(n9381));
  jand g09126(.dina(b57 ), .dinb(b56 ), .dout(n9382));
  jand g09127(.dina(n8804), .dinb(n8803), .dout(n9383));
  jor  g09128(.dina(n9383), .dinb(n9382), .dout(n9384));
  jxor g09129(.dina(b58 ), .dinb(b57 ), .dout(n9385));
  jnot g09130(.din(n9385), .dout(n9386));
  jxor g09131(.dina(n9386), .dinb(n9384), .dout(n9387));
  jor  g09132(.dina(n9387), .dinb(n264), .dout(n9388));
  jor  g09133(.dina(n284), .dinb(n8789), .dout(n9389));
  jnot g09134(.din(b58 ), .dout(n9390));
  jor  g09135(.dina(n269), .dinb(n9390), .dout(n9391));
  jor  g09136(.dina(n271), .dinb(n8809), .dout(n9392));
  jand g09137(.dina(n9392), .dinb(n9391), .dout(n9393));
  jand g09138(.dina(n9393), .dinb(n9389), .dout(n9394));
  jand g09139(.dina(n9394), .dinb(n9388), .dout(n9395));
  jxor g09140(.dina(n9395), .dinb(n260), .dout(n9396));
  jxor g09141(.dina(n9396), .dinb(n9381), .dout(n9397));
  jxor g09142(.dina(n9397), .dinb(n9086), .dout(f58 ));
  jand g09143(.dina(n9396), .dinb(n9381), .dout(n9399));
  jand g09144(.dina(n9397), .dinb(n9086), .dout(n9400));
  jor  g09145(.dina(n9400), .dinb(n9399), .dout(n9401));
  jand g09146(.dina(n9379), .dinb(n9098), .dout(n9402));
  jand g09147(.dina(n9380), .dinb(n9089), .dout(n9403));
  jor  g09148(.dina(n9403), .dinb(n9402), .dout(n9404));
  jand g09149(.dina(b58 ), .dinb(b57 ), .dout(n9405));
  jand g09150(.dina(n9385), .dinb(n9384), .dout(n9406));
  jor  g09151(.dina(n9406), .dinb(n9405), .dout(n9407));
  jxor g09152(.dina(b59 ), .dinb(b58 ), .dout(n9408));
  jnot g09153(.din(n9408), .dout(n9409));
  jxor g09154(.dina(n9409), .dinb(n9407), .dout(n9410));
  jor  g09155(.dina(n9410), .dinb(n264), .dout(n9411));
  jor  g09156(.dina(n284), .dinb(n8809), .dout(n9412));
  jnot g09157(.din(b59 ), .dout(n9413));
  jor  g09158(.dina(n269), .dinb(n9413), .dout(n9414));
  jor  g09159(.dina(n271), .dinb(n9390), .dout(n9415));
  jand g09160(.dina(n9415), .dinb(n9414), .dout(n9416));
  jand g09161(.dina(n9416), .dinb(n9412), .dout(n9417));
  jand g09162(.dina(n9417), .dinb(n9411), .dout(n9418));
  jxor g09163(.dina(n9418), .dinb(n260), .dout(n9419));
  jor  g09164(.dina(n8786), .dinb(n402), .dout(n9420));
  jor  g09165(.dina(n371), .dinb(n7960), .dout(n9421));
  jor  g09166(.dina(n405), .dinb(n8231), .dout(n9422));
  jor  g09167(.dina(n332), .dinb(n8789), .dout(n9423));
  jand g09168(.dina(n9423), .dinb(n9422), .dout(n9424));
  jand g09169(.dina(n9424), .dinb(n9421), .dout(n9425));
  jand g09170(.dina(n9425), .dinb(n9420), .dout(n9426));
  jxor g09171(.dina(n9426), .dinb(a5 ), .dout(n9427));
  jnot g09172(.din(n9427), .dout(n9428));
  jand g09173(.dina(n9377), .dinb(n9110), .dout(n9429));
  jand g09174(.dina(n9378), .dinb(n9101), .dout(n9430));
  jor  g09175(.dina(n9430), .dinb(n9429), .dout(n9431));
  jor  g09176(.dina(n7680), .dinb(n528), .dout(n9432));
  jor  g09177(.dina(n490), .dinb(n7149), .dout(n9433));
  jor  g09178(.dina(n531), .dinb(n7411), .dout(n9434));
  jor  g09179(.dina(n533), .dinb(n7683), .dout(n9435));
  jand g09180(.dina(n9435), .dinb(n9434), .dout(n9436));
  jand g09181(.dina(n9436), .dinb(n9433), .dout(n9437));
  jand g09182(.dina(n9437), .dinb(n9432), .dout(n9438));
  jxor g09183(.dina(n9438), .dinb(a8 ), .dout(n9439));
  jnot g09184(.din(n9439), .dout(n9440));
  jnot g09185(.din(n9123), .dout(n9441));
  jand g09186(.dina(n9375), .dinb(n9441), .dout(n9442));
  jnot g09187(.din(n9442), .dout(n9443));
  jor  g09188(.dina(n9376), .dinb(n9115), .dout(n9444));
  jand g09189(.dina(n9444), .dinb(n9443), .dout(n9445));
  jand g09190(.dina(n9373), .dinb(n9135), .dout(n9446));
  jand g09191(.dina(n9374), .dinb(n9126), .dout(n9447));
  jor  g09192(.dina(n9447), .dinb(n9446), .dout(n9448));
  jor  g09193(.dina(n6349), .dinb(n974), .dout(n9449));
  jor  g09194(.dina(n908), .dinb(n5862), .dout(n9450));
  jor  g09195(.dina(n977), .dinb(n6106), .dout(n9451));
  jor  g09196(.dina(n979), .dinb(n6352), .dout(n9452));
  jand g09197(.dina(n9452), .dinb(n9451), .dout(n9453));
  jand g09198(.dina(n9453), .dinb(n9450), .dout(n9454));
  jand g09199(.dina(n9454), .dinb(n9449), .dout(n9455));
  jxor g09200(.dina(n9455), .dinb(a14 ), .dout(n9456));
  jnot g09201(.din(n9456), .dout(n9457));
  jor  g09202(.dina(n9371), .dinb(n9363), .dout(n9458));
  jnot g09203(.din(n9458), .dout(n9459));
  jand g09204(.dina(n9372), .dinb(n9139), .dout(n9460));
  jor  g09205(.dina(n9460), .dinb(n9459), .dout(n9461));
  jnot g09206(.din(n9161), .dout(n9462));
  jnot g09207(.din(n9052), .dout(n9463));
  jor  g09208(.dina(n9463), .dinb(n8880), .dout(n9464));
  jand g09209(.dina(n9464), .dinb(n9462), .dout(n9465));
  jxor g09210(.dina(n9352), .dinb(n9465), .dout(n9466));
  jor  g09211(.dina(n9361), .dinb(n9466), .dout(n9467));
  jnot g09212(.din(n9467), .dout(n9468));
  jxor g09213(.dina(n9361), .dinb(n9466), .dout(n9469));
  jand g09214(.dina(n9469), .dinb(n9160), .dout(n9470));
  jor  g09215(.dina(n9470), .dinb(n9468), .dout(n9471));
  jnot g09216(.din(n9342), .dout(n9472));
  jor  g09217(.dina(n9350), .dinb(n9472), .dout(n9473));
  jor  g09218(.dina(n9351), .dinb(n9465), .dout(n9474));
  jand g09219(.dina(n9474), .dinb(n9473), .dout(n9475));
  jor  g09220(.dina(n9340), .dinb(n9332), .dout(n9476));
  jnot g09221(.din(n9476), .dout(n9477));
  jand g09222(.dina(n9341), .dinb(n9170), .dout(n9478));
  jor  g09223(.dina(n9478), .dinb(n9477), .dout(n9479));
  jand g09224(.dina(n9329), .dinb(n9182), .dout(n9480));
  jand g09225(.dina(n9330), .dinb(n9173), .dout(n9481));
  jor  g09226(.dina(n9481), .dinb(n9480), .dout(n9482));
  jor  g09227(.dina(n3052), .dinb(n2784), .dout(n9483));
  jor  g09228(.dina(n2661), .dinb(n2870), .dout(n9484));
  jor  g09229(.dina(n2787), .dinb(n3035), .dout(n9485));
  jor  g09230(.dina(n2789), .dinb(n3055), .dout(n9486));
  jand g09231(.dina(n9486), .dinb(n9485), .dout(n9487));
  jand g09232(.dina(n9487), .dinb(n9484), .dout(n9488));
  jand g09233(.dina(n9488), .dinb(n9483), .dout(n9489));
  jxor g09234(.dina(n9489), .dinb(a29 ), .dout(n9490));
  jnot g09235(.din(n9490), .dout(n9491));
  jor  g09236(.dina(n9327), .dinb(n9319), .dout(n9492));
  jand g09237(.dina(n9328), .dinb(n9187), .dout(n9493));
  jnot g09238(.din(n9493), .dout(n9494));
  jand g09239(.dina(n9494), .dinb(n9492), .dout(n9495));
  jnot g09240(.din(n9495), .dout(n9496));
  jor  g09241(.dina(n9316), .dinb(n9308), .dout(n9497));
  jand g09242(.dina(n9317), .dinb(n9192), .dout(n9498));
  jnot g09243(.din(n9498), .dout(n9499));
  jand g09244(.dina(n9499), .dinb(n9497), .dout(n9500));
  jnot g09245(.din(n9500), .dout(n9501));
  jor  g09246(.dina(n9305), .dinb(n9297), .dout(n9502));
  jand g09247(.dina(n9306), .dinb(n9195), .dout(n9503));
  jnot g09248(.din(n9503), .dout(n9504));
  jand g09249(.dina(n9504), .dinb(n9502), .dout(n9505));
  jnot g09250(.din(n9505), .dout(n9506));
  jor  g09251(.dina(n4415), .dinb(n1864), .dout(n9507));
  jor  g09252(.dina(n4272), .dinb(n1620), .dout(n9508));
  jor  g09253(.dina(n4418), .dinb(n1742), .dout(n9509));
  jor  g09254(.dina(n4420), .dinb(n1867), .dout(n9510));
  jand g09255(.dina(n9510), .dinb(n9509), .dout(n9511));
  jand g09256(.dina(n9511), .dinb(n9508), .dout(n9512));
  jand g09257(.dina(n9512), .dinb(n9507), .dout(n9513));
  jxor g09258(.dina(n9513), .dinb(a38 ), .dout(n9514));
  jnot g09259(.din(n9514), .dout(n9515));
  jor  g09260(.dina(n9294), .dinb(n9286), .dout(n9516));
  jand g09261(.dina(n9295), .dinb(n9198), .dout(n9517));
  jnot g09262(.din(n9517), .dout(n9518));
  jand g09263(.dina(n9518), .dinb(n9516), .dout(n9519));
  jnot g09264(.din(n9519), .dout(n9520));
  jor  g09265(.dina(n5096), .dinb(n1417), .dout(n9521));
  jor  g09266(.dina(n4904), .dinb(n1290), .dout(n9522));
  jor  g09267(.dina(n5099), .dinb(n1400), .dout(n9523));
  jor  g09268(.dina(n5101), .dinb(n1420), .dout(n9524));
  jand g09269(.dina(n9524), .dinb(n9523), .dout(n9525));
  jand g09270(.dina(n9525), .dinb(n9522), .dout(n9526));
  jand g09271(.dina(n9526), .dinb(n9521), .dout(n9527));
  jxor g09272(.dina(n9527), .dinb(a41 ), .dout(n9528));
  jnot g09273(.din(n9528), .dout(n9529));
  jor  g09274(.dina(n9283), .dinb(n9275), .dout(n9530));
  jand g09275(.dina(n9284), .dinb(n9201), .dout(n9531));
  jnot g09276(.din(n9531), .dout(n9532));
  jand g09277(.dina(n9532), .dinb(n9530), .dout(n9533));
  jnot g09278(.din(n9533), .dout(n9534));
  jor  g09279(.dina(n5739), .dinb(n1190), .dout(n9535));
  jor  g09280(.dina(n5574), .dinb(n939), .dout(n9536));
  jor  g09281(.dina(n5742), .dinb(n1022), .dout(n9537));
  jor  g09282(.dina(n5744), .dinb(n1193), .dout(n9538));
  jand g09283(.dina(n9538), .dinb(n9537), .dout(n9539));
  jand g09284(.dina(n9539), .dinb(n9536), .dout(n9540));
  jand g09285(.dina(n9540), .dinb(n9535), .dout(n9541));
  jxor g09286(.dina(n9541), .dinb(a44 ), .dout(n9542));
  jnot g09287(.din(n9542), .dout(n9543));
  jor  g09288(.dina(n9272), .dinb(n9264), .dout(n9544));
  jand g09289(.dina(n9273), .dinb(n9204), .dout(n9545));
  jnot g09290(.din(n9545), .dout(n9546));
  jand g09291(.dina(n9546), .dinb(n9544), .dout(n9547));
  jnot g09292(.din(n9547), .dout(n9548));
  jor  g09293(.dina(n9261), .dinb(n9253), .dout(n9549));
  jand g09294(.dina(n9262), .dinb(n9207), .dout(n9550));
  jnot g09295(.din(n9550), .dout(n9551));
  jand g09296(.dina(n9551), .dinb(n9549), .dout(n9552));
  jnot g09297(.din(n9552), .dout(n9553));
  jor  g09298(.dina(n7266), .dinb(n644), .dout(n9554));
  jor  g09299(.dina(n7021), .dinb(n564), .dout(n9555));
  jor  g09300(.dina(n7269), .dinb(n627), .dout(n9556));
  jor  g09301(.dina(n7271), .dinb(n647), .dout(n9557));
  jand g09302(.dina(n9557), .dinb(n9556), .dout(n9558));
  jand g09303(.dina(n9558), .dinb(n9555), .dout(n9559));
  jand g09304(.dina(n9559), .dinb(n9554), .dout(n9560));
  jxor g09305(.dina(n9560), .dinb(a50 ), .dout(n9561));
  jnot g09306(.din(n9561), .dout(n9562));
  jand g09307(.dina(n9250), .dinb(n9221), .dout(n9563));
  jand g09308(.dina(n9251), .dinb(n9212), .dout(n9564));
  jor  g09309(.dina(n9564), .dinb(n9563), .dout(n9565));
  jor  g09310(.dina(n8125), .dinb(n509), .dout(n9566));
  jor  g09311(.dina(n7846), .dinb(n395), .dout(n9567));
  jor  g09312(.dina(n8128), .dinb(n431), .dout(n9568));
  jor  g09313(.dina(n8130), .dinb(n512), .dout(n9569));
  jand g09314(.dina(n9569), .dinb(n9568), .dout(n9570));
  jand g09315(.dina(n9570), .dinb(n9567), .dout(n9571));
  jand g09316(.dina(n9571), .dinb(n9566), .dout(n9572));
  jxor g09317(.dina(n9572), .dinb(a53 ), .dout(n9573));
  jnot g09318(.din(n9573), .dout(n9574));
  jand g09319(.dina(n9248), .dinb(n9234), .dout(n9575));
  jand g09320(.dina(n9249), .dinb(n9225), .dout(n9576));
  jor  g09321(.dina(n9576), .dinb(n9575), .dout(n9577));
  jor  g09322(.dina(n8978), .dinb(n354), .dout(n9578));
  jor  g09323(.dina(n8677), .dinb(n299), .dout(n9579));
  jor  g09324(.dina(n8981), .dinb(n322), .dout(n9580));
  jor  g09325(.dina(n8983), .dinb(n357), .dout(n9581));
  jand g09326(.dina(n9581), .dinb(n9580), .dout(n9582));
  jand g09327(.dina(n9582), .dinb(n9579), .dout(n9583));
  jand g09328(.dina(n9583), .dinb(n9578), .dout(n9584));
  jxor g09329(.dina(n9584), .dinb(a56 ), .dout(n9585));
  jnot g09330(.din(n9585), .dout(n9586));
  jnot g09331(.din(n9247), .dout(n9587));
  jand g09332(.dina(n8992), .dinb(a59 ), .dout(n9588));
  jand g09333(.dina(n9588), .dinb(n9587), .dout(n9589));
  jnot g09334(.din(n9589), .dout(n9590));
  jand g09335(.dina(n9590), .dinb(a59 ), .dout(n9591));
  jor  g09336(.dina(n9241), .dinb(n9237), .dout(n9592));
  jor  g09337(.dina(n9592), .dinb(n8990), .dout(n9593));
  jnot g09338(.din(n9593), .dout(n9594));
  jand g09339(.dina(n9594), .dinb(b0 ), .dout(n9595));
  jand g09340(.dina(n9238), .dinb(b2 ), .dout(n9596));
  jand g09341(.dina(n9242), .dinb(b1 ), .dout(n9597));
  jand g09342(.dina(n9244), .dinb(n375), .dout(n9598));
  jor  g09343(.dina(n9598), .dinb(n9597), .dout(n9599));
  jor  g09344(.dina(n9599), .dinb(n9596), .dout(n9600));
  jor  g09345(.dina(n9600), .dinb(n9595), .dout(n9601));
  jxor g09346(.dina(n9601), .dinb(n9591), .dout(n9602));
  jxor g09347(.dina(n9602), .dinb(n9586), .dout(n9603));
  jxor g09348(.dina(n9603), .dinb(n9577), .dout(n9604));
  jxor g09349(.dina(n9604), .dinb(n9574), .dout(n9605));
  jxor g09350(.dina(n9605), .dinb(n9565), .dout(n9606));
  jxor g09351(.dina(n9606), .dinb(n9562), .dout(n9607));
  jxor g09352(.dina(n9607), .dinb(n9553), .dout(n9608));
  jnot g09353(.din(n9608), .dout(n9609));
  jor  g09354(.dina(n6490), .dinb(n855), .dout(n9610));
  jor  g09355(.dina(n6262), .dinb(n758), .dout(n9611));
  jor  g09356(.dina(n6493), .dinb(n778), .dout(n9612));
  jor  g09357(.dina(n6495), .dinb(n858), .dout(n9613));
  jand g09358(.dina(n9613), .dinb(n9612), .dout(n9614));
  jand g09359(.dina(n9614), .dinb(n9611), .dout(n9615));
  jand g09360(.dina(n9615), .dinb(n9610), .dout(n9616));
  jxor g09361(.dina(n9616), .dinb(a47 ), .dout(n9617));
  jxor g09362(.dina(n9617), .dinb(n9609), .dout(n9618));
  jxor g09363(.dina(n9618), .dinb(n9548), .dout(n9619));
  jxor g09364(.dina(n9619), .dinb(n9543), .dout(n9620));
  jxor g09365(.dina(n9620), .dinb(n9534), .dout(n9621));
  jxor g09366(.dina(n9621), .dinb(n9529), .dout(n9622));
  jxor g09367(.dina(n9622), .dinb(n9520), .dout(n9623));
  jxor g09368(.dina(n9623), .dinb(n9515), .dout(n9624));
  jxor g09369(.dina(n9624), .dinb(n9506), .dout(n9625));
  jnot g09370(.din(n9625), .dout(n9626));
  jor  g09371(.dina(n3849), .dinb(n2145), .dout(n9627));
  jor  g09372(.dina(n3689), .dinb(n1887), .dout(n9628));
  jor  g09373(.dina(n3852), .dinb(n2010), .dout(n9629));
  jor  g09374(.dina(n3854), .dinb(n2148), .dout(n9630));
  jand g09375(.dina(n9630), .dinb(n9629), .dout(n9631));
  jand g09376(.dina(n9631), .dinb(n9628), .dout(n9632));
  jand g09377(.dina(n9632), .dinb(n9627), .dout(n9633));
  jxor g09378(.dina(n9633), .dinb(a35 ), .dout(n9634));
  jxor g09379(.dina(n9634), .dinb(n9626), .dout(n9635));
  jxor g09380(.dina(n9635), .dinb(n9501), .dout(n9636));
  jnot g09381(.din(n9636), .dout(n9637));
  jor  g09382(.dina(n3301), .dinb(n2576), .dout(n9638));
  jor  g09383(.dina(n3136), .dinb(n2407), .dout(n9639));
  jor  g09384(.dina(n3304), .dinb(n2559), .dout(n9640));
  jor  g09385(.dina(n3306), .dinb(n2579), .dout(n9641));
  jand g09386(.dina(n9641), .dinb(n9640), .dout(n9642));
  jand g09387(.dina(n9642), .dinb(n9639), .dout(n9643));
  jand g09388(.dina(n9643), .dinb(n9638), .dout(n9644));
  jxor g09389(.dina(n9644), .dinb(a32 ), .dout(n9645));
  jxor g09390(.dina(n9645), .dinb(n9637), .dout(n9646));
  jxor g09391(.dina(n9646), .dinb(n9496), .dout(n9647));
  jxor g09392(.dina(n9647), .dinb(n9491), .dout(n9648));
  jxor g09393(.dina(n9648), .dinb(n9482), .dout(n9649));
  jnot g09394(.din(n9649), .dout(n9650));
  jor  g09395(.dina(n3585), .dinb(n2319), .dout(n9651));
  jor  g09396(.dina(n2224), .dinb(n3230), .dout(n9652));
  jor  g09397(.dina(n2322), .dinb(n3403), .dout(n9653));
  jor  g09398(.dina(n2324), .dinb(n3588), .dout(n9654));
  jand g09399(.dina(n9654), .dinb(n9653), .dout(n9655));
  jand g09400(.dina(n9655), .dinb(n9652), .dout(n9656));
  jand g09401(.dina(n9656), .dinb(n9651), .dout(n9657));
  jxor g09402(.dina(n9657), .dinb(a26 ), .dout(n9658));
  jxor g09403(.dina(n9658), .dinb(n9650), .dout(n9659));
  jxor g09404(.dina(n9659), .dinb(n9479), .dout(n9660));
  jor  g09405(.dina(n4337), .dinb(n1939), .dout(n9661));
  jor  g09406(.dina(n1827), .dinb(n3942), .dout(n9662));
  jor  g09407(.dina(n1942), .dinb(n4140), .dout(n9663));
  jor  g09408(.dina(n1944), .dinb(n4340), .dout(n9664));
  jand g09409(.dina(n9664), .dinb(n9663), .dout(n9665));
  jand g09410(.dina(n9665), .dinb(n9662), .dout(n9666));
  jand g09411(.dina(n9666), .dinb(n9661), .dout(n9667));
  jxor g09412(.dina(n9667), .dinb(a23 ), .dout(n9668));
  jxor g09413(.dina(n9668), .dinb(n9660), .dout(n9669));
  jnot g09414(.din(n9669), .dout(n9670));
  jxor g09415(.dina(n9670), .dinb(n9475), .dout(n9671));
  jor  g09416(.dina(n4971), .dinb(n1566), .dout(n9672));
  jor  g09417(.dina(n1489), .dinb(n4537), .dout(n9673));
  jor  g09418(.dina(n1569), .dinb(n4557), .dout(n9674));
  jor  g09419(.dina(n1571), .dinb(n4974), .dout(n9675));
  jand g09420(.dina(n9675), .dinb(n9674), .dout(n9676));
  jand g09421(.dina(n9676), .dinb(n9673), .dout(n9677));
  jand g09422(.dina(n9677), .dinb(n9672), .dout(n9678));
  jxor g09423(.dina(n9678), .dinb(a20 ), .dout(n9679));
  jxor g09424(.dina(n9679), .dinb(n9671), .dout(n9680));
  jxor g09425(.dina(n9680), .dinb(n9471), .dout(n9681));
  jor  g09426(.dina(n5425), .dinb(n1245), .dout(n9682));
  jor  g09427(.dina(n1165), .dinb(n4994), .dout(n9683));
  jor  g09428(.dina(n1248), .dinb(n5408), .dout(n9684));
  jor  g09429(.dina(n1250), .dinb(n5428), .dout(n9685));
  jand g09430(.dina(n9685), .dinb(n9684), .dout(n9686));
  jand g09431(.dina(n9686), .dinb(n9683), .dout(n9687));
  jand g09432(.dina(n9687), .dinb(n9682), .dout(n9688));
  jxor g09433(.dina(n9688), .dinb(a17 ), .dout(n9689));
  jnot g09434(.din(n9689), .dout(n9690));
  jxor g09435(.dina(n9690), .dinb(n9681), .dout(n9691));
  jxor g09436(.dina(n9691), .dinb(n9461), .dout(n9692));
  jxor g09437(.dina(n9692), .dinb(n9457), .dout(n9693));
  jxor g09438(.dina(n9693), .dinb(n9448), .dout(n9694));
  jor  g09439(.dina(n7126), .dinb(n706), .dout(n9695));
  jor  g09440(.dina(n683), .dinb(n6372), .dout(n9696));
  jor  g09441(.dina(n709), .dinb(n6867), .dout(n9697));
  jor  g09442(.dina(n711), .dinb(n7129), .dout(n9698));
  jand g09443(.dina(n9698), .dinb(n9697), .dout(n9699));
  jand g09444(.dina(n9699), .dinb(n9696), .dout(n9700));
  jand g09445(.dina(n9700), .dinb(n9695), .dout(n9701));
  jxor g09446(.dina(n9701), .dinb(a11 ), .dout(n9702));
  jxor g09447(.dina(n9702), .dinb(n9694), .dout(n9703));
  jxor g09448(.dina(n9703), .dinb(n9445), .dout(n9704));
  jxor g09449(.dina(n9704), .dinb(n9440), .dout(n9705));
  jxor g09450(.dina(n9705), .dinb(n9431), .dout(n9706));
  jxor g09451(.dina(n9706), .dinb(n9428), .dout(n9707));
  jxor g09452(.dina(n9707), .dinb(n9419), .dout(n9708));
  jxor g09453(.dina(n9708), .dinb(n9404), .dout(n9709));
  jxor g09454(.dina(n9709), .dinb(n9401), .dout(f59 ));
  jand g09455(.dina(n9708), .dinb(n9404), .dout(n9711));
  jand g09456(.dina(n9709), .dinb(n9401), .dout(n9712));
  jor  g09457(.dina(n9712), .dinb(n9711), .dout(n9713));
  jand g09458(.dina(n9706), .dinb(n9428), .dout(n9714));
  jand g09459(.dina(n9707), .dinb(n9419), .dout(n9715));
  jor  g09460(.dina(n9715), .dinb(n9714), .dout(n9716));
  jand g09461(.dina(b59 ), .dinb(b58 ), .dout(n9717));
  jand g09462(.dina(n9408), .dinb(n9407), .dout(n9718));
  jor  g09463(.dina(n9718), .dinb(n9717), .dout(n9719));
  jxor g09464(.dina(b60 ), .dinb(b59 ), .dout(n9720));
  jnot g09465(.din(n9720), .dout(n9721));
  jxor g09466(.dina(n9721), .dinb(n9719), .dout(n9722));
  jor  g09467(.dina(n9722), .dinb(n264), .dout(n9723));
  jor  g09468(.dina(n284), .dinb(n9390), .dout(n9724));
  jnot g09469(.din(b60 ), .dout(n9725));
  jor  g09470(.dina(n269), .dinb(n9725), .dout(n9726));
  jor  g09471(.dina(n271), .dinb(n9413), .dout(n9727));
  jand g09472(.dina(n9727), .dinb(n9726), .dout(n9728));
  jand g09473(.dina(n9728), .dinb(n9724), .dout(n9729));
  jand g09474(.dina(n9729), .dinb(n9723), .dout(n9730));
  jxor g09475(.dina(n9730), .dinb(n260), .dout(n9731));
  jor  g09476(.dina(n8806), .dinb(n402), .dout(n9732));
  jor  g09477(.dina(n371), .dinb(n8231), .dout(n9733));
  jor  g09478(.dina(n405), .dinb(n8789), .dout(n9734));
  jor  g09479(.dina(n332), .dinb(n8809), .dout(n9735));
  jand g09480(.dina(n9735), .dinb(n9734), .dout(n9736));
  jand g09481(.dina(n9736), .dinb(n9733), .dout(n9737));
  jand g09482(.dina(n9737), .dinb(n9732), .dout(n9738));
  jxor g09483(.dina(n9738), .dinb(a5 ), .dout(n9739));
  jnot g09484(.din(n9739), .dout(n9740));
  jand g09485(.dina(n9704), .dinb(n9440), .dout(n9741));
  jand g09486(.dina(n9705), .dinb(n9431), .dout(n9742));
  jor  g09487(.dina(n9742), .dinb(n9741), .dout(n9743));
  jor  g09488(.dina(n7957), .dinb(n528), .dout(n9744));
  jor  g09489(.dina(n490), .dinb(n7411), .dout(n9745));
  jor  g09490(.dina(n531), .dinb(n7683), .dout(n9746));
  jor  g09491(.dina(n533), .dinb(n7960), .dout(n9747));
  jand g09492(.dina(n9747), .dinb(n9746), .dout(n9748));
  jand g09493(.dina(n9748), .dinb(n9745), .dout(n9749));
  jand g09494(.dina(n9749), .dinb(n9744), .dout(n9750));
  jxor g09495(.dina(n9750), .dinb(a8 ), .dout(n9751));
  jnot g09496(.din(n9751), .dout(n9752));
  jnot g09497(.din(n9694), .dout(n9753));
  jor  g09498(.dina(n9702), .dinb(n9753), .dout(n9754));
  jor  g09499(.dina(n9703), .dinb(n9445), .dout(n9755));
  jand g09500(.dina(n9755), .dinb(n9754), .dout(n9756));
  jor  g09501(.dina(n7146), .dinb(n706), .dout(n9757));
  jor  g09502(.dina(n683), .dinb(n6867), .dout(n9758));
  jor  g09503(.dina(n709), .dinb(n7129), .dout(n9759));
  jor  g09504(.dina(n711), .dinb(n7149), .dout(n9760));
  jand g09505(.dina(n9760), .dinb(n9759), .dout(n9761));
  jand g09506(.dina(n9761), .dinb(n9758), .dout(n9762));
  jand g09507(.dina(n9762), .dinb(n9757), .dout(n9763));
  jxor g09508(.dina(n9763), .dinb(a11 ), .dout(n9764));
  jand g09509(.dina(n9692), .dinb(n9457), .dout(n9765));
  jand g09510(.dina(n9693), .dinb(n9448), .dout(n9766));
  jor  g09511(.dina(n9766), .dinb(n9765), .dout(n9767));
  jor  g09512(.dina(n6369), .dinb(n974), .dout(n9768));
  jor  g09513(.dina(n908), .dinb(n6106), .dout(n9769));
  jor  g09514(.dina(n977), .dinb(n6352), .dout(n9770));
  jor  g09515(.dina(n979), .dinb(n6372), .dout(n9771));
  jand g09516(.dina(n9771), .dinb(n9770), .dout(n9772));
  jand g09517(.dina(n9772), .dinb(n9769), .dout(n9773));
  jand g09518(.dina(n9773), .dinb(n9768), .dout(n9774));
  jxor g09519(.dina(n9774), .dinb(a14 ), .dout(n9775));
  jnot g09520(.din(n9775), .dout(n9776));
  jand g09521(.dina(n9690), .dinb(n9681), .dout(n9777));
  jand g09522(.dina(n9691), .dinb(n9461), .dout(n9778));
  jor  g09523(.dina(n9778), .dinb(n9777), .dout(n9779));
  jor  g09524(.dina(n5859), .dinb(n1245), .dout(n9780));
  jor  g09525(.dina(n1165), .dinb(n5408), .dout(n9781));
  jor  g09526(.dina(n1248), .dinb(n5428), .dout(n9782));
  jor  g09527(.dina(n1250), .dinb(n5862), .dout(n9783));
  jand g09528(.dina(n9783), .dinb(n9782), .dout(n9784));
  jand g09529(.dina(n9784), .dinb(n9781), .dout(n9785));
  jand g09530(.dina(n9785), .dinb(n9780), .dout(n9786));
  jxor g09531(.dina(n9786), .dinb(a17 ), .dout(n9787));
  jnot g09532(.din(n9787), .dout(n9788));
  jor  g09533(.dina(n9679), .dinb(n9671), .dout(n9789));
  jnot g09534(.din(n9789), .dout(n9790));
  jand g09535(.dina(n9680), .dinb(n9471), .dout(n9791));
  jor  g09536(.dina(n9791), .dinb(n9790), .dout(n9792));
  jnot g09537(.din(n9660), .dout(n9793));
  jor  g09538(.dina(n9668), .dinb(n9793), .dout(n9794));
  jor  g09539(.dina(n9669), .dinb(n9475), .dout(n9795));
  jand g09540(.dina(n9795), .dinb(n9794), .dout(n9796));
  jor  g09541(.dina(n9658), .dinb(n9650), .dout(n9797));
  jnot g09542(.din(n9797), .dout(n9798));
  jand g09543(.dina(n9659), .dinb(n9479), .dout(n9799));
  jor  g09544(.dina(n9799), .dinb(n9798), .dout(n9800));
  jor  g09545(.dina(n3939), .dinb(n2319), .dout(n9801));
  jor  g09546(.dina(n2224), .dinb(n3403), .dout(n9802));
  jor  g09547(.dina(n2322), .dinb(n3588), .dout(n9803));
  jor  g09548(.dina(n2324), .dinb(n3942), .dout(n9804));
  jand g09549(.dina(n9804), .dinb(n9803), .dout(n9805));
  jand g09550(.dina(n9805), .dinb(n9802), .dout(n9806));
  jand g09551(.dina(n9806), .dinb(n9801), .dout(n9807));
  jxor g09552(.dina(n9807), .dinb(a26 ), .dout(n9808));
  jnot g09553(.din(n9808), .dout(n9809));
  jand g09554(.dina(n9647), .dinb(n9491), .dout(n9810));
  jand g09555(.dina(n9648), .dinb(n9482), .dout(n9811));
  jor  g09556(.dina(n9811), .dinb(n9810), .dout(n9812));
  jor  g09557(.dina(n9645), .dinb(n9637), .dout(n9813));
  jand g09558(.dina(n9646), .dinb(n9496), .dout(n9814));
  jnot g09559(.din(n9814), .dout(n9815));
  jand g09560(.dina(n9815), .dinb(n9813), .dout(n9816));
  jnot g09561(.din(n9816), .dout(n9817));
  jor  g09562(.dina(n9634), .dinb(n9626), .dout(n9818));
  jand g09563(.dina(n9635), .dinb(n9501), .dout(n9819));
  jnot g09564(.din(n9819), .dout(n9820));
  jand g09565(.dina(n9820), .dinb(n9818), .dout(n9821));
  jnot g09566(.din(n9821), .dout(n9822));
  jand g09567(.dina(n9623), .dinb(n9515), .dout(n9823));
  jand g09568(.dina(n9624), .dinb(n9506), .dout(n9824));
  jor  g09569(.dina(n9824), .dinb(n9823), .dout(n9825));
  jand g09570(.dina(n9621), .dinb(n9529), .dout(n9826));
  jand g09571(.dina(n9622), .dinb(n9520), .dout(n9827));
  jor  g09572(.dina(n9827), .dinb(n9826), .dout(n9828));
  jor  g09573(.dina(n5096), .dinb(n1617), .dout(n9829));
  jor  g09574(.dina(n4904), .dinb(n1400), .dout(n9830));
  jor  g09575(.dina(n5099), .dinb(n1420), .dout(n9831));
  jor  g09576(.dina(n5101), .dinb(n1620), .dout(n9832));
  jand g09577(.dina(n9832), .dinb(n9831), .dout(n9833));
  jand g09578(.dina(n9833), .dinb(n9830), .dout(n9834));
  jand g09579(.dina(n9834), .dinb(n9829), .dout(n9835));
  jxor g09580(.dina(n9835), .dinb(a41 ), .dout(n9836));
  jnot g09581(.din(n9836), .dout(n9837));
  jand g09582(.dina(n9619), .dinb(n9543), .dout(n9838));
  jand g09583(.dina(n9620), .dinb(n9534), .dout(n9839));
  jor  g09584(.dina(n9839), .dinb(n9838), .dout(n9840));
  jor  g09585(.dina(n5739), .dinb(n1287), .dout(n9841));
  jor  g09586(.dina(n5574), .dinb(n1022), .dout(n9842));
  jor  g09587(.dina(n5742), .dinb(n1193), .dout(n9843));
  jor  g09588(.dina(n5744), .dinb(n1290), .dout(n9844));
  jand g09589(.dina(n9844), .dinb(n9843), .dout(n9845));
  jand g09590(.dina(n9845), .dinb(n9842), .dout(n9846));
  jand g09591(.dina(n9846), .dinb(n9841), .dout(n9847));
  jxor g09592(.dina(n9847), .dinb(a44 ), .dout(n9848));
  jnot g09593(.din(n9848), .dout(n9849));
  jor  g09594(.dina(n9617), .dinb(n9609), .dout(n9850));
  jand g09595(.dina(n9618), .dinb(n9548), .dout(n9851));
  jnot g09596(.din(n9851), .dout(n9852));
  jand g09597(.dina(n9852), .dinb(n9850), .dout(n9853));
  jnot g09598(.din(n9853), .dout(n9854));
  jor  g09599(.dina(n6490), .dinb(n936), .dout(n9855));
  jor  g09600(.dina(n6262), .dinb(n778), .dout(n9856));
  jor  g09601(.dina(n6493), .dinb(n858), .dout(n9857));
  jor  g09602(.dina(n6495), .dinb(n939), .dout(n9858));
  jand g09603(.dina(n9858), .dinb(n9857), .dout(n9859));
  jand g09604(.dina(n9859), .dinb(n9856), .dout(n9860));
  jand g09605(.dina(n9860), .dinb(n9855), .dout(n9861));
  jxor g09606(.dina(n9861), .dinb(a47 ), .dout(n9862));
  jnot g09607(.din(n9862), .dout(n9863));
  jand g09608(.dina(n9606), .dinb(n9562), .dout(n9864));
  jand g09609(.dina(n9607), .dinb(n9553), .dout(n9865));
  jor  g09610(.dina(n9865), .dinb(n9864), .dout(n9866));
  jor  g09611(.dina(n7266), .dinb(n755), .dout(n9867));
  jor  g09612(.dina(n7021), .dinb(n627), .dout(n9868));
  jor  g09613(.dina(n7269), .dinb(n647), .dout(n9869));
  jor  g09614(.dina(n7271), .dinb(n758), .dout(n9870));
  jand g09615(.dina(n9870), .dinb(n9869), .dout(n9871));
  jand g09616(.dina(n9871), .dinb(n9868), .dout(n9872));
  jand g09617(.dina(n9872), .dinb(n9867), .dout(n9873));
  jxor g09618(.dina(n9873), .dinb(a50 ), .dout(n9874));
  jnot g09619(.din(n9874), .dout(n9875));
  jand g09620(.dina(n9604), .dinb(n9574), .dout(n9876));
  jand g09621(.dina(n9605), .dinb(n9565), .dout(n9877));
  jor  g09622(.dina(n9877), .dinb(n9876), .dout(n9878));
  jor  g09623(.dina(n8125), .dinb(n561), .dout(n9879));
  jor  g09624(.dina(n7846), .dinb(n431), .dout(n9880));
  jor  g09625(.dina(n8128), .dinb(n512), .dout(n9881));
  jor  g09626(.dina(n8130), .dinb(n564), .dout(n9882));
  jand g09627(.dina(n9882), .dinb(n9881), .dout(n9883));
  jand g09628(.dina(n9883), .dinb(n9880), .dout(n9884));
  jand g09629(.dina(n9884), .dinb(n9879), .dout(n9885));
  jxor g09630(.dina(n9885), .dinb(a53 ), .dout(n9886));
  jnot g09631(.din(n9886), .dout(n9887));
  jand g09632(.dina(n9602), .dinb(n9586), .dout(n9888));
  jand g09633(.dina(n9603), .dinb(n9577), .dout(n9889));
  jor  g09634(.dina(n9889), .dinb(n9888), .dout(n9890));
  jnot g09635(.din(n9244), .dout(n9891));
  jor  g09636(.dina(n9891), .dinb(n296), .dout(n9892));
  jor  g09637(.dina(n9593), .dinb(n267), .dout(n9893));
  jnot g09638(.din(n9242), .dout(n9894));
  jor  g09639(.dina(n9894), .dinb(n279), .dout(n9895));
  jnot g09640(.din(n9238), .dout(n9896));
  jor  g09641(.dina(n9896), .dinb(n299), .dout(n9897));
  jand g09642(.dina(n9897), .dinb(n9895), .dout(n9898));
  jand g09643(.dina(n9898), .dinb(n9893), .dout(n9899));
  jand g09644(.dina(n9899), .dinb(n9892), .dout(n9900));
  jxor g09645(.dina(n9900), .dinb(a59 ), .dout(n9901));
  jnot g09646(.din(n9901), .dout(n9902));
  jxor g09647(.dina(a60 ), .dinb(a59 ), .dout(n9903));
  jand g09648(.dina(n9903), .dinb(b0 ), .dout(n9904));
  jnot g09649(.din(n9904), .dout(n9905));
  jor  g09650(.dina(n9601), .dinb(n9590), .dout(n9906));
  jxor g09651(.dina(n9906), .dinb(n9905), .dout(n9907));
  jxor g09652(.dina(n9907), .dinb(n9902), .dout(n9908));
  jnot g09653(.din(n9908), .dout(n9909));
  jor  g09654(.dina(n8978), .dinb(n392), .dout(n9910));
  jor  g09655(.dina(n8677), .dinb(n322), .dout(n9911));
  jor  g09656(.dina(n8981), .dinb(n357), .dout(n9912));
  jor  g09657(.dina(n8983), .dinb(n395), .dout(n9913));
  jand g09658(.dina(n9913), .dinb(n9912), .dout(n9914));
  jand g09659(.dina(n9914), .dinb(n9911), .dout(n9915));
  jand g09660(.dina(n9915), .dinb(n9910), .dout(n9916));
  jxor g09661(.dina(n9916), .dinb(a56 ), .dout(n9917));
  jxor g09662(.dina(n9917), .dinb(n9909), .dout(n9918));
  jxor g09663(.dina(n9918), .dinb(n9890), .dout(n9919));
  jxor g09664(.dina(n9919), .dinb(n9887), .dout(n9920));
  jxor g09665(.dina(n9920), .dinb(n9878), .dout(n9921));
  jxor g09666(.dina(n9921), .dinb(n9875), .dout(n9922));
  jxor g09667(.dina(n9922), .dinb(n9866), .dout(n9923));
  jxor g09668(.dina(n9923), .dinb(n9863), .dout(n9924));
  jxor g09669(.dina(n9924), .dinb(n9854), .dout(n9925));
  jxor g09670(.dina(n9925), .dinb(n9849), .dout(n9926));
  jxor g09671(.dina(n9926), .dinb(n9840), .dout(n9927));
  jxor g09672(.dina(n9927), .dinb(n9837), .dout(n9928));
  jxor g09673(.dina(n9928), .dinb(n9828), .dout(n9929));
  jnot g09674(.din(n9929), .dout(n9930));
  jor  g09675(.dina(n4415), .dinb(n1884), .dout(n9931));
  jor  g09676(.dina(n4272), .dinb(n1742), .dout(n9932));
  jor  g09677(.dina(n4418), .dinb(n1867), .dout(n9933));
  jor  g09678(.dina(n4420), .dinb(n1887), .dout(n9934));
  jand g09679(.dina(n9934), .dinb(n9933), .dout(n9935));
  jand g09680(.dina(n9935), .dinb(n9932), .dout(n9936));
  jand g09681(.dina(n9936), .dinb(n9931), .dout(n9937));
  jxor g09682(.dina(n9937), .dinb(a38 ), .dout(n9938));
  jxor g09683(.dina(n9938), .dinb(n9930), .dout(n9939));
  jxor g09684(.dina(n9939), .dinb(n9825), .dout(n9940));
  jnot g09685(.din(n9940), .dout(n9941));
  jor  g09686(.dina(n3849), .dinb(n2404), .dout(n9942));
  jor  g09687(.dina(n3689), .dinb(n2010), .dout(n9943));
  jor  g09688(.dina(n3852), .dinb(n2148), .dout(n9944));
  jor  g09689(.dina(n3854), .dinb(n2407), .dout(n9945));
  jand g09690(.dina(n9945), .dinb(n9944), .dout(n9946));
  jand g09691(.dina(n9946), .dinb(n9943), .dout(n9947));
  jand g09692(.dina(n9947), .dinb(n9942), .dout(n9948));
  jxor g09693(.dina(n9948), .dinb(a35 ), .dout(n9949));
  jxor g09694(.dina(n9949), .dinb(n9941), .dout(n9950));
  jxor g09695(.dina(n9950), .dinb(n9822), .dout(n9951));
  jnot g09696(.din(n9951), .dout(n9952));
  jor  g09697(.dina(n3301), .dinb(n2867), .dout(n9953));
  jor  g09698(.dina(n3136), .dinb(n2559), .dout(n9954));
  jor  g09699(.dina(n3304), .dinb(n2579), .dout(n9955));
  jor  g09700(.dina(n3306), .dinb(n2870), .dout(n9956));
  jand g09701(.dina(n9956), .dinb(n9955), .dout(n9957));
  jand g09702(.dina(n9957), .dinb(n9954), .dout(n9958));
  jand g09703(.dina(n9958), .dinb(n9953), .dout(n9959));
  jxor g09704(.dina(n9959), .dinb(a32 ), .dout(n9960));
  jxor g09705(.dina(n9960), .dinb(n9952), .dout(n9961));
  jxor g09706(.dina(n9961), .dinb(n9817), .dout(n9962));
  jnot g09707(.din(n9962), .dout(n9963));
  jor  g09708(.dina(n3227), .dinb(n2784), .dout(n9964));
  jor  g09709(.dina(n2661), .dinb(n3035), .dout(n9965));
  jor  g09710(.dina(n2787), .dinb(n3055), .dout(n9966));
  jor  g09711(.dina(n2789), .dinb(n3230), .dout(n9967));
  jand g09712(.dina(n9967), .dinb(n9966), .dout(n9968));
  jand g09713(.dina(n9968), .dinb(n9965), .dout(n9969));
  jand g09714(.dina(n9969), .dinb(n9964), .dout(n9970));
  jxor g09715(.dina(n9970), .dinb(a29 ), .dout(n9971));
  jxor g09716(.dina(n9971), .dinb(n9963), .dout(n9972));
  jxor g09717(.dina(n9972), .dinb(n9812), .dout(n9973));
  jxor g09718(.dina(n9973), .dinb(n9809), .dout(n9974));
  jxor g09719(.dina(n9974), .dinb(n9800), .dout(n9975));
  jor  g09720(.dina(n4534), .dinb(n1939), .dout(n9976));
  jor  g09721(.dina(n1827), .dinb(n4140), .dout(n9977));
  jor  g09722(.dina(n1942), .dinb(n4340), .dout(n9978));
  jor  g09723(.dina(n1944), .dinb(n4537), .dout(n9979));
  jand g09724(.dina(n9979), .dinb(n9978), .dout(n9980));
  jand g09725(.dina(n9980), .dinb(n9977), .dout(n9981));
  jand g09726(.dina(n9981), .dinb(n9976), .dout(n9982));
  jxor g09727(.dina(n9982), .dinb(a23 ), .dout(n9983));
  jxor g09728(.dina(n9983), .dinb(n9975), .dout(n9984));
  jnot g09729(.din(n9984), .dout(n9985));
  jxor g09730(.dina(n9985), .dinb(n9796), .dout(n9986));
  jor  g09731(.dina(n4991), .dinb(n1566), .dout(n9987));
  jor  g09732(.dina(n1489), .dinb(n4557), .dout(n9988));
  jor  g09733(.dina(n1569), .dinb(n4974), .dout(n9989));
  jor  g09734(.dina(n1571), .dinb(n4994), .dout(n9990));
  jand g09735(.dina(n9990), .dinb(n9989), .dout(n9991));
  jand g09736(.dina(n9991), .dinb(n9988), .dout(n9992));
  jand g09737(.dina(n9992), .dinb(n9987), .dout(n9993));
  jxor g09738(.dina(n9993), .dinb(a20 ), .dout(n9994));
  jxor g09739(.dina(n9994), .dinb(n9986), .dout(n9995));
  jxor g09740(.dina(n9995), .dinb(n9792), .dout(n9996));
  jxor g09741(.dina(n9996), .dinb(n9788), .dout(n9997));
  jxor g09742(.dina(n9997), .dinb(n9779), .dout(n9998));
  jxor g09743(.dina(n9998), .dinb(n9776), .dout(n9999));
  jxor g09744(.dina(n9999), .dinb(n9767), .dout(n10000));
  jxor g09745(.dina(n10000), .dinb(n9764), .dout(n10001));
  jxor g09746(.dina(n10001), .dinb(n9756), .dout(n10002));
  jxor g09747(.dina(n10002), .dinb(n9752), .dout(n10003));
  jxor g09748(.dina(n10003), .dinb(n9743), .dout(n10004));
  jxor g09749(.dina(n10004), .dinb(n9740), .dout(n10005));
  jxor g09750(.dina(n10005), .dinb(n9731), .dout(n10006));
  jxor g09751(.dina(n10006), .dinb(n9716), .dout(n10007));
  jxor g09752(.dina(n10007), .dinb(n9713), .dout(f60 ));
  jand g09753(.dina(n10004), .dinb(n9740), .dout(n10009));
  jand g09754(.dina(n10005), .dinb(n9731), .dout(n10010));
  jor  g09755(.dina(n10010), .dinb(n10009), .dout(n10011));
  jand g09756(.dina(n10002), .dinb(n9752), .dout(n10012));
  jand g09757(.dina(n10003), .dinb(n9743), .dout(n10013));
  jor  g09758(.dina(n10013), .dinb(n10012), .dout(n10014));
  jnot g09759(.din(n9764), .dout(n10015));
  jand g09760(.dina(n10000), .dinb(n10015), .dout(n10016));
  jnot g09761(.din(n10016), .dout(n10017));
  jor  g09762(.dina(n10001), .dinb(n9756), .dout(n10018));
  jand g09763(.dina(n10018), .dinb(n10017), .dout(n10019));
  jor  g09764(.dina(n7408), .dinb(n706), .dout(n10020));
  jor  g09765(.dina(n683), .dinb(n7129), .dout(n10021));
  jor  g09766(.dina(n709), .dinb(n7149), .dout(n10022));
  jor  g09767(.dina(n711), .dinb(n7411), .dout(n10023));
  jand g09768(.dina(n10023), .dinb(n10022), .dout(n10024));
  jand g09769(.dina(n10024), .dinb(n10021), .dout(n10025));
  jand g09770(.dina(n10025), .dinb(n10020), .dout(n10026));
  jxor g09771(.dina(n10026), .dinb(a11 ), .dout(n10027));
  jand g09772(.dina(n9998), .dinb(n9776), .dout(n10028));
  jand g09773(.dina(n9999), .dinb(n9767), .dout(n10029));
  jor  g09774(.dina(n10029), .dinb(n10028), .dout(n10030));
  jor  g09775(.dina(n6864), .dinb(n974), .dout(n10031));
  jor  g09776(.dina(n908), .dinb(n6352), .dout(n10032));
  jor  g09777(.dina(n977), .dinb(n6372), .dout(n10033));
  jor  g09778(.dina(n979), .dinb(n6867), .dout(n10034));
  jand g09779(.dina(n10034), .dinb(n10033), .dout(n10035));
  jand g09780(.dina(n10035), .dinb(n10032), .dout(n10036));
  jand g09781(.dina(n10036), .dinb(n10031), .dout(n10037));
  jxor g09782(.dina(n10037), .dinb(a14 ), .dout(n10038));
  jnot g09783(.din(n10038), .dout(n10039));
  jand g09784(.dina(n9996), .dinb(n9788), .dout(n10040));
  jand g09785(.dina(n9997), .dinb(n9779), .dout(n10041));
  jor  g09786(.dina(n10041), .dinb(n10040), .dout(n10042));
  jor  g09787(.dina(n6103), .dinb(n1245), .dout(n10043));
  jor  g09788(.dina(n1165), .dinb(n5428), .dout(n10044));
  jor  g09789(.dina(n1248), .dinb(n5862), .dout(n10045));
  jor  g09790(.dina(n1250), .dinb(n6106), .dout(n10046));
  jand g09791(.dina(n10046), .dinb(n10045), .dout(n10047));
  jand g09792(.dina(n10047), .dinb(n10044), .dout(n10048));
  jand g09793(.dina(n10048), .dinb(n10043), .dout(n10049));
  jxor g09794(.dina(n10049), .dinb(a17 ), .dout(n10050));
  jnot g09795(.din(n10050), .dout(n10051));
  jor  g09796(.dina(n9994), .dinb(n9986), .dout(n10052));
  jnot g09797(.din(n10052), .dout(n10053));
  jand g09798(.dina(n9995), .dinb(n9792), .dout(n10054));
  jor  g09799(.dina(n10054), .dinb(n10053), .dout(n10055));
  jnot g09800(.din(n9975), .dout(n10056));
  jor  g09801(.dina(n9983), .dinb(n10056), .dout(n10057));
  jnot g09802(.din(n10057), .dout(n10058));
  jnot g09803(.din(n9794), .dout(n10059));
  jnot g09804(.din(n9473), .dout(n10060));
  jand g09805(.dina(n9352), .dinb(n9166), .dout(n10061));
  jor  g09806(.dina(n10061), .dinb(n10060), .dout(n10062));
  jand g09807(.dina(n9670), .dinb(n10062), .dout(n10063));
  jor  g09808(.dina(n10063), .dinb(n10059), .dout(n10064));
  jand g09809(.dina(n9985), .dinb(n10064), .dout(n10065));
  jor  g09810(.dina(n10065), .dinb(n10058), .dout(n10066));
  jand g09811(.dina(n9973), .dinb(n9809), .dout(n10067));
  jand g09812(.dina(n9974), .dinb(n9800), .dout(n10068));
  jor  g09813(.dina(n10068), .dinb(n10067), .dout(n10069));
  jor  g09814(.dina(n9971), .dinb(n9963), .dout(n10070));
  jand g09815(.dina(n9972), .dinb(n9812), .dout(n10071));
  jnot g09816(.din(n10071), .dout(n10072));
  jand g09817(.dina(n10072), .dinb(n10070), .dout(n10073));
  jnot g09818(.din(n10073), .dout(n10074));
  jor  g09819(.dina(n3400), .dinb(n2784), .dout(n10075));
  jor  g09820(.dina(n2661), .dinb(n3055), .dout(n10076));
  jor  g09821(.dina(n2787), .dinb(n3230), .dout(n10077));
  jor  g09822(.dina(n2789), .dinb(n3403), .dout(n10078));
  jand g09823(.dina(n10078), .dinb(n10077), .dout(n10079));
  jand g09824(.dina(n10079), .dinb(n10076), .dout(n10080));
  jand g09825(.dina(n10080), .dinb(n10075), .dout(n10081));
  jxor g09826(.dina(n10081), .dinb(a29 ), .dout(n10082));
  jnot g09827(.din(n10082), .dout(n10083));
  jor  g09828(.dina(n9960), .dinb(n9952), .dout(n10084));
  jand g09829(.dina(n9961), .dinb(n9817), .dout(n10085));
  jnot g09830(.din(n10085), .dout(n10086));
  jand g09831(.dina(n10086), .dinb(n10084), .dout(n10087));
  jnot g09832(.din(n10087), .dout(n10088));
  jor  g09833(.dina(n9949), .dinb(n9941), .dout(n10089));
  jand g09834(.dina(n9950), .dinb(n9822), .dout(n10090));
  jnot g09835(.din(n10090), .dout(n10091));
  jand g09836(.dina(n10091), .dinb(n10089), .dout(n10092));
  jnot g09837(.din(n10092), .dout(n10093));
  jor  g09838(.dina(n9938), .dinb(n9930), .dout(n10094));
  jand g09839(.dina(n9939), .dinb(n9825), .dout(n10095));
  jnot g09840(.din(n10095), .dout(n10096));
  jand g09841(.dina(n10096), .dinb(n10094), .dout(n10097));
  jnot g09842(.din(n10097), .dout(n10098));
  jand g09843(.dina(n9927), .dinb(n9837), .dout(n10099));
  jand g09844(.dina(n9928), .dinb(n9828), .dout(n10100));
  jor  g09845(.dina(n10100), .dinb(n10099), .dout(n10101));
  jand g09846(.dina(n9925), .dinb(n9849), .dout(n10102));
  jand g09847(.dina(n9926), .dinb(n9840), .dout(n10103));
  jor  g09848(.dina(n10103), .dinb(n10102), .dout(n10104));
  jand g09849(.dina(n9923), .dinb(n9863), .dout(n10105));
  jand g09850(.dina(n9924), .dinb(n9854), .dout(n10106));
  jor  g09851(.dina(n10106), .dinb(n10105), .dout(n10107));
  jand g09852(.dina(n9921), .dinb(n9875), .dout(n10108));
  jand g09853(.dina(n9922), .dinb(n9866), .dout(n10109));
  jor  g09854(.dina(n10109), .dinb(n10108), .dout(n10110));
  jand g09855(.dina(n9919), .dinb(n9887), .dout(n10111));
  jand g09856(.dina(n9920), .dinb(n9878), .dout(n10112));
  jor  g09857(.dina(n10112), .dinb(n10111), .dout(n10113));
  jor  g09858(.dina(n9917), .dinb(n9909), .dout(n10114));
  jand g09859(.dina(n9918), .dinb(n9890), .dout(n10115));
  jnot g09860(.din(n10115), .dout(n10116));
  jand g09861(.dina(n10116), .dinb(n10114), .dout(n10117));
  jnot g09862(.din(n10117), .dout(n10118));
  jor  g09863(.dina(n8978), .dinb(n428), .dout(n10119));
  jor  g09864(.dina(n8677), .dinb(n357), .dout(n10120));
  jor  g09865(.dina(n8981), .dinb(n395), .dout(n10121));
  jor  g09866(.dina(n8983), .dinb(n431), .dout(n10122));
  jand g09867(.dina(n10122), .dinb(n10121), .dout(n10123));
  jand g09868(.dina(n10123), .dinb(n10120), .dout(n10124));
  jand g09869(.dina(n10124), .dinb(n10119), .dout(n10125));
  jxor g09870(.dina(n10125), .dinb(a56 ), .dout(n10126));
  jnot g09871(.din(n10126), .dout(n10127));
  jnot g09872(.din(n9906), .dout(n10128));
  jand g09873(.dina(n10128), .dinb(n9904), .dout(n10129));
  jand g09874(.dina(n9907), .dinb(n9902), .dout(n10130));
  jor  g09875(.dina(n10130), .dinb(n10129), .dout(n10131));
  jor  g09876(.dina(n9891), .dinb(n319), .dout(n10132));
  jor  g09877(.dina(n9593), .dinb(n279), .dout(n10133));
  jor  g09878(.dina(n9894), .dinb(n299), .dout(n10134));
  jor  g09879(.dina(n9896), .dinb(n322), .dout(n10135));
  jand g09880(.dina(n10135), .dinb(n10134), .dout(n10136));
  jand g09881(.dina(n10136), .dinb(n10133), .dout(n10137));
  jand g09882(.dina(n10137), .dinb(n10132), .dout(n10138));
  jxor g09883(.dina(n10138), .dinb(a59 ), .dout(n10139));
  jnot g09884(.din(n10139), .dout(n10140));
  jand g09885(.dina(n9904), .dinb(a62 ), .dout(n10141));
  jxor g09886(.dina(a62 ), .dinb(a61 ), .dout(n10142));
  jnot g09887(.din(n10142), .dout(n10143));
  jand g09888(.dina(n10143), .dinb(n9903), .dout(n10144));
  jand g09889(.dina(n10144), .dinb(b1 ), .dout(n10145));
  jnot g09890(.din(n9903), .dout(n10146));
  jxor g09891(.dina(a61 ), .dinb(a60 ), .dout(n10147));
  jand g09892(.dina(n10147), .dinb(n10146), .dout(n10148));
  jand g09893(.dina(n10148), .dinb(b0 ), .dout(n10149));
  jand g09894(.dina(n10142), .dinb(n9903), .dout(n10150));
  jand g09895(.dina(n10150), .dinb(n338), .dout(n10151));
  jor  g09896(.dina(n10151), .dinb(n10149), .dout(n10152));
  jor  g09897(.dina(n10152), .dinb(n10145), .dout(n10153));
  jxor g09898(.dina(n10153), .dinb(n10141), .dout(n10154));
  jxor g09899(.dina(n10154), .dinb(n10140), .dout(n10155));
  jxor g09900(.dina(n10155), .dinb(n10131), .dout(n10156));
  jxor g09901(.dina(n10156), .dinb(n10127), .dout(n10157));
  jxor g09902(.dina(n10157), .dinb(n10118), .dout(n10158));
  jnot g09903(.din(n10158), .dout(n10159));
  jor  g09904(.dina(n8125), .dinb(n624), .dout(n10160));
  jor  g09905(.dina(n7846), .dinb(n512), .dout(n10161));
  jor  g09906(.dina(n8128), .dinb(n564), .dout(n10162));
  jor  g09907(.dina(n8130), .dinb(n627), .dout(n10163));
  jand g09908(.dina(n10163), .dinb(n10162), .dout(n10164));
  jand g09909(.dina(n10164), .dinb(n10161), .dout(n10165));
  jand g09910(.dina(n10165), .dinb(n10160), .dout(n10166));
  jxor g09911(.dina(n10166), .dinb(a53 ), .dout(n10167));
  jxor g09912(.dina(n10167), .dinb(n10159), .dout(n10168));
  jxor g09913(.dina(n10168), .dinb(n10113), .dout(n10169));
  jnot g09914(.din(n10169), .dout(n10170));
  jor  g09915(.dina(n7266), .dinb(n775), .dout(n10171));
  jor  g09916(.dina(n7021), .dinb(n647), .dout(n10172));
  jor  g09917(.dina(n7269), .dinb(n758), .dout(n10173));
  jor  g09918(.dina(n7271), .dinb(n778), .dout(n10174));
  jand g09919(.dina(n10174), .dinb(n10173), .dout(n10175));
  jand g09920(.dina(n10175), .dinb(n10172), .dout(n10176));
  jand g09921(.dina(n10176), .dinb(n10171), .dout(n10177));
  jxor g09922(.dina(n10177), .dinb(a50 ), .dout(n10178));
  jxor g09923(.dina(n10178), .dinb(n10170), .dout(n10179));
  jxor g09924(.dina(n10179), .dinb(n10110), .dout(n10180));
  jnot g09925(.din(n10180), .dout(n10181));
  jor  g09926(.dina(n6490), .dinb(n1019), .dout(n10182));
  jor  g09927(.dina(n6262), .dinb(n858), .dout(n10183));
  jor  g09928(.dina(n6493), .dinb(n939), .dout(n10184));
  jor  g09929(.dina(n6495), .dinb(n1022), .dout(n10185));
  jand g09930(.dina(n10185), .dinb(n10184), .dout(n10186));
  jand g09931(.dina(n10186), .dinb(n10183), .dout(n10187));
  jand g09932(.dina(n10187), .dinb(n10182), .dout(n10188));
  jxor g09933(.dina(n10188), .dinb(a47 ), .dout(n10189));
  jxor g09934(.dina(n10189), .dinb(n10181), .dout(n10190));
  jxor g09935(.dina(n10190), .dinb(n10107), .dout(n10191));
  jnot g09936(.din(n10191), .dout(n10192));
  jor  g09937(.dina(n5739), .dinb(n1397), .dout(n10193));
  jor  g09938(.dina(n5574), .dinb(n1193), .dout(n10194));
  jor  g09939(.dina(n5742), .dinb(n1290), .dout(n10195));
  jor  g09940(.dina(n5744), .dinb(n1400), .dout(n10196));
  jand g09941(.dina(n10196), .dinb(n10195), .dout(n10197));
  jand g09942(.dina(n10197), .dinb(n10194), .dout(n10198));
  jand g09943(.dina(n10198), .dinb(n10193), .dout(n10199));
  jxor g09944(.dina(n10199), .dinb(a44 ), .dout(n10200));
  jxor g09945(.dina(n10200), .dinb(n10192), .dout(n10201));
  jxor g09946(.dina(n10201), .dinb(n10104), .dout(n10202));
  jnot g09947(.din(n10202), .dout(n10203));
  jor  g09948(.dina(n5096), .dinb(n1739), .dout(n10204));
  jor  g09949(.dina(n4904), .dinb(n1420), .dout(n10205));
  jor  g09950(.dina(n5099), .dinb(n1620), .dout(n10206));
  jor  g09951(.dina(n5101), .dinb(n1742), .dout(n10207));
  jand g09952(.dina(n10207), .dinb(n10206), .dout(n10208));
  jand g09953(.dina(n10208), .dinb(n10205), .dout(n10209));
  jand g09954(.dina(n10209), .dinb(n10204), .dout(n10210));
  jxor g09955(.dina(n10210), .dinb(a41 ), .dout(n10211));
  jxor g09956(.dina(n10211), .dinb(n10203), .dout(n10212));
  jxor g09957(.dina(n10212), .dinb(n10101), .dout(n10213));
  jnot g09958(.din(n10213), .dout(n10214));
  jor  g09959(.dina(n4415), .dinb(n2007), .dout(n10215));
  jor  g09960(.dina(n4272), .dinb(n1867), .dout(n10216));
  jor  g09961(.dina(n4418), .dinb(n1887), .dout(n10217));
  jor  g09962(.dina(n4420), .dinb(n2010), .dout(n10218));
  jand g09963(.dina(n10218), .dinb(n10217), .dout(n10219));
  jand g09964(.dina(n10219), .dinb(n10216), .dout(n10220));
  jand g09965(.dina(n10220), .dinb(n10215), .dout(n10221));
  jxor g09966(.dina(n10221), .dinb(a38 ), .dout(n10222));
  jxor g09967(.dina(n10222), .dinb(n10214), .dout(n10223));
  jxor g09968(.dina(n10223), .dinb(n10098), .dout(n10224));
  jnot g09969(.din(n10224), .dout(n10225));
  jor  g09970(.dina(n3849), .dinb(n2556), .dout(n10226));
  jor  g09971(.dina(n3689), .dinb(n2148), .dout(n10227));
  jor  g09972(.dina(n3852), .dinb(n2407), .dout(n10228));
  jor  g09973(.dina(n3854), .dinb(n2559), .dout(n10229));
  jand g09974(.dina(n10229), .dinb(n10228), .dout(n10230));
  jand g09975(.dina(n10230), .dinb(n10227), .dout(n10231));
  jand g09976(.dina(n10231), .dinb(n10226), .dout(n10232));
  jxor g09977(.dina(n10232), .dinb(a35 ), .dout(n10233));
  jxor g09978(.dina(n10233), .dinb(n10225), .dout(n10234));
  jxor g09979(.dina(n10234), .dinb(n10093), .dout(n10235));
  jnot g09980(.din(n10235), .dout(n10236));
  jor  g09981(.dina(n3032), .dinb(n3301), .dout(n10237));
  jor  g09982(.dina(n3136), .dinb(n2579), .dout(n10238));
  jor  g09983(.dina(n3304), .dinb(n2870), .dout(n10239));
  jor  g09984(.dina(n3306), .dinb(n3035), .dout(n10240));
  jand g09985(.dina(n10240), .dinb(n10239), .dout(n10241));
  jand g09986(.dina(n10241), .dinb(n10238), .dout(n10242));
  jand g09987(.dina(n10242), .dinb(n10237), .dout(n10243));
  jxor g09988(.dina(n10243), .dinb(a32 ), .dout(n10244));
  jxor g09989(.dina(n10244), .dinb(n10236), .dout(n10245));
  jxor g09990(.dina(n10245), .dinb(n10088), .dout(n10246));
  jxor g09991(.dina(n10246), .dinb(n10083), .dout(n10247));
  jxor g09992(.dina(n10247), .dinb(n10074), .dout(n10248));
  jnot g09993(.din(n10248), .dout(n10249));
  jor  g09994(.dina(n4137), .dinb(n2319), .dout(n10250));
  jor  g09995(.dina(n2224), .dinb(n3588), .dout(n10251));
  jor  g09996(.dina(n2322), .dinb(n3942), .dout(n10252));
  jor  g09997(.dina(n2324), .dinb(n4140), .dout(n10253));
  jand g09998(.dina(n10253), .dinb(n10252), .dout(n10254));
  jand g09999(.dina(n10254), .dinb(n10251), .dout(n10255));
  jand g10000(.dina(n10255), .dinb(n10250), .dout(n10256));
  jxor g10001(.dina(n10256), .dinb(a26 ), .dout(n10257));
  jxor g10002(.dina(n10257), .dinb(n10249), .dout(n10258));
  jxor g10003(.dina(n10258), .dinb(n10069), .dout(n10259));
  jor  g10004(.dina(n4554), .dinb(n1939), .dout(n10260));
  jor  g10005(.dina(n1827), .dinb(n4340), .dout(n10261));
  jor  g10006(.dina(n1942), .dinb(n4537), .dout(n10262));
  jor  g10007(.dina(n1944), .dinb(n4557), .dout(n10263));
  jand g10008(.dina(n10263), .dinb(n10262), .dout(n10264));
  jand g10009(.dina(n10264), .dinb(n10261), .dout(n10265));
  jand g10010(.dina(n10265), .dinb(n10260), .dout(n10266));
  jxor g10011(.dina(n10266), .dinb(a23 ), .dout(n10267));
  jxor g10012(.dina(n10267), .dinb(n10259), .dout(n10268));
  jxor g10013(.dina(n10268), .dinb(n10066), .dout(n10269));
  jor  g10014(.dina(n5405), .dinb(n1566), .dout(n10270));
  jor  g10015(.dina(n1489), .dinb(n4974), .dout(n10271));
  jor  g10016(.dina(n1569), .dinb(n4994), .dout(n10272));
  jor  g10017(.dina(n1571), .dinb(n5408), .dout(n10273));
  jand g10018(.dina(n10273), .dinb(n10272), .dout(n10274));
  jand g10019(.dina(n10274), .dinb(n10271), .dout(n10275));
  jand g10020(.dina(n10275), .dinb(n10270), .dout(n10276));
  jxor g10021(.dina(n10276), .dinb(a20 ), .dout(n10277));
  jxor g10022(.dina(n10277), .dinb(n10269), .dout(n10278));
  jxor g10023(.dina(n10278), .dinb(n10055), .dout(n10279));
  jxor g10024(.dina(n10279), .dinb(n10051), .dout(n10280));
  jxor g10025(.dina(n10280), .dinb(n10042), .dout(n10281));
  jxor g10026(.dina(n10281), .dinb(n10039), .dout(n10282));
  jxor g10027(.dina(n10282), .dinb(n10030), .dout(n10283));
  jxor g10028(.dina(n10283), .dinb(n10027), .dout(n10284));
  jnot g10029(.din(n10284), .dout(n10285));
  jxor g10030(.dina(n10285), .dinb(n10019), .dout(n10286));
  jor  g10031(.dina(n8228), .dinb(n528), .dout(n10287));
  jor  g10032(.dina(n490), .dinb(n7683), .dout(n10288));
  jor  g10033(.dina(n531), .dinb(n7960), .dout(n10289));
  jor  g10034(.dina(n533), .dinb(n8231), .dout(n10290));
  jand g10035(.dina(n10290), .dinb(n10289), .dout(n10291));
  jand g10036(.dina(n10291), .dinb(n10288), .dout(n10292));
  jand g10037(.dina(n10292), .dinb(n10287), .dout(n10293));
  jxor g10038(.dina(n10293), .dinb(a8 ), .dout(n10294));
  jxor g10039(.dina(n10294), .dinb(n10286), .dout(n10295));
  jxor g10040(.dina(n10295), .dinb(n10014), .dout(n10296));
  jor  g10041(.dina(n9387), .dinb(n402), .dout(n10297));
  jor  g10042(.dina(n371), .dinb(n8789), .dout(n10298));
  jor  g10043(.dina(n405), .dinb(n8809), .dout(n10299));
  jor  g10044(.dina(n332), .dinb(n9390), .dout(n10300));
  jand g10045(.dina(n10300), .dinb(n10299), .dout(n10301));
  jand g10046(.dina(n10301), .dinb(n10298), .dout(n10302));
  jand g10047(.dina(n10302), .dinb(n10297), .dout(n10303));
  jxor g10048(.dina(n10303), .dinb(a5 ), .dout(n10304));
  jxor g10049(.dina(n10304), .dinb(n10296), .dout(n10305));
  jand g10050(.dina(b60 ), .dinb(b59 ), .dout(n10306));
  jand g10051(.dina(n9720), .dinb(n9719), .dout(n10307));
  jor  g10052(.dina(n10307), .dinb(n10306), .dout(n10308));
  jxor g10053(.dina(b61 ), .dinb(b60 ), .dout(n10309));
  jnot g10054(.din(n10309), .dout(n10310));
  jxor g10055(.dina(n10310), .dinb(n10308), .dout(n10311));
  jor  g10056(.dina(n10311), .dinb(n264), .dout(n10312));
  jor  g10057(.dina(n284), .dinb(n9413), .dout(n10313));
  jnot g10058(.din(b61 ), .dout(n10314));
  jor  g10059(.dina(n269), .dinb(n10314), .dout(n10315));
  jor  g10060(.dina(n271), .dinb(n9725), .dout(n10316));
  jand g10061(.dina(n10316), .dinb(n10315), .dout(n10317));
  jand g10062(.dina(n10317), .dinb(n10313), .dout(n10318));
  jand g10063(.dina(n10318), .dinb(n10312), .dout(n10319));
  jxor g10064(.dina(n10319), .dinb(a2 ), .dout(n10320));
  jxor g10065(.dina(n10320), .dinb(n10305), .dout(n10321));
  jxor g10066(.dina(n10321), .dinb(n10011), .dout(n10322));
  jand g10067(.dina(n10006), .dinb(n9716), .dout(n10323));
  jand g10068(.dina(n10007), .dinb(n9713), .dout(n10324));
  jor  g10069(.dina(n10324), .dinb(n10323), .dout(n10325));
  jxor g10070(.dina(n10325), .dinb(n10322), .dout(f61 ));
  jand g10071(.dina(n10321), .dinb(n10011), .dout(n10327));
  jand g10072(.dina(n10325), .dinb(n10322), .dout(n10328));
  jor  g10073(.dina(n10328), .dinb(n10327), .dout(n10329));
  jor  g10074(.dina(n10294), .dinb(n10286), .dout(n10330));
  jnot g10075(.din(n10330), .dout(n10331));
  jand g10076(.dina(n10295), .dinb(n10014), .dout(n10332));
  jor  g10077(.dina(n10332), .dinb(n10331), .dout(n10333));
  jnot g10078(.din(n10027), .dout(n10334));
  jand g10079(.dina(n10283), .dinb(n10334), .dout(n10335));
  jnot g10080(.din(n10335), .dout(n10336));
  jor  g10081(.dina(n10284), .dinb(n10019), .dout(n10337));
  jand g10082(.dina(n10337), .dinb(n10336), .dout(n10338));
  jor  g10083(.dina(n7680), .dinb(n706), .dout(n10339));
  jor  g10084(.dina(n683), .dinb(n7149), .dout(n10340));
  jor  g10085(.dina(n709), .dinb(n7411), .dout(n10341));
  jor  g10086(.dina(n711), .dinb(n7683), .dout(n10342));
  jand g10087(.dina(n10342), .dinb(n10341), .dout(n10343));
  jand g10088(.dina(n10343), .dinb(n10340), .dout(n10344));
  jand g10089(.dina(n10344), .dinb(n10339), .dout(n10345));
  jxor g10090(.dina(n10345), .dinb(a11 ), .dout(n10346));
  jand g10091(.dina(n10281), .dinb(n10039), .dout(n10347));
  jand g10092(.dina(n10282), .dinb(n10030), .dout(n10348));
  jor  g10093(.dina(n10348), .dinb(n10347), .dout(n10349));
  jand g10094(.dina(n10279), .dinb(n10051), .dout(n10350));
  jand g10095(.dina(n10280), .dinb(n10042), .dout(n10351));
  jor  g10096(.dina(n10351), .dinb(n10350), .dout(n10352));
  jor  g10097(.dina(n6349), .dinb(n1245), .dout(n10353));
  jor  g10098(.dina(n1165), .dinb(n5862), .dout(n10354));
  jor  g10099(.dina(n1248), .dinb(n6106), .dout(n10355));
  jor  g10100(.dina(n1250), .dinb(n6352), .dout(n10356));
  jand g10101(.dina(n10356), .dinb(n10355), .dout(n10357));
  jand g10102(.dina(n10357), .dinb(n10354), .dout(n10358));
  jand g10103(.dina(n10358), .dinb(n10353), .dout(n10359));
  jxor g10104(.dina(n10359), .dinb(a17 ), .dout(n10360));
  jnot g10105(.din(n10360), .dout(n10361));
  jor  g10106(.dina(n10277), .dinb(n10269), .dout(n10362));
  jnot g10107(.din(n10362), .dout(n10363));
  jand g10108(.dina(n10278), .dinb(n10055), .dout(n10364));
  jor  g10109(.dina(n10364), .dinb(n10363), .dout(n10365));
  jnot g10110(.din(n10259), .dout(n10366));
  jor  g10111(.dina(n10267), .dinb(n10366), .dout(n10367));
  jnot g10112(.din(n10367), .dout(n10368));
  jnot g10113(.din(n10268), .dout(n10369));
  jand g10114(.dina(n10369), .dinb(n10066), .dout(n10370));
  jor  g10115(.dina(n10370), .dinb(n10368), .dout(n10371));
  jor  g10116(.dina(n10257), .dinb(n10249), .dout(n10372));
  jnot g10117(.din(n10372), .dout(n10373));
  jand g10118(.dina(n10258), .dinb(n10069), .dout(n10374));
  jor  g10119(.dina(n10374), .dinb(n10373), .dout(n10375));
  jand g10120(.dina(n10246), .dinb(n10083), .dout(n10376));
  jand g10121(.dina(n10247), .dinb(n10074), .dout(n10377));
  jor  g10122(.dina(n10377), .dinb(n10376), .dout(n10378));
  jor  g10123(.dina(n10244), .dinb(n10236), .dout(n10379));
  jand g10124(.dina(n10245), .dinb(n10088), .dout(n10380));
  jnot g10125(.din(n10380), .dout(n10381));
  jand g10126(.dina(n10381), .dinb(n10379), .dout(n10382));
  jnot g10127(.din(n10382), .dout(n10383));
  jor  g10128(.dina(n10233), .dinb(n10225), .dout(n10384));
  jand g10129(.dina(n10234), .dinb(n10093), .dout(n10385));
  jnot g10130(.din(n10385), .dout(n10386));
  jand g10131(.dina(n10386), .dinb(n10384), .dout(n10387));
  jnot g10132(.din(n10387), .dout(n10388));
  jor  g10133(.dina(n10222), .dinb(n10214), .dout(n10389));
  jand g10134(.dina(n10223), .dinb(n10098), .dout(n10390));
  jnot g10135(.din(n10390), .dout(n10391));
  jand g10136(.dina(n10391), .dinb(n10389), .dout(n10392));
  jnot g10137(.din(n10392), .dout(n10393));
  jor  g10138(.dina(n10211), .dinb(n10203), .dout(n10394));
  jand g10139(.dina(n10212), .dinb(n10101), .dout(n10395));
  jnot g10140(.din(n10395), .dout(n10396));
  jand g10141(.dina(n10396), .dinb(n10394), .dout(n10397));
  jnot g10142(.din(n10397), .dout(n10398));
  jor  g10143(.dina(n5096), .dinb(n1864), .dout(n10399));
  jor  g10144(.dina(n4904), .dinb(n1620), .dout(n10400));
  jor  g10145(.dina(n5099), .dinb(n1742), .dout(n10401));
  jor  g10146(.dina(n5101), .dinb(n1867), .dout(n10402));
  jand g10147(.dina(n10402), .dinb(n10401), .dout(n10403));
  jand g10148(.dina(n10403), .dinb(n10400), .dout(n10404));
  jand g10149(.dina(n10404), .dinb(n10399), .dout(n10405));
  jxor g10150(.dina(n10405), .dinb(a41 ), .dout(n10406));
  jnot g10151(.din(n10406), .dout(n10407));
  jor  g10152(.dina(n10200), .dinb(n10192), .dout(n10408));
  jand g10153(.dina(n10201), .dinb(n10104), .dout(n10409));
  jnot g10154(.din(n10409), .dout(n10410));
  jand g10155(.dina(n10410), .dinb(n10408), .dout(n10411));
  jnot g10156(.din(n10411), .dout(n10412));
  jor  g10157(.dina(n5739), .dinb(n1417), .dout(n10413));
  jor  g10158(.dina(n5574), .dinb(n1290), .dout(n10414));
  jor  g10159(.dina(n5742), .dinb(n1400), .dout(n10415));
  jor  g10160(.dina(n5744), .dinb(n1420), .dout(n10416));
  jand g10161(.dina(n10416), .dinb(n10415), .dout(n10417));
  jand g10162(.dina(n10417), .dinb(n10414), .dout(n10418));
  jand g10163(.dina(n10418), .dinb(n10413), .dout(n10419));
  jxor g10164(.dina(n10419), .dinb(a44 ), .dout(n10420));
  jnot g10165(.din(n10420), .dout(n10421));
  jor  g10166(.dina(n10189), .dinb(n10181), .dout(n10422));
  jand g10167(.dina(n10190), .dinb(n10107), .dout(n10423));
  jnot g10168(.din(n10423), .dout(n10424));
  jand g10169(.dina(n10424), .dinb(n10422), .dout(n10425));
  jnot g10170(.din(n10425), .dout(n10426));
  jor  g10171(.dina(n6490), .dinb(n1190), .dout(n10427));
  jor  g10172(.dina(n6262), .dinb(n939), .dout(n10428));
  jor  g10173(.dina(n6493), .dinb(n1022), .dout(n10429));
  jor  g10174(.dina(n6495), .dinb(n1193), .dout(n10430));
  jand g10175(.dina(n10430), .dinb(n10429), .dout(n10431));
  jand g10176(.dina(n10431), .dinb(n10428), .dout(n10432));
  jand g10177(.dina(n10432), .dinb(n10427), .dout(n10433));
  jxor g10178(.dina(n10433), .dinb(a47 ), .dout(n10434));
  jnot g10179(.din(n10434), .dout(n10435));
  jor  g10180(.dina(n10178), .dinb(n10170), .dout(n10436));
  jand g10181(.dina(n10179), .dinb(n10110), .dout(n10437));
  jnot g10182(.din(n10437), .dout(n10438));
  jand g10183(.dina(n10438), .dinb(n10436), .dout(n10439));
  jnot g10184(.din(n10439), .dout(n10440));
  jor  g10185(.dina(n10167), .dinb(n10159), .dout(n10441));
  jand g10186(.dina(n10168), .dinb(n10113), .dout(n10442));
  jnot g10187(.din(n10442), .dout(n10443));
  jand g10188(.dina(n10443), .dinb(n10441), .dout(n10444));
  jnot g10189(.din(n10444), .dout(n10445));
  jor  g10190(.dina(n8125), .dinb(n644), .dout(n10446));
  jor  g10191(.dina(n7846), .dinb(n564), .dout(n10447));
  jor  g10192(.dina(n8128), .dinb(n627), .dout(n10448));
  jor  g10193(.dina(n8130), .dinb(n647), .dout(n10449));
  jand g10194(.dina(n10449), .dinb(n10448), .dout(n10450));
  jand g10195(.dina(n10450), .dinb(n10447), .dout(n10451));
  jand g10196(.dina(n10451), .dinb(n10446), .dout(n10452));
  jxor g10197(.dina(n10452), .dinb(a53 ), .dout(n10453));
  jnot g10198(.din(n10453), .dout(n10454));
  jand g10199(.dina(n10156), .dinb(n10127), .dout(n10455));
  jand g10200(.dina(n10157), .dinb(n10118), .dout(n10456));
  jor  g10201(.dina(n10456), .dinb(n10455), .dout(n10457));
  jor  g10202(.dina(n8978), .dinb(n509), .dout(n10458));
  jor  g10203(.dina(n8677), .dinb(n395), .dout(n10459));
  jor  g10204(.dina(n8981), .dinb(n431), .dout(n10460));
  jor  g10205(.dina(n8983), .dinb(n512), .dout(n10461));
  jand g10206(.dina(n10461), .dinb(n10460), .dout(n10462));
  jand g10207(.dina(n10462), .dinb(n10459), .dout(n10463));
  jand g10208(.dina(n10463), .dinb(n10458), .dout(n10464));
  jxor g10209(.dina(n10464), .dinb(a56 ), .dout(n10465));
  jnot g10210(.din(n10465), .dout(n10466));
  jand g10211(.dina(n10154), .dinb(n10140), .dout(n10467));
  jand g10212(.dina(n10155), .dinb(n10131), .dout(n10468));
  jor  g10213(.dina(n10468), .dinb(n10467), .dout(n10469));
  jor  g10214(.dina(n9891), .dinb(n354), .dout(n10470));
  jor  g10215(.dina(n9593), .dinb(n299), .dout(n10471));
  jor  g10216(.dina(n9894), .dinb(n322), .dout(n10472));
  jor  g10217(.dina(n9896), .dinb(n357), .dout(n10473));
  jand g10218(.dina(n10473), .dinb(n10472), .dout(n10474));
  jand g10219(.dina(n10474), .dinb(n10471), .dout(n10475));
  jand g10220(.dina(n10475), .dinb(n10470), .dout(n10476));
  jxor g10221(.dina(n10476), .dinb(a59 ), .dout(n10477));
  jnot g10222(.din(n10477), .dout(n10478));
  jnot g10223(.din(n10153), .dout(n10479));
  jand g10224(.dina(n9905), .dinb(a62 ), .dout(n10480));
  jand g10225(.dina(n10480), .dinb(n10479), .dout(n10481));
  jnot g10226(.din(n10481), .dout(n10482));
  jand g10227(.dina(n10482), .dinb(a62 ), .dout(n10483));
  jor  g10228(.dina(n10147), .dinb(n10143), .dout(n10484));
  jor  g10229(.dina(n10484), .dinb(n9903), .dout(n10485));
  jnot g10230(.din(n10485), .dout(n10486));
  jand g10231(.dina(n10486), .dinb(b0 ), .dout(n10487));
  jand g10232(.dina(n10144), .dinb(b2 ), .dout(n10488));
  jand g10233(.dina(n10148), .dinb(b1 ), .dout(n10489));
  jand g10234(.dina(n10150), .dinb(n375), .dout(n10490));
  jor  g10235(.dina(n10490), .dinb(n10489), .dout(n10491));
  jor  g10236(.dina(n10491), .dinb(n10488), .dout(n10492));
  jor  g10237(.dina(n10492), .dinb(n10487), .dout(n10493));
  jxor g10238(.dina(n10493), .dinb(n10483), .dout(n10494));
  jxor g10239(.dina(n10494), .dinb(n10478), .dout(n10495));
  jxor g10240(.dina(n10495), .dinb(n10469), .dout(n10496));
  jxor g10241(.dina(n10496), .dinb(n10466), .dout(n10497));
  jxor g10242(.dina(n10497), .dinb(n10457), .dout(n10498));
  jxor g10243(.dina(n10498), .dinb(n10454), .dout(n10499));
  jxor g10244(.dina(n10499), .dinb(n10445), .dout(n10500));
  jnot g10245(.din(n10500), .dout(n10501));
  jor  g10246(.dina(n7266), .dinb(n855), .dout(n10502));
  jor  g10247(.dina(n7021), .dinb(n758), .dout(n10503));
  jor  g10248(.dina(n7269), .dinb(n778), .dout(n10504));
  jor  g10249(.dina(n7271), .dinb(n858), .dout(n10505));
  jand g10250(.dina(n10505), .dinb(n10504), .dout(n10506));
  jand g10251(.dina(n10506), .dinb(n10503), .dout(n10507));
  jand g10252(.dina(n10507), .dinb(n10502), .dout(n10508));
  jxor g10253(.dina(n10508), .dinb(a50 ), .dout(n10509));
  jxor g10254(.dina(n10509), .dinb(n10501), .dout(n10510));
  jxor g10255(.dina(n10510), .dinb(n10440), .dout(n10511));
  jxor g10256(.dina(n10511), .dinb(n10435), .dout(n10512));
  jxor g10257(.dina(n10512), .dinb(n10426), .dout(n10513));
  jxor g10258(.dina(n10513), .dinb(n10421), .dout(n10514));
  jxor g10259(.dina(n10514), .dinb(n10412), .dout(n10515));
  jxor g10260(.dina(n10515), .dinb(n10407), .dout(n10516));
  jxor g10261(.dina(n10516), .dinb(n10398), .dout(n10517));
  jnot g10262(.din(n10517), .dout(n10518));
  jor  g10263(.dina(n4415), .dinb(n2145), .dout(n10519));
  jor  g10264(.dina(n4272), .dinb(n1887), .dout(n10520));
  jor  g10265(.dina(n4418), .dinb(n2010), .dout(n10521));
  jor  g10266(.dina(n4420), .dinb(n2148), .dout(n10522));
  jand g10267(.dina(n10522), .dinb(n10521), .dout(n10523));
  jand g10268(.dina(n10523), .dinb(n10520), .dout(n10524));
  jand g10269(.dina(n10524), .dinb(n10519), .dout(n10525));
  jxor g10270(.dina(n10525), .dinb(a38 ), .dout(n10526));
  jxor g10271(.dina(n10526), .dinb(n10518), .dout(n10527));
  jxor g10272(.dina(n10527), .dinb(n10393), .dout(n10528));
  jnot g10273(.din(n10528), .dout(n10529));
  jor  g10274(.dina(n3849), .dinb(n2576), .dout(n10530));
  jor  g10275(.dina(n3689), .dinb(n2407), .dout(n10531));
  jor  g10276(.dina(n3852), .dinb(n2559), .dout(n10532));
  jor  g10277(.dina(n3854), .dinb(n2579), .dout(n10533));
  jand g10278(.dina(n10533), .dinb(n10532), .dout(n10534));
  jand g10279(.dina(n10534), .dinb(n10531), .dout(n10535));
  jand g10280(.dina(n10535), .dinb(n10530), .dout(n10536));
  jxor g10281(.dina(n10536), .dinb(a35 ), .dout(n10537));
  jxor g10282(.dina(n10537), .dinb(n10529), .dout(n10538));
  jxor g10283(.dina(n10538), .dinb(n10388), .dout(n10539));
  jnot g10284(.din(n10539), .dout(n10540));
  jor  g10285(.dina(n3052), .dinb(n3301), .dout(n10541));
  jor  g10286(.dina(n3136), .dinb(n2870), .dout(n10542));
  jor  g10287(.dina(n3304), .dinb(n3035), .dout(n10543));
  jor  g10288(.dina(n3306), .dinb(n3055), .dout(n10544));
  jand g10289(.dina(n10544), .dinb(n10543), .dout(n10545));
  jand g10290(.dina(n10545), .dinb(n10542), .dout(n10546));
  jand g10291(.dina(n10546), .dinb(n10541), .dout(n10547));
  jxor g10292(.dina(n10547), .dinb(a32 ), .dout(n10548));
  jxor g10293(.dina(n10548), .dinb(n10540), .dout(n10549));
  jxor g10294(.dina(n10549), .dinb(n10383), .dout(n10550));
  jnot g10295(.din(n10550), .dout(n10551));
  jor  g10296(.dina(n3585), .dinb(n2784), .dout(n10552));
  jor  g10297(.dina(n2661), .dinb(n3230), .dout(n10553));
  jor  g10298(.dina(n2787), .dinb(n3403), .dout(n10554));
  jor  g10299(.dina(n2789), .dinb(n3588), .dout(n10555));
  jand g10300(.dina(n10555), .dinb(n10554), .dout(n10556));
  jand g10301(.dina(n10556), .dinb(n10553), .dout(n10557));
  jand g10302(.dina(n10557), .dinb(n10552), .dout(n10558));
  jxor g10303(.dina(n10558), .dinb(a29 ), .dout(n10559));
  jxor g10304(.dina(n10559), .dinb(n10551), .dout(n10560));
  jxor g10305(.dina(n10560), .dinb(n10378), .dout(n10561));
  jnot g10306(.din(n10561), .dout(n10562));
  jor  g10307(.dina(n4337), .dinb(n2319), .dout(n10563));
  jor  g10308(.dina(n2224), .dinb(n3942), .dout(n10564));
  jor  g10309(.dina(n2322), .dinb(n4140), .dout(n10565));
  jor  g10310(.dina(n2324), .dinb(n4340), .dout(n10566));
  jand g10311(.dina(n10566), .dinb(n10565), .dout(n10567));
  jand g10312(.dina(n10567), .dinb(n10564), .dout(n10568));
  jand g10313(.dina(n10568), .dinb(n10563), .dout(n10569));
  jxor g10314(.dina(n10569), .dinb(a26 ), .dout(n10570));
  jxor g10315(.dina(n10570), .dinb(n10562), .dout(n10571));
  jxor g10316(.dina(n10571), .dinb(n10375), .dout(n10572));
  jnot g10317(.din(n10572), .dout(n10573));
  jor  g10318(.dina(n4971), .dinb(n1939), .dout(n10574));
  jor  g10319(.dina(n1827), .dinb(n4537), .dout(n10575));
  jor  g10320(.dina(n1942), .dinb(n4557), .dout(n10576));
  jor  g10321(.dina(n1944), .dinb(n4974), .dout(n10577));
  jand g10322(.dina(n10577), .dinb(n10576), .dout(n10578));
  jand g10323(.dina(n10578), .dinb(n10575), .dout(n10579));
  jand g10324(.dina(n10579), .dinb(n10574), .dout(n10580));
  jxor g10325(.dina(n10580), .dinb(a23 ), .dout(n10581));
  jxor g10326(.dina(n10581), .dinb(n10573), .dout(n10582));
  jxor g10327(.dina(n10582), .dinb(n10371), .dout(n10583));
  jor  g10328(.dina(n5425), .dinb(n1566), .dout(n10584));
  jor  g10329(.dina(n1489), .dinb(n4994), .dout(n10585));
  jor  g10330(.dina(n1569), .dinb(n5408), .dout(n10586));
  jor  g10331(.dina(n1571), .dinb(n5428), .dout(n10587));
  jand g10332(.dina(n10587), .dinb(n10586), .dout(n10588));
  jand g10333(.dina(n10588), .dinb(n10585), .dout(n10589));
  jand g10334(.dina(n10589), .dinb(n10584), .dout(n10590));
  jxor g10335(.dina(n10590), .dinb(a20 ), .dout(n10591));
  jnot g10336(.din(n10591), .dout(n10592));
  jxor g10337(.dina(n10592), .dinb(n10583), .dout(n10593));
  jxor g10338(.dina(n10593), .dinb(n10365), .dout(n10594));
  jxor g10339(.dina(n10594), .dinb(n10361), .dout(n10595));
  jxor g10340(.dina(n10595), .dinb(n10352), .dout(n10596));
  jor  g10341(.dina(n7126), .dinb(n974), .dout(n10597));
  jor  g10342(.dina(n908), .dinb(n6372), .dout(n10598));
  jor  g10343(.dina(n977), .dinb(n6867), .dout(n10599));
  jor  g10344(.dina(n979), .dinb(n7129), .dout(n10600));
  jand g10345(.dina(n10600), .dinb(n10599), .dout(n10601));
  jand g10346(.dina(n10601), .dinb(n10598), .dout(n10602));
  jand g10347(.dina(n10602), .dinb(n10597), .dout(n10603));
  jxor g10348(.dina(n10603), .dinb(a14 ), .dout(n10604));
  jnot g10349(.din(n10604), .dout(n10605));
  jxor g10350(.dina(n10605), .dinb(n10596), .dout(n10606));
  jxor g10351(.dina(n10606), .dinb(n10349), .dout(n10607));
  jxor g10352(.dina(n10607), .dinb(n10346), .dout(n10608));
  jxor g10353(.dina(n10608), .dinb(n10338), .dout(n10609));
  jor  g10354(.dina(n8786), .dinb(n528), .dout(n10610));
  jor  g10355(.dina(n490), .dinb(n7960), .dout(n10611));
  jor  g10356(.dina(n531), .dinb(n8231), .dout(n10612));
  jor  g10357(.dina(n533), .dinb(n8789), .dout(n10613));
  jand g10358(.dina(n10613), .dinb(n10612), .dout(n10614));
  jand g10359(.dina(n10614), .dinb(n10611), .dout(n10615));
  jand g10360(.dina(n10615), .dinb(n10610), .dout(n10616));
  jxor g10361(.dina(n10616), .dinb(a8 ), .dout(n10617));
  jxor g10362(.dina(n10617), .dinb(n10609), .dout(n10618));
  jor  g10363(.dina(n9410), .dinb(n402), .dout(n10619));
  jor  g10364(.dina(n371), .dinb(n8809), .dout(n10620));
  jor  g10365(.dina(n405), .dinb(n9390), .dout(n10621));
  jor  g10366(.dina(n332), .dinb(n9413), .dout(n10622));
  jand g10367(.dina(n10622), .dinb(n10621), .dout(n10623));
  jand g10368(.dina(n10623), .dinb(n10620), .dout(n10624));
  jand g10369(.dina(n10624), .dinb(n10619), .dout(n10625));
  jxor g10370(.dina(n10625), .dinb(a5 ), .dout(n10626));
  jxor g10371(.dina(n10626), .dinb(n10618), .dout(n10627));
  jxor g10372(.dina(n10627), .dinb(n10333), .dout(n10628));
  jand g10373(.dina(b61 ), .dinb(b60 ), .dout(n10629));
  jand g10374(.dina(n10309), .dinb(n10308), .dout(n10630));
  jor  g10375(.dina(n10630), .dinb(n10629), .dout(n10631));
  jxor g10376(.dina(b62 ), .dinb(b61 ), .dout(n10632));
  jnot g10377(.din(n10632), .dout(n10633));
  jxor g10378(.dina(n10633), .dinb(n10631), .dout(n10634));
  jor  g10379(.dina(n10634), .dinb(n264), .dout(n10635));
  jor  g10380(.dina(n284), .dinb(n9725), .dout(n10636));
  jnot g10381(.din(b62 ), .dout(n10637));
  jor  g10382(.dina(n269), .dinb(n10637), .dout(n10638));
  jor  g10383(.dina(n271), .dinb(n10314), .dout(n10639));
  jand g10384(.dina(n10639), .dinb(n10638), .dout(n10640));
  jand g10385(.dina(n10640), .dinb(n10636), .dout(n10641));
  jand g10386(.dina(n10641), .dinb(n10635), .dout(n10642));
  jxor g10387(.dina(n10642), .dinb(n260), .dout(n10643));
  jxor g10388(.dina(n10643), .dinb(n10628), .dout(n10644));
  jnot g10389(.din(n10296), .dout(n10645));
  jor  g10390(.dina(n10304), .dinb(n10645), .dout(n10646));
  jnot g10391(.din(n10646), .dout(n10647));
  jand g10392(.dina(n10304), .dinb(n10645), .dout(n10648));
  jnot g10393(.din(n10648), .dout(n10649));
  jxor g10394(.dina(n10319), .dinb(n260), .dout(n10650));
  jand g10395(.dina(n10650), .dinb(n10649), .dout(n10651));
  jor  g10396(.dina(n10651), .dinb(n10647), .dout(n10652));
  jxor g10397(.dina(n10652), .dinb(n10644), .dout(n10653));
  jxor g10398(.dina(n10653), .dinb(n10329), .dout(f62 ));
  jand g10399(.dina(n10652), .dinb(n10644), .dout(n10655));
  jand g10400(.dina(n10653), .dinb(n10329), .dout(n10656));
  jor  g10401(.dina(n10656), .dinb(n10655), .dout(n10657));
  jand g10402(.dina(n10627), .dinb(n10333), .dout(n10658));
  jand g10403(.dina(n10643), .dinb(n10628), .dout(n10659));
  jor  g10404(.dina(n10659), .dinb(n10658), .dout(n10660));
  jor  g10405(.dina(n9722), .dinb(n402), .dout(n10661));
  jor  g10406(.dina(n371), .dinb(n9390), .dout(n10662));
  jor  g10407(.dina(n405), .dinb(n9413), .dout(n10663));
  jor  g10408(.dina(n332), .dinb(n9725), .dout(n10664));
  jand g10409(.dina(n10664), .dinb(n10663), .dout(n10665));
  jand g10410(.dina(n10665), .dinb(n10662), .dout(n10666));
  jand g10411(.dina(n10666), .dinb(n10661), .dout(n10667));
  jxor g10412(.dina(n10667), .dinb(n364), .dout(n10668));
  jnot g10413(.din(n10668), .dout(n10669));
  jnot g10414(.din(n10346), .dout(n10670));
  jand g10415(.dina(n10607), .dinb(n10670), .dout(n10671));
  jnot g10416(.din(n10671), .dout(n10672));
  jor  g10417(.dina(n10608), .dinb(n10338), .dout(n10673));
  jand g10418(.dina(n10673), .dinb(n10672), .dout(n10674));
  jand g10419(.dina(n10605), .dinb(n10596), .dout(n10675));
  jand g10420(.dina(n10606), .dinb(n10349), .dout(n10676));
  jor  g10421(.dina(n10676), .dinb(n10675), .dout(n10677));
  jor  g10422(.dina(n7146), .dinb(n974), .dout(n10678));
  jor  g10423(.dina(n908), .dinb(n6867), .dout(n10679));
  jor  g10424(.dina(n977), .dinb(n7129), .dout(n10680));
  jor  g10425(.dina(n979), .dinb(n7149), .dout(n10681));
  jand g10426(.dina(n10681), .dinb(n10680), .dout(n10682));
  jand g10427(.dina(n10682), .dinb(n10679), .dout(n10683));
  jand g10428(.dina(n10683), .dinb(n10678), .dout(n10684));
  jxor g10429(.dina(n10684), .dinb(a14 ), .dout(n10685));
  jnot g10430(.din(n10685), .dout(n10686));
  jand g10431(.dina(n10594), .dinb(n10361), .dout(n10687));
  jand g10432(.dina(n10595), .dinb(n10352), .dout(n10688));
  jor  g10433(.dina(n10688), .dinb(n10687), .dout(n10689));
  jor  g10434(.dina(n6369), .dinb(n1245), .dout(n10690));
  jor  g10435(.dina(n1165), .dinb(n6106), .dout(n10691));
  jor  g10436(.dina(n1248), .dinb(n6352), .dout(n10692));
  jor  g10437(.dina(n1250), .dinb(n6372), .dout(n10693));
  jand g10438(.dina(n10693), .dinb(n10692), .dout(n10694));
  jand g10439(.dina(n10694), .dinb(n10691), .dout(n10695));
  jand g10440(.dina(n10695), .dinb(n10690), .dout(n10696));
  jxor g10441(.dina(n10696), .dinb(a17 ), .dout(n10697));
  jnot g10442(.din(n10697), .dout(n10698));
  jand g10443(.dina(n10592), .dinb(n10583), .dout(n10699));
  jand g10444(.dina(n10593), .dinb(n10365), .dout(n10700));
  jor  g10445(.dina(n10700), .dinb(n10699), .dout(n10701));
  jor  g10446(.dina(n5859), .dinb(n1566), .dout(n10702));
  jor  g10447(.dina(n1489), .dinb(n5408), .dout(n10703));
  jor  g10448(.dina(n1569), .dinb(n5428), .dout(n10704));
  jor  g10449(.dina(n1571), .dinb(n5862), .dout(n10705));
  jand g10450(.dina(n10705), .dinb(n10704), .dout(n10706));
  jand g10451(.dina(n10706), .dinb(n10703), .dout(n10707));
  jand g10452(.dina(n10707), .dinb(n10702), .dout(n10708));
  jxor g10453(.dina(n10708), .dinb(a20 ), .dout(n10709));
  jnot g10454(.din(n10709), .dout(n10710));
  jor  g10455(.dina(n10581), .dinb(n10573), .dout(n10711));
  jnot g10456(.din(n10711), .dout(n10712));
  jand g10457(.dina(n10582), .dinb(n10371), .dout(n10713));
  jor  g10458(.dina(n10713), .dinb(n10712), .dout(n10714));
  jor  g10459(.dina(n4991), .dinb(n1939), .dout(n10715));
  jor  g10460(.dina(n1827), .dinb(n4557), .dout(n10716));
  jor  g10461(.dina(n1942), .dinb(n4974), .dout(n10717));
  jor  g10462(.dina(n1944), .dinb(n4994), .dout(n10718));
  jand g10463(.dina(n10718), .dinb(n10717), .dout(n10719));
  jand g10464(.dina(n10719), .dinb(n10716), .dout(n10720));
  jand g10465(.dina(n10720), .dinb(n10715), .dout(n10721));
  jxor g10466(.dina(n10721), .dinb(a23 ), .dout(n10722));
  jnot g10467(.din(n10722), .dout(n10723));
  jor  g10468(.dina(n10570), .dinb(n10562), .dout(n10724));
  jnot g10469(.din(n10724), .dout(n10725));
  jand g10470(.dina(n10571), .dinb(n10375), .dout(n10726));
  jor  g10471(.dina(n10726), .dinb(n10725), .dout(n10727));
  jor  g10472(.dina(n10559), .dinb(n10551), .dout(n10728));
  jand g10473(.dina(n10560), .dinb(n10378), .dout(n10729));
  jnot g10474(.din(n10729), .dout(n10730));
  jand g10475(.dina(n10730), .dinb(n10728), .dout(n10731));
  jor  g10476(.dina(n3939), .dinb(n2784), .dout(n10732));
  jor  g10477(.dina(n2661), .dinb(n3403), .dout(n10733));
  jor  g10478(.dina(n2787), .dinb(n3588), .dout(n10734));
  jor  g10479(.dina(n2789), .dinb(n3942), .dout(n10735));
  jand g10480(.dina(n10735), .dinb(n10734), .dout(n10736));
  jand g10481(.dina(n10736), .dinb(n10733), .dout(n10737));
  jand g10482(.dina(n10737), .dinb(n10732), .dout(n10738));
  jxor g10483(.dina(n10738), .dinb(a29 ), .dout(n10739));
  jnot g10484(.din(n10739), .dout(n10740));
  jor  g10485(.dina(n10548), .dinb(n10540), .dout(n10741));
  jand g10486(.dina(n10549), .dinb(n10383), .dout(n10742));
  jnot g10487(.din(n10742), .dout(n10743));
  jand g10488(.dina(n10743), .dinb(n10741), .dout(n10744));
  jnot g10489(.din(n10744), .dout(n10745));
  jor  g10490(.dina(n10526), .dinb(n10518), .dout(n10746));
  jand g10491(.dina(n10527), .dinb(n10393), .dout(n10747));
  jnot g10492(.din(n10747), .dout(n10748));
  jand g10493(.dina(n10748), .dinb(n10746), .dout(n10749));
  jnot g10494(.din(n10749), .dout(n10750));
  jand g10495(.dina(n10515), .dinb(n10407), .dout(n10751));
  jand g10496(.dina(n10516), .dinb(n10398), .dout(n10752));
  jor  g10497(.dina(n10752), .dinb(n10751), .dout(n10753));
  jand g10498(.dina(n10513), .dinb(n10421), .dout(n10754));
  jand g10499(.dina(n10514), .dinb(n10412), .dout(n10755));
  jor  g10500(.dina(n10755), .dinb(n10754), .dout(n10756));
  jor  g10501(.dina(n5739), .dinb(n1617), .dout(n10757));
  jor  g10502(.dina(n5574), .dinb(n1400), .dout(n10758));
  jor  g10503(.dina(n5742), .dinb(n1420), .dout(n10759));
  jor  g10504(.dina(n5744), .dinb(n1620), .dout(n10760));
  jand g10505(.dina(n10760), .dinb(n10759), .dout(n10761));
  jand g10506(.dina(n10761), .dinb(n10758), .dout(n10762));
  jand g10507(.dina(n10762), .dinb(n10757), .dout(n10763));
  jxor g10508(.dina(n10763), .dinb(a44 ), .dout(n10764));
  jnot g10509(.din(n10764), .dout(n10765));
  jand g10510(.dina(n10511), .dinb(n10435), .dout(n10766));
  jand g10511(.dina(n10512), .dinb(n10426), .dout(n10767));
  jor  g10512(.dina(n10767), .dinb(n10766), .dout(n10768));
  jor  g10513(.dina(n10509), .dinb(n10501), .dout(n10769));
  jand g10514(.dina(n10510), .dinb(n10440), .dout(n10770));
  jnot g10515(.din(n10770), .dout(n10771));
  jand g10516(.dina(n10771), .dinb(n10769), .dout(n10772));
  jnot g10517(.din(n10772), .dout(n10773));
  jand g10518(.dina(n10498), .dinb(n10454), .dout(n10774));
  jand g10519(.dina(n10499), .dinb(n10445), .dout(n10775));
  jor  g10520(.dina(n10775), .dinb(n10774), .dout(n10776));
  jor  g10521(.dina(n8125), .dinb(n755), .dout(n10777));
  jor  g10522(.dina(n7846), .dinb(n627), .dout(n10778));
  jor  g10523(.dina(n8128), .dinb(n647), .dout(n10779));
  jor  g10524(.dina(n8130), .dinb(n758), .dout(n10780));
  jand g10525(.dina(n10780), .dinb(n10779), .dout(n10781));
  jand g10526(.dina(n10781), .dinb(n10778), .dout(n10782));
  jand g10527(.dina(n10782), .dinb(n10777), .dout(n10783));
  jxor g10528(.dina(n10783), .dinb(a53 ), .dout(n10784));
  jnot g10529(.din(n10784), .dout(n10785));
  jand g10530(.dina(n10496), .dinb(n10466), .dout(n10786));
  jand g10531(.dina(n10497), .dinb(n10457), .dout(n10787));
  jor  g10532(.dina(n10787), .dinb(n10786), .dout(n10788));
  jand g10533(.dina(n10494), .dinb(n10478), .dout(n10789));
  jand g10534(.dina(n10495), .dinb(n10469), .dout(n10790));
  jor  g10535(.dina(n10790), .dinb(n10789), .dout(n10791));
  jor  g10536(.dina(n9891), .dinb(n392), .dout(n10792));
  jor  g10537(.dina(n9593), .dinb(n322), .dout(n10793));
  jor  g10538(.dina(n9894), .dinb(n357), .dout(n10794));
  jor  g10539(.dina(n9896), .dinb(n395), .dout(n10795));
  jand g10540(.dina(n10795), .dinb(n10794), .dout(n10796));
  jand g10541(.dina(n10796), .dinb(n10793), .dout(n10797));
  jand g10542(.dina(n10797), .dinb(n10792), .dout(n10798));
  jxor g10543(.dina(n10798), .dinb(a59 ), .dout(n10799));
  jnot g10544(.din(n10799), .dout(n10800));
  jxor g10545(.dina(a63 ), .dinb(a62 ), .dout(n10801));
  jand g10546(.dina(n10801), .dinb(b0 ), .dout(n10802));
  jnot g10547(.din(n10802), .dout(n10803));
  jor  g10548(.dina(n10493), .dinb(n10482), .dout(n10804));
  jxor g10549(.dina(n10804), .dinb(n10803), .dout(n10805));
  jnot g10550(.din(n10150), .dout(n10806));
  jor  g10551(.dina(n10806), .dinb(n296), .dout(n10807));
  jor  g10552(.dina(n10485), .dinb(n267), .dout(n10808));
  jnot g10553(.din(n10148), .dout(n10809));
  jor  g10554(.dina(n10809), .dinb(n279), .dout(n10810));
  jnot g10555(.din(n10144), .dout(n10811));
  jor  g10556(.dina(n10811), .dinb(n299), .dout(n10812));
  jand g10557(.dina(n10812), .dinb(n10810), .dout(n10813));
  jand g10558(.dina(n10813), .dinb(n10808), .dout(n10814));
  jand g10559(.dina(n10814), .dinb(n10807), .dout(n10815));
  jxor g10560(.dina(n10815), .dinb(a62 ), .dout(n10816));
  jnot g10561(.din(n10816), .dout(n10817));
  jxor g10562(.dina(n10817), .dinb(n10805), .dout(n10818));
  jxor g10563(.dina(n10818), .dinb(n10800), .dout(n10819));
  jxor g10564(.dina(n10819), .dinb(n10791), .dout(n10820));
  jnot g10565(.din(n10820), .dout(n10821));
  jor  g10566(.dina(n8978), .dinb(n561), .dout(n10822));
  jor  g10567(.dina(n8677), .dinb(n431), .dout(n10823));
  jor  g10568(.dina(n8981), .dinb(n512), .dout(n10824));
  jor  g10569(.dina(n8983), .dinb(n564), .dout(n10825));
  jand g10570(.dina(n10825), .dinb(n10824), .dout(n10826));
  jand g10571(.dina(n10826), .dinb(n10823), .dout(n10827));
  jand g10572(.dina(n10827), .dinb(n10822), .dout(n10828));
  jxor g10573(.dina(n10828), .dinb(a56 ), .dout(n10829));
  jxor g10574(.dina(n10829), .dinb(n10821), .dout(n10830));
  jxor g10575(.dina(n10830), .dinb(n10788), .dout(n10831));
  jxor g10576(.dina(n10831), .dinb(n10785), .dout(n10832));
  jxor g10577(.dina(n10832), .dinb(n10776), .dout(n10833));
  jnot g10578(.din(n10833), .dout(n10834));
  jor  g10579(.dina(n7266), .dinb(n936), .dout(n10835));
  jor  g10580(.dina(n7021), .dinb(n778), .dout(n10836));
  jor  g10581(.dina(n7269), .dinb(n858), .dout(n10837));
  jor  g10582(.dina(n7271), .dinb(n939), .dout(n10838));
  jand g10583(.dina(n10838), .dinb(n10837), .dout(n10839));
  jand g10584(.dina(n10839), .dinb(n10836), .dout(n10840));
  jand g10585(.dina(n10840), .dinb(n10835), .dout(n10841));
  jxor g10586(.dina(n10841), .dinb(a50 ), .dout(n10842));
  jxor g10587(.dina(n10842), .dinb(n10834), .dout(n10843));
  jxor g10588(.dina(n10843), .dinb(n10773), .dout(n10844));
  jnot g10589(.din(n10844), .dout(n10845));
  jor  g10590(.dina(n6490), .dinb(n1287), .dout(n10846));
  jor  g10591(.dina(n6262), .dinb(n1022), .dout(n10847));
  jor  g10592(.dina(n6493), .dinb(n1193), .dout(n10848));
  jor  g10593(.dina(n6495), .dinb(n1290), .dout(n10849));
  jand g10594(.dina(n10849), .dinb(n10848), .dout(n10850));
  jand g10595(.dina(n10850), .dinb(n10847), .dout(n10851));
  jand g10596(.dina(n10851), .dinb(n10846), .dout(n10852));
  jxor g10597(.dina(n10852), .dinb(a47 ), .dout(n10853));
  jxor g10598(.dina(n10853), .dinb(n10845), .dout(n10854));
  jxor g10599(.dina(n10854), .dinb(n10768), .dout(n10855));
  jxor g10600(.dina(n10855), .dinb(n10765), .dout(n10856));
  jxor g10601(.dina(n10856), .dinb(n10756), .dout(n10857));
  jnot g10602(.din(n10857), .dout(n10858));
  jor  g10603(.dina(n5096), .dinb(n1884), .dout(n10859));
  jor  g10604(.dina(n4904), .dinb(n1742), .dout(n10860));
  jor  g10605(.dina(n5099), .dinb(n1867), .dout(n10861));
  jor  g10606(.dina(n5101), .dinb(n1887), .dout(n10862));
  jand g10607(.dina(n10862), .dinb(n10861), .dout(n10863));
  jand g10608(.dina(n10863), .dinb(n10860), .dout(n10864));
  jand g10609(.dina(n10864), .dinb(n10859), .dout(n10865));
  jxor g10610(.dina(n10865), .dinb(a41 ), .dout(n10866));
  jxor g10611(.dina(n10866), .dinb(n10858), .dout(n10867));
  jxor g10612(.dina(n10867), .dinb(n10753), .dout(n10868));
  jnot g10613(.din(n10868), .dout(n10869));
  jor  g10614(.dina(n4415), .dinb(n2404), .dout(n10870));
  jor  g10615(.dina(n4272), .dinb(n2010), .dout(n10871));
  jor  g10616(.dina(n4418), .dinb(n2148), .dout(n10872));
  jor  g10617(.dina(n4420), .dinb(n2407), .dout(n10873));
  jand g10618(.dina(n10873), .dinb(n10872), .dout(n10874));
  jand g10619(.dina(n10874), .dinb(n10871), .dout(n10875));
  jand g10620(.dina(n10875), .dinb(n10870), .dout(n10876));
  jxor g10621(.dina(n10876), .dinb(a38 ), .dout(n10877));
  jxor g10622(.dina(n10877), .dinb(n10869), .dout(n10878));
  jxor g10623(.dina(n10878), .dinb(n10750), .dout(n10879));
  jnot g10624(.din(n10879), .dout(n10880));
  jor  g10625(.dina(n3849), .dinb(n2867), .dout(n10881));
  jor  g10626(.dina(n3689), .dinb(n2559), .dout(n10882));
  jor  g10627(.dina(n3852), .dinb(n2579), .dout(n10883));
  jor  g10628(.dina(n3854), .dinb(n2870), .dout(n10884));
  jand g10629(.dina(n10884), .dinb(n10883), .dout(n10885));
  jand g10630(.dina(n10885), .dinb(n10882), .dout(n10886));
  jand g10631(.dina(n10886), .dinb(n10881), .dout(n10887));
  jxor g10632(.dina(n10887), .dinb(a35 ), .dout(n10888));
  jxor g10633(.dina(n10888), .dinb(n10880), .dout(n10889));
  jnot g10634(.din(n10889), .dout(n10890));
  jor  g10635(.dina(n10537), .dinb(n10529), .dout(n10891));
  jand g10636(.dina(n10538), .dinb(n10388), .dout(n10892));
  jnot g10637(.din(n10892), .dout(n10893));
  jand g10638(.dina(n10893), .dinb(n10891), .dout(n10894));
  jxor g10639(.dina(n10894), .dinb(n10890), .dout(n10895));
  jnot g10640(.din(n10895), .dout(n10896));
  jor  g10641(.dina(n3227), .dinb(n3301), .dout(n10897));
  jor  g10642(.dina(n3136), .dinb(n3035), .dout(n10898));
  jor  g10643(.dina(n3304), .dinb(n3055), .dout(n10899));
  jor  g10644(.dina(n3306), .dinb(n3230), .dout(n10900));
  jand g10645(.dina(n10900), .dinb(n10899), .dout(n10901));
  jand g10646(.dina(n10901), .dinb(n10898), .dout(n10902));
  jand g10647(.dina(n10902), .dinb(n10897), .dout(n10903));
  jxor g10648(.dina(n10903), .dinb(a32 ), .dout(n10904));
  jxor g10649(.dina(n10904), .dinb(n10896), .dout(n10905));
  jxor g10650(.dina(n10905), .dinb(n10745), .dout(n10906));
  jxor g10651(.dina(n10906), .dinb(n10740), .dout(n10907));
  jxor g10652(.dina(n10907), .dinb(n10731), .dout(n10908));
  jor  g10653(.dina(n4534), .dinb(n2319), .dout(n10909));
  jor  g10654(.dina(n2224), .dinb(n4140), .dout(n10910));
  jor  g10655(.dina(n2322), .dinb(n4340), .dout(n10911));
  jor  g10656(.dina(n2324), .dinb(n4537), .dout(n10912));
  jand g10657(.dina(n10912), .dinb(n10911), .dout(n10913));
  jand g10658(.dina(n10913), .dinb(n10910), .dout(n10914));
  jand g10659(.dina(n10914), .dinb(n10909), .dout(n10915));
  jxor g10660(.dina(n10915), .dinb(a26 ), .dout(n10916));
  jxor g10661(.dina(n10916), .dinb(n10908), .dout(n10917));
  jxor g10662(.dina(n10917), .dinb(n10727), .dout(n10918));
  jxor g10663(.dina(n10918), .dinb(n10723), .dout(n10919));
  jxor g10664(.dina(n10919), .dinb(n10714), .dout(n10920));
  jxor g10665(.dina(n10920), .dinb(n10710), .dout(n10921));
  jxor g10666(.dina(n10921), .dinb(n10701), .dout(n10922));
  jxor g10667(.dina(n10922), .dinb(n10698), .dout(n10923));
  jxor g10668(.dina(n10923), .dinb(n10689), .dout(n10924));
  jxor g10669(.dina(n10924), .dinb(n10686), .dout(n10925));
  jnot g10670(.din(n10925), .dout(n10926));
  jxor g10671(.dina(n10926), .dinb(n10677), .dout(n10927));
  jor  g10672(.dina(n7957), .dinb(n706), .dout(n10928));
  jor  g10673(.dina(n683), .dinb(n7411), .dout(n10929));
  jor  g10674(.dina(n709), .dinb(n7683), .dout(n10930));
  jor  g10675(.dina(n711), .dinb(n7960), .dout(n10931));
  jand g10676(.dina(n10931), .dinb(n10930), .dout(n10932));
  jand g10677(.dina(n10932), .dinb(n10929), .dout(n10933));
  jand g10678(.dina(n10933), .dinb(n10928), .dout(n10934));
  jxor g10679(.dina(n10934), .dinb(a11 ), .dout(n10935));
  jxor g10680(.dina(n10935), .dinb(n10927), .dout(n10936));
  jxor g10681(.dina(n10936), .dinb(n10674), .dout(n10937));
  jor  g10682(.dina(n8806), .dinb(n528), .dout(n10938));
  jor  g10683(.dina(n490), .dinb(n8231), .dout(n10939));
  jor  g10684(.dina(n531), .dinb(n8789), .dout(n10940));
  jor  g10685(.dina(n533), .dinb(n8809), .dout(n10941));
  jand g10686(.dina(n10941), .dinb(n10940), .dout(n10942));
  jand g10687(.dina(n10942), .dinb(n10939), .dout(n10943));
  jand g10688(.dina(n10943), .dinb(n10938), .dout(n10944));
  jxor g10689(.dina(n10944), .dinb(a8 ), .dout(n10945));
  jxor g10690(.dina(n10945), .dinb(n10937), .dout(n10946));
  jxor g10691(.dina(n10946), .dinb(n10669), .dout(n10947));
  jnot g10692(.din(n10609), .dout(n10948));
  jor  g10693(.dina(n10617), .dinb(n10948), .dout(n10949));
  jand g10694(.dina(n10617), .dinb(n10948), .dout(n10950));
  jor  g10695(.dina(n10626), .dinb(n10950), .dout(n10951));
  jand g10696(.dina(n10951), .dinb(n10949), .dout(n10952));
  jand g10697(.dina(n10952), .dinb(n10947), .dout(n10953));
  jor  g10698(.dina(n10952), .dinb(n10947), .dout(n10954));
  jnot g10699(.din(n10954), .dout(n10955));
  jor  g10700(.dina(n10955), .dinb(n10953), .dout(n10956));
  jand g10701(.dina(b62 ), .dinb(b61 ), .dout(n10957));
  jand g10702(.dina(n10632), .dinb(n10631), .dout(n10958));
  jor  g10703(.dina(n10958), .dinb(n10957), .dout(n10959));
  jxor g10704(.dina(b63 ), .dinb(n10637), .dout(n10960));
  jxor g10705(.dina(n10960), .dinb(n10959), .dout(n10961));
  jor  g10706(.dina(n10961), .dinb(n264), .dout(n10962));
  jor  g10707(.dina(n284), .dinb(n10314), .dout(n10963));
  jnot g10708(.din(b63 ), .dout(n10964));
  jor  g10709(.dina(n269), .dinb(n10964), .dout(n10965));
  jor  g10710(.dina(n271), .dinb(n10637), .dout(n10966));
  jand g10711(.dina(n10966), .dinb(n10965), .dout(n10967));
  jand g10712(.dina(n10967), .dinb(n10963), .dout(n10968));
  jand g10713(.dina(n10968), .dinb(n10962), .dout(n10969));
  jxor g10714(.dina(n10969), .dinb(a2 ), .dout(n10970));
  jxor g10715(.dina(n10970), .dinb(n10956), .dout(n10971));
  jxor g10716(.dina(n10971), .dinb(n10660), .dout(n10972));
  jxor g10717(.dina(n10972), .dinb(n10657), .dout(f63 ));
  jand g10718(.dina(n10971), .dinb(n10660), .dout(n10974));
  jand g10719(.dina(n10972), .dinb(n10657), .dout(n10975));
  jor  g10720(.dina(n10975), .dinb(n10974), .dout(n10976));
  jxor g10721(.dina(n10959), .dinb(b62 ), .dout(n10977));
  jor  g10722(.dina(n10977), .dinb(n10960), .dout(n10978));
  jor  g10723(.dina(n10978), .dinb(n264), .dout(n10979));
  jor  g10724(.dina(n284), .dinb(n10637), .dout(n10980));
  jor  g10725(.dina(n271), .dinb(n10964), .dout(n10981));
  jand g10726(.dina(n10981), .dinb(n10980), .dout(n10982));
  jand g10727(.dina(n10982), .dinb(n10979), .dout(n10983));
  jxor g10728(.dina(n10983), .dinb(n260), .dout(n10984));
  jor  g10729(.dina(n10945), .dinb(n10937), .dout(n10985));
  jnot g10730(.din(n10985), .dout(n10986));
  jand g10731(.dina(n10946), .dinb(n10668), .dout(n10987));
  jor  g10732(.dina(n10987), .dinb(n10986), .dout(n10988));
  jor  g10733(.dina(n10311), .dinb(n402), .dout(n10989));
  jor  g10734(.dina(n371), .dinb(n9413), .dout(n10990));
  jor  g10735(.dina(n405), .dinb(n9725), .dout(n10991));
  jor  g10736(.dina(n332), .dinb(n10314), .dout(n10992));
  jand g10737(.dina(n10992), .dinb(n10991), .dout(n10993));
  jand g10738(.dina(n10993), .dinb(n10990), .dout(n10994));
  jand g10739(.dina(n10994), .dinb(n10989), .dout(n10995));
  jxor g10740(.dina(n10995), .dinb(n364), .dout(n10996));
  jor  g10741(.dina(n10935), .dinb(n10927), .dout(n10997));
  jnot g10742(.din(n10936), .dout(n10998));
  jor  g10743(.dina(n10998), .dinb(n10674), .dout(n10999));
  jand g10744(.dina(n10999), .dinb(n10997), .dout(n11000));
  jor  g10745(.dina(n8228), .dinb(n706), .dout(n11001));
  jor  g10746(.dina(n683), .dinb(n7683), .dout(n11002));
  jor  g10747(.dina(n709), .dinb(n7960), .dout(n11003));
  jor  g10748(.dina(n711), .dinb(n8231), .dout(n11004));
  jand g10749(.dina(n11004), .dinb(n11003), .dout(n11005));
  jand g10750(.dina(n11005), .dinb(n11002), .dout(n11006));
  jand g10751(.dina(n11006), .dinb(n11001), .dout(n11007));
  jxor g10752(.dina(n11007), .dinb(a11 ), .dout(n11008));
  jnot g10753(.din(n11008), .dout(n11009));
  jand g10754(.dina(n10924), .dinb(n10686), .dout(n11010));
  jand g10755(.dina(n10925), .dinb(n10677), .dout(n11011));
  jor  g10756(.dina(n11011), .dinb(n11010), .dout(n11012));
  jor  g10757(.dina(n7408), .dinb(n974), .dout(n11013));
  jor  g10758(.dina(n908), .dinb(n7129), .dout(n11014));
  jor  g10759(.dina(n977), .dinb(n7149), .dout(n11015));
  jor  g10760(.dina(n979), .dinb(n7411), .dout(n11016));
  jand g10761(.dina(n11016), .dinb(n11015), .dout(n11017));
  jand g10762(.dina(n11017), .dinb(n11014), .dout(n11018));
  jand g10763(.dina(n11018), .dinb(n11013), .dout(n11019));
  jxor g10764(.dina(n11019), .dinb(a14 ), .dout(n11020));
  jnot g10765(.din(n11020), .dout(n11021));
  jand g10766(.dina(n10922), .dinb(n10698), .dout(n11022));
  jand g10767(.dina(n10923), .dinb(n10689), .dout(n11023));
  jor  g10768(.dina(n11023), .dinb(n11022), .dout(n11024));
  jor  g10769(.dina(n6864), .dinb(n1245), .dout(n11025));
  jor  g10770(.dina(n1165), .dinb(n6352), .dout(n11026));
  jor  g10771(.dina(n1248), .dinb(n6372), .dout(n11027));
  jor  g10772(.dina(n1250), .dinb(n6867), .dout(n11028));
  jand g10773(.dina(n11028), .dinb(n11027), .dout(n11029));
  jand g10774(.dina(n11029), .dinb(n11026), .dout(n11030));
  jand g10775(.dina(n11030), .dinb(n11025), .dout(n11031));
  jxor g10776(.dina(n11031), .dinb(a17 ), .dout(n11032));
  jnot g10777(.din(n11032), .dout(n11033));
  jand g10778(.dina(n10920), .dinb(n10710), .dout(n11034));
  jand g10779(.dina(n10921), .dinb(n10701), .dout(n11035));
  jor  g10780(.dina(n11035), .dinb(n11034), .dout(n11036));
  jor  g10781(.dina(n6103), .dinb(n1566), .dout(n11037));
  jor  g10782(.dina(n1489), .dinb(n5428), .dout(n11038));
  jor  g10783(.dina(n1569), .dinb(n5862), .dout(n11039));
  jor  g10784(.dina(n1571), .dinb(n6106), .dout(n11040));
  jand g10785(.dina(n11040), .dinb(n11039), .dout(n11041));
  jand g10786(.dina(n11041), .dinb(n11038), .dout(n11042));
  jand g10787(.dina(n11042), .dinb(n11037), .dout(n11043));
  jxor g10788(.dina(n11043), .dinb(a20 ), .dout(n11044));
  jnot g10789(.din(n11044), .dout(n11045));
  jand g10790(.dina(n10918), .dinb(n10723), .dout(n11046));
  jand g10791(.dina(n10919), .dinb(n10714), .dout(n11047));
  jor  g10792(.dina(n11047), .dinb(n11046), .dout(n11048));
  jor  g10793(.dina(n5405), .dinb(n1939), .dout(n11049));
  jor  g10794(.dina(n1827), .dinb(n4974), .dout(n11050));
  jor  g10795(.dina(n1942), .dinb(n4994), .dout(n11051));
  jor  g10796(.dina(n1944), .dinb(n5408), .dout(n11052));
  jand g10797(.dina(n11052), .dinb(n11051), .dout(n11053));
  jand g10798(.dina(n11053), .dinb(n11050), .dout(n11054));
  jand g10799(.dina(n11054), .dinb(n11049), .dout(n11055));
  jxor g10800(.dina(n11055), .dinb(a23 ), .dout(n11056));
  jnot g10801(.din(n11056), .dout(n11057));
  jor  g10802(.dina(n10916), .dinb(n10908), .dout(n11058));
  jnot g10803(.din(n11058), .dout(n11059));
  jand g10804(.dina(n10917), .dinb(n10727), .dout(n11060));
  jor  g10805(.dina(n11060), .dinb(n11059), .dout(n11061));
  jand g10806(.dina(n10906), .dinb(n10740), .dout(n11062));
  jnot g10807(.din(n11062), .dout(n11063));
  jnot g10808(.din(n10907), .dout(n11064));
  jor  g10809(.dina(n11064), .dinb(n10731), .dout(n11065));
  jand g10810(.dina(n11065), .dinb(n11063), .dout(n11066));
  jor  g10811(.dina(n10904), .dinb(n10896), .dout(n11067));
  jand g10812(.dina(n10905), .dinb(n10745), .dout(n11068));
  jnot g10813(.din(n11068), .dout(n11069));
  jand g10814(.dina(n11069), .dinb(n11067), .dout(n11070));
  jor  g10815(.dina(n10877), .dinb(n10869), .dout(n11071));
  jand g10816(.dina(n10878), .dinb(n10750), .dout(n11072));
  jnot g10817(.din(n11072), .dout(n11073));
  jand g10818(.dina(n11073), .dinb(n11071), .dout(n11074));
  jnot g10819(.din(n11074), .dout(n11075));
  jor  g10820(.dina(n10866), .dinb(n10858), .dout(n11076));
  jand g10821(.dina(n10867), .dinb(n10753), .dout(n11077));
  jnot g10822(.din(n11077), .dout(n11078));
  jand g10823(.dina(n11078), .dinb(n11076), .dout(n11079));
  jnot g10824(.din(n11079), .dout(n11080));
  jand g10825(.dina(n10855), .dinb(n10765), .dout(n11081));
  jand g10826(.dina(n10856), .dinb(n10756), .dout(n11082));
  jor  g10827(.dina(n11082), .dinb(n11081), .dout(n11083));
  jor  g10828(.dina(n10842), .dinb(n10834), .dout(n11084));
  jand g10829(.dina(n10843), .dinb(n10773), .dout(n11085));
  jnot g10830(.din(n11085), .dout(n11086));
  jand g10831(.dina(n11086), .dinb(n11084), .dout(n11087));
  jnot g10832(.din(n11087), .dout(n11088));
  jor  g10833(.dina(n10829), .dinb(n10821), .dout(n11089));
  jand g10834(.dina(n10830), .dinb(n10788), .dout(n11090));
  jnot g10835(.din(n11090), .dout(n11091));
  jand g10836(.dina(n11091), .dinb(n11089), .dout(n11092));
  jnot g10837(.din(n11092), .dout(n11093));
  jand g10838(.dina(n10818), .dinb(n10800), .dout(n11094));
  jand g10839(.dina(n10819), .dinb(n10791), .dout(n11095));
  jor  g10840(.dina(n11095), .dinb(n11094), .dout(n11096));
  jor  g10841(.dina(n10806), .dinb(n319), .dout(n11097));
  jor  g10842(.dina(n10485), .dinb(n279), .dout(n11098));
  jor  g10843(.dina(n10809), .dinb(n299), .dout(n11099));
  jor  g10844(.dina(n10811), .dinb(n322), .dout(n11100));
  jand g10845(.dina(n11100), .dinb(n11099), .dout(n11101));
  jand g10846(.dina(n11101), .dinb(n11098), .dout(n11102));
  jand g10847(.dina(n11102), .dinb(n11097), .dout(n11103));
  jxor g10848(.dina(n11103), .dinb(a62 ), .dout(n11104));
  jnot g10849(.din(n11104), .dout(n11105));
  jand g10850(.dina(n10801), .dinb(b1 ), .dout(n11106));
  jand g10851(.dina(a63 ), .dinb(a62 ), .dout(n11107));
  jand g10852(.dina(n11107), .dinb(b0 ), .dout(n11108));
  jor  g10853(.dina(n11108), .dinb(n11106), .dout(n11109));
  jxor g10854(.dina(n11109), .dinb(n11105), .dout(n11110));
  jand g10855(.dina(n10804), .dinb(n10803), .dout(n11111));
  jnot g10856(.din(n11111), .dout(n11112));
  jand g10857(.dina(n10817), .dinb(n11112), .dout(n11116));
  jxor g10858(.dina(n11116), .dinb(n11110), .dout(n11117));
  jnot g10859(.din(n11117), .dout(n11118));
  jor  g10860(.dina(n9891), .dinb(n428), .dout(n11119));
  jor  g10861(.dina(n9593), .dinb(n357), .dout(n11120));
  jor  g10862(.dina(n9894), .dinb(n395), .dout(n11121));
  jor  g10863(.dina(n9896), .dinb(n431), .dout(n11122));
  jand g10864(.dina(n11122), .dinb(n11121), .dout(n11123));
  jand g10865(.dina(n11123), .dinb(n11120), .dout(n11124));
  jand g10866(.dina(n11124), .dinb(n11119), .dout(n11125));
  jxor g10867(.dina(n11125), .dinb(a59 ), .dout(n11126));
  jxor g10868(.dina(n11126), .dinb(n11118), .dout(n11127));
  jxor g10869(.dina(n11127), .dinb(n11096), .dout(n11128));
  jnot g10870(.din(n11128), .dout(n11129));
  jor  g10871(.dina(n8978), .dinb(n624), .dout(n11130));
  jor  g10872(.dina(n8677), .dinb(n512), .dout(n11131));
  jor  g10873(.dina(n8981), .dinb(n564), .dout(n11132));
  jor  g10874(.dina(n8983), .dinb(n627), .dout(n11133));
  jand g10875(.dina(n11133), .dinb(n11132), .dout(n11134));
  jand g10876(.dina(n11134), .dinb(n11131), .dout(n11135));
  jand g10877(.dina(n11135), .dinb(n11130), .dout(n11136));
  jxor g10878(.dina(n11136), .dinb(a56 ), .dout(n11137));
  jxor g10879(.dina(n11137), .dinb(n11129), .dout(n11138));
  jxor g10880(.dina(n11138), .dinb(n11093), .dout(n11139));
  jnot g10881(.din(n11139), .dout(n11140));
  jor  g10882(.dina(n8125), .dinb(n775), .dout(n11141));
  jor  g10883(.dina(n7846), .dinb(n647), .dout(n11142));
  jor  g10884(.dina(n8128), .dinb(n758), .dout(n11143));
  jor  g10885(.dina(n8130), .dinb(n778), .dout(n11144));
  jand g10886(.dina(n11144), .dinb(n11143), .dout(n11145));
  jand g10887(.dina(n11145), .dinb(n11142), .dout(n11146));
  jand g10888(.dina(n11146), .dinb(n11141), .dout(n11147));
  jxor g10889(.dina(n11147), .dinb(a53 ), .dout(n11148));
  jxor g10890(.dina(n11148), .dinb(n11140), .dout(n11149));
  jand g10891(.dina(n10831), .dinb(n10785), .dout(n11150));
  jand g10892(.dina(n10832), .dinb(n10776), .dout(n11151));
  jor  g10893(.dina(n11151), .dinb(n11150), .dout(n11152));
  jxor g10894(.dina(n11152), .dinb(n11149), .dout(n11153));
  jnot g10895(.din(n11153), .dout(n11154));
  jor  g10896(.dina(n7266), .dinb(n1019), .dout(n11155));
  jor  g10897(.dina(n7021), .dinb(n858), .dout(n11156));
  jor  g10898(.dina(n7269), .dinb(n939), .dout(n11157));
  jor  g10899(.dina(n7271), .dinb(n1022), .dout(n11158));
  jand g10900(.dina(n11158), .dinb(n11157), .dout(n11159));
  jand g10901(.dina(n11159), .dinb(n11156), .dout(n11160));
  jand g10902(.dina(n11160), .dinb(n11155), .dout(n11161));
  jxor g10903(.dina(n11161), .dinb(a50 ), .dout(n11162));
  jxor g10904(.dina(n11162), .dinb(n11154), .dout(n11163));
  jxor g10905(.dina(n11163), .dinb(n11088), .dout(n11164));
  jnot g10906(.din(n11164), .dout(n11165));
  jor  g10907(.dina(n6490), .dinb(n1397), .dout(n11166));
  jor  g10908(.dina(n6262), .dinb(n1193), .dout(n11167));
  jor  g10909(.dina(n6493), .dinb(n1290), .dout(n11168));
  jor  g10910(.dina(n6495), .dinb(n1400), .dout(n11169));
  jand g10911(.dina(n11169), .dinb(n11168), .dout(n11170));
  jand g10912(.dina(n11170), .dinb(n11167), .dout(n11171));
  jand g10913(.dina(n11171), .dinb(n11166), .dout(n11172));
  jxor g10914(.dina(n11172), .dinb(a47 ), .dout(n11173));
  jxor g10915(.dina(n11173), .dinb(n11165), .dout(n11174));
  jnot g10916(.din(n11174), .dout(n11175));
  jor  g10917(.dina(n10853), .dinb(n10845), .dout(n11176));
  jand g10918(.dina(n10854), .dinb(n10768), .dout(n11177));
  jnot g10919(.din(n11177), .dout(n11178));
  jand g10920(.dina(n11178), .dinb(n11176), .dout(n11179));
  jxor g10921(.dina(n11179), .dinb(n11175), .dout(n11180));
  jnot g10922(.din(n11180), .dout(n11181));
  jor  g10923(.dina(n5739), .dinb(n1739), .dout(n11182));
  jor  g10924(.dina(n5574), .dinb(n1420), .dout(n11183));
  jor  g10925(.dina(n5742), .dinb(n1620), .dout(n11184));
  jor  g10926(.dina(n5744), .dinb(n1742), .dout(n11185));
  jand g10927(.dina(n11185), .dinb(n11184), .dout(n11186));
  jand g10928(.dina(n11186), .dinb(n11183), .dout(n11187));
  jand g10929(.dina(n11187), .dinb(n11182), .dout(n11188));
  jxor g10930(.dina(n11188), .dinb(a44 ), .dout(n11189));
  jxor g10931(.dina(n11189), .dinb(n11181), .dout(n11190));
  jxor g10932(.dina(n11190), .dinb(n11083), .dout(n11191));
  jnot g10933(.din(n11191), .dout(n11192));
  jor  g10934(.dina(n5096), .dinb(n2007), .dout(n11193));
  jor  g10935(.dina(n4904), .dinb(n1867), .dout(n11194));
  jor  g10936(.dina(n5099), .dinb(n1887), .dout(n11195));
  jor  g10937(.dina(n5101), .dinb(n2010), .dout(n11196));
  jand g10938(.dina(n11196), .dinb(n11195), .dout(n11197));
  jand g10939(.dina(n11197), .dinb(n11194), .dout(n11198));
  jand g10940(.dina(n11198), .dinb(n11193), .dout(n11199));
  jxor g10941(.dina(n11199), .dinb(a41 ), .dout(n11200));
  jxor g10942(.dina(n11200), .dinb(n11192), .dout(n11201));
  jxor g10943(.dina(n11201), .dinb(n11080), .dout(n11202));
  jnot g10944(.din(n11202), .dout(n11203));
  jor  g10945(.dina(n4415), .dinb(n2556), .dout(n11204));
  jor  g10946(.dina(n4272), .dinb(n2148), .dout(n11205));
  jor  g10947(.dina(n4418), .dinb(n2407), .dout(n11206));
  jor  g10948(.dina(n4420), .dinb(n2559), .dout(n11207));
  jand g10949(.dina(n11207), .dinb(n11206), .dout(n11208));
  jand g10950(.dina(n11208), .dinb(n11205), .dout(n11209));
  jand g10951(.dina(n11209), .dinb(n11204), .dout(n11210));
  jxor g10952(.dina(n11210), .dinb(a38 ), .dout(n11211));
  jxor g10953(.dina(n11211), .dinb(n11203), .dout(n11212));
  jxor g10954(.dina(n11212), .dinb(n11075), .dout(n11213));
  jnot g10955(.din(n11213), .dout(n11214));
  jor  g10956(.dina(n3849), .dinb(n3032), .dout(n11215));
  jor  g10957(.dina(n3689), .dinb(n2579), .dout(n11216));
  jor  g10958(.dina(n3852), .dinb(n2870), .dout(n11217));
  jor  g10959(.dina(n3854), .dinb(n3035), .dout(n11218));
  jand g10960(.dina(n11218), .dinb(n11217), .dout(n11219));
  jand g10961(.dina(n11219), .dinb(n11216), .dout(n11220));
  jand g10962(.dina(n11220), .dinb(n11215), .dout(n11221));
  jxor g10963(.dina(n11221), .dinb(a35 ), .dout(n11222));
  jxor g10964(.dina(n11222), .dinb(n11214), .dout(n11223));
  jnot g10965(.din(n11223), .dout(n11224));
  jor  g10966(.dina(n10888), .dinb(n10880), .dout(n11225));
  jor  g10967(.dina(n10894), .dinb(n10890), .dout(n11226));
  jand g10968(.dina(n11226), .dinb(n11225), .dout(n11227));
  jxor g10969(.dina(n11227), .dinb(n11224), .dout(n11228));
  jnot g10970(.din(n11228), .dout(n11229));
  jor  g10971(.dina(n3400), .dinb(n3301), .dout(n11230));
  jor  g10972(.dina(n3136), .dinb(n3055), .dout(n11231));
  jor  g10973(.dina(n3304), .dinb(n3230), .dout(n11232));
  jor  g10974(.dina(n3306), .dinb(n3403), .dout(n11233));
  jand g10975(.dina(n11233), .dinb(n11232), .dout(n11234));
  jand g10976(.dina(n11234), .dinb(n11231), .dout(n11235));
  jand g10977(.dina(n11235), .dinb(n11230), .dout(n11236));
  jxor g10978(.dina(n11236), .dinb(a32 ), .dout(n11237));
  jxor g10979(.dina(n11237), .dinb(n11229), .dout(n11238));
  jxor g10980(.dina(n11238), .dinb(n11070), .dout(n11239));
  jor  g10981(.dina(n4137), .dinb(n2784), .dout(n11240));
  jor  g10982(.dina(n2661), .dinb(n3588), .dout(n11241));
  jor  g10983(.dina(n2787), .dinb(n3942), .dout(n11242));
  jor  g10984(.dina(n2789), .dinb(n4140), .dout(n11243));
  jand g10985(.dina(n11243), .dinb(n11242), .dout(n11244));
  jand g10986(.dina(n11244), .dinb(n11241), .dout(n11245));
  jand g10987(.dina(n11245), .dinb(n11240), .dout(n11246));
  jxor g10988(.dina(n11246), .dinb(a29 ), .dout(n11247));
  jxor g10989(.dina(n11247), .dinb(n11239), .dout(n11248));
  jxor g10990(.dina(n11248), .dinb(n11066), .dout(n11249));
  jor  g10991(.dina(n4554), .dinb(n2319), .dout(n11250));
  jor  g10992(.dina(n2224), .dinb(n4340), .dout(n11251));
  jor  g10993(.dina(n2322), .dinb(n4537), .dout(n11252));
  jor  g10994(.dina(n2324), .dinb(n4557), .dout(n11253));
  jand g10995(.dina(n11253), .dinb(n11252), .dout(n11254));
  jand g10996(.dina(n11254), .dinb(n11251), .dout(n11255));
  jand g10997(.dina(n11255), .dinb(n11250), .dout(n11256));
  jxor g10998(.dina(n11256), .dinb(a26 ), .dout(n11257));
  jxor g10999(.dina(n11257), .dinb(n11249), .dout(n11258));
  jxor g11000(.dina(n11258), .dinb(n11061), .dout(n11259));
  jxor g11001(.dina(n11259), .dinb(n11057), .dout(n11260));
  jxor g11002(.dina(n11260), .dinb(n11048), .dout(n11261));
  jxor g11003(.dina(n11261), .dinb(n11045), .dout(n11262));
  jxor g11004(.dina(n11262), .dinb(n11036), .dout(n11263));
  jxor g11005(.dina(n11263), .dinb(n11033), .dout(n11264));
  jxor g11006(.dina(n11264), .dinb(n11024), .dout(n11265));
  jxor g11007(.dina(n11265), .dinb(n11021), .dout(n11266));
  jxor g11008(.dina(n11266), .dinb(n11012), .dout(n11267));
  jxor g11009(.dina(n11267), .dinb(n11009), .dout(n11268));
  jxor g11010(.dina(n11268), .dinb(n11000), .dout(n11269));
  jor  g11011(.dina(n9387), .dinb(n528), .dout(n11270));
  jor  g11012(.dina(n490), .dinb(n8789), .dout(n11271));
  jor  g11013(.dina(n531), .dinb(n8809), .dout(n11272));
  jor  g11014(.dina(n533), .dinb(n9390), .dout(n11273));
  jand g11015(.dina(n11273), .dinb(n11272), .dout(n11274));
  jand g11016(.dina(n11274), .dinb(n11271), .dout(n11275));
  jand g11017(.dina(n11275), .dinb(n11270), .dout(n11276));
  jxor g11018(.dina(n11276), .dinb(a8 ), .dout(n11277));
  jxor g11019(.dina(n11277), .dinb(n11269), .dout(n11278));
  jxor g11020(.dina(n11278), .dinb(n10996), .dout(n11279));
  jxor g11021(.dina(n11279), .dinb(n10988), .dout(n11280));
  jxor g11022(.dina(n11280), .dinb(n10984), .dout(n11281));
  jnot g11023(.din(n10953), .dout(n11282));
  jxor g11024(.dina(n10969), .dinb(n260), .dout(n11283));
  jand g11025(.dina(n11283), .dinb(n11282), .dout(n11284));
  jor  g11026(.dina(n11284), .dinb(n10955), .dout(n11285));
  jxor g11027(.dina(n11285), .dinb(n11281), .dout(n11286));
  jxor g11028(.dina(n11286), .dinb(n10976), .dout(f64 ));
  jand g11029(.dina(n11279), .dinb(n10988), .dout(n11288));
  jand g11030(.dina(n11280), .dinb(n10984), .dout(n11289));
  jor  g11031(.dina(n11289), .dinb(n11288), .dout(n11290));
  jor  g11032(.dina(n11277), .dinb(n11269), .dout(n11291));
  jand g11033(.dina(n11278), .dinb(n10996), .dout(n11292));
  jnot g11034(.din(n11292), .dout(n11293));
  jand g11035(.dina(n11293), .dinb(n11291), .dout(n11294));
  jnot g11036(.din(n11294), .dout(n11295));
  jor  g11037(.dina(n10959), .dinb(b62 ), .dout(n11296));
  jor  g11038(.dina(n264), .dinb(n10964), .dout(n11297));
  jnot g11039(.din(n11297), .dout(n11298));
  jand g11040(.dina(n11298), .dinb(n11296), .dout(n11299));
  jnot g11041(.din(n11299), .dout(n11300));
  jor  g11042(.dina(n284), .dinb(n10964), .dout(n11301));
  jand g11043(.dina(n11301), .dinb(a2 ), .dout(n11302));
  jand g11044(.dina(n11302), .dinb(n11300), .dout(n11303));
  jand g11045(.dina(n11299), .dinb(n260), .dout(n11304));
  jor  g11046(.dina(n11304), .dinb(n11303), .dout(n11305));
  jxor g11047(.dina(n11305), .dinb(n11295), .dout(n11306));
  jand g11048(.dina(n11267), .dinb(n11009), .dout(n11307));
  jnot g11049(.din(n11000), .dout(n11308));
  jand g11050(.dina(n11268), .dinb(n11308), .dout(n11309));
  jor  g11051(.dina(n11309), .dinb(n11307), .dout(n11310));
  jnot g11052(.din(n11310), .dout(n11311));
  jand g11053(.dina(n11265), .dinb(n11021), .dout(n11312));
  jand g11054(.dina(n11266), .dinb(n11012), .dout(n11313));
  jor  g11055(.dina(n11313), .dinb(n11312), .dout(n11314));
  jand g11056(.dina(n11263), .dinb(n11033), .dout(n11315));
  jand g11057(.dina(n11264), .dinb(n11024), .dout(n11316));
  jor  g11058(.dina(n11316), .dinb(n11315), .dout(n11317));
  jnot g11059(.din(n11317), .dout(n11318));
  jor  g11060(.dina(n7126), .dinb(n1245), .dout(n11319));
  jor  g11061(.dina(n1165), .dinb(n6372), .dout(n11320));
  jor  g11062(.dina(n1248), .dinb(n6867), .dout(n11321));
  jor  g11063(.dina(n1250), .dinb(n7129), .dout(n11322));
  jand g11064(.dina(n11322), .dinb(n11321), .dout(n11323));
  jand g11065(.dina(n11323), .dinb(n11320), .dout(n11324));
  jand g11066(.dina(n11324), .dinb(n11319), .dout(n11325));
  jxor g11067(.dina(n11325), .dinb(a17 ), .dout(n11326));
  jnot g11068(.din(n11326), .dout(n11327));
  jand g11069(.dina(n11261), .dinb(n11045), .dout(n11328));
  jand g11070(.dina(n11262), .dinb(n11036), .dout(n11329));
  jor  g11071(.dina(n11329), .dinb(n11328), .dout(n11330));
  jor  g11072(.dina(n6349), .dinb(n1566), .dout(n11331));
  jor  g11073(.dina(n1489), .dinb(n5862), .dout(n11332));
  jor  g11074(.dina(n1569), .dinb(n6106), .dout(n11333));
  jor  g11075(.dina(n1571), .dinb(n6352), .dout(n11334));
  jand g11076(.dina(n11334), .dinb(n11333), .dout(n11335));
  jand g11077(.dina(n11335), .dinb(n11332), .dout(n11336));
  jand g11078(.dina(n11336), .dinb(n11331), .dout(n11337));
  jxor g11079(.dina(n11337), .dinb(a20 ), .dout(n11338));
  jnot g11080(.din(n11338), .dout(n11339));
  jand g11081(.dina(n11259), .dinb(n11057), .dout(n11340));
  jand g11082(.dina(n11260), .dinb(n11048), .dout(n11341));
  jor  g11083(.dina(n11341), .dinb(n11340), .dout(n11342));
  jor  g11084(.dina(n11257), .dinb(n11249), .dout(n11343));
  jand g11085(.dina(n11258), .dinb(n11061), .dout(n11344));
  jnot g11086(.din(n11344), .dout(n11345));
  jand g11087(.dina(n11345), .dinb(n11343), .dout(n11346));
  jor  g11088(.dina(n11247), .dinb(n11239), .dout(n11347));
  jnot g11089(.din(n11248), .dout(n11348));
  jor  g11090(.dina(n11348), .dinb(n11066), .dout(n11349));
  jand g11091(.dina(n11349), .dinb(n11347), .dout(n11350));
  jor  g11092(.dina(n11237), .dinb(n11229), .dout(n11351));
  jnot g11093(.din(n11238), .dout(n11352));
  jor  g11094(.dina(n11352), .dinb(n11070), .dout(n11353));
  jand g11095(.dina(n11353), .dinb(n11351), .dout(n11354));
  jor  g11096(.dina(n11222), .dinb(n11214), .dout(n11355));
  jor  g11097(.dina(n11227), .dinb(n11224), .dout(n11356));
  jand g11098(.dina(n11356), .dinb(n11355), .dout(n11357));
  jnot g11099(.din(n11357), .dout(n11358));
  jor  g11100(.dina(n11211), .dinb(n11203), .dout(n11359));
  jand g11101(.dina(n11212), .dinb(n11075), .dout(n11360));
  jnot g11102(.din(n11360), .dout(n11361));
  jand g11103(.dina(n11361), .dinb(n11359), .dout(n11362));
  jnot g11104(.din(n11362), .dout(n11363));
  jor  g11105(.dina(n11200), .dinb(n11192), .dout(n11364));
  jand g11106(.dina(n11201), .dinb(n11080), .dout(n11365));
  jnot g11107(.din(n11365), .dout(n11366));
  jand g11108(.dina(n11366), .dinb(n11364), .dout(n11367));
  jnot g11109(.din(n11367), .dout(n11368));
  jor  g11110(.dina(n11189), .dinb(n11181), .dout(n11369));
  jand g11111(.dina(n11190), .dinb(n11083), .dout(n11370));
  jnot g11112(.din(n11370), .dout(n11371));
  jand g11113(.dina(n11371), .dinb(n11369), .dout(n11372));
  jnot g11114(.din(n11372), .dout(n11373));
  jor  g11115(.dina(n5739), .dinb(n1864), .dout(n11374));
  jor  g11116(.dina(n5574), .dinb(n1620), .dout(n11375));
  jor  g11117(.dina(n5742), .dinb(n1742), .dout(n11376));
  jor  g11118(.dina(n5744), .dinb(n1867), .dout(n11377));
  jand g11119(.dina(n11377), .dinb(n11376), .dout(n11378));
  jand g11120(.dina(n11378), .dinb(n11375), .dout(n11379));
  jand g11121(.dina(n11379), .dinb(n11374), .dout(n11380));
  jxor g11122(.dina(n11380), .dinb(a44 ), .dout(n11381));
  jnot g11123(.din(n11381), .dout(n11382));
  jor  g11124(.dina(n11173), .dinb(n11165), .dout(n11383));
  jor  g11125(.dina(n11179), .dinb(n11175), .dout(n11384));
  jand g11126(.dina(n11384), .dinb(n11383), .dout(n11385));
  jnot g11127(.din(n11385), .dout(n11386));
  jor  g11128(.dina(n11162), .dinb(n11154), .dout(n11387));
  jand g11129(.dina(n11163), .dinb(n11088), .dout(n11388));
  jnot g11130(.din(n11388), .dout(n11389));
  jand g11131(.dina(n11389), .dinb(n11387), .dout(n11390));
  jnot g11132(.din(n11390), .dout(n11391));
  jor  g11133(.dina(n7266), .dinb(n1190), .dout(n11392));
  jor  g11134(.dina(n7021), .dinb(n939), .dout(n11393));
  jor  g11135(.dina(n7269), .dinb(n1022), .dout(n11394));
  jor  g11136(.dina(n7271), .dinb(n1193), .dout(n11395));
  jand g11137(.dina(n11395), .dinb(n11394), .dout(n11396));
  jand g11138(.dina(n11396), .dinb(n11393), .dout(n11397));
  jand g11139(.dina(n11397), .dinb(n11392), .dout(n11398));
  jxor g11140(.dina(n11398), .dinb(a50 ), .dout(n11399));
  jnot g11141(.din(n11399), .dout(n11400));
  jor  g11142(.dina(n11148), .dinb(n11140), .dout(n11401));
  jand g11143(.dina(n11152), .dinb(n11149), .dout(n11402));
  jnot g11144(.din(n11402), .dout(n11403));
  jand g11145(.dina(n11403), .dinb(n11401), .dout(n11404));
  jnot g11146(.din(n11404), .dout(n11405));
  jor  g11147(.dina(n11137), .dinb(n11129), .dout(n11406));
  jand g11148(.dina(n11138), .dinb(n11093), .dout(n11407));
  jnot g11149(.din(n11407), .dout(n11408));
  jand g11150(.dina(n11408), .dinb(n11406), .dout(n11409));
  jnot g11151(.din(n11409), .dout(n11410));
  jor  g11152(.dina(n8978), .dinb(n644), .dout(n11411));
  jor  g11153(.dina(n8677), .dinb(n564), .dout(n11412));
  jor  g11154(.dina(n8981), .dinb(n627), .dout(n11413));
  jor  g11155(.dina(n8983), .dinb(n647), .dout(n11414));
  jand g11156(.dina(n11414), .dinb(n11413), .dout(n11415));
  jand g11157(.dina(n11415), .dinb(n11412), .dout(n11416));
  jand g11158(.dina(n11416), .dinb(n11411), .dout(n11417));
  jxor g11159(.dina(n11417), .dinb(a56 ), .dout(n11418));
  jnot g11160(.din(n11418), .dout(n11419));
  jor  g11161(.dina(n11126), .dinb(n11118), .dout(n11420));
  jand g11162(.dina(n11127), .dinb(n11096), .dout(n11421));
  jnot g11163(.din(n11421), .dout(n11422));
  jand g11164(.dina(n11422), .dinb(n11420), .dout(n11423));
  jnot g11165(.din(n11423), .dout(n11424));
  jand g11166(.dina(n11109), .dinb(n11105), .dout(n11425));
  jand g11167(.dina(n11116), .dinb(n11110), .dout(n11426));
  jor  g11168(.dina(n11426), .dinb(n11425), .dout(n11427));
  jor  g11169(.dina(n10806), .dinb(n354), .dout(n11428));
  jor  g11170(.dina(n10485), .dinb(n299), .dout(n11429));
  jor  g11171(.dina(n10809), .dinb(n322), .dout(n11430));
  jor  g11172(.dina(n10811), .dinb(n357), .dout(n11431));
  jand g11173(.dina(n11431), .dinb(n11430), .dout(n11432));
  jand g11174(.dina(n11432), .dinb(n11429), .dout(n11433));
  jand g11175(.dina(n11433), .dinb(n11428), .dout(n11434));
  jxor g11176(.dina(n11434), .dinb(a62 ), .dout(n11435));
  jnot g11177(.din(n11435), .dout(n11436));
  jand g11178(.dina(n10801), .dinb(b2 ), .dout(n11437));
  jand g11179(.dina(n11107), .dinb(b1 ), .dout(n11438));
  jor  g11180(.dina(n11438), .dinb(n11437), .dout(n11439));
  jxor g11181(.dina(n11439), .dinb(n11436), .dout(n11440));
  jxor g11182(.dina(n11440), .dinb(n11427), .dout(n11441));
  jnot g11183(.din(n11441), .dout(n11442));
  jor  g11184(.dina(n9891), .dinb(n509), .dout(n11443));
  jor  g11185(.dina(n9593), .dinb(n395), .dout(n11444));
  jor  g11186(.dina(n9894), .dinb(n431), .dout(n11445));
  jor  g11187(.dina(n9896), .dinb(n512), .dout(n11446));
  jand g11188(.dina(n11446), .dinb(n11445), .dout(n11447));
  jand g11189(.dina(n11447), .dinb(n11444), .dout(n11448));
  jand g11190(.dina(n11448), .dinb(n11443), .dout(n11449));
  jxor g11191(.dina(n11449), .dinb(a59 ), .dout(n11450));
  jxor g11192(.dina(n11450), .dinb(n11442), .dout(n11451));
  jxor g11193(.dina(n11451), .dinb(n11424), .dout(n11452));
  jxor g11194(.dina(n11452), .dinb(n11419), .dout(n11453));
  jxor g11195(.dina(n11453), .dinb(n11410), .dout(n11454));
  jnot g11196(.din(n11454), .dout(n11455));
  jor  g11197(.dina(n8125), .dinb(n855), .dout(n11456));
  jor  g11198(.dina(n7846), .dinb(n758), .dout(n11457));
  jor  g11199(.dina(n8128), .dinb(n778), .dout(n11458));
  jor  g11200(.dina(n8130), .dinb(n858), .dout(n11459));
  jand g11201(.dina(n11459), .dinb(n11458), .dout(n11460));
  jand g11202(.dina(n11460), .dinb(n11457), .dout(n11461));
  jand g11203(.dina(n11461), .dinb(n11456), .dout(n11462));
  jxor g11204(.dina(n11462), .dinb(a53 ), .dout(n11463));
  jxor g11205(.dina(n11463), .dinb(n11455), .dout(n11464));
  jxor g11206(.dina(n11464), .dinb(n11405), .dout(n11465));
  jxor g11207(.dina(n11465), .dinb(n11400), .dout(n11466));
  jxor g11208(.dina(n11466), .dinb(n11391), .dout(n11467));
  jnot g11209(.din(n11467), .dout(n11468));
  jor  g11210(.dina(n6490), .dinb(n1417), .dout(n11469));
  jor  g11211(.dina(n6262), .dinb(n1290), .dout(n11470));
  jor  g11212(.dina(n6493), .dinb(n1400), .dout(n11471));
  jor  g11213(.dina(n6495), .dinb(n1420), .dout(n11472));
  jand g11214(.dina(n11472), .dinb(n11471), .dout(n11473));
  jand g11215(.dina(n11473), .dinb(n11470), .dout(n11474));
  jand g11216(.dina(n11474), .dinb(n11469), .dout(n11475));
  jxor g11217(.dina(n11475), .dinb(a47 ), .dout(n11476));
  jxor g11218(.dina(n11476), .dinb(n11468), .dout(n11477));
  jxor g11219(.dina(n11477), .dinb(n11386), .dout(n11478));
  jxor g11220(.dina(n11478), .dinb(n11382), .dout(n11479));
  jxor g11221(.dina(n11479), .dinb(n11373), .dout(n11480));
  jnot g11222(.din(n11480), .dout(n11481));
  jor  g11223(.dina(n5096), .dinb(n2145), .dout(n11482));
  jor  g11224(.dina(n4904), .dinb(n1887), .dout(n11483));
  jor  g11225(.dina(n5099), .dinb(n2010), .dout(n11484));
  jor  g11226(.dina(n5101), .dinb(n2148), .dout(n11485));
  jand g11227(.dina(n11485), .dinb(n11484), .dout(n11486));
  jand g11228(.dina(n11486), .dinb(n11483), .dout(n11487));
  jand g11229(.dina(n11487), .dinb(n11482), .dout(n11488));
  jxor g11230(.dina(n11488), .dinb(a41 ), .dout(n11489));
  jxor g11231(.dina(n11489), .dinb(n11481), .dout(n11490));
  jxor g11232(.dina(n11490), .dinb(n11368), .dout(n11491));
  jnot g11233(.din(n11491), .dout(n11492));
  jor  g11234(.dina(n4415), .dinb(n2576), .dout(n11493));
  jor  g11235(.dina(n4272), .dinb(n2407), .dout(n11494));
  jor  g11236(.dina(n4418), .dinb(n2559), .dout(n11495));
  jor  g11237(.dina(n4420), .dinb(n2579), .dout(n11496));
  jand g11238(.dina(n11496), .dinb(n11495), .dout(n11497));
  jand g11239(.dina(n11497), .dinb(n11494), .dout(n11498));
  jand g11240(.dina(n11498), .dinb(n11493), .dout(n11499));
  jxor g11241(.dina(n11499), .dinb(a38 ), .dout(n11500));
  jxor g11242(.dina(n11500), .dinb(n11492), .dout(n11501));
  jxor g11243(.dina(n11501), .dinb(n11363), .dout(n11502));
  jnot g11244(.din(n11502), .dout(n11503));
  jor  g11245(.dina(n3849), .dinb(n3052), .dout(n11504));
  jor  g11246(.dina(n3689), .dinb(n2870), .dout(n11505));
  jor  g11247(.dina(n3852), .dinb(n3035), .dout(n11506));
  jor  g11248(.dina(n3854), .dinb(n3055), .dout(n11507));
  jand g11249(.dina(n11507), .dinb(n11506), .dout(n11508));
  jand g11250(.dina(n11508), .dinb(n11505), .dout(n11509));
  jand g11251(.dina(n11509), .dinb(n11504), .dout(n11510));
  jxor g11252(.dina(n11510), .dinb(a35 ), .dout(n11511));
  jxor g11253(.dina(n11511), .dinb(n11503), .dout(n11512));
  jxor g11254(.dina(n11512), .dinb(n11358), .dout(n11513));
  jnot g11255(.din(n11513), .dout(n11514));
  jor  g11256(.dina(n3585), .dinb(n3301), .dout(n11515));
  jor  g11257(.dina(n3136), .dinb(n3230), .dout(n11516));
  jor  g11258(.dina(n3304), .dinb(n3403), .dout(n11517));
  jor  g11259(.dina(n3306), .dinb(n3588), .dout(n11518));
  jand g11260(.dina(n11518), .dinb(n11517), .dout(n11519));
  jand g11261(.dina(n11519), .dinb(n11516), .dout(n11520));
  jand g11262(.dina(n11520), .dinb(n11515), .dout(n11521));
  jxor g11263(.dina(n11521), .dinb(a32 ), .dout(n11522));
  jxor g11264(.dina(n11522), .dinb(n11514), .dout(n11523));
  jxor g11265(.dina(n11523), .dinb(n11354), .dout(n11524));
  jor  g11266(.dina(n4337), .dinb(n2784), .dout(n11525));
  jor  g11267(.dina(n2661), .dinb(n3942), .dout(n11526));
  jor  g11268(.dina(n2787), .dinb(n4140), .dout(n11527));
  jor  g11269(.dina(n2789), .dinb(n4340), .dout(n11528));
  jand g11270(.dina(n11528), .dinb(n11527), .dout(n11529));
  jand g11271(.dina(n11529), .dinb(n11526), .dout(n11530));
  jand g11272(.dina(n11530), .dinb(n11525), .dout(n11531));
  jxor g11273(.dina(n11531), .dinb(a29 ), .dout(n11532));
  jxor g11274(.dina(n11532), .dinb(n11524), .dout(n11533));
  jxor g11275(.dina(n11533), .dinb(n11350), .dout(n11534));
  jor  g11276(.dina(n4971), .dinb(n2319), .dout(n11535));
  jor  g11277(.dina(n2224), .dinb(n4537), .dout(n11536));
  jor  g11278(.dina(n2322), .dinb(n4557), .dout(n11537));
  jor  g11279(.dina(n2324), .dinb(n4974), .dout(n11538));
  jand g11280(.dina(n11538), .dinb(n11537), .dout(n11539));
  jand g11281(.dina(n11539), .dinb(n11536), .dout(n11540));
  jand g11282(.dina(n11540), .dinb(n11535), .dout(n11541));
  jxor g11283(.dina(n11541), .dinb(a26 ), .dout(n11542));
  jxor g11284(.dina(n11542), .dinb(n11534), .dout(n11543));
  jxor g11285(.dina(n11543), .dinb(n11346), .dout(n11544));
  jor  g11286(.dina(n5425), .dinb(n1939), .dout(n11545));
  jor  g11287(.dina(n1827), .dinb(n4994), .dout(n11546));
  jor  g11288(.dina(n1942), .dinb(n5408), .dout(n11547));
  jor  g11289(.dina(n1944), .dinb(n5428), .dout(n11548));
  jand g11290(.dina(n11548), .dinb(n11547), .dout(n11549));
  jand g11291(.dina(n11549), .dinb(n11546), .dout(n11550));
  jand g11292(.dina(n11550), .dinb(n11545), .dout(n11551));
  jxor g11293(.dina(n11551), .dinb(a23 ), .dout(n11552));
  jxor g11294(.dina(n11552), .dinb(n11544), .dout(n11553));
  jxor g11295(.dina(n11553), .dinb(n11342), .dout(n11554));
  jxor g11296(.dina(n11554), .dinb(n11339), .dout(n11555));
  jxor g11297(.dina(n11555), .dinb(n11330), .dout(n11556));
  jxor g11298(.dina(n11556), .dinb(n11327), .dout(n11557));
  jxor g11299(.dina(n11557), .dinb(n11318), .dout(n11558));
  jor  g11300(.dina(n7680), .dinb(n974), .dout(n11559));
  jor  g11301(.dina(n908), .dinb(n7149), .dout(n11560));
  jor  g11302(.dina(n977), .dinb(n7411), .dout(n11561));
  jor  g11303(.dina(n979), .dinb(n7683), .dout(n11562));
  jand g11304(.dina(n11562), .dinb(n11561), .dout(n11563));
  jand g11305(.dina(n11563), .dinb(n11560), .dout(n11564));
  jand g11306(.dina(n11564), .dinb(n11559), .dout(n11565));
  jxor g11307(.dina(n11565), .dinb(a14 ), .dout(n11566));
  jxor g11308(.dina(n11566), .dinb(n11558), .dout(n11567));
  jxor g11309(.dina(n11567), .dinb(n11314), .dout(n11568));
  jor  g11310(.dina(n8786), .dinb(n706), .dout(n11569));
  jor  g11311(.dina(n683), .dinb(n7960), .dout(n11570));
  jor  g11312(.dina(n709), .dinb(n8231), .dout(n11571));
  jor  g11313(.dina(n711), .dinb(n8789), .dout(n11572));
  jand g11314(.dina(n11572), .dinb(n11571), .dout(n11573));
  jand g11315(.dina(n11573), .dinb(n11570), .dout(n11574));
  jand g11316(.dina(n11574), .dinb(n11569), .dout(n11575));
  jxor g11317(.dina(n11575), .dinb(a11 ), .dout(n11576));
  jxor g11318(.dina(n11576), .dinb(n11568), .dout(n11577));
  jor  g11319(.dina(n9410), .dinb(n528), .dout(n11578));
  jor  g11320(.dina(n490), .dinb(n8809), .dout(n11579));
  jor  g11321(.dina(n531), .dinb(n9390), .dout(n11580));
  jor  g11322(.dina(n533), .dinb(n9413), .dout(n11581));
  jand g11323(.dina(n11581), .dinb(n11580), .dout(n11582));
  jand g11324(.dina(n11582), .dinb(n11579), .dout(n11583));
  jand g11325(.dina(n11583), .dinb(n11578), .dout(n11584));
  jxor g11326(.dina(n11584), .dinb(a8 ), .dout(n11585));
  jxor g11327(.dina(n11585), .dinb(n11577), .dout(n11586));
  jxor g11328(.dina(n11586), .dinb(n11311), .dout(n11587));
  jor  g11329(.dina(n10634), .dinb(n402), .dout(n11588));
  jor  g11330(.dina(n371), .dinb(n9725), .dout(n11589));
  jor  g11331(.dina(n405), .dinb(n10314), .dout(n11590));
  jor  g11332(.dina(n332), .dinb(n10637), .dout(n11591));
  jand g11333(.dina(n11591), .dinb(n11590), .dout(n11592));
  jand g11334(.dina(n11592), .dinb(n11589), .dout(n11593));
  jand g11335(.dina(n11593), .dinb(n11588), .dout(n11594));
  jxor g11336(.dina(n11594), .dinb(a5 ), .dout(n11595));
  jxor g11337(.dina(n11595), .dinb(n11587), .dout(n11596));
  jxor g11338(.dina(n11596), .dinb(n11306), .dout(n11597));
  jxor g11339(.dina(n11597), .dinb(n11290), .dout(n11598));
  jand g11340(.dina(n11285), .dinb(n11281), .dout(n11599));
  jand g11341(.dina(n11286), .dinb(n10976), .dout(n11600));
  jor  g11342(.dina(n11600), .dinb(n11599), .dout(n11601));
  jxor g11343(.dina(n11601), .dinb(n11598), .dout(f65 ));
  jor  g11344(.dina(n8806), .dinb(n706), .dout(n11603));
  jor  g11345(.dina(n683), .dinb(n8231), .dout(n11604));
  jor  g11346(.dina(n709), .dinb(n8789), .dout(n11605));
  jor  g11347(.dina(n711), .dinb(n8809), .dout(n11606));
  jand g11348(.dina(n11606), .dinb(n11605), .dout(n11607));
  jand g11349(.dina(n11607), .dinb(n11604), .dout(n11608));
  jand g11350(.dina(n11608), .dinb(n11603), .dout(n11609));
  jxor g11351(.dina(n11609), .dinb(a11 ), .dout(n11610));
  jor  g11352(.dina(n11566), .dinb(n11558), .dout(n11611));
  jand g11353(.dina(n11567), .dinb(n11314), .dout(n11612));
  jnot g11354(.din(n11612), .dout(n11613));
  jand g11355(.dina(n11613), .dinb(n11611), .dout(n11614));
  jxor g11356(.dina(n11614), .dinb(n11610), .dout(n11615));
  jor  g11357(.dina(n7146), .dinb(n1245), .dout(n11616));
  jor  g11358(.dina(n1165), .dinb(n6867), .dout(n11617));
  jor  g11359(.dina(n1248), .dinb(n7129), .dout(n11618));
  jor  g11360(.dina(n1250), .dinb(n7149), .dout(n11619));
  jand g11361(.dina(n11619), .dinb(n11618), .dout(n11620));
  jand g11362(.dina(n11620), .dinb(n11617), .dout(n11621));
  jand g11363(.dina(n11621), .dinb(n11616), .dout(n11622));
  jxor g11364(.dina(n11622), .dinb(a17 ), .dout(n11623));
  jnot g11365(.din(n11623), .dout(n11624));
  jand g11366(.dina(n11554), .dinb(n11339), .dout(n11625));
  jand g11367(.dina(n11555), .dinb(n11330), .dout(n11626));
  jor  g11368(.dina(n11626), .dinb(n11625), .dout(n11627));
  jxor g11369(.dina(n11627), .dinb(n11624), .dout(n11628));
  jor  g11370(.dina(n6369), .dinb(n1566), .dout(n11629));
  jor  g11371(.dina(n1489), .dinb(n6106), .dout(n11630));
  jor  g11372(.dina(n1569), .dinb(n6352), .dout(n11631));
  jor  g11373(.dina(n1571), .dinb(n6372), .dout(n11632));
  jand g11374(.dina(n11632), .dinb(n11631), .dout(n11633));
  jand g11375(.dina(n11633), .dinb(n11630), .dout(n11634));
  jand g11376(.dina(n11634), .dinb(n11629), .dout(n11635));
  jxor g11377(.dina(n11635), .dinb(a20 ), .dout(n11636));
  jor  g11378(.dina(n11552), .dinb(n11544), .dout(n11637));
  jand g11379(.dina(n11553), .dinb(n11342), .dout(n11638));
  jnot g11380(.din(n11638), .dout(n11639));
  jand g11381(.dina(n11639), .dinb(n11637), .dout(n11640));
  jxor g11382(.dina(n11640), .dinb(n11636), .dout(n11641));
  jor  g11383(.dina(n4991), .dinb(n2319), .dout(n11642));
  jor  g11384(.dina(n2224), .dinb(n4557), .dout(n11643));
  jor  g11385(.dina(n2322), .dinb(n4974), .dout(n11644));
  jor  g11386(.dina(n2324), .dinb(n4994), .dout(n11645));
  jand g11387(.dina(n11645), .dinb(n11644), .dout(n11646));
  jand g11388(.dina(n11646), .dinb(n11643), .dout(n11647));
  jand g11389(.dina(n11647), .dinb(n11642), .dout(n11648));
  jxor g11390(.dina(n11648), .dinb(a26 ), .dout(n11649));
  jor  g11391(.dina(n11532), .dinb(n11524), .dout(n11650));
  jnot g11392(.din(n11350), .dout(n11651));
  jand g11393(.dina(n11533), .dinb(n11651), .dout(n11652));
  jnot g11394(.din(n11652), .dout(n11653));
  jand g11395(.dina(n11653), .dinb(n11650), .dout(n11654));
  jxor g11396(.dina(n11654), .dinb(n11649), .dout(n11655));
  jor  g11397(.dina(n11522), .dinb(n11514), .dout(n11656));
  jnot g11398(.din(n11354), .dout(n11657));
  jand g11399(.dina(n11523), .dinb(n11657), .dout(n11658));
  jnot g11400(.din(n11658), .dout(n11659));
  jand g11401(.dina(n11659), .dinb(n11656), .dout(n11660));
  jor  g11402(.dina(n4534), .dinb(n2784), .dout(n11661));
  jor  g11403(.dina(n2661), .dinb(n4140), .dout(n11662));
  jor  g11404(.dina(n2787), .dinb(n4340), .dout(n11663));
  jor  g11405(.dina(n2789), .dinb(n4537), .dout(n11664));
  jand g11406(.dina(n11664), .dinb(n11663), .dout(n11665));
  jand g11407(.dina(n11665), .dinb(n11662), .dout(n11666));
  jand g11408(.dina(n11666), .dinb(n11661), .dout(n11667));
  jxor g11409(.dina(n11667), .dinb(a29 ), .dout(n11668));
  jxor g11410(.dina(n11668), .dinb(n11660), .dout(n11669));
  jor  g11411(.dina(n11511), .dinb(n11503), .dout(n11670));
  jand g11412(.dina(n11512), .dinb(n11358), .dout(n11671));
  jnot g11413(.din(n11671), .dout(n11672));
  jand g11414(.dina(n11672), .dinb(n11670), .dout(n11673));
  jor  g11415(.dina(n3939), .dinb(n3301), .dout(n11674));
  jor  g11416(.dina(n3136), .dinb(n3403), .dout(n11675));
  jor  g11417(.dina(n3304), .dinb(n3588), .dout(n11676));
  jor  g11418(.dina(n3306), .dinb(n3942), .dout(n11677));
  jand g11419(.dina(n11677), .dinb(n11676), .dout(n11678));
  jand g11420(.dina(n11678), .dinb(n11675), .dout(n11679));
  jand g11421(.dina(n11679), .dinb(n11674), .dout(n11680));
  jxor g11422(.dina(n11680), .dinb(a32 ), .dout(n11681));
  jxor g11423(.dina(n11681), .dinb(n11673), .dout(n11682));
  jor  g11424(.dina(n11489), .dinb(n11481), .dout(n11683));
  jand g11425(.dina(n11490), .dinb(n11368), .dout(n11684));
  jnot g11426(.din(n11684), .dout(n11685));
  jand g11427(.dina(n11685), .dinb(n11683), .dout(n11686));
  jnot g11428(.din(n11686), .dout(n11687));
  jand g11429(.dina(n11478), .dinb(n11382), .dout(n11688));
  jand g11430(.dina(n11479), .dinb(n11373), .dout(n11689));
  jor  g11431(.dina(n11689), .dinb(n11688), .dout(n11690));
  jand g11432(.dina(n11465), .dinb(n11400), .dout(n11691));
  jand g11433(.dina(n11466), .dinb(n11391), .dout(n11692));
  jor  g11434(.dina(n11692), .dinb(n11691), .dout(n11693));
  jor  g11435(.dina(n11463), .dinb(n11455), .dout(n11694));
  jand g11436(.dina(n11464), .dinb(n11405), .dout(n11695));
  jnot g11437(.din(n11695), .dout(n11696));
  jand g11438(.dina(n11696), .dinb(n11694), .dout(n11697));
  jand g11439(.dina(n11452), .dinb(n11419), .dout(n11698));
  jand g11440(.dina(n11453), .dinb(n11410), .dout(n11699));
  jor  g11441(.dina(n11699), .dinb(n11698), .dout(n11700));
  jor  g11442(.dina(n8978), .dinb(n755), .dout(n11701));
  jor  g11443(.dina(n8677), .dinb(n627), .dout(n11702));
  jor  g11444(.dina(n8981), .dinb(n647), .dout(n11703));
  jor  g11445(.dina(n8983), .dinb(n758), .dout(n11704));
  jand g11446(.dina(n11704), .dinb(n11703), .dout(n11705));
  jand g11447(.dina(n11705), .dinb(n11702), .dout(n11706));
  jand g11448(.dina(n11706), .dinb(n11701), .dout(n11707));
  jxor g11449(.dina(n11707), .dinb(a56 ), .dout(n11708));
  jnot g11450(.din(n11708), .dout(n11709));
  jor  g11451(.dina(n11450), .dinb(n11442), .dout(n11710));
  jand g11452(.dina(n11451), .dinb(n11424), .dout(n11711));
  jnot g11453(.din(n11711), .dout(n11712));
  jand g11454(.dina(n11712), .dinb(n11710), .dout(n11713));
  jnot g11455(.din(n11713), .dout(n11714));
  jand g11456(.dina(n11439), .dinb(n11436), .dout(n11715));
  jand g11457(.dina(n11440), .dinb(n11427), .dout(n11716));
  jor  g11458(.dina(n11716), .dinb(n11715), .dout(n11717));
  jand g11459(.dina(n10801), .dinb(b3 ), .dout(n11718));
  jand g11460(.dina(n11107), .dinb(b2 ), .dout(n11719));
  jor  g11461(.dina(n11719), .dinb(n11718), .dout(n11720));
  jxor g11462(.dina(n11720), .dinb(a2 ), .dout(n11721));
  jnot g11463(.din(n11721), .dout(n11722));
  jor  g11464(.dina(n10806), .dinb(n392), .dout(n11723));
  jor  g11465(.dina(n10485), .dinb(n322), .dout(n11724));
  jor  g11466(.dina(n10809), .dinb(n357), .dout(n11725));
  jor  g11467(.dina(n10811), .dinb(n395), .dout(n11726));
  jand g11468(.dina(n11726), .dinb(n11725), .dout(n11727));
  jand g11469(.dina(n11727), .dinb(n11724), .dout(n11728));
  jand g11470(.dina(n11728), .dinb(n11723), .dout(n11729));
  jxor g11471(.dina(n11729), .dinb(a62 ), .dout(n11730));
  jxor g11472(.dina(n11730), .dinb(n11722), .dout(n11731));
  jxor g11473(.dina(n11731), .dinb(n11717), .dout(n11732));
  jor  g11474(.dina(n9891), .dinb(n561), .dout(n11733));
  jor  g11475(.dina(n9593), .dinb(n431), .dout(n11734));
  jor  g11476(.dina(n9894), .dinb(n512), .dout(n11735));
  jor  g11477(.dina(n9896), .dinb(n564), .dout(n11736));
  jand g11478(.dina(n11736), .dinb(n11735), .dout(n11737));
  jand g11479(.dina(n11737), .dinb(n11734), .dout(n11738));
  jand g11480(.dina(n11738), .dinb(n11733), .dout(n11739));
  jxor g11481(.dina(n11739), .dinb(a59 ), .dout(n11740));
  jnot g11482(.din(n11740), .dout(n11741));
  jxor g11483(.dina(n11741), .dinb(n11732), .dout(n11742));
  jxor g11484(.dina(n11742), .dinb(n11714), .dout(n11743));
  jxor g11485(.dina(n11743), .dinb(n11709), .dout(n11744));
  jxor g11486(.dina(n11744), .dinb(n11700), .dout(n11745));
  jor  g11487(.dina(n8125), .dinb(n936), .dout(n11746));
  jor  g11488(.dina(n7846), .dinb(n778), .dout(n11747));
  jor  g11489(.dina(n8128), .dinb(n858), .dout(n11748));
  jor  g11490(.dina(n8130), .dinb(n939), .dout(n11749));
  jand g11491(.dina(n11749), .dinb(n11748), .dout(n11750));
  jand g11492(.dina(n11750), .dinb(n11747), .dout(n11751));
  jand g11493(.dina(n11751), .dinb(n11746), .dout(n11752));
  jxor g11494(.dina(n11752), .dinb(a53 ), .dout(n11753));
  jnot g11495(.din(n11753), .dout(n11754));
  jxor g11496(.dina(n11754), .dinb(n11745), .dout(n11755));
  jnot g11497(.din(n11755), .dout(n11756));
  jxor g11498(.dina(n11756), .dinb(n11697), .dout(n11757));
  jor  g11499(.dina(n7266), .dinb(n1287), .dout(n11758));
  jor  g11500(.dina(n7021), .dinb(n1022), .dout(n11759));
  jor  g11501(.dina(n7269), .dinb(n1193), .dout(n11760));
  jor  g11502(.dina(n7271), .dinb(n1290), .dout(n11761));
  jand g11503(.dina(n11761), .dinb(n11760), .dout(n11762));
  jand g11504(.dina(n11762), .dinb(n11759), .dout(n11763));
  jand g11505(.dina(n11763), .dinb(n11758), .dout(n11764));
  jxor g11506(.dina(n11764), .dinb(a50 ), .dout(n11765));
  jnot g11507(.din(n11765), .dout(n11766));
  jxor g11508(.dina(n11766), .dinb(n11757), .dout(n11767));
  jxor g11509(.dina(n11767), .dinb(n11693), .dout(n11768));
  jnot g11510(.din(n11768), .dout(n11769));
  jor  g11511(.dina(n6490), .dinb(n1617), .dout(n11770));
  jor  g11512(.dina(n6262), .dinb(n1400), .dout(n11771));
  jor  g11513(.dina(n6493), .dinb(n1420), .dout(n11772));
  jor  g11514(.dina(n6495), .dinb(n1620), .dout(n11773));
  jand g11515(.dina(n11773), .dinb(n11772), .dout(n11774));
  jand g11516(.dina(n11774), .dinb(n11771), .dout(n11775));
  jand g11517(.dina(n11775), .dinb(n11770), .dout(n11776));
  jxor g11518(.dina(n11776), .dinb(a47 ), .dout(n11777));
  jxor g11519(.dina(n11777), .dinb(n11769), .dout(n11778));
  jnot g11520(.din(n11778), .dout(n11779));
  jor  g11521(.dina(n11476), .dinb(n11468), .dout(n11780));
  jand g11522(.dina(n11477), .dinb(n11386), .dout(n11781));
  jnot g11523(.din(n11781), .dout(n11782));
  jand g11524(.dina(n11782), .dinb(n11780), .dout(n11783));
  jxor g11525(.dina(n11783), .dinb(n11779), .dout(n11784));
  jor  g11526(.dina(n5739), .dinb(n1884), .dout(n11785));
  jor  g11527(.dina(n5574), .dinb(n1742), .dout(n11786));
  jor  g11528(.dina(n5742), .dinb(n1867), .dout(n11787));
  jor  g11529(.dina(n5744), .dinb(n1887), .dout(n11788));
  jand g11530(.dina(n11788), .dinb(n11787), .dout(n11789));
  jand g11531(.dina(n11789), .dinb(n11786), .dout(n11790));
  jand g11532(.dina(n11790), .dinb(n11785), .dout(n11791));
  jxor g11533(.dina(n11791), .dinb(a44 ), .dout(n11792));
  jnot g11534(.din(n11792), .dout(n11793));
  jxor g11535(.dina(n11793), .dinb(n11784), .dout(n11794));
  jxor g11536(.dina(n11794), .dinb(n11690), .dout(n11795));
  jor  g11537(.dina(n5096), .dinb(n2404), .dout(n11796));
  jor  g11538(.dina(n4904), .dinb(n2010), .dout(n11797));
  jor  g11539(.dina(n5099), .dinb(n2148), .dout(n11798));
  jor  g11540(.dina(n5101), .dinb(n2407), .dout(n11799));
  jand g11541(.dina(n11799), .dinb(n11798), .dout(n11800));
  jand g11542(.dina(n11800), .dinb(n11797), .dout(n11801));
  jand g11543(.dina(n11801), .dinb(n11796), .dout(n11802));
  jxor g11544(.dina(n11802), .dinb(a41 ), .dout(n11803));
  jnot g11545(.din(n11803), .dout(n11804));
  jxor g11546(.dina(n11804), .dinb(n11795), .dout(n11805));
  jxor g11547(.dina(n11805), .dinb(n11687), .dout(n11806));
  jnot g11548(.din(n11806), .dout(n11807));
  jor  g11549(.dina(n4415), .dinb(n2867), .dout(n11808));
  jor  g11550(.dina(n4272), .dinb(n2559), .dout(n11809));
  jor  g11551(.dina(n4418), .dinb(n2579), .dout(n11810));
  jor  g11552(.dina(n4420), .dinb(n2870), .dout(n11811));
  jand g11553(.dina(n11811), .dinb(n11810), .dout(n11812));
  jand g11554(.dina(n11812), .dinb(n11809), .dout(n11813));
  jand g11555(.dina(n11813), .dinb(n11808), .dout(n11814));
  jxor g11556(.dina(n11814), .dinb(a38 ), .dout(n11815));
  jxor g11557(.dina(n11815), .dinb(n11807), .dout(n11816));
  jnot g11558(.din(n11816), .dout(n11817));
  jor  g11559(.dina(n11500), .dinb(n11492), .dout(n11818));
  jand g11560(.dina(n11501), .dinb(n11363), .dout(n11819));
  jnot g11561(.din(n11819), .dout(n11820));
  jand g11562(.dina(n11820), .dinb(n11818), .dout(n11821));
  jxor g11563(.dina(n11821), .dinb(n11817), .dout(n11822));
  jor  g11564(.dina(n3849), .dinb(n3227), .dout(n11823));
  jor  g11565(.dina(n3689), .dinb(n3035), .dout(n11824));
  jor  g11566(.dina(n3852), .dinb(n3055), .dout(n11825));
  jor  g11567(.dina(n3854), .dinb(n3230), .dout(n11826));
  jand g11568(.dina(n11826), .dinb(n11825), .dout(n11827));
  jand g11569(.dina(n11827), .dinb(n11824), .dout(n11828));
  jand g11570(.dina(n11828), .dinb(n11823), .dout(n11829));
  jxor g11571(.dina(n11829), .dinb(a35 ), .dout(n11830));
  jnot g11572(.din(n11830), .dout(n11831));
  jxor g11573(.dina(n11831), .dinb(n11822), .dout(n11832));
  jxor g11574(.dina(n11832), .dinb(n11682), .dout(n11833));
  jxor g11575(.dina(n11833), .dinb(n11669), .dout(n11834));
  jxor g11576(.dina(n11834), .dinb(n11655), .dout(n11835));
  jor  g11577(.dina(n11542), .dinb(n11534), .dout(n11836));
  jnot g11578(.din(n11346), .dout(n11837));
  jand g11579(.dina(n11543), .dinb(n11837), .dout(n11838));
  jnot g11580(.din(n11838), .dout(n11839));
  jand g11581(.dina(n11839), .dinb(n11836), .dout(n11840));
  jor  g11582(.dina(n5859), .dinb(n1939), .dout(n11841));
  jor  g11583(.dina(n1827), .dinb(n5408), .dout(n11842));
  jor  g11584(.dina(n1942), .dinb(n5428), .dout(n11843));
  jor  g11585(.dina(n1944), .dinb(n5862), .dout(n11844));
  jand g11586(.dina(n11844), .dinb(n11843), .dout(n11845));
  jand g11587(.dina(n11845), .dinb(n11842), .dout(n11846));
  jand g11588(.dina(n11846), .dinb(n11841), .dout(n11847));
  jxor g11589(.dina(n11847), .dinb(a23 ), .dout(n11848));
  jxor g11590(.dina(n11848), .dinb(n11840), .dout(n11849));
  jxor g11591(.dina(n11849), .dinb(n11835), .dout(n11850));
  jxor g11592(.dina(n11850), .dinb(n11641), .dout(n11851));
  jxor g11593(.dina(n11851), .dinb(n11628), .dout(n11852));
  jand g11594(.dina(n11556), .dinb(n11327), .dout(n11853));
  jand g11595(.dina(n11557), .dinb(n11317), .dout(n11854));
  jor  g11596(.dina(n11854), .dinb(n11853), .dout(n11855));
  jnot g11597(.din(n11855), .dout(n11856));
  jor  g11598(.dina(n7957), .dinb(n974), .dout(n11857));
  jor  g11599(.dina(n908), .dinb(n7411), .dout(n11858));
  jor  g11600(.dina(n977), .dinb(n7683), .dout(n11859));
  jor  g11601(.dina(n979), .dinb(n7960), .dout(n11860));
  jand g11602(.dina(n11860), .dinb(n11859), .dout(n11861));
  jand g11603(.dina(n11861), .dinb(n11858), .dout(n11862));
  jand g11604(.dina(n11862), .dinb(n11857), .dout(n11863));
  jxor g11605(.dina(n11863), .dinb(a14 ), .dout(n11864));
  jxor g11606(.dina(n11864), .dinb(n11856), .dout(n11865));
  jxor g11607(.dina(n11865), .dinb(n11852), .dout(n11866));
  jnot g11608(.din(n11866), .dout(n11867));
  jxor g11609(.dina(n11867), .dinb(n11615), .dout(n11868));
  jor  g11610(.dina(n9722), .dinb(n528), .dout(n11869));
  jor  g11611(.dina(n490), .dinb(n9390), .dout(n11870));
  jor  g11612(.dina(n531), .dinb(n9413), .dout(n11871));
  jor  g11613(.dina(n533), .dinb(n9725), .dout(n11872));
  jand g11614(.dina(n11872), .dinb(n11871), .dout(n11873));
  jand g11615(.dina(n11873), .dinb(n11870), .dout(n11874));
  jand g11616(.dina(n11874), .dinb(n11869), .dout(n11875));
  jxor g11617(.dina(n11875), .dinb(a8 ), .dout(n11876));
  jnot g11618(.din(n11876), .dout(n11877));
  jnot g11619(.din(n11568), .dout(n11878));
  jor  g11620(.dina(n11576), .dinb(n11878), .dout(n11879));
  jand g11621(.dina(n11576), .dinb(n11878), .dout(n11880));
  jor  g11622(.dina(n11585), .dinb(n11880), .dout(n11881));
  jand g11623(.dina(n11881), .dinb(n11879), .dout(n11882));
  jxor g11624(.dina(n11882), .dinb(n11877), .dout(n11883));
  jxor g11625(.dina(n11883), .dinb(n11868), .dout(n11884));
  jor  g11626(.dina(n10961), .dinb(n402), .dout(n11885));
  jor  g11627(.dina(n371), .dinb(n10314), .dout(n11886));
  jor  g11628(.dina(n405), .dinb(n10637), .dout(n11887));
  jor  g11629(.dina(n332), .dinb(n10964), .dout(n11888));
  jand g11630(.dina(n11888), .dinb(n11887), .dout(n11889));
  jand g11631(.dina(n11889), .dinb(n11886), .dout(n11890));
  jand g11632(.dina(n11890), .dinb(n11885), .dout(n11891));
  jxor g11633(.dina(n11891), .dinb(a5 ), .dout(n11892));
  jnot g11634(.din(n11892), .dout(n11893));
  jor  g11635(.dina(n11586), .dinb(n11310), .dout(n11894));
  jand g11636(.dina(n11586), .dinb(n11310), .dout(n11895));
  jnot g11637(.din(n11595), .dout(n11896));
  jor  g11638(.dina(n11896), .dinb(n11895), .dout(n11897));
  jand g11639(.dina(n11897), .dinb(n11894), .dout(n11898));
  jxor g11640(.dina(n11898), .dinb(n11893), .dout(n11899));
  jxor g11641(.dina(n11899), .dinb(n11884), .dout(n11900));
  jor  g11642(.dina(n11305), .dinb(n11295), .dout(n11901));
  jand g11643(.dina(n11305), .dinb(n11295), .dout(n11902));
  jor  g11644(.dina(n11596), .dinb(n11902), .dout(n11903));
  jand g11645(.dina(n11903), .dinb(n11901), .dout(n11904));
  jxor g11646(.dina(n11904), .dinb(n11900), .dout(n11905));
  jand g11647(.dina(n11597), .dinb(n11290), .dout(n11906));
  jand g11648(.dina(n11601), .dinb(n11598), .dout(n11907));
  jor  g11649(.dina(n11907), .dinb(n11906), .dout(n11908));
  jxor g11650(.dina(n11908), .dinb(n11905), .dout(f66 ));
  jand g11651(.dina(n11904), .dinb(n11900), .dout(n11910));
  jand g11652(.dina(n11908), .dinb(n11905), .dout(n11911));
  jor  g11653(.dina(n11911), .dinb(n11910), .dout(n11912));
  jand g11654(.dina(n11898), .dinb(n11893), .dout(n11913));
  jand g11655(.dina(n11899), .dinb(n11884), .dout(n11914));
  jor  g11656(.dina(n11914), .dinb(n11913), .dout(n11915));
  jor  g11657(.dina(n8228), .dinb(n974), .dout(n11916));
  jor  g11658(.dina(n908), .dinb(n7683), .dout(n11917));
  jor  g11659(.dina(n977), .dinb(n7960), .dout(n11918));
  jor  g11660(.dina(n979), .dinb(n8231), .dout(n11919));
  jand g11661(.dina(n11919), .dinb(n11918), .dout(n11920));
  jand g11662(.dina(n11920), .dinb(n11917), .dout(n11921));
  jand g11663(.dina(n11921), .dinb(n11916), .dout(n11922));
  jxor g11664(.dina(n11922), .dinb(a14 ), .dout(n11923));
  jnot g11665(.din(n11923), .dout(n11924));
  jand g11666(.dina(n11627), .dinb(n11624), .dout(n11925));
  jand g11667(.dina(n11851), .dinb(n11628), .dout(n11926));
  jor  g11668(.dina(n11926), .dinb(n11925), .dout(n11927));
  jxor g11669(.dina(n11927), .dinb(n11924), .dout(n11928));
  jor  g11670(.dina(n6864), .dinb(n1566), .dout(n11929));
  jor  g11671(.dina(n1489), .dinb(n6352), .dout(n11930));
  jor  g11672(.dina(n1569), .dinb(n6372), .dout(n11931));
  jor  g11673(.dina(n1571), .dinb(n6867), .dout(n11932));
  jand g11674(.dina(n11932), .dinb(n11931), .dout(n11933));
  jand g11675(.dina(n11933), .dinb(n11930), .dout(n11934));
  jand g11676(.dina(n11934), .dinb(n11929), .dout(n11935));
  jxor g11677(.dina(n11935), .dinb(a20 ), .dout(n11936));
  jor  g11678(.dina(n11848), .dinb(n11840), .dout(n11937));
  jand g11679(.dina(n11849), .dinb(n11835), .dout(n11938));
  jnot g11680(.din(n11938), .dout(n11939));
  jand g11681(.dina(n11939), .dinb(n11937), .dout(n11940));
  jxor g11682(.dina(n11940), .dinb(n11936), .dout(n11941));
  jor  g11683(.dina(n5405), .dinb(n2319), .dout(n11942));
  jor  g11684(.dina(n2224), .dinb(n4974), .dout(n11943));
  jor  g11685(.dina(n2322), .dinb(n4994), .dout(n11944));
  jor  g11686(.dina(n2324), .dinb(n5408), .dout(n11945));
  jand g11687(.dina(n11945), .dinb(n11944), .dout(n11946));
  jand g11688(.dina(n11946), .dinb(n11943), .dout(n11947));
  jand g11689(.dina(n11947), .dinb(n11942), .dout(n11948));
  jxor g11690(.dina(n11948), .dinb(a26 ), .dout(n11949));
  jor  g11691(.dina(n11668), .dinb(n11660), .dout(n11950));
  jand g11692(.dina(n11833), .dinb(n11669), .dout(n11951));
  jnot g11693(.din(n11951), .dout(n11952));
  jand g11694(.dina(n11952), .dinb(n11950), .dout(n11953));
  jxor g11695(.dina(n11953), .dinb(n11949), .dout(n11954));
  jor  g11696(.dina(n4137), .dinb(n3301), .dout(n11955));
  jor  g11697(.dina(n3136), .dinb(n3588), .dout(n11956));
  jor  g11698(.dina(n3304), .dinb(n3942), .dout(n11957));
  jor  g11699(.dina(n3306), .dinb(n4140), .dout(n11958));
  jand g11700(.dina(n11958), .dinb(n11957), .dout(n11959));
  jand g11701(.dina(n11959), .dinb(n11956), .dout(n11960));
  jand g11702(.dina(n11960), .dinb(n11955), .dout(n11961));
  jxor g11703(.dina(n11961), .dinb(a32 ), .dout(n11962));
  jnot g11704(.din(n11821), .dout(n11963));
  jand g11705(.dina(n11963), .dinb(n11816), .dout(n11964));
  jnot g11706(.din(n11964), .dout(n11965));
  jand g11707(.dina(n11821), .dinb(n11817), .dout(n11966));
  jor  g11708(.dina(n11830), .dinb(n11966), .dout(n11967));
  jand g11709(.dina(n11967), .dinb(n11965), .dout(n11968));
  jxor g11710(.dina(n11968), .dinb(n11962), .dout(n11969));
  jor  g11711(.dina(n3849), .dinb(n3400), .dout(n11970));
  jor  g11712(.dina(n3689), .dinb(n3055), .dout(n11971));
  jor  g11713(.dina(n3852), .dinb(n3230), .dout(n11972));
  jor  g11714(.dina(n3854), .dinb(n3403), .dout(n11973));
  jand g11715(.dina(n11973), .dinb(n11972), .dout(n11974));
  jand g11716(.dina(n11974), .dinb(n11971), .dout(n11975));
  jand g11717(.dina(n11975), .dinb(n11970), .dout(n11976));
  jxor g11718(.dina(n11976), .dinb(a35 ), .dout(n11977));
  jand g11719(.dina(n11805), .dinb(n11687), .dout(n11978));
  jnot g11720(.din(n11978), .dout(n11979));
  jor  g11721(.dina(n11815), .dinb(n11807), .dout(n11980));
  jand g11722(.dina(n11980), .dinb(n11979), .dout(n11981));
  jor  g11723(.dina(n5739), .dinb(n2007), .dout(n11982));
  jor  g11724(.dina(n5574), .dinb(n1867), .dout(n11983));
  jor  g11725(.dina(n5742), .dinb(n1887), .dout(n11984));
  jor  g11726(.dina(n5744), .dinb(n2010), .dout(n11985));
  jand g11727(.dina(n11985), .dinb(n11984), .dout(n11986));
  jand g11728(.dina(n11986), .dinb(n11983), .dout(n11987));
  jand g11729(.dina(n11987), .dinb(n11982), .dout(n11988));
  jxor g11730(.dina(n11988), .dinb(a44 ), .dout(n11989));
  jnot g11731(.din(n11989), .dout(n11990));
  jand g11732(.dina(n11767), .dinb(n11693), .dout(n11991));
  jnot g11733(.din(n11991), .dout(n11992));
  jor  g11734(.dina(n11777), .dinb(n11769), .dout(n11993));
  jand g11735(.dina(n11993), .dinb(n11992), .dout(n11994));
  jnot g11736(.din(n11994), .dout(n11995));
  jand g11737(.dina(n11720), .dinb(a2 ), .dout(n11996));
  jnot g11738(.din(n11996), .dout(n11997));
  jor  g11739(.dina(n11730), .dinb(n11722), .dout(n11998));
  jand g11740(.dina(n11998), .dinb(n11997), .dout(n11999));
  jnot g11741(.din(n11999), .dout(n12000));
  jor  g11742(.dina(n10806), .dinb(n428), .dout(n12001));
  jor  g11743(.dina(n10485), .dinb(n357), .dout(n12002));
  jor  g11744(.dina(n10809), .dinb(n395), .dout(n12003));
  jor  g11745(.dina(n10811), .dinb(n431), .dout(n12004));
  jand g11746(.dina(n12004), .dinb(n12003), .dout(n12005));
  jand g11747(.dina(n12005), .dinb(n12002), .dout(n12006));
  jand g11748(.dina(n12006), .dinb(n12001), .dout(n12007));
  jxor g11749(.dina(n12007), .dinb(a62 ), .dout(n12008));
  jnot g11750(.din(n12008), .dout(n12009));
  jand g11751(.dina(n10801), .dinb(b4 ), .dout(n12010));
  jand g11752(.dina(n11107), .dinb(b3 ), .dout(n12011));
  jor  g11753(.dina(n12011), .dinb(n12010), .dout(n12012));
  jxor g11754(.dina(n12012), .dinb(a2 ), .dout(n12013));
  jxor g11755(.dina(n12013), .dinb(n12009), .dout(n12014));
  jxor g11756(.dina(n12014), .dinb(n12000), .dout(n12015));
  jor  g11757(.dina(n9891), .dinb(n624), .dout(n12016));
  jor  g11758(.dina(n9593), .dinb(n512), .dout(n12017));
  jor  g11759(.dina(n9894), .dinb(n564), .dout(n12018));
  jor  g11760(.dina(n9896), .dinb(n627), .dout(n12019));
  jand g11761(.dina(n12019), .dinb(n12018), .dout(n12020));
  jand g11762(.dina(n12020), .dinb(n12017), .dout(n12021));
  jand g11763(.dina(n12021), .dinb(n12016), .dout(n12022));
  jxor g11764(.dina(n12022), .dinb(a59 ), .dout(n12023));
  jnot g11765(.din(n12023), .dout(n12024));
  jxor g11766(.dina(n12024), .dinb(n12015), .dout(n12025));
  jor  g11767(.dina(n11731), .dinb(n11717), .dout(n12026));
  jand g11768(.dina(n11731), .dinb(n11717), .dout(n12027));
  jor  g11769(.dina(n11741), .dinb(n12027), .dout(n12028));
  jand g11770(.dina(n12028), .dinb(n12026), .dout(n12029));
  jxor g11771(.dina(n12029), .dinb(n12025), .dout(n12030));
  jnot g11772(.din(n12030), .dout(n12031));
  jor  g11773(.dina(n8978), .dinb(n775), .dout(n12032));
  jor  g11774(.dina(n8677), .dinb(n647), .dout(n12033));
  jor  g11775(.dina(n8981), .dinb(n758), .dout(n12034));
  jor  g11776(.dina(n8983), .dinb(n778), .dout(n12035));
  jand g11777(.dina(n12035), .dinb(n12034), .dout(n12036));
  jand g11778(.dina(n12036), .dinb(n12033), .dout(n12037));
  jand g11779(.dina(n12037), .dinb(n12032), .dout(n12038));
  jxor g11780(.dina(n12038), .dinb(a56 ), .dout(n12039));
  jxor g11781(.dina(n12039), .dinb(n12031), .dout(n12040));
  jand g11782(.dina(n11742), .dinb(n11714), .dout(n12041));
  jand g11783(.dina(n11743), .dinb(n11709), .dout(n12042));
  jor  g11784(.dina(n12042), .dinb(n12041), .dout(n12043));
  jxor g11785(.dina(n12043), .dinb(n12040), .dout(n12044));
  jor  g11786(.dina(n8125), .dinb(n1019), .dout(n12045));
  jor  g11787(.dina(n7846), .dinb(n858), .dout(n12046));
  jor  g11788(.dina(n8128), .dinb(n939), .dout(n12047));
  jor  g11789(.dina(n8130), .dinb(n1022), .dout(n12048));
  jand g11790(.dina(n12048), .dinb(n12047), .dout(n12049));
  jand g11791(.dina(n12049), .dinb(n12046), .dout(n12050));
  jand g11792(.dina(n12050), .dinb(n12045), .dout(n12051));
  jxor g11793(.dina(n12051), .dinb(a53 ), .dout(n12052));
  jnot g11794(.din(n12052), .dout(n12053));
  jxor g11795(.dina(n12053), .dinb(n12044), .dout(n12054));
  jor  g11796(.dina(n11744), .dinb(n11700), .dout(n12055));
  jand g11797(.dina(n11744), .dinb(n11700), .dout(n12056));
  jor  g11798(.dina(n11754), .dinb(n12056), .dout(n12057));
  jand g11799(.dina(n12057), .dinb(n12055), .dout(n12058));
  jxor g11800(.dina(n12058), .dinb(n12054), .dout(n12059));
  jor  g11801(.dina(n7266), .dinb(n1397), .dout(n12060));
  jor  g11802(.dina(n7021), .dinb(n1193), .dout(n12061));
  jor  g11803(.dina(n7269), .dinb(n1290), .dout(n12062));
  jor  g11804(.dina(n7271), .dinb(n1400), .dout(n12063));
  jand g11805(.dina(n12063), .dinb(n12062), .dout(n12064));
  jand g11806(.dina(n12064), .dinb(n12061), .dout(n12065));
  jand g11807(.dina(n12065), .dinb(n12060), .dout(n12066));
  jxor g11808(.dina(n12066), .dinb(a50 ), .dout(n12067));
  jnot g11809(.din(n12067), .dout(n12068));
  jxor g11810(.dina(n12068), .dinb(n12059), .dout(n12069));
  jand g11811(.dina(n11756), .dinb(n11697), .dout(n12070));
  jnot g11812(.din(n12070), .dout(n12071));
  jnot g11813(.din(n11697), .dout(n12072));
  jand g11814(.dina(n11755), .dinb(n12072), .dout(n12073));
  jor  g11815(.dina(n11766), .dinb(n12073), .dout(n12074));
  jand g11816(.dina(n12074), .dinb(n12071), .dout(n12075));
  jxor g11817(.dina(n12075), .dinb(n12069), .dout(n12076));
  jor  g11818(.dina(n6490), .dinb(n1739), .dout(n12077));
  jor  g11819(.dina(n6262), .dinb(n1420), .dout(n12078));
  jor  g11820(.dina(n6493), .dinb(n1620), .dout(n12079));
  jor  g11821(.dina(n6495), .dinb(n1742), .dout(n12080));
  jand g11822(.dina(n12080), .dinb(n12079), .dout(n12081));
  jand g11823(.dina(n12081), .dinb(n12078), .dout(n12082));
  jand g11824(.dina(n12082), .dinb(n12077), .dout(n12083));
  jxor g11825(.dina(n12083), .dinb(a47 ), .dout(n12084));
  jnot g11826(.din(n12084), .dout(n12085));
  jxor g11827(.dina(n12085), .dinb(n12076), .dout(n12086));
  jxor g11828(.dina(n12086), .dinb(n11995), .dout(n12087));
  jxor g11829(.dina(n12087), .dinb(n11990), .dout(n12088));
  jnot g11830(.din(n12088), .dout(n12089));
  jnot g11831(.din(n11783), .dout(n12090));
  jand g11832(.dina(n12090), .dinb(n11778), .dout(n12091));
  jnot g11833(.din(n12091), .dout(n12092));
  jand g11834(.dina(n11783), .dinb(n11779), .dout(n12093));
  jor  g11835(.dina(n11792), .dinb(n12093), .dout(n12094));
  jand g11836(.dina(n12094), .dinb(n12092), .dout(n12095));
  jxor g11837(.dina(n12095), .dinb(n12089), .dout(n12096));
  jor  g11838(.dina(n5096), .dinb(n2556), .dout(n12097));
  jor  g11839(.dina(n4904), .dinb(n2148), .dout(n12098));
  jor  g11840(.dina(n5099), .dinb(n2407), .dout(n12099));
  jor  g11841(.dina(n5101), .dinb(n2559), .dout(n12100));
  jand g11842(.dina(n12100), .dinb(n12099), .dout(n12101));
  jand g11843(.dina(n12101), .dinb(n12098), .dout(n12102));
  jand g11844(.dina(n12102), .dinb(n12097), .dout(n12103));
  jxor g11845(.dina(n12103), .dinb(a41 ), .dout(n12104));
  jnot g11846(.din(n12104), .dout(n12105));
  jxor g11847(.dina(n12105), .dinb(n12096), .dout(n12106));
  jnot g11848(.din(n11690), .dout(n12107));
  jnot g11849(.din(n11794), .dout(n12108));
  jand g11850(.dina(n12108), .dinb(n12107), .dout(n12109));
  jnot g11851(.din(n12109), .dout(n12110));
  jand g11852(.dina(n11794), .dinb(n11690), .dout(n12111));
  jor  g11853(.dina(n11804), .dinb(n12111), .dout(n12112));
  jand g11854(.dina(n12112), .dinb(n12110), .dout(n12113));
  jxor g11855(.dina(n12113), .dinb(n12106), .dout(n12114));
  jnot g11856(.din(n12114), .dout(n12115));
  jor  g11857(.dina(n4415), .dinb(n3032), .dout(n12116));
  jor  g11858(.dina(n4272), .dinb(n2579), .dout(n12117));
  jor  g11859(.dina(n4418), .dinb(n2870), .dout(n12118));
  jor  g11860(.dina(n4420), .dinb(n3035), .dout(n12119));
  jand g11861(.dina(n12119), .dinb(n12118), .dout(n12120));
  jand g11862(.dina(n12120), .dinb(n12117), .dout(n12121));
  jand g11863(.dina(n12121), .dinb(n12116), .dout(n12122));
  jxor g11864(.dina(n12122), .dinb(a38 ), .dout(n12123));
  jxor g11865(.dina(n12123), .dinb(n12115), .dout(n12124));
  jxor g11866(.dina(n12124), .dinb(n11981), .dout(n12125));
  jxor g11867(.dina(n12125), .dinb(n11977), .dout(n12126));
  jxor g11868(.dina(n12126), .dinb(n11969), .dout(n12127));
  jor  g11869(.dina(n11681), .dinb(n11673), .dout(n12128));
  jand g11870(.dina(n11832), .dinb(n11682), .dout(n12129));
  jnot g11871(.din(n12129), .dout(n12130));
  jand g11872(.dina(n12130), .dinb(n12128), .dout(n12131));
  jor  g11873(.dina(n4554), .dinb(n2784), .dout(n12132));
  jor  g11874(.dina(n2661), .dinb(n4340), .dout(n12133));
  jor  g11875(.dina(n2787), .dinb(n4537), .dout(n12134));
  jor  g11876(.dina(n2789), .dinb(n4557), .dout(n12135));
  jand g11877(.dina(n12135), .dinb(n12134), .dout(n12136));
  jand g11878(.dina(n12136), .dinb(n12133), .dout(n12137));
  jand g11879(.dina(n12137), .dinb(n12132), .dout(n12138));
  jxor g11880(.dina(n12138), .dinb(a29 ), .dout(n12139));
  jxor g11881(.dina(n12139), .dinb(n12131), .dout(n12140));
  jxor g11882(.dina(n12140), .dinb(n12127), .dout(n12141));
  jxor g11883(.dina(n12141), .dinb(n11954), .dout(n12142));
  jor  g11884(.dina(n6103), .dinb(n1939), .dout(n12143));
  jor  g11885(.dina(n1827), .dinb(n5428), .dout(n12144));
  jor  g11886(.dina(n1942), .dinb(n5862), .dout(n12145));
  jor  g11887(.dina(n1944), .dinb(n6106), .dout(n12146));
  jand g11888(.dina(n12146), .dinb(n12145), .dout(n12147));
  jand g11889(.dina(n12147), .dinb(n12144), .dout(n12148));
  jand g11890(.dina(n12148), .dinb(n12143), .dout(n12149));
  jxor g11891(.dina(n12149), .dinb(a23 ), .dout(n12150));
  jor  g11892(.dina(n11654), .dinb(n11649), .dout(n12151));
  jand g11893(.dina(n11834), .dinb(n11655), .dout(n12152));
  jnot g11894(.din(n12152), .dout(n12153));
  jand g11895(.dina(n12153), .dinb(n12151), .dout(n12154));
  jxor g11896(.dina(n12154), .dinb(n12150), .dout(n12155));
  jxor g11897(.dina(n12155), .dinb(n12142), .dout(n12156));
  jxor g11898(.dina(n12156), .dinb(n11941), .dout(n12157));
  jor  g11899(.dina(n7408), .dinb(n1245), .dout(n12158));
  jor  g11900(.dina(n1165), .dinb(n7129), .dout(n12159));
  jor  g11901(.dina(n1248), .dinb(n7149), .dout(n12160));
  jor  g11902(.dina(n1250), .dinb(n7411), .dout(n12161));
  jand g11903(.dina(n12161), .dinb(n12160), .dout(n12162));
  jand g11904(.dina(n12162), .dinb(n12159), .dout(n12163));
  jand g11905(.dina(n12163), .dinb(n12158), .dout(n12164));
  jxor g11906(.dina(n12164), .dinb(a17 ), .dout(n12165));
  jor  g11907(.dina(n11640), .dinb(n11636), .dout(n12166));
  jand g11908(.dina(n11850), .dinb(n11641), .dout(n12167));
  jnot g11909(.din(n12167), .dout(n12168));
  jand g11910(.dina(n12168), .dinb(n12166), .dout(n12169));
  jxor g11911(.dina(n12169), .dinb(n12165), .dout(n12170));
  jxor g11912(.dina(n12170), .dinb(n12157), .dout(n12171));
  jxor g11913(.dina(n12171), .dinb(n11928), .dout(n12172));
  jor  g11914(.dina(n11864), .dinb(n11856), .dout(n12173));
  jand g11915(.dina(n11865), .dinb(n11852), .dout(n12174));
  jnot g11916(.din(n12174), .dout(n12175));
  jand g11917(.dina(n12175), .dinb(n12173), .dout(n12176));
  jor  g11918(.dina(n9387), .dinb(n706), .dout(n12177));
  jor  g11919(.dina(n683), .dinb(n8789), .dout(n12178));
  jor  g11920(.dina(n709), .dinb(n8809), .dout(n12179));
  jor  g11921(.dina(n711), .dinb(n9390), .dout(n12180));
  jand g11922(.dina(n12180), .dinb(n12179), .dout(n12181));
  jand g11923(.dina(n12181), .dinb(n12178), .dout(n12182));
  jand g11924(.dina(n12182), .dinb(n12177), .dout(n12183));
  jxor g11925(.dina(n12183), .dinb(a11 ), .dout(n12184));
  jxor g11926(.dina(n12184), .dinb(n12176), .dout(n12185));
  jxor g11927(.dina(n12185), .dinb(n12172), .dout(n12186));
  jor  g11928(.dina(n10311), .dinb(n528), .dout(n12187));
  jor  g11929(.dina(n490), .dinb(n9413), .dout(n12188));
  jor  g11930(.dina(n531), .dinb(n9725), .dout(n12189));
  jor  g11931(.dina(n533), .dinb(n10314), .dout(n12190));
  jand g11932(.dina(n12190), .dinb(n12189), .dout(n12191));
  jand g11933(.dina(n12191), .dinb(n12188), .dout(n12192));
  jand g11934(.dina(n12192), .dinb(n12187), .dout(n12193));
  jxor g11935(.dina(n12193), .dinb(a8 ), .dout(n12194));
  jand g11936(.dina(n11614), .dinb(n11610), .dout(n12195));
  jor  g11937(.dina(n11614), .dinb(n11610), .dout(n12196));
  jand g11938(.dina(n11867), .dinb(n12196), .dout(n12197));
  jor  g11939(.dina(n12197), .dinb(n12195), .dout(n12198));
  jxor g11940(.dina(n12198), .dinb(n12194), .dout(n12199));
  jxor g11941(.dina(n12199), .dinb(n12186), .dout(n12200));
  jor  g11942(.dina(n11882), .dinb(n11876), .dout(n12201));
  jor  g11943(.dina(n11883), .dinb(n11868), .dout(n12202));
  jand g11944(.dina(n12202), .dinb(n12201), .dout(n12203));
  jor  g11945(.dina(n10978), .dinb(n402), .dout(n12204));
  jor  g11946(.dina(n371), .dinb(n10637), .dout(n12205));
  jor  g11947(.dina(n405), .dinb(n10964), .dout(n12206));
  jand g11948(.dina(n12206), .dinb(n12205), .dout(n12207));
  jand g11949(.dina(n12207), .dinb(n12204), .dout(n12208));
  jxor g11950(.dina(n12208), .dinb(a5 ), .dout(n12209));
  jxor g11951(.dina(n12209), .dinb(n12203), .dout(n12210));
  jxor g11952(.dina(n12210), .dinb(n12200), .dout(n12211));
  jxor g11953(.dina(n12211), .dinb(n11915), .dout(n12212));
  jxor g11954(.dina(n12212), .dinb(n11912), .dout(f67 ));
  jand g11955(.dina(n12211), .dinb(n11915), .dout(n12214));
  jand g11956(.dina(n12212), .dinb(n11912), .dout(n12215));
  jor  g11957(.dina(n12215), .dinb(n12214), .dout(n12216));
  jor  g11958(.dina(n12209), .dinb(n12203), .dout(n12217));
  jnot g11959(.din(n12217), .dout(n12218));
  jand g11960(.dina(n12210), .dinb(n12200), .dout(n12219));
  jor  g11961(.dina(n12219), .dinb(n12218), .dout(n12220));
  jor  g11962(.dina(n9410), .dinb(n706), .dout(n12221));
  jor  g11963(.dina(n683), .dinb(n8809), .dout(n12222));
  jor  g11964(.dina(n709), .dinb(n9390), .dout(n12223));
  jor  g11965(.dina(n711), .dinb(n9413), .dout(n12224));
  jand g11966(.dina(n12224), .dinb(n12223), .dout(n12225));
  jand g11967(.dina(n12225), .dinb(n12222), .dout(n12226));
  jand g11968(.dina(n12226), .dinb(n12221), .dout(n12227));
  jxor g11969(.dina(n12227), .dinb(a11 ), .dout(n12228));
  jnot g11970(.din(n12228), .dout(n12229));
  jand g11971(.dina(n11927), .dinb(n11924), .dout(n12230));
  jand g11972(.dina(n12171), .dinb(n11928), .dout(n12231));
  jor  g11973(.dina(n12231), .dinb(n12230), .dout(n12232));
  jxor g11974(.dina(n12232), .dinb(n12229), .dout(n12233));
  jor  g11975(.dina(n11940), .dinb(n11936), .dout(n12234));
  jand g11976(.dina(n12156), .dinb(n11941), .dout(n12235));
  jnot g11977(.din(n12235), .dout(n12236));
  jand g11978(.dina(n12236), .dinb(n12234), .dout(n12237));
  jor  g11979(.dina(n7680), .dinb(n1245), .dout(n12238));
  jor  g11980(.dina(n1165), .dinb(n7149), .dout(n12239));
  jor  g11981(.dina(n1248), .dinb(n7411), .dout(n12240));
  jor  g11982(.dina(n1250), .dinb(n7683), .dout(n12241));
  jand g11983(.dina(n12241), .dinb(n12240), .dout(n12242));
  jand g11984(.dina(n12242), .dinb(n12239), .dout(n12243));
  jand g11985(.dina(n12243), .dinb(n12238), .dout(n12244));
  jxor g11986(.dina(n12244), .dinb(a17 ), .dout(n12245));
  jxor g11987(.dina(n12245), .dinb(n12237), .dout(n12246));
  jor  g11988(.dina(n6349), .dinb(n1939), .dout(n12247));
  jor  g11989(.dina(n1827), .dinb(n5862), .dout(n12248));
  jor  g11990(.dina(n1942), .dinb(n6106), .dout(n12249));
  jor  g11991(.dina(n1944), .dinb(n6352), .dout(n12250));
  jand g11992(.dina(n12250), .dinb(n12249), .dout(n12251));
  jand g11993(.dina(n12251), .dinb(n12248), .dout(n12252));
  jand g11994(.dina(n12252), .dinb(n12247), .dout(n12253));
  jxor g11995(.dina(n12253), .dinb(a23 ), .dout(n12254));
  jor  g11996(.dina(n11953), .dinb(n11949), .dout(n12255));
  jand g11997(.dina(n12141), .dinb(n11954), .dout(n12256));
  jnot g11998(.din(n12256), .dout(n12257));
  jand g11999(.dina(n12257), .dinb(n12255), .dout(n12258));
  jxor g12000(.dina(n12258), .dinb(n12254), .dout(n12259));
  jor  g12001(.dina(n12139), .dinb(n12131), .dout(n12260));
  jand g12002(.dina(n12140), .dinb(n12127), .dout(n12261));
  jnot g12003(.din(n12261), .dout(n12262));
  jand g12004(.dina(n12262), .dinb(n12260), .dout(n12263));
  jor  g12005(.dina(n5425), .dinb(n2319), .dout(n12264));
  jor  g12006(.dina(n2224), .dinb(n4994), .dout(n12265));
  jor  g12007(.dina(n2322), .dinb(n5408), .dout(n12266));
  jor  g12008(.dina(n2324), .dinb(n5428), .dout(n12267));
  jand g12009(.dina(n12267), .dinb(n12266), .dout(n12268));
  jand g12010(.dina(n12268), .dinb(n12265), .dout(n12269));
  jand g12011(.dina(n12269), .dinb(n12264), .dout(n12270));
  jxor g12012(.dina(n12270), .dinb(a26 ), .dout(n12271));
  jxor g12013(.dina(n12271), .dinb(n12263), .dout(n12272));
  jor  g12014(.dina(n4971), .dinb(n2784), .dout(n12273));
  jor  g12015(.dina(n2661), .dinb(n4537), .dout(n12274));
  jor  g12016(.dina(n2787), .dinb(n4557), .dout(n12275));
  jor  g12017(.dina(n2789), .dinb(n4974), .dout(n12276));
  jand g12018(.dina(n12276), .dinb(n12275), .dout(n12277));
  jand g12019(.dina(n12277), .dinb(n12274), .dout(n12278));
  jand g12020(.dina(n12278), .dinb(n12273), .dout(n12279));
  jxor g12021(.dina(n12279), .dinb(a29 ), .dout(n12280));
  jor  g12022(.dina(n11968), .dinb(n11962), .dout(n12281));
  jand g12023(.dina(n12126), .dinb(n11969), .dout(n12282));
  jnot g12024(.din(n12282), .dout(n12283));
  jand g12025(.dina(n12283), .dinb(n12281), .dout(n12284));
  jxor g12026(.dina(n12284), .dinb(n12280), .dout(n12285));
  jor  g12027(.dina(n4337), .dinb(n3301), .dout(n12286));
  jor  g12028(.dina(n3136), .dinb(n3942), .dout(n12287));
  jor  g12029(.dina(n3304), .dinb(n4140), .dout(n12288));
  jor  g12030(.dina(n3306), .dinb(n4340), .dout(n12289));
  jand g12031(.dina(n12289), .dinb(n12288), .dout(n12290));
  jand g12032(.dina(n12290), .dinb(n12287), .dout(n12291));
  jand g12033(.dina(n12291), .dinb(n12286), .dout(n12292));
  jxor g12034(.dina(n12292), .dinb(a32 ), .dout(n12293));
  jnot g12035(.din(n12293), .dout(n12294));
  jnot g12036(.din(n11981), .dout(n12295));
  jor  g12037(.dina(n12124), .dinb(n12295), .dout(n12296));
  jnot g12038(.din(n11977), .dout(n12297));
  jand g12039(.dina(n12124), .dinb(n12295), .dout(n12298));
  jor  g12040(.dina(n12298), .dinb(n12297), .dout(n12299));
  jand g12041(.dina(n12299), .dinb(n12296), .dout(n12300));
  jxor g12042(.dina(n12300), .dinb(n12294), .dout(n12301));
  jor  g12043(.dina(n12095), .dinb(n12089), .dout(n12302));
  jand g12044(.dina(n12095), .dinb(n12089), .dout(n12303));
  jor  g12045(.dina(n12104), .dinb(n12303), .dout(n12304));
  jand g12046(.dina(n12304), .dinb(n12302), .dout(n12305));
  jnot g12047(.din(n12305), .dout(n12306));
  jand g12048(.dina(n12086), .dinb(n11995), .dout(n12307));
  jand g12049(.dina(n12087), .dinb(n11990), .dout(n12308));
  jor  g12050(.dina(n12308), .dinb(n12307), .dout(n12309));
  jand g12051(.dina(n12043), .dinb(n12040), .dout(n12310));
  jnot g12052(.din(n12310), .dout(n12311));
  jnot g12053(.din(n12040), .dout(n12312));
  jnot g12054(.din(n12043), .dout(n12313));
  jand g12055(.dina(n12313), .dinb(n12312), .dout(n12314));
  jor  g12056(.dina(n12052), .dinb(n12314), .dout(n12315));
  jand g12057(.dina(n12315), .dinb(n12311), .dout(n12316));
  jnot g12058(.din(n12316), .dout(n12317));
  jor  g12059(.dina(n8125), .dinb(n1190), .dout(n12318));
  jor  g12060(.dina(n7846), .dinb(n939), .dout(n12319));
  jor  g12061(.dina(n8128), .dinb(n1022), .dout(n12320));
  jor  g12062(.dina(n8130), .dinb(n1193), .dout(n12321));
  jand g12063(.dina(n12321), .dinb(n12320), .dout(n12322));
  jand g12064(.dina(n12322), .dinb(n12319), .dout(n12323));
  jand g12065(.dina(n12323), .dinb(n12318), .dout(n12324));
  jxor g12066(.dina(n12324), .dinb(a53 ), .dout(n12325));
  jand g12067(.dina(n12029), .dinb(n12025), .dout(n12326));
  jnot g12068(.din(n12326), .dout(n12327));
  jor  g12069(.dina(n12039), .dinb(n12031), .dout(n12328));
  jand g12070(.dina(n12328), .dinb(n12327), .dout(n12329));
  jand g12071(.dina(n12012), .dinb(a2 ), .dout(n12330));
  jand g12072(.dina(n12013), .dinb(n12009), .dout(n12331));
  jor  g12073(.dina(n12331), .dinb(n12330), .dout(n12332));
  jor  g12074(.dina(n10806), .dinb(n509), .dout(n12333));
  jor  g12075(.dina(n10485), .dinb(n395), .dout(n12334));
  jor  g12076(.dina(n10809), .dinb(n431), .dout(n12335));
  jor  g12077(.dina(n10811), .dinb(n512), .dout(n12336));
  jand g12078(.dina(n12336), .dinb(n12335), .dout(n12337));
  jand g12079(.dina(n12337), .dinb(n12334), .dout(n12338));
  jand g12080(.dina(n12338), .dinb(n12333), .dout(n12339));
  jxor g12081(.dina(n12339), .dinb(a62 ), .dout(n12340));
  jnot g12082(.din(n12340), .dout(n12341));
  jand g12083(.dina(n10801), .dinb(b5 ), .dout(n12342));
  jand g12084(.dina(n11107), .dinb(b4 ), .dout(n12343));
  jor  g12085(.dina(n12343), .dinb(n12342), .dout(n12344));
  jxor g12086(.dina(n12344), .dinb(a2 ), .dout(n12345));
  jxor g12087(.dina(n12345), .dinb(n12341), .dout(n12346));
  jxor g12088(.dina(n12346), .dinb(n12332), .dout(n12347));
  jnot g12089(.din(n12347), .dout(n12348));
  jor  g12090(.dina(n9891), .dinb(n644), .dout(n12349));
  jor  g12091(.dina(n9593), .dinb(n564), .dout(n12350));
  jor  g12092(.dina(n9894), .dinb(n627), .dout(n12351));
  jor  g12093(.dina(n9896), .dinb(n647), .dout(n12352));
  jand g12094(.dina(n12352), .dinb(n12351), .dout(n12353));
  jand g12095(.dina(n12353), .dinb(n12350), .dout(n12354));
  jand g12096(.dina(n12354), .dinb(n12349), .dout(n12355));
  jxor g12097(.dina(n12355), .dinb(a59 ), .dout(n12356));
  jxor g12098(.dina(n12356), .dinb(n12348), .dout(n12357));
  jnot g12099(.din(n12014), .dout(n12358));
  jand g12100(.dina(n12358), .dinb(n11999), .dout(n12359));
  jnot g12101(.din(n12359), .dout(n12360));
  jand g12102(.dina(n12014), .dinb(n12000), .dout(n12361));
  jor  g12103(.dina(n12024), .dinb(n12361), .dout(n12362));
  jand g12104(.dina(n12362), .dinb(n12360), .dout(n12363));
  jxor g12105(.dina(n12363), .dinb(n12357), .dout(n12364));
  jor  g12106(.dina(n8978), .dinb(n855), .dout(n12365));
  jor  g12107(.dina(n8677), .dinb(n758), .dout(n12366));
  jor  g12108(.dina(n8981), .dinb(n778), .dout(n12367));
  jor  g12109(.dina(n8983), .dinb(n858), .dout(n12368));
  jand g12110(.dina(n12368), .dinb(n12367), .dout(n12369));
  jand g12111(.dina(n12369), .dinb(n12366), .dout(n12370));
  jand g12112(.dina(n12370), .dinb(n12365), .dout(n12371));
  jxor g12113(.dina(n12371), .dinb(a56 ), .dout(n12372));
  jnot g12114(.din(n12372), .dout(n12373));
  jxor g12115(.dina(n12373), .dinb(n12364), .dout(n12374));
  jxor g12116(.dina(n12374), .dinb(n12329), .dout(n12375));
  jxor g12117(.dina(n12375), .dinb(n12325), .dout(n12376));
  jxor g12118(.dina(n12376), .dinb(n12317), .dout(n12377));
  jnot g12119(.din(n12377), .dout(n12378));
  jor  g12120(.dina(n7266), .dinb(n1417), .dout(n12379));
  jor  g12121(.dina(n7021), .dinb(n1290), .dout(n12380));
  jor  g12122(.dina(n7269), .dinb(n1400), .dout(n12381));
  jor  g12123(.dina(n7271), .dinb(n1420), .dout(n12382));
  jand g12124(.dina(n12382), .dinb(n12381), .dout(n12383));
  jand g12125(.dina(n12383), .dinb(n12380), .dout(n12384));
  jand g12126(.dina(n12384), .dinb(n12379), .dout(n12385));
  jxor g12127(.dina(n12385), .dinb(a50 ), .dout(n12386));
  jxor g12128(.dina(n12386), .dinb(n12378), .dout(n12387));
  jnot g12129(.din(n12054), .dout(n12388));
  jnot g12130(.din(n12058), .dout(n12389));
  jand g12131(.dina(n12389), .dinb(n12388), .dout(n12390));
  jnot g12132(.din(n12390), .dout(n12391));
  jand g12133(.dina(n12058), .dinb(n12054), .dout(n12392));
  jor  g12134(.dina(n12068), .dinb(n12392), .dout(n12393));
  jand g12135(.dina(n12393), .dinb(n12391), .dout(n12394));
  jxor g12136(.dina(n12394), .dinb(n12387), .dout(n12395));
  jor  g12137(.dina(n6490), .dinb(n1864), .dout(n12396));
  jor  g12138(.dina(n6262), .dinb(n1620), .dout(n12397));
  jor  g12139(.dina(n6493), .dinb(n1742), .dout(n12398));
  jor  g12140(.dina(n6495), .dinb(n1867), .dout(n12399));
  jand g12141(.dina(n12399), .dinb(n12398), .dout(n12400));
  jand g12142(.dina(n12400), .dinb(n12397), .dout(n12401));
  jand g12143(.dina(n12401), .dinb(n12396), .dout(n12402));
  jxor g12144(.dina(n12402), .dinb(a47 ), .dout(n12403));
  jnot g12145(.din(n12403), .dout(n12404));
  jxor g12146(.dina(n12404), .dinb(n12395), .dout(n12405));
  jnot g12147(.din(n12069), .dout(n12406));
  jnot g12148(.din(n12075), .dout(n12407));
  jand g12149(.dina(n12407), .dinb(n12406), .dout(n12408));
  jnot g12150(.din(n12408), .dout(n12409));
  jand g12151(.dina(n12075), .dinb(n12069), .dout(n12410));
  jor  g12152(.dina(n12085), .dinb(n12410), .dout(n12411));
  jand g12153(.dina(n12411), .dinb(n12409), .dout(n12412));
  jxor g12154(.dina(n12412), .dinb(n12405), .dout(n12413));
  jor  g12155(.dina(n5739), .dinb(n2145), .dout(n12414));
  jor  g12156(.dina(n5574), .dinb(n1887), .dout(n12415));
  jor  g12157(.dina(n5742), .dinb(n2010), .dout(n12416));
  jor  g12158(.dina(n5744), .dinb(n2148), .dout(n12417));
  jand g12159(.dina(n12417), .dinb(n12416), .dout(n12418));
  jand g12160(.dina(n12418), .dinb(n12415), .dout(n12419));
  jand g12161(.dina(n12419), .dinb(n12414), .dout(n12420));
  jxor g12162(.dina(n12420), .dinb(a44 ), .dout(n12421));
  jnot g12163(.din(n12421), .dout(n12422));
  jxor g12164(.dina(n12422), .dinb(n12413), .dout(n12423));
  jxor g12165(.dina(n12423), .dinb(n12309), .dout(n12424));
  jor  g12166(.dina(n5096), .dinb(n2576), .dout(n12425));
  jor  g12167(.dina(n4904), .dinb(n2407), .dout(n12426));
  jor  g12168(.dina(n5099), .dinb(n2559), .dout(n12427));
  jor  g12169(.dina(n5101), .dinb(n2579), .dout(n12428));
  jand g12170(.dina(n12428), .dinb(n12427), .dout(n12429));
  jand g12171(.dina(n12429), .dinb(n12426), .dout(n12430));
  jand g12172(.dina(n12430), .dinb(n12425), .dout(n12431));
  jxor g12173(.dina(n12431), .dinb(a41 ), .dout(n12432));
  jnot g12174(.din(n12432), .dout(n12433));
  jxor g12175(.dina(n12433), .dinb(n12424), .dout(n12434));
  jxor g12176(.dina(n12434), .dinb(n12306), .dout(n12435));
  jnot g12177(.din(n12435), .dout(n12436));
  jor  g12178(.dina(n4415), .dinb(n3052), .dout(n12437));
  jor  g12179(.dina(n4272), .dinb(n2870), .dout(n12438));
  jor  g12180(.dina(n4418), .dinb(n3035), .dout(n12439));
  jor  g12181(.dina(n4420), .dinb(n3055), .dout(n12440));
  jand g12182(.dina(n12440), .dinb(n12439), .dout(n12441));
  jand g12183(.dina(n12441), .dinb(n12438), .dout(n12442));
  jand g12184(.dina(n12442), .dinb(n12437), .dout(n12443));
  jxor g12185(.dina(n12443), .dinb(a38 ), .dout(n12444));
  jxor g12186(.dina(n12444), .dinb(n12436), .dout(n12445));
  jnot g12187(.din(n12445), .dout(n12446));
  jand g12188(.dina(n12113), .dinb(n12106), .dout(n12447));
  jnot g12189(.din(n12447), .dout(n12448));
  jor  g12190(.dina(n12123), .dinb(n12115), .dout(n12449));
  jand g12191(.dina(n12449), .dinb(n12448), .dout(n12450));
  jxor g12192(.dina(n12450), .dinb(n12446), .dout(n12451));
  jor  g12193(.dina(n3585), .dinb(n3849), .dout(n12452));
  jor  g12194(.dina(n3689), .dinb(n3230), .dout(n12453));
  jor  g12195(.dina(n3852), .dinb(n3403), .dout(n12454));
  jor  g12196(.dina(n3854), .dinb(n3588), .dout(n12455));
  jand g12197(.dina(n12455), .dinb(n12454), .dout(n12456));
  jand g12198(.dina(n12456), .dinb(n12453), .dout(n12457));
  jand g12199(.dina(n12457), .dinb(n12452), .dout(n12458));
  jxor g12200(.dina(n12458), .dinb(a35 ), .dout(n12459));
  jnot g12201(.din(n12459), .dout(n12460));
  jxor g12202(.dina(n12460), .dinb(n12451), .dout(n12461));
  jxor g12203(.dina(n12461), .dinb(n12301), .dout(n12462));
  jxor g12204(.dina(n12462), .dinb(n12285), .dout(n12463));
  jxor g12205(.dina(n12463), .dinb(n12272), .dout(n12464));
  jxor g12206(.dina(n12464), .dinb(n12259), .dout(n12465));
  jor  g12207(.dina(n7126), .dinb(n1566), .dout(n12466));
  jor  g12208(.dina(n1489), .dinb(n6372), .dout(n12467));
  jor  g12209(.dina(n1569), .dinb(n6867), .dout(n12468));
  jor  g12210(.dina(n1571), .dinb(n7129), .dout(n12469));
  jand g12211(.dina(n12469), .dinb(n12468), .dout(n12470));
  jand g12212(.dina(n12470), .dinb(n12467), .dout(n12471));
  jand g12213(.dina(n12471), .dinb(n12466), .dout(n12472));
  jxor g12214(.dina(n12472), .dinb(a20 ), .dout(n12473));
  jor  g12215(.dina(n12154), .dinb(n12150), .dout(n12474));
  jand g12216(.dina(n12155), .dinb(n12142), .dout(n12475));
  jnot g12217(.din(n12475), .dout(n12476));
  jand g12218(.dina(n12476), .dinb(n12474), .dout(n12477));
  jxor g12219(.dina(n12477), .dinb(n12473), .dout(n12478));
  jxor g12220(.dina(n12478), .dinb(n12465), .dout(n12479));
  jxor g12221(.dina(n12479), .dinb(n12246), .dout(n12480));
  jor  g12222(.dina(n8786), .dinb(n974), .dout(n12481));
  jor  g12223(.dina(n908), .dinb(n7960), .dout(n12482));
  jor  g12224(.dina(n977), .dinb(n8231), .dout(n12483));
  jor  g12225(.dina(n979), .dinb(n8789), .dout(n12484));
  jand g12226(.dina(n12484), .dinb(n12483), .dout(n12485));
  jand g12227(.dina(n12485), .dinb(n12482), .dout(n12486));
  jand g12228(.dina(n12486), .dinb(n12481), .dout(n12487));
  jxor g12229(.dina(n12487), .dinb(a14 ), .dout(n12488));
  jor  g12230(.dina(n12169), .dinb(n12165), .dout(n12489));
  jand g12231(.dina(n12170), .dinb(n12157), .dout(n12490));
  jnot g12232(.din(n12490), .dout(n12491));
  jand g12233(.dina(n12491), .dinb(n12489), .dout(n12492));
  jxor g12234(.dina(n12492), .dinb(n12488), .dout(n12493));
  jxor g12235(.dina(n12493), .dinb(n12480), .dout(n12494));
  jxor g12236(.dina(n12494), .dinb(n12233), .dout(n12495));
  jnot g12237(.din(n12495), .dout(n12496));
  jor  g12238(.dina(n12184), .dinb(n12176), .dout(n12497));
  jnot g12239(.din(n12497), .dout(n12498));
  jand g12240(.dina(n12185), .dinb(n12172), .dout(n12499));
  jor  g12241(.dina(n12499), .dinb(n12498), .dout(n12500));
  jor  g12242(.dina(n10634), .dinb(n528), .dout(n12501));
  jor  g12243(.dina(n490), .dinb(n9725), .dout(n12502));
  jor  g12244(.dina(n531), .dinb(n10314), .dout(n12503));
  jor  g12245(.dina(n533), .dinb(n10637), .dout(n12504));
  jand g12246(.dina(n12504), .dinb(n12503), .dout(n12505));
  jand g12247(.dina(n12505), .dinb(n12502), .dout(n12506));
  jand g12248(.dina(n12506), .dinb(n12501), .dout(n12507));
  jxor g12249(.dina(n12507), .dinb(a8 ), .dout(n12508));
  jxor g12250(.dina(n12508), .dinb(n12500), .dout(n12509));
  jxor g12251(.dina(n12509), .dinb(n12496), .dout(n12510));
  jnot g12252(.din(n12194), .dout(n12511));
  jnot g12253(.din(n12198), .dout(n12512));
  jand g12254(.dina(n12512), .dinb(n12511), .dout(n12513));
  jand g12255(.dina(n12199), .dinb(n12186), .dout(n12514));
  jor  g12256(.dina(n12514), .dinb(n12513), .dout(n12515));
  jnot g12257(.din(n12515), .dout(n12516));
  jnot g12258(.din(n371), .dout(n12517));
  jand g12259(.dina(n11296), .dinb(n339), .dout(n12518));
  jor  g12260(.dina(n12518), .dinb(n12517), .dout(n12519));
  jand g12261(.dina(n12519), .dinb(b63 ), .dout(n12520));
  jxor g12262(.dina(n12520), .dinb(n364), .dout(n12521));
  jxor g12263(.dina(n12521), .dinb(n12516), .dout(n12522));
  jxor g12264(.dina(n12522), .dinb(n12510), .dout(n12523));
  jxor g12265(.dina(n12523), .dinb(n12220), .dout(n12524));
  jxor g12266(.dina(n12524), .dinb(n12216), .dout(f68 ));
  jand g12267(.dina(n12523), .dinb(n12220), .dout(n12526));
  jand g12268(.dina(n12524), .dinb(n12216), .dout(n12527));
  jor  g12269(.dina(n12527), .dinb(n12526), .dout(n12528));
  jor  g12270(.dina(n12521), .dinb(n12516), .dout(n12529));
  jnot g12271(.din(n12529), .dout(n12530));
  jand g12272(.dina(n12522), .dinb(n12510), .dout(n12531));
  jor  g12273(.dina(n12531), .dinb(n12530), .dout(n12532));
  jnot g12274(.din(n12500), .dout(n12533));
  jor  g12275(.dina(n12508), .dinb(n12533), .dout(n12534));
  jor  g12276(.dina(n12509), .dinb(n12496), .dout(n12535));
  jand g12277(.dina(n12535), .dinb(n12534), .dout(n12536));
  jor  g12278(.dina(n10961), .dinb(n528), .dout(n12537));
  jor  g12279(.dina(n490), .dinb(n10314), .dout(n12538));
  jor  g12280(.dina(n531), .dinb(n10637), .dout(n12539));
  jor  g12281(.dina(n533), .dinb(n10964), .dout(n12540));
  jand g12282(.dina(n12540), .dinb(n12539), .dout(n12541));
  jand g12283(.dina(n12541), .dinb(n12538), .dout(n12542));
  jand g12284(.dina(n12542), .dinb(n12537), .dout(n12543));
  jxor g12285(.dina(n12543), .dinb(a8 ), .dout(n12544));
  jxor g12286(.dina(n12544), .dinb(n12536), .dout(n12545));
  jor  g12287(.dina(n9722), .dinb(n706), .dout(n12546));
  jor  g12288(.dina(n683), .dinb(n9390), .dout(n12547));
  jor  g12289(.dina(n709), .dinb(n9413), .dout(n12548));
  jor  g12290(.dina(n711), .dinb(n9725), .dout(n12549));
  jand g12291(.dina(n12549), .dinb(n12548), .dout(n12550));
  jand g12292(.dina(n12550), .dinb(n12547), .dout(n12551));
  jand g12293(.dina(n12551), .dinb(n12546), .dout(n12552));
  jxor g12294(.dina(n12552), .dinb(a11 ), .dout(n12553));
  jnot g12295(.din(n12553), .dout(n12554));
  jand g12296(.dina(n12232), .dinb(n12229), .dout(n12555));
  jand g12297(.dina(n12494), .dinb(n12233), .dout(n12556));
  jor  g12298(.dina(n12556), .dinb(n12555), .dout(n12557));
  jxor g12299(.dina(n12557), .dinb(n12554), .dout(n12558));
  jor  g12300(.dina(n8806), .dinb(n974), .dout(n12559));
  jor  g12301(.dina(n908), .dinb(n8231), .dout(n12560));
  jor  g12302(.dina(n977), .dinb(n8789), .dout(n12561));
  jor  g12303(.dina(n979), .dinb(n8809), .dout(n12562));
  jand g12304(.dina(n12562), .dinb(n12561), .dout(n12563));
  jand g12305(.dina(n12563), .dinb(n12560), .dout(n12564));
  jand g12306(.dina(n12564), .dinb(n12559), .dout(n12565));
  jxor g12307(.dina(n12565), .dinb(a14 ), .dout(n12566));
  jor  g12308(.dina(n12492), .dinb(n12488), .dout(n12567));
  jand g12309(.dina(n12493), .dinb(n12480), .dout(n12568));
  jnot g12310(.din(n12568), .dout(n12569));
  jand g12311(.dina(n12569), .dinb(n12567), .dout(n12570));
  jxor g12312(.dina(n12570), .dinb(n12566), .dout(n12571));
  jor  g12313(.dina(n7146), .dinb(n1566), .dout(n12572));
  jor  g12314(.dina(n1489), .dinb(n6867), .dout(n12573));
  jor  g12315(.dina(n1569), .dinb(n7129), .dout(n12574));
  jor  g12316(.dina(n1571), .dinb(n7149), .dout(n12575));
  jand g12317(.dina(n12575), .dinb(n12574), .dout(n12576));
  jand g12318(.dina(n12576), .dinb(n12573), .dout(n12577));
  jand g12319(.dina(n12577), .dinb(n12572), .dout(n12578));
  jxor g12320(.dina(n12578), .dinb(a20 ), .dout(n12579));
  jor  g12321(.dina(n12477), .dinb(n12473), .dout(n12580));
  jand g12322(.dina(n12478), .dinb(n12465), .dout(n12581));
  jnot g12323(.din(n12581), .dout(n12582));
  jand g12324(.dina(n12582), .dinb(n12580), .dout(n12583));
  jxor g12325(.dina(n12583), .dinb(n12579), .dout(n12584));
  jor  g12326(.dina(n6369), .dinb(n1939), .dout(n12585));
  jor  g12327(.dina(n1827), .dinb(n6106), .dout(n12586));
  jor  g12328(.dina(n1942), .dinb(n6352), .dout(n12587));
  jor  g12329(.dina(n1944), .dinb(n6372), .dout(n12588));
  jand g12330(.dina(n12588), .dinb(n12587), .dout(n12589));
  jand g12331(.dina(n12589), .dinb(n12586), .dout(n12590));
  jand g12332(.dina(n12590), .dinb(n12585), .dout(n12591));
  jxor g12333(.dina(n12591), .dinb(a23 ), .dout(n12592));
  jor  g12334(.dina(n12258), .dinb(n12254), .dout(n12593));
  jand g12335(.dina(n12464), .dinb(n12259), .dout(n12594));
  jnot g12336(.din(n12594), .dout(n12595));
  jand g12337(.dina(n12595), .dinb(n12593), .dout(n12596));
  jxor g12338(.dina(n12596), .dinb(n12592), .dout(n12597));
  jor  g12339(.dina(n4991), .dinb(n2784), .dout(n12598));
  jor  g12340(.dina(n2661), .dinb(n4557), .dout(n12599));
  jor  g12341(.dina(n2787), .dinb(n4974), .dout(n12600));
  jor  g12342(.dina(n2789), .dinb(n4994), .dout(n12601));
  jand g12343(.dina(n12601), .dinb(n12600), .dout(n12602));
  jand g12344(.dina(n12602), .dinb(n12599), .dout(n12603));
  jand g12345(.dina(n12603), .dinb(n12598), .dout(n12604));
  jxor g12346(.dina(n12604), .dinb(a29 ), .dout(n12605));
  jand g12347(.dina(n12284), .dinb(n12280), .dout(n12606));
  jor  g12348(.dina(n12284), .dinb(n12280), .dout(n12607));
  jnot g12349(.din(n12462), .dout(n12608));
  jand g12350(.dina(n12608), .dinb(n12607), .dout(n12609));
  jor  g12351(.dina(n12609), .dinb(n12606), .dout(n12610));
  jxor g12352(.dina(n12610), .dinb(n12605), .dout(n12611));
  jor  g12353(.dina(n3939), .dinb(n3849), .dout(n12612));
  jor  g12354(.dina(n3689), .dinb(n3403), .dout(n12613));
  jor  g12355(.dina(n3852), .dinb(n3588), .dout(n12614));
  jor  g12356(.dina(n3854), .dinb(n3942), .dout(n12615));
  jand g12357(.dina(n12615), .dinb(n12614), .dout(n12616));
  jand g12358(.dina(n12616), .dinb(n12613), .dout(n12617));
  jand g12359(.dina(n12617), .dinb(n12612), .dout(n12618));
  jxor g12360(.dina(n12618), .dinb(a35 ), .dout(n12619));
  jnot g12361(.din(n12619), .dout(n12620));
  jand g12362(.dina(n12434), .dinb(n12306), .dout(n12621));
  jnot g12363(.din(n12621), .dout(n12622));
  jor  g12364(.dina(n12444), .dinb(n12436), .dout(n12623));
  jand g12365(.dina(n12623), .dinb(n12622), .dout(n12624));
  jnot g12366(.din(n12624), .dout(n12625));
  jor  g12367(.dina(n4415), .dinb(n3227), .dout(n12626));
  jor  g12368(.dina(n4272), .dinb(n3035), .dout(n12627));
  jor  g12369(.dina(n4418), .dinb(n3055), .dout(n12628));
  jor  g12370(.dina(n4420), .dinb(n3230), .dout(n12629));
  jand g12371(.dina(n12629), .dinb(n12628), .dout(n12630));
  jand g12372(.dina(n12630), .dinb(n12627), .dout(n12631));
  jand g12373(.dina(n12631), .dinb(n12626), .dout(n12632));
  jxor g12374(.dina(n12632), .dinb(a38 ), .dout(n12633));
  jor  g12375(.dina(n6490), .dinb(n1884), .dout(n12634));
  jor  g12376(.dina(n6262), .dinb(n1742), .dout(n12635));
  jor  g12377(.dina(n6493), .dinb(n1867), .dout(n12636));
  jor  g12378(.dina(n6495), .dinb(n1887), .dout(n12637));
  jand g12379(.dina(n12637), .dinb(n12636), .dout(n12638));
  jand g12380(.dina(n12638), .dinb(n12635), .dout(n12639));
  jand g12381(.dina(n12639), .dinb(n12634), .dout(n12640));
  jxor g12382(.dina(n12640), .dinb(a47 ), .dout(n12641));
  jnot g12383(.din(n12641), .dout(n12642));
  jand g12384(.dina(n12376), .dinb(n12317), .dout(n12643));
  jnot g12385(.din(n12643), .dout(n12644));
  jor  g12386(.dina(n12386), .dinb(n12378), .dout(n12645));
  jand g12387(.dina(n12645), .dinb(n12644), .dout(n12646));
  jnot g12388(.din(n12646), .dout(n12647));
  jor  g12389(.dina(n8978), .dinb(n936), .dout(n12648));
  jor  g12390(.dina(n8677), .dinb(n778), .dout(n12649));
  jor  g12391(.dina(n8981), .dinb(n858), .dout(n12650));
  jor  g12392(.dina(n8983), .dinb(n939), .dout(n12651));
  jand g12393(.dina(n12651), .dinb(n12650), .dout(n12652));
  jand g12394(.dina(n12652), .dinb(n12649), .dout(n12653));
  jand g12395(.dina(n12653), .dinb(n12648), .dout(n12654));
  jxor g12396(.dina(n12654), .dinb(a56 ), .dout(n12655));
  jnot g12397(.din(n12655), .dout(n12656));
  jand g12398(.dina(n12346), .dinb(n12332), .dout(n12657));
  jnot g12399(.din(n12657), .dout(n12658));
  jor  g12400(.dina(n12356), .dinb(n12348), .dout(n12659));
  jand g12401(.dina(n12659), .dinb(n12658), .dout(n12660));
  jnot g12402(.din(n12660), .dout(n12661));
  jor  g12403(.dina(n9891), .dinb(n755), .dout(n12662));
  jor  g12404(.dina(n9593), .dinb(n627), .dout(n12663));
  jor  g12405(.dina(n9894), .dinb(n647), .dout(n12664));
  jor  g12406(.dina(n9896), .dinb(n758), .dout(n12665));
  jand g12407(.dina(n12665), .dinb(n12664), .dout(n12666));
  jand g12408(.dina(n12666), .dinb(n12663), .dout(n12667));
  jand g12409(.dina(n12667), .dinb(n12662), .dout(n12668));
  jxor g12410(.dina(n12668), .dinb(a59 ), .dout(n12669));
  jnot g12411(.din(n12669), .dout(n12670));
  jand g12412(.dina(n12344), .dinb(a2 ), .dout(n12671));
  jand g12413(.dina(n12345), .dinb(n12341), .dout(n12672));
  jor  g12414(.dina(n12672), .dinb(n12671), .dout(n12673));
  jxor g12415(.dina(a5 ), .dinb(a2 ), .dout(n12674));
  jand g12416(.dina(n10801), .dinb(b6 ), .dout(n12675));
  jand g12417(.dina(n11107), .dinb(b5 ), .dout(n12676));
  jor  g12418(.dina(n12676), .dinb(n12675), .dout(n12677));
  jxor g12419(.dina(n12677), .dinb(n12674), .dout(n12678));
  jxor g12420(.dina(n12678), .dinb(n12673), .dout(n12679));
  jnot g12421(.din(n12679), .dout(n12680));
  jor  g12422(.dina(n10806), .dinb(n561), .dout(n12681));
  jor  g12423(.dina(n10485), .dinb(n431), .dout(n12682));
  jor  g12424(.dina(n10809), .dinb(n512), .dout(n12683));
  jor  g12425(.dina(n10811), .dinb(n564), .dout(n12684));
  jand g12426(.dina(n12684), .dinb(n12683), .dout(n12685));
  jand g12427(.dina(n12685), .dinb(n12682), .dout(n12686));
  jand g12428(.dina(n12686), .dinb(n12681), .dout(n12687));
  jxor g12429(.dina(n12687), .dinb(a62 ), .dout(n12688));
  jxor g12430(.dina(n12688), .dinb(n12680), .dout(n12689));
  jxor g12431(.dina(n12689), .dinb(n12670), .dout(n12690));
  jxor g12432(.dina(n12690), .dinb(n12661), .dout(n12691));
  jxor g12433(.dina(n12691), .dinb(n12656), .dout(n12692));
  jor  g12434(.dina(n12363), .dinb(n12357), .dout(n12693));
  jand g12435(.dina(n12363), .dinb(n12357), .dout(n12694));
  jor  g12436(.dina(n12373), .dinb(n12694), .dout(n12695));
  jand g12437(.dina(n12695), .dinb(n12693), .dout(n12696));
  jxor g12438(.dina(n12696), .dinb(n12692), .dout(n12697));
  jnot g12439(.din(n12697), .dout(n12698));
  jor  g12440(.dina(n8125), .dinb(n1287), .dout(n12699));
  jor  g12441(.dina(n7846), .dinb(n1022), .dout(n12700));
  jor  g12442(.dina(n8128), .dinb(n1193), .dout(n12701));
  jor  g12443(.dina(n8130), .dinb(n1290), .dout(n12702));
  jand g12444(.dina(n12702), .dinb(n12701), .dout(n12703));
  jand g12445(.dina(n12703), .dinb(n12700), .dout(n12704));
  jand g12446(.dina(n12704), .dinb(n12699), .dout(n12705));
  jxor g12447(.dina(n12705), .dinb(a53 ), .dout(n12706));
  jxor g12448(.dina(n12706), .dinb(n12698), .dout(n12707));
  jnot g12449(.din(n12329), .dout(n12708));
  jor  g12450(.dina(n12374), .dinb(n12708), .dout(n12709));
  jnot g12451(.din(n12325), .dout(n12710));
  jand g12452(.dina(n12374), .dinb(n12708), .dout(n12711));
  jor  g12453(.dina(n12711), .dinb(n12710), .dout(n12712));
  jand g12454(.dina(n12712), .dinb(n12709), .dout(n12713));
  jxor g12455(.dina(n12713), .dinb(n12707), .dout(n12714));
  jnot g12456(.din(n12714), .dout(n12715));
  jor  g12457(.dina(n7266), .dinb(n1617), .dout(n12716));
  jor  g12458(.dina(n7021), .dinb(n1400), .dout(n12717));
  jor  g12459(.dina(n7269), .dinb(n1420), .dout(n12718));
  jor  g12460(.dina(n7271), .dinb(n1620), .dout(n12719));
  jand g12461(.dina(n12719), .dinb(n12718), .dout(n12720));
  jand g12462(.dina(n12720), .dinb(n12717), .dout(n12721));
  jand g12463(.dina(n12721), .dinb(n12716), .dout(n12722));
  jxor g12464(.dina(n12722), .dinb(a50 ), .dout(n12723));
  jxor g12465(.dina(n12723), .dinb(n12715), .dout(n12724));
  jxor g12466(.dina(n12724), .dinb(n12647), .dout(n12725));
  jxor g12467(.dina(n12725), .dinb(n12642), .dout(n12726));
  jor  g12468(.dina(n12394), .dinb(n12387), .dout(n12727));
  jand g12469(.dina(n12394), .dinb(n12387), .dout(n12728));
  jor  g12470(.dina(n12404), .dinb(n12728), .dout(n12729));
  jand g12471(.dina(n12729), .dinb(n12727), .dout(n12730));
  jxor g12472(.dina(n12730), .dinb(n12726), .dout(n12731));
  jnot g12473(.din(n12731), .dout(n12732));
  jor  g12474(.dina(n5739), .dinb(n2404), .dout(n12733));
  jor  g12475(.dina(n5574), .dinb(n2010), .dout(n12734));
  jor  g12476(.dina(n5742), .dinb(n2148), .dout(n12735));
  jor  g12477(.dina(n5744), .dinb(n2407), .dout(n12736));
  jand g12478(.dina(n12736), .dinb(n12735), .dout(n12737));
  jand g12479(.dina(n12737), .dinb(n12734), .dout(n12738));
  jand g12480(.dina(n12738), .dinb(n12733), .dout(n12739));
  jxor g12481(.dina(n12739), .dinb(a44 ), .dout(n12740));
  jxor g12482(.dina(n12740), .dinb(n12732), .dout(n12741));
  jnot g12483(.din(n12405), .dout(n12742));
  jnot g12484(.din(n12412), .dout(n12743));
  jand g12485(.dina(n12743), .dinb(n12742), .dout(n12744));
  jnot g12486(.din(n12744), .dout(n12745));
  jand g12487(.dina(n12412), .dinb(n12405), .dout(n12746));
  jor  g12488(.dina(n12422), .dinb(n12746), .dout(n12747));
  jand g12489(.dina(n12747), .dinb(n12745), .dout(n12748));
  jxor g12490(.dina(n12748), .dinb(n12741), .dout(n12749));
  jnot g12491(.din(n12749), .dout(n12750));
  jor  g12492(.dina(n5096), .dinb(n2867), .dout(n12751));
  jor  g12493(.dina(n4904), .dinb(n2559), .dout(n12752));
  jor  g12494(.dina(n5099), .dinb(n2579), .dout(n12753));
  jor  g12495(.dina(n5101), .dinb(n2870), .dout(n12754));
  jand g12496(.dina(n12754), .dinb(n12753), .dout(n12755));
  jand g12497(.dina(n12755), .dinb(n12752), .dout(n12756));
  jand g12498(.dina(n12756), .dinb(n12751), .dout(n12757));
  jxor g12499(.dina(n12757), .dinb(a41 ), .dout(n12758));
  jxor g12500(.dina(n12758), .dinb(n12750), .dout(n12759));
  jnot g12501(.din(n12759), .dout(n12760));
  jnot g12502(.din(n12309), .dout(n12761));
  jnot g12503(.din(n12423), .dout(n12762));
  jand g12504(.dina(n12762), .dinb(n12761), .dout(n12763));
  jnot g12505(.din(n12763), .dout(n12764));
  jand g12506(.dina(n12423), .dinb(n12309), .dout(n12765));
  jor  g12507(.dina(n12433), .dinb(n12765), .dout(n12766));
  jand g12508(.dina(n12766), .dinb(n12764), .dout(n12767));
  jxor g12509(.dina(n12767), .dinb(n12760), .dout(n12768));
  jxor g12510(.dina(n12768), .dinb(n12633), .dout(n12769));
  jxor g12511(.dina(n12769), .dinb(n12625), .dout(n12770));
  jxor g12512(.dina(n12770), .dinb(n12620), .dout(n12771));
  jnot g12513(.din(n12771), .dout(n12772));
  jnot g12514(.din(n12450), .dout(n12773));
  jand g12515(.dina(n12773), .dinb(n12445), .dout(n12774));
  jnot g12516(.din(n12774), .dout(n12775));
  jand g12517(.dina(n12450), .dinb(n12446), .dout(n12776));
  jor  g12518(.dina(n12459), .dinb(n12776), .dout(n12777));
  jand g12519(.dina(n12777), .dinb(n12775), .dout(n12778));
  jxor g12520(.dina(n12778), .dinb(n12772), .dout(n12779));
  jor  g12521(.dina(n4534), .dinb(n3301), .dout(n12780));
  jor  g12522(.dina(n3136), .dinb(n4140), .dout(n12781));
  jor  g12523(.dina(n3304), .dinb(n4340), .dout(n12782));
  jor  g12524(.dina(n3306), .dinb(n4537), .dout(n12783));
  jand g12525(.dina(n12783), .dinb(n12782), .dout(n12784));
  jand g12526(.dina(n12784), .dinb(n12781), .dout(n12785));
  jand g12527(.dina(n12785), .dinb(n12780), .dout(n12786));
  jxor g12528(.dina(n12786), .dinb(a32 ), .dout(n12787));
  jnot g12529(.din(n12787), .dout(n12788));
  jor  g12530(.dina(n12300), .dinb(n12294), .dout(n12789));
  jand g12531(.dina(n12300), .dinb(n12294), .dout(n12790));
  jor  g12532(.dina(n12461), .dinb(n12790), .dout(n12791));
  jand g12533(.dina(n12791), .dinb(n12789), .dout(n12792));
  jxor g12534(.dina(n12792), .dinb(n12788), .dout(n12793));
  jxor g12535(.dina(n12793), .dinb(n12779), .dout(n12794));
  jxor g12536(.dina(n12794), .dinb(n12611), .dout(n12795));
  jor  g12537(.dina(n12271), .dinb(n12263), .dout(n12796));
  jand g12538(.dina(n12463), .dinb(n12272), .dout(n12797));
  jnot g12539(.din(n12797), .dout(n12798));
  jand g12540(.dina(n12798), .dinb(n12796), .dout(n12799));
  jor  g12541(.dina(n5859), .dinb(n2319), .dout(n12800));
  jor  g12542(.dina(n2224), .dinb(n5408), .dout(n12801));
  jor  g12543(.dina(n2322), .dinb(n5428), .dout(n12802));
  jor  g12544(.dina(n2324), .dinb(n5862), .dout(n12803));
  jand g12545(.dina(n12803), .dinb(n12802), .dout(n12804));
  jand g12546(.dina(n12804), .dinb(n12801), .dout(n12805));
  jand g12547(.dina(n12805), .dinb(n12800), .dout(n12806));
  jxor g12548(.dina(n12806), .dinb(a26 ), .dout(n12807));
  jxor g12549(.dina(n12807), .dinb(n12799), .dout(n12808));
  jxor g12550(.dina(n12808), .dinb(n12795), .dout(n12809));
  jxor g12551(.dina(n12809), .dinb(n12597), .dout(n12810));
  jxor g12552(.dina(n12810), .dinb(n12584), .dout(n12811));
  jor  g12553(.dina(n12245), .dinb(n12237), .dout(n12812));
  jand g12554(.dina(n12479), .dinb(n12246), .dout(n12813));
  jnot g12555(.din(n12813), .dout(n12814));
  jand g12556(.dina(n12814), .dinb(n12812), .dout(n12815));
  jor  g12557(.dina(n7957), .dinb(n1245), .dout(n12816));
  jor  g12558(.dina(n1165), .dinb(n7411), .dout(n12817));
  jor  g12559(.dina(n1248), .dinb(n7683), .dout(n12818));
  jor  g12560(.dina(n1250), .dinb(n7960), .dout(n12819));
  jand g12561(.dina(n12819), .dinb(n12818), .dout(n12820));
  jand g12562(.dina(n12820), .dinb(n12817), .dout(n12821));
  jand g12563(.dina(n12821), .dinb(n12816), .dout(n12822));
  jxor g12564(.dina(n12822), .dinb(a17 ), .dout(n12823));
  jxor g12565(.dina(n12823), .dinb(n12815), .dout(n12824));
  jxor g12566(.dina(n12824), .dinb(n12811), .dout(n12825));
  jxor g12567(.dina(n12825), .dinb(n12571), .dout(n12826));
  jxor g12568(.dina(n12826), .dinb(n12558), .dout(n12827));
  jxor g12569(.dina(n12827), .dinb(n12545), .dout(n12828));
  jxor g12570(.dina(n12828), .dinb(n12532), .dout(n12829));
  jxor g12571(.dina(n12829), .dinb(n12528), .dout(f69 ));
  jand g12572(.dina(n12828), .dinb(n12532), .dout(n12831));
  jand g12573(.dina(n12829), .dinb(n12528), .dout(n12832));
  jor  g12574(.dina(n12832), .dinb(n12831), .dout(n12833));
  jor  g12575(.dina(n12544), .dinb(n12536), .dout(n12834));
  jand g12576(.dina(n12827), .dinb(n12545), .dout(n12835));
  jnot g12577(.din(n12835), .dout(n12836));
  jand g12578(.dina(n12836), .dinb(n12834), .dout(n12837));
  jnot g12579(.din(n12837), .dout(n12838));
  jor  g12580(.dina(n10978), .dinb(n528), .dout(n12839));
  jor  g12581(.dina(n490), .dinb(n10637), .dout(n12840));
  jor  g12582(.dina(n531), .dinb(n10964), .dout(n12841));
  jand g12583(.dina(n12841), .dinb(n12840), .dout(n12842));
  jand g12584(.dina(n12842), .dinb(n12839), .dout(n12843));
  jxor g12585(.dina(n12843), .dinb(a8 ), .dout(n12844));
  jnot g12586(.din(n12844), .dout(n12845));
  jnot g12587(.din(n12557), .dout(n12846));
  jand g12588(.dina(n12846), .dinb(n12553), .dout(n12847));
  jnot g12589(.din(n12847), .dout(n12848));
  jand g12590(.dina(n12557), .dinb(n12554), .dout(n12849));
  jor  g12591(.dina(n12826), .dinb(n12849), .dout(n12850));
  jand g12592(.dina(n12850), .dinb(n12848), .dout(n12851));
  jxor g12593(.dina(n12851), .dinb(n12845), .dout(n12852));
  jor  g12594(.dina(n10311), .dinb(n706), .dout(n12853));
  jor  g12595(.dina(n683), .dinb(n9413), .dout(n12854));
  jor  g12596(.dina(n709), .dinb(n9725), .dout(n12855));
  jor  g12597(.dina(n711), .dinb(n10314), .dout(n12856));
  jand g12598(.dina(n12856), .dinb(n12855), .dout(n12857));
  jand g12599(.dina(n12857), .dinb(n12854), .dout(n12858));
  jand g12600(.dina(n12858), .dinb(n12853), .dout(n12859));
  jxor g12601(.dina(n12859), .dinb(a11 ), .dout(n12860));
  jand g12602(.dina(n12570), .dinb(n12566), .dout(n12861));
  jnot g12603(.din(n12861), .dout(n12862));
  jnot g12604(.din(n12566), .dout(n12863));
  jnot g12605(.din(n12570), .dout(n12864));
  jand g12606(.dina(n12864), .dinb(n12863), .dout(n12865));
  jor  g12607(.dina(n12825), .dinb(n12865), .dout(n12866));
  jand g12608(.dina(n12866), .dinb(n12862), .dout(n12867));
  jxor g12609(.dina(n12867), .dinb(n12860), .dout(n12868));
  jor  g12610(.dina(n12823), .dinb(n12815), .dout(n12869));
  jnot g12611(.din(n12869), .dout(n12870));
  jand g12612(.dina(n12824), .dinb(n12811), .dout(n12871));
  jor  g12613(.dina(n12871), .dinb(n12870), .dout(n12872));
  jor  g12614(.dina(n9387), .dinb(n974), .dout(n12873));
  jor  g12615(.dina(n908), .dinb(n8789), .dout(n12874));
  jor  g12616(.dina(n977), .dinb(n8809), .dout(n12875));
  jor  g12617(.dina(n979), .dinb(n9390), .dout(n12876));
  jand g12618(.dina(n12876), .dinb(n12875), .dout(n12877));
  jand g12619(.dina(n12877), .dinb(n12874), .dout(n12878));
  jand g12620(.dina(n12878), .dinb(n12873), .dout(n12879));
  jxor g12621(.dina(n12879), .dinb(a14 ), .dout(n12880));
  jxor g12622(.dina(n12880), .dinb(n12872), .dout(n12881));
  jor  g12623(.dina(n8228), .dinb(n1245), .dout(n12882));
  jor  g12624(.dina(n1165), .dinb(n7683), .dout(n12883));
  jor  g12625(.dina(n1248), .dinb(n7960), .dout(n12884));
  jor  g12626(.dina(n1250), .dinb(n8231), .dout(n12885));
  jand g12627(.dina(n12885), .dinb(n12884), .dout(n12886));
  jand g12628(.dina(n12886), .dinb(n12883), .dout(n12887));
  jand g12629(.dina(n12887), .dinb(n12882), .dout(n12888));
  jxor g12630(.dina(n12888), .dinb(a17 ), .dout(n12889));
  jor  g12631(.dina(n12583), .dinb(n12579), .dout(n12890));
  jand g12632(.dina(n12810), .dinb(n12584), .dout(n12891));
  jnot g12633(.din(n12891), .dout(n12892));
  jand g12634(.dina(n12892), .dinb(n12890), .dout(n12893));
  jxor g12635(.dina(n12893), .dinb(n12889), .dout(n12894));
  jor  g12636(.dina(n7408), .dinb(n1566), .dout(n12895));
  jor  g12637(.dina(n1489), .dinb(n7129), .dout(n12896));
  jor  g12638(.dina(n1569), .dinb(n7149), .dout(n12897));
  jor  g12639(.dina(n1571), .dinb(n7411), .dout(n12898));
  jand g12640(.dina(n12898), .dinb(n12897), .dout(n12899));
  jand g12641(.dina(n12899), .dinb(n12896), .dout(n12900));
  jand g12642(.dina(n12900), .dinb(n12895), .dout(n12901));
  jxor g12643(.dina(n12901), .dinb(a20 ), .dout(n12902));
  jor  g12644(.dina(n12596), .dinb(n12592), .dout(n12903));
  jand g12645(.dina(n12809), .dinb(n12597), .dout(n12904));
  jnot g12646(.din(n12904), .dout(n12905));
  jand g12647(.dina(n12905), .dinb(n12903), .dout(n12906));
  jxor g12648(.dina(n12906), .dinb(n12902), .dout(n12907));
  jnot g12649(.din(n12605), .dout(n12908));
  jnot g12650(.din(n12610), .dout(n12909));
  jand g12651(.dina(n12909), .dinb(n12908), .dout(n12910));
  jand g12652(.dina(n12794), .dinb(n12611), .dout(n12911));
  jor  g12653(.dina(n12911), .dinb(n12910), .dout(n12912));
  jnot g12654(.din(n12912), .dout(n12913));
  jor  g12655(.dina(n6103), .dinb(n2319), .dout(n12914));
  jor  g12656(.dina(n2224), .dinb(n5428), .dout(n12915));
  jor  g12657(.dina(n2322), .dinb(n5862), .dout(n12916));
  jor  g12658(.dina(n2324), .dinb(n6106), .dout(n12917));
  jand g12659(.dina(n12917), .dinb(n12916), .dout(n12918));
  jand g12660(.dina(n12918), .dinb(n12915), .dout(n12919));
  jand g12661(.dina(n12919), .dinb(n12914), .dout(n12920));
  jxor g12662(.dina(n12920), .dinb(a26 ), .dout(n12921));
  jxor g12663(.dina(n12921), .dinb(n12913), .dout(n12922));
  jor  g12664(.dina(n5405), .dinb(n2784), .dout(n12923));
  jor  g12665(.dina(n2661), .dinb(n4974), .dout(n12924));
  jor  g12666(.dina(n2787), .dinb(n4994), .dout(n12925));
  jor  g12667(.dina(n2789), .dinb(n5408), .dout(n12926));
  jand g12668(.dina(n12926), .dinb(n12925), .dout(n12927));
  jand g12669(.dina(n12927), .dinb(n12924), .dout(n12928));
  jand g12670(.dina(n12928), .dinb(n12923), .dout(n12929));
  jxor g12671(.dina(n12929), .dinb(a29 ), .dout(n12930));
  jnot g12672(.din(n12930), .dout(n12931));
  jand g12673(.dina(n12792), .dinb(n12788), .dout(n12932));
  jand g12674(.dina(n12793), .dinb(n12779), .dout(n12933));
  jor  g12675(.dina(n12933), .dinb(n12932), .dout(n12934));
  jxor g12676(.dina(n12934), .dinb(n12931), .dout(n12935));
  jor  g12677(.dina(n4554), .dinb(n3301), .dout(n12936));
  jor  g12678(.dina(n3136), .dinb(n4340), .dout(n12937));
  jor  g12679(.dina(n3304), .dinb(n4537), .dout(n12938));
  jor  g12680(.dina(n3306), .dinb(n4557), .dout(n12939));
  jand g12681(.dina(n12939), .dinb(n12938), .dout(n12940));
  jand g12682(.dina(n12940), .dinb(n12937), .dout(n12941));
  jand g12683(.dina(n12941), .dinb(n12936), .dout(n12942));
  jxor g12684(.dina(n12942), .dinb(a32 ), .dout(n12943));
  jand g12685(.dina(n12770), .dinb(n12620), .dout(n12944));
  jnot g12686(.din(n12944), .dout(n12945));
  jor  g12687(.dina(n12778), .dinb(n12772), .dout(n12946));
  jand g12688(.dina(n12946), .dinb(n12945), .dout(n12947));
  jxor g12689(.dina(n12947), .dinb(n12943), .dout(n12948));
  jor  g12690(.dina(n4137), .dinb(n3849), .dout(n12949));
  jor  g12691(.dina(n3689), .dinb(n3588), .dout(n12950));
  jor  g12692(.dina(n3852), .dinb(n3942), .dout(n12951));
  jor  g12693(.dina(n3854), .dinb(n4140), .dout(n12952));
  jand g12694(.dina(n12952), .dinb(n12951), .dout(n12953));
  jand g12695(.dina(n12953), .dinb(n12950), .dout(n12954));
  jand g12696(.dina(n12954), .dinb(n12949), .dout(n12955));
  jxor g12697(.dina(n12955), .dinb(a35 ), .dout(n12956));
  jnot g12698(.din(n12956), .dout(n12957));
  jor  g12699(.dina(n12768), .dinb(n12633), .dout(n12958));
  jand g12700(.dina(n12769), .dinb(n12625), .dout(n12959));
  jnot g12701(.din(n12959), .dout(n12960));
  jand g12702(.dina(n12960), .dinb(n12958), .dout(n12961));
  jnot g12703(.din(n12961), .dout(n12962));
  jor  g12704(.dina(n4415), .dinb(n3400), .dout(n12963));
  jor  g12705(.dina(n4272), .dinb(n3055), .dout(n12964));
  jor  g12706(.dina(n4418), .dinb(n3230), .dout(n12965));
  jor  g12707(.dina(n4420), .dinb(n3403), .dout(n12966));
  jand g12708(.dina(n12966), .dinb(n12965), .dout(n12967));
  jand g12709(.dina(n12967), .dinb(n12964), .dout(n12968));
  jand g12710(.dina(n12968), .dinb(n12963), .dout(n12969));
  jxor g12711(.dina(n12969), .dinb(a38 ), .dout(n12970));
  jnot g12712(.din(n12970), .dout(n12971));
  jor  g12713(.dina(n12740), .dinb(n12732), .dout(n12972));
  jand g12714(.dina(n12748), .dinb(n12741), .dout(n12973));
  jnot g12715(.din(n12973), .dout(n12974));
  jand g12716(.dina(n12974), .dinb(n12972), .dout(n12975));
  jnot g12717(.din(n12975), .dout(n12976));
  jand g12718(.dina(n12725), .dinb(n12642), .dout(n12977));
  jand g12719(.dina(n12730), .dinb(n12726), .dout(n12978));
  jor  g12720(.dina(n12978), .dinb(n12977), .dout(n12979));
  jor  g12721(.dina(n12723), .dinb(n12715), .dout(n12980));
  jand g12722(.dina(n12724), .dinb(n12647), .dout(n12981));
  jnot g12723(.din(n12981), .dout(n12982));
  jand g12724(.dina(n12982), .dinb(n12980), .dout(n12983));
  jnot g12725(.din(n12983), .dout(n12984));
  jor  g12726(.dina(n12706), .dinb(n12698), .dout(n12985));
  jand g12727(.dina(n12713), .dinb(n12707), .dout(n12986));
  jnot g12728(.din(n12986), .dout(n12987));
  jand g12729(.dina(n12987), .dinb(n12985), .dout(n12988));
  jnot g12730(.din(n12988), .dout(n12989));
  jand g12731(.dina(n12691), .dinb(n12656), .dout(n12990));
  jand g12732(.dina(n12696), .dinb(n12692), .dout(n12991));
  jor  g12733(.dina(n12991), .dinb(n12990), .dout(n12992));
  jand g12734(.dina(n12689), .dinb(n12670), .dout(n12993));
  jand g12735(.dina(n12690), .dinb(n12661), .dout(n12994));
  jor  g12736(.dina(n12994), .dinb(n12993), .dout(n12995));
  jand g12737(.dina(n12678), .dinb(n12673), .dout(n12996));
  jnot g12738(.din(n12996), .dout(n12997));
  jor  g12739(.dina(n12688), .dinb(n12680), .dout(n12998));
  jand g12740(.dina(n12998), .dinb(n12997), .dout(n12999));
  jnot g12741(.din(n12999), .dout(n13000));
  jand g12742(.dina(n364), .dinb(n260), .dout(n13001));
  jand g12743(.dina(n12677), .dinb(n12674), .dout(n13002));
  jor  g12744(.dina(n13002), .dinb(n13001), .dout(n13003));
  jand g12745(.dina(n10801), .dinb(b7 ), .dout(n13004));
  jand g12746(.dina(n11107), .dinb(b6 ), .dout(n13005));
  jor  g12747(.dina(n13005), .dinb(n13004), .dout(n13006));
  jnot g12748(.din(n13006), .dout(n13007));
  jxor g12749(.dina(n13007), .dinb(n13003), .dout(n13008));
  jnot g12750(.din(n13008), .dout(n13009));
  jor  g12751(.dina(n10806), .dinb(n624), .dout(n13010));
  jor  g12752(.dina(n10485), .dinb(n512), .dout(n13011));
  jor  g12753(.dina(n10809), .dinb(n564), .dout(n13012));
  jor  g12754(.dina(n10811), .dinb(n627), .dout(n13013));
  jand g12755(.dina(n13013), .dinb(n13012), .dout(n13014));
  jand g12756(.dina(n13014), .dinb(n13011), .dout(n13015));
  jand g12757(.dina(n13015), .dinb(n13010), .dout(n13016));
  jxor g12758(.dina(n13016), .dinb(a62 ), .dout(n13017));
  jxor g12759(.dina(n13017), .dinb(n13009), .dout(n13018));
  jxor g12760(.dina(n13018), .dinb(n13000), .dout(n13019));
  jor  g12761(.dina(n9891), .dinb(n775), .dout(n13020));
  jor  g12762(.dina(n9593), .dinb(n647), .dout(n13021));
  jor  g12763(.dina(n9894), .dinb(n758), .dout(n13022));
  jor  g12764(.dina(n9896), .dinb(n778), .dout(n13023));
  jand g12765(.dina(n13023), .dinb(n13022), .dout(n13024));
  jand g12766(.dina(n13024), .dinb(n13021), .dout(n13025));
  jand g12767(.dina(n13025), .dinb(n13020), .dout(n13026));
  jxor g12768(.dina(n13026), .dinb(a59 ), .dout(n13027));
  jnot g12769(.din(n13027), .dout(n13028));
  jxor g12770(.dina(n13028), .dinb(n13019), .dout(n13029));
  jxor g12771(.dina(n13029), .dinb(n12995), .dout(n13030));
  jor  g12772(.dina(n8978), .dinb(n1019), .dout(n13031));
  jor  g12773(.dina(n8677), .dinb(n858), .dout(n13032));
  jor  g12774(.dina(n8981), .dinb(n939), .dout(n13033));
  jor  g12775(.dina(n8983), .dinb(n1022), .dout(n13034));
  jand g12776(.dina(n13034), .dinb(n13033), .dout(n13035));
  jand g12777(.dina(n13035), .dinb(n13032), .dout(n13036));
  jand g12778(.dina(n13036), .dinb(n13031), .dout(n13037));
  jxor g12779(.dina(n13037), .dinb(a56 ), .dout(n13038));
  jnot g12780(.din(n13038), .dout(n13039));
  jxor g12781(.dina(n13039), .dinb(n13030), .dout(n13040));
  jxor g12782(.dina(n13040), .dinb(n12992), .dout(n13041));
  jor  g12783(.dina(n8125), .dinb(n1397), .dout(n13042));
  jor  g12784(.dina(n7846), .dinb(n1193), .dout(n13043));
  jor  g12785(.dina(n8128), .dinb(n1290), .dout(n13044));
  jor  g12786(.dina(n8130), .dinb(n1400), .dout(n13045));
  jand g12787(.dina(n13045), .dinb(n13044), .dout(n13046));
  jand g12788(.dina(n13046), .dinb(n13043), .dout(n13047));
  jand g12789(.dina(n13047), .dinb(n13042), .dout(n13048));
  jxor g12790(.dina(n13048), .dinb(a53 ), .dout(n13049));
  jnot g12791(.din(n13049), .dout(n13050));
  jxor g12792(.dina(n13050), .dinb(n13041), .dout(n13051));
  jxor g12793(.dina(n13051), .dinb(n12989), .dout(n13052));
  jor  g12794(.dina(n7266), .dinb(n1739), .dout(n13053));
  jor  g12795(.dina(n7021), .dinb(n1420), .dout(n13054));
  jor  g12796(.dina(n7269), .dinb(n1620), .dout(n13055));
  jor  g12797(.dina(n7271), .dinb(n1742), .dout(n13056));
  jand g12798(.dina(n13056), .dinb(n13055), .dout(n13057));
  jand g12799(.dina(n13057), .dinb(n13054), .dout(n13058));
  jand g12800(.dina(n13058), .dinb(n13053), .dout(n13059));
  jxor g12801(.dina(n13059), .dinb(a50 ), .dout(n13060));
  jnot g12802(.din(n13060), .dout(n13061));
  jxor g12803(.dina(n13061), .dinb(n13052), .dout(n13062));
  jxor g12804(.dina(n13062), .dinb(n12984), .dout(n13063));
  jor  g12805(.dina(n6490), .dinb(n2007), .dout(n13064));
  jor  g12806(.dina(n6262), .dinb(n1867), .dout(n13065));
  jor  g12807(.dina(n6493), .dinb(n1887), .dout(n13066));
  jor  g12808(.dina(n6495), .dinb(n2010), .dout(n13067));
  jand g12809(.dina(n13067), .dinb(n13066), .dout(n13068));
  jand g12810(.dina(n13068), .dinb(n13065), .dout(n13069));
  jand g12811(.dina(n13069), .dinb(n13064), .dout(n13070));
  jxor g12812(.dina(n13070), .dinb(a47 ), .dout(n13071));
  jnot g12813(.din(n13071), .dout(n13072));
  jxor g12814(.dina(n13072), .dinb(n13063), .dout(n13073));
  jxor g12815(.dina(n13073), .dinb(n12979), .dout(n13074));
  jor  g12816(.dina(n5739), .dinb(n2556), .dout(n13075));
  jor  g12817(.dina(n5574), .dinb(n2148), .dout(n13076));
  jor  g12818(.dina(n5742), .dinb(n2407), .dout(n13077));
  jor  g12819(.dina(n5744), .dinb(n2559), .dout(n13078));
  jand g12820(.dina(n13078), .dinb(n13077), .dout(n13079));
  jand g12821(.dina(n13079), .dinb(n13076), .dout(n13080));
  jand g12822(.dina(n13080), .dinb(n13075), .dout(n13081));
  jxor g12823(.dina(n13081), .dinb(a44 ), .dout(n13082));
  jnot g12824(.din(n13082), .dout(n13083));
  jxor g12825(.dina(n13083), .dinb(n13074), .dout(n13084));
  jxor g12826(.dina(n13084), .dinb(n12976), .dout(n13085));
  jnot g12827(.din(n13085), .dout(n13086));
  jor  g12828(.dina(n5096), .dinb(n3032), .dout(n13087));
  jor  g12829(.dina(n4904), .dinb(n2579), .dout(n13088));
  jor  g12830(.dina(n5099), .dinb(n2870), .dout(n13089));
  jor  g12831(.dina(n5101), .dinb(n3035), .dout(n13090));
  jand g12832(.dina(n13090), .dinb(n13089), .dout(n13091));
  jand g12833(.dina(n13091), .dinb(n13088), .dout(n13092));
  jand g12834(.dina(n13092), .dinb(n13087), .dout(n13093));
  jxor g12835(.dina(n13093), .dinb(a41 ), .dout(n13094));
  jxor g12836(.dina(n13094), .dinb(n13086), .dout(n13095));
  jand g12837(.dina(n12758), .dinb(n12750), .dout(n13096));
  jnot g12838(.din(n13096), .dout(n13097));
  jnot g12839(.din(n12758), .dout(n13098));
  jand g12840(.dina(n13098), .dinb(n12749), .dout(n13099));
  jor  g12841(.dina(n12767), .dinb(n13099), .dout(n13100));
  jand g12842(.dina(n13100), .dinb(n13097), .dout(n13101));
  jxor g12843(.dina(n13101), .dinb(n13095), .dout(n13102));
  jxor g12844(.dina(n13102), .dinb(n12971), .dout(n13103));
  jxor g12845(.dina(n13103), .dinb(n12962), .dout(n13104));
  jxor g12846(.dina(n13104), .dinb(n12957), .dout(n13105));
  jxor g12847(.dina(n13105), .dinb(n12948), .dout(n13106));
  jxor g12848(.dina(n13106), .dinb(n12935), .dout(n13107));
  jxor g12849(.dina(n13107), .dinb(n12922), .dout(n13108));
  jor  g12850(.dina(n6864), .dinb(n1939), .dout(n13109));
  jor  g12851(.dina(n1827), .dinb(n6352), .dout(n13110));
  jor  g12852(.dina(n1942), .dinb(n6372), .dout(n13111));
  jor  g12853(.dina(n1944), .dinb(n6867), .dout(n13112));
  jand g12854(.dina(n13112), .dinb(n13111), .dout(n13113));
  jand g12855(.dina(n13113), .dinb(n13110), .dout(n13114));
  jand g12856(.dina(n13114), .dinb(n13109), .dout(n13115));
  jxor g12857(.dina(n13115), .dinb(a23 ), .dout(n13116));
  jor  g12858(.dina(n12807), .dinb(n12799), .dout(n13117));
  jand g12859(.dina(n12808), .dinb(n12795), .dout(n13118));
  jnot g12860(.din(n13118), .dout(n13119));
  jand g12861(.dina(n13119), .dinb(n13117), .dout(n13120));
  jxor g12862(.dina(n13120), .dinb(n13116), .dout(n13121));
  jxor g12863(.dina(n13121), .dinb(n13108), .dout(n13122));
  jxor g12864(.dina(n13122), .dinb(n12907), .dout(n13123));
  jxor g12865(.dina(n13123), .dinb(n12894), .dout(n13124));
  jxor g12866(.dina(n13124), .dinb(n12881), .dout(n13125));
  jxor g12867(.dina(n13125), .dinb(n12868), .dout(n13126));
  jxor g12868(.dina(n13126), .dinb(n12852), .dout(n13127));
  jxor g12869(.dina(n13127), .dinb(n12838), .dout(n13128));
  jxor g12870(.dina(n13128), .dinb(n12833), .dout(f70 ));
  jand g12871(.dina(n13127), .dinb(n12838), .dout(n13130));
  jand g12872(.dina(n13128), .dinb(n12833), .dout(n13131));
  jor  g12873(.dina(n13131), .dinb(n13130), .dout(n13132));
  jor  g12874(.dina(n8786), .dinb(n1245), .dout(n13133));
  jor  g12875(.dina(n1165), .dinb(n7960), .dout(n13134));
  jor  g12876(.dina(n1248), .dinb(n8231), .dout(n13135));
  jor  g12877(.dina(n1250), .dinb(n8789), .dout(n13136));
  jand g12878(.dina(n13136), .dinb(n13135), .dout(n13137));
  jand g12879(.dina(n13137), .dinb(n13134), .dout(n13138));
  jand g12880(.dina(n13138), .dinb(n13133), .dout(n13139));
  jxor g12881(.dina(n13139), .dinb(a17 ), .dout(n13140));
  jor  g12882(.dina(n12906), .dinb(n12902), .dout(n13141));
  jand g12883(.dina(n13122), .dinb(n12907), .dout(n13142));
  jnot g12884(.din(n13142), .dout(n13143));
  jand g12885(.dina(n13143), .dinb(n13141), .dout(n13144));
  jxor g12886(.dina(n13144), .dinb(n13140), .dout(n13145));
  jor  g12887(.dina(n7126), .dinb(n1939), .dout(n13146));
  jor  g12888(.dina(n1827), .dinb(n6372), .dout(n13147));
  jor  g12889(.dina(n1942), .dinb(n6867), .dout(n13148));
  jor  g12890(.dina(n1944), .dinb(n7129), .dout(n13149));
  jand g12891(.dina(n13149), .dinb(n13148), .dout(n13150));
  jand g12892(.dina(n13150), .dinb(n13147), .dout(n13151));
  jand g12893(.dina(n13151), .dinb(n13146), .dout(n13152));
  jxor g12894(.dina(n13152), .dinb(a23 ), .dout(n13153));
  jor  g12895(.dina(n12921), .dinb(n12913), .dout(n13154));
  jand g12896(.dina(n13107), .dinb(n12922), .dout(n13155));
  jnot g12897(.din(n13155), .dout(n13156));
  jand g12898(.dina(n13156), .dinb(n13154), .dout(n13157));
  jxor g12899(.dina(n13157), .dinb(n13153), .dout(n13158));
  jor  g12900(.dina(n6349), .dinb(n2319), .dout(n13159));
  jor  g12901(.dina(n2224), .dinb(n5862), .dout(n13160));
  jor  g12902(.dina(n2322), .dinb(n6106), .dout(n13161));
  jor  g12903(.dina(n2324), .dinb(n6352), .dout(n13162));
  jand g12904(.dina(n13162), .dinb(n13161), .dout(n13163));
  jand g12905(.dina(n13163), .dinb(n13160), .dout(n13164));
  jand g12906(.dina(n13164), .dinb(n13159), .dout(n13165));
  jxor g12907(.dina(n13165), .dinb(a26 ), .dout(n13166));
  jnot g12908(.din(n13166), .dout(n13167));
  jand g12909(.dina(n12934), .dinb(n12931), .dout(n13168));
  jand g12910(.dina(n13106), .dinb(n12935), .dout(n13169));
  jor  g12911(.dina(n13169), .dinb(n13168), .dout(n13170));
  jxor g12912(.dina(n13170), .dinb(n13167), .dout(n13171));
  jor  g12913(.dina(n4971), .dinb(n3301), .dout(n13172));
  jor  g12914(.dina(n3136), .dinb(n4537), .dout(n13173));
  jor  g12915(.dina(n3304), .dinb(n4557), .dout(n13174));
  jor  g12916(.dina(n3306), .dinb(n4974), .dout(n13175));
  jand g12917(.dina(n13175), .dinb(n13174), .dout(n13176));
  jand g12918(.dina(n13176), .dinb(n13173), .dout(n13177));
  jand g12919(.dina(n13177), .dinb(n13172), .dout(n13178));
  jxor g12920(.dina(n13178), .dinb(a32 ), .dout(n13179));
  jnot g12921(.din(n13179), .dout(n13180));
  jor  g12922(.dina(n13103), .dinb(n12962), .dout(n13181));
  jand g12923(.dina(n13103), .dinb(n12962), .dout(n13182));
  jor  g12924(.dina(n13182), .dinb(n12957), .dout(n13183));
  jand g12925(.dina(n13183), .dinb(n13181), .dout(n13184));
  jxor g12926(.dina(n13184), .dinb(n13180), .dout(n13185));
  jand g12927(.dina(n13101), .dinb(n13095), .dout(n13186));
  jand g12928(.dina(n13102), .dinb(n12971), .dout(n13187));
  jor  g12929(.dina(n13187), .dinb(n13186), .dout(n13188));
  jor  g12930(.dina(n7266), .dinb(n1864), .dout(n13189));
  jor  g12931(.dina(n7021), .dinb(n1620), .dout(n13190));
  jor  g12932(.dina(n7269), .dinb(n1742), .dout(n13191));
  jor  g12933(.dina(n7271), .dinb(n1867), .dout(n13192));
  jand g12934(.dina(n13192), .dinb(n13191), .dout(n13193));
  jand g12935(.dina(n13193), .dinb(n13190), .dout(n13194));
  jand g12936(.dina(n13194), .dinb(n13189), .dout(n13195));
  jxor g12937(.dina(n13195), .dinb(a50 ), .dout(n13196));
  jnot g12938(.din(n13196), .dout(n13197));
  jor  g12939(.dina(n9891), .dinb(n855), .dout(n13198));
  jor  g12940(.dina(n9593), .dinb(n758), .dout(n13199));
  jor  g12941(.dina(n9894), .dinb(n778), .dout(n13200));
  jor  g12942(.dina(n9896), .dinb(n858), .dout(n13201));
  jand g12943(.dina(n13201), .dinb(n13200), .dout(n13202));
  jand g12944(.dina(n13202), .dinb(n13199), .dout(n13203));
  jand g12945(.dina(n13203), .dinb(n13198), .dout(n13204));
  jxor g12946(.dina(n13204), .dinb(a59 ), .dout(n13205));
  jnot g12947(.din(n13205), .dout(n13206));
  jor  g12948(.dina(n10806), .dinb(n644), .dout(n13207));
  jor  g12949(.dina(n10485), .dinb(n564), .dout(n13208));
  jor  g12950(.dina(n10809), .dinb(n627), .dout(n13209));
  jor  g12951(.dina(n10811), .dinb(n647), .dout(n13210));
  jand g12952(.dina(n13210), .dinb(n13209), .dout(n13211));
  jand g12953(.dina(n13211), .dinb(n13208), .dout(n13212));
  jand g12954(.dina(n13212), .dinb(n13207), .dout(n13213));
  jxor g12955(.dina(n13213), .dinb(a62 ), .dout(n13214));
  jnot g12956(.din(n13214), .dout(n13215));
  jand g12957(.dina(n13007), .dinb(n13003), .dout(n13216));
  jnot g12958(.din(n13216), .dout(n13217));
  jor  g12959(.dina(n13017), .dinb(n13009), .dout(n13218));
  jand g12960(.dina(n13218), .dinb(n13217), .dout(n13219));
  jnot g12961(.din(n13219), .dout(n13220));
  jand g12962(.dina(n10801), .dinb(b8 ), .dout(n13221));
  jand g12963(.dina(n11107), .dinb(b7 ), .dout(n13222));
  jor  g12964(.dina(n13222), .dinb(n13221), .dout(n13223));
  jnot g12965(.din(n13223), .dout(n13224));
  jxor g12966(.dina(n13224), .dinb(n13006), .dout(n13225));
  jxor g12967(.dina(n13225), .dinb(n13220), .dout(n13226));
  jxor g12968(.dina(n13226), .dinb(n13215), .dout(n13227));
  jxor g12969(.dina(n13227), .dinb(n13206), .dout(n13228));
  jor  g12970(.dina(n13018), .dinb(n13000), .dout(n13229));
  jand g12971(.dina(n13018), .dinb(n13000), .dout(n13230));
  jor  g12972(.dina(n13028), .dinb(n13230), .dout(n13231));
  jand g12973(.dina(n13231), .dinb(n13229), .dout(n13232));
  jxor g12974(.dina(n13232), .dinb(n13228), .dout(n13233));
  jor  g12975(.dina(n8978), .dinb(n1190), .dout(n13234));
  jor  g12976(.dina(n8677), .dinb(n939), .dout(n13235));
  jor  g12977(.dina(n8981), .dinb(n1022), .dout(n13236));
  jor  g12978(.dina(n8983), .dinb(n1193), .dout(n13237));
  jand g12979(.dina(n13237), .dinb(n13236), .dout(n13238));
  jand g12980(.dina(n13238), .dinb(n13235), .dout(n13239));
  jand g12981(.dina(n13239), .dinb(n13234), .dout(n13240));
  jxor g12982(.dina(n13240), .dinb(a56 ), .dout(n13241));
  jnot g12983(.din(n13241), .dout(n13242));
  jxor g12984(.dina(n13242), .dinb(n13233), .dout(n13243));
  jnot g12985(.din(n12995), .dout(n13244));
  jnot g12986(.din(n13029), .dout(n13245));
  jand g12987(.dina(n13245), .dinb(n13244), .dout(n13246));
  jnot g12988(.din(n13246), .dout(n13247));
  jand g12989(.dina(n13029), .dinb(n12995), .dout(n13248));
  jor  g12990(.dina(n13039), .dinb(n13248), .dout(n13249));
  jand g12991(.dina(n13249), .dinb(n13247), .dout(n13250));
  jxor g12992(.dina(n13250), .dinb(n13243), .dout(n13251));
  jnot g12993(.din(n13251), .dout(n13252));
  jor  g12994(.dina(n8125), .dinb(n1417), .dout(n13253));
  jor  g12995(.dina(n7846), .dinb(n1290), .dout(n13254));
  jor  g12996(.dina(n8128), .dinb(n1400), .dout(n13255));
  jor  g12997(.dina(n8130), .dinb(n1420), .dout(n13256));
  jand g12998(.dina(n13256), .dinb(n13255), .dout(n13257));
  jand g12999(.dina(n13257), .dinb(n13254), .dout(n13258));
  jand g13000(.dina(n13258), .dinb(n13253), .dout(n13259));
  jxor g13001(.dina(n13259), .dinb(a53 ), .dout(n13260));
  jxor g13002(.dina(n13260), .dinb(n13252), .dout(n13261));
  jnot g13003(.din(n12992), .dout(n13262));
  jnot g13004(.din(n13040), .dout(n13263));
  jand g13005(.dina(n13263), .dinb(n13262), .dout(n13264));
  jnot g13006(.din(n13264), .dout(n13265));
  jand g13007(.dina(n13040), .dinb(n12992), .dout(n13266));
  jor  g13008(.dina(n13050), .dinb(n13266), .dout(n13267));
  jand g13009(.dina(n13267), .dinb(n13265), .dout(n13268));
  jxor g13010(.dina(n13268), .dinb(n13261), .dout(n13269));
  jxor g13011(.dina(n13269), .dinb(n13197), .dout(n13270));
  jnot g13012(.din(n13051), .dout(n13271));
  jand g13013(.dina(n13271), .dinb(n12988), .dout(n13272));
  jnot g13014(.din(n13272), .dout(n13273));
  jand g13015(.dina(n13051), .dinb(n12989), .dout(n13274));
  jor  g13016(.dina(n13061), .dinb(n13274), .dout(n13275));
  jand g13017(.dina(n13275), .dinb(n13273), .dout(n13276));
  jxor g13018(.dina(n13276), .dinb(n13270), .dout(n13277));
  jor  g13019(.dina(n6490), .dinb(n2145), .dout(n13278));
  jor  g13020(.dina(n6262), .dinb(n1887), .dout(n13279));
  jor  g13021(.dina(n6493), .dinb(n2010), .dout(n13280));
  jor  g13022(.dina(n6495), .dinb(n2148), .dout(n13281));
  jand g13023(.dina(n13281), .dinb(n13280), .dout(n13282));
  jand g13024(.dina(n13282), .dinb(n13279), .dout(n13283));
  jand g13025(.dina(n13283), .dinb(n13278), .dout(n13284));
  jxor g13026(.dina(n13284), .dinb(a47 ), .dout(n13285));
  jnot g13027(.din(n13285), .dout(n13286));
  jxor g13028(.dina(n13286), .dinb(n13277), .dout(n13287));
  jnot g13029(.din(n13062), .dout(n13288));
  jand g13030(.dina(n13288), .dinb(n12983), .dout(n13289));
  jnot g13031(.din(n13289), .dout(n13290));
  jand g13032(.dina(n13062), .dinb(n12984), .dout(n13291));
  jor  g13033(.dina(n13072), .dinb(n13291), .dout(n13292));
  jand g13034(.dina(n13292), .dinb(n13290), .dout(n13293));
  jxor g13035(.dina(n13293), .dinb(n13287), .dout(n13294));
  jor  g13036(.dina(n5739), .dinb(n2576), .dout(n13295));
  jor  g13037(.dina(n5574), .dinb(n2407), .dout(n13296));
  jor  g13038(.dina(n5742), .dinb(n2559), .dout(n13297));
  jor  g13039(.dina(n5744), .dinb(n2579), .dout(n13298));
  jand g13040(.dina(n13298), .dinb(n13297), .dout(n13299));
  jand g13041(.dina(n13299), .dinb(n13296), .dout(n13300));
  jand g13042(.dina(n13300), .dinb(n13295), .dout(n13301));
  jxor g13043(.dina(n13301), .dinb(a44 ), .dout(n13302));
  jnot g13044(.din(n13302), .dout(n13303));
  jxor g13045(.dina(n13303), .dinb(n13294), .dout(n13304));
  jnot g13046(.din(n12979), .dout(n13305));
  jnot g13047(.din(n13073), .dout(n13306));
  jand g13048(.dina(n13306), .dinb(n13305), .dout(n13307));
  jnot g13049(.din(n13307), .dout(n13308));
  jand g13050(.dina(n13073), .dinb(n12979), .dout(n13309));
  jor  g13051(.dina(n13083), .dinb(n13309), .dout(n13310));
  jand g13052(.dina(n13310), .dinb(n13308), .dout(n13311));
  jxor g13053(.dina(n13311), .dinb(n13304), .dout(n13312));
  jnot g13054(.din(n13312), .dout(n13313));
  jor  g13055(.dina(n5096), .dinb(n3052), .dout(n13314));
  jor  g13056(.dina(n4904), .dinb(n2870), .dout(n13315));
  jor  g13057(.dina(n5099), .dinb(n3035), .dout(n13316));
  jor  g13058(.dina(n5101), .dinb(n3055), .dout(n13317));
  jand g13059(.dina(n13317), .dinb(n13316), .dout(n13318));
  jand g13060(.dina(n13318), .dinb(n13315), .dout(n13319));
  jand g13061(.dina(n13319), .dinb(n13314), .dout(n13320));
  jxor g13062(.dina(n13320), .dinb(a41 ), .dout(n13321));
  jxor g13063(.dina(n13321), .dinb(n13313), .dout(n13322));
  jand g13064(.dina(n13084), .dinb(n12976), .dout(n13323));
  jnot g13065(.din(n13323), .dout(n13324));
  jor  g13066(.dina(n13094), .dinb(n13086), .dout(n13325));
  jand g13067(.dina(n13325), .dinb(n13324), .dout(n13326));
  jnot g13068(.din(n13326), .dout(n13327));
  jxor g13069(.dina(n13327), .dinb(n13322), .dout(n13328));
  jnot g13070(.din(n13328), .dout(n13329));
  jor  g13071(.dina(n4415), .dinb(n3585), .dout(n13330));
  jor  g13072(.dina(n4272), .dinb(n3230), .dout(n13331));
  jor  g13073(.dina(n4418), .dinb(n3403), .dout(n13332));
  jor  g13074(.dina(n4420), .dinb(n3588), .dout(n13333));
  jand g13075(.dina(n13333), .dinb(n13332), .dout(n13334));
  jand g13076(.dina(n13334), .dinb(n13331), .dout(n13335));
  jand g13077(.dina(n13335), .dinb(n13330), .dout(n13336));
  jxor g13078(.dina(n13336), .dinb(a38 ), .dout(n13337));
  jxor g13079(.dina(n13337), .dinb(n13329), .dout(n13338));
  jxor g13080(.dina(n13338), .dinb(n13188), .dout(n13339));
  jnot g13081(.din(n13339), .dout(n13340));
  jor  g13082(.dina(n4337), .dinb(n3849), .dout(n13341));
  jor  g13083(.dina(n3689), .dinb(n3942), .dout(n13342));
  jor  g13084(.dina(n3852), .dinb(n4140), .dout(n13343));
  jor  g13085(.dina(n3854), .dinb(n4340), .dout(n13344));
  jand g13086(.dina(n13344), .dinb(n13343), .dout(n13345));
  jand g13087(.dina(n13345), .dinb(n13342), .dout(n13346));
  jand g13088(.dina(n13346), .dinb(n13341), .dout(n13347));
  jxor g13089(.dina(n13347), .dinb(a35 ), .dout(n13348));
  jxor g13090(.dina(n13348), .dinb(n13340), .dout(n13349));
  jxor g13091(.dina(n13349), .dinb(n13185), .dout(n13350));
  jor  g13092(.dina(n5425), .dinb(n2784), .dout(n13351));
  jor  g13093(.dina(n2661), .dinb(n4994), .dout(n13352));
  jor  g13094(.dina(n2787), .dinb(n5408), .dout(n13353));
  jor  g13095(.dina(n2789), .dinb(n5428), .dout(n13354));
  jand g13096(.dina(n13354), .dinb(n13353), .dout(n13355));
  jand g13097(.dina(n13355), .dinb(n13352), .dout(n13356));
  jand g13098(.dina(n13356), .dinb(n13351), .dout(n13357));
  jxor g13099(.dina(n13357), .dinb(a29 ), .dout(n13358));
  jand g13100(.dina(n12947), .dinb(n12943), .dout(n13359));
  jor  g13101(.dina(n12947), .dinb(n12943), .dout(n13360));
  jnot g13102(.din(n13105), .dout(n13361));
  jand g13103(.dina(n13361), .dinb(n13360), .dout(n13362));
  jor  g13104(.dina(n13362), .dinb(n13359), .dout(n13363));
  jxor g13105(.dina(n13363), .dinb(n13358), .dout(n13364));
  jxor g13106(.dina(n13364), .dinb(n13350), .dout(n13365));
  jxor g13107(.dina(n13365), .dinb(n13171), .dout(n13366));
  jxor g13108(.dina(n13366), .dinb(n13158), .dout(n13367));
  jor  g13109(.dina(n13120), .dinb(n13116), .dout(n13368));
  jand g13110(.dina(n13121), .dinb(n13108), .dout(n13369));
  jnot g13111(.din(n13369), .dout(n13370));
  jand g13112(.dina(n13370), .dinb(n13368), .dout(n13371));
  jor  g13113(.dina(n7680), .dinb(n1566), .dout(n13372));
  jor  g13114(.dina(n1489), .dinb(n7149), .dout(n13373));
  jor  g13115(.dina(n1569), .dinb(n7411), .dout(n13374));
  jor  g13116(.dina(n1571), .dinb(n7683), .dout(n13375));
  jand g13117(.dina(n13375), .dinb(n13374), .dout(n13376));
  jand g13118(.dina(n13376), .dinb(n13373), .dout(n13377));
  jand g13119(.dina(n13377), .dinb(n13372), .dout(n13378));
  jxor g13120(.dina(n13378), .dinb(a20 ), .dout(n13379));
  jxor g13121(.dina(n13379), .dinb(n13371), .dout(n13380));
  jxor g13122(.dina(n13380), .dinb(n13367), .dout(n13381));
  jnot g13123(.din(n13381), .dout(n13382));
  jxor g13124(.dina(n13382), .dinb(n13145), .dout(n13383));
  jor  g13125(.dina(n9410), .dinb(n974), .dout(n13384));
  jor  g13126(.dina(n908), .dinb(n8809), .dout(n13385));
  jor  g13127(.dina(n977), .dinb(n9390), .dout(n13386));
  jor  g13128(.dina(n979), .dinb(n9413), .dout(n13387));
  jand g13129(.dina(n13387), .dinb(n13386), .dout(n13388));
  jand g13130(.dina(n13388), .dinb(n13385), .dout(n13389));
  jand g13131(.dina(n13389), .dinb(n13384), .dout(n13390));
  jxor g13132(.dina(n13390), .dinb(a14 ), .dout(n13391));
  jor  g13133(.dina(n12893), .dinb(n12889), .dout(n13392));
  jand g13134(.dina(n13123), .dinb(n12894), .dout(n13393));
  jnot g13135(.din(n13393), .dout(n13394));
  jand g13136(.dina(n13394), .dinb(n13392), .dout(n13395));
  jxor g13137(.dina(n13395), .dinb(n13391), .dout(n13396));
  jxor g13138(.dina(n13396), .dinb(n13383), .dout(n13397));
  jnot g13139(.din(n12872), .dout(n13398));
  jor  g13140(.dina(n12880), .dinb(n13398), .dout(n13399));
  jnot g13141(.din(n13124), .dout(n13400));
  jor  g13142(.dina(n13400), .dinb(n12881), .dout(n13401));
  jand g13143(.dina(n13401), .dinb(n13399), .dout(n13402));
  jor  g13144(.dina(n10634), .dinb(n706), .dout(n13403));
  jor  g13145(.dina(n683), .dinb(n9725), .dout(n13404));
  jor  g13146(.dina(n709), .dinb(n10314), .dout(n13405));
  jor  g13147(.dina(n711), .dinb(n10637), .dout(n13406));
  jand g13148(.dina(n13406), .dinb(n13405), .dout(n13407));
  jand g13149(.dina(n13407), .dinb(n13404), .dout(n13408));
  jand g13150(.dina(n13408), .dinb(n13403), .dout(n13409));
  jxor g13151(.dina(n13409), .dinb(a11 ), .dout(n13410));
  jnot g13152(.din(n13410), .dout(n13411));
  jxor g13153(.dina(n13411), .dinb(n13402), .dout(n13412));
  jxor g13154(.dina(n13412), .dinb(n13397), .dout(n13413));
  jnot g13155(.din(n12860), .dout(n13414));
  jand g13156(.dina(n12867), .dinb(n13414), .dout(n13415));
  jnot g13157(.din(n13415), .dout(n13416));
  jor  g13158(.dina(n13125), .dinb(n12868), .dout(n13417));
  jand g13159(.dina(n13417), .dinb(n13416), .dout(n13418));
  jand g13160(.dina(n11296), .dinb(n458), .dout(n13419));
  jor  g13161(.dina(n13419), .dinb(n491), .dout(n13420));
  jand g13162(.dina(n13420), .dinb(b63 ), .dout(n13421));
  jxor g13163(.dina(n13421), .dinb(n483), .dout(n13422));
  jxor g13164(.dina(n13422), .dinb(n13418), .dout(n13423));
  jxor g13165(.dina(n13423), .dinb(n13413), .dout(n13424));
  jor  g13166(.dina(n12851), .dinb(n12845), .dout(n13425));
  jand g13167(.dina(n12851), .dinb(n12845), .dout(n13426));
  jor  g13168(.dina(n13126), .dinb(n13426), .dout(n13427));
  jand g13169(.dina(n13427), .dinb(n13425), .dout(n13428));
  jxor g13170(.dina(n13428), .dinb(n13424), .dout(n13429));
  jxor g13171(.dina(n13429), .dinb(n13132), .dout(f71 ));
  jand g13172(.dina(n13428), .dinb(n13424), .dout(n13431));
  jand g13173(.dina(n13429), .dinb(n13132), .dout(n13432));
  jor  g13174(.dina(n13432), .dinb(n13431), .dout(n13433));
  jor  g13175(.dina(n13422), .dinb(n13418), .dout(n13434));
  jnot g13176(.din(n13434), .dout(n13435));
  jand g13177(.dina(n13423), .dinb(n13413), .dout(n13436));
  jor  g13178(.dina(n13436), .dinb(n13435), .dout(n13437));
  jor  g13179(.dina(n8806), .dinb(n1245), .dout(n13438));
  jor  g13180(.dina(n1165), .dinb(n8231), .dout(n13439));
  jor  g13181(.dina(n1248), .dinb(n8789), .dout(n13440));
  jor  g13182(.dina(n1250), .dinb(n8809), .dout(n13441));
  jand g13183(.dina(n13441), .dinb(n13440), .dout(n13442));
  jand g13184(.dina(n13442), .dinb(n13439), .dout(n13443));
  jand g13185(.dina(n13443), .dinb(n13438), .dout(n13444));
  jxor g13186(.dina(n13444), .dinb(a17 ), .dout(n13445));
  jand g13187(.dina(n13144), .dinb(n13140), .dout(n13446));
  jor  g13188(.dina(n13144), .dinb(n13140), .dout(n13447));
  jand g13189(.dina(n13382), .dinb(n13447), .dout(n13448));
  jor  g13190(.dina(n13448), .dinb(n13446), .dout(n13449));
  jxor g13191(.dina(n13449), .dinb(n13445), .dout(n13450));
  jor  g13192(.dina(n7146), .dinb(n1939), .dout(n13451));
  jor  g13193(.dina(n1827), .dinb(n6867), .dout(n13452));
  jor  g13194(.dina(n1942), .dinb(n7129), .dout(n13453));
  jor  g13195(.dina(n1944), .dinb(n7149), .dout(n13454));
  jand g13196(.dina(n13454), .dinb(n13453), .dout(n13455));
  jand g13197(.dina(n13455), .dinb(n13452), .dout(n13456));
  jand g13198(.dina(n13456), .dinb(n13451), .dout(n13457));
  jxor g13199(.dina(n13457), .dinb(a23 ), .dout(n13458));
  jor  g13200(.dina(n13157), .dinb(n13153), .dout(n13459));
  jand g13201(.dina(n13366), .dinb(n13158), .dout(n13460));
  jnot g13202(.din(n13460), .dout(n13461));
  jand g13203(.dina(n13461), .dinb(n13459), .dout(n13462));
  jxor g13204(.dina(n13462), .dinb(n13458), .dout(n13463));
  jor  g13205(.dina(n6369), .dinb(n2319), .dout(n13464));
  jor  g13206(.dina(n2224), .dinb(n6106), .dout(n13465));
  jor  g13207(.dina(n2322), .dinb(n6352), .dout(n13466));
  jor  g13208(.dina(n2324), .dinb(n6372), .dout(n13467));
  jand g13209(.dina(n13467), .dinb(n13466), .dout(n13468));
  jand g13210(.dina(n13468), .dinb(n13465), .dout(n13469));
  jand g13211(.dina(n13469), .dinb(n13464), .dout(n13470));
  jxor g13212(.dina(n13470), .dinb(a26 ), .dout(n13471));
  jnot g13213(.din(n13471), .dout(n13472));
  jand g13214(.dina(n13170), .dinb(n13167), .dout(n13473));
  jand g13215(.dina(n13365), .dinb(n13171), .dout(n13474));
  jor  g13216(.dina(n13474), .dinb(n13473), .dout(n13475));
  jxor g13217(.dina(n13475), .dinb(n13472), .dout(n13476));
  jnot g13218(.din(n13358), .dout(n13477));
  jnot g13219(.din(n13363), .dout(n13478));
  jand g13220(.dina(n13478), .dinb(n13477), .dout(n13479));
  jand g13221(.dina(n13364), .dinb(n13350), .dout(n13480));
  jor  g13222(.dina(n13480), .dinb(n13479), .dout(n13481));
  jnot g13223(.din(n13481), .dout(n13482));
  jor  g13224(.dina(n5859), .dinb(n2784), .dout(n13483));
  jor  g13225(.dina(n2661), .dinb(n5408), .dout(n13484));
  jor  g13226(.dina(n2787), .dinb(n5428), .dout(n13485));
  jor  g13227(.dina(n2789), .dinb(n5862), .dout(n13486));
  jand g13228(.dina(n13486), .dinb(n13485), .dout(n13487));
  jand g13229(.dina(n13487), .dinb(n13484), .dout(n13488));
  jand g13230(.dina(n13488), .dinb(n13483), .dout(n13489));
  jxor g13231(.dina(n13489), .dinb(a29 ), .dout(n13490));
  jxor g13232(.dina(n13490), .dinb(n13482), .dout(n13491));
  jand g13233(.dina(n13338), .dinb(n13188), .dout(n13492));
  jnot g13234(.din(n13492), .dout(n13493));
  jor  g13235(.dina(n13348), .dinb(n13340), .dout(n13494));
  jand g13236(.dina(n13494), .dinb(n13493), .dout(n13495));
  jnot g13237(.din(n13495), .dout(n13496));
  jor  g13238(.dina(n4415), .dinb(n3939), .dout(n13497));
  jor  g13239(.dina(n4272), .dinb(n3403), .dout(n13498));
  jor  g13240(.dina(n4418), .dinb(n3588), .dout(n13499));
  jor  g13241(.dina(n4420), .dinb(n3942), .dout(n13500));
  jand g13242(.dina(n13500), .dinb(n13499), .dout(n13501));
  jand g13243(.dina(n13501), .dinb(n13498), .dout(n13502));
  jand g13244(.dina(n13502), .dinb(n13497), .dout(n13503));
  jxor g13245(.dina(n13503), .dinb(a38 ), .dout(n13504));
  jnot g13246(.din(n13504), .dout(n13505));
  jand g13247(.dina(n13311), .dinb(n13304), .dout(n13506));
  jnot g13248(.din(n13506), .dout(n13507));
  jor  g13249(.dina(n13321), .dinb(n13313), .dout(n13508));
  jand g13250(.dina(n13508), .dinb(n13507), .dout(n13509));
  jnot g13251(.din(n13509), .dout(n13510));
  jor  g13252(.dina(n5096), .dinb(n3227), .dout(n13511));
  jor  g13253(.dina(n4904), .dinb(n3035), .dout(n13512));
  jor  g13254(.dina(n5099), .dinb(n3055), .dout(n13513));
  jor  g13255(.dina(n5101), .dinb(n3230), .dout(n13514));
  jand g13256(.dina(n13514), .dinb(n13513), .dout(n13515));
  jand g13257(.dina(n13515), .dinb(n13512), .dout(n13516));
  jand g13258(.dina(n13516), .dinb(n13511), .dout(n13517));
  jxor g13259(.dina(n13517), .dinb(a41 ), .dout(n13518));
  jor  g13260(.dina(n6490), .dinb(n2404), .dout(n13519));
  jor  g13261(.dina(n6262), .dinb(n2010), .dout(n13520));
  jor  g13262(.dina(n6493), .dinb(n2148), .dout(n13521));
  jor  g13263(.dina(n6495), .dinb(n2407), .dout(n13522));
  jand g13264(.dina(n13522), .dinb(n13521), .dout(n13523));
  jand g13265(.dina(n13523), .dinb(n13520), .dout(n13524));
  jand g13266(.dina(n13524), .dinb(n13519), .dout(n13525));
  jxor g13267(.dina(n13525), .dinb(a47 ), .dout(n13526));
  jnot g13268(.din(n13526), .dout(n13527));
  jand g13269(.dina(n13268), .dinb(n13261), .dout(n13528));
  jand g13270(.dina(n13269), .dinb(n13197), .dout(n13529));
  jor  g13271(.dina(n13529), .dinb(n13528), .dout(n13530));
  jor  g13272(.dina(n7266), .dinb(n1884), .dout(n13531));
  jor  g13273(.dina(n7021), .dinb(n1742), .dout(n13532));
  jor  g13274(.dina(n7269), .dinb(n1867), .dout(n13533));
  jor  g13275(.dina(n7271), .dinb(n1887), .dout(n13534));
  jand g13276(.dina(n13534), .dinb(n13533), .dout(n13535));
  jand g13277(.dina(n13535), .dinb(n13532), .dout(n13536));
  jand g13278(.dina(n13536), .dinb(n13531), .dout(n13537));
  jxor g13279(.dina(n13537), .dinb(a50 ), .dout(n13538));
  jnot g13280(.din(n13538), .dout(n13539));
  jand g13281(.dina(n13250), .dinb(n13243), .dout(n13540));
  jnot g13282(.din(n13540), .dout(n13541));
  jor  g13283(.dina(n13260), .dinb(n13252), .dout(n13542));
  jand g13284(.dina(n13542), .dinb(n13541), .dout(n13543));
  jnot g13285(.din(n13543), .dout(n13544));
  jand g13286(.dina(n13226), .dinb(n13215), .dout(n13545));
  jand g13287(.dina(n13227), .dinb(n13206), .dout(n13546));
  jor  g13288(.dina(n13546), .dinb(n13545), .dout(n13547));
  jor  g13289(.dina(n9891), .dinb(n936), .dout(n13548));
  jor  g13290(.dina(n9593), .dinb(n778), .dout(n13549));
  jor  g13291(.dina(n9894), .dinb(n858), .dout(n13550));
  jor  g13292(.dina(n9896), .dinb(n939), .dout(n13551));
  jand g13293(.dina(n13551), .dinb(n13550), .dout(n13552));
  jand g13294(.dina(n13552), .dinb(n13549), .dout(n13553));
  jand g13295(.dina(n13553), .dinb(n13548), .dout(n13554));
  jxor g13296(.dina(n13554), .dinb(a59 ), .dout(n13555));
  jnot g13297(.din(n13555), .dout(n13556));
  jor  g13298(.dina(n10806), .dinb(n755), .dout(n13557));
  jor  g13299(.dina(n10485), .dinb(n627), .dout(n13558));
  jor  g13300(.dina(n10809), .dinb(n647), .dout(n13559));
  jor  g13301(.dina(n10811), .dinb(n758), .dout(n13560));
  jand g13302(.dina(n13560), .dinb(n13559), .dout(n13561));
  jand g13303(.dina(n13561), .dinb(n13558), .dout(n13562));
  jand g13304(.dina(n13562), .dinb(n13557), .dout(n13563));
  jxor g13305(.dina(n13563), .dinb(a62 ), .dout(n13564));
  jnot g13306(.din(n13564), .dout(n13565));
  jand g13307(.dina(n13224), .dinb(n13006), .dout(n13566));
  jand g13308(.dina(n13225), .dinb(n13220), .dout(n13567));
  jor  g13309(.dina(n13567), .dinb(n13566), .dout(n13568));
  jxor g13310(.dina(n13223), .dinb(n483), .dout(n13569));
  jand g13311(.dina(n10801), .dinb(b9 ), .dout(n13570));
  jand g13312(.dina(n11107), .dinb(b8 ), .dout(n13571));
  jor  g13313(.dina(n13571), .dinb(n13570), .dout(n13572));
  jxor g13314(.dina(n13572), .dinb(n13569), .dout(n13573));
  jxor g13315(.dina(n13573), .dinb(n13568), .dout(n13574));
  jxor g13316(.dina(n13574), .dinb(n13565), .dout(n13575));
  jxor g13317(.dina(n13575), .dinb(n13556), .dout(n13576));
  jxor g13318(.dina(n13576), .dinb(n13547), .dout(n13577));
  jnot g13319(.din(n13577), .dout(n13578));
  jor  g13320(.dina(n8978), .dinb(n1287), .dout(n13579));
  jor  g13321(.dina(n8677), .dinb(n1022), .dout(n13580));
  jor  g13322(.dina(n8981), .dinb(n1193), .dout(n13581));
  jor  g13323(.dina(n8983), .dinb(n1290), .dout(n13582));
  jand g13324(.dina(n13582), .dinb(n13581), .dout(n13583));
  jand g13325(.dina(n13583), .dinb(n13580), .dout(n13584));
  jand g13326(.dina(n13584), .dinb(n13579), .dout(n13585));
  jxor g13327(.dina(n13585), .dinb(a56 ), .dout(n13586));
  jxor g13328(.dina(n13586), .dinb(n13578), .dout(n13587));
  jnot g13329(.din(n13228), .dout(n13588));
  jnot g13330(.din(n13232), .dout(n13589));
  jand g13331(.dina(n13589), .dinb(n13588), .dout(n13590));
  jnot g13332(.din(n13590), .dout(n13591));
  jand g13333(.dina(n13232), .dinb(n13228), .dout(n13592));
  jor  g13334(.dina(n13242), .dinb(n13592), .dout(n13593));
  jand g13335(.dina(n13593), .dinb(n13591), .dout(n13594));
  jxor g13336(.dina(n13594), .dinb(n13587), .dout(n13595));
  jnot g13337(.din(n13595), .dout(n13596));
  jor  g13338(.dina(n8125), .dinb(n1617), .dout(n13597));
  jor  g13339(.dina(n7846), .dinb(n1400), .dout(n13598));
  jor  g13340(.dina(n8128), .dinb(n1420), .dout(n13599));
  jor  g13341(.dina(n8130), .dinb(n1620), .dout(n13600));
  jand g13342(.dina(n13600), .dinb(n13599), .dout(n13601));
  jand g13343(.dina(n13601), .dinb(n13598), .dout(n13602));
  jand g13344(.dina(n13602), .dinb(n13597), .dout(n13603));
  jxor g13345(.dina(n13603), .dinb(a53 ), .dout(n13604));
  jxor g13346(.dina(n13604), .dinb(n13596), .dout(n13605));
  jxor g13347(.dina(n13605), .dinb(n13544), .dout(n13606));
  jxor g13348(.dina(n13606), .dinb(n13539), .dout(n13607));
  jxor g13349(.dina(n13607), .dinb(n13530), .dout(n13608));
  jxor g13350(.dina(n13608), .dinb(n13527), .dout(n13609));
  jor  g13351(.dina(n13276), .dinb(n13270), .dout(n13610));
  jand g13352(.dina(n13276), .dinb(n13270), .dout(n13611));
  jor  g13353(.dina(n13286), .dinb(n13611), .dout(n13612));
  jand g13354(.dina(n13612), .dinb(n13610), .dout(n13613));
  jxor g13355(.dina(n13613), .dinb(n13609), .dout(n13614));
  jnot g13356(.din(n13614), .dout(n13615));
  jor  g13357(.dina(n5739), .dinb(n2867), .dout(n13616));
  jor  g13358(.dina(n5574), .dinb(n2559), .dout(n13617));
  jor  g13359(.dina(n5742), .dinb(n2579), .dout(n13618));
  jor  g13360(.dina(n5744), .dinb(n2870), .dout(n13619));
  jand g13361(.dina(n13619), .dinb(n13618), .dout(n13620));
  jand g13362(.dina(n13620), .dinb(n13617), .dout(n13621));
  jand g13363(.dina(n13621), .dinb(n13616), .dout(n13622));
  jxor g13364(.dina(n13622), .dinb(a44 ), .dout(n13623));
  jxor g13365(.dina(n13623), .dinb(n13615), .dout(n13624));
  jnot g13366(.din(n13287), .dout(n13625));
  jnot g13367(.din(n13293), .dout(n13626));
  jand g13368(.dina(n13626), .dinb(n13625), .dout(n13627));
  jnot g13369(.din(n13627), .dout(n13628));
  jand g13370(.dina(n13293), .dinb(n13287), .dout(n13629));
  jor  g13371(.dina(n13303), .dinb(n13629), .dout(n13630));
  jand g13372(.dina(n13630), .dinb(n13628), .dout(n13631));
  jnot g13373(.din(n13631), .dout(n13632));
  jxor g13374(.dina(n13632), .dinb(n13624), .dout(n13633));
  jxor g13375(.dina(n13633), .dinb(n13518), .dout(n13634));
  jxor g13376(.dina(n13634), .dinb(n13510), .dout(n13635));
  jxor g13377(.dina(n13635), .dinb(n13505), .dout(n13636));
  jnot g13378(.din(n13636), .dout(n13637));
  jand g13379(.dina(n13327), .dinb(n13322), .dout(n13638));
  jnot g13380(.din(n13638), .dout(n13639));
  jnot g13381(.din(n13322), .dout(n13640));
  jand g13382(.dina(n13326), .dinb(n13640), .dout(n13641));
  jor  g13383(.dina(n13337), .dinb(n13641), .dout(n13642));
  jand g13384(.dina(n13642), .dinb(n13639), .dout(n13643));
  jxor g13385(.dina(n13643), .dinb(n13637), .dout(n13644));
  jnot g13386(.din(n13644), .dout(n13645));
  jor  g13387(.dina(n4534), .dinb(n3849), .dout(n13646));
  jor  g13388(.dina(n3689), .dinb(n4140), .dout(n13647));
  jor  g13389(.dina(n3852), .dinb(n4340), .dout(n13648));
  jor  g13390(.dina(n3854), .dinb(n4537), .dout(n13649));
  jand g13391(.dina(n13649), .dinb(n13648), .dout(n13650));
  jand g13392(.dina(n13650), .dinb(n13647), .dout(n13651));
  jand g13393(.dina(n13651), .dinb(n13646), .dout(n13652));
  jxor g13394(.dina(n13652), .dinb(a35 ), .dout(n13653));
  jxor g13395(.dina(n13653), .dinb(n13645), .dout(n13654));
  jxor g13396(.dina(n13654), .dinb(n13496), .dout(n13655));
  jand g13397(.dina(n13184), .dinb(n13180), .dout(n13656));
  jand g13398(.dina(n13349), .dinb(n13185), .dout(n13657));
  jor  g13399(.dina(n13657), .dinb(n13656), .dout(n13658));
  jnot g13400(.din(n13658), .dout(n13659));
  jor  g13401(.dina(n4991), .dinb(n3301), .dout(n13660));
  jor  g13402(.dina(n3136), .dinb(n4557), .dout(n13661));
  jor  g13403(.dina(n3304), .dinb(n4974), .dout(n13662));
  jor  g13404(.dina(n3306), .dinb(n4994), .dout(n13663));
  jand g13405(.dina(n13663), .dinb(n13662), .dout(n13664));
  jand g13406(.dina(n13664), .dinb(n13661), .dout(n13665));
  jand g13407(.dina(n13665), .dinb(n13660), .dout(n13666));
  jxor g13408(.dina(n13666), .dinb(a32 ), .dout(n13667));
  jxor g13409(.dina(n13667), .dinb(n13659), .dout(n13668));
  jxor g13410(.dina(n13668), .dinb(n13655), .dout(n13669));
  jxor g13411(.dina(n13669), .dinb(n13491), .dout(n13670));
  jxor g13412(.dina(n13670), .dinb(n13476), .dout(n13671));
  jnot g13413(.din(n13671), .dout(n13672));
  jxor g13414(.dina(n13672), .dinb(n13463), .dout(n13673));
  jnot g13415(.din(n13673), .dout(n13674));
  jor  g13416(.dina(n13379), .dinb(n13371), .dout(n13675));
  jand g13417(.dina(n13380), .dinb(n13367), .dout(n13676));
  jnot g13418(.din(n13676), .dout(n13677));
  jand g13419(.dina(n13677), .dinb(n13675), .dout(n13678));
  jor  g13420(.dina(n7957), .dinb(n1566), .dout(n13679));
  jor  g13421(.dina(n1489), .dinb(n7411), .dout(n13680));
  jor  g13422(.dina(n1569), .dinb(n7683), .dout(n13681));
  jor  g13423(.dina(n1571), .dinb(n7960), .dout(n13682));
  jand g13424(.dina(n13682), .dinb(n13681), .dout(n13683));
  jand g13425(.dina(n13683), .dinb(n13680), .dout(n13684));
  jand g13426(.dina(n13684), .dinb(n13679), .dout(n13685));
  jxor g13427(.dina(n13685), .dinb(a20 ), .dout(n13686));
  jxor g13428(.dina(n13686), .dinb(n13678), .dout(n13687));
  jxor g13429(.dina(n13687), .dinb(n13674), .dout(n13688));
  jxor g13430(.dina(n13688), .dinb(n13450), .dout(n13689));
  jor  g13431(.dina(n13395), .dinb(n13391), .dout(n13690));
  jnot g13432(.din(n13396), .dout(n13691));
  jor  g13433(.dina(n13691), .dinb(n13383), .dout(n13692));
  jand g13434(.dina(n13692), .dinb(n13690), .dout(n13693));
  jor  g13435(.dina(n9722), .dinb(n974), .dout(n13694));
  jor  g13436(.dina(n908), .dinb(n9390), .dout(n13695));
  jor  g13437(.dina(n977), .dinb(n9413), .dout(n13696));
  jor  g13438(.dina(n979), .dinb(n9725), .dout(n13697));
  jand g13439(.dina(n13697), .dinb(n13696), .dout(n13698));
  jand g13440(.dina(n13698), .dinb(n13695), .dout(n13699));
  jand g13441(.dina(n13699), .dinb(n13694), .dout(n13700));
  jxor g13442(.dina(n13700), .dinb(a14 ), .dout(n13701));
  jxor g13443(.dina(n13701), .dinb(n13693), .dout(n13702));
  jxor g13444(.dina(n13702), .dinb(n13689), .dout(n13703));
  jor  g13445(.dina(n13410), .dinb(n13402), .dout(n13704));
  jor  g13446(.dina(n13412), .dinb(n13397), .dout(n13705));
  jand g13447(.dina(n13705), .dinb(n13704), .dout(n13706));
  jor  g13448(.dina(n10961), .dinb(n706), .dout(n13707));
  jor  g13449(.dina(n683), .dinb(n10314), .dout(n13708));
  jor  g13450(.dina(n709), .dinb(n10637), .dout(n13709));
  jor  g13451(.dina(n711), .dinb(n10964), .dout(n13710));
  jand g13452(.dina(n13710), .dinb(n13709), .dout(n13711));
  jand g13453(.dina(n13711), .dinb(n13708), .dout(n13712));
  jand g13454(.dina(n13712), .dinb(n13707), .dout(n13713));
  jxor g13455(.dina(n13713), .dinb(a11 ), .dout(n13714));
  jxor g13456(.dina(n13714), .dinb(n13706), .dout(n13715));
  jxor g13457(.dina(n13715), .dinb(n13703), .dout(n13716));
  jxor g13458(.dina(n13716), .dinb(n13437), .dout(n13717));
  jxor g13459(.dina(n13717), .dinb(n13433), .dout(f72 ));
  jand g13460(.dina(n13716), .dinb(n13437), .dout(n13719));
  jand g13461(.dina(n13717), .dinb(n13433), .dout(n13720));
  jor  g13462(.dina(n13720), .dinb(n13719), .dout(n13721));
  jor  g13463(.dina(n13714), .dinb(n13706), .dout(n13722));
  jnot g13464(.din(n13722), .dout(n13723));
  jand g13465(.dina(n13715), .dinb(n13703), .dout(n13724));
  jor  g13466(.dina(n13724), .dinb(n13723), .dout(n13725));
  jor  g13467(.dina(n10311), .dinb(n974), .dout(n13726));
  jor  g13468(.dina(n908), .dinb(n9413), .dout(n13727));
  jor  g13469(.dina(n977), .dinb(n9725), .dout(n13728));
  jor  g13470(.dina(n979), .dinb(n10314), .dout(n13729));
  jand g13471(.dina(n13729), .dinb(n13728), .dout(n13730));
  jand g13472(.dina(n13730), .dinb(n13727), .dout(n13731));
  jand g13473(.dina(n13731), .dinb(n13726), .dout(n13732));
  jxor g13474(.dina(n13732), .dinb(a14 ), .dout(n13733));
  jnot g13475(.din(n13733), .dout(n13734));
  jnot g13476(.din(n13445), .dout(n13735));
  jnot g13477(.din(n13449), .dout(n13736));
  jand g13478(.dina(n13736), .dinb(n13735), .dout(n13737));
  jand g13479(.dina(n13688), .dinb(n13450), .dout(n13738));
  jor  g13480(.dina(n13738), .dinb(n13737), .dout(n13739));
  jxor g13481(.dina(n13739), .dinb(n13734), .dout(n13740));
  jor  g13482(.dina(n8228), .dinb(n1566), .dout(n13741));
  jor  g13483(.dina(n1489), .dinb(n7683), .dout(n13742));
  jor  g13484(.dina(n1569), .dinb(n7960), .dout(n13743));
  jor  g13485(.dina(n1571), .dinb(n8231), .dout(n13744));
  jand g13486(.dina(n13744), .dinb(n13743), .dout(n13745));
  jand g13487(.dina(n13745), .dinb(n13742), .dout(n13746));
  jand g13488(.dina(n13746), .dinb(n13741), .dout(n13747));
  jxor g13489(.dina(n13747), .dinb(a20 ), .dout(n13748));
  jnot g13490(.din(n13748), .dout(n13749));
  jand g13491(.dina(n13462), .dinb(n13458), .dout(n13750));
  jnot g13492(.din(n13750), .dout(n13751));
  jnot g13493(.din(n13458), .dout(n13752));
  jnot g13494(.din(n13462), .dout(n13753));
  jand g13495(.dina(n13753), .dinb(n13752), .dout(n13754));
  jor  g13496(.dina(n13671), .dinb(n13754), .dout(n13755));
  jand g13497(.dina(n13755), .dinb(n13751), .dout(n13756));
  jxor g13498(.dina(n13756), .dinb(n13749), .dout(n13757));
  jor  g13499(.dina(n7408), .dinb(n1939), .dout(n13758));
  jor  g13500(.dina(n1827), .dinb(n7129), .dout(n13759));
  jor  g13501(.dina(n1942), .dinb(n7149), .dout(n13760));
  jor  g13502(.dina(n1944), .dinb(n7411), .dout(n13761));
  jand g13503(.dina(n13761), .dinb(n13760), .dout(n13762));
  jand g13504(.dina(n13762), .dinb(n13759), .dout(n13763));
  jand g13505(.dina(n13763), .dinb(n13758), .dout(n13764));
  jxor g13506(.dina(n13764), .dinb(a23 ), .dout(n13765));
  jnot g13507(.din(n13765), .dout(n13766));
  jand g13508(.dina(n13475), .dinb(n13472), .dout(n13767));
  jand g13509(.dina(n13670), .dinb(n13476), .dout(n13768));
  jor  g13510(.dina(n13768), .dinb(n13767), .dout(n13769));
  jxor g13511(.dina(n13769), .dinb(n13766), .dout(n13770));
  jor  g13512(.dina(n13667), .dinb(n13659), .dout(n13771));
  jand g13513(.dina(n13668), .dinb(n13655), .dout(n13772));
  jnot g13514(.din(n13772), .dout(n13773));
  jand g13515(.dina(n13773), .dinb(n13771), .dout(n13774));
  jor  g13516(.dina(n6103), .dinb(n2784), .dout(n13775));
  jor  g13517(.dina(n2661), .dinb(n5428), .dout(n13776));
  jor  g13518(.dina(n2787), .dinb(n5862), .dout(n13777));
  jor  g13519(.dina(n2789), .dinb(n6106), .dout(n13778));
  jand g13520(.dina(n13778), .dinb(n13777), .dout(n13779));
  jand g13521(.dina(n13779), .dinb(n13776), .dout(n13780));
  jand g13522(.dina(n13780), .dinb(n13775), .dout(n13781));
  jxor g13523(.dina(n13781), .dinb(a29 ), .dout(n13782));
  jxor g13524(.dina(n13782), .dinb(n13774), .dout(n13783));
  jor  g13525(.dina(n5405), .dinb(n3301), .dout(n13784));
  jor  g13526(.dina(n3136), .dinb(n4974), .dout(n13785));
  jor  g13527(.dina(n3304), .dinb(n4994), .dout(n13786));
  jor  g13528(.dina(n3306), .dinb(n5408), .dout(n13787));
  jand g13529(.dina(n13787), .dinb(n13786), .dout(n13788));
  jand g13530(.dina(n13788), .dinb(n13785), .dout(n13789));
  jand g13531(.dina(n13789), .dinb(n13784), .dout(n13790));
  jxor g13532(.dina(n13790), .dinb(a32 ), .dout(n13791));
  jor  g13533(.dina(n13653), .dinb(n13645), .dout(n13792));
  jand g13534(.dina(n13654), .dinb(n13496), .dout(n13793));
  jnot g13535(.din(n13793), .dout(n13794));
  jand g13536(.dina(n13794), .dinb(n13792), .dout(n13795));
  jxor g13537(.dina(n13795), .dinb(n13791), .dout(n13796));
  jor  g13538(.dina(n4554), .dinb(n3849), .dout(n13797));
  jor  g13539(.dina(n3689), .dinb(n4340), .dout(n13798));
  jor  g13540(.dina(n3852), .dinb(n4537), .dout(n13799));
  jor  g13541(.dina(n3854), .dinb(n4557), .dout(n13800));
  jand g13542(.dina(n13800), .dinb(n13799), .dout(n13801));
  jand g13543(.dina(n13801), .dinb(n13798), .dout(n13802));
  jand g13544(.dina(n13802), .dinb(n13797), .dout(n13803));
  jxor g13545(.dina(n13803), .dinb(a35 ), .dout(n13804));
  jnot g13546(.din(n13804), .dout(n13805));
  jand g13547(.dina(n13635), .dinb(n13505), .dout(n13806));
  jnot g13548(.din(n13806), .dout(n13807));
  jor  g13549(.dina(n13643), .dinb(n13637), .dout(n13808));
  jand g13550(.dina(n13808), .dinb(n13807), .dout(n13809));
  jnot g13551(.din(n13809), .dout(n13810));
  jor  g13552(.dina(n4137), .dinb(n4415), .dout(n13811));
  jor  g13553(.dina(n4272), .dinb(n3588), .dout(n13812));
  jor  g13554(.dina(n4418), .dinb(n3942), .dout(n13813));
  jor  g13555(.dina(n4420), .dinb(n4140), .dout(n13814));
  jand g13556(.dina(n13814), .dinb(n13813), .dout(n13815));
  jand g13557(.dina(n13815), .dinb(n13812), .dout(n13816));
  jand g13558(.dina(n13816), .dinb(n13811), .dout(n13817));
  jxor g13559(.dina(n13817), .dinb(a38 ), .dout(n13818));
  jnot g13560(.din(n13818), .dout(n13819));
  jor  g13561(.dina(n13633), .dinb(n13518), .dout(n13820));
  jand g13562(.dina(n13634), .dinb(n13510), .dout(n13821));
  jnot g13563(.din(n13821), .dout(n13822));
  jand g13564(.dina(n13822), .dinb(n13820), .dout(n13823));
  jnot g13565(.din(n13823), .dout(n13824));
  jor  g13566(.dina(n5096), .dinb(n3400), .dout(n13825));
  jor  g13567(.dina(n4904), .dinb(n3055), .dout(n13826));
  jor  g13568(.dina(n5099), .dinb(n3230), .dout(n13827));
  jor  g13569(.dina(n5101), .dinb(n3403), .dout(n13828));
  jand g13570(.dina(n13828), .dinb(n13827), .dout(n13829));
  jand g13571(.dina(n13829), .dinb(n13826), .dout(n13830));
  jand g13572(.dina(n13830), .dinb(n13825), .dout(n13831));
  jxor g13573(.dina(n13831), .dinb(a41 ), .dout(n13832));
  jnot g13574(.din(n13832), .dout(n13833));
  jand g13575(.dina(n13608), .dinb(n13527), .dout(n13834));
  jand g13576(.dina(n13613), .dinb(n13609), .dout(n13835));
  jor  g13577(.dina(n13835), .dinb(n13834), .dout(n13836));
  jand g13578(.dina(n13606), .dinb(n13539), .dout(n13837));
  jand g13579(.dina(n13607), .dinb(n13530), .dout(n13838));
  jor  g13580(.dina(n13838), .dinb(n13837), .dout(n13839));
  jor  g13581(.dina(n13604), .dinb(n13596), .dout(n13840));
  jand g13582(.dina(n13605), .dinb(n13544), .dout(n13841));
  jnot g13583(.din(n13841), .dout(n13842));
  jand g13584(.dina(n13842), .dinb(n13840), .dout(n13843));
  jnot g13585(.din(n13843), .dout(n13844));
  jor  g13586(.dina(n13586), .dinb(n13578), .dout(n13845));
  jand g13587(.dina(n13594), .dinb(n13587), .dout(n13846));
  jnot g13588(.din(n13846), .dout(n13847));
  jand g13589(.dina(n13847), .dinb(n13845), .dout(n13848));
  jnot g13590(.din(n13848), .dout(n13849));
  jand g13591(.dina(n13575), .dinb(n13556), .dout(n13850));
  jand g13592(.dina(n13576), .dinb(n13547), .dout(n13851));
  jor  g13593(.dina(n13851), .dinb(n13850), .dout(n13852));
  jor  g13594(.dina(n9891), .dinb(n1019), .dout(n13853));
  jor  g13595(.dina(n9593), .dinb(n858), .dout(n13854));
  jor  g13596(.dina(n9894), .dinb(n939), .dout(n13855));
  jor  g13597(.dina(n9896), .dinb(n1022), .dout(n13856));
  jand g13598(.dina(n13856), .dinb(n13855), .dout(n13857));
  jand g13599(.dina(n13857), .dinb(n13854), .dout(n13858));
  jand g13600(.dina(n13858), .dinb(n13853), .dout(n13859));
  jxor g13601(.dina(n13859), .dinb(a59 ), .dout(n13860));
  jnot g13602(.din(n13860), .dout(n13861));
  jand g13603(.dina(n13573), .dinb(n13568), .dout(n13862));
  jand g13604(.dina(n13574), .dinb(n13565), .dout(n13863));
  jor  g13605(.dina(n13863), .dinb(n13862), .dout(n13864));
  jor  g13606(.dina(n10806), .dinb(n775), .dout(n13865));
  jor  g13607(.dina(n10485), .dinb(n647), .dout(n13866));
  jor  g13608(.dina(n10809), .dinb(n758), .dout(n13867));
  jor  g13609(.dina(n10811), .dinb(n778), .dout(n13868));
  jand g13610(.dina(n13868), .dinb(n13867), .dout(n13869));
  jand g13611(.dina(n13869), .dinb(n13866), .dout(n13870));
  jand g13612(.dina(n13870), .dinb(n13865), .dout(n13871));
  jxor g13613(.dina(n13871), .dinb(a62 ), .dout(n13872));
  jand g13614(.dina(n13223), .dinb(n483), .dout(n13873));
  jand g13615(.dina(n13572), .dinb(n13569), .dout(n13874));
  jor  g13616(.dina(n13874), .dinb(n13873), .dout(n13875));
  jand g13617(.dina(n10801), .dinb(b10 ), .dout(n13876));
  jand g13618(.dina(n11107), .dinb(b9 ), .dout(n13877));
  jor  g13619(.dina(n13877), .dinb(n13876), .dout(n13878));
  jxor g13620(.dina(n13878), .dinb(n13875), .dout(n13879));
  jxor g13621(.dina(n13879), .dinb(n13872), .dout(n13880));
  jxor g13622(.dina(n13880), .dinb(n13864), .dout(n13881));
  jxor g13623(.dina(n13881), .dinb(n13861), .dout(n13882));
  jxor g13624(.dina(n13882), .dinb(n13852), .dout(n13883));
  jor  g13625(.dina(n8978), .dinb(n1397), .dout(n13884));
  jor  g13626(.dina(n8677), .dinb(n1193), .dout(n13885));
  jor  g13627(.dina(n8981), .dinb(n1290), .dout(n13886));
  jor  g13628(.dina(n8983), .dinb(n1400), .dout(n13887));
  jand g13629(.dina(n13887), .dinb(n13886), .dout(n13888));
  jand g13630(.dina(n13888), .dinb(n13885), .dout(n13889));
  jand g13631(.dina(n13889), .dinb(n13884), .dout(n13890));
  jxor g13632(.dina(n13890), .dinb(a56 ), .dout(n13891));
  jnot g13633(.din(n13891), .dout(n13892));
  jxor g13634(.dina(n13892), .dinb(n13883), .dout(n13893));
  jxor g13635(.dina(n13893), .dinb(n13849), .dout(n13894));
  jor  g13636(.dina(n8125), .dinb(n1739), .dout(n13895));
  jor  g13637(.dina(n7846), .dinb(n1420), .dout(n13896));
  jor  g13638(.dina(n8128), .dinb(n1620), .dout(n13897));
  jor  g13639(.dina(n8130), .dinb(n1742), .dout(n13898));
  jand g13640(.dina(n13898), .dinb(n13897), .dout(n13899));
  jand g13641(.dina(n13899), .dinb(n13896), .dout(n13900));
  jand g13642(.dina(n13900), .dinb(n13895), .dout(n13901));
  jxor g13643(.dina(n13901), .dinb(a53 ), .dout(n13902));
  jnot g13644(.din(n13902), .dout(n13903));
  jxor g13645(.dina(n13903), .dinb(n13894), .dout(n13904));
  jxor g13646(.dina(n13904), .dinb(n13844), .dout(n13905));
  jor  g13647(.dina(n7266), .dinb(n2007), .dout(n13906));
  jor  g13648(.dina(n7021), .dinb(n1867), .dout(n13907));
  jor  g13649(.dina(n7269), .dinb(n1887), .dout(n13908));
  jor  g13650(.dina(n7271), .dinb(n2010), .dout(n13909));
  jand g13651(.dina(n13909), .dinb(n13908), .dout(n13910));
  jand g13652(.dina(n13910), .dinb(n13907), .dout(n13911));
  jand g13653(.dina(n13911), .dinb(n13906), .dout(n13912));
  jxor g13654(.dina(n13912), .dinb(a50 ), .dout(n13913));
  jnot g13655(.din(n13913), .dout(n13914));
  jxor g13656(.dina(n13914), .dinb(n13905), .dout(n13915));
  jxor g13657(.dina(n13915), .dinb(n13839), .dout(n13916));
  jor  g13658(.dina(n6490), .dinb(n2556), .dout(n13917));
  jor  g13659(.dina(n6262), .dinb(n2148), .dout(n13918));
  jor  g13660(.dina(n6493), .dinb(n2407), .dout(n13919));
  jor  g13661(.dina(n6495), .dinb(n2559), .dout(n13920));
  jand g13662(.dina(n13920), .dinb(n13919), .dout(n13921));
  jand g13663(.dina(n13921), .dinb(n13918), .dout(n13922));
  jand g13664(.dina(n13922), .dinb(n13917), .dout(n13923));
  jxor g13665(.dina(n13923), .dinb(a47 ), .dout(n13924));
  jnot g13666(.din(n13924), .dout(n13925));
  jxor g13667(.dina(n13925), .dinb(n13916), .dout(n13926));
  jxor g13668(.dina(n13926), .dinb(n13836), .dout(n13927));
  jnot g13669(.din(n13927), .dout(n13928));
  jor  g13670(.dina(n5739), .dinb(n3032), .dout(n13929));
  jor  g13671(.dina(n5574), .dinb(n2579), .dout(n13930));
  jor  g13672(.dina(n5742), .dinb(n2870), .dout(n13931));
  jor  g13673(.dina(n5744), .dinb(n3035), .dout(n13932));
  jand g13674(.dina(n13932), .dinb(n13931), .dout(n13933));
  jand g13675(.dina(n13933), .dinb(n13930), .dout(n13934));
  jand g13676(.dina(n13934), .dinb(n13929), .dout(n13935));
  jxor g13677(.dina(n13935), .dinb(a44 ), .dout(n13936));
  jxor g13678(.dina(n13936), .dinb(n13928), .dout(n13937));
  jand g13679(.dina(n13623), .dinb(n13615), .dout(n13938));
  jnot g13680(.din(n13938), .dout(n13939));
  jnot g13681(.din(n13623), .dout(n13940));
  jand g13682(.dina(n13940), .dinb(n13614), .dout(n13941));
  jor  g13683(.dina(n13631), .dinb(n13941), .dout(n13942));
  jand g13684(.dina(n13942), .dinb(n13939), .dout(n13943));
  jxor g13685(.dina(n13943), .dinb(n13937), .dout(n13944));
  jxor g13686(.dina(n13944), .dinb(n13833), .dout(n13945));
  jxor g13687(.dina(n13945), .dinb(n13824), .dout(n13946));
  jxor g13688(.dina(n13946), .dinb(n13819), .dout(n13947));
  jxor g13689(.dina(n13947), .dinb(n13810), .dout(n13948));
  jxor g13690(.dina(n13948), .dinb(n13805), .dout(n13949));
  jxor g13691(.dina(n13949), .dinb(n13796), .dout(n13950));
  jxor g13692(.dina(n13950), .dinb(n13783), .dout(n13951));
  jor  g13693(.dina(n6864), .dinb(n2319), .dout(n13952));
  jor  g13694(.dina(n2224), .dinb(n6352), .dout(n13953));
  jor  g13695(.dina(n2322), .dinb(n6372), .dout(n13954));
  jor  g13696(.dina(n2324), .dinb(n6867), .dout(n13955));
  jand g13697(.dina(n13955), .dinb(n13954), .dout(n13956));
  jand g13698(.dina(n13956), .dinb(n13953), .dout(n13957));
  jand g13699(.dina(n13957), .dinb(n13952), .dout(n13958));
  jxor g13700(.dina(n13958), .dinb(a26 ), .dout(n13959));
  jor  g13701(.dina(n13490), .dinb(n13482), .dout(n13960));
  jand g13702(.dina(n13669), .dinb(n13491), .dout(n13961));
  jnot g13703(.din(n13961), .dout(n13962));
  jand g13704(.dina(n13962), .dinb(n13960), .dout(n13963));
  jxor g13705(.dina(n13963), .dinb(n13959), .dout(n13964));
  jxor g13706(.dina(n13964), .dinb(n13951), .dout(n13965));
  jxor g13707(.dina(n13965), .dinb(n13770), .dout(n13966));
  jxor g13708(.dina(n13966), .dinb(n13757), .dout(n13967));
  jor  g13709(.dina(n13686), .dinb(n13678), .dout(n13968));
  jand g13710(.dina(n13687), .dinb(n13674), .dout(n13969));
  jnot g13711(.din(n13969), .dout(n13970));
  jand g13712(.dina(n13970), .dinb(n13968), .dout(n13971));
  jor  g13713(.dina(n9387), .dinb(n1245), .dout(n13972));
  jor  g13714(.dina(n1165), .dinb(n8789), .dout(n13973));
  jor  g13715(.dina(n1248), .dinb(n8809), .dout(n13974));
  jor  g13716(.dina(n1250), .dinb(n9390), .dout(n13975));
  jand g13717(.dina(n13975), .dinb(n13974), .dout(n13976));
  jand g13718(.dina(n13976), .dinb(n13973), .dout(n13977));
  jand g13719(.dina(n13977), .dinb(n13972), .dout(n13978));
  jxor g13720(.dina(n13978), .dinb(a17 ), .dout(n13979));
  jxor g13721(.dina(n13979), .dinb(n13971), .dout(n13980));
  jxor g13722(.dina(n13980), .dinb(n13967), .dout(n13981));
  jxor g13723(.dina(n13981), .dinb(n13740), .dout(n13982));
  jor  g13724(.dina(n13701), .dinb(n13693), .dout(n13983));
  jnot g13725(.din(n13689), .dout(n13984));
  jnot g13726(.din(n13702), .dout(n13985));
  jor  g13727(.dina(n13985), .dinb(n13984), .dout(n13986));
  jand g13728(.dina(n13986), .dinb(n13983), .dout(n13987));
  jor  g13729(.dina(n10978), .dinb(n706), .dout(n13988));
  jor  g13730(.dina(n683), .dinb(n10637), .dout(n13989));
  jor  g13731(.dina(n709), .dinb(n10964), .dout(n13990));
  jand g13732(.dina(n13990), .dinb(n13989), .dout(n13991));
  jand g13733(.dina(n13991), .dinb(n13988), .dout(n13992));
  jxor g13734(.dina(n13992), .dinb(a11 ), .dout(n13993));
  jxor g13735(.dina(n13993), .dinb(n13987), .dout(n13994));
  jxor g13736(.dina(n13994), .dinb(n13982), .dout(n13995));
  jxor g13737(.dina(n13995), .dinb(n13725), .dout(n13996));
  jxor g13738(.dina(n13996), .dinb(n13721), .dout(f73 ));
  jand g13739(.dina(n13995), .dinb(n13725), .dout(n13998));
  jand g13740(.dina(n13996), .dinb(n13721), .dout(n13999));
  jor  g13741(.dina(n13999), .dinb(n13998), .dout(n14000));
  jor  g13742(.dina(n13993), .dinb(n13987), .dout(n14001));
  jnot g13743(.din(n14001), .dout(n14002));
  jand g13744(.dina(n13994), .dinb(n13982), .dout(n14003));
  jor  g13745(.dina(n14003), .dinb(n14002), .dout(n14004));
  jor  g13746(.dina(n13979), .dinb(n13971), .dout(n14005));
  jand g13747(.dina(n13980), .dinb(n13967), .dout(n14006));
  jnot g13748(.din(n14006), .dout(n14007));
  jand g13749(.dina(n14007), .dinb(n14005), .dout(n14008));
  jor  g13750(.dina(n10634), .dinb(n974), .dout(n14009));
  jor  g13751(.dina(n908), .dinb(n9725), .dout(n14010));
  jor  g13752(.dina(n977), .dinb(n10314), .dout(n14011));
  jor  g13753(.dina(n979), .dinb(n10637), .dout(n14012));
  jand g13754(.dina(n14012), .dinb(n14011), .dout(n14013));
  jand g13755(.dina(n14013), .dinb(n14010), .dout(n14014));
  jand g13756(.dina(n14014), .dinb(n14009), .dout(n14015));
  jxor g13757(.dina(n14015), .dinb(a14 ), .dout(n14016));
  jxor g13758(.dina(n14016), .dinb(n14008), .dout(n14017));
  jor  g13759(.dina(n9410), .dinb(n1245), .dout(n14018));
  jor  g13760(.dina(n1165), .dinb(n8809), .dout(n14019));
  jor  g13761(.dina(n1248), .dinb(n9390), .dout(n14020));
  jor  g13762(.dina(n1250), .dinb(n9413), .dout(n14021));
  jand g13763(.dina(n14021), .dinb(n14020), .dout(n14022));
  jand g13764(.dina(n14022), .dinb(n14019), .dout(n14023));
  jand g13765(.dina(n14023), .dinb(n14018), .dout(n14024));
  jxor g13766(.dina(n14024), .dinb(a17 ), .dout(n14025));
  jnot g13767(.din(n14025), .dout(n14026));
  jand g13768(.dina(n13756), .dinb(n13749), .dout(n14027));
  jand g13769(.dina(n13966), .dinb(n13757), .dout(n14028));
  jor  g13770(.dina(n14028), .dinb(n14027), .dout(n14029));
  jxor g13771(.dina(n14029), .dinb(n14026), .dout(n14030));
  jor  g13772(.dina(n8786), .dinb(n1566), .dout(n14031));
  jor  g13773(.dina(n1489), .dinb(n7960), .dout(n14032));
  jor  g13774(.dina(n1569), .dinb(n8231), .dout(n14033));
  jor  g13775(.dina(n1571), .dinb(n8789), .dout(n14034));
  jand g13776(.dina(n14034), .dinb(n14033), .dout(n14035));
  jand g13777(.dina(n14035), .dinb(n14032), .dout(n14036));
  jand g13778(.dina(n14036), .dinb(n14031), .dout(n14037));
  jxor g13779(.dina(n14037), .dinb(a20 ), .dout(n14038));
  jnot g13780(.din(n14038), .dout(n14039));
  jand g13781(.dina(n13769), .dinb(n13766), .dout(n14040));
  jand g13782(.dina(n13965), .dinb(n13770), .dout(n14041));
  jor  g13783(.dina(n14041), .dinb(n14040), .dout(n14042));
  jxor g13784(.dina(n14042), .dinb(n14039), .dout(n14043));
  jor  g13785(.dina(n13782), .dinb(n13774), .dout(n14044));
  jand g13786(.dina(n13950), .dinb(n13783), .dout(n14045));
  jnot g13787(.din(n14045), .dout(n14046));
  jand g13788(.dina(n14046), .dinb(n14044), .dout(n14047));
  jor  g13789(.dina(n7126), .dinb(n2319), .dout(n14048));
  jor  g13790(.dina(n2224), .dinb(n6372), .dout(n14049));
  jor  g13791(.dina(n2322), .dinb(n6867), .dout(n14050));
  jor  g13792(.dina(n2324), .dinb(n7129), .dout(n14051));
  jand g13793(.dina(n14051), .dinb(n14050), .dout(n14052));
  jand g13794(.dina(n14052), .dinb(n14049), .dout(n14053));
  jand g13795(.dina(n14053), .dinb(n14048), .dout(n14054));
  jxor g13796(.dina(n14054), .dinb(a26 ), .dout(n14055));
  jxor g13797(.dina(n14055), .dinb(n14047), .dout(n14056));
  jor  g13798(.dina(n6349), .dinb(n2784), .dout(n14057));
  jor  g13799(.dina(n2661), .dinb(n5862), .dout(n14058));
  jor  g13800(.dina(n2787), .dinb(n6106), .dout(n14059));
  jor  g13801(.dina(n2789), .dinb(n6352), .dout(n14060));
  jand g13802(.dina(n14060), .dinb(n14059), .dout(n14061));
  jand g13803(.dina(n14061), .dinb(n14058), .dout(n14062));
  jand g13804(.dina(n14062), .dinb(n14057), .dout(n14063));
  jxor g13805(.dina(n14063), .dinb(a29 ), .dout(n14064));
  jand g13806(.dina(n13795), .dinb(n13791), .dout(n14065));
  jor  g13807(.dina(n13795), .dinb(n13791), .dout(n14066));
  jnot g13808(.din(n13949), .dout(n14067));
  jand g13809(.dina(n14067), .dinb(n14066), .dout(n14068));
  jor  g13810(.dina(n14068), .dinb(n14065), .dout(n14069));
  jxor g13811(.dina(n14069), .dinb(n14064), .dout(n14070));
  jor  g13812(.dina(n5425), .dinb(n3301), .dout(n14071));
  jor  g13813(.dina(n3136), .dinb(n4994), .dout(n14072));
  jor  g13814(.dina(n3304), .dinb(n5408), .dout(n14073));
  jor  g13815(.dina(n3306), .dinb(n5428), .dout(n14074));
  jand g13816(.dina(n14074), .dinb(n14073), .dout(n14075));
  jand g13817(.dina(n14075), .dinb(n14072), .dout(n14076));
  jand g13818(.dina(n14076), .dinb(n14071), .dout(n14077));
  jxor g13819(.dina(n14077), .dinb(a32 ), .dout(n14078));
  jnot g13820(.din(n14078), .dout(n14079));
  jor  g13821(.dina(n13947), .dinb(n13810), .dout(n14080));
  jand g13822(.dina(n13947), .dinb(n13810), .dout(n14081));
  jor  g13823(.dina(n14081), .dinb(n13805), .dout(n14082));
  jand g13824(.dina(n14082), .dinb(n14080), .dout(n14083));
  jxor g13825(.dina(n14083), .dinb(n14079), .dout(n14084));
  jor  g13826(.dina(n4971), .dinb(n3849), .dout(n14085));
  jor  g13827(.dina(n3689), .dinb(n4537), .dout(n14086));
  jor  g13828(.dina(n3852), .dinb(n4557), .dout(n14087));
  jor  g13829(.dina(n3854), .dinb(n4974), .dout(n14088));
  jand g13830(.dina(n14088), .dinb(n14087), .dout(n14089));
  jand g13831(.dina(n14089), .dinb(n14086), .dout(n14090));
  jand g13832(.dina(n14090), .dinb(n14085), .dout(n14091));
  jxor g13833(.dina(n14091), .dinb(a35 ), .dout(n14092));
  jnot g13834(.din(n14092), .dout(n14093));
  jand g13835(.dina(n13945), .dinb(n13824), .dout(n14094));
  jand g13836(.dina(n13946), .dinb(n13819), .dout(n14095));
  jor  g13837(.dina(n14095), .dinb(n14094), .dout(n14096));
  jand g13838(.dina(n13943), .dinb(n13937), .dout(n14097));
  jand g13839(.dina(n13944), .dinb(n13833), .dout(n14098));
  jor  g13840(.dina(n14098), .dinb(n14097), .dout(n14099));
  jor  g13841(.dina(n7266), .dinb(n2145), .dout(n14100));
  jor  g13842(.dina(n7021), .dinb(n1887), .dout(n14101));
  jor  g13843(.dina(n7269), .dinb(n2010), .dout(n14102));
  jor  g13844(.dina(n7271), .dinb(n2148), .dout(n14103));
  jand g13845(.dina(n14103), .dinb(n14102), .dout(n14104));
  jand g13846(.dina(n14104), .dinb(n14101), .dout(n14105));
  jand g13847(.dina(n14105), .dinb(n14100), .dout(n14106));
  jxor g13848(.dina(n14106), .dinb(a50 ), .dout(n14107));
  jnot g13849(.din(n14107), .dout(n14108));
  jor  g13850(.dina(n8125), .dinb(n1864), .dout(n14109));
  jor  g13851(.dina(n7846), .dinb(n1620), .dout(n14110));
  jor  g13852(.dina(n8128), .dinb(n1742), .dout(n14111));
  jor  g13853(.dina(n8130), .dinb(n1867), .dout(n14112));
  jand g13854(.dina(n14112), .dinb(n14111), .dout(n14113));
  jand g13855(.dina(n14113), .dinb(n14110), .dout(n14114));
  jand g13856(.dina(n14114), .dinb(n14109), .dout(n14115));
  jxor g13857(.dina(n14115), .dinb(a53 ), .dout(n14116));
  jnot g13858(.din(n14116), .dout(n14117));
  jor  g13859(.dina(n9891), .dinb(n1190), .dout(n14118));
  jor  g13860(.dina(n9593), .dinb(n939), .dout(n14119));
  jor  g13861(.dina(n9894), .dinb(n1022), .dout(n14120));
  jor  g13862(.dina(n9896), .dinb(n1193), .dout(n14121));
  jand g13863(.dina(n14121), .dinb(n14120), .dout(n14122));
  jand g13864(.dina(n14122), .dinb(n14119), .dout(n14123));
  jand g13865(.dina(n14123), .dinb(n14118), .dout(n14124));
  jxor g13866(.dina(n14124), .dinb(a59 ), .dout(n14125));
  jor  g13867(.dina(n10806), .dinb(n855), .dout(n14126));
  jor  g13868(.dina(n10485), .dinb(n758), .dout(n14127));
  jor  g13869(.dina(n10809), .dinb(n778), .dout(n14128));
  jor  g13870(.dina(n10811), .dinb(n858), .dout(n14129));
  jand g13871(.dina(n14129), .dinb(n14128), .dout(n14130));
  jand g13872(.dina(n14130), .dinb(n14127), .dout(n14131));
  jand g13873(.dina(n14131), .dinb(n14126), .dout(n14132));
  jxor g13874(.dina(n14132), .dinb(a62 ), .dout(n14133));
  jnot g13875(.din(n13878), .dout(n14134));
  jand g13876(.dina(n10801), .dinb(b11 ), .dout(n14135));
  jand g13877(.dina(n11107), .dinb(b10 ), .dout(n14136));
  jor  g13878(.dina(n14136), .dinb(n14135), .dout(n14137));
  jxor g13879(.dina(n14137), .dinb(n14134), .dout(n14138));
  jor  g13880(.dina(n14134), .dinb(n13875), .dout(n14139));
  jnot g13881(.din(n13872), .dout(n14140));
  jand g13882(.dina(n14134), .dinb(n13875), .dout(n14141));
  jor  g13883(.dina(n14141), .dinb(n14140), .dout(n14142));
  jand g13884(.dina(n14142), .dinb(n14139), .dout(n14143));
  jxor g13885(.dina(n14143), .dinb(n14138), .dout(n14144));
  jxor g13886(.dina(n14144), .dinb(n14133), .dout(n14145));
  jxor g13887(.dina(n14145), .dinb(n14125), .dout(n14146));
  jor  g13888(.dina(n13880), .dinb(n13864), .dout(n14147));
  jand g13889(.dina(n13880), .dinb(n13864), .dout(n14148));
  jor  g13890(.dina(n14148), .dinb(n13861), .dout(n14149));
  jand g13891(.dina(n14149), .dinb(n14147), .dout(n14150));
  jxor g13892(.dina(n14150), .dinb(n14146), .dout(n14151));
  jnot g13893(.din(n14151), .dout(n14152));
  jor  g13894(.dina(n8978), .dinb(n1417), .dout(n14153));
  jor  g13895(.dina(n8677), .dinb(n1290), .dout(n14154));
  jor  g13896(.dina(n8981), .dinb(n1400), .dout(n14155));
  jor  g13897(.dina(n8983), .dinb(n1420), .dout(n14156));
  jand g13898(.dina(n14156), .dinb(n14155), .dout(n14157));
  jand g13899(.dina(n14157), .dinb(n14154), .dout(n14158));
  jand g13900(.dina(n14158), .dinb(n14153), .dout(n14159));
  jxor g13901(.dina(n14159), .dinb(a56 ), .dout(n14160));
  jxor g13902(.dina(n14160), .dinb(n14152), .dout(n14161));
  jnot g13903(.din(n13852), .dout(n14162));
  jnot g13904(.din(n13882), .dout(n14163));
  jand g13905(.dina(n14163), .dinb(n14162), .dout(n14164));
  jnot g13906(.din(n14164), .dout(n14165));
  jand g13907(.dina(n13882), .dinb(n13852), .dout(n14166));
  jor  g13908(.dina(n13892), .dinb(n14166), .dout(n14167));
  jand g13909(.dina(n14167), .dinb(n14165), .dout(n14168));
  jxor g13910(.dina(n14168), .dinb(n14161), .dout(n14169));
  jxor g13911(.dina(n14169), .dinb(n14117), .dout(n14170));
  jnot g13912(.din(n13893), .dout(n14171));
  jand g13913(.dina(n14171), .dinb(n13848), .dout(n14172));
  jnot g13914(.din(n14172), .dout(n14173));
  jand g13915(.dina(n13893), .dinb(n13849), .dout(n14174));
  jor  g13916(.dina(n13903), .dinb(n14174), .dout(n14175));
  jand g13917(.dina(n14175), .dinb(n14173), .dout(n14176));
  jxor g13918(.dina(n14176), .dinb(n14170), .dout(n14177));
  jxor g13919(.dina(n14177), .dinb(n14108), .dout(n14178));
  jnot g13920(.din(n13904), .dout(n14179));
  jand g13921(.dina(n14179), .dinb(n13843), .dout(n14180));
  jnot g13922(.din(n14180), .dout(n14181));
  jand g13923(.dina(n13904), .dinb(n13844), .dout(n14182));
  jor  g13924(.dina(n13914), .dinb(n14182), .dout(n14183));
  jand g13925(.dina(n14183), .dinb(n14181), .dout(n14184));
  jxor g13926(.dina(n14184), .dinb(n14178), .dout(n14185));
  jor  g13927(.dina(n6490), .dinb(n2576), .dout(n14186));
  jor  g13928(.dina(n6262), .dinb(n2407), .dout(n14187));
  jor  g13929(.dina(n6493), .dinb(n2559), .dout(n14188));
  jor  g13930(.dina(n6495), .dinb(n2579), .dout(n14189));
  jand g13931(.dina(n14189), .dinb(n14188), .dout(n14190));
  jand g13932(.dina(n14190), .dinb(n14187), .dout(n14191));
  jand g13933(.dina(n14191), .dinb(n14186), .dout(n14192));
  jxor g13934(.dina(n14192), .dinb(a47 ), .dout(n14193));
  jnot g13935(.din(n14193), .dout(n14194));
  jxor g13936(.dina(n14194), .dinb(n14185), .dout(n14195));
  jnot g13937(.din(n13839), .dout(n14196));
  jnot g13938(.din(n13915), .dout(n14197));
  jand g13939(.dina(n14197), .dinb(n14196), .dout(n14198));
  jnot g13940(.din(n14198), .dout(n14199));
  jand g13941(.dina(n13915), .dinb(n13839), .dout(n14200));
  jor  g13942(.dina(n13925), .dinb(n14200), .dout(n14201));
  jand g13943(.dina(n14201), .dinb(n14199), .dout(n14202));
  jxor g13944(.dina(n14202), .dinb(n14195), .dout(n14203));
  jnot g13945(.din(n14203), .dout(n14204));
  jor  g13946(.dina(n5739), .dinb(n3052), .dout(n14205));
  jor  g13947(.dina(n5574), .dinb(n2870), .dout(n14206));
  jor  g13948(.dina(n5742), .dinb(n3035), .dout(n14207));
  jor  g13949(.dina(n5744), .dinb(n3055), .dout(n14208));
  jand g13950(.dina(n14208), .dinb(n14207), .dout(n14209));
  jand g13951(.dina(n14209), .dinb(n14206), .dout(n14210));
  jand g13952(.dina(n14210), .dinb(n14205), .dout(n14211));
  jxor g13953(.dina(n14211), .dinb(a44 ), .dout(n14212));
  jxor g13954(.dina(n14212), .dinb(n14204), .dout(n14213));
  jand g13955(.dina(n13926), .dinb(n13836), .dout(n14214));
  jnot g13956(.din(n14214), .dout(n14215));
  jor  g13957(.dina(n13936), .dinb(n13928), .dout(n14216));
  jand g13958(.dina(n14216), .dinb(n14215), .dout(n14217));
  jnot g13959(.din(n14217), .dout(n14218));
  jxor g13960(.dina(n14218), .dinb(n14213), .dout(n14219));
  jnot g13961(.din(n14219), .dout(n14220));
  jor  g13962(.dina(n5096), .dinb(n3585), .dout(n14221));
  jor  g13963(.dina(n4904), .dinb(n3230), .dout(n14222));
  jor  g13964(.dina(n5099), .dinb(n3403), .dout(n14223));
  jor  g13965(.dina(n5101), .dinb(n3588), .dout(n14224));
  jand g13966(.dina(n14224), .dinb(n14223), .dout(n14225));
  jand g13967(.dina(n14225), .dinb(n14222), .dout(n14226));
  jand g13968(.dina(n14226), .dinb(n14221), .dout(n14227));
  jxor g13969(.dina(n14227), .dinb(a41 ), .dout(n14228));
  jxor g13970(.dina(n14228), .dinb(n14220), .dout(n14229));
  jxor g13971(.dina(n14229), .dinb(n14099), .dout(n14230));
  jnot g13972(.din(n14230), .dout(n14231));
  jor  g13973(.dina(n4337), .dinb(n4415), .dout(n14232));
  jor  g13974(.dina(n4272), .dinb(n3942), .dout(n14233));
  jor  g13975(.dina(n4418), .dinb(n4140), .dout(n14234));
  jor  g13976(.dina(n4420), .dinb(n4340), .dout(n14235));
  jand g13977(.dina(n14235), .dinb(n14234), .dout(n14236));
  jand g13978(.dina(n14236), .dinb(n14233), .dout(n14237));
  jand g13979(.dina(n14237), .dinb(n14232), .dout(n14238));
  jxor g13980(.dina(n14238), .dinb(a38 ), .dout(n14239));
  jxor g13981(.dina(n14239), .dinb(n14231), .dout(n14240));
  jxor g13982(.dina(n14240), .dinb(n14096), .dout(n14241));
  jxor g13983(.dina(n14241), .dinb(n14093), .dout(n14242));
  jxor g13984(.dina(n14242), .dinb(n14084), .dout(n14243));
  jxor g13985(.dina(n14243), .dinb(n14070), .dout(n14244));
  jxor g13986(.dina(n14244), .dinb(n14056), .dout(n14245));
  jor  g13987(.dina(n13963), .dinb(n13959), .dout(n14246));
  jand g13988(.dina(n13964), .dinb(n13951), .dout(n14247));
  jnot g13989(.din(n14247), .dout(n14248));
  jand g13990(.dina(n14248), .dinb(n14246), .dout(n14249));
  jor  g13991(.dina(n7680), .dinb(n1939), .dout(n14250));
  jor  g13992(.dina(n1827), .dinb(n7149), .dout(n14251));
  jor  g13993(.dina(n1942), .dinb(n7411), .dout(n14252));
  jor  g13994(.dina(n1944), .dinb(n7683), .dout(n14253));
  jand g13995(.dina(n14253), .dinb(n14252), .dout(n14254));
  jand g13996(.dina(n14254), .dinb(n14251), .dout(n14255));
  jand g13997(.dina(n14255), .dinb(n14250), .dout(n14256));
  jxor g13998(.dina(n14256), .dinb(a23 ), .dout(n14257));
  jxor g13999(.dina(n14257), .dinb(n14249), .dout(n14258));
  jxor g14000(.dina(n14258), .dinb(n14245), .dout(n14259));
  jxor g14001(.dina(n14259), .dinb(n14043), .dout(n14260));
  jxor g14002(.dina(n14260), .dinb(n14030), .dout(n14261));
  jxor g14003(.dina(n14261), .dinb(n14017), .dout(n14262));
  jand g14004(.dina(n13739), .dinb(n13734), .dout(n14263));
  jand g14005(.dina(n13981), .dinb(n13740), .dout(n14264));
  jor  g14006(.dina(n14264), .dinb(n14263), .dout(n14265));
  jnot g14007(.din(n14265), .dout(n14266));
  jand g14008(.dina(n11296), .dinb(n601), .dout(n14267));
  jor  g14009(.dina(n14267), .dinb(n684), .dout(n14268));
  jand g14010(.dina(n14268), .dinb(b63 ), .dout(n14269));
  jxor g14011(.dina(n14269), .dinb(n678), .dout(n14270));
  jxor g14012(.dina(n14270), .dinb(n14266), .dout(n14271));
  jxor g14013(.dina(n14271), .dinb(n14262), .dout(n14272));
  jxor g14014(.dina(n14272), .dinb(n14004), .dout(n14273));
  jxor g14015(.dina(n14273), .dinb(n14000), .dout(f74 ));
  jand g14016(.dina(n14272), .dinb(n14004), .dout(n14275));
  jand g14017(.dina(n14273), .dinb(n14000), .dout(n14276));
  jor  g14018(.dina(n14276), .dinb(n14275), .dout(n14277));
  jor  g14019(.dina(n14270), .dinb(n14266), .dout(n14278));
  jand g14020(.dina(n14271), .dinb(n14262), .dout(n14279));
  jnot g14021(.din(n14279), .dout(n14280));
  jand g14022(.dina(n14280), .dinb(n14278), .dout(n14281));
  jnot g14023(.din(n14281), .dout(n14282));
  jor  g14024(.dina(n8806), .dinb(n1566), .dout(n14283));
  jor  g14025(.dina(n1489), .dinb(n8231), .dout(n14284));
  jor  g14026(.dina(n1569), .dinb(n8789), .dout(n14285));
  jor  g14027(.dina(n1571), .dinb(n8809), .dout(n14286));
  jand g14028(.dina(n14286), .dinb(n14285), .dout(n14287));
  jand g14029(.dina(n14287), .dinb(n14284), .dout(n14288));
  jand g14030(.dina(n14288), .dinb(n14283), .dout(n14289));
  jxor g14031(.dina(n14289), .dinb(a20 ), .dout(n14290));
  jnot g14032(.din(n14290), .dout(n14291));
  jand g14033(.dina(n14042), .dinb(n14039), .dout(n14292));
  jand g14034(.dina(n14259), .dinb(n14043), .dout(n14293));
  jor  g14035(.dina(n14293), .dinb(n14292), .dout(n14294));
  jxor g14036(.dina(n14294), .dinb(n14291), .dout(n14295));
  jor  g14037(.dina(n7146), .dinb(n2319), .dout(n14296));
  jor  g14038(.dina(n2224), .dinb(n6867), .dout(n14297));
  jor  g14039(.dina(n2322), .dinb(n7129), .dout(n14298));
  jor  g14040(.dina(n2324), .dinb(n7149), .dout(n14299));
  jand g14041(.dina(n14299), .dinb(n14298), .dout(n14300));
  jand g14042(.dina(n14300), .dinb(n14297), .dout(n14301));
  jand g14043(.dina(n14301), .dinb(n14296), .dout(n14302));
  jxor g14044(.dina(n14302), .dinb(a26 ), .dout(n14303));
  jor  g14045(.dina(n14055), .dinb(n14047), .dout(n14304));
  jand g14046(.dina(n14244), .dinb(n14056), .dout(n14305));
  jnot g14047(.din(n14305), .dout(n14306));
  jand g14048(.dina(n14306), .dinb(n14304), .dout(n14307));
  jxor g14049(.dina(n14307), .dinb(n14303), .dout(n14308));
  jor  g14050(.dina(n4991), .dinb(n3849), .dout(n14309));
  jor  g14051(.dina(n3689), .dinb(n4557), .dout(n14310));
  jor  g14052(.dina(n3852), .dinb(n4974), .dout(n14311));
  jor  g14053(.dina(n3854), .dinb(n4994), .dout(n14312));
  jand g14054(.dina(n14312), .dinb(n14311), .dout(n14313));
  jand g14055(.dina(n14313), .dinb(n14310), .dout(n14314));
  jand g14056(.dina(n14314), .dinb(n14309), .dout(n14315));
  jxor g14057(.dina(n14315), .dinb(a35 ), .dout(n14316));
  jnot g14058(.din(n14316), .dout(n14317));
  jand g14059(.dina(n14229), .dinb(n14099), .dout(n14318));
  jnot g14060(.din(n14318), .dout(n14319));
  jor  g14061(.dina(n14239), .dinb(n14231), .dout(n14320));
  jand g14062(.dina(n14320), .dinb(n14319), .dout(n14321));
  jnot g14063(.din(n14321), .dout(n14322));
  jor  g14064(.dina(n5096), .dinb(n3939), .dout(n14323));
  jor  g14065(.dina(n4904), .dinb(n3403), .dout(n14324));
  jor  g14066(.dina(n5099), .dinb(n3588), .dout(n14325));
  jor  g14067(.dina(n5101), .dinb(n3942), .dout(n14326));
  jand g14068(.dina(n14326), .dinb(n14325), .dout(n14327));
  jand g14069(.dina(n14327), .dinb(n14324), .dout(n14328));
  jand g14070(.dina(n14328), .dinb(n14323), .dout(n14329));
  jxor g14071(.dina(n14329), .dinb(a41 ), .dout(n14330));
  jnot g14072(.din(n14330), .dout(n14331));
  jand g14073(.dina(n14202), .dinb(n14195), .dout(n14332));
  jnot g14074(.din(n14332), .dout(n14333));
  jor  g14075(.dina(n14212), .dinb(n14204), .dout(n14334));
  jand g14076(.dina(n14334), .dinb(n14333), .dout(n14335));
  jnot g14077(.din(n14335), .dout(n14336));
  jor  g14078(.dina(n5739), .dinb(n3227), .dout(n14337));
  jor  g14079(.dina(n5574), .dinb(n3035), .dout(n14338));
  jor  g14080(.dina(n5742), .dinb(n3055), .dout(n14339));
  jor  g14081(.dina(n5744), .dinb(n3230), .dout(n14340));
  jand g14082(.dina(n14340), .dinb(n14339), .dout(n14341));
  jand g14083(.dina(n14341), .dinb(n14338), .dout(n14342));
  jand g14084(.dina(n14342), .dinb(n14337), .dout(n14343));
  jxor g14085(.dina(n14343), .dinb(a44 ), .dout(n14344));
  jand g14086(.dina(n14176), .dinb(n14170), .dout(n14345));
  jand g14087(.dina(n14177), .dinb(n14108), .dout(n14346));
  jor  g14088(.dina(n14346), .dinb(n14345), .dout(n14347));
  jor  g14089(.dina(n7266), .dinb(n2404), .dout(n14348));
  jor  g14090(.dina(n7021), .dinb(n2010), .dout(n14349));
  jor  g14091(.dina(n7269), .dinb(n2148), .dout(n14350));
  jor  g14092(.dina(n7271), .dinb(n2407), .dout(n14351));
  jand g14093(.dina(n14351), .dinb(n14350), .dout(n14352));
  jand g14094(.dina(n14352), .dinb(n14349), .dout(n14353));
  jand g14095(.dina(n14353), .dinb(n14348), .dout(n14354));
  jxor g14096(.dina(n14354), .dinb(a50 ), .dout(n14355));
  jnot g14097(.din(n14355), .dout(n14356));
  jand g14098(.dina(n14168), .dinb(n14161), .dout(n14357));
  jand g14099(.dina(n14169), .dinb(n14117), .dout(n14358));
  jor  g14100(.dina(n14358), .dinb(n14357), .dout(n14359));
  jor  g14101(.dina(n8125), .dinb(n1884), .dout(n14360));
  jor  g14102(.dina(n7846), .dinb(n1742), .dout(n14361));
  jor  g14103(.dina(n8128), .dinb(n1867), .dout(n14362));
  jor  g14104(.dina(n8130), .dinb(n1887), .dout(n14363));
  jand g14105(.dina(n14363), .dinb(n14362), .dout(n14364));
  jand g14106(.dina(n14364), .dinb(n14361), .dout(n14365));
  jand g14107(.dina(n14365), .dinb(n14360), .dout(n14366));
  jxor g14108(.dina(n14366), .dinb(a53 ), .dout(n14367));
  jnot g14109(.din(n14367), .dout(n14368));
  jand g14110(.dina(n14150), .dinb(n14146), .dout(n14369));
  jnot g14111(.din(n14369), .dout(n14370));
  jor  g14112(.dina(n14160), .dinb(n14152), .dout(n14371));
  jand g14113(.dina(n14371), .dinb(n14370), .dout(n14372));
  jnot g14114(.din(n14372), .dout(n14373));
  jor  g14115(.dina(n9891), .dinb(n1287), .dout(n14374));
  jor  g14116(.dina(n9593), .dinb(n1022), .dout(n14375));
  jor  g14117(.dina(n9894), .dinb(n1193), .dout(n14376));
  jor  g14118(.dina(n9896), .dinb(n1290), .dout(n14377));
  jand g14119(.dina(n14377), .dinb(n14376), .dout(n14378));
  jand g14120(.dina(n14378), .dinb(n14375), .dout(n14379));
  jand g14121(.dina(n14379), .dinb(n14374), .dout(n14380));
  jxor g14122(.dina(n14380), .dinb(a59 ), .dout(n14381));
  jnot g14123(.din(n14381), .dout(n14382));
  jand g14124(.dina(n14137), .dinb(n14134), .dout(n14383));
  jand g14125(.dina(n14143), .dinb(n14138), .dout(n14384));
  jor  g14126(.dina(n14384), .dinb(n14383), .dout(n14385));
  jor  g14127(.dina(n10806), .dinb(n936), .dout(n14386));
  jor  g14128(.dina(n10485), .dinb(n778), .dout(n14387));
  jor  g14129(.dina(n10809), .dinb(n858), .dout(n14388));
  jor  g14130(.dina(n10811), .dinb(n939), .dout(n14389));
  jand g14131(.dina(n14389), .dinb(n14388), .dout(n14390));
  jand g14132(.dina(n14390), .dinb(n14387), .dout(n14391));
  jand g14133(.dina(n14391), .dinb(n14386), .dout(n14392));
  jxor g14134(.dina(n14392), .dinb(a62 ), .dout(n14393));
  jnot g14135(.din(n14393), .dout(n14394));
  jxor g14136(.dina(n13878), .dinb(n678), .dout(n14395));
  jand g14137(.dina(n10801), .dinb(b12 ), .dout(n14396));
  jand g14138(.dina(n11107), .dinb(b11 ), .dout(n14397));
  jor  g14139(.dina(n14397), .dinb(n14396), .dout(n14398));
  jxor g14140(.dina(n14398), .dinb(n14395), .dout(n14399));
  jxor g14141(.dina(n14399), .dinb(n14394), .dout(n14400));
  jxor g14142(.dina(n14400), .dinb(n14385), .dout(n14401));
  jxor g14143(.dina(n14401), .dinb(n14382), .dout(n14402));
  jnot g14144(.din(n14133), .dout(n14403));
  jor  g14145(.dina(n14144), .dinb(n14403), .dout(n14404));
  jnot g14146(.din(n14125), .dout(n14405));
  jand g14147(.dina(n14144), .dinb(n14403), .dout(n14406));
  jor  g14148(.dina(n14406), .dinb(n14405), .dout(n14407));
  jand g14149(.dina(n14407), .dinb(n14404), .dout(n14408));
  jxor g14150(.dina(n14408), .dinb(n14402), .dout(n14409));
  jnot g14151(.din(n14409), .dout(n14410));
  jor  g14152(.dina(n8978), .dinb(n1617), .dout(n14411));
  jor  g14153(.dina(n8677), .dinb(n1400), .dout(n14412));
  jor  g14154(.dina(n8981), .dinb(n1420), .dout(n14413));
  jor  g14155(.dina(n8983), .dinb(n1620), .dout(n14414));
  jand g14156(.dina(n14414), .dinb(n14413), .dout(n14415));
  jand g14157(.dina(n14415), .dinb(n14412), .dout(n14416));
  jand g14158(.dina(n14416), .dinb(n14411), .dout(n14417));
  jxor g14159(.dina(n14417), .dinb(a56 ), .dout(n14418));
  jxor g14160(.dina(n14418), .dinb(n14410), .dout(n14419));
  jxor g14161(.dina(n14419), .dinb(n14373), .dout(n14420));
  jxor g14162(.dina(n14420), .dinb(n14368), .dout(n14421));
  jxor g14163(.dina(n14421), .dinb(n14359), .dout(n14422));
  jxor g14164(.dina(n14422), .dinb(n14356), .dout(n14423));
  jxor g14165(.dina(n14423), .dinb(n14347), .dout(n14424));
  jnot g14166(.din(n14424), .dout(n14425));
  jor  g14167(.dina(n6490), .dinb(n2867), .dout(n14426));
  jor  g14168(.dina(n6262), .dinb(n2559), .dout(n14427));
  jor  g14169(.dina(n6493), .dinb(n2579), .dout(n14428));
  jor  g14170(.dina(n6495), .dinb(n2870), .dout(n14429));
  jand g14171(.dina(n14429), .dinb(n14428), .dout(n14430));
  jand g14172(.dina(n14430), .dinb(n14427), .dout(n14431));
  jand g14173(.dina(n14431), .dinb(n14426), .dout(n14432));
  jxor g14174(.dina(n14432), .dinb(a47 ), .dout(n14433));
  jxor g14175(.dina(n14433), .dinb(n14425), .dout(n14434));
  jor  g14176(.dina(n14184), .dinb(n14178), .dout(n14435));
  jand g14177(.dina(n14184), .dinb(n14178), .dout(n14436));
  jor  g14178(.dina(n14194), .dinb(n14436), .dout(n14437));
  jand g14179(.dina(n14437), .dinb(n14435), .dout(n14438));
  jnot g14180(.din(n14438), .dout(n14439));
  jxor g14181(.dina(n14439), .dinb(n14434), .dout(n14440));
  jxor g14182(.dina(n14440), .dinb(n14344), .dout(n14441));
  jxor g14183(.dina(n14441), .dinb(n14336), .dout(n14442));
  jxor g14184(.dina(n14442), .dinb(n14331), .dout(n14443));
  jnot g14185(.din(n14443), .dout(n14444));
  jand g14186(.dina(n14218), .dinb(n14213), .dout(n14445));
  jnot g14187(.din(n14445), .dout(n14446));
  jnot g14188(.din(n14213), .dout(n14447));
  jand g14189(.dina(n14217), .dinb(n14447), .dout(n14448));
  jor  g14190(.dina(n14228), .dinb(n14448), .dout(n14449));
  jand g14191(.dina(n14449), .dinb(n14446), .dout(n14450));
  jxor g14192(.dina(n14450), .dinb(n14444), .dout(n14451));
  jnot g14193(.din(n14451), .dout(n14452));
  jor  g14194(.dina(n4534), .dinb(n4415), .dout(n14453));
  jor  g14195(.dina(n4272), .dinb(n4140), .dout(n14454));
  jor  g14196(.dina(n4418), .dinb(n4340), .dout(n14455));
  jor  g14197(.dina(n4420), .dinb(n4537), .dout(n14456));
  jand g14198(.dina(n14456), .dinb(n14455), .dout(n14457));
  jand g14199(.dina(n14457), .dinb(n14454), .dout(n14458));
  jand g14200(.dina(n14458), .dinb(n14453), .dout(n14459));
  jxor g14201(.dina(n14459), .dinb(a38 ), .dout(n14460));
  jxor g14202(.dina(n14460), .dinb(n14452), .dout(n14461));
  jxor g14203(.dina(n14461), .dinb(n14322), .dout(n14462));
  jxor g14204(.dina(n14462), .dinb(n14317), .dout(n14463));
  jor  g14205(.dina(n14240), .dinb(n14096), .dout(n14464));
  jand g14206(.dina(n14240), .dinb(n14096), .dout(n14465));
  jor  g14207(.dina(n14465), .dinb(n14093), .dout(n14466));
  jand g14208(.dina(n14466), .dinb(n14464), .dout(n14467));
  jxor g14209(.dina(n14467), .dinb(n14463), .dout(n14468));
  jor  g14210(.dina(n5859), .dinb(n3301), .dout(n14469));
  jor  g14211(.dina(n3136), .dinb(n5408), .dout(n14470));
  jor  g14212(.dina(n3304), .dinb(n5428), .dout(n14471));
  jor  g14213(.dina(n3306), .dinb(n5862), .dout(n14472));
  jand g14214(.dina(n14472), .dinb(n14471), .dout(n14473));
  jand g14215(.dina(n14473), .dinb(n14470), .dout(n14474));
  jand g14216(.dina(n14474), .dinb(n14469), .dout(n14475));
  jxor g14217(.dina(n14475), .dinb(a32 ), .dout(n14476));
  jnot g14218(.din(n14476), .dout(n14477));
  jor  g14219(.dina(n14083), .dinb(n14079), .dout(n14478));
  jand g14220(.dina(n14083), .dinb(n14079), .dout(n14479));
  jor  g14221(.dina(n14242), .dinb(n14479), .dout(n14480));
  jand g14222(.dina(n14480), .dinb(n14478), .dout(n14481));
  jxor g14223(.dina(n14481), .dinb(n14477), .dout(n14482));
  jxor g14224(.dina(n14482), .dinb(n14468), .dout(n14483));
  jnot g14225(.din(n14064), .dout(n14484));
  jnot g14226(.din(n14069), .dout(n14485));
  jand g14227(.dina(n14485), .dinb(n14484), .dout(n14486));
  jand g14228(.dina(n14243), .dinb(n14070), .dout(n14487));
  jor  g14229(.dina(n14487), .dinb(n14486), .dout(n14488));
  jnot g14230(.din(n14488), .dout(n14489));
  jor  g14231(.dina(n6369), .dinb(n2784), .dout(n14490));
  jor  g14232(.dina(n2661), .dinb(n6106), .dout(n14491));
  jor  g14233(.dina(n2787), .dinb(n6352), .dout(n14492));
  jor  g14234(.dina(n2789), .dinb(n6372), .dout(n14493));
  jand g14235(.dina(n14493), .dinb(n14492), .dout(n14494));
  jand g14236(.dina(n14494), .dinb(n14491), .dout(n14495));
  jand g14237(.dina(n14495), .dinb(n14490), .dout(n14496));
  jxor g14238(.dina(n14496), .dinb(a29 ), .dout(n14497));
  jxor g14239(.dina(n14497), .dinb(n14489), .dout(n14498));
  jxor g14240(.dina(n14498), .dinb(n14483), .dout(n14499));
  jxor g14241(.dina(n14499), .dinb(n14308), .dout(n14500));
  jor  g14242(.dina(n14257), .dinb(n14249), .dout(n14501));
  jand g14243(.dina(n14258), .dinb(n14245), .dout(n14502));
  jnot g14244(.din(n14502), .dout(n14503));
  jand g14245(.dina(n14503), .dinb(n14501), .dout(n14504));
  jor  g14246(.dina(n7957), .dinb(n1939), .dout(n14505));
  jor  g14247(.dina(n1827), .dinb(n7411), .dout(n14506));
  jor  g14248(.dina(n1942), .dinb(n7683), .dout(n14507));
  jor  g14249(.dina(n1944), .dinb(n7960), .dout(n14508));
  jand g14250(.dina(n14508), .dinb(n14507), .dout(n14509));
  jand g14251(.dina(n14509), .dinb(n14506), .dout(n14510));
  jand g14252(.dina(n14510), .dinb(n14505), .dout(n14511));
  jxor g14253(.dina(n14511), .dinb(a23 ), .dout(n14512));
  jxor g14254(.dina(n14512), .dinb(n14504), .dout(n14513));
  jxor g14255(.dina(n14513), .dinb(n14500), .dout(n14514));
  jxor g14256(.dina(n14514), .dinb(n14295), .dout(n14515));
  jand g14257(.dina(n14029), .dinb(n14026), .dout(n14516));
  jand g14258(.dina(n14260), .dinb(n14030), .dout(n14517));
  jor  g14259(.dina(n14517), .dinb(n14516), .dout(n14518));
  jnot g14260(.din(n14518), .dout(n14519));
  jor  g14261(.dina(n9722), .dinb(n1245), .dout(n14520));
  jor  g14262(.dina(n1165), .dinb(n9390), .dout(n14521));
  jor  g14263(.dina(n1248), .dinb(n9413), .dout(n14522));
  jor  g14264(.dina(n1250), .dinb(n9725), .dout(n14523));
  jand g14265(.dina(n14523), .dinb(n14522), .dout(n14524));
  jand g14266(.dina(n14524), .dinb(n14521), .dout(n14525));
  jand g14267(.dina(n14525), .dinb(n14520), .dout(n14526));
  jxor g14268(.dina(n14526), .dinb(a17 ), .dout(n14527));
  jxor g14269(.dina(n14527), .dinb(n14519), .dout(n14528));
  jxor g14270(.dina(n14528), .dinb(n14515), .dout(n14529));
  jor  g14271(.dina(n14016), .dinb(n14008), .dout(n14530));
  jand g14272(.dina(n14261), .dinb(n14017), .dout(n14531));
  jnot g14273(.din(n14531), .dout(n14532));
  jand g14274(.dina(n14532), .dinb(n14530), .dout(n14533));
  jor  g14275(.dina(n10961), .dinb(n974), .dout(n14534));
  jor  g14276(.dina(n908), .dinb(n10314), .dout(n14535));
  jor  g14277(.dina(n977), .dinb(n10637), .dout(n14536));
  jor  g14278(.dina(n979), .dinb(n10964), .dout(n14537));
  jand g14279(.dina(n14537), .dinb(n14536), .dout(n14538));
  jand g14280(.dina(n14538), .dinb(n14535), .dout(n14539));
  jand g14281(.dina(n14539), .dinb(n14534), .dout(n14540));
  jxor g14282(.dina(n14540), .dinb(a14 ), .dout(n14541));
  jxor g14283(.dina(n14541), .dinb(n14533), .dout(n14542));
  jxor g14284(.dina(n14542), .dinb(n14529), .dout(n14543));
  jxor g14285(.dina(n14543), .dinb(n14282), .dout(n14544));
  jxor g14286(.dina(n14544), .dinb(n14277), .dout(f75 ));
  jand g14287(.dina(n14543), .dinb(n14282), .dout(n14546));
  jand g14288(.dina(n14544), .dinb(n14277), .dout(n14547));
  jor  g14289(.dina(n14547), .dinb(n14546), .dout(n14548));
  jor  g14290(.dina(n14541), .dinb(n14533), .dout(n14549));
  jand g14291(.dina(n14542), .dinb(n14529), .dout(n14550));
  jnot g14292(.din(n14550), .dout(n14551));
  jand g14293(.dina(n14551), .dinb(n14549), .dout(n14552));
  jnot g14294(.din(n14552), .dout(n14553));
  jor  g14295(.dina(n10311), .dinb(n1245), .dout(n14554));
  jor  g14296(.dina(n1165), .dinb(n9413), .dout(n14555));
  jor  g14297(.dina(n1248), .dinb(n9725), .dout(n14556));
  jor  g14298(.dina(n1250), .dinb(n10314), .dout(n14557));
  jand g14299(.dina(n14557), .dinb(n14556), .dout(n14558));
  jand g14300(.dina(n14558), .dinb(n14555), .dout(n14559));
  jand g14301(.dina(n14559), .dinb(n14554), .dout(n14560));
  jxor g14302(.dina(n14560), .dinb(a17 ), .dout(n14561));
  jnot g14303(.din(n14561), .dout(n14562));
  jand g14304(.dina(n14294), .dinb(n14291), .dout(n14563));
  jand g14305(.dina(n14514), .dinb(n14295), .dout(n14564));
  jor  g14306(.dina(n14564), .dinb(n14563), .dout(n14565));
  jxor g14307(.dina(n14565), .dinb(n14562), .dout(n14566));
  jor  g14308(.dina(n14497), .dinb(n14489), .dout(n14567));
  jand g14309(.dina(n14498), .dinb(n14483), .dout(n14568));
  jnot g14310(.din(n14568), .dout(n14569));
  jand g14311(.dina(n14569), .dinb(n14567), .dout(n14570));
  jor  g14312(.dina(n7408), .dinb(n2319), .dout(n14571));
  jor  g14313(.dina(n2224), .dinb(n7129), .dout(n14572));
  jor  g14314(.dina(n2322), .dinb(n7149), .dout(n14573));
  jor  g14315(.dina(n2324), .dinb(n7411), .dout(n14574));
  jand g14316(.dina(n14574), .dinb(n14573), .dout(n14575));
  jand g14317(.dina(n14575), .dinb(n14572), .dout(n14576));
  jand g14318(.dina(n14576), .dinb(n14571), .dout(n14577));
  jxor g14319(.dina(n14577), .dinb(a26 ), .dout(n14578));
  jxor g14320(.dina(n14578), .dinb(n14570), .dout(n14579));
  jand g14321(.dina(n14462), .dinb(n14317), .dout(n14580));
  jand g14322(.dina(n14467), .dinb(n14463), .dout(n14581));
  jor  g14323(.dina(n14581), .dinb(n14580), .dout(n14582));
  jnot g14324(.din(n14582), .dout(n14583));
  jor  g14325(.dina(n6103), .dinb(n3301), .dout(n14584));
  jor  g14326(.dina(n3136), .dinb(n5428), .dout(n14585));
  jor  g14327(.dina(n3304), .dinb(n5862), .dout(n14586));
  jor  g14328(.dina(n3306), .dinb(n6106), .dout(n14587));
  jand g14329(.dina(n14587), .dinb(n14586), .dout(n14588));
  jand g14330(.dina(n14588), .dinb(n14585), .dout(n14589));
  jand g14331(.dina(n14589), .dinb(n14584), .dout(n14590));
  jxor g14332(.dina(n14590), .dinb(a32 ), .dout(n14591));
  jxor g14333(.dina(n14591), .dinb(n14583), .dout(n14592));
  jor  g14334(.dina(n14460), .dinb(n14452), .dout(n14593));
  jand g14335(.dina(n14461), .dinb(n14322), .dout(n14594));
  jnot g14336(.din(n14594), .dout(n14595));
  jand g14337(.dina(n14595), .dinb(n14593), .dout(n14596));
  jnot g14338(.din(n14596), .dout(n14597));
  jor  g14339(.dina(n4554), .dinb(n4415), .dout(n14598));
  jor  g14340(.dina(n4272), .dinb(n4340), .dout(n14599));
  jor  g14341(.dina(n4418), .dinb(n4537), .dout(n14600));
  jor  g14342(.dina(n4420), .dinb(n4557), .dout(n14601));
  jand g14343(.dina(n14601), .dinb(n14600), .dout(n14602));
  jand g14344(.dina(n14602), .dinb(n14599), .dout(n14603));
  jand g14345(.dina(n14603), .dinb(n14598), .dout(n14604));
  jxor g14346(.dina(n14604), .dinb(a38 ), .dout(n14605));
  jnot g14347(.din(n14605), .dout(n14606));
  jand g14348(.dina(n14442), .dinb(n14331), .dout(n14607));
  jnot g14349(.din(n14607), .dout(n14608));
  jor  g14350(.dina(n14450), .dinb(n14444), .dout(n14609));
  jand g14351(.dina(n14609), .dinb(n14608), .dout(n14610));
  jnot g14352(.din(n14610), .dout(n14611));
  jor  g14353(.dina(n5096), .dinb(n4137), .dout(n14612));
  jor  g14354(.dina(n4904), .dinb(n3588), .dout(n14613));
  jor  g14355(.dina(n5099), .dinb(n3942), .dout(n14614));
  jor  g14356(.dina(n5101), .dinb(n4140), .dout(n14615));
  jand g14357(.dina(n14615), .dinb(n14614), .dout(n14616));
  jand g14358(.dina(n14616), .dinb(n14613), .dout(n14617));
  jand g14359(.dina(n14617), .dinb(n14612), .dout(n14618));
  jxor g14360(.dina(n14618), .dinb(a41 ), .dout(n14619));
  jnot g14361(.din(n14619), .dout(n14620));
  jor  g14362(.dina(n14440), .dinb(n14344), .dout(n14621));
  jand g14363(.dina(n14441), .dinb(n14336), .dout(n14622));
  jnot g14364(.din(n14622), .dout(n14623));
  jand g14365(.dina(n14623), .dinb(n14621), .dout(n14624));
  jnot g14366(.din(n14624), .dout(n14625));
  jor  g14367(.dina(n5739), .dinb(n3400), .dout(n14626));
  jor  g14368(.dina(n5574), .dinb(n3055), .dout(n14627));
  jor  g14369(.dina(n5742), .dinb(n3230), .dout(n14628));
  jor  g14370(.dina(n5744), .dinb(n3403), .dout(n14629));
  jand g14371(.dina(n14629), .dinb(n14628), .dout(n14630));
  jand g14372(.dina(n14630), .dinb(n14627), .dout(n14631));
  jand g14373(.dina(n14631), .dinb(n14626), .dout(n14632));
  jxor g14374(.dina(n14632), .dinb(a44 ), .dout(n14633));
  jnot g14375(.din(n14633), .dout(n14634));
  jor  g14376(.dina(n6490), .dinb(n3032), .dout(n14635));
  jor  g14377(.dina(n6262), .dinb(n2579), .dout(n14636));
  jor  g14378(.dina(n6493), .dinb(n2870), .dout(n14637));
  jor  g14379(.dina(n6495), .dinb(n3035), .dout(n14638));
  jand g14380(.dina(n14638), .dinb(n14637), .dout(n14639));
  jand g14381(.dina(n14639), .dinb(n14636), .dout(n14640));
  jand g14382(.dina(n14640), .dinb(n14635), .dout(n14641));
  jxor g14383(.dina(n14641), .dinb(a47 ), .dout(n14642));
  jnot g14384(.din(n14642), .dout(n14643));
  jand g14385(.dina(n14422), .dinb(n14356), .dout(n14644));
  jand g14386(.dina(n14423), .dinb(n14347), .dout(n14645));
  jor  g14387(.dina(n14645), .dinb(n14644), .dout(n14646));
  jand g14388(.dina(n14420), .dinb(n14368), .dout(n14647));
  jand g14389(.dina(n14421), .dinb(n14359), .dout(n14648));
  jor  g14390(.dina(n14648), .dinb(n14647), .dout(n14649));
  jor  g14391(.dina(n14418), .dinb(n14410), .dout(n14650));
  jand g14392(.dina(n14419), .dinb(n14373), .dout(n14651));
  jnot g14393(.din(n14651), .dout(n14652));
  jand g14394(.dina(n14652), .dinb(n14650), .dout(n14653));
  jnot g14395(.din(n14653), .dout(n14654));
  jand g14396(.dina(n14401), .dinb(n14382), .dout(n14655));
  jand g14397(.dina(n14408), .dinb(n14402), .dout(n14656));
  jor  g14398(.dina(n14656), .dinb(n14655), .dout(n14657));
  jand g14399(.dina(n14399), .dinb(n14394), .dout(n14658));
  jand g14400(.dina(n14400), .dinb(n14385), .dout(n14659));
  jor  g14401(.dina(n14659), .dinb(n14658), .dout(n14660));
  jor  g14402(.dina(n10806), .dinb(n1019), .dout(n14661));
  jor  g14403(.dina(n10485), .dinb(n858), .dout(n14662));
  jor  g14404(.dina(n10809), .dinb(n939), .dout(n14663));
  jor  g14405(.dina(n10811), .dinb(n1022), .dout(n14664));
  jand g14406(.dina(n14664), .dinb(n14663), .dout(n14665));
  jand g14407(.dina(n14665), .dinb(n14662), .dout(n14666));
  jand g14408(.dina(n14666), .dinb(n14661), .dout(n14667));
  jxor g14409(.dina(n14667), .dinb(a62 ), .dout(n14668));
  jnot g14410(.din(n14668), .dout(n14669));
  jand g14411(.dina(n13878), .dinb(n678), .dout(n14670));
  jand g14412(.dina(n14398), .dinb(n14395), .dout(n14671));
  jor  g14413(.dina(n14671), .dinb(n14670), .dout(n14672));
  jand g14414(.dina(n10801), .dinb(b13 ), .dout(n14673));
  jand g14415(.dina(n11107), .dinb(b12 ), .dout(n14674));
  jor  g14416(.dina(n14674), .dinb(n14673), .dout(n14675));
  jnot g14417(.din(n14675), .dout(n14676));
  jxor g14418(.dina(n14676), .dinb(n14672), .dout(n14677));
  jxor g14419(.dina(n14677), .dinb(n14669), .dout(n14678));
  jxor g14420(.dina(n14678), .dinb(n14660), .dout(n14679));
  jor  g14421(.dina(n9891), .dinb(n1397), .dout(n14680));
  jor  g14422(.dina(n9593), .dinb(n1193), .dout(n14681));
  jor  g14423(.dina(n9894), .dinb(n1290), .dout(n14682));
  jor  g14424(.dina(n9896), .dinb(n1400), .dout(n14683));
  jand g14425(.dina(n14683), .dinb(n14682), .dout(n14684));
  jand g14426(.dina(n14684), .dinb(n14681), .dout(n14685));
  jand g14427(.dina(n14685), .dinb(n14680), .dout(n14686));
  jxor g14428(.dina(n14686), .dinb(a59 ), .dout(n14687));
  jnot g14429(.din(n14687), .dout(n14688));
  jxor g14430(.dina(n14688), .dinb(n14679), .dout(n14689));
  jxor g14431(.dina(n14689), .dinb(n14657), .dout(n14690));
  jor  g14432(.dina(n8978), .dinb(n1739), .dout(n14691));
  jor  g14433(.dina(n8677), .dinb(n1420), .dout(n14692));
  jor  g14434(.dina(n8981), .dinb(n1620), .dout(n14693));
  jor  g14435(.dina(n8983), .dinb(n1742), .dout(n14694));
  jand g14436(.dina(n14694), .dinb(n14693), .dout(n14695));
  jand g14437(.dina(n14695), .dinb(n14692), .dout(n14696));
  jand g14438(.dina(n14696), .dinb(n14691), .dout(n14697));
  jxor g14439(.dina(n14697), .dinb(a56 ), .dout(n14698));
  jnot g14440(.din(n14698), .dout(n14699));
  jxor g14441(.dina(n14699), .dinb(n14690), .dout(n14700));
  jxor g14442(.dina(n14700), .dinb(n14654), .dout(n14701));
  jor  g14443(.dina(n8125), .dinb(n2007), .dout(n14702));
  jor  g14444(.dina(n7846), .dinb(n1867), .dout(n14703));
  jor  g14445(.dina(n8128), .dinb(n1887), .dout(n14704));
  jor  g14446(.dina(n8130), .dinb(n2010), .dout(n14705));
  jand g14447(.dina(n14705), .dinb(n14704), .dout(n14706));
  jand g14448(.dina(n14706), .dinb(n14703), .dout(n14707));
  jand g14449(.dina(n14707), .dinb(n14702), .dout(n14708));
  jxor g14450(.dina(n14708), .dinb(a53 ), .dout(n14709));
  jnot g14451(.din(n14709), .dout(n14710));
  jxor g14452(.dina(n14710), .dinb(n14701), .dout(n14711));
  jxor g14453(.dina(n14711), .dinb(n14649), .dout(n14712));
  jnot g14454(.din(n14712), .dout(n14713));
  jor  g14455(.dina(n7266), .dinb(n2556), .dout(n14714));
  jor  g14456(.dina(n7021), .dinb(n2148), .dout(n14715));
  jor  g14457(.dina(n7269), .dinb(n2407), .dout(n14716));
  jor  g14458(.dina(n7271), .dinb(n2559), .dout(n14717));
  jand g14459(.dina(n14717), .dinb(n14716), .dout(n14718));
  jand g14460(.dina(n14718), .dinb(n14715), .dout(n14719));
  jand g14461(.dina(n14719), .dinb(n14714), .dout(n14720));
  jxor g14462(.dina(n14720), .dinb(a50 ), .dout(n14721));
  jxor g14463(.dina(n14721), .dinb(n14713), .dout(n14722));
  jxor g14464(.dina(n14722), .dinb(n14646), .dout(n14723));
  jxor g14465(.dina(n14723), .dinb(n14643), .dout(n14724));
  jand g14466(.dina(n14433), .dinb(n14425), .dout(n14725));
  jnot g14467(.din(n14725), .dout(n14726));
  jnot g14468(.din(n14433), .dout(n14727));
  jand g14469(.dina(n14727), .dinb(n14424), .dout(n14728));
  jor  g14470(.dina(n14438), .dinb(n14728), .dout(n14729));
  jand g14471(.dina(n14729), .dinb(n14726), .dout(n14730));
  jxor g14472(.dina(n14730), .dinb(n14724), .dout(n14731));
  jxor g14473(.dina(n14731), .dinb(n14634), .dout(n14732));
  jxor g14474(.dina(n14732), .dinb(n14625), .dout(n14733));
  jxor g14475(.dina(n14733), .dinb(n14620), .dout(n14734));
  jxor g14476(.dina(n14734), .dinb(n14611), .dout(n14735));
  jxor g14477(.dina(n14735), .dinb(n14606), .dout(n14736));
  jxor g14478(.dina(n14736), .dinb(n14597), .dout(n14737));
  jor  g14479(.dina(n5405), .dinb(n3849), .dout(n14738));
  jor  g14480(.dina(n3689), .dinb(n4974), .dout(n14739));
  jor  g14481(.dina(n3852), .dinb(n4994), .dout(n14740));
  jor  g14482(.dina(n3854), .dinb(n5408), .dout(n14741));
  jand g14483(.dina(n14741), .dinb(n14740), .dout(n14742));
  jand g14484(.dina(n14742), .dinb(n14739), .dout(n14743));
  jand g14485(.dina(n14743), .dinb(n14738), .dout(n14744));
  jxor g14486(.dina(n14744), .dinb(a35 ), .dout(n14745));
  jnot g14487(.din(n14745), .dout(n14746));
  jxor g14488(.dina(n14746), .dinb(n14737), .dout(n14747));
  jxor g14489(.dina(n14747), .dinb(n14592), .dout(n14748));
  jor  g14490(.dina(n6864), .dinb(n2784), .dout(n14749));
  jor  g14491(.dina(n2661), .dinb(n6352), .dout(n14750));
  jor  g14492(.dina(n2787), .dinb(n6372), .dout(n14751));
  jor  g14493(.dina(n2789), .dinb(n6867), .dout(n14752));
  jand g14494(.dina(n14752), .dinb(n14751), .dout(n14753));
  jand g14495(.dina(n14753), .dinb(n14750), .dout(n14754));
  jand g14496(.dina(n14754), .dinb(n14749), .dout(n14755));
  jxor g14497(.dina(n14755), .dinb(a29 ), .dout(n14756));
  jnot g14498(.din(n14756), .dout(n14757));
  jand g14499(.dina(n14481), .dinb(n14477), .dout(n14758));
  jand g14500(.dina(n14482), .dinb(n14468), .dout(n14759));
  jor  g14501(.dina(n14759), .dinb(n14758), .dout(n14760));
  jxor g14502(.dina(n14760), .dinb(n14757), .dout(n14761));
  jxor g14503(.dina(n14761), .dinb(n14748), .dout(n14762));
  jnot g14504(.din(n14762), .dout(n14763));
  jxor g14505(.dina(n14763), .dinb(n14579), .dout(n14764));
  jnot g14506(.din(n14764), .dout(n14765));
  jor  g14507(.dina(n8228), .dinb(n1939), .dout(n14766));
  jor  g14508(.dina(n1827), .dinb(n7683), .dout(n14767));
  jor  g14509(.dina(n1942), .dinb(n7960), .dout(n14768));
  jor  g14510(.dina(n1944), .dinb(n8231), .dout(n14769));
  jand g14511(.dina(n14769), .dinb(n14768), .dout(n14770));
  jand g14512(.dina(n14770), .dinb(n14767), .dout(n14771));
  jand g14513(.dina(n14771), .dinb(n14766), .dout(n14772));
  jxor g14514(.dina(n14772), .dinb(a23 ), .dout(n14773));
  jor  g14515(.dina(n14307), .dinb(n14303), .dout(n14774));
  jand g14516(.dina(n14499), .dinb(n14308), .dout(n14775));
  jnot g14517(.din(n14775), .dout(n14776));
  jand g14518(.dina(n14776), .dinb(n14774), .dout(n14777));
  jxor g14519(.dina(n14777), .dinb(n14773), .dout(n14778));
  jxor g14520(.dina(n14778), .dinb(n14765), .dout(n14779));
  jor  g14521(.dina(n14512), .dinb(n14504), .dout(n14780));
  jand g14522(.dina(n14513), .dinb(n14500), .dout(n14781));
  jnot g14523(.din(n14781), .dout(n14782));
  jand g14524(.dina(n14782), .dinb(n14780), .dout(n14783));
  jor  g14525(.dina(n9387), .dinb(n1566), .dout(n14784));
  jor  g14526(.dina(n1489), .dinb(n8789), .dout(n14785));
  jor  g14527(.dina(n1569), .dinb(n8809), .dout(n14786));
  jor  g14528(.dina(n1571), .dinb(n9390), .dout(n14787));
  jand g14529(.dina(n14787), .dinb(n14786), .dout(n14788));
  jand g14530(.dina(n14788), .dinb(n14785), .dout(n14789));
  jand g14531(.dina(n14789), .dinb(n14784), .dout(n14790));
  jxor g14532(.dina(n14790), .dinb(a20 ), .dout(n14791));
  jxor g14533(.dina(n14791), .dinb(n14783), .dout(n14792));
  jxor g14534(.dina(n14792), .dinb(n14779), .dout(n14793));
  jxor g14535(.dina(n14793), .dinb(n14566), .dout(n14794));
  jor  g14536(.dina(n14527), .dinb(n14519), .dout(n14795));
  jand g14537(.dina(n14528), .dinb(n14515), .dout(n14796));
  jnot g14538(.din(n14796), .dout(n14797));
  jand g14539(.dina(n14797), .dinb(n14795), .dout(n14798));
  jor  g14540(.dina(n10978), .dinb(n974), .dout(n14799));
  jor  g14541(.dina(n908), .dinb(n10637), .dout(n14800));
  jor  g14542(.dina(n977), .dinb(n10964), .dout(n14801));
  jand g14543(.dina(n14801), .dinb(n14800), .dout(n14802));
  jand g14544(.dina(n14802), .dinb(n14799), .dout(n14803));
  jxor g14545(.dina(n14803), .dinb(a14 ), .dout(n14804));
  jxor g14546(.dina(n14804), .dinb(n14798), .dout(n14805));
  jxor g14547(.dina(n14805), .dinb(n14794), .dout(n14806));
  jxor g14548(.dina(n14806), .dinb(n14553), .dout(n14807));
  jxor g14549(.dina(n14807), .dinb(n14548), .dout(f76 ));
  jand g14550(.dina(n14806), .dinb(n14553), .dout(n14809));
  jand g14551(.dina(n14807), .dinb(n14548), .dout(n14810));
  jor  g14552(.dina(n14810), .dinb(n14809), .dout(n14811));
  jor  g14553(.dina(n14804), .dinb(n14798), .dout(n14812));
  jand g14554(.dina(n14805), .dinb(n14794), .dout(n14813));
  jnot g14555(.din(n14813), .dout(n14814));
  jand g14556(.dina(n14814), .dinb(n14812), .dout(n14815));
  jnot g14557(.din(n14815), .dout(n14816));
  jor  g14558(.dina(n9410), .dinb(n1566), .dout(n14817));
  jor  g14559(.dina(n1489), .dinb(n8809), .dout(n14818));
  jor  g14560(.dina(n1569), .dinb(n9390), .dout(n14819));
  jor  g14561(.dina(n1571), .dinb(n9413), .dout(n14820));
  jand g14562(.dina(n14820), .dinb(n14819), .dout(n14821));
  jand g14563(.dina(n14821), .dinb(n14818), .dout(n14822));
  jand g14564(.dina(n14822), .dinb(n14817), .dout(n14823));
  jxor g14565(.dina(n14823), .dinb(a20 ), .dout(n14824));
  jor  g14566(.dina(n14777), .dinb(n14773), .dout(n14825));
  jand g14567(.dina(n14778), .dinb(n14765), .dout(n14826));
  jnot g14568(.din(n14826), .dout(n14827));
  jand g14569(.dina(n14827), .dinb(n14825), .dout(n14828));
  jxor g14570(.dina(n14828), .dinb(n14824), .dout(n14829));
  jor  g14571(.dina(n8786), .dinb(n1939), .dout(n14830));
  jor  g14572(.dina(n1827), .dinb(n7960), .dout(n14831));
  jor  g14573(.dina(n1942), .dinb(n8231), .dout(n14832));
  jor  g14574(.dina(n1944), .dinb(n8789), .dout(n14833));
  jand g14575(.dina(n14833), .dinb(n14832), .dout(n14834));
  jand g14576(.dina(n14834), .dinb(n14831), .dout(n14835));
  jand g14577(.dina(n14835), .dinb(n14830), .dout(n14836));
  jxor g14578(.dina(n14836), .dinb(a23 ), .dout(n14837));
  jnot g14579(.din(n14837), .dout(n14838));
  jand g14580(.dina(n14578), .dinb(n14570), .dout(n14839));
  jnot g14581(.din(n14839), .dout(n14840));
  jnot g14582(.din(n14570), .dout(n14841));
  jnot g14583(.din(n14578), .dout(n14842));
  jand g14584(.dina(n14842), .dinb(n14841), .dout(n14843));
  jor  g14585(.dina(n14762), .dinb(n14843), .dout(n14844));
  jand g14586(.dina(n14844), .dinb(n14840), .dout(n14845));
  jxor g14587(.dina(n14845), .dinb(n14838), .dout(n14846));
  jnot g14588(.din(n14846), .dout(n14847));
  jor  g14589(.dina(n7680), .dinb(n2319), .dout(n14848));
  jor  g14590(.dina(n2224), .dinb(n7149), .dout(n14849));
  jor  g14591(.dina(n2322), .dinb(n7411), .dout(n14850));
  jor  g14592(.dina(n2324), .dinb(n7683), .dout(n14851));
  jand g14593(.dina(n14851), .dinb(n14850), .dout(n14852));
  jand g14594(.dina(n14852), .dinb(n14849), .dout(n14853));
  jand g14595(.dina(n14853), .dinb(n14848), .dout(n14854));
  jxor g14596(.dina(n14854), .dinb(a26 ), .dout(n14855));
  jand g14597(.dina(n14760), .dinb(n14757), .dout(n14856));
  jand g14598(.dina(n14761), .dinb(n14748), .dout(n14857));
  jor  g14599(.dina(n14857), .dinb(n14856), .dout(n14858));
  jnot g14600(.din(n14858), .dout(n14859));
  jxor g14601(.dina(n14859), .dinb(n14855), .dout(n14860));
  jor  g14602(.dina(n14591), .dinb(n14583), .dout(n14861));
  jand g14603(.dina(n14747), .dinb(n14592), .dout(n14862));
  jnot g14604(.din(n14862), .dout(n14863));
  jand g14605(.dina(n14863), .dinb(n14861), .dout(n14864));
  jor  g14606(.dina(n7126), .dinb(n2784), .dout(n14865));
  jor  g14607(.dina(n2661), .dinb(n6372), .dout(n14866));
  jor  g14608(.dina(n2787), .dinb(n6867), .dout(n14867));
  jor  g14609(.dina(n2789), .dinb(n7129), .dout(n14868));
  jand g14610(.dina(n14868), .dinb(n14867), .dout(n14869));
  jand g14611(.dina(n14869), .dinb(n14866), .dout(n14870));
  jand g14612(.dina(n14870), .dinb(n14865), .dout(n14871));
  jxor g14613(.dina(n14871), .dinb(a29 ), .dout(n14872));
  jxor g14614(.dina(n14872), .dinb(n14864), .dout(n14873));
  jor  g14615(.dina(n6349), .dinb(n3301), .dout(n14874));
  jor  g14616(.dina(n3136), .dinb(n5862), .dout(n14875));
  jor  g14617(.dina(n3304), .dinb(n6106), .dout(n14876));
  jor  g14618(.dina(n3306), .dinb(n6352), .dout(n14877));
  jand g14619(.dina(n14877), .dinb(n14876), .dout(n14878));
  jand g14620(.dina(n14878), .dinb(n14875), .dout(n14879));
  jand g14621(.dina(n14879), .dinb(n14874), .dout(n14880));
  jxor g14622(.dina(n14880), .dinb(a32 ), .dout(n14881));
  jnot g14623(.din(n14881), .dout(n14882));
  jor  g14624(.dina(n14736), .dinb(n14597), .dout(n14883));
  jand g14625(.dina(n14736), .dinb(n14597), .dout(n14884));
  jor  g14626(.dina(n14746), .dinb(n14884), .dout(n14885));
  jand g14627(.dina(n14885), .dinb(n14883), .dout(n14886));
  jxor g14628(.dina(n14886), .dinb(n14882), .dout(n14887));
  jor  g14629(.dina(n5425), .dinb(n3849), .dout(n14888));
  jor  g14630(.dina(n3689), .dinb(n4994), .dout(n14889));
  jor  g14631(.dina(n3852), .dinb(n5408), .dout(n14890));
  jor  g14632(.dina(n3854), .dinb(n5428), .dout(n14891));
  jand g14633(.dina(n14891), .dinb(n14890), .dout(n14892));
  jand g14634(.dina(n14892), .dinb(n14889), .dout(n14893));
  jand g14635(.dina(n14893), .dinb(n14888), .dout(n14894));
  jxor g14636(.dina(n14894), .dinb(a35 ), .dout(n14895));
  jnot g14637(.din(n14895), .dout(n14896));
  jand g14638(.dina(n14734), .dinb(n14611), .dout(n14897));
  jand g14639(.dina(n14735), .dinb(n14606), .dout(n14898));
  jor  g14640(.dina(n14898), .dinb(n14897), .dout(n14899));
  jor  g14641(.dina(n4971), .dinb(n4415), .dout(n14900));
  jor  g14642(.dina(n4272), .dinb(n4537), .dout(n14901));
  jor  g14643(.dina(n4418), .dinb(n4557), .dout(n14902));
  jor  g14644(.dina(n4420), .dinb(n4974), .dout(n14903));
  jand g14645(.dina(n14903), .dinb(n14902), .dout(n14904));
  jand g14646(.dina(n14904), .dinb(n14901), .dout(n14905));
  jand g14647(.dina(n14905), .dinb(n14900), .dout(n14906));
  jxor g14648(.dina(n14906), .dinb(a38 ), .dout(n14907));
  jnot g14649(.din(n14907), .dout(n14908));
  jand g14650(.dina(n14732), .dinb(n14625), .dout(n14909));
  jand g14651(.dina(n14733), .dinb(n14620), .dout(n14910));
  jor  g14652(.dina(n14910), .dinb(n14909), .dout(n14911));
  jand g14653(.dina(n14730), .dinb(n14724), .dout(n14912));
  jand g14654(.dina(n14731), .dinb(n14634), .dout(n14913));
  jor  g14655(.dina(n14913), .dinb(n14912), .dout(n14914));
  jand g14656(.dina(n14722), .dinb(n14646), .dout(n14915));
  jand g14657(.dina(n14723), .dinb(n14643), .dout(n14916));
  jor  g14658(.dina(n14916), .dinb(n14915), .dout(n14917));
  jor  g14659(.dina(n6490), .dinb(n3052), .dout(n14918));
  jor  g14660(.dina(n6262), .dinb(n2870), .dout(n14919));
  jor  g14661(.dina(n6493), .dinb(n3035), .dout(n14920));
  jor  g14662(.dina(n6495), .dinb(n3055), .dout(n14921));
  jand g14663(.dina(n14921), .dinb(n14920), .dout(n14922));
  jand g14664(.dina(n14922), .dinb(n14919), .dout(n14923));
  jand g14665(.dina(n14923), .dinb(n14918), .dout(n14924));
  jxor g14666(.dina(n14924), .dinb(a47 ), .dout(n14925));
  jnot g14667(.din(n14925), .dout(n14926));
  jand g14668(.dina(n14711), .dinb(n14649), .dout(n14927));
  jnot g14669(.din(n14927), .dout(n14928));
  jor  g14670(.dina(n14721), .dinb(n14713), .dout(n14929));
  jand g14671(.dina(n14929), .dinb(n14928), .dout(n14930));
  jnot g14672(.din(n14930), .dout(n14931));
  jor  g14673(.dina(n8125), .dinb(n2145), .dout(n14932));
  jor  g14674(.dina(n7846), .dinb(n1887), .dout(n14933));
  jor  g14675(.dina(n8128), .dinb(n2010), .dout(n14934));
  jor  g14676(.dina(n8130), .dinb(n2148), .dout(n14935));
  jand g14677(.dina(n14935), .dinb(n14934), .dout(n14936));
  jand g14678(.dina(n14936), .dinb(n14933), .dout(n14937));
  jand g14679(.dina(n14937), .dinb(n14932), .dout(n14938));
  jxor g14680(.dina(n14938), .dinb(a53 ), .dout(n14939));
  jnot g14681(.din(n14939), .dout(n14940));
  jand g14682(.dina(n14676), .dinb(n14672), .dout(n14941));
  jand g14683(.dina(n14677), .dinb(n14669), .dout(n14942));
  jor  g14684(.dina(n14942), .dinb(n14941), .dout(n14943));
  jand g14685(.dina(n10801), .dinb(b14 ), .dout(n14944));
  jand g14686(.dina(n11107), .dinb(b13 ), .dout(n14945));
  jor  g14687(.dina(n14945), .dinb(n14944), .dout(n14946));
  jxor g14688(.dina(n14946), .dinb(n14676), .dout(n14947));
  jnot g14689(.din(n14947), .dout(n14948));
  jor  g14690(.dina(n10806), .dinb(n1190), .dout(n14949));
  jor  g14691(.dina(n10485), .dinb(n939), .dout(n14950));
  jor  g14692(.dina(n10809), .dinb(n1022), .dout(n14951));
  jor  g14693(.dina(n10811), .dinb(n1193), .dout(n14952));
  jand g14694(.dina(n14952), .dinb(n14951), .dout(n14953));
  jand g14695(.dina(n14953), .dinb(n14950), .dout(n14954));
  jand g14696(.dina(n14954), .dinb(n14949), .dout(n14955));
  jxor g14697(.dina(n14955), .dinb(a62 ), .dout(n14956));
  jxor g14698(.dina(n14956), .dinb(n14948), .dout(n14957));
  jxor g14699(.dina(n14957), .dinb(n14943), .dout(n14958));
  jor  g14700(.dina(n9891), .dinb(n1417), .dout(n14959));
  jor  g14701(.dina(n9593), .dinb(n1290), .dout(n14960));
  jor  g14702(.dina(n9894), .dinb(n1400), .dout(n14961));
  jor  g14703(.dina(n9896), .dinb(n1420), .dout(n14962));
  jand g14704(.dina(n14962), .dinb(n14961), .dout(n14963));
  jand g14705(.dina(n14963), .dinb(n14960), .dout(n14964));
  jand g14706(.dina(n14964), .dinb(n14959), .dout(n14965));
  jxor g14707(.dina(n14965), .dinb(a59 ), .dout(n14966));
  jnot g14708(.din(n14966), .dout(n14967));
  jxor g14709(.dina(n14967), .dinb(n14958), .dout(n14968));
  jnot g14710(.din(n14660), .dout(n14969));
  jnot g14711(.din(n14678), .dout(n14970));
  jand g14712(.dina(n14970), .dinb(n14969), .dout(n14971));
  jnot g14713(.din(n14971), .dout(n14972));
  jand g14714(.dina(n14678), .dinb(n14660), .dout(n14973));
  jor  g14715(.dina(n14688), .dinb(n14973), .dout(n14974));
  jand g14716(.dina(n14974), .dinb(n14972), .dout(n14975));
  jxor g14717(.dina(n14975), .dinb(n14968), .dout(n14976));
  jnot g14718(.din(n14976), .dout(n14977));
  jor  g14719(.dina(n8978), .dinb(n1864), .dout(n14978));
  jor  g14720(.dina(n8677), .dinb(n1620), .dout(n14979));
  jor  g14721(.dina(n8981), .dinb(n1742), .dout(n14980));
  jor  g14722(.dina(n8983), .dinb(n1867), .dout(n14981));
  jand g14723(.dina(n14981), .dinb(n14980), .dout(n14982));
  jand g14724(.dina(n14982), .dinb(n14979), .dout(n14983));
  jand g14725(.dina(n14983), .dinb(n14978), .dout(n14984));
  jxor g14726(.dina(n14984), .dinb(a56 ), .dout(n14985));
  jxor g14727(.dina(n14985), .dinb(n14977), .dout(n14986));
  jnot g14728(.din(n14657), .dout(n14987));
  jnot g14729(.din(n14689), .dout(n14988));
  jand g14730(.dina(n14988), .dinb(n14987), .dout(n14989));
  jnot g14731(.din(n14989), .dout(n14990));
  jand g14732(.dina(n14689), .dinb(n14657), .dout(n14991));
  jor  g14733(.dina(n14699), .dinb(n14991), .dout(n14992));
  jand g14734(.dina(n14992), .dinb(n14990), .dout(n14993));
  jxor g14735(.dina(n14993), .dinb(n14986), .dout(n14994));
  jxor g14736(.dina(n14994), .dinb(n14940), .dout(n14995));
  jnot g14737(.din(n14700), .dout(n14996));
  jand g14738(.dina(n14996), .dinb(n14653), .dout(n14997));
  jnot g14739(.din(n14997), .dout(n14998));
  jand g14740(.dina(n14700), .dinb(n14654), .dout(n14999));
  jor  g14741(.dina(n14710), .dinb(n14999), .dout(n15000));
  jand g14742(.dina(n15000), .dinb(n14998), .dout(n15001));
  jxor g14743(.dina(n15001), .dinb(n14995), .dout(n15002));
  jor  g14744(.dina(n7266), .dinb(n2576), .dout(n15003));
  jor  g14745(.dina(n7021), .dinb(n2407), .dout(n15004));
  jor  g14746(.dina(n7269), .dinb(n2559), .dout(n15005));
  jor  g14747(.dina(n7271), .dinb(n2579), .dout(n15006));
  jand g14748(.dina(n15006), .dinb(n15005), .dout(n15007));
  jand g14749(.dina(n15007), .dinb(n15004), .dout(n15008));
  jand g14750(.dina(n15008), .dinb(n15003), .dout(n15009));
  jxor g14751(.dina(n15009), .dinb(a50 ), .dout(n15010));
  jnot g14752(.din(n15010), .dout(n15011));
  jxor g14753(.dina(n15011), .dinb(n15002), .dout(n15012));
  jxor g14754(.dina(n15012), .dinb(n14931), .dout(n15013));
  jxor g14755(.dina(n15013), .dinb(n14926), .dout(n15014));
  jxor g14756(.dina(n15014), .dinb(n14917), .dout(n15015));
  jor  g14757(.dina(n5739), .dinb(n3585), .dout(n15016));
  jor  g14758(.dina(n5574), .dinb(n3230), .dout(n15017));
  jor  g14759(.dina(n5742), .dinb(n3403), .dout(n15018));
  jor  g14760(.dina(n5744), .dinb(n3588), .dout(n15019));
  jand g14761(.dina(n15019), .dinb(n15018), .dout(n15020));
  jand g14762(.dina(n15020), .dinb(n15017), .dout(n15021));
  jand g14763(.dina(n15021), .dinb(n15016), .dout(n15022));
  jxor g14764(.dina(n15022), .dinb(a44 ), .dout(n15023));
  jnot g14765(.din(n15023), .dout(n15024));
  jxor g14766(.dina(n15024), .dinb(n15015), .dout(n15025));
  jxor g14767(.dina(n15025), .dinb(n14914), .dout(n15026));
  jnot g14768(.din(n15026), .dout(n15027));
  jor  g14769(.dina(n5096), .dinb(n4337), .dout(n15028));
  jor  g14770(.dina(n4904), .dinb(n3942), .dout(n15029));
  jor  g14771(.dina(n5099), .dinb(n4140), .dout(n15030));
  jor  g14772(.dina(n5101), .dinb(n4340), .dout(n15031));
  jand g14773(.dina(n15031), .dinb(n15030), .dout(n15032));
  jand g14774(.dina(n15032), .dinb(n15029), .dout(n15033));
  jand g14775(.dina(n15033), .dinb(n15028), .dout(n15034));
  jxor g14776(.dina(n15034), .dinb(a41 ), .dout(n15035));
  jxor g14777(.dina(n15035), .dinb(n15027), .dout(n15036));
  jxor g14778(.dina(n15036), .dinb(n14911), .dout(n15037));
  jxor g14779(.dina(n15037), .dinb(n14908), .dout(n15038));
  jxor g14780(.dina(n15038), .dinb(n14899), .dout(n15039));
  jxor g14781(.dina(n15039), .dinb(n14896), .dout(n15040));
  jxor g14782(.dina(n15040), .dinb(n14887), .dout(n15041));
  jxor g14783(.dina(n15041), .dinb(n14873), .dout(n15042));
  jnot g14784(.din(n15042), .dout(n15043));
  jxor g14785(.dina(n15043), .dinb(n14860), .dout(n15044));
  jxor g14786(.dina(n15044), .dinb(n14847), .dout(n15045));
  jxor g14787(.dina(n15045), .dinb(n14829), .dout(n15046));
  jor  g14788(.dina(n14791), .dinb(n14783), .dout(n15047));
  jand g14789(.dina(n14792), .dinb(n14779), .dout(n15048));
  jnot g14790(.din(n15048), .dout(n15049));
  jand g14791(.dina(n15049), .dinb(n15047), .dout(n15050));
  jor  g14792(.dina(n10634), .dinb(n1245), .dout(n15051));
  jor  g14793(.dina(n1165), .dinb(n9725), .dout(n15052));
  jor  g14794(.dina(n1248), .dinb(n10314), .dout(n15053));
  jor  g14795(.dina(n1250), .dinb(n10637), .dout(n15054));
  jand g14796(.dina(n15054), .dinb(n15053), .dout(n15055));
  jand g14797(.dina(n15055), .dinb(n15052), .dout(n15056));
  jand g14798(.dina(n15056), .dinb(n15051), .dout(n15057));
  jxor g14799(.dina(n15057), .dinb(a17 ), .dout(n15058));
  jxor g14800(.dina(n15058), .dinb(n15050), .dout(n15059));
  jxor g14801(.dina(n15059), .dinb(n15046), .dout(n15060));
  jand g14802(.dina(n14565), .dinb(n14562), .dout(n15061));
  jand g14803(.dina(n14793), .dinb(n14566), .dout(n15062));
  jor  g14804(.dina(n15062), .dinb(n15061), .dout(n15063));
  jnot g14805(.din(n15063), .dout(n15064));
  jnot g14806(.din(a14 ), .dout(n15065));
  jand g14807(.dina(n11296), .dinb(n815), .dout(n15066));
  jor  g14808(.dina(n15066), .dinb(n909), .dout(n15067));
  jand g14809(.dina(n15067), .dinb(b63 ), .dout(n15068));
  jxor g14810(.dina(n15068), .dinb(n15065), .dout(n15069));
  jxor g14811(.dina(n15069), .dinb(n15064), .dout(n15070));
  jxor g14812(.dina(n15070), .dinb(n15060), .dout(n15071));
  jxor g14813(.dina(n15071), .dinb(n14816), .dout(n15072));
  jxor g14814(.dina(n15072), .dinb(n14811), .dout(f77 ));
  jor  g14815(.dina(n15069), .dinb(n15064), .dout(n15074));
  jand g14816(.dina(n15070), .dinb(n15060), .dout(n15075));
  jnot g14817(.din(n15075), .dout(n15076));
  jand g14818(.dina(n15076), .dinb(n15074), .dout(n15077));
  jnot g14819(.din(n15077), .dout(n15078));
  jor  g14820(.dina(n9722), .dinb(n1566), .dout(n15079));
  jor  g14821(.dina(n1489), .dinb(n9390), .dout(n15080));
  jor  g14822(.dina(n1569), .dinb(n9413), .dout(n15081));
  jor  g14823(.dina(n1571), .dinb(n9725), .dout(n15082));
  jand g14824(.dina(n15082), .dinb(n15081), .dout(n15083));
  jand g14825(.dina(n15083), .dinb(n15080), .dout(n15084));
  jand g14826(.dina(n15084), .dinb(n15079), .dout(n15085));
  jxor g14827(.dina(n15085), .dinb(a20 ), .dout(n15086));
  jor  g14828(.dina(n14828), .dinb(n14824), .dout(n15087));
  jand g14829(.dina(n15045), .dinb(n14829), .dout(n15088));
  jnot g14830(.din(n15088), .dout(n15089));
  jand g14831(.dina(n15089), .dinb(n15087), .dout(n15090));
  jxor g14832(.dina(n15090), .dinb(n15086), .dout(n15091));
  jand g14833(.dina(n14845), .dinb(n14838), .dout(n15092));
  jnot g14834(.din(n15092), .dout(n15093));
  jor  g14835(.dina(n15044), .dinb(n14847), .dout(n15094));
  jand g14836(.dina(n15094), .dinb(n15093), .dout(n15095));
  jor  g14837(.dina(n8806), .dinb(n1939), .dout(n15096));
  jor  g14838(.dina(n1827), .dinb(n8231), .dout(n15097));
  jor  g14839(.dina(n1942), .dinb(n8789), .dout(n15098));
  jor  g14840(.dina(n1944), .dinb(n8809), .dout(n15099));
  jand g14841(.dina(n15099), .dinb(n15098), .dout(n15100));
  jand g14842(.dina(n15100), .dinb(n15097), .dout(n15101));
  jand g14843(.dina(n15101), .dinb(n15096), .dout(n15102));
  jxor g14844(.dina(n15102), .dinb(a23 ), .dout(n15103));
  jxor g14845(.dina(n15103), .dinb(n15095), .dout(n15104));
  jor  g14846(.dina(n7957), .dinb(n2319), .dout(n15105));
  jor  g14847(.dina(n2224), .dinb(n7411), .dout(n15106));
  jor  g14848(.dina(n2322), .dinb(n7683), .dout(n15107));
  jor  g14849(.dina(n2324), .dinb(n7960), .dout(n15108));
  jand g14850(.dina(n15108), .dinb(n15107), .dout(n15109));
  jand g14851(.dina(n15109), .dinb(n15106), .dout(n15110));
  jand g14852(.dina(n15110), .dinb(n15105), .dout(n15111));
  jxor g14853(.dina(n15111), .dinb(a26 ), .dout(n15112));
  jnot g14854(.din(n15112), .dout(n15113));
  jand g14855(.dina(n14859), .dinb(n14855), .dout(n15114));
  jnot g14856(.din(n15114), .dout(n15115));
  jnot g14857(.din(n14855), .dout(n15116));
  jand g14858(.dina(n14858), .dinb(n15116), .dout(n15117));
  jor  g14859(.dina(n15042), .dinb(n15117), .dout(n15118));
  jand g14860(.dina(n15118), .dinb(n15115), .dout(n15119));
  jxor g14861(.dina(n15119), .dinb(n15113), .dout(n15120));
  jor  g14862(.dina(n7146), .dinb(n2784), .dout(n15121));
  jor  g14863(.dina(n2661), .dinb(n6867), .dout(n15122));
  jor  g14864(.dina(n2787), .dinb(n7129), .dout(n15123));
  jor  g14865(.dina(n2789), .dinb(n7149), .dout(n15124));
  jand g14866(.dina(n15124), .dinb(n15123), .dout(n15125));
  jand g14867(.dina(n15125), .dinb(n15122), .dout(n15126));
  jand g14868(.dina(n15126), .dinb(n15121), .dout(n15127));
  jxor g14869(.dina(n15127), .dinb(a29 ), .dout(n15128));
  jnot g14870(.din(n15128), .dout(n15129));
  jand g14871(.dina(n14872), .dinb(n14864), .dout(n15130));
  jnot g14872(.din(n15130), .dout(n15131));
  jnot g14873(.din(n14864), .dout(n15132));
  jnot g14874(.din(n14872), .dout(n15133));
  jand g14875(.dina(n15133), .dinb(n15132), .dout(n15134));
  jor  g14876(.dina(n15041), .dinb(n15134), .dout(n15135));
  jand g14877(.dina(n15135), .dinb(n15131), .dout(n15136));
  jxor g14878(.dina(n15136), .dinb(n15129), .dout(n15137));
  jand g14879(.dina(n15036), .dinb(n14911), .dout(n15138));
  jand g14880(.dina(n15037), .dinb(n14908), .dout(n15139));
  jor  g14881(.dina(n15139), .dinb(n15138), .dout(n15140));
  jor  g14882(.dina(n4991), .dinb(n4415), .dout(n15141));
  jor  g14883(.dina(n4272), .dinb(n4557), .dout(n15142));
  jor  g14884(.dina(n4418), .dinb(n4974), .dout(n15143));
  jor  g14885(.dina(n4420), .dinb(n4994), .dout(n15144));
  jand g14886(.dina(n15144), .dinb(n15143), .dout(n15145));
  jand g14887(.dina(n15145), .dinb(n15142), .dout(n15146));
  jand g14888(.dina(n15146), .dinb(n15141), .dout(n15147));
  jxor g14889(.dina(n15147), .dinb(a38 ), .dout(n15148));
  jnot g14890(.din(n15148), .dout(n15149));
  jand g14891(.dina(n15025), .dinb(n14914), .dout(n15150));
  jnot g14892(.din(n15150), .dout(n15151));
  jor  g14893(.dina(n15035), .dinb(n15027), .dout(n15152));
  jand g14894(.dina(n15152), .dinb(n15151), .dout(n15153));
  jnot g14895(.din(n15153), .dout(n15154));
  jor  g14896(.dina(n5739), .dinb(n3939), .dout(n15155));
  jor  g14897(.dina(n5574), .dinb(n3403), .dout(n15156));
  jor  g14898(.dina(n5742), .dinb(n3588), .dout(n15157));
  jor  g14899(.dina(n5744), .dinb(n3942), .dout(n15158));
  jand g14900(.dina(n15158), .dinb(n15157), .dout(n15159));
  jand g14901(.dina(n15159), .dinb(n15156), .dout(n15160));
  jand g14902(.dina(n15160), .dinb(n15155), .dout(n15161));
  jxor g14903(.dina(n15161), .dinb(a44 ), .dout(n15162));
  jnot g14904(.din(n15162), .dout(n15163));
  jand g14905(.dina(n15012), .dinb(n14931), .dout(n15164));
  jand g14906(.dina(n15013), .dinb(n14926), .dout(n15165));
  jor  g14907(.dina(n15165), .dinb(n15164), .dout(n15166));
  jand g14908(.dina(n14993), .dinb(n14986), .dout(n15167));
  jand g14909(.dina(n14994), .dinb(n14940), .dout(n15168));
  jor  g14910(.dina(n15168), .dinb(n15167), .dout(n15169));
  jor  g14911(.dina(n8125), .dinb(n2404), .dout(n15170));
  jor  g14912(.dina(n7846), .dinb(n2010), .dout(n15171));
  jor  g14913(.dina(n8128), .dinb(n2148), .dout(n15172));
  jor  g14914(.dina(n8130), .dinb(n2407), .dout(n15173));
  jand g14915(.dina(n15173), .dinb(n15172), .dout(n15174));
  jand g14916(.dina(n15174), .dinb(n15171), .dout(n15175));
  jand g14917(.dina(n15175), .dinb(n15170), .dout(n15176));
  jxor g14918(.dina(n15176), .dinb(a53 ), .dout(n15177));
  jand g14919(.dina(n14975), .dinb(n14968), .dout(n15178));
  jnot g14920(.din(n15178), .dout(n15179));
  jor  g14921(.dina(n14985), .dinb(n14977), .dout(n15180));
  jand g14922(.dina(n15180), .dinb(n15179), .dout(n15181));
  jand g14923(.dina(n14946), .dinb(n14676), .dout(n15182));
  jnot g14924(.din(n15182), .dout(n15183));
  jor  g14925(.dina(n14956), .dinb(n14948), .dout(n15184));
  jand g14926(.dina(n15184), .dinb(n15183), .dout(n15185));
  jnot g14927(.din(n15185), .dout(n15186));
  jor  g14928(.dina(n10806), .dinb(n1287), .dout(n15187));
  jor  g14929(.dina(n10485), .dinb(n1022), .dout(n15188));
  jor  g14930(.dina(n10809), .dinb(n1193), .dout(n15189));
  jor  g14931(.dina(n10811), .dinb(n1290), .dout(n15190));
  jand g14932(.dina(n15190), .dinb(n15189), .dout(n15191));
  jand g14933(.dina(n15191), .dinb(n15188), .dout(n15192));
  jand g14934(.dina(n15192), .dinb(n15187), .dout(n15193));
  jxor g14935(.dina(n15193), .dinb(a62 ), .dout(n15194));
  jnot g14936(.din(n15194), .dout(n15195));
  jand g14937(.dina(n10801), .dinb(b15 ), .dout(n15196));
  jand g14938(.dina(n11107), .dinb(b14 ), .dout(n15197));
  jor  g14939(.dina(n15197), .dinb(n15196), .dout(n15198));
  jxor g14940(.dina(n15198), .dinb(n15065), .dout(n15199));
  jxor g14941(.dina(n15199), .dinb(n14675), .dout(n15200));
  jxor g14942(.dina(n15200), .dinb(n15195), .dout(n15201));
  jxor g14943(.dina(n15201), .dinb(n15186), .dout(n15202));
  jnot g14944(.din(n15202), .dout(n15203));
  jor  g14945(.dina(n9891), .dinb(n1617), .dout(n15204));
  jor  g14946(.dina(n9593), .dinb(n1400), .dout(n15205));
  jor  g14947(.dina(n9894), .dinb(n1420), .dout(n15206));
  jor  g14948(.dina(n9896), .dinb(n1620), .dout(n15207));
  jand g14949(.dina(n15207), .dinb(n15206), .dout(n15208));
  jand g14950(.dina(n15208), .dinb(n15205), .dout(n15209));
  jand g14951(.dina(n15209), .dinb(n15204), .dout(n15210));
  jxor g14952(.dina(n15210), .dinb(a59 ), .dout(n15211));
  jxor g14953(.dina(n15211), .dinb(n15203), .dout(n15212));
  jor  g14954(.dina(n14957), .dinb(n14943), .dout(n15213));
  jand g14955(.dina(n14957), .dinb(n14943), .dout(n15214));
  jor  g14956(.dina(n14967), .dinb(n15214), .dout(n15215));
  jand g14957(.dina(n15215), .dinb(n15213), .dout(n15216));
  jxor g14958(.dina(n15216), .dinb(n15212), .dout(n15217));
  jnot g14959(.din(n15217), .dout(n15218));
  jor  g14960(.dina(n8978), .dinb(n1884), .dout(n15219));
  jor  g14961(.dina(n8677), .dinb(n1742), .dout(n15220));
  jor  g14962(.dina(n8981), .dinb(n1867), .dout(n15221));
  jor  g14963(.dina(n8983), .dinb(n1887), .dout(n15222));
  jand g14964(.dina(n15222), .dinb(n15221), .dout(n15223));
  jand g14965(.dina(n15223), .dinb(n15220), .dout(n15224));
  jand g14966(.dina(n15224), .dinb(n15219), .dout(n15225));
  jxor g14967(.dina(n15225), .dinb(a56 ), .dout(n15226));
  jxor g14968(.dina(n15226), .dinb(n15218), .dout(n15227));
  jxor g14969(.dina(n15227), .dinb(n15181), .dout(n15228));
  jxor g14970(.dina(n15228), .dinb(n15177), .dout(n15229));
  jxor g14971(.dina(n15229), .dinb(n15169), .dout(n15230));
  jnot g14972(.din(n15230), .dout(n15231));
  jor  g14973(.dina(n7266), .dinb(n2867), .dout(n15232));
  jor  g14974(.dina(n7021), .dinb(n2559), .dout(n15233));
  jor  g14975(.dina(n7269), .dinb(n2579), .dout(n15234));
  jor  g14976(.dina(n7271), .dinb(n2870), .dout(n15235));
  jand g14977(.dina(n15235), .dinb(n15234), .dout(n15236));
  jand g14978(.dina(n15236), .dinb(n15233), .dout(n15237));
  jand g14979(.dina(n15237), .dinb(n15232), .dout(n15238));
  jxor g14980(.dina(n15238), .dinb(a50 ), .dout(n15239));
  jxor g14981(.dina(n15239), .dinb(n15231), .dout(n15240));
  jor  g14982(.dina(n15001), .dinb(n14995), .dout(n15241));
  jand g14983(.dina(n15001), .dinb(n14995), .dout(n15242));
  jor  g14984(.dina(n15011), .dinb(n15242), .dout(n15243));
  jand g14985(.dina(n15243), .dinb(n15241), .dout(n15244));
  jxor g14986(.dina(n15244), .dinb(n15240), .dout(n15245));
  jnot g14987(.din(n15245), .dout(n15246));
  jor  g14988(.dina(n6490), .dinb(n3227), .dout(n15247));
  jor  g14989(.dina(n6262), .dinb(n3035), .dout(n15248));
  jor  g14990(.dina(n6493), .dinb(n3055), .dout(n15249));
  jor  g14991(.dina(n6495), .dinb(n3230), .dout(n15250));
  jand g14992(.dina(n15250), .dinb(n15249), .dout(n15251));
  jand g14993(.dina(n15251), .dinb(n15248), .dout(n15252));
  jand g14994(.dina(n15252), .dinb(n15247), .dout(n15253));
  jxor g14995(.dina(n15253), .dinb(a47 ), .dout(n15254));
  jxor g14996(.dina(n15254), .dinb(n15246), .dout(n15255));
  jxor g14997(.dina(n15255), .dinb(n15166), .dout(n15256));
  jxor g14998(.dina(n15256), .dinb(n15163), .dout(n15257));
  jnot g14999(.din(n14917), .dout(n15258));
  jnot g15000(.din(n15014), .dout(n15259));
  jand g15001(.dina(n15259), .dinb(n15258), .dout(n15260));
  jnot g15002(.din(n15260), .dout(n15261));
  jand g15003(.dina(n15014), .dinb(n14917), .dout(n15262));
  jor  g15004(.dina(n15024), .dinb(n15262), .dout(n15263));
  jand g15005(.dina(n15263), .dinb(n15261), .dout(n15264));
  jxor g15006(.dina(n15264), .dinb(n15257), .dout(n15265));
  jnot g15007(.din(n15265), .dout(n15266));
  jor  g15008(.dina(n5096), .dinb(n4534), .dout(n15267));
  jor  g15009(.dina(n4904), .dinb(n4140), .dout(n15268));
  jor  g15010(.dina(n5099), .dinb(n4340), .dout(n15269));
  jor  g15011(.dina(n5101), .dinb(n4537), .dout(n15270));
  jand g15012(.dina(n15270), .dinb(n15269), .dout(n15271));
  jand g15013(.dina(n15271), .dinb(n15268), .dout(n15272));
  jand g15014(.dina(n15272), .dinb(n15267), .dout(n15273));
  jxor g15015(.dina(n15273), .dinb(a41 ), .dout(n15274));
  jxor g15016(.dina(n15274), .dinb(n15266), .dout(n15275));
  jxor g15017(.dina(n15275), .dinb(n15154), .dout(n15276));
  jxor g15018(.dina(n15276), .dinb(n15149), .dout(n15277));
  jxor g15019(.dina(n15277), .dinb(n15140), .dout(n15278));
  jnot g15020(.din(n15278), .dout(n15279));
  jor  g15021(.dina(n5859), .dinb(n3849), .dout(n15280));
  jor  g15022(.dina(n3689), .dinb(n5408), .dout(n15281));
  jor  g15023(.dina(n3852), .dinb(n5428), .dout(n15282));
  jor  g15024(.dina(n3854), .dinb(n5862), .dout(n15283));
  jand g15025(.dina(n15283), .dinb(n15282), .dout(n15284));
  jand g15026(.dina(n15284), .dinb(n15281), .dout(n15285));
  jand g15027(.dina(n15285), .dinb(n15280), .dout(n15286));
  jxor g15028(.dina(n15286), .dinb(a35 ), .dout(n15287));
  jxor g15029(.dina(n15287), .dinb(n15279), .dout(n15288));
  jor  g15030(.dina(n15038), .dinb(n14899), .dout(n15289));
  jand g15031(.dina(n15038), .dinb(n14899), .dout(n15290));
  jor  g15032(.dina(n15290), .dinb(n14896), .dout(n15291));
  jand g15033(.dina(n15291), .dinb(n15289), .dout(n15292));
  jxor g15034(.dina(n15292), .dinb(n15288), .dout(n15293));
  jor  g15035(.dina(n6369), .dinb(n3301), .dout(n15294));
  jor  g15036(.dina(n3136), .dinb(n6106), .dout(n15295));
  jor  g15037(.dina(n3304), .dinb(n6352), .dout(n15296));
  jor  g15038(.dina(n3306), .dinb(n6372), .dout(n15297));
  jand g15039(.dina(n15297), .dinb(n15296), .dout(n15298));
  jand g15040(.dina(n15298), .dinb(n15295), .dout(n15299));
  jand g15041(.dina(n15299), .dinb(n15294), .dout(n15300));
  jxor g15042(.dina(n15300), .dinb(a32 ), .dout(n15301));
  jnot g15043(.din(n15301), .dout(n15302));
  jor  g15044(.dina(n14886), .dinb(n14882), .dout(n15303));
  jand g15045(.dina(n14886), .dinb(n14882), .dout(n15304));
  jor  g15046(.dina(n15040), .dinb(n15304), .dout(n15305));
  jand g15047(.dina(n15305), .dinb(n15303), .dout(n15306));
  jxor g15048(.dina(n15306), .dinb(n15302), .dout(n15307));
  jxor g15049(.dina(n15307), .dinb(n15293), .dout(n15308));
  jxor g15050(.dina(n15308), .dinb(n15137), .dout(n15309));
  jxor g15051(.dina(n15309), .dinb(n15120), .dout(n15310));
  jxor g15052(.dina(n15310), .dinb(n15104), .dout(n15311));
  jxor g15053(.dina(n15311), .dinb(n15091), .dout(n15312));
  jor  g15054(.dina(n15058), .dinb(n15050), .dout(n15313));
  jand g15055(.dina(n15059), .dinb(n15046), .dout(n15314));
  jnot g15056(.din(n15314), .dout(n15315));
  jand g15057(.dina(n15315), .dinb(n15313), .dout(n15316));
  jor  g15058(.dina(n10961), .dinb(n1245), .dout(n15317));
  jor  g15059(.dina(n1165), .dinb(n10314), .dout(n15318));
  jor  g15060(.dina(n1248), .dinb(n10637), .dout(n15319));
  jor  g15061(.dina(n1250), .dinb(n10964), .dout(n15320));
  jand g15062(.dina(n15320), .dinb(n15319), .dout(n15321));
  jand g15063(.dina(n15321), .dinb(n15318), .dout(n15322));
  jand g15064(.dina(n15322), .dinb(n15317), .dout(n15323));
  jxor g15065(.dina(n15323), .dinb(a17 ), .dout(n15324));
  jxor g15066(.dina(n15324), .dinb(n15316), .dout(n15325));
  jxor g15067(.dina(n15325), .dinb(n15312), .dout(n15326));
  jxor g15068(.dina(n15326), .dinb(n15078), .dout(n15327));
  jand g15069(.dina(n15071), .dinb(n14816), .dout(n15328));
  jand g15070(.dina(n15072), .dinb(n14811), .dout(n15329));
  jor  g15071(.dina(n15329), .dinb(n15328), .dout(n15330));
  jxor g15072(.dina(n15330), .dinb(n15327), .dout(f78 ));
  jor  g15073(.dina(n15324), .dinb(n15316), .dout(n15332));
  jand g15074(.dina(n15325), .dinb(n15312), .dout(n15333));
  jnot g15075(.din(n15333), .dout(n15334));
  jand g15076(.dina(n15334), .dinb(n15332), .dout(n15335));
  jnot g15077(.din(n15335), .dout(n15336));
  jor  g15078(.dina(n15090), .dinb(n15086), .dout(n15337));
  jand g15079(.dina(n15311), .dinb(n15091), .dout(n15338));
  jnot g15080(.din(n15338), .dout(n15339));
  jand g15081(.dina(n15339), .dinb(n15337), .dout(n15340));
  jor  g15082(.dina(n10978), .dinb(n1245), .dout(n15341));
  jor  g15083(.dina(n1165), .dinb(n10637), .dout(n15342));
  jor  g15084(.dina(n1248), .dinb(n10964), .dout(n15343));
  jand g15085(.dina(n15343), .dinb(n15342), .dout(n15344));
  jand g15086(.dina(n15344), .dinb(n15341), .dout(n15345));
  jxor g15087(.dina(n15345), .dinb(a17 ), .dout(n15346));
  jxor g15088(.dina(n15346), .dinb(n15340), .dout(n15347));
  jor  g15089(.dina(n10311), .dinb(n1566), .dout(n15348));
  jor  g15090(.dina(n1489), .dinb(n9413), .dout(n15349));
  jor  g15091(.dina(n1569), .dinb(n9725), .dout(n15350));
  jor  g15092(.dina(n1571), .dinb(n10314), .dout(n15351));
  jand g15093(.dina(n15351), .dinb(n15350), .dout(n15352));
  jand g15094(.dina(n15352), .dinb(n15349), .dout(n15353));
  jand g15095(.dina(n15353), .dinb(n15348), .dout(n15354));
  jxor g15096(.dina(n15354), .dinb(a20 ), .dout(n15355));
  jnot g15097(.din(n15355), .dout(n15356));
  jand g15098(.dina(n15103), .dinb(n15095), .dout(n15357));
  jnot g15099(.din(n15357), .dout(n15358));
  jnot g15100(.din(n15095), .dout(n15359));
  jnot g15101(.din(n15103), .dout(n15360));
  jand g15102(.dina(n15360), .dinb(n15359), .dout(n15361));
  jor  g15103(.dina(n15310), .dinb(n15361), .dout(n15362));
  jand g15104(.dina(n15362), .dinb(n15358), .dout(n15363));
  jxor g15105(.dina(n15363), .dinb(n15356), .dout(n15364));
  jand g15106(.dina(n15119), .dinb(n15113), .dout(n15365));
  jand g15107(.dina(n15309), .dinb(n15120), .dout(n15366));
  jor  g15108(.dina(n15366), .dinb(n15365), .dout(n15367));
  jnot g15109(.din(n15367), .dout(n15368));
  jor  g15110(.dina(n9387), .dinb(n1939), .dout(n15369));
  jor  g15111(.dina(n1827), .dinb(n8789), .dout(n15370));
  jor  g15112(.dina(n1942), .dinb(n8809), .dout(n15371));
  jor  g15113(.dina(n1944), .dinb(n9390), .dout(n15372));
  jand g15114(.dina(n15372), .dinb(n15371), .dout(n15373));
  jand g15115(.dina(n15373), .dinb(n15370), .dout(n15374));
  jand g15116(.dina(n15374), .dinb(n15369), .dout(n15375));
  jxor g15117(.dina(n15375), .dinb(a23 ), .dout(n15376));
  jxor g15118(.dina(n15376), .dinb(n15368), .dout(n15377));
  jor  g15119(.dina(n8228), .dinb(n2319), .dout(n15378));
  jor  g15120(.dina(n2224), .dinb(n7683), .dout(n15379));
  jor  g15121(.dina(n2322), .dinb(n7960), .dout(n15380));
  jor  g15122(.dina(n2324), .dinb(n8231), .dout(n15381));
  jand g15123(.dina(n15381), .dinb(n15380), .dout(n15382));
  jand g15124(.dina(n15382), .dinb(n15379), .dout(n15383));
  jand g15125(.dina(n15383), .dinb(n15378), .dout(n15384));
  jxor g15126(.dina(n15384), .dinb(a26 ), .dout(n15385));
  jnot g15127(.din(n15385), .dout(n15386));
  jand g15128(.dina(n15136), .dinb(n15129), .dout(n15387));
  jand g15129(.dina(n15308), .dinb(n15137), .dout(n15388));
  jor  g15130(.dina(n15388), .dinb(n15387), .dout(n15389));
  jxor g15131(.dina(n15389), .dinb(n15386), .dout(n15390));
  jor  g15132(.dina(n6864), .dinb(n3301), .dout(n15391));
  jor  g15133(.dina(n3136), .dinb(n6352), .dout(n15392));
  jor  g15134(.dina(n3304), .dinb(n6372), .dout(n15393));
  jor  g15135(.dina(n3306), .dinb(n6867), .dout(n15394));
  jand g15136(.dina(n15394), .dinb(n15393), .dout(n15395));
  jand g15137(.dina(n15395), .dinb(n15392), .dout(n15396));
  jand g15138(.dina(n15396), .dinb(n15391), .dout(n15397));
  jxor g15139(.dina(n15397), .dinb(a32 ), .dout(n15398));
  jor  g15140(.dina(n15287), .dinb(n15279), .dout(n15399));
  jand g15141(.dina(n15292), .dinb(n15288), .dout(n15400));
  jnot g15142(.din(n15400), .dout(n15401));
  jand g15143(.dina(n15401), .dinb(n15399), .dout(n15402));
  jxor g15144(.dina(n15402), .dinb(n15398), .dout(n15403));
  jand g15145(.dina(n15276), .dinb(n15149), .dout(n15404));
  jand g15146(.dina(n15277), .dinb(n15140), .dout(n15405));
  jor  g15147(.dina(n15405), .dinb(n15404), .dout(n15406));
  jor  g15148(.dina(n15274), .dinb(n15266), .dout(n15407));
  jand g15149(.dina(n15275), .dinb(n15154), .dout(n15408));
  jnot g15150(.din(n15408), .dout(n15409));
  jand g15151(.dina(n15409), .dinb(n15407), .dout(n15410));
  jnot g15152(.din(n15410), .dout(n15411));
  jor  g15153(.dina(n5096), .dinb(n4554), .dout(n15412));
  jor  g15154(.dina(n4904), .dinb(n4340), .dout(n15413));
  jor  g15155(.dina(n5099), .dinb(n4537), .dout(n15414));
  jor  g15156(.dina(n5101), .dinb(n4557), .dout(n15415));
  jand g15157(.dina(n15415), .dinb(n15414), .dout(n15416));
  jand g15158(.dina(n15416), .dinb(n15413), .dout(n15417));
  jand g15159(.dina(n15417), .dinb(n15412), .dout(n15418));
  jxor g15160(.dina(n15418), .dinb(a41 ), .dout(n15419));
  jnot g15161(.din(n15419), .dout(n15420));
  jand g15162(.dina(n15256), .dinb(n15163), .dout(n15421));
  jand g15163(.dina(n15264), .dinb(n15257), .dout(n15422));
  jor  g15164(.dina(n15422), .dinb(n15421), .dout(n15423));
  jor  g15165(.dina(n5739), .dinb(n4137), .dout(n15424));
  jor  g15166(.dina(n5574), .dinb(n3588), .dout(n15425));
  jor  g15167(.dina(n5742), .dinb(n3942), .dout(n15426));
  jor  g15168(.dina(n5744), .dinb(n4140), .dout(n15427));
  jand g15169(.dina(n15427), .dinb(n15426), .dout(n15428));
  jand g15170(.dina(n15428), .dinb(n15425), .dout(n15429));
  jand g15171(.dina(n15429), .dinb(n15424), .dout(n15430));
  jxor g15172(.dina(n15430), .dinb(a44 ), .dout(n15431));
  jnot g15173(.din(n15431), .dout(n15432));
  jor  g15174(.dina(n15254), .dinb(n15246), .dout(n15433));
  jand g15175(.dina(n15255), .dinb(n15166), .dout(n15434));
  jnot g15176(.din(n15434), .dout(n15435));
  jand g15177(.dina(n15435), .dinb(n15433), .dout(n15436));
  jnot g15178(.din(n15436), .dout(n15437));
  jor  g15179(.dina(n15239), .dinb(n15231), .dout(n15438));
  jand g15180(.dina(n15244), .dinb(n15240), .dout(n15439));
  jnot g15181(.din(n15439), .dout(n15440));
  jand g15182(.dina(n15440), .dinb(n15438), .dout(n15441));
  jnot g15183(.din(n15441), .dout(n15442));
  jor  g15184(.dina(n8125), .dinb(n2556), .dout(n15443));
  jor  g15185(.dina(n7846), .dinb(n2148), .dout(n15444));
  jor  g15186(.dina(n8128), .dinb(n2407), .dout(n15445));
  jor  g15187(.dina(n8130), .dinb(n2559), .dout(n15446));
  jand g15188(.dina(n15446), .dinb(n15445), .dout(n15447));
  jand g15189(.dina(n15447), .dinb(n15444), .dout(n15448));
  jand g15190(.dina(n15448), .dinb(n15443), .dout(n15449));
  jxor g15191(.dina(n15449), .dinb(a53 ), .dout(n15450));
  jnot g15192(.din(n15450), .dout(n15451));
  jor  g15193(.dina(n15211), .dinb(n15203), .dout(n15452));
  jand g15194(.dina(n15216), .dinb(n15212), .dout(n15453));
  jnot g15195(.din(n15453), .dout(n15454));
  jand g15196(.dina(n15454), .dinb(n15452), .dout(n15455));
  jnot g15197(.din(n15455), .dout(n15456));
  jand g15198(.dina(n15200), .dinb(n15195), .dout(n15457));
  jand g15199(.dina(n15201), .dinb(n15186), .dout(n15458));
  jor  g15200(.dina(n15458), .dinb(n15457), .dout(n15459));
  jand g15201(.dina(n15198), .dinb(n15065), .dout(n15460));
  jand g15202(.dina(n15199), .dinb(n14675), .dout(n15461));
  jor  g15203(.dina(n15461), .dinb(n15460), .dout(n15462));
  jand g15204(.dina(n10801), .dinb(b16 ), .dout(n15463));
  jand g15205(.dina(n11107), .dinb(b15 ), .dout(n15464));
  jor  g15206(.dina(n15464), .dinb(n15463), .dout(n15465));
  jnot g15207(.din(n15465), .dout(n15466));
  jxor g15208(.dina(n15466), .dinb(n15462), .dout(n15467));
  jnot g15209(.din(n15467), .dout(n15468));
  jor  g15210(.dina(n10806), .dinb(n1397), .dout(n15469));
  jor  g15211(.dina(n10485), .dinb(n1193), .dout(n15470));
  jor  g15212(.dina(n10809), .dinb(n1290), .dout(n15471));
  jor  g15213(.dina(n10811), .dinb(n1400), .dout(n15472));
  jand g15214(.dina(n15472), .dinb(n15471), .dout(n15473));
  jand g15215(.dina(n15473), .dinb(n15470), .dout(n15474));
  jand g15216(.dina(n15474), .dinb(n15469), .dout(n15475));
  jxor g15217(.dina(n15475), .dinb(a62 ), .dout(n15476));
  jxor g15218(.dina(n15476), .dinb(n15468), .dout(n15477));
  jxor g15219(.dina(n15477), .dinb(n15459), .dout(n15478));
  jor  g15220(.dina(n9891), .dinb(n1739), .dout(n15479));
  jor  g15221(.dina(n9593), .dinb(n1420), .dout(n15480));
  jor  g15222(.dina(n9894), .dinb(n1620), .dout(n15481));
  jor  g15223(.dina(n9896), .dinb(n1742), .dout(n15482));
  jand g15224(.dina(n15482), .dinb(n15481), .dout(n15483));
  jand g15225(.dina(n15483), .dinb(n15480), .dout(n15484));
  jand g15226(.dina(n15484), .dinb(n15479), .dout(n15485));
  jxor g15227(.dina(n15485), .dinb(a59 ), .dout(n15486));
  jnot g15228(.din(n15486), .dout(n15487));
  jxor g15229(.dina(n15487), .dinb(n15478), .dout(n15488));
  jxor g15230(.dina(n15488), .dinb(n15456), .dout(n15489));
  jor  g15231(.dina(n8978), .dinb(n2007), .dout(n15490));
  jor  g15232(.dina(n8677), .dinb(n1867), .dout(n15491));
  jor  g15233(.dina(n8981), .dinb(n1887), .dout(n15492));
  jor  g15234(.dina(n8983), .dinb(n2010), .dout(n15493));
  jand g15235(.dina(n15493), .dinb(n15492), .dout(n15494));
  jand g15236(.dina(n15494), .dinb(n15491), .dout(n15495));
  jand g15237(.dina(n15495), .dinb(n15490), .dout(n15496));
  jxor g15238(.dina(n15496), .dinb(a56 ), .dout(n15497));
  jnot g15239(.din(n15497), .dout(n15498));
  jxor g15240(.dina(n15498), .dinb(n15489), .dout(n15499));
  jand g15241(.dina(n15226), .dinb(n15218), .dout(n15500));
  jnot g15242(.din(n15226), .dout(n15501));
  jand g15243(.dina(n15501), .dinb(n15217), .dout(n15502));
  jnot g15244(.din(n15502), .dout(n15503));
  jand g15245(.dina(n15503), .dinb(n15181), .dout(n15504));
  jor  g15246(.dina(n15504), .dinb(n15500), .dout(n15505));
  jnot g15247(.din(n15505), .dout(n15506));
  jxor g15248(.dina(n15506), .dinb(n15499), .dout(n15507));
  jxor g15249(.dina(n15507), .dinb(n15451), .dout(n15508));
  jnot g15250(.din(n15508), .dout(n15509));
  jor  g15251(.dina(n15228), .dinb(n15177), .dout(n15510));
  jand g15252(.dina(n15229), .dinb(n15169), .dout(n15511));
  jnot g15253(.din(n15511), .dout(n15512));
  jand g15254(.dina(n15512), .dinb(n15510), .dout(n15513));
  jxor g15255(.dina(n15513), .dinb(n15509), .dout(n15514));
  jnot g15256(.din(n15514), .dout(n15515));
  jor  g15257(.dina(n7266), .dinb(n3032), .dout(n15516));
  jor  g15258(.dina(n7021), .dinb(n2579), .dout(n15517));
  jor  g15259(.dina(n7269), .dinb(n2870), .dout(n15518));
  jor  g15260(.dina(n7271), .dinb(n3035), .dout(n15519));
  jand g15261(.dina(n15519), .dinb(n15518), .dout(n15520));
  jand g15262(.dina(n15520), .dinb(n15517), .dout(n15521));
  jand g15263(.dina(n15521), .dinb(n15516), .dout(n15522));
  jxor g15264(.dina(n15522), .dinb(a50 ), .dout(n15523));
  jxor g15265(.dina(n15523), .dinb(n15515), .dout(n15524));
  jxor g15266(.dina(n15524), .dinb(n15442), .dout(n15525));
  jnot g15267(.din(n15525), .dout(n15526));
  jor  g15268(.dina(n6490), .dinb(n3400), .dout(n15527));
  jor  g15269(.dina(n6262), .dinb(n3055), .dout(n15528));
  jor  g15270(.dina(n6493), .dinb(n3230), .dout(n15529));
  jor  g15271(.dina(n6495), .dinb(n3403), .dout(n15530));
  jand g15272(.dina(n15530), .dinb(n15529), .dout(n15531));
  jand g15273(.dina(n15531), .dinb(n15528), .dout(n15532));
  jand g15274(.dina(n15532), .dinb(n15527), .dout(n15533));
  jxor g15275(.dina(n15533), .dinb(a47 ), .dout(n15534));
  jxor g15276(.dina(n15534), .dinb(n15526), .dout(n15535));
  jxor g15277(.dina(n15535), .dinb(n15437), .dout(n15536));
  jxor g15278(.dina(n15536), .dinb(n15432), .dout(n15537));
  jxor g15279(.dina(n15537), .dinb(n15423), .dout(n15538));
  jxor g15280(.dina(n15538), .dinb(n15420), .dout(n15539));
  jxor g15281(.dina(n15539), .dinb(n15411), .dout(n15540));
  jor  g15282(.dina(n5405), .dinb(n4415), .dout(n15541));
  jor  g15283(.dina(n4272), .dinb(n4974), .dout(n15542));
  jor  g15284(.dina(n4418), .dinb(n4994), .dout(n15543));
  jor  g15285(.dina(n4420), .dinb(n5408), .dout(n15544));
  jand g15286(.dina(n15544), .dinb(n15543), .dout(n15545));
  jand g15287(.dina(n15545), .dinb(n15542), .dout(n15546));
  jand g15288(.dina(n15546), .dinb(n15541), .dout(n15547));
  jxor g15289(.dina(n15547), .dinb(a38 ), .dout(n15548));
  jnot g15290(.din(n15548), .dout(n15549));
  jxor g15291(.dina(n15549), .dinb(n15540), .dout(n15550));
  jxor g15292(.dina(n15550), .dinb(n15406), .dout(n15551));
  jor  g15293(.dina(n6103), .dinb(n3849), .dout(n15552));
  jor  g15294(.dina(n3689), .dinb(n5428), .dout(n15553));
  jor  g15295(.dina(n3852), .dinb(n5862), .dout(n15554));
  jor  g15296(.dina(n3854), .dinb(n6106), .dout(n15555));
  jand g15297(.dina(n15555), .dinb(n15554), .dout(n15556));
  jand g15298(.dina(n15556), .dinb(n15553), .dout(n15557));
  jand g15299(.dina(n15557), .dinb(n15552), .dout(n15558));
  jxor g15300(.dina(n15558), .dinb(a35 ), .dout(n15559));
  jnot g15301(.din(n15559), .dout(n15560));
  jxor g15302(.dina(n15560), .dinb(n15551), .dout(n15561));
  jxor g15303(.dina(n15561), .dinb(n15403), .dout(n15562));
  jor  g15304(.dina(n7408), .dinb(n2784), .dout(n15563));
  jor  g15305(.dina(n2661), .dinb(n7129), .dout(n15564));
  jor  g15306(.dina(n2787), .dinb(n7149), .dout(n15565));
  jor  g15307(.dina(n2789), .dinb(n7411), .dout(n15566));
  jand g15308(.dina(n15566), .dinb(n15565), .dout(n15567));
  jand g15309(.dina(n15567), .dinb(n15564), .dout(n15568));
  jand g15310(.dina(n15568), .dinb(n15563), .dout(n15569));
  jxor g15311(.dina(n15569), .dinb(a29 ), .dout(n15570));
  jnot g15312(.din(n15570), .dout(n15571));
  jand g15313(.dina(n15306), .dinb(n15302), .dout(n15572));
  jand g15314(.dina(n15307), .dinb(n15293), .dout(n15573));
  jor  g15315(.dina(n15573), .dinb(n15572), .dout(n15574));
  jxor g15316(.dina(n15574), .dinb(n15571), .dout(n15575));
  jxor g15317(.dina(n15575), .dinb(n15562), .dout(n15576));
  jxor g15318(.dina(n15576), .dinb(n15390), .dout(n15577));
  jxor g15319(.dina(n15577), .dinb(n15377), .dout(n15578));
  jxor g15320(.dina(n15578), .dinb(n15364), .dout(n15579));
  jxor g15321(.dina(n15579), .dinb(n15347), .dout(n15580));
  jxor g15322(.dina(n15580), .dinb(n15336), .dout(n15581));
  jand g15323(.dina(n15326), .dinb(n15078), .dout(n15582));
  jand g15324(.dina(n15330), .dinb(n15327), .dout(n15583));
  jor  g15325(.dina(n15583), .dinb(n15582), .dout(n15584));
  jxor g15326(.dina(n15584), .dinb(n15581), .dout(f79 ));
  jand g15327(.dina(n15580), .dinb(n15336), .dout(n15586));
  jand g15328(.dina(n15584), .dinb(n15581), .dout(n15587));
  jor  g15329(.dina(n15587), .dinb(n15586), .dout(n15588));
  jor  g15330(.dina(n10634), .dinb(n1566), .dout(n15589));
  jor  g15331(.dina(n1489), .dinb(n9725), .dout(n15590));
  jor  g15332(.dina(n1569), .dinb(n10314), .dout(n15591));
  jor  g15333(.dina(n1571), .dinb(n10637), .dout(n15592));
  jand g15334(.dina(n15592), .dinb(n15591), .dout(n15593));
  jand g15335(.dina(n15593), .dinb(n15590), .dout(n15594));
  jand g15336(.dina(n15594), .dinb(n15589), .dout(n15595));
  jxor g15337(.dina(n15595), .dinb(a20 ), .dout(n15596));
  jor  g15338(.dina(n15376), .dinb(n15368), .dout(n15597));
  jand g15339(.dina(n15577), .dinb(n15377), .dout(n15598));
  jnot g15340(.din(n15598), .dout(n15599));
  jand g15341(.dina(n15599), .dinb(n15597), .dout(n15600));
  jxor g15342(.dina(n15600), .dinb(n15596), .dout(n15601));
  jor  g15343(.dina(n8786), .dinb(n2319), .dout(n15602));
  jor  g15344(.dina(n2224), .dinb(n7960), .dout(n15603));
  jor  g15345(.dina(n2322), .dinb(n8231), .dout(n15604));
  jor  g15346(.dina(n2324), .dinb(n8789), .dout(n15605));
  jand g15347(.dina(n15605), .dinb(n15604), .dout(n15606));
  jand g15348(.dina(n15606), .dinb(n15603), .dout(n15607));
  jand g15349(.dina(n15607), .dinb(n15602), .dout(n15608));
  jxor g15350(.dina(n15608), .dinb(a26 ), .dout(n15609));
  jnot g15351(.din(n15609), .dout(n15610));
  jand g15352(.dina(n15574), .dinb(n15571), .dout(n15611));
  jand g15353(.dina(n15575), .dinb(n15562), .dout(n15612));
  jor  g15354(.dina(n15612), .dinb(n15611), .dout(n15613));
  jxor g15355(.dina(n15613), .dinb(n15610), .dout(n15614));
  jor  g15356(.dina(n7126), .dinb(n3301), .dout(n15615));
  jor  g15357(.dina(n3136), .dinb(n6372), .dout(n15616));
  jor  g15358(.dina(n3304), .dinb(n6867), .dout(n15617));
  jor  g15359(.dina(n3306), .dinb(n7129), .dout(n15618));
  jand g15360(.dina(n15618), .dinb(n15617), .dout(n15619));
  jand g15361(.dina(n15619), .dinb(n15616), .dout(n15620));
  jand g15362(.dina(n15620), .dinb(n15615), .dout(n15621));
  jxor g15363(.dina(n15621), .dinb(a32 ), .dout(n15622));
  jnot g15364(.din(n15622), .dout(n15623));
  jnot g15365(.din(n15406), .dout(n15624));
  jnot g15366(.din(n15550), .dout(n15625));
  jand g15367(.dina(n15625), .dinb(n15624), .dout(n15626));
  jnot g15368(.din(n15626), .dout(n15627));
  jand g15369(.dina(n15550), .dinb(n15406), .dout(n15628));
  jor  g15370(.dina(n15560), .dinb(n15628), .dout(n15629));
  jand g15371(.dina(n15629), .dinb(n15627), .dout(n15630));
  jxor g15372(.dina(n15630), .dinb(n15623), .dout(n15631));
  jor  g15373(.dina(n5425), .dinb(n4415), .dout(n15632));
  jor  g15374(.dina(n4272), .dinb(n4994), .dout(n15633));
  jor  g15375(.dina(n4418), .dinb(n5408), .dout(n15634));
  jor  g15376(.dina(n4420), .dinb(n5428), .dout(n15635));
  jand g15377(.dina(n15635), .dinb(n15634), .dout(n15636));
  jand g15378(.dina(n15636), .dinb(n15633), .dout(n15637));
  jand g15379(.dina(n15637), .dinb(n15632), .dout(n15638));
  jxor g15380(.dina(n15638), .dinb(a38 ), .dout(n15639));
  jnot g15381(.din(n15639), .dout(n15640));
  jand g15382(.dina(n15537), .dinb(n15423), .dout(n15641));
  jand g15383(.dina(n15538), .dinb(n15420), .dout(n15642));
  jor  g15384(.dina(n15642), .dinb(n15641), .dout(n15643));
  jor  g15385(.dina(n4971), .dinb(n5096), .dout(n15644));
  jor  g15386(.dina(n4904), .dinb(n4537), .dout(n15645));
  jor  g15387(.dina(n5099), .dinb(n4557), .dout(n15646));
  jor  g15388(.dina(n5101), .dinb(n4974), .dout(n15647));
  jand g15389(.dina(n15647), .dinb(n15646), .dout(n15648));
  jand g15390(.dina(n15648), .dinb(n15645), .dout(n15649));
  jand g15391(.dina(n15649), .dinb(n15644), .dout(n15650));
  jxor g15392(.dina(n15650), .dinb(a41 ), .dout(n15651));
  jnot g15393(.din(n15651), .dout(n15652));
  jand g15394(.dina(n15535), .dinb(n15437), .dout(n15653));
  jand g15395(.dina(n15536), .dinb(n15432), .dout(n15654));
  jor  g15396(.dina(n15654), .dinb(n15653), .dout(n15655));
  jor  g15397(.dina(n5739), .dinb(n4337), .dout(n15656));
  jor  g15398(.dina(n5574), .dinb(n3942), .dout(n15657));
  jor  g15399(.dina(n5742), .dinb(n4140), .dout(n15658));
  jor  g15400(.dina(n5744), .dinb(n4340), .dout(n15659));
  jand g15401(.dina(n15659), .dinb(n15658), .dout(n15660));
  jand g15402(.dina(n15660), .dinb(n15657), .dout(n15661));
  jand g15403(.dina(n15661), .dinb(n15656), .dout(n15662));
  jxor g15404(.dina(n15662), .dinb(a44 ), .dout(n15663));
  jnot g15405(.din(n15663), .dout(n15664));
  jand g15406(.dina(n15524), .dinb(n15442), .dout(n15665));
  jnot g15407(.din(n15665), .dout(n15666));
  jor  g15408(.dina(n15534), .dinb(n15526), .dout(n15667));
  jand g15409(.dina(n15667), .dinb(n15666), .dout(n15668));
  jnot g15410(.din(n15668), .dout(n15669));
  jor  g15411(.dina(n7266), .dinb(n3052), .dout(n15670));
  jor  g15412(.dina(n7021), .dinb(n2870), .dout(n15671));
  jor  g15413(.dina(n7269), .dinb(n3035), .dout(n15672));
  jor  g15414(.dina(n7271), .dinb(n3055), .dout(n15673));
  jand g15415(.dina(n15673), .dinb(n15672), .dout(n15674));
  jand g15416(.dina(n15674), .dinb(n15671), .dout(n15675));
  jand g15417(.dina(n15675), .dinb(n15670), .dout(n15676));
  jxor g15418(.dina(n15676), .dinb(a50 ), .dout(n15677));
  jnot g15419(.din(n15677), .dout(n15678));
  jand g15420(.dina(n15506), .dinb(n15499), .dout(n15679));
  jand g15421(.dina(n15507), .dinb(n15451), .dout(n15680));
  jor  g15422(.dina(n15680), .dinb(n15679), .dout(n15681));
  jor  g15423(.dina(n8978), .dinb(n2145), .dout(n15682));
  jor  g15424(.dina(n8677), .dinb(n1887), .dout(n15683));
  jor  g15425(.dina(n8981), .dinb(n2010), .dout(n15684));
  jor  g15426(.dina(n8983), .dinb(n2148), .dout(n15685));
  jand g15427(.dina(n15685), .dinb(n15684), .dout(n15686));
  jand g15428(.dina(n15686), .dinb(n15683), .dout(n15687));
  jand g15429(.dina(n15687), .dinb(n15682), .dout(n15688));
  jxor g15430(.dina(n15688), .dinb(a56 ), .dout(n15689));
  jnot g15431(.din(n15689), .dout(n15690));
  jand g15432(.dina(n15466), .dinb(n15462), .dout(n15691));
  jnot g15433(.din(n15691), .dout(n15692));
  jor  g15434(.dina(n15476), .dinb(n15468), .dout(n15693));
  jand g15435(.dina(n15693), .dinb(n15692), .dout(n15694));
  jnot g15436(.din(n15694), .dout(n15695));
  jor  g15437(.dina(n10806), .dinb(n1417), .dout(n15696));
  jor  g15438(.dina(n10485), .dinb(n1290), .dout(n15697));
  jor  g15439(.dina(n10809), .dinb(n1400), .dout(n15698));
  jor  g15440(.dina(n10811), .dinb(n1420), .dout(n15699));
  jand g15441(.dina(n15699), .dinb(n15698), .dout(n15700));
  jand g15442(.dina(n15700), .dinb(n15697), .dout(n15701));
  jand g15443(.dina(n15701), .dinb(n15696), .dout(n15702));
  jxor g15444(.dina(n15702), .dinb(a62 ), .dout(n15703));
  jnot g15445(.din(n15703), .dout(n15704));
  jand g15446(.dina(n10801), .dinb(b17 ), .dout(n15705));
  jand g15447(.dina(n11107), .dinb(b16 ), .dout(n15706));
  jor  g15448(.dina(n15706), .dinb(n15705), .dout(n15707));
  jnot g15449(.din(n15707), .dout(n15708));
  jxor g15450(.dina(n15708), .dinb(n15465), .dout(n15709));
  jxor g15451(.dina(n15709), .dinb(n15704), .dout(n15710));
  jxor g15452(.dina(n15710), .dinb(n15695), .dout(n15711));
  jnot g15453(.din(n15711), .dout(n15712));
  jor  g15454(.dina(n9891), .dinb(n1864), .dout(n15713));
  jor  g15455(.dina(n9593), .dinb(n1620), .dout(n15714));
  jor  g15456(.dina(n9894), .dinb(n1742), .dout(n15715));
  jor  g15457(.dina(n9896), .dinb(n1867), .dout(n15716));
  jand g15458(.dina(n15716), .dinb(n15715), .dout(n15717));
  jand g15459(.dina(n15717), .dinb(n15714), .dout(n15718));
  jand g15460(.dina(n15718), .dinb(n15713), .dout(n15719));
  jxor g15461(.dina(n15719), .dinb(a59 ), .dout(n15720));
  jxor g15462(.dina(n15720), .dinb(n15712), .dout(n15721));
  jor  g15463(.dina(n15477), .dinb(n15459), .dout(n15722));
  jand g15464(.dina(n15477), .dinb(n15459), .dout(n15723));
  jor  g15465(.dina(n15487), .dinb(n15723), .dout(n15724));
  jand g15466(.dina(n15724), .dinb(n15722), .dout(n15725));
  jxor g15467(.dina(n15725), .dinb(n15721), .dout(n15726));
  jxor g15468(.dina(n15726), .dinb(n15690), .dout(n15727));
  jnot g15469(.din(n15488), .dout(n15728));
  jand g15470(.dina(n15728), .dinb(n15455), .dout(n15729));
  jnot g15471(.din(n15729), .dout(n15730));
  jand g15472(.dina(n15488), .dinb(n15456), .dout(n15731));
  jor  g15473(.dina(n15498), .dinb(n15731), .dout(n15732));
  jand g15474(.dina(n15732), .dinb(n15730), .dout(n15733));
  jxor g15475(.dina(n15733), .dinb(n15727), .dout(n15734));
  jor  g15476(.dina(n8125), .dinb(n2576), .dout(n15735));
  jor  g15477(.dina(n7846), .dinb(n2407), .dout(n15736));
  jor  g15478(.dina(n8128), .dinb(n2559), .dout(n15737));
  jor  g15479(.dina(n8130), .dinb(n2579), .dout(n15738));
  jand g15480(.dina(n15738), .dinb(n15737), .dout(n15739));
  jand g15481(.dina(n15739), .dinb(n15736), .dout(n15740));
  jand g15482(.dina(n15740), .dinb(n15735), .dout(n15741));
  jxor g15483(.dina(n15741), .dinb(a53 ), .dout(n15742));
  jnot g15484(.din(n15742), .dout(n15743));
  jxor g15485(.dina(n15743), .dinb(n15734), .dout(n15744));
  jxor g15486(.dina(n15744), .dinb(n15681), .dout(n15745));
  jxor g15487(.dina(n15745), .dinb(n15678), .dout(n15746));
  jnot g15488(.din(n15746), .dout(n15747));
  jnot g15489(.din(n15513), .dout(n15748));
  jand g15490(.dina(n15748), .dinb(n15508), .dout(n15749));
  jnot g15491(.din(n15749), .dout(n15750));
  jand g15492(.dina(n15513), .dinb(n15509), .dout(n15751));
  jor  g15493(.dina(n15523), .dinb(n15751), .dout(n15752));
  jand g15494(.dina(n15752), .dinb(n15750), .dout(n15753));
  jxor g15495(.dina(n15753), .dinb(n15747), .dout(n15754));
  jnot g15496(.din(n15754), .dout(n15755));
  jor  g15497(.dina(n6490), .dinb(n3585), .dout(n15756));
  jor  g15498(.dina(n6262), .dinb(n3230), .dout(n15757));
  jor  g15499(.dina(n6493), .dinb(n3403), .dout(n15758));
  jor  g15500(.dina(n6495), .dinb(n3588), .dout(n15759));
  jand g15501(.dina(n15759), .dinb(n15758), .dout(n15760));
  jand g15502(.dina(n15760), .dinb(n15757), .dout(n15761));
  jand g15503(.dina(n15761), .dinb(n15756), .dout(n15762));
  jxor g15504(.dina(n15762), .dinb(a47 ), .dout(n15763));
  jxor g15505(.dina(n15763), .dinb(n15755), .dout(n15764));
  jxor g15506(.dina(n15764), .dinb(n15669), .dout(n15765));
  jxor g15507(.dina(n15765), .dinb(n15664), .dout(n15766));
  jxor g15508(.dina(n15766), .dinb(n15655), .dout(n15767));
  jxor g15509(.dina(n15767), .dinb(n15652), .dout(n15768));
  jxor g15510(.dina(n15768), .dinb(n15643), .dout(n15769));
  jxor g15511(.dina(n15769), .dinb(n15640), .dout(n15770));
  jor  g15512(.dina(n15539), .dinb(n15411), .dout(n15771));
  jand g15513(.dina(n15539), .dinb(n15411), .dout(n15772));
  jor  g15514(.dina(n15549), .dinb(n15772), .dout(n15773));
  jand g15515(.dina(n15773), .dinb(n15771), .dout(n15774));
  jxor g15516(.dina(n15774), .dinb(n15770), .dout(n15775));
  jor  g15517(.dina(n6349), .dinb(n3849), .dout(n15776));
  jor  g15518(.dina(n3689), .dinb(n5862), .dout(n15777));
  jor  g15519(.dina(n3852), .dinb(n6106), .dout(n15778));
  jor  g15520(.dina(n3854), .dinb(n6352), .dout(n15779));
  jand g15521(.dina(n15779), .dinb(n15778), .dout(n15780));
  jand g15522(.dina(n15780), .dinb(n15777), .dout(n15781));
  jand g15523(.dina(n15781), .dinb(n15776), .dout(n15782));
  jxor g15524(.dina(n15782), .dinb(a35 ), .dout(n15783));
  jnot g15525(.din(n15783), .dout(n15784));
  jxor g15526(.dina(n15784), .dinb(n15775), .dout(n15785));
  jxor g15527(.dina(n15785), .dinb(n15631), .dout(n15786));
  jor  g15528(.dina(n7680), .dinb(n2784), .dout(n15787));
  jor  g15529(.dina(n2661), .dinb(n7149), .dout(n15788));
  jor  g15530(.dina(n2787), .dinb(n7411), .dout(n15789));
  jor  g15531(.dina(n2789), .dinb(n7683), .dout(n15790));
  jand g15532(.dina(n15790), .dinb(n15789), .dout(n15791));
  jand g15533(.dina(n15791), .dinb(n15788), .dout(n15792));
  jand g15534(.dina(n15792), .dinb(n15787), .dout(n15793));
  jxor g15535(.dina(n15793), .dinb(a29 ), .dout(n15794));
  jor  g15536(.dina(n15402), .dinb(n15398), .dout(n15795));
  jand g15537(.dina(n15561), .dinb(n15403), .dout(n15796));
  jnot g15538(.din(n15796), .dout(n15797));
  jand g15539(.dina(n15797), .dinb(n15795), .dout(n15798));
  jxor g15540(.dina(n15798), .dinb(n15794), .dout(n15799));
  jxor g15541(.dina(n15799), .dinb(n15786), .dout(n15800));
  jxor g15542(.dina(n15800), .dinb(n15614), .dout(n15801));
  jor  g15543(.dina(n9410), .dinb(n1939), .dout(n15802));
  jor  g15544(.dina(n1827), .dinb(n8809), .dout(n15803));
  jor  g15545(.dina(n1942), .dinb(n9390), .dout(n15804));
  jor  g15546(.dina(n1944), .dinb(n9413), .dout(n15805));
  jand g15547(.dina(n15805), .dinb(n15804), .dout(n15806));
  jand g15548(.dina(n15806), .dinb(n15803), .dout(n15807));
  jand g15549(.dina(n15807), .dinb(n15802), .dout(n15808));
  jxor g15550(.dina(n15808), .dinb(a23 ), .dout(n15809));
  jnot g15551(.din(n15809), .dout(n15810));
  jand g15552(.dina(n15389), .dinb(n15386), .dout(n15811));
  jand g15553(.dina(n15576), .dinb(n15390), .dout(n15812));
  jor  g15554(.dina(n15812), .dinb(n15811), .dout(n15813));
  jxor g15555(.dina(n15813), .dinb(n15810), .dout(n15814));
  jxor g15556(.dina(n15814), .dinb(n15801), .dout(n15815));
  jxor g15557(.dina(n15815), .dinb(n15601), .dout(n15816));
  jand g15558(.dina(n15363), .dinb(n15356), .dout(n15817));
  jand g15559(.dina(n15578), .dinb(n15364), .dout(n15818));
  jor  g15560(.dina(n15818), .dinb(n15817), .dout(n15819));
  jnot g15561(.din(n15819), .dout(n15820));
  jnot g15562(.din(a17 ), .dout(n15821));
  jand g15563(.dina(n11296), .dinb(n1090), .dout(n15822));
  jor  g15564(.dina(n15822), .dinb(n1166), .dout(n15823));
  jand g15565(.dina(n15823), .dinb(b63 ), .dout(n15824));
  jxor g15566(.dina(n15824), .dinb(n15821), .dout(n15825));
  jxor g15567(.dina(n15825), .dinb(n15820), .dout(n15826));
  jxor g15568(.dina(n15826), .dinb(n15816), .dout(n15827));
  jand g15569(.dina(n15346), .dinb(n15340), .dout(n15828));
  jnot g15570(.din(n15828), .dout(n15829));
  jnot g15571(.din(n15340), .dout(n15830));
  jnot g15572(.din(n15346), .dout(n15831));
  jand g15573(.dina(n15831), .dinb(n15830), .dout(n15832));
  jor  g15574(.dina(n15579), .dinb(n15832), .dout(n15833));
  jand g15575(.dina(n15833), .dinb(n15829), .dout(n15834));
  jxor g15576(.dina(n15834), .dinb(n15827), .dout(n15835));
  jxor g15577(.dina(n15835), .dinb(n15588), .dout(f80 ));
  jand g15578(.dina(n15834), .dinb(n15827), .dout(n15837));
  jand g15579(.dina(n15835), .dinb(n15588), .dout(n15838));
  jor  g15580(.dina(n15838), .dinb(n15837), .dout(n15839));
  jor  g15581(.dina(n15825), .dinb(n15820), .dout(n15840));
  jand g15582(.dina(n15826), .dinb(n15816), .dout(n15841));
  jnot g15583(.din(n15841), .dout(n15842));
  jand g15584(.dina(n15842), .dinb(n15840), .dout(n15843));
  jnot g15585(.din(n15843), .dout(n15844));
  jor  g15586(.dina(n15600), .dinb(n15596), .dout(n15845));
  jand g15587(.dina(n15815), .dinb(n15601), .dout(n15846));
  jnot g15588(.din(n15846), .dout(n15847));
  jand g15589(.dina(n15847), .dinb(n15845), .dout(n15848));
  jor  g15590(.dina(n10961), .dinb(n1566), .dout(n15849));
  jor  g15591(.dina(n1489), .dinb(n10314), .dout(n15850));
  jor  g15592(.dina(n1569), .dinb(n10637), .dout(n15851));
  jor  g15593(.dina(n1571), .dinb(n10964), .dout(n15852));
  jand g15594(.dina(n15852), .dinb(n15851), .dout(n15853));
  jand g15595(.dina(n15853), .dinb(n15850), .dout(n15854));
  jand g15596(.dina(n15854), .dinb(n15849), .dout(n15855));
  jxor g15597(.dina(n15855), .dinb(a20 ), .dout(n15856));
  jxor g15598(.dina(n15856), .dinb(n15848), .dout(n15857));
  jor  g15599(.dina(n9722), .dinb(n1939), .dout(n15858));
  jor  g15600(.dina(n1827), .dinb(n9390), .dout(n15859));
  jor  g15601(.dina(n1942), .dinb(n9413), .dout(n15860));
  jor  g15602(.dina(n1944), .dinb(n9725), .dout(n15861));
  jand g15603(.dina(n15861), .dinb(n15860), .dout(n15862));
  jand g15604(.dina(n15862), .dinb(n15859), .dout(n15863));
  jand g15605(.dina(n15863), .dinb(n15858), .dout(n15864));
  jxor g15606(.dina(n15864), .dinb(a23 ), .dout(n15865));
  jnot g15607(.din(n15865), .dout(n15866));
  jand g15608(.dina(n15813), .dinb(n15810), .dout(n15867));
  jand g15609(.dina(n15814), .dinb(n15801), .dout(n15868));
  jor  g15610(.dina(n15868), .dinb(n15867), .dout(n15869));
  jxor g15611(.dina(n15869), .dinb(n15866), .dout(n15870));
  jor  g15612(.dina(n7957), .dinb(n2784), .dout(n15871));
  jor  g15613(.dina(n2661), .dinb(n7411), .dout(n15872));
  jor  g15614(.dina(n2787), .dinb(n7683), .dout(n15873));
  jor  g15615(.dina(n2789), .dinb(n7960), .dout(n15874));
  jand g15616(.dina(n15874), .dinb(n15873), .dout(n15875));
  jand g15617(.dina(n15875), .dinb(n15872), .dout(n15876));
  jand g15618(.dina(n15876), .dinb(n15871), .dout(n15877));
  jxor g15619(.dina(n15877), .dinb(a29 ), .dout(n15878));
  jor  g15620(.dina(n15798), .dinb(n15794), .dout(n15879));
  jand g15621(.dina(n15799), .dinb(n15786), .dout(n15880));
  jnot g15622(.din(n15880), .dout(n15881));
  jand g15623(.dina(n15881), .dinb(n15879), .dout(n15882));
  jxor g15624(.dina(n15882), .dinb(n15878), .dout(n15883));
  jand g15625(.dina(n15768), .dinb(n15643), .dout(n15884));
  jand g15626(.dina(n15769), .dinb(n15640), .dout(n15885));
  jor  g15627(.dina(n15885), .dinb(n15884), .dout(n15886));
  jand g15628(.dina(n15766), .dinb(n15655), .dout(n15887));
  jand g15629(.dina(n15767), .dinb(n15652), .dout(n15888));
  jor  g15630(.dina(n15888), .dinb(n15887), .dout(n15889));
  jor  g15631(.dina(n4991), .dinb(n5096), .dout(n15890));
  jor  g15632(.dina(n4904), .dinb(n4557), .dout(n15891));
  jor  g15633(.dina(n5099), .dinb(n4974), .dout(n15892));
  jor  g15634(.dina(n5101), .dinb(n4994), .dout(n15893));
  jand g15635(.dina(n15893), .dinb(n15892), .dout(n15894));
  jand g15636(.dina(n15894), .dinb(n15891), .dout(n15895));
  jand g15637(.dina(n15895), .dinb(n15890), .dout(n15896));
  jxor g15638(.dina(n15896), .dinb(a41 ), .dout(n15897));
  jnot g15639(.din(n15897), .dout(n15898));
  jand g15640(.dina(n15764), .dinb(n15669), .dout(n15899));
  jand g15641(.dina(n15765), .dinb(n15664), .dout(n15900));
  jor  g15642(.dina(n15900), .dinb(n15899), .dout(n15901));
  jor  g15643(.dina(n6490), .dinb(n3939), .dout(n15902));
  jor  g15644(.dina(n6262), .dinb(n3403), .dout(n15903));
  jor  g15645(.dina(n6493), .dinb(n3588), .dout(n15904));
  jor  g15646(.dina(n6495), .dinb(n3942), .dout(n15905));
  jand g15647(.dina(n15905), .dinb(n15904), .dout(n15906));
  jand g15648(.dina(n15906), .dinb(n15903), .dout(n15907));
  jand g15649(.dina(n15907), .dinb(n15902), .dout(n15908));
  jxor g15650(.dina(n15908), .dinb(a47 ), .dout(n15909));
  jnot g15651(.din(n15909), .dout(n15910));
  jand g15652(.dina(n15725), .dinb(n15721), .dout(n15911));
  jand g15653(.dina(n15726), .dinb(n15690), .dout(n15912));
  jor  g15654(.dina(n15912), .dinb(n15911), .dout(n15913));
  jand g15655(.dina(n15710), .dinb(n15695), .dout(n15914));
  jnot g15656(.din(n15914), .dout(n15915));
  jor  g15657(.dina(n15720), .dinb(n15712), .dout(n15916));
  jand g15658(.dina(n15916), .dinb(n15915), .dout(n15917));
  jnot g15659(.din(n15917), .dout(n15918));
  jor  g15660(.dina(n9891), .dinb(n1884), .dout(n15919));
  jor  g15661(.dina(n9593), .dinb(n1742), .dout(n15920));
  jor  g15662(.dina(n9894), .dinb(n1867), .dout(n15921));
  jor  g15663(.dina(n9896), .dinb(n1887), .dout(n15922));
  jand g15664(.dina(n15922), .dinb(n15921), .dout(n15923));
  jand g15665(.dina(n15923), .dinb(n15920), .dout(n15924));
  jand g15666(.dina(n15924), .dinb(n15919), .dout(n15925));
  jxor g15667(.dina(n15925), .dinb(a59 ), .dout(n15926));
  jnot g15668(.din(n15926), .dout(n15927));
  jand g15669(.dina(n15708), .dinb(n15465), .dout(n15928));
  jand g15670(.dina(n15709), .dinb(n15704), .dout(n15929));
  jor  g15671(.dina(n15929), .dinb(n15928), .dout(n15930));
  jor  g15672(.dina(n10806), .dinb(n1617), .dout(n15931));
  jor  g15673(.dina(n10485), .dinb(n1400), .dout(n15932));
  jor  g15674(.dina(n10809), .dinb(n1420), .dout(n15933));
  jor  g15675(.dina(n10811), .dinb(n1620), .dout(n15934));
  jand g15676(.dina(n15934), .dinb(n15933), .dout(n15935));
  jand g15677(.dina(n15935), .dinb(n15932), .dout(n15936));
  jand g15678(.dina(n15936), .dinb(n15931), .dout(n15937));
  jxor g15679(.dina(n15937), .dinb(a62 ), .dout(n15938));
  jnot g15680(.din(n15938), .dout(n15939));
  jand g15681(.dina(n10801), .dinb(b18 ), .dout(n15940));
  jand g15682(.dina(n11107), .dinb(b17 ), .dout(n15941));
  jor  g15683(.dina(n15941), .dinb(n15940), .dout(n15942));
  jxor g15684(.dina(n15942), .dinb(n15821), .dout(n15943));
  jxor g15685(.dina(n15943), .dinb(n15707), .dout(n15944));
  jxor g15686(.dina(n15944), .dinb(n15939), .dout(n15945));
  jxor g15687(.dina(n15945), .dinb(n15930), .dout(n15946));
  jxor g15688(.dina(n15946), .dinb(n15927), .dout(n15947));
  jxor g15689(.dina(n15947), .dinb(n15918), .dout(n15948));
  jnot g15690(.din(n15948), .dout(n15949));
  jor  g15691(.dina(n8978), .dinb(n2404), .dout(n15950));
  jor  g15692(.dina(n8677), .dinb(n2010), .dout(n15951));
  jor  g15693(.dina(n8981), .dinb(n2148), .dout(n15952));
  jor  g15694(.dina(n8983), .dinb(n2407), .dout(n15953));
  jand g15695(.dina(n15953), .dinb(n15952), .dout(n15954));
  jand g15696(.dina(n15954), .dinb(n15951), .dout(n15955));
  jand g15697(.dina(n15955), .dinb(n15950), .dout(n15956));
  jxor g15698(.dina(n15956), .dinb(a56 ), .dout(n15957));
  jxor g15699(.dina(n15957), .dinb(n15949), .dout(n15958));
  jxor g15700(.dina(n15958), .dinb(n15913), .dout(n15959));
  jnot g15701(.din(n15959), .dout(n15960));
  jor  g15702(.dina(n8125), .dinb(n2867), .dout(n15961));
  jor  g15703(.dina(n7846), .dinb(n2559), .dout(n15962));
  jor  g15704(.dina(n8128), .dinb(n2579), .dout(n15963));
  jor  g15705(.dina(n8130), .dinb(n2870), .dout(n15964));
  jand g15706(.dina(n15964), .dinb(n15963), .dout(n15965));
  jand g15707(.dina(n15965), .dinb(n15962), .dout(n15966));
  jand g15708(.dina(n15966), .dinb(n15961), .dout(n15967));
  jxor g15709(.dina(n15967), .dinb(a53 ), .dout(n15968));
  jxor g15710(.dina(n15968), .dinb(n15960), .dout(n15969));
  jor  g15711(.dina(n15733), .dinb(n15727), .dout(n15970));
  jand g15712(.dina(n15733), .dinb(n15727), .dout(n15971));
  jor  g15713(.dina(n15743), .dinb(n15971), .dout(n15972));
  jand g15714(.dina(n15972), .dinb(n15970), .dout(n15973));
  jxor g15715(.dina(n15973), .dinb(n15969), .dout(n15974));
  jor  g15716(.dina(n7266), .dinb(n3227), .dout(n15975));
  jor  g15717(.dina(n7021), .dinb(n3035), .dout(n15976));
  jor  g15718(.dina(n7269), .dinb(n3055), .dout(n15977));
  jor  g15719(.dina(n7271), .dinb(n3230), .dout(n15978));
  jand g15720(.dina(n15978), .dinb(n15977), .dout(n15979));
  jand g15721(.dina(n15979), .dinb(n15976), .dout(n15980));
  jand g15722(.dina(n15980), .dinb(n15975), .dout(n15981));
  jxor g15723(.dina(n15981), .dinb(a50 ), .dout(n15982));
  jnot g15724(.din(n15982), .dout(n15983));
  jand g15725(.dina(n15744), .dinb(n15681), .dout(n15984));
  jand g15726(.dina(n15745), .dinb(n15678), .dout(n15985));
  jor  g15727(.dina(n15985), .dinb(n15984), .dout(n15986));
  jxor g15728(.dina(n15986), .dinb(n15983), .dout(n15987));
  jxor g15729(.dina(n15987), .dinb(n15974), .dout(n15988));
  jxor g15730(.dina(n15988), .dinb(n15910), .dout(n15989));
  jnot g15731(.din(n15989), .dout(n15990));
  jor  g15732(.dina(n15753), .dinb(n15747), .dout(n15991));
  jand g15733(.dina(n15753), .dinb(n15747), .dout(n15992));
  jor  g15734(.dina(n15763), .dinb(n15992), .dout(n15993));
  jand g15735(.dina(n15993), .dinb(n15991), .dout(n15994));
  jxor g15736(.dina(n15994), .dinb(n15990), .dout(n15995));
  jnot g15737(.din(n15995), .dout(n15996));
  jor  g15738(.dina(n5739), .dinb(n4534), .dout(n15997));
  jor  g15739(.dina(n5574), .dinb(n4140), .dout(n15998));
  jor  g15740(.dina(n5742), .dinb(n4340), .dout(n15999));
  jor  g15741(.dina(n5744), .dinb(n4537), .dout(n16000));
  jand g15742(.dina(n16000), .dinb(n15999), .dout(n16001));
  jand g15743(.dina(n16001), .dinb(n15998), .dout(n16002));
  jand g15744(.dina(n16002), .dinb(n15997), .dout(n16003));
  jxor g15745(.dina(n16003), .dinb(a44 ), .dout(n16004));
  jxor g15746(.dina(n16004), .dinb(n15996), .dout(n16005));
  jxor g15747(.dina(n16005), .dinb(n15901), .dout(n16006));
  jxor g15748(.dina(n16006), .dinb(n15898), .dout(n16007));
  jxor g15749(.dina(n16007), .dinb(n15889), .dout(n16008));
  jnot g15750(.din(n16008), .dout(n16009));
  jor  g15751(.dina(n5859), .dinb(n4415), .dout(n16010));
  jor  g15752(.dina(n4272), .dinb(n5408), .dout(n16011));
  jor  g15753(.dina(n4418), .dinb(n5428), .dout(n16012));
  jor  g15754(.dina(n4420), .dinb(n5862), .dout(n16013));
  jand g15755(.dina(n16013), .dinb(n16012), .dout(n16014));
  jand g15756(.dina(n16014), .dinb(n16011), .dout(n16015));
  jand g15757(.dina(n16015), .dinb(n16010), .dout(n16016));
  jxor g15758(.dina(n16016), .dinb(a38 ), .dout(n16017));
  jxor g15759(.dina(n16017), .dinb(n16009), .dout(n16018));
  jxor g15760(.dina(n16018), .dinb(n15886), .dout(n16019));
  jnot g15761(.din(n16019), .dout(n16020));
  jor  g15762(.dina(n6369), .dinb(n3849), .dout(n16021));
  jor  g15763(.dina(n3689), .dinb(n6106), .dout(n16022));
  jor  g15764(.dina(n3852), .dinb(n6352), .dout(n16023));
  jor  g15765(.dina(n3854), .dinb(n6372), .dout(n16024));
  jand g15766(.dina(n16024), .dinb(n16023), .dout(n16025));
  jand g15767(.dina(n16025), .dinb(n16022), .dout(n16026));
  jand g15768(.dina(n16026), .dinb(n16021), .dout(n16027));
  jxor g15769(.dina(n16027), .dinb(a35 ), .dout(n16028));
  jxor g15770(.dina(n16028), .dinb(n16020), .dout(n16029));
  jor  g15771(.dina(n15774), .dinb(n15770), .dout(n16030));
  jand g15772(.dina(n15774), .dinb(n15770), .dout(n16031));
  jor  g15773(.dina(n15784), .dinb(n16031), .dout(n16032));
  jand g15774(.dina(n16032), .dinb(n16030), .dout(n16033));
  jxor g15775(.dina(n16033), .dinb(n16029), .dout(n16034));
  jor  g15776(.dina(n7146), .dinb(n3301), .dout(n16035));
  jor  g15777(.dina(n3136), .dinb(n6867), .dout(n16036));
  jor  g15778(.dina(n3304), .dinb(n7129), .dout(n16037));
  jor  g15779(.dina(n3306), .dinb(n7149), .dout(n16038));
  jand g15780(.dina(n16038), .dinb(n16037), .dout(n16039));
  jand g15781(.dina(n16039), .dinb(n16036), .dout(n16040));
  jand g15782(.dina(n16040), .dinb(n16035), .dout(n16041));
  jxor g15783(.dina(n16041), .dinb(a32 ), .dout(n16042));
  jnot g15784(.din(n16042), .dout(n16043));
  jand g15785(.dina(n15630), .dinb(n15623), .dout(n16044));
  jand g15786(.dina(n15785), .dinb(n15631), .dout(n16045));
  jor  g15787(.dina(n16045), .dinb(n16044), .dout(n16046));
  jxor g15788(.dina(n16046), .dinb(n16043), .dout(n16047));
  jxor g15789(.dina(n16047), .dinb(n16034), .dout(n16048));
  jnot g15790(.din(n16048), .dout(n16049));
  jxor g15791(.dina(n16049), .dinb(n15883), .dout(n16050));
  jnot g15792(.din(n16050), .dout(n16051));
  jor  g15793(.dina(n8806), .dinb(n2319), .dout(n16052));
  jor  g15794(.dina(n2224), .dinb(n8231), .dout(n16053));
  jor  g15795(.dina(n2322), .dinb(n8789), .dout(n16054));
  jor  g15796(.dina(n2324), .dinb(n8809), .dout(n16055));
  jand g15797(.dina(n16055), .dinb(n16054), .dout(n16056));
  jand g15798(.dina(n16056), .dinb(n16053), .dout(n16057));
  jand g15799(.dina(n16057), .dinb(n16052), .dout(n16058));
  jxor g15800(.dina(n16058), .dinb(a26 ), .dout(n16059));
  jnot g15801(.din(n16059), .dout(n16060));
  jand g15802(.dina(n15613), .dinb(n15610), .dout(n16061));
  jand g15803(.dina(n15800), .dinb(n15614), .dout(n16062));
  jor  g15804(.dina(n16062), .dinb(n16061), .dout(n16063));
  jxor g15805(.dina(n16063), .dinb(n16060), .dout(n16064));
  jxor g15806(.dina(n16064), .dinb(n16051), .dout(n16065));
  jxor g15807(.dina(n16065), .dinb(n15870), .dout(n16066));
  jxor g15808(.dina(n16066), .dinb(n15857), .dout(n16067));
  jxor g15809(.dina(n16067), .dinb(n15844), .dout(n16068));
  jxor g15810(.dina(n16068), .dinb(n15839), .dout(f81 ));
  jand g15811(.dina(n16067), .dinb(n15844), .dout(n16070));
  jand g15812(.dina(n16068), .dinb(n15839), .dout(n16071));
  jor  g15813(.dina(n16071), .dinb(n16070), .dout(n16072));
  jor  g15814(.dina(n15856), .dinb(n15848), .dout(n16073));
  jand g15815(.dina(n16066), .dinb(n15857), .dout(n16074));
  jnot g15816(.din(n16074), .dout(n16075));
  jand g15817(.dina(n16075), .dinb(n16073), .dout(n16076));
  jnot g15818(.din(n16076), .dout(n16077));
  jor  g15819(.dina(n10978), .dinb(n1566), .dout(n16078));
  jor  g15820(.dina(n1489), .dinb(n10637), .dout(n16079));
  jor  g15821(.dina(n1569), .dinb(n10964), .dout(n16080));
  jand g15822(.dina(n16080), .dinb(n16079), .dout(n16081));
  jand g15823(.dina(n16081), .dinb(n16078), .dout(n16082));
  jxor g15824(.dina(n16082), .dinb(a20 ), .dout(n16083));
  jnot g15825(.din(n16083), .dout(n16084));
  jnot g15826(.din(n15869), .dout(n16085));
  jand g15827(.dina(n16085), .dinb(n15865), .dout(n16086));
  jnot g15828(.din(n16086), .dout(n16087));
  jand g15829(.dina(n15869), .dinb(n15866), .dout(n16088));
  jor  g15830(.dina(n16065), .dinb(n16088), .dout(n16089));
  jand g15831(.dina(n16089), .dinb(n16087), .dout(n16090));
  jxor g15832(.dina(n16090), .dinb(n16084), .dout(n16091));
  jor  g15833(.dina(n10311), .dinb(n1939), .dout(n16092));
  jor  g15834(.dina(n1827), .dinb(n9413), .dout(n16093));
  jor  g15835(.dina(n1942), .dinb(n9725), .dout(n16094));
  jor  g15836(.dina(n1944), .dinb(n10314), .dout(n16095));
  jand g15837(.dina(n16095), .dinb(n16094), .dout(n16096));
  jand g15838(.dina(n16096), .dinb(n16093), .dout(n16097));
  jand g15839(.dina(n16097), .dinb(n16092), .dout(n16098));
  jxor g15840(.dina(n16098), .dinb(a23 ), .dout(n16099));
  jnot g15841(.din(n16063), .dout(n16100));
  jand g15842(.dina(n16100), .dinb(n16059), .dout(n16101));
  jnot g15843(.din(n16101), .dout(n16102));
  jand g15844(.dina(n16063), .dinb(n16060), .dout(n16103));
  jor  g15845(.dina(n16103), .dinb(n16051), .dout(n16104));
  jand g15846(.dina(n16104), .dinb(n16102), .dout(n16105));
  jnot g15847(.din(n16105), .dout(n16106));
  jxor g15848(.dina(n16106), .dinb(n16099), .dout(n16107));
  jor  g15849(.dina(n9387), .dinb(n2319), .dout(n16108));
  jor  g15850(.dina(n2224), .dinb(n8789), .dout(n16109));
  jor  g15851(.dina(n2322), .dinb(n8809), .dout(n16110));
  jor  g15852(.dina(n2324), .dinb(n9390), .dout(n16111));
  jand g15853(.dina(n16111), .dinb(n16110), .dout(n16112));
  jand g15854(.dina(n16112), .dinb(n16109), .dout(n16113));
  jand g15855(.dina(n16113), .dinb(n16108), .dout(n16114));
  jxor g15856(.dina(n16114), .dinb(a26 ), .dout(n16115));
  jand g15857(.dina(n15882), .dinb(n15878), .dout(n16116));
  jor  g15858(.dina(n15882), .dinb(n15878), .dout(n16117));
  jand g15859(.dina(n16049), .dinb(n16117), .dout(n16118));
  jor  g15860(.dina(n16118), .dinb(n16116), .dout(n16119));
  jxor g15861(.dina(n16119), .dinb(n16115), .dout(n16120));
  jor  g15862(.dina(n8228), .dinb(n2784), .dout(n16121));
  jor  g15863(.dina(n2661), .dinb(n7683), .dout(n16122));
  jor  g15864(.dina(n2787), .dinb(n7960), .dout(n16123));
  jor  g15865(.dina(n2789), .dinb(n8231), .dout(n16124));
  jand g15866(.dina(n16124), .dinb(n16123), .dout(n16125));
  jand g15867(.dina(n16125), .dinb(n16122), .dout(n16126));
  jand g15868(.dina(n16126), .dinb(n16121), .dout(n16127));
  jxor g15869(.dina(n16127), .dinb(a29 ), .dout(n16128));
  jnot g15870(.din(n16128), .dout(n16129));
  jand g15871(.dina(n16046), .dinb(n16043), .dout(n16130));
  jnot g15872(.din(n16046), .dout(n16131));
  jand g15873(.dina(n16131), .dinb(n16042), .dout(n16132));
  jnot g15874(.din(n16132), .dout(n16133));
  jand g15875(.dina(n16133), .dinb(n16034), .dout(n16134));
  jor  g15876(.dina(n16134), .dinb(n16130), .dout(n16135));
  jxor g15877(.dina(n16135), .dinb(n16129), .dout(n16136));
  jor  g15878(.dina(n7408), .dinb(n3301), .dout(n16137));
  jor  g15879(.dina(n3136), .dinb(n7129), .dout(n16138));
  jor  g15880(.dina(n3304), .dinb(n7149), .dout(n16139));
  jor  g15881(.dina(n3306), .dinb(n7411), .dout(n16140));
  jand g15882(.dina(n16140), .dinb(n16139), .dout(n16141));
  jand g15883(.dina(n16141), .dinb(n16138), .dout(n16142));
  jand g15884(.dina(n16142), .dinb(n16137), .dout(n16143));
  jxor g15885(.dina(n16143), .dinb(a32 ), .dout(n16144));
  jor  g15886(.dina(n16028), .dinb(n16020), .dout(n16145));
  jand g15887(.dina(n16033), .dinb(n16029), .dout(n16146));
  jnot g15888(.din(n16146), .dout(n16147));
  jand g15889(.dina(n16147), .dinb(n16145), .dout(n16148));
  jxor g15890(.dina(n16148), .dinb(n16144), .dout(n16149));
  jor  g15891(.dina(n16017), .dinb(n16009), .dout(n16150));
  jand g15892(.dina(n16018), .dinb(n15886), .dout(n16151));
  jnot g15893(.din(n16151), .dout(n16152));
  jand g15894(.dina(n16152), .dinb(n16150), .dout(n16153));
  jnot g15895(.din(n16153), .dout(n16154));
  jand g15896(.dina(n16006), .dinb(n15898), .dout(n16155));
  jand g15897(.dina(n16007), .dinb(n15889), .dout(n16156));
  jor  g15898(.dina(n16156), .dinb(n16155), .dout(n16157));
  jor  g15899(.dina(n16004), .dinb(n15996), .dout(n16158));
  jand g15900(.dina(n16005), .dinb(n15901), .dout(n16159));
  jnot g15901(.din(n16159), .dout(n16160));
  jand g15902(.dina(n16160), .dinb(n16158), .dout(n16161));
  jnot g15903(.din(n16161), .dout(n16162));
  jor  g15904(.dina(n5739), .dinb(n4554), .dout(n16163));
  jor  g15905(.dina(n5574), .dinb(n4340), .dout(n16164));
  jor  g15906(.dina(n5742), .dinb(n4537), .dout(n16165));
  jor  g15907(.dina(n5744), .dinb(n4557), .dout(n16166));
  jand g15908(.dina(n16166), .dinb(n16165), .dout(n16167));
  jand g15909(.dina(n16167), .dinb(n16164), .dout(n16168));
  jand g15910(.dina(n16168), .dinb(n16163), .dout(n16169));
  jxor g15911(.dina(n16169), .dinb(a44 ), .dout(n16170));
  jnot g15912(.din(n16170), .dout(n16171));
  jand g15913(.dina(n15988), .dinb(n15910), .dout(n16172));
  jnot g15914(.din(n16172), .dout(n16173));
  jor  g15915(.dina(n15994), .dinb(n15990), .dout(n16174));
  jand g15916(.dina(n16174), .dinb(n16173), .dout(n16175));
  jnot g15917(.din(n16175), .dout(n16176));
  jand g15918(.dina(n15986), .dinb(n15983), .dout(n16177));
  jand g15919(.dina(n15987), .dinb(n15974), .dout(n16178));
  jor  g15920(.dina(n16178), .dinb(n16177), .dout(n16179));
  jor  g15921(.dina(n15968), .dinb(n15960), .dout(n16180));
  jand g15922(.dina(n15973), .dinb(n15969), .dout(n16181));
  jnot g15923(.din(n16181), .dout(n16182));
  jand g15924(.dina(n16182), .dinb(n16180), .dout(n16183));
  jnot g15925(.din(n16183), .dout(n16184));
  jor  g15926(.dina(n8978), .dinb(n2556), .dout(n16185));
  jor  g15927(.dina(n8677), .dinb(n2148), .dout(n16186));
  jor  g15928(.dina(n8981), .dinb(n2407), .dout(n16187));
  jor  g15929(.dina(n8983), .dinb(n2559), .dout(n16188));
  jand g15930(.dina(n16188), .dinb(n16187), .dout(n16189));
  jand g15931(.dina(n16189), .dinb(n16186), .dout(n16190));
  jand g15932(.dina(n16190), .dinb(n16185), .dout(n16191));
  jxor g15933(.dina(n16191), .dinb(a56 ), .dout(n16192));
  jnot g15934(.din(n16192), .dout(n16193));
  jand g15935(.dina(n15946), .dinb(n15927), .dout(n16194));
  jand g15936(.dina(n15947), .dinb(n15918), .dout(n16195));
  jor  g15937(.dina(n16195), .dinb(n16194), .dout(n16196));
  jand g15938(.dina(n15942), .dinb(n15821), .dout(n16197));
  jand g15939(.dina(n15943), .dinb(n15707), .dout(n16198));
  jor  g15940(.dina(n16198), .dinb(n16197), .dout(n16199));
  jand g15941(.dina(n10801), .dinb(b19 ), .dout(n16200));
  jand g15942(.dina(n11107), .dinb(b18 ), .dout(n16201));
  jor  g15943(.dina(n16201), .dinb(n16200), .dout(n16202));
  jnot g15944(.din(n16202), .dout(n16203));
  jxor g15945(.dina(n16203), .dinb(n16199), .dout(n16204));
  jnot g15946(.din(n16204), .dout(n16205));
  jor  g15947(.dina(n10806), .dinb(n1739), .dout(n16206));
  jor  g15948(.dina(n10485), .dinb(n1420), .dout(n16207));
  jor  g15949(.dina(n10809), .dinb(n1620), .dout(n16208));
  jor  g15950(.dina(n10811), .dinb(n1742), .dout(n16209));
  jand g15951(.dina(n16209), .dinb(n16208), .dout(n16210));
  jand g15952(.dina(n16210), .dinb(n16207), .dout(n16211));
  jand g15953(.dina(n16211), .dinb(n16206), .dout(n16212));
  jxor g15954(.dina(n16212), .dinb(a62 ), .dout(n16213));
  jxor g15955(.dina(n16213), .dinb(n16205), .dout(n16214));
  jand g15956(.dina(n15944), .dinb(n15939), .dout(n16215));
  jand g15957(.dina(n15945), .dinb(n15930), .dout(n16216));
  jor  g15958(.dina(n16216), .dinb(n16215), .dout(n16217));
  jxor g15959(.dina(n16217), .dinb(n16214), .dout(n16218));
  jnot g15960(.din(n16218), .dout(n16219));
  jor  g15961(.dina(n9891), .dinb(n2007), .dout(n16220));
  jor  g15962(.dina(n9593), .dinb(n1867), .dout(n16221));
  jor  g15963(.dina(n9894), .dinb(n1887), .dout(n16222));
  jor  g15964(.dina(n9896), .dinb(n2010), .dout(n16223));
  jand g15965(.dina(n16223), .dinb(n16222), .dout(n16224));
  jand g15966(.dina(n16224), .dinb(n16221), .dout(n16225));
  jand g15967(.dina(n16225), .dinb(n16220), .dout(n16226));
  jxor g15968(.dina(n16226), .dinb(a59 ), .dout(n16227));
  jxor g15969(.dina(n16227), .dinb(n16219), .dout(n16228));
  jxor g15970(.dina(n16228), .dinb(n16196), .dout(n16229));
  jxor g15971(.dina(n16229), .dinb(n16193), .dout(n16230));
  jnot g15972(.din(n16230), .dout(n16231));
  jor  g15973(.dina(n15957), .dinb(n15949), .dout(n16232));
  jand g15974(.dina(n15958), .dinb(n15913), .dout(n16233));
  jnot g15975(.din(n16233), .dout(n16234));
  jand g15976(.dina(n16234), .dinb(n16232), .dout(n16235));
  jxor g15977(.dina(n16235), .dinb(n16231), .dout(n16236));
  jor  g15978(.dina(n8125), .dinb(n3032), .dout(n16237));
  jor  g15979(.dina(n7846), .dinb(n2579), .dout(n16238));
  jor  g15980(.dina(n8128), .dinb(n2870), .dout(n16239));
  jor  g15981(.dina(n8130), .dinb(n3035), .dout(n16240));
  jand g15982(.dina(n16240), .dinb(n16239), .dout(n16241));
  jand g15983(.dina(n16241), .dinb(n16238), .dout(n16242));
  jand g15984(.dina(n16242), .dinb(n16237), .dout(n16243));
  jxor g15985(.dina(n16243), .dinb(a53 ), .dout(n16244));
  jnot g15986(.din(n16244), .dout(n16245));
  jxor g15987(.dina(n16245), .dinb(n16236), .dout(n16246));
  jxor g15988(.dina(n16246), .dinb(n16184), .dout(n16247));
  jor  g15989(.dina(n7266), .dinb(n3400), .dout(n16248));
  jor  g15990(.dina(n7021), .dinb(n3055), .dout(n16249));
  jor  g15991(.dina(n7269), .dinb(n3230), .dout(n16250));
  jor  g15992(.dina(n7271), .dinb(n3403), .dout(n16251));
  jand g15993(.dina(n16251), .dinb(n16250), .dout(n16252));
  jand g15994(.dina(n16252), .dinb(n16249), .dout(n16253));
  jand g15995(.dina(n16253), .dinb(n16248), .dout(n16254));
  jxor g15996(.dina(n16254), .dinb(a50 ), .dout(n16255));
  jnot g15997(.din(n16255), .dout(n16256));
  jxor g15998(.dina(n16256), .dinb(n16247), .dout(n16257));
  jxor g15999(.dina(n16257), .dinb(n16179), .dout(n16258));
  jnot g16000(.din(n16258), .dout(n16259));
  jor  g16001(.dina(n6490), .dinb(n4137), .dout(n16260));
  jor  g16002(.dina(n6262), .dinb(n3588), .dout(n16261));
  jor  g16003(.dina(n6493), .dinb(n3942), .dout(n16262));
  jor  g16004(.dina(n6495), .dinb(n4140), .dout(n16263));
  jand g16005(.dina(n16263), .dinb(n16262), .dout(n16264));
  jand g16006(.dina(n16264), .dinb(n16261), .dout(n16265));
  jand g16007(.dina(n16265), .dinb(n16260), .dout(n16266));
  jxor g16008(.dina(n16266), .dinb(a47 ), .dout(n16267));
  jxor g16009(.dina(n16267), .dinb(n16259), .dout(n16268));
  jxor g16010(.dina(n16268), .dinb(n16176), .dout(n16269));
  jxor g16011(.dina(n16269), .dinb(n16171), .dout(n16270));
  jxor g16012(.dina(n16270), .dinb(n16162), .dout(n16271));
  jor  g16013(.dina(n5405), .dinb(n5096), .dout(n16272));
  jor  g16014(.dina(n4904), .dinb(n4974), .dout(n16273));
  jor  g16015(.dina(n5099), .dinb(n4994), .dout(n16274));
  jor  g16016(.dina(n5101), .dinb(n5408), .dout(n16275));
  jand g16017(.dina(n16275), .dinb(n16274), .dout(n16276));
  jand g16018(.dina(n16276), .dinb(n16273), .dout(n16277));
  jand g16019(.dina(n16277), .dinb(n16272), .dout(n16278));
  jxor g16020(.dina(n16278), .dinb(a41 ), .dout(n16279));
  jnot g16021(.din(n16279), .dout(n16280));
  jxor g16022(.dina(n16280), .dinb(n16271), .dout(n16281));
  jxor g16023(.dina(n16281), .dinb(n16157), .dout(n16282));
  jor  g16024(.dina(n6103), .dinb(n4415), .dout(n16283));
  jor  g16025(.dina(n4272), .dinb(n5428), .dout(n16284));
  jor  g16026(.dina(n4418), .dinb(n5862), .dout(n16285));
  jor  g16027(.dina(n4420), .dinb(n6106), .dout(n16286));
  jand g16028(.dina(n16286), .dinb(n16285), .dout(n16287));
  jand g16029(.dina(n16287), .dinb(n16284), .dout(n16288));
  jand g16030(.dina(n16288), .dinb(n16283), .dout(n16289));
  jxor g16031(.dina(n16289), .dinb(a38 ), .dout(n16290));
  jnot g16032(.din(n16290), .dout(n16291));
  jxor g16033(.dina(n16291), .dinb(n16282), .dout(n16292));
  jxor g16034(.dina(n16292), .dinb(n16154), .dout(n16293));
  jor  g16035(.dina(n6864), .dinb(n3849), .dout(n16294));
  jor  g16036(.dina(n3689), .dinb(n6352), .dout(n16295));
  jor  g16037(.dina(n3852), .dinb(n6372), .dout(n16296));
  jor  g16038(.dina(n3854), .dinb(n6867), .dout(n16297));
  jand g16039(.dina(n16297), .dinb(n16296), .dout(n16298));
  jand g16040(.dina(n16298), .dinb(n16295), .dout(n16299));
  jand g16041(.dina(n16299), .dinb(n16294), .dout(n16300));
  jxor g16042(.dina(n16300), .dinb(a35 ), .dout(n16301));
  jnot g16043(.din(n16301), .dout(n16302));
  jxor g16044(.dina(n16302), .dinb(n16293), .dout(n16303));
  jxor g16045(.dina(n16303), .dinb(n16149), .dout(n16304));
  jxor g16046(.dina(n16304), .dinb(n16136), .dout(n16305));
  jxor g16047(.dina(n16305), .dinb(n16120), .dout(n16306));
  jxor g16048(.dina(n16306), .dinb(n16107), .dout(n16307));
  jxor g16049(.dina(n16307), .dinb(n16091), .dout(n16308));
  jxor g16050(.dina(n16308), .dinb(n16077), .dout(n16309));
  jxor g16051(.dina(n16309), .dinb(n16072), .dout(f82 ));
  jand g16052(.dina(n16308), .dinb(n16077), .dout(n16311));
  jand g16053(.dina(n16309), .dinb(n16072), .dout(n16312));
  jor  g16054(.dina(n16312), .dinb(n16311), .dout(n16313));
  jand g16055(.dina(n16090), .dinb(n16084), .dout(n16314));
  jand g16056(.dina(n16307), .dinb(n16091), .dout(n16315));
  jor  g16057(.dina(n16315), .dinb(n16314), .dout(n16316));
  jor  g16058(.dina(n9410), .dinb(n2319), .dout(n16317));
  jor  g16059(.dina(n2224), .dinb(n8809), .dout(n16318));
  jor  g16060(.dina(n2322), .dinb(n9390), .dout(n16319));
  jor  g16061(.dina(n2324), .dinb(n9413), .dout(n16320));
  jand g16062(.dina(n16320), .dinb(n16319), .dout(n16321));
  jand g16063(.dina(n16321), .dinb(n16318), .dout(n16322));
  jand g16064(.dina(n16322), .dinb(n16317), .dout(n16323));
  jxor g16065(.dina(n16323), .dinb(a26 ), .dout(n16324));
  jnot g16066(.din(n16324), .dout(n16325));
  jand g16067(.dina(n16135), .dinb(n16129), .dout(n16326));
  jand g16068(.dina(n16304), .dinb(n16136), .dout(n16327));
  jor  g16069(.dina(n16327), .dinb(n16326), .dout(n16328));
  jxor g16070(.dina(n16328), .dinb(n16325), .dout(n16329));
  jor  g16071(.dina(n7680), .dinb(n3301), .dout(n16330));
  jor  g16072(.dina(n3136), .dinb(n7149), .dout(n16331));
  jor  g16073(.dina(n3304), .dinb(n7411), .dout(n16332));
  jor  g16074(.dina(n3306), .dinb(n7683), .dout(n16333));
  jand g16075(.dina(n16333), .dinb(n16332), .dout(n16334));
  jand g16076(.dina(n16334), .dinb(n16331), .dout(n16335));
  jand g16077(.dina(n16335), .dinb(n16330), .dout(n16336));
  jxor g16078(.dina(n16336), .dinb(a32 ), .dout(n16337));
  jnot g16079(.din(n16337), .dout(n16338));
  jnot g16080(.din(n16292), .dout(n16339));
  jand g16081(.dina(n16339), .dinb(n16153), .dout(n16340));
  jnot g16082(.din(n16340), .dout(n16341));
  jand g16083(.dina(n16292), .dinb(n16154), .dout(n16342));
  jor  g16084(.dina(n16302), .dinb(n16342), .dout(n16343));
  jand g16085(.dina(n16343), .dinb(n16341), .dout(n16344));
  jxor g16086(.dina(n16344), .dinb(n16338), .dout(n16345));
  jor  g16087(.dina(n5425), .dinb(n5096), .dout(n16346));
  jor  g16088(.dina(n4904), .dinb(n4994), .dout(n16347));
  jor  g16089(.dina(n5099), .dinb(n5408), .dout(n16348));
  jor  g16090(.dina(n5101), .dinb(n5428), .dout(n16349));
  jand g16091(.dina(n16349), .dinb(n16348), .dout(n16350));
  jand g16092(.dina(n16350), .dinb(n16347), .dout(n16351));
  jand g16093(.dina(n16351), .dinb(n16346), .dout(n16352));
  jxor g16094(.dina(n16352), .dinb(a41 ), .dout(n16353));
  jnot g16095(.din(n16353), .dout(n16354));
  jand g16096(.dina(n16268), .dinb(n16176), .dout(n16355));
  jand g16097(.dina(n16269), .dinb(n16171), .dout(n16356));
  jor  g16098(.dina(n16356), .dinb(n16355), .dout(n16357));
  jor  g16099(.dina(n5739), .dinb(n4971), .dout(n16358));
  jor  g16100(.dina(n5574), .dinb(n4537), .dout(n16359));
  jor  g16101(.dina(n5742), .dinb(n4557), .dout(n16360));
  jor  g16102(.dina(n5744), .dinb(n4974), .dout(n16361));
  jand g16103(.dina(n16361), .dinb(n16360), .dout(n16362));
  jand g16104(.dina(n16362), .dinb(n16359), .dout(n16363));
  jand g16105(.dina(n16363), .dinb(n16358), .dout(n16364));
  jxor g16106(.dina(n16364), .dinb(a44 ), .dout(n16365));
  jnot g16107(.din(n16365), .dout(n16366));
  jand g16108(.dina(n16257), .dinb(n16179), .dout(n16367));
  jnot g16109(.din(n16367), .dout(n16368));
  jor  g16110(.dina(n16267), .dinb(n16259), .dout(n16369));
  jand g16111(.dina(n16369), .dinb(n16368), .dout(n16370));
  jnot g16112(.din(n16370), .dout(n16371));
  jor  g16113(.dina(n6490), .dinb(n4337), .dout(n16372));
  jor  g16114(.dina(n6262), .dinb(n3942), .dout(n16373));
  jor  g16115(.dina(n6493), .dinb(n4140), .dout(n16374));
  jor  g16116(.dina(n6495), .dinb(n4340), .dout(n16375));
  jand g16117(.dina(n16375), .dinb(n16374), .dout(n16376));
  jand g16118(.dina(n16376), .dinb(n16373), .dout(n16377));
  jand g16119(.dina(n16377), .dinb(n16372), .dout(n16378));
  jxor g16120(.dina(n16378), .dinb(a47 ), .dout(n16379));
  jnot g16121(.din(n16379), .dout(n16380));
  jor  g16122(.dina(n7266), .dinb(n3585), .dout(n16381));
  jor  g16123(.dina(n7021), .dinb(n3230), .dout(n16382));
  jor  g16124(.dina(n7269), .dinb(n3403), .dout(n16383));
  jor  g16125(.dina(n7271), .dinb(n3588), .dout(n16384));
  jand g16126(.dina(n16384), .dinb(n16383), .dout(n16385));
  jand g16127(.dina(n16385), .dinb(n16382), .dout(n16386));
  jand g16128(.dina(n16386), .dinb(n16381), .dout(n16387));
  jxor g16129(.dina(n16387), .dinb(a50 ), .dout(n16388));
  jnot g16130(.din(n16388), .dout(n16389));
  jor  g16131(.dina(n8125), .dinb(n3052), .dout(n16390));
  jor  g16132(.dina(n7846), .dinb(n2870), .dout(n16391));
  jor  g16133(.dina(n8128), .dinb(n3035), .dout(n16392));
  jor  g16134(.dina(n8130), .dinb(n3055), .dout(n16393));
  jand g16135(.dina(n16393), .dinb(n16392), .dout(n16394));
  jand g16136(.dina(n16394), .dinb(n16391), .dout(n16395));
  jand g16137(.dina(n16395), .dinb(n16390), .dout(n16396));
  jxor g16138(.dina(n16396), .dinb(a53 ), .dout(n16397));
  jnot g16139(.din(n16397), .dout(n16398));
  jand g16140(.dina(n16228), .dinb(n16196), .dout(n16399));
  jand g16141(.dina(n16229), .dinb(n16193), .dout(n16400));
  jor  g16142(.dina(n16400), .dinb(n16399), .dout(n16401));
  jor  g16143(.dina(n9891), .dinb(n2145), .dout(n16402));
  jor  g16144(.dina(n9593), .dinb(n1887), .dout(n16403));
  jor  g16145(.dina(n9894), .dinb(n2010), .dout(n16404));
  jor  g16146(.dina(n9896), .dinb(n2148), .dout(n16405));
  jand g16147(.dina(n16405), .dinb(n16404), .dout(n16406));
  jand g16148(.dina(n16406), .dinb(n16403), .dout(n16407));
  jand g16149(.dina(n16407), .dinb(n16402), .dout(n16408));
  jxor g16150(.dina(n16408), .dinb(a59 ), .dout(n16409));
  jnot g16151(.din(n16409), .dout(n16410));
  jand g16152(.dina(n16203), .dinb(n16199), .dout(n16411));
  jnot g16153(.din(n16411), .dout(n16412));
  jor  g16154(.dina(n16213), .dinb(n16205), .dout(n16413));
  jand g16155(.dina(n16413), .dinb(n16412), .dout(n16414));
  jnot g16156(.din(n16414), .dout(n16415));
  jand g16157(.dina(n10801), .dinb(b20 ), .dout(n16416));
  jand g16158(.dina(n11107), .dinb(b19 ), .dout(n16417));
  jor  g16159(.dina(n16417), .dinb(n16416), .dout(n16418));
  jnot g16160(.din(n16418), .dout(n16419));
  jxor g16161(.dina(n16419), .dinb(n16202), .dout(n16420));
  jnot g16162(.din(n16420), .dout(n16421));
  jor  g16163(.dina(n10806), .dinb(n1864), .dout(n16422));
  jor  g16164(.dina(n10485), .dinb(n1620), .dout(n16423));
  jor  g16165(.dina(n10809), .dinb(n1742), .dout(n16424));
  jor  g16166(.dina(n10811), .dinb(n1867), .dout(n16425));
  jand g16167(.dina(n16425), .dinb(n16424), .dout(n16426));
  jand g16168(.dina(n16426), .dinb(n16423), .dout(n16427));
  jand g16169(.dina(n16427), .dinb(n16422), .dout(n16428));
  jxor g16170(.dina(n16428), .dinb(a62 ), .dout(n16429));
  jxor g16171(.dina(n16429), .dinb(n16421), .dout(n16430));
  jxor g16172(.dina(n16430), .dinb(n16415), .dout(n16431));
  jxor g16173(.dina(n16431), .dinb(n16410), .dout(n16432));
  jand g16174(.dina(n16217), .dinb(n16214), .dout(n16433));
  jnot g16175(.din(n16433), .dout(n16434));
  jnot g16176(.din(n16214), .dout(n16435));
  jnot g16177(.din(n16217), .dout(n16436));
  jand g16178(.dina(n16436), .dinb(n16435), .dout(n16437));
  jor  g16179(.dina(n16227), .dinb(n16437), .dout(n16438));
  jand g16180(.dina(n16438), .dinb(n16434), .dout(n16439));
  jnot g16181(.din(n16439), .dout(n16440));
  jxor g16182(.dina(n16440), .dinb(n16432), .dout(n16441));
  jnot g16183(.din(n16441), .dout(n16442));
  jor  g16184(.dina(n8978), .dinb(n2576), .dout(n16443));
  jor  g16185(.dina(n8677), .dinb(n2407), .dout(n16444));
  jor  g16186(.dina(n8981), .dinb(n2559), .dout(n16445));
  jor  g16187(.dina(n8983), .dinb(n2579), .dout(n16446));
  jand g16188(.dina(n16446), .dinb(n16445), .dout(n16447));
  jand g16189(.dina(n16447), .dinb(n16444), .dout(n16448));
  jand g16190(.dina(n16448), .dinb(n16443), .dout(n16449));
  jxor g16191(.dina(n16449), .dinb(a56 ), .dout(n16450));
  jxor g16192(.dina(n16450), .dinb(n16442), .dout(n16451));
  jxor g16193(.dina(n16451), .dinb(n16401), .dout(n16452));
  jxor g16194(.dina(n16452), .dinb(n16398), .dout(n16453));
  jnot g16195(.din(n16453), .dout(n16454));
  jnot g16196(.din(n16235), .dout(n16455));
  jand g16197(.dina(n16455), .dinb(n16230), .dout(n16456));
  jnot g16198(.din(n16456), .dout(n16457));
  jand g16199(.dina(n16235), .dinb(n16231), .dout(n16458));
  jor  g16200(.dina(n16244), .dinb(n16458), .dout(n16459));
  jand g16201(.dina(n16459), .dinb(n16457), .dout(n16460));
  jxor g16202(.dina(n16460), .dinb(n16454), .dout(n16461));
  jxor g16203(.dina(n16461), .dinb(n16389), .dout(n16462));
  jnot g16204(.din(n16246), .dout(n16463));
  jand g16205(.dina(n16463), .dinb(n16183), .dout(n16464));
  jnot g16206(.din(n16464), .dout(n16465));
  jand g16207(.dina(n16246), .dinb(n16184), .dout(n16466));
  jor  g16208(.dina(n16256), .dinb(n16466), .dout(n16467));
  jand g16209(.dina(n16467), .dinb(n16465), .dout(n16468));
  jxor g16210(.dina(n16468), .dinb(n16462), .dout(n16469));
  jxor g16211(.dina(n16469), .dinb(n16380), .dout(n16470));
  jxor g16212(.dina(n16470), .dinb(n16371), .dout(n16471));
  jxor g16213(.dina(n16471), .dinb(n16366), .dout(n16472));
  jxor g16214(.dina(n16472), .dinb(n16357), .dout(n16473));
  jxor g16215(.dina(n16473), .dinb(n16354), .dout(n16474));
  jor  g16216(.dina(n16270), .dinb(n16162), .dout(n16475));
  jand g16217(.dina(n16270), .dinb(n16162), .dout(n16476));
  jor  g16218(.dina(n16280), .dinb(n16476), .dout(n16477));
  jand g16219(.dina(n16477), .dinb(n16475), .dout(n16478));
  jxor g16220(.dina(n16478), .dinb(n16474), .dout(n16479));
  jor  g16221(.dina(n6349), .dinb(n4415), .dout(n16480));
  jor  g16222(.dina(n4272), .dinb(n5862), .dout(n16481));
  jor  g16223(.dina(n4418), .dinb(n6106), .dout(n16482));
  jor  g16224(.dina(n4420), .dinb(n6352), .dout(n16483));
  jand g16225(.dina(n16483), .dinb(n16482), .dout(n16484));
  jand g16226(.dina(n16484), .dinb(n16481), .dout(n16485));
  jand g16227(.dina(n16485), .dinb(n16480), .dout(n16486));
  jxor g16228(.dina(n16486), .dinb(a38 ), .dout(n16487));
  jnot g16229(.din(n16487), .dout(n16488));
  jxor g16230(.dina(n16488), .dinb(n16479), .dout(n16489));
  jnot g16231(.din(n16157), .dout(n16490));
  jnot g16232(.din(n16281), .dout(n16491));
  jand g16233(.dina(n16491), .dinb(n16490), .dout(n16492));
  jnot g16234(.din(n16492), .dout(n16493));
  jand g16235(.dina(n16281), .dinb(n16157), .dout(n16494));
  jor  g16236(.dina(n16291), .dinb(n16494), .dout(n16495));
  jand g16237(.dina(n16495), .dinb(n16493), .dout(n16496));
  jxor g16238(.dina(n16496), .dinb(n16489), .dout(n16497));
  jnot g16239(.din(n16497), .dout(n16498));
  jor  g16240(.dina(n7126), .dinb(n3849), .dout(n16499));
  jor  g16241(.dina(n3689), .dinb(n6372), .dout(n16500));
  jor  g16242(.dina(n3852), .dinb(n6867), .dout(n16501));
  jor  g16243(.dina(n3854), .dinb(n7129), .dout(n16502));
  jand g16244(.dina(n16502), .dinb(n16501), .dout(n16503));
  jand g16245(.dina(n16503), .dinb(n16500), .dout(n16504));
  jand g16246(.dina(n16504), .dinb(n16499), .dout(n16505));
  jxor g16247(.dina(n16505), .dinb(a35 ), .dout(n16506));
  jxor g16248(.dina(n16506), .dinb(n16498), .dout(n16507));
  jxor g16249(.dina(n16507), .dinb(n16345), .dout(n16508));
  jor  g16250(.dina(n8786), .dinb(n2784), .dout(n16509));
  jor  g16251(.dina(n2661), .dinb(n7960), .dout(n16510));
  jor  g16252(.dina(n2787), .dinb(n8231), .dout(n16511));
  jor  g16253(.dina(n2789), .dinb(n8789), .dout(n16512));
  jand g16254(.dina(n16512), .dinb(n16511), .dout(n16513));
  jand g16255(.dina(n16513), .dinb(n16510), .dout(n16514));
  jand g16256(.dina(n16514), .dinb(n16509), .dout(n16515));
  jxor g16257(.dina(n16515), .dinb(a29 ), .dout(n16516));
  jor  g16258(.dina(n16148), .dinb(n16144), .dout(n16517));
  jand g16259(.dina(n16303), .dinb(n16149), .dout(n16518));
  jnot g16260(.din(n16518), .dout(n16519));
  jand g16261(.dina(n16519), .dinb(n16517), .dout(n16520));
  jxor g16262(.dina(n16520), .dinb(n16516), .dout(n16521));
  jxor g16263(.dina(n16521), .dinb(n16508), .dout(n16522));
  jxor g16264(.dina(n16522), .dinb(n16329), .dout(n16523));
  jor  g16265(.dina(n10634), .dinb(n1939), .dout(n16524));
  jor  g16266(.dina(n1827), .dinb(n9725), .dout(n16525));
  jor  g16267(.dina(n1942), .dinb(n10314), .dout(n16526));
  jor  g16268(.dina(n1944), .dinb(n10637), .dout(n16527));
  jand g16269(.dina(n16527), .dinb(n16526), .dout(n16528));
  jand g16270(.dina(n16528), .dinb(n16525), .dout(n16529));
  jand g16271(.dina(n16529), .dinb(n16524), .dout(n16530));
  jxor g16272(.dina(n16530), .dinb(a23 ), .dout(n16531));
  jnot g16273(.din(n16531), .dout(n16532));
  jnot g16274(.din(n16115), .dout(n16533));
  jnot g16275(.din(n16119), .dout(n16534));
  jand g16276(.dina(n16534), .dinb(n16533), .dout(n16535));
  jand g16277(.dina(n16305), .dinb(n16120), .dout(n16536));
  jor  g16278(.dina(n16536), .dinb(n16535), .dout(n16537));
  jxor g16279(.dina(n16537), .dinb(n16532), .dout(n16538));
  jxor g16280(.dina(n16538), .dinb(n16523), .dout(n16539));
  jnot g16281(.din(a20 ), .dout(n16540));
  jand g16282(.dina(n11296), .dinb(n1345), .dout(n16541));
  jor  g16283(.dina(n16541), .dinb(n1490), .dout(n16542));
  jand g16284(.dina(n16542), .dinb(b63 ), .dout(n16543));
  jxor g16285(.dina(n16543), .dinb(n16540), .dout(n16544));
  jnot g16286(.din(n16544), .dout(n16545));
  jand g16287(.dina(n16106), .dinb(n16099), .dout(n16546));
  jnot g16288(.din(n16546), .dout(n16547));
  jnot g16289(.din(n16099), .dout(n16548));
  jand g16290(.dina(n16105), .dinb(n16548), .dout(n16549));
  jor  g16291(.dina(n16306), .dinb(n16549), .dout(n16550));
  jand g16292(.dina(n16550), .dinb(n16547), .dout(n16551));
  jxor g16293(.dina(n16551), .dinb(n16545), .dout(n16552));
  jxor g16294(.dina(n16552), .dinb(n16539), .dout(n16553));
  jxor g16295(.dina(n16553), .dinb(n16316), .dout(n16554));
  jxor g16296(.dina(n16554), .dinb(n16313), .dout(f83 ));
  jand g16297(.dina(n16551), .dinb(n16545), .dout(n16556));
  jand g16298(.dina(n16552), .dinb(n16539), .dout(n16557));
  jor  g16299(.dina(n16557), .dinb(n16556), .dout(n16558));
  jor  g16300(.dina(n9722), .dinb(n2319), .dout(n16559));
  jor  g16301(.dina(n2224), .dinb(n9390), .dout(n16560));
  jor  g16302(.dina(n2322), .dinb(n9413), .dout(n16561));
  jor  g16303(.dina(n2324), .dinb(n9725), .dout(n16562));
  jand g16304(.dina(n16562), .dinb(n16561), .dout(n16563));
  jand g16305(.dina(n16563), .dinb(n16560), .dout(n16564));
  jand g16306(.dina(n16564), .dinb(n16559), .dout(n16565));
  jxor g16307(.dina(n16565), .dinb(a26 ), .dout(n16566));
  jnot g16308(.din(n16566), .dout(n16567));
  jand g16309(.dina(n16328), .dinb(n16325), .dout(n16568));
  jand g16310(.dina(n16522), .dinb(n16329), .dout(n16569));
  jor  g16311(.dina(n16569), .dinb(n16568), .dout(n16570));
  jxor g16312(.dina(n16570), .dinb(n16567), .dout(n16571));
  jor  g16313(.dina(n7957), .dinb(n3301), .dout(n16572));
  jor  g16314(.dina(n3136), .dinb(n7411), .dout(n16573));
  jor  g16315(.dina(n3304), .dinb(n7683), .dout(n16574));
  jor  g16316(.dina(n3306), .dinb(n7960), .dout(n16575));
  jand g16317(.dina(n16575), .dinb(n16574), .dout(n16576));
  jand g16318(.dina(n16576), .dinb(n16573), .dout(n16577));
  jand g16319(.dina(n16577), .dinb(n16572), .dout(n16578));
  jxor g16320(.dina(n16578), .dinb(a32 ), .dout(n16579));
  jnot g16321(.din(n16579), .dout(n16580));
  jand g16322(.dina(n16344), .dinb(n16338), .dout(n16581));
  jand g16323(.dina(n16507), .dinb(n16345), .dout(n16582));
  jor  g16324(.dina(n16582), .dinb(n16581), .dout(n16583));
  jxor g16325(.dina(n16583), .dinb(n16580), .dout(n16584));
  jnot g16326(.din(n16584), .dout(n16585));
  jand g16327(.dina(n16496), .dinb(n16489), .dout(n16586));
  jnot g16328(.din(n16586), .dout(n16587));
  jor  g16329(.dina(n16506), .dinb(n16498), .dout(n16588));
  jand g16330(.dina(n16588), .dinb(n16587), .dout(n16589));
  jand g16331(.dina(n16472), .dinb(n16357), .dout(n16590));
  jand g16332(.dina(n16473), .dinb(n16354), .dout(n16591));
  jor  g16333(.dina(n16591), .dinb(n16590), .dout(n16592));
  jand g16334(.dina(n16470), .dinb(n16371), .dout(n16593));
  jand g16335(.dina(n16471), .dinb(n16366), .dout(n16594));
  jor  g16336(.dina(n16594), .dinb(n16593), .dout(n16595));
  jand g16337(.dina(n16468), .dinb(n16462), .dout(n16596));
  jand g16338(.dina(n16469), .dinb(n16380), .dout(n16597));
  jor  g16339(.dina(n16597), .dinb(n16596), .dout(n16598));
  jor  g16340(.dina(n16460), .dinb(n16454), .dout(n16599));
  jand g16341(.dina(n16461), .dinb(n16389), .dout(n16600));
  jnot g16342(.din(n16600), .dout(n16601));
  jand g16343(.dina(n16601), .dinb(n16599), .dout(n16602));
  jnot g16344(.din(n16602), .dout(n16603));
  jor  g16345(.dina(n7266), .dinb(n3939), .dout(n16604));
  jor  g16346(.dina(n7021), .dinb(n3403), .dout(n16605));
  jor  g16347(.dina(n7269), .dinb(n3588), .dout(n16606));
  jor  g16348(.dina(n7271), .dinb(n3942), .dout(n16607));
  jand g16349(.dina(n16607), .dinb(n16606), .dout(n16608));
  jand g16350(.dina(n16608), .dinb(n16605), .dout(n16609));
  jand g16351(.dina(n16609), .dinb(n16604), .dout(n16610));
  jxor g16352(.dina(n16610), .dinb(a50 ), .dout(n16611));
  jnot g16353(.din(n16611), .dout(n16612));
  jand g16354(.dina(n16440), .dinb(n16432), .dout(n16613));
  jnot g16355(.din(n16613), .dout(n16614));
  jnot g16356(.din(n16432), .dout(n16615));
  jand g16357(.dina(n16439), .dinb(n16615), .dout(n16616));
  jor  g16358(.dina(n16450), .dinb(n16616), .dout(n16617));
  jand g16359(.dina(n16617), .dinb(n16614), .dout(n16618));
  jnot g16360(.din(n16618), .dout(n16619));
  jand g16361(.dina(n16430), .dinb(n16415), .dout(n16620));
  jand g16362(.dina(n16431), .dinb(n16410), .dout(n16621));
  jor  g16363(.dina(n16621), .dinb(n16620), .dout(n16622));
  jor  g16364(.dina(n9891), .dinb(n2404), .dout(n16623));
  jor  g16365(.dina(n9593), .dinb(n2010), .dout(n16624));
  jor  g16366(.dina(n9894), .dinb(n2148), .dout(n16625));
  jor  g16367(.dina(n9896), .dinb(n2407), .dout(n16626));
  jand g16368(.dina(n16626), .dinb(n16625), .dout(n16627));
  jand g16369(.dina(n16627), .dinb(n16624), .dout(n16628));
  jand g16370(.dina(n16628), .dinb(n16623), .dout(n16629));
  jxor g16371(.dina(n16629), .dinb(a59 ), .dout(n16630));
  jnot g16372(.din(n16630), .dout(n16631));
  jand g16373(.dina(n16419), .dinb(n16202), .dout(n16632));
  jnot g16374(.din(n16632), .dout(n16633));
  jor  g16375(.dina(n16429), .dinb(n16421), .dout(n16634));
  jand g16376(.dina(n16634), .dinb(n16633), .dout(n16635));
  jnot g16377(.din(n16635), .dout(n16636));
  jand g16378(.dina(n10801), .dinb(b21 ), .dout(n16637));
  jand g16379(.dina(n11107), .dinb(b20 ), .dout(n16638));
  jor  g16380(.dina(n16638), .dinb(n16637), .dout(n16639));
  jxor g16381(.dina(n16639), .dinb(n16540), .dout(n16640));
  jxor g16382(.dina(n16640), .dinb(n16418), .dout(n16641));
  jnot g16383(.din(n16641), .dout(n16642));
  jor  g16384(.dina(n10806), .dinb(n1884), .dout(n16643));
  jor  g16385(.dina(n10485), .dinb(n1742), .dout(n16644));
  jor  g16386(.dina(n10809), .dinb(n1867), .dout(n16645));
  jor  g16387(.dina(n10811), .dinb(n1887), .dout(n16646));
  jand g16388(.dina(n16646), .dinb(n16645), .dout(n16647));
  jand g16389(.dina(n16647), .dinb(n16644), .dout(n16648));
  jand g16390(.dina(n16648), .dinb(n16643), .dout(n16649));
  jxor g16391(.dina(n16649), .dinb(a62 ), .dout(n16650));
  jxor g16392(.dina(n16650), .dinb(n16642), .dout(n16651));
  jxor g16393(.dina(n16651), .dinb(n16636), .dout(n16652));
  jxor g16394(.dina(n16652), .dinb(n16631), .dout(n16653));
  jxor g16395(.dina(n16653), .dinb(n16622), .dout(n16654));
  jnot g16396(.din(n16654), .dout(n16655));
  jor  g16397(.dina(n8978), .dinb(n2867), .dout(n16656));
  jor  g16398(.dina(n8677), .dinb(n2559), .dout(n16657));
  jor  g16399(.dina(n8981), .dinb(n2579), .dout(n16658));
  jor  g16400(.dina(n8983), .dinb(n2870), .dout(n16659));
  jand g16401(.dina(n16659), .dinb(n16658), .dout(n16660));
  jand g16402(.dina(n16660), .dinb(n16657), .dout(n16661));
  jand g16403(.dina(n16661), .dinb(n16656), .dout(n16662));
  jxor g16404(.dina(n16662), .dinb(a56 ), .dout(n16663));
  jxor g16405(.dina(n16663), .dinb(n16655), .dout(n16664));
  jxor g16406(.dina(n16664), .dinb(n16619), .dout(n16665));
  jor  g16407(.dina(n8125), .dinb(n3227), .dout(n16666));
  jor  g16408(.dina(n7846), .dinb(n3035), .dout(n16667));
  jor  g16409(.dina(n8128), .dinb(n3055), .dout(n16668));
  jor  g16410(.dina(n8130), .dinb(n3230), .dout(n16669));
  jand g16411(.dina(n16669), .dinb(n16668), .dout(n16670));
  jand g16412(.dina(n16670), .dinb(n16667), .dout(n16671));
  jand g16413(.dina(n16671), .dinb(n16666), .dout(n16672));
  jxor g16414(.dina(n16672), .dinb(a53 ), .dout(n16673));
  jnot g16415(.din(n16673), .dout(n16674));
  jand g16416(.dina(n16451), .dinb(n16401), .dout(n16675));
  jand g16417(.dina(n16452), .dinb(n16398), .dout(n16676));
  jor  g16418(.dina(n16676), .dinb(n16675), .dout(n16677));
  jxor g16419(.dina(n16677), .dinb(n16674), .dout(n16678));
  jxor g16420(.dina(n16678), .dinb(n16665), .dout(n16679));
  jxor g16421(.dina(n16679), .dinb(n16612), .dout(n16680));
  jxor g16422(.dina(n16680), .dinb(n16603), .dout(n16681));
  jnot g16423(.din(n16681), .dout(n16682));
  jor  g16424(.dina(n6490), .dinb(n4534), .dout(n16683));
  jor  g16425(.dina(n6262), .dinb(n4140), .dout(n16684));
  jor  g16426(.dina(n6493), .dinb(n4340), .dout(n16685));
  jor  g16427(.dina(n6495), .dinb(n4537), .dout(n16686));
  jand g16428(.dina(n16686), .dinb(n16685), .dout(n16687));
  jand g16429(.dina(n16687), .dinb(n16684), .dout(n16688));
  jand g16430(.dina(n16688), .dinb(n16683), .dout(n16689));
  jxor g16431(.dina(n16689), .dinb(a47 ), .dout(n16690));
  jxor g16432(.dina(n16690), .dinb(n16682), .dout(n16691));
  jxor g16433(.dina(n16691), .dinb(n16598), .dout(n16692));
  jnot g16434(.din(n16692), .dout(n16693));
  jor  g16435(.dina(n5739), .dinb(n4991), .dout(n16694));
  jor  g16436(.dina(n5574), .dinb(n4557), .dout(n16695));
  jor  g16437(.dina(n5742), .dinb(n4974), .dout(n16696));
  jor  g16438(.dina(n5744), .dinb(n4994), .dout(n16697));
  jand g16439(.dina(n16697), .dinb(n16696), .dout(n16698));
  jand g16440(.dina(n16698), .dinb(n16695), .dout(n16699));
  jand g16441(.dina(n16699), .dinb(n16694), .dout(n16700));
  jxor g16442(.dina(n16700), .dinb(a44 ), .dout(n16701));
  jxor g16443(.dina(n16701), .dinb(n16693), .dout(n16702));
  jxor g16444(.dina(n16702), .dinb(n16595), .dout(n16703));
  jnot g16445(.din(n16703), .dout(n16704));
  jor  g16446(.dina(n5859), .dinb(n5096), .dout(n16705));
  jor  g16447(.dina(n4904), .dinb(n5408), .dout(n16706));
  jor  g16448(.dina(n5099), .dinb(n5428), .dout(n16707));
  jor  g16449(.dina(n5101), .dinb(n5862), .dout(n16708));
  jand g16450(.dina(n16708), .dinb(n16707), .dout(n16709));
  jand g16451(.dina(n16709), .dinb(n16706), .dout(n16710));
  jand g16452(.dina(n16710), .dinb(n16705), .dout(n16711));
  jxor g16453(.dina(n16711), .dinb(a41 ), .dout(n16712));
  jxor g16454(.dina(n16712), .dinb(n16704), .dout(n16713));
  jxor g16455(.dina(n16713), .dinb(n16592), .dout(n16714));
  jnot g16456(.din(n16714), .dout(n16715));
  jor  g16457(.dina(n6369), .dinb(n4415), .dout(n16716));
  jor  g16458(.dina(n4272), .dinb(n6106), .dout(n16717));
  jor  g16459(.dina(n4418), .dinb(n6352), .dout(n16718));
  jor  g16460(.dina(n4420), .dinb(n6372), .dout(n16719));
  jand g16461(.dina(n16719), .dinb(n16718), .dout(n16720));
  jand g16462(.dina(n16720), .dinb(n16717), .dout(n16721));
  jand g16463(.dina(n16721), .dinb(n16716), .dout(n16722));
  jxor g16464(.dina(n16722), .dinb(a38 ), .dout(n16723));
  jxor g16465(.dina(n16723), .dinb(n16715), .dout(n16724));
  jor  g16466(.dina(n16478), .dinb(n16474), .dout(n16725));
  jand g16467(.dina(n16478), .dinb(n16474), .dout(n16726));
  jor  g16468(.dina(n16488), .dinb(n16726), .dout(n16727));
  jand g16469(.dina(n16727), .dinb(n16725), .dout(n16728));
  jxor g16470(.dina(n16728), .dinb(n16724), .dout(n16729));
  jnot g16471(.din(n16729), .dout(n16730));
  jor  g16472(.dina(n7146), .dinb(n3849), .dout(n16731));
  jor  g16473(.dina(n3689), .dinb(n6867), .dout(n16732));
  jor  g16474(.dina(n3852), .dinb(n7129), .dout(n16733));
  jor  g16475(.dina(n3854), .dinb(n7149), .dout(n16734));
  jand g16476(.dina(n16734), .dinb(n16733), .dout(n16735));
  jand g16477(.dina(n16735), .dinb(n16732), .dout(n16736));
  jand g16478(.dina(n16736), .dinb(n16731), .dout(n16737));
  jxor g16479(.dina(n16737), .dinb(a35 ), .dout(n16738));
  jxor g16480(.dina(n16738), .dinb(n16730), .dout(n16739));
  jxor g16481(.dina(n16739), .dinb(n16589), .dout(n16740));
  jxor g16482(.dina(n16740), .dinb(n16585), .dout(n16741));
  jor  g16483(.dina(n16520), .dinb(n16516), .dout(n16742));
  jand g16484(.dina(n16521), .dinb(n16508), .dout(n16743));
  jnot g16485(.din(n16743), .dout(n16744));
  jand g16486(.dina(n16744), .dinb(n16742), .dout(n16745));
  jor  g16487(.dina(n8806), .dinb(n2784), .dout(n16746));
  jor  g16488(.dina(n2661), .dinb(n8231), .dout(n16747));
  jor  g16489(.dina(n2787), .dinb(n8789), .dout(n16748));
  jor  g16490(.dina(n2789), .dinb(n8809), .dout(n16749));
  jand g16491(.dina(n16749), .dinb(n16748), .dout(n16750));
  jand g16492(.dina(n16750), .dinb(n16747), .dout(n16751));
  jand g16493(.dina(n16751), .dinb(n16746), .dout(n16752));
  jxor g16494(.dina(n16752), .dinb(a29 ), .dout(n16753));
  jxor g16495(.dina(n16753), .dinb(n16745), .dout(n16754));
  jxor g16496(.dina(n16754), .dinb(n16741), .dout(n16755));
  jxor g16497(.dina(n16755), .dinb(n16571), .dout(n16756));
  jand g16498(.dina(n16537), .dinb(n16532), .dout(n16757));
  jand g16499(.dina(n16538), .dinb(n16523), .dout(n16758));
  jor  g16500(.dina(n16758), .dinb(n16757), .dout(n16759));
  jnot g16501(.din(n16759), .dout(n16760));
  jor  g16502(.dina(n10961), .dinb(n1939), .dout(n16761));
  jor  g16503(.dina(n1827), .dinb(n10314), .dout(n16762));
  jor  g16504(.dina(n1942), .dinb(n10637), .dout(n16763));
  jor  g16505(.dina(n1944), .dinb(n10964), .dout(n16764));
  jand g16506(.dina(n16764), .dinb(n16763), .dout(n16765));
  jand g16507(.dina(n16765), .dinb(n16762), .dout(n16766));
  jand g16508(.dina(n16766), .dinb(n16761), .dout(n16767));
  jxor g16509(.dina(n16767), .dinb(a23 ), .dout(n16768));
  jxor g16510(.dina(n16768), .dinb(n16760), .dout(n16769));
  jxor g16511(.dina(n16769), .dinb(n16756), .dout(n16770));
  jxor g16512(.dina(n16770), .dinb(n16558), .dout(n16771));
  jand g16513(.dina(n16553), .dinb(n16316), .dout(n16772));
  jand g16514(.dina(n16554), .dinb(n16313), .dout(n16773));
  jor  g16515(.dina(n16773), .dinb(n16772), .dout(n16774));
  jxor g16516(.dina(n16774), .dinb(n16771), .dout(f84 ));
  jand g16517(.dina(n16570), .dinb(n16567), .dout(n16776));
  jand g16518(.dina(n16755), .dinb(n16571), .dout(n16777));
  jor  g16519(.dina(n16777), .dinb(n16776), .dout(n16778));
  jnot g16520(.din(n16778), .dout(n16779));
  jor  g16521(.dina(n10978), .dinb(n1939), .dout(n16780));
  jor  g16522(.dina(n1827), .dinb(n10637), .dout(n16781));
  jor  g16523(.dina(n1942), .dinb(n10964), .dout(n16782));
  jand g16524(.dina(n16782), .dinb(n16781), .dout(n16783));
  jand g16525(.dina(n16783), .dinb(n16780), .dout(n16784));
  jxor g16526(.dina(n16784), .dinb(a23 ), .dout(n16785));
  jxor g16527(.dina(n16785), .dinb(n16779), .dout(n16786));
  jor  g16528(.dina(n10311), .dinb(n2319), .dout(n16787));
  jor  g16529(.dina(n2224), .dinb(n9413), .dout(n16788));
  jor  g16530(.dina(n2322), .dinb(n9725), .dout(n16789));
  jor  g16531(.dina(n2324), .dinb(n10314), .dout(n16790));
  jand g16532(.dina(n16790), .dinb(n16789), .dout(n16791));
  jand g16533(.dina(n16791), .dinb(n16788), .dout(n16792));
  jand g16534(.dina(n16792), .dinb(n16787), .dout(n16793));
  jxor g16535(.dina(n16793), .dinb(a26 ), .dout(n16794));
  jor  g16536(.dina(n16753), .dinb(n16745), .dout(n16795));
  jand g16537(.dina(n16754), .dinb(n16741), .dout(n16796));
  jnot g16538(.din(n16796), .dout(n16797));
  jand g16539(.dina(n16797), .dinb(n16795), .dout(n16798));
  jxor g16540(.dina(n16798), .dinb(n16794), .dout(n16799));
  jand g16541(.dina(n16583), .dinb(n16580), .dout(n16800));
  jnot g16542(.din(n16800), .dout(n16801));
  jor  g16543(.dina(n16740), .dinb(n16585), .dout(n16802));
  jand g16544(.dina(n16802), .dinb(n16801), .dout(n16803));
  jor  g16545(.dina(n9387), .dinb(n2784), .dout(n16804));
  jor  g16546(.dina(n2661), .dinb(n8789), .dout(n16805));
  jor  g16547(.dina(n2787), .dinb(n8809), .dout(n16806));
  jor  g16548(.dina(n2789), .dinb(n9390), .dout(n16807));
  jand g16549(.dina(n16807), .dinb(n16806), .dout(n16808));
  jand g16550(.dina(n16808), .dinb(n16805), .dout(n16809));
  jand g16551(.dina(n16809), .dinb(n16804), .dout(n16810));
  jxor g16552(.dina(n16810), .dinb(a29 ), .dout(n16811));
  jxor g16553(.dina(n16811), .dinb(n16803), .dout(n16812));
  jor  g16554(.dina(n8228), .dinb(n3301), .dout(n16813));
  jor  g16555(.dina(n3136), .dinb(n7683), .dout(n16814));
  jor  g16556(.dina(n3304), .dinb(n7960), .dout(n16815));
  jor  g16557(.dina(n3306), .dinb(n8231), .dout(n16816));
  jand g16558(.dina(n16816), .dinb(n16815), .dout(n16817));
  jand g16559(.dina(n16817), .dinb(n16814), .dout(n16818));
  jand g16560(.dina(n16818), .dinb(n16813), .dout(n16819));
  jxor g16561(.dina(n16819), .dinb(a32 ), .dout(n16820));
  jand g16562(.dina(n16738), .dinb(n16730), .dout(n16821));
  jnot g16563(.din(n16738), .dout(n16822));
  jand g16564(.dina(n16822), .dinb(n16729), .dout(n16823));
  jnot g16565(.din(n16823), .dout(n16824));
  jand g16566(.dina(n16824), .dinb(n16589), .dout(n16825));
  jor  g16567(.dina(n16825), .dinb(n16821), .dout(n16826));
  jxor g16568(.dina(n16826), .dinb(n16820), .dout(n16827));
  jor  g16569(.dina(n16723), .dinb(n16715), .dout(n16828));
  jand g16570(.dina(n16728), .dinb(n16724), .dout(n16829));
  jnot g16571(.din(n16829), .dout(n16830));
  jand g16572(.dina(n16830), .dinb(n16828), .dout(n16831));
  jnot g16573(.din(n16831), .dout(n16832));
  jor  g16574(.dina(n16712), .dinb(n16704), .dout(n16833));
  jand g16575(.dina(n16713), .dinb(n16592), .dout(n16834));
  jnot g16576(.din(n16834), .dout(n16835));
  jand g16577(.dina(n16835), .dinb(n16833), .dout(n16836));
  jnot g16578(.din(n16836), .dout(n16837));
  jor  g16579(.dina(n16701), .dinb(n16693), .dout(n16838));
  jand g16580(.dina(n16702), .dinb(n16595), .dout(n16839));
  jnot g16581(.din(n16839), .dout(n16840));
  jand g16582(.dina(n16840), .dinb(n16838), .dout(n16841));
  jnot g16583(.din(n16841), .dout(n16842));
  jor  g16584(.dina(n16690), .dinb(n16682), .dout(n16843));
  jand g16585(.dina(n16691), .dinb(n16598), .dout(n16844));
  jnot g16586(.din(n16844), .dout(n16845));
  jand g16587(.dina(n16845), .dinb(n16843), .dout(n16846));
  jnot g16588(.din(n16846), .dout(n16847));
  jor  g16589(.dina(n6490), .dinb(n4554), .dout(n16848));
  jor  g16590(.dina(n6262), .dinb(n4340), .dout(n16849));
  jor  g16591(.dina(n6493), .dinb(n4537), .dout(n16850));
  jor  g16592(.dina(n6495), .dinb(n4557), .dout(n16851));
  jand g16593(.dina(n16851), .dinb(n16850), .dout(n16852));
  jand g16594(.dina(n16852), .dinb(n16849), .dout(n16853));
  jand g16595(.dina(n16853), .dinb(n16848), .dout(n16854));
  jxor g16596(.dina(n16854), .dinb(a47 ), .dout(n16855));
  jnot g16597(.din(n16855), .dout(n16856));
  jand g16598(.dina(n16679), .dinb(n16612), .dout(n16857));
  jand g16599(.dina(n16680), .dinb(n16603), .dout(n16858));
  jor  g16600(.dina(n16858), .dinb(n16857), .dout(n16859));
  jand g16601(.dina(n16677), .dinb(n16674), .dout(n16860));
  jand g16602(.dina(n16678), .dinb(n16665), .dout(n16861));
  jor  g16603(.dina(n16861), .dinb(n16860), .dout(n16862));
  jor  g16604(.dina(n16663), .dinb(n16655), .dout(n16863));
  jand g16605(.dina(n16664), .dinb(n16619), .dout(n16864));
  jnot g16606(.din(n16864), .dout(n16865));
  jand g16607(.dina(n16865), .dinb(n16863), .dout(n16866));
  jnot g16608(.din(n16866), .dout(n16867));
  jand g16609(.dina(n16652), .dinb(n16631), .dout(n16868));
  jand g16610(.dina(n16653), .dinb(n16622), .dout(n16869));
  jor  g16611(.dina(n16869), .dinb(n16868), .dout(n16870));
  jor  g16612(.dina(n9891), .dinb(n2556), .dout(n16871));
  jor  g16613(.dina(n9593), .dinb(n2148), .dout(n16872));
  jor  g16614(.dina(n9894), .dinb(n2407), .dout(n16873));
  jor  g16615(.dina(n9896), .dinb(n2559), .dout(n16874));
  jand g16616(.dina(n16874), .dinb(n16873), .dout(n16875));
  jand g16617(.dina(n16875), .dinb(n16872), .dout(n16876));
  jand g16618(.dina(n16876), .dinb(n16871), .dout(n16877));
  jxor g16619(.dina(n16877), .dinb(a59 ), .dout(n16878));
  jnot g16620(.din(n16878), .dout(n16879));
  jor  g16621(.dina(n16650), .dinb(n16642), .dout(n16880));
  jand g16622(.dina(n16651), .dinb(n16636), .dout(n16881));
  jnot g16623(.din(n16881), .dout(n16882));
  jand g16624(.dina(n16882), .dinb(n16880), .dout(n16883));
  jnot g16625(.din(n16883), .dout(n16884));
  jand g16626(.dina(n16639), .dinb(n16540), .dout(n16885));
  jand g16627(.dina(n16640), .dinb(n16418), .dout(n16886));
  jor  g16628(.dina(n16886), .dinb(n16885), .dout(n16887));
  jand g16629(.dina(n10801), .dinb(b22 ), .dout(n16888));
  jand g16630(.dina(n11107), .dinb(b21 ), .dout(n16889));
  jor  g16631(.dina(n16889), .dinb(n16888), .dout(n16890));
  jnot g16632(.din(n16890), .dout(n16891));
  jxor g16633(.dina(n16891), .dinb(n16887), .dout(n16892));
  jnot g16634(.din(n16892), .dout(n16893));
  jor  g16635(.dina(n10806), .dinb(n2007), .dout(n16894));
  jor  g16636(.dina(n10485), .dinb(n1867), .dout(n16895));
  jor  g16637(.dina(n10809), .dinb(n1887), .dout(n16896));
  jor  g16638(.dina(n10811), .dinb(n2010), .dout(n16897));
  jand g16639(.dina(n16897), .dinb(n16896), .dout(n16898));
  jand g16640(.dina(n16898), .dinb(n16895), .dout(n16899));
  jand g16641(.dina(n16899), .dinb(n16894), .dout(n16900));
  jxor g16642(.dina(n16900), .dinb(a62 ), .dout(n16901));
  jxor g16643(.dina(n16901), .dinb(n16893), .dout(n16902));
  jxor g16644(.dina(n16902), .dinb(n16884), .dout(n16903));
  jxor g16645(.dina(n16903), .dinb(n16879), .dout(n16904));
  jxor g16646(.dina(n16904), .dinb(n16870), .dout(n16905));
  jor  g16647(.dina(n8978), .dinb(n3032), .dout(n16906));
  jor  g16648(.dina(n8677), .dinb(n2579), .dout(n16907));
  jor  g16649(.dina(n8981), .dinb(n2870), .dout(n16908));
  jor  g16650(.dina(n8983), .dinb(n3035), .dout(n16909));
  jand g16651(.dina(n16909), .dinb(n16908), .dout(n16910));
  jand g16652(.dina(n16910), .dinb(n16907), .dout(n16911));
  jand g16653(.dina(n16911), .dinb(n16906), .dout(n16912));
  jxor g16654(.dina(n16912), .dinb(a56 ), .dout(n16913));
  jnot g16655(.din(n16913), .dout(n16914));
  jxor g16656(.dina(n16914), .dinb(n16905), .dout(n16915));
  jxor g16657(.dina(n16915), .dinb(n16867), .dout(n16916));
  jor  g16658(.dina(n8125), .dinb(n3400), .dout(n16917));
  jor  g16659(.dina(n7846), .dinb(n3055), .dout(n16918));
  jor  g16660(.dina(n8128), .dinb(n3230), .dout(n16919));
  jor  g16661(.dina(n8130), .dinb(n3403), .dout(n16920));
  jand g16662(.dina(n16920), .dinb(n16919), .dout(n16921));
  jand g16663(.dina(n16921), .dinb(n16918), .dout(n16922));
  jand g16664(.dina(n16922), .dinb(n16917), .dout(n16923));
  jxor g16665(.dina(n16923), .dinb(a53 ), .dout(n16924));
  jnot g16666(.din(n16924), .dout(n16925));
  jxor g16667(.dina(n16925), .dinb(n16916), .dout(n16926));
  jxor g16668(.dina(n16926), .dinb(n16862), .dout(n16927));
  jnot g16669(.din(n16927), .dout(n16928));
  jor  g16670(.dina(n7266), .dinb(n4137), .dout(n16929));
  jor  g16671(.dina(n7021), .dinb(n3588), .dout(n16930));
  jor  g16672(.dina(n7269), .dinb(n3942), .dout(n16931));
  jor  g16673(.dina(n7271), .dinb(n4140), .dout(n16932));
  jand g16674(.dina(n16932), .dinb(n16931), .dout(n16933));
  jand g16675(.dina(n16933), .dinb(n16930), .dout(n16934));
  jand g16676(.dina(n16934), .dinb(n16929), .dout(n16935));
  jxor g16677(.dina(n16935), .dinb(a50 ), .dout(n16936));
  jxor g16678(.dina(n16936), .dinb(n16928), .dout(n16937));
  jxor g16679(.dina(n16937), .dinb(n16859), .dout(n16938));
  jxor g16680(.dina(n16938), .dinb(n16856), .dout(n16939));
  jxor g16681(.dina(n16939), .dinb(n16847), .dout(n16940));
  jor  g16682(.dina(n5405), .dinb(n5739), .dout(n16941));
  jor  g16683(.dina(n5574), .dinb(n4974), .dout(n16942));
  jor  g16684(.dina(n5742), .dinb(n4994), .dout(n16943));
  jor  g16685(.dina(n5744), .dinb(n5408), .dout(n16944));
  jand g16686(.dina(n16944), .dinb(n16943), .dout(n16945));
  jand g16687(.dina(n16945), .dinb(n16942), .dout(n16946));
  jand g16688(.dina(n16946), .dinb(n16941), .dout(n16947));
  jxor g16689(.dina(n16947), .dinb(a44 ), .dout(n16948));
  jnot g16690(.din(n16948), .dout(n16949));
  jxor g16691(.dina(n16949), .dinb(n16940), .dout(n16950));
  jxor g16692(.dina(n16950), .dinb(n16842), .dout(n16951));
  jor  g16693(.dina(n6103), .dinb(n5096), .dout(n16952));
  jor  g16694(.dina(n4904), .dinb(n5428), .dout(n16953));
  jor  g16695(.dina(n5099), .dinb(n5862), .dout(n16954));
  jor  g16696(.dina(n5101), .dinb(n6106), .dout(n16955));
  jand g16697(.dina(n16955), .dinb(n16954), .dout(n16956));
  jand g16698(.dina(n16956), .dinb(n16953), .dout(n16957));
  jand g16699(.dina(n16957), .dinb(n16952), .dout(n16958));
  jxor g16700(.dina(n16958), .dinb(a41 ), .dout(n16959));
  jnot g16701(.din(n16959), .dout(n16960));
  jxor g16702(.dina(n16960), .dinb(n16951), .dout(n16961));
  jxor g16703(.dina(n16961), .dinb(n16837), .dout(n16962));
  jor  g16704(.dina(n6864), .dinb(n4415), .dout(n16963));
  jor  g16705(.dina(n4272), .dinb(n6352), .dout(n16964));
  jor  g16706(.dina(n4418), .dinb(n6372), .dout(n16965));
  jor  g16707(.dina(n4420), .dinb(n6867), .dout(n16966));
  jand g16708(.dina(n16966), .dinb(n16965), .dout(n16967));
  jand g16709(.dina(n16967), .dinb(n16964), .dout(n16968));
  jand g16710(.dina(n16968), .dinb(n16963), .dout(n16969));
  jxor g16711(.dina(n16969), .dinb(a38 ), .dout(n16970));
  jnot g16712(.din(n16970), .dout(n16971));
  jxor g16713(.dina(n16971), .dinb(n16962), .dout(n16972));
  jxor g16714(.dina(n16972), .dinb(n16832), .dout(n16973));
  jor  g16715(.dina(n7408), .dinb(n3849), .dout(n16974));
  jor  g16716(.dina(n3689), .dinb(n7129), .dout(n16975));
  jor  g16717(.dina(n3852), .dinb(n7149), .dout(n16976));
  jor  g16718(.dina(n3854), .dinb(n7411), .dout(n16977));
  jand g16719(.dina(n16977), .dinb(n16976), .dout(n16978));
  jand g16720(.dina(n16978), .dinb(n16975), .dout(n16979));
  jand g16721(.dina(n16979), .dinb(n16974), .dout(n16980));
  jxor g16722(.dina(n16980), .dinb(a35 ), .dout(n16981));
  jnot g16723(.din(n16981), .dout(n16982));
  jxor g16724(.dina(n16982), .dinb(n16973), .dout(n16983));
  jxor g16725(.dina(n16983), .dinb(n16827), .dout(n16984));
  jxor g16726(.dina(n16984), .dinb(n16812), .dout(n16985));
  jxor g16727(.dina(n16985), .dinb(n16799), .dout(n16986));
  jnot g16728(.din(n16986), .dout(n16987));
  jxor g16729(.dina(n16987), .dinb(n16786), .dout(n16988));
  jor  g16730(.dina(n16768), .dinb(n16760), .dout(n16989));
  jand g16731(.dina(n16769), .dinb(n16756), .dout(n16990));
  jnot g16732(.din(n16990), .dout(n16991));
  jand g16733(.dina(n16991), .dinb(n16989), .dout(n16992));
  jxor g16734(.dina(n16992), .dinb(n16988), .dout(n16993));
  jand g16735(.dina(n16770), .dinb(n16558), .dout(n16994));
  jand g16736(.dina(n16774), .dinb(n16771), .dout(n16995));
  jor  g16737(.dina(n16995), .dinb(n16994), .dout(n16996));
  jxor g16738(.dina(n16996), .dinb(n16993), .dout(f85 ));
  jor  g16739(.dina(n16992), .dinb(n16988), .dout(n16998));
  jnot g16740(.din(n16998), .dout(n16999));
  jand g16741(.dina(n16996), .dinb(n16993), .dout(n17000));
  jor  g16742(.dina(n17000), .dinb(n16999), .dout(n17001));
  jor  g16743(.dina(n16798), .dinb(n16794), .dout(n17002));
  jand g16744(.dina(n16985), .dinb(n16799), .dout(n17003));
  jnot g16745(.din(n17003), .dout(n17004));
  jand g16746(.dina(n17004), .dinb(n17002), .dout(n17005));
  jnot g16747(.din(a23 ), .dout(n17006));
  jand g16748(.dina(n11296), .dinb(n1690), .dout(n17007));
  jor  g16749(.dina(n17007), .dinb(n1828), .dout(n17008));
  jand g16750(.dina(n17008), .dinb(b63 ), .dout(n17009));
  jxor g16751(.dina(n17009), .dinb(n17006), .dout(n17010));
  jxor g16752(.dina(n17010), .dinb(n17005), .dout(n17011));
  jor  g16753(.dina(n10634), .dinb(n2319), .dout(n17012));
  jor  g16754(.dina(n2224), .dinb(n9725), .dout(n17013));
  jor  g16755(.dina(n2322), .dinb(n10314), .dout(n17014));
  jor  g16756(.dina(n2324), .dinb(n10637), .dout(n17015));
  jand g16757(.dina(n17015), .dinb(n17014), .dout(n17016));
  jand g16758(.dina(n17016), .dinb(n17013), .dout(n17017));
  jand g16759(.dina(n17017), .dinb(n17012), .dout(n17018));
  jxor g16760(.dina(n17018), .dinb(a26 ), .dout(n17019));
  jor  g16761(.dina(n16811), .dinb(n16803), .dout(n17020));
  jand g16762(.dina(n16984), .dinb(n16812), .dout(n17021));
  jnot g16763(.din(n17021), .dout(n17022));
  jand g16764(.dina(n17022), .dinb(n17020), .dout(n17023));
  jxor g16765(.dina(n17023), .dinb(n17019), .dout(n17024));
  jor  g16766(.dina(n9410), .dinb(n2784), .dout(n17025));
  jor  g16767(.dina(n2661), .dinb(n8809), .dout(n17026));
  jor  g16768(.dina(n2787), .dinb(n9390), .dout(n17027));
  jor  g16769(.dina(n2789), .dinb(n9413), .dout(n17028));
  jand g16770(.dina(n17028), .dinb(n17027), .dout(n17029));
  jand g16771(.dina(n17029), .dinb(n17026), .dout(n17030));
  jand g16772(.dina(n17030), .dinb(n17025), .dout(n17031));
  jxor g16773(.dina(n17031), .dinb(a29 ), .dout(n17032));
  jnot g16774(.din(n17032), .dout(n17033));
  jnot g16775(.din(n16820), .dout(n17034));
  jnot g16776(.din(n16826), .dout(n17035));
  jand g16777(.dina(n17035), .dinb(n17034), .dout(n17036));
  jand g16778(.dina(n16983), .dinb(n16827), .dout(n17037));
  jor  g16779(.dina(n17037), .dinb(n17036), .dout(n17038));
  jxor g16780(.dina(n17038), .dinb(n17033), .dout(n17039));
  jor  g16781(.dina(n8786), .dinb(n3301), .dout(n17040));
  jor  g16782(.dina(n3136), .dinb(n7960), .dout(n17041));
  jor  g16783(.dina(n3304), .dinb(n8231), .dout(n17042));
  jor  g16784(.dina(n3306), .dinb(n8789), .dout(n17043));
  jand g16785(.dina(n17043), .dinb(n17042), .dout(n17044));
  jand g16786(.dina(n17044), .dinb(n17041), .dout(n17045));
  jand g16787(.dina(n17045), .dinb(n17040), .dout(n17046));
  jxor g16788(.dina(n17046), .dinb(a32 ), .dout(n17047));
  jnot g16789(.din(n16972), .dout(n17048));
  jand g16790(.dina(n17048), .dinb(n16831), .dout(n17049));
  jnot g16791(.din(n17049), .dout(n17050));
  jand g16792(.dina(n16972), .dinb(n16832), .dout(n17051));
  jor  g16793(.dina(n16982), .dinb(n17051), .dout(n17052));
  jand g16794(.dina(n17052), .dinb(n17050), .dout(n17053));
  jnot g16795(.din(n17053), .dout(n17054));
  jxor g16796(.dina(n17054), .dinb(n17047), .dout(n17055));
  jor  g16797(.dina(n7680), .dinb(n3849), .dout(n17056));
  jor  g16798(.dina(n3689), .dinb(n7149), .dout(n17057));
  jor  g16799(.dina(n3852), .dinb(n7411), .dout(n17058));
  jor  g16800(.dina(n3854), .dinb(n7683), .dout(n17059));
  jand g16801(.dina(n17059), .dinb(n17058), .dout(n17060));
  jand g16802(.dina(n17060), .dinb(n17057), .dout(n17061));
  jand g16803(.dina(n17061), .dinb(n17056), .dout(n17062));
  jxor g16804(.dina(n17062), .dinb(a35 ), .dout(n17063));
  jnot g16805(.din(n17063), .dout(n17064));
  jor  g16806(.dina(n5425), .dinb(n5739), .dout(n17065));
  jor  g16807(.dina(n5574), .dinb(n4994), .dout(n17066));
  jor  g16808(.dina(n5742), .dinb(n5408), .dout(n17067));
  jor  g16809(.dina(n5744), .dinb(n5428), .dout(n17068));
  jand g16810(.dina(n17068), .dinb(n17067), .dout(n17069));
  jand g16811(.dina(n17069), .dinb(n17066), .dout(n17070));
  jand g16812(.dina(n17070), .dinb(n17065), .dout(n17071));
  jxor g16813(.dina(n17071), .dinb(a44 ), .dout(n17072));
  jnot g16814(.din(n17072), .dout(n17073));
  jand g16815(.dina(n16937), .dinb(n16859), .dout(n17074));
  jand g16816(.dina(n16938), .dinb(n16856), .dout(n17075));
  jor  g16817(.dina(n17075), .dinb(n17074), .dout(n17076));
  jor  g16818(.dina(n6490), .dinb(n4971), .dout(n17077));
  jor  g16819(.dina(n6262), .dinb(n4537), .dout(n17078));
  jor  g16820(.dina(n6493), .dinb(n4557), .dout(n17079));
  jor  g16821(.dina(n6495), .dinb(n4974), .dout(n17080));
  jand g16822(.dina(n17080), .dinb(n17079), .dout(n17081));
  jand g16823(.dina(n17081), .dinb(n17078), .dout(n17082));
  jand g16824(.dina(n17082), .dinb(n17077), .dout(n17083));
  jxor g16825(.dina(n17083), .dinb(a47 ), .dout(n17084));
  jnot g16826(.din(n17084), .dout(n17085));
  jand g16827(.dina(n16926), .dinb(n16862), .dout(n17086));
  jnot g16828(.din(n17086), .dout(n17087));
  jor  g16829(.dina(n16936), .dinb(n16928), .dout(n17088));
  jand g16830(.dina(n17088), .dinb(n17087), .dout(n17089));
  jnot g16831(.din(n17089), .dout(n17090));
  jor  g16832(.dina(n8125), .dinb(n3585), .dout(n17091));
  jor  g16833(.dina(n7846), .dinb(n3230), .dout(n17092));
  jor  g16834(.dina(n8128), .dinb(n3403), .dout(n17093));
  jor  g16835(.dina(n8130), .dinb(n3588), .dout(n17094));
  jand g16836(.dina(n17094), .dinb(n17093), .dout(n17095));
  jand g16837(.dina(n17095), .dinb(n17092), .dout(n17096));
  jand g16838(.dina(n17096), .dinb(n17091), .dout(n17097));
  jxor g16839(.dina(n17097), .dinb(a53 ), .dout(n17098));
  jnot g16840(.din(n17098), .dout(n17099));
  jand g16841(.dina(n16902), .dinb(n16884), .dout(n17100));
  jand g16842(.dina(n16903), .dinb(n16879), .dout(n17101));
  jor  g16843(.dina(n17101), .dinb(n17100), .dout(n17102));
  jand g16844(.dina(n16891), .dinb(n16887), .dout(n17103));
  jnot g16845(.din(n17103), .dout(n17104));
  jor  g16846(.dina(n16901), .dinb(n16893), .dout(n17105));
  jand g16847(.dina(n17105), .dinb(n17104), .dout(n17106));
  jnot g16848(.din(n17106), .dout(n17107));
  jand g16849(.dina(n10801), .dinb(b23 ), .dout(n17108));
  jand g16850(.dina(n11107), .dinb(b22 ), .dout(n17109));
  jor  g16851(.dina(n17109), .dinb(n17108), .dout(n17110));
  jnot g16852(.din(n17110), .dout(n17111));
  jxor g16853(.dina(n17111), .dinb(n16890), .dout(n17112));
  jnot g16854(.din(n17112), .dout(n17113));
  jor  g16855(.dina(n10806), .dinb(n2145), .dout(n17114));
  jor  g16856(.dina(n10485), .dinb(n1887), .dout(n17115));
  jor  g16857(.dina(n10809), .dinb(n2010), .dout(n17116));
  jor  g16858(.dina(n10811), .dinb(n2148), .dout(n17117));
  jand g16859(.dina(n17117), .dinb(n17116), .dout(n17118));
  jand g16860(.dina(n17118), .dinb(n17115), .dout(n17119));
  jand g16861(.dina(n17119), .dinb(n17114), .dout(n17120));
  jxor g16862(.dina(n17120), .dinb(a62 ), .dout(n17121));
  jxor g16863(.dina(n17121), .dinb(n17113), .dout(n17122));
  jxor g16864(.dina(n17122), .dinb(n17107), .dout(n17123));
  jor  g16865(.dina(n9891), .dinb(n2576), .dout(n17124));
  jor  g16866(.dina(n9593), .dinb(n2407), .dout(n17125));
  jor  g16867(.dina(n9894), .dinb(n2559), .dout(n17126));
  jor  g16868(.dina(n9896), .dinb(n2579), .dout(n17127));
  jand g16869(.dina(n17127), .dinb(n17126), .dout(n17128));
  jand g16870(.dina(n17128), .dinb(n17125), .dout(n17129));
  jand g16871(.dina(n17129), .dinb(n17124), .dout(n17130));
  jxor g16872(.dina(n17130), .dinb(a59 ), .dout(n17131));
  jnot g16873(.din(n17131), .dout(n17132));
  jxor g16874(.dina(n17132), .dinb(n17123), .dout(n17133));
  jxor g16875(.dina(n17133), .dinb(n17102), .dout(n17134));
  jnot g16876(.din(n17134), .dout(n17135));
  jor  g16877(.dina(n8978), .dinb(n3052), .dout(n17136));
  jor  g16878(.dina(n8677), .dinb(n2870), .dout(n17137));
  jor  g16879(.dina(n8981), .dinb(n3035), .dout(n17138));
  jor  g16880(.dina(n8983), .dinb(n3055), .dout(n17139));
  jand g16881(.dina(n17139), .dinb(n17138), .dout(n17140));
  jand g16882(.dina(n17140), .dinb(n17137), .dout(n17141));
  jand g16883(.dina(n17141), .dinb(n17136), .dout(n17142));
  jxor g16884(.dina(n17142), .dinb(a56 ), .dout(n17143));
  jxor g16885(.dina(n17143), .dinb(n17135), .dout(n17144));
  jor  g16886(.dina(n16904), .dinb(n16870), .dout(n17145));
  jand g16887(.dina(n16904), .dinb(n16870), .dout(n17146));
  jor  g16888(.dina(n16914), .dinb(n17146), .dout(n17147));
  jand g16889(.dina(n17147), .dinb(n17145), .dout(n17148));
  jxor g16890(.dina(n17148), .dinb(n17144), .dout(n17149));
  jxor g16891(.dina(n17149), .dinb(n17099), .dout(n17150));
  jnot g16892(.din(n16915), .dout(n17151));
  jand g16893(.dina(n17151), .dinb(n16866), .dout(n17152));
  jnot g16894(.din(n17152), .dout(n17153));
  jand g16895(.dina(n16915), .dinb(n16867), .dout(n17154));
  jor  g16896(.dina(n16925), .dinb(n17154), .dout(n17155));
  jand g16897(.dina(n17155), .dinb(n17153), .dout(n17156));
  jxor g16898(.dina(n17156), .dinb(n17150), .dout(n17157));
  jor  g16899(.dina(n7266), .dinb(n4337), .dout(n17158));
  jor  g16900(.dina(n7021), .dinb(n3942), .dout(n17159));
  jor  g16901(.dina(n7269), .dinb(n4140), .dout(n17160));
  jor  g16902(.dina(n7271), .dinb(n4340), .dout(n17161));
  jand g16903(.dina(n17161), .dinb(n17160), .dout(n17162));
  jand g16904(.dina(n17162), .dinb(n17159), .dout(n17163));
  jand g16905(.dina(n17163), .dinb(n17158), .dout(n17164));
  jxor g16906(.dina(n17164), .dinb(a50 ), .dout(n17165));
  jnot g16907(.din(n17165), .dout(n17166));
  jxor g16908(.dina(n17166), .dinb(n17157), .dout(n17167));
  jxor g16909(.dina(n17167), .dinb(n17090), .dout(n17168));
  jxor g16910(.dina(n17168), .dinb(n17085), .dout(n17169));
  jxor g16911(.dina(n17169), .dinb(n17076), .dout(n17170));
  jxor g16912(.dina(n17170), .dinb(n17073), .dout(n17171));
  jor  g16913(.dina(n16939), .dinb(n16847), .dout(n17172));
  jand g16914(.dina(n16939), .dinb(n16847), .dout(n17173));
  jor  g16915(.dina(n16949), .dinb(n17173), .dout(n17174));
  jand g16916(.dina(n17174), .dinb(n17172), .dout(n17175));
  jxor g16917(.dina(n17175), .dinb(n17171), .dout(n17176));
  jor  g16918(.dina(n6349), .dinb(n5096), .dout(n17177));
  jor  g16919(.dina(n4904), .dinb(n5862), .dout(n17178));
  jor  g16920(.dina(n5099), .dinb(n6106), .dout(n17179));
  jor  g16921(.dina(n5101), .dinb(n6352), .dout(n17180));
  jand g16922(.dina(n17180), .dinb(n17179), .dout(n17181));
  jand g16923(.dina(n17181), .dinb(n17178), .dout(n17182));
  jand g16924(.dina(n17182), .dinb(n17177), .dout(n17183));
  jxor g16925(.dina(n17183), .dinb(a41 ), .dout(n17184));
  jnot g16926(.din(n17184), .dout(n17185));
  jxor g16927(.dina(n17185), .dinb(n17176), .dout(n17186));
  jnot g16928(.din(n16950), .dout(n17187));
  jand g16929(.dina(n17187), .dinb(n16841), .dout(n17188));
  jnot g16930(.din(n17188), .dout(n17189));
  jand g16931(.dina(n16950), .dinb(n16842), .dout(n17190));
  jor  g16932(.dina(n16960), .dinb(n17190), .dout(n17191));
  jand g16933(.dina(n17191), .dinb(n17189), .dout(n17192));
  jxor g16934(.dina(n17192), .dinb(n17186), .dout(n17193));
  jnot g16935(.din(n17193), .dout(n17194));
  jor  g16936(.dina(n7126), .dinb(n4415), .dout(n17195));
  jor  g16937(.dina(n4272), .dinb(n6372), .dout(n17196));
  jor  g16938(.dina(n4418), .dinb(n6867), .dout(n17197));
  jor  g16939(.dina(n4420), .dinb(n7129), .dout(n17198));
  jand g16940(.dina(n17198), .dinb(n17197), .dout(n17199));
  jand g16941(.dina(n17199), .dinb(n17196), .dout(n17200));
  jand g16942(.dina(n17200), .dinb(n17195), .dout(n17201));
  jxor g16943(.dina(n17201), .dinb(a38 ), .dout(n17202));
  jxor g16944(.dina(n17202), .dinb(n17194), .dout(n17203));
  jnot g16945(.din(n16961), .dout(n17204));
  jand g16946(.dina(n17204), .dinb(n16836), .dout(n17205));
  jnot g16947(.din(n17205), .dout(n17206));
  jand g16948(.dina(n16961), .dinb(n16837), .dout(n17207));
  jor  g16949(.dina(n16971), .dinb(n17207), .dout(n17208));
  jand g16950(.dina(n17208), .dinb(n17206), .dout(n17209));
  jxor g16951(.dina(n17209), .dinb(n17203), .dout(n17210));
  jxor g16952(.dina(n17210), .dinb(n17064), .dout(n17211));
  jxor g16953(.dina(n17211), .dinb(n17055), .dout(n17212));
  jxor g16954(.dina(n17212), .dinb(n17039), .dout(n17213));
  jxor g16955(.dina(n17213), .dinb(n17024), .dout(n17214));
  jxor g16956(.dina(n17214), .dinb(n17011), .dout(n17215));
  jand g16957(.dina(n16785), .dinb(n16779), .dout(n17216));
  jnot g16958(.din(n17216), .dout(n17217));
  jnot g16959(.din(n16785), .dout(n17218));
  jand g16960(.dina(n17218), .dinb(n16778), .dout(n17219));
  jor  g16961(.dina(n16986), .dinb(n17219), .dout(n17220));
  jand g16962(.dina(n17220), .dinb(n17217), .dout(n17221));
  jxor g16963(.dina(n17221), .dinb(n17215), .dout(n17222));
  jxor g16964(.dina(n17222), .dinb(n17001), .dout(f86 ));
  jand g16965(.dina(n17221), .dinb(n17215), .dout(n17224));
  jand g16966(.dina(n17222), .dinb(n17001), .dout(n17225));
  jor  g16967(.dina(n17225), .dinb(n17224), .dout(n17226));
  jor  g16968(.dina(n17010), .dinb(n17005), .dout(n17227));
  jand g16969(.dina(n17214), .dinb(n17011), .dout(n17228));
  jnot g16970(.din(n17228), .dout(n17229));
  jand g16971(.dina(n17229), .dinb(n17227), .dout(n17230));
  jnot g16972(.din(n17230), .dout(n17231));
  jand g16973(.dina(n17038), .dinb(n17033), .dout(n17232));
  jand g16974(.dina(n17212), .dinb(n17039), .dout(n17233));
  jor  g16975(.dina(n17233), .dinb(n17232), .dout(n17234));
  jnot g16976(.din(n17234), .dout(n17235));
  jor  g16977(.dina(n9722), .dinb(n2784), .dout(n17236));
  jor  g16978(.dina(n2661), .dinb(n9390), .dout(n17237));
  jor  g16979(.dina(n2787), .dinb(n9413), .dout(n17238));
  jor  g16980(.dina(n2789), .dinb(n9725), .dout(n17239));
  jand g16981(.dina(n17239), .dinb(n17238), .dout(n17240));
  jand g16982(.dina(n17240), .dinb(n17237), .dout(n17241));
  jand g16983(.dina(n17241), .dinb(n17236), .dout(n17242));
  jxor g16984(.dina(n17242), .dinb(a29 ), .dout(n17243));
  jxor g16985(.dina(n17243), .dinb(n17235), .dout(n17244));
  jor  g16986(.dina(n8806), .dinb(n3301), .dout(n17245));
  jor  g16987(.dina(n3136), .dinb(n8231), .dout(n17246));
  jor  g16988(.dina(n3304), .dinb(n8789), .dout(n17247));
  jor  g16989(.dina(n3306), .dinb(n8809), .dout(n17248));
  jand g16990(.dina(n17248), .dinb(n17247), .dout(n17249));
  jand g16991(.dina(n17249), .dinb(n17246), .dout(n17250));
  jand g16992(.dina(n17250), .dinb(n17245), .dout(n17251));
  jxor g16993(.dina(n17251), .dinb(a32 ), .dout(n17252));
  jnot g16994(.din(n17252), .dout(n17253));
  jand g16995(.dina(n17054), .dinb(n17047), .dout(n17254));
  jnot g16996(.din(n17254), .dout(n17255));
  jnot g16997(.din(n17047), .dout(n17256));
  jand g16998(.dina(n17053), .dinb(n17256), .dout(n17257));
  jor  g16999(.dina(n17211), .dinb(n17257), .dout(n17258));
  jand g17000(.dina(n17258), .dinb(n17255), .dout(n17259));
  jxor g17001(.dina(n17259), .dinb(n17253), .dout(n17260));
  jor  g17002(.dina(n7957), .dinb(n3849), .dout(n17261));
  jor  g17003(.dina(n3689), .dinb(n7411), .dout(n17262));
  jor  g17004(.dina(n3852), .dinb(n7683), .dout(n17263));
  jor  g17005(.dina(n3854), .dinb(n7960), .dout(n17264));
  jand g17006(.dina(n17264), .dinb(n17263), .dout(n17265));
  jand g17007(.dina(n17265), .dinb(n17262), .dout(n17266));
  jand g17008(.dina(n17266), .dinb(n17261), .dout(n17267));
  jxor g17009(.dina(n17267), .dinb(a35 ), .dout(n17268));
  jand g17010(.dina(n17192), .dinb(n17186), .dout(n17269));
  jnot g17011(.din(n17269), .dout(n17270));
  jor  g17012(.dina(n17202), .dinb(n17194), .dout(n17271));
  jand g17013(.dina(n17271), .dinb(n17270), .dout(n17272));
  jand g17014(.dina(n17169), .dinb(n17076), .dout(n17273));
  jand g17015(.dina(n17170), .dinb(n17073), .dout(n17274));
  jor  g17016(.dina(n17274), .dinb(n17273), .dout(n17275));
  jor  g17017(.dina(n5859), .dinb(n5739), .dout(n17276));
  jor  g17018(.dina(n5574), .dinb(n5408), .dout(n17277));
  jor  g17019(.dina(n5742), .dinb(n5428), .dout(n17278));
  jor  g17020(.dina(n5744), .dinb(n5862), .dout(n17279));
  jand g17021(.dina(n17279), .dinb(n17278), .dout(n17280));
  jand g17022(.dina(n17280), .dinb(n17277), .dout(n17281));
  jand g17023(.dina(n17281), .dinb(n17276), .dout(n17282));
  jxor g17024(.dina(n17282), .dinb(a44 ), .dout(n17283));
  jnot g17025(.din(n17283), .dout(n17284));
  jand g17026(.dina(n17167), .dinb(n17090), .dout(n17285));
  jand g17027(.dina(n17168), .dinb(n17085), .dout(n17286));
  jor  g17028(.dina(n17286), .dinb(n17285), .dout(n17287));
  jand g17029(.dina(n17148), .dinb(n17144), .dout(n17288));
  jand g17030(.dina(n17149), .dinb(n17099), .dout(n17289));
  jor  g17031(.dina(n17289), .dinb(n17288), .dout(n17290));
  jor  g17032(.dina(n9891), .dinb(n2867), .dout(n17291));
  jor  g17033(.dina(n9593), .dinb(n2559), .dout(n17292));
  jor  g17034(.dina(n9894), .dinb(n2579), .dout(n17293));
  jor  g17035(.dina(n9896), .dinb(n2870), .dout(n17294));
  jand g17036(.dina(n17294), .dinb(n17293), .dout(n17295));
  jand g17037(.dina(n17295), .dinb(n17292), .dout(n17296));
  jand g17038(.dina(n17296), .dinb(n17291), .dout(n17297));
  jxor g17039(.dina(n17297), .dinb(a59 ), .dout(n17298));
  jnot g17040(.din(n17298), .dout(n17299));
  jand g17041(.dina(n17111), .dinb(n16890), .dout(n17300));
  jnot g17042(.din(n17300), .dout(n17301));
  jor  g17043(.dina(n17121), .dinb(n17113), .dout(n17302));
  jand g17044(.dina(n17302), .dinb(n17301), .dout(n17303));
  jnot g17045(.din(n17303), .dout(n17304));
  jand g17046(.dina(n10801), .dinb(b24 ), .dout(n17305));
  jand g17047(.dina(n11107), .dinb(b23 ), .dout(n17306));
  jor  g17048(.dina(n17306), .dinb(n17305), .dout(n17307));
  jxor g17049(.dina(n17307), .dinb(n17006), .dout(n17308));
  jxor g17050(.dina(n17308), .dinb(n17110), .dout(n17309));
  jnot g17051(.din(n17309), .dout(n17310));
  jor  g17052(.dina(n10806), .dinb(n2404), .dout(n17311));
  jor  g17053(.dina(n10485), .dinb(n2010), .dout(n17312));
  jor  g17054(.dina(n10809), .dinb(n2148), .dout(n17313));
  jor  g17055(.dina(n10811), .dinb(n2407), .dout(n17314));
  jand g17056(.dina(n17314), .dinb(n17313), .dout(n17315));
  jand g17057(.dina(n17315), .dinb(n17312), .dout(n17316));
  jand g17058(.dina(n17316), .dinb(n17311), .dout(n17317));
  jxor g17059(.dina(n17317), .dinb(a62 ), .dout(n17318));
  jxor g17060(.dina(n17318), .dinb(n17310), .dout(n17319));
  jxor g17061(.dina(n17319), .dinb(n17304), .dout(n17320));
  jxor g17062(.dina(n17320), .dinb(n17299), .dout(n17321));
  jor  g17063(.dina(n17122), .dinb(n17107), .dout(n17322));
  jand g17064(.dina(n17122), .dinb(n17107), .dout(n17323));
  jor  g17065(.dina(n17132), .dinb(n17323), .dout(n17324));
  jand g17066(.dina(n17324), .dinb(n17322), .dout(n17325));
  jxor g17067(.dina(n17325), .dinb(n17321), .dout(n17326));
  jor  g17068(.dina(n8978), .dinb(n3227), .dout(n17327));
  jor  g17069(.dina(n8677), .dinb(n3035), .dout(n17328));
  jor  g17070(.dina(n8981), .dinb(n3055), .dout(n17329));
  jor  g17071(.dina(n8983), .dinb(n3230), .dout(n17330));
  jand g17072(.dina(n17330), .dinb(n17329), .dout(n17331));
  jand g17073(.dina(n17331), .dinb(n17328), .dout(n17332));
  jand g17074(.dina(n17332), .dinb(n17327), .dout(n17333));
  jxor g17075(.dina(n17333), .dinb(a56 ), .dout(n17334));
  jand g17076(.dina(n17133), .dinb(n17102), .dout(n17335));
  jnot g17077(.din(n17335), .dout(n17336));
  jor  g17078(.dina(n17143), .dinb(n17135), .dout(n17337));
  jand g17079(.dina(n17337), .dinb(n17336), .dout(n17338));
  jxor g17080(.dina(n17338), .dinb(n17334), .dout(n17339));
  jxor g17081(.dina(n17339), .dinb(n17326), .dout(n17340));
  jnot g17082(.din(n17340), .dout(n17341));
  jor  g17083(.dina(n8125), .dinb(n3939), .dout(n17342));
  jor  g17084(.dina(n7846), .dinb(n3403), .dout(n17343));
  jor  g17085(.dina(n8128), .dinb(n3588), .dout(n17344));
  jor  g17086(.dina(n8130), .dinb(n3942), .dout(n17345));
  jand g17087(.dina(n17345), .dinb(n17344), .dout(n17346));
  jand g17088(.dina(n17346), .dinb(n17343), .dout(n17347));
  jand g17089(.dina(n17347), .dinb(n17342), .dout(n17348));
  jxor g17090(.dina(n17348), .dinb(a53 ), .dout(n17349));
  jxor g17091(.dina(n17349), .dinb(n17341), .dout(n17350));
  jxor g17092(.dina(n17350), .dinb(n17290), .dout(n17351));
  jnot g17093(.din(n17351), .dout(n17352));
  jor  g17094(.dina(n7266), .dinb(n4534), .dout(n17353));
  jor  g17095(.dina(n7021), .dinb(n4140), .dout(n17354));
  jor  g17096(.dina(n7269), .dinb(n4340), .dout(n17355));
  jor  g17097(.dina(n7271), .dinb(n4537), .dout(n17356));
  jand g17098(.dina(n17356), .dinb(n17355), .dout(n17357));
  jand g17099(.dina(n17357), .dinb(n17354), .dout(n17358));
  jand g17100(.dina(n17358), .dinb(n17353), .dout(n17359));
  jxor g17101(.dina(n17359), .dinb(a50 ), .dout(n17360));
  jxor g17102(.dina(n17360), .dinb(n17352), .dout(n17361));
  jor  g17103(.dina(n17156), .dinb(n17150), .dout(n17362));
  jand g17104(.dina(n17156), .dinb(n17150), .dout(n17363));
  jor  g17105(.dina(n17166), .dinb(n17363), .dout(n17364));
  jand g17106(.dina(n17364), .dinb(n17362), .dout(n17365));
  jxor g17107(.dina(n17365), .dinb(n17361), .dout(n17366));
  jnot g17108(.din(n17366), .dout(n17367));
  jor  g17109(.dina(n6490), .dinb(n4991), .dout(n17368));
  jor  g17110(.dina(n6262), .dinb(n4557), .dout(n17369));
  jor  g17111(.dina(n6493), .dinb(n4974), .dout(n17370));
  jor  g17112(.dina(n6495), .dinb(n4994), .dout(n17371));
  jand g17113(.dina(n17371), .dinb(n17370), .dout(n17372));
  jand g17114(.dina(n17372), .dinb(n17369), .dout(n17373));
  jand g17115(.dina(n17373), .dinb(n17368), .dout(n17374));
  jxor g17116(.dina(n17374), .dinb(a47 ), .dout(n17375));
  jxor g17117(.dina(n17375), .dinb(n17367), .dout(n17376));
  jxor g17118(.dina(n17376), .dinb(n17287), .dout(n17377));
  jxor g17119(.dina(n17377), .dinb(n17284), .dout(n17378));
  jxor g17120(.dina(n17378), .dinb(n17275), .dout(n17379));
  jnot g17121(.din(n17379), .dout(n17380));
  jor  g17122(.dina(n6369), .dinb(n5096), .dout(n17381));
  jor  g17123(.dina(n4904), .dinb(n6106), .dout(n17382));
  jor  g17124(.dina(n5099), .dinb(n6352), .dout(n17383));
  jor  g17125(.dina(n5101), .dinb(n6372), .dout(n17384));
  jand g17126(.dina(n17384), .dinb(n17383), .dout(n17385));
  jand g17127(.dina(n17385), .dinb(n17382), .dout(n17386));
  jand g17128(.dina(n17386), .dinb(n17381), .dout(n17387));
  jxor g17129(.dina(n17387), .dinb(a41 ), .dout(n17388));
  jxor g17130(.dina(n17388), .dinb(n17380), .dout(n17389));
  jor  g17131(.dina(n17175), .dinb(n17171), .dout(n17390));
  jand g17132(.dina(n17175), .dinb(n17171), .dout(n17391));
  jor  g17133(.dina(n17185), .dinb(n17391), .dout(n17392));
  jand g17134(.dina(n17392), .dinb(n17390), .dout(n17393));
  jxor g17135(.dina(n17393), .dinb(n17389), .dout(n17394));
  jnot g17136(.din(n17394), .dout(n17395));
  jor  g17137(.dina(n7146), .dinb(n4415), .dout(n17396));
  jor  g17138(.dina(n4272), .dinb(n6867), .dout(n17397));
  jor  g17139(.dina(n4418), .dinb(n7129), .dout(n17398));
  jor  g17140(.dina(n4420), .dinb(n7149), .dout(n17399));
  jand g17141(.dina(n17399), .dinb(n17398), .dout(n17400));
  jand g17142(.dina(n17400), .dinb(n17397), .dout(n17401));
  jand g17143(.dina(n17401), .dinb(n17396), .dout(n17402));
  jxor g17144(.dina(n17402), .dinb(a38 ), .dout(n17403));
  jxor g17145(.dina(n17403), .dinb(n17395), .dout(n17404));
  jxor g17146(.dina(n17404), .dinb(n17272), .dout(n17405));
  jxor g17147(.dina(n17405), .dinb(n17268), .dout(n17406));
  jor  g17148(.dina(n17209), .dinb(n17203), .dout(n17407));
  jand g17149(.dina(n17209), .dinb(n17203), .dout(n17408));
  jor  g17150(.dina(n17408), .dinb(n17064), .dout(n17409));
  jand g17151(.dina(n17409), .dinb(n17407), .dout(n17410));
  jxor g17152(.dina(n17410), .dinb(n17406), .dout(n17411));
  jxor g17153(.dina(n17411), .dinb(n17260), .dout(n17412));
  jxor g17154(.dina(n17412), .dinb(n17244), .dout(n17413));
  jor  g17155(.dina(n17023), .dinb(n17019), .dout(n17414));
  jand g17156(.dina(n17213), .dinb(n17024), .dout(n17415));
  jnot g17157(.din(n17415), .dout(n17416));
  jand g17158(.dina(n17416), .dinb(n17414), .dout(n17417));
  jor  g17159(.dina(n10961), .dinb(n2319), .dout(n17418));
  jor  g17160(.dina(n2224), .dinb(n10314), .dout(n17419));
  jor  g17161(.dina(n2322), .dinb(n10637), .dout(n17420));
  jor  g17162(.dina(n2324), .dinb(n10964), .dout(n17421));
  jand g17163(.dina(n17421), .dinb(n17420), .dout(n17422));
  jand g17164(.dina(n17422), .dinb(n17419), .dout(n17423));
  jand g17165(.dina(n17423), .dinb(n17418), .dout(n17424));
  jxor g17166(.dina(n17424), .dinb(a26 ), .dout(n17425));
  jxor g17167(.dina(n17425), .dinb(n17417), .dout(n17426));
  jxor g17168(.dina(n17426), .dinb(n17413), .dout(n17427));
  jxor g17169(.dina(n17427), .dinb(n17231), .dout(n17428));
  jxor g17170(.dina(n17428), .dinb(n17226), .dout(f87 ));
  jand g17171(.dina(n17427), .dinb(n17231), .dout(n17430));
  jand g17172(.dina(n17428), .dinb(n17226), .dout(n17431));
  jor  g17173(.dina(n17431), .dinb(n17430), .dout(n17432));
  jor  g17174(.dina(n17425), .dinb(n17417), .dout(n17433));
  jand g17175(.dina(n17426), .dinb(n17413), .dout(n17434));
  jnot g17176(.din(n17434), .dout(n17435));
  jand g17177(.dina(n17435), .dinb(n17433), .dout(n17436));
  jnot g17178(.din(n17436), .dout(n17437));
  jor  g17179(.dina(n17405), .dinb(n17268), .dout(n17438));
  jand g17180(.dina(n17410), .dinb(n17406), .dout(n17439));
  jnot g17181(.din(n17439), .dout(n17440));
  jand g17182(.dina(n17440), .dinb(n17438), .dout(n17441));
  jor  g17183(.dina(n9387), .dinb(n3301), .dout(n17442));
  jor  g17184(.dina(n3136), .dinb(n8789), .dout(n17443));
  jor  g17185(.dina(n3304), .dinb(n8809), .dout(n17444));
  jor  g17186(.dina(n3306), .dinb(n9390), .dout(n17445));
  jand g17187(.dina(n17445), .dinb(n17444), .dout(n17446));
  jand g17188(.dina(n17446), .dinb(n17443), .dout(n17447));
  jand g17189(.dina(n17447), .dinb(n17442), .dout(n17448));
  jxor g17190(.dina(n17448), .dinb(a32 ), .dout(n17449));
  jxor g17191(.dina(n17449), .dinb(n17441), .dout(n17450));
  jor  g17192(.dina(n8228), .dinb(n3849), .dout(n17451));
  jor  g17193(.dina(n3689), .dinb(n7683), .dout(n17452));
  jor  g17194(.dina(n3852), .dinb(n7960), .dout(n17453));
  jor  g17195(.dina(n3854), .dinb(n8231), .dout(n17454));
  jand g17196(.dina(n17454), .dinb(n17453), .dout(n17455));
  jand g17197(.dina(n17455), .dinb(n17452), .dout(n17456));
  jand g17198(.dina(n17456), .dinb(n17451), .dout(n17457));
  jxor g17199(.dina(n17457), .dinb(a35 ), .dout(n17458));
  jnot g17200(.din(n17458), .dout(n17459));
  jor  g17201(.dina(n17388), .dinb(n17380), .dout(n17460));
  jand g17202(.dina(n17393), .dinb(n17389), .dout(n17461));
  jnot g17203(.din(n17461), .dout(n17462));
  jand g17204(.dina(n17462), .dinb(n17460), .dout(n17463));
  jnot g17205(.din(n17463), .dout(n17464));
  jand g17206(.dina(n17377), .dinb(n17284), .dout(n17465));
  jand g17207(.dina(n17378), .dinb(n17275), .dout(n17466));
  jor  g17208(.dina(n17466), .dinb(n17465), .dout(n17467));
  jor  g17209(.dina(n17375), .dinb(n17367), .dout(n17468));
  jand g17210(.dina(n17376), .dinb(n17287), .dout(n17469));
  jnot g17211(.din(n17469), .dout(n17470));
  jand g17212(.dina(n17470), .dinb(n17468), .dout(n17471));
  jnot g17213(.din(n17471), .dout(n17472));
  jor  g17214(.dina(n17360), .dinb(n17352), .dout(n17473));
  jand g17215(.dina(n17365), .dinb(n17361), .dout(n17474));
  jnot g17216(.din(n17474), .dout(n17475));
  jand g17217(.dina(n17475), .dinb(n17473), .dout(n17476));
  jnot g17218(.din(n17476), .dout(n17477));
  jor  g17219(.dina(n7266), .dinb(n4554), .dout(n17478));
  jor  g17220(.dina(n7021), .dinb(n4340), .dout(n17479));
  jor  g17221(.dina(n7269), .dinb(n4537), .dout(n17480));
  jor  g17222(.dina(n7271), .dinb(n4557), .dout(n17481));
  jand g17223(.dina(n17481), .dinb(n17480), .dout(n17482));
  jand g17224(.dina(n17482), .dinb(n17479), .dout(n17483));
  jand g17225(.dina(n17483), .dinb(n17478), .dout(n17484));
  jxor g17226(.dina(n17484), .dinb(a50 ), .dout(n17485));
  jnot g17227(.din(n17485), .dout(n17486));
  jor  g17228(.dina(n17349), .dinb(n17341), .dout(n17487));
  jand g17229(.dina(n17350), .dinb(n17290), .dout(n17488));
  jnot g17230(.din(n17488), .dout(n17489));
  jand g17231(.dina(n17489), .dinb(n17487), .dout(n17490));
  jnot g17232(.din(n17490), .dout(n17491));
  jor  g17233(.dina(n17338), .dinb(n17334), .dout(n17492));
  jand g17234(.dina(n17339), .dinb(n17326), .dout(n17493));
  jnot g17235(.din(n17493), .dout(n17494));
  jand g17236(.dina(n17494), .dinb(n17492), .dout(n17495));
  jnot g17237(.din(n17495), .dout(n17496));
  jand g17238(.dina(n17320), .dinb(n17299), .dout(n17497));
  jand g17239(.dina(n17325), .dinb(n17321), .dout(n17498));
  jor  g17240(.dina(n17498), .dinb(n17497), .dout(n17499));
  jor  g17241(.dina(n17318), .dinb(n17310), .dout(n17500));
  jand g17242(.dina(n17319), .dinb(n17304), .dout(n17501));
  jnot g17243(.din(n17501), .dout(n17502));
  jand g17244(.dina(n17502), .dinb(n17500), .dout(n17503));
  jnot g17245(.din(n17503), .dout(n17504));
  jand g17246(.dina(n17307), .dinb(n17006), .dout(n17505));
  jand g17247(.dina(n17308), .dinb(n17110), .dout(n17506));
  jor  g17248(.dina(n17506), .dinb(n17505), .dout(n17507));
  jand g17249(.dina(n10801), .dinb(b25 ), .dout(n17508));
  jand g17250(.dina(n11107), .dinb(b24 ), .dout(n17509));
  jor  g17251(.dina(n17509), .dinb(n17508), .dout(n17510));
  jnot g17252(.din(n17510), .dout(n17511));
  jxor g17253(.dina(n17511), .dinb(n17507), .dout(n17512));
  jnot g17254(.din(n17512), .dout(n17513));
  jor  g17255(.dina(n10806), .dinb(n2556), .dout(n17514));
  jor  g17256(.dina(n10485), .dinb(n2148), .dout(n17515));
  jor  g17257(.dina(n10809), .dinb(n2407), .dout(n17516));
  jor  g17258(.dina(n10811), .dinb(n2559), .dout(n17517));
  jand g17259(.dina(n17517), .dinb(n17516), .dout(n17518));
  jand g17260(.dina(n17518), .dinb(n17515), .dout(n17519));
  jand g17261(.dina(n17519), .dinb(n17514), .dout(n17520));
  jxor g17262(.dina(n17520), .dinb(a62 ), .dout(n17521));
  jxor g17263(.dina(n17521), .dinb(n17513), .dout(n17522));
  jxor g17264(.dina(n17522), .dinb(n17504), .dout(n17523));
  jor  g17265(.dina(n9891), .dinb(n3032), .dout(n17524));
  jor  g17266(.dina(n9593), .dinb(n2579), .dout(n17525));
  jor  g17267(.dina(n9894), .dinb(n2870), .dout(n17526));
  jor  g17268(.dina(n9896), .dinb(n3035), .dout(n17527));
  jand g17269(.dina(n17527), .dinb(n17526), .dout(n17528));
  jand g17270(.dina(n17528), .dinb(n17525), .dout(n17529));
  jand g17271(.dina(n17529), .dinb(n17524), .dout(n17530));
  jxor g17272(.dina(n17530), .dinb(a59 ), .dout(n17531));
  jnot g17273(.din(n17531), .dout(n17532));
  jxor g17274(.dina(n17532), .dinb(n17523), .dout(n17533));
  jxor g17275(.dina(n17533), .dinb(n17499), .dout(n17534));
  jor  g17276(.dina(n8978), .dinb(n3400), .dout(n17535));
  jor  g17277(.dina(n8677), .dinb(n3055), .dout(n17536));
  jor  g17278(.dina(n8981), .dinb(n3230), .dout(n17537));
  jor  g17279(.dina(n8983), .dinb(n3403), .dout(n17538));
  jand g17280(.dina(n17538), .dinb(n17537), .dout(n17539));
  jand g17281(.dina(n17539), .dinb(n17536), .dout(n17540));
  jand g17282(.dina(n17540), .dinb(n17535), .dout(n17541));
  jxor g17283(.dina(n17541), .dinb(a56 ), .dout(n17542));
  jnot g17284(.din(n17542), .dout(n17543));
  jxor g17285(.dina(n17543), .dinb(n17534), .dout(n17544));
  jxor g17286(.dina(n17544), .dinb(n17496), .dout(n17545));
  jnot g17287(.din(n17545), .dout(n17546));
  jor  g17288(.dina(n8125), .dinb(n4137), .dout(n17547));
  jor  g17289(.dina(n7846), .dinb(n3588), .dout(n17548));
  jor  g17290(.dina(n8128), .dinb(n3942), .dout(n17549));
  jor  g17291(.dina(n8130), .dinb(n4140), .dout(n17550));
  jand g17292(.dina(n17550), .dinb(n17549), .dout(n17551));
  jand g17293(.dina(n17551), .dinb(n17548), .dout(n17552));
  jand g17294(.dina(n17552), .dinb(n17547), .dout(n17553));
  jxor g17295(.dina(n17553), .dinb(a53 ), .dout(n17554));
  jxor g17296(.dina(n17554), .dinb(n17546), .dout(n17555));
  jxor g17297(.dina(n17555), .dinb(n17491), .dout(n17556));
  jxor g17298(.dina(n17556), .dinb(n17486), .dout(n17557));
  jxor g17299(.dina(n17557), .dinb(n17477), .dout(n17558));
  jor  g17300(.dina(n6490), .dinb(n5405), .dout(n17559));
  jor  g17301(.dina(n6262), .dinb(n4974), .dout(n17560));
  jor  g17302(.dina(n6493), .dinb(n4994), .dout(n17561));
  jor  g17303(.dina(n6495), .dinb(n5408), .dout(n17562));
  jand g17304(.dina(n17562), .dinb(n17561), .dout(n17563));
  jand g17305(.dina(n17563), .dinb(n17560), .dout(n17564));
  jand g17306(.dina(n17564), .dinb(n17559), .dout(n17565));
  jxor g17307(.dina(n17565), .dinb(a47 ), .dout(n17566));
  jnot g17308(.din(n17566), .dout(n17567));
  jxor g17309(.dina(n17567), .dinb(n17558), .dout(n17568));
  jxor g17310(.dina(n17568), .dinb(n17472), .dout(n17569));
  jor  g17311(.dina(n6103), .dinb(n5739), .dout(n17570));
  jor  g17312(.dina(n5574), .dinb(n5428), .dout(n17571));
  jor  g17313(.dina(n5742), .dinb(n5862), .dout(n17572));
  jor  g17314(.dina(n5744), .dinb(n6106), .dout(n17573));
  jand g17315(.dina(n17573), .dinb(n17572), .dout(n17574));
  jand g17316(.dina(n17574), .dinb(n17571), .dout(n17575));
  jand g17317(.dina(n17575), .dinb(n17570), .dout(n17576));
  jxor g17318(.dina(n17576), .dinb(a44 ), .dout(n17577));
  jnot g17319(.din(n17577), .dout(n17578));
  jxor g17320(.dina(n17578), .dinb(n17569), .dout(n17579));
  jxor g17321(.dina(n17579), .dinb(n17467), .dout(n17580));
  jor  g17322(.dina(n6864), .dinb(n5096), .dout(n17581));
  jor  g17323(.dina(n4904), .dinb(n6352), .dout(n17582));
  jor  g17324(.dina(n5099), .dinb(n6372), .dout(n17583));
  jor  g17325(.dina(n5101), .dinb(n6867), .dout(n17584));
  jand g17326(.dina(n17584), .dinb(n17583), .dout(n17585));
  jand g17327(.dina(n17585), .dinb(n17582), .dout(n17586));
  jand g17328(.dina(n17586), .dinb(n17581), .dout(n17587));
  jxor g17329(.dina(n17587), .dinb(a41 ), .dout(n17588));
  jnot g17330(.din(n17588), .dout(n17589));
  jxor g17331(.dina(n17589), .dinb(n17580), .dout(n17590));
  jxor g17332(.dina(n17590), .dinb(n17464), .dout(n17591));
  jor  g17333(.dina(n7408), .dinb(n4415), .dout(n17592));
  jor  g17334(.dina(n4272), .dinb(n7129), .dout(n17593));
  jor  g17335(.dina(n4418), .dinb(n7149), .dout(n17594));
  jor  g17336(.dina(n4420), .dinb(n7411), .dout(n17595));
  jand g17337(.dina(n17595), .dinb(n17594), .dout(n17596));
  jand g17338(.dina(n17596), .dinb(n17593), .dout(n17597));
  jand g17339(.dina(n17597), .dinb(n17592), .dout(n17598));
  jxor g17340(.dina(n17598), .dinb(a38 ), .dout(n17599));
  jnot g17341(.din(n17599), .dout(n17600));
  jxor g17342(.dina(n17600), .dinb(n17591), .dout(n17601));
  jand g17343(.dina(n17403), .dinb(n17395), .dout(n17602));
  jnot g17344(.din(n17403), .dout(n17603));
  jand g17345(.dina(n17603), .dinb(n17394), .dout(n17604));
  jnot g17346(.din(n17604), .dout(n17605));
  jand g17347(.dina(n17605), .dinb(n17272), .dout(n17606));
  jor  g17348(.dina(n17606), .dinb(n17602), .dout(n17607));
  jnot g17349(.din(n17607), .dout(n17608));
  jxor g17350(.dina(n17608), .dinb(n17601), .dout(n17609));
  jxor g17351(.dina(n17609), .dinb(n17459), .dout(n17610));
  jxor g17352(.dina(n17610), .dinb(n17450), .dout(n17611));
  jor  g17353(.dina(n10311), .dinb(n2784), .dout(n17612));
  jor  g17354(.dina(n2661), .dinb(n9413), .dout(n17613));
  jor  g17355(.dina(n2787), .dinb(n9725), .dout(n17614));
  jor  g17356(.dina(n2789), .dinb(n10314), .dout(n17615));
  jand g17357(.dina(n17615), .dinb(n17614), .dout(n17616));
  jand g17358(.dina(n17616), .dinb(n17613), .dout(n17617));
  jand g17359(.dina(n17617), .dinb(n17612), .dout(n17618));
  jxor g17360(.dina(n17618), .dinb(a29 ), .dout(n17619));
  jnot g17361(.din(n17619), .dout(n17620));
  jand g17362(.dina(n17259), .dinb(n17253), .dout(n17621));
  jand g17363(.dina(n17411), .dinb(n17260), .dout(n17622));
  jor  g17364(.dina(n17622), .dinb(n17621), .dout(n17623));
  jxor g17365(.dina(n17623), .dinb(n17620), .dout(n17624));
  jxor g17366(.dina(n17624), .dinb(n17611), .dout(n17625));
  jor  g17367(.dina(n17243), .dinb(n17235), .dout(n17626));
  jand g17368(.dina(n17412), .dinb(n17244), .dout(n17627));
  jnot g17369(.din(n17627), .dout(n17628));
  jand g17370(.dina(n17628), .dinb(n17626), .dout(n17629));
  jor  g17371(.dina(n10978), .dinb(n2319), .dout(n17630));
  jor  g17372(.dina(n2224), .dinb(n10637), .dout(n17631));
  jor  g17373(.dina(n2322), .dinb(n10964), .dout(n17632));
  jand g17374(.dina(n17632), .dinb(n17631), .dout(n17633));
  jand g17375(.dina(n17633), .dinb(n17630), .dout(n17634));
  jxor g17376(.dina(n17634), .dinb(a26 ), .dout(n17635));
  jxor g17377(.dina(n17635), .dinb(n17629), .dout(n17636));
  jxor g17378(.dina(n17636), .dinb(n17625), .dout(n17637));
  jxor g17379(.dina(n17637), .dinb(n17437), .dout(n17638));
  jxor g17380(.dina(n17638), .dinb(n17432), .dout(f88 ));
  jand g17381(.dina(n17637), .dinb(n17437), .dout(n17640));
  jand g17382(.dina(n17638), .dinb(n17432), .dout(n17641));
  jor  g17383(.dina(n17641), .dinb(n17640), .dout(n17642));
  jor  g17384(.dina(n17635), .dinb(n17629), .dout(n17643));
  jand g17385(.dina(n17636), .dinb(n17625), .dout(n17644));
  jnot g17386(.din(n17644), .dout(n17645));
  jand g17387(.dina(n17645), .dinb(n17643), .dout(n17646));
  jnot g17388(.din(n17646), .dout(n17647));
  jor  g17389(.dina(n10634), .dinb(n2784), .dout(n17648));
  jor  g17390(.dina(n2661), .dinb(n9725), .dout(n17649));
  jor  g17391(.dina(n2787), .dinb(n10314), .dout(n17650));
  jor  g17392(.dina(n2789), .dinb(n10637), .dout(n17651));
  jand g17393(.dina(n17651), .dinb(n17650), .dout(n17652));
  jand g17394(.dina(n17652), .dinb(n17649), .dout(n17653));
  jand g17395(.dina(n17653), .dinb(n17648), .dout(n17654));
  jxor g17396(.dina(n17654), .dinb(a29 ), .dout(n17655));
  jor  g17397(.dina(n17449), .dinb(n17441), .dout(n17656));
  jand g17398(.dina(n17610), .dinb(n17450), .dout(n17657));
  jnot g17399(.din(n17657), .dout(n17658));
  jand g17400(.dina(n17658), .dinb(n17656), .dout(n17659));
  jxor g17401(.dina(n17659), .dinb(n17655), .dout(n17660));
  jor  g17402(.dina(n9410), .dinb(n3301), .dout(n17661));
  jor  g17403(.dina(n3136), .dinb(n8809), .dout(n17662));
  jor  g17404(.dina(n3304), .dinb(n9390), .dout(n17663));
  jor  g17405(.dina(n3306), .dinb(n9413), .dout(n17664));
  jand g17406(.dina(n17664), .dinb(n17663), .dout(n17665));
  jand g17407(.dina(n17665), .dinb(n17662), .dout(n17666));
  jand g17408(.dina(n17666), .dinb(n17661), .dout(n17667));
  jxor g17409(.dina(n17667), .dinb(a32 ), .dout(n17668));
  jand g17410(.dina(n17608), .dinb(n17601), .dout(n17669));
  jand g17411(.dina(n17609), .dinb(n17459), .dout(n17670));
  jor  g17412(.dina(n17670), .dinb(n17669), .dout(n17671));
  jnot g17413(.din(n17671), .dout(n17672));
  jxor g17414(.dina(n17672), .dinb(n17668), .dout(n17673));
  jor  g17415(.dina(n8786), .dinb(n3849), .dout(n17674));
  jor  g17416(.dina(n3689), .dinb(n7960), .dout(n17675));
  jor  g17417(.dina(n3852), .dinb(n8231), .dout(n17676));
  jor  g17418(.dina(n3854), .dinb(n8789), .dout(n17677));
  jand g17419(.dina(n17677), .dinb(n17676), .dout(n17678));
  jand g17420(.dina(n17678), .dinb(n17675), .dout(n17679));
  jand g17421(.dina(n17679), .dinb(n17674), .dout(n17680));
  jxor g17422(.dina(n17680), .dinb(a35 ), .dout(n17681));
  jnot g17423(.din(n17681), .dout(n17682));
  jor  g17424(.dina(n7680), .dinb(n4415), .dout(n17683));
  jor  g17425(.dina(n4272), .dinb(n7149), .dout(n17684));
  jor  g17426(.dina(n4418), .dinb(n7411), .dout(n17685));
  jor  g17427(.dina(n4420), .dinb(n7683), .dout(n17686));
  jand g17428(.dina(n17686), .dinb(n17685), .dout(n17687));
  jand g17429(.dina(n17687), .dinb(n17684), .dout(n17688));
  jand g17430(.dina(n17688), .dinb(n17683), .dout(n17689));
  jxor g17431(.dina(n17689), .dinb(a38 ), .dout(n17690));
  jnot g17432(.din(n17690), .dout(n17691));
  jor  g17433(.dina(n6490), .dinb(n5425), .dout(n17692));
  jor  g17434(.dina(n6262), .dinb(n4994), .dout(n17693));
  jor  g17435(.dina(n6493), .dinb(n5408), .dout(n17694));
  jor  g17436(.dina(n6495), .dinb(n5428), .dout(n17695));
  jand g17437(.dina(n17695), .dinb(n17694), .dout(n17696));
  jand g17438(.dina(n17696), .dinb(n17693), .dout(n17697));
  jand g17439(.dina(n17697), .dinb(n17692), .dout(n17698));
  jxor g17440(.dina(n17698), .dinb(a47 ), .dout(n17699));
  jnot g17441(.din(n17699), .dout(n17700));
  jand g17442(.dina(n17555), .dinb(n17491), .dout(n17701));
  jand g17443(.dina(n17556), .dinb(n17486), .dout(n17702));
  jor  g17444(.dina(n17702), .dinb(n17701), .dout(n17703));
  jor  g17445(.dina(n7266), .dinb(n4971), .dout(n17704));
  jor  g17446(.dina(n7021), .dinb(n4537), .dout(n17705));
  jor  g17447(.dina(n7269), .dinb(n4557), .dout(n17706));
  jor  g17448(.dina(n7271), .dinb(n4974), .dout(n17707));
  jand g17449(.dina(n17707), .dinb(n17706), .dout(n17708));
  jand g17450(.dina(n17708), .dinb(n17705), .dout(n17709));
  jand g17451(.dina(n17709), .dinb(n17704), .dout(n17710));
  jxor g17452(.dina(n17710), .dinb(a50 ), .dout(n17711));
  jnot g17453(.din(n17711), .dout(n17712));
  jand g17454(.dina(n17544), .dinb(n17496), .dout(n17713));
  jnot g17455(.din(n17713), .dout(n17714));
  jor  g17456(.dina(n17554), .dinb(n17546), .dout(n17715));
  jand g17457(.dina(n17715), .dinb(n17714), .dout(n17716));
  jnot g17458(.din(n17716), .dout(n17717));
  jor  g17459(.dina(n8978), .dinb(n3585), .dout(n17718));
  jor  g17460(.dina(n8677), .dinb(n3230), .dout(n17719));
  jor  g17461(.dina(n8981), .dinb(n3403), .dout(n17720));
  jor  g17462(.dina(n8983), .dinb(n3588), .dout(n17721));
  jand g17463(.dina(n17721), .dinb(n17720), .dout(n17722));
  jand g17464(.dina(n17722), .dinb(n17719), .dout(n17723));
  jand g17465(.dina(n17723), .dinb(n17718), .dout(n17724));
  jxor g17466(.dina(n17724), .dinb(a56 ), .dout(n17725));
  jnot g17467(.din(n17725), .dout(n17726));
  jor  g17468(.dina(n9891), .dinb(n3052), .dout(n17727));
  jor  g17469(.dina(n9593), .dinb(n2870), .dout(n17728));
  jor  g17470(.dina(n9894), .dinb(n3035), .dout(n17729));
  jor  g17471(.dina(n9896), .dinb(n3055), .dout(n17730));
  jand g17472(.dina(n17730), .dinb(n17729), .dout(n17731));
  jand g17473(.dina(n17731), .dinb(n17728), .dout(n17732));
  jand g17474(.dina(n17732), .dinb(n17727), .dout(n17733));
  jxor g17475(.dina(n17733), .dinb(a59 ), .dout(n17734));
  jnot g17476(.din(n17734), .dout(n17735));
  jand g17477(.dina(n17511), .dinb(n17507), .dout(n17736));
  jnot g17478(.din(n17736), .dout(n17737));
  jor  g17479(.dina(n17521), .dinb(n17513), .dout(n17738));
  jand g17480(.dina(n17738), .dinb(n17737), .dout(n17739));
  jnot g17481(.din(n17739), .dout(n17740));
  jand g17482(.dina(n10801), .dinb(b26 ), .dout(n17741));
  jand g17483(.dina(n11107), .dinb(b25 ), .dout(n17742));
  jor  g17484(.dina(n17742), .dinb(n17741), .dout(n17743));
  jnot g17485(.din(n17743), .dout(n17744));
  jxor g17486(.dina(n17744), .dinb(n17510), .dout(n17745));
  jnot g17487(.din(n17745), .dout(n17746));
  jor  g17488(.dina(n10806), .dinb(n2576), .dout(n17747));
  jor  g17489(.dina(n10485), .dinb(n2407), .dout(n17748));
  jor  g17490(.dina(n10809), .dinb(n2559), .dout(n17749));
  jor  g17491(.dina(n10811), .dinb(n2579), .dout(n17750));
  jand g17492(.dina(n17750), .dinb(n17749), .dout(n17751));
  jand g17493(.dina(n17751), .dinb(n17748), .dout(n17752));
  jand g17494(.dina(n17752), .dinb(n17747), .dout(n17753));
  jxor g17495(.dina(n17753), .dinb(a62 ), .dout(n17754));
  jxor g17496(.dina(n17754), .dinb(n17746), .dout(n17755));
  jxor g17497(.dina(n17755), .dinb(n17740), .dout(n17756));
  jxor g17498(.dina(n17756), .dinb(n17735), .dout(n17757));
  jor  g17499(.dina(n17522), .dinb(n17504), .dout(n17758));
  jand g17500(.dina(n17522), .dinb(n17504), .dout(n17759));
  jor  g17501(.dina(n17532), .dinb(n17759), .dout(n17760));
  jand g17502(.dina(n17760), .dinb(n17758), .dout(n17761));
  jxor g17503(.dina(n17761), .dinb(n17757), .dout(n17762));
  jxor g17504(.dina(n17762), .dinb(n17726), .dout(n17763));
  jnot g17505(.din(n17499), .dout(n17764));
  jnot g17506(.din(n17533), .dout(n17765));
  jand g17507(.dina(n17765), .dinb(n17764), .dout(n17766));
  jnot g17508(.din(n17766), .dout(n17767));
  jand g17509(.dina(n17533), .dinb(n17499), .dout(n17768));
  jor  g17510(.dina(n17543), .dinb(n17768), .dout(n17769));
  jand g17511(.dina(n17769), .dinb(n17767), .dout(n17770));
  jxor g17512(.dina(n17770), .dinb(n17763), .dout(n17771));
  jor  g17513(.dina(n8125), .dinb(n4337), .dout(n17772));
  jor  g17514(.dina(n7846), .dinb(n3942), .dout(n17773));
  jor  g17515(.dina(n8128), .dinb(n4140), .dout(n17774));
  jor  g17516(.dina(n8130), .dinb(n4340), .dout(n17775));
  jand g17517(.dina(n17775), .dinb(n17774), .dout(n17776));
  jand g17518(.dina(n17776), .dinb(n17773), .dout(n17777));
  jand g17519(.dina(n17777), .dinb(n17772), .dout(n17778));
  jxor g17520(.dina(n17778), .dinb(a53 ), .dout(n17779));
  jnot g17521(.din(n17779), .dout(n17780));
  jxor g17522(.dina(n17780), .dinb(n17771), .dout(n17781));
  jxor g17523(.dina(n17781), .dinb(n17717), .dout(n17782));
  jxor g17524(.dina(n17782), .dinb(n17712), .dout(n17783));
  jxor g17525(.dina(n17783), .dinb(n17703), .dout(n17784));
  jxor g17526(.dina(n17784), .dinb(n17700), .dout(n17785));
  jor  g17527(.dina(n17557), .dinb(n17477), .dout(n17786));
  jand g17528(.dina(n17557), .dinb(n17477), .dout(n17787));
  jor  g17529(.dina(n17567), .dinb(n17787), .dout(n17788));
  jand g17530(.dina(n17788), .dinb(n17786), .dout(n17789));
  jxor g17531(.dina(n17789), .dinb(n17785), .dout(n17790));
  jor  g17532(.dina(n6349), .dinb(n5739), .dout(n17791));
  jor  g17533(.dina(n5574), .dinb(n5862), .dout(n17792));
  jor  g17534(.dina(n5742), .dinb(n6106), .dout(n17793));
  jor  g17535(.dina(n5744), .dinb(n6352), .dout(n17794));
  jand g17536(.dina(n17794), .dinb(n17793), .dout(n17795));
  jand g17537(.dina(n17795), .dinb(n17792), .dout(n17796));
  jand g17538(.dina(n17796), .dinb(n17791), .dout(n17797));
  jxor g17539(.dina(n17797), .dinb(a44 ), .dout(n17798));
  jnot g17540(.din(n17798), .dout(n17799));
  jxor g17541(.dina(n17799), .dinb(n17790), .dout(n17800));
  jnot g17542(.din(n17568), .dout(n17801));
  jand g17543(.dina(n17801), .dinb(n17471), .dout(n17802));
  jnot g17544(.din(n17802), .dout(n17803));
  jand g17545(.dina(n17568), .dinb(n17472), .dout(n17804));
  jor  g17546(.dina(n17578), .dinb(n17804), .dout(n17805));
  jand g17547(.dina(n17805), .dinb(n17803), .dout(n17806));
  jxor g17548(.dina(n17806), .dinb(n17800), .dout(n17807));
  jnot g17549(.din(n17807), .dout(n17808));
  jor  g17550(.dina(n7126), .dinb(n5096), .dout(n17809));
  jor  g17551(.dina(n4904), .dinb(n6372), .dout(n17810));
  jor  g17552(.dina(n5099), .dinb(n6867), .dout(n17811));
  jor  g17553(.dina(n5101), .dinb(n7129), .dout(n17812));
  jand g17554(.dina(n17812), .dinb(n17811), .dout(n17813));
  jand g17555(.dina(n17813), .dinb(n17810), .dout(n17814));
  jand g17556(.dina(n17814), .dinb(n17809), .dout(n17815));
  jxor g17557(.dina(n17815), .dinb(a41 ), .dout(n17816));
  jxor g17558(.dina(n17816), .dinb(n17808), .dout(n17817));
  jnot g17559(.din(n17467), .dout(n17818));
  jnot g17560(.din(n17579), .dout(n17819));
  jand g17561(.dina(n17819), .dinb(n17818), .dout(n17820));
  jnot g17562(.din(n17820), .dout(n17821));
  jand g17563(.dina(n17579), .dinb(n17467), .dout(n17822));
  jor  g17564(.dina(n17589), .dinb(n17822), .dout(n17823));
  jand g17565(.dina(n17823), .dinb(n17821), .dout(n17824));
  jxor g17566(.dina(n17824), .dinb(n17817), .dout(n17825));
  jxor g17567(.dina(n17825), .dinb(n17691), .dout(n17826));
  jnot g17568(.din(n17590), .dout(n17827));
  jand g17569(.dina(n17827), .dinb(n17463), .dout(n17828));
  jnot g17570(.din(n17828), .dout(n17829));
  jand g17571(.dina(n17590), .dinb(n17464), .dout(n17830));
  jor  g17572(.dina(n17600), .dinb(n17830), .dout(n17831));
  jand g17573(.dina(n17831), .dinb(n17829), .dout(n17832));
  jxor g17574(.dina(n17832), .dinb(n17826), .dout(n17833));
  jxor g17575(.dina(n17833), .dinb(n17682), .dout(n17834));
  jxor g17576(.dina(n17834), .dinb(n17673), .dout(n17835));
  jxor g17577(.dina(n17835), .dinb(n17660), .dout(n17836));
  jand g17578(.dina(n17623), .dinb(n17620), .dout(n17837));
  jand g17579(.dina(n17624), .dinb(n17611), .dout(n17838));
  jor  g17580(.dina(n17838), .dinb(n17837), .dout(n17839));
  jnot g17581(.din(n17839), .dout(n17840));
  jnot g17582(.din(a26 ), .dout(n17841));
  jand g17583(.dina(n11296), .dinb(n2076), .dout(n17842));
  jor  g17584(.dina(n17842), .dinb(n2225), .dout(n17843));
  jand g17585(.dina(n17843), .dinb(b63 ), .dout(n17844));
  jxor g17586(.dina(n17844), .dinb(n17841), .dout(n17845));
  jxor g17587(.dina(n17845), .dinb(n17840), .dout(n17846));
  jxor g17588(.dina(n17846), .dinb(n17836), .dout(n17847));
  jxor g17589(.dina(n17847), .dinb(n17647), .dout(n17848));
  jxor g17590(.dina(n17848), .dinb(n17642), .dout(f89 ));
  jor  g17591(.dina(n17845), .dinb(n17840), .dout(n17850));
  jand g17592(.dina(n17846), .dinb(n17836), .dout(n17851));
  jnot g17593(.din(n17851), .dout(n17852));
  jand g17594(.dina(n17852), .dinb(n17850), .dout(n17853));
  jnot g17595(.din(n17853), .dout(n17854));
  jand g17596(.dina(n17824), .dinb(n17817), .dout(n17855));
  jand g17597(.dina(n17825), .dinb(n17691), .dout(n17856));
  jor  g17598(.dina(n17856), .dinb(n17855), .dout(n17857));
  jor  g17599(.dina(n7957), .dinb(n4415), .dout(n17858));
  jor  g17600(.dina(n4272), .dinb(n7411), .dout(n17859));
  jor  g17601(.dina(n4418), .dinb(n7683), .dout(n17860));
  jor  g17602(.dina(n4420), .dinb(n7960), .dout(n17861));
  jand g17603(.dina(n17861), .dinb(n17860), .dout(n17862));
  jand g17604(.dina(n17862), .dinb(n17859), .dout(n17863));
  jand g17605(.dina(n17863), .dinb(n17858), .dout(n17864));
  jxor g17606(.dina(n17864), .dinb(a38 ), .dout(n17865));
  jand g17607(.dina(n17806), .dinb(n17800), .dout(n17866));
  jnot g17608(.din(n17866), .dout(n17867));
  jor  g17609(.dina(n17816), .dinb(n17808), .dout(n17868));
  jand g17610(.dina(n17868), .dinb(n17867), .dout(n17869));
  jand g17611(.dina(n17783), .dinb(n17703), .dout(n17870));
  jand g17612(.dina(n17784), .dinb(n17700), .dout(n17871));
  jor  g17613(.dina(n17871), .dinb(n17870), .dout(n17872));
  jor  g17614(.dina(n6490), .dinb(n5859), .dout(n17873));
  jor  g17615(.dina(n6262), .dinb(n5408), .dout(n17874));
  jor  g17616(.dina(n6493), .dinb(n5428), .dout(n17875));
  jor  g17617(.dina(n6495), .dinb(n5862), .dout(n17876));
  jand g17618(.dina(n17876), .dinb(n17875), .dout(n17877));
  jand g17619(.dina(n17877), .dinb(n17874), .dout(n17878));
  jand g17620(.dina(n17878), .dinb(n17873), .dout(n17879));
  jxor g17621(.dina(n17879), .dinb(a47 ), .dout(n17880));
  jnot g17622(.din(n17880), .dout(n17881));
  jand g17623(.dina(n17781), .dinb(n17717), .dout(n17882));
  jand g17624(.dina(n17782), .dinb(n17712), .dout(n17883));
  jor  g17625(.dina(n17883), .dinb(n17882), .dout(n17884));
  jand g17626(.dina(n17761), .dinb(n17757), .dout(n17885));
  jand g17627(.dina(n17762), .dinb(n17726), .dout(n17886));
  jor  g17628(.dina(n17886), .dinb(n17885), .dout(n17887));
  jor  g17629(.dina(n9891), .dinb(n3227), .dout(n17888));
  jor  g17630(.dina(n9593), .dinb(n3035), .dout(n17889));
  jor  g17631(.dina(n9894), .dinb(n3055), .dout(n17890));
  jor  g17632(.dina(n9896), .dinb(n3230), .dout(n17891));
  jand g17633(.dina(n17891), .dinb(n17890), .dout(n17892));
  jand g17634(.dina(n17892), .dinb(n17889), .dout(n17893));
  jand g17635(.dina(n17893), .dinb(n17888), .dout(n17894));
  jxor g17636(.dina(n17894), .dinb(a59 ), .dout(n17895));
  jnot g17637(.din(n17895), .dout(n17896));
  jand g17638(.dina(n17755), .dinb(n17740), .dout(n17897));
  jand g17639(.dina(n17756), .dinb(n17735), .dout(n17898));
  jor  g17640(.dina(n17898), .dinb(n17897), .dout(n17899));
  jxor g17641(.dina(n17899), .dinb(n17896), .dout(n17900));
  jand g17642(.dina(n17744), .dinb(n17510), .dout(n17901));
  jnot g17643(.din(n17901), .dout(n17902));
  jor  g17644(.dina(n17754), .dinb(n17746), .dout(n17903));
  jand g17645(.dina(n17903), .dinb(n17902), .dout(n17904));
  jnot g17646(.din(n17904), .dout(n17905));
  jand g17647(.dina(n10801), .dinb(b27 ), .dout(n17906));
  jand g17648(.dina(n11107), .dinb(b26 ), .dout(n17907));
  jor  g17649(.dina(n17907), .dinb(n17906), .dout(n17908));
  jxor g17650(.dina(n17908), .dinb(n17841), .dout(n17909));
  jxor g17651(.dina(n17909), .dinb(n17743), .dout(n17910));
  jxor g17652(.dina(n17910), .dinb(n17905), .dout(n17911));
  jor  g17653(.dina(n10806), .dinb(n2867), .dout(n17912));
  jor  g17654(.dina(n10485), .dinb(n2559), .dout(n17913));
  jor  g17655(.dina(n10809), .dinb(n2579), .dout(n17914));
  jor  g17656(.dina(n10811), .dinb(n2870), .dout(n17915));
  jand g17657(.dina(n17915), .dinb(n17914), .dout(n17916));
  jand g17658(.dina(n17916), .dinb(n17913), .dout(n17917));
  jand g17659(.dina(n17917), .dinb(n17912), .dout(n17918));
  jxor g17660(.dina(n17918), .dinb(a62 ), .dout(n17919));
  jnot g17661(.din(n17919), .dout(n17920));
  jxor g17662(.dina(n17920), .dinb(n17911), .dout(n17921));
  jxor g17663(.dina(n17921), .dinb(n17900), .dout(n17922));
  jnot g17664(.din(n17922), .dout(n17923));
  jor  g17665(.dina(n8978), .dinb(n3939), .dout(n17924));
  jor  g17666(.dina(n8677), .dinb(n3403), .dout(n17925));
  jor  g17667(.dina(n8981), .dinb(n3588), .dout(n17926));
  jor  g17668(.dina(n8983), .dinb(n3942), .dout(n17927));
  jand g17669(.dina(n17927), .dinb(n17926), .dout(n17928));
  jand g17670(.dina(n17928), .dinb(n17925), .dout(n17929));
  jand g17671(.dina(n17929), .dinb(n17924), .dout(n17930));
  jxor g17672(.dina(n17930), .dinb(a56 ), .dout(n17931));
  jxor g17673(.dina(n17931), .dinb(n17923), .dout(n17932));
  jxor g17674(.dina(n17932), .dinb(n17887), .dout(n17933));
  jnot g17675(.din(n17933), .dout(n17934));
  jor  g17676(.dina(n8125), .dinb(n4534), .dout(n17935));
  jor  g17677(.dina(n7846), .dinb(n4140), .dout(n17936));
  jor  g17678(.dina(n8128), .dinb(n4340), .dout(n17937));
  jor  g17679(.dina(n8130), .dinb(n4537), .dout(n17938));
  jand g17680(.dina(n17938), .dinb(n17937), .dout(n17939));
  jand g17681(.dina(n17939), .dinb(n17936), .dout(n17940));
  jand g17682(.dina(n17940), .dinb(n17935), .dout(n17941));
  jxor g17683(.dina(n17941), .dinb(a53 ), .dout(n17942));
  jxor g17684(.dina(n17942), .dinb(n17934), .dout(n17943));
  jor  g17685(.dina(n17770), .dinb(n17763), .dout(n17944));
  jand g17686(.dina(n17770), .dinb(n17763), .dout(n17945));
  jor  g17687(.dina(n17780), .dinb(n17945), .dout(n17946));
  jand g17688(.dina(n17946), .dinb(n17944), .dout(n17947));
  jxor g17689(.dina(n17947), .dinb(n17943), .dout(n17948));
  jnot g17690(.din(n17948), .dout(n17949));
  jor  g17691(.dina(n7266), .dinb(n4991), .dout(n17950));
  jor  g17692(.dina(n7021), .dinb(n4557), .dout(n17951));
  jor  g17693(.dina(n7269), .dinb(n4974), .dout(n17952));
  jor  g17694(.dina(n7271), .dinb(n4994), .dout(n17953));
  jand g17695(.dina(n17953), .dinb(n17952), .dout(n17954));
  jand g17696(.dina(n17954), .dinb(n17951), .dout(n17955));
  jand g17697(.dina(n17955), .dinb(n17950), .dout(n17956));
  jxor g17698(.dina(n17956), .dinb(a50 ), .dout(n17957));
  jxor g17699(.dina(n17957), .dinb(n17949), .dout(n17958));
  jxor g17700(.dina(n17958), .dinb(n17884), .dout(n17959));
  jxor g17701(.dina(n17959), .dinb(n17881), .dout(n17960));
  jxor g17702(.dina(n17960), .dinb(n17872), .dout(n17961));
  jnot g17703(.din(n17961), .dout(n17962));
  jor  g17704(.dina(n6369), .dinb(n5739), .dout(n17963));
  jor  g17705(.dina(n5574), .dinb(n6106), .dout(n17964));
  jor  g17706(.dina(n5742), .dinb(n6352), .dout(n17965));
  jor  g17707(.dina(n5744), .dinb(n6372), .dout(n17966));
  jand g17708(.dina(n17966), .dinb(n17965), .dout(n17967));
  jand g17709(.dina(n17967), .dinb(n17964), .dout(n17968));
  jand g17710(.dina(n17968), .dinb(n17963), .dout(n17969));
  jxor g17711(.dina(n17969), .dinb(a44 ), .dout(n17970));
  jxor g17712(.dina(n17970), .dinb(n17962), .dout(n17971));
  jor  g17713(.dina(n17789), .dinb(n17785), .dout(n17972));
  jand g17714(.dina(n17789), .dinb(n17785), .dout(n17973));
  jor  g17715(.dina(n17799), .dinb(n17973), .dout(n17974));
  jand g17716(.dina(n17974), .dinb(n17972), .dout(n17975));
  jxor g17717(.dina(n17975), .dinb(n17971), .dout(n17976));
  jnot g17718(.din(n17976), .dout(n17977));
  jor  g17719(.dina(n7146), .dinb(n5096), .dout(n17978));
  jor  g17720(.dina(n4904), .dinb(n6867), .dout(n17979));
  jor  g17721(.dina(n5099), .dinb(n7129), .dout(n17980));
  jor  g17722(.dina(n5101), .dinb(n7149), .dout(n17981));
  jand g17723(.dina(n17981), .dinb(n17980), .dout(n17982));
  jand g17724(.dina(n17982), .dinb(n17979), .dout(n17983));
  jand g17725(.dina(n17983), .dinb(n17978), .dout(n17984));
  jxor g17726(.dina(n17984), .dinb(a41 ), .dout(n17985));
  jxor g17727(.dina(n17985), .dinb(n17977), .dout(n17986));
  jxor g17728(.dina(n17986), .dinb(n17869), .dout(n17987));
  jxor g17729(.dina(n17987), .dinb(n17865), .dout(n17988));
  jxor g17730(.dina(n17988), .dinb(n17857), .dout(n17989));
  jnot g17731(.din(n17989), .dout(n17990));
  jor  g17732(.dina(n8806), .dinb(n3849), .dout(n17991));
  jor  g17733(.dina(n3689), .dinb(n8231), .dout(n17992));
  jor  g17734(.dina(n3852), .dinb(n8789), .dout(n17993));
  jor  g17735(.dina(n3854), .dinb(n8809), .dout(n17994));
  jand g17736(.dina(n17994), .dinb(n17993), .dout(n17995));
  jand g17737(.dina(n17995), .dinb(n17992), .dout(n17996));
  jand g17738(.dina(n17996), .dinb(n17991), .dout(n17997));
  jxor g17739(.dina(n17997), .dinb(a35 ), .dout(n17998));
  jxor g17740(.dina(n17998), .dinb(n17990), .dout(n17999));
  jor  g17741(.dina(n17832), .dinb(n17826), .dout(n18000));
  jand g17742(.dina(n17832), .dinb(n17826), .dout(n18001));
  jor  g17743(.dina(n18001), .dinb(n17682), .dout(n18002));
  jand g17744(.dina(n18002), .dinb(n18000), .dout(n18003));
  jxor g17745(.dina(n18003), .dinb(n17999), .dout(n18004));
  jor  g17746(.dina(n9722), .dinb(n3301), .dout(n18005));
  jor  g17747(.dina(n3136), .dinb(n9390), .dout(n18006));
  jor  g17748(.dina(n3304), .dinb(n9413), .dout(n18007));
  jor  g17749(.dina(n3306), .dinb(n9725), .dout(n18008));
  jand g17750(.dina(n18008), .dinb(n18007), .dout(n18009));
  jand g17751(.dina(n18009), .dinb(n18006), .dout(n18010));
  jand g17752(.dina(n18010), .dinb(n18005), .dout(n18011));
  jxor g17753(.dina(n18011), .dinb(a32 ), .dout(n18012));
  jnot g17754(.din(n18012), .dout(n18013));
  jand g17755(.dina(n17672), .dinb(n17668), .dout(n18014));
  jnot g17756(.din(n18014), .dout(n18015));
  jnot g17757(.din(n17668), .dout(n18016));
  jand g17758(.dina(n17671), .dinb(n18016), .dout(n18017));
  jor  g17759(.dina(n17834), .dinb(n18017), .dout(n18018));
  jand g17760(.dina(n18018), .dinb(n18015), .dout(n18019));
  jxor g17761(.dina(n18019), .dinb(n18013), .dout(n18020));
  jxor g17762(.dina(n18020), .dinb(n18004), .dout(n18021));
  jor  g17763(.dina(n17659), .dinb(n17655), .dout(n18022));
  jand g17764(.dina(n17835), .dinb(n17660), .dout(n18023));
  jnot g17765(.din(n18023), .dout(n18024));
  jand g17766(.dina(n18024), .dinb(n18022), .dout(n18025));
  jor  g17767(.dina(n10961), .dinb(n2784), .dout(n18026));
  jor  g17768(.dina(n2661), .dinb(n10314), .dout(n18027));
  jor  g17769(.dina(n2787), .dinb(n10637), .dout(n18028));
  jor  g17770(.dina(n2789), .dinb(n10964), .dout(n18029));
  jand g17771(.dina(n18029), .dinb(n18028), .dout(n18030));
  jand g17772(.dina(n18030), .dinb(n18027), .dout(n18031));
  jand g17773(.dina(n18031), .dinb(n18026), .dout(n18032));
  jxor g17774(.dina(n18032), .dinb(a29 ), .dout(n18033));
  jxor g17775(.dina(n18033), .dinb(n18025), .dout(n18034));
  jxor g17776(.dina(n18034), .dinb(n18021), .dout(n18035));
  jxor g17777(.dina(n18035), .dinb(n17854), .dout(n18036));
  jand g17778(.dina(n17847), .dinb(n17647), .dout(n18037));
  jand g17779(.dina(n17848), .dinb(n17642), .dout(n18038));
  jor  g17780(.dina(n18038), .dinb(n18037), .dout(n18039));
  jxor g17781(.dina(n18039), .dinb(n18036), .dout(f90 ));
  jor  g17782(.dina(n18033), .dinb(n18025), .dout(n18041));
  jand g17783(.dina(n18034), .dinb(n18021), .dout(n18042));
  jnot g17784(.din(n18042), .dout(n18043));
  jand g17785(.dina(n18043), .dinb(n18041), .dout(n18044));
  jnot g17786(.din(n18044), .dout(n18045));
  jand g17787(.dina(n18019), .dinb(n18013), .dout(n18046));
  jand g17788(.dina(n18020), .dinb(n18004), .dout(n18047));
  jor  g17789(.dina(n18047), .dinb(n18046), .dout(n18048));
  jnot g17790(.din(n18048), .dout(n18049));
  jor  g17791(.dina(n10978), .dinb(n2784), .dout(n18050));
  jor  g17792(.dina(n2661), .dinb(n10637), .dout(n18051));
  jor  g17793(.dina(n2787), .dinb(n10964), .dout(n18052));
  jand g17794(.dina(n18052), .dinb(n18051), .dout(n18053));
  jand g17795(.dina(n18053), .dinb(n18050), .dout(n18054));
  jxor g17796(.dina(n18054), .dinb(a29 ), .dout(n18055));
  jxor g17797(.dina(n18055), .dinb(n18049), .dout(n18056));
  jor  g17798(.dina(n10311), .dinb(n3301), .dout(n18057));
  jor  g17799(.dina(n3136), .dinb(n9413), .dout(n18058));
  jor  g17800(.dina(n3304), .dinb(n9725), .dout(n18059));
  jor  g17801(.dina(n3306), .dinb(n10314), .dout(n18060));
  jand g17802(.dina(n18060), .dinb(n18059), .dout(n18061));
  jand g17803(.dina(n18061), .dinb(n18058), .dout(n18062));
  jand g17804(.dina(n18062), .dinb(n18057), .dout(n18063));
  jxor g17805(.dina(n18063), .dinb(a32 ), .dout(n18064));
  jor  g17806(.dina(n17998), .dinb(n17990), .dout(n18065));
  jand g17807(.dina(n18003), .dinb(n17999), .dout(n18066));
  jnot g17808(.din(n18066), .dout(n18067));
  jand g17809(.dina(n18067), .dinb(n18065), .dout(n18068));
  jxor g17810(.dina(n18068), .dinb(n18064), .dout(n18069));
  jor  g17811(.dina(n17987), .dinb(n17865), .dout(n18070));
  jand g17812(.dina(n17988), .dinb(n17857), .dout(n18071));
  jnot g17813(.din(n18071), .dout(n18072));
  jand g17814(.dina(n18072), .dinb(n18070), .dout(n18073));
  jnot g17815(.din(n18073), .dout(n18074));
  jor  g17816(.dina(n8228), .dinb(n4415), .dout(n18075));
  jor  g17817(.dina(n4272), .dinb(n7683), .dout(n18076));
  jor  g17818(.dina(n4418), .dinb(n7960), .dout(n18077));
  jor  g17819(.dina(n4420), .dinb(n8231), .dout(n18078));
  jand g17820(.dina(n18078), .dinb(n18077), .dout(n18079));
  jand g17821(.dina(n18079), .dinb(n18076), .dout(n18080));
  jand g17822(.dina(n18080), .dinb(n18075), .dout(n18081));
  jxor g17823(.dina(n18081), .dinb(a38 ), .dout(n18082));
  jnot g17824(.din(n18082), .dout(n18083));
  jor  g17825(.dina(n17970), .dinb(n17962), .dout(n18084));
  jand g17826(.dina(n17975), .dinb(n17971), .dout(n18085));
  jnot g17827(.din(n18085), .dout(n18086));
  jand g17828(.dina(n18086), .dinb(n18084), .dout(n18087));
  jnot g17829(.din(n18087), .dout(n18088));
  jand g17830(.dina(n17959), .dinb(n17881), .dout(n18089));
  jand g17831(.dina(n17960), .dinb(n17872), .dout(n18090));
  jor  g17832(.dina(n18090), .dinb(n18089), .dout(n18091));
  jor  g17833(.dina(n17957), .dinb(n17949), .dout(n18092));
  jand g17834(.dina(n17958), .dinb(n17884), .dout(n18093));
  jnot g17835(.din(n18093), .dout(n18094));
  jand g17836(.dina(n18094), .dinb(n18092), .dout(n18095));
  jnot g17837(.din(n18095), .dout(n18096));
  jor  g17838(.dina(n17942), .dinb(n17934), .dout(n18097));
  jand g17839(.dina(n17947), .dinb(n17943), .dout(n18098));
  jnot g17840(.din(n18098), .dout(n18099));
  jand g17841(.dina(n18099), .dinb(n18097), .dout(n18100));
  jnot g17842(.din(n18100), .dout(n18101));
  jor  g17843(.dina(n8125), .dinb(n4554), .dout(n18102));
  jor  g17844(.dina(n7846), .dinb(n4340), .dout(n18103));
  jor  g17845(.dina(n8128), .dinb(n4537), .dout(n18104));
  jor  g17846(.dina(n8130), .dinb(n4557), .dout(n18105));
  jand g17847(.dina(n18105), .dinb(n18104), .dout(n18106));
  jand g17848(.dina(n18106), .dinb(n18103), .dout(n18107));
  jand g17849(.dina(n18107), .dinb(n18102), .dout(n18108));
  jxor g17850(.dina(n18108), .dinb(a53 ), .dout(n18109));
  jnot g17851(.din(n18109), .dout(n18110));
  jor  g17852(.dina(n17931), .dinb(n17923), .dout(n18111));
  jand g17853(.dina(n17932), .dinb(n17887), .dout(n18112));
  jnot g17854(.din(n18112), .dout(n18113));
  jand g17855(.dina(n18113), .dinb(n18111), .dout(n18114));
  jnot g17856(.din(n18114), .dout(n18115));
  jor  g17857(.dina(n8978), .dinb(n4137), .dout(n18116));
  jor  g17858(.dina(n8677), .dinb(n3588), .dout(n18117));
  jor  g17859(.dina(n8981), .dinb(n3942), .dout(n18118));
  jor  g17860(.dina(n8983), .dinb(n4140), .dout(n18119));
  jand g17861(.dina(n18119), .dinb(n18118), .dout(n18120));
  jand g17862(.dina(n18120), .dinb(n18117), .dout(n18121));
  jand g17863(.dina(n18121), .dinb(n18116), .dout(n18122));
  jxor g17864(.dina(n18122), .dinb(a56 ), .dout(n18123));
  jnot g17865(.din(n18123), .dout(n18124));
  jand g17866(.dina(n17899), .dinb(n17896), .dout(n18125));
  jand g17867(.dina(n17921), .dinb(n17900), .dout(n18126));
  jor  g17868(.dina(n18126), .dinb(n18125), .dout(n18127));
  jand g17869(.dina(n17908), .dinb(n17841), .dout(n18128));
  jand g17870(.dina(n17909), .dinb(n17743), .dout(n18129));
  jor  g17871(.dina(n18129), .dinb(n18128), .dout(n18130));
  jand g17872(.dina(n10801), .dinb(b28 ), .dout(n18131));
  jand g17873(.dina(n11107), .dinb(b27 ), .dout(n18132));
  jor  g17874(.dina(n18132), .dinb(n18131), .dout(n18133));
  jnot g17875(.din(n18133), .dout(n18134));
  jxor g17876(.dina(n18134), .dinb(n18130), .dout(n18135));
  jnot g17877(.din(n18135), .dout(n18136));
  jor  g17878(.dina(n10806), .dinb(n3032), .dout(n18137));
  jor  g17879(.dina(n10485), .dinb(n2579), .dout(n18138));
  jor  g17880(.dina(n10809), .dinb(n2870), .dout(n18139));
  jor  g17881(.dina(n10811), .dinb(n3035), .dout(n18140));
  jand g17882(.dina(n18140), .dinb(n18139), .dout(n18141));
  jand g17883(.dina(n18141), .dinb(n18138), .dout(n18142));
  jand g17884(.dina(n18142), .dinb(n18137), .dout(n18143));
  jxor g17885(.dina(n18143), .dinb(a62 ), .dout(n18144));
  jxor g17886(.dina(n18144), .dinb(n18136), .dout(n18145));
  jor  g17887(.dina(n17910), .dinb(n17905), .dout(n18146));
  jand g17888(.dina(n17910), .dinb(n17905), .dout(n18147));
  jor  g17889(.dina(n17920), .dinb(n18147), .dout(n18148));
  jand g17890(.dina(n18148), .dinb(n18146), .dout(n18149));
  jxor g17891(.dina(n18149), .dinb(n18145), .dout(n18150));
  jor  g17892(.dina(n9891), .dinb(n3400), .dout(n18151));
  jor  g17893(.dina(n9593), .dinb(n3055), .dout(n18152));
  jor  g17894(.dina(n9894), .dinb(n3230), .dout(n18153));
  jor  g17895(.dina(n9896), .dinb(n3403), .dout(n18154));
  jand g17896(.dina(n18154), .dinb(n18153), .dout(n18155));
  jand g17897(.dina(n18155), .dinb(n18152), .dout(n18156));
  jand g17898(.dina(n18156), .dinb(n18151), .dout(n18157));
  jxor g17899(.dina(n18157), .dinb(a59 ), .dout(n18158));
  jnot g17900(.din(n18158), .dout(n18159));
  jxor g17901(.dina(n18159), .dinb(n18150), .dout(n18160));
  jxor g17902(.dina(n18160), .dinb(n18127), .dout(n18161));
  jxor g17903(.dina(n18161), .dinb(n18124), .dout(n18162));
  jxor g17904(.dina(n18162), .dinb(n18115), .dout(n18163));
  jxor g17905(.dina(n18163), .dinb(n18110), .dout(n18164));
  jxor g17906(.dina(n18164), .dinb(n18101), .dout(n18165));
  jor  g17907(.dina(n7266), .dinb(n5405), .dout(n18166));
  jor  g17908(.dina(n7021), .dinb(n4974), .dout(n18167));
  jor  g17909(.dina(n7269), .dinb(n4994), .dout(n18168));
  jor  g17910(.dina(n7271), .dinb(n5408), .dout(n18169));
  jand g17911(.dina(n18169), .dinb(n18168), .dout(n18170));
  jand g17912(.dina(n18170), .dinb(n18167), .dout(n18171));
  jand g17913(.dina(n18171), .dinb(n18166), .dout(n18172));
  jxor g17914(.dina(n18172), .dinb(a50 ), .dout(n18173));
  jnot g17915(.din(n18173), .dout(n18174));
  jxor g17916(.dina(n18174), .dinb(n18165), .dout(n18175));
  jxor g17917(.dina(n18175), .dinb(n18096), .dout(n18176));
  jor  g17918(.dina(n6103), .dinb(n6490), .dout(n18177));
  jor  g17919(.dina(n6262), .dinb(n5428), .dout(n18178));
  jor  g17920(.dina(n6493), .dinb(n5862), .dout(n18179));
  jor  g17921(.dina(n6495), .dinb(n6106), .dout(n18180));
  jand g17922(.dina(n18180), .dinb(n18179), .dout(n18181));
  jand g17923(.dina(n18181), .dinb(n18178), .dout(n18182));
  jand g17924(.dina(n18182), .dinb(n18177), .dout(n18183));
  jxor g17925(.dina(n18183), .dinb(a47 ), .dout(n18184));
  jnot g17926(.din(n18184), .dout(n18185));
  jxor g17927(.dina(n18185), .dinb(n18176), .dout(n18186));
  jxor g17928(.dina(n18186), .dinb(n18091), .dout(n18187));
  jor  g17929(.dina(n6864), .dinb(n5739), .dout(n18188));
  jor  g17930(.dina(n5574), .dinb(n6352), .dout(n18189));
  jor  g17931(.dina(n5742), .dinb(n6372), .dout(n18190));
  jor  g17932(.dina(n5744), .dinb(n6867), .dout(n18191));
  jand g17933(.dina(n18191), .dinb(n18190), .dout(n18192));
  jand g17934(.dina(n18192), .dinb(n18189), .dout(n18193));
  jand g17935(.dina(n18193), .dinb(n18188), .dout(n18194));
  jxor g17936(.dina(n18194), .dinb(a44 ), .dout(n18195));
  jnot g17937(.din(n18195), .dout(n18196));
  jxor g17938(.dina(n18196), .dinb(n18187), .dout(n18197));
  jxor g17939(.dina(n18197), .dinb(n18088), .dout(n18198));
  jor  g17940(.dina(n7408), .dinb(n5096), .dout(n18199));
  jor  g17941(.dina(n4904), .dinb(n7129), .dout(n18200));
  jor  g17942(.dina(n5099), .dinb(n7149), .dout(n18201));
  jor  g17943(.dina(n5101), .dinb(n7411), .dout(n18202));
  jand g17944(.dina(n18202), .dinb(n18201), .dout(n18203));
  jand g17945(.dina(n18203), .dinb(n18200), .dout(n18204));
  jand g17946(.dina(n18204), .dinb(n18199), .dout(n18205));
  jxor g17947(.dina(n18205), .dinb(a41 ), .dout(n18206));
  jnot g17948(.din(n18206), .dout(n18207));
  jxor g17949(.dina(n18207), .dinb(n18198), .dout(n18208));
  jand g17950(.dina(n17985), .dinb(n17977), .dout(n18209));
  jnot g17951(.din(n17985), .dout(n18210));
  jand g17952(.dina(n18210), .dinb(n17976), .dout(n18211));
  jnot g17953(.din(n18211), .dout(n18212));
  jand g17954(.dina(n18212), .dinb(n17869), .dout(n18213));
  jor  g17955(.dina(n18213), .dinb(n18209), .dout(n18214));
  jnot g17956(.din(n18214), .dout(n18215));
  jxor g17957(.dina(n18215), .dinb(n18208), .dout(n18216));
  jxor g17958(.dina(n18216), .dinb(n18083), .dout(n18217));
  jxor g17959(.dina(n18217), .dinb(n18074), .dout(n18218));
  jor  g17960(.dina(n9387), .dinb(n3849), .dout(n18219));
  jor  g17961(.dina(n3689), .dinb(n8789), .dout(n18220));
  jor  g17962(.dina(n3852), .dinb(n8809), .dout(n18221));
  jor  g17963(.dina(n3854), .dinb(n9390), .dout(n18222));
  jand g17964(.dina(n18222), .dinb(n18221), .dout(n18223));
  jand g17965(.dina(n18223), .dinb(n18220), .dout(n18224));
  jand g17966(.dina(n18224), .dinb(n18219), .dout(n18225));
  jxor g17967(.dina(n18225), .dinb(a35 ), .dout(n18226));
  jnot g17968(.din(n18226), .dout(n18227));
  jxor g17969(.dina(n18227), .dinb(n18218), .dout(n18228));
  jxor g17970(.dina(n18228), .dinb(n18069), .dout(n18229));
  jxor g17971(.dina(n18229), .dinb(n18056), .dout(n18230));
  jxor g17972(.dina(n18230), .dinb(n18045), .dout(n18231));
  jand g17973(.dina(n18035), .dinb(n17854), .dout(n18232));
  jand g17974(.dina(n18039), .dinb(n18036), .dout(n18233));
  jor  g17975(.dina(n18233), .dinb(n18232), .dout(n18234));
  jxor g17976(.dina(n18234), .dinb(n18231), .dout(f91 ));
  jand g17977(.dina(n18230), .dinb(n18045), .dout(n18236));
  jand g17978(.dina(n18234), .dinb(n18231), .dout(n18237));
  jor  g17979(.dina(n18237), .dinb(n18236), .dout(n18238));
  jor  g17980(.dina(n18055), .dinb(n18049), .dout(n18239));
  jand g17981(.dina(n18229), .dinb(n18056), .dout(n18240));
  jnot g17982(.din(n18240), .dout(n18241));
  jand g17983(.dina(n18241), .dinb(n18239), .dout(n18242));
  jnot g17984(.din(n18242), .dout(n18243));
  jor  g17985(.dina(n10634), .dinb(n3301), .dout(n18244));
  jor  g17986(.dina(n3136), .dinb(n9725), .dout(n18245));
  jor  g17987(.dina(n3304), .dinb(n10314), .dout(n18246));
  jor  g17988(.dina(n3306), .dinb(n10637), .dout(n18247));
  jand g17989(.dina(n18247), .dinb(n18246), .dout(n18248));
  jand g17990(.dina(n18248), .dinb(n18245), .dout(n18249));
  jand g17991(.dina(n18249), .dinb(n18244), .dout(n18250));
  jxor g17992(.dina(n18250), .dinb(a32 ), .dout(n18251));
  jnot g17993(.din(n18251), .dout(n18252));
  jor  g17994(.dina(n18217), .dinb(n18074), .dout(n18253));
  jand g17995(.dina(n18217), .dinb(n18074), .dout(n18254));
  jor  g17996(.dina(n18227), .dinb(n18254), .dout(n18255));
  jand g17997(.dina(n18255), .dinb(n18253), .dout(n18256));
  jxor g17998(.dina(n18256), .dinb(n18252), .dout(n18257));
  jand g17999(.dina(n18215), .dinb(n18208), .dout(n18258));
  jand g18000(.dina(n18216), .dinb(n18083), .dout(n18259));
  jor  g18001(.dina(n18259), .dinb(n18258), .dout(n18260));
  jor  g18002(.dina(n8786), .dinb(n4415), .dout(n18261));
  jor  g18003(.dina(n4272), .dinb(n7960), .dout(n18262));
  jor  g18004(.dina(n4418), .dinb(n8231), .dout(n18263));
  jor  g18005(.dina(n4420), .dinb(n8789), .dout(n18264));
  jand g18006(.dina(n18264), .dinb(n18263), .dout(n18265));
  jand g18007(.dina(n18265), .dinb(n18262), .dout(n18266));
  jand g18008(.dina(n18266), .dinb(n18261), .dout(n18267));
  jxor g18009(.dina(n18267), .dinb(a38 ), .dout(n18268));
  jnot g18010(.din(n18268), .dout(n18269));
  jor  g18011(.dina(n7680), .dinb(n5096), .dout(n18270));
  jor  g18012(.dina(n4904), .dinb(n7149), .dout(n18271));
  jor  g18013(.dina(n5099), .dinb(n7411), .dout(n18272));
  jor  g18014(.dina(n5101), .dinb(n7683), .dout(n18273));
  jand g18015(.dina(n18273), .dinb(n18272), .dout(n18274));
  jand g18016(.dina(n18274), .dinb(n18271), .dout(n18275));
  jand g18017(.dina(n18275), .dinb(n18270), .dout(n18276));
  jxor g18018(.dina(n18276), .dinb(a41 ), .dout(n18277));
  jnot g18019(.din(n18277), .dout(n18278));
  jor  g18020(.dina(n7266), .dinb(n5425), .dout(n18279));
  jor  g18021(.dina(n7021), .dinb(n4994), .dout(n18280));
  jor  g18022(.dina(n7269), .dinb(n5408), .dout(n18281));
  jor  g18023(.dina(n7271), .dinb(n5428), .dout(n18282));
  jand g18024(.dina(n18282), .dinb(n18281), .dout(n18283));
  jand g18025(.dina(n18283), .dinb(n18280), .dout(n18284));
  jand g18026(.dina(n18284), .dinb(n18279), .dout(n18285));
  jxor g18027(.dina(n18285), .dinb(a50 ), .dout(n18286));
  jnot g18028(.din(n18286), .dout(n18287));
  jand g18029(.dina(n18162), .dinb(n18115), .dout(n18288));
  jand g18030(.dina(n18163), .dinb(n18110), .dout(n18289));
  jor  g18031(.dina(n18289), .dinb(n18288), .dout(n18290));
  jor  g18032(.dina(n8125), .dinb(n4971), .dout(n18291));
  jor  g18033(.dina(n7846), .dinb(n4537), .dout(n18292));
  jor  g18034(.dina(n8128), .dinb(n4557), .dout(n18293));
  jor  g18035(.dina(n8130), .dinb(n4974), .dout(n18294));
  jand g18036(.dina(n18294), .dinb(n18293), .dout(n18295));
  jand g18037(.dina(n18295), .dinb(n18292), .dout(n18296));
  jand g18038(.dina(n18296), .dinb(n18291), .dout(n18297));
  jxor g18039(.dina(n18297), .dinb(a53 ), .dout(n18298));
  jnot g18040(.din(n18298), .dout(n18299));
  jand g18041(.dina(n18160), .dinb(n18127), .dout(n18300));
  jand g18042(.dina(n18161), .dinb(n18124), .dout(n18301));
  jor  g18043(.dina(n18301), .dinb(n18300), .dout(n18302));
  jor  g18044(.dina(n9891), .dinb(n3585), .dout(n18303));
  jor  g18045(.dina(n9593), .dinb(n3230), .dout(n18304));
  jor  g18046(.dina(n9894), .dinb(n3403), .dout(n18305));
  jor  g18047(.dina(n9896), .dinb(n3588), .dout(n18306));
  jand g18048(.dina(n18306), .dinb(n18305), .dout(n18307));
  jand g18049(.dina(n18307), .dinb(n18304), .dout(n18308));
  jand g18050(.dina(n18308), .dinb(n18303), .dout(n18309));
  jxor g18051(.dina(n18309), .dinb(a59 ), .dout(n18310));
  jnot g18052(.din(n18310), .dout(n18311));
  jor  g18053(.dina(n10806), .dinb(n3052), .dout(n18312));
  jor  g18054(.dina(n10485), .dinb(n2870), .dout(n18313));
  jor  g18055(.dina(n10809), .dinb(n3035), .dout(n18314));
  jor  g18056(.dina(n10811), .dinb(n3055), .dout(n18315));
  jand g18057(.dina(n18315), .dinb(n18314), .dout(n18316));
  jand g18058(.dina(n18316), .dinb(n18313), .dout(n18317));
  jand g18059(.dina(n18317), .dinb(n18312), .dout(n18318));
  jxor g18060(.dina(n18318), .dinb(a62 ), .dout(n18319));
  jnot g18061(.din(n18319), .dout(n18320));
  jand g18062(.dina(n18134), .dinb(n18130), .dout(n18321));
  jnot g18063(.din(n18321), .dout(n18322));
  jor  g18064(.dina(n18144), .dinb(n18136), .dout(n18323));
  jand g18065(.dina(n18323), .dinb(n18322), .dout(n18324));
  jnot g18066(.din(n18324), .dout(n18325));
  jand g18067(.dina(n10801), .dinb(b29 ), .dout(n18326));
  jand g18068(.dina(n11107), .dinb(b28 ), .dout(n18327));
  jor  g18069(.dina(n18327), .dinb(n18326), .dout(n18328));
  jnot g18070(.din(n18328), .dout(n18329));
  jxor g18071(.dina(n18329), .dinb(n18133), .dout(n18330));
  jxor g18072(.dina(n18330), .dinb(n18325), .dout(n18331));
  jxor g18073(.dina(n18331), .dinb(n18320), .dout(n18332));
  jxor g18074(.dina(n18332), .dinb(n18311), .dout(n18333));
  jor  g18075(.dina(n18149), .dinb(n18145), .dout(n18334));
  jand g18076(.dina(n18149), .dinb(n18145), .dout(n18335));
  jor  g18077(.dina(n18159), .dinb(n18335), .dout(n18336));
  jand g18078(.dina(n18336), .dinb(n18334), .dout(n18337));
  jxor g18079(.dina(n18337), .dinb(n18333), .dout(n18338));
  jor  g18080(.dina(n8978), .dinb(n4337), .dout(n18339));
  jor  g18081(.dina(n8677), .dinb(n3942), .dout(n18340));
  jor  g18082(.dina(n8981), .dinb(n4140), .dout(n18341));
  jor  g18083(.dina(n8983), .dinb(n4340), .dout(n18342));
  jand g18084(.dina(n18342), .dinb(n18341), .dout(n18343));
  jand g18085(.dina(n18343), .dinb(n18340), .dout(n18344));
  jand g18086(.dina(n18344), .dinb(n18339), .dout(n18345));
  jxor g18087(.dina(n18345), .dinb(a56 ), .dout(n18346));
  jnot g18088(.din(n18346), .dout(n18347));
  jxor g18089(.dina(n18347), .dinb(n18338), .dout(n18348));
  jxor g18090(.dina(n18348), .dinb(n18302), .dout(n18349));
  jxor g18091(.dina(n18349), .dinb(n18299), .dout(n18350));
  jxor g18092(.dina(n18350), .dinb(n18290), .dout(n18351));
  jxor g18093(.dina(n18351), .dinb(n18287), .dout(n18352));
  jor  g18094(.dina(n18164), .dinb(n18101), .dout(n18353));
  jand g18095(.dina(n18164), .dinb(n18101), .dout(n18354));
  jor  g18096(.dina(n18174), .dinb(n18354), .dout(n18355));
  jand g18097(.dina(n18355), .dinb(n18353), .dout(n18356));
  jxor g18098(.dina(n18356), .dinb(n18352), .dout(n18357));
  jor  g18099(.dina(n6349), .dinb(n6490), .dout(n18358));
  jor  g18100(.dina(n6262), .dinb(n5862), .dout(n18359));
  jor  g18101(.dina(n6493), .dinb(n6106), .dout(n18360));
  jor  g18102(.dina(n6495), .dinb(n6352), .dout(n18361));
  jand g18103(.dina(n18361), .dinb(n18360), .dout(n18362));
  jand g18104(.dina(n18362), .dinb(n18359), .dout(n18363));
  jand g18105(.dina(n18363), .dinb(n18358), .dout(n18364));
  jxor g18106(.dina(n18364), .dinb(a47 ), .dout(n18365));
  jnot g18107(.din(n18365), .dout(n18366));
  jxor g18108(.dina(n18366), .dinb(n18357), .dout(n18367));
  jnot g18109(.din(n18175), .dout(n18368));
  jand g18110(.dina(n18368), .dinb(n18095), .dout(n18369));
  jnot g18111(.din(n18369), .dout(n18370));
  jand g18112(.dina(n18175), .dinb(n18096), .dout(n18371));
  jor  g18113(.dina(n18185), .dinb(n18371), .dout(n18372));
  jand g18114(.dina(n18372), .dinb(n18370), .dout(n18373));
  jxor g18115(.dina(n18373), .dinb(n18367), .dout(n18374));
  jnot g18116(.din(n18374), .dout(n18375));
  jor  g18117(.dina(n7126), .dinb(n5739), .dout(n18376));
  jor  g18118(.dina(n5574), .dinb(n6372), .dout(n18377));
  jor  g18119(.dina(n5742), .dinb(n6867), .dout(n18378));
  jor  g18120(.dina(n5744), .dinb(n7129), .dout(n18379));
  jand g18121(.dina(n18379), .dinb(n18378), .dout(n18380));
  jand g18122(.dina(n18380), .dinb(n18377), .dout(n18381));
  jand g18123(.dina(n18381), .dinb(n18376), .dout(n18382));
  jxor g18124(.dina(n18382), .dinb(a44 ), .dout(n18383));
  jxor g18125(.dina(n18383), .dinb(n18375), .dout(n18384));
  jnot g18126(.din(n18091), .dout(n18385));
  jnot g18127(.din(n18186), .dout(n18386));
  jand g18128(.dina(n18386), .dinb(n18385), .dout(n18387));
  jnot g18129(.din(n18387), .dout(n18388));
  jand g18130(.dina(n18186), .dinb(n18091), .dout(n18389));
  jor  g18131(.dina(n18196), .dinb(n18389), .dout(n18390));
  jand g18132(.dina(n18390), .dinb(n18388), .dout(n18391));
  jxor g18133(.dina(n18391), .dinb(n18384), .dout(n18392));
  jxor g18134(.dina(n18392), .dinb(n18278), .dout(n18393));
  jnot g18135(.din(n18197), .dout(n18394));
  jand g18136(.dina(n18394), .dinb(n18087), .dout(n18395));
  jnot g18137(.din(n18395), .dout(n18396));
  jand g18138(.dina(n18197), .dinb(n18088), .dout(n18397));
  jor  g18139(.dina(n18207), .dinb(n18397), .dout(n18398));
  jand g18140(.dina(n18398), .dinb(n18396), .dout(n18399));
  jxor g18141(.dina(n18399), .dinb(n18393), .dout(n18400));
  jxor g18142(.dina(n18400), .dinb(n18269), .dout(n18401));
  jxor g18143(.dina(n18401), .dinb(n18260), .dout(n18402));
  jor  g18144(.dina(n9410), .dinb(n3849), .dout(n18403));
  jor  g18145(.dina(n3689), .dinb(n8809), .dout(n18404));
  jor  g18146(.dina(n3852), .dinb(n9390), .dout(n18405));
  jor  g18147(.dina(n3854), .dinb(n9413), .dout(n18406));
  jand g18148(.dina(n18406), .dinb(n18405), .dout(n18407));
  jand g18149(.dina(n18407), .dinb(n18404), .dout(n18408));
  jand g18150(.dina(n18408), .dinb(n18403), .dout(n18409));
  jxor g18151(.dina(n18409), .dinb(a35 ), .dout(n18410));
  jnot g18152(.din(n18410), .dout(n18411));
  jxor g18153(.dina(n18411), .dinb(n18402), .dout(n18412));
  jxor g18154(.dina(n18412), .dinb(n18257), .dout(n18413));
  jor  g18155(.dina(n18068), .dinb(n18064), .dout(n18414));
  jand g18156(.dina(n18228), .dinb(n18069), .dout(n18415));
  jnot g18157(.din(n18415), .dout(n18416));
  jand g18158(.dina(n18416), .dinb(n18414), .dout(n18417));
  jnot g18159(.din(a29 ), .dout(n18418));
  jand g18160(.dina(n11296), .dinb(n2482), .dout(n18419));
  jor  g18161(.dina(n18419), .dinb(n2662), .dout(n18420));
  jand g18162(.dina(n18420), .dinb(b63 ), .dout(n18421));
  jxor g18163(.dina(n18421), .dinb(n18418), .dout(n18422));
  jxor g18164(.dina(n18422), .dinb(n18417), .dout(n18423));
  jxor g18165(.dina(n18423), .dinb(n18413), .dout(n18424));
  jxor g18166(.dina(n18424), .dinb(n18243), .dout(n18425));
  jxor g18167(.dina(n18425), .dinb(n18238), .dout(f92 ));
  jand g18168(.dina(n18424), .dinb(n18243), .dout(n18427));
  jand g18169(.dina(n18425), .dinb(n18238), .dout(n18428));
  jor  g18170(.dina(n18428), .dinb(n18427), .dout(n18429));
  jor  g18171(.dina(n18422), .dinb(n18417), .dout(n18430));
  jand g18172(.dina(n18423), .dinb(n18413), .dout(n18431));
  jnot g18173(.din(n18431), .dout(n18432));
  jand g18174(.dina(n18432), .dinb(n18430), .dout(n18433));
  jnot g18175(.din(n18433), .dout(n18434));
  jand g18176(.dina(n18399), .dinb(n18393), .dout(n18435));
  jand g18177(.dina(n18400), .dinb(n18269), .dout(n18436));
  jor  g18178(.dina(n18436), .dinb(n18435), .dout(n18437));
  jand g18179(.dina(n18391), .dinb(n18384), .dout(n18438));
  jand g18180(.dina(n18392), .dinb(n18278), .dout(n18439));
  jor  g18181(.dina(n18439), .dinb(n18438), .dout(n18440));
  jor  g18182(.dina(n7957), .dinb(n5096), .dout(n18441));
  jor  g18183(.dina(n4904), .dinb(n7411), .dout(n18442));
  jor  g18184(.dina(n5099), .dinb(n7683), .dout(n18443));
  jor  g18185(.dina(n5101), .dinb(n7960), .dout(n18444));
  jand g18186(.dina(n18444), .dinb(n18443), .dout(n18445));
  jand g18187(.dina(n18445), .dinb(n18442), .dout(n18446));
  jand g18188(.dina(n18446), .dinb(n18441), .dout(n18447));
  jxor g18189(.dina(n18447), .dinb(a41 ), .dout(n18448));
  jand g18190(.dina(n18373), .dinb(n18367), .dout(n18449));
  jnot g18191(.din(n18449), .dout(n18450));
  jor  g18192(.dina(n18383), .dinb(n18375), .dout(n18451));
  jand g18193(.dina(n18451), .dinb(n18450), .dout(n18452));
  jand g18194(.dina(n18350), .dinb(n18290), .dout(n18453));
  jand g18195(.dina(n18351), .dinb(n18287), .dout(n18454));
  jor  g18196(.dina(n18454), .dinb(n18453), .dout(n18455));
  jor  g18197(.dina(n7266), .dinb(n5859), .dout(n18456));
  jor  g18198(.dina(n7021), .dinb(n5408), .dout(n18457));
  jor  g18199(.dina(n7269), .dinb(n5428), .dout(n18458));
  jor  g18200(.dina(n7271), .dinb(n5862), .dout(n18459));
  jand g18201(.dina(n18459), .dinb(n18458), .dout(n18460));
  jand g18202(.dina(n18460), .dinb(n18457), .dout(n18461));
  jand g18203(.dina(n18461), .dinb(n18456), .dout(n18462));
  jxor g18204(.dina(n18462), .dinb(a50 ), .dout(n18463));
  jnot g18205(.din(n18463), .dout(n18464));
  jand g18206(.dina(n18348), .dinb(n18302), .dout(n18465));
  jand g18207(.dina(n18349), .dinb(n18299), .dout(n18466));
  jor  g18208(.dina(n18466), .dinb(n18465), .dout(n18467));
  jand g18209(.dina(n18331), .dinb(n18320), .dout(n18468));
  jand g18210(.dina(n18332), .dinb(n18311), .dout(n18469));
  jor  g18211(.dina(n18469), .dinb(n18468), .dout(n18470));
  jor  g18212(.dina(n9891), .dinb(n3939), .dout(n18471));
  jor  g18213(.dina(n9593), .dinb(n3403), .dout(n18472));
  jor  g18214(.dina(n9894), .dinb(n3588), .dout(n18473));
  jor  g18215(.dina(n9896), .dinb(n3942), .dout(n18474));
  jand g18216(.dina(n18474), .dinb(n18473), .dout(n18475));
  jand g18217(.dina(n18475), .dinb(n18472), .dout(n18476));
  jand g18218(.dina(n18476), .dinb(n18471), .dout(n18477));
  jxor g18219(.dina(n18477), .dinb(a59 ), .dout(n18478));
  jnot g18220(.din(n18478), .dout(n18479));
  jor  g18221(.dina(n10806), .dinb(n3227), .dout(n18480));
  jor  g18222(.dina(n10485), .dinb(n3035), .dout(n18481));
  jor  g18223(.dina(n10809), .dinb(n3055), .dout(n18482));
  jor  g18224(.dina(n10811), .dinb(n3230), .dout(n18483));
  jand g18225(.dina(n18483), .dinb(n18482), .dout(n18484));
  jand g18226(.dina(n18484), .dinb(n18481), .dout(n18485));
  jand g18227(.dina(n18485), .dinb(n18480), .dout(n18486));
  jxor g18228(.dina(n18486), .dinb(a62 ), .dout(n18487));
  jnot g18229(.din(n18487), .dout(n18488));
  jand g18230(.dina(n18329), .dinb(n18133), .dout(n18489));
  jand g18231(.dina(n18330), .dinb(n18325), .dout(n18490));
  jor  g18232(.dina(n18490), .dinb(n18489), .dout(n18491));
  jand g18233(.dina(n10801), .dinb(b30 ), .dout(n18492));
  jand g18234(.dina(n11107), .dinb(b29 ), .dout(n18493));
  jor  g18235(.dina(n18493), .dinb(n18492), .dout(n18494));
  jxor g18236(.dina(n18494), .dinb(n18418), .dout(n18495));
  jxor g18237(.dina(n18495), .dinb(n18328), .dout(n18496));
  jxor g18238(.dina(n18496), .dinb(n18491), .dout(n18497));
  jxor g18239(.dina(n18497), .dinb(n18488), .dout(n18498));
  jxor g18240(.dina(n18498), .dinb(n18479), .dout(n18499));
  jxor g18241(.dina(n18499), .dinb(n18470), .dout(n18500));
  jnot g18242(.din(n18500), .dout(n18501));
  jor  g18243(.dina(n8978), .dinb(n4534), .dout(n18502));
  jor  g18244(.dina(n8677), .dinb(n4140), .dout(n18503));
  jor  g18245(.dina(n8981), .dinb(n4340), .dout(n18504));
  jor  g18246(.dina(n8983), .dinb(n4537), .dout(n18505));
  jand g18247(.dina(n18505), .dinb(n18504), .dout(n18506));
  jand g18248(.dina(n18506), .dinb(n18503), .dout(n18507));
  jand g18249(.dina(n18507), .dinb(n18502), .dout(n18508));
  jxor g18250(.dina(n18508), .dinb(a56 ), .dout(n18509));
  jxor g18251(.dina(n18509), .dinb(n18501), .dout(n18510));
  jor  g18252(.dina(n18337), .dinb(n18333), .dout(n18511));
  jand g18253(.dina(n18337), .dinb(n18333), .dout(n18512));
  jor  g18254(.dina(n18347), .dinb(n18512), .dout(n18513));
  jand g18255(.dina(n18513), .dinb(n18511), .dout(n18514));
  jxor g18256(.dina(n18514), .dinb(n18510), .dout(n18515));
  jnot g18257(.din(n18515), .dout(n18516));
  jor  g18258(.dina(n8125), .dinb(n4991), .dout(n18517));
  jor  g18259(.dina(n7846), .dinb(n4557), .dout(n18518));
  jor  g18260(.dina(n8128), .dinb(n4974), .dout(n18519));
  jor  g18261(.dina(n8130), .dinb(n4994), .dout(n18520));
  jand g18262(.dina(n18520), .dinb(n18519), .dout(n18521));
  jand g18263(.dina(n18521), .dinb(n18518), .dout(n18522));
  jand g18264(.dina(n18522), .dinb(n18517), .dout(n18523));
  jxor g18265(.dina(n18523), .dinb(a53 ), .dout(n18524));
  jxor g18266(.dina(n18524), .dinb(n18516), .dout(n18525));
  jxor g18267(.dina(n18525), .dinb(n18467), .dout(n18526));
  jxor g18268(.dina(n18526), .dinb(n18464), .dout(n18527));
  jxor g18269(.dina(n18527), .dinb(n18455), .dout(n18528));
  jnot g18270(.din(n18528), .dout(n18529));
  jor  g18271(.dina(n6369), .dinb(n6490), .dout(n18530));
  jor  g18272(.dina(n6262), .dinb(n6106), .dout(n18531));
  jor  g18273(.dina(n6493), .dinb(n6352), .dout(n18532));
  jor  g18274(.dina(n6495), .dinb(n6372), .dout(n18533));
  jand g18275(.dina(n18533), .dinb(n18532), .dout(n18534));
  jand g18276(.dina(n18534), .dinb(n18531), .dout(n18535));
  jand g18277(.dina(n18535), .dinb(n18530), .dout(n18536));
  jxor g18278(.dina(n18536), .dinb(a47 ), .dout(n18537));
  jxor g18279(.dina(n18537), .dinb(n18529), .dout(n18538));
  jor  g18280(.dina(n18356), .dinb(n18352), .dout(n18539));
  jand g18281(.dina(n18356), .dinb(n18352), .dout(n18540));
  jor  g18282(.dina(n18366), .dinb(n18540), .dout(n18541));
  jand g18283(.dina(n18541), .dinb(n18539), .dout(n18542));
  jxor g18284(.dina(n18542), .dinb(n18538), .dout(n18543));
  jnot g18285(.din(n18543), .dout(n18544));
  jor  g18286(.dina(n7146), .dinb(n5739), .dout(n18545));
  jor  g18287(.dina(n5574), .dinb(n6867), .dout(n18546));
  jor  g18288(.dina(n5742), .dinb(n7129), .dout(n18547));
  jor  g18289(.dina(n5744), .dinb(n7149), .dout(n18548));
  jand g18290(.dina(n18548), .dinb(n18547), .dout(n18549));
  jand g18291(.dina(n18549), .dinb(n18546), .dout(n18550));
  jand g18292(.dina(n18550), .dinb(n18545), .dout(n18551));
  jxor g18293(.dina(n18551), .dinb(a44 ), .dout(n18552));
  jxor g18294(.dina(n18552), .dinb(n18544), .dout(n18553));
  jxor g18295(.dina(n18553), .dinb(n18452), .dout(n18554));
  jxor g18296(.dina(n18554), .dinb(n18448), .dout(n18555));
  jxor g18297(.dina(n18555), .dinb(n18440), .dout(n18556));
  jnot g18298(.din(n18556), .dout(n18557));
  jor  g18299(.dina(n8806), .dinb(n4415), .dout(n18558));
  jor  g18300(.dina(n4272), .dinb(n8231), .dout(n18559));
  jor  g18301(.dina(n4418), .dinb(n8789), .dout(n18560));
  jor  g18302(.dina(n4420), .dinb(n8809), .dout(n18561));
  jand g18303(.dina(n18561), .dinb(n18560), .dout(n18562));
  jand g18304(.dina(n18562), .dinb(n18559), .dout(n18563));
  jand g18305(.dina(n18563), .dinb(n18558), .dout(n18564));
  jxor g18306(.dina(n18564), .dinb(a38 ), .dout(n18565));
  jxor g18307(.dina(n18565), .dinb(n18557), .dout(n18566));
  jxor g18308(.dina(n18566), .dinb(n18437), .dout(n18567));
  jnot g18309(.din(n18567), .dout(n18568));
  jor  g18310(.dina(n9722), .dinb(n3849), .dout(n18569));
  jor  g18311(.dina(n3689), .dinb(n9390), .dout(n18570));
  jor  g18312(.dina(n3852), .dinb(n9413), .dout(n18571));
  jor  g18313(.dina(n3854), .dinb(n9725), .dout(n18572));
  jand g18314(.dina(n18572), .dinb(n18571), .dout(n18573));
  jand g18315(.dina(n18573), .dinb(n18570), .dout(n18574));
  jand g18316(.dina(n18574), .dinb(n18569), .dout(n18575));
  jxor g18317(.dina(n18575), .dinb(a35 ), .dout(n18576));
  jxor g18318(.dina(n18576), .dinb(n18568), .dout(n18577));
  jor  g18319(.dina(n18401), .dinb(n18260), .dout(n18578));
  jand g18320(.dina(n18401), .dinb(n18260), .dout(n18579));
  jor  g18321(.dina(n18411), .dinb(n18579), .dout(n18580));
  jand g18322(.dina(n18580), .dinb(n18578), .dout(n18581));
  jxor g18323(.dina(n18581), .dinb(n18577), .dout(n18582));
  jand g18324(.dina(n18256), .dinb(n18252), .dout(n18583));
  jand g18325(.dina(n18412), .dinb(n18257), .dout(n18584));
  jor  g18326(.dina(n18584), .dinb(n18583), .dout(n18585));
  jnot g18327(.din(n18585), .dout(n18586));
  jor  g18328(.dina(n10961), .dinb(n3301), .dout(n18587));
  jor  g18329(.dina(n3136), .dinb(n10314), .dout(n18588));
  jor  g18330(.dina(n3304), .dinb(n10637), .dout(n18589));
  jor  g18331(.dina(n3306), .dinb(n10964), .dout(n18590));
  jand g18332(.dina(n18590), .dinb(n18589), .dout(n18591));
  jand g18333(.dina(n18591), .dinb(n18588), .dout(n18592));
  jand g18334(.dina(n18592), .dinb(n18587), .dout(n18593));
  jxor g18335(.dina(n18593), .dinb(a32 ), .dout(n18594));
  jxor g18336(.dina(n18594), .dinb(n18586), .dout(n18595));
  jxor g18337(.dina(n18595), .dinb(n18582), .dout(n18596));
  jxor g18338(.dina(n18596), .dinb(n18434), .dout(n18597));
  jxor g18339(.dina(n18597), .dinb(n18429), .dout(f93 ));
  jand g18340(.dina(n18596), .dinb(n18434), .dout(n18599));
  jand g18341(.dina(n18597), .dinb(n18429), .dout(n18600));
  jor  g18342(.dina(n18600), .dinb(n18599), .dout(n18601));
  jor  g18343(.dina(n18594), .dinb(n18586), .dout(n18602));
  jand g18344(.dina(n18595), .dinb(n18582), .dout(n18603));
  jnot g18345(.din(n18603), .dout(n18604));
  jand g18346(.dina(n18604), .dinb(n18602), .dout(n18605));
  jnot g18347(.din(n18605), .dout(n18606));
  jor  g18348(.dina(n18576), .dinb(n18568), .dout(n18607));
  jand g18349(.dina(n18581), .dinb(n18577), .dout(n18608));
  jnot g18350(.din(n18608), .dout(n18609));
  jand g18351(.dina(n18609), .dinb(n18607), .dout(n18610));
  jor  g18352(.dina(n10978), .dinb(n3301), .dout(n18611));
  jor  g18353(.dina(n3136), .dinb(n10637), .dout(n18612));
  jor  g18354(.dina(n3304), .dinb(n10964), .dout(n18613));
  jand g18355(.dina(n18613), .dinb(n18612), .dout(n18614));
  jand g18356(.dina(n18614), .dinb(n18611), .dout(n18615));
  jxor g18357(.dina(n18615), .dinb(a32 ), .dout(n18616));
  jxor g18358(.dina(n18616), .dinb(n18610), .dout(n18617));
  jor  g18359(.dina(n18565), .dinb(n18557), .dout(n18618));
  jand g18360(.dina(n18566), .dinb(n18437), .dout(n18619));
  jnot g18361(.din(n18619), .dout(n18620));
  jand g18362(.dina(n18620), .dinb(n18618), .dout(n18621));
  jnot g18363(.din(n18621), .dout(n18622));
  jor  g18364(.dina(n18554), .dinb(n18448), .dout(n18623));
  jand g18365(.dina(n18555), .dinb(n18440), .dout(n18624));
  jnot g18366(.din(n18624), .dout(n18625));
  jand g18367(.dina(n18625), .dinb(n18623), .dout(n18626));
  jnot g18368(.din(n18626), .dout(n18627));
  jor  g18369(.dina(n8228), .dinb(n5096), .dout(n18628));
  jor  g18370(.dina(n4904), .dinb(n7683), .dout(n18629));
  jor  g18371(.dina(n5099), .dinb(n7960), .dout(n18630));
  jor  g18372(.dina(n5101), .dinb(n8231), .dout(n18631));
  jand g18373(.dina(n18631), .dinb(n18630), .dout(n18632));
  jand g18374(.dina(n18632), .dinb(n18629), .dout(n18633));
  jand g18375(.dina(n18633), .dinb(n18628), .dout(n18634));
  jxor g18376(.dina(n18634), .dinb(a41 ), .dout(n18635));
  jnot g18377(.din(n18635), .dout(n18636));
  jor  g18378(.dina(n18537), .dinb(n18529), .dout(n18637));
  jand g18379(.dina(n18542), .dinb(n18538), .dout(n18638));
  jnot g18380(.din(n18638), .dout(n18639));
  jand g18381(.dina(n18639), .dinb(n18637), .dout(n18640));
  jnot g18382(.din(n18640), .dout(n18641));
  jand g18383(.dina(n18526), .dinb(n18464), .dout(n18642));
  jand g18384(.dina(n18527), .dinb(n18455), .dout(n18643));
  jor  g18385(.dina(n18643), .dinb(n18642), .dout(n18644));
  jor  g18386(.dina(n18524), .dinb(n18516), .dout(n18645));
  jand g18387(.dina(n18525), .dinb(n18467), .dout(n18646));
  jnot g18388(.din(n18646), .dout(n18647));
  jand g18389(.dina(n18647), .dinb(n18645), .dout(n18648));
  jnot g18390(.din(n18648), .dout(n18649));
  jor  g18391(.dina(n18509), .dinb(n18501), .dout(n18650));
  jand g18392(.dina(n18514), .dinb(n18510), .dout(n18651));
  jnot g18393(.din(n18651), .dout(n18652));
  jand g18394(.dina(n18652), .dinb(n18650), .dout(n18653));
  jnot g18395(.din(n18653), .dout(n18654));
  jor  g18396(.dina(n8978), .dinb(n4554), .dout(n18655));
  jor  g18397(.dina(n8677), .dinb(n4340), .dout(n18656));
  jor  g18398(.dina(n8981), .dinb(n4537), .dout(n18657));
  jor  g18399(.dina(n8983), .dinb(n4557), .dout(n18658));
  jand g18400(.dina(n18658), .dinb(n18657), .dout(n18659));
  jand g18401(.dina(n18659), .dinb(n18656), .dout(n18660));
  jand g18402(.dina(n18660), .dinb(n18655), .dout(n18661));
  jxor g18403(.dina(n18661), .dinb(a56 ), .dout(n18662));
  jnot g18404(.din(n18662), .dout(n18663));
  jand g18405(.dina(n18498), .dinb(n18479), .dout(n18664));
  jand g18406(.dina(n18499), .dinb(n18470), .dout(n18665));
  jor  g18407(.dina(n18665), .dinb(n18664), .dout(n18666));
  jor  g18408(.dina(n9891), .dinb(n4137), .dout(n18667));
  jor  g18409(.dina(n9593), .dinb(n3588), .dout(n18668));
  jor  g18410(.dina(n9894), .dinb(n3942), .dout(n18669));
  jor  g18411(.dina(n9896), .dinb(n4140), .dout(n18670));
  jand g18412(.dina(n18670), .dinb(n18669), .dout(n18671));
  jand g18413(.dina(n18671), .dinb(n18668), .dout(n18672));
  jand g18414(.dina(n18672), .dinb(n18667), .dout(n18673));
  jxor g18415(.dina(n18673), .dinb(a59 ), .dout(n18674));
  jnot g18416(.din(n18674), .dout(n18675));
  jand g18417(.dina(n18496), .dinb(n18491), .dout(n18676));
  jand g18418(.dina(n18497), .dinb(n18488), .dout(n18677));
  jor  g18419(.dina(n18677), .dinb(n18676), .dout(n18678));
  jand g18420(.dina(n18494), .dinb(n18418), .dout(n18679));
  jor  g18421(.dina(n18494), .dinb(n18418), .dout(n18680));
  jand g18422(.dina(n18680), .dinb(n18328), .dout(n18681));
  jor  g18423(.dina(n18681), .dinb(n18679), .dout(n18682));
  jand g18424(.dina(n10801), .dinb(b31 ), .dout(n18683));
  jand g18425(.dina(n11107), .dinb(b30 ), .dout(n18684));
  jor  g18426(.dina(n18684), .dinb(n18683), .dout(n18685));
  jnot g18427(.din(n18685), .dout(n18686));
  jxor g18428(.dina(n18686), .dinb(n18682), .dout(n18687));
  jnot g18429(.din(n18687), .dout(n18688));
  jor  g18430(.dina(n10806), .dinb(n3400), .dout(n18689));
  jor  g18431(.dina(n10485), .dinb(n3055), .dout(n18690));
  jor  g18432(.dina(n10809), .dinb(n3230), .dout(n18691));
  jor  g18433(.dina(n10811), .dinb(n3403), .dout(n18692));
  jand g18434(.dina(n18692), .dinb(n18691), .dout(n18693));
  jand g18435(.dina(n18693), .dinb(n18690), .dout(n18694));
  jand g18436(.dina(n18694), .dinb(n18689), .dout(n18695));
  jxor g18437(.dina(n18695), .dinb(a62 ), .dout(n18696));
  jxor g18438(.dina(n18696), .dinb(n18688), .dout(n18697));
  jxor g18439(.dina(n18697), .dinb(n18678), .dout(n18698));
  jxor g18440(.dina(n18698), .dinb(n18675), .dout(n18699));
  jxor g18441(.dina(n18699), .dinb(n18666), .dout(n18700));
  jxor g18442(.dina(n18700), .dinb(n18663), .dout(n18701));
  jxor g18443(.dina(n18701), .dinb(n18654), .dout(n18702));
  jor  g18444(.dina(n8125), .dinb(n5405), .dout(n18703));
  jor  g18445(.dina(n7846), .dinb(n4974), .dout(n18704));
  jor  g18446(.dina(n8128), .dinb(n4994), .dout(n18705));
  jor  g18447(.dina(n8130), .dinb(n5408), .dout(n18706));
  jand g18448(.dina(n18706), .dinb(n18705), .dout(n18707));
  jand g18449(.dina(n18707), .dinb(n18704), .dout(n18708));
  jand g18450(.dina(n18708), .dinb(n18703), .dout(n18709));
  jxor g18451(.dina(n18709), .dinb(a53 ), .dout(n18710));
  jnot g18452(.din(n18710), .dout(n18711));
  jxor g18453(.dina(n18711), .dinb(n18702), .dout(n18712));
  jxor g18454(.dina(n18712), .dinb(n18649), .dout(n18713));
  jor  g18455(.dina(n7266), .dinb(n6103), .dout(n18714));
  jor  g18456(.dina(n7021), .dinb(n5428), .dout(n18715));
  jor  g18457(.dina(n7269), .dinb(n5862), .dout(n18716));
  jor  g18458(.dina(n7271), .dinb(n6106), .dout(n18717));
  jand g18459(.dina(n18717), .dinb(n18716), .dout(n18718));
  jand g18460(.dina(n18718), .dinb(n18715), .dout(n18719));
  jand g18461(.dina(n18719), .dinb(n18714), .dout(n18720));
  jxor g18462(.dina(n18720), .dinb(a50 ), .dout(n18721));
  jnot g18463(.din(n18721), .dout(n18722));
  jxor g18464(.dina(n18722), .dinb(n18713), .dout(n18723));
  jxor g18465(.dina(n18723), .dinb(n18644), .dout(n18724));
  jor  g18466(.dina(n6864), .dinb(n6490), .dout(n18725));
  jor  g18467(.dina(n6262), .dinb(n6352), .dout(n18726));
  jor  g18468(.dina(n6493), .dinb(n6372), .dout(n18727));
  jor  g18469(.dina(n6495), .dinb(n6867), .dout(n18728));
  jand g18470(.dina(n18728), .dinb(n18727), .dout(n18729));
  jand g18471(.dina(n18729), .dinb(n18726), .dout(n18730));
  jand g18472(.dina(n18730), .dinb(n18725), .dout(n18731));
  jxor g18473(.dina(n18731), .dinb(a47 ), .dout(n18732));
  jnot g18474(.din(n18732), .dout(n18733));
  jxor g18475(.dina(n18733), .dinb(n18724), .dout(n18734));
  jxor g18476(.dina(n18734), .dinb(n18641), .dout(n18735));
  jor  g18477(.dina(n7408), .dinb(n5739), .dout(n18736));
  jor  g18478(.dina(n5574), .dinb(n7129), .dout(n18737));
  jor  g18479(.dina(n5742), .dinb(n7149), .dout(n18738));
  jor  g18480(.dina(n5744), .dinb(n7411), .dout(n18739));
  jand g18481(.dina(n18739), .dinb(n18738), .dout(n18740));
  jand g18482(.dina(n18740), .dinb(n18737), .dout(n18741));
  jand g18483(.dina(n18741), .dinb(n18736), .dout(n18742));
  jxor g18484(.dina(n18742), .dinb(a44 ), .dout(n18743));
  jnot g18485(.din(n18743), .dout(n18744));
  jxor g18486(.dina(n18744), .dinb(n18735), .dout(n18745));
  jand g18487(.dina(n18552), .dinb(n18544), .dout(n18746));
  jnot g18488(.din(n18552), .dout(n18747));
  jand g18489(.dina(n18747), .dinb(n18543), .dout(n18748));
  jnot g18490(.din(n18748), .dout(n18749));
  jand g18491(.dina(n18749), .dinb(n18452), .dout(n18750));
  jor  g18492(.dina(n18750), .dinb(n18746), .dout(n18751));
  jnot g18493(.din(n18751), .dout(n18752));
  jxor g18494(.dina(n18752), .dinb(n18745), .dout(n18753));
  jxor g18495(.dina(n18753), .dinb(n18636), .dout(n18754));
  jxor g18496(.dina(n18754), .dinb(n18627), .dout(n18755));
  jor  g18497(.dina(n9387), .dinb(n4415), .dout(n18756));
  jor  g18498(.dina(n4272), .dinb(n8789), .dout(n18757));
  jor  g18499(.dina(n4418), .dinb(n8809), .dout(n18758));
  jor  g18500(.dina(n4420), .dinb(n9390), .dout(n18759));
  jand g18501(.dina(n18759), .dinb(n18758), .dout(n18760));
  jand g18502(.dina(n18760), .dinb(n18757), .dout(n18761));
  jand g18503(.dina(n18761), .dinb(n18756), .dout(n18762));
  jxor g18504(.dina(n18762), .dinb(a38 ), .dout(n18763));
  jnot g18505(.din(n18763), .dout(n18764));
  jxor g18506(.dina(n18764), .dinb(n18755), .dout(n18765));
  jxor g18507(.dina(n18765), .dinb(n18622), .dout(n18766));
  jnot g18508(.din(n18766), .dout(n18767));
  jor  g18509(.dina(n10311), .dinb(n3849), .dout(n18768));
  jor  g18510(.dina(n3689), .dinb(n9413), .dout(n18769));
  jor  g18511(.dina(n3852), .dinb(n9725), .dout(n18770));
  jor  g18512(.dina(n3854), .dinb(n10314), .dout(n18771));
  jand g18513(.dina(n18771), .dinb(n18770), .dout(n18772));
  jand g18514(.dina(n18772), .dinb(n18769), .dout(n18773));
  jand g18515(.dina(n18773), .dinb(n18768), .dout(n18774));
  jxor g18516(.dina(n18774), .dinb(a35 ), .dout(n18775));
  jxor g18517(.dina(n18775), .dinb(n18767), .dout(n18776));
  jxor g18518(.dina(n18776), .dinb(n18617), .dout(n18777));
  jxor g18519(.dina(n18777), .dinb(n18606), .dout(n18778));
  jxor g18520(.dina(n18778), .dinb(n18601), .dout(f94 ));
  jand g18521(.dina(n18777), .dinb(n18606), .dout(n18780));
  jand g18522(.dina(n18778), .dinb(n18601), .dout(n18781));
  jor  g18523(.dina(n18781), .dinb(n18780), .dout(n18782));
  jor  g18524(.dina(n18616), .dinb(n18610), .dout(n18783));
  jand g18525(.dina(n18776), .dinb(n18617), .dout(n18784));
  jnot g18526(.din(n18784), .dout(n18785));
  jand g18527(.dina(n18785), .dinb(n18783), .dout(n18786));
  jnot g18528(.din(n18786), .dout(n18787));
  jand g18529(.dina(n18765), .dinb(n18622), .dout(n18788));
  jnot g18530(.din(n18788), .dout(n18789));
  jor  g18531(.dina(n18775), .dinb(n18767), .dout(n18790));
  jand g18532(.dina(n18790), .dinb(n18789), .dout(n18791));
  jnot g18533(.din(a32 ), .dout(n18792));
  jand g18534(.dina(n11296), .dinb(n2941), .dout(n18793));
  jor  g18535(.dina(n18793), .dinb(n3137), .dout(n18794));
  jand g18536(.dina(n18794), .dinb(b63 ), .dout(n18795));
  jxor g18537(.dina(n18795), .dinb(n18792), .dout(n18796));
  jxor g18538(.dina(n18796), .dinb(n18791), .dout(n18797));
  jand g18539(.dina(n18752), .dinb(n18745), .dout(n18798));
  jand g18540(.dina(n18753), .dinb(n18636), .dout(n18799));
  jor  g18541(.dina(n18799), .dinb(n18798), .dout(n18800));
  jor  g18542(.dina(n8786), .dinb(n5096), .dout(n18801));
  jor  g18543(.dina(n4904), .dinb(n7960), .dout(n18802));
  jor  g18544(.dina(n5099), .dinb(n8231), .dout(n18803));
  jor  g18545(.dina(n5101), .dinb(n8789), .dout(n18804));
  jand g18546(.dina(n18804), .dinb(n18803), .dout(n18805));
  jand g18547(.dina(n18805), .dinb(n18802), .dout(n18806));
  jand g18548(.dina(n18806), .dinb(n18801), .dout(n18807));
  jxor g18549(.dina(n18807), .dinb(a41 ), .dout(n18808));
  jnot g18550(.din(n18808), .dout(n18809));
  jor  g18551(.dina(n7680), .dinb(n5739), .dout(n18810));
  jor  g18552(.dina(n5574), .dinb(n7149), .dout(n18811));
  jor  g18553(.dina(n5742), .dinb(n7411), .dout(n18812));
  jor  g18554(.dina(n5744), .dinb(n7683), .dout(n18813));
  jand g18555(.dina(n18813), .dinb(n18812), .dout(n18814));
  jand g18556(.dina(n18814), .dinb(n18811), .dout(n18815));
  jand g18557(.dina(n18815), .dinb(n18810), .dout(n18816));
  jxor g18558(.dina(n18816), .dinb(a44 ), .dout(n18817));
  jnot g18559(.din(n18817), .dout(n18818));
  jor  g18560(.dina(n8125), .dinb(n5425), .dout(n18819));
  jor  g18561(.dina(n7846), .dinb(n4994), .dout(n18820));
  jor  g18562(.dina(n8128), .dinb(n5408), .dout(n18821));
  jor  g18563(.dina(n8130), .dinb(n5428), .dout(n18822));
  jand g18564(.dina(n18822), .dinb(n18821), .dout(n18823));
  jand g18565(.dina(n18823), .dinb(n18820), .dout(n18824));
  jand g18566(.dina(n18824), .dinb(n18819), .dout(n18825));
  jxor g18567(.dina(n18825), .dinb(a53 ), .dout(n18826));
  jnot g18568(.din(n18826), .dout(n18827));
  jand g18569(.dina(n18699), .dinb(n18666), .dout(n18828));
  jand g18570(.dina(n18700), .dinb(n18663), .dout(n18829));
  jor  g18571(.dina(n18829), .dinb(n18828), .dout(n18830));
  jor  g18572(.dina(n8978), .dinb(n4971), .dout(n18831));
  jor  g18573(.dina(n8677), .dinb(n4537), .dout(n18832));
  jor  g18574(.dina(n8981), .dinb(n4557), .dout(n18833));
  jor  g18575(.dina(n8983), .dinb(n4974), .dout(n18834));
  jand g18576(.dina(n18834), .dinb(n18833), .dout(n18835));
  jand g18577(.dina(n18835), .dinb(n18832), .dout(n18836));
  jand g18578(.dina(n18836), .dinb(n18831), .dout(n18837));
  jxor g18579(.dina(n18837), .dinb(a56 ), .dout(n18838));
  jnot g18580(.din(n18838), .dout(n18839));
  jand g18581(.dina(n18697), .dinb(n18678), .dout(n18840));
  jand g18582(.dina(n18698), .dinb(n18675), .dout(n18841));
  jor  g18583(.dina(n18841), .dinb(n18840), .dout(n18842));
  jor  g18584(.dina(n9891), .dinb(n4337), .dout(n18843));
  jor  g18585(.dina(n9593), .dinb(n3942), .dout(n18844));
  jor  g18586(.dina(n9894), .dinb(n4140), .dout(n18845));
  jor  g18587(.dina(n9896), .dinb(n4340), .dout(n18846));
  jand g18588(.dina(n18846), .dinb(n18845), .dout(n18847));
  jand g18589(.dina(n18847), .dinb(n18844), .dout(n18848));
  jand g18590(.dina(n18848), .dinb(n18843), .dout(n18849));
  jxor g18591(.dina(n18849), .dinb(a59 ), .dout(n18850));
  jnot g18592(.din(n18850), .dout(n18851));
  jand g18593(.dina(n18686), .dinb(n18682), .dout(n18852));
  jnot g18594(.din(n18852), .dout(n18853));
  jor  g18595(.dina(n18696), .dinb(n18688), .dout(n18854));
  jand g18596(.dina(n18854), .dinb(n18853), .dout(n18855));
  jnot g18597(.din(n18855), .dout(n18856));
  jand g18598(.dina(n10801), .dinb(b32 ), .dout(n18857));
  jand g18599(.dina(n11107), .dinb(b31 ), .dout(n18858));
  jor  g18600(.dina(n18858), .dinb(n18857), .dout(n18859));
  jnot g18601(.din(n18859), .dout(n18860));
  jxor g18602(.dina(n18860), .dinb(n18685), .dout(n18861));
  jxor g18603(.dina(n18861), .dinb(n18856), .dout(n18862));
  jnot g18604(.din(n18862), .dout(n18863));
  jor  g18605(.dina(n10806), .dinb(n3585), .dout(n18864));
  jor  g18606(.dina(n10485), .dinb(n3230), .dout(n18865));
  jor  g18607(.dina(n10809), .dinb(n3403), .dout(n18866));
  jor  g18608(.dina(n10811), .dinb(n3588), .dout(n18867));
  jand g18609(.dina(n18867), .dinb(n18866), .dout(n18868));
  jand g18610(.dina(n18868), .dinb(n18865), .dout(n18869));
  jand g18611(.dina(n18869), .dinb(n18864), .dout(n18870));
  jxor g18612(.dina(n18870), .dinb(a62 ), .dout(n18871));
  jxor g18613(.dina(n18871), .dinb(n18863), .dout(n18872));
  jxor g18614(.dina(n18872), .dinb(n18851), .dout(n18873));
  jxor g18615(.dina(n18873), .dinb(n18842), .dout(n18874));
  jxor g18616(.dina(n18874), .dinb(n18839), .dout(n18875));
  jxor g18617(.dina(n18875), .dinb(n18830), .dout(n18876));
  jxor g18618(.dina(n18876), .dinb(n18827), .dout(n18877));
  jor  g18619(.dina(n18701), .dinb(n18654), .dout(n18878));
  jand g18620(.dina(n18701), .dinb(n18654), .dout(n18879));
  jor  g18621(.dina(n18711), .dinb(n18879), .dout(n18880));
  jand g18622(.dina(n18880), .dinb(n18878), .dout(n18881));
  jxor g18623(.dina(n18881), .dinb(n18877), .dout(n18882));
  jor  g18624(.dina(n7266), .dinb(n6349), .dout(n18883));
  jor  g18625(.dina(n7021), .dinb(n5862), .dout(n18884));
  jor  g18626(.dina(n7269), .dinb(n6106), .dout(n18885));
  jor  g18627(.dina(n7271), .dinb(n6352), .dout(n18886));
  jand g18628(.dina(n18886), .dinb(n18885), .dout(n18887));
  jand g18629(.dina(n18887), .dinb(n18884), .dout(n18888));
  jand g18630(.dina(n18888), .dinb(n18883), .dout(n18889));
  jxor g18631(.dina(n18889), .dinb(a50 ), .dout(n18890));
  jnot g18632(.din(n18890), .dout(n18891));
  jxor g18633(.dina(n18891), .dinb(n18882), .dout(n18892));
  jnot g18634(.din(n18712), .dout(n18893));
  jand g18635(.dina(n18893), .dinb(n18648), .dout(n18894));
  jnot g18636(.din(n18894), .dout(n18895));
  jand g18637(.dina(n18712), .dinb(n18649), .dout(n18896));
  jor  g18638(.dina(n18722), .dinb(n18896), .dout(n18897));
  jand g18639(.dina(n18897), .dinb(n18895), .dout(n18898));
  jxor g18640(.dina(n18898), .dinb(n18892), .dout(n18899));
  jnot g18641(.din(n18899), .dout(n18900));
  jor  g18642(.dina(n7126), .dinb(n6490), .dout(n18901));
  jor  g18643(.dina(n6262), .dinb(n6372), .dout(n18902));
  jor  g18644(.dina(n6493), .dinb(n6867), .dout(n18903));
  jor  g18645(.dina(n6495), .dinb(n7129), .dout(n18904));
  jand g18646(.dina(n18904), .dinb(n18903), .dout(n18905));
  jand g18647(.dina(n18905), .dinb(n18902), .dout(n18906));
  jand g18648(.dina(n18906), .dinb(n18901), .dout(n18907));
  jxor g18649(.dina(n18907), .dinb(a47 ), .dout(n18908));
  jxor g18650(.dina(n18908), .dinb(n18900), .dout(n18909));
  jnot g18651(.din(n18644), .dout(n18910));
  jnot g18652(.din(n18723), .dout(n18911));
  jand g18653(.dina(n18911), .dinb(n18910), .dout(n18912));
  jnot g18654(.din(n18912), .dout(n18913));
  jand g18655(.dina(n18723), .dinb(n18644), .dout(n18914));
  jor  g18656(.dina(n18733), .dinb(n18914), .dout(n18915));
  jand g18657(.dina(n18915), .dinb(n18913), .dout(n18916));
  jxor g18658(.dina(n18916), .dinb(n18909), .dout(n18917));
  jxor g18659(.dina(n18917), .dinb(n18818), .dout(n18918));
  jnot g18660(.din(n18734), .dout(n18919));
  jand g18661(.dina(n18919), .dinb(n18640), .dout(n18920));
  jnot g18662(.din(n18920), .dout(n18921));
  jand g18663(.dina(n18734), .dinb(n18641), .dout(n18922));
  jor  g18664(.dina(n18744), .dinb(n18922), .dout(n18923));
  jand g18665(.dina(n18923), .dinb(n18921), .dout(n18924));
  jxor g18666(.dina(n18924), .dinb(n18918), .dout(n18925));
  jxor g18667(.dina(n18925), .dinb(n18809), .dout(n18926));
  jxor g18668(.dina(n18926), .dinb(n18800), .dout(n18927));
  jor  g18669(.dina(n9410), .dinb(n4415), .dout(n18928));
  jor  g18670(.dina(n4272), .dinb(n8809), .dout(n18929));
  jor  g18671(.dina(n4418), .dinb(n9390), .dout(n18930));
  jor  g18672(.dina(n4420), .dinb(n9413), .dout(n18931));
  jand g18673(.dina(n18931), .dinb(n18930), .dout(n18932));
  jand g18674(.dina(n18932), .dinb(n18929), .dout(n18933));
  jand g18675(.dina(n18933), .dinb(n18928), .dout(n18934));
  jxor g18676(.dina(n18934), .dinb(a38 ), .dout(n18935));
  jnot g18677(.din(n18935), .dout(n18936));
  jxor g18678(.dina(n18936), .dinb(n18927), .dout(n18937));
  jor  g18679(.dina(n18754), .dinb(n18627), .dout(n18938));
  jand g18680(.dina(n18754), .dinb(n18627), .dout(n18939));
  jor  g18681(.dina(n18764), .dinb(n18939), .dout(n18940));
  jand g18682(.dina(n18940), .dinb(n18938), .dout(n18941));
  jxor g18683(.dina(n18941), .dinb(n18937), .dout(n18942));
  jor  g18684(.dina(n10634), .dinb(n3849), .dout(n18943));
  jor  g18685(.dina(n3689), .dinb(n9725), .dout(n18944));
  jor  g18686(.dina(n3852), .dinb(n10314), .dout(n18945));
  jor  g18687(.dina(n3854), .dinb(n10637), .dout(n18946));
  jand g18688(.dina(n18946), .dinb(n18945), .dout(n18947));
  jand g18689(.dina(n18947), .dinb(n18944), .dout(n18948));
  jand g18690(.dina(n18948), .dinb(n18943), .dout(n18949));
  jxor g18691(.dina(n18949), .dinb(a35 ), .dout(n18950));
  jnot g18692(.din(n18950), .dout(n18951));
  jxor g18693(.dina(n18951), .dinb(n18942), .dout(n18952));
  jxor g18694(.dina(n18952), .dinb(n18797), .dout(n18953));
  jxor g18695(.dina(n18953), .dinb(n18787), .dout(n18954));
  jxor g18696(.dina(n18954), .dinb(n18782), .dout(f95 ));
  jand g18697(.dina(n18953), .dinb(n18787), .dout(n18956));
  jand g18698(.dina(n18954), .dinb(n18782), .dout(n18957));
  jor  g18699(.dina(n18957), .dinb(n18956), .dout(n18958));
  jor  g18700(.dina(n18796), .dinb(n18791), .dout(n18959));
  jand g18701(.dina(n18952), .dinb(n18797), .dout(n18960));
  jnot g18702(.din(n18960), .dout(n18961));
  jand g18703(.dina(n18961), .dinb(n18959), .dout(n18962));
  jnot g18704(.din(n18962), .dout(n18963));
  jand g18705(.dina(n18924), .dinb(n18918), .dout(n18964));
  jand g18706(.dina(n18925), .dinb(n18809), .dout(n18965));
  jor  g18707(.dina(n18965), .dinb(n18964), .dout(n18966));
  jand g18708(.dina(n18916), .dinb(n18909), .dout(n18967));
  jand g18709(.dina(n18917), .dinb(n18818), .dout(n18968));
  jor  g18710(.dina(n18968), .dinb(n18967), .dout(n18969));
  jor  g18711(.dina(n7957), .dinb(n5739), .dout(n18970));
  jor  g18712(.dina(n5574), .dinb(n7411), .dout(n18971));
  jor  g18713(.dina(n5742), .dinb(n7683), .dout(n18972));
  jor  g18714(.dina(n5744), .dinb(n7960), .dout(n18973));
  jand g18715(.dina(n18973), .dinb(n18972), .dout(n18974));
  jand g18716(.dina(n18974), .dinb(n18971), .dout(n18975));
  jand g18717(.dina(n18975), .dinb(n18970), .dout(n18976));
  jxor g18718(.dina(n18976), .dinb(a44 ), .dout(n18977));
  jand g18719(.dina(n18898), .dinb(n18892), .dout(n18978));
  jnot g18720(.din(n18978), .dout(n18979));
  jor  g18721(.dina(n18908), .dinb(n18900), .dout(n18980));
  jand g18722(.dina(n18980), .dinb(n18979), .dout(n18981));
  jand g18723(.dina(n18875), .dinb(n18830), .dout(n18982));
  jand g18724(.dina(n18876), .dinb(n18827), .dout(n18983));
  jor  g18725(.dina(n18983), .dinb(n18982), .dout(n18984));
  jand g18726(.dina(n18873), .dinb(n18842), .dout(n18985));
  jand g18727(.dina(n18874), .dinb(n18839), .dout(n18986));
  jor  g18728(.dina(n18986), .dinb(n18985), .dout(n18987));
  jor  g18729(.dina(n18871), .dinb(n18863), .dout(n18988));
  jand g18730(.dina(n18872), .dinb(n18851), .dout(n18989));
  jnot g18731(.din(n18989), .dout(n18990));
  jand g18732(.dina(n18990), .dinb(n18988), .dout(n18991));
  jnot g18733(.din(n18991), .dout(n18992));
  jor  g18734(.dina(n9891), .dinb(n4534), .dout(n18993));
  jor  g18735(.dina(n9593), .dinb(n4140), .dout(n18994));
  jor  g18736(.dina(n9894), .dinb(n4340), .dout(n18995));
  jor  g18737(.dina(n9896), .dinb(n4537), .dout(n18996));
  jand g18738(.dina(n18996), .dinb(n18995), .dout(n18997));
  jand g18739(.dina(n18997), .dinb(n18994), .dout(n18998));
  jand g18740(.dina(n18998), .dinb(n18993), .dout(n18999));
  jxor g18741(.dina(n18999), .dinb(a59 ), .dout(n19000));
  jnot g18742(.din(n19000), .dout(n19001));
  jor  g18743(.dina(n10806), .dinb(n3939), .dout(n19002));
  jor  g18744(.dina(n10485), .dinb(n3403), .dout(n19003));
  jor  g18745(.dina(n10809), .dinb(n3588), .dout(n19004));
  jor  g18746(.dina(n10811), .dinb(n3942), .dout(n19005));
  jand g18747(.dina(n19005), .dinb(n19004), .dout(n19006));
  jand g18748(.dina(n19006), .dinb(n19003), .dout(n19007));
  jand g18749(.dina(n19007), .dinb(n19002), .dout(n19008));
  jxor g18750(.dina(n19008), .dinb(a62 ), .dout(n19009));
  jnot g18751(.din(n19009), .dout(n19010));
  jand g18752(.dina(n18860), .dinb(n18685), .dout(n19011));
  jand g18753(.dina(n18861), .dinb(n18856), .dout(n19012));
  jor  g18754(.dina(n19012), .dinb(n19011), .dout(n19013));
  jand g18755(.dina(n10801), .dinb(b33 ), .dout(n19014));
  jand g18756(.dina(n11107), .dinb(b32 ), .dout(n19015));
  jor  g18757(.dina(n19015), .dinb(n19014), .dout(n19016));
  jxor g18758(.dina(n19016), .dinb(n18792), .dout(n19017));
  jxor g18759(.dina(n19017), .dinb(n18859), .dout(n19018));
  jxor g18760(.dina(n19018), .dinb(n19013), .dout(n19019));
  jxor g18761(.dina(n19019), .dinb(n19010), .dout(n19020));
  jxor g18762(.dina(n19020), .dinb(n19001), .dout(n19021));
  jxor g18763(.dina(n19021), .dinb(n18992), .dout(n19022));
  jnot g18764(.din(n19022), .dout(n19023));
  jor  g18765(.dina(n8978), .dinb(n4991), .dout(n19024));
  jor  g18766(.dina(n8677), .dinb(n4557), .dout(n19025));
  jor  g18767(.dina(n8981), .dinb(n4974), .dout(n19026));
  jor  g18768(.dina(n8983), .dinb(n4994), .dout(n19027));
  jand g18769(.dina(n19027), .dinb(n19026), .dout(n19028));
  jand g18770(.dina(n19028), .dinb(n19025), .dout(n19029));
  jand g18771(.dina(n19029), .dinb(n19024), .dout(n19030));
  jxor g18772(.dina(n19030), .dinb(a56 ), .dout(n19031));
  jxor g18773(.dina(n19031), .dinb(n19023), .dout(n19032));
  jxor g18774(.dina(n19032), .dinb(n18987), .dout(n19033));
  jnot g18775(.din(n19033), .dout(n19034));
  jor  g18776(.dina(n8125), .dinb(n5859), .dout(n19035));
  jor  g18777(.dina(n7846), .dinb(n5408), .dout(n19036));
  jor  g18778(.dina(n8128), .dinb(n5428), .dout(n19037));
  jor  g18779(.dina(n8130), .dinb(n5862), .dout(n19038));
  jand g18780(.dina(n19038), .dinb(n19037), .dout(n19039));
  jand g18781(.dina(n19039), .dinb(n19036), .dout(n19040));
  jand g18782(.dina(n19040), .dinb(n19035), .dout(n19041));
  jxor g18783(.dina(n19041), .dinb(a53 ), .dout(n19042));
  jxor g18784(.dina(n19042), .dinb(n19034), .dout(n19043));
  jxor g18785(.dina(n19043), .dinb(n18984), .dout(n19044));
  jnot g18786(.din(n19044), .dout(n19045));
  jor  g18787(.dina(n7266), .dinb(n6369), .dout(n19046));
  jor  g18788(.dina(n7021), .dinb(n6106), .dout(n19047));
  jor  g18789(.dina(n7269), .dinb(n6352), .dout(n19048));
  jor  g18790(.dina(n7271), .dinb(n6372), .dout(n19049));
  jand g18791(.dina(n19049), .dinb(n19048), .dout(n19050));
  jand g18792(.dina(n19050), .dinb(n19047), .dout(n19051));
  jand g18793(.dina(n19051), .dinb(n19046), .dout(n19052));
  jxor g18794(.dina(n19052), .dinb(a50 ), .dout(n19053));
  jxor g18795(.dina(n19053), .dinb(n19045), .dout(n19054));
  jor  g18796(.dina(n18881), .dinb(n18877), .dout(n19055));
  jand g18797(.dina(n18881), .dinb(n18877), .dout(n19056));
  jor  g18798(.dina(n18891), .dinb(n19056), .dout(n19057));
  jand g18799(.dina(n19057), .dinb(n19055), .dout(n19058));
  jxor g18800(.dina(n19058), .dinb(n19054), .dout(n19059));
  jnot g18801(.din(n19059), .dout(n19060));
  jor  g18802(.dina(n7146), .dinb(n6490), .dout(n19061));
  jor  g18803(.dina(n6262), .dinb(n6867), .dout(n19062));
  jor  g18804(.dina(n6493), .dinb(n7129), .dout(n19063));
  jor  g18805(.dina(n6495), .dinb(n7149), .dout(n19064));
  jand g18806(.dina(n19064), .dinb(n19063), .dout(n19065));
  jand g18807(.dina(n19065), .dinb(n19062), .dout(n19066));
  jand g18808(.dina(n19066), .dinb(n19061), .dout(n19067));
  jxor g18809(.dina(n19067), .dinb(a47 ), .dout(n19068));
  jxor g18810(.dina(n19068), .dinb(n19060), .dout(n19069));
  jxor g18811(.dina(n19069), .dinb(n18981), .dout(n19070));
  jxor g18812(.dina(n19070), .dinb(n18977), .dout(n19071));
  jxor g18813(.dina(n19071), .dinb(n18969), .dout(n19072));
  jnot g18814(.din(n19072), .dout(n19073));
  jor  g18815(.dina(n8806), .dinb(n5096), .dout(n19074));
  jor  g18816(.dina(n4904), .dinb(n8231), .dout(n19075));
  jor  g18817(.dina(n5099), .dinb(n8789), .dout(n19076));
  jor  g18818(.dina(n5101), .dinb(n8809), .dout(n19077));
  jand g18819(.dina(n19077), .dinb(n19076), .dout(n19078));
  jand g18820(.dina(n19078), .dinb(n19075), .dout(n19079));
  jand g18821(.dina(n19079), .dinb(n19074), .dout(n19080));
  jxor g18822(.dina(n19080), .dinb(a41 ), .dout(n19081));
  jxor g18823(.dina(n19081), .dinb(n19073), .dout(n19082));
  jxor g18824(.dina(n19082), .dinb(n18966), .dout(n19083));
  jnot g18825(.din(n19083), .dout(n19084));
  jor  g18826(.dina(n9722), .dinb(n4415), .dout(n19085));
  jor  g18827(.dina(n4272), .dinb(n9390), .dout(n19086));
  jor  g18828(.dina(n4418), .dinb(n9413), .dout(n19087));
  jor  g18829(.dina(n4420), .dinb(n9725), .dout(n19088));
  jand g18830(.dina(n19088), .dinb(n19087), .dout(n19089));
  jand g18831(.dina(n19089), .dinb(n19086), .dout(n19090));
  jand g18832(.dina(n19090), .dinb(n19085), .dout(n19091));
  jxor g18833(.dina(n19091), .dinb(a38 ), .dout(n19092));
  jxor g18834(.dina(n19092), .dinb(n19084), .dout(n19093));
  jor  g18835(.dina(n18926), .dinb(n18800), .dout(n19094));
  jand g18836(.dina(n18926), .dinb(n18800), .dout(n19095));
  jor  g18837(.dina(n18936), .dinb(n19095), .dout(n19096));
  jand g18838(.dina(n19096), .dinb(n19094), .dout(n19097));
  jxor g18839(.dina(n19097), .dinb(n19093), .dout(n19098));
  jor  g18840(.dina(n10961), .dinb(n3849), .dout(n19099));
  jor  g18841(.dina(n3689), .dinb(n10314), .dout(n19100));
  jor  g18842(.dina(n3852), .dinb(n10637), .dout(n19101));
  jor  g18843(.dina(n3854), .dinb(n10964), .dout(n19102));
  jand g18844(.dina(n19102), .dinb(n19101), .dout(n19103));
  jand g18845(.dina(n19103), .dinb(n19100), .dout(n19104));
  jand g18846(.dina(n19104), .dinb(n19099), .dout(n19105));
  jxor g18847(.dina(n19105), .dinb(a35 ), .dout(n19106));
  jnot g18848(.din(n19106), .dout(n19107));
  jnot g18849(.din(n18937), .dout(n19108));
  jnot g18850(.din(n18941), .dout(n19109));
  jand g18851(.dina(n19109), .dinb(n19108), .dout(n19110));
  jnot g18852(.din(n19110), .dout(n19111));
  jand g18853(.dina(n18941), .dinb(n18937), .dout(n19112));
  jor  g18854(.dina(n18951), .dinb(n19112), .dout(n19113));
  jand g18855(.dina(n19113), .dinb(n19111), .dout(n19114));
  jxor g18856(.dina(n19114), .dinb(n19107), .dout(n19115));
  jxor g18857(.dina(n19115), .dinb(n19098), .dout(n19116));
  jxor g18858(.dina(n19116), .dinb(n18963), .dout(n19117));
  jxor g18859(.dina(n19117), .dinb(n18958), .dout(f96 ));
  jand g18860(.dina(n19116), .dinb(n18963), .dout(n19119));
  jand g18861(.dina(n19117), .dinb(n18958), .dout(n19120));
  jor  g18862(.dina(n19120), .dinb(n19119), .dout(n19121));
  jand g18863(.dina(n19114), .dinb(n19107), .dout(n19122));
  jand g18864(.dina(n19115), .dinb(n19098), .dout(n19123));
  jor  g18865(.dina(n19123), .dinb(n19122), .dout(n19124));
  jor  g18866(.dina(n19092), .dinb(n19084), .dout(n19125));
  jand g18867(.dina(n19097), .dinb(n19093), .dout(n19126));
  jnot g18868(.din(n19126), .dout(n19127));
  jand g18869(.dina(n19127), .dinb(n19125), .dout(n19128));
  jor  g18870(.dina(n10978), .dinb(n3849), .dout(n19129));
  jor  g18871(.dina(n3689), .dinb(n10637), .dout(n19130));
  jor  g18872(.dina(n3852), .dinb(n10964), .dout(n19131));
  jand g18873(.dina(n19131), .dinb(n19130), .dout(n19132));
  jand g18874(.dina(n19132), .dinb(n19129), .dout(n19133));
  jxor g18875(.dina(n19133), .dinb(a35 ), .dout(n19134));
  jxor g18876(.dina(n19134), .dinb(n19128), .dout(n19135));
  jor  g18877(.dina(n19081), .dinb(n19073), .dout(n19136));
  jand g18878(.dina(n19082), .dinb(n18966), .dout(n19137));
  jnot g18879(.din(n19137), .dout(n19138));
  jand g18880(.dina(n19138), .dinb(n19136), .dout(n19139));
  jnot g18881(.din(n19139), .dout(n19140));
  jor  g18882(.dina(n19070), .dinb(n18977), .dout(n19141));
  jand g18883(.dina(n19071), .dinb(n18969), .dout(n19142));
  jnot g18884(.din(n19142), .dout(n19143));
  jand g18885(.dina(n19143), .dinb(n19141), .dout(n19144));
  jnot g18886(.din(n19144), .dout(n19145));
  jor  g18887(.dina(n8228), .dinb(n5739), .dout(n19146));
  jor  g18888(.dina(n5574), .dinb(n7683), .dout(n19147));
  jor  g18889(.dina(n5742), .dinb(n7960), .dout(n19148));
  jor  g18890(.dina(n5744), .dinb(n8231), .dout(n19149));
  jand g18891(.dina(n19149), .dinb(n19148), .dout(n19150));
  jand g18892(.dina(n19150), .dinb(n19147), .dout(n19151));
  jand g18893(.dina(n19151), .dinb(n19146), .dout(n19152));
  jxor g18894(.dina(n19152), .dinb(a44 ), .dout(n19153));
  jnot g18895(.din(n19153), .dout(n19154));
  jor  g18896(.dina(n19053), .dinb(n19045), .dout(n19155));
  jand g18897(.dina(n19058), .dinb(n19054), .dout(n19156));
  jnot g18898(.din(n19156), .dout(n19157));
  jand g18899(.dina(n19157), .dinb(n19155), .dout(n19158));
  jnot g18900(.din(n19158), .dout(n19159));
  jor  g18901(.dina(n19042), .dinb(n19034), .dout(n19160));
  jand g18902(.dina(n19043), .dinb(n18984), .dout(n19161));
  jnot g18903(.din(n19161), .dout(n19162));
  jand g18904(.dina(n19162), .dinb(n19160), .dout(n19163));
  jnot g18905(.din(n19163), .dout(n19164));
  jor  g18906(.dina(n19031), .dinb(n19023), .dout(n19165));
  jand g18907(.dina(n19032), .dinb(n18987), .dout(n19166));
  jnot g18908(.din(n19166), .dout(n19167));
  jand g18909(.dina(n19167), .dinb(n19165), .dout(n19168));
  jnot g18910(.din(n19168), .dout(n19169));
  jand g18911(.dina(n19020), .dinb(n19001), .dout(n19170));
  jand g18912(.dina(n19021), .dinb(n18992), .dout(n19171));
  jor  g18913(.dina(n19171), .dinb(n19170), .dout(n19172));
  jor  g18914(.dina(n9891), .dinb(n4554), .dout(n19173));
  jor  g18915(.dina(n9593), .dinb(n4340), .dout(n19174));
  jor  g18916(.dina(n9894), .dinb(n4537), .dout(n19175));
  jor  g18917(.dina(n9896), .dinb(n4557), .dout(n19176));
  jand g18918(.dina(n19176), .dinb(n19175), .dout(n19177));
  jand g18919(.dina(n19177), .dinb(n19174), .dout(n19178));
  jand g18920(.dina(n19178), .dinb(n19173), .dout(n19179));
  jxor g18921(.dina(n19179), .dinb(a59 ), .dout(n19180));
  jnot g18922(.din(n19180), .dout(n19181));
  jand g18923(.dina(n19018), .dinb(n19013), .dout(n19182));
  jand g18924(.dina(n19019), .dinb(n19010), .dout(n19183));
  jor  g18925(.dina(n19183), .dinb(n19182), .dout(n19184));
  jand g18926(.dina(n19016), .dinb(n18792), .dout(n19185));
  jor  g18927(.dina(n19016), .dinb(n18792), .dout(n19186));
  jand g18928(.dina(n19186), .dinb(n18859), .dout(n19187));
  jor  g18929(.dina(n19187), .dinb(n19185), .dout(n19188));
  jand g18930(.dina(n10801), .dinb(b34 ), .dout(n19189));
  jand g18931(.dina(n11107), .dinb(b33 ), .dout(n19190));
  jor  g18932(.dina(n19190), .dinb(n19189), .dout(n19191));
  jnot g18933(.din(n19191), .dout(n19192));
  jxor g18934(.dina(n19192), .dinb(n19188), .dout(n19193));
  jnot g18935(.din(n19193), .dout(n19194));
  jor  g18936(.dina(n10806), .dinb(n4137), .dout(n19195));
  jor  g18937(.dina(n10485), .dinb(n3588), .dout(n19196));
  jor  g18938(.dina(n10809), .dinb(n3942), .dout(n19197));
  jor  g18939(.dina(n10811), .dinb(n4140), .dout(n19198));
  jand g18940(.dina(n19198), .dinb(n19197), .dout(n19199));
  jand g18941(.dina(n19199), .dinb(n19196), .dout(n19200));
  jand g18942(.dina(n19200), .dinb(n19195), .dout(n19201));
  jxor g18943(.dina(n19201), .dinb(a62 ), .dout(n19202));
  jxor g18944(.dina(n19202), .dinb(n19194), .dout(n19203));
  jxor g18945(.dina(n19203), .dinb(n19184), .dout(n19204));
  jxor g18946(.dina(n19204), .dinb(n19181), .dout(n19205));
  jxor g18947(.dina(n19205), .dinb(n19172), .dout(n19206));
  jor  g18948(.dina(n8978), .dinb(n5405), .dout(n19207));
  jor  g18949(.dina(n8677), .dinb(n4974), .dout(n19208));
  jor  g18950(.dina(n8981), .dinb(n4994), .dout(n19209));
  jor  g18951(.dina(n8983), .dinb(n5408), .dout(n19210));
  jand g18952(.dina(n19210), .dinb(n19209), .dout(n19211));
  jand g18953(.dina(n19211), .dinb(n19208), .dout(n19212));
  jand g18954(.dina(n19212), .dinb(n19207), .dout(n19213));
  jxor g18955(.dina(n19213), .dinb(a56 ), .dout(n19214));
  jnot g18956(.din(n19214), .dout(n19215));
  jxor g18957(.dina(n19215), .dinb(n19206), .dout(n19216));
  jxor g18958(.dina(n19216), .dinb(n19169), .dout(n19217));
  jor  g18959(.dina(n8125), .dinb(n6103), .dout(n19218));
  jor  g18960(.dina(n7846), .dinb(n5428), .dout(n19219));
  jor  g18961(.dina(n8128), .dinb(n5862), .dout(n19220));
  jor  g18962(.dina(n8130), .dinb(n6106), .dout(n19221));
  jand g18963(.dina(n19221), .dinb(n19220), .dout(n19222));
  jand g18964(.dina(n19222), .dinb(n19219), .dout(n19223));
  jand g18965(.dina(n19223), .dinb(n19218), .dout(n19224));
  jxor g18966(.dina(n19224), .dinb(a53 ), .dout(n19225));
  jnot g18967(.din(n19225), .dout(n19226));
  jxor g18968(.dina(n19226), .dinb(n19217), .dout(n19227));
  jxor g18969(.dina(n19227), .dinb(n19164), .dout(n19228));
  jor  g18970(.dina(n6864), .dinb(n7266), .dout(n19229));
  jor  g18971(.dina(n7021), .dinb(n6352), .dout(n19230));
  jor  g18972(.dina(n7269), .dinb(n6372), .dout(n19231));
  jor  g18973(.dina(n7271), .dinb(n6867), .dout(n19232));
  jand g18974(.dina(n19232), .dinb(n19231), .dout(n19233));
  jand g18975(.dina(n19233), .dinb(n19230), .dout(n19234));
  jand g18976(.dina(n19234), .dinb(n19229), .dout(n19235));
  jxor g18977(.dina(n19235), .dinb(a50 ), .dout(n19236));
  jnot g18978(.din(n19236), .dout(n19237));
  jxor g18979(.dina(n19237), .dinb(n19228), .dout(n19238));
  jxor g18980(.dina(n19238), .dinb(n19159), .dout(n19239));
  jor  g18981(.dina(n7408), .dinb(n6490), .dout(n19240));
  jor  g18982(.dina(n6262), .dinb(n7129), .dout(n19241));
  jor  g18983(.dina(n6493), .dinb(n7149), .dout(n19242));
  jor  g18984(.dina(n6495), .dinb(n7411), .dout(n19243));
  jand g18985(.dina(n19243), .dinb(n19242), .dout(n19244));
  jand g18986(.dina(n19244), .dinb(n19241), .dout(n19245));
  jand g18987(.dina(n19245), .dinb(n19240), .dout(n19246));
  jxor g18988(.dina(n19246), .dinb(a47 ), .dout(n19247));
  jnot g18989(.din(n19247), .dout(n19248));
  jxor g18990(.dina(n19248), .dinb(n19239), .dout(n19249));
  jand g18991(.dina(n19068), .dinb(n19060), .dout(n19250));
  jnot g18992(.din(n19068), .dout(n19251));
  jand g18993(.dina(n19251), .dinb(n19059), .dout(n19252));
  jnot g18994(.din(n19252), .dout(n19253));
  jand g18995(.dina(n19253), .dinb(n18981), .dout(n19254));
  jor  g18996(.dina(n19254), .dinb(n19250), .dout(n19255));
  jnot g18997(.din(n19255), .dout(n19256));
  jxor g18998(.dina(n19256), .dinb(n19249), .dout(n19257));
  jxor g18999(.dina(n19257), .dinb(n19154), .dout(n19258));
  jxor g19000(.dina(n19258), .dinb(n19145), .dout(n19259));
  jor  g19001(.dina(n9387), .dinb(n5096), .dout(n19260));
  jor  g19002(.dina(n4904), .dinb(n8789), .dout(n19261));
  jor  g19003(.dina(n5099), .dinb(n8809), .dout(n19262));
  jor  g19004(.dina(n5101), .dinb(n9390), .dout(n19263));
  jand g19005(.dina(n19263), .dinb(n19262), .dout(n19264));
  jand g19006(.dina(n19264), .dinb(n19261), .dout(n19265));
  jand g19007(.dina(n19265), .dinb(n19260), .dout(n19266));
  jxor g19008(.dina(n19266), .dinb(a41 ), .dout(n19267));
  jnot g19009(.din(n19267), .dout(n19268));
  jxor g19010(.dina(n19268), .dinb(n19259), .dout(n19269));
  jxor g19011(.dina(n19269), .dinb(n19140), .dout(n19270));
  jnot g19012(.din(n19270), .dout(n19271));
  jor  g19013(.dina(n10311), .dinb(n4415), .dout(n19272));
  jor  g19014(.dina(n4272), .dinb(n9413), .dout(n19273));
  jor  g19015(.dina(n4418), .dinb(n9725), .dout(n19274));
  jor  g19016(.dina(n4420), .dinb(n10314), .dout(n19275));
  jand g19017(.dina(n19275), .dinb(n19274), .dout(n19276));
  jand g19018(.dina(n19276), .dinb(n19273), .dout(n19277));
  jand g19019(.dina(n19277), .dinb(n19272), .dout(n19278));
  jxor g19020(.dina(n19278), .dinb(a38 ), .dout(n19279));
  jxor g19021(.dina(n19279), .dinb(n19271), .dout(n19280));
  jxor g19022(.dina(n19280), .dinb(n19135), .dout(n19281));
  jxor g19023(.dina(n19281), .dinb(n19124), .dout(n19282));
  jxor g19024(.dina(n19282), .dinb(n19121), .dout(f97 ));
  jand g19025(.dina(n19281), .dinb(n19124), .dout(n19284));
  jand g19026(.dina(n19282), .dinb(n19121), .dout(n19285));
  jor  g19027(.dina(n19285), .dinb(n19284), .dout(n19286));
  jor  g19028(.dina(n19134), .dinb(n19128), .dout(n19287));
  jand g19029(.dina(n19280), .dinb(n19135), .dout(n19288));
  jnot g19030(.din(n19288), .dout(n19289));
  jand g19031(.dina(n19289), .dinb(n19287), .dout(n19290));
  jnot g19032(.din(n19290), .dout(n19291));
  jand g19033(.dina(n19269), .dinb(n19140), .dout(n19292));
  jnot g19034(.din(n19292), .dout(n19293));
  jor  g19035(.dina(n19279), .dinb(n19271), .dout(n19294));
  jand g19036(.dina(n19294), .dinb(n19293), .dout(n19295));
  jnot g19037(.din(a35 ), .dout(n19296));
  jand g19038(.dina(n11296), .dinb(n3480), .dout(n19297));
  jor  g19039(.dina(n19297), .dinb(n3690), .dout(n19298));
  jand g19040(.dina(n19298), .dinb(b63 ), .dout(n19299));
  jxor g19041(.dina(n19299), .dinb(n19296), .dout(n19300));
  jxor g19042(.dina(n19300), .dinb(n19295), .dout(n19301));
  jand g19043(.dina(n19256), .dinb(n19249), .dout(n19302));
  jand g19044(.dina(n19257), .dinb(n19154), .dout(n19303));
  jor  g19045(.dina(n19303), .dinb(n19302), .dout(n19304));
  jor  g19046(.dina(n8786), .dinb(n5739), .dout(n19305));
  jor  g19047(.dina(n5574), .dinb(n7960), .dout(n19306));
  jor  g19048(.dina(n5742), .dinb(n8231), .dout(n19307));
  jor  g19049(.dina(n5744), .dinb(n8789), .dout(n19308));
  jand g19050(.dina(n19308), .dinb(n19307), .dout(n19309));
  jand g19051(.dina(n19309), .dinb(n19306), .dout(n19310));
  jand g19052(.dina(n19310), .dinb(n19305), .dout(n19311));
  jxor g19053(.dina(n19311), .dinb(a44 ), .dout(n19312));
  jnot g19054(.din(n19312), .dout(n19313));
  jor  g19055(.dina(n7680), .dinb(n6490), .dout(n19314));
  jor  g19056(.dina(n6262), .dinb(n7149), .dout(n19315));
  jor  g19057(.dina(n6493), .dinb(n7411), .dout(n19316));
  jor  g19058(.dina(n6495), .dinb(n7683), .dout(n19317));
  jand g19059(.dina(n19317), .dinb(n19316), .dout(n19318));
  jand g19060(.dina(n19318), .dinb(n19315), .dout(n19319));
  jand g19061(.dina(n19319), .dinb(n19314), .dout(n19320));
  jxor g19062(.dina(n19320), .dinb(a47 ), .dout(n19321));
  jnot g19063(.din(n19321), .dout(n19322));
  jor  g19064(.dina(n8978), .dinb(n5425), .dout(n19323));
  jor  g19065(.dina(n8677), .dinb(n4994), .dout(n19324));
  jor  g19066(.dina(n8981), .dinb(n5408), .dout(n19325));
  jor  g19067(.dina(n8983), .dinb(n5428), .dout(n19326));
  jand g19068(.dina(n19326), .dinb(n19325), .dout(n19327));
  jand g19069(.dina(n19327), .dinb(n19324), .dout(n19328));
  jand g19070(.dina(n19328), .dinb(n19323), .dout(n19329));
  jxor g19071(.dina(n19329), .dinb(a56 ), .dout(n19330));
  jnot g19072(.din(n19330), .dout(n19331));
  jand g19073(.dina(n19203), .dinb(n19184), .dout(n19332));
  jand g19074(.dina(n19204), .dinb(n19181), .dout(n19333));
  jor  g19075(.dina(n19333), .dinb(n19332), .dout(n19334));
  jor  g19076(.dina(n9891), .dinb(n4971), .dout(n19335));
  jor  g19077(.dina(n9593), .dinb(n4537), .dout(n19336));
  jor  g19078(.dina(n9894), .dinb(n4557), .dout(n19337));
  jor  g19079(.dina(n9896), .dinb(n4974), .dout(n19338));
  jand g19080(.dina(n19338), .dinb(n19337), .dout(n19339));
  jand g19081(.dina(n19339), .dinb(n19336), .dout(n19340));
  jand g19082(.dina(n19340), .dinb(n19335), .dout(n19341));
  jxor g19083(.dina(n19341), .dinb(a59 ), .dout(n19342));
  jnot g19084(.din(n19342), .dout(n19343));
  jand g19085(.dina(n19192), .dinb(n19188), .dout(n19344));
  jnot g19086(.din(n19344), .dout(n19345));
  jor  g19087(.dina(n19202), .dinb(n19194), .dout(n19346));
  jand g19088(.dina(n19346), .dinb(n19345), .dout(n19347));
  jnot g19089(.din(n19347), .dout(n19348));
  jand g19090(.dina(n10801), .dinb(b35 ), .dout(n19349));
  jand g19091(.dina(n11107), .dinb(b34 ), .dout(n19350));
  jor  g19092(.dina(n19350), .dinb(n19349), .dout(n19351));
  jnot g19093(.din(n19351), .dout(n19352));
  jxor g19094(.dina(n19352), .dinb(n19191), .dout(n19353));
  jxor g19095(.dina(n19353), .dinb(n19348), .dout(n19354));
  jnot g19096(.din(n19354), .dout(n19355));
  jor  g19097(.dina(n10806), .dinb(n4337), .dout(n19356));
  jor  g19098(.dina(n10485), .dinb(n3942), .dout(n19357));
  jor  g19099(.dina(n10809), .dinb(n4140), .dout(n19358));
  jor  g19100(.dina(n10811), .dinb(n4340), .dout(n19359));
  jand g19101(.dina(n19359), .dinb(n19358), .dout(n19360));
  jand g19102(.dina(n19360), .dinb(n19357), .dout(n19361));
  jand g19103(.dina(n19361), .dinb(n19356), .dout(n19362));
  jxor g19104(.dina(n19362), .dinb(a62 ), .dout(n19363));
  jxor g19105(.dina(n19363), .dinb(n19355), .dout(n19364));
  jxor g19106(.dina(n19364), .dinb(n19343), .dout(n19365));
  jxor g19107(.dina(n19365), .dinb(n19334), .dout(n19366));
  jxor g19108(.dina(n19366), .dinb(n19331), .dout(n19367));
  jor  g19109(.dina(n19205), .dinb(n19172), .dout(n19368));
  jand g19110(.dina(n19205), .dinb(n19172), .dout(n19369));
  jor  g19111(.dina(n19215), .dinb(n19369), .dout(n19370));
  jand g19112(.dina(n19370), .dinb(n19368), .dout(n19371));
  jxor g19113(.dina(n19371), .dinb(n19367), .dout(n19372));
  jor  g19114(.dina(n8125), .dinb(n6349), .dout(n19373));
  jor  g19115(.dina(n7846), .dinb(n5862), .dout(n19374));
  jor  g19116(.dina(n8128), .dinb(n6106), .dout(n19375));
  jor  g19117(.dina(n8130), .dinb(n6352), .dout(n19376));
  jand g19118(.dina(n19376), .dinb(n19375), .dout(n19377));
  jand g19119(.dina(n19377), .dinb(n19374), .dout(n19378));
  jand g19120(.dina(n19378), .dinb(n19373), .dout(n19379));
  jxor g19121(.dina(n19379), .dinb(a53 ), .dout(n19380));
  jnot g19122(.din(n19380), .dout(n19381));
  jxor g19123(.dina(n19381), .dinb(n19372), .dout(n19382));
  jnot g19124(.din(n19216), .dout(n19383));
  jand g19125(.dina(n19383), .dinb(n19168), .dout(n19384));
  jnot g19126(.din(n19384), .dout(n19385));
  jand g19127(.dina(n19216), .dinb(n19169), .dout(n19386));
  jor  g19128(.dina(n19226), .dinb(n19386), .dout(n19387));
  jand g19129(.dina(n19387), .dinb(n19385), .dout(n19388));
  jxor g19130(.dina(n19388), .dinb(n19382), .dout(n19389));
  jnot g19131(.din(n19389), .dout(n19390));
  jor  g19132(.dina(n7126), .dinb(n7266), .dout(n19391));
  jor  g19133(.dina(n7021), .dinb(n6372), .dout(n19392));
  jor  g19134(.dina(n7269), .dinb(n6867), .dout(n19393));
  jor  g19135(.dina(n7271), .dinb(n7129), .dout(n19394));
  jand g19136(.dina(n19394), .dinb(n19393), .dout(n19395));
  jand g19137(.dina(n19395), .dinb(n19392), .dout(n19396));
  jand g19138(.dina(n19396), .dinb(n19391), .dout(n19397));
  jxor g19139(.dina(n19397), .dinb(a50 ), .dout(n19398));
  jxor g19140(.dina(n19398), .dinb(n19390), .dout(n19399));
  jnot g19141(.din(n19227), .dout(n19400));
  jand g19142(.dina(n19400), .dinb(n19163), .dout(n19401));
  jnot g19143(.din(n19401), .dout(n19402));
  jand g19144(.dina(n19227), .dinb(n19164), .dout(n19403));
  jor  g19145(.dina(n19237), .dinb(n19403), .dout(n19404));
  jand g19146(.dina(n19404), .dinb(n19402), .dout(n19405));
  jxor g19147(.dina(n19405), .dinb(n19399), .dout(n19406));
  jxor g19148(.dina(n19406), .dinb(n19322), .dout(n19407));
  jnot g19149(.din(n19238), .dout(n19408));
  jand g19150(.dina(n19408), .dinb(n19158), .dout(n19409));
  jnot g19151(.din(n19409), .dout(n19410));
  jand g19152(.dina(n19238), .dinb(n19159), .dout(n19411));
  jor  g19153(.dina(n19248), .dinb(n19411), .dout(n19412));
  jand g19154(.dina(n19412), .dinb(n19410), .dout(n19413));
  jxor g19155(.dina(n19413), .dinb(n19407), .dout(n19414));
  jxor g19156(.dina(n19414), .dinb(n19313), .dout(n19415));
  jxor g19157(.dina(n19415), .dinb(n19304), .dout(n19416));
  jor  g19158(.dina(n9410), .dinb(n5096), .dout(n19417));
  jor  g19159(.dina(n4904), .dinb(n8809), .dout(n19418));
  jor  g19160(.dina(n5099), .dinb(n9390), .dout(n19419));
  jor  g19161(.dina(n5101), .dinb(n9413), .dout(n19420));
  jand g19162(.dina(n19420), .dinb(n19419), .dout(n19421));
  jand g19163(.dina(n19421), .dinb(n19418), .dout(n19422));
  jand g19164(.dina(n19422), .dinb(n19417), .dout(n19423));
  jxor g19165(.dina(n19423), .dinb(a41 ), .dout(n19424));
  jnot g19166(.din(n19424), .dout(n19425));
  jxor g19167(.dina(n19425), .dinb(n19416), .dout(n19426));
  jor  g19168(.dina(n19258), .dinb(n19145), .dout(n19427));
  jand g19169(.dina(n19258), .dinb(n19145), .dout(n19428));
  jor  g19170(.dina(n19268), .dinb(n19428), .dout(n19429));
  jand g19171(.dina(n19429), .dinb(n19427), .dout(n19430));
  jxor g19172(.dina(n19430), .dinb(n19426), .dout(n19431));
  jor  g19173(.dina(n10634), .dinb(n4415), .dout(n19432));
  jor  g19174(.dina(n4272), .dinb(n9725), .dout(n19433));
  jor  g19175(.dina(n4418), .dinb(n10314), .dout(n19434));
  jor  g19176(.dina(n4420), .dinb(n10637), .dout(n19435));
  jand g19177(.dina(n19435), .dinb(n19434), .dout(n19436));
  jand g19178(.dina(n19436), .dinb(n19433), .dout(n19437));
  jand g19179(.dina(n19437), .dinb(n19432), .dout(n19438));
  jxor g19180(.dina(n19438), .dinb(a38 ), .dout(n19439));
  jnot g19181(.din(n19439), .dout(n19440));
  jxor g19182(.dina(n19440), .dinb(n19431), .dout(n19441));
  jxor g19183(.dina(n19441), .dinb(n19301), .dout(n19442));
  jxor g19184(.dina(n19442), .dinb(n19291), .dout(n19443));
  jxor g19185(.dina(n19443), .dinb(n19286), .dout(f98 ));
  jand g19186(.dina(n19442), .dinb(n19291), .dout(n19445));
  jand g19187(.dina(n19443), .dinb(n19286), .dout(n19446));
  jor  g19188(.dina(n19446), .dinb(n19445), .dout(n19447));
  jand g19189(.dina(n19413), .dinb(n19407), .dout(n19448));
  jand g19190(.dina(n19414), .dinb(n19313), .dout(n19449));
  jor  g19191(.dina(n19449), .dinb(n19448), .dout(n19450));
  jand g19192(.dina(n19405), .dinb(n19399), .dout(n19451));
  jand g19193(.dina(n19406), .dinb(n19322), .dout(n19452));
  jor  g19194(.dina(n19452), .dinb(n19451), .dout(n19453));
  jor  g19195(.dina(n7957), .dinb(n6490), .dout(n19454));
  jor  g19196(.dina(n6262), .dinb(n7411), .dout(n19455));
  jor  g19197(.dina(n6493), .dinb(n7683), .dout(n19456));
  jor  g19198(.dina(n6495), .dinb(n7960), .dout(n19457));
  jand g19199(.dina(n19457), .dinb(n19456), .dout(n19458));
  jand g19200(.dina(n19458), .dinb(n19455), .dout(n19459));
  jand g19201(.dina(n19459), .dinb(n19454), .dout(n19460));
  jxor g19202(.dina(n19460), .dinb(a47 ), .dout(n19461));
  jnot g19203(.din(n19461), .dout(n19462));
  jand g19204(.dina(n19388), .dinb(n19382), .dout(n19463));
  jnot g19205(.din(n19463), .dout(n19464));
  jor  g19206(.dina(n19398), .dinb(n19390), .dout(n19465));
  jand g19207(.dina(n19465), .dinb(n19464), .dout(n19466));
  jnot g19208(.din(n19466), .dout(n19467));
  jand g19209(.dina(n19365), .dinb(n19334), .dout(n19468));
  jand g19210(.dina(n19366), .dinb(n19331), .dout(n19469));
  jor  g19211(.dina(n19469), .dinb(n19468), .dout(n19470));
  jor  g19212(.dina(n8978), .dinb(n5859), .dout(n19471));
  jor  g19213(.dina(n8677), .dinb(n5408), .dout(n19472));
  jor  g19214(.dina(n8981), .dinb(n5428), .dout(n19473));
  jor  g19215(.dina(n8983), .dinb(n5862), .dout(n19474));
  jand g19216(.dina(n19474), .dinb(n19473), .dout(n19475));
  jand g19217(.dina(n19475), .dinb(n19472), .dout(n19476));
  jand g19218(.dina(n19476), .dinb(n19471), .dout(n19477));
  jxor g19219(.dina(n19477), .dinb(a56 ), .dout(n19478));
  jnot g19220(.din(n19478), .dout(n19479));
  jor  g19221(.dina(n19363), .dinb(n19355), .dout(n19480));
  jand g19222(.dina(n19364), .dinb(n19343), .dout(n19481));
  jnot g19223(.din(n19481), .dout(n19482));
  jand g19224(.dina(n19482), .dinb(n19480), .dout(n19483));
  jnot g19225(.din(n19483), .dout(n19484));
  jand g19226(.dina(n19352), .dinb(n19191), .dout(n19485));
  jand g19227(.dina(n19353), .dinb(n19348), .dout(n19486));
  jor  g19228(.dina(n19486), .dinb(n19485), .dout(n19487));
  jxor g19229(.dina(n19351), .dinb(n19296), .dout(n19488));
  jand g19230(.dina(n10801), .dinb(b36 ), .dout(n19489));
  jand g19231(.dina(n11107), .dinb(b35 ), .dout(n19490));
  jor  g19232(.dina(n19490), .dinb(n19489), .dout(n19491));
  jxor g19233(.dina(n19491), .dinb(n19488), .dout(n19492));
  jxor g19234(.dina(n19492), .dinb(n19487), .dout(n19493));
  jnot g19235(.din(n19493), .dout(n19494));
  jor  g19236(.dina(n10806), .dinb(n4534), .dout(n19495));
  jor  g19237(.dina(n10485), .dinb(n4140), .dout(n19496));
  jor  g19238(.dina(n10809), .dinb(n4340), .dout(n19497));
  jor  g19239(.dina(n10811), .dinb(n4537), .dout(n19498));
  jand g19240(.dina(n19498), .dinb(n19497), .dout(n19499));
  jand g19241(.dina(n19499), .dinb(n19496), .dout(n19500));
  jand g19242(.dina(n19500), .dinb(n19495), .dout(n19501));
  jxor g19243(.dina(n19501), .dinb(a62 ), .dout(n19502));
  jxor g19244(.dina(n19502), .dinb(n19494), .dout(n19503));
  jnot g19245(.din(n19503), .dout(n19504));
  jor  g19246(.dina(n9891), .dinb(n4991), .dout(n19505));
  jor  g19247(.dina(n9593), .dinb(n4557), .dout(n19506));
  jor  g19248(.dina(n9894), .dinb(n4974), .dout(n19507));
  jor  g19249(.dina(n9896), .dinb(n4994), .dout(n19508));
  jand g19250(.dina(n19508), .dinb(n19507), .dout(n19509));
  jand g19251(.dina(n19509), .dinb(n19506), .dout(n19510));
  jand g19252(.dina(n19510), .dinb(n19505), .dout(n19511));
  jxor g19253(.dina(n19511), .dinb(a59 ), .dout(n19512));
  jxor g19254(.dina(n19512), .dinb(n19504), .dout(n19513));
  jxor g19255(.dina(n19513), .dinb(n19484), .dout(n19514));
  jxor g19256(.dina(n19514), .dinb(n19479), .dout(n19515));
  jxor g19257(.dina(n19515), .dinb(n19470), .dout(n19516));
  jnot g19258(.din(n19516), .dout(n19517));
  jor  g19259(.dina(n8125), .dinb(n6369), .dout(n19518));
  jor  g19260(.dina(n7846), .dinb(n6106), .dout(n19519));
  jor  g19261(.dina(n8128), .dinb(n6352), .dout(n19520));
  jor  g19262(.dina(n8130), .dinb(n6372), .dout(n19521));
  jand g19263(.dina(n19521), .dinb(n19520), .dout(n19522));
  jand g19264(.dina(n19522), .dinb(n19519), .dout(n19523));
  jand g19265(.dina(n19523), .dinb(n19518), .dout(n19524));
  jxor g19266(.dina(n19524), .dinb(a53 ), .dout(n19525));
  jxor g19267(.dina(n19525), .dinb(n19517), .dout(n19526));
  jor  g19268(.dina(n19371), .dinb(n19367), .dout(n19527));
  jand g19269(.dina(n19371), .dinb(n19367), .dout(n19528));
  jor  g19270(.dina(n19381), .dinb(n19528), .dout(n19529));
  jand g19271(.dina(n19529), .dinb(n19527), .dout(n19530));
  jxor g19272(.dina(n19530), .dinb(n19526), .dout(n19531));
  jnot g19273(.din(n19531), .dout(n19532));
  jor  g19274(.dina(n7146), .dinb(n7266), .dout(n19533));
  jor  g19275(.dina(n7021), .dinb(n6867), .dout(n19534));
  jor  g19276(.dina(n7269), .dinb(n7129), .dout(n19535));
  jor  g19277(.dina(n7271), .dinb(n7149), .dout(n19536));
  jand g19278(.dina(n19536), .dinb(n19535), .dout(n19537));
  jand g19279(.dina(n19537), .dinb(n19534), .dout(n19538));
  jand g19280(.dina(n19538), .dinb(n19533), .dout(n19539));
  jxor g19281(.dina(n19539), .dinb(a50 ), .dout(n19540));
  jxor g19282(.dina(n19540), .dinb(n19532), .dout(n19541));
  jxor g19283(.dina(n19541), .dinb(n19467), .dout(n19542));
  jxor g19284(.dina(n19542), .dinb(n19462), .dout(n19543));
  jxor g19285(.dina(n19543), .dinb(n19453), .dout(n19544));
  jnot g19286(.din(n19544), .dout(n19545));
  jor  g19287(.dina(n8806), .dinb(n5739), .dout(n19546));
  jor  g19288(.dina(n5574), .dinb(n8231), .dout(n19547));
  jor  g19289(.dina(n5742), .dinb(n8789), .dout(n19548));
  jor  g19290(.dina(n5744), .dinb(n8809), .dout(n19549));
  jand g19291(.dina(n19549), .dinb(n19548), .dout(n19550));
  jand g19292(.dina(n19550), .dinb(n19547), .dout(n19551));
  jand g19293(.dina(n19551), .dinb(n19546), .dout(n19552));
  jxor g19294(.dina(n19552), .dinb(a44 ), .dout(n19553));
  jxor g19295(.dina(n19553), .dinb(n19545), .dout(n19554));
  jxor g19296(.dina(n19554), .dinb(n19450), .dout(n19555));
  jnot g19297(.din(n19555), .dout(n19556));
  jor  g19298(.dina(n9722), .dinb(n5096), .dout(n19557));
  jor  g19299(.dina(n4904), .dinb(n9390), .dout(n19558));
  jor  g19300(.dina(n5099), .dinb(n9413), .dout(n19559));
  jor  g19301(.dina(n5101), .dinb(n9725), .dout(n19560));
  jand g19302(.dina(n19560), .dinb(n19559), .dout(n19561));
  jand g19303(.dina(n19561), .dinb(n19558), .dout(n19562));
  jand g19304(.dina(n19562), .dinb(n19557), .dout(n19563));
  jxor g19305(.dina(n19563), .dinb(a41 ), .dout(n19564));
  jxor g19306(.dina(n19564), .dinb(n19556), .dout(n19565));
  jor  g19307(.dina(n19415), .dinb(n19304), .dout(n19566));
  jand g19308(.dina(n19415), .dinb(n19304), .dout(n19567));
  jor  g19309(.dina(n19425), .dinb(n19567), .dout(n19568));
  jand g19310(.dina(n19568), .dinb(n19566), .dout(n19569));
  jxor g19311(.dina(n19569), .dinb(n19565), .dout(n19570));
  jnot g19312(.din(n19570), .dout(n19571));
  jor  g19313(.dina(n10961), .dinb(n4415), .dout(n19572));
  jor  g19314(.dina(n4272), .dinb(n10314), .dout(n19573));
  jor  g19315(.dina(n4418), .dinb(n10637), .dout(n19574));
  jor  g19316(.dina(n4420), .dinb(n10964), .dout(n19575));
  jand g19317(.dina(n19575), .dinb(n19574), .dout(n19576));
  jand g19318(.dina(n19576), .dinb(n19573), .dout(n19577));
  jand g19319(.dina(n19577), .dinb(n19572), .dout(n19578));
  jxor g19320(.dina(n19578), .dinb(a38 ), .dout(n19579));
  jxor g19321(.dina(n19579), .dinb(n19571), .dout(n19580));
  jnot g19322(.din(n19426), .dout(n19581));
  jnot g19323(.din(n19430), .dout(n19582));
  jand g19324(.dina(n19582), .dinb(n19581), .dout(n19583));
  jnot g19325(.din(n19583), .dout(n19584));
  jand g19326(.dina(n19430), .dinb(n19426), .dout(n19585));
  jor  g19327(.dina(n19440), .dinb(n19585), .dout(n19586));
  jand g19328(.dina(n19586), .dinb(n19584), .dout(n19587));
  jxor g19329(.dina(n19587), .dinb(n19580), .dout(n19588));
  jnot g19330(.din(n19588), .dout(n19589));
  jor  g19331(.dina(n19300), .dinb(n19295), .dout(n19590));
  jand g19332(.dina(n19441), .dinb(n19301), .dout(n19591));
  jnot g19333(.din(n19591), .dout(n19592));
  jand g19334(.dina(n19592), .dinb(n19590), .dout(n19593));
  jxor g19335(.dina(n19593), .dinb(n19589), .dout(n19594));
  jxor g19336(.dina(n19594), .dinb(n19447), .dout(f99 ));
  jor  g19337(.dina(n19579), .dinb(n19571), .dout(n19596));
  jand g19338(.dina(n19587), .dinb(n19580), .dout(n19597));
  jnot g19339(.din(n19597), .dout(n19598));
  jand g19340(.dina(n19598), .dinb(n19596), .dout(n19599));
  jnot g19341(.din(n19599), .dout(n19600));
  jor  g19342(.dina(n19564), .dinb(n19556), .dout(n19601));
  jand g19343(.dina(n19569), .dinb(n19565), .dout(n19602));
  jnot g19344(.din(n19602), .dout(n19603));
  jand g19345(.dina(n19603), .dinb(n19601), .dout(n19604));
  jor  g19346(.dina(n10978), .dinb(n4415), .dout(n19605));
  jor  g19347(.dina(n4272), .dinb(n10637), .dout(n19606));
  jor  g19348(.dina(n4418), .dinb(n10964), .dout(n19607));
  jand g19349(.dina(n19607), .dinb(n19606), .dout(n19608));
  jand g19350(.dina(n19608), .dinb(n19605), .dout(n19609));
  jxor g19351(.dina(n19609), .dinb(a38 ), .dout(n19610));
  jxor g19352(.dina(n19610), .dinb(n19604), .dout(n19611));
  jor  g19353(.dina(n19553), .dinb(n19545), .dout(n19612));
  jand g19354(.dina(n19554), .dinb(n19450), .dout(n19613));
  jnot g19355(.din(n19613), .dout(n19614));
  jand g19356(.dina(n19614), .dinb(n19612), .dout(n19615));
  jnot g19357(.din(n19615), .dout(n19616));
  jand g19358(.dina(n19542), .dinb(n19462), .dout(n19617));
  jand g19359(.dina(n19543), .dinb(n19453), .dout(n19618));
  jor  g19360(.dina(n19618), .dinb(n19617), .dout(n19619));
  jor  g19361(.dina(n8228), .dinb(n6490), .dout(n19620));
  jor  g19362(.dina(n6262), .dinb(n7683), .dout(n19621));
  jor  g19363(.dina(n6493), .dinb(n7960), .dout(n19622));
  jor  g19364(.dina(n6495), .dinb(n8231), .dout(n19623));
  jand g19365(.dina(n19623), .dinb(n19622), .dout(n19624));
  jand g19366(.dina(n19624), .dinb(n19621), .dout(n19625));
  jand g19367(.dina(n19625), .dinb(n19620), .dout(n19626));
  jxor g19368(.dina(n19626), .dinb(a47 ), .dout(n19627));
  jnot g19369(.din(n19627), .dout(n19628));
  jor  g19370(.dina(n19540), .dinb(n19532), .dout(n19629));
  jand g19371(.dina(n19541), .dinb(n19467), .dout(n19630));
  jnot g19372(.din(n19630), .dout(n19631));
  jand g19373(.dina(n19631), .dinb(n19629), .dout(n19632));
  jnot g19374(.din(n19632), .dout(n19633));
  jor  g19375(.dina(n19525), .dinb(n19517), .dout(n19634));
  jand g19376(.dina(n19530), .dinb(n19526), .dout(n19635));
  jnot g19377(.din(n19635), .dout(n19636));
  jand g19378(.dina(n19636), .dinb(n19634), .dout(n19637));
  jnot g19379(.din(n19637), .dout(n19638));
  jand g19380(.dina(n19514), .dinb(n19479), .dout(n19639));
  jand g19381(.dina(n19515), .dinb(n19470), .dout(n19640));
  jor  g19382(.dina(n19640), .dinb(n19639), .dout(n19641));
  jor  g19383(.dina(n19512), .dinb(n19504), .dout(n19642));
  jand g19384(.dina(n19513), .dinb(n19484), .dout(n19643));
  jnot g19385(.din(n19643), .dout(n19644));
  jand g19386(.dina(n19644), .dinb(n19642), .dout(n19645));
  jand g19387(.dina(n19492), .dinb(n19487), .dout(n19646));
  jnot g19388(.din(n19646), .dout(n19647));
  jor  g19389(.dina(n19502), .dinb(n19494), .dout(n19648));
  jand g19390(.dina(n19648), .dinb(n19647), .dout(n19649));
  jor  g19391(.dina(n10806), .dinb(n4554), .dout(n19650));
  jor  g19392(.dina(n10485), .dinb(n4340), .dout(n19651));
  jor  g19393(.dina(n10809), .dinb(n4537), .dout(n19652));
  jor  g19394(.dina(n10811), .dinb(n4557), .dout(n19653));
  jand g19395(.dina(n19653), .dinb(n19652), .dout(n19654));
  jand g19396(.dina(n19654), .dinb(n19651), .dout(n19655));
  jand g19397(.dina(n19655), .dinb(n19650), .dout(n19656));
  jxor g19398(.dina(n19656), .dinb(a62 ), .dout(n19657));
  jnot g19399(.din(n19657), .dout(n19658));
  jand g19400(.dina(n19351), .dinb(n19296), .dout(n19659));
  jand g19401(.dina(n19491), .dinb(n19488), .dout(n19660));
  jor  g19402(.dina(n19660), .dinb(n19659), .dout(n19661));
  jand g19403(.dina(n10801), .dinb(b37 ), .dout(n19662));
  jand g19404(.dina(n11107), .dinb(b36 ), .dout(n19663));
  jor  g19405(.dina(n19663), .dinb(n19662), .dout(n19664));
  jnot g19406(.din(n19664), .dout(n19665));
  jxor g19407(.dina(n19665), .dinb(n19661), .dout(n19666));
  jxor g19408(.dina(n19666), .dinb(n19658), .dout(n19667));
  jnot g19409(.din(n19667), .dout(n19668));
  jxor g19410(.dina(n19668), .dinb(n19649), .dout(n19669));
  jor  g19411(.dina(n9891), .dinb(n5405), .dout(n19670));
  jor  g19412(.dina(n9593), .dinb(n4974), .dout(n19671));
  jor  g19413(.dina(n9894), .dinb(n4994), .dout(n19672));
  jor  g19414(.dina(n9896), .dinb(n5408), .dout(n19673));
  jand g19415(.dina(n19673), .dinb(n19672), .dout(n19674));
  jand g19416(.dina(n19674), .dinb(n19671), .dout(n19675));
  jand g19417(.dina(n19675), .dinb(n19670), .dout(n19676));
  jxor g19418(.dina(n19676), .dinb(a59 ), .dout(n19677));
  jnot g19419(.din(n19677), .dout(n19678));
  jxor g19420(.dina(n19678), .dinb(n19669), .dout(n19679));
  jnot g19421(.din(n19679), .dout(n19680));
  jxor g19422(.dina(n19680), .dinb(n19645), .dout(n19681));
  jor  g19423(.dina(n8978), .dinb(n6103), .dout(n19682));
  jor  g19424(.dina(n8677), .dinb(n5428), .dout(n19683));
  jor  g19425(.dina(n8981), .dinb(n5862), .dout(n19684));
  jor  g19426(.dina(n8983), .dinb(n6106), .dout(n19685));
  jand g19427(.dina(n19685), .dinb(n19684), .dout(n19686));
  jand g19428(.dina(n19686), .dinb(n19683), .dout(n19687));
  jand g19429(.dina(n19687), .dinb(n19682), .dout(n19688));
  jxor g19430(.dina(n19688), .dinb(a56 ), .dout(n19689));
  jnot g19431(.din(n19689), .dout(n19690));
  jxor g19432(.dina(n19690), .dinb(n19681), .dout(n19691));
  jxor g19433(.dina(n19691), .dinb(n19641), .dout(n19692));
  jor  g19434(.dina(n8125), .dinb(n6864), .dout(n19693));
  jor  g19435(.dina(n7846), .dinb(n6352), .dout(n19694));
  jor  g19436(.dina(n8128), .dinb(n6372), .dout(n19695));
  jor  g19437(.dina(n8130), .dinb(n6867), .dout(n19696));
  jand g19438(.dina(n19696), .dinb(n19695), .dout(n19697));
  jand g19439(.dina(n19697), .dinb(n19694), .dout(n19698));
  jand g19440(.dina(n19698), .dinb(n19693), .dout(n19699));
  jxor g19441(.dina(n19699), .dinb(a53 ), .dout(n19700));
  jnot g19442(.din(n19700), .dout(n19701));
  jxor g19443(.dina(n19701), .dinb(n19692), .dout(n19702));
  jxor g19444(.dina(n19702), .dinb(n19638), .dout(n19703));
  jor  g19445(.dina(n7408), .dinb(n7266), .dout(n19704));
  jor  g19446(.dina(n7021), .dinb(n7129), .dout(n19705));
  jor  g19447(.dina(n7269), .dinb(n7149), .dout(n19706));
  jor  g19448(.dina(n7271), .dinb(n7411), .dout(n19707));
  jand g19449(.dina(n19707), .dinb(n19706), .dout(n19708));
  jand g19450(.dina(n19708), .dinb(n19705), .dout(n19709));
  jand g19451(.dina(n19709), .dinb(n19704), .dout(n19710));
  jxor g19452(.dina(n19710), .dinb(a50 ), .dout(n19711));
  jnot g19453(.din(n19711), .dout(n19712));
  jxor g19454(.dina(n19712), .dinb(n19703), .dout(n19713));
  jxor g19455(.dina(n19713), .dinb(n19633), .dout(n19714));
  jxor g19456(.dina(n19714), .dinb(n19628), .dout(n19715));
  jxor g19457(.dina(n19715), .dinb(n19619), .dout(n19716));
  jor  g19458(.dina(n9387), .dinb(n5739), .dout(n19717));
  jor  g19459(.dina(n5574), .dinb(n8789), .dout(n19718));
  jor  g19460(.dina(n5742), .dinb(n8809), .dout(n19719));
  jor  g19461(.dina(n5744), .dinb(n9390), .dout(n19720));
  jand g19462(.dina(n19720), .dinb(n19719), .dout(n19721));
  jand g19463(.dina(n19721), .dinb(n19718), .dout(n19722));
  jand g19464(.dina(n19722), .dinb(n19717), .dout(n19723));
  jxor g19465(.dina(n19723), .dinb(a44 ), .dout(n19724));
  jnot g19466(.din(n19724), .dout(n19725));
  jxor g19467(.dina(n19725), .dinb(n19716), .dout(n19726));
  jxor g19468(.dina(n19726), .dinb(n19616), .dout(n19727));
  jnot g19469(.din(n19727), .dout(n19728));
  jor  g19470(.dina(n10311), .dinb(n5096), .dout(n19729));
  jor  g19471(.dina(n4904), .dinb(n9413), .dout(n19730));
  jor  g19472(.dina(n5099), .dinb(n9725), .dout(n19731));
  jor  g19473(.dina(n5101), .dinb(n10314), .dout(n19732));
  jand g19474(.dina(n19732), .dinb(n19731), .dout(n19733));
  jand g19475(.dina(n19733), .dinb(n19730), .dout(n19734));
  jand g19476(.dina(n19734), .dinb(n19729), .dout(n19735));
  jxor g19477(.dina(n19735), .dinb(a41 ), .dout(n19736));
  jxor g19478(.dina(n19736), .dinb(n19728), .dout(n19737));
  jxor g19479(.dina(n19737), .dinb(n19611), .dout(n19738));
  jxor g19480(.dina(n19738), .dinb(n19600), .dout(n19739));
  jor  g19481(.dina(n19593), .dinb(n19589), .dout(n19740));
  jnot g19482(.din(n19740), .dout(n19741));
  jand g19483(.dina(n19594), .dinb(n19447), .dout(n19742));
  jor  g19484(.dina(n19742), .dinb(n19741), .dout(n19743));
  jxor g19485(.dina(n19743), .dinb(n19739), .dout(f100 ));
  jand g19486(.dina(n19738), .dinb(n19600), .dout(n19745));
  jand g19487(.dina(n19743), .dinb(n19739), .dout(n19746));
  jor  g19488(.dina(n19746), .dinb(n19745), .dout(n19747));
  jor  g19489(.dina(n19610), .dinb(n19604), .dout(n19748));
  jand g19490(.dina(n19737), .dinb(n19611), .dout(n19749));
  jnot g19491(.din(n19749), .dout(n19750));
  jand g19492(.dina(n19750), .dinb(n19748), .dout(n19751));
  jnot g19493(.din(n19751), .dout(n19752));
  jand g19494(.dina(n19726), .dinb(n19616), .dout(n19753));
  jnot g19495(.din(n19753), .dout(n19754));
  jor  g19496(.dina(n19736), .dinb(n19728), .dout(n19755));
  jand g19497(.dina(n19755), .dinb(n19754), .dout(n19756));
  jnot g19498(.din(a38 ), .dout(n19757));
  jand g19499(.dina(n11296), .dinb(n4059), .dout(n19758));
  jor  g19500(.dina(n19758), .dinb(n4273), .dout(n19759));
  jand g19501(.dina(n19759), .dinb(b63 ), .dout(n19760));
  jxor g19502(.dina(n19760), .dinb(n19757), .dout(n19761));
  jxor g19503(.dina(n19761), .dinb(n19756), .dout(n19762));
  jand g19504(.dina(n19713), .dinb(n19633), .dout(n19763));
  jand g19505(.dina(n19714), .dinb(n19628), .dout(n19764));
  jor  g19506(.dina(n19764), .dinb(n19763), .dout(n19765));
  jor  g19507(.dina(n8786), .dinb(n6490), .dout(n19766));
  jor  g19508(.dina(n6262), .dinb(n7960), .dout(n19767));
  jor  g19509(.dina(n6493), .dinb(n8231), .dout(n19768));
  jor  g19510(.dina(n6495), .dinb(n8789), .dout(n19769));
  jand g19511(.dina(n19769), .dinb(n19768), .dout(n19770));
  jand g19512(.dina(n19770), .dinb(n19767), .dout(n19771));
  jand g19513(.dina(n19771), .dinb(n19766), .dout(n19772));
  jxor g19514(.dina(n19772), .dinb(a47 ), .dout(n19773));
  jnot g19515(.din(n19773), .dout(n19774));
  jor  g19516(.dina(n7680), .dinb(n7266), .dout(n19775));
  jor  g19517(.dina(n7021), .dinb(n7149), .dout(n19776));
  jor  g19518(.dina(n7269), .dinb(n7411), .dout(n19777));
  jor  g19519(.dina(n7271), .dinb(n7683), .dout(n19778));
  jand g19520(.dina(n19778), .dinb(n19777), .dout(n19779));
  jand g19521(.dina(n19779), .dinb(n19776), .dout(n19780));
  jand g19522(.dina(n19780), .dinb(n19775), .dout(n19781));
  jxor g19523(.dina(n19781), .dinb(a50 ), .dout(n19782));
  jnot g19524(.din(n19782), .dout(n19783));
  jor  g19525(.dina(n9891), .dinb(n5425), .dout(n19784));
  jor  g19526(.dina(n9593), .dinb(n4994), .dout(n19785));
  jor  g19527(.dina(n9894), .dinb(n5408), .dout(n19786));
  jor  g19528(.dina(n9896), .dinb(n5428), .dout(n19787));
  jand g19529(.dina(n19787), .dinb(n19786), .dout(n19788));
  jand g19530(.dina(n19788), .dinb(n19785), .dout(n19789));
  jand g19531(.dina(n19789), .dinb(n19784), .dout(n19790));
  jxor g19532(.dina(n19790), .dinb(a59 ), .dout(n19791));
  jnot g19533(.din(n19791), .dout(n19792));
  jor  g19534(.dina(n10806), .dinb(n4971), .dout(n19793));
  jor  g19535(.dina(n10485), .dinb(n4537), .dout(n19794));
  jor  g19536(.dina(n10809), .dinb(n4557), .dout(n19795));
  jor  g19537(.dina(n10811), .dinb(n4974), .dout(n19796));
  jand g19538(.dina(n19796), .dinb(n19795), .dout(n19797));
  jand g19539(.dina(n19797), .dinb(n19794), .dout(n19798));
  jand g19540(.dina(n19798), .dinb(n19793), .dout(n19799));
  jxor g19541(.dina(n19799), .dinb(a62 ), .dout(n19800));
  jnot g19542(.din(n19800), .dout(n19801));
  jand g19543(.dina(n10801), .dinb(b38 ), .dout(n19802));
  jand g19544(.dina(n11107), .dinb(b37 ), .dout(n19803));
  jor  g19545(.dina(n19803), .dinb(n19802), .dout(n19804));
  jxor g19546(.dina(n19804), .dinb(n19665), .dout(n19805));
  jor  g19547(.dina(n19665), .dinb(n19661), .dout(n19806));
  jand g19548(.dina(n19665), .dinb(n19661), .dout(n19807));
  jor  g19549(.dina(n19807), .dinb(n19658), .dout(n19808));
  jand g19550(.dina(n19808), .dinb(n19806), .dout(n19809));
  jxor g19551(.dina(n19809), .dinb(n19805), .dout(n19810));
  jxor g19552(.dina(n19810), .dinb(n19801), .dout(n19811));
  jxor g19553(.dina(n19811), .dinb(n19792), .dout(n19812));
  jand g19554(.dina(n19668), .dinb(n19649), .dout(n19813));
  jnot g19555(.din(n19813), .dout(n19814));
  jnot g19556(.din(n19649), .dout(n19815));
  jand g19557(.dina(n19667), .dinb(n19815), .dout(n19816));
  jor  g19558(.dina(n19678), .dinb(n19816), .dout(n19817));
  jand g19559(.dina(n19817), .dinb(n19814), .dout(n19818));
  jxor g19560(.dina(n19818), .dinb(n19812), .dout(n19819));
  jor  g19561(.dina(n8978), .dinb(n6349), .dout(n19820));
  jor  g19562(.dina(n8677), .dinb(n5862), .dout(n19821));
  jor  g19563(.dina(n8981), .dinb(n6106), .dout(n19822));
  jor  g19564(.dina(n8983), .dinb(n6352), .dout(n19823));
  jand g19565(.dina(n19823), .dinb(n19822), .dout(n19824));
  jand g19566(.dina(n19824), .dinb(n19821), .dout(n19825));
  jand g19567(.dina(n19825), .dinb(n19820), .dout(n19826));
  jxor g19568(.dina(n19826), .dinb(a56 ), .dout(n19827));
  jnot g19569(.din(n19827), .dout(n19828));
  jxor g19570(.dina(n19828), .dinb(n19819), .dout(n19829));
  jand g19571(.dina(n19680), .dinb(n19645), .dout(n19830));
  jnot g19572(.din(n19830), .dout(n19831));
  jnot g19573(.din(n19645), .dout(n19832));
  jand g19574(.dina(n19679), .dinb(n19832), .dout(n19833));
  jor  g19575(.dina(n19690), .dinb(n19833), .dout(n19834));
  jand g19576(.dina(n19834), .dinb(n19831), .dout(n19835));
  jxor g19577(.dina(n19835), .dinb(n19829), .dout(n19836));
  jnot g19578(.din(n19836), .dout(n19837));
  jor  g19579(.dina(n8125), .dinb(n7126), .dout(n19838));
  jor  g19580(.dina(n7846), .dinb(n6372), .dout(n19839));
  jor  g19581(.dina(n8128), .dinb(n6867), .dout(n19840));
  jor  g19582(.dina(n8130), .dinb(n7129), .dout(n19841));
  jand g19583(.dina(n19841), .dinb(n19840), .dout(n19842));
  jand g19584(.dina(n19842), .dinb(n19839), .dout(n19843));
  jand g19585(.dina(n19843), .dinb(n19838), .dout(n19844));
  jxor g19586(.dina(n19844), .dinb(a53 ), .dout(n19845));
  jxor g19587(.dina(n19845), .dinb(n19837), .dout(n19846));
  jnot g19588(.din(n19641), .dout(n19847));
  jnot g19589(.din(n19691), .dout(n19848));
  jand g19590(.dina(n19848), .dinb(n19847), .dout(n19849));
  jnot g19591(.din(n19849), .dout(n19850));
  jand g19592(.dina(n19691), .dinb(n19641), .dout(n19851));
  jor  g19593(.dina(n19701), .dinb(n19851), .dout(n19852));
  jand g19594(.dina(n19852), .dinb(n19850), .dout(n19853));
  jxor g19595(.dina(n19853), .dinb(n19846), .dout(n19854));
  jxor g19596(.dina(n19854), .dinb(n19783), .dout(n19855));
  jnot g19597(.din(n19702), .dout(n19856));
  jand g19598(.dina(n19856), .dinb(n19637), .dout(n19857));
  jnot g19599(.din(n19857), .dout(n19858));
  jand g19600(.dina(n19702), .dinb(n19638), .dout(n19859));
  jor  g19601(.dina(n19712), .dinb(n19859), .dout(n19860));
  jand g19602(.dina(n19860), .dinb(n19858), .dout(n19861));
  jxor g19603(.dina(n19861), .dinb(n19855), .dout(n19862));
  jxor g19604(.dina(n19862), .dinb(n19774), .dout(n19863));
  jxor g19605(.dina(n19863), .dinb(n19765), .dout(n19864));
  jor  g19606(.dina(n9410), .dinb(n5739), .dout(n19865));
  jor  g19607(.dina(n5574), .dinb(n8809), .dout(n19866));
  jor  g19608(.dina(n5742), .dinb(n9390), .dout(n19867));
  jor  g19609(.dina(n5744), .dinb(n9413), .dout(n19868));
  jand g19610(.dina(n19868), .dinb(n19867), .dout(n19869));
  jand g19611(.dina(n19869), .dinb(n19866), .dout(n19870));
  jand g19612(.dina(n19870), .dinb(n19865), .dout(n19871));
  jxor g19613(.dina(n19871), .dinb(a44 ), .dout(n19872));
  jnot g19614(.din(n19872), .dout(n19873));
  jxor g19615(.dina(n19873), .dinb(n19864), .dout(n19874));
  jnot g19616(.din(n19619), .dout(n19875));
  jnot g19617(.din(n19715), .dout(n19876));
  jand g19618(.dina(n19876), .dinb(n19875), .dout(n19877));
  jnot g19619(.din(n19877), .dout(n19878));
  jand g19620(.dina(n19715), .dinb(n19619), .dout(n19879));
  jor  g19621(.dina(n19725), .dinb(n19879), .dout(n19880));
  jand g19622(.dina(n19880), .dinb(n19878), .dout(n19881));
  jxor g19623(.dina(n19881), .dinb(n19874), .dout(n19882));
  jor  g19624(.dina(n10634), .dinb(n5096), .dout(n19883));
  jor  g19625(.dina(n4904), .dinb(n9725), .dout(n19884));
  jor  g19626(.dina(n5099), .dinb(n10314), .dout(n19885));
  jor  g19627(.dina(n5101), .dinb(n10637), .dout(n19886));
  jand g19628(.dina(n19886), .dinb(n19885), .dout(n19887));
  jand g19629(.dina(n19887), .dinb(n19884), .dout(n19888));
  jand g19630(.dina(n19888), .dinb(n19883), .dout(n19889));
  jxor g19631(.dina(n19889), .dinb(a41 ), .dout(n19890));
  jnot g19632(.din(n19890), .dout(n19891));
  jxor g19633(.dina(n19891), .dinb(n19882), .dout(n19892));
  jxor g19634(.dina(n19892), .dinb(n19762), .dout(n19893));
  jxor g19635(.dina(n19893), .dinb(n19752), .dout(n19894));
  jxor g19636(.dina(n19894), .dinb(n19747), .dout(f101 ));
  jand g19637(.dina(n19893), .dinb(n19752), .dout(n19896));
  jand g19638(.dina(n19894), .dinb(n19747), .dout(n19897));
  jor  g19639(.dina(n19897), .dinb(n19896), .dout(n19898));
  jand g19640(.dina(n19861), .dinb(n19855), .dout(n19899));
  jand g19641(.dina(n19862), .dinb(n19774), .dout(n19900));
  jor  g19642(.dina(n19900), .dinb(n19899), .dout(n19901));
  jand g19643(.dina(n19853), .dinb(n19846), .dout(n19902));
  jand g19644(.dina(n19854), .dinb(n19783), .dout(n19903));
  jor  g19645(.dina(n19903), .dinb(n19902), .dout(n19904));
  jor  g19646(.dina(n7957), .dinb(n7266), .dout(n19905));
  jor  g19647(.dina(n7021), .dinb(n7411), .dout(n19906));
  jor  g19648(.dina(n7269), .dinb(n7683), .dout(n19907));
  jor  g19649(.dina(n7271), .dinb(n7960), .dout(n19908));
  jand g19650(.dina(n19908), .dinb(n19907), .dout(n19909));
  jand g19651(.dina(n19909), .dinb(n19906), .dout(n19910));
  jand g19652(.dina(n19910), .dinb(n19905), .dout(n19911));
  jxor g19653(.dina(n19911), .dinb(a50 ), .dout(n19912));
  jnot g19654(.din(n19912), .dout(n19913));
  jand g19655(.dina(n19835), .dinb(n19829), .dout(n19914));
  jnot g19656(.din(n19914), .dout(n19915));
  jor  g19657(.dina(n19845), .dinb(n19837), .dout(n19916));
  jand g19658(.dina(n19916), .dinb(n19915), .dout(n19917));
  jnot g19659(.din(n19917), .dout(n19918));
  jor  g19660(.dina(n8978), .dinb(n6369), .dout(n19919));
  jor  g19661(.dina(n8677), .dinb(n6106), .dout(n19920));
  jor  g19662(.dina(n8981), .dinb(n6352), .dout(n19921));
  jor  g19663(.dina(n8983), .dinb(n6372), .dout(n19922));
  jand g19664(.dina(n19922), .dinb(n19921), .dout(n19923));
  jand g19665(.dina(n19923), .dinb(n19920), .dout(n19924));
  jand g19666(.dina(n19924), .dinb(n19919), .dout(n19925));
  jxor g19667(.dina(n19925), .dinb(a56 ), .dout(n19926));
  jnot g19668(.din(n19926), .dout(n19927));
  jand g19669(.dina(n19810), .dinb(n19801), .dout(n19928));
  jand g19670(.dina(n19811), .dinb(n19792), .dout(n19929));
  jor  g19671(.dina(n19929), .dinb(n19928), .dout(n19930));
  jor  g19672(.dina(n9891), .dinb(n5859), .dout(n19931));
  jor  g19673(.dina(n9593), .dinb(n5408), .dout(n19932));
  jor  g19674(.dina(n9894), .dinb(n5428), .dout(n19933));
  jor  g19675(.dina(n9896), .dinb(n5862), .dout(n19934));
  jand g19676(.dina(n19934), .dinb(n19933), .dout(n19935));
  jand g19677(.dina(n19935), .dinb(n19932), .dout(n19936));
  jand g19678(.dina(n19936), .dinb(n19931), .dout(n19937));
  jxor g19679(.dina(n19937), .dinb(a59 ), .dout(n19938));
  jnot g19680(.din(n19938), .dout(n19939));
  jand g19681(.dina(n19804), .dinb(n19665), .dout(n19940));
  jand g19682(.dina(n19809), .dinb(n19805), .dout(n19941));
  jor  g19683(.dina(n19941), .dinb(n19940), .dout(n19942));
  jxor g19684(.dina(n19664), .dinb(n19757), .dout(n19943));
  jand g19685(.dina(n10801), .dinb(b39 ), .dout(n19944));
  jand g19686(.dina(n11107), .dinb(b38 ), .dout(n19945));
  jor  g19687(.dina(n19945), .dinb(n19944), .dout(n19946));
  jxor g19688(.dina(n19946), .dinb(n19943), .dout(n19947));
  jxor g19689(.dina(n19947), .dinb(n19942), .dout(n19948));
  jor  g19690(.dina(n10806), .dinb(n4991), .dout(n19949));
  jor  g19691(.dina(n10485), .dinb(n4557), .dout(n19950));
  jor  g19692(.dina(n10809), .dinb(n4974), .dout(n19951));
  jor  g19693(.dina(n10811), .dinb(n4994), .dout(n19952));
  jand g19694(.dina(n19952), .dinb(n19951), .dout(n19953));
  jand g19695(.dina(n19953), .dinb(n19950), .dout(n19954));
  jand g19696(.dina(n19954), .dinb(n19949), .dout(n19955));
  jxor g19697(.dina(n19955), .dinb(a62 ), .dout(n19956));
  jnot g19698(.din(n19956), .dout(n19957));
  jxor g19699(.dina(n19957), .dinb(n19948), .dout(n19958));
  jxor g19700(.dina(n19958), .dinb(n19939), .dout(n19959));
  jxor g19701(.dina(n19959), .dinb(n19930), .dout(n19960));
  jxor g19702(.dina(n19960), .dinb(n19927), .dout(n19961));
  jnot g19703(.din(n19812), .dout(n19962));
  jnot g19704(.din(n19818), .dout(n19963));
  jand g19705(.dina(n19963), .dinb(n19962), .dout(n19964));
  jnot g19706(.din(n19964), .dout(n19965));
  jand g19707(.dina(n19818), .dinb(n19812), .dout(n19966));
  jor  g19708(.dina(n19828), .dinb(n19966), .dout(n19967));
  jand g19709(.dina(n19967), .dinb(n19965), .dout(n19968));
  jxor g19710(.dina(n19968), .dinb(n19961), .dout(n19969));
  jnot g19711(.din(n19969), .dout(n19970));
  jor  g19712(.dina(n8125), .dinb(n7146), .dout(n19971));
  jor  g19713(.dina(n7846), .dinb(n6867), .dout(n19972));
  jor  g19714(.dina(n8128), .dinb(n7129), .dout(n19973));
  jor  g19715(.dina(n8130), .dinb(n7149), .dout(n19974));
  jand g19716(.dina(n19974), .dinb(n19973), .dout(n19975));
  jand g19717(.dina(n19975), .dinb(n19972), .dout(n19976));
  jand g19718(.dina(n19976), .dinb(n19971), .dout(n19977));
  jxor g19719(.dina(n19977), .dinb(a53 ), .dout(n19978));
  jxor g19720(.dina(n19978), .dinb(n19970), .dout(n19979));
  jxor g19721(.dina(n19979), .dinb(n19918), .dout(n19980));
  jxor g19722(.dina(n19980), .dinb(n19913), .dout(n19981));
  jxor g19723(.dina(n19981), .dinb(n19904), .dout(n19982));
  jnot g19724(.din(n19982), .dout(n19983));
  jor  g19725(.dina(n8806), .dinb(n6490), .dout(n19984));
  jor  g19726(.dina(n6262), .dinb(n8231), .dout(n19985));
  jor  g19727(.dina(n6493), .dinb(n8789), .dout(n19986));
  jor  g19728(.dina(n6495), .dinb(n8809), .dout(n19987));
  jand g19729(.dina(n19987), .dinb(n19986), .dout(n19988));
  jand g19730(.dina(n19988), .dinb(n19985), .dout(n19989));
  jand g19731(.dina(n19989), .dinb(n19984), .dout(n19990));
  jxor g19732(.dina(n19990), .dinb(a47 ), .dout(n19991));
  jxor g19733(.dina(n19991), .dinb(n19983), .dout(n19992));
  jxor g19734(.dina(n19992), .dinb(n19901), .dout(n19993));
  jnot g19735(.din(n19993), .dout(n19994));
  jor  g19736(.dina(n9722), .dinb(n5739), .dout(n19995));
  jor  g19737(.dina(n5574), .dinb(n9390), .dout(n19996));
  jor  g19738(.dina(n5742), .dinb(n9413), .dout(n19997));
  jor  g19739(.dina(n5744), .dinb(n9725), .dout(n19998));
  jand g19740(.dina(n19998), .dinb(n19997), .dout(n19999));
  jand g19741(.dina(n19999), .dinb(n19996), .dout(n20000));
  jand g19742(.dina(n20000), .dinb(n19995), .dout(n20001));
  jxor g19743(.dina(n20001), .dinb(a44 ), .dout(n20002));
  jxor g19744(.dina(n20002), .dinb(n19994), .dout(n20003));
  jor  g19745(.dina(n19863), .dinb(n19765), .dout(n20004));
  jand g19746(.dina(n19863), .dinb(n19765), .dout(n20005));
  jor  g19747(.dina(n19873), .dinb(n20005), .dout(n20006));
  jand g19748(.dina(n20006), .dinb(n20004), .dout(n20007));
  jxor g19749(.dina(n20007), .dinb(n20003), .dout(n20008));
  jnot g19750(.din(n20008), .dout(n20009));
  jor  g19751(.dina(n10961), .dinb(n5096), .dout(n20010));
  jor  g19752(.dina(n4904), .dinb(n10314), .dout(n20011));
  jor  g19753(.dina(n5099), .dinb(n10637), .dout(n20012));
  jor  g19754(.dina(n5101), .dinb(n10964), .dout(n20013));
  jand g19755(.dina(n20013), .dinb(n20012), .dout(n20014));
  jand g19756(.dina(n20014), .dinb(n20011), .dout(n20015));
  jand g19757(.dina(n20015), .dinb(n20010), .dout(n20016));
  jxor g19758(.dina(n20016), .dinb(a41 ), .dout(n20017));
  jxor g19759(.dina(n20017), .dinb(n20009), .dout(n20018));
  jnot g19760(.din(n19874), .dout(n20019));
  jnot g19761(.din(n19881), .dout(n20020));
  jand g19762(.dina(n20020), .dinb(n20019), .dout(n20021));
  jnot g19763(.din(n20021), .dout(n20022));
  jand g19764(.dina(n19881), .dinb(n19874), .dout(n20023));
  jor  g19765(.dina(n19891), .dinb(n20023), .dout(n20024));
  jand g19766(.dina(n20024), .dinb(n20022), .dout(n20025));
  jxor g19767(.dina(n20025), .dinb(n20018), .dout(n20026));
  jnot g19768(.din(n20026), .dout(n20027));
  jor  g19769(.dina(n19761), .dinb(n19756), .dout(n20028));
  jand g19770(.dina(n19892), .dinb(n19762), .dout(n20029));
  jnot g19771(.din(n20029), .dout(n20030));
  jand g19772(.dina(n20030), .dinb(n20028), .dout(n20031));
  jxor g19773(.dina(n20031), .dinb(n20027), .dout(n20032));
  jxor g19774(.dina(n20032), .dinb(n19898), .dout(f102 ));
  jor  g19775(.dina(n20017), .dinb(n20009), .dout(n20034));
  jand g19776(.dina(n20025), .dinb(n20018), .dout(n20035));
  jnot g19777(.din(n20035), .dout(n20036));
  jand g19778(.dina(n20036), .dinb(n20034), .dout(n20037));
  jnot g19779(.din(n20037), .dout(n20038));
  jor  g19780(.dina(n20002), .dinb(n19994), .dout(n20039));
  jand g19781(.dina(n20007), .dinb(n20003), .dout(n20040));
  jnot g19782(.din(n20040), .dout(n20041));
  jand g19783(.dina(n20041), .dinb(n20039), .dout(n20042));
  jor  g19784(.dina(n10978), .dinb(n5096), .dout(n20043));
  jor  g19785(.dina(n4904), .dinb(n10637), .dout(n20044));
  jor  g19786(.dina(n5099), .dinb(n10964), .dout(n20045));
  jand g19787(.dina(n20045), .dinb(n20044), .dout(n20046));
  jand g19788(.dina(n20046), .dinb(n20043), .dout(n20047));
  jxor g19789(.dina(n20047), .dinb(a41 ), .dout(n20048));
  jxor g19790(.dina(n20048), .dinb(n20042), .dout(n20049));
  jor  g19791(.dina(n19991), .dinb(n19983), .dout(n20050));
  jand g19792(.dina(n19992), .dinb(n19901), .dout(n20051));
  jnot g19793(.din(n20051), .dout(n20052));
  jand g19794(.dina(n20052), .dinb(n20050), .dout(n20053));
  jnot g19795(.din(n20053), .dout(n20054));
  jand g19796(.dina(n19980), .dinb(n19913), .dout(n20055));
  jand g19797(.dina(n19981), .dinb(n19904), .dout(n20056));
  jor  g19798(.dina(n20056), .dinb(n20055), .dout(n20057));
  jor  g19799(.dina(n8228), .dinb(n7266), .dout(n20058));
  jor  g19800(.dina(n7021), .dinb(n7683), .dout(n20059));
  jor  g19801(.dina(n7269), .dinb(n7960), .dout(n20060));
  jor  g19802(.dina(n7271), .dinb(n8231), .dout(n20061));
  jand g19803(.dina(n20061), .dinb(n20060), .dout(n20062));
  jand g19804(.dina(n20062), .dinb(n20059), .dout(n20063));
  jand g19805(.dina(n20063), .dinb(n20058), .dout(n20064));
  jxor g19806(.dina(n20064), .dinb(a50 ), .dout(n20065));
  jnot g19807(.din(n20065), .dout(n20066));
  jor  g19808(.dina(n19978), .dinb(n19970), .dout(n20067));
  jand g19809(.dina(n19979), .dinb(n19918), .dout(n20068));
  jnot g19810(.din(n20068), .dout(n20069));
  jand g19811(.dina(n20069), .dinb(n20067), .dout(n20070));
  jnot g19812(.din(n20070), .dout(n20071));
  jand g19813(.dina(n19960), .dinb(n19927), .dout(n20072));
  jand g19814(.dina(n19968), .dinb(n19961), .dout(n20073));
  jor  g19815(.dina(n20073), .dinb(n20072), .dout(n20074));
  jand g19816(.dina(n19958), .dinb(n19939), .dout(n20075));
  jand g19817(.dina(n19959), .dinb(n19930), .dout(n20076));
  jor  g19818(.dina(n20076), .dinb(n20075), .dout(n20077));
  jand g19819(.dina(n19664), .dinb(n19757), .dout(n20078));
  jand g19820(.dina(n19946), .dinb(n19943), .dout(n20079));
  jor  g19821(.dina(n20079), .dinb(n20078), .dout(n20080));
  jand g19822(.dina(n10801), .dinb(b40 ), .dout(n20081));
  jand g19823(.dina(n11107), .dinb(b39 ), .dout(n20082));
  jor  g19824(.dina(n20082), .dinb(n20081), .dout(n20083));
  jnot g19825(.din(n20083), .dout(n20084));
  jxor g19826(.dina(n20084), .dinb(n20080), .dout(n20085));
  jnot g19827(.din(n20085), .dout(n20086));
  jor  g19828(.dina(n10806), .dinb(n5405), .dout(n20087));
  jor  g19829(.dina(n10485), .dinb(n4974), .dout(n20088));
  jor  g19830(.dina(n10809), .dinb(n4994), .dout(n20089));
  jor  g19831(.dina(n10811), .dinb(n5408), .dout(n20090));
  jand g19832(.dina(n20090), .dinb(n20089), .dout(n20091));
  jand g19833(.dina(n20091), .dinb(n20088), .dout(n20092));
  jand g19834(.dina(n20092), .dinb(n20087), .dout(n20093));
  jxor g19835(.dina(n20093), .dinb(a62 ), .dout(n20094));
  jxor g19836(.dina(n20094), .dinb(n20086), .dout(n20095));
  jor  g19837(.dina(n19947), .dinb(n19942), .dout(n20096));
  jand g19838(.dina(n19947), .dinb(n19942), .dout(n20097));
  jor  g19839(.dina(n19957), .dinb(n20097), .dout(n20098));
  jand g19840(.dina(n20098), .dinb(n20096), .dout(n20099));
  jxor g19841(.dina(n20099), .dinb(n20095), .dout(n20100));
  jor  g19842(.dina(n9891), .dinb(n6103), .dout(n20101));
  jor  g19843(.dina(n9593), .dinb(n5428), .dout(n20102));
  jor  g19844(.dina(n9894), .dinb(n5862), .dout(n20103));
  jor  g19845(.dina(n9896), .dinb(n6106), .dout(n20104));
  jand g19846(.dina(n20104), .dinb(n20103), .dout(n20105));
  jand g19847(.dina(n20105), .dinb(n20102), .dout(n20106));
  jand g19848(.dina(n20106), .dinb(n20101), .dout(n20107));
  jxor g19849(.dina(n20107), .dinb(a59 ), .dout(n20108));
  jnot g19850(.din(n20108), .dout(n20109));
  jxor g19851(.dina(n20109), .dinb(n20100), .dout(n20110));
  jxor g19852(.dina(n20110), .dinb(n20077), .dout(n20111));
  jor  g19853(.dina(n8978), .dinb(n6864), .dout(n20112));
  jor  g19854(.dina(n8677), .dinb(n6352), .dout(n20113));
  jor  g19855(.dina(n8981), .dinb(n6372), .dout(n20114));
  jor  g19856(.dina(n8983), .dinb(n6867), .dout(n20115));
  jand g19857(.dina(n20115), .dinb(n20114), .dout(n20116));
  jand g19858(.dina(n20116), .dinb(n20113), .dout(n20117));
  jand g19859(.dina(n20117), .dinb(n20112), .dout(n20118));
  jxor g19860(.dina(n20118), .dinb(a56 ), .dout(n20119));
  jnot g19861(.din(n20119), .dout(n20120));
  jxor g19862(.dina(n20120), .dinb(n20111), .dout(n20121));
  jxor g19863(.dina(n20121), .dinb(n20074), .dout(n20122));
  jor  g19864(.dina(n8125), .dinb(n7408), .dout(n20123));
  jor  g19865(.dina(n7846), .dinb(n7129), .dout(n20124));
  jor  g19866(.dina(n8128), .dinb(n7149), .dout(n20125));
  jor  g19867(.dina(n8130), .dinb(n7411), .dout(n20126));
  jand g19868(.dina(n20126), .dinb(n20125), .dout(n20127));
  jand g19869(.dina(n20127), .dinb(n20124), .dout(n20128));
  jand g19870(.dina(n20128), .dinb(n20123), .dout(n20129));
  jxor g19871(.dina(n20129), .dinb(a53 ), .dout(n20130));
  jnot g19872(.din(n20130), .dout(n20131));
  jxor g19873(.dina(n20131), .dinb(n20122), .dout(n20132));
  jxor g19874(.dina(n20132), .dinb(n20071), .dout(n20133));
  jxor g19875(.dina(n20133), .dinb(n20066), .dout(n20134));
  jxor g19876(.dina(n20134), .dinb(n20057), .dout(n20135));
  jor  g19877(.dina(n9387), .dinb(n6490), .dout(n20136));
  jor  g19878(.dina(n6262), .dinb(n8789), .dout(n20137));
  jor  g19879(.dina(n6493), .dinb(n8809), .dout(n20138));
  jor  g19880(.dina(n6495), .dinb(n9390), .dout(n20139));
  jand g19881(.dina(n20139), .dinb(n20138), .dout(n20140));
  jand g19882(.dina(n20140), .dinb(n20137), .dout(n20141));
  jand g19883(.dina(n20141), .dinb(n20136), .dout(n20142));
  jxor g19884(.dina(n20142), .dinb(a47 ), .dout(n20143));
  jnot g19885(.din(n20143), .dout(n20144));
  jxor g19886(.dina(n20144), .dinb(n20135), .dout(n20145));
  jxor g19887(.dina(n20145), .dinb(n20054), .dout(n20146));
  jnot g19888(.din(n20146), .dout(n20147));
  jor  g19889(.dina(n10311), .dinb(n5739), .dout(n20148));
  jor  g19890(.dina(n5574), .dinb(n9413), .dout(n20149));
  jor  g19891(.dina(n5742), .dinb(n9725), .dout(n20150));
  jor  g19892(.dina(n5744), .dinb(n10314), .dout(n20151));
  jand g19893(.dina(n20151), .dinb(n20150), .dout(n20152));
  jand g19894(.dina(n20152), .dinb(n20149), .dout(n20153));
  jand g19895(.dina(n20153), .dinb(n20148), .dout(n20154));
  jxor g19896(.dina(n20154), .dinb(a44 ), .dout(n20155));
  jxor g19897(.dina(n20155), .dinb(n20147), .dout(n20156));
  jxor g19898(.dina(n20156), .dinb(n20049), .dout(n20157));
  jxor g19899(.dina(n20157), .dinb(n20038), .dout(n20158));
  jor  g19900(.dina(n20031), .dinb(n20027), .dout(n20159));
  jnot g19901(.din(n20159), .dout(n20160));
  jand g19902(.dina(n20032), .dinb(n19898), .dout(n20161));
  jor  g19903(.dina(n20161), .dinb(n20160), .dout(n20162));
  jxor g19904(.dina(n20162), .dinb(n20158), .dout(f103 ));
  jand g19905(.dina(n20157), .dinb(n20038), .dout(n20164));
  jand g19906(.dina(n20162), .dinb(n20158), .dout(n20165));
  jor  g19907(.dina(n20165), .dinb(n20164), .dout(n20166));
  jor  g19908(.dina(n20048), .dinb(n20042), .dout(n20167));
  jand g19909(.dina(n20156), .dinb(n20049), .dout(n20168));
  jnot g19910(.din(n20168), .dout(n20169));
  jand g19911(.dina(n20169), .dinb(n20167), .dout(n20170));
  jnot g19912(.din(n20170), .dout(n20171));
  jand g19913(.dina(n20145), .dinb(n20054), .dout(n20172));
  jnot g19914(.din(n20172), .dout(n20173));
  jor  g19915(.dina(n20155), .dinb(n20147), .dout(n20174));
  jand g19916(.dina(n20174), .dinb(n20173), .dout(n20175));
  jnot g19917(.din(a41 ), .dout(n20176));
  jand g19918(.dina(n11296), .dinb(n4670), .dout(n20177));
  jor  g19919(.dina(n20177), .dinb(n4905), .dout(n20178));
  jand g19920(.dina(n20178), .dinb(b63 ), .dout(n20179));
  jxor g19921(.dina(n20179), .dinb(n20176), .dout(n20180));
  jxor g19922(.dina(n20180), .dinb(n20175), .dout(n20181));
  jand g19923(.dina(n20132), .dinb(n20071), .dout(n20182));
  jand g19924(.dina(n20133), .dinb(n20066), .dout(n20183));
  jor  g19925(.dina(n20183), .dinb(n20182), .dout(n20184));
  jor  g19926(.dina(n8786), .dinb(n7266), .dout(n20185));
  jor  g19927(.dina(n7021), .dinb(n7960), .dout(n20186));
  jor  g19928(.dina(n7269), .dinb(n8231), .dout(n20187));
  jor  g19929(.dina(n7271), .dinb(n8789), .dout(n20188));
  jand g19930(.dina(n20188), .dinb(n20187), .dout(n20189));
  jand g19931(.dina(n20189), .dinb(n20186), .dout(n20190));
  jand g19932(.dina(n20190), .dinb(n20185), .dout(n20191));
  jxor g19933(.dina(n20191), .dinb(a50 ), .dout(n20192));
  jnot g19934(.din(n20192), .dout(n20193));
  jor  g19935(.dina(n7680), .dinb(n8125), .dout(n20194));
  jor  g19936(.dina(n7846), .dinb(n7149), .dout(n20195));
  jor  g19937(.dina(n8128), .dinb(n7411), .dout(n20196));
  jor  g19938(.dina(n8130), .dinb(n7683), .dout(n20197));
  jand g19939(.dina(n20197), .dinb(n20196), .dout(n20198));
  jand g19940(.dina(n20198), .dinb(n20195), .dout(n20199));
  jand g19941(.dina(n20199), .dinb(n20194), .dout(n20200));
  jxor g19942(.dina(n20200), .dinb(a53 ), .dout(n20201));
  jnot g19943(.din(n20201), .dout(n20202));
  jor  g19944(.dina(n9891), .dinb(n6349), .dout(n20203));
  jor  g19945(.dina(n9593), .dinb(n5862), .dout(n20204));
  jor  g19946(.dina(n9894), .dinb(n6106), .dout(n20205));
  jor  g19947(.dina(n9896), .dinb(n6352), .dout(n20206));
  jand g19948(.dina(n20206), .dinb(n20205), .dout(n20207));
  jand g19949(.dina(n20207), .dinb(n20204), .dout(n20208));
  jand g19950(.dina(n20208), .dinb(n20203), .dout(n20209));
  jxor g19951(.dina(n20209), .dinb(a59 ), .dout(n20210));
  jnot g19952(.din(n20210), .dout(n20211));
  jor  g19953(.dina(n10806), .dinb(n5425), .dout(n20212));
  jor  g19954(.dina(n10485), .dinb(n4994), .dout(n20213));
  jor  g19955(.dina(n10809), .dinb(n5408), .dout(n20214));
  jor  g19956(.dina(n10811), .dinb(n5428), .dout(n20215));
  jand g19957(.dina(n20215), .dinb(n20214), .dout(n20216));
  jand g19958(.dina(n20216), .dinb(n20213), .dout(n20217));
  jand g19959(.dina(n20217), .dinb(n20212), .dout(n20218));
  jxor g19960(.dina(n20218), .dinb(a62 ), .dout(n20219));
  jnot g19961(.din(n20219), .dout(n20220));
  jand g19962(.dina(n20084), .dinb(n20080), .dout(n20221));
  jnot g19963(.din(n20221), .dout(n20222));
  jor  g19964(.dina(n20094), .dinb(n20086), .dout(n20223));
  jand g19965(.dina(n20223), .dinb(n20222), .dout(n20224));
  jnot g19966(.din(n20224), .dout(n20225));
  jand g19967(.dina(n10801), .dinb(b41 ), .dout(n20226));
  jand g19968(.dina(n11107), .dinb(b40 ), .dout(n20227));
  jor  g19969(.dina(n20227), .dinb(n20226), .dout(n20228));
  jxor g19970(.dina(n20228), .dinb(n20084), .dout(n20229));
  jxor g19971(.dina(n20229), .dinb(n20225), .dout(n20230));
  jxor g19972(.dina(n20230), .dinb(n20220), .dout(n20231));
  jxor g19973(.dina(n20231), .dinb(n20211), .dout(n20232));
  jor  g19974(.dina(n20099), .dinb(n20095), .dout(n20233));
  jand g19975(.dina(n20099), .dinb(n20095), .dout(n20234));
  jor  g19976(.dina(n20109), .dinb(n20234), .dout(n20235));
  jand g19977(.dina(n20235), .dinb(n20233), .dout(n20236));
  jxor g19978(.dina(n20236), .dinb(n20232), .dout(n20237));
  jnot g19979(.din(n20237), .dout(n20238));
  jor  g19980(.dina(n8978), .dinb(n7126), .dout(n20239));
  jor  g19981(.dina(n8677), .dinb(n6372), .dout(n20240));
  jor  g19982(.dina(n8981), .dinb(n6867), .dout(n20241));
  jor  g19983(.dina(n8983), .dinb(n7129), .dout(n20242));
  jand g19984(.dina(n20242), .dinb(n20241), .dout(n20243));
  jand g19985(.dina(n20243), .dinb(n20240), .dout(n20244));
  jand g19986(.dina(n20244), .dinb(n20239), .dout(n20245));
  jxor g19987(.dina(n20245), .dinb(a56 ), .dout(n20246));
  jxor g19988(.dina(n20246), .dinb(n20238), .dout(n20247));
  jnot g19989(.din(n20077), .dout(n20248));
  jnot g19990(.din(n20110), .dout(n20249));
  jand g19991(.dina(n20249), .dinb(n20248), .dout(n20250));
  jnot g19992(.din(n20250), .dout(n20251));
  jand g19993(.dina(n20110), .dinb(n20077), .dout(n20252));
  jor  g19994(.dina(n20120), .dinb(n20252), .dout(n20253));
  jand g19995(.dina(n20253), .dinb(n20251), .dout(n20254));
  jxor g19996(.dina(n20254), .dinb(n20247), .dout(n20255));
  jxor g19997(.dina(n20255), .dinb(n20202), .dout(n20256));
  jnot g19998(.din(n20074), .dout(n20257));
  jnot g19999(.din(n20121), .dout(n20258));
  jand g20000(.dina(n20258), .dinb(n20257), .dout(n20259));
  jnot g20001(.din(n20259), .dout(n20260));
  jand g20002(.dina(n20121), .dinb(n20074), .dout(n20261));
  jor  g20003(.dina(n20131), .dinb(n20261), .dout(n20262));
  jand g20004(.dina(n20262), .dinb(n20260), .dout(n20263));
  jxor g20005(.dina(n20263), .dinb(n20256), .dout(n20264));
  jxor g20006(.dina(n20264), .dinb(n20193), .dout(n20265));
  jxor g20007(.dina(n20265), .dinb(n20184), .dout(n20266));
  jor  g20008(.dina(n9410), .dinb(n6490), .dout(n20267));
  jor  g20009(.dina(n6262), .dinb(n8809), .dout(n20268));
  jor  g20010(.dina(n6493), .dinb(n9390), .dout(n20269));
  jor  g20011(.dina(n6495), .dinb(n9413), .dout(n20270));
  jand g20012(.dina(n20270), .dinb(n20269), .dout(n20271));
  jand g20013(.dina(n20271), .dinb(n20268), .dout(n20272));
  jand g20014(.dina(n20272), .dinb(n20267), .dout(n20273));
  jxor g20015(.dina(n20273), .dinb(a47 ), .dout(n20274));
  jnot g20016(.din(n20274), .dout(n20275));
  jxor g20017(.dina(n20275), .dinb(n20266), .dout(n20276));
  jnot g20018(.din(n20057), .dout(n20277));
  jnot g20019(.din(n20134), .dout(n20278));
  jand g20020(.dina(n20278), .dinb(n20277), .dout(n20279));
  jnot g20021(.din(n20279), .dout(n20280));
  jand g20022(.dina(n20134), .dinb(n20057), .dout(n20281));
  jor  g20023(.dina(n20144), .dinb(n20281), .dout(n20282));
  jand g20024(.dina(n20282), .dinb(n20280), .dout(n20283));
  jxor g20025(.dina(n20283), .dinb(n20276), .dout(n20284));
  jor  g20026(.dina(n10634), .dinb(n5739), .dout(n20285));
  jor  g20027(.dina(n5574), .dinb(n9725), .dout(n20286));
  jor  g20028(.dina(n5742), .dinb(n10314), .dout(n20287));
  jor  g20029(.dina(n5744), .dinb(n10637), .dout(n20288));
  jand g20030(.dina(n20288), .dinb(n20287), .dout(n20289));
  jand g20031(.dina(n20289), .dinb(n20286), .dout(n20290));
  jand g20032(.dina(n20290), .dinb(n20285), .dout(n20291));
  jxor g20033(.dina(n20291), .dinb(a44 ), .dout(n20292));
  jnot g20034(.din(n20292), .dout(n20293));
  jxor g20035(.dina(n20293), .dinb(n20284), .dout(n20294));
  jxor g20036(.dina(n20294), .dinb(n20181), .dout(n20295));
  jxor g20037(.dina(n20295), .dinb(n20171), .dout(n20296));
  jxor g20038(.dina(n20296), .dinb(n20166), .dout(f104 ));
  jand g20039(.dina(n20295), .dinb(n20171), .dout(n20298));
  jand g20040(.dina(n20296), .dinb(n20166), .dout(n20299));
  jor  g20041(.dina(n20299), .dinb(n20298), .dout(n20300));
  jand g20042(.dina(n20263), .dinb(n20256), .dout(n20301));
  jand g20043(.dina(n20264), .dinb(n20193), .dout(n20302));
  jor  g20044(.dina(n20302), .dinb(n20301), .dout(n20303));
  jor  g20045(.dina(n8806), .dinb(n7266), .dout(n20304));
  jor  g20046(.dina(n7021), .dinb(n8231), .dout(n20305));
  jor  g20047(.dina(n7269), .dinb(n8789), .dout(n20306));
  jor  g20048(.dina(n7271), .dinb(n8809), .dout(n20307));
  jand g20049(.dina(n20307), .dinb(n20306), .dout(n20308));
  jand g20050(.dina(n20308), .dinb(n20305), .dout(n20309));
  jand g20051(.dina(n20309), .dinb(n20304), .dout(n20310));
  jxor g20052(.dina(n20310), .dinb(a50 ), .dout(n20311));
  jnot g20053(.din(n20311), .dout(n20312));
  jand g20054(.dina(n20254), .dinb(n20247), .dout(n20313));
  jand g20055(.dina(n20255), .dinb(n20202), .dout(n20314));
  jor  g20056(.dina(n20314), .dinb(n20313), .dout(n20315));
  jor  g20057(.dina(n7957), .dinb(n8125), .dout(n20316));
  jor  g20058(.dina(n7846), .dinb(n7411), .dout(n20317));
  jor  g20059(.dina(n8128), .dinb(n7683), .dout(n20318));
  jor  g20060(.dina(n8130), .dinb(n7960), .dout(n20319));
  jand g20061(.dina(n20319), .dinb(n20318), .dout(n20320));
  jand g20062(.dina(n20320), .dinb(n20317), .dout(n20321));
  jand g20063(.dina(n20321), .dinb(n20316), .dout(n20322));
  jxor g20064(.dina(n20322), .dinb(a53 ), .dout(n20323));
  jnot g20065(.din(n20323), .dout(n20324));
  jand g20066(.dina(n20236), .dinb(n20232), .dout(n20325));
  jnot g20067(.din(n20325), .dout(n20326));
  jor  g20068(.dina(n20246), .dinb(n20238), .dout(n20327));
  jand g20069(.dina(n20327), .dinb(n20326), .dout(n20328));
  jnot g20070(.din(n20328), .dout(n20329));
  jor  g20071(.dina(n8978), .dinb(n7146), .dout(n20330));
  jor  g20072(.dina(n8677), .dinb(n6867), .dout(n20331));
  jor  g20073(.dina(n8981), .dinb(n7129), .dout(n20332));
  jor  g20074(.dina(n8983), .dinb(n7149), .dout(n20333));
  jand g20075(.dina(n20333), .dinb(n20332), .dout(n20334));
  jand g20076(.dina(n20334), .dinb(n20331), .dout(n20335));
  jand g20077(.dina(n20335), .dinb(n20330), .dout(n20336));
  jxor g20078(.dina(n20336), .dinb(a56 ), .dout(n20337));
  jnot g20079(.din(n20337), .dout(n20338));
  jand g20080(.dina(n20230), .dinb(n20220), .dout(n20339));
  jand g20081(.dina(n20231), .dinb(n20211), .dout(n20340));
  jor  g20082(.dina(n20340), .dinb(n20339), .dout(n20341));
  jand g20083(.dina(n20228), .dinb(n20084), .dout(n20342));
  jand g20084(.dina(n20229), .dinb(n20225), .dout(n20343));
  jor  g20085(.dina(n20343), .dinb(n20342), .dout(n20344));
  jxor g20086(.dina(n20083), .dinb(n20176), .dout(n20345));
  jand g20087(.dina(n10801), .dinb(b42 ), .dout(n20346));
  jand g20088(.dina(n11107), .dinb(b41 ), .dout(n20347));
  jor  g20089(.dina(n20347), .dinb(n20346), .dout(n20348));
  jxor g20090(.dina(n20348), .dinb(n20345), .dout(n20349));
  jnot g20091(.din(n20349), .dout(n20350));
  jor  g20092(.dina(n10806), .dinb(n5859), .dout(n20351));
  jor  g20093(.dina(n10485), .dinb(n5408), .dout(n20352));
  jor  g20094(.dina(n10809), .dinb(n5428), .dout(n20353));
  jor  g20095(.dina(n10811), .dinb(n5862), .dout(n20354));
  jand g20096(.dina(n20354), .dinb(n20353), .dout(n20355));
  jand g20097(.dina(n20355), .dinb(n20352), .dout(n20356));
  jand g20098(.dina(n20356), .dinb(n20351), .dout(n20357));
  jxor g20099(.dina(n20357), .dinb(a62 ), .dout(n20358));
  jxor g20100(.dina(n20358), .dinb(n20350), .dout(n20359));
  jxor g20101(.dina(n20359), .dinb(n20344), .dout(n20360));
  jnot g20102(.din(n20360), .dout(n20361));
  jor  g20103(.dina(n9891), .dinb(n6369), .dout(n20362));
  jor  g20104(.dina(n9593), .dinb(n6106), .dout(n20363));
  jor  g20105(.dina(n9894), .dinb(n6352), .dout(n20364));
  jor  g20106(.dina(n9896), .dinb(n6372), .dout(n20365));
  jand g20107(.dina(n20365), .dinb(n20364), .dout(n20366));
  jand g20108(.dina(n20366), .dinb(n20363), .dout(n20367));
  jand g20109(.dina(n20367), .dinb(n20362), .dout(n20368));
  jxor g20110(.dina(n20368), .dinb(a59 ), .dout(n20369));
  jxor g20111(.dina(n20369), .dinb(n20361), .dout(n20370));
  jxor g20112(.dina(n20370), .dinb(n20341), .dout(n20371));
  jxor g20113(.dina(n20371), .dinb(n20338), .dout(n20372));
  jxor g20114(.dina(n20372), .dinb(n20329), .dout(n20373));
  jxor g20115(.dina(n20373), .dinb(n20324), .dout(n20374));
  jxor g20116(.dina(n20374), .dinb(n20315), .dout(n20375));
  jxor g20117(.dina(n20375), .dinb(n20312), .dout(n20376));
  jxor g20118(.dina(n20376), .dinb(n20303), .dout(n20377));
  jnot g20119(.din(n20377), .dout(n20378));
  jor  g20120(.dina(n9722), .dinb(n6490), .dout(n20379));
  jor  g20121(.dina(n6262), .dinb(n9390), .dout(n20380));
  jor  g20122(.dina(n6493), .dinb(n9413), .dout(n20381));
  jor  g20123(.dina(n6495), .dinb(n9725), .dout(n20382));
  jand g20124(.dina(n20382), .dinb(n20381), .dout(n20383));
  jand g20125(.dina(n20383), .dinb(n20380), .dout(n20384));
  jand g20126(.dina(n20384), .dinb(n20379), .dout(n20385));
  jxor g20127(.dina(n20385), .dinb(a47 ), .dout(n20386));
  jxor g20128(.dina(n20386), .dinb(n20378), .dout(n20387));
  jor  g20129(.dina(n20265), .dinb(n20184), .dout(n20388));
  jand g20130(.dina(n20265), .dinb(n20184), .dout(n20389));
  jor  g20131(.dina(n20275), .dinb(n20389), .dout(n20390));
  jand g20132(.dina(n20390), .dinb(n20388), .dout(n20391));
  jxor g20133(.dina(n20391), .dinb(n20387), .dout(n20392));
  jnot g20134(.din(n20392), .dout(n20393));
  jor  g20135(.dina(n10961), .dinb(n5739), .dout(n20394));
  jor  g20136(.dina(n5574), .dinb(n10314), .dout(n20395));
  jor  g20137(.dina(n5742), .dinb(n10637), .dout(n20396));
  jor  g20138(.dina(n5744), .dinb(n10964), .dout(n20397));
  jand g20139(.dina(n20397), .dinb(n20396), .dout(n20398));
  jand g20140(.dina(n20398), .dinb(n20395), .dout(n20399));
  jand g20141(.dina(n20399), .dinb(n20394), .dout(n20400));
  jxor g20142(.dina(n20400), .dinb(a44 ), .dout(n20401));
  jxor g20143(.dina(n20401), .dinb(n20393), .dout(n20402));
  jnot g20144(.din(n20276), .dout(n20403));
  jnot g20145(.din(n20283), .dout(n20404));
  jand g20146(.dina(n20404), .dinb(n20403), .dout(n20405));
  jnot g20147(.din(n20405), .dout(n20406));
  jand g20148(.dina(n20283), .dinb(n20276), .dout(n20407));
  jor  g20149(.dina(n20293), .dinb(n20407), .dout(n20408));
  jand g20150(.dina(n20408), .dinb(n20406), .dout(n20409));
  jxor g20151(.dina(n20409), .dinb(n20402), .dout(n20410));
  jnot g20152(.din(n20410), .dout(n20411));
  jor  g20153(.dina(n20180), .dinb(n20175), .dout(n20412));
  jand g20154(.dina(n20294), .dinb(n20181), .dout(n20413));
  jnot g20155(.din(n20413), .dout(n20414));
  jand g20156(.dina(n20414), .dinb(n20412), .dout(n20415));
  jxor g20157(.dina(n20415), .dinb(n20411), .dout(n20416));
  jxor g20158(.dina(n20416), .dinb(n20300), .dout(f105 ));
  jor  g20159(.dina(n20401), .dinb(n20393), .dout(n20418));
  jand g20160(.dina(n20409), .dinb(n20402), .dout(n20419));
  jnot g20161(.din(n20419), .dout(n20420));
  jand g20162(.dina(n20420), .dinb(n20418), .dout(n20421));
  jnot g20163(.din(n20421), .dout(n20422));
  jor  g20164(.dina(n20386), .dinb(n20378), .dout(n20423));
  jand g20165(.dina(n20391), .dinb(n20387), .dout(n20424));
  jnot g20166(.din(n20424), .dout(n20425));
  jand g20167(.dina(n20425), .dinb(n20423), .dout(n20426));
  jor  g20168(.dina(n10978), .dinb(n5739), .dout(n20427));
  jor  g20169(.dina(n5574), .dinb(n10637), .dout(n20428));
  jor  g20170(.dina(n5742), .dinb(n10964), .dout(n20429));
  jand g20171(.dina(n20429), .dinb(n20428), .dout(n20430));
  jand g20172(.dina(n20430), .dinb(n20427), .dout(n20431));
  jxor g20173(.dina(n20431), .dinb(a44 ), .dout(n20432));
  jxor g20174(.dina(n20432), .dinb(n20426), .dout(n20433));
  jor  g20175(.dina(n10311), .dinb(n6490), .dout(n20434));
  jor  g20176(.dina(n6262), .dinb(n9413), .dout(n20435));
  jor  g20177(.dina(n6493), .dinb(n9725), .dout(n20436));
  jor  g20178(.dina(n6495), .dinb(n10314), .dout(n20437));
  jand g20179(.dina(n20437), .dinb(n20436), .dout(n20438));
  jand g20180(.dina(n20438), .dinb(n20435), .dout(n20439));
  jand g20181(.dina(n20439), .dinb(n20434), .dout(n20440));
  jxor g20182(.dina(n20440), .dinb(a47 ), .dout(n20441));
  jnot g20183(.din(n20441), .dout(n20442));
  jand g20184(.dina(n20375), .dinb(n20312), .dout(n20443));
  jand g20185(.dina(n20376), .dinb(n20303), .dout(n20444));
  jor  g20186(.dina(n20444), .dinb(n20443), .dout(n20445));
  jor  g20187(.dina(n9387), .dinb(n7266), .dout(n20446));
  jor  g20188(.dina(n7021), .dinb(n8789), .dout(n20447));
  jor  g20189(.dina(n7269), .dinb(n8809), .dout(n20448));
  jor  g20190(.dina(n7271), .dinb(n9390), .dout(n20449));
  jand g20191(.dina(n20449), .dinb(n20448), .dout(n20450));
  jand g20192(.dina(n20450), .dinb(n20447), .dout(n20451));
  jand g20193(.dina(n20451), .dinb(n20446), .dout(n20452));
  jxor g20194(.dina(n20452), .dinb(a50 ), .dout(n20453));
  jnot g20195(.din(n20453), .dout(n20454));
  jand g20196(.dina(n20373), .dinb(n20324), .dout(n20455));
  jand g20197(.dina(n20374), .dinb(n20315), .dout(n20456));
  jor  g20198(.dina(n20456), .dinb(n20455), .dout(n20457));
  jand g20199(.dina(n20371), .dinb(n20338), .dout(n20458));
  jand g20200(.dina(n20372), .dinb(n20329), .dout(n20459));
  jor  g20201(.dina(n20459), .dinb(n20458), .dout(n20460));
  jor  g20202(.dina(n20369), .dinb(n20361), .dout(n20461));
  jand g20203(.dina(n20370), .dinb(n20341), .dout(n20462));
  jnot g20204(.din(n20462), .dout(n20463));
  jand g20205(.dina(n20463), .dinb(n20461), .dout(n20464));
  jnot g20206(.din(n20464), .dout(n20465));
  jor  g20207(.dina(n20358), .dinb(n20350), .dout(n20466));
  jand g20208(.dina(n20359), .dinb(n20344), .dout(n20467));
  jnot g20209(.din(n20467), .dout(n20468));
  jand g20210(.dina(n20468), .dinb(n20466), .dout(n20469));
  jnot g20211(.din(n20469), .dout(n20470));
  jor  g20212(.dina(n10806), .dinb(n6103), .dout(n20471));
  jor  g20213(.dina(n10485), .dinb(n5428), .dout(n20472));
  jor  g20214(.dina(n10809), .dinb(n5862), .dout(n20473));
  jor  g20215(.dina(n10811), .dinb(n6106), .dout(n20474));
  jand g20216(.dina(n20474), .dinb(n20473), .dout(n20475));
  jand g20217(.dina(n20475), .dinb(n20472), .dout(n20476));
  jand g20218(.dina(n20476), .dinb(n20471), .dout(n20477));
  jxor g20219(.dina(n20477), .dinb(a62 ), .dout(n20478));
  jnot g20220(.din(n20478), .dout(n20479));
  jand g20221(.dina(n20083), .dinb(n20176), .dout(n20480));
  jand g20222(.dina(n20348), .dinb(n20345), .dout(n20481));
  jor  g20223(.dina(n20481), .dinb(n20480), .dout(n20482));
  jand g20224(.dina(n10801), .dinb(b43 ), .dout(n20483));
  jand g20225(.dina(n11107), .dinb(b42 ), .dout(n20484));
  jor  g20226(.dina(n20484), .dinb(n20483), .dout(n20485));
  jnot g20227(.din(n20485), .dout(n20486));
  jxor g20228(.dina(n20486), .dinb(n20482), .dout(n20487));
  jxor g20229(.dina(n20487), .dinb(n20479), .dout(n20488));
  jxor g20230(.dina(n20488), .dinb(n20470), .dout(n20489));
  jor  g20231(.dina(n9891), .dinb(n6864), .dout(n20490));
  jor  g20232(.dina(n9593), .dinb(n6352), .dout(n20491));
  jor  g20233(.dina(n9894), .dinb(n6372), .dout(n20492));
  jor  g20234(.dina(n9896), .dinb(n6867), .dout(n20493));
  jand g20235(.dina(n20493), .dinb(n20492), .dout(n20494));
  jand g20236(.dina(n20494), .dinb(n20491), .dout(n20495));
  jand g20237(.dina(n20495), .dinb(n20490), .dout(n20496));
  jxor g20238(.dina(n20496), .dinb(a59 ), .dout(n20497));
  jnot g20239(.din(n20497), .dout(n20498));
  jxor g20240(.dina(n20498), .dinb(n20489), .dout(n20499));
  jxor g20241(.dina(n20499), .dinb(n20465), .dout(n20500));
  jor  g20242(.dina(n8978), .dinb(n7408), .dout(n20501));
  jor  g20243(.dina(n8677), .dinb(n7129), .dout(n20502));
  jor  g20244(.dina(n8981), .dinb(n7149), .dout(n20503));
  jor  g20245(.dina(n8983), .dinb(n7411), .dout(n20504));
  jand g20246(.dina(n20504), .dinb(n20503), .dout(n20505));
  jand g20247(.dina(n20505), .dinb(n20502), .dout(n20506));
  jand g20248(.dina(n20506), .dinb(n20501), .dout(n20507));
  jxor g20249(.dina(n20507), .dinb(a56 ), .dout(n20508));
  jnot g20250(.din(n20508), .dout(n20509));
  jxor g20251(.dina(n20509), .dinb(n20500), .dout(n20510));
  jxor g20252(.dina(n20510), .dinb(n20460), .dout(n20511));
  jor  g20253(.dina(n8228), .dinb(n8125), .dout(n20512));
  jor  g20254(.dina(n7846), .dinb(n7683), .dout(n20513));
  jor  g20255(.dina(n8128), .dinb(n7960), .dout(n20514));
  jor  g20256(.dina(n8130), .dinb(n8231), .dout(n20515));
  jand g20257(.dina(n20515), .dinb(n20514), .dout(n20516));
  jand g20258(.dina(n20516), .dinb(n20513), .dout(n20517));
  jand g20259(.dina(n20517), .dinb(n20512), .dout(n20518));
  jxor g20260(.dina(n20518), .dinb(a53 ), .dout(n20519));
  jnot g20261(.din(n20519), .dout(n20520));
  jxor g20262(.dina(n20520), .dinb(n20511), .dout(n20521));
  jxor g20263(.dina(n20521), .dinb(n20457), .dout(n20522));
  jxor g20264(.dina(n20522), .dinb(n20454), .dout(n20523));
  jxor g20265(.dina(n20523), .dinb(n20445), .dout(n20524));
  jxor g20266(.dina(n20524), .dinb(n20442), .dout(n20525));
  jxor g20267(.dina(n20525), .dinb(n20433), .dout(n20526));
  jxor g20268(.dina(n20526), .dinb(n20422), .dout(n20527));
  jor  g20269(.dina(n20415), .dinb(n20411), .dout(n20528));
  jnot g20270(.din(n20528), .dout(n20529));
  jand g20271(.dina(n20416), .dinb(n20300), .dout(n20530));
  jor  g20272(.dina(n20530), .dinb(n20529), .dout(n20531));
  jxor g20273(.dina(n20531), .dinb(n20527), .dout(f106 ));
  jand g20274(.dina(n20526), .dinb(n20422), .dout(n20533));
  jand g20275(.dina(n20531), .dinb(n20527), .dout(n20534));
  jor  g20276(.dina(n20534), .dinb(n20533), .dout(n20535));
  jnot g20277(.din(a44 ), .dout(n20536));
  jand g20278(.dina(n11296), .dinb(n5298), .dout(n20537));
  jor  g20279(.dina(n20537), .dinb(n5575), .dout(n20538));
  jand g20280(.dina(n20538), .dinb(b63 ), .dout(n20539));
  jxor g20281(.dina(n20539), .dinb(n20536), .dout(n20540));
  jnot g20282(.din(n20540), .dout(n20541));
  jor  g20283(.dina(n20523), .dinb(n20445), .dout(n20542));
  jand g20284(.dina(n20523), .dinb(n20445), .dout(n20543));
  jor  g20285(.dina(n20543), .dinb(n20442), .dout(n20544));
  jand g20286(.dina(n20544), .dinb(n20542), .dout(n20545));
  jxor g20287(.dina(n20545), .dinb(n20541), .dout(n20546));
  jor  g20288(.dina(n10634), .dinb(n6490), .dout(n20547));
  jor  g20289(.dina(n6262), .dinb(n9725), .dout(n20548));
  jor  g20290(.dina(n6493), .dinb(n10314), .dout(n20549));
  jor  g20291(.dina(n6495), .dinb(n10637), .dout(n20550));
  jand g20292(.dina(n20550), .dinb(n20549), .dout(n20551));
  jand g20293(.dina(n20551), .dinb(n20548), .dout(n20552));
  jand g20294(.dina(n20552), .dinb(n20547), .dout(n20553));
  jxor g20295(.dina(n20553), .dinb(a47 ), .dout(n20554));
  jnot g20296(.din(n20554), .dout(n20555));
  jand g20297(.dina(n20521), .dinb(n20457), .dout(n20556));
  jand g20298(.dina(n20522), .dinb(n20454), .dout(n20557));
  jor  g20299(.dina(n20557), .dinb(n20556), .dout(n20558));
  jor  g20300(.dina(n8786), .dinb(n8125), .dout(n20559));
  jor  g20301(.dina(n7846), .dinb(n7960), .dout(n20560));
  jor  g20302(.dina(n8128), .dinb(n8231), .dout(n20561));
  jor  g20303(.dina(n8130), .dinb(n8789), .dout(n20562));
  jand g20304(.dina(n20562), .dinb(n20561), .dout(n20563));
  jand g20305(.dina(n20563), .dinb(n20560), .dout(n20564));
  jand g20306(.dina(n20564), .dinb(n20559), .dout(n20565));
  jxor g20307(.dina(n20565), .dinb(a53 ), .dout(n20566));
  jnot g20308(.din(n20566), .dout(n20567));
  jor  g20309(.dina(n8978), .dinb(n7680), .dout(n20568));
  jor  g20310(.dina(n8677), .dinb(n7149), .dout(n20569));
  jor  g20311(.dina(n8981), .dinb(n7411), .dout(n20570));
  jor  g20312(.dina(n8983), .dinb(n7683), .dout(n20571));
  jand g20313(.dina(n20571), .dinb(n20570), .dout(n20572));
  jand g20314(.dina(n20572), .dinb(n20569), .dout(n20573));
  jand g20315(.dina(n20573), .dinb(n20568), .dout(n20574));
  jxor g20316(.dina(n20574), .dinb(a56 ), .dout(n20575));
  jnot g20317(.din(n20575), .dout(n20576));
  jor  g20318(.dina(n9891), .dinb(n7126), .dout(n20577));
  jor  g20319(.dina(n9593), .dinb(n6372), .dout(n20578));
  jor  g20320(.dina(n9894), .dinb(n6867), .dout(n20579));
  jor  g20321(.dina(n9896), .dinb(n7129), .dout(n20580));
  jand g20322(.dina(n20580), .dinb(n20579), .dout(n20581));
  jand g20323(.dina(n20581), .dinb(n20578), .dout(n20582));
  jand g20324(.dina(n20582), .dinb(n20577), .dout(n20583));
  jxor g20325(.dina(n20583), .dinb(a59 ), .dout(n20584));
  jnot g20326(.din(n20584), .dout(n20585));
  jand g20327(.dina(n20486), .dinb(n20482), .dout(n20586));
  jand g20328(.dina(n20487), .dinb(n20479), .dout(n20587));
  jor  g20329(.dina(n20587), .dinb(n20586), .dout(n20588));
  jand g20330(.dina(n10801), .dinb(b44 ), .dout(n20589));
  jand g20331(.dina(n11107), .dinb(b43 ), .dout(n20590));
  jor  g20332(.dina(n20590), .dinb(n20589), .dout(n20591));
  jxor g20333(.dina(n20591), .dinb(n20486), .dout(n20592));
  jnot g20334(.din(n20592), .dout(n20593));
  jor  g20335(.dina(n10806), .dinb(n6349), .dout(n20594));
  jor  g20336(.dina(n10485), .dinb(n5862), .dout(n20595));
  jor  g20337(.dina(n10809), .dinb(n6106), .dout(n20596));
  jor  g20338(.dina(n10811), .dinb(n6352), .dout(n20597));
  jand g20339(.dina(n20597), .dinb(n20596), .dout(n20598));
  jand g20340(.dina(n20598), .dinb(n20595), .dout(n20599));
  jand g20341(.dina(n20599), .dinb(n20594), .dout(n20600));
  jxor g20342(.dina(n20600), .dinb(a62 ), .dout(n20601));
  jxor g20343(.dina(n20601), .dinb(n20593), .dout(n20602));
  jxor g20344(.dina(n20602), .dinb(n20588), .dout(n20603));
  jxor g20345(.dina(n20603), .dinb(n20585), .dout(n20604));
  jor  g20346(.dina(n20488), .dinb(n20470), .dout(n20605));
  jand g20347(.dina(n20488), .dinb(n20470), .dout(n20606));
  jor  g20348(.dina(n20498), .dinb(n20606), .dout(n20607));
  jand g20349(.dina(n20607), .dinb(n20605), .dout(n20608));
  jxor g20350(.dina(n20608), .dinb(n20604), .dout(n20609));
  jxor g20351(.dina(n20609), .dinb(n20576), .dout(n20610));
  jnot g20352(.din(n20499), .dout(n20611));
  jand g20353(.dina(n20611), .dinb(n20464), .dout(n20612));
  jnot g20354(.din(n20612), .dout(n20613));
  jand g20355(.dina(n20499), .dinb(n20465), .dout(n20614));
  jor  g20356(.dina(n20509), .dinb(n20614), .dout(n20615));
  jand g20357(.dina(n20615), .dinb(n20613), .dout(n20616));
  jxor g20358(.dina(n20616), .dinb(n20610), .dout(n20617));
  jxor g20359(.dina(n20617), .dinb(n20567), .dout(n20618));
  jnot g20360(.din(n20460), .dout(n20619));
  jnot g20361(.din(n20510), .dout(n20620));
  jand g20362(.dina(n20620), .dinb(n20619), .dout(n20621));
  jnot g20363(.din(n20621), .dout(n20622));
  jand g20364(.dina(n20510), .dinb(n20460), .dout(n20623));
  jor  g20365(.dina(n20520), .dinb(n20623), .dout(n20624));
  jand g20366(.dina(n20624), .dinb(n20622), .dout(n20625));
  jxor g20367(.dina(n20625), .dinb(n20618), .dout(n20626));
  jor  g20368(.dina(n9410), .dinb(n7266), .dout(n20627));
  jor  g20369(.dina(n7021), .dinb(n8809), .dout(n20628));
  jor  g20370(.dina(n7269), .dinb(n9390), .dout(n20629));
  jor  g20371(.dina(n7271), .dinb(n9413), .dout(n20630));
  jand g20372(.dina(n20630), .dinb(n20629), .dout(n20631));
  jand g20373(.dina(n20631), .dinb(n20628), .dout(n20632));
  jand g20374(.dina(n20632), .dinb(n20627), .dout(n20633));
  jxor g20375(.dina(n20633), .dinb(a50 ), .dout(n20634));
  jnot g20376(.din(n20634), .dout(n20635));
  jxor g20377(.dina(n20635), .dinb(n20626), .dout(n20636));
  jxor g20378(.dina(n20636), .dinb(n20558), .dout(n20637));
  jxor g20379(.dina(n20637), .dinb(n20555), .dout(n20638));
  jxor g20380(.dina(n20638), .dinb(n20546), .dout(n20639));
  jand g20381(.dina(n20432), .dinb(n20426), .dout(n20640));
  jnot g20382(.din(n20640), .dout(n20641));
  jnot g20383(.din(n20426), .dout(n20642));
  jnot g20384(.din(n20432), .dout(n20643));
  jand g20385(.dina(n20643), .dinb(n20642), .dout(n20644));
  jor  g20386(.dina(n20525), .dinb(n20644), .dout(n20645));
  jand g20387(.dina(n20645), .dinb(n20641), .dout(n20646));
  jxor g20388(.dina(n20646), .dinb(n20639), .dout(n20647));
  jxor g20389(.dina(n20647), .dinb(n20535), .dout(f107 ));
  jand g20390(.dina(n20646), .dinb(n20639), .dout(n20649));
  jand g20391(.dina(n20647), .dinb(n20535), .dout(n20650));
  jor  g20392(.dina(n20650), .dinb(n20649), .dout(n20651));
  jor  g20393(.dina(n9722), .dinb(n7266), .dout(n20652));
  jor  g20394(.dina(n7021), .dinb(n9390), .dout(n20653));
  jor  g20395(.dina(n7269), .dinb(n9413), .dout(n20654));
  jor  g20396(.dina(n7271), .dinb(n9725), .dout(n20655));
  jand g20397(.dina(n20655), .dinb(n20654), .dout(n20656));
  jand g20398(.dina(n20656), .dinb(n20653), .dout(n20657));
  jand g20399(.dina(n20657), .dinb(n20652), .dout(n20658));
  jxor g20400(.dina(n20658), .dinb(a50 ), .dout(n20659));
  jnot g20401(.din(n20659), .dout(n20660));
  jand g20402(.dina(n20616), .dinb(n20610), .dout(n20661));
  jand g20403(.dina(n20617), .dinb(n20567), .dout(n20662));
  jor  g20404(.dina(n20662), .dinb(n20661), .dout(n20663));
  jor  g20405(.dina(n8806), .dinb(n8125), .dout(n20664));
  jor  g20406(.dina(n7846), .dinb(n8231), .dout(n20665));
  jor  g20407(.dina(n8128), .dinb(n8789), .dout(n20666));
  jor  g20408(.dina(n8130), .dinb(n8809), .dout(n20667));
  jand g20409(.dina(n20667), .dinb(n20666), .dout(n20668));
  jand g20410(.dina(n20668), .dinb(n20665), .dout(n20669));
  jand g20411(.dina(n20669), .dinb(n20664), .dout(n20670));
  jxor g20412(.dina(n20670), .dinb(a53 ), .dout(n20671));
  jnot g20413(.din(n20671), .dout(n20672));
  jand g20414(.dina(n20608), .dinb(n20604), .dout(n20673));
  jand g20415(.dina(n20609), .dinb(n20576), .dout(n20674));
  jor  g20416(.dina(n20674), .dinb(n20673), .dout(n20675));
  jor  g20417(.dina(n8978), .dinb(n7957), .dout(n20676));
  jor  g20418(.dina(n8677), .dinb(n7411), .dout(n20677));
  jor  g20419(.dina(n8981), .dinb(n7683), .dout(n20678));
  jor  g20420(.dina(n8983), .dinb(n7960), .dout(n20679));
  jand g20421(.dina(n20679), .dinb(n20678), .dout(n20680));
  jand g20422(.dina(n20680), .dinb(n20677), .dout(n20681));
  jand g20423(.dina(n20681), .dinb(n20676), .dout(n20682));
  jxor g20424(.dina(n20682), .dinb(a56 ), .dout(n20683));
  jnot g20425(.din(n20683), .dout(n20684));
  jand g20426(.dina(n20602), .dinb(n20588), .dout(n20685));
  jand g20427(.dina(n20603), .dinb(n20585), .dout(n20686));
  jor  g20428(.dina(n20686), .dinb(n20685), .dout(n20687));
  jor  g20429(.dina(n9891), .dinb(n7146), .dout(n20688));
  jor  g20430(.dina(n9593), .dinb(n6867), .dout(n20689));
  jor  g20431(.dina(n9894), .dinb(n7129), .dout(n20690));
  jor  g20432(.dina(n9896), .dinb(n7149), .dout(n20691));
  jand g20433(.dina(n20691), .dinb(n20690), .dout(n20692));
  jand g20434(.dina(n20692), .dinb(n20689), .dout(n20693));
  jand g20435(.dina(n20693), .dinb(n20688), .dout(n20694));
  jxor g20436(.dina(n20694), .dinb(a59 ), .dout(n20695));
  jnot g20437(.din(n20695), .dout(n20696));
  jor  g20438(.dina(n10806), .dinb(n6369), .dout(n20697));
  jor  g20439(.dina(n10485), .dinb(n6106), .dout(n20698));
  jor  g20440(.dina(n10809), .dinb(n6352), .dout(n20699));
  jor  g20441(.dina(n10811), .dinb(n6372), .dout(n20700));
  jand g20442(.dina(n20700), .dinb(n20699), .dout(n20701));
  jand g20443(.dina(n20701), .dinb(n20698), .dout(n20702));
  jand g20444(.dina(n20702), .dinb(n20697), .dout(n20703));
  jxor g20445(.dina(n20703), .dinb(a62 ), .dout(n20704));
  jnot g20446(.din(n20704), .dout(n20705));
  jand g20447(.dina(n20591), .dinb(n20486), .dout(n20706));
  jnot g20448(.din(n20706), .dout(n20707));
  jor  g20449(.dina(n20601), .dinb(n20593), .dout(n20708));
  jand g20450(.dina(n20708), .dinb(n20707), .dout(n20709));
  jnot g20451(.din(n20709), .dout(n20710));
  jand g20452(.dina(n10801), .dinb(b45 ), .dout(n20711));
  jand g20453(.dina(n11107), .dinb(b44 ), .dout(n20712));
  jor  g20454(.dina(n20712), .dinb(n20711), .dout(n20713));
  jxor g20455(.dina(n20713), .dinb(n20536), .dout(n20714));
  jxor g20456(.dina(n20714), .dinb(n20485), .dout(n20715));
  jxor g20457(.dina(n20715), .dinb(n20710), .dout(n20716));
  jxor g20458(.dina(n20716), .dinb(n20705), .dout(n20717));
  jxor g20459(.dina(n20717), .dinb(n20696), .dout(n20718));
  jxor g20460(.dina(n20718), .dinb(n20687), .dout(n20719));
  jxor g20461(.dina(n20719), .dinb(n20684), .dout(n20720));
  jxor g20462(.dina(n20720), .dinb(n20675), .dout(n20721));
  jxor g20463(.dina(n20721), .dinb(n20672), .dout(n20722));
  jxor g20464(.dina(n20722), .dinb(n20663), .dout(n20723));
  jxor g20465(.dina(n20723), .dinb(n20660), .dout(n20724));
  jor  g20466(.dina(n20625), .dinb(n20618), .dout(n20725));
  jand g20467(.dina(n20625), .dinb(n20618), .dout(n20726));
  jor  g20468(.dina(n20635), .dinb(n20726), .dout(n20727));
  jand g20469(.dina(n20727), .dinb(n20725), .dout(n20728));
  jxor g20470(.dina(n20728), .dinb(n20724), .dout(n20729));
  jnot g20471(.din(n20729), .dout(n20730));
  jor  g20472(.dina(n10961), .dinb(n6490), .dout(n20731));
  jor  g20473(.dina(n6262), .dinb(n10314), .dout(n20732));
  jor  g20474(.dina(n6493), .dinb(n10637), .dout(n20733));
  jor  g20475(.dina(n6495), .dinb(n10964), .dout(n20734));
  jand g20476(.dina(n20734), .dinb(n20733), .dout(n20735));
  jand g20477(.dina(n20735), .dinb(n20732), .dout(n20736));
  jand g20478(.dina(n20736), .dinb(n20731), .dout(n20737));
  jxor g20479(.dina(n20737), .dinb(a47 ), .dout(n20738));
  jxor g20480(.dina(n20738), .dinb(n20730), .dout(n20739));
  jor  g20481(.dina(n20636), .dinb(n20558), .dout(n20740));
  jand g20482(.dina(n20636), .dinb(n20558), .dout(n20741));
  jor  g20483(.dina(n20741), .dinb(n20555), .dout(n20742));
  jand g20484(.dina(n20742), .dinb(n20740), .dout(n20743));
  jxor g20485(.dina(n20743), .dinb(n20739), .dout(n20744));
  jand g20486(.dina(n20545), .dinb(n20541), .dout(n20745));
  jand g20487(.dina(n20638), .dinb(n20546), .dout(n20746));
  jor  g20488(.dina(n20746), .dinb(n20745), .dout(n20747));
  jxor g20489(.dina(n20747), .dinb(n20744), .dout(n20748));
  jxor g20490(.dina(n20748), .dinb(n20651), .dout(f108 ));
  jor  g20491(.dina(n20738), .dinb(n20730), .dout(n20750));
  jand g20492(.dina(n20743), .dinb(n20739), .dout(n20751));
  jnot g20493(.din(n20751), .dout(n20752));
  jand g20494(.dina(n20752), .dinb(n20750), .dout(n20753));
  jnot g20495(.din(n20753), .dout(n20754));
  jand g20496(.dina(n20723), .dinb(n20660), .dout(n20755));
  jand g20497(.dina(n20728), .dinb(n20724), .dout(n20756));
  jor  g20498(.dina(n20756), .dinb(n20755), .dout(n20757));
  jnot g20499(.din(n20757), .dout(n20758));
  jor  g20500(.dina(n10978), .dinb(n6490), .dout(n20759));
  jor  g20501(.dina(n6262), .dinb(n10637), .dout(n20760));
  jor  g20502(.dina(n6493), .dinb(n10964), .dout(n20761));
  jand g20503(.dina(n20761), .dinb(n20760), .dout(n20762));
  jand g20504(.dina(n20762), .dinb(n20759), .dout(n20763));
  jxor g20505(.dina(n20763), .dinb(a47 ), .dout(n20764));
  jxor g20506(.dina(n20764), .dinb(n20758), .dout(n20765));
  jor  g20507(.dina(n10311), .dinb(n7266), .dout(n20766));
  jor  g20508(.dina(n7021), .dinb(n9413), .dout(n20767));
  jor  g20509(.dina(n7269), .dinb(n9725), .dout(n20768));
  jor  g20510(.dina(n7271), .dinb(n10314), .dout(n20769));
  jand g20511(.dina(n20769), .dinb(n20768), .dout(n20770));
  jand g20512(.dina(n20770), .dinb(n20767), .dout(n20771));
  jand g20513(.dina(n20771), .dinb(n20766), .dout(n20772));
  jxor g20514(.dina(n20772), .dinb(a50 ), .dout(n20773));
  jnot g20515(.din(n20773), .dout(n20774));
  jand g20516(.dina(n20721), .dinb(n20672), .dout(n20775));
  jand g20517(.dina(n20722), .dinb(n20663), .dout(n20776));
  jor  g20518(.dina(n20776), .dinb(n20775), .dout(n20777));
  jor  g20519(.dina(n9387), .dinb(n8125), .dout(n20778));
  jor  g20520(.dina(n7846), .dinb(n8789), .dout(n20779));
  jor  g20521(.dina(n8128), .dinb(n8809), .dout(n20780));
  jor  g20522(.dina(n8130), .dinb(n9390), .dout(n20781));
  jand g20523(.dina(n20781), .dinb(n20780), .dout(n20782));
  jand g20524(.dina(n20782), .dinb(n20779), .dout(n20783));
  jand g20525(.dina(n20783), .dinb(n20778), .dout(n20784));
  jxor g20526(.dina(n20784), .dinb(a53 ), .dout(n20785));
  jnot g20527(.din(n20785), .dout(n20786));
  jand g20528(.dina(n20719), .dinb(n20684), .dout(n20787));
  jand g20529(.dina(n20720), .dinb(n20675), .dout(n20788));
  jor  g20530(.dina(n20788), .dinb(n20787), .dout(n20789));
  jand g20531(.dina(n20717), .dinb(n20696), .dout(n20790));
  jand g20532(.dina(n20718), .dinb(n20687), .dout(n20791));
  jor  g20533(.dina(n20791), .dinb(n20790), .dout(n20792));
  jor  g20534(.dina(n9891), .dinb(n7408), .dout(n20793));
  jor  g20535(.dina(n9593), .dinb(n7129), .dout(n20794));
  jor  g20536(.dina(n9894), .dinb(n7149), .dout(n20795));
  jor  g20537(.dina(n9896), .dinb(n7411), .dout(n20796));
  jand g20538(.dina(n20796), .dinb(n20795), .dout(n20797));
  jand g20539(.dina(n20797), .dinb(n20794), .dout(n20798));
  jand g20540(.dina(n20798), .dinb(n20793), .dout(n20799));
  jxor g20541(.dina(n20799), .dinb(a59 ), .dout(n20800));
  jnot g20542(.din(n20800), .dout(n20801));
  jand g20543(.dina(n20715), .dinb(n20710), .dout(n20802));
  jand g20544(.dina(n20716), .dinb(n20705), .dout(n20803));
  jor  g20545(.dina(n20803), .dinb(n20802), .dout(n20804));
  jand g20546(.dina(n20713), .dinb(n20536), .dout(n20805));
  jor  g20547(.dina(n20713), .dinb(n20536), .dout(n20806));
  jand g20548(.dina(n20806), .dinb(n20485), .dout(n20807));
  jor  g20549(.dina(n20807), .dinb(n20805), .dout(n20808));
  jand g20550(.dina(n10801), .dinb(b46 ), .dout(n20809));
  jand g20551(.dina(n11107), .dinb(b45 ), .dout(n20810));
  jor  g20552(.dina(n20810), .dinb(n20809), .dout(n20811));
  jnot g20553(.din(n20811), .dout(n20812));
  jxor g20554(.dina(n20812), .dinb(n20808), .dout(n20813));
  jnot g20555(.din(n20813), .dout(n20814));
  jor  g20556(.dina(n10806), .dinb(n6864), .dout(n20815));
  jor  g20557(.dina(n10485), .dinb(n6352), .dout(n20816));
  jor  g20558(.dina(n10809), .dinb(n6372), .dout(n20817));
  jor  g20559(.dina(n10811), .dinb(n6867), .dout(n20818));
  jand g20560(.dina(n20818), .dinb(n20817), .dout(n20819));
  jand g20561(.dina(n20819), .dinb(n20816), .dout(n20820));
  jand g20562(.dina(n20820), .dinb(n20815), .dout(n20821));
  jxor g20563(.dina(n20821), .dinb(a62 ), .dout(n20822));
  jxor g20564(.dina(n20822), .dinb(n20814), .dout(n20823));
  jxor g20565(.dina(n20823), .dinb(n20804), .dout(n20824));
  jxor g20566(.dina(n20824), .dinb(n20801), .dout(n20825));
  jxor g20567(.dina(n20825), .dinb(n20792), .dout(n20826));
  jor  g20568(.dina(n8978), .dinb(n8228), .dout(n20827));
  jor  g20569(.dina(n8677), .dinb(n7683), .dout(n20828));
  jor  g20570(.dina(n8981), .dinb(n7960), .dout(n20829));
  jor  g20571(.dina(n8983), .dinb(n8231), .dout(n20830));
  jand g20572(.dina(n20830), .dinb(n20829), .dout(n20831));
  jand g20573(.dina(n20831), .dinb(n20828), .dout(n20832));
  jand g20574(.dina(n20832), .dinb(n20827), .dout(n20833));
  jxor g20575(.dina(n20833), .dinb(a56 ), .dout(n20834));
  jnot g20576(.din(n20834), .dout(n20835));
  jxor g20577(.dina(n20835), .dinb(n20826), .dout(n20836));
  jxor g20578(.dina(n20836), .dinb(n20789), .dout(n20837));
  jxor g20579(.dina(n20837), .dinb(n20786), .dout(n20838));
  jxor g20580(.dina(n20838), .dinb(n20777), .dout(n20839));
  jxor g20581(.dina(n20839), .dinb(n20774), .dout(n20840));
  jxor g20582(.dina(n20840), .dinb(n20765), .dout(n20841));
  jxor g20583(.dina(n20841), .dinb(n20754), .dout(n20842));
  jand g20584(.dina(n20747), .dinb(n20744), .dout(n20843));
  jand g20585(.dina(n20748), .dinb(n20651), .dout(n20844));
  jor  g20586(.dina(n20844), .dinb(n20843), .dout(n20845));
  jxor g20587(.dina(n20845), .dinb(n20842), .dout(f109 ));
  jnot g20588(.din(a47 ), .dout(n20847));
  jand g20589(.dina(n11296), .dinb(n5977), .dout(n20848));
  jor  g20590(.dina(n20848), .dinb(n6263), .dout(n20849));
  jand g20591(.dina(n20849), .dinb(b63 ), .dout(n20850));
  jxor g20592(.dina(n20850), .dinb(n20847), .dout(n20851));
  jnot g20593(.din(n20851), .dout(n20852));
  jor  g20594(.dina(n20838), .dinb(n20777), .dout(n20853));
  jand g20595(.dina(n20838), .dinb(n20777), .dout(n20854));
  jor  g20596(.dina(n20854), .dinb(n20774), .dout(n20855));
  jand g20597(.dina(n20855), .dinb(n20853), .dout(n20856));
  jxor g20598(.dina(n20856), .dinb(n20852), .dout(n20857));
  jor  g20599(.dina(n10634), .dinb(n7266), .dout(n20858));
  jor  g20600(.dina(n7021), .dinb(n9725), .dout(n20859));
  jor  g20601(.dina(n7269), .dinb(n10314), .dout(n20860));
  jor  g20602(.dina(n7271), .dinb(n10637), .dout(n20861));
  jand g20603(.dina(n20861), .dinb(n20860), .dout(n20862));
  jand g20604(.dina(n20862), .dinb(n20859), .dout(n20863));
  jand g20605(.dina(n20863), .dinb(n20858), .dout(n20864));
  jxor g20606(.dina(n20864), .dinb(a50 ), .dout(n20865));
  jnot g20607(.din(n20865), .dout(n20866));
  jand g20608(.dina(n20836), .dinb(n20789), .dout(n20867));
  jand g20609(.dina(n20837), .dinb(n20786), .dout(n20868));
  jor  g20610(.dina(n20868), .dinb(n20867), .dout(n20869));
  jor  g20611(.dina(n8786), .dinb(n8978), .dout(n20870));
  jor  g20612(.dina(n8677), .dinb(n7960), .dout(n20871));
  jor  g20613(.dina(n8981), .dinb(n8231), .dout(n20872));
  jor  g20614(.dina(n8983), .dinb(n8789), .dout(n20873));
  jand g20615(.dina(n20873), .dinb(n20872), .dout(n20874));
  jand g20616(.dina(n20874), .dinb(n20871), .dout(n20875));
  jand g20617(.dina(n20875), .dinb(n20870), .dout(n20876));
  jxor g20618(.dina(n20876), .dinb(a56 ), .dout(n20877));
  jnot g20619(.din(n20877), .dout(n20878));
  jand g20620(.dina(n20823), .dinb(n20804), .dout(n20879));
  jand g20621(.dina(n20824), .dinb(n20801), .dout(n20880));
  jor  g20622(.dina(n20880), .dinb(n20879), .dout(n20881));
  jor  g20623(.dina(n9891), .dinb(n7680), .dout(n20882));
  jor  g20624(.dina(n9593), .dinb(n7149), .dout(n20883));
  jor  g20625(.dina(n9894), .dinb(n7411), .dout(n20884));
  jor  g20626(.dina(n9896), .dinb(n7683), .dout(n20885));
  jand g20627(.dina(n20885), .dinb(n20884), .dout(n20886));
  jand g20628(.dina(n20886), .dinb(n20883), .dout(n20887));
  jand g20629(.dina(n20887), .dinb(n20882), .dout(n20888));
  jxor g20630(.dina(n20888), .dinb(a59 ), .dout(n20889));
  jnot g20631(.din(n20889), .dout(n20890));
  jor  g20632(.dina(n10806), .dinb(n7126), .dout(n20891));
  jor  g20633(.dina(n10485), .dinb(n6372), .dout(n20892));
  jor  g20634(.dina(n10809), .dinb(n6867), .dout(n20893));
  jor  g20635(.dina(n10811), .dinb(n7129), .dout(n20894));
  jand g20636(.dina(n20894), .dinb(n20893), .dout(n20895));
  jand g20637(.dina(n20895), .dinb(n20892), .dout(n20896));
  jand g20638(.dina(n20896), .dinb(n20891), .dout(n20897));
  jxor g20639(.dina(n20897), .dinb(a62 ), .dout(n20898));
  jnot g20640(.din(n20898), .dout(n20899));
  jand g20641(.dina(n20812), .dinb(n20808), .dout(n20900));
  jnot g20642(.din(n20900), .dout(n20901));
  jor  g20643(.dina(n20822), .dinb(n20814), .dout(n20902));
  jand g20644(.dina(n20902), .dinb(n20901), .dout(n20903));
  jnot g20645(.din(n20903), .dout(n20904));
  jand g20646(.dina(n10801), .dinb(b47 ), .dout(n20905));
  jand g20647(.dina(n11107), .dinb(b46 ), .dout(n20906));
  jor  g20648(.dina(n20906), .dinb(n20905), .dout(n20907));
  jnot g20649(.din(n20907), .dout(n20908));
  jxor g20650(.dina(n20908), .dinb(n20811), .dout(n20909));
  jxor g20651(.dina(n20909), .dinb(n20904), .dout(n20910));
  jxor g20652(.dina(n20910), .dinb(n20899), .dout(n20911));
  jxor g20653(.dina(n20911), .dinb(n20890), .dout(n20912));
  jxor g20654(.dina(n20912), .dinb(n20881), .dout(n20913));
  jxor g20655(.dina(n20913), .dinb(n20878), .dout(n20914));
  jor  g20656(.dina(n20825), .dinb(n20792), .dout(n20915));
  jand g20657(.dina(n20825), .dinb(n20792), .dout(n20916));
  jor  g20658(.dina(n20835), .dinb(n20916), .dout(n20917));
  jand g20659(.dina(n20917), .dinb(n20915), .dout(n20918));
  jxor g20660(.dina(n20918), .dinb(n20914), .dout(n20919));
  jor  g20661(.dina(n9410), .dinb(n8125), .dout(n20920));
  jor  g20662(.dina(n7846), .dinb(n8809), .dout(n20921));
  jor  g20663(.dina(n8128), .dinb(n9390), .dout(n20922));
  jor  g20664(.dina(n8130), .dinb(n9413), .dout(n20923));
  jand g20665(.dina(n20923), .dinb(n20922), .dout(n20924));
  jand g20666(.dina(n20924), .dinb(n20921), .dout(n20925));
  jand g20667(.dina(n20925), .dinb(n20920), .dout(n20926));
  jxor g20668(.dina(n20926), .dinb(a53 ), .dout(n20927));
  jnot g20669(.din(n20927), .dout(n20928));
  jxor g20670(.dina(n20928), .dinb(n20919), .dout(n20929));
  jxor g20671(.dina(n20929), .dinb(n20869), .dout(n20930));
  jxor g20672(.dina(n20930), .dinb(n20866), .dout(n20931));
  jxor g20673(.dina(n20931), .dinb(n20857), .dout(n20932));
  jand g20674(.dina(n20764), .dinb(n20758), .dout(n20933));
  jnot g20675(.din(n20933), .dout(n20934));
  jnot g20676(.din(n20764), .dout(n20935));
  jand g20677(.dina(n20935), .dinb(n20757), .dout(n20936));
  jor  g20678(.dina(n20840), .dinb(n20936), .dout(n20937));
  jand g20679(.dina(n20937), .dinb(n20934), .dout(n20938));
  jxor g20680(.dina(n20938), .dinb(n20932), .dout(n20939));
  jand g20681(.dina(n20841), .dinb(n20754), .dout(n20940));
  jand g20682(.dina(n20845), .dinb(n20842), .dout(n20941));
  jor  g20683(.dina(n20941), .dinb(n20940), .dout(n20942));
  jxor g20684(.dina(n20942), .dinb(n20939), .dout(f110 ));
  jor  g20685(.dina(n9722), .dinb(n8125), .dout(n20944));
  jor  g20686(.dina(n7846), .dinb(n9390), .dout(n20945));
  jor  g20687(.dina(n8128), .dinb(n9413), .dout(n20946));
  jor  g20688(.dina(n8130), .dinb(n9725), .dout(n20947));
  jand g20689(.dina(n20947), .dinb(n20946), .dout(n20948));
  jand g20690(.dina(n20948), .dinb(n20945), .dout(n20949));
  jand g20691(.dina(n20949), .dinb(n20944), .dout(n20950));
  jxor g20692(.dina(n20950), .dinb(a53 ), .dout(n20951));
  jnot g20693(.din(n20951), .dout(n20952));
  jand g20694(.dina(n20912), .dinb(n20881), .dout(n20953));
  jand g20695(.dina(n20913), .dinb(n20878), .dout(n20954));
  jor  g20696(.dina(n20954), .dinb(n20953), .dout(n20955));
  jor  g20697(.dina(n8806), .dinb(n8978), .dout(n20956));
  jor  g20698(.dina(n8677), .dinb(n8231), .dout(n20957));
  jor  g20699(.dina(n8981), .dinb(n8789), .dout(n20958));
  jor  g20700(.dina(n8983), .dinb(n8809), .dout(n20959));
  jand g20701(.dina(n20959), .dinb(n20958), .dout(n20960));
  jand g20702(.dina(n20960), .dinb(n20957), .dout(n20961));
  jand g20703(.dina(n20961), .dinb(n20956), .dout(n20962));
  jxor g20704(.dina(n20962), .dinb(a56 ), .dout(n20963));
  jnot g20705(.din(n20963), .dout(n20964));
  jand g20706(.dina(n20910), .dinb(n20899), .dout(n20965));
  jand g20707(.dina(n20911), .dinb(n20890), .dout(n20966));
  jor  g20708(.dina(n20966), .dinb(n20965), .dout(n20967));
  jor  g20709(.dina(n9891), .dinb(n7957), .dout(n20968));
  jor  g20710(.dina(n9593), .dinb(n7411), .dout(n20969));
  jor  g20711(.dina(n9894), .dinb(n7683), .dout(n20970));
  jor  g20712(.dina(n9896), .dinb(n7960), .dout(n20971));
  jand g20713(.dina(n20971), .dinb(n20970), .dout(n20972));
  jand g20714(.dina(n20972), .dinb(n20969), .dout(n20973));
  jand g20715(.dina(n20973), .dinb(n20968), .dout(n20974));
  jxor g20716(.dina(n20974), .dinb(a59 ), .dout(n20975));
  jnot g20717(.din(n20975), .dout(n20976));
  jand g20718(.dina(n20908), .dinb(n20811), .dout(n20977));
  jand g20719(.dina(n20909), .dinb(n20904), .dout(n20978));
  jor  g20720(.dina(n20978), .dinb(n20977), .dout(n20979));
  jor  g20721(.dina(n10806), .dinb(n7146), .dout(n20980));
  jor  g20722(.dina(n10485), .dinb(n6867), .dout(n20981));
  jor  g20723(.dina(n10809), .dinb(n7129), .dout(n20982));
  jor  g20724(.dina(n10811), .dinb(n7149), .dout(n20983));
  jand g20725(.dina(n20983), .dinb(n20982), .dout(n20984));
  jand g20726(.dina(n20984), .dinb(n20981), .dout(n20985));
  jand g20727(.dina(n20985), .dinb(n20980), .dout(n20986));
  jxor g20728(.dina(n20986), .dinb(a62 ), .dout(n20987));
  jnot g20729(.din(n20987), .dout(n20988));
  jxor g20730(.dina(n20907), .dinb(n20847), .dout(n20989));
  jand g20731(.dina(n10801), .dinb(b48 ), .dout(n20990));
  jand g20732(.dina(n11107), .dinb(b47 ), .dout(n20991));
  jor  g20733(.dina(n20991), .dinb(n20990), .dout(n20992));
  jxor g20734(.dina(n20992), .dinb(n20989), .dout(n20993));
  jxor g20735(.dina(n20993), .dinb(n20988), .dout(n20994));
  jxor g20736(.dina(n20994), .dinb(n20979), .dout(n20995));
  jxor g20737(.dina(n20995), .dinb(n20976), .dout(n20996));
  jxor g20738(.dina(n20996), .dinb(n20967), .dout(n20997));
  jxor g20739(.dina(n20997), .dinb(n20964), .dout(n20998));
  jxor g20740(.dina(n20998), .dinb(n20955), .dout(n20999));
  jxor g20741(.dina(n20999), .dinb(n20952), .dout(n21000));
  jor  g20742(.dina(n20918), .dinb(n20914), .dout(n21001));
  jand g20743(.dina(n20918), .dinb(n20914), .dout(n21002));
  jor  g20744(.dina(n20928), .dinb(n21002), .dout(n21003));
  jand g20745(.dina(n21003), .dinb(n21001), .dout(n21004));
  jxor g20746(.dina(n21004), .dinb(n21000), .dout(n21005));
  jnot g20747(.din(n21005), .dout(n21006));
  jor  g20748(.dina(n10961), .dinb(n7266), .dout(n21007));
  jor  g20749(.dina(n7021), .dinb(n10314), .dout(n21008));
  jor  g20750(.dina(n7269), .dinb(n10637), .dout(n21009));
  jor  g20751(.dina(n7271), .dinb(n10964), .dout(n21010));
  jand g20752(.dina(n21010), .dinb(n21009), .dout(n21011));
  jand g20753(.dina(n21011), .dinb(n21008), .dout(n21012));
  jand g20754(.dina(n21012), .dinb(n21007), .dout(n21013));
  jxor g20755(.dina(n21013), .dinb(a50 ), .dout(n21014));
  jxor g20756(.dina(n21014), .dinb(n21006), .dout(n21015));
  jor  g20757(.dina(n20929), .dinb(n20869), .dout(n21016));
  jand g20758(.dina(n20929), .dinb(n20869), .dout(n21017));
  jor  g20759(.dina(n21017), .dinb(n20866), .dout(n21018));
  jand g20760(.dina(n21018), .dinb(n21016), .dout(n21019));
  jxor g20761(.dina(n21019), .dinb(n21015), .dout(n21020));
  jor  g20762(.dina(n20856), .dinb(n20852), .dout(n21021));
  jand g20763(.dina(n20856), .dinb(n20852), .dout(n21022));
  jor  g20764(.dina(n20931), .dinb(n21022), .dout(n21023));
  jand g20765(.dina(n21023), .dinb(n21021), .dout(n21024));
  jxor g20766(.dina(n21024), .dinb(n21020), .dout(n21025));
  jand g20767(.dina(n20938), .dinb(n20932), .dout(n21026));
  jand g20768(.dina(n20942), .dinb(n20939), .dout(n21027));
  jor  g20769(.dina(n21027), .dinb(n21026), .dout(n21028));
  jxor g20770(.dina(n21028), .dinb(n21025), .dout(f111 ));
  jor  g20771(.dina(n21014), .dinb(n21006), .dout(n21030));
  jand g20772(.dina(n21019), .dinb(n21015), .dout(n21031));
  jnot g20773(.din(n21031), .dout(n21032));
  jand g20774(.dina(n21032), .dinb(n21030), .dout(n21033));
  jnot g20775(.din(n21033), .dout(n21034));
  jand g20776(.dina(n20999), .dinb(n20952), .dout(n21035));
  jand g20777(.dina(n21004), .dinb(n21000), .dout(n21036));
  jor  g20778(.dina(n21036), .dinb(n21035), .dout(n21037));
  jor  g20779(.dina(n10311), .dinb(n8125), .dout(n21038));
  jor  g20780(.dina(n7846), .dinb(n9413), .dout(n21039));
  jor  g20781(.dina(n8128), .dinb(n9725), .dout(n21040));
  jor  g20782(.dina(n8130), .dinb(n10314), .dout(n21041));
  jand g20783(.dina(n21041), .dinb(n21040), .dout(n21042));
  jand g20784(.dina(n21042), .dinb(n21039), .dout(n21043));
  jand g20785(.dina(n21043), .dinb(n21038), .dout(n21044));
  jxor g20786(.dina(n21044), .dinb(a53 ), .dout(n21045));
  jnot g20787(.din(n21045), .dout(n21046));
  jand g20788(.dina(n20997), .dinb(n20964), .dout(n21047));
  jand g20789(.dina(n20998), .dinb(n20955), .dout(n21048));
  jor  g20790(.dina(n21048), .dinb(n21047), .dout(n21049));
  jor  g20791(.dina(n9387), .dinb(n8978), .dout(n21050));
  jor  g20792(.dina(n8677), .dinb(n8789), .dout(n21051));
  jor  g20793(.dina(n8981), .dinb(n8809), .dout(n21052));
  jor  g20794(.dina(n8983), .dinb(n9390), .dout(n21053));
  jand g20795(.dina(n21053), .dinb(n21052), .dout(n21054));
  jand g20796(.dina(n21054), .dinb(n21051), .dout(n21055));
  jand g20797(.dina(n21055), .dinb(n21050), .dout(n21056));
  jxor g20798(.dina(n21056), .dinb(a56 ), .dout(n21057));
  jnot g20799(.din(n21057), .dout(n21058));
  jand g20800(.dina(n20995), .dinb(n20976), .dout(n21059));
  jand g20801(.dina(n20996), .dinb(n20967), .dout(n21060));
  jor  g20802(.dina(n21060), .dinb(n21059), .dout(n21061));
  jor  g20803(.dina(n9891), .dinb(n8228), .dout(n21062));
  jor  g20804(.dina(n9593), .dinb(n7683), .dout(n21063));
  jor  g20805(.dina(n9894), .dinb(n7960), .dout(n21064));
  jor  g20806(.dina(n9896), .dinb(n8231), .dout(n21065));
  jand g20807(.dina(n21065), .dinb(n21064), .dout(n21066));
  jand g20808(.dina(n21066), .dinb(n21063), .dout(n21067));
  jand g20809(.dina(n21067), .dinb(n21062), .dout(n21068));
  jxor g20810(.dina(n21068), .dinb(a59 ), .dout(n21069));
  jnot g20811(.din(n21069), .dout(n21070));
  jand g20812(.dina(n20993), .dinb(n20988), .dout(n21071));
  jand g20813(.dina(n20994), .dinb(n20979), .dout(n21072));
  jor  g20814(.dina(n21072), .dinb(n21071), .dout(n21073));
  jand g20815(.dina(n20907), .dinb(n20847), .dout(n21074));
  jand g20816(.dina(n20992), .dinb(n20989), .dout(n21075));
  jor  g20817(.dina(n21075), .dinb(n21074), .dout(n21076));
  jand g20818(.dina(n10801), .dinb(b49 ), .dout(n21077));
  jand g20819(.dina(n11107), .dinb(b48 ), .dout(n21078));
  jor  g20820(.dina(n21078), .dinb(n21077), .dout(n21079));
  jnot g20821(.din(n21079), .dout(n21080));
  jxor g20822(.dina(n21080), .dinb(n21076), .dout(n21081));
  jnot g20823(.din(n21081), .dout(n21082));
  jor  g20824(.dina(n10806), .dinb(n7408), .dout(n21083));
  jor  g20825(.dina(n10485), .dinb(n7129), .dout(n21084));
  jor  g20826(.dina(n10809), .dinb(n7149), .dout(n21085));
  jor  g20827(.dina(n10811), .dinb(n7411), .dout(n21086));
  jand g20828(.dina(n21086), .dinb(n21085), .dout(n21087));
  jand g20829(.dina(n21087), .dinb(n21084), .dout(n21088));
  jand g20830(.dina(n21088), .dinb(n21083), .dout(n21089));
  jxor g20831(.dina(n21089), .dinb(a62 ), .dout(n21090));
  jxor g20832(.dina(n21090), .dinb(n21082), .dout(n21091));
  jxor g20833(.dina(n21091), .dinb(n21073), .dout(n21092));
  jxor g20834(.dina(n21092), .dinb(n21070), .dout(n21093));
  jxor g20835(.dina(n21093), .dinb(n21061), .dout(n21094));
  jxor g20836(.dina(n21094), .dinb(n21058), .dout(n21095));
  jxor g20837(.dina(n21095), .dinb(n21049), .dout(n21096));
  jxor g20838(.dina(n21096), .dinb(n21046), .dout(n21097));
  jxor g20839(.dina(n21097), .dinb(n21037), .dout(n21098));
  jor  g20840(.dina(n10978), .dinb(n7266), .dout(n21099));
  jor  g20841(.dina(n7021), .dinb(n10637), .dout(n21100));
  jor  g20842(.dina(n7269), .dinb(n10964), .dout(n21101));
  jand g20843(.dina(n21101), .dinb(n21100), .dout(n21102));
  jand g20844(.dina(n21102), .dinb(n21099), .dout(n21103));
  jxor g20845(.dina(n21103), .dinb(a50 ), .dout(n21104));
  jnot g20846(.din(n21104), .dout(n21105));
  jxor g20847(.dina(n21105), .dinb(n21098), .dout(n21106));
  jxor g20848(.dina(n21106), .dinb(n21034), .dout(n21107));
  jand g20849(.dina(n21024), .dinb(n21020), .dout(n21108));
  jand g20850(.dina(n21028), .dinb(n21025), .dout(n21109));
  jor  g20851(.dina(n21109), .dinb(n21108), .dout(n21110));
  jxor g20852(.dina(n21110), .dinb(n21107), .dout(f112 ));
  jand g20853(.dina(n21095), .dinb(n21049), .dout(n21112));
  jand g20854(.dina(n21096), .dinb(n21046), .dout(n21113));
  jor  g20855(.dina(n21113), .dinb(n21112), .dout(n21114));
  jnot g20856(.din(n21114), .dout(n21115));
  jnot g20857(.din(a50 ), .dout(n21116));
  jand g20858(.dina(n11296), .dinb(n6728), .dout(n21117));
  jor  g20859(.dina(n21117), .dinb(n7022), .dout(n21118));
  jand g20860(.dina(n21118), .dinb(b63 ), .dout(n21119));
  jxor g20861(.dina(n21119), .dinb(n21116), .dout(n21120));
  jxor g20862(.dina(n21120), .dinb(n21115), .dout(n21121));
  jand g20863(.dina(n21093), .dinb(n21061), .dout(n21122));
  jand g20864(.dina(n21094), .dinb(n21058), .dout(n21123));
  jor  g20865(.dina(n21123), .dinb(n21122), .dout(n21124));
  jand g20866(.dina(n21091), .dinb(n21073), .dout(n21125));
  jand g20867(.dina(n21092), .dinb(n21070), .dout(n21126));
  jor  g20868(.dina(n21126), .dinb(n21125), .dout(n21127));
  jand g20869(.dina(n21080), .dinb(n21076), .dout(n21128));
  jnot g20870(.din(n21128), .dout(n21129));
  jor  g20871(.dina(n21090), .dinb(n21082), .dout(n21130));
  jand g20872(.dina(n21130), .dinb(n21129), .dout(n21131));
  jnot g20873(.din(n21131), .dout(n21132));
  jor  g20874(.dina(n10806), .dinb(n7680), .dout(n21133));
  jor  g20875(.dina(n10485), .dinb(n7149), .dout(n21134));
  jor  g20876(.dina(n10809), .dinb(n7411), .dout(n21135));
  jor  g20877(.dina(n10811), .dinb(n7683), .dout(n21136));
  jand g20878(.dina(n21136), .dinb(n21135), .dout(n21137));
  jand g20879(.dina(n21137), .dinb(n21134), .dout(n21138));
  jand g20880(.dina(n21138), .dinb(n21133), .dout(n21139));
  jxor g20881(.dina(n21139), .dinb(a62 ), .dout(n21140));
  jnot g20882(.din(n21140), .dout(n21141));
  jand g20883(.dina(n10801), .dinb(b50 ), .dout(n21142));
  jand g20884(.dina(n11107), .dinb(b49 ), .dout(n21143));
  jor  g20885(.dina(n21143), .dinb(n21142), .dout(n21144));
  jxor g20886(.dina(n21144), .dinb(n21080), .dout(n21145));
  jxor g20887(.dina(n21145), .dinb(n21141), .dout(n21146));
  jxor g20888(.dina(n21146), .dinb(n21132), .dout(n21147));
  jnot g20889(.din(n21147), .dout(n21148));
  jor  g20890(.dina(n9891), .dinb(n8786), .dout(n21149));
  jor  g20891(.dina(n9593), .dinb(n7960), .dout(n21150));
  jor  g20892(.dina(n9894), .dinb(n8231), .dout(n21151));
  jor  g20893(.dina(n9896), .dinb(n8789), .dout(n21152));
  jand g20894(.dina(n21152), .dinb(n21151), .dout(n21153));
  jand g20895(.dina(n21153), .dinb(n21150), .dout(n21154));
  jand g20896(.dina(n21154), .dinb(n21149), .dout(n21155));
  jxor g20897(.dina(n21155), .dinb(a59 ), .dout(n21156));
  jxor g20898(.dina(n21156), .dinb(n21148), .dout(n21157));
  jxor g20899(.dina(n21157), .dinb(n21127), .dout(n21158));
  jor  g20900(.dina(n9410), .dinb(n8978), .dout(n21159));
  jor  g20901(.dina(n8677), .dinb(n8809), .dout(n21160));
  jor  g20902(.dina(n8981), .dinb(n9390), .dout(n21161));
  jor  g20903(.dina(n8983), .dinb(n9413), .dout(n21162));
  jand g20904(.dina(n21162), .dinb(n21161), .dout(n21163));
  jand g20905(.dina(n21163), .dinb(n21160), .dout(n21164));
  jand g20906(.dina(n21164), .dinb(n21159), .dout(n21165));
  jxor g20907(.dina(n21165), .dinb(a56 ), .dout(n21166));
  jnot g20908(.din(n21166), .dout(n21167));
  jxor g20909(.dina(n21167), .dinb(n21158), .dout(n21168));
  jxor g20910(.dina(n21168), .dinb(n21124), .dout(n21169));
  jor  g20911(.dina(n10634), .dinb(n8125), .dout(n21170));
  jor  g20912(.dina(n7846), .dinb(n9725), .dout(n21171));
  jor  g20913(.dina(n8128), .dinb(n10314), .dout(n21172));
  jor  g20914(.dina(n8130), .dinb(n10637), .dout(n21173));
  jand g20915(.dina(n21173), .dinb(n21172), .dout(n21174));
  jand g20916(.dina(n21174), .dinb(n21171), .dout(n21175));
  jand g20917(.dina(n21175), .dinb(n21170), .dout(n21176));
  jxor g20918(.dina(n21176), .dinb(a53 ), .dout(n21177));
  jnot g20919(.din(n21177), .dout(n21178));
  jxor g20920(.dina(n21178), .dinb(n21169), .dout(n21179));
  jxor g20921(.dina(n21179), .dinb(n21121), .dout(n21180));
  jor  g20922(.dina(n21097), .dinb(n21037), .dout(n21181));
  jand g20923(.dina(n21097), .dinb(n21037), .dout(n21182));
  jor  g20924(.dina(n21105), .dinb(n21182), .dout(n21183));
  jand g20925(.dina(n21183), .dinb(n21181), .dout(n21184));
  jxor g20926(.dina(n21184), .dinb(n21180), .dout(n21185));
  jand g20927(.dina(n21106), .dinb(n21034), .dout(n21186));
  jand g20928(.dina(n21110), .dinb(n21107), .dout(n21187));
  jor  g20929(.dina(n21187), .dinb(n21186), .dout(n21188));
  jxor g20930(.dina(n21188), .dinb(n21185), .dout(f113 ));
  jor  g20931(.dina(n9722), .dinb(n8978), .dout(n21190));
  jor  g20932(.dina(n8677), .dinb(n9390), .dout(n21191));
  jor  g20933(.dina(n8981), .dinb(n9413), .dout(n21192));
  jor  g20934(.dina(n8983), .dinb(n9725), .dout(n21193));
  jand g20935(.dina(n21193), .dinb(n21192), .dout(n21194));
  jand g20936(.dina(n21194), .dinb(n21191), .dout(n21195));
  jand g20937(.dina(n21195), .dinb(n21190), .dout(n21196));
  jxor g20938(.dina(n21196), .dinb(a56 ), .dout(n21197));
  jnot g20939(.din(n21197), .dout(n21198));
  jand g20940(.dina(n21146), .dinb(n21132), .dout(n21199));
  jnot g20941(.din(n21199), .dout(n21200));
  jor  g20942(.dina(n21156), .dinb(n21148), .dout(n21201));
  jand g20943(.dina(n21201), .dinb(n21200), .dout(n21202));
  jnot g20944(.din(n21202), .dout(n21203));
  jor  g20945(.dina(n9891), .dinb(n8806), .dout(n21204));
  jor  g20946(.dina(n9593), .dinb(n8231), .dout(n21205));
  jor  g20947(.dina(n9894), .dinb(n8789), .dout(n21206));
  jor  g20948(.dina(n9896), .dinb(n8809), .dout(n21207));
  jand g20949(.dina(n21207), .dinb(n21206), .dout(n21208));
  jand g20950(.dina(n21208), .dinb(n21205), .dout(n21209));
  jand g20951(.dina(n21209), .dinb(n21204), .dout(n21210));
  jxor g20952(.dina(n21210), .dinb(a59 ), .dout(n21211));
  jnot g20953(.din(n21211), .dout(n21212));
  jor  g20954(.dina(n10806), .dinb(n7957), .dout(n21213));
  jor  g20955(.dina(n10485), .dinb(n7411), .dout(n21214));
  jor  g20956(.dina(n10809), .dinb(n7683), .dout(n21215));
  jor  g20957(.dina(n10811), .dinb(n7960), .dout(n21216));
  jand g20958(.dina(n21216), .dinb(n21215), .dout(n21217));
  jand g20959(.dina(n21217), .dinb(n21214), .dout(n21218));
  jand g20960(.dina(n21218), .dinb(n21213), .dout(n21219));
  jxor g20961(.dina(n21219), .dinb(a62 ), .dout(n21220));
  jnot g20962(.din(n21220), .dout(n21221));
  jand g20963(.dina(n21144), .dinb(n21080), .dout(n21222));
  jand g20964(.dina(n21145), .dinb(n21141), .dout(n21223));
  jor  g20965(.dina(n21223), .dinb(n21222), .dout(n21224));
  jand g20966(.dina(n10801), .dinb(b51 ), .dout(n21225));
  jand g20967(.dina(n11107), .dinb(b50 ), .dout(n21226));
  jor  g20968(.dina(n21226), .dinb(n21225), .dout(n21227));
  jxor g20969(.dina(n21227), .dinb(n21116), .dout(n21228));
  jxor g20970(.dina(n21228), .dinb(n21079), .dout(n21229));
  jxor g20971(.dina(n21229), .dinb(n21224), .dout(n21230));
  jxor g20972(.dina(n21230), .dinb(n21221), .dout(n21231));
  jxor g20973(.dina(n21231), .dinb(n21212), .dout(n21232));
  jxor g20974(.dina(n21232), .dinb(n21203), .dout(n21233));
  jxor g20975(.dina(n21233), .dinb(n21198), .dout(n21234));
  jor  g20976(.dina(n21157), .dinb(n21127), .dout(n21235));
  jand g20977(.dina(n21157), .dinb(n21127), .dout(n21236));
  jor  g20978(.dina(n21167), .dinb(n21236), .dout(n21237));
  jand g20979(.dina(n21237), .dinb(n21235), .dout(n21238));
  jxor g20980(.dina(n21238), .dinb(n21234), .dout(n21239));
  jnot g20981(.din(n21239), .dout(n21240));
  jor  g20982(.dina(n10961), .dinb(n8125), .dout(n21241));
  jor  g20983(.dina(n7846), .dinb(n10314), .dout(n21242));
  jor  g20984(.dina(n8128), .dinb(n10637), .dout(n21243));
  jor  g20985(.dina(n8130), .dinb(n10964), .dout(n21244));
  jand g20986(.dina(n21244), .dinb(n21243), .dout(n21245));
  jand g20987(.dina(n21245), .dinb(n21242), .dout(n21246));
  jand g20988(.dina(n21246), .dinb(n21241), .dout(n21247));
  jxor g20989(.dina(n21247), .dinb(a53 ), .dout(n21248));
  jxor g20990(.dina(n21248), .dinb(n21240), .dout(n21249));
  jnot g20991(.din(n21124), .dout(n21250));
  jnot g20992(.din(n21168), .dout(n21251));
  jand g20993(.dina(n21251), .dinb(n21250), .dout(n21252));
  jnot g20994(.din(n21252), .dout(n21253));
  jand g20995(.dina(n21168), .dinb(n21124), .dout(n21254));
  jor  g20996(.dina(n21178), .dinb(n21254), .dout(n21255));
  jand g20997(.dina(n21255), .dinb(n21253), .dout(n21256));
  jxor g20998(.dina(n21256), .dinb(n21249), .dout(n21257));
  jand g20999(.dina(n21120), .dinb(n21115), .dout(n21258));
  jnot g21000(.din(n21258), .dout(n21259));
  jnot g21001(.din(n21120), .dout(n21260));
  jand g21002(.dina(n21260), .dinb(n21114), .dout(n21261));
  jor  g21003(.dina(n21179), .dinb(n21261), .dout(n21262));
  jand g21004(.dina(n21262), .dinb(n21259), .dout(n21263));
  jxor g21005(.dina(n21263), .dinb(n21257), .dout(n21264));
  jand g21006(.dina(n21184), .dinb(n21180), .dout(n21265));
  jand g21007(.dina(n21188), .dinb(n21185), .dout(n21266));
  jor  g21008(.dina(n21266), .dinb(n21265), .dout(n21267));
  jxor g21009(.dina(n21267), .dinb(n21264), .dout(f114 ));
  jor  g21010(.dina(n21248), .dinb(n21240), .dout(n21269));
  jand g21011(.dina(n21256), .dinb(n21249), .dout(n21270));
  jnot g21012(.din(n21270), .dout(n21271));
  jand g21013(.dina(n21271), .dinb(n21269), .dout(n21272));
  jnot g21014(.din(n21272), .dout(n21273));
  jand g21015(.dina(n21233), .dinb(n21198), .dout(n21274));
  jand g21016(.dina(n21238), .dinb(n21234), .dout(n21275));
  jor  g21017(.dina(n21275), .dinb(n21274), .dout(n21276));
  jor  g21018(.dina(n10311), .dinb(n8978), .dout(n21277));
  jor  g21019(.dina(n8677), .dinb(n9413), .dout(n21278));
  jor  g21020(.dina(n8981), .dinb(n9725), .dout(n21279));
  jor  g21021(.dina(n8983), .dinb(n10314), .dout(n21280));
  jand g21022(.dina(n21280), .dinb(n21279), .dout(n21281));
  jand g21023(.dina(n21281), .dinb(n21278), .dout(n21282));
  jand g21024(.dina(n21282), .dinb(n21277), .dout(n21283));
  jxor g21025(.dina(n21283), .dinb(a56 ), .dout(n21284));
  jnot g21026(.din(n21284), .dout(n21285));
  jand g21027(.dina(n21231), .dinb(n21212), .dout(n21286));
  jand g21028(.dina(n21232), .dinb(n21203), .dout(n21287));
  jor  g21029(.dina(n21287), .dinb(n21286), .dout(n21288));
  jor  g21030(.dina(n9387), .dinb(n9891), .dout(n21289));
  jor  g21031(.dina(n9593), .dinb(n8789), .dout(n21290));
  jor  g21032(.dina(n9894), .dinb(n8809), .dout(n21291));
  jor  g21033(.dina(n9896), .dinb(n9390), .dout(n21292));
  jand g21034(.dina(n21292), .dinb(n21291), .dout(n21293));
  jand g21035(.dina(n21293), .dinb(n21290), .dout(n21294));
  jand g21036(.dina(n21294), .dinb(n21289), .dout(n21295));
  jxor g21037(.dina(n21295), .dinb(a59 ), .dout(n21296));
  jnot g21038(.din(n21296), .dout(n21297));
  jand g21039(.dina(n21229), .dinb(n21224), .dout(n21298));
  jand g21040(.dina(n21230), .dinb(n21221), .dout(n21299));
  jor  g21041(.dina(n21299), .dinb(n21298), .dout(n21300));
  jand g21042(.dina(n21227), .dinb(n21116), .dout(n21301));
  jand g21043(.dina(n21228), .dinb(n21079), .dout(n21302));
  jor  g21044(.dina(n21302), .dinb(n21301), .dout(n21303));
  jand g21045(.dina(n10801), .dinb(b52 ), .dout(n21304));
  jand g21046(.dina(n11107), .dinb(b51 ), .dout(n21305));
  jor  g21047(.dina(n21305), .dinb(n21304), .dout(n21306));
  jnot g21048(.din(n21306), .dout(n21307));
  jxor g21049(.dina(n21307), .dinb(n21303), .dout(n21308));
  jnot g21050(.din(n21308), .dout(n21309));
  jor  g21051(.dina(n10806), .dinb(n8228), .dout(n21310));
  jor  g21052(.dina(n10485), .dinb(n7683), .dout(n21311));
  jor  g21053(.dina(n10809), .dinb(n7960), .dout(n21312));
  jor  g21054(.dina(n10811), .dinb(n8231), .dout(n21313));
  jand g21055(.dina(n21313), .dinb(n21312), .dout(n21314));
  jand g21056(.dina(n21314), .dinb(n21311), .dout(n21315));
  jand g21057(.dina(n21315), .dinb(n21310), .dout(n21316));
  jxor g21058(.dina(n21316), .dinb(a62 ), .dout(n21317));
  jxor g21059(.dina(n21317), .dinb(n21309), .dout(n21318));
  jxor g21060(.dina(n21318), .dinb(n21300), .dout(n21319));
  jxor g21061(.dina(n21319), .dinb(n21297), .dout(n21320));
  jxor g21062(.dina(n21320), .dinb(n21288), .dout(n21321));
  jxor g21063(.dina(n21321), .dinb(n21285), .dout(n21322));
  jxor g21064(.dina(n21322), .dinb(n21276), .dout(n21323));
  jor  g21065(.dina(n10978), .dinb(n8125), .dout(n21324));
  jor  g21066(.dina(n7846), .dinb(n10637), .dout(n21325));
  jor  g21067(.dina(n8128), .dinb(n10964), .dout(n21326));
  jand g21068(.dina(n21326), .dinb(n21325), .dout(n21327));
  jand g21069(.dina(n21327), .dinb(n21324), .dout(n21328));
  jxor g21070(.dina(n21328), .dinb(a53 ), .dout(n21329));
  jnot g21071(.din(n21329), .dout(n21330));
  jxor g21072(.dina(n21330), .dinb(n21323), .dout(n21331));
  jxor g21073(.dina(n21331), .dinb(n21273), .dout(n21332));
  jand g21074(.dina(n21263), .dinb(n21257), .dout(n21333));
  jand g21075(.dina(n21267), .dinb(n21264), .dout(n21334));
  jor  g21076(.dina(n21334), .dinb(n21333), .dout(n21335));
  jxor g21077(.dina(n21335), .dinb(n21332), .dout(f115 ));
  jand g21078(.dina(n21320), .dinb(n21288), .dout(n21337));
  jand g21079(.dina(n21321), .dinb(n21285), .dout(n21338));
  jor  g21080(.dina(n21338), .dinb(n21337), .dout(n21339));
  jnot g21081(.din(n21339), .dout(n21340));
  jnot g21082(.din(a53 ), .dout(n21341));
  jand g21083(.dina(n11296), .dinb(n7521), .dout(n21342));
  jor  g21084(.dina(n21342), .dinb(n7847), .dout(n21343));
  jand g21085(.dina(n21343), .dinb(b63 ), .dout(n21344));
  jxor g21086(.dina(n21344), .dinb(n21341), .dout(n21345));
  jxor g21087(.dina(n21345), .dinb(n21340), .dout(n21346));
  jand g21088(.dina(n21318), .dinb(n21300), .dout(n21347));
  jand g21089(.dina(n21319), .dinb(n21297), .dout(n21348));
  jor  g21090(.dina(n21348), .dinb(n21347), .dout(n21349));
  jor  g21091(.dina(n9410), .dinb(n9891), .dout(n21350));
  jor  g21092(.dina(n9593), .dinb(n8809), .dout(n21351));
  jor  g21093(.dina(n9894), .dinb(n9390), .dout(n21352));
  jor  g21094(.dina(n9896), .dinb(n9413), .dout(n21353));
  jand g21095(.dina(n21353), .dinb(n21352), .dout(n21354));
  jand g21096(.dina(n21354), .dinb(n21351), .dout(n21355));
  jand g21097(.dina(n21355), .dinb(n21350), .dout(n21356));
  jxor g21098(.dina(n21356), .dinb(a59 ), .dout(n21357));
  jnot g21099(.din(n21357), .dout(n21358));
  jor  g21100(.dina(n10806), .dinb(n8786), .dout(n21359));
  jor  g21101(.dina(n10485), .dinb(n7960), .dout(n21360));
  jor  g21102(.dina(n10809), .dinb(n8231), .dout(n21361));
  jor  g21103(.dina(n10811), .dinb(n8789), .dout(n21362));
  jand g21104(.dina(n21362), .dinb(n21361), .dout(n21363));
  jand g21105(.dina(n21363), .dinb(n21360), .dout(n21364));
  jand g21106(.dina(n21364), .dinb(n21359), .dout(n21365));
  jxor g21107(.dina(n21365), .dinb(a62 ), .dout(n21366));
  jnot g21108(.din(n21366), .dout(n21367));
  jand g21109(.dina(n21307), .dinb(n21303), .dout(n21368));
  jnot g21110(.din(n21368), .dout(n21369));
  jor  g21111(.dina(n21317), .dinb(n21309), .dout(n21370));
  jand g21112(.dina(n21370), .dinb(n21369), .dout(n21371));
  jnot g21113(.din(n21371), .dout(n21372));
  jand g21114(.dina(n10801), .dinb(b53 ), .dout(n21373));
  jand g21115(.dina(n11107), .dinb(b52 ), .dout(n21374));
  jor  g21116(.dina(n21374), .dinb(n21373), .dout(n21375));
  jxor g21117(.dina(n21375), .dinb(n21307), .dout(n21376));
  jxor g21118(.dina(n21376), .dinb(n21372), .dout(n21377));
  jxor g21119(.dina(n21377), .dinb(n21367), .dout(n21378));
  jxor g21120(.dina(n21378), .dinb(n21358), .dout(n21379));
  jxor g21121(.dina(n21379), .dinb(n21349), .dout(n21380));
  jor  g21122(.dina(n10634), .dinb(n8978), .dout(n21381));
  jor  g21123(.dina(n8677), .dinb(n9725), .dout(n21382));
  jor  g21124(.dina(n8981), .dinb(n10314), .dout(n21383));
  jor  g21125(.dina(n8983), .dinb(n10637), .dout(n21384));
  jand g21126(.dina(n21384), .dinb(n21383), .dout(n21385));
  jand g21127(.dina(n21385), .dinb(n21382), .dout(n21386));
  jand g21128(.dina(n21386), .dinb(n21381), .dout(n21387));
  jxor g21129(.dina(n21387), .dinb(a56 ), .dout(n21388));
  jnot g21130(.din(n21388), .dout(n21389));
  jxor g21131(.dina(n21389), .dinb(n21380), .dout(n21390));
  jxor g21132(.dina(n21390), .dinb(n21346), .dout(n21391));
  jor  g21133(.dina(n21322), .dinb(n21276), .dout(n21392));
  jand g21134(.dina(n21322), .dinb(n21276), .dout(n21393));
  jor  g21135(.dina(n21330), .dinb(n21393), .dout(n21394));
  jand g21136(.dina(n21394), .dinb(n21392), .dout(n21395));
  jxor g21137(.dina(n21395), .dinb(n21391), .dout(n21396));
  jand g21138(.dina(n21331), .dinb(n21273), .dout(n21397));
  jand g21139(.dina(n21335), .dinb(n21332), .dout(n21398));
  jor  g21140(.dina(n21398), .dinb(n21397), .dout(n21399));
  jxor g21141(.dina(n21399), .dinb(n21396), .dout(f116 ));
  jand g21142(.dina(n21395), .dinb(n21391), .dout(n21401));
  jand g21143(.dina(n21399), .dinb(n21396), .dout(n21402));
  jor  g21144(.dina(n21402), .dinb(n21401), .dout(n21403));
  jor  g21145(.dina(n10961), .dinb(n8978), .dout(n21404));
  jor  g21146(.dina(n8677), .dinb(n10314), .dout(n21405));
  jor  g21147(.dina(n8981), .dinb(n10637), .dout(n21406));
  jor  g21148(.dina(n8983), .dinb(n10964), .dout(n21407));
  jand g21149(.dina(n21407), .dinb(n21406), .dout(n21408));
  jand g21150(.dina(n21408), .dinb(n21405), .dout(n21409));
  jand g21151(.dina(n21409), .dinb(n21404), .dout(n21410));
  jxor g21152(.dina(n21410), .dinb(a56 ), .dout(n21411));
  jnot g21153(.din(n21411), .dout(n21412));
  jnot g21154(.din(n21349), .dout(n21413));
  jnot g21155(.din(n21379), .dout(n21414));
  jand g21156(.dina(n21414), .dinb(n21413), .dout(n21415));
  jnot g21157(.din(n21415), .dout(n21416));
  jand g21158(.dina(n21379), .dinb(n21349), .dout(n21417));
  jor  g21159(.dina(n21389), .dinb(n21417), .dout(n21418));
  jand g21160(.dina(n21418), .dinb(n21416), .dout(n21419));
  jxor g21161(.dina(n21419), .dinb(n21412), .dout(n21420));
  jand g21162(.dina(n21377), .dinb(n21367), .dout(n21421));
  jand g21163(.dina(n21378), .dinb(n21358), .dout(n21422));
  jor  g21164(.dina(n21422), .dinb(n21421), .dout(n21423));
  jor  g21165(.dina(n9722), .dinb(n9891), .dout(n21424));
  jor  g21166(.dina(n9593), .dinb(n9390), .dout(n21425));
  jor  g21167(.dina(n9894), .dinb(n9413), .dout(n21426));
  jor  g21168(.dina(n9896), .dinb(n9725), .dout(n21427));
  jand g21169(.dina(n21427), .dinb(n21426), .dout(n21428));
  jand g21170(.dina(n21428), .dinb(n21425), .dout(n21429));
  jand g21171(.dina(n21429), .dinb(n21424), .dout(n21430));
  jxor g21172(.dina(n21430), .dinb(a59 ), .dout(n21431));
  jnot g21173(.din(n21431), .dout(n21432));
  jnot g21174(.din(n21375), .dout(n21433));
  jand g21175(.dina(n21433), .dinb(n21306), .dout(n21434));
  jand g21176(.dina(n21376), .dinb(n21372), .dout(n21435));
  jor  g21177(.dina(n21435), .dinb(n21434), .dout(n21436));
  jxor g21178(.dina(n21375), .dinb(n21341), .dout(n21437));
  jand g21179(.dina(n10801), .dinb(b54 ), .dout(n21438));
  jand g21180(.dina(n11107), .dinb(b53 ), .dout(n21439));
  jor  g21181(.dina(n21439), .dinb(n21438), .dout(n21440));
  jxor g21182(.dina(n21440), .dinb(n21437), .dout(n21441));
  jnot g21183(.din(n21441), .dout(n21442));
  jor  g21184(.dina(n10806), .dinb(n8806), .dout(n21443));
  jor  g21185(.dina(n10485), .dinb(n8231), .dout(n21444));
  jor  g21186(.dina(n10809), .dinb(n8789), .dout(n21445));
  jor  g21187(.dina(n10811), .dinb(n8809), .dout(n21446));
  jand g21188(.dina(n21446), .dinb(n21445), .dout(n21447));
  jand g21189(.dina(n21447), .dinb(n21444), .dout(n21448));
  jand g21190(.dina(n21448), .dinb(n21443), .dout(n21449));
  jxor g21191(.dina(n21449), .dinb(a62 ), .dout(n21450));
  jxor g21192(.dina(n21450), .dinb(n21442), .dout(n21451));
  jxor g21193(.dina(n21451), .dinb(n21436), .dout(n21452));
  jxor g21194(.dina(n21452), .dinb(n21432), .dout(n21453));
  jxor g21195(.dina(n21453), .dinb(n21423), .dout(n21454));
  jxor g21196(.dina(n21454), .dinb(n21420), .dout(n21455));
  jand g21197(.dina(n21345), .dinb(n21340), .dout(n21456));
  jnot g21198(.din(n21456), .dout(n21457));
  jnot g21199(.din(n21345), .dout(n21458));
  jand g21200(.dina(n21458), .dinb(n21339), .dout(n21459));
  jor  g21201(.dina(n21390), .dinb(n21459), .dout(n21460));
  jand g21202(.dina(n21460), .dinb(n21457), .dout(n21461));
  jxor g21203(.dina(n21461), .dinb(n21455), .dout(n21462));
  jxor g21204(.dina(n21462), .dinb(n21403), .dout(f117 ));
  jand g21205(.dina(n21461), .dinb(n21455), .dout(n21464));
  jand g21206(.dina(n21462), .dinb(n21403), .dout(n21465));
  jor  g21207(.dina(n21465), .dinb(n21464), .dout(n21466));
  jand g21208(.dina(n21419), .dinb(n21412), .dout(n21467));
  jand g21209(.dina(n21454), .dinb(n21420), .dout(n21468));
  jor  g21210(.dina(n21468), .dinb(n21467), .dout(n21469));
  jand g21211(.dina(n21452), .dinb(n21432), .dout(n21470));
  jand g21212(.dina(n21453), .dinb(n21423), .dout(n21471));
  jor  g21213(.dina(n21471), .dinb(n21470), .dout(n21472));
  jor  g21214(.dina(n10311), .dinb(n9891), .dout(n21473));
  jor  g21215(.dina(n9593), .dinb(n9413), .dout(n21474));
  jor  g21216(.dina(n9894), .dinb(n9725), .dout(n21475));
  jor  g21217(.dina(n9896), .dinb(n10314), .dout(n21476));
  jand g21218(.dina(n21476), .dinb(n21475), .dout(n21477));
  jand g21219(.dina(n21477), .dinb(n21474), .dout(n21478));
  jand g21220(.dina(n21478), .dinb(n21473), .dout(n21479));
  jxor g21221(.dina(n21479), .dinb(a59 ), .dout(n21480));
  jnot g21222(.din(n21480), .dout(n21481));
  jor  g21223(.dina(n21450), .dinb(n21442), .dout(n21482));
  jand g21224(.dina(n21451), .dinb(n21436), .dout(n21483));
  jnot g21225(.din(n21483), .dout(n21484));
  jand g21226(.dina(n21484), .dinb(n21482), .dout(n21485));
  jnot g21227(.din(n21485), .dout(n21486));
  jand g21228(.dina(n21375), .dinb(n21341), .dout(n21487));
  jand g21229(.dina(n21440), .dinb(n21437), .dout(n21488));
  jor  g21230(.dina(n21488), .dinb(n21487), .dout(n21489));
  jand g21231(.dina(n10801), .dinb(b55 ), .dout(n21490));
  jand g21232(.dina(n11107), .dinb(b54 ), .dout(n21491));
  jor  g21233(.dina(n21491), .dinb(n21490), .dout(n21492));
  jnot g21234(.din(n21492), .dout(n21493));
  jxor g21235(.dina(n21493), .dinb(n21489), .dout(n21494));
  jnot g21236(.din(n21494), .dout(n21495));
  jor  g21237(.dina(n10806), .dinb(n9387), .dout(n21496));
  jor  g21238(.dina(n10485), .dinb(n8789), .dout(n21497));
  jor  g21239(.dina(n10809), .dinb(n8809), .dout(n21498));
  jor  g21240(.dina(n10811), .dinb(n9390), .dout(n21499));
  jand g21241(.dina(n21499), .dinb(n21498), .dout(n21500));
  jand g21242(.dina(n21500), .dinb(n21497), .dout(n21501));
  jand g21243(.dina(n21501), .dinb(n21496), .dout(n21502));
  jxor g21244(.dina(n21502), .dinb(a62 ), .dout(n21503));
  jxor g21245(.dina(n21503), .dinb(n21495), .dout(n21504));
  jxor g21246(.dina(n21504), .dinb(n21486), .dout(n21505));
  jxor g21247(.dina(n21505), .dinb(n21481), .dout(n21506));
  jxor g21248(.dina(n21506), .dinb(n21472), .dout(n21507));
  jor  g21249(.dina(n10978), .dinb(n8978), .dout(n21508));
  jor  g21250(.dina(n8677), .dinb(n10637), .dout(n21509));
  jor  g21251(.dina(n8981), .dinb(n10964), .dout(n21510));
  jand g21252(.dina(n21510), .dinb(n21509), .dout(n21511));
  jand g21253(.dina(n21511), .dinb(n21508), .dout(n21512));
  jxor g21254(.dina(n21512), .dinb(a56 ), .dout(n21513));
  jnot g21255(.din(n21513), .dout(n21514));
  jxor g21256(.dina(n21514), .dinb(n21507), .dout(n21515));
  jxor g21257(.dina(n21515), .dinb(n21469), .dout(n21516));
  jxor g21258(.dina(n21516), .dinb(n21466), .dout(f118 ));
  jand g21259(.dina(n21504), .dinb(n21486), .dout(n21518));
  jand g21260(.dina(n21505), .dinb(n21481), .dout(n21519));
  jor  g21261(.dina(n21519), .dinb(n21518), .dout(n21520));
  jnot g21262(.din(n21520), .dout(n21521));
  jnot g21263(.din(a56 ), .dout(n21522));
  jand g21264(.dina(n11296), .dinb(n8368), .dout(n21523));
  jor  g21265(.dina(n21523), .dinb(n8678), .dout(n21524));
  jand g21266(.dina(n21524), .dinb(b63 ), .dout(n21525));
  jxor g21267(.dina(n21525), .dinb(n21522), .dout(n21526));
  jxor g21268(.dina(n21526), .dinb(n21521), .dout(n21527));
  jand g21269(.dina(n21493), .dinb(n21489), .dout(n21528));
  jnot g21270(.din(n21528), .dout(n21529));
  jor  g21271(.dina(n21503), .dinb(n21495), .dout(n21530));
  jand g21272(.dina(n21530), .dinb(n21529), .dout(n21531));
  jnot g21273(.din(n21531), .dout(n21532));
  jor  g21274(.dina(n10806), .dinb(n9410), .dout(n21533));
  jor  g21275(.dina(n10485), .dinb(n8809), .dout(n21534));
  jor  g21276(.dina(n10809), .dinb(n9390), .dout(n21535));
  jor  g21277(.dina(n10811), .dinb(n9413), .dout(n21536));
  jand g21278(.dina(n21536), .dinb(n21535), .dout(n21537));
  jand g21279(.dina(n21537), .dinb(n21534), .dout(n21538));
  jand g21280(.dina(n21538), .dinb(n21533), .dout(n21539));
  jxor g21281(.dina(n21539), .dinb(a62 ), .dout(n21540));
  jnot g21282(.din(n21540), .dout(n21541));
  jand g21283(.dina(n10801), .dinb(b56 ), .dout(n21542));
  jand g21284(.dina(n11107), .dinb(b55 ), .dout(n21543));
  jor  g21285(.dina(n21543), .dinb(n21542), .dout(n21544));
  jxor g21286(.dina(n21544), .dinb(n21493), .dout(n21545));
  jxor g21287(.dina(n21545), .dinb(n21541), .dout(n21546));
  jxor g21288(.dina(n21546), .dinb(n21532), .dout(n21547));
  jor  g21289(.dina(n10634), .dinb(n9891), .dout(n21548));
  jor  g21290(.dina(n9593), .dinb(n9725), .dout(n21549));
  jor  g21291(.dina(n9894), .dinb(n10314), .dout(n21550));
  jor  g21292(.dina(n9896), .dinb(n10637), .dout(n21551));
  jand g21293(.dina(n21551), .dinb(n21550), .dout(n21552));
  jand g21294(.dina(n21552), .dinb(n21549), .dout(n21553));
  jand g21295(.dina(n21553), .dinb(n21548), .dout(n21554));
  jxor g21296(.dina(n21554), .dinb(a59 ), .dout(n21555));
  jnot g21297(.din(n21555), .dout(n21556));
  jxor g21298(.dina(n21556), .dinb(n21547), .dout(n21557));
  jxor g21299(.dina(n21557), .dinb(n21527), .dout(n21558));
  jor  g21300(.dina(n21506), .dinb(n21472), .dout(n21559));
  jand g21301(.dina(n21506), .dinb(n21472), .dout(n21560));
  jor  g21302(.dina(n21514), .dinb(n21560), .dout(n21561));
  jand g21303(.dina(n21561), .dinb(n21559), .dout(n21562));
  jxor g21304(.dina(n21562), .dinb(n21558), .dout(n21563));
  jand g21305(.dina(n21515), .dinb(n21469), .dout(n21564));
  jand g21306(.dina(n21516), .dinb(n21466), .dout(n21565));
  jor  g21307(.dina(n21565), .dinb(n21564), .dout(n21566));
  jxor g21308(.dina(n21566), .dinb(n21563), .dout(f119 ));
  jand g21309(.dina(n21544), .dinb(n21493), .dout(n21568));
  jand g21310(.dina(n21545), .dinb(n21541), .dout(n21569));
  jor  g21311(.dina(n21569), .dinb(n21568), .dout(n21570));
  jand g21312(.dina(n10801), .dinb(b57 ), .dout(n21571));
  jand g21313(.dina(n11107), .dinb(b56 ), .dout(n21572));
  jor  g21314(.dina(n21572), .dinb(n21571), .dout(n21573));
  jxor g21315(.dina(n21573), .dinb(n21522), .dout(n21574));
  jxor g21316(.dina(n21574), .dinb(n21492), .dout(n21575));
  jxor g21317(.dina(n21575), .dinb(n21570), .dout(n21576));
  jnot g21318(.din(n21576), .dout(n21577));
  jor  g21319(.dina(n10806), .dinb(n9722), .dout(n21578));
  jor  g21320(.dina(n10485), .dinb(n9390), .dout(n21579));
  jor  g21321(.dina(n10809), .dinb(n9413), .dout(n21580));
  jor  g21322(.dina(n10811), .dinb(n9725), .dout(n21581));
  jand g21323(.dina(n21581), .dinb(n21580), .dout(n21582));
  jand g21324(.dina(n21582), .dinb(n21579), .dout(n21583));
  jand g21325(.dina(n21583), .dinb(n21578), .dout(n21584));
  jxor g21326(.dina(n21584), .dinb(a62 ), .dout(n21585));
  jxor g21327(.dina(n21585), .dinb(n21577), .dout(n21586));
  jor  g21328(.dina(n10961), .dinb(n9891), .dout(n21587));
  jor  g21329(.dina(n9593), .dinb(n10314), .dout(n21588));
  jor  g21330(.dina(n9894), .dinb(n10637), .dout(n21589));
  jor  g21331(.dina(n9896), .dinb(n10964), .dout(n21590));
  jand g21332(.dina(n21590), .dinb(n21589), .dout(n21591));
  jand g21333(.dina(n21591), .dinb(n21588), .dout(n21592));
  jand g21334(.dina(n21592), .dinb(n21587), .dout(n21593));
  jxor g21335(.dina(n21593), .dinb(a59 ), .dout(n21594));
  jnot g21336(.din(n21594), .dout(n21595));
  jnot g21337(.din(n21546), .dout(n21596));
  jand g21338(.dina(n21596), .dinb(n21531), .dout(n21597));
  jnot g21339(.din(n21597), .dout(n21598));
  jand g21340(.dina(n21546), .dinb(n21532), .dout(n21599));
  jor  g21341(.dina(n21556), .dinb(n21599), .dout(n21600));
  jand g21342(.dina(n21600), .dinb(n21598), .dout(n21601));
  jxor g21343(.dina(n21601), .dinb(n21595), .dout(n21602));
  jxor g21344(.dina(n21602), .dinb(n21586), .dout(n21603));
  jand g21345(.dina(n21526), .dinb(n21521), .dout(n21604));
  jnot g21346(.din(n21604), .dout(n21605));
  jnot g21347(.din(n21526), .dout(n21606));
  jand g21348(.dina(n21606), .dinb(n21520), .dout(n21607));
  jor  g21349(.dina(n21557), .dinb(n21607), .dout(n21608));
  jand g21350(.dina(n21608), .dinb(n21605), .dout(n21609));
  jxor g21351(.dina(n21609), .dinb(n21603), .dout(n21610));
  jand g21352(.dina(n21562), .dinb(n21558), .dout(n21611));
  jand g21353(.dina(n21566), .dinb(n21563), .dout(n21612));
  jor  g21354(.dina(n21612), .dinb(n21611), .dout(n21613));
  jxor g21355(.dina(n21613), .dinb(n21610), .dout(f120 ));
  jand g21356(.dina(n21601), .dinb(n21595), .dout(n21615));
  jand g21357(.dina(n21602), .dinb(n21586), .dout(n21616));
  jor  g21358(.dina(n21616), .dinb(n21615), .dout(n21617));
  jand g21359(.dina(n21575), .dinb(n21570), .dout(n21618));
  jnot g21360(.din(n21618), .dout(n21619));
  jor  g21361(.dina(n21585), .dinb(n21577), .dout(n21620));
  jand g21362(.dina(n21620), .dinb(n21619), .dout(n21621));
  jand g21363(.dina(n21573), .dinb(n21522), .dout(n21622));
  jand g21364(.dina(n21574), .dinb(n21492), .dout(n21623));
  jor  g21365(.dina(n21623), .dinb(n21622), .dout(n21624));
  jand g21366(.dina(n10801), .dinb(b58 ), .dout(n21625));
  jand g21367(.dina(n11107), .dinb(b57 ), .dout(n21626));
  jor  g21368(.dina(n21626), .dinb(n21625), .dout(n21627));
  jnot g21369(.din(n21627), .dout(n21628));
  jxor g21370(.dina(n21628), .dinb(n21624), .dout(n21629));
  jor  g21371(.dina(n10311), .dinb(n10806), .dout(n21630));
  jor  g21372(.dina(n10485), .dinb(n9413), .dout(n21631));
  jor  g21373(.dina(n10809), .dinb(n9725), .dout(n21632));
  jor  g21374(.dina(n10811), .dinb(n10314), .dout(n21633));
  jand g21375(.dina(n21633), .dinb(n21632), .dout(n21634));
  jand g21376(.dina(n21634), .dinb(n21631), .dout(n21635));
  jand g21377(.dina(n21635), .dinb(n21630), .dout(n21636));
  jxor g21378(.dina(n21636), .dinb(a62 ), .dout(n21637));
  jnot g21379(.din(n21637), .dout(n21638));
  jxor g21380(.dina(n21638), .dinb(n21629), .dout(n21639));
  jxor g21381(.dina(n21639), .dinb(n21621), .dout(n21640));
  jor  g21382(.dina(n10978), .dinb(n9891), .dout(n21641));
  jor  g21383(.dina(n9593), .dinb(n10637), .dout(n21642));
  jor  g21384(.dina(n9894), .dinb(n10964), .dout(n21643));
  jand g21385(.dina(n21643), .dinb(n21642), .dout(n21644));
  jand g21386(.dina(n21644), .dinb(n21641), .dout(n21645));
  jxor g21387(.dina(n21645), .dinb(a59 ), .dout(n21646));
  jxor g21388(.dina(n21646), .dinb(n21640), .dout(n21647));
  jxor g21389(.dina(n21647), .dinb(n21617), .dout(n21648));
  jand g21390(.dina(n21609), .dinb(n21603), .dout(n21649));
  jand g21391(.dina(n21613), .dinb(n21610), .dout(n21650));
  jor  g21392(.dina(n21650), .dinb(n21649), .dout(n21651));
  jxor g21393(.dina(n21651), .dinb(n21648), .dout(f121 ));
  jand g21394(.dina(n21647), .dinb(n21617), .dout(n21653));
  jand g21395(.dina(n21651), .dinb(n21648), .dout(n21654));
  jor  g21396(.dina(n21654), .dinb(n21653), .dout(n21655));
  jand g21397(.dina(n21628), .dinb(n21624), .dout(n21656));
  jand g21398(.dina(n21638), .dinb(n21629), .dout(n21657));
  jor  g21399(.dina(n21657), .dinb(n21656), .dout(n21658));
  jand g21400(.dina(n10801), .dinb(b59 ), .dout(n21659));
  jand g21401(.dina(n11107), .dinb(b58 ), .dout(n21660));
  jor  g21402(.dina(n21660), .dinb(n21659), .dout(n21661));
  jnot g21403(.din(n21661), .dout(n21662));
  jxor g21404(.dina(n21662), .dinb(n21627), .dout(n21663));
  jxor g21405(.dina(n21663), .dinb(n21658), .dout(n21664));
  jor  g21406(.dina(n10634), .dinb(n10806), .dout(n21665));
  jor  g21407(.dina(n10485), .dinb(n9725), .dout(n21666));
  jor  g21408(.dina(n10809), .dinb(n10314), .dout(n21667));
  jor  g21409(.dina(n10811), .dinb(n10637), .dout(n21668));
  jand g21410(.dina(n21668), .dinb(n21667), .dout(n21669));
  jand g21411(.dina(n21669), .dinb(n21666), .dout(n21670));
  jand g21412(.dina(n21670), .dinb(n21665), .dout(n21671));
  jxor g21413(.dina(n21671), .dinb(a62 ), .dout(n21672));
  jnot g21414(.din(a59 ), .dout(n21673));
  jand g21415(.dina(n11296), .dinb(n9244), .dout(n21674));
  jor  g21416(.dina(n21674), .dinb(n9594), .dout(n21675));
  jand g21417(.dina(n21675), .dinb(b63 ), .dout(n21676));
  jxor g21418(.dina(n21676), .dinb(n21673), .dout(n21677));
  jxor g21419(.dina(n21677), .dinb(n21672), .dout(n21678));
  jxor g21420(.dina(n21678), .dinb(n21664), .dout(n21679));
  jnot g21421(.din(n21621), .dout(n21680));
  jor  g21422(.dina(n21639), .dinb(n21680), .dout(n21681));
  jand g21423(.dina(n21639), .dinb(n21680), .dout(n21682));
  jnot g21424(.din(n21646), .dout(n21683));
  jor  g21425(.dina(n21683), .dinb(n21682), .dout(n21684));
  jand g21426(.dina(n21684), .dinb(n21681), .dout(n21685));
  jxor g21427(.dina(n21685), .dinb(n21679), .dout(n21686));
  jxor g21428(.dina(n21686), .dinb(n21655), .dout(f122 ));
  jand g21429(.dina(n21685), .dinb(n21679), .dout(n21688));
  jand g21430(.dina(n21686), .dinb(n21655), .dout(n21689));
  jor  g21431(.dina(n21689), .dinb(n21688), .dout(n21690));
  jnot g21432(.din(n21672), .dout(n21691));
  jnot g21433(.din(n21677), .dout(n21692));
  jand g21434(.dina(n21692), .dinb(n21691), .dout(n21693));
  jand g21435(.dina(n21678), .dinb(n21664), .dout(n21694));
  jor  g21436(.dina(n21694), .dinb(n21693), .dout(n21695));
  jand g21437(.dina(n21662), .dinb(n21627), .dout(n21696));
  jand g21438(.dina(n21663), .dinb(n21658), .dout(n21697));
  jor  g21439(.dina(n21697), .dinb(n21696), .dout(n21698));
  jxor g21440(.dina(n21661), .dinb(n21673), .dout(n21699));
  jand g21441(.dina(n10801), .dinb(b60 ), .dout(n21700));
  jand g21442(.dina(n11107), .dinb(b59 ), .dout(n21701));
  jor  g21443(.dina(n21701), .dinb(n21700), .dout(n21702));
  jxor g21444(.dina(n21702), .dinb(n21699), .dout(n21703));
  jor  g21445(.dina(n10961), .dinb(n10806), .dout(n21704));
  jor  g21446(.dina(n10485), .dinb(n10314), .dout(n21705));
  jor  g21447(.dina(n10809), .dinb(n10637), .dout(n21706));
  jor  g21448(.dina(n10811), .dinb(n10964), .dout(n21707));
  jand g21449(.dina(n21707), .dinb(n21706), .dout(n21708));
  jand g21450(.dina(n21708), .dinb(n21705), .dout(n21709));
  jand g21451(.dina(n21709), .dinb(n21704), .dout(n21710));
  jxor g21452(.dina(n21710), .dinb(a62 ), .dout(n21711));
  jnot g21453(.din(n21711), .dout(n21712));
  jxor g21454(.dina(n21712), .dinb(n21703), .dout(n21713));
  jxor g21455(.dina(n21713), .dinb(n21698), .dout(n21714));
  jxor g21456(.dina(n21714), .dinb(n21695), .dout(n21715));
  jxor g21457(.dina(n21715), .dinb(n21690), .dout(f123 ));
  jand g21458(.dina(n21714), .dinb(n21695), .dout(n21717));
  jand g21459(.dina(n21715), .dinb(n21690), .dout(n21718));
  jor  g21460(.dina(n21718), .dinb(n21717), .dout(n21719));
  jand g21461(.dina(n21712), .dinb(n21703), .dout(n21720));
  jand g21462(.dina(n21713), .dinb(n21698), .dout(n21721));
  jor  g21463(.dina(n21721), .dinb(n21720), .dout(n21722));
  jand g21464(.dina(n21661), .dinb(n21673), .dout(n21723));
  jand g21465(.dina(n21702), .dinb(n21699), .dout(n21724));
  jor  g21466(.dina(n21724), .dinb(n21723), .dout(n21725));
  jand g21467(.dina(n10801), .dinb(b61 ), .dout(n21726));
  jand g21468(.dina(n11107), .dinb(b60 ), .dout(n21727));
  jor  g21469(.dina(n21727), .dinb(n21726), .dout(n21728));
  jnot g21470(.din(n21728), .dout(n21729));
  jxor g21471(.dina(n21729), .dinb(n21725), .dout(n21730));
  jor  g21472(.dina(n10978), .dinb(n10806), .dout(n21731));
  jor  g21473(.dina(n10485), .dinb(n10637), .dout(n21732));
  jor  g21474(.dina(n10809), .dinb(n10964), .dout(n21733));
  jand g21475(.dina(n21733), .dinb(n21732), .dout(n21734));
  jand g21476(.dina(n21734), .dinb(n21731), .dout(n21735));
  jxor g21477(.dina(n21735), .dinb(a62 ), .dout(n21736));
  jnot g21478(.din(n21736), .dout(n21737));
  jxor g21479(.dina(n21737), .dinb(n21730), .dout(n21738));
  jxor g21480(.dina(n21738), .dinb(n21722), .dout(n21739));
  jxor g21481(.dina(n21739), .dinb(n21719), .dout(f124 ));
  jand g21482(.dina(n21738), .dinb(n21722), .dout(n21741));
  jand g21483(.dina(n21739), .dinb(n21719), .dout(n21742));
  jor  g21484(.dina(n21742), .dinb(n21741), .dout(n21743));
  jand g21485(.dina(n21729), .dinb(n21725), .dout(n21744));
  jand g21486(.dina(n21737), .dinb(n21730), .dout(n21745));
  jor  g21487(.dina(n21745), .dinb(n21744), .dout(n21746));
  jand g21488(.dina(n10801), .dinb(b62 ), .dout(n21747));
  jand g21489(.dina(n11107), .dinb(b61 ), .dout(n21748));
  jor  g21490(.dina(n21748), .dinb(n21747), .dout(n21749));
  jxor g21491(.dina(n21749), .dinb(n21729), .dout(n21750));
  jnot g21492(.din(a62 ), .dout(n21751));
  jand g21493(.dina(n11296), .dinb(n10150), .dout(n21752));
  jor  g21494(.dina(n21752), .dinb(n10486), .dout(n21753));
  jand g21495(.dina(n21753), .dinb(b63 ), .dout(n21754));
  jxor g21496(.dina(n21754), .dinb(n21751), .dout(n21755));
  jnot g21497(.din(n21755), .dout(n21756));
  jxor g21498(.dina(n21756), .dinb(n21750), .dout(n21757));
  jxor g21499(.dina(n21757), .dinb(n21746), .dout(n21758));
  jxor g21500(.dina(n21758), .dinb(n21743), .dout(f125 ));
  jand g21501(.dina(n21757), .dinb(n21746), .dout(n21760));
  jand g21502(.dina(n21758), .dinb(n21743), .dout(n21761));
  jor  g21503(.dina(n21761), .dinb(n21760), .dout(n21762));
  jand g21504(.dina(n21749), .dinb(n21729), .dout(n21763));
  jand g21505(.dina(n21756), .dinb(n21750), .dout(n21764));
  jor  g21506(.dina(n21764), .dinb(n21763), .dout(n21765));
  jand g21507(.dina(b63 ), .dinb(a63 ), .dout(n21766));
  jand g21508(.dina(n10964), .dinb(a62 ), .dout(n21767));
  jor  g21509(.dina(n21767), .dinb(n21766), .dout(n21768));
  jand g21510(.dina(b62 ), .dinb(a62 ), .dout(n21769));
  jand g21511(.dina(n21769), .dinb(n11107), .dout(n21770));
  jnot g21512(.din(n21770), .dout(n21771));
  jand g21513(.dina(n21771), .dinb(n21768), .dout(n21772));
  jxor g21514(.dina(n21772), .dinb(n21729), .dout(n21773));
  jxor g21515(.dina(n21773), .dinb(n21765), .dout(n21774));
  jxor g21516(.dina(n21774), .dinb(n21762), .dout(f126 ));
  jand g21517(.dina(n21773), .dinb(n21765), .dout(n21776));
  jand g21518(.dina(n21774), .dinb(n21762), .dout(n21777));
  jor  g21519(.dina(n21777), .dinb(n21776), .dout(n21778));
  jnot g21520(.din(n21766), .dout(n21779));
  jor  g21521(.dina(n21772), .dinb(n21729), .dout(n21780));
  jnot g21522(.din(n21780), .dout(n21781));
  jor  g21523(.dina(n21781), .dinb(n21779), .dout(n21782));
  jand g21524(.dina(n21766), .dinb(a62 ), .dout(n21783));
  jor  g21525(.dina(n21783), .dinb(n21780), .dout(n21784));
  jand g21526(.dina(n21784), .dinb(n21782), .dout(n21785));
  jxor g21527(.dina(n21785), .dinb(n21778), .dout(f127 ));
endmodule


