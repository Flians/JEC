// Benchmark "top" written by ABC on Wed May 27 23:36:46 2020

module top ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , a16 ,
    a17 , a18 , a19 , a20 , a21 , a22 , a23 , a24 ,
    a25 , a26 , a27 , a28 , a29 , a30 , a31 , a32 ,
    a33 , a34 , a35 , a36 , a37 , a38 , a39 , a40 ,
    a41 , a42 , a43 , a44 , a45 , a46 , a47 , a48 ,
    a49 , a50 , a51 , a52 , a53 , a54 , a55 , a56 ,
    a57 , a58 , a59 , a60 , a61 , a62 , a63 , a64 ,
    a65 , a66 , a67 , a68 , a69 , a70 , a71 , a72 ,
    a73 , a74 , a75 , a76 , a77 , a78 , a79 , a80 ,
    a81 , a82 , a83 , a84 , a85 , a86 , a87 , a88 ,
    a89 , a90 , a91 , a92 , a93 , a94 , a95 , a96 ,
    a97 , a98 , a99 , a100 , a101 , a102 , a103 ,
    a104 , a105 , a106 , a107 , a108 , a109 , a110 ,
    a111 , a112 , a113 , a114 , a115 , a116 , a117 ,
    a118 , a119 , a120 , a121 , a122 , a123 , a124 ,
    a125 , a126 , a127 , shift0 , shift1 , shift2 ,
    shift3 , shift4 , shift5 , shift6 ,
    result0 , result1 , result2 , result3 , result4 ,
    result5 , result6 , result7 , result8 , result9 ,
    result10 , result11 , result12 , result13 , result14 ,
    result15 , result16 , result17 , result18 , result19 ,
    result20 , result21 , result22 , result23 , result24 ,
    result25 , result26 , result27 , result28 , result29 ,
    result30 , result31 , result32 , result33 , result34 ,
    result35 , result36 , result37 , result38 , result39 ,
    result40 , result41 , result42 , result43 , result44 ,
    result45 , result46 , result47 , result48 , result49 ,
    result50 , result51 , result52 , result53 , result54 ,
    result55 , result56 , result57 , result58 , result59 ,
    result60 , result61 , result62 , result63 , result64 ,
    result65 , result66 , result67 , result68 , result69 ,
    result70 , result71 , result72 , result73 , result74 ,
    result75 , result76 , result77 , result78 , result79 ,
    result80 , result81 , result82 , result83 , result84 ,
    result85 , result86 , result87 , result88 , result89 ,
    result90 , result91 , result92 , result93 , result94 ,
    result95 , result96 , result97 , result98 , result99 ,
    result100 , result101 , result102 , result103 ,
    result104 , result105 , result106 , result107 ,
    result108 , result109 , result110 , result111 ,
    result112 , result113 , result114 , result115 ,
    result116 , result117 , result118 , result119 ,
    result120 , result121 , result122 , result123 ,
    result124 , result125 , result126 , result127   );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    a16 , a17 , a18 , a19 , a20 , a21 , a22 , a23 ,
    a24 , a25 , a26 , a27 , a28 , a29 , a30 , a31 ,
    a32 , a33 , a34 , a35 , a36 , a37 , a38 , a39 ,
    a40 , a41 , a42 , a43 , a44 , a45 , a46 , a47 ,
    a48 , a49 , a50 , a51 , a52 , a53 , a54 , a55 ,
    a56 , a57 , a58 , a59 , a60 , a61 , a62 , a63 ,
    a64 , a65 , a66 , a67 , a68 , a69 , a70 , a71 ,
    a72 , a73 , a74 , a75 , a76 , a77 , a78 , a79 ,
    a80 , a81 , a82 , a83 , a84 , a85 , a86 , a87 ,
    a88 , a89 , a90 , a91 , a92 , a93 , a94 , a95 ,
    a96 , a97 , a98 , a99 , a100 , a101 , a102 ,
    a103 , a104 , a105 , a106 , a107 , a108 , a109 ,
    a110 , a111 , a112 , a113 , a114 , a115 , a116 ,
    a117 , a118 , a119 , a120 , a121 , a122 , a123 ,
    a124 , a125 , a126 , a127 , shift0 , shift1 ,
    shift2 , shift3 , shift4 , shift5 , shift6 ;
  output result0 , result1 , result2 , result3 , result4 ,
    result5 , result6 , result7 , result8 , result9 ,
    result10 , result11 , result12 , result13 , result14 ,
    result15 , result16 , result17 , result18 , result19 ,
    result20 , result21 , result22 , result23 , result24 ,
    result25 , result26 , result27 , result28 , result29 ,
    result30 , result31 , result32 , result33 , result34 ,
    result35 , result36 , result37 , result38 , result39 ,
    result40 , result41 , result42 , result43 , result44 ,
    result45 , result46 , result47 , result48 , result49 ,
    result50 , result51 , result52 , result53 , result54 ,
    result55 , result56 , result57 , result58 , result59 ,
    result60 , result61 , result62 , result63 , result64 ,
    result65 , result66 , result67 , result68 , result69 ,
    result70 , result71 , result72 , result73 , result74 ,
    result75 , result76 , result77 , result78 , result79 ,
    result80 , result81 , result82 , result83 , result84 ,
    result85 , result86 , result87 , result88 , result89 ,
    result90 , result91 , result92 , result93 , result94 ,
    result95 , result96 , result97 , result98 , result99 ,
    result100 , result101 , result102 , result103 ,
    result104 , result105 , result106 , result107 ,
    result108 , result109 , result110 , result111 ,
    result112 , result113 , result114 , result115 ,
    result116 , result117 , result118 , result119 ,
    result120 , result121 , result122 , result123 ,
    result124 , result125 , result126 , result127 ;
  wire n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n639, n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
    n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
    n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
    n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
    n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
    n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
    n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
    n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
    n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2367, n2368,
    n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
    n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501, n2503, n2504, n2505, n2506,
    n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
    n2634, n2635, n2636, n2637, n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
    n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2758, n2759, n2760, n2761,
    n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
    n2772, n2773, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2923, n2924, n2925, n2926, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
    n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3030, n3031, n3033, n3034, n3036, n3037, n3039, n3040,
    n3042, n3043, n3045, n3046, n3048, n3049, n3051, n3052, n3054, n3055,
    n3057, n3058, n3060, n3061, n3063, n3064, n3066, n3067, n3069, n3070,
    n3072, n3073, n3075, n3076, n3078, n3079, n3081, n3082, n3084, n3085,
    n3087, n3088, n3090, n3091, n3093, n3094, n3096, n3097, n3099, n3100,
    n3102, n3103, n3105, n3106, n3108, n3109, n3111, n3112, n3114, n3115,
    n3117, n3118, n3120, n3121, n3123, n3124, n3126, n3127, n3129, n3130,
    n3132, n3133, n3135, n3136, n3138, n3139, n3141, n3142, n3144, n3145,
    n3147, n3148, n3150, n3151, n3153, n3154, n3156, n3157, n3159, n3160,
    n3162, n3163, n3165, n3166, n3168, n3169, n3171, n3172, n3174, n3175,
    n3177, n3178, n3180, n3181, n3183, n3184, n3186, n3187, n3189, n3190,
    n3192, n3193, n3195, n3196, n3198, n3199, n3201, n3202, n3204, n3205,
    n3207, n3208, n3210, n3211, n3213, n3214, n3216, n3217, n3219, n3220;
  jnot g0000(.din(shift6 ), .dout(n263));
  jnot g0001(.din(shift4 ), .dout(n264));
  jand g0002(.dina(shift5 ), .dinb(n264), .dout(n265));
  jnot g0003(.din(shift3 ), .dout(n266));
  jand g0004(.dina(n266), .dinb(shift2 ), .dout(n267));
  jor  g0005(.dina(shift0 ), .dinb(a28 ), .dout(n268));
  jnot g0006(.din(shift0 ), .dout(n269));
  jor  g0007(.dina(n269), .dinb(a27 ), .dout(n270));
  jand g0008(.dina(n270), .dinb(n268), .dout(n271));
  jor  g0009(.dina(n271), .dinb(shift1 ), .dout(n272));
  jnot g0010(.din(shift1 ), .dout(n273));
  jor  g0011(.dina(shift0 ), .dinb(a26 ), .dout(n274));
  jor  g0012(.dina(n269), .dinb(a25 ), .dout(n275));
  jand g0013(.dina(n275), .dinb(n274), .dout(n276));
  jor  g0014(.dina(n276), .dinb(n273), .dout(n277));
  jand g0015(.dina(n277), .dinb(n272), .dout(n278));
  jand g0016(.dina(n278), .dinb(n267), .dout(n279));
  jnot g0017(.din(shift2 ), .dout(n280));
  jand g0018(.dina(shift3 ), .dinb(n280), .dout(n281));
  jor  g0019(.dina(shift0 ), .dinb(a24 ), .dout(n282));
  jor  g0020(.dina(n269), .dinb(a23 ), .dout(n283));
  jand g0021(.dina(n283), .dinb(n282), .dout(n284));
  jor  g0022(.dina(n284), .dinb(shift1 ), .dout(n285));
  jor  g0023(.dina(shift0 ), .dinb(a22 ), .dout(n286));
  jor  g0024(.dina(n269), .dinb(a21 ), .dout(n287));
  jand g0025(.dina(n287), .dinb(n286), .dout(n288));
  jor  g0026(.dina(n288), .dinb(n273), .dout(n289));
  jand g0027(.dina(n289), .dinb(n285), .dout(n290));
  jand g0028(.dina(n290), .dinb(n281), .dout(n291));
  jand g0029(.dina(shift3 ), .dinb(shift2 ), .dout(n292));
  jor  g0030(.dina(shift0 ), .dinb(a20 ), .dout(n293));
  jor  g0031(.dina(n269), .dinb(a19 ), .dout(n294));
  jand g0032(.dina(n294), .dinb(n293), .dout(n295));
  jor  g0033(.dina(n295), .dinb(shift1 ), .dout(n296));
  jor  g0034(.dina(shift0 ), .dinb(a18 ), .dout(n297));
  jor  g0035(.dina(n269), .dinb(a17 ), .dout(n298));
  jand g0036(.dina(n298), .dinb(n297), .dout(n299));
  jor  g0037(.dina(n299), .dinb(n273), .dout(n300));
  jand g0038(.dina(n300), .dinb(n296), .dout(n301));
  jand g0039(.dina(n301), .dinb(n292), .dout(n302));
  jor  g0040(.dina(n302), .dinb(n291), .dout(n303));
  jand g0041(.dina(n266), .dinb(n280), .dout(n304));
  jor  g0042(.dina(shift0 ), .dinb(a32 ), .dout(n305));
  jor  g0043(.dina(n269), .dinb(a31 ), .dout(n306));
  jand g0044(.dina(n306), .dinb(n305), .dout(n307));
  jor  g0045(.dina(n307), .dinb(shift1 ), .dout(n308));
  jor  g0046(.dina(shift0 ), .dinb(a30 ), .dout(n309));
  jor  g0047(.dina(n269), .dinb(a29 ), .dout(n310));
  jand g0048(.dina(n310), .dinb(n309), .dout(n311));
  jor  g0049(.dina(n311), .dinb(n273), .dout(n312));
  jand g0050(.dina(n312), .dinb(n308), .dout(n313));
  jand g0051(.dina(n313), .dinb(n304), .dout(n314));
  jor  g0052(.dina(n314), .dinb(n303), .dout(n315));
  jor  g0053(.dina(n315), .dinb(n279), .dout(n316));
  jand g0054(.dina(n316), .dinb(n265), .dout(n317));
  jnot g0055(.din(shift5 ), .dout(n318));
  jand g0056(.dina(n318), .dinb(shift4 ), .dout(n319));
  jor  g0057(.dina(shift0 ), .dinb(a36 ), .dout(n320));
  jor  g0058(.dina(n269), .dinb(a35 ), .dout(n321));
  jand g0059(.dina(n321), .dinb(n320), .dout(n322));
  jor  g0060(.dina(n322), .dinb(shift1 ), .dout(n323));
  jor  g0061(.dina(shift0 ), .dinb(a34 ), .dout(n324));
  jor  g0062(.dina(n269), .dinb(a33 ), .dout(n325));
  jand g0063(.dina(n325), .dinb(n324), .dout(n326));
  jor  g0064(.dina(n326), .dinb(n273), .dout(n327));
  jand g0065(.dina(n327), .dinb(n323), .dout(n328));
  jand g0066(.dina(n328), .dinb(n292), .dout(n329));
  jor  g0067(.dina(shift0 ), .dinb(a40 ), .dout(n330));
  jor  g0068(.dina(n269), .dinb(a39 ), .dout(n331));
  jand g0069(.dina(n331), .dinb(n330), .dout(n332));
  jand g0070(.dina(n332), .dinb(n273), .dout(n333));
  jor  g0071(.dina(shift0 ), .dinb(a38 ), .dout(n334));
  jor  g0072(.dina(n269), .dinb(a37 ), .dout(n335));
  jand g0073(.dina(n335), .dinb(n334), .dout(n336));
  jand g0074(.dina(n336), .dinb(shift1 ), .dout(n337));
  jor  g0075(.dina(n337), .dinb(n333), .dout(n338));
  jand g0076(.dina(n338), .dinb(n281), .dout(n339));
  jor  g0077(.dina(shift0 ), .dinb(a44 ), .dout(n340));
  jor  g0078(.dina(n269), .dinb(a43 ), .dout(n341));
  jand g0079(.dina(n341), .dinb(n340), .dout(n342));
  jor  g0080(.dina(n342), .dinb(shift1 ), .dout(n343));
  jor  g0081(.dina(shift0 ), .dinb(a42 ), .dout(n344));
  jor  g0082(.dina(n269), .dinb(a41 ), .dout(n345));
  jand g0083(.dina(n345), .dinb(n344), .dout(n346));
  jor  g0084(.dina(n346), .dinb(n273), .dout(n347));
  jand g0085(.dina(n347), .dinb(n343), .dout(n348));
  jand g0086(.dina(n348), .dinb(n267), .dout(n349));
  jor  g0087(.dina(n349), .dinb(n339), .dout(n350));
  jor  g0088(.dina(shift0 ), .dinb(a48 ), .dout(n351));
  jor  g0089(.dina(n269), .dinb(a47 ), .dout(n352));
  jand g0090(.dina(n352), .dinb(n351), .dout(n353));
  jor  g0091(.dina(n353), .dinb(shift1 ), .dout(n354));
  jor  g0092(.dina(shift0 ), .dinb(a46 ), .dout(n355));
  jor  g0093(.dina(n269), .dinb(a45 ), .dout(n356));
  jand g0094(.dina(n356), .dinb(n355), .dout(n357));
  jor  g0095(.dina(n357), .dinb(n273), .dout(n358));
  jand g0096(.dina(n358), .dinb(n354), .dout(n359));
  jand g0097(.dina(n359), .dinb(n304), .dout(n360));
  jor  g0098(.dina(n360), .dinb(n350), .dout(n361));
  jor  g0099(.dina(n361), .dinb(n329), .dout(n362));
  jand g0100(.dina(n362), .dinb(n319), .dout(n363));
  jand g0101(.dina(n318), .dinb(n264), .dout(n364));
  jor  g0102(.dina(shift0 ), .dinb(a64 ), .dout(n365));
  jor  g0103(.dina(n269), .dinb(a63 ), .dout(n366));
  jand g0104(.dina(n366), .dinb(n365), .dout(n367));
  jor  g0105(.dina(n367), .dinb(shift1 ), .dout(n368));
  jor  g0106(.dina(shift0 ), .dinb(a62 ), .dout(n369));
  jor  g0107(.dina(n269), .dinb(a61 ), .dout(n370));
  jand g0108(.dina(n370), .dinb(n369), .dout(n371));
  jor  g0109(.dina(n371), .dinb(n273), .dout(n372));
  jand g0110(.dina(n372), .dinb(n368), .dout(n373));
  jand g0111(.dina(n373), .dinb(n304), .dout(n374));
  jor  g0112(.dina(shift0 ), .dinb(a56 ), .dout(n375));
  jor  g0113(.dina(n269), .dinb(a55 ), .dout(n376));
  jand g0114(.dina(n376), .dinb(n375), .dout(n377));
  jor  g0115(.dina(n377), .dinb(shift1 ), .dout(n378));
  jor  g0116(.dina(shift0 ), .dinb(a54 ), .dout(n379));
  jor  g0117(.dina(n269), .dinb(a53 ), .dout(n380));
  jand g0118(.dina(n380), .dinb(n379), .dout(n381));
  jor  g0119(.dina(n381), .dinb(n273), .dout(n382));
  jand g0120(.dina(n382), .dinb(n378), .dout(n383));
  jand g0121(.dina(n383), .dinb(n281), .dout(n384));
  jor  g0122(.dina(shift0 ), .dinb(a60 ), .dout(n385));
  jor  g0123(.dina(n269), .dinb(a59 ), .dout(n386));
  jand g0124(.dina(n386), .dinb(n385), .dout(n387));
  jor  g0125(.dina(n387), .dinb(shift1 ), .dout(n388));
  jor  g0126(.dina(shift0 ), .dinb(a58 ), .dout(n389));
  jor  g0127(.dina(n269), .dinb(a57 ), .dout(n390));
  jand g0128(.dina(n390), .dinb(n389), .dout(n391));
  jor  g0129(.dina(n391), .dinb(n273), .dout(n392));
  jand g0130(.dina(n392), .dinb(n388), .dout(n393));
  jand g0131(.dina(n393), .dinb(n267), .dout(n394));
  jor  g0132(.dina(n394), .dinb(n384), .dout(n395));
  jor  g0133(.dina(shift0 ), .dinb(a52 ), .dout(n396));
  jor  g0134(.dina(n269), .dinb(a51 ), .dout(n397));
  jand g0135(.dina(n397), .dinb(n396), .dout(n398));
  jor  g0136(.dina(n398), .dinb(shift1 ), .dout(n399));
  jor  g0137(.dina(shift0 ), .dinb(a50 ), .dout(n400));
  jor  g0138(.dina(n269), .dinb(a49 ), .dout(n401));
  jand g0139(.dina(n401), .dinb(n400), .dout(n402));
  jor  g0140(.dina(n402), .dinb(n273), .dout(n403));
  jand g0141(.dina(n403), .dinb(n399), .dout(n404));
  jand g0142(.dina(n404), .dinb(n292), .dout(n405));
  jor  g0143(.dina(n405), .dinb(n395), .dout(n406));
  jor  g0144(.dina(n406), .dinb(n374), .dout(n407));
  jand g0145(.dina(n407), .dinb(n364), .dout(n408));
  jor  g0146(.dina(n408), .dinb(n363), .dout(n409));
  jand g0147(.dina(shift5 ), .dinb(shift4 ), .dout(n410));
  jor  g0148(.dina(shift0 ), .dinb(a12 ), .dout(n411));
  jor  g0149(.dina(n269), .dinb(a11 ), .dout(n412));
  jand g0150(.dina(n412), .dinb(n411), .dout(n413));
  jor  g0151(.dina(n413), .dinb(shift1 ), .dout(n414));
  jor  g0152(.dina(shift0 ), .dinb(a10 ), .dout(n415));
  jor  g0153(.dina(n269), .dinb(a9 ), .dout(n416));
  jand g0154(.dina(n416), .dinb(n415), .dout(n417));
  jor  g0155(.dina(n417), .dinb(n273), .dout(n418));
  jand g0156(.dina(n418), .dinb(n414), .dout(n419));
  jand g0157(.dina(n419), .dinb(n267), .dout(n420));
  jor  g0158(.dina(shift0 ), .dinb(a8 ), .dout(n421));
  jor  g0159(.dina(n269), .dinb(a7 ), .dout(n422));
  jand g0160(.dina(n422), .dinb(n421), .dout(n423));
  jor  g0161(.dina(n423), .dinb(shift1 ), .dout(n424));
  jor  g0162(.dina(shift0 ), .dinb(a6 ), .dout(n425));
  jor  g0163(.dina(n269), .dinb(a5 ), .dout(n426));
  jand g0164(.dina(n426), .dinb(n425), .dout(n427));
  jor  g0165(.dina(n427), .dinb(n273), .dout(n428));
  jand g0166(.dina(n428), .dinb(n424), .dout(n429));
  jand g0167(.dina(n429), .dinb(n281), .dout(n430));
  jor  g0168(.dina(shift0 ), .dinb(a4 ), .dout(n431));
  jor  g0169(.dina(n269), .dinb(a3 ), .dout(n432));
  jand g0170(.dina(n432), .dinb(n431), .dout(n433));
  jor  g0171(.dina(n433), .dinb(shift1 ), .dout(n434));
  jor  g0172(.dina(shift0 ), .dinb(a2 ), .dout(n435));
  jor  g0173(.dina(n269), .dinb(a1 ), .dout(n436));
  jand g0174(.dina(n436), .dinb(n435), .dout(n437));
  jor  g0175(.dina(n437), .dinb(n273), .dout(n438));
  jand g0176(.dina(n438), .dinb(n434), .dout(n439));
  jand g0177(.dina(n439), .dinb(n292), .dout(n440));
  jor  g0178(.dina(n440), .dinb(n430), .dout(n441));
  jor  g0179(.dina(shift0 ), .dinb(a16 ), .dout(n442));
  jor  g0180(.dina(n269), .dinb(a15 ), .dout(n443));
  jand g0181(.dina(n443), .dinb(n442), .dout(n444));
  jor  g0182(.dina(n444), .dinb(shift1 ), .dout(n445));
  jor  g0183(.dina(shift0 ), .dinb(a14 ), .dout(n446));
  jor  g0184(.dina(n269), .dinb(a13 ), .dout(n447));
  jand g0185(.dina(n447), .dinb(n446), .dout(n448));
  jor  g0186(.dina(n448), .dinb(n273), .dout(n449));
  jand g0187(.dina(n449), .dinb(n445), .dout(n450));
  jand g0188(.dina(n450), .dinb(n304), .dout(n451));
  jor  g0189(.dina(n451), .dinb(n441), .dout(n452));
  jor  g0190(.dina(n452), .dinb(n420), .dout(n453));
  jand g0191(.dina(n453), .dinb(n410), .dout(n454));
  jor  g0192(.dina(n454), .dinb(n409), .dout(n455));
  jor  g0193(.dina(n455), .dinb(n317), .dout(n456));
  jor  g0194(.dina(n456), .dinb(n263), .dout(n457));
  jor  g0195(.dina(shift0 ), .dinb(a68 ), .dout(n458));
  jor  g0196(.dina(n269), .dinb(a67 ), .dout(n459));
  jand g0197(.dina(n459), .dinb(n458), .dout(n460));
  jor  g0198(.dina(n460), .dinb(shift1 ), .dout(n461));
  jor  g0199(.dina(shift0 ), .dinb(a66 ), .dout(n462));
  jor  g0200(.dina(n269), .dinb(a65 ), .dout(n463));
  jand g0201(.dina(n463), .dinb(n462), .dout(n464));
  jor  g0202(.dina(n464), .dinb(n273), .dout(n465));
  jand g0203(.dina(n465), .dinb(n461), .dout(n466));
  jand g0204(.dina(n466), .dinb(n292), .dout(n467));
  jor  g0205(.dina(shift0 ), .dinb(a72 ), .dout(n468));
  jor  g0206(.dina(n269), .dinb(a71 ), .dout(n469));
  jand g0207(.dina(n469), .dinb(n468), .dout(n470));
  jor  g0208(.dina(n470), .dinb(shift1 ), .dout(n471));
  jor  g0209(.dina(shift0 ), .dinb(a70 ), .dout(n472));
  jor  g0210(.dina(n269), .dinb(a69 ), .dout(n473));
  jand g0211(.dina(n473), .dinb(n472), .dout(n474));
  jor  g0212(.dina(n474), .dinb(n273), .dout(n475));
  jand g0213(.dina(n475), .dinb(n471), .dout(n476));
  jand g0214(.dina(n476), .dinb(n281), .dout(n477));
  jor  g0215(.dina(shift0 ), .dinb(a76 ), .dout(n478));
  jor  g0216(.dina(n269), .dinb(a75 ), .dout(n479));
  jand g0217(.dina(n479), .dinb(n478), .dout(n480));
  jor  g0218(.dina(n480), .dinb(shift1 ), .dout(n481));
  jor  g0219(.dina(shift0 ), .dinb(a74 ), .dout(n482));
  jor  g0220(.dina(n269), .dinb(a73 ), .dout(n483));
  jand g0221(.dina(n483), .dinb(n482), .dout(n484));
  jor  g0222(.dina(n484), .dinb(n273), .dout(n485));
  jand g0223(.dina(n485), .dinb(n481), .dout(n486));
  jand g0224(.dina(n486), .dinb(n267), .dout(n487));
  jor  g0225(.dina(n487), .dinb(n477), .dout(n488));
  jor  g0226(.dina(shift0 ), .dinb(a80 ), .dout(n489));
  jor  g0227(.dina(n269), .dinb(a79 ), .dout(n490));
  jand g0228(.dina(n490), .dinb(n489), .dout(n491));
  jor  g0229(.dina(n491), .dinb(shift1 ), .dout(n492));
  jor  g0230(.dina(shift0 ), .dinb(a78 ), .dout(n493));
  jor  g0231(.dina(n269), .dinb(a77 ), .dout(n494));
  jand g0232(.dina(n494), .dinb(n493), .dout(n495));
  jor  g0233(.dina(n495), .dinb(n273), .dout(n496));
  jand g0234(.dina(n496), .dinb(n492), .dout(n497));
  jand g0235(.dina(n497), .dinb(n304), .dout(n498));
  jor  g0236(.dina(n498), .dinb(n488), .dout(n499));
  jor  g0237(.dina(n499), .dinb(n467), .dout(n500));
  jand g0238(.dina(n500), .dinb(n410), .dout(n501));
  jor  g0239(.dina(shift0 ), .dinb(a100 ), .dout(n502));
  jor  g0240(.dina(n269), .dinb(a99 ), .dout(n503));
  jand g0241(.dina(n503), .dinb(n502), .dout(n504));
  jor  g0242(.dina(n504), .dinb(shift1 ), .dout(n505));
  jor  g0243(.dina(shift0 ), .dinb(a98 ), .dout(n506));
  jor  g0244(.dina(n269), .dinb(a97 ), .dout(n507));
  jand g0245(.dina(n507), .dinb(n506), .dout(n508));
  jor  g0246(.dina(n508), .dinb(n273), .dout(n509));
  jand g0247(.dina(n509), .dinb(n505), .dout(n510));
  jand g0248(.dina(n510), .dinb(n292), .dout(n511));
  jor  g0249(.dina(shift0 ), .dinb(a104 ), .dout(n512));
  jor  g0250(.dina(n269), .dinb(a103 ), .dout(n513));
  jand g0251(.dina(n513), .dinb(n512), .dout(n514));
  jor  g0252(.dina(n514), .dinb(shift1 ), .dout(n515));
  jor  g0253(.dina(shift0 ), .dinb(a102 ), .dout(n516));
  jor  g0254(.dina(n269), .dinb(a101 ), .dout(n517));
  jand g0255(.dina(n517), .dinb(n516), .dout(n518));
  jor  g0256(.dina(n518), .dinb(n273), .dout(n519));
  jand g0257(.dina(n519), .dinb(n515), .dout(n520));
  jand g0258(.dina(n520), .dinb(n281), .dout(n521));
  jor  g0259(.dina(shift0 ), .dinb(a108 ), .dout(n522));
  jor  g0260(.dina(n269), .dinb(a107 ), .dout(n523));
  jand g0261(.dina(n523), .dinb(n522), .dout(n524));
  jor  g0262(.dina(n524), .dinb(shift1 ), .dout(n525));
  jor  g0263(.dina(shift0 ), .dinb(a106 ), .dout(n526));
  jor  g0264(.dina(n269), .dinb(a105 ), .dout(n527));
  jand g0265(.dina(n527), .dinb(n526), .dout(n528));
  jor  g0266(.dina(n528), .dinb(n273), .dout(n529));
  jand g0267(.dina(n529), .dinb(n525), .dout(n530));
  jand g0268(.dina(n530), .dinb(n267), .dout(n531));
  jor  g0269(.dina(n531), .dinb(n521), .dout(n532));
  jor  g0270(.dina(shift0 ), .dinb(a112 ), .dout(n533));
  jor  g0271(.dina(n269), .dinb(a111 ), .dout(n534));
  jand g0272(.dina(n534), .dinb(n533), .dout(n535));
  jor  g0273(.dina(n535), .dinb(shift1 ), .dout(n536));
  jor  g0274(.dina(shift0 ), .dinb(a110 ), .dout(n537));
  jor  g0275(.dina(n269), .dinb(a109 ), .dout(n538));
  jand g0276(.dina(n538), .dinb(n537), .dout(n539));
  jor  g0277(.dina(n539), .dinb(n273), .dout(n540));
  jand g0278(.dina(n540), .dinb(n536), .dout(n541));
  jand g0279(.dina(n541), .dinb(n304), .dout(n542));
  jor  g0280(.dina(n542), .dinb(n532), .dout(n543));
  jor  g0281(.dina(n543), .dinb(n511), .dout(n544));
  jand g0282(.dina(n544), .dinb(n319), .dout(n545));
  jor  g0283(.dina(shift0 ), .dinb(a92 ), .dout(n546));
  jor  g0284(.dina(n269), .dinb(a91 ), .dout(n547));
  jand g0285(.dina(n547), .dinb(n546), .dout(n548));
  jor  g0286(.dina(n548), .dinb(shift1 ), .dout(n549));
  jor  g0287(.dina(shift0 ), .dinb(a90 ), .dout(n550));
  jor  g0288(.dina(n269), .dinb(a89 ), .dout(n551));
  jand g0289(.dina(n551), .dinb(n550), .dout(n552));
  jor  g0290(.dina(n552), .dinb(n273), .dout(n553));
  jand g0291(.dina(n553), .dinb(n549), .dout(n554));
  jand g0292(.dina(n554), .dinb(n267), .dout(n555));
  jor  g0293(.dina(shift0 ), .dinb(a88 ), .dout(n556));
  jor  g0294(.dina(n269), .dinb(a87 ), .dout(n557));
  jand g0295(.dina(n557), .dinb(n556), .dout(n558));
  jor  g0296(.dina(n558), .dinb(shift1 ), .dout(n559));
  jor  g0297(.dina(shift0 ), .dinb(a86 ), .dout(n560));
  jor  g0298(.dina(n269), .dinb(a85 ), .dout(n561));
  jand g0299(.dina(n561), .dinb(n560), .dout(n562));
  jor  g0300(.dina(n562), .dinb(n273), .dout(n563));
  jand g0301(.dina(n563), .dinb(n559), .dout(n564));
  jand g0302(.dina(n564), .dinb(n281), .dout(n565));
  jor  g0303(.dina(shift0 ), .dinb(a84 ), .dout(n566));
  jor  g0304(.dina(n269), .dinb(a83 ), .dout(n567));
  jand g0305(.dina(n567), .dinb(n566), .dout(n568));
  jor  g0306(.dina(n568), .dinb(shift1 ), .dout(n569));
  jor  g0307(.dina(shift0 ), .dinb(a82 ), .dout(n570));
  jor  g0308(.dina(n269), .dinb(a81 ), .dout(n571));
  jand g0309(.dina(n571), .dinb(n570), .dout(n572));
  jor  g0310(.dina(n572), .dinb(n273), .dout(n573));
  jand g0311(.dina(n573), .dinb(n569), .dout(n574));
  jand g0312(.dina(n574), .dinb(n292), .dout(n575));
  jor  g0313(.dina(n575), .dinb(n565), .dout(n576));
  jor  g0314(.dina(shift0 ), .dinb(a96 ), .dout(n577));
  jor  g0315(.dina(n269), .dinb(a95 ), .dout(n578));
  jand g0316(.dina(n578), .dinb(n577), .dout(n579));
  jor  g0317(.dina(n579), .dinb(shift1 ), .dout(n580));
  jor  g0318(.dina(shift0 ), .dinb(a94 ), .dout(n581));
  jor  g0319(.dina(n269), .dinb(a93 ), .dout(n582));
  jand g0320(.dina(n582), .dinb(n581), .dout(n583));
  jor  g0321(.dina(n583), .dinb(n273), .dout(n584));
  jand g0322(.dina(n584), .dinb(n580), .dout(n585));
  jand g0323(.dina(n585), .dinb(n304), .dout(n586));
  jor  g0324(.dina(n586), .dinb(n576), .dout(n587));
  jor  g0325(.dina(n587), .dinb(n555), .dout(n588));
  jand g0326(.dina(n588), .dinb(n265), .dout(n589));
  jor  g0327(.dina(n589), .dinb(n545), .dout(n590));
  jor  g0328(.dina(shift0 ), .dinb(a124 ), .dout(n591));
  jor  g0329(.dina(n269), .dinb(a123 ), .dout(n592));
  jand g0330(.dina(n592), .dinb(n591), .dout(n593));
  jor  g0331(.dina(n593), .dinb(shift1 ), .dout(n594));
  jor  g0332(.dina(shift0 ), .dinb(a122 ), .dout(n595));
  jor  g0333(.dina(n269), .dinb(a121 ), .dout(n596));
  jand g0334(.dina(n596), .dinb(n595), .dout(n597));
  jor  g0335(.dina(n597), .dinb(n273), .dout(n598));
  jand g0336(.dina(n598), .dinb(n594), .dout(n599));
  jand g0337(.dina(n599), .dinb(n267), .dout(n600));
  jor  g0338(.dina(shift0 ), .dinb(a120 ), .dout(n601));
  jor  g0339(.dina(n269), .dinb(a119 ), .dout(n602));
  jand g0340(.dina(n602), .dinb(n601), .dout(n603));
  jor  g0341(.dina(n603), .dinb(shift1 ), .dout(n604));
  jor  g0342(.dina(shift0 ), .dinb(a118 ), .dout(n605));
  jor  g0343(.dina(n269), .dinb(a117 ), .dout(n606));
  jand g0344(.dina(n606), .dinb(n605), .dout(n607));
  jor  g0345(.dina(n607), .dinb(n273), .dout(n608));
  jand g0346(.dina(n608), .dinb(n604), .dout(n609));
  jand g0347(.dina(n609), .dinb(n281), .dout(n610));
  jor  g0348(.dina(shift0 ), .dinb(a116 ), .dout(n611));
  jor  g0349(.dina(n269), .dinb(a115 ), .dout(n612));
  jand g0350(.dina(n612), .dinb(n611), .dout(n613));
  jor  g0351(.dina(n613), .dinb(shift1 ), .dout(n614));
  jor  g0352(.dina(shift0 ), .dinb(a114 ), .dout(n615));
  jor  g0353(.dina(n269), .dinb(a113 ), .dout(n616));
  jand g0354(.dina(n616), .dinb(n615), .dout(n617));
  jor  g0355(.dina(n617), .dinb(n273), .dout(n618));
  jand g0356(.dina(n618), .dinb(n614), .dout(n619));
  jand g0357(.dina(n619), .dinb(n292), .dout(n620));
  jor  g0358(.dina(n620), .dinb(n610), .dout(n621));
  jor  g0359(.dina(shift0 ), .dinb(a0 ), .dout(n622));
  jor  g0360(.dina(n269), .dinb(a127 ), .dout(n623));
  jand g0361(.dina(n623), .dinb(n622), .dout(n624));
  jor  g0362(.dina(n624), .dinb(shift1 ), .dout(n625));
  jor  g0363(.dina(shift0 ), .dinb(a126 ), .dout(n626));
  jor  g0364(.dina(n269), .dinb(a125 ), .dout(n627));
  jand g0365(.dina(n627), .dinb(n626), .dout(n628));
  jor  g0366(.dina(n628), .dinb(n273), .dout(n629));
  jand g0367(.dina(n629), .dinb(n625), .dout(n630));
  jand g0368(.dina(n630), .dinb(n304), .dout(n631));
  jor  g0369(.dina(n631), .dinb(n621), .dout(n632));
  jor  g0370(.dina(n632), .dinb(n600), .dout(n633));
  jand g0371(.dina(n633), .dinb(n364), .dout(n634));
  jor  g0372(.dina(n634), .dinb(n590), .dout(n635));
  jor  g0373(.dina(n635), .dinb(n501), .dout(n636));
  jor  g0374(.dina(n636), .dinb(shift6 ), .dout(n637));
  jand g0375(.dina(n637), .dinb(n457), .dout(result0 ));
  jor  g0376(.dina(shift0 ), .dinb(a61 ), .dout(n639));
  jor  g0377(.dina(n269), .dinb(a60 ), .dout(n640));
  jand g0378(.dina(n640), .dinb(n639), .dout(n641));
  jand g0379(.dina(n641), .dinb(n273), .dout(n642));
  jor  g0380(.dina(shift0 ), .dinb(a59 ), .dout(n643));
  jor  g0381(.dina(n269), .dinb(a58 ), .dout(n644));
  jand g0382(.dina(n644), .dinb(n643), .dout(n645));
  jand g0383(.dina(n645), .dinb(shift1 ), .dout(n646));
  jor  g0384(.dina(n646), .dinb(n642), .dout(n647));
  jand g0385(.dina(n647), .dinb(n267), .dout(n648));
  jor  g0386(.dina(shift0 ), .dinb(a57 ), .dout(n649));
  jor  g0387(.dina(n269), .dinb(a56 ), .dout(n650));
  jand g0388(.dina(n650), .dinb(n649), .dout(n651));
  jand g0389(.dina(n651), .dinb(n273), .dout(n652));
  jor  g0390(.dina(shift0 ), .dinb(a55 ), .dout(n653));
  jor  g0391(.dina(n269), .dinb(a54 ), .dout(n654));
  jand g0392(.dina(n654), .dinb(n653), .dout(n655));
  jand g0393(.dina(n655), .dinb(shift1 ), .dout(n656));
  jor  g0394(.dina(n656), .dinb(n652), .dout(n657));
  jand g0395(.dina(n657), .dinb(n281), .dout(n658));
  jor  g0396(.dina(shift0 ), .dinb(a53 ), .dout(n659));
  jor  g0397(.dina(n269), .dinb(a52 ), .dout(n660));
  jand g0398(.dina(n660), .dinb(n659), .dout(n661));
  jand g0399(.dina(n661), .dinb(n273), .dout(n662));
  jor  g0400(.dina(shift0 ), .dinb(a51 ), .dout(n663));
  jor  g0401(.dina(n269), .dinb(a50 ), .dout(n664));
  jand g0402(.dina(n664), .dinb(n663), .dout(n665));
  jand g0403(.dina(n665), .dinb(shift1 ), .dout(n666));
  jor  g0404(.dina(n666), .dinb(n662), .dout(n667));
  jand g0405(.dina(n667), .dinb(n292), .dout(n668));
  jor  g0406(.dina(n668), .dinb(n658), .dout(n669));
  jor  g0407(.dina(shift0 ), .dinb(a65 ), .dout(n670));
  jor  g0408(.dina(n269), .dinb(a64 ), .dout(n671));
  jand g0409(.dina(n671), .dinb(n670), .dout(n672));
  jand g0410(.dina(n672), .dinb(n273), .dout(n673));
  jor  g0411(.dina(shift0 ), .dinb(a63 ), .dout(n674));
  jor  g0412(.dina(n269), .dinb(a62 ), .dout(n675));
  jand g0413(.dina(n675), .dinb(n674), .dout(n676));
  jand g0414(.dina(n676), .dinb(shift1 ), .dout(n677));
  jor  g0415(.dina(n677), .dinb(n673), .dout(n678));
  jand g0416(.dina(n678), .dinb(n304), .dout(n679));
  jor  g0417(.dina(n679), .dinb(n669), .dout(n680));
  jor  g0418(.dina(n680), .dinb(n648), .dout(n681));
  jand g0419(.dina(n681), .dinb(n364), .dout(n682));
  jor  g0420(.dina(shift0 ), .dinb(a21 ), .dout(n683));
  jor  g0421(.dina(n269), .dinb(a20 ), .dout(n684));
  jand g0422(.dina(n684), .dinb(n683), .dout(n685));
  jand g0423(.dina(n685), .dinb(n273), .dout(n686));
  jor  g0424(.dina(shift0 ), .dinb(a19 ), .dout(n687));
  jor  g0425(.dina(n269), .dinb(a18 ), .dout(n688));
  jand g0426(.dina(n688), .dinb(n687), .dout(n689));
  jand g0427(.dina(n689), .dinb(shift1 ), .dout(n690));
  jor  g0428(.dina(n690), .dinb(n686), .dout(n691));
  jand g0429(.dina(n691), .dinb(n292), .dout(n692));
  jor  g0430(.dina(shift0 ), .dinb(a25 ), .dout(n693));
  jor  g0431(.dina(n269), .dinb(a24 ), .dout(n694));
  jand g0432(.dina(n694), .dinb(n693), .dout(n695));
  jand g0433(.dina(n695), .dinb(n273), .dout(n696));
  jor  g0434(.dina(shift0 ), .dinb(a23 ), .dout(n697));
  jor  g0435(.dina(n269), .dinb(a22 ), .dout(n698));
  jand g0436(.dina(n698), .dinb(n697), .dout(n699));
  jand g0437(.dina(n699), .dinb(shift1 ), .dout(n700));
  jor  g0438(.dina(n700), .dinb(n696), .dout(n701));
  jand g0439(.dina(n701), .dinb(n281), .dout(n702));
  jor  g0440(.dina(shift0 ), .dinb(a29 ), .dout(n703));
  jor  g0441(.dina(n269), .dinb(a28 ), .dout(n704));
  jand g0442(.dina(n704), .dinb(n703), .dout(n705));
  jand g0443(.dina(n705), .dinb(n273), .dout(n706));
  jor  g0444(.dina(shift0 ), .dinb(a27 ), .dout(n707));
  jor  g0445(.dina(n269), .dinb(a26 ), .dout(n708));
  jand g0446(.dina(n708), .dinb(n707), .dout(n709));
  jand g0447(.dina(n709), .dinb(shift1 ), .dout(n710));
  jor  g0448(.dina(n710), .dinb(n706), .dout(n711));
  jand g0449(.dina(n711), .dinb(n267), .dout(n712));
  jor  g0450(.dina(n712), .dinb(n702), .dout(n713));
  jor  g0451(.dina(shift0 ), .dinb(a33 ), .dout(n714));
  jor  g0452(.dina(n269), .dinb(a32 ), .dout(n715));
  jand g0453(.dina(n715), .dinb(n714), .dout(n716));
  jand g0454(.dina(n716), .dinb(n273), .dout(n717));
  jor  g0455(.dina(shift0 ), .dinb(a31 ), .dout(n718));
  jor  g0456(.dina(n269), .dinb(a30 ), .dout(n719));
  jand g0457(.dina(n719), .dinb(n718), .dout(n720));
  jand g0458(.dina(n720), .dinb(shift1 ), .dout(n721));
  jor  g0459(.dina(n721), .dinb(n717), .dout(n722));
  jand g0460(.dina(n722), .dinb(n304), .dout(n723));
  jor  g0461(.dina(n723), .dinb(n713), .dout(n724));
  jor  g0462(.dina(n724), .dinb(n692), .dout(n725));
  jand g0463(.dina(n725), .dinb(n265), .dout(n726));
  jor  g0464(.dina(shift0 ), .dinb(a17 ), .dout(n727));
  jor  g0465(.dina(n269), .dinb(a16 ), .dout(n728));
  jand g0466(.dina(n728), .dinb(n727), .dout(n729));
  jand g0467(.dina(n729), .dinb(n273), .dout(n730));
  jor  g0468(.dina(shift0 ), .dinb(a15 ), .dout(n731));
  jor  g0469(.dina(n269), .dinb(a14 ), .dout(n732));
  jand g0470(.dina(n732), .dinb(n731), .dout(n733));
  jand g0471(.dina(n733), .dinb(shift1 ), .dout(n734));
  jor  g0472(.dina(n734), .dinb(n730), .dout(n735));
  jand g0473(.dina(n735), .dinb(n304), .dout(n736));
  jor  g0474(.dina(shift0 ), .dinb(a9 ), .dout(n737));
  jor  g0475(.dina(n269), .dinb(a8 ), .dout(n738));
  jand g0476(.dina(n738), .dinb(n737), .dout(n739));
  jand g0477(.dina(n739), .dinb(n273), .dout(n740));
  jor  g0478(.dina(shift0 ), .dinb(a7 ), .dout(n741));
  jor  g0479(.dina(n269), .dinb(a6 ), .dout(n742));
  jand g0480(.dina(n742), .dinb(n741), .dout(n743));
  jand g0481(.dina(n743), .dinb(shift1 ), .dout(n744));
  jor  g0482(.dina(n744), .dinb(n740), .dout(n745));
  jand g0483(.dina(n745), .dinb(n281), .dout(n746));
  jor  g0484(.dina(shift0 ), .dinb(a5 ), .dout(n747));
  jor  g0485(.dina(n269), .dinb(a4 ), .dout(n748));
  jand g0486(.dina(n748), .dinb(n747), .dout(n749));
  jand g0487(.dina(n749), .dinb(n273), .dout(n750));
  jor  g0488(.dina(shift0 ), .dinb(a3 ), .dout(n751));
  jor  g0489(.dina(n269), .dinb(a2 ), .dout(n752));
  jand g0490(.dina(n752), .dinb(n751), .dout(n753));
  jand g0491(.dina(n753), .dinb(shift1 ), .dout(n754));
  jor  g0492(.dina(n754), .dinb(n750), .dout(n755));
  jand g0493(.dina(n755), .dinb(n292), .dout(n756));
  jor  g0494(.dina(n756), .dinb(n746), .dout(n757));
  jor  g0495(.dina(shift0 ), .dinb(a13 ), .dout(n758));
  jor  g0496(.dina(n269), .dinb(a12 ), .dout(n759));
  jand g0497(.dina(n759), .dinb(n758), .dout(n760));
  jand g0498(.dina(n760), .dinb(n273), .dout(n761));
  jor  g0499(.dina(shift0 ), .dinb(a11 ), .dout(n762));
  jor  g0500(.dina(n269), .dinb(a10 ), .dout(n763));
  jand g0501(.dina(n763), .dinb(n762), .dout(n764));
  jand g0502(.dina(n764), .dinb(shift1 ), .dout(n765));
  jor  g0503(.dina(n765), .dinb(n761), .dout(n766));
  jand g0504(.dina(n766), .dinb(n267), .dout(n767));
  jor  g0505(.dina(n767), .dinb(n757), .dout(n768));
  jor  g0506(.dina(n768), .dinb(n736), .dout(n769));
  jand g0507(.dina(n769), .dinb(n410), .dout(n770));
  jor  g0508(.dina(n770), .dinb(n726), .dout(n771));
  jor  g0509(.dina(shift0 ), .dinb(a37 ), .dout(n772));
  jor  g0510(.dina(n269), .dinb(a36 ), .dout(n773));
  jand g0511(.dina(n773), .dinb(n772), .dout(n774));
  jand g0512(.dina(n774), .dinb(n273), .dout(n775));
  jor  g0513(.dina(shift0 ), .dinb(a35 ), .dout(n776));
  jor  g0514(.dina(n269), .dinb(a34 ), .dout(n777));
  jand g0515(.dina(n777), .dinb(n776), .dout(n778));
  jand g0516(.dina(n778), .dinb(shift1 ), .dout(n779));
  jor  g0517(.dina(n779), .dinb(n775), .dout(n780));
  jand g0518(.dina(n780), .dinb(n292), .dout(n781));
  jor  g0519(.dina(shift0 ), .dinb(a39 ), .dout(n782));
  jor  g0520(.dina(n269), .dinb(a38 ), .dout(n783));
  jand g0521(.dina(n783), .dinb(n782), .dout(n784));
  jor  g0522(.dina(n784), .dinb(n273), .dout(n785));
  jor  g0523(.dina(shift0 ), .dinb(a41 ), .dout(n786));
  jor  g0524(.dina(n269), .dinb(a40 ), .dout(n787));
  jand g0525(.dina(n787), .dinb(n786), .dout(n788));
  jor  g0526(.dina(n788), .dinb(shift1 ), .dout(n789));
  jand g0527(.dina(n789), .dinb(n785), .dout(n790));
  jand g0528(.dina(n790), .dinb(n281), .dout(n791));
  jor  g0529(.dina(shift0 ), .dinb(a45 ), .dout(n792));
  jor  g0530(.dina(n269), .dinb(a44 ), .dout(n793));
  jand g0531(.dina(n793), .dinb(n792), .dout(n794));
  jor  g0532(.dina(n794), .dinb(shift1 ), .dout(n795));
  jor  g0533(.dina(shift0 ), .dinb(a43 ), .dout(n796));
  jor  g0534(.dina(n269), .dinb(a42 ), .dout(n797));
  jand g0535(.dina(n797), .dinb(n796), .dout(n798));
  jor  g0536(.dina(n798), .dinb(n273), .dout(n799));
  jand g0537(.dina(n799), .dinb(n795), .dout(n800));
  jand g0538(.dina(n800), .dinb(n267), .dout(n801));
  jor  g0539(.dina(n801), .dinb(n791), .dout(n802));
  jor  g0540(.dina(shift0 ), .dinb(a49 ), .dout(n803));
  jor  g0541(.dina(n269), .dinb(a48 ), .dout(n804));
  jand g0542(.dina(n804), .dinb(n803), .dout(n805));
  jand g0543(.dina(n805), .dinb(n273), .dout(n806));
  jor  g0544(.dina(shift0 ), .dinb(a47 ), .dout(n807));
  jor  g0545(.dina(n269), .dinb(a46 ), .dout(n808));
  jand g0546(.dina(n808), .dinb(n807), .dout(n809));
  jand g0547(.dina(n809), .dinb(shift1 ), .dout(n810));
  jor  g0548(.dina(n810), .dinb(n806), .dout(n811));
  jand g0549(.dina(n811), .dinb(n304), .dout(n812));
  jor  g0550(.dina(n812), .dinb(n802), .dout(n813));
  jor  g0551(.dina(n813), .dinb(n781), .dout(n814));
  jand g0552(.dina(n814), .dinb(n319), .dout(n815));
  jor  g0553(.dina(n815), .dinb(n771), .dout(n816));
  jor  g0554(.dina(n816), .dinb(n682), .dout(n817));
  jor  g0555(.dina(n817), .dinb(n263), .dout(n818));
  jor  g0556(.dina(shift0 ), .dinb(a69 ), .dout(n819));
  jor  g0557(.dina(n269), .dinb(a68 ), .dout(n820));
  jand g0558(.dina(n820), .dinb(n819), .dout(n821));
  jand g0559(.dina(n821), .dinb(n273), .dout(n822));
  jor  g0560(.dina(shift0 ), .dinb(a67 ), .dout(n823));
  jor  g0561(.dina(n269), .dinb(a66 ), .dout(n824));
  jand g0562(.dina(n824), .dinb(n823), .dout(n825));
  jand g0563(.dina(n825), .dinb(shift1 ), .dout(n826));
  jor  g0564(.dina(n826), .dinb(n822), .dout(n827));
  jand g0565(.dina(n827), .dinb(n292), .dout(n828));
  jor  g0566(.dina(shift0 ), .dinb(a73 ), .dout(n829));
  jor  g0567(.dina(n269), .dinb(a72 ), .dout(n830));
  jand g0568(.dina(n830), .dinb(n829), .dout(n831));
  jand g0569(.dina(n831), .dinb(n273), .dout(n832));
  jor  g0570(.dina(shift0 ), .dinb(a71 ), .dout(n833));
  jor  g0571(.dina(n269), .dinb(a70 ), .dout(n834));
  jand g0572(.dina(n834), .dinb(n833), .dout(n835));
  jand g0573(.dina(n835), .dinb(shift1 ), .dout(n836));
  jor  g0574(.dina(n836), .dinb(n832), .dout(n837));
  jand g0575(.dina(n837), .dinb(n281), .dout(n838));
  jor  g0576(.dina(shift0 ), .dinb(a77 ), .dout(n839));
  jor  g0577(.dina(n269), .dinb(a76 ), .dout(n840));
  jand g0578(.dina(n840), .dinb(n839), .dout(n841));
  jand g0579(.dina(n841), .dinb(n273), .dout(n842));
  jor  g0580(.dina(shift0 ), .dinb(a75 ), .dout(n843));
  jor  g0581(.dina(n269), .dinb(a74 ), .dout(n844));
  jand g0582(.dina(n844), .dinb(n843), .dout(n845));
  jand g0583(.dina(n845), .dinb(shift1 ), .dout(n846));
  jor  g0584(.dina(n846), .dinb(n842), .dout(n847));
  jand g0585(.dina(n847), .dinb(n267), .dout(n848));
  jor  g0586(.dina(n848), .dinb(n838), .dout(n849));
  jor  g0587(.dina(shift0 ), .dinb(a81 ), .dout(n850));
  jor  g0588(.dina(n269), .dinb(a80 ), .dout(n851));
  jand g0589(.dina(n851), .dinb(n850), .dout(n852));
  jand g0590(.dina(n852), .dinb(n273), .dout(n853));
  jor  g0591(.dina(shift0 ), .dinb(a79 ), .dout(n854));
  jor  g0592(.dina(n269), .dinb(a78 ), .dout(n855));
  jand g0593(.dina(n855), .dinb(n854), .dout(n856));
  jand g0594(.dina(n856), .dinb(shift1 ), .dout(n857));
  jor  g0595(.dina(n857), .dinb(n853), .dout(n858));
  jand g0596(.dina(n858), .dinb(n304), .dout(n859));
  jor  g0597(.dina(n859), .dinb(n849), .dout(n860));
  jor  g0598(.dina(n860), .dinb(n828), .dout(n861));
  jand g0599(.dina(n861), .dinb(n410), .dout(n862));
  jor  g0600(.dina(shift0 ), .dinb(a101 ), .dout(n863));
  jor  g0601(.dina(n269), .dinb(a100 ), .dout(n864));
  jand g0602(.dina(n864), .dinb(n863), .dout(n865));
  jand g0603(.dina(n865), .dinb(n273), .dout(n866));
  jor  g0604(.dina(shift0 ), .dinb(a99 ), .dout(n867));
  jor  g0605(.dina(n269), .dinb(a98 ), .dout(n868));
  jand g0606(.dina(n868), .dinb(n867), .dout(n869));
  jand g0607(.dina(n869), .dinb(shift1 ), .dout(n870));
  jor  g0608(.dina(n870), .dinb(n866), .dout(n871));
  jand g0609(.dina(n871), .dinb(n292), .dout(n872));
  jor  g0610(.dina(shift0 ), .dinb(a105 ), .dout(n873));
  jor  g0611(.dina(n269), .dinb(a104 ), .dout(n874));
  jand g0612(.dina(n874), .dinb(n873), .dout(n875));
  jand g0613(.dina(n875), .dinb(n273), .dout(n876));
  jor  g0614(.dina(shift0 ), .dinb(a103 ), .dout(n877));
  jor  g0615(.dina(n269), .dinb(a102 ), .dout(n878));
  jand g0616(.dina(n878), .dinb(n877), .dout(n879));
  jand g0617(.dina(n879), .dinb(shift1 ), .dout(n880));
  jor  g0618(.dina(n880), .dinb(n876), .dout(n881));
  jand g0619(.dina(n881), .dinb(n281), .dout(n882));
  jor  g0620(.dina(shift0 ), .dinb(a109 ), .dout(n883));
  jor  g0621(.dina(n269), .dinb(a108 ), .dout(n884));
  jand g0622(.dina(n884), .dinb(n883), .dout(n885));
  jand g0623(.dina(n885), .dinb(n273), .dout(n886));
  jor  g0624(.dina(shift0 ), .dinb(a107 ), .dout(n887));
  jor  g0625(.dina(n269), .dinb(a106 ), .dout(n888));
  jand g0626(.dina(n888), .dinb(n887), .dout(n889));
  jand g0627(.dina(n889), .dinb(shift1 ), .dout(n890));
  jor  g0628(.dina(n890), .dinb(n886), .dout(n891));
  jand g0629(.dina(n891), .dinb(n267), .dout(n892));
  jor  g0630(.dina(n892), .dinb(n882), .dout(n893));
  jor  g0631(.dina(shift0 ), .dinb(a113 ), .dout(n894));
  jor  g0632(.dina(n269), .dinb(a112 ), .dout(n895));
  jand g0633(.dina(n895), .dinb(n894), .dout(n896));
  jand g0634(.dina(n896), .dinb(n273), .dout(n897));
  jor  g0635(.dina(shift0 ), .dinb(a111 ), .dout(n898));
  jor  g0636(.dina(n269), .dinb(a110 ), .dout(n899));
  jand g0637(.dina(n899), .dinb(n898), .dout(n900));
  jand g0638(.dina(n900), .dinb(shift1 ), .dout(n901));
  jor  g0639(.dina(n901), .dinb(n897), .dout(n902));
  jand g0640(.dina(n902), .dinb(n304), .dout(n903));
  jor  g0641(.dina(n903), .dinb(n893), .dout(n904));
  jor  g0642(.dina(n904), .dinb(n872), .dout(n905));
  jand g0643(.dina(n905), .dinb(n319), .dout(n906));
  jor  g0644(.dina(shift0 ), .dinb(a85 ), .dout(n907));
  jor  g0645(.dina(n269), .dinb(a84 ), .dout(n908));
  jand g0646(.dina(n908), .dinb(n907), .dout(n909));
  jand g0647(.dina(n909), .dinb(n273), .dout(n910));
  jor  g0648(.dina(shift0 ), .dinb(a83 ), .dout(n911));
  jor  g0649(.dina(n269), .dinb(a82 ), .dout(n912));
  jand g0650(.dina(n912), .dinb(n911), .dout(n913));
  jand g0651(.dina(n913), .dinb(shift1 ), .dout(n914));
  jor  g0652(.dina(n914), .dinb(n910), .dout(n915));
  jand g0653(.dina(n915), .dinb(n292), .dout(n916));
  jor  g0654(.dina(shift0 ), .dinb(a89 ), .dout(n917));
  jor  g0655(.dina(n269), .dinb(a88 ), .dout(n918));
  jand g0656(.dina(n918), .dinb(n917), .dout(n919));
  jand g0657(.dina(n919), .dinb(n273), .dout(n920));
  jor  g0658(.dina(shift0 ), .dinb(a87 ), .dout(n921));
  jor  g0659(.dina(n269), .dinb(a86 ), .dout(n922));
  jand g0660(.dina(n922), .dinb(n921), .dout(n923));
  jand g0661(.dina(n923), .dinb(shift1 ), .dout(n924));
  jor  g0662(.dina(n924), .dinb(n920), .dout(n925));
  jand g0663(.dina(n925), .dinb(n281), .dout(n926));
  jor  g0664(.dina(shift0 ), .dinb(a93 ), .dout(n927));
  jor  g0665(.dina(n269), .dinb(a92 ), .dout(n928));
  jand g0666(.dina(n928), .dinb(n927), .dout(n929));
  jand g0667(.dina(n929), .dinb(n273), .dout(n930));
  jor  g0668(.dina(shift0 ), .dinb(a91 ), .dout(n931));
  jor  g0669(.dina(n269), .dinb(a90 ), .dout(n932));
  jand g0670(.dina(n932), .dinb(n931), .dout(n933));
  jand g0671(.dina(n933), .dinb(shift1 ), .dout(n934));
  jor  g0672(.dina(n934), .dinb(n930), .dout(n935));
  jand g0673(.dina(n935), .dinb(n267), .dout(n936));
  jor  g0674(.dina(n936), .dinb(n926), .dout(n937));
  jor  g0675(.dina(shift0 ), .dinb(a97 ), .dout(n938));
  jor  g0676(.dina(n269), .dinb(a96 ), .dout(n939));
  jand g0677(.dina(n939), .dinb(n938), .dout(n940));
  jand g0678(.dina(n940), .dinb(n273), .dout(n941));
  jor  g0679(.dina(shift0 ), .dinb(a95 ), .dout(n942));
  jor  g0680(.dina(n269), .dinb(a94 ), .dout(n943));
  jand g0681(.dina(n943), .dinb(n942), .dout(n944));
  jand g0682(.dina(n944), .dinb(shift1 ), .dout(n945));
  jor  g0683(.dina(n945), .dinb(n941), .dout(n946));
  jand g0684(.dina(n946), .dinb(n304), .dout(n947));
  jor  g0685(.dina(n947), .dinb(n937), .dout(n948));
  jor  g0686(.dina(n948), .dinb(n916), .dout(n949));
  jand g0687(.dina(n949), .dinb(n265), .dout(n950));
  jor  g0688(.dina(n950), .dinb(n906), .dout(n951));
  jor  g0689(.dina(shift0 ), .dinb(a125 ), .dout(n952));
  jor  g0690(.dina(n269), .dinb(a124 ), .dout(n953));
  jand g0691(.dina(n953), .dinb(n952), .dout(n954));
  jand g0692(.dina(n954), .dinb(n273), .dout(n955));
  jor  g0693(.dina(shift0 ), .dinb(a123 ), .dout(n956));
  jor  g0694(.dina(n269), .dinb(a122 ), .dout(n957));
  jand g0695(.dina(n957), .dinb(n956), .dout(n958));
  jand g0696(.dina(n958), .dinb(shift1 ), .dout(n959));
  jor  g0697(.dina(n959), .dinb(n955), .dout(n960));
  jand g0698(.dina(n960), .dinb(n267), .dout(n961));
  jor  g0699(.dina(shift0 ), .dinb(a121 ), .dout(n962));
  jor  g0700(.dina(n269), .dinb(a120 ), .dout(n963));
  jand g0701(.dina(n963), .dinb(n962), .dout(n964));
  jand g0702(.dina(n964), .dinb(n273), .dout(n965));
  jor  g0703(.dina(shift0 ), .dinb(a119 ), .dout(n966));
  jor  g0704(.dina(n269), .dinb(a118 ), .dout(n967));
  jand g0705(.dina(n967), .dinb(n966), .dout(n968));
  jand g0706(.dina(n968), .dinb(shift1 ), .dout(n969));
  jor  g0707(.dina(n969), .dinb(n965), .dout(n970));
  jand g0708(.dina(n970), .dinb(n281), .dout(n971));
  jor  g0709(.dina(shift0 ), .dinb(a117 ), .dout(n972));
  jor  g0710(.dina(n269), .dinb(a116 ), .dout(n973));
  jand g0711(.dina(n973), .dinb(n972), .dout(n974));
  jand g0712(.dina(n974), .dinb(n273), .dout(n975));
  jor  g0713(.dina(shift0 ), .dinb(a115 ), .dout(n976));
  jor  g0714(.dina(n269), .dinb(a114 ), .dout(n977));
  jand g0715(.dina(n977), .dinb(n976), .dout(n978));
  jand g0716(.dina(n978), .dinb(shift1 ), .dout(n979));
  jor  g0717(.dina(n979), .dinb(n975), .dout(n980));
  jand g0718(.dina(n980), .dinb(n292), .dout(n981));
  jor  g0719(.dina(n981), .dinb(n971), .dout(n982));
  jor  g0720(.dina(shift0 ), .dinb(a1 ), .dout(n983));
  jor  g0721(.dina(n269), .dinb(a0 ), .dout(n984));
  jand g0722(.dina(n984), .dinb(n983), .dout(n985));
  jand g0723(.dina(n985), .dinb(n273), .dout(n986));
  jor  g0724(.dina(shift0 ), .dinb(a127 ), .dout(n987));
  jor  g0725(.dina(n269), .dinb(a126 ), .dout(n988));
  jand g0726(.dina(n988), .dinb(n987), .dout(n989));
  jand g0727(.dina(n989), .dinb(shift1 ), .dout(n990));
  jor  g0728(.dina(n990), .dinb(n986), .dout(n991));
  jand g0729(.dina(n991), .dinb(n304), .dout(n992));
  jor  g0730(.dina(n992), .dinb(n982), .dout(n993));
  jor  g0731(.dina(n993), .dinb(n961), .dout(n994));
  jand g0732(.dina(n994), .dinb(n364), .dout(n995));
  jor  g0733(.dina(n995), .dinb(n951), .dout(n996));
  jor  g0734(.dina(n996), .dinb(n862), .dout(n997));
  jor  g0735(.dina(n997), .dinb(shift6 ), .dout(n998));
  jand g0736(.dina(n998), .dinb(n818), .dout(result1 ));
  jor  g0737(.dina(n357), .dinb(shift1 ), .dout(n1000));
  jor  g0738(.dina(n342), .dinb(n273), .dout(n1001));
  jand g0739(.dina(n1001), .dinb(n1000), .dout(n1002));
  jand g0740(.dina(n1002), .dinb(n267), .dout(n1003));
  jor  g0741(.dina(n332), .dinb(n273), .dout(n1004));
  jor  g0742(.dina(n346), .dinb(shift1 ), .dout(n1005));
  jand g0743(.dina(n1005), .dinb(n1004), .dout(n1006));
  jand g0744(.dina(n1006), .dinb(n281), .dout(n1007));
  jor  g0745(.dina(n322), .dinb(n273), .dout(n1008));
  jor  g0746(.dina(n336), .dinb(shift1 ), .dout(n1009));
  jand g0747(.dina(n1009), .dinb(n1008), .dout(n1010));
  jand g0748(.dina(n1010), .dinb(n292), .dout(n1011));
  jor  g0749(.dina(n1011), .dinb(n1007), .dout(n1012));
  jor  g0750(.dina(n353), .dinb(n273), .dout(n1013));
  jor  g0751(.dina(n402), .dinb(shift1 ), .dout(n1014));
  jand g0752(.dina(n1014), .dinb(n1013), .dout(n1015));
  jand g0753(.dina(n1015), .dinb(n304), .dout(n1016));
  jor  g0754(.dina(n1016), .dinb(n1012), .dout(n1017));
  jor  g0755(.dina(n1017), .dinb(n1003), .dout(n1018));
  jand g0756(.dina(n1018), .dinb(n319), .dout(n1019));
  jor  g0757(.dina(n295), .dinb(n273), .dout(n1020));
  jor  g0758(.dina(n288), .dinb(shift1 ), .dout(n1021));
  jand g0759(.dina(n1021), .dinb(n1020), .dout(n1022));
  jand g0760(.dina(n1022), .dinb(n292), .dout(n1023));
  jor  g0761(.dina(n284), .dinb(n273), .dout(n1024));
  jor  g0762(.dina(n276), .dinb(shift1 ), .dout(n1025));
  jand g0763(.dina(n1025), .dinb(n1024), .dout(n1026));
  jand g0764(.dina(n1026), .dinb(n281), .dout(n1027));
  jor  g0765(.dina(n271), .dinb(n273), .dout(n1028));
  jor  g0766(.dina(n311), .dinb(shift1 ), .dout(n1029));
  jand g0767(.dina(n1029), .dinb(n1028), .dout(n1030));
  jand g0768(.dina(n1030), .dinb(n267), .dout(n1031));
  jor  g0769(.dina(n1031), .dinb(n1027), .dout(n1032));
  jor  g0770(.dina(n307), .dinb(n273), .dout(n1033));
  jor  g0771(.dina(n326), .dinb(shift1 ), .dout(n1034));
  jand g0772(.dina(n1034), .dinb(n1033), .dout(n1035));
  jand g0773(.dina(n1035), .dinb(n304), .dout(n1036));
  jor  g0774(.dina(n1036), .dinb(n1032), .dout(n1037));
  jor  g0775(.dina(n1037), .dinb(n1023), .dout(n1038));
  jand g0776(.dina(n1038), .dinb(n265), .dout(n1039));
  jor  g0777(.dina(n444), .dinb(n273), .dout(n1040));
  jor  g0778(.dina(n299), .dinb(shift1 ), .dout(n1041));
  jand g0779(.dina(n1041), .dinb(n1040), .dout(n1042));
  jand g0780(.dina(n1042), .dinb(n304), .dout(n1043));
  jor  g0781(.dina(n423), .dinb(n273), .dout(n1044));
  jor  g0782(.dina(n417), .dinb(shift1 ), .dout(n1045));
  jand g0783(.dina(n1045), .dinb(n1044), .dout(n1046));
  jand g0784(.dina(n1046), .dinb(n281), .dout(n1047));
  jor  g0785(.dina(n413), .dinb(n273), .dout(n1048));
  jor  g0786(.dina(n448), .dinb(shift1 ), .dout(n1049));
  jand g0787(.dina(n1049), .dinb(n1048), .dout(n1050));
  jand g0788(.dina(n1050), .dinb(n267), .dout(n1051));
  jor  g0789(.dina(n1051), .dinb(n1047), .dout(n1052));
  jor  g0790(.dina(n433), .dinb(n273), .dout(n1053));
  jor  g0791(.dina(n427), .dinb(shift1 ), .dout(n1054));
  jand g0792(.dina(n1054), .dinb(n1053), .dout(n1055));
  jand g0793(.dina(n1055), .dinb(n292), .dout(n1056));
  jor  g0794(.dina(n1056), .dinb(n1052), .dout(n1057));
  jor  g0795(.dina(n1057), .dinb(n1043), .dout(n1058));
  jand g0796(.dina(n1058), .dinb(n410), .dout(n1059));
  jor  g0797(.dina(n1059), .dinb(n1039), .dout(n1060));
  jor  g0798(.dina(n398), .dinb(n273), .dout(n1061));
  jor  g0799(.dina(n381), .dinb(shift1 ), .dout(n1062));
  jand g0800(.dina(n1062), .dinb(n1061), .dout(n1063));
  jand g0801(.dina(n1063), .dinb(n292), .dout(n1064));
  jor  g0802(.dina(n377), .dinb(n273), .dout(n1065));
  jor  g0803(.dina(n391), .dinb(shift1 ), .dout(n1066));
  jand g0804(.dina(n1066), .dinb(n1065), .dout(n1067));
  jand g0805(.dina(n1067), .dinb(n281), .dout(n1068));
  jor  g0806(.dina(n387), .dinb(n273), .dout(n1069));
  jor  g0807(.dina(n371), .dinb(shift1 ), .dout(n1070));
  jand g0808(.dina(n1070), .dinb(n1069), .dout(n1071));
  jand g0809(.dina(n1071), .dinb(n267), .dout(n1072));
  jor  g0810(.dina(n1072), .dinb(n1068), .dout(n1073));
  jor  g0811(.dina(n367), .dinb(n273), .dout(n1074));
  jor  g0812(.dina(n464), .dinb(shift1 ), .dout(n1075));
  jand g0813(.dina(n1075), .dinb(n1074), .dout(n1076));
  jand g0814(.dina(n1076), .dinb(n304), .dout(n1077));
  jor  g0815(.dina(n1077), .dinb(n1073), .dout(n1078));
  jor  g0816(.dina(n1078), .dinb(n1064), .dout(n1079));
  jand g0817(.dina(n1079), .dinb(n364), .dout(n1080));
  jor  g0818(.dina(n1080), .dinb(n1060), .dout(n1081));
  jor  g0819(.dina(n1081), .dinb(n1019), .dout(n1082));
  jor  g0820(.dina(n1082), .dinb(n263), .dout(n1083));
  jor  g0821(.dina(n480), .dinb(n273), .dout(n1084));
  jor  g0822(.dina(n495), .dinb(shift1 ), .dout(n1085));
  jand g0823(.dina(n1085), .dinb(n1084), .dout(n1086));
  jand g0824(.dina(n1086), .dinb(n267), .dout(n1087));
  jor  g0825(.dina(n470), .dinb(n273), .dout(n1088));
  jor  g0826(.dina(n484), .dinb(shift1 ), .dout(n1089));
  jand g0827(.dina(n1089), .dinb(n1088), .dout(n1090));
  jand g0828(.dina(n1090), .dinb(n281), .dout(n1091));
  jor  g0829(.dina(n460), .dinb(n273), .dout(n1092));
  jor  g0830(.dina(n474), .dinb(shift1 ), .dout(n1093));
  jand g0831(.dina(n1093), .dinb(n1092), .dout(n1094));
  jand g0832(.dina(n1094), .dinb(n292), .dout(n1095));
  jor  g0833(.dina(n1095), .dinb(n1091), .dout(n1096));
  jor  g0834(.dina(n491), .dinb(n273), .dout(n1097));
  jor  g0835(.dina(n572), .dinb(shift1 ), .dout(n1098));
  jand g0836(.dina(n1098), .dinb(n1097), .dout(n1099));
  jand g0837(.dina(n1099), .dinb(n304), .dout(n1100));
  jor  g0838(.dina(n1100), .dinb(n1096), .dout(n1101));
  jor  g0839(.dina(n1101), .dinb(n1087), .dout(n1102));
  jand g0840(.dina(n1102), .dinb(n410), .dout(n1103));
  jor  g0841(.dina(n535), .dinb(n273), .dout(n1104));
  jor  g0842(.dina(n617), .dinb(shift1 ), .dout(n1105));
  jand g0843(.dina(n1105), .dinb(n1104), .dout(n1106));
  jand g0844(.dina(n1106), .dinb(n304), .dout(n1107));
  jor  g0845(.dina(n514), .dinb(n273), .dout(n1108));
  jor  g0846(.dina(n528), .dinb(shift1 ), .dout(n1109));
  jand g0847(.dina(n1109), .dinb(n1108), .dout(n1110));
  jand g0848(.dina(n1110), .dinb(n281), .dout(n1111));
  jor  g0849(.dina(n504), .dinb(n273), .dout(n1112));
  jor  g0850(.dina(n518), .dinb(shift1 ), .dout(n1113));
  jand g0851(.dina(n1113), .dinb(n1112), .dout(n1114));
  jand g0852(.dina(n1114), .dinb(n292), .dout(n1115));
  jor  g0853(.dina(n1115), .dinb(n1111), .dout(n1116));
  jor  g0854(.dina(n524), .dinb(n273), .dout(n1117));
  jor  g0855(.dina(n539), .dinb(shift1 ), .dout(n1118));
  jand g0856(.dina(n1118), .dinb(n1117), .dout(n1119));
  jand g0857(.dina(n1119), .dinb(n267), .dout(n1120));
  jor  g0858(.dina(n1120), .dinb(n1116), .dout(n1121));
  jor  g0859(.dina(n1121), .dinb(n1107), .dout(n1122));
  jand g0860(.dina(n1122), .dinb(n319), .dout(n1123));
  jor  g0861(.dina(n624), .dinb(n273), .dout(n1124));
  jor  g0862(.dina(n437), .dinb(shift1 ), .dout(n1125));
  jand g0863(.dina(n1125), .dinb(n1124), .dout(n1126));
  jand g0864(.dina(n1126), .dinb(n304), .dout(n1127));
  jor  g0865(.dina(n603), .dinb(n273), .dout(n1128));
  jor  g0866(.dina(n597), .dinb(shift1 ), .dout(n1129));
  jand g0867(.dina(n1129), .dinb(n1128), .dout(n1130));
  jand g0868(.dina(n1130), .dinb(n281), .dout(n1131));
  jor  g0869(.dina(n593), .dinb(n273), .dout(n1132));
  jor  g0870(.dina(n628), .dinb(shift1 ), .dout(n1133));
  jand g0871(.dina(n1133), .dinb(n1132), .dout(n1134));
  jand g0872(.dina(n1134), .dinb(n267), .dout(n1135));
  jor  g0873(.dina(n1135), .dinb(n1131), .dout(n1136));
  jor  g0874(.dina(n613), .dinb(n273), .dout(n1137));
  jor  g0875(.dina(n607), .dinb(shift1 ), .dout(n1138));
  jand g0876(.dina(n1138), .dinb(n1137), .dout(n1139));
  jand g0877(.dina(n1139), .dinb(n292), .dout(n1140));
  jor  g0878(.dina(n1140), .dinb(n1136), .dout(n1141));
  jor  g0879(.dina(n1141), .dinb(n1127), .dout(n1142));
  jand g0880(.dina(n1142), .dinb(n364), .dout(n1143));
  jor  g0881(.dina(n1143), .dinb(n1123), .dout(n1144));
  jor  g0882(.dina(n568), .dinb(n273), .dout(n1145));
  jor  g0883(.dina(n562), .dinb(shift1 ), .dout(n1146));
  jand g0884(.dina(n1146), .dinb(n1145), .dout(n1147));
  jand g0885(.dina(n1147), .dinb(n292), .dout(n1148));
  jor  g0886(.dina(n558), .dinb(n273), .dout(n1149));
  jor  g0887(.dina(n552), .dinb(shift1 ), .dout(n1150));
  jand g0888(.dina(n1150), .dinb(n1149), .dout(n1151));
  jand g0889(.dina(n1151), .dinb(n281), .dout(n1152));
  jor  g0890(.dina(n548), .dinb(n273), .dout(n1153));
  jor  g0891(.dina(n583), .dinb(shift1 ), .dout(n1154));
  jand g0892(.dina(n1154), .dinb(n1153), .dout(n1155));
  jand g0893(.dina(n1155), .dinb(n267), .dout(n1156));
  jor  g0894(.dina(n1156), .dinb(n1152), .dout(n1157));
  jor  g0895(.dina(n579), .dinb(n273), .dout(n1158));
  jor  g0896(.dina(n508), .dinb(shift1 ), .dout(n1159));
  jand g0897(.dina(n1159), .dinb(n1158), .dout(n1160));
  jand g0898(.dina(n1160), .dinb(n304), .dout(n1161));
  jor  g0899(.dina(n1161), .dinb(n1157), .dout(n1162));
  jor  g0900(.dina(n1162), .dinb(n1148), .dout(n1163));
  jand g0901(.dina(n1163), .dinb(n265), .dout(n1164));
  jor  g0902(.dina(n1164), .dinb(n1144), .dout(n1165));
  jor  g0903(.dina(n1165), .dinb(n1103), .dout(n1166));
  jor  g0904(.dina(n1166), .dinb(shift6 ), .dout(n1167));
  jand g0905(.dina(n1167), .dinb(n1083), .dout(result2 ));
  jand g0906(.dina(n661), .dinb(shift1 ), .dout(n1169));
  jand g0907(.dina(n655), .dinb(n273), .dout(n1170));
  jor  g0908(.dina(n1170), .dinb(n1169), .dout(n1171));
  jand g0909(.dina(n1171), .dinb(n292), .dout(n1172));
  jand g0910(.dina(n651), .dinb(shift1 ), .dout(n1173));
  jand g0911(.dina(n645), .dinb(n273), .dout(n1174));
  jor  g0912(.dina(n1174), .dinb(n1173), .dout(n1175));
  jand g0913(.dina(n1175), .dinb(n281), .dout(n1176));
  jand g0914(.dina(n641), .dinb(shift1 ), .dout(n1177));
  jand g0915(.dina(n676), .dinb(n273), .dout(n1178));
  jor  g0916(.dina(n1178), .dinb(n1177), .dout(n1179));
  jand g0917(.dina(n1179), .dinb(n267), .dout(n1180));
  jor  g0918(.dina(n1180), .dinb(n1176), .dout(n1181));
  jand g0919(.dina(n672), .dinb(shift1 ), .dout(n1182));
  jand g0920(.dina(n825), .dinb(n273), .dout(n1183));
  jor  g0921(.dina(n1183), .dinb(n1182), .dout(n1184));
  jand g0922(.dina(n1184), .dinb(n304), .dout(n1185));
  jor  g0923(.dina(n1185), .dinb(n1181), .dout(n1186));
  jor  g0924(.dina(n1186), .dinb(n1172), .dout(n1187));
  jand g0925(.dina(n1187), .dinb(n364), .dout(n1188));
  jand g0926(.dina(n716), .dinb(shift1 ), .dout(n1189));
  jand g0927(.dina(n778), .dinb(n273), .dout(n1190));
  jor  g0928(.dina(n1190), .dinb(n1189), .dout(n1191));
  jand g0929(.dina(n1191), .dinb(n304), .dout(n1192));
  jand g0930(.dina(n695), .dinb(shift1 ), .dout(n1193));
  jand g0931(.dina(n709), .dinb(n273), .dout(n1194));
  jor  g0932(.dina(n1194), .dinb(n1193), .dout(n1195));
  jand g0933(.dina(n1195), .dinb(n281), .dout(n1196));
  jand g0934(.dina(n685), .dinb(shift1 ), .dout(n1197));
  jand g0935(.dina(n699), .dinb(n273), .dout(n1198));
  jor  g0936(.dina(n1198), .dinb(n1197), .dout(n1199));
  jand g0937(.dina(n1199), .dinb(n292), .dout(n1200));
  jor  g0938(.dina(n1200), .dinb(n1196), .dout(n1201));
  jand g0939(.dina(n705), .dinb(shift1 ), .dout(n1202));
  jand g0940(.dina(n720), .dinb(n273), .dout(n1203));
  jor  g0941(.dina(n1203), .dinb(n1202), .dout(n1204));
  jand g0942(.dina(n1204), .dinb(n267), .dout(n1205));
  jor  g0943(.dina(n1205), .dinb(n1201), .dout(n1206));
  jor  g0944(.dina(n1206), .dinb(n1192), .dout(n1207));
  jand g0945(.dina(n1207), .dinb(n265), .dout(n1208));
  jand g0946(.dina(n729), .dinb(shift1 ), .dout(n1209));
  jand g0947(.dina(n689), .dinb(n273), .dout(n1210));
  jor  g0948(.dina(n1210), .dinb(n1209), .dout(n1211));
  jand g0949(.dina(n1211), .dinb(n304), .dout(n1212));
  jand g0950(.dina(n739), .dinb(shift1 ), .dout(n1213));
  jand g0951(.dina(n764), .dinb(n273), .dout(n1214));
  jor  g0952(.dina(n1214), .dinb(n1213), .dout(n1215));
  jand g0953(.dina(n1215), .dinb(n281), .dout(n1216));
  jand g0954(.dina(n760), .dinb(shift1 ), .dout(n1217));
  jand g0955(.dina(n733), .dinb(n273), .dout(n1218));
  jor  g0956(.dina(n1218), .dinb(n1217), .dout(n1219));
  jand g0957(.dina(n1219), .dinb(n267), .dout(n1220));
  jor  g0958(.dina(n1220), .dinb(n1216), .dout(n1221));
  jand g0959(.dina(n749), .dinb(shift1 ), .dout(n1222));
  jand g0960(.dina(n743), .dinb(n273), .dout(n1223));
  jor  g0961(.dina(n1223), .dinb(n1222), .dout(n1224));
  jand g0962(.dina(n1224), .dinb(n292), .dout(n1225));
  jor  g0963(.dina(n1225), .dinb(n1221), .dout(n1226));
  jor  g0964(.dina(n1226), .dinb(n1212), .dout(n1227));
  jand g0965(.dina(n1227), .dinb(n410), .dout(n1228));
  jor  g0966(.dina(n1228), .dinb(n1208), .dout(n1229));
  jand g0967(.dina(n774), .dinb(shift1 ), .dout(n1230));
  jand g0968(.dina(n784), .dinb(n273), .dout(n1231));
  jor  g0969(.dina(n1231), .dinb(n1230), .dout(n1232));
  jand g0970(.dina(n1232), .dinb(n292), .dout(n1233));
  jand g0971(.dina(n788), .dinb(shift1 ), .dout(n1234));
  jand g0972(.dina(n798), .dinb(n273), .dout(n1235));
  jor  g0973(.dina(n1235), .dinb(n1234), .dout(n1236));
  jand g0974(.dina(n1236), .dinb(n281), .dout(n1237));
  jor  g0975(.dina(n809), .dinb(shift1 ), .dout(n1238));
  jor  g0976(.dina(n794), .dinb(n273), .dout(n1239));
  jand g0977(.dina(n1239), .dinb(n1238), .dout(n1240));
  jand g0978(.dina(n1240), .dinb(n267), .dout(n1241));
  jor  g0979(.dina(n1241), .dinb(n1237), .dout(n1242));
  jand g0980(.dina(n805), .dinb(shift1 ), .dout(n1243));
  jand g0981(.dina(n665), .dinb(n273), .dout(n1244));
  jor  g0982(.dina(n1244), .dinb(n1243), .dout(n1245));
  jand g0983(.dina(n1245), .dinb(n304), .dout(n1246));
  jor  g0984(.dina(n1246), .dinb(n1242), .dout(n1247));
  jor  g0985(.dina(n1247), .dinb(n1233), .dout(n1248));
  jand g0986(.dina(n1248), .dinb(n319), .dout(n1249));
  jor  g0987(.dina(n1249), .dinb(n1229), .dout(n1250));
  jor  g0988(.dina(n1250), .dinb(n1188), .dout(n1251));
  jor  g0989(.dina(n1251), .dinb(n263), .dout(n1252));
  jand g0990(.dina(n896), .dinb(shift1 ), .dout(n1253));
  jand g0991(.dina(n978), .dinb(n273), .dout(n1254));
  jor  g0992(.dina(n1254), .dinb(n1253), .dout(n1255));
  jand g0993(.dina(n1255), .dinb(n304), .dout(n1256));
  jand g0994(.dina(n875), .dinb(shift1 ), .dout(n1257));
  jand g0995(.dina(n889), .dinb(n273), .dout(n1258));
  jor  g0996(.dina(n1258), .dinb(n1257), .dout(n1259));
  jand g0997(.dina(n1259), .dinb(n281), .dout(n1260));
  jand g0998(.dina(n885), .dinb(shift1 ), .dout(n1261));
  jand g0999(.dina(n900), .dinb(n273), .dout(n1262));
  jor  g1000(.dina(n1262), .dinb(n1261), .dout(n1263));
  jand g1001(.dina(n1263), .dinb(n267), .dout(n1264));
  jor  g1002(.dina(n1264), .dinb(n1260), .dout(n1265));
  jand g1003(.dina(n865), .dinb(shift1 ), .dout(n1266));
  jand g1004(.dina(n879), .dinb(n273), .dout(n1267));
  jor  g1005(.dina(n1267), .dinb(n1266), .dout(n1268));
  jand g1006(.dina(n1268), .dinb(n292), .dout(n1269));
  jor  g1007(.dina(n1269), .dinb(n1265), .dout(n1270));
  jor  g1008(.dina(n1270), .dinb(n1256), .dout(n1271));
  jand g1009(.dina(n1271), .dinb(n319), .dout(n1272));
  jand g1010(.dina(n852), .dinb(shift1 ), .dout(n1273));
  jand g1011(.dina(n913), .dinb(n273), .dout(n1274));
  jor  g1012(.dina(n1274), .dinb(n1273), .dout(n1275));
  jand g1013(.dina(n1275), .dinb(n304), .dout(n1276));
  jand g1014(.dina(n831), .dinb(shift1 ), .dout(n1277));
  jand g1015(.dina(n845), .dinb(n273), .dout(n1278));
  jor  g1016(.dina(n1278), .dinb(n1277), .dout(n1279));
  jand g1017(.dina(n1279), .dinb(n281), .dout(n1280));
  jand g1018(.dina(n841), .dinb(shift1 ), .dout(n1281));
  jand g1019(.dina(n856), .dinb(n273), .dout(n1282));
  jor  g1020(.dina(n1282), .dinb(n1281), .dout(n1283));
  jand g1021(.dina(n1283), .dinb(n267), .dout(n1284));
  jor  g1022(.dina(n1284), .dinb(n1280), .dout(n1285));
  jand g1023(.dina(n821), .dinb(shift1 ), .dout(n1286));
  jand g1024(.dina(n835), .dinb(n273), .dout(n1287));
  jor  g1025(.dina(n1287), .dinb(n1286), .dout(n1288));
  jand g1026(.dina(n1288), .dinb(n292), .dout(n1289));
  jor  g1027(.dina(n1289), .dinb(n1285), .dout(n1290));
  jor  g1028(.dina(n1290), .dinb(n1276), .dout(n1291));
  jand g1029(.dina(n1291), .dinb(n410), .dout(n1292));
  jand g1030(.dina(n974), .dinb(shift1 ), .dout(n1293));
  jand g1031(.dina(n968), .dinb(n273), .dout(n1294));
  jor  g1032(.dina(n1294), .dinb(n1293), .dout(n1295));
  jand g1033(.dina(n1295), .dinb(n292), .dout(n1296));
  jand g1034(.dina(n964), .dinb(shift1 ), .dout(n1297));
  jand g1035(.dina(n958), .dinb(n273), .dout(n1298));
  jor  g1036(.dina(n1298), .dinb(n1297), .dout(n1299));
  jand g1037(.dina(n1299), .dinb(n281), .dout(n1300));
  jand g1038(.dina(n954), .dinb(shift1 ), .dout(n1301));
  jand g1039(.dina(n989), .dinb(n273), .dout(n1302));
  jor  g1040(.dina(n1302), .dinb(n1301), .dout(n1303));
  jand g1041(.dina(n1303), .dinb(n267), .dout(n1304));
  jor  g1042(.dina(n1304), .dinb(n1300), .dout(n1305));
  jand g1043(.dina(n985), .dinb(shift1 ), .dout(n1306));
  jand g1044(.dina(n753), .dinb(n273), .dout(n1307));
  jor  g1045(.dina(n1307), .dinb(n1306), .dout(n1308));
  jand g1046(.dina(n1308), .dinb(n304), .dout(n1309));
  jor  g1047(.dina(n1309), .dinb(n1305), .dout(n1310));
  jor  g1048(.dina(n1310), .dinb(n1296), .dout(n1311));
  jand g1049(.dina(n1311), .dinb(n364), .dout(n1312));
  jor  g1050(.dina(n1312), .dinb(n1292), .dout(n1313));
  jand g1051(.dina(n940), .dinb(shift1 ), .dout(n1314));
  jand g1052(.dina(n869), .dinb(n273), .dout(n1315));
  jor  g1053(.dina(n1315), .dinb(n1314), .dout(n1316));
  jand g1054(.dina(n1316), .dinb(n304), .dout(n1317));
  jand g1055(.dina(n919), .dinb(shift1 ), .dout(n1318));
  jand g1056(.dina(n933), .dinb(n273), .dout(n1319));
  jor  g1057(.dina(n1319), .dinb(n1318), .dout(n1320));
  jand g1058(.dina(n1320), .dinb(n281), .dout(n1321));
  jand g1059(.dina(n929), .dinb(shift1 ), .dout(n1322));
  jand g1060(.dina(n944), .dinb(n273), .dout(n1323));
  jor  g1061(.dina(n1323), .dinb(n1322), .dout(n1324));
  jand g1062(.dina(n1324), .dinb(n267), .dout(n1325));
  jor  g1063(.dina(n1325), .dinb(n1321), .dout(n1326));
  jand g1064(.dina(n909), .dinb(shift1 ), .dout(n1327));
  jand g1065(.dina(n923), .dinb(n273), .dout(n1328));
  jor  g1066(.dina(n1328), .dinb(n1327), .dout(n1329));
  jand g1067(.dina(n1329), .dinb(n292), .dout(n1330));
  jor  g1068(.dina(n1330), .dinb(n1326), .dout(n1331));
  jor  g1069(.dina(n1331), .dinb(n1317), .dout(n1332));
  jand g1070(.dina(n1332), .dinb(n265), .dout(n1333));
  jor  g1071(.dina(n1333), .dinb(n1313), .dout(n1334));
  jor  g1072(.dina(n1334), .dinb(n1272), .dout(n1335));
  jor  g1073(.dina(n1335), .dinb(shift6 ), .dout(n1336));
  jand g1074(.dina(n1336), .dinb(n1252), .dout(result3 ));
  jand g1075(.dina(n383), .dinb(n292), .dout(n1338));
  jand g1076(.dina(n393), .dinb(n281), .dout(n1339));
  jand g1077(.dina(n373), .dinb(n267), .dout(n1340));
  jor  g1078(.dina(n1340), .dinb(n1339), .dout(n1341));
  jand g1079(.dina(n466), .dinb(n304), .dout(n1342));
  jor  g1080(.dina(n1342), .dinb(n1341), .dout(n1343));
  jor  g1081(.dina(n1343), .dinb(n1338), .dout(n1344));
  jand g1082(.dina(n1344), .dinb(n364), .dout(n1345));
  jand g1083(.dina(n450), .dinb(n267), .dout(n1346));
  jand g1084(.dina(n419), .dinb(n281), .dout(n1347));
  jand g1085(.dina(n429), .dinb(n292), .dout(n1348));
  jor  g1086(.dina(n1348), .dinb(n1347), .dout(n1349));
  jand g1087(.dina(n304), .dinb(n301), .dout(n1350));
  jor  g1088(.dina(n1350), .dinb(n1349), .dout(n1351));
  jor  g1089(.dina(n1351), .dinb(n1346), .dout(n1352));
  jand g1090(.dina(n1352), .dinb(n410), .dout(n1353));
  jand g1091(.dina(n328), .dinb(n304), .dout(n1354));
  jand g1092(.dina(n281), .dinb(n278), .dout(n1355));
  jand g1093(.dina(n292), .dinb(n290), .dout(n1356));
  jor  g1094(.dina(n1356), .dinb(n1355), .dout(n1357));
  jand g1095(.dina(n313), .dinb(n267), .dout(n1358));
  jor  g1096(.dina(n1358), .dinb(n1357), .dout(n1359));
  jor  g1097(.dina(n1359), .dinb(n1354), .dout(n1360));
  jand g1098(.dina(n1360), .dinb(n265), .dout(n1361));
  jor  g1099(.dina(n1361), .dinb(n1353), .dout(n1362));
  jand g1100(.dina(n359), .dinb(n267), .dout(n1363));
  jand g1101(.dina(n348), .dinb(n281), .dout(n1364));
  jand g1102(.dina(n338), .dinb(n292), .dout(n1365));
  jor  g1103(.dina(n1365), .dinb(n1364), .dout(n1366));
  jand g1104(.dina(n404), .dinb(n304), .dout(n1367));
  jor  g1105(.dina(n1367), .dinb(n1366), .dout(n1368));
  jor  g1106(.dina(n1368), .dinb(n1363), .dout(n1369));
  jand g1107(.dina(n1369), .dinb(n319), .dout(n1370));
  jor  g1108(.dina(n1370), .dinb(n1362), .dout(n1371));
  jor  g1109(.dina(n1371), .dinb(n1345), .dout(n1372));
  jor  g1110(.dina(n1372), .dinb(n263), .dout(n1373));
  jand g1111(.dina(n585), .dinb(n267), .dout(n1374));
  jand g1112(.dina(n554), .dinb(n281), .dout(n1375));
  jand g1113(.dina(n564), .dinb(n292), .dout(n1376));
  jor  g1114(.dina(n1376), .dinb(n1375), .dout(n1377));
  jand g1115(.dina(n510), .dinb(n304), .dout(n1378));
  jor  g1116(.dina(n1378), .dinb(n1377), .dout(n1379));
  jor  g1117(.dina(n1379), .dinb(n1374), .dout(n1380));
  jand g1118(.dina(n1380), .dinb(n265), .dout(n1381));
  jand g1119(.dina(n619), .dinb(n304), .dout(n1382));
  jand g1120(.dina(n530), .dinb(n281), .dout(n1383));
  jand g1121(.dina(n541), .dinb(n267), .dout(n1384));
  jor  g1122(.dina(n1384), .dinb(n1383), .dout(n1385));
  jand g1123(.dina(n520), .dinb(n292), .dout(n1386));
  jor  g1124(.dina(n1386), .dinb(n1385), .dout(n1387));
  jor  g1125(.dina(n1387), .dinb(n1382), .dout(n1388));
  jand g1126(.dina(n1388), .dinb(n319), .dout(n1389));
  jand g1127(.dina(n439), .dinb(n304), .dout(n1390));
  jand g1128(.dina(n599), .dinb(n281), .dout(n1391));
  jand g1129(.dina(n609), .dinb(n292), .dout(n1392));
  jor  g1130(.dina(n1392), .dinb(n1391), .dout(n1393));
  jand g1131(.dina(n630), .dinb(n267), .dout(n1394));
  jor  g1132(.dina(n1394), .dinb(n1393), .dout(n1395));
  jor  g1133(.dina(n1395), .dinb(n1390), .dout(n1396));
  jand g1134(.dina(n1396), .dinb(n364), .dout(n1397));
  jor  g1135(.dina(n1397), .dinb(n1389), .dout(n1398));
  jand g1136(.dina(n574), .dinb(n304), .dout(n1399));
  jand g1137(.dina(n486), .dinb(n281), .dout(n1400));
  jand g1138(.dina(n497), .dinb(n267), .dout(n1401));
  jor  g1139(.dina(n1401), .dinb(n1400), .dout(n1402));
  jand g1140(.dina(n476), .dinb(n292), .dout(n1403));
  jor  g1141(.dina(n1403), .dinb(n1402), .dout(n1404));
  jor  g1142(.dina(n1404), .dinb(n1399), .dout(n1405));
  jand g1143(.dina(n1405), .dinb(n410), .dout(n1406));
  jor  g1144(.dina(n1406), .dinb(n1398), .dout(n1407));
  jor  g1145(.dina(n1407), .dinb(n1381), .dout(n1408));
  jor  g1146(.dina(n1408), .dinb(shift6 ), .dout(n1409));
  jand g1147(.dina(n1409), .dinb(n1373), .dout(result4 ));
  jand g1148(.dina(n667), .dinb(n304), .dout(n1411));
  jand g1149(.dina(n800), .dinb(n281), .dout(n1412));
  jand g1150(.dina(n790), .dinb(n292), .dout(n1413));
  jor  g1151(.dina(n1413), .dinb(n1412), .dout(n1414));
  jand g1152(.dina(n811), .dinb(n267), .dout(n1415));
  jor  g1153(.dina(n1415), .dinb(n1414), .dout(n1416));
  jor  g1154(.dina(n1416), .dinb(n1411), .dout(n1417));
  jand g1155(.dina(n1417), .dinb(n319), .dout(n1418));
  jand g1156(.dina(n745), .dinb(n292), .dout(n1419));
  jand g1157(.dina(n766), .dinb(n281), .dout(n1420));
  jand g1158(.dina(n735), .dinb(n267), .dout(n1421));
  jor  g1159(.dina(n1421), .dinb(n1420), .dout(n1422));
  jand g1160(.dina(n691), .dinb(n304), .dout(n1423));
  jor  g1161(.dina(n1423), .dinb(n1422), .dout(n1424));
  jor  g1162(.dina(n1424), .dinb(n1419), .dout(n1425));
  jand g1163(.dina(n1425), .dinb(n410), .dout(n1426));
  jand g1164(.dina(n701), .dinb(n292), .dout(n1427));
  jand g1165(.dina(n711), .dinb(n281), .dout(n1428));
  jand g1166(.dina(n722), .dinb(n267), .dout(n1429));
  jor  g1167(.dina(n1429), .dinb(n1428), .dout(n1430));
  jand g1168(.dina(n780), .dinb(n304), .dout(n1431));
  jor  g1169(.dina(n1431), .dinb(n1430), .dout(n1432));
  jor  g1170(.dina(n1432), .dinb(n1427), .dout(n1433));
  jand g1171(.dina(n1433), .dinb(n265), .dout(n1434));
  jor  g1172(.dina(n1434), .dinb(n1426), .dout(n1435));
  jand g1173(.dina(n827), .dinb(n304), .dout(n1436));
  jand g1174(.dina(n647), .dinb(n281), .dout(n1437));
  jand g1175(.dina(n678), .dinb(n267), .dout(n1438));
  jor  g1176(.dina(n1438), .dinb(n1437), .dout(n1439));
  jand g1177(.dina(n657), .dinb(n292), .dout(n1440));
  jor  g1178(.dina(n1440), .dinb(n1439), .dout(n1441));
  jor  g1179(.dina(n1441), .dinb(n1436), .dout(n1442));
  jand g1180(.dina(n1442), .dinb(n364), .dout(n1443));
  jor  g1181(.dina(n1443), .dinb(n1435), .dout(n1444));
  jor  g1182(.dina(n1444), .dinb(n1418), .dout(n1445));
  jor  g1183(.dina(n1445), .dinb(n263), .dout(n1446));
  jand g1184(.dina(n837), .dinb(n292), .dout(n1447));
  jand g1185(.dina(n847), .dinb(n281), .dout(n1448));
  jand g1186(.dina(n858), .dinb(n267), .dout(n1449));
  jor  g1187(.dina(n1449), .dinb(n1448), .dout(n1450));
  jand g1188(.dina(n915), .dinb(n304), .dout(n1451));
  jor  g1189(.dina(n1451), .dinb(n1450), .dout(n1452));
  jor  g1190(.dina(n1452), .dinb(n1447), .dout(n1453));
  jand g1191(.dina(n1453), .dinb(n410), .dout(n1454));
  jand g1192(.dina(n980), .dinb(n304), .dout(n1455));
  jand g1193(.dina(n891), .dinb(n281), .dout(n1456));
  jand g1194(.dina(n881), .dinb(n292), .dout(n1457));
  jor  g1195(.dina(n1457), .dinb(n1456), .dout(n1458));
  jand g1196(.dina(n902), .dinb(n267), .dout(n1459));
  jor  g1197(.dina(n1459), .dinb(n1458), .dout(n1460));
  jor  g1198(.dina(n1460), .dinb(n1455), .dout(n1461));
  jand g1199(.dina(n1461), .dinb(n319), .dout(n1462));
  jand g1200(.dina(n871), .dinb(n304), .dout(n1463));
  jand g1201(.dina(n935), .dinb(n281), .dout(n1464));
  jand g1202(.dina(n925), .dinb(n292), .dout(n1465));
  jor  g1203(.dina(n1465), .dinb(n1464), .dout(n1466));
  jand g1204(.dina(n946), .dinb(n267), .dout(n1467));
  jor  g1205(.dina(n1467), .dinb(n1466), .dout(n1468));
  jor  g1206(.dina(n1468), .dinb(n1463), .dout(n1469));
  jand g1207(.dina(n1469), .dinb(n265), .dout(n1470));
  jor  g1208(.dina(n1470), .dinb(n1462), .dout(n1471));
  jand g1209(.dina(n755), .dinb(n304), .dout(n1472));
  jand g1210(.dina(n960), .dinb(n281), .dout(n1473));
  jand g1211(.dina(n970), .dinb(n292), .dout(n1474));
  jor  g1212(.dina(n1474), .dinb(n1473), .dout(n1475));
  jand g1213(.dina(n991), .dinb(n267), .dout(n1476));
  jor  g1214(.dina(n1476), .dinb(n1475), .dout(n1477));
  jor  g1215(.dina(n1477), .dinb(n1472), .dout(n1478));
  jand g1216(.dina(n1478), .dinb(n364), .dout(n1479));
  jor  g1217(.dina(n1479), .dinb(n1471), .dout(n1480));
  jor  g1218(.dina(n1480), .dinb(n1454), .dout(n1481));
  jor  g1219(.dina(n1481), .dinb(shift6 ), .dout(n1482));
  jand g1220(.dina(n1482), .dinb(n1446), .dout(result5 ));
  jand g1221(.dina(n1010), .dinb(n304), .dout(n1484));
  jand g1222(.dina(n1030), .dinb(n281), .dout(n1485));
  jand g1223(.dina(n1026), .dinb(n292), .dout(n1486));
  jor  g1224(.dina(n1486), .dinb(n1485), .dout(n1487));
  jand g1225(.dina(n1035), .dinb(n267), .dout(n1488));
  jor  g1226(.dina(n1488), .dinb(n1487), .dout(n1489));
  jor  g1227(.dina(n1489), .dinb(n1484), .dout(n1490));
  jand g1228(.dina(n1490), .dinb(n265), .dout(n1491));
  jand g1229(.dina(n1042), .dinb(n267), .dout(n1492));
  jand g1230(.dina(n1050), .dinb(n281), .dout(n1493));
  jand g1231(.dina(n1046), .dinb(n292), .dout(n1494));
  jor  g1232(.dina(n1494), .dinb(n1493), .dout(n1495));
  jand g1233(.dina(n1022), .dinb(n304), .dout(n1496));
  jor  g1234(.dina(n1496), .dinb(n1495), .dout(n1497));
  jor  g1235(.dina(n1497), .dinb(n1492), .dout(n1498));
  jand g1236(.dina(n1498), .dinb(n410), .dout(n1499));
  jand g1237(.dina(n1076), .dinb(n267), .dout(n1500));
  jand g1238(.dina(n1071), .dinb(n281), .dout(n1501));
  jand g1239(.dina(n1067), .dinb(n292), .dout(n1502));
  jor  g1240(.dina(n1502), .dinb(n1501), .dout(n1503));
  jand g1241(.dina(n1094), .dinb(n304), .dout(n1504));
  jor  g1242(.dina(n1504), .dinb(n1503), .dout(n1505));
  jor  g1243(.dina(n1505), .dinb(n1500), .dout(n1506));
  jand g1244(.dina(n1506), .dinb(n364), .dout(n1507));
  jor  g1245(.dina(n1507), .dinb(n1499), .dout(n1508));
  jand g1246(.dina(n1063), .dinb(n304), .dout(n1509));
  jand g1247(.dina(n1002), .dinb(n281), .dout(n1510));
  jand g1248(.dina(n1015), .dinb(n267), .dout(n1511));
  jor  g1249(.dina(n1511), .dinb(n1510), .dout(n1512));
  jand g1250(.dina(n1006), .dinb(n292), .dout(n1513));
  jor  g1251(.dina(n1513), .dinb(n1512), .dout(n1514));
  jor  g1252(.dina(n1514), .dinb(n1509), .dout(n1515));
  jand g1253(.dina(n1515), .dinb(n319), .dout(n1516));
  jor  g1254(.dina(n1516), .dinb(n1508), .dout(n1517));
  jor  g1255(.dina(n1517), .dinb(n1491), .dout(n1518));
  jor  g1256(.dina(n1518), .dinb(n263), .dout(n1519));
  jand g1257(.dina(n1147), .dinb(n304), .dout(n1520));
  jand g1258(.dina(n1086), .dinb(n281), .dout(n1521));
  jand g1259(.dina(n1099), .dinb(n267), .dout(n1522));
  jor  g1260(.dina(n1522), .dinb(n1521), .dout(n1523));
  jand g1261(.dina(n1090), .dinb(n292), .dout(n1524));
  jor  g1262(.dina(n1524), .dinb(n1523), .dout(n1525));
  jor  g1263(.dina(n1525), .dinb(n1520), .dout(n1526));
  jand g1264(.dina(n1526), .dinb(n410), .dout(n1527));
  jand g1265(.dina(n1106), .dinb(n267), .dout(n1528));
  jand g1266(.dina(n1119), .dinb(n281), .dout(n1529));
  jand g1267(.dina(n1110), .dinb(n292), .dout(n1530));
  jor  g1268(.dina(n1530), .dinb(n1529), .dout(n1531));
  jand g1269(.dina(n1139), .dinb(n304), .dout(n1532));
  jor  g1270(.dina(n1532), .dinb(n1531), .dout(n1533));
  jor  g1271(.dina(n1533), .dinb(n1528), .dout(n1534));
  jand g1272(.dina(n1534), .dinb(n319), .dout(n1535));
  jand g1273(.dina(n1055), .dinb(n304), .dout(n1536));
  jand g1274(.dina(n1134), .dinb(n281), .dout(n1537));
  jand g1275(.dina(n1126), .dinb(n267), .dout(n1538));
  jor  g1276(.dina(n1538), .dinb(n1537), .dout(n1539));
  jand g1277(.dina(n1130), .dinb(n292), .dout(n1540));
  jor  g1278(.dina(n1540), .dinb(n1539), .dout(n1541));
  jor  g1279(.dina(n1541), .dinb(n1536), .dout(n1542));
  jand g1280(.dina(n1542), .dinb(n364), .dout(n1543));
  jor  g1281(.dina(n1543), .dinb(n1535), .dout(n1544));
  jand g1282(.dina(n1151), .dinb(n292), .dout(n1545));
  jand g1283(.dina(n1155), .dinb(n281), .dout(n1546));
  jand g1284(.dina(n1160), .dinb(n267), .dout(n1547));
  jor  g1285(.dina(n1547), .dinb(n1546), .dout(n1548));
  jand g1286(.dina(n1114), .dinb(n304), .dout(n1549));
  jor  g1287(.dina(n1549), .dinb(n1548), .dout(n1550));
  jor  g1288(.dina(n1550), .dinb(n1545), .dout(n1551));
  jand g1289(.dina(n1551), .dinb(n265), .dout(n1552));
  jor  g1290(.dina(n1552), .dinb(n1544), .dout(n1553));
  jor  g1291(.dina(n1553), .dinb(n1527), .dout(n1554));
  jor  g1292(.dina(n1554), .dinb(shift6 ), .dout(n1555));
  jand g1293(.dina(n1555), .dinb(n1519), .dout(result6 ));
  jand g1294(.dina(n1191), .dinb(n267), .dout(n1557));
  jand g1295(.dina(n1204), .dinb(n281), .dout(n1558));
  jand g1296(.dina(n1195), .dinb(n292), .dout(n1559));
  jor  g1297(.dina(n1559), .dinb(n1558), .dout(n1560));
  jand g1298(.dina(n1232), .dinb(n304), .dout(n1561));
  jor  g1299(.dina(n1561), .dinb(n1560), .dout(n1562));
  jor  g1300(.dina(n1562), .dinb(n1557), .dout(n1563));
  jand g1301(.dina(n1563), .dinb(n265), .dout(n1564));
  jand g1302(.dina(n1199), .dinb(n304), .dout(n1565));
  jand g1303(.dina(n1219), .dinb(n281), .dout(n1566));
  jand g1304(.dina(n1211), .dinb(n267), .dout(n1567));
  jor  g1305(.dina(n1567), .dinb(n1566), .dout(n1568));
  jand g1306(.dina(n1215), .dinb(n292), .dout(n1569));
  jor  g1307(.dina(n1569), .dinb(n1568), .dout(n1570));
  jor  g1308(.dina(n1570), .dinb(n1565), .dout(n1571));
  jand g1309(.dina(n1571), .dinb(n410), .dout(n1572));
  jand g1310(.dina(n1184), .dinb(n267), .dout(n1573));
  jand g1311(.dina(n1179), .dinb(n281), .dout(n1574));
  jand g1312(.dina(n1175), .dinb(n292), .dout(n1575));
  jor  g1313(.dina(n1575), .dinb(n1574), .dout(n1576));
  jand g1314(.dina(n1288), .dinb(n304), .dout(n1577));
  jor  g1315(.dina(n1577), .dinb(n1576), .dout(n1578));
  jor  g1316(.dina(n1578), .dinb(n1573), .dout(n1579));
  jand g1317(.dina(n1579), .dinb(n364), .dout(n1580));
  jor  g1318(.dina(n1580), .dinb(n1572), .dout(n1581));
  jand g1319(.dina(n1240), .dinb(n281), .dout(n1582));
  jand g1320(.dina(n1171), .dinb(n304), .dout(n1583));
  jand g1321(.dina(n1236), .dinb(n292), .dout(n1584));
  jor  g1322(.dina(n1584), .dinb(n1583), .dout(n1585));
  jand g1323(.dina(n1245), .dinb(n267), .dout(n1586));
  jor  g1324(.dina(n1586), .dinb(n1585), .dout(n1587));
  jor  g1325(.dina(n1587), .dinb(n1582), .dout(n1588));
  jand g1326(.dina(n1588), .dinb(n319), .dout(n1589));
  jor  g1327(.dina(n1589), .dinb(n1581), .dout(n1590));
  jor  g1328(.dina(n1590), .dinb(n1564), .dout(n1591));
  jor  g1329(.dina(n1591), .dinb(n263), .dout(n1592));
  jand g1330(.dina(n1329), .dinb(n304), .dout(n1593));
  jand g1331(.dina(n1283), .dinb(n281), .dout(n1594));
  jand g1332(.dina(n1279), .dinb(n292), .dout(n1595));
  jor  g1333(.dina(n1595), .dinb(n1594), .dout(n1596));
  jand g1334(.dina(n1275), .dinb(n267), .dout(n1597));
  jor  g1335(.dina(n1597), .dinb(n1596), .dout(n1598));
  jor  g1336(.dina(n1598), .dinb(n1593), .dout(n1599));
  jand g1337(.dina(n1599), .dinb(n410), .dout(n1600));
  jand g1338(.dina(n1255), .dinb(n267), .dout(n1601));
  jand g1339(.dina(n1263), .dinb(n281), .dout(n1602));
  jand g1340(.dina(n1259), .dinb(n292), .dout(n1603));
  jor  g1341(.dina(n1603), .dinb(n1602), .dout(n1604));
  jand g1342(.dina(n1295), .dinb(n304), .dout(n1605));
  jor  g1343(.dina(n1605), .dinb(n1604), .dout(n1606));
  jor  g1344(.dina(n1606), .dinb(n1601), .dout(n1607));
  jand g1345(.dina(n1607), .dinb(n319), .dout(n1608));
  jand g1346(.dina(n1268), .dinb(n304), .dout(n1609));
  jand g1347(.dina(n1324), .dinb(n281), .dout(n1610));
  jand g1348(.dina(n1316), .dinb(n267), .dout(n1611));
  jor  g1349(.dina(n1611), .dinb(n1610), .dout(n1612));
  jand g1350(.dina(n1320), .dinb(n292), .dout(n1613));
  jor  g1351(.dina(n1613), .dinb(n1612), .dout(n1614));
  jor  g1352(.dina(n1614), .dinb(n1609), .dout(n1615));
  jand g1353(.dina(n1615), .dinb(n265), .dout(n1616));
  jor  g1354(.dina(n1616), .dinb(n1608), .dout(n1617));
  jand g1355(.dina(n1308), .dinb(n267), .dout(n1618));
  jand g1356(.dina(n1303), .dinb(n281), .dout(n1619));
  jand g1357(.dina(n1299), .dinb(n292), .dout(n1620));
  jor  g1358(.dina(n1620), .dinb(n1619), .dout(n1621));
  jand g1359(.dina(n1224), .dinb(n304), .dout(n1622));
  jor  g1360(.dina(n1622), .dinb(n1621), .dout(n1623));
  jor  g1361(.dina(n1623), .dinb(n1618), .dout(n1624));
  jand g1362(.dina(n1624), .dinb(n364), .dout(n1625));
  jor  g1363(.dina(n1625), .dinb(n1617), .dout(n1626));
  jor  g1364(.dina(n1626), .dinb(n1600), .dout(n1627));
  jor  g1365(.dina(n1627), .dinb(shift6 ), .dout(n1628));
  jand g1366(.dina(n1628), .dinb(n1592), .dout(result7 ));
  jand g1367(.dina(n292), .dinb(n278), .dout(n1630));
  jand g1368(.dina(n313), .dinb(n281), .dout(n1631));
  jand g1369(.dina(n328), .dinb(n267), .dout(n1632));
  jor  g1370(.dina(n1632), .dinb(n1631), .dout(n1633));
  jand g1371(.dina(n338), .dinb(n304), .dout(n1634));
  jor  g1372(.dina(n1634), .dinb(n1633), .dout(n1635));
  jor  g1373(.dina(n1635), .dinb(n1630), .dout(n1636));
  jand g1374(.dina(n1636), .dinb(n265), .dout(n1637));
  jand g1375(.dina(n304), .dinb(n290), .dout(n1638));
  jand g1376(.dina(n450), .dinb(n281), .dout(n1639));
  jand g1377(.dina(n301), .dinb(n267), .dout(n1640));
  jor  g1378(.dina(n1640), .dinb(n1639), .dout(n1641));
  jand g1379(.dina(n419), .dinb(n292), .dout(n1642));
  jor  g1380(.dina(n1642), .dinb(n1641), .dout(n1643));
  jor  g1381(.dina(n1643), .dinb(n1638), .dout(n1644));
  jand g1382(.dina(n1644), .dinb(n410), .dout(n1645));
  jand g1383(.dina(n476), .dinb(n304), .dout(n1646));
  jand g1384(.dina(n373), .dinb(n281), .dout(n1647));
  jand g1385(.dina(n393), .dinb(n292), .dout(n1648));
  jor  g1386(.dina(n1648), .dinb(n1647), .dout(n1649));
  jand g1387(.dina(n466), .dinb(n267), .dout(n1650));
  jor  g1388(.dina(n1650), .dinb(n1649), .dout(n1651));
  jor  g1389(.dina(n1651), .dinb(n1646), .dout(n1652));
  jand g1390(.dina(n1652), .dinb(n364), .dout(n1653));
  jor  g1391(.dina(n1653), .dinb(n1645), .dout(n1654));
  jand g1392(.dina(n348), .dinb(n292), .dout(n1655));
  jand g1393(.dina(n359), .dinb(n281), .dout(n1656));
  jand g1394(.dina(n404), .dinb(n267), .dout(n1657));
  jor  g1395(.dina(n1657), .dinb(n1656), .dout(n1658));
  jand g1396(.dina(n383), .dinb(n304), .dout(n1659));
  jor  g1397(.dina(n1659), .dinb(n1658), .dout(n1660));
  jor  g1398(.dina(n1660), .dinb(n1655), .dout(n1661));
  jand g1399(.dina(n1661), .dinb(n319), .dout(n1662));
  jor  g1400(.dina(n1662), .dinb(n1654), .dout(n1663));
  jor  g1401(.dina(n1663), .dinb(n1637), .dout(n1664));
  jor  g1402(.dina(n1664), .dinb(n263), .dout(n1665));
  jand g1403(.dina(n486), .dinb(n292), .dout(n1666));
  jand g1404(.dina(n497), .dinb(n281), .dout(n1667));
  jand g1405(.dina(n574), .dinb(n267), .dout(n1668));
  jor  g1406(.dina(n1668), .dinb(n1667), .dout(n1669));
  jand g1407(.dina(n564), .dinb(n304), .dout(n1670));
  jor  g1408(.dina(n1670), .dinb(n1669), .dout(n1671));
  jor  g1409(.dina(n1671), .dinb(n1666), .dout(n1672));
  jand g1410(.dina(n1672), .dinb(n410), .dout(n1673));
  jand g1411(.dina(n609), .dinb(n304), .dout(n1674));
  jand g1412(.dina(n541), .dinb(n281), .dout(n1675));
  jand g1413(.dina(n530), .dinb(n292), .dout(n1676));
  jor  g1414(.dina(n1676), .dinb(n1675), .dout(n1677));
  jand g1415(.dina(n619), .dinb(n267), .dout(n1678));
  jor  g1416(.dina(n1678), .dinb(n1677), .dout(n1679));
  jor  g1417(.dina(n1679), .dinb(n1674), .dout(n1680));
  jand g1418(.dina(n1680), .dinb(n319), .dout(n1681));
  jand g1419(.dina(n439), .dinb(n267), .dout(n1682));
  jand g1420(.dina(n630), .dinb(n281), .dout(n1683));
  jand g1421(.dina(n599), .dinb(n292), .dout(n1684));
  jor  g1422(.dina(n1684), .dinb(n1683), .dout(n1685));
  jand g1423(.dina(n429), .dinb(n304), .dout(n1686));
  jor  g1424(.dina(n1686), .dinb(n1685), .dout(n1687));
  jor  g1425(.dina(n1687), .dinb(n1682), .dout(n1688));
  jand g1426(.dina(n1688), .dinb(n364), .dout(n1689));
  jor  g1427(.dina(n1689), .dinb(n1681), .dout(n1690));
  jand g1428(.dina(n554), .dinb(n292), .dout(n1691));
  jand g1429(.dina(n585), .dinb(n281), .dout(n1692));
  jand g1430(.dina(n510), .dinb(n267), .dout(n1693));
  jor  g1431(.dina(n1693), .dinb(n1692), .dout(n1694));
  jand g1432(.dina(n520), .dinb(n304), .dout(n1695));
  jor  g1433(.dina(n1695), .dinb(n1694), .dout(n1696));
  jor  g1434(.dina(n1696), .dinb(n1691), .dout(n1697));
  jand g1435(.dina(n1697), .dinb(n265), .dout(n1698));
  jor  g1436(.dina(n1698), .dinb(n1690), .dout(n1699));
  jor  g1437(.dina(n1699), .dinb(n1673), .dout(n1700));
  jor  g1438(.dina(n1700), .dinb(shift6 ), .dout(n1701));
  jand g1439(.dina(n1701), .dinb(n1665), .dout(result8 ));
  jand g1440(.dina(n647), .dinb(n292), .dout(n1703));
  jand g1441(.dina(n678), .dinb(n281), .dout(n1704));
  jand g1442(.dina(n827), .dinb(n267), .dout(n1705));
  jor  g1443(.dina(n1705), .dinb(n1704), .dout(n1706));
  jand g1444(.dina(n837), .dinb(n304), .dout(n1707));
  jor  g1445(.dina(n1707), .dinb(n1706), .dout(n1708));
  jor  g1446(.dina(n1708), .dinb(n1703), .dout(n1709));
  jand g1447(.dina(n1709), .dinb(n364), .dout(n1710));
  jand g1448(.dina(n701), .dinb(n304), .dout(n1711));
  jand g1449(.dina(n735), .dinb(n281), .dout(n1712));
  jand g1450(.dina(n766), .dinb(n292), .dout(n1713));
  jor  g1451(.dina(n1713), .dinb(n1712), .dout(n1714));
  jand g1452(.dina(n691), .dinb(n267), .dout(n1715));
  jor  g1453(.dina(n1715), .dinb(n1714), .dout(n1716));
  jor  g1454(.dina(n1716), .dinb(n1711), .dout(n1717));
  jand g1455(.dina(n1717), .dinb(n410), .dout(n1718));
  jand g1456(.dina(n711), .dinb(n292), .dout(n1719));
  jand g1457(.dina(n722), .dinb(n281), .dout(n1720));
  jand g1458(.dina(n780), .dinb(n267), .dout(n1721));
  jor  g1459(.dina(n1721), .dinb(n1720), .dout(n1722));
  jand g1460(.dina(n790), .dinb(n304), .dout(n1723));
  jor  g1461(.dina(n1723), .dinb(n1722), .dout(n1724));
  jor  g1462(.dina(n1724), .dinb(n1719), .dout(n1725));
  jand g1463(.dina(n1725), .dinb(n265), .dout(n1726));
  jor  g1464(.dina(n1726), .dinb(n1718), .dout(n1727));
  jand g1465(.dina(n800), .dinb(n292), .dout(n1728));
  jand g1466(.dina(n811), .dinb(n281), .dout(n1729));
  jand g1467(.dina(n667), .dinb(n267), .dout(n1730));
  jor  g1468(.dina(n1730), .dinb(n1729), .dout(n1731));
  jand g1469(.dina(n657), .dinb(n304), .dout(n1732));
  jor  g1470(.dina(n1732), .dinb(n1731), .dout(n1733));
  jor  g1471(.dina(n1733), .dinb(n1728), .dout(n1734));
  jand g1472(.dina(n1734), .dinb(n319), .dout(n1735));
  jor  g1473(.dina(n1735), .dinb(n1727), .dout(n1736));
  jor  g1474(.dina(n1736), .dinb(n1710), .dout(n1737));
  jor  g1475(.dina(n1737), .dinb(n263), .dout(n1738));
  jand g1476(.dina(n881), .dinb(n304), .dout(n1739));
  jand g1477(.dina(n946), .dinb(n281), .dout(n1740));
  jand g1478(.dina(n935), .dinb(n292), .dout(n1741));
  jor  g1479(.dina(n1741), .dinb(n1740), .dout(n1742));
  jand g1480(.dina(n871), .dinb(n267), .dout(n1743));
  jor  g1481(.dina(n1743), .dinb(n1742), .dout(n1744));
  jor  g1482(.dina(n1744), .dinb(n1739), .dout(n1745));
  jand g1483(.dina(n1745), .dinb(n265), .dout(n1746));
  jand g1484(.dina(n891), .dinb(n292), .dout(n1747));
  jand g1485(.dina(n902), .dinb(n281), .dout(n1748));
  jand g1486(.dina(n980), .dinb(n267), .dout(n1749));
  jor  g1487(.dina(n1749), .dinb(n1748), .dout(n1750));
  jand g1488(.dina(n970), .dinb(n304), .dout(n1751));
  jor  g1489(.dina(n1751), .dinb(n1750), .dout(n1752));
  jor  g1490(.dina(n1752), .dinb(n1747), .dout(n1753));
  jand g1491(.dina(n1753), .dinb(n319), .dout(n1754));
  jand g1492(.dina(n960), .dinb(n292), .dout(n1755));
  jand g1493(.dina(n991), .dinb(n281), .dout(n1756));
  jand g1494(.dina(n755), .dinb(n267), .dout(n1757));
  jor  g1495(.dina(n1757), .dinb(n1756), .dout(n1758));
  jand g1496(.dina(n745), .dinb(n304), .dout(n1759));
  jor  g1497(.dina(n1759), .dinb(n1758), .dout(n1760));
  jor  g1498(.dina(n1760), .dinb(n1755), .dout(n1761));
  jand g1499(.dina(n1761), .dinb(n364), .dout(n1762));
  jor  g1500(.dina(n1762), .dinb(n1754), .dout(n1763));
  jand g1501(.dina(n847), .dinb(n292), .dout(n1764));
  jand g1502(.dina(n858), .dinb(n281), .dout(n1765));
  jand g1503(.dina(n915), .dinb(n267), .dout(n1766));
  jor  g1504(.dina(n1766), .dinb(n1765), .dout(n1767));
  jand g1505(.dina(n925), .dinb(n304), .dout(n1768));
  jor  g1506(.dina(n1768), .dinb(n1767), .dout(n1769));
  jor  g1507(.dina(n1769), .dinb(n1764), .dout(n1770));
  jand g1508(.dina(n1770), .dinb(n410), .dout(n1771));
  jor  g1509(.dina(n1771), .dinb(n1763), .dout(n1772));
  jor  g1510(.dina(n1772), .dinb(n1746), .dout(n1773));
  jor  g1511(.dina(n1773), .dinb(shift6 ), .dout(n1774));
  jand g1512(.dina(n1774), .dinb(n1738), .dout(result9 ));
  jand g1513(.dina(n1067), .dinb(n304), .dout(n1776));
  jand g1514(.dina(n1015), .dinb(n281), .dout(n1777));
  jand g1515(.dina(n1002), .dinb(n292), .dout(n1778));
  jor  g1516(.dina(n1778), .dinb(n1777), .dout(n1779));
  jand g1517(.dina(n1063), .dinb(n267), .dout(n1780));
  jor  g1518(.dina(n1780), .dinb(n1779), .dout(n1781));
  jor  g1519(.dina(n1781), .dinb(n1776), .dout(n1782));
  jand g1520(.dina(n1782), .dinb(n319), .dout(n1783));
  jand g1521(.dina(n1022), .dinb(n267), .dout(n1784));
  jand g1522(.dina(n1042), .dinb(n281), .dout(n1785));
  jand g1523(.dina(n1050), .dinb(n292), .dout(n1786));
  jor  g1524(.dina(n1786), .dinb(n1785), .dout(n1787));
  jand g1525(.dina(n1026), .dinb(n304), .dout(n1788));
  jor  g1526(.dina(n1788), .dinb(n1787), .dout(n1789));
  jor  g1527(.dina(n1789), .dinb(n1784), .dout(n1790));
  jand g1528(.dina(n1790), .dinb(n410), .dout(n1791));
  jand g1529(.dina(n1010), .dinb(n267), .dout(n1792));
  jand g1530(.dina(n1035), .dinb(n281), .dout(n1793));
  jand g1531(.dina(n1030), .dinb(n292), .dout(n1794));
  jor  g1532(.dina(n1794), .dinb(n1793), .dout(n1795));
  jand g1533(.dina(n1006), .dinb(n304), .dout(n1796));
  jor  g1534(.dina(n1796), .dinb(n1795), .dout(n1797));
  jor  g1535(.dina(n1797), .dinb(n1792), .dout(n1798));
  jand g1536(.dina(n1798), .dinb(n265), .dout(n1799));
  jor  g1537(.dina(n1799), .dinb(n1791), .dout(n1800));
  jand g1538(.dina(n1090), .dinb(n304), .dout(n1801));
  jand g1539(.dina(n1076), .dinb(n281), .dout(n1802));
  jand g1540(.dina(n1071), .dinb(n292), .dout(n1803));
  jor  g1541(.dina(n1803), .dinb(n1802), .dout(n1804));
  jand g1542(.dina(n1094), .dinb(n267), .dout(n1805));
  jor  g1543(.dina(n1805), .dinb(n1804), .dout(n1806));
  jor  g1544(.dina(n1806), .dinb(n1801), .dout(n1807));
  jand g1545(.dina(n1807), .dinb(n364), .dout(n1808));
  jor  g1546(.dina(n1808), .dinb(n1800), .dout(n1809));
  jor  g1547(.dina(n1809), .dinb(n1783), .dout(n1810));
  jor  g1548(.dina(n1810), .dinb(n263), .dout(n1811));
  jand g1549(.dina(n1046), .dinb(n304), .dout(n1812));
  jand g1550(.dina(n1126), .dinb(n281), .dout(n1813));
  jand g1551(.dina(n1055), .dinb(n267), .dout(n1814));
  jor  g1552(.dina(n1814), .dinb(n1813), .dout(n1815));
  jand g1553(.dina(n1134), .dinb(n292), .dout(n1816));
  jor  g1554(.dina(n1816), .dinb(n1815), .dout(n1817));
  jor  g1555(.dina(n1817), .dinb(n1812), .dout(n1818));
  jand g1556(.dina(n1818), .dinb(n364), .dout(n1819));
  jand g1557(.dina(n1119), .dinb(n292), .dout(n1820));
  jand g1558(.dina(n1106), .dinb(n281), .dout(n1821));
  jand g1559(.dina(n1139), .dinb(n267), .dout(n1822));
  jor  g1560(.dina(n1822), .dinb(n1821), .dout(n1823));
  jand g1561(.dina(n1130), .dinb(n304), .dout(n1824));
  jor  g1562(.dina(n1824), .dinb(n1823), .dout(n1825));
  jor  g1563(.dina(n1825), .dinb(n1820), .dout(n1826));
  jand g1564(.dina(n1826), .dinb(n319), .dout(n1827));
  jand g1565(.dina(n1110), .dinb(n304), .dout(n1828));
  jand g1566(.dina(n1160), .dinb(n281), .dout(n1829));
  jand g1567(.dina(n1114), .dinb(n267), .dout(n1830));
  jor  g1568(.dina(n1830), .dinb(n1829), .dout(n1831));
  jand g1569(.dina(n1155), .dinb(n292), .dout(n1832));
  jor  g1570(.dina(n1832), .dinb(n1831), .dout(n1833));
  jor  g1571(.dina(n1833), .dinb(n1828), .dout(n1834));
  jand g1572(.dina(n1834), .dinb(n265), .dout(n1835));
  jor  g1573(.dina(n1835), .dinb(n1827), .dout(n1836));
  jand g1574(.dina(n1151), .dinb(n304), .dout(n1837));
  jand g1575(.dina(n1099), .dinb(n281), .dout(n1838));
  jand g1576(.dina(n1086), .dinb(n292), .dout(n1839));
  jor  g1577(.dina(n1839), .dinb(n1838), .dout(n1840));
  jand g1578(.dina(n1147), .dinb(n267), .dout(n1841));
  jor  g1579(.dina(n1841), .dinb(n1840), .dout(n1842));
  jor  g1580(.dina(n1842), .dinb(n1837), .dout(n1843));
  jand g1581(.dina(n1843), .dinb(n410), .dout(n1844));
  jor  g1582(.dina(n1844), .dinb(n1836), .dout(n1845));
  jor  g1583(.dina(n1845), .dinb(n1819), .dout(n1846));
  jor  g1584(.dina(n1846), .dinb(shift6 ), .dout(n1847));
  jand g1585(.dina(n1847), .dinb(n1811), .dout(result10 ));
  jand g1586(.dina(n1245), .dinb(n281), .dout(n1849));
  jand g1587(.dina(n1171), .dinb(n267), .dout(n1850));
  jand g1588(.dina(n1240), .dinb(n292), .dout(n1851));
  jor  g1589(.dina(n1851), .dinb(n1850), .dout(n1852));
  jand g1590(.dina(n1175), .dinb(n304), .dout(n1853));
  jor  g1591(.dina(n1853), .dinb(n1852), .dout(n1854));
  jor  g1592(.dina(n1854), .dinb(n1849), .dout(n1855));
  jand g1593(.dina(n1855), .dinb(n319), .dout(n1856));
  jand g1594(.dina(n1195), .dinb(n304), .dout(n1857));
  jand g1595(.dina(n1211), .dinb(n281), .dout(n1858));
  jand g1596(.dina(n1219), .dinb(n292), .dout(n1859));
  jor  g1597(.dina(n1859), .dinb(n1858), .dout(n1860));
  jand g1598(.dina(n1199), .dinb(n267), .dout(n1861));
  jor  g1599(.dina(n1861), .dinb(n1860), .dout(n1862));
  jor  g1600(.dina(n1862), .dinb(n1857), .dout(n1863));
  jand g1601(.dina(n1863), .dinb(n410), .dout(n1864));
  jand g1602(.dina(n1236), .dinb(n304), .dout(n1865));
  jand g1603(.dina(n1191), .dinb(n281), .dout(n1866));
  jand g1604(.dina(n1204), .dinb(n292), .dout(n1867));
  jor  g1605(.dina(n1867), .dinb(n1866), .dout(n1868));
  jand g1606(.dina(n1232), .dinb(n267), .dout(n1869));
  jor  g1607(.dina(n1869), .dinb(n1868), .dout(n1870));
  jor  g1608(.dina(n1870), .dinb(n1865), .dout(n1871));
  jand g1609(.dina(n1871), .dinb(n265), .dout(n1872));
  jor  g1610(.dina(n1872), .dinb(n1864), .dout(n1873));
  jand g1611(.dina(n1279), .dinb(n304), .dout(n1874));
  jand g1612(.dina(n1184), .dinb(n281), .dout(n1875));
  jand g1613(.dina(n1288), .dinb(n267), .dout(n1876));
  jor  g1614(.dina(n1876), .dinb(n1875), .dout(n1877));
  jand g1615(.dina(n1179), .dinb(n292), .dout(n1878));
  jor  g1616(.dina(n1878), .dinb(n1877), .dout(n1879));
  jor  g1617(.dina(n1879), .dinb(n1874), .dout(n1880));
  jand g1618(.dina(n1880), .dinb(n364), .dout(n1881));
  jor  g1619(.dina(n1881), .dinb(n1873), .dout(n1882));
  jor  g1620(.dina(n1882), .dinb(n1856), .dout(n1883));
  jor  g1621(.dina(n1883), .dinb(n263), .dout(n1884));
  jand g1622(.dina(n1320), .dinb(n304), .dout(n1885));
  jand g1623(.dina(n1275), .dinb(n281), .dout(n1886));
  jand g1624(.dina(n1283), .dinb(n292), .dout(n1887));
  jor  g1625(.dina(n1887), .dinb(n1886), .dout(n1888));
  jand g1626(.dina(n1329), .dinb(n267), .dout(n1889));
  jor  g1627(.dina(n1889), .dinb(n1888), .dout(n1890));
  jor  g1628(.dina(n1890), .dinb(n1885), .dout(n1891));
  jand g1629(.dina(n1891), .dinb(n410), .dout(n1892));
  jand g1630(.dina(n1299), .dinb(n304), .dout(n1893));
  jand g1631(.dina(n1255), .dinb(n281), .dout(n1894));
  jand g1632(.dina(n1263), .dinb(n292), .dout(n1895));
  jor  g1633(.dina(n1895), .dinb(n1894), .dout(n1896));
  jand g1634(.dina(n1295), .dinb(n267), .dout(n1897));
  jor  g1635(.dina(n1897), .dinb(n1896), .dout(n1898));
  jor  g1636(.dina(n1898), .dinb(n1893), .dout(n1899));
  jand g1637(.dina(n1899), .dinb(n319), .dout(n1900));
  jand g1638(.dina(n1259), .dinb(n304), .dout(n1901));
  jand g1639(.dina(n1316), .dinb(n281), .dout(n1902));
  jand g1640(.dina(n1324), .dinb(n292), .dout(n1903));
  jor  g1641(.dina(n1903), .dinb(n1902), .dout(n1904));
  jand g1642(.dina(n1268), .dinb(n267), .dout(n1905));
  jor  g1643(.dina(n1905), .dinb(n1904), .dout(n1906));
  jor  g1644(.dina(n1906), .dinb(n1901), .dout(n1907));
  jand g1645(.dina(n1907), .dinb(n265), .dout(n1908));
  jor  g1646(.dina(n1908), .dinb(n1900), .dout(n1909));
  jand g1647(.dina(n1303), .dinb(n292), .dout(n1910));
  jand g1648(.dina(n1308), .dinb(n281), .dout(n1911));
  jand g1649(.dina(n1224), .dinb(n267), .dout(n1912));
  jor  g1650(.dina(n1912), .dinb(n1911), .dout(n1913));
  jand g1651(.dina(n1215), .dinb(n304), .dout(n1914));
  jor  g1652(.dina(n1914), .dinb(n1913), .dout(n1915));
  jor  g1653(.dina(n1915), .dinb(n1910), .dout(n1916));
  jand g1654(.dina(n1916), .dinb(n364), .dout(n1917));
  jor  g1655(.dina(n1917), .dinb(n1909), .dout(n1918));
  jor  g1656(.dina(n1918), .dinb(n1892), .dout(n1919));
  jor  g1657(.dina(n1919), .dinb(shift6 ), .dout(n1920));
  jand g1658(.dina(n1920), .dinb(n1884), .dout(result11 ));
  jand g1659(.dina(n348), .dinb(n304), .dout(n1922));
  jand g1660(.dina(n328), .dinb(n281), .dout(n1923));
  jand g1661(.dina(n313), .dinb(n292), .dout(n1924));
  jor  g1662(.dina(n1924), .dinb(n1923), .dout(n1925));
  jand g1663(.dina(n338), .dinb(n267), .dout(n1926));
  jor  g1664(.dina(n1926), .dinb(n1925), .dout(n1927));
  jor  g1665(.dina(n1927), .dinb(n1922), .dout(n1928));
  jand g1666(.dina(n1928), .dinb(n265), .dout(n1929));
  jand g1667(.dina(n304), .dinb(n278), .dout(n1930));
  jand g1668(.dina(n301), .dinb(n281), .dout(n1931));
  jand g1669(.dina(n450), .dinb(n292), .dout(n1932));
  jor  g1670(.dina(n1932), .dinb(n1931), .dout(n1933));
  jand g1671(.dina(n290), .dinb(n267), .dout(n1934));
  jor  g1672(.dina(n1934), .dinb(n1933), .dout(n1935));
  jor  g1673(.dina(n1935), .dinb(n1930), .dout(n1936));
  jand g1674(.dina(n1936), .dinb(n410), .dout(n1937));
  jand g1675(.dina(n486), .dinb(n304), .dout(n1938));
  jand g1676(.dina(n466), .dinb(n281), .dout(n1939));
  jand g1677(.dina(n476), .dinb(n267), .dout(n1940));
  jor  g1678(.dina(n1940), .dinb(n1939), .dout(n1941));
  jand g1679(.dina(n373), .dinb(n292), .dout(n1942));
  jor  g1680(.dina(n1942), .dinb(n1941), .dout(n1943));
  jor  g1681(.dina(n1943), .dinb(n1938), .dout(n1944));
  jand g1682(.dina(n1944), .dinb(n364), .dout(n1945));
  jor  g1683(.dina(n1945), .dinb(n1937), .dout(n1946));
  jand g1684(.dina(n393), .dinb(n304), .dout(n1947));
  jand g1685(.dina(n404), .dinb(n281), .dout(n1948));
  jand g1686(.dina(n383), .dinb(n267), .dout(n1949));
  jor  g1687(.dina(n1949), .dinb(n1948), .dout(n1950));
  jand g1688(.dina(n359), .dinb(n292), .dout(n1951));
  jor  g1689(.dina(n1951), .dinb(n1950), .dout(n1952));
  jor  g1690(.dina(n1952), .dinb(n1947), .dout(n1953));
  jand g1691(.dina(n1953), .dinb(n319), .dout(n1954));
  jor  g1692(.dina(n1954), .dinb(n1946), .dout(n1955));
  jor  g1693(.dina(n1955), .dinb(n1929), .dout(n1956));
  jor  g1694(.dina(n1956), .dinb(n263), .dout(n1957));
  jand g1695(.dina(n419), .dinb(n304), .dout(n1958));
  jand g1696(.dina(n439), .dinb(n281), .dout(n1959));
  jand g1697(.dina(n630), .dinb(n292), .dout(n1960));
  jor  g1698(.dina(n1960), .dinb(n1959), .dout(n1961));
  jand g1699(.dina(n429), .dinb(n267), .dout(n1962));
  jor  g1700(.dina(n1962), .dinb(n1961), .dout(n1963));
  jor  g1701(.dina(n1963), .dinb(n1958), .dout(n1964));
  jand g1702(.dina(n1964), .dinb(n364), .dout(n1965));
  jand g1703(.dina(n599), .dinb(n304), .dout(n1966));
  jand g1704(.dina(n619), .dinb(n281), .dout(n1967));
  jand g1705(.dina(n609), .dinb(n267), .dout(n1968));
  jor  g1706(.dina(n1968), .dinb(n1967), .dout(n1969));
  jand g1707(.dina(n541), .dinb(n292), .dout(n1970));
  jor  g1708(.dina(n1970), .dinb(n1969), .dout(n1971));
  jor  g1709(.dina(n1971), .dinb(n1966), .dout(n1972));
  jand g1710(.dina(n1972), .dinb(n319), .dout(n1973));
  jand g1711(.dina(n530), .dinb(n304), .dout(n1974));
  jand g1712(.dina(n510), .dinb(n281), .dout(n1975));
  jand g1713(.dina(n585), .dinb(n292), .dout(n1976));
  jor  g1714(.dina(n1976), .dinb(n1975), .dout(n1977));
  jand g1715(.dina(n520), .dinb(n267), .dout(n1978));
  jor  g1716(.dina(n1978), .dinb(n1977), .dout(n1979));
  jor  g1717(.dina(n1979), .dinb(n1974), .dout(n1980));
  jand g1718(.dina(n1980), .dinb(n265), .dout(n1981));
  jor  g1719(.dina(n1981), .dinb(n1973), .dout(n1982));
  jand g1720(.dina(n554), .dinb(n304), .dout(n1983));
  jand g1721(.dina(n574), .dinb(n281), .dout(n1984));
  jand g1722(.dina(n564), .dinb(n267), .dout(n1985));
  jor  g1723(.dina(n1985), .dinb(n1984), .dout(n1986));
  jand g1724(.dina(n497), .dinb(n292), .dout(n1987));
  jor  g1725(.dina(n1987), .dinb(n1986), .dout(n1988));
  jor  g1726(.dina(n1988), .dinb(n1983), .dout(n1989));
  jand g1727(.dina(n1989), .dinb(n410), .dout(n1990));
  jor  g1728(.dina(n1990), .dinb(n1982), .dout(n1991));
  jor  g1729(.dina(n1991), .dinb(n1965), .dout(n1992));
  jor  g1730(.dina(n1992), .dinb(shift6 ), .dout(n1993));
  jand g1731(.dina(n1993), .dinb(n1957), .dout(result12 ));
  jand g1732(.dina(n790), .dinb(n267), .dout(n1995));
  jand g1733(.dina(n780), .dinb(n281), .dout(n1996));
  jand g1734(.dina(n722), .dinb(n292), .dout(n1997));
  jor  g1735(.dina(n1997), .dinb(n1996), .dout(n1998));
  jand g1736(.dina(n800), .dinb(n304), .dout(n1999));
  jor  g1737(.dina(n1999), .dinb(n1998), .dout(n2000));
  jor  g1738(.dina(n2000), .dinb(n1995), .dout(n2001));
  jand g1739(.dina(n2001), .dinb(n265), .dout(n2002));
  jand g1740(.dina(n711), .dinb(n304), .dout(n2003));
  jand g1741(.dina(n691), .dinb(n281), .dout(n2004));
  jand g1742(.dina(n735), .dinb(n292), .dout(n2005));
  jor  g1743(.dina(n2005), .dinb(n2004), .dout(n2006));
  jand g1744(.dina(n701), .dinb(n267), .dout(n2007));
  jor  g1745(.dina(n2007), .dinb(n2006), .dout(n2008));
  jor  g1746(.dina(n2008), .dinb(n2003), .dout(n2009));
  jand g1747(.dina(n2009), .dinb(n410), .dout(n2010));
  jand g1748(.dina(n847), .dinb(n304), .dout(n2011));
  jand g1749(.dina(n827), .dinb(n281), .dout(n2012));
  jand g1750(.dina(n678), .dinb(n292), .dout(n2013));
  jor  g1751(.dina(n2013), .dinb(n2012), .dout(n2014));
  jand g1752(.dina(n837), .dinb(n267), .dout(n2015));
  jor  g1753(.dina(n2015), .dinb(n2014), .dout(n2016));
  jor  g1754(.dina(n2016), .dinb(n2011), .dout(n2017));
  jand g1755(.dina(n2017), .dinb(n364), .dout(n2018));
  jor  g1756(.dina(n2018), .dinb(n2010), .dout(n2019));
  jand g1757(.dina(n657), .dinb(n267), .dout(n2020));
  jand g1758(.dina(n667), .dinb(n281), .dout(n2021));
  jand g1759(.dina(n811), .dinb(n292), .dout(n2022));
  jor  g1760(.dina(n2022), .dinb(n2021), .dout(n2023));
  jand g1761(.dina(n647), .dinb(n304), .dout(n2024));
  jor  g1762(.dina(n2024), .dinb(n2023), .dout(n2025));
  jor  g1763(.dina(n2025), .dinb(n2020), .dout(n2026));
  jand g1764(.dina(n2026), .dinb(n319), .dout(n2027));
  jor  g1765(.dina(n2027), .dinb(n2019), .dout(n2028));
  jor  g1766(.dina(n2028), .dinb(n2002), .dout(n2029));
  jor  g1767(.dina(n2029), .dinb(n263), .dout(n2030));
  jand g1768(.dina(n935), .dinb(n304), .dout(n2031));
  jand g1769(.dina(n915), .dinb(n281), .dout(n2032));
  jand g1770(.dina(n925), .dinb(n267), .dout(n2033));
  jor  g1771(.dina(n2033), .dinb(n2032), .dout(n2034));
  jand g1772(.dina(n858), .dinb(n292), .dout(n2035));
  jor  g1773(.dina(n2035), .dinb(n2034), .dout(n2036));
  jor  g1774(.dina(n2036), .dinb(n2031), .dout(n2037));
  jand g1775(.dina(n2037), .dinb(n410), .dout(n2038));
  jand g1776(.dina(n960), .dinb(n304), .dout(n2039));
  jand g1777(.dina(n980), .dinb(n281), .dout(n2040));
  jand g1778(.dina(n902), .dinb(n292), .dout(n2041));
  jor  g1779(.dina(n2041), .dinb(n2040), .dout(n2042));
  jand g1780(.dina(n970), .dinb(n267), .dout(n2043));
  jor  g1781(.dina(n2043), .dinb(n2042), .dout(n2044));
  jor  g1782(.dina(n2044), .dinb(n2039), .dout(n2045));
  jand g1783(.dina(n2045), .dinb(n319), .dout(n2046));
  jand g1784(.dina(n766), .dinb(n304), .dout(n2047));
  jand g1785(.dina(n755), .dinb(n281), .dout(n2048));
  jand g1786(.dina(n991), .dinb(n292), .dout(n2049));
  jor  g1787(.dina(n2049), .dinb(n2048), .dout(n2050));
  jand g1788(.dina(n745), .dinb(n267), .dout(n2051));
  jor  g1789(.dina(n2051), .dinb(n2050), .dout(n2052));
  jor  g1790(.dina(n2052), .dinb(n2047), .dout(n2053));
  jand g1791(.dina(n2053), .dinb(n364), .dout(n2054));
  jor  g1792(.dina(n2054), .dinb(n2046), .dout(n2055));
  jand g1793(.dina(n881), .dinb(n267), .dout(n2056));
  jand g1794(.dina(n871), .dinb(n281), .dout(n2057));
  jand g1795(.dina(n946), .dinb(n292), .dout(n2058));
  jor  g1796(.dina(n2058), .dinb(n2057), .dout(n2059));
  jand g1797(.dina(n891), .dinb(n304), .dout(n2060));
  jor  g1798(.dina(n2060), .dinb(n2059), .dout(n2061));
  jor  g1799(.dina(n2061), .dinb(n2056), .dout(n2062));
  jand g1800(.dina(n2062), .dinb(n265), .dout(n2063));
  jor  g1801(.dina(n2063), .dinb(n2055), .dout(n2064));
  jor  g1802(.dina(n2064), .dinb(n2038), .dout(n2065));
  jor  g1803(.dina(n2065), .dinb(shift6 ), .dout(n2066));
  jand g1804(.dina(n2066), .dinb(n2030), .dout(result13 ));
  jand g1805(.dina(n1071), .dinb(n304), .dout(n2068));
  jand g1806(.dina(n1063), .dinb(n281), .dout(n2069));
  jand g1807(.dina(n1067), .dinb(n267), .dout(n2070));
  jor  g1808(.dina(n2070), .dinb(n2069), .dout(n2071));
  jand g1809(.dina(n1015), .dinb(n292), .dout(n2072));
  jor  g1810(.dina(n2072), .dinb(n2071), .dout(n2073));
  jor  g1811(.dina(n2073), .dinb(n2068), .dout(n2074));
  jand g1812(.dina(n2074), .dinb(n319), .dout(n2075));
  jand g1813(.dina(n1042), .dinb(n292), .dout(n2076));
  jand g1814(.dina(n1022), .dinb(n281), .dout(n2077));
  jand g1815(.dina(n1026), .dinb(n267), .dout(n2078));
  jor  g1816(.dina(n2078), .dinb(n2077), .dout(n2079));
  jand g1817(.dina(n1030), .dinb(n304), .dout(n2080));
  jor  g1818(.dina(n2080), .dinb(n2079), .dout(n2081));
  jor  g1819(.dina(n2081), .dinb(n2076), .dout(n2082));
  jand g1820(.dina(n2082), .dinb(n410), .dout(n2083));
  jand g1821(.dina(n1086), .dinb(n304), .dout(n2084));
  jand g1822(.dina(n1094), .dinb(n281), .dout(n2085));
  jand g1823(.dina(n1076), .dinb(n292), .dout(n2086));
  jor  g1824(.dina(n2086), .dinb(n2085), .dout(n2087));
  jand g1825(.dina(n1090), .dinb(n267), .dout(n2088));
  jor  g1826(.dina(n2088), .dinb(n2087), .dout(n2089));
  jor  g1827(.dina(n2089), .dinb(n2084), .dout(n2090));
  jand g1828(.dina(n2090), .dinb(n364), .dout(n2091));
  jor  g1829(.dina(n2091), .dinb(n2083), .dout(n2092));
  jand g1830(.dina(n1006), .dinb(n267), .dout(n2093));
  jand g1831(.dina(n1010), .dinb(n281), .dout(n2094));
  jand g1832(.dina(n1035), .dinb(n292), .dout(n2095));
  jor  g1833(.dina(n2095), .dinb(n2094), .dout(n2096));
  jand g1834(.dina(n1002), .dinb(n304), .dout(n2097));
  jor  g1835(.dina(n2097), .dinb(n2096), .dout(n2098));
  jor  g1836(.dina(n2098), .dinb(n2093), .dout(n2099));
  jand g1837(.dina(n2099), .dinb(n265), .dout(n2100));
  jor  g1838(.dina(n2100), .dinb(n2092), .dout(n2101));
  jor  g1839(.dina(n2101), .dinb(n2075), .dout(n2102));
  jor  g1840(.dina(n2102), .dinb(n263), .dout(n2103));
  jand g1841(.dina(n1160), .dinb(n292), .dout(n2104));
  jand g1842(.dina(n1114), .dinb(n281), .dout(n2105));
  jand g1843(.dina(n1110), .dinb(n267), .dout(n2106));
  jor  g1844(.dina(n2106), .dinb(n2105), .dout(n2107));
  jand g1845(.dina(n1119), .dinb(n304), .dout(n2108));
  jor  g1846(.dina(n2108), .dinb(n2107), .dout(n2109));
  jor  g1847(.dina(n2109), .dinb(n2104), .dout(n2110));
  jand g1848(.dina(n2110), .dinb(n265), .dout(n2111));
  jand g1849(.dina(n1134), .dinb(n304), .dout(n2112));
  jand g1850(.dina(n1139), .dinb(n281), .dout(n2113));
  jand g1851(.dina(n1130), .dinb(n267), .dout(n2114));
  jor  g1852(.dina(n2114), .dinb(n2113), .dout(n2115));
  jand g1853(.dina(n1106), .dinb(n292), .dout(n2116));
  jor  g1854(.dina(n2116), .dinb(n2115), .dout(n2117));
  jor  g1855(.dina(n2117), .dinb(n2112), .dout(n2118));
  jand g1856(.dina(n2118), .dinb(n319), .dout(n2119));
  jand g1857(.dina(n1050), .dinb(n304), .dout(n2120));
  jand g1858(.dina(n1055), .dinb(n281), .dout(n2121));
  jand g1859(.dina(n1126), .dinb(n292), .dout(n2122));
  jor  g1860(.dina(n2122), .dinb(n2121), .dout(n2123));
  jand g1861(.dina(n1046), .dinb(n267), .dout(n2124));
  jor  g1862(.dina(n2124), .dinb(n2123), .dout(n2125));
  jor  g1863(.dina(n2125), .dinb(n2120), .dout(n2126));
  jand g1864(.dina(n2126), .dinb(n364), .dout(n2127));
  jor  g1865(.dina(n2127), .dinb(n2119), .dout(n2128));
  jand g1866(.dina(n1099), .dinb(n292), .dout(n2129));
  jand g1867(.dina(n1147), .dinb(n281), .dout(n2130));
  jand g1868(.dina(n1151), .dinb(n267), .dout(n2131));
  jor  g1869(.dina(n2131), .dinb(n2130), .dout(n2132));
  jand g1870(.dina(n1155), .dinb(n304), .dout(n2133));
  jor  g1871(.dina(n2133), .dinb(n2132), .dout(n2134));
  jor  g1872(.dina(n2134), .dinb(n2129), .dout(n2135));
  jand g1873(.dina(n2135), .dinb(n410), .dout(n2136));
  jor  g1874(.dina(n2136), .dinb(n2128), .dout(n2137));
  jor  g1875(.dina(n2137), .dinb(n2111), .dout(n2138));
  jor  g1876(.dina(n2138), .dinb(shift6 ), .dout(n2139));
  jand g1877(.dina(n2139), .dinb(n2103), .dout(result14 ));
  jand g1878(.dina(n1175), .dinb(n267), .dout(n2141));
  jand g1879(.dina(n1171), .dinb(n281), .dout(n2142));
  jand g1880(.dina(n1245), .dinb(n292), .dout(n2143));
  jor  g1881(.dina(n2143), .dinb(n2142), .dout(n2144));
  jand g1882(.dina(n1179), .dinb(n304), .dout(n2145));
  jor  g1883(.dina(n2145), .dinb(n2144), .dout(n2146));
  jor  g1884(.dina(n2146), .dinb(n2141), .dout(n2147));
  jand g1885(.dina(n2147), .dinb(n319), .dout(n2148));
  jand g1886(.dina(n1204), .dinb(n304), .dout(n2149));
  jand g1887(.dina(n1199), .dinb(n281), .dout(n2150));
  jand g1888(.dina(n1211), .dinb(n292), .dout(n2151));
  jor  g1889(.dina(n2151), .dinb(n2150), .dout(n2152));
  jand g1890(.dina(n1195), .dinb(n267), .dout(n2153));
  jor  g1891(.dina(n2153), .dinb(n2152), .dout(n2154));
  jor  g1892(.dina(n2154), .dinb(n2149), .dout(n2155));
  jand g1893(.dina(n2155), .dinb(n410), .dout(n2156));
  jand g1894(.dina(n1236), .dinb(n267), .dout(n2157));
  jand g1895(.dina(n1232), .dinb(n281), .dout(n2158));
  jand g1896(.dina(n1191), .dinb(n292), .dout(n2159));
  jor  g1897(.dina(n2159), .dinb(n2158), .dout(n2160));
  jand g1898(.dina(n1240), .dinb(n304), .dout(n2161));
  jor  g1899(.dina(n2161), .dinb(n2160), .dout(n2162));
  jor  g1900(.dina(n2162), .dinb(n2157), .dout(n2163));
  jand g1901(.dina(n2163), .dinb(n265), .dout(n2164));
  jor  g1902(.dina(n2164), .dinb(n2156), .dout(n2165));
  jand g1903(.dina(n1184), .dinb(n292), .dout(n2166));
  jand g1904(.dina(n1288), .dinb(n281), .dout(n2167));
  jand g1905(.dina(n1279), .dinb(n267), .dout(n2168));
  jor  g1906(.dina(n2168), .dinb(n2167), .dout(n2169));
  jand g1907(.dina(n1283), .dinb(n304), .dout(n2170));
  jor  g1908(.dina(n2170), .dinb(n2169), .dout(n2171));
  jor  g1909(.dina(n2171), .dinb(n2166), .dout(n2172));
  jand g1910(.dina(n2172), .dinb(n364), .dout(n2173));
  jor  g1911(.dina(n2173), .dinb(n2165), .dout(n2174));
  jor  g1912(.dina(n2174), .dinb(n2148), .dout(n2175));
  jor  g1913(.dina(n2175), .dinb(n263), .dout(n2176));
  jand g1914(.dina(n1219), .dinb(n304), .dout(n2177));
  jand g1915(.dina(n1224), .dinb(n281), .dout(n2178));
  jand g1916(.dina(n1308), .dinb(n292), .dout(n2179));
  jor  g1917(.dina(n2179), .dinb(n2178), .dout(n2180));
  jand g1918(.dina(n1215), .dinb(n267), .dout(n2181));
  jor  g1919(.dina(n2181), .dinb(n2180), .dout(n2182));
  jor  g1920(.dina(n2182), .dinb(n2177), .dout(n2183));
  jand g1921(.dina(n2183), .dinb(n364), .dout(n2184));
  jand g1922(.dina(n1303), .dinb(n304), .dout(n2185));
  jand g1923(.dina(n1295), .dinb(n281), .dout(n2186));
  jand g1924(.dina(n1299), .dinb(n267), .dout(n2187));
  jor  g1925(.dina(n2187), .dinb(n2186), .dout(n2188));
  jand g1926(.dina(n1255), .dinb(n292), .dout(n2189));
  jor  g1927(.dina(n2189), .dinb(n2188), .dout(n2190));
  jor  g1928(.dina(n2190), .dinb(n2185), .dout(n2191));
  jand g1929(.dina(n2191), .dinb(n319), .dout(n2192));
  jand g1930(.dina(n1263), .dinb(n304), .dout(n2193));
  jand g1931(.dina(n1268), .dinb(n281), .dout(n2194));
  jand g1932(.dina(n1259), .dinb(n267), .dout(n2195));
  jor  g1933(.dina(n2195), .dinb(n2194), .dout(n2196));
  jand g1934(.dina(n1316), .dinb(n292), .dout(n2197));
  jor  g1935(.dina(n2197), .dinb(n2196), .dout(n2198));
  jor  g1936(.dina(n2198), .dinb(n2193), .dout(n2199));
  jand g1937(.dina(n2199), .dinb(n265), .dout(n2200));
  jor  g1938(.dina(n2200), .dinb(n2192), .dout(n2201));
  jand g1939(.dina(n1320), .dinb(n267), .dout(n2202));
  jand g1940(.dina(n1329), .dinb(n281), .dout(n2203));
  jand g1941(.dina(n1275), .dinb(n292), .dout(n2204));
  jor  g1942(.dina(n2204), .dinb(n2203), .dout(n2205));
  jand g1943(.dina(n1324), .dinb(n304), .dout(n2206));
  jor  g1944(.dina(n2206), .dinb(n2205), .dout(n2207));
  jor  g1945(.dina(n2207), .dinb(n2202), .dout(n2208));
  jand g1946(.dina(n2208), .dinb(n410), .dout(n2209));
  jor  g1947(.dina(n2209), .dinb(n2201), .dout(n2210));
  jor  g1948(.dina(n2210), .dinb(n2184), .dout(n2211));
  jor  g1949(.dina(n2211), .dinb(shift6 ), .dout(n2212));
  jand g1950(.dina(n2212), .dinb(n2176), .dout(result15 ));
  jand g1951(.dina(n407), .dinb(n319), .dout(n2214));
  jand g1952(.dina(n362), .dinb(n265), .dout(n2215));
  jand g1953(.dina(n410), .dinb(n316), .dout(n2216));
  jor  g1954(.dina(n2216), .dinb(n2215), .dout(n2217));
  jand g1955(.dina(n500), .dinb(n364), .dout(n2218));
  jor  g1956(.dina(n2218), .dinb(n2217), .dout(n2219));
  jor  g1957(.dina(n2219), .dinb(n2214), .dout(n2220));
  jor  g1958(.dina(n2220), .dinb(n263), .dout(n2221));
  jand g1959(.dina(n588), .dinb(n410), .dout(n2222));
  jand g1960(.dina(n633), .dinb(n319), .dout(n2223));
  jand g1961(.dina(n544), .dinb(n265), .dout(n2224));
  jor  g1962(.dina(n2224), .dinb(n2223), .dout(n2225));
  jand g1963(.dina(n453), .dinb(n364), .dout(n2226));
  jor  g1964(.dina(n2226), .dinb(n2225), .dout(n2227));
  jor  g1965(.dina(n2227), .dinb(n2222), .dout(n2228));
  jor  g1966(.dina(n2228), .dinb(shift6 ), .dout(n2229));
  jand g1967(.dina(n2229), .dinb(n2221), .dout(result16 ));
  jand g1968(.dina(n814), .dinb(n265), .dout(n2231));
  jand g1969(.dina(n725), .dinb(n410), .dout(n2232));
  jand g1970(.dina(n861), .dinb(n364), .dout(n2233));
  jor  g1971(.dina(n2233), .dinb(n2232), .dout(n2234));
  jand g1972(.dina(n681), .dinb(n319), .dout(n2235));
  jor  g1973(.dina(n2235), .dinb(n2234), .dout(n2236));
  jor  g1974(.dina(n2236), .dinb(n2231), .dout(n2237));
  jor  g1975(.dina(n2237), .dinb(n263), .dout(n2238));
  jand g1976(.dina(n769), .dinb(n364), .dout(n2239));
  jand g1977(.dina(n994), .dinb(n319), .dout(n2240));
  jand g1978(.dina(n905), .dinb(n265), .dout(n2241));
  jor  g1979(.dina(n2241), .dinb(n2240), .dout(n2242));
  jand g1980(.dina(n949), .dinb(n410), .dout(n2243));
  jor  g1981(.dina(n2243), .dinb(n2242), .dout(n2244));
  jor  g1982(.dina(n2244), .dinb(n2239), .dout(n2245));
  jor  g1983(.dina(n2245), .dinb(shift6 ), .dout(n2246));
  jand g1984(.dina(n2246), .dinb(n2238), .dout(result17 ));
  jand g1985(.dina(n1102), .dinb(n364), .dout(n2248));
  jand g1986(.dina(n1038), .dinb(n410), .dout(n2249));
  jand g1987(.dina(n1018), .dinb(n265), .dout(n2250));
  jor  g1988(.dina(n2250), .dinb(n2249), .dout(n2251));
  jand g1989(.dina(n1079), .dinb(n319), .dout(n2252));
  jor  g1990(.dina(n2252), .dinb(n2251), .dout(n2253));
  jor  g1991(.dina(n2253), .dinb(n2248), .dout(n2254));
  jor  g1992(.dina(n2254), .dinb(n263), .dout(n2255));
  jand g1993(.dina(n1058), .dinb(n364), .dout(n2256));
  jand g1994(.dina(n1142), .dinb(n319), .dout(n2257));
  jand g1995(.dina(n1122), .dinb(n265), .dout(n2258));
  jor  g1996(.dina(n2258), .dinb(n2257), .dout(n2259));
  jand g1997(.dina(n1163), .dinb(n410), .dout(n2260));
  jor  g1998(.dina(n2260), .dinb(n2259), .dout(n2261));
  jor  g1999(.dina(n2261), .dinb(n2256), .dout(n2262));
  jor  g2000(.dina(n2262), .dinb(shift6 ), .dout(n2263));
  jand g2001(.dina(n2263), .dinb(n2255), .dout(result18 ));
  jand g2002(.dina(n1187), .dinb(n319), .dout(n2265));
  jand g2003(.dina(n1248), .dinb(n265), .dout(n2266));
  jand g2004(.dina(n1207), .dinb(n410), .dout(n2267));
  jor  g2005(.dina(n2267), .dinb(n2266), .dout(n2268));
  jand g2006(.dina(n1291), .dinb(n364), .dout(n2269));
  jor  g2007(.dina(n2269), .dinb(n2268), .dout(n2270));
  jor  g2008(.dina(n2270), .dinb(n2265), .dout(n2271));
  jor  g2009(.dina(n2271), .dinb(n263), .dout(n2272));
  jand g2010(.dina(n1271), .dinb(n265), .dout(n2273));
  jand g2011(.dina(n1227), .dinb(n364), .dout(n2274));
  jand g2012(.dina(n1311), .dinb(n319), .dout(n2275));
  jor  g2013(.dina(n2275), .dinb(n2274), .dout(n2276));
  jand g2014(.dina(n1332), .dinb(n410), .dout(n2277));
  jor  g2015(.dina(n2277), .dinb(n2276), .dout(n2278));
  jor  g2016(.dina(n2278), .dinb(n2273), .dout(n2279));
  jor  g2017(.dina(n2279), .dinb(shift6 ), .dout(n2280));
  jand g2018(.dina(n2280), .dinb(n2272), .dout(result19 ));
  jand g2019(.dina(n1405), .dinb(n364), .dout(n2282));
  jand g2020(.dina(n1344), .dinb(n319), .dout(n2283));
  jand g2021(.dina(n1360), .dinb(n410), .dout(n2284));
  jor  g2022(.dina(n2284), .dinb(n2283), .dout(n2285));
  jand g2023(.dina(n1369), .dinb(n265), .dout(n2286));
  jor  g2024(.dina(n2286), .dinb(n2285), .dout(n2287));
  jor  g2025(.dina(n2287), .dinb(n2282), .dout(n2288));
  jor  g2026(.dina(n2288), .dinb(n263), .dout(n2289));
  jand g2027(.dina(n1380), .dinb(n410), .dout(n2290));
  jand g2028(.dina(n1396), .dinb(n319), .dout(n2291));
  jand g2029(.dina(n1388), .dinb(n265), .dout(n2292));
  jor  g2030(.dina(n2292), .dinb(n2291), .dout(n2293));
  jand g2031(.dina(n1352), .dinb(n364), .dout(n2294));
  jor  g2032(.dina(n2294), .dinb(n2293), .dout(n2295));
  jor  g2033(.dina(n2295), .dinb(n2290), .dout(n2296));
  jor  g2034(.dina(n2296), .dinb(shift6 ), .dout(n2297));
  jand g2035(.dina(n2297), .dinb(n2289), .dout(result20 ));
  jand g2036(.dina(n1417), .dinb(n265), .dout(n2299));
  jand g2037(.dina(n1442), .dinb(n319), .dout(n2300));
  jand g2038(.dina(n1433), .dinb(n410), .dout(n2301));
  jor  g2039(.dina(n2301), .dinb(n2300), .dout(n2302));
  jand g2040(.dina(n1453), .dinb(n364), .dout(n2303));
  jor  g2041(.dina(n2303), .dinb(n2302), .dout(n2304));
  jor  g2042(.dina(n2304), .dinb(n2299), .dout(n2305));
  jor  g2043(.dina(n2305), .dinb(n263), .dout(n2306));
  jand g2044(.dina(n1469), .dinb(n410), .dout(n2307));
  jand g2045(.dina(n1478), .dinb(n319), .dout(n2308));
  jand g2046(.dina(n1425), .dinb(n364), .dout(n2309));
  jor  g2047(.dina(n2309), .dinb(n2308), .dout(n2310));
  jand g2048(.dina(n1461), .dinb(n265), .dout(n2311));
  jor  g2049(.dina(n2311), .dinb(n2310), .dout(n2312));
  jor  g2050(.dina(n2312), .dinb(n2307), .dout(n2313));
  jor  g2051(.dina(n2313), .dinb(shift6 ), .dout(n2314));
  jand g2052(.dina(n2314), .dinb(n2306), .dout(result21 ));
  jand g2053(.dina(n1515), .dinb(n265), .dout(n2316));
  jand g2054(.dina(n1506), .dinb(n319), .dout(n2317));
  jand g2055(.dina(n1490), .dinb(n410), .dout(n2318));
  jor  g2056(.dina(n2318), .dinb(n2317), .dout(n2319));
  jand g2057(.dina(n1526), .dinb(n364), .dout(n2320));
  jor  g2058(.dina(n2320), .dinb(n2319), .dout(n2321));
  jor  g2059(.dina(n2321), .dinb(n2316), .dout(n2322));
  jor  g2060(.dina(n2322), .dinb(n263), .dout(n2323));
  jand g2061(.dina(n1551), .dinb(n410), .dout(n2324));
  jand g2062(.dina(n1542), .dinb(n319), .dout(n2325));
  jand g2063(.dina(n1534), .dinb(n265), .dout(n2326));
  jor  g2064(.dina(n2326), .dinb(n2325), .dout(n2327));
  jand g2065(.dina(n1498), .dinb(n364), .dout(n2328));
  jor  g2066(.dina(n2328), .dinb(n2327), .dout(n2329));
  jor  g2067(.dina(n2329), .dinb(n2324), .dout(n2330));
  jor  g2068(.dina(n2330), .dinb(shift6 ), .dout(n2331));
  jand g2069(.dina(n2331), .dinb(n2323), .dout(result22 ));
  jand g2070(.dina(n1588), .dinb(n265), .dout(n2333));
  jand g2071(.dina(n1599), .dinb(n364), .dout(n2334));
  jand g2072(.dina(n1579), .dinb(n319), .dout(n2335));
  jor  g2073(.dina(n2335), .dinb(n2334), .dout(n2336));
  jand g2074(.dina(n1563), .dinb(n410), .dout(n2337));
  jor  g2075(.dina(n2337), .dinb(n2336), .dout(n2338));
  jor  g2076(.dina(n2338), .dinb(n2333), .dout(n2339));
  jor  g2077(.dina(n2339), .dinb(n263), .dout(n2340));
  jand g2078(.dina(n1615), .dinb(n410), .dout(n2341));
  jand g2079(.dina(n1607), .dinb(n265), .dout(n2342));
  jand g2080(.dina(n1624), .dinb(n319), .dout(n2343));
  jor  g2081(.dina(n2343), .dinb(n2342), .dout(n2344));
  jand g2082(.dina(n1571), .dinb(n364), .dout(n2345));
  jor  g2083(.dina(n2345), .dinb(n2344), .dout(n2346));
  jor  g2084(.dina(n2346), .dinb(n2341), .dout(n2347));
  jor  g2085(.dina(n2347), .dinb(shift6 ), .dout(n2348));
  jand g2086(.dina(n2348), .dinb(n2340), .dout(result23 ));
  jand g2087(.dina(n1661), .dinb(n265), .dout(n2350));
  jand g2088(.dina(n1672), .dinb(n364), .dout(n2351));
  jand g2089(.dina(n1652), .dinb(n319), .dout(n2352));
  jor  g2090(.dina(n2352), .dinb(n2351), .dout(n2353));
  jand g2091(.dina(n1636), .dinb(n410), .dout(n2354));
  jor  g2092(.dina(n2354), .dinb(n2353), .dout(n2355));
  jor  g2093(.dina(n2355), .dinb(n2350), .dout(n2356));
  jor  g2094(.dina(n2356), .dinb(n263), .dout(n2357));
  jand g2095(.dina(n1688), .dinb(n319), .dout(n2358));
  jand g2096(.dina(n1680), .dinb(n265), .dout(n2359));
  jand g2097(.dina(n1644), .dinb(n364), .dout(n2360));
  jor  g2098(.dina(n2360), .dinb(n2359), .dout(n2361));
  jand g2099(.dina(n1697), .dinb(n410), .dout(n2362));
  jor  g2100(.dina(n2362), .dinb(n2361), .dout(n2363));
  jor  g2101(.dina(n2363), .dinb(n2358), .dout(n2364));
  jor  g2102(.dina(n2364), .dinb(shift6 ), .dout(n2365));
  jand g2103(.dina(n2365), .dinb(n2357), .dout(result24 ));
  jand g2104(.dina(n1725), .dinb(n410), .dout(n2367));
  jand g2105(.dina(n1770), .dinb(n364), .dout(n2368));
  jand g2106(.dina(n1709), .dinb(n319), .dout(n2369));
  jor  g2107(.dina(n2369), .dinb(n2368), .dout(n2370));
  jand g2108(.dina(n1734), .dinb(n265), .dout(n2371));
  jor  g2109(.dina(n2371), .dinb(n2370), .dout(n2372));
  jor  g2110(.dina(n2372), .dinb(n2367), .dout(n2373));
  jor  g2111(.dina(n2373), .dinb(n263), .dout(n2374));
  jand g2112(.dina(n1761), .dinb(n319), .dout(n2375));
  jand g2113(.dina(n1753), .dinb(n265), .dout(n2376));
  jand g2114(.dina(n1717), .dinb(n364), .dout(n2377));
  jor  g2115(.dina(n2377), .dinb(n2376), .dout(n2378));
  jand g2116(.dina(n1745), .dinb(n410), .dout(n2379));
  jor  g2117(.dina(n2379), .dinb(n2378), .dout(n2380));
  jor  g2118(.dina(n2380), .dinb(n2375), .dout(n2381));
  jor  g2119(.dina(n2381), .dinb(shift6 ), .dout(n2382));
  jand g2120(.dina(n2382), .dinb(n2374), .dout(result25 ));
  jand g2121(.dina(n1807), .dinb(n319), .dout(n2384));
  jand g2122(.dina(n1843), .dinb(n364), .dout(n2385));
  jand g2123(.dina(n1798), .dinb(n410), .dout(n2386));
  jor  g2124(.dina(n2386), .dinb(n2385), .dout(n2387));
  jand g2125(.dina(n1782), .dinb(n265), .dout(n2388));
  jor  g2126(.dina(n2388), .dinb(n2387), .dout(n2389));
  jor  g2127(.dina(n2389), .dinb(n2384), .dout(n2390));
  jor  g2128(.dina(n2390), .dinb(n263), .dout(n2391));
  jand g2129(.dina(n1834), .dinb(n410), .dout(n2392));
  jand g2130(.dina(n1818), .dinb(n319), .dout(n2393));
  jand g2131(.dina(n1826), .dinb(n265), .dout(n2394));
  jor  g2132(.dina(n2394), .dinb(n2393), .dout(n2395));
  jand g2133(.dina(n1790), .dinb(n364), .dout(n2396));
  jor  g2134(.dina(n2396), .dinb(n2395), .dout(n2397));
  jor  g2135(.dina(n2397), .dinb(n2392), .dout(n2398));
  jor  g2136(.dina(n2398), .dinb(shift6 ), .dout(n2399));
  jand g2137(.dina(n2399), .dinb(n2391), .dout(result26 ));
  jand g2138(.dina(n1855), .dinb(n265), .dout(n2401));
  jand g2139(.dina(n1891), .dinb(n364), .dout(n2402));
  jand g2140(.dina(n1871), .dinb(n410), .dout(n2403));
  jor  g2141(.dina(n2403), .dinb(n2402), .dout(n2404));
  jand g2142(.dina(n1880), .dinb(n319), .dout(n2405));
  jor  g2143(.dina(n2405), .dinb(n2404), .dout(n2406));
  jor  g2144(.dina(n2406), .dinb(n2401), .dout(n2407));
  jor  g2145(.dina(n2407), .dinb(n263), .dout(n2408));
  jand g2146(.dina(n1907), .dinb(n410), .dout(n2409));
  jand g2147(.dina(n1916), .dinb(n319), .dout(n2410));
  jand g2148(.dina(n1899), .dinb(n265), .dout(n2411));
  jor  g2149(.dina(n2411), .dinb(n2410), .dout(n2412));
  jand g2150(.dina(n1863), .dinb(n364), .dout(n2413));
  jor  g2151(.dina(n2413), .dinb(n2412), .dout(n2414));
  jor  g2152(.dina(n2414), .dinb(n2409), .dout(n2415));
  jor  g2153(.dina(n2415), .dinb(shift6 ), .dout(n2416));
  jand g2154(.dina(n2416), .dinb(n2408), .dout(result27 ));
  jand g2155(.dina(n1953), .dinb(n265), .dout(n2418));
  jand g2156(.dina(n1989), .dinb(n364), .dout(n2419));
  jand g2157(.dina(n1944), .dinb(n319), .dout(n2420));
  jor  g2158(.dina(n2420), .dinb(n2419), .dout(n2421));
  jand g2159(.dina(n1928), .dinb(n410), .dout(n2422));
  jor  g2160(.dina(n2422), .dinb(n2421), .dout(n2423));
  jor  g2161(.dina(n2423), .dinb(n2418), .dout(n2424));
  jor  g2162(.dina(n2424), .dinb(n263), .dout(n2425));
  jand g2163(.dina(n1972), .dinb(n265), .dout(n2426));
  jand g2164(.dina(n1964), .dinb(n319), .dout(n2427));
  jand g2165(.dina(n1936), .dinb(n364), .dout(n2428));
  jor  g2166(.dina(n2428), .dinb(n2427), .dout(n2429));
  jand g2167(.dina(n1980), .dinb(n410), .dout(n2430));
  jor  g2168(.dina(n2430), .dinb(n2429), .dout(n2431));
  jor  g2169(.dina(n2431), .dinb(n2426), .dout(n2432));
  jor  g2170(.dina(n2432), .dinb(shift6 ), .dout(n2433));
  jand g2171(.dina(n2433), .dinb(n2425), .dout(result28 ));
  jand g2172(.dina(n2017), .dinb(n319), .dout(n2435));
  jand g2173(.dina(n2037), .dinb(n364), .dout(n2436));
  jand g2174(.dina(n2001), .dinb(n410), .dout(n2437));
  jor  g2175(.dina(n2437), .dinb(n2436), .dout(n2438));
  jand g2176(.dina(n2026), .dinb(n265), .dout(n2439));
  jor  g2177(.dina(n2439), .dinb(n2438), .dout(n2440));
  jor  g2178(.dina(n2440), .dinb(n2435), .dout(n2441));
  jor  g2179(.dina(n2441), .dinb(n263), .dout(n2442));
  jand g2180(.dina(n2062), .dinb(n410), .dout(n2443));
  jand g2181(.dina(n2053), .dinb(n319), .dout(n2444));
  jand g2182(.dina(n2045), .dinb(n265), .dout(n2445));
  jor  g2183(.dina(n2445), .dinb(n2444), .dout(n2446));
  jand g2184(.dina(n2009), .dinb(n364), .dout(n2447));
  jor  g2185(.dina(n2447), .dinb(n2446), .dout(n2448));
  jor  g2186(.dina(n2448), .dinb(n2443), .dout(n2449));
  jor  g2187(.dina(n2449), .dinb(shift6 ), .dout(n2450));
  jand g2188(.dina(n2450), .dinb(n2442), .dout(result29 ));
  jand g2189(.dina(n2090), .dinb(n319), .dout(n2452));
  jand g2190(.dina(n2135), .dinb(n364), .dout(n2453));
  jand g2191(.dina(n2099), .dinb(n410), .dout(n2454));
  jor  g2192(.dina(n2454), .dinb(n2453), .dout(n2455));
  jand g2193(.dina(n2074), .dinb(n265), .dout(n2456));
  jor  g2194(.dina(n2456), .dinb(n2455), .dout(n2457));
  jor  g2195(.dina(n2457), .dinb(n2452), .dout(n2458));
  jor  g2196(.dina(n2458), .dinb(n263), .dout(n2459));
  jand g2197(.dina(n2082), .dinb(n364), .dout(n2460));
  jand g2198(.dina(n2126), .dinb(n319), .dout(n2461));
  jand g2199(.dina(n2118), .dinb(n265), .dout(n2462));
  jor  g2200(.dina(n2462), .dinb(n2461), .dout(n2463));
  jand g2201(.dina(n2110), .dinb(n410), .dout(n2464));
  jor  g2202(.dina(n2464), .dinb(n2463), .dout(n2465));
  jor  g2203(.dina(n2465), .dinb(n2460), .dout(n2466));
  jor  g2204(.dina(n2466), .dinb(shift6 ), .dout(n2467));
  jand g2205(.dina(n2467), .dinb(n2459), .dout(result30 ));
  jand g2206(.dina(n2147), .dinb(n265), .dout(n2469));
  jand g2207(.dina(n2208), .dinb(n364), .dout(n2470));
  jand g2208(.dina(n2163), .dinb(n410), .dout(n2471));
  jor  g2209(.dina(n2471), .dinb(n2470), .dout(n2472));
  jand g2210(.dina(n2172), .dinb(n319), .dout(n2473));
  jor  g2211(.dina(n2473), .dinb(n2472), .dout(n2474));
  jor  g2212(.dina(n2474), .dinb(n2469), .dout(n2475));
  jor  g2213(.dina(n2475), .dinb(n263), .dout(n2476));
  jand g2214(.dina(n2191), .dinb(n265), .dout(n2477));
  jand g2215(.dina(n2183), .dinb(n319), .dout(n2478));
  jand g2216(.dina(n2155), .dinb(n364), .dout(n2479));
  jor  g2217(.dina(n2479), .dinb(n2478), .dout(n2480));
  jand g2218(.dina(n2199), .dinb(n410), .dout(n2481));
  jor  g2219(.dina(n2481), .dinb(n2480), .dout(n2482));
  jor  g2220(.dina(n2482), .dinb(n2477), .dout(n2483));
  jor  g2221(.dina(n2483), .dinb(shift6 ), .dout(n2484));
  jand g2222(.dina(n2484), .dinb(n2476), .dout(result31 ));
  jand g2223(.dina(n500), .dinb(n319), .dout(n2486));
  jand g2224(.dina(n410), .dinb(n362), .dout(n2487));
  jand g2225(.dina(n588), .dinb(n364), .dout(n2488));
  jor  g2226(.dina(n2488), .dinb(n2487), .dout(n2489));
  jand g2227(.dina(n407), .dinb(n265), .dout(n2490));
  jor  g2228(.dina(n2490), .dinb(n2489), .dout(n2491));
  jor  g2229(.dina(n2491), .dinb(n2486), .dout(n2492));
  jor  g2230(.dina(n2492), .dinb(n263), .dout(n2493));
  jand g2231(.dina(n633), .dinb(n265), .dout(n2494));
  jand g2232(.dina(n453), .dinb(n319), .dout(n2495));
  jand g2233(.dina(n364), .dinb(n316), .dout(n2496));
  jor  g2234(.dina(n2496), .dinb(n2495), .dout(n2497));
  jand g2235(.dina(n544), .dinb(n410), .dout(n2498));
  jor  g2236(.dina(n2498), .dinb(n2497), .dout(n2499));
  jor  g2237(.dina(n2499), .dinb(n2494), .dout(n2500));
  jor  g2238(.dina(n2500), .dinb(shift6 ), .dout(n2501));
  jand g2239(.dina(n2501), .dinb(n2493), .dout(result32 ));
  jand g2240(.dina(n861), .dinb(n319), .dout(n2503));
  jand g2241(.dina(n949), .dinb(n364), .dout(n2504));
  jand g2242(.dina(n814), .dinb(n410), .dout(n2505));
  jor  g2243(.dina(n2505), .dinb(n2504), .dout(n2506));
  jand g2244(.dina(n681), .dinb(n265), .dout(n2507));
  jor  g2245(.dina(n2507), .dinb(n2506), .dout(n2508));
  jor  g2246(.dina(n2508), .dinb(n2503), .dout(n2509));
  jor  g2247(.dina(n2509), .dinb(n263), .dout(n2510));
  jand g2248(.dina(n994), .dinb(n265), .dout(n2511));
  jand g2249(.dina(n769), .dinb(n319), .dout(n2512));
  jand g2250(.dina(n725), .dinb(n364), .dout(n2513));
  jor  g2251(.dina(n2513), .dinb(n2512), .dout(n2514));
  jand g2252(.dina(n905), .dinb(n410), .dout(n2515));
  jor  g2253(.dina(n2515), .dinb(n2514), .dout(n2516));
  jor  g2254(.dina(n2516), .dinb(n2511), .dout(n2517));
  jor  g2255(.dina(n2517), .dinb(shift6 ), .dout(n2518));
  jand g2256(.dina(n2518), .dinb(n2510), .dout(result33 ));
  jand g2257(.dina(n1079), .dinb(n265), .dout(n2520));
  jand g2258(.dina(n1163), .dinb(n364), .dout(n2521));
  jand g2259(.dina(n1102), .dinb(n319), .dout(n2522));
  jor  g2260(.dina(n2522), .dinb(n2521), .dout(n2523));
  jand g2261(.dina(n1018), .dinb(n410), .dout(n2524));
  jor  g2262(.dina(n2524), .dinb(n2523), .dout(n2525));
  jor  g2263(.dina(n2525), .dinb(n2520), .dout(n2526));
  jor  g2264(.dina(n2526), .dinb(n263), .dout(n2527));
  jand g2265(.dina(n1122), .dinb(n410), .dout(n2528));
  jand g2266(.dina(n1058), .dinb(n319), .dout(n2529));
  jand g2267(.dina(n1142), .dinb(n265), .dout(n2530));
  jor  g2268(.dina(n2530), .dinb(n2529), .dout(n2531));
  jand g2269(.dina(n1038), .dinb(n364), .dout(n2532));
  jor  g2270(.dina(n2532), .dinb(n2531), .dout(n2533));
  jor  g2271(.dina(n2533), .dinb(n2528), .dout(n2534));
  jor  g2272(.dina(n2534), .dinb(shift6 ), .dout(n2535));
  jand g2273(.dina(n2535), .dinb(n2527), .dout(result34 ));
  jand g2274(.dina(n1187), .dinb(n265), .dout(n2537));
  jand g2275(.dina(n1291), .dinb(n319), .dout(n2538));
  jand g2276(.dina(n1332), .dinb(n364), .dout(n2539));
  jor  g2277(.dina(n2539), .dinb(n2538), .dout(n2540));
  jand g2278(.dina(n1248), .dinb(n410), .dout(n2541));
  jor  g2279(.dina(n2541), .dinb(n2540), .dout(n2542));
  jor  g2280(.dina(n2542), .dinb(n2537), .dout(n2543));
  jor  g2281(.dina(n2543), .dinb(n263), .dout(n2544));
  jand g2282(.dina(n1271), .dinb(n410), .dout(n2545));
  jand g2283(.dina(n1227), .dinb(n319), .dout(n2546));
  jand g2284(.dina(n1311), .dinb(n265), .dout(n2547));
  jor  g2285(.dina(n2547), .dinb(n2546), .dout(n2548));
  jand g2286(.dina(n1207), .dinb(n364), .dout(n2549));
  jor  g2287(.dina(n2549), .dinb(n2548), .dout(n2550));
  jor  g2288(.dina(n2550), .dinb(n2545), .dout(n2551));
  jor  g2289(.dina(n2551), .dinb(shift6 ), .dout(n2552));
  jand g2290(.dina(n2552), .dinb(n2544), .dout(result35 ));
  jand g2291(.dina(n1405), .dinb(n319), .dout(n2554));
  jand g2292(.dina(n1369), .dinb(n410), .dout(n2555));
  jand g2293(.dina(n1380), .dinb(n364), .dout(n2556));
  jor  g2294(.dina(n2556), .dinb(n2555), .dout(n2557));
  jand g2295(.dina(n1344), .dinb(n265), .dout(n2558));
  jor  g2296(.dina(n2558), .dinb(n2557), .dout(n2559));
  jor  g2297(.dina(n2559), .dinb(n2554), .dout(n2560));
  jor  g2298(.dina(n2560), .dinb(n263), .dout(n2561));
  jand g2299(.dina(n1396), .dinb(n265), .dout(n2562));
  jand g2300(.dina(n1352), .dinb(n319), .dout(n2563));
  jand g2301(.dina(n1360), .dinb(n364), .dout(n2564));
  jor  g2302(.dina(n2564), .dinb(n2563), .dout(n2565));
  jand g2303(.dina(n1388), .dinb(n410), .dout(n2566));
  jor  g2304(.dina(n2566), .dinb(n2565), .dout(n2567));
  jor  g2305(.dina(n2567), .dinb(n2562), .dout(n2568));
  jor  g2306(.dina(n2568), .dinb(shift6 ), .dout(n2569));
  jand g2307(.dina(n2569), .dinb(n2561), .dout(result36 ));
  jand g2308(.dina(n1453), .dinb(n319), .dout(n2571));
  jand g2309(.dina(n1417), .dinb(n410), .dout(n2572));
  jand g2310(.dina(n1469), .dinb(n364), .dout(n2573));
  jor  g2311(.dina(n2573), .dinb(n2572), .dout(n2574));
  jand g2312(.dina(n1442), .dinb(n265), .dout(n2575));
  jor  g2313(.dina(n2575), .dinb(n2574), .dout(n2576));
  jor  g2314(.dina(n2576), .dinb(n2571), .dout(n2577));
  jor  g2315(.dina(n2577), .dinb(n263), .dout(n2578));
  jand g2316(.dina(n1461), .dinb(n410), .dout(n2579));
  jand g2317(.dina(n1425), .dinb(n319), .dout(n2580));
  jand g2318(.dina(n1433), .dinb(n364), .dout(n2581));
  jor  g2319(.dina(n2581), .dinb(n2580), .dout(n2582));
  jand g2320(.dina(n1478), .dinb(n265), .dout(n2583));
  jor  g2321(.dina(n2583), .dinb(n2582), .dout(n2584));
  jor  g2322(.dina(n2584), .dinb(n2579), .dout(n2585));
  jor  g2323(.dina(n2585), .dinb(shift6 ), .dout(n2586));
  jand g2324(.dina(n2586), .dinb(n2578), .dout(result37 ));
  jand g2325(.dina(n1506), .dinb(n265), .dout(n2588));
  jand g2326(.dina(n1515), .dinb(n410), .dout(n2589));
  jand g2327(.dina(n1551), .dinb(n364), .dout(n2590));
  jor  g2328(.dina(n2590), .dinb(n2589), .dout(n2591));
  jand g2329(.dina(n1526), .dinb(n319), .dout(n2592));
  jor  g2330(.dina(n2592), .dinb(n2591), .dout(n2593));
  jor  g2331(.dina(n2593), .dinb(n2588), .dout(n2594));
  jor  g2332(.dina(n2594), .dinb(n263), .dout(n2595));
  jand g2333(.dina(n1534), .dinb(n410), .dout(n2596));
  jand g2334(.dina(n1498), .dinb(n319), .dout(n2597));
  jand g2335(.dina(n1542), .dinb(n265), .dout(n2598));
  jor  g2336(.dina(n2598), .dinb(n2597), .dout(n2599));
  jand g2337(.dina(n1490), .dinb(n364), .dout(n2600));
  jor  g2338(.dina(n2600), .dinb(n2599), .dout(n2601));
  jor  g2339(.dina(n2601), .dinb(n2596), .dout(n2602));
  jor  g2340(.dina(n2602), .dinb(shift6 ), .dout(n2603));
  jand g2341(.dina(n2603), .dinb(n2595), .dout(result38 ));
  jand g2342(.dina(n1588), .dinb(n410), .dout(n2605));
  jand g2343(.dina(n1599), .dinb(n319), .dout(n2606));
  jand g2344(.dina(n1579), .dinb(n265), .dout(n2607));
  jor  g2345(.dina(n2607), .dinb(n2606), .dout(n2608));
  jand g2346(.dina(n1615), .dinb(n364), .dout(n2609));
  jor  g2347(.dina(n2609), .dinb(n2608), .dout(n2610));
  jor  g2348(.dina(n2610), .dinb(n2605), .dout(n2611));
  jor  g2349(.dina(n2611), .dinb(n263), .dout(n2612));
  jand g2350(.dina(n1571), .dinb(n319), .dout(n2613));
  jand g2351(.dina(n1607), .dinb(n410), .dout(n2614));
  jand g2352(.dina(n1563), .dinb(n364), .dout(n2615));
  jor  g2353(.dina(n2615), .dinb(n2614), .dout(n2616));
  jand g2354(.dina(n1624), .dinb(n265), .dout(n2617));
  jor  g2355(.dina(n2617), .dinb(n2616), .dout(n2618));
  jor  g2356(.dina(n2618), .dinb(n2613), .dout(n2619));
  jor  g2357(.dina(n2619), .dinb(shift6 ), .dout(n2620));
  jand g2358(.dina(n2620), .dinb(n2612), .dout(result39 ));
  jand g2359(.dina(n1661), .dinb(n410), .dout(n2622));
  jand g2360(.dina(n1672), .dinb(n319), .dout(n2623));
  jand g2361(.dina(n1697), .dinb(n364), .dout(n2624));
  jor  g2362(.dina(n2624), .dinb(n2623), .dout(n2625));
  jand g2363(.dina(n1652), .dinb(n265), .dout(n2626));
  jor  g2364(.dina(n2626), .dinb(n2625), .dout(n2627));
  jor  g2365(.dina(n2627), .dinb(n2622), .dout(n2628));
  jor  g2366(.dina(n2628), .dinb(n263), .dout(n2629));
  jand g2367(.dina(n1688), .dinb(n265), .dout(n2630));
  jand g2368(.dina(n1680), .dinb(n410), .dout(n2631));
  jand g2369(.dina(n1636), .dinb(n364), .dout(n2632));
  jor  g2370(.dina(n2632), .dinb(n2631), .dout(n2633));
  jand g2371(.dina(n1644), .dinb(n319), .dout(n2634));
  jor  g2372(.dina(n2634), .dinb(n2633), .dout(n2635));
  jor  g2373(.dina(n2635), .dinb(n2630), .dout(n2636));
  jor  g2374(.dina(n2636), .dinb(shift6 ), .dout(n2637));
  jand g2375(.dina(n2637), .dinb(n2629), .dout(result40 ));
  jand g2376(.dina(n1709), .dinb(n265), .dout(n2639));
  jand g2377(.dina(n1770), .dinb(n319), .dout(n2640));
  jand g2378(.dina(n1745), .dinb(n364), .dout(n2641));
  jor  g2379(.dina(n2641), .dinb(n2640), .dout(n2642));
  jand g2380(.dina(n1734), .dinb(n410), .dout(n2643));
  jor  g2381(.dina(n2643), .dinb(n2642), .dout(n2644));
  jor  g2382(.dina(n2644), .dinb(n2639), .dout(n2645));
  jor  g2383(.dina(n2645), .dinb(n263), .dout(n2646));
  jand g2384(.dina(n1717), .dinb(n319), .dout(n2647));
  jand g2385(.dina(n1753), .dinb(n410), .dout(n2648));
  jand g2386(.dina(n1725), .dinb(n364), .dout(n2649));
  jor  g2387(.dina(n2649), .dinb(n2648), .dout(n2650));
  jand g2388(.dina(n1761), .dinb(n265), .dout(n2651));
  jor  g2389(.dina(n2651), .dinb(n2650), .dout(n2652));
  jor  g2390(.dina(n2652), .dinb(n2647), .dout(n2653));
  jor  g2391(.dina(n2653), .dinb(shift6 ), .dout(n2654));
  jand g2392(.dina(n2654), .dinb(n2646), .dout(result41 ));
  jand g2393(.dina(n1782), .dinb(n410), .dout(n2656));
  jand g2394(.dina(n1843), .dinb(n319), .dout(n2657));
  jand g2395(.dina(n1834), .dinb(n364), .dout(n2658));
  jor  g2396(.dina(n2658), .dinb(n2657), .dout(n2659));
  jand g2397(.dina(n1807), .dinb(n265), .dout(n2660));
  jor  g2398(.dina(n2660), .dinb(n2659), .dout(n2661));
  jor  g2399(.dina(n2661), .dinb(n2656), .dout(n2662));
  jor  g2400(.dina(n2662), .dinb(n263), .dout(n2663));
  jand g2401(.dina(n1818), .dinb(n265), .dout(n2664));
  jand g2402(.dina(n1790), .dinb(n319), .dout(n2665));
  jand g2403(.dina(n1798), .dinb(n364), .dout(n2666));
  jor  g2404(.dina(n2666), .dinb(n2665), .dout(n2667));
  jand g2405(.dina(n1826), .dinb(n410), .dout(n2668));
  jor  g2406(.dina(n2668), .dinb(n2667), .dout(n2669));
  jor  g2407(.dina(n2669), .dinb(n2664), .dout(n2670));
  jor  g2408(.dina(n2670), .dinb(shift6 ), .dout(n2671));
  jand g2409(.dina(n2671), .dinb(n2663), .dout(result42 ));
  jand g2410(.dina(n1907), .dinb(n364), .dout(n2673));
  jand g2411(.dina(n1891), .dinb(n319), .dout(n2674));
  jand g2412(.dina(n1880), .dinb(n265), .dout(n2675));
  jor  g2413(.dina(n2675), .dinb(n2674), .dout(n2676));
  jand g2414(.dina(n1855), .dinb(n410), .dout(n2677));
  jor  g2415(.dina(n2677), .dinb(n2676), .dout(n2678));
  jor  g2416(.dina(n2678), .dinb(n2673), .dout(n2679));
  jor  g2417(.dina(n2679), .dinb(n263), .dout(n2680));
  jand g2418(.dina(n1871), .dinb(n364), .dout(n2681));
  jand g2419(.dina(n1863), .dinb(n319), .dout(n2682));
  jand g2420(.dina(n1916), .dinb(n265), .dout(n2683));
  jor  g2421(.dina(n2683), .dinb(n2682), .dout(n2684));
  jand g2422(.dina(n1899), .dinb(n410), .dout(n2685));
  jor  g2423(.dina(n2685), .dinb(n2684), .dout(n2686));
  jor  g2424(.dina(n2686), .dinb(n2681), .dout(n2687));
  jor  g2425(.dina(n2687), .dinb(shift6 ), .dout(n2688));
  jand g2426(.dina(n2688), .dinb(n2680), .dout(result43 ));
  jand g2427(.dina(n1953), .dinb(n410), .dout(n2690));
  jand g2428(.dina(n1989), .dinb(n319), .dout(n2691));
  jand g2429(.dina(n1980), .dinb(n364), .dout(n2692));
  jor  g2430(.dina(n2692), .dinb(n2691), .dout(n2693));
  jand g2431(.dina(n1944), .dinb(n265), .dout(n2694));
  jor  g2432(.dina(n2694), .dinb(n2693), .dout(n2695));
  jor  g2433(.dina(n2695), .dinb(n2690), .dout(n2696));
  jor  g2434(.dina(n2696), .dinb(n263), .dout(n2697));
  jand g2435(.dina(n1964), .dinb(n265), .dout(n2698));
  jand g2436(.dina(n1936), .dinb(n319), .dout(n2699));
  jand g2437(.dina(n1928), .dinb(n364), .dout(n2700));
  jor  g2438(.dina(n2700), .dinb(n2699), .dout(n2701));
  jand g2439(.dina(n1972), .dinb(n410), .dout(n2702));
  jor  g2440(.dina(n2702), .dinb(n2701), .dout(n2703));
  jor  g2441(.dina(n2703), .dinb(n2698), .dout(n2704));
  jor  g2442(.dina(n2704), .dinb(shift6 ), .dout(n2705));
  jand g2443(.dina(n2705), .dinb(n2697), .dout(result44 ));
  jand g2444(.dina(n2017), .dinb(n265), .dout(n2707));
  jand g2445(.dina(n2037), .dinb(n319), .dout(n2708));
  jand g2446(.dina(n2062), .dinb(n364), .dout(n2709));
  jor  g2447(.dina(n2709), .dinb(n2708), .dout(n2710));
  jand g2448(.dina(n2026), .dinb(n410), .dout(n2711));
  jor  g2449(.dina(n2711), .dinb(n2710), .dout(n2712));
  jor  g2450(.dina(n2712), .dinb(n2707), .dout(n2713));
  jor  g2451(.dina(n2713), .dinb(n263), .dout(n2714));
  jand g2452(.dina(n2045), .dinb(n410), .dout(n2715));
  jand g2453(.dina(n2009), .dinb(n319), .dout(n2716));
  jand g2454(.dina(n2053), .dinb(n265), .dout(n2717));
  jor  g2455(.dina(n2717), .dinb(n2716), .dout(n2718));
  jand g2456(.dina(n2001), .dinb(n364), .dout(n2719));
  jor  g2457(.dina(n2719), .dinb(n2718), .dout(n2720));
  jor  g2458(.dina(n2720), .dinb(n2715), .dout(n2721));
  jor  g2459(.dina(n2721), .dinb(shift6 ), .dout(n2722));
  jand g2460(.dina(n2722), .dinb(n2714), .dout(result45 ));
  jand g2461(.dina(n2110), .dinb(n364), .dout(n2724));
  jand g2462(.dina(n2135), .dinb(n319), .dout(n2725));
  jand g2463(.dina(n2090), .dinb(n265), .dout(n2726));
  jor  g2464(.dina(n2726), .dinb(n2725), .dout(n2727));
  jand g2465(.dina(n2074), .dinb(n410), .dout(n2728));
  jor  g2466(.dina(n2728), .dinb(n2727), .dout(n2729));
  jor  g2467(.dina(n2729), .dinb(n2724), .dout(n2730));
  jor  g2468(.dina(n2730), .dinb(n263), .dout(n2731));
  jand g2469(.dina(n2118), .dinb(n410), .dout(n2732));
  jand g2470(.dina(n2082), .dinb(n319), .dout(n2733));
  jand g2471(.dina(n2099), .dinb(n364), .dout(n2734));
  jor  g2472(.dina(n2734), .dinb(n2733), .dout(n2735));
  jand g2473(.dina(n2126), .dinb(n265), .dout(n2736));
  jor  g2474(.dina(n2736), .dinb(n2735), .dout(n2737));
  jor  g2475(.dina(n2737), .dinb(n2732), .dout(n2738));
  jor  g2476(.dina(n2738), .dinb(shift6 ), .dout(n2739));
  jand g2477(.dina(n2739), .dinb(n2731), .dout(result46 ));
  jand g2478(.dina(n2172), .dinb(n265), .dout(n2741));
  jand g2479(.dina(n2208), .dinb(n319), .dout(n2742));
  jand g2480(.dina(n2199), .dinb(n364), .dout(n2743));
  jor  g2481(.dina(n2743), .dinb(n2742), .dout(n2744));
  jand g2482(.dina(n2147), .dinb(n410), .dout(n2745));
  jor  g2483(.dina(n2745), .dinb(n2744), .dout(n2746));
  jor  g2484(.dina(n2746), .dinb(n2741), .dout(n2747));
  jor  g2485(.dina(n2747), .dinb(n263), .dout(n2748));
  jand g2486(.dina(n2191), .dinb(n410), .dout(n2749));
  jand g2487(.dina(n2155), .dinb(n319), .dout(n2750));
  jand g2488(.dina(n2163), .dinb(n364), .dout(n2751));
  jor  g2489(.dina(n2751), .dinb(n2750), .dout(n2752));
  jand g2490(.dina(n2183), .dinb(n265), .dout(n2753));
  jor  g2491(.dina(n2753), .dinb(n2752), .dout(n2754));
  jor  g2492(.dina(n2754), .dinb(n2749), .dout(n2755));
  jor  g2493(.dina(n2755), .dinb(shift6 ), .dout(n2756));
  jand g2494(.dina(n2756), .dinb(n2748), .dout(result47 ));
  jand g2495(.dina(n410), .dinb(n407), .dout(n2758));
  jand g2496(.dina(n544), .dinb(n364), .dout(n2759));
  jand g2497(.dina(n588), .dinb(n319), .dout(n2760));
  jor  g2498(.dina(n2760), .dinb(n2759), .dout(n2761));
  jand g2499(.dina(n500), .dinb(n265), .dout(n2762));
  jor  g2500(.dina(n2762), .dinb(n2761), .dout(n2763));
  jor  g2501(.dina(n2763), .dinb(n2758), .dout(n2764));
  jor  g2502(.dina(n2764), .dinb(n263), .dout(n2765));
  jand g2503(.dina(n453), .dinb(n265), .dout(n2766));
  jand g2504(.dina(n319), .dinb(n316), .dout(n2767));
  jand g2505(.dina(n364), .dinb(n362), .dout(n2768));
  jor  g2506(.dina(n2768), .dinb(n2767), .dout(n2769));
  jand g2507(.dina(n633), .dinb(n410), .dout(n2770));
  jor  g2508(.dina(n2770), .dinb(n2769), .dout(n2771));
  jor  g2509(.dina(n2771), .dinb(n2766), .dout(n2772));
  jor  g2510(.dina(n2772), .dinb(shift6 ), .dout(n2773));
  jand g2511(.dina(n2773), .dinb(n2765), .dout(result48 ));
  jand g2512(.dina(n861), .dinb(n265), .dout(n2775));
  jand g2513(.dina(n949), .dinb(n319), .dout(n2776));
  jand g2514(.dina(n905), .dinb(n364), .dout(n2777));
  jor  g2515(.dina(n2777), .dinb(n2776), .dout(n2778));
  jand g2516(.dina(n681), .dinb(n410), .dout(n2779));
  jor  g2517(.dina(n2779), .dinb(n2778), .dout(n2780));
  jor  g2518(.dina(n2780), .dinb(n2775), .dout(n2781));
  jor  g2519(.dina(n2781), .dinb(n263), .dout(n2782));
  jand g2520(.dina(n994), .dinb(n410), .dout(n2783));
  jand g2521(.dina(n725), .dinb(n319), .dout(n2784));
  jand g2522(.dina(n769), .dinb(n265), .dout(n2785));
  jor  g2523(.dina(n2785), .dinb(n2784), .dout(n2786));
  jand g2524(.dina(n814), .dinb(n364), .dout(n2787));
  jor  g2525(.dina(n2787), .dinb(n2786), .dout(n2788));
  jor  g2526(.dina(n2788), .dinb(n2783), .dout(n2789));
  jor  g2527(.dina(n2789), .dinb(shift6 ), .dout(n2790));
  jand g2528(.dina(n2790), .dinb(n2782), .dout(result49 ));
  jand g2529(.dina(n1079), .dinb(n410), .dout(n2792));
  jand g2530(.dina(n1163), .dinb(n319), .dout(n2793));
  jand g2531(.dina(n1102), .dinb(n265), .dout(n2794));
  jor  g2532(.dina(n2794), .dinb(n2793), .dout(n2795));
  jand g2533(.dina(n1122), .dinb(n364), .dout(n2796));
  jor  g2534(.dina(n2796), .dinb(n2795), .dout(n2797));
  jor  g2535(.dina(n2797), .dinb(n2792), .dout(n2798));
  jor  g2536(.dina(n2798), .dinb(n263), .dout(n2799));
  jand g2537(.dina(n1018), .dinb(n364), .dout(n2800));
  jand g2538(.dina(n1038), .dinb(n319), .dout(n2801));
  jand g2539(.dina(n1058), .dinb(n265), .dout(n2802));
  jor  g2540(.dina(n2802), .dinb(n2801), .dout(n2803));
  jand g2541(.dina(n1142), .dinb(n410), .dout(n2804));
  jor  g2542(.dina(n2804), .dinb(n2803), .dout(n2805));
  jor  g2543(.dina(n2805), .dinb(n2800), .dout(n2806));
  jor  g2544(.dina(n2806), .dinb(shift6 ), .dout(n2807));
  jand g2545(.dina(n2807), .dinb(n2799), .dout(result50 ));
  jand g2546(.dina(n1187), .dinb(n410), .dout(n2809));
  jand g2547(.dina(n1332), .dinb(n319), .dout(n2810));
  jand g2548(.dina(n1291), .dinb(n265), .dout(n2811));
  jor  g2549(.dina(n2811), .dinb(n2810), .dout(n2812));
  jand g2550(.dina(n1271), .dinb(n364), .dout(n2813));
  jor  g2551(.dina(n2813), .dinb(n2812), .dout(n2814));
  jor  g2552(.dina(n2814), .dinb(n2809), .dout(n2815));
  jor  g2553(.dina(n2815), .dinb(n263), .dout(n2816));
  jand g2554(.dina(n1248), .dinb(n364), .dout(n2817));
  jand g2555(.dina(n1227), .dinb(n265), .dout(n2818));
  jand g2556(.dina(n1207), .dinb(n319), .dout(n2819));
  jor  g2557(.dina(n2819), .dinb(n2818), .dout(n2820));
  jand g2558(.dina(n1311), .dinb(n410), .dout(n2821));
  jor  g2559(.dina(n2821), .dinb(n2820), .dout(n2822));
  jor  g2560(.dina(n2822), .dinb(n2817), .dout(n2823));
  jor  g2561(.dina(n2823), .dinb(shift6 ), .dout(n2824));
  jand g2562(.dina(n2824), .dinb(n2816), .dout(result51 ));
  jand g2563(.dina(n1380), .dinb(n319), .dout(n2826));
  jand g2564(.dina(n1344), .dinb(n410), .dout(n2827));
  jand g2565(.dina(n1388), .dinb(n364), .dout(n2828));
  jor  g2566(.dina(n2828), .dinb(n2827), .dout(n2829));
  jand g2567(.dina(n1405), .dinb(n265), .dout(n2830));
  jor  g2568(.dina(n2830), .dinb(n2829), .dout(n2831));
  jor  g2569(.dina(n2831), .dinb(n2826), .dout(n2832));
  jor  g2570(.dina(n2832), .dinb(n263), .dout(n2833));
  jand g2571(.dina(n1360), .dinb(n319), .dout(n2834));
  jand g2572(.dina(n1352), .dinb(n265), .dout(n2835));
  jand g2573(.dina(n1396), .dinb(n410), .dout(n2836));
  jor  g2574(.dina(n2836), .dinb(n2835), .dout(n2837));
  jand g2575(.dina(n1369), .dinb(n364), .dout(n2838));
  jor  g2576(.dina(n2838), .dinb(n2837), .dout(n2839));
  jor  g2577(.dina(n2839), .dinb(n2834), .dout(n2840));
  jor  g2578(.dina(n2840), .dinb(shift6 ), .dout(n2841));
  jand g2579(.dina(n2841), .dinb(n2833), .dout(result52 ));
  jand g2580(.dina(n1453), .dinb(n265), .dout(n2843));
  jand g2581(.dina(n1442), .dinb(n410), .dout(n2844));
  jand g2582(.dina(n1469), .dinb(n319), .dout(n2845));
  jor  g2583(.dina(n2845), .dinb(n2844), .dout(n2846));
  jand g2584(.dina(n1461), .dinb(n364), .dout(n2847));
  jor  g2585(.dina(n2847), .dinb(n2846), .dout(n2848));
  jor  g2586(.dina(n2848), .dinb(n2843), .dout(n2849));
  jor  g2587(.dina(n2849), .dinb(n263), .dout(n2850));
  jand g2588(.dina(n1417), .dinb(n364), .dout(n2851));
  jand g2589(.dina(n1425), .dinb(n265), .dout(n2852));
  jand g2590(.dina(n1433), .dinb(n319), .dout(n2853));
  jor  g2591(.dina(n2853), .dinb(n2852), .dout(n2854));
  jand g2592(.dina(n1478), .dinb(n410), .dout(n2855));
  jor  g2593(.dina(n2855), .dinb(n2854), .dout(n2856));
  jor  g2594(.dina(n2856), .dinb(n2851), .dout(n2857));
  jor  g2595(.dina(n2857), .dinb(shift6 ), .dout(n2858));
  jand g2596(.dina(n2858), .dinb(n2850), .dout(result53 ));
  jand g2597(.dina(n1534), .dinb(n364), .dout(n2860));
  jand g2598(.dina(n1506), .dinb(n410), .dout(n2861));
  jand g2599(.dina(n1551), .dinb(n319), .dout(n2862));
  jor  g2600(.dina(n2862), .dinb(n2861), .dout(n2863));
  jand g2601(.dina(n1526), .dinb(n265), .dout(n2864));
  jor  g2602(.dina(n2864), .dinb(n2863), .dout(n2865));
  jor  g2603(.dina(n2865), .dinb(n2860), .dout(n2866));
  jor  g2604(.dina(n2866), .dinb(n263), .dout(n2867));
  jand g2605(.dina(n1515), .dinb(n364), .dout(n2868));
  jand g2606(.dina(n1498), .dinb(n265), .dout(n2869));
  jand g2607(.dina(n1542), .dinb(n410), .dout(n2870));
  jor  g2608(.dina(n2870), .dinb(n2869), .dout(n2871));
  jand g2609(.dina(n1490), .dinb(n319), .dout(n2872));
  jor  g2610(.dina(n2872), .dinb(n2871), .dout(n2873));
  jor  g2611(.dina(n2873), .dinb(n2868), .dout(n2874));
  jor  g2612(.dina(n2874), .dinb(shift6 ), .dout(n2875));
  jand g2613(.dina(n2875), .dinb(n2867), .dout(result54 ));
  jand g2614(.dina(n1579), .dinb(n410), .dout(n2877));
  jand g2615(.dina(n1615), .dinb(n319), .dout(n2878));
  jand g2616(.dina(n1599), .dinb(n265), .dout(n2879));
  jor  g2617(.dina(n2879), .dinb(n2878), .dout(n2880));
  jand g2618(.dina(n1607), .dinb(n364), .dout(n2881));
  jor  g2619(.dina(n2881), .dinb(n2880), .dout(n2882));
  jor  g2620(.dina(n2882), .dinb(n2877), .dout(n2883));
  jor  g2621(.dina(n2883), .dinb(n263), .dout(n2884));
  jand g2622(.dina(n1571), .dinb(n265), .dout(n2885));
  jand g2623(.dina(n1563), .dinb(n319), .dout(n2886));
  jand g2624(.dina(n1624), .dinb(n410), .dout(n2887));
  jor  g2625(.dina(n2887), .dinb(n2886), .dout(n2888));
  jand g2626(.dina(n1588), .dinb(n364), .dout(n2889));
  jor  g2627(.dina(n2889), .dinb(n2888), .dout(n2890));
  jor  g2628(.dina(n2890), .dinb(n2885), .dout(n2891));
  jor  g2629(.dina(n2891), .dinb(shift6 ), .dout(n2892));
  jand g2630(.dina(n2892), .dinb(n2884), .dout(result55 ));
  jand g2631(.dina(n1680), .dinb(n364), .dout(n2894));
  jand g2632(.dina(n1697), .dinb(n319), .dout(n2895));
  jand g2633(.dina(n1672), .dinb(n265), .dout(n2896));
  jor  g2634(.dina(n2896), .dinb(n2895), .dout(n2897));
  jand g2635(.dina(n1652), .dinb(n410), .dout(n2898));
  jor  g2636(.dina(n2898), .dinb(n2897), .dout(n2899));
  jor  g2637(.dina(n2899), .dinb(n2894), .dout(n2900));
  jor  g2638(.dina(n2900), .dinb(n263), .dout(n2901));
  jand g2639(.dina(n1688), .dinb(n410), .dout(n2902));
  jand g2640(.dina(n1636), .dinb(n319), .dout(n2903));
  jand g2641(.dina(n1644), .dinb(n265), .dout(n2904));
  jor  g2642(.dina(n2904), .dinb(n2903), .dout(n2905));
  jand g2643(.dina(n1661), .dinb(n364), .dout(n2906));
  jor  g2644(.dina(n2906), .dinb(n2905), .dout(n2907));
  jor  g2645(.dina(n2907), .dinb(n2902), .dout(n2908));
  jor  g2646(.dina(n2908), .dinb(shift6 ), .dout(n2909));
  jand g2647(.dina(n2909), .dinb(n2901), .dout(result56 ));
  jand g2648(.dina(n1770), .dinb(n265), .dout(n2911));
  jand g2649(.dina(n1745), .dinb(n319), .dout(n2912));
  jand g2650(.dina(n1753), .dinb(n364), .dout(n2913));
  jor  g2651(.dina(n2913), .dinb(n2912), .dout(n2914));
  jand g2652(.dina(n1709), .dinb(n410), .dout(n2915));
  jor  g2653(.dina(n2915), .dinb(n2914), .dout(n2916));
  jor  g2654(.dina(n2916), .dinb(n2911), .dout(n2917));
  jor  g2655(.dina(n2917), .dinb(n263), .dout(n2918));
  jand g2656(.dina(n1717), .dinb(n265), .dout(n2919));
  jand g2657(.dina(n1725), .dinb(n319), .dout(n2920));
  jand g2658(.dina(n1761), .dinb(n410), .dout(n2921));
  jor  g2659(.dina(n2921), .dinb(n2920), .dout(n2922));
  jand g2660(.dina(n1734), .dinb(n364), .dout(n2923));
  jor  g2661(.dina(n2923), .dinb(n2922), .dout(n2924));
  jor  g2662(.dina(n2924), .dinb(n2919), .dout(n2925));
  jor  g2663(.dina(n2925), .dinb(shift6 ), .dout(n2926));
  jand g2664(.dina(n2926), .dinb(n2918), .dout(result57 ));
  jand g2665(.dina(n1807), .dinb(n410), .dout(n2928));
  jand g2666(.dina(n1834), .dinb(n319), .dout(n2929));
  jand g2667(.dina(n1843), .dinb(n265), .dout(n2930));
  jor  g2668(.dina(n2930), .dinb(n2929), .dout(n2931));
  jand g2669(.dina(n1826), .dinb(n364), .dout(n2932));
  jor  g2670(.dina(n2932), .dinb(n2931), .dout(n2933));
  jor  g2671(.dina(n2933), .dinb(n2928), .dout(n2934));
  jor  g2672(.dina(n2934), .dinb(n263), .dout(n2935));
  jand g2673(.dina(n1818), .dinb(n410), .dout(n2936));
  jand g2674(.dina(n1790), .dinb(n265), .dout(n2937));
  jand g2675(.dina(n1798), .dinb(n319), .dout(n2938));
  jor  g2676(.dina(n2938), .dinb(n2937), .dout(n2939));
  jand g2677(.dina(n1782), .dinb(n364), .dout(n2940));
  jor  g2678(.dina(n2940), .dinb(n2939), .dout(n2941));
  jor  g2679(.dina(n2941), .dinb(n2936), .dout(n2942));
  jor  g2680(.dina(n2942), .dinb(shift6 ), .dout(n2943));
  jand g2681(.dina(n2943), .dinb(n2935), .dout(result58 ));
  jand g2682(.dina(n1899), .dinb(n364), .dout(n2945));
  jand g2683(.dina(n1907), .dinb(n319), .dout(n2946));
  jand g2684(.dina(n1891), .dinb(n265), .dout(n2947));
  jor  g2685(.dina(n2947), .dinb(n2946), .dout(n2948));
  jand g2686(.dina(n1880), .dinb(n410), .dout(n2949));
  jor  g2687(.dina(n2949), .dinb(n2948), .dout(n2950));
  jor  g2688(.dina(n2950), .dinb(n2945), .dout(n2951));
  jor  g2689(.dina(n2951), .dinb(n263), .dout(n2952));
  jand g2690(.dina(n1871), .dinb(n319), .dout(n2953));
  jand g2691(.dina(n1863), .dinb(n265), .dout(n2954));
  jand g2692(.dina(n1916), .dinb(n410), .dout(n2955));
  jor  g2693(.dina(n2955), .dinb(n2954), .dout(n2956));
  jand g2694(.dina(n1855), .dinb(n364), .dout(n2957));
  jor  g2695(.dina(n2957), .dinb(n2956), .dout(n2958));
  jor  g2696(.dina(n2958), .dinb(n2953), .dout(n2959));
  jor  g2697(.dina(n2959), .dinb(shift6 ), .dout(n2960));
  jand g2698(.dina(n2960), .dinb(n2952), .dout(result59 ));
  jand g2699(.dina(n1989), .dinb(n265), .dout(n2962));
  jand g2700(.dina(n1980), .dinb(n319), .dout(n2963));
  jand g2701(.dina(n1972), .dinb(n364), .dout(n2964));
  jor  g2702(.dina(n2964), .dinb(n2963), .dout(n2965));
  jand g2703(.dina(n1944), .dinb(n410), .dout(n2966));
  jor  g2704(.dina(n2966), .dinb(n2965), .dout(n2967));
  jor  g2705(.dina(n2967), .dinb(n2962), .dout(n2968));
  jor  g2706(.dina(n2968), .dinb(n263), .dout(n2969));
  jand g2707(.dina(n1928), .dinb(n319), .dout(n2970));
  jand g2708(.dina(n1936), .dinb(n265), .dout(n2971));
  jand g2709(.dina(n1964), .dinb(n410), .dout(n2972));
  jor  g2710(.dina(n2972), .dinb(n2971), .dout(n2973));
  jand g2711(.dina(n1953), .dinb(n364), .dout(n2974));
  jor  g2712(.dina(n2974), .dinb(n2973), .dout(n2975));
  jor  g2713(.dina(n2975), .dinb(n2970), .dout(n2976));
  jor  g2714(.dina(n2976), .dinb(shift6 ), .dout(n2977));
  jand g2715(.dina(n2977), .dinb(n2969), .dout(result60 ));
  jand g2716(.dina(n2037), .dinb(n265), .dout(n2979));
  jand g2717(.dina(n2062), .dinb(n319), .dout(n2980));
  jand g2718(.dina(n2045), .dinb(n364), .dout(n2981));
  jor  g2719(.dina(n2981), .dinb(n2980), .dout(n2982));
  jand g2720(.dina(n2017), .dinb(n410), .dout(n2983));
  jor  g2721(.dina(n2983), .dinb(n2982), .dout(n2984));
  jor  g2722(.dina(n2984), .dinb(n2979), .dout(n2985));
  jor  g2723(.dina(n2985), .dinb(n263), .dout(n2986));
  jand g2724(.dina(n2026), .dinb(n364), .dout(n2987));
  jand g2725(.dina(n2009), .dinb(n265), .dout(n2988));
  jand g2726(.dina(n2053), .dinb(n410), .dout(n2989));
  jor  g2727(.dina(n2989), .dinb(n2988), .dout(n2990));
  jand g2728(.dina(n2001), .dinb(n319), .dout(n2991));
  jor  g2729(.dina(n2991), .dinb(n2990), .dout(n2992));
  jor  g2730(.dina(n2992), .dinb(n2987), .dout(n2993));
  jor  g2731(.dina(n2993), .dinb(shift6 ), .dout(n2994));
  jand g2732(.dina(n2994), .dinb(n2986), .dout(result61 ));
  jand g2733(.dina(n2118), .dinb(n364), .dout(n2996));
  jand g2734(.dina(n2110), .dinb(n319), .dout(n2997));
  jand g2735(.dina(n2135), .dinb(n265), .dout(n2998));
  jor  g2736(.dina(n2998), .dinb(n2997), .dout(n2999));
  jand g2737(.dina(n2090), .dinb(n410), .dout(n3000));
  jor  g2738(.dina(n3000), .dinb(n2999), .dout(n3001));
  jor  g2739(.dina(n3001), .dinb(n2996), .dout(n3002));
  jor  g2740(.dina(n3002), .dinb(n263), .dout(n3003));
  jand g2741(.dina(n2126), .dinb(n410), .dout(n3004));
  jand g2742(.dina(n2082), .dinb(n265), .dout(n3005));
  jand g2743(.dina(n2099), .dinb(n319), .dout(n3006));
  jor  g2744(.dina(n3006), .dinb(n3005), .dout(n3007));
  jand g2745(.dina(n2074), .dinb(n364), .dout(n3008));
  jor  g2746(.dina(n3008), .dinb(n3007), .dout(n3009));
  jor  g2747(.dina(n3009), .dinb(n3004), .dout(n3010));
  jor  g2748(.dina(n3010), .dinb(shift6 ), .dout(n3011));
  jand g2749(.dina(n3011), .dinb(n3003), .dout(result62 ));
  jand g2750(.dina(n2191), .dinb(n364), .dout(n3013));
  jand g2751(.dina(n2199), .dinb(n319), .dout(n3014));
  jand g2752(.dina(n2208), .dinb(n265), .dout(n3015));
  jor  g2753(.dina(n3015), .dinb(n3014), .dout(n3016));
  jand g2754(.dina(n2172), .dinb(n410), .dout(n3017));
  jor  g2755(.dina(n3017), .dinb(n3016), .dout(n3018));
  jor  g2756(.dina(n3018), .dinb(n3013), .dout(n3019));
  jor  g2757(.dina(n3019), .dinb(n263), .dout(n3020));
  jand g2758(.dina(n2147), .dinb(n364), .dout(n3021));
  jand g2759(.dina(n2155), .dinb(n265), .dout(n3022));
  jand g2760(.dina(n2183), .dinb(n410), .dout(n3023));
  jor  g2761(.dina(n3023), .dinb(n3022), .dout(n3024));
  jand g2762(.dina(n2163), .dinb(n319), .dout(n3025));
  jor  g2763(.dina(n3025), .dinb(n3024), .dout(n3026));
  jor  g2764(.dina(n3026), .dinb(n3021), .dout(n3027));
  jor  g2765(.dina(n3027), .dinb(shift6 ), .dout(n3028));
  jand g2766(.dina(n3028), .dinb(n3020), .dout(result63 ));
  jor  g2767(.dina(n636), .dinb(n263), .dout(n3030));
  jor  g2768(.dina(n456), .dinb(shift6 ), .dout(n3031));
  jand g2769(.dina(n3031), .dinb(n3030), .dout(result64 ));
  jor  g2770(.dina(n997), .dinb(n263), .dout(n3033));
  jor  g2771(.dina(n817), .dinb(shift6 ), .dout(n3034));
  jand g2772(.dina(n3034), .dinb(n3033), .dout(result65 ));
  jor  g2773(.dina(n1166), .dinb(n263), .dout(n3036));
  jor  g2774(.dina(n1082), .dinb(shift6 ), .dout(n3037));
  jand g2775(.dina(n3037), .dinb(n3036), .dout(result66 ));
  jor  g2776(.dina(n1335), .dinb(n263), .dout(n3039));
  jor  g2777(.dina(n1251), .dinb(shift6 ), .dout(n3040));
  jand g2778(.dina(n3040), .dinb(n3039), .dout(result67 ));
  jor  g2779(.dina(n1408), .dinb(n263), .dout(n3042));
  jor  g2780(.dina(n1372), .dinb(shift6 ), .dout(n3043));
  jand g2781(.dina(n3043), .dinb(n3042), .dout(result68 ));
  jor  g2782(.dina(n1481), .dinb(n263), .dout(n3045));
  jor  g2783(.dina(n1445), .dinb(shift6 ), .dout(n3046));
  jand g2784(.dina(n3046), .dinb(n3045), .dout(result69 ));
  jor  g2785(.dina(n1554), .dinb(n263), .dout(n3048));
  jor  g2786(.dina(n1518), .dinb(shift6 ), .dout(n3049));
  jand g2787(.dina(n3049), .dinb(n3048), .dout(result70 ));
  jor  g2788(.dina(n1627), .dinb(n263), .dout(n3051));
  jor  g2789(.dina(n1591), .dinb(shift6 ), .dout(n3052));
  jand g2790(.dina(n3052), .dinb(n3051), .dout(result71 ));
  jor  g2791(.dina(n1700), .dinb(n263), .dout(n3054));
  jor  g2792(.dina(n1664), .dinb(shift6 ), .dout(n3055));
  jand g2793(.dina(n3055), .dinb(n3054), .dout(result72 ));
  jor  g2794(.dina(n1773), .dinb(n263), .dout(n3057));
  jor  g2795(.dina(n1737), .dinb(shift6 ), .dout(n3058));
  jand g2796(.dina(n3058), .dinb(n3057), .dout(result73 ));
  jor  g2797(.dina(n1846), .dinb(n263), .dout(n3060));
  jor  g2798(.dina(n1810), .dinb(shift6 ), .dout(n3061));
  jand g2799(.dina(n3061), .dinb(n3060), .dout(result74 ));
  jor  g2800(.dina(n1919), .dinb(n263), .dout(n3063));
  jor  g2801(.dina(n1883), .dinb(shift6 ), .dout(n3064));
  jand g2802(.dina(n3064), .dinb(n3063), .dout(result75 ));
  jor  g2803(.dina(n1992), .dinb(n263), .dout(n3066));
  jor  g2804(.dina(n1956), .dinb(shift6 ), .dout(n3067));
  jand g2805(.dina(n3067), .dinb(n3066), .dout(result76 ));
  jor  g2806(.dina(n2065), .dinb(n263), .dout(n3069));
  jor  g2807(.dina(n2029), .dinb(shift6 ), .dout(n3070));
  jand g2808(.dina(n3070), .dinb(n3069), .dout(result77 ));
  jor  g2809(.dina(n2138), .dinb(n263), .dout(n3072));
  jor  g2810(.dina(n2102), .dinb(shift6 ), .dout(n3073));
  jand g2811(.dina(n3073), .dinb(n3072), .dout(result78 ));
  jor  g2812(.dina(n2211), .dinb(n263), .dout(n3075));
  jor  g2813(.dina(n2175), .dinb(shift6 ), .dout(n3076));
  jand g2814(.dina(n3076), .dinb(n3075), .dout(result79 ));
  jor  g2815(.dina(n2228), .dinb(n263), .dout(n3078));
  jor  g2816(.dina(n2220), .dinb(shift6 ), .dout(n3079));
  jand g2817(.dina(n3079), .dinb(n3078), .dout(result80 ));
  jor  g2818(.dina(n2245), .dinb(n263), .dout(n3081));
  jor  g2819(.dina(n2237), .dinb(shift6 ), .dout(n3082));
  jand g2820(.dina(n3082), .dinb(n3081), .dout(result81 ));
  jor  g2821(.dina(n2262), .dinb(n263), .dout(n3084));
  jor  g2822(.dina(n2254), .dinb(shift6 ), .dout(n3085));
  jand g2823(.dina(n3085), .dinb(n3084), .dout(result82 ));
  jor  g2824(.dina(n2279), .dinb(n263), .dout(n3087));
  jor  g2825(.dina(n2271), .dinb(shift6 ), .dout(n3088));
  jand g2826(.dina(n3088), .dinb(n3087), .dout(result83 ));
  jor  g2827(.dina(n2296), .dinb(n263), .dout(n3090));
  jor  g2828(.dina(n2288), .dinb(shift6 ), .dout(n3091));
  jand g2829(.dina(n3091), .dinb(n3090), .dout(result84 ));
  jor  g2830(.dina(n2313), .dinb(n263), .dout(n3093));
  jor  g2831(.dina(n2305), .dinb(shift6 ), .dout(n3094));
  jand g2832(.dina(n3094), .dinb(n3093), .dout(result85 ));
  jor  g2833(.dina(n2330), .dinb(n263), .dout(n3096));
  jor  g2834(.dina(n2322), .dinb(shift6 ), .dout(n3097));
  jand g2835(.dina(n3097), .dinb(n3096), .dout(result86 ));
  jor  g2836(.dina(n2347), .dinb(n263), .dout(n3099));
  jor  g2837(.dina(n2339), .dinb(shift6 ), .dout(n3100));
  jand g2838(.dina(n3100), .dinb(n3099), .dout(result87 ));
  jor  g2839(.dina(n2364), .dinb(n263), .dout(n3102));
  jor  g2840(.dina(n2356), .dinb(shift6 ), .dout(n3103));
  jand g2841(.dina(n3103), .dinb(n3102), .dout(result88 ));
  jor  g2842(.dina(n2381), .dinb(n263), .dout(n3105));
  jor  g2843(.dina(n2373), .dinb(shift6 ), .dout(n3106));
  jand g2844(.dina(n3106), .dinb(n3105), .dout(result89 ));
  jor  g2845(.dina(n2398), .dinb(n263), .dout(n3108));
  jor  g2846(.dina(n2390), .dinb(shift6 ), .dout(n3109));
  jand g2847(.dina(n3109), .dinb(n3108), .dout(result90 ));
  jor  g2848(.dina(n2415), .dinb(n263), .dout(n3111));
  jor  g2849(.dina(n2407), .dinb(shift6 ), .dout(n3112));
  jand g2850(.dina(n3112), .dinb(n3111), .dout(result91 ));
  jor  g2851(.dina(n2432), .dinb(n263), .dout(n3114));
  jor  g2852(.dina(n2424), .dinb(shift6 ), .dout(n3115));
  jand g2853(.dina(n3115), .dinb(n3114), .dout(result92 ));
  jor  g2854(.dina(n2449), .dinb(n263), .dout(n3117));
  jor  g2855(.dina(n2441), .dinb(shift6 ), .dout(n3118));
  jand g2856(.dina(n3118), .dinb(n3117), .dout(result93 ));
  jor  g2857(.dina(n2466), .dinb(n263), .dout(n3120));
  jor  g2858(.dina(n2458), .dinb(shift6 ), .dout(n3121));
  jand g2859(.dina(n3121), .dinb(n3120), .dout(result94 ));
  jor  g2860(.dina(n2483), .dinb(n263), .dout(n3123));
  jor  g2861(.dina(n2475), .dinb(shift6 ), .dout(n3124));
  jand g2862(.dina(n3124), .dinb(n3123), .dout(result95 ));
  jor  g2863(.dina(n2500), .dinb(n263), .dout(n3126));
  jor  g2864(.dina(n2492), .dinb(shift6 ), .dout(n3127));
  jand g2865(.dina(n3127), .dinb(n3126), .dout(result96 ));
  jor  g2866(.dina(n2517), .dinb(n263), .dout(n3129));
  jor  g2867(.dina(n2509), .dinb(shift6 ), .dout(n3130));
  jand g2868(.dina(n3130), .dinb(n3129), .dout(result97 ));
  jor  g2869(.dina(n2534), .dinb(n263), .dout(n3132));
  jor  g2870(.dina(n2526), .dinb(shift6 ), .dout(n3133));
  jand g2871(.dina(n3133), .dinb(n3132), .dout(result98 ));
  jor  g2872(.dina(n2551), .dinb(n263), .dout(n3135));
  jor  g2873(.dina(n2543), .dinb(shift6 ), .dout(n3136));
  jand g2874(.dina(n3136), .dinb(n3135), .dout(result99 ));
  jor  g2875(.dina(n2568), .dinb(n263), .dout(n3138));
  jor  g2876(.dina(n2560), .dinb(shift6 ), .dout(n3139));
  jand g2877(.dina(n3139), .dinb(n3138), .dout(result100 ));
  jor  g2878(.dina(n2585), .dinb(n263), .dout(n3141));
  jor  g2879(.dina(n2577), .dinb(shift6 ), .dout(n3142));
  jand g2880(.dina(n3142), .dinb(n3141), .dout(result101 ));
  jor  g2881(.dina(n2602), .dinb(n263), .dout(n3144));
  jor  g2882(.dina(n2594), .dinb(shift6 ), .dout(n3145));
  jand g2883(.dina(n3145), .dinb(n3144), .dout(result102 ));
  jor  g2884(.dina(n2619), .dinb(n263), .dout(n3147));
  jor  g2885(.dina(n2611), .dinb(shift6 ), .dout(n3148));
  jand g2886(.dina(n3148), .dinb(n3147), .dout(result103 ));
  jor  g2887(.dina(n2636), .dinb(n263), .dout(n3150));
  jor  g2888(.dina(n2628), .dinb(shift6 ), .dout(n3151));
  jand g2889(.dina(n3151), .dinb(n3150), .dout(result104 ));
  jor  g2890(.dina(n2653), .dinb(n263), .dout(n3153));
  jor  g2891(.dina(n2645), .dinb(shift6 ), .dout(n3154));
  jand g2892(.dina(n3154), .dinb(n3153), .dout(result105 ));
  jor  g2893(.dina(n2670), .dinb(n263), .dout(n3156));
  jor  g2894(.dina(n2662), .dinb(shift6 ), .dout(n3157));
  jand g2895(.dina(n3157), .dinb(n3156), .dout(result106 ));
  jor  g2896(.dina(n2687), .dinb(n263), .dout(n3159));
  jor  g2897(.dina(n2679), .dinb(shift6 ), .dout(n3160));
  jand g2898(.dina(n3160), .dinb(n3159), .dout(result107 ));
  jor  g2899(.dina(n2704), .dinb(n263), .dout(n3162));
  jor  g2900(.dina(n2696), .dinb(shift6 ), .dout(n3163));
  jand g2901(.dina(n3163), .dinb(n3162), .dout(result108 ));
  jor  g2902(.dina(n2721), .dinb(n263), .dout(n3165));
  jor  g2903(.dina(n2713), .dinb(shift6 ), .dout(n3166));
  jand g2904(.dina(n3166), .dinb(n3165), .dout(result109 ));
  jor  g2905(.dina(n2738), .dinb(n263), .dout(n3168));
  jor  g2906(.dina(n2730), .dinb(shift6 ), .dout(n3169));
  jand g2907(.dina(n3169), .dinb(n3168), .dout(result110 ));
  jor  g2908(.dina(n2755), .dinb(n263), .dout(n3171));
  jor  g2909(.dina(n2747), .dinb(shift6 ), .dout(n3172));
  jand g2910(.dina(n3172), .dinb(n3171), .dout(result111 ));
  jor  g2911(.dina(n2772), .dinb(n263), .dout(n3174));
  jor  g2912(.dina(n2764), .dinb(shift6 ), .dout(n3175));
  jand g2913(.dina(n3175), .dinb(n3174), .dout(result112 ));
  jor  g2914(.dina(n2789), .dinb(n263), .dout(n3177));
  jor  g2915(.dina(n2781), .dinb(shift6 ), .dout(n3178));
  jand g2916(.dina(n3178), .dinb(n3177), .dout(result113 ));
  jor  g2917(.dina(n2806), .dinb(n263), .dout(n3180));
  jor  g2918(.dina(n2798), .dinb(shift6 ), .dout(n3181));
  jand g2919(.dina(n3181), .dinb(n3180), .dout(result114 ));
  jor  g2920(.dina(n2823), .dinb(n263), .dout(n3183));
  jor  g2921(.dina(n2815), .dinb(shift6 ), .dout(n3184));
  jand g2922(.dina(n3184), .dinb(n3183), .dout(result115 ));
  jor  g2923(.dina(n2840), .dinb(n263), .dout(n3186));
  jor  g2924(.dina(n2832), .dinb(shift6 ), .dout(n3187));
  jand g2925(.dina(n3187), .dinb(n3186), .dout(result116 ));
  jor  g2926(.dina(n2857), .dinb(n263), .dout(n3189));
  jor  g2927(.dina(n2849), .dinb(shift6 ), .dout(n3190));
  jand g2928(.dina(n3190), .dinb(n3189), .dout(result117 ));
  jor  g2929(.dina(n2874), .dinb(n263), .dout(n3192));
  jor  g2930(.dina(n2866), .dinb(shift6 ), .dout(n3193));
  jand g2931(.dina(n3193), .dinb(n3192), .dout(result118 ));
  jor  g2932(.dina(n2891), .dinb(n263), .dout(n3195));
  jor  g2933(.dina(n2883), .dinb(shift6 ), .dout(n3196));
  jand g2934(.dina(n3196), .dinb(n3195), .dout(result119 ));
  jor  g2935(.dina(n2908), .dinb(n263), .dout(n3198));
  jor  g2936(.dina(n2900), .dinb(shift6 ), .dout(n3199));
  jand g2937(.dina(n3199), .dinb(n3198), .dout(result120 ));
  jor  g2938(.dina(n2925), .dinb(n263), .dout(n3201));
  jor  g2939(.dina(n2917), .dinb(shift6 ), .dout(n3202));
  jand g2940(.dina(n3202), .dinb(n3201), .dout(result121 ));
  jor  g2941(.dina(n2942), .dinb(n263), .dout(n3204));
  jor  g2942(.dina(n2934), .dinb(shift6 ), .dout(n3205));
  jand g2943(.dina(n3205), .dinb(n3204), .dout(result122 ));
  jor  g2944(.dina(n2959), .dinb(n263), .dout(n3207));
  jor  g2945(.dina(n2951), .dinb(shift6 ), .dout(n3208));
  jand g2946(.dina(n3208), .dinb(n3207), .dout(result123 ));
  jor  g2947(.dina(n2976), .dinb(n263), .dout(n3210));
  jor  g2948(.dina(n2968), .dinb(shift6 ), .dout(n3211));
  jand g2949(.dina(n3211), .dinb(n3210), .dout(result124 ));
  jor  g2950(.dina(n2993), .dinb(n263), .dout(n3213));
  jor  g2951(.dina(n2985), .dinb(shift6 ), .dout(n3214));
  jand g2952(.dina(n3214), .dinb(n3213), .dout(result125 ));
  jor  g2953(.dina(n3010), .dinb(n263), .dout(n3216));
  jor  g2954(.dina(n3002), .dinb(shift6 ), .dout(n3217));
  jand g2955(.dina(n3217), .dinb(n3216), .dout(result126 ));
  jor  g2956(.dina(n3027), .dinb(n263), .dout(n3219));
  jor  g2957(.dina(n3019), .dinb(shift6 ), .dout(n3220));
  jand g2958(.dina(n3220), .dinb(n3219), .dout(result127 ));
endmodule


