/*

c432:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jdff: 329
	jand: 111
	jor: 110

Summary:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jdff: 329
	jand: 111
	jor: 110

The maximum logic level gap of any gate:
	c432: 8
*/

module rf_c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n43;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n150;
	wire n151;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n217;
	wire n218;
	wire n219;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n235;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n244;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n262;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G4gat_0;
	wire[2:0] w_G8gat_0;
	wire[2:0] w_G11gat_0;
	wire[2:0] w_G14gat_0;
	wire[2:0] w_G17gat_0;
	wire[2:0] w_G21gat_0;
	wire[1:0] w_G21gat_1;
	wire[1:0] w_G24gat_0;
	wire[1:0] w_G27gat_0;
	wire[1:0] w_G30gat_0;
	wire[2:0] w_G34gat_0;
	wire[2:0] w_G37gat_0;
	wire[1:0] w_G40gat_0;
	wire[2:0] w_G43gat_0;
	wire[1:0] w_G43gat_1;
	wire[1:0] w_G47gat_0;
	wire[2:0] w_G50gat_0;
	wire[1:0] w_G53gat_0;
	wire[2:0] w_G56gat_0;
	wire[2:0] w_G60gat_0;
	wire[2:0] w_G63gat_0;
	wire[1:0] w_G66gat_0;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G73gat_0;
	wire[1:0] w_G76gat_0;
	wire[1:0] w_G79gat_0;
	wire[2:0] w_G82gat_0;
	wire[2:0] w_G86gat_0;
	wire[1:0] w_G86gat_1;
	wire[2:0] w_G89gat_0;
	wire[2:0] w_G92gat_0;
	wire[2:0] w_G95gat_0;
	wire[2:0] w_G99gat_0;
	wire[2:0] w_G102gat_0;
	wire[1:0] w_G105gat_0;
	wire[2:0] w_G108gat_0;
	wire[2:0] w_G112gat_0;
	wire[1:0] w_G115gat_0;
	wire[2:0] w_G223gat_0;
	wire[2:0] w_G223gat_1;
	wire[2:0] w_G223gat_2;
	wire[1:0] w_G223gat_3;
	wire G223gat_fa_;
	wire[2:0] w_G329gat_0;
	wire[2:0] w_G329gat_1;
	wire[2:0] w_G329gat_2;
	wire[2:0] w_G329gat_3;
	wire[2:0] w_G329gat_4;
	wire[2:0] w_G329gat_5;
	wire w_G329gat_6;
	wire G329gat_fa_;
	wire[2:0] w_G370gat_0;
	wire[2:0] w_G370gat_1;
	wire w_G370gat_2;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire[1:0] w_n43_0;
	wire[1:0] w_n44_0;
	wire[1:0] w_n47_0;
	wire[1:0] w_n52_0;
	wire[1:0] w_n53_0;
	wire[1:0] w_n56_0;
	wire[1:0] w_n58_0;
	wire[1:0] w_n61_0;
	wire[1:0] w_n63_0;
	wire[1:0] w_n69_0;
	wire[1:0] w_n71_0;
	wire[1:0] w_n72_0;
	wire[1:0] w_n73_0;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[1:0] w_n79_0;
	wire[1:0] w_n82_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n87_0;
	wire[1:0] w_n89_0;
	wire[2:0] w_n94_0;
	wire[2:0] w_n94_1;
	wire[2:0] w_n94_2;
	wire[2:0] w_n94_3;
	wire[1:0] w_n94_4;
	wire[1:0] w_n96_0;
	wire[1:0] w_n98_0;
	wire[1:0] w_n100_0;
	wire[1:0] w_n107_0;
	wire[1:0] w_n109_0;
	wire[2:0] w_n114_0;
	wire[1:0] w_n115_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n121_0;
	wire[1:0] w_n123_0;
	wire[2:0] w_n126_0;
	wire[1:0] w_n128_0;
	wire[2:0] w_n130_0;
	wire[1:0] w_n132_0;
	wire[1:0] w_n139_0;
	wire[1:0] w_n141_0;
	wire[1:0] w_n142_0;
	wire[1:0] w_n145_0;
	wire[1:0] w_n146_0;
	wire[1:0] w_n147_0;
	wire[1:0] w_n150_0;
	wire[1:0] w_n151_0;
	wire[1:0] w_n154_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n159_0;
	wire[1:0] w_n164_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n174_0;
	wire[1:0] w_n177_0;
	wire[2:0] w_n182_0;
	wire[2:0] w_n182_1;
	wire[2:0] w_n182_2;
	wire[1:0] w_n182_3;
	wire[1:0] w_n184_0;
	wire[1:0] w_n188_0;
	wire[1:0] w_n191_0;
	wire[1:0] w_n193_0;
	wire[1:0] w_n197_0;
	wire[1:0] w_n198_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n205_0;
	wire[1:0] w_n217_0;
	wire[1:0] w_n219_0;
	wire[1:0] w_n222_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n231_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n260_0;
	wire[2:0] w_n271_0;
	wire[2:0] w_n271_1;
	wire[2:0] w_n271_2;
	wire[1:0] w_n271_3;
	wire[1:0] w_n274_0;
	wire[1:0] w_n281_0;
	wire[1:0] w_n283_0;
	wire[1:0] w_n286_0;
	wire[1:0] w_n290_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n296_0;
	wire[1:0] w_n303_0;
	wire[1:0] w_n305_0;
	wire[1:0] w_n313_0;
	wire[1:0] w_n314_0;
	wire[2:0] w_n317_0;
	wire[1:0] w_n319_0;
	wire w_dff_B_XtHeAfHt3_1;
	wire w_dff_B_mU4a1R0G9_1;
	wire w_dff_B_rtAp55pV5_1;
	wire w_dff_B_zXWR4QiJ6_0;
	wire w_dff_B_nHXfgPoY1_0;
	wire w_dff_B_bNEI4rL86_0;
	wire w_dff_B_IMDGVjcC1_0;
	wire w_dff_B_aRJZPg1J1_0;
	wire w_dff_B_iDU98mng5_1;
	wire w_dff_A_WEGfJ7D77_0;
	wire w_dff_B_2fu6BJoY9_0;
	wire w_dff_B_yGPvgfJt3_0;
	wire w_dff_B_9Xu2oV544_0;
	wire w_dff_B_nTjcGx367_0;
	wire w_dff_B_XsdkV8eb0_0;
	wire w_dff_A_CPVisDct8_0;
	wire w_dff_B_Cy7OM6LL8_1;
	wire w_dff_B_Tz57h5cV9_0;
	wire w_dff_B_vvFGQoVh3_0;
	wire w_dff_B_LZ0A1fIT9_0;
	wire w_dff_B_Fgsm36Nb6_0;
	wire w_dff_B_dr6xUBbA2_0;
	wire w_dff_A_ZCGVbZ6j3_0;
	wire w_dff_A_hPDd8nNh7_0;
	wire w_dff_A_62pZ9gad9_0;
	wire w_dff_A_LP1iDE6J0_0;
	wire w_dff_A_lX0tC26d5_0;
	wire w_dff_A_6NAHzLAd6_0;
	wire w_dff_A_w4LmiAQl5_0;
	wire w_dff_B_5YqJoV4e2_1;
	wire w_dff_B_k5ymrU9g7_1;
	wire w_dff_B_MXFl03cr1_1;
	wire w_dff_B_6vj4xBQp7_1;
	wire w_dff_B_VsfiNflG8_1;
	wire w_dff_B_SLaXVEXg4_1;
	wire w_dff_B_a73vCTRQ3_1;
	wire w_dff_B_H0wA1PPA9_1;
	wire w_dff_B_y6aSXzkD7_1;
	wire w_dff_B_CH96FsCJ4_1;
	wire w_dff_B_VbQXb5dF0_1;
	wire w_dff_B_AVqRZJd08_1;
	wire w_dff_B_CHTtVXaK8_1;
	wire w_dff_B_Vvdh6JPd3_1;
	wire w_dff_B_9t1Ri9rA7_1;
	wire w_dff_B_29msO7Ij6_1;
	wire w_dff_B_TP2ysv185_1;
	wire w_dff_B_kOZLYA213_1;
	wire w_dff_B_4CizjBJQ7_1;
	wire w_dff_B_7d2hg9nE5_1;
	wire w_dff_B_t64QZ5Sx5_1;
	wire w_dff_B_stNHmWmI6_1;
	wire w_dff_B_ElDv60aw7_1;
	wire w_dff_B_1fsV7m6g8_1;
	wire w_dff_B_dXfHzVvI2_1;
	wire w_dff_B_YuoYgjBp9_1;
	wire w_dff_B_Le00bwyL1_1;
	wire w_dff_B_FissYN5J5_0;
	wire w_dff_B_9gYMrj778_0;
	wire w_dff_B_cwhqTbIK1_0;
	wire w_dff_A_uSygbgaG4_1;
	wire w_dff_A_lX7HOrsH8_1;
	wire w_dff_A_UIBVQYQS0_1;
	wire w_dff_A_QGG2jtbD0_1;
	wire w_dff_A_PSVXGahE5_1;
	wire w_dff_A_401m6pOU5_1;
	wire w_dff_B_JYpo5TJY7_1;
	wire w_dff_B_WNoS3vJn2_0;
	wire w_dff_B_xXpzcbdI5_0;
	wire w_dff_B_5pVV6fYM3_0;
	wire w_dff_B_nwK4xXoc8_0;
	wire w_dff_B_LU7xsRHL2_0;
	wire w_dff_B_PJdAhUWv3_1;
	wire w_dff_B_N0MoOT9q2_0;
	wire w_dff_B_Wmb5Vblx7_0;
	wire w_dff_B_1tvf18FW4_0;
	wire w_dff_B_rOrn4pq43_0;
	wire w_dff_A_fy0OtTh78_0;
	wire w_dff_A_06P2op1q6_0;
	wire w_dff_A_Auye3inr6_0;
	wire w_dff_A_VfJ30puZ9_0;
	wire w_dff_A_ZtLsp5To9_0;
	wire w_dff_A_Io8wu6CR0_0;
	wire w_dff_A_mDAUDbsT8_0;
	wire w_dff_A_dmfuDBAc4_0;
	wire w_dff_A_fakqwGEj0_0;
	wire w_dff_A_qMYvcXrW2_0;
	wire w_dff_A_lHtqvvXo0_0;
	wire w_dff_A_RDuB9J604_0;
	wire w_dff_A_KiXnnO0H1_0;
	wire w_dff_A_rRNuASCT2_0;
	wire w_dff_A_k3ABFhLk2_0;
	wire w_dff_A_TWJ76dEY2_0;
	wire w_dff_A_EOkWvfXL5_0;
	wire w_dff_A_elp8uBYG5_0;
	wire w_dff_B_0pQmMgYh3_0;
	wire w_dff_B_Ei3srVPx3_0;
	wire w_dff_B_FfSBo8dk2_0;
	wire w_dff_B_3GouIE3F3_0;
	wire w_dff_B_zut9mmyo8_0;
	wire w_dff_B_GD1r0xmC1_0;
	wire w_dff_B_8MFLnt5m9_1;
	wire w_dff_B_VWnVZ5F89_1;
	wire w_dff_B_ErEIblJx5_1;
	wire w_dff_A_jAzNkW4y0_0;
	wire w_dff_A_Z94B9Lvk9_0;
	wire w_dff_A_hwgTDZLm7_0;
	wire w_dff_A_xhCE7X622_0;
	wire w_dff_A_nkxJFDy28_0;
	wire w_dff_A_HQnMQAMg9_0;
	wire w_dff_A_Wh1RiAQx6_0;
	wire w_dff_A_UjGwj7CU3_0;
	wire w_dff_A_ALys9RFq4_0;
	wire w_dff_A_31UNmNVu2_0;
	wire w_dff_A_CYPpKWXV4_0;
	wire w_dff_B_qg7mWGb20_2;
	wire w_dff_B_MW5gfkNF4_2;
	wire w_dff_B_rsVgH1GT7_2;
	wire w_dff_B_o2BQCpRe8_2;
	wire w_dff_B_Ak0plN7W2_2;
	wire w_dff_B_2qaQWBAQ4_2;
	wire w_dff_B_yjhHwxmA9_2;
	wire w_dff_B_fFVjhWS68_2;
	wire w_dff_B_woW1UOno0_2;
	wire w_dff_B_ivtfX5JB3_2;
	wire w_dff_B_Vqrr3Xeq4_2;
	wire w_dff_B_hfXbhLSj7_2;
	wire w_dff_B_TqRYiniu7_2;
	wire w_dff_B_tiu2edyZ9_2;
	wire w_dff_B_FyFM8Ygp2_1;
	wire w_dff_B_eNrwTtNg3_1;
	wire w_dff_B_yggQB6Ys8_1;
	wire w_dff_B_U0MpGuxn5_1;
	wire w_dff_B_NYlgNJl09_1;
	wire w_dff_B_x5QkcuRc4_1;
	wire w_dff_B_HcES8P0P0_1;
	wire w_dff_B_ppmixOzB9_1;
	wire w_dff_B_vmiTmYiF4_1;
	wire w_dff_B_OYUCZ4l41_1;
	wire w_dff_B_aHMr6rBz7_1;
	wire w_dff_B_QLbN3OC24_1;
	wire w_dff_B_AM95yKvk0_1;
	wire w_dff_B_CHp7zuqa4_1;
	wire w_dff_B_Y2xHbUVu2_1;
	wire w_dff_B_laHDFc1W2_1;
	wire w_dff_B_kGyIrKsw1_1;
	wire w_dff_B_KgFU634u2_1;
	wire w_dff_B_My7Aav3g5_1;
	wire w_dff_B_ngP0PGs45_1;
	wire w_dff_B_I2tvJizq0_1;
	wire w_dff_B_moXcOpP59_1;
	wire w_dff_B_CxDoqWCF9_1;
	wire w_dff_B_bQ8DlPv90_1;
	wire w_dff_B_NKML2GtR0_1;
	wire w_dff_B_9K2odaVq1_1;
	wire w_dff_A_zbikquwd1_0;
	wire w_dff_A_QVn7yNck3_0;
	wire w_dff_A_n0TYYcXN6_0;
	wire w_dff_A_ECPX5BkF9_0;
	wire w_dff_A_A6r9DdmE6_0;
	wire w_dff_A_aR5lBUSR9_0;
	wire w_dff_B_EMSPp0NZ0_2;
	wire w_dff_B_hQvT0f3E4_2;
	wire w_dff_B_25WKhGGk9_2;
	wire w_dff_B_mh33z2Yd4_2;
	wire w_dff_B_uQoBKJ9X1_2;
	wire w_dff_B_5kEo7zCX8_2;
	wire w_dff_B_9kmsZGCh0_2;
	wire w_dff_B_pXCl8kXn9_2;
	wire w_dff_B_k24UfNbR5_2;
	wire w_dff_B_izS80gCz9_2;
	wire w_dff_B_kemnXx8M0_2;
	wire w_dff_B_R3jnqyQA0_2;
	wire w_dff_B_4HksJLIe0_2;
	wire w_dff_A_uViN6cTm4_0;
	wire w_dff_A_nnKjElT53_0;
	wire w_dff_A_vbNNgIQg3_0;
	wire w_dff_A_Ah0ngBQz4_0;
	wire w_dff_A_Qbd9lZ5L1_0;
	wire w_dff_A_0CZK0CXH3_0;
	wire w_dff_A_r845OfmA6_0;
	wire w_dff_A_eCkCE2r60_0;
	wire w_dff_A_Laa5sYIB7_0;
	wire w_dff_A_360d4E9j8_0;
	wire w_dff_A_6lc62de52_0;
	wire w_dff_A_r64e4DY39_0;
	wire w_dff_B_VBOZ7g2j6_2;
	wire w_dff_B_eV0S1xYl3_2;
	wire w_dff_B_KPEBxuUq7_2;
	wire w_dff_B_CEDaHPVs2_2;
	wire w_dff_B_cqlO6qAm3_2;
	wire w_dff_B_ZBpyvRCx3_2;
	wire w_dff_B_bi592kgC7_2;
	wire w_dff_B_l1YZ9jLP0_2;
	wire w_dff_B_uG2bxopE2_2;
	wire w_dff_B_3BRfc02z0_2;
	wire w_dff_B_dh96HMii8_2;
	wire w_dff_B_yLoxZPxV0_2;
	wire w_dff_B_dCAN8GhJ7_2;
	wire w_dff_A_6tWAUU271_0;
	wire w_dff_A_6WZoJxMl3_0;
	wire w_dff_A_2Eqx7S8l2_0;
	wire w_dff_A_PYtGB0pE4_0;
	wire w_dff_A_pVQUDdVA1_0;
	wire w_dff_A_FVGC99NZ8_0;
	wire w_dff_A_4TF5M3ij0_0;
	wire w_dff_A_7kQZIIpO5_0;
	wire w_dff_A_K3LifHUO9_0;
	wire w_dff_A_1bHFImJt9_0;
	wire w_dff_A_JQPDQPyt7_0;
	wire w_dff_A_0jaXmlQm8_0;
	wire w_dff_B_30JJ7VWd1_1;
	wire w_dff_A_0Kr7sAnf0_0;
	wire w_dff_A_3FKVdAia8_0;
	wire w_dff_A_6dUHppkX9_0;
	wire w_dff_A_caFBgMjP5_0;
	wire w_dff_A_Cg9vU7Wc4_0;
	wire w_dff_A_GeqVoK4M6_0;
	wire w_dff_A_hTuuCm4F8_0;
	wire w_dff_A_s5PcXhe91_0;
	wire w_dff_A_Zd29BN252_0;
	wire w_dff_A_2sWQGN515_0;
	wire w_dff_A_OJmXFrQB0_0;
	wire w_dff_A_RISmnG7W4_0;
	wire w_dff_B_sda6iCdK6_1;
	wire w_dff_B_8UbO43Uq1_1;
	wire w_dff_B_KDKRnPY56_1;
	wire w_dff_B_bLrzaVhU1_1;
	wire w_dff_B_yRRxXC9F0_1;
	wire w_dff_B_6pAiUECP2_1;
	wire w_dff_A_uOjPQsTM7_0;
	wire w_dff_A_FhGZDlhD1_0;
	wire w_dff_A_Sz5H8gib4_0;
	wire w_dff_A_y5ZGbqtw9_0;
	wire w_dff_B_5Z31j0s29_2;
	wire w_dff_A_qRBfRAPu7_0;
	wire w_dff_A_PefwWC5e3_0;
	wire w_dff_A_Py2NcyGQ4_0;
	wire w_dff_A_g0hdhvdd4_0;
	wire w_dff_A_PuumVz3v9_0;
	wire w_dff_A_H9jgYljp9_0;
	wire w_dff_A_FbOkL3oh9_0;
	wire w_dff_A_LB8qNsp02_0;
	wire w_dff_A_N6GA9OXz6_0;
	wire w_dff_A_7jkH8cLA8_0;
	wire w_dff_A_yDCvhztt5_0;
	wire w_dff_A_SXewAdwv0_0;
	wire w_dff_A_tgyV8E6r7_0;
	wire w_dff_A_1Jq4nkXF1_0;
	wire w_dff_A_yJLP9fDB7_0;
	wire w_dff_A_bIl8ee3p0_0;
	wire w_dff_A_WQ2gkHU33_0;
	wire w_dff_A_CZVKhSoJ6_0;
	wire w_dff_A_lPNB9SXU5_0;
	wire w_dff_A_7Ts3aUSM7_0;
	wire w_dff_A_f1iMwhNx3_0;
	wire w_dff_A_FZkAdwT63_0;
	wire w_dff_A_KANBbx909_0;
	wire w_dff_B_MIhgDrZp5_2;
	wire w_dff_B_QuZuGzNj1_2;
	wire w_dff_B_vuG75snK7_2;
	wire w_dff_B_AbNuQma71_2;
	wire w_dff_B_Zkvwf1hd9_2;
	wire w_dff_B_1k3jrDMp1_2;
	wire w_dff_B_3eMPSOt68_2;
	wire w_dff_B_jGDwblWz6_2;
	wire w_dff_B_bcqC3Odf5_2;
	wire w_dff_B_UNxknqTt3_2;
	wire w_dff_B_QNKmPUo10_2;
	wire w_dff_B_V9oMdfJU2_2;
	wire w_dff_B_lDNCmbYg3_2;
	wire w_dff_B_R2JwCoqq6_2;
	wire w_dff_A_g6hg80xF5_1;
	wire w_dff_A_6uNmkRof2_1;
	wire w_dff_A_T4EavMuv3_1;
	wire w_dff_A_iDTa47vb4_1;
	wire w_dff_A_Sd3vZQAW8_0;
	wire w_dff_A_TWd66Ggc0_0;
	wire w_dff_A_ZFkON3pV8_0;
	wire w_dff_A_tC9e8ZTm8_0;
	wire w_dff_A_Tv1nYxhP5_0;
	wire w_dff_A_HK2fndwt2_0;
	wire w_dff_A_HeeEoTy64_0;
	wire w_dff_A_n5GzK4zV6_1;
	wire w_dff_A_DoLX5AFt6_1;
	wire w_dff_A_YaurMj0r3_1;
	wire w_dff_A_F6Ecdgn17_1;
	wire w_dff_A_O5uDvHnT1_1;
	wire w_dff_A_4wpWuhcS5_1;
	wire w_dff_A_U2myqVlw1_2;
	wire w_dff_A_r1PolYoN8_0;
	wire w_dff_A_npYM2eh68_0;
	wire w_dff_A_vxUEi8dk1_0;
	wire w_dff_A_oDi1ha292_0;
	wire w_dff_A_LP3ezWcE7_0;
	wire w_dff_A_5IA7FVEp8_0;
	wire w_dff_A_rUXUmbIs5_0;
	wire w_dff_A_WfCN4ii01_0;
	wire w_dff_A_FEVZJuwM1_0;
	wire w_dff_A_qrQbfMeW7_0;
	wire w_dff_A_LDgfQkT33_0;
	wire w_dff_A_Rn7gZ7Wo9_0;
	wire w_dff_A_ILLmIjGa0_0;
	wire w_dff_A_ThmFGEWB0_0;
	wire w_dff_A_IbJyhUjl3_0;
	wire w_dff_A_drZFLKzm1_0;
	wire w_dff_A_DHS1iso26_0;
	wire w_dff_A_BntL2tG77_0;
	wire w_dff_A_PCOFOU9c5_0;
	wire w_dff_A_6BlOj4PO6_1;
	wire w_dff_A_gJ9QO1IN4_0;
	wire w_dff_A_YyOfjQmG0_0;
	wire w_dff_A_VNlNLTow8_0;
	wire w_dff_A_ei14NpkH3_0;
	wire w_dff_A_nXsGjgZx3_0;
	wire w_dff_A_PEk6LAkq2_0;
	wire w_dff_A_geYzOqFe7_0;
	wire w_dff_A_OewmXfb11_0;
	wire w_dff_A_HoXvt9rV9_0;
	wire w_dff_A_4pRC4xYS3_0;
	wire w_dff_A_mWAVF39O0_0;
	wire w_dff_A_zFdNpgDY2_0;
	wire w_dff_A_iURVVgb10_1;
	wire w_dff_A_6oMFTJmt9_0;
	wire w_dff_A_Z3cxfR5c0_0;
	wire w_dff_A_T4u4e5Ml8_0;
	wire w_dff_A_zyEgun1U8_0;
	wire w_dff_A_l0pFLbh48_0;
	wire w_dff_A_C8M0FakO9_1;
	wire w_dff_A_gmAmFeKr4_0;
	jnot g000(.din(w_G76gat_0[1]),.dout(n43),.clk(gclk));
	jand g001(.dina(w_G82gat_0[2]),.dinb(w_n43_0[1]),.dout(n44),.clk(gclk));
	jnot g002(.din(w_G24gat_0[1]),.dout(n45),.clk(gclk));
	jand g003(.dina(w_G30gat_0[1]),.dinb(n45),.dout(n46),.clk(gclk));
	jnot g004(.din(w_G11gat_0[2]),.dout(n47),.clk(gclk));
	jand g005(.dina(w_G17gat_0[2]),.dinb(w_n47_0[1]),.dout(n48),.clk(gclk));
	jor g006(.dina(n48),.dinb(n46),.dout(n49),.clk(gclk));
	jor g007(.dina(n49),.dinb(w_n44_0[1]),.dout(n50),.clk(gclk));
	jnot g008(.din(w_G37gat_0[2]),.dout(n51),.clk(gclk));
	jand g009(.dina(w_G43gat_1[1]),.dinb(n51),.dout(n52),.clk(gclk));
	jnot g010(.din(w_G63gat_0[2]),.dout(n53),.clk(gclk));
	jand g011(.dina(w_G69gat_0[2]),.dinb(w_n53_0[1]),.dout(n54),.clk(gclk));
	jor g012(.dina(n54),.dinb(w_n52_0[1]),.dout(n55),.clk(gclk));
	jnot g013(.din(w_G102gat_0[2]),.dout(n56),.clk(gclk));
	jand g014(.dina(w_G108gat_0[2]),.dinb(w_n56_0[1]),.dout(n57),.clk(gclk));
	jnot g015(.din(w_G50gat_0[2]),.dout(n58),.clk(gclk));
	jand g016(.dina(w_G56gat_0[2]),.dinb(w_n58_0[1]),.dout(n59),.clk(gclk));
	jor g017(.dina(n59),.dinb(n57),.dout(n60),.clk(gclk));
	jnot g018(.din(w_G89gat_0[2]),.dout(n61),.clk(gclk));
	jand g019(.dina(w_G95gat_0[2]),.dinb(w_n61_0[1]),.dout(n62),.clk(gclk));
	jnot g020(.din(w_G1gat_0[2]),.dout(n63),.clk(gclk));
	jand g021(.dina(w_G4gat_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jor g022(.dina(n64),.dinb(n62),.dout(n65),.clk(gclk));
	jor g023(.dina(n65),.dinb(n60),.dout(n66),.clk(gclk));
	jor g024(.dina(n66),.dinb(n55),.dout(n67),.clk(gclk));
	jor g025(.dina(n67),.dinb(n50),.dout(G223gat_fa_),.clk(gclk));
	jnot g026(.din(w_G112gat_0[2]),.dout(n69),.clk(gclk));
	jnot g027(.din(w_n44_0[0]),.dout(n70),.clk(gclk));
	jnot g028(.din(w_G30gat_0[0]),.dout(n71),.clk(gclk));
	jor g029(.dina(w_n71_0[1]),.dinb(w_G24gat_0[0]),.dout(n72),.clk(gclk));
	jnot g030(.din(w_G17gat_0[1]),.dout(n73),.clk(gclk));
	jor g031(.dina(w_n73_0[1]),.dinb(w_G11gat_0[1]),.dout(n74),.clk(gclk));
	jand g032(.dina(n74),.dinb(w_n72_0[1]),.dout(n75),.clk(gclk));
	jand g033(.dina(n75),.dinb(n70),.dout(n76),.clk(gclk));
	jnot g034(.din(w_G43gat_1[0]),.dout(n77),.clk(gclk));
	jor g035(.dina(w_n77_0[1]),.dinb(w_G37gat_0[1]),.dout(n78),.clk(gclk));
	jnot g036(.din(w_G69gat_0[1]),.dout(n79),.clk(gclk));
	jor g037(.dina(w_n79_0[1]),.dinb(w_G63gat_0[1]),.dout(n80),.clk(gclk));
	jand g038(.dina(n80),.dinb(w_n78_0[1]),.dout(n81),.clk(gclk));
	jnot g039(.din(w_G108gat_0[1]),.dout(n82),.clk(gclk));
	jor g040(.dina(w_n82_0[1]),.dinb(w_G102gat_0[1]),.dout(n83),.clk(gclk));
	jnot g041(.din(w_G56gat_0[1]),.dout(n84),.clk(gclk));
	jor g042(.dina(w_n84_0[1]),.dinb(w_G50gat_0[1]),.dout(n85),.clk(gclk));
	jand g043(.dina(n85),.dinb(n83),.dout(n86),.clk(gclk));
	jnot g044(.din(w_G95gat_0[1]),.dout(n87),.clk(gclk));
	jor g045(.dina(w_n87_0[1]),.dinb(w_G89gat_0[1]),.dout(n88),.clk(gclk));
	jnot g046(.din(w_G4gat_0[1]),.dout(n89),.clk(gclk));
	jor g047(.dina(w_n89_0[1]),.dinb(w_G1gat_0[1]),.dout(n90),.clk(gclk));
	jand g048(.dina(n90),.dinb(n88),.dout(n91),.clk(gclk));
	jand g049(.dina(n91),.dinb(n86),.dout(n92),.clk(gclk));
	jand g050(.dina(n92),.dinb(n81),.dout(n93),.clk(gclk));
	jand g051(.dina(n93),.dinb(n76),.dout(n94),.clk(gclk));
	jor g052(.dina(w_n94_4[1]),.dinb(w_n56_0[0]),.dout(n95),.clk(gclk));
	jand g053(.dina(n95),.dinb(w_G108gat_0[0]),.dout(n96),.clk(gclk));
	jand g054(.dina(w_n96_0[1]),.dinb(w_n69_0[1]),.dout(n97),.clk(gclk));
	jnot g055(.din(w_G8gat_0[2]),.dout(n98),.clk(gclk));
	jor g056(.dina(w_n94_4[0]),.dinb(w_n63_0[0]),.dout(n99),.clk(gclk));
	jand g057(.dina(n99),.dinb(w_G4gat_0[0]),.dout(n100),.clk(gclk));
	jand g058(.dina(w_n100_0[1]),.dinb(w_n98_0[1]),.dout(n101),.clk(gclk));
	jor g059(.dina(n101),.dinb(n97),.dout(n102),.clk(gclk));
	jnot g060(.din(w_G99gat_0[2]),.dout(n103),.clk(gclk));
	jor g061(.dina(w_n94_3[2]),.dinb(w_n61_0[0]),.dout(n104),.clk(gclk));
	jand g062(.dina(n104),.dinb(w_G95gat_0[0]),.dout(n105),.clk(gclk));
	jand g063(.dina(n105),.dinb(n103),.dout(n106),.clk(gclk));
	jnot g064(.din(w_G73gat_0[2]),.dout(n107),.clk(gclk));
	jor g065(.dina(w_n94_3[1]),.dinb(w_n53_0[0]),.dout(n108),.clk(gclk));
	jand g066(.dina(n108),.dinb(w_G69gat_0[0]),.dout(n109),.clk(gclk));
	jand g067(.dina(w_n109_0[1]),.dinb(w_n107_0[1]),.dout(n110),.clk(gclk));
	jor g068(.dina(n110),.dinb(n106),.dout(n111),.clk(gclk));
	jor g069(.dina(n111),.dinb(n102),.dout(n112),.clk(gclk));
	jxor g070(.dina(w_n94_3[0]),.dinb(w_n72_0[0]),.dout(n113),.clk(gclk));
	jor g071(.dina(n113),.dinb(w_n71_0[0]),.dout(n114),.clk(gclk));
	jor g072(.dina(w_n114_0[2]),.dinb(w_G34gat_0[2]),.dout(n115),.clk(gclk));
	jnot g073(.din(w_n115_0[1]),.dout(n116),.clk(gclk));
	jnot g074(.din(w_G60gat_0[2]),.dout(n117),.clk(gclk));
	jor g075(.dina(w_n94_2[2]),.dinb(w_n58_0[0]),.dout(n118),.clk(gclk));
	jand g076(.dina(n118),.dinb(w_G56gat_0[0]),.dout(n119),.clk(gclk));
	jand g077(.dina(w_n119_0[1]),.dinb(n117),.dout(n120),.clk(gclk));
	jxor g078(.dina(w_n94_2[1]),.dinb(w_n52_0[0]),.dout(n121),.clk(gclk));
	jnot g079(.din(w_G47gat_0[1]),.dout(n122),.clk(gclk));
	jand g080(.dina(n122),.dinb(w_G43gat_0[2]),.dout(n123),.clk(gclk));
	jand g081(.dina(w_n123_0[1]),.dinb(w_n121_0[1]),.dout(n124),.clk(gclk));
	jor g082(.dina(n124),.dinb(n120),.dout(n125),.clk(gclk));
	jnot g083(.din(w_G86gat_1[1]),.dout(n126),.clk(gclk));
	jor g084(.dina(w_n94_2[0]),.dinb(w_n43_0[0]),.dout(n127),.clk(gclk));
	jand g085(.dina(n127),.dinb(w_G82gat_0[1]),.dout(n128),.clk(gclk));
	jand g086(.dina(w_n128_0[1]),.dinb(w_n126_0[2]),.dout(n129),.clk(gclk));
	jnot g087(.din(w_G21gat_1[1]),.dout(n130),.clk(gclk));
	jor g088(.dina(w_n94_1[2]),.dinb(w_n47_0[0]),.dout(n131),.clk(gclk));
	jand g089(.dina(n131),.dinb(w_G17gat_0[0]),.dout(n132),.clk(gclk));
	jand g090(.dina(w_n132_0[1]),.dinb(w_n130_0[2]),.dout(n133),.clk(gclk));
	jor g091(.dina(n133),.dinb(n129),.dout(n134),.clk(gclk));
	jor g092(.dina(n134),.dinb(n125),.dout(n135),.clk(gclk));
	jor g093(.dina(n135),.dinb(n116),.dout(n136),.clk(gclk));
	jor g094(.dina(n136),.dinb(n112),.dout(G329gat_fa_),.clk(gclk));
	jand g095(.dina(w_G223gat_3[1]),.dinb(w_G89gat_0[0]),.dout(n138),.clk(gclk));
	jor g096(.dina(n138),.dinb(w_n87_0[0]),.dout(n139),.clk(gclk));
	jand g097(.dina(w_G329gat_6),.dinb(w_G99gat_0[1]),.dout(n140),.clk(gclk));
	jor g098(.dina(n140),.dinb(w_n139_0[1]),.dout(n141),.clk(gclk));
	jor g099(.dina(w_n141_0[1]),.dinb(w_G105gat_0[1]),.dout(n142),.clk(gclk));
	jnot g100(.din(w_n142_0[1]),.dout(n143),.clk(gclk));
	jand g101(.dina(w_G223gat_3[0]),.dinb(w_G50gat_0[0]),.dout(n144),.clk(gclk));
	jor g102(.dina(n144),.dinb(w_n84_0[0]),.dout(n145),.clk(gclk));
	jor g103(.dina(w_n145_0[1]),.dinb(w_G60gat_0[1]),.dout(n146),.clk(gclk));
	jand g104(.dina(w_G329gat_5[2]),.dinb(w_n146_0[1]),.dout(n147),.clk(gclk));
	jnot g105(.din(w_n147_0[1]),.dout(n148),.clk(gclk));
	jnot g106(.din(w_G66gat_0[1]),.dout(n150),.clk(gclk));
	jand g107(.dina(w_n119_0[0]),.dinb(w_n150_0[1]),.dout(n151),.clk(gclk));
	jand g108(.dina(w_n151_0[1]),.dinb(n148),.dout(n153),.clk(gclk));
	jnot g109(.din(w_G79gat_0[1]),.dout(n154),.clk(gclk));
	jand g110(.dina(w_G223gat_2[2]),.dinb(w_G102gat_0[0]),.dout(n155),.clk(gclk));
	jor g111(.dina(n155),.dinb(w_n82_0[0]),.dout(n156),.clk(gclk));
	jor g112(.dina(w_n156_0[1]),.dinb(w_G112gat_0[1]),.dout(n157),.clk(gclk));
	jand g113(.dina(w_G223gat_2[1]),.dinb(w_G1gat_0[0]),.dout(n158),.clk(gclk));
	jor g114(.dina(n158),.dinb(w_n89_0[0]),.dout(n159),.clk(gclk));
	jor g115(.dina(w_n159_0[1]),.dinb(w_G8gat_0[1]),.dout(n160),.clk(gclk));
	jand g116(.dina(n160),.dinb(n157),.dout(n161),.clk(gclk));
	jor g117(.dina(w_n139_0[0]),.dinb(w_G99gat_0[0]),.dout(n162),.clk(gclk));
	jand g118(.dina(w_G223gat_2[0]),.dinb(w_G63gat_0[0]),.dout(n163),.clk(gclk));
	jor g119(.dina(n163),.dinb(w_n79_0[0]),.dout(n164),.clk(gclk));
	jor g120(.dina(w_n164_0[1]),.dinb(w_G73gat_0[1]),.dout(n165),.clk(gclk));
	jand g121(.dina(n165),.dinb(n162),.dout(n166),.clk(gclk));
	jand g122(.dina(n166),.dinb(n161),.dout(n167),.clk(gclk));
	jxor g123(.dina(w_n94_1[1]),.dinb(w_n78_0[0]),.dout(n168),.clk(gclk));
	jnot g124(.din(w_n123_0[0]),.dout(n169),.clk(gclk));
	jor g125(.dina(n169),.dinb(n168),.dout(n170),.clk(gclk));
	jand g126(.dina(w_n170_0[1]),.dinb(w_n146_0[0]),.dout(n171),.clk(gclk));
	jnot g127(.din(w_G82gat_0[0]),.dout(n172),.clk(gclk));
	jand g128(.dina(w_G223gat_1[2]),.dinb(w_G76gat_0[0]),.dout(n173),.clk(gclk));
	jor g129(.dina(n173),.dinb(w_dff_B_6pAiUECP2_1),.dout(n174),.clk(gclk));
	jor g130(.dina(w_n174_0[1]),.dinb(w_G86gat_1[0]),.dout(n175),.clk(gclk));
	jand g131(.dina(w_G223gat_1[1]),.dinb(w_G11gat_0[0]),.dout(n176),.clk(gclk));
	jor g132(.dina(n176),.dinb(w_n73_0[0]),.dout(n177),.clk(gclk));
	jor g133(.dina(w_n177_0[1]),.dinb(w_G21gat_1[0]),.dout(n178),.clk(gclk));
	jand g134(.dina(n178),.dinb(n175),.dout(n179),.clk(gclk));
	jand g135(.dina(n179),.dinb(n171),.dout(n180),.clk(gclk));
	jand g136(.dina(n180),.dinb(w_n115_0[0]),.dout(n181),.clk(gclk));
	jand g137(.dina(n181),.dinb(w_dff_B_30JJ7VWd1_1),.dout(n182),.clk(gclk));
	jor g138(.dina(w_n182_3[1]),.dinb(w_n107_0[0]),.dout(n183),.clk(gclk));
	jand g139(.dina(n183),.dinb(w_n109_0[0]),.dout(n184),.clk(gclk));
	jand g140(.dina(w_n184_0[1]),.dinb(w_n154_0[1]),.dout(n185),.clk(gclk));
	jor g141(.dina(n185),.dinb(n153),.dout(n186),.clk(gclk));
	jor g142(.dina(n186),.dinb(n143),.dout(n187),.clk(gclk));
	jand g143(.dina(w_G329gat_5[1]),.dinb(w_n170_0[0]),.dout(n188),.clk(gclk));
	jnot g144(.din(w_n188_0[1]),.dout(n189),.clk(gclk));
	jnot g145(.din(w_G53gat_0[1]),.dout(n191),.clk(gclk));
	jand g146(.dina(w_n191_0[1]),.dinb(w_G43gat_0[1]),.dout(n192),.clk(gclk));
	jand g147(.dina(n192),.dinb(w_n121_0[0]),.dout(n193),.clk(gclk));
	jand g148(.dina(w_n193_0[1]),.dinb(n189),.dout(n195),.clk(gclk));
	jor g149(.dina(w_n182_3[0]),.dinb(w_n130_0[1]),.dout(n196),.clk(gclk));
	jand g150(.dina(n196),.dinb(w_n132_0[0]),.dout(n197),.clk(gclk));
	jnot g151(.din(w_G27gat_0[1]),.dout(n198),.clk(gclk));
	jor g152(.dina(w_G329gat_5[0]),.dinb(w_G21gat_0[2]),.dout(n199),.clk(gclk));
	jand g153(.dina(n199),.dinb(w_n198_0[1]),.dout(n200),.clk(gclk));
	jand g154(.dina(n200),.dinb(w_n197_0[1]),.dout(n201),.clk(gclk));
	jor g155(.dina(n201),.dinb(n195),.dout(n202),.clk(gclk));
	jor g156(.dina(w_n182_2[2]),.dinb(w_n126_0[1]),.dout(n203),.clk(gclk));
	jand g157(.dina(n203),.dinb(w_n128_0[0]),.dout(n204),.clk(gclk));
	jnot g158(.din(w_G92gat_0[2]),.dout(n205),.clk(gclk));
	jor g159(.dina(w_G329gat_4[2]),.dinb(w_G86gat_0[2]),.dout(n206),.clk(gclk));
	jand g160(.dina(n206),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jand g161(.dina(n207),.dinb(w_n204_0[1]),.dout(n208),.clk(gclk));
	jnot g162(.din(w_G14gat_0[2]),.dout(n209),.clk(gclk));
	jor g163(.dina(w_n182_2[1]),.dinb(w_n98_0[0]),.dout(n210),.clk(gclk));
	jand g164(.dina(n210),.dinb(w_n100_0[0]),.dout(n211),.clk(gclk));
	jand g165(.dina(n211),.dinb(w_dff_B_9K2odaVq1_1),.dout(n212),.clk(gclk));
	jor g166(.dina(n212),.dinb(n208),.dout(n213),.clk(gclk));
	jnot g167(.din(w_G34gat_0[1]),.dout(n214),.clk(gclk));
	jor g168(.dina(w_n182_2[0]),.dinb(w_dff_B_QLbN3OC24_1),.dout(n215),.clk(gclk));
	jnot g169(.din(w_G40gat_0[1]),.dout(n217),.clk(gclk));
	jnot g170(.din(w_n114_0[1]),.dout(n218),.clk(gclk));
	jand g171(.dina(n218),.dinb(w_n217_0[1]),.dout(n219),.clk(gclk));
	jand g172(.dina(w_n219_0[1]),.dinb(n215),.dout(n221),.clk(gclk));
	jnot g173(.din(w_G115gat_0[1]),.dout(n222),.clk(gclk));
	jor g174(.dina(w_n182_1[2]),.dinb(w_n69_0[0]),.dout(n223),.clk(gclk));
	jand g175(.dina(n223),.dinb(w_n96_0[0]),.dout(n224),.clk(gclk));
	jand g176(.dina(w_n224_0[1]),.dinb(w_n222_0[1]),.dout(n225),.clk(gclk));
	jor g177(.dina(n225),.dinb(w_dff_B_ErEIblJx5_1),.dout(n226),.clk(gclk));
	jor g178(.dina(n226),.dinb(n213),.dout(n227),.clk(gclk));
	jor g179(.dina(n227),.dinb(w_dff_B_VWnVZ5F89_1),.dout(n228),.clk(gclk));
	jor g180(.dina(n228),.dinb(w_dff_B_8MFLnt5m9_1),.dout(G370gat_fa_),.clk(gclk));
	jand g181(.dina(w_G329gat_4[1]),.dinb(w_G8gat_0[0]),.dout(n230),.clk(gclk));
	jor g182(.dina(n230),.dinb(w_n159_0[0]),.dout(n231),.clk(gclk));
	jand g183(.dina(w_G370gat_2),.dinb(w_G14gat_0[1]),.dout(n232),.clk(gclk));
	jor g184(.dina(n232),.dinb(w_n231_0[1]),.dout(n233),.clk(gclk));
	jnot g185(.din(w_n151_0[0]),.dout(n235),.clk(gclk));
	jor g186(.dina(w_dff_B_rOrn4pq43_0),.dinb(w_n147_0[0]),.dout(n237),.clk(gclk));
	jand g187(.dina(w_G329gat_4[0]),.dinb(w_G73gat_0[0]),.dout(n238),.clk(gclk));
	jor g188(.dina(n238),.dinb(w_n164_0[0]),.dout(n239),.clk(gclk));
	jor g189(.dina(n239),.dinb(w_G79gat_0[0]),.dout(n240),.clk(gclk));
	jand g190(.dina(n240),.dinb(w_dff_B_PJdAhUWv3_1),.dout(n241),.clk(gclk));
	jand g191(.dina(n241),.dinb(w_n142_0[0]),.dout(n242),.clk(gclk));
	jnot g192(.din(w_n193_0[0]),.dout(n244),.clk(gclk));
	jor g193(.dina(w_dff_B_LU7xsRHL2_0),.dinb(w_n188_0[0]),.dout(n246),.clk(gclk));
	jand g194(.dina(w_G329gat_3[2]),.dinb(w_G21gat_0[1]),.dout(n247),.clk(gclk));
	jor g195(.dina(n247),.dinb(w_n177_0[0]),.dout(n248),.clk(gclk));
	jand g196(.dina(w_n182_1[1]),.dinb(w_n130_0[0]),.dout(n249),.clk(gclk));
	jor g197(.dina(n249),.dinb(w_G27gat_0[0]),.dout(n250),.clk(gclk));
	jor g198(.dina(n250),.dinb(n248),.dout(n251),.clk(gclk));
	jand g199(.dina(n251),.dinb(w_dff_B_JYpo5TJY7_1),.dout(n252),.clk(gclk));
	jand g200(.dina(w_G329gat_3[1]),.dinb(w_G86gat_0[1]),.dout(n253),.clk(gclk));
	jor g201(.dina(n253),.dinb(w_n174_0[0]),.dout(n254),.clk(gclk));
	jand g202(.dina(w_n182_1[0]),.dinb(w_n126_0[0]),.dout(n255),.clk(gclk));
	jor g203(.dina(n255),.dinb(w_G92gat_0[1]),.dout(n256),.clk(gclk));
	jor g204(.dina(n256),.dinb(w_n254_0[1]),.dout(n257),.clk(gclk));
	jor g205(.dina(w_n231_0[0]),.dinb(w_G14gat_0[0]),.dout(n258),.clk(gclk));
	jand g206(.dina(n258),.dinb(n257),.dout(n259),.clk(gclk));
	jand g207(.dina(w_G329gat_3[0]),.dinb(w_G34gat_0[0]),.dout(n260),.clk(gclk));
	jnot g208(.din(w_n219_0[0]),.dout(n262),.clk(gclk));
	jor g209(.dina(w_dff_B_cwhqTbIK1_0),.dinb(w_n260_0[1]),.dout(n264),.clk(gclk));
	jand g210(.dina(w_G329gat_2[2]),.dinb(w_G112gat_0[0]),.dout(n265),.clk(gclk));
	jor g211(.dina(n265),.dinb(w_n156_0[0]),.dout(n266),.clk(gclk));
	jor g212(.dina(n266),.dinb(w_G115gat_0[0]),.dout(n267),.clk(gclk));
	jand g213(.dina(n267),.dinb(w_dff_B_Le00bwyL1_1),.dout(n268),.clk(gclk));
	jand g214(.dina(n268),.dinb(n259),.dout(n269),.clk(gclk));
	jand g215(.dina(n269),.dinb(w_dff_B_YuoYgjBp9_1),.dout(n270),.clk(gclk));
	jand g216(.dina(n270),.dinb(w_dff_B_dXfHzVvI2_1),.dout(n271),.clk(gclk));
	jor g217(.dina(w_n271_3[1]),.dinb(w_n150_0[0]),.dout(n272),.clk(gclk));
	jand g218(.dina(w_G329gat_2[1]),.dinb(w_G60gat_0[0]),.dout(n273),.clk(gclk));
	jor g219(.dina(n273),.dinb(w_n145_0[0]),.dout(n274),.clk(gclk));
	jnot g220(.din(w_n274_0[1]),.dout(n275),.clk(gclk));
	jand g221(.dina(w_dff_B_aRJZPg1J1_0),.dinb(n272),.dout(n276),.clk(gclk));
	jor g222(.dina(w_n271_3[0]),.dinb(w_n191_0[0]),.dout(n277),.clk(gclk));
	jand g223(.dina(w_G329gat_2[0]),.dinb(w_G47gat_0[0]),.dout(n278),.clk(gclk));
	jand g224(.dina(w_G223gat_1[0]),.dinb(w_G37gat_0[0]),.dout(n279),.clk(gclk));
	jor g225(.dina(n279),.dinb(w_n77_0[0]),.dout(n280),.clk(gclk));
	jor g226(.dina(w_dff_B_GD1r0xmC1_0),.dinb(n278),.dout(n281),.clk(gclk));
	jnot g227(.din(w_n281_0[1]),.dout(n282),.clk(gclk));
	jand g228(.dina(w_dff_B_dr6xUBbA2_0),.dinb(n277),.dout(n283),.clk(gclk));
	jor g229(.dina(w_n283_0[1]),.dinb(n276),.dout(n284),.clk(gclk));
	jor g230(.dina(w_n271_2[2]),.dinb(w_n198_0[0]),.dout(n285),.clk(gclk));
	jand g231(.dina(n285),.dinb(w_n197_0[0]),.dout(n286),.clk(gclk));
	jor g232(.dina(w_n271_2[1]),.dinb(w_n217_0[0]),.dout(n287),.clk(gclk));
	jor g233(.dina(w_n114_0[0]),.dinb(w_n260_0[0]),.dout(n290),.clk(gclk));
	jnot g234(.din(w_n290_0[1]),.dout(n291),.clk(gclk));
	jand g235(.dina(w_dff_B_XsdkV8eb0_0),.dinb(n287),.dout(n292),.clk(gclk));
	jor g236(.dina(n292),.dinb(w_n286_0[1]),.dout(n293),.clk(gclk));
	jor g237(.dina(w_n293_0[1]),.dinb(n284),.dout(G430gat_fa_),.clk(gclk));
	jor g238(.dina(w_n271_2[0]),.dinb(w_n205_0[0]),.dout(n295),.clk(gclk));
	jand g239(.dina(n295),.dinb(w_n204_0[0]),.dout(n296),.clk(gclk));
	jor g240(.dina(w_n271_1[2]),.dinb(w_n222_0[0]),.dout(n297),.clk(gclk));
	jand g241(.dina(n297),.dinb(w_n224_0[0]),.dout(n298),.clk(gclk));
	jor g242(.dina(n298),.dinb(w_n296_0[1]),.dout(n299),.clk(gclk));
	jnot g243(.din(w_n141_0[0]),.dout(n300),.clk(gclk));
	jnot g244(.din(w_G105gat_0[0]),.dout(n301),.clk(gclk));
	jor g245(.dina(w_n271_1[1]),.dinb(w_dff_B_1fsV7m6g8_1),.dout(n302),.clk(gclk));
	jand g246(.dina(n302),.dinb(w_dff_B_VsfiNflG8_1),.dout(n303),.clk(gclk));
	jor g247(.dina(w_n271_1[0]),.dinb(w_n154_0[0]),.dout(n304),.clk(gclk));
	jand g248(.dina(n304),.dinb(w_n184_0[0]),.dout(n305),.clk(gclk));
	jor g249(.dina(w_n305_0[1]),.dinb(w_n303_0[1]),.dout(n306),.clk(gclk));
	jor g250(.dina(n306),.dinb(n299),.dout(n307),.clk(gclk));
	jor g251(.dina(n307),.dinb(w_G430gat_0),.dout(n308),.clk(gclk));
	jand g252(.dina(n308),.dinb(w_dff_B_rtAp55pV5_1),.dout(G421gat),.clk(gclk));
	jand g253(.dina(w_G370gat_1[2]),.dinb(w_G66gat_0[0]),.dout(n310),.clk(gclk));
	jor g254(.dina(w_n274_0[0]),.dinb(n310),.dout(n311),.clk(gclk));
	jand g255(.dina(w_G370gat_1[1]),.dinb(w_G53gat_0[0]),.dout(n312),.clk(gclk));
	jor g256(.dina(w_n281_0[0]),.dinb(n312),.dout(n313),.clk(gclk));
	jand g257(.dina(w_n313_0[1]),.dinb(n311),.dout(n314),.clk(gclk));
	jand g258(.dina(w_n296_0[0]),.dinb(w_n314_0[1]),.dout(n315),.clk(gclk));
	jand g259(.dina(w_G370gat_1[0]),.dinb(w_G40gat_0[0]),.dout(n316),.clk(gclk));
	jor g260(.dina(w_n290_0[0]),.dinb(n316),.dout(n317),.clk(gclk));
	jand g261(.dina(w_n305_0[0]),.dinb(w_n317_0[2]),.dout(n318),.clk(gclk));
	jand g262(.dina(n318),.dinb(w_n314_0[0]),.dout(n319),.clk(gclk));
	jor g263(.dina(w_n319_0[1]),.dinb(w_n293_0[0]),.dout(n320),.clk(gclk));
	jor g264(.dina(n320),.dinb(w_dff_B_iDU98mng5_1),.dout(G431gat),.clk(gclk));
	jand g265(.dina(w_G370gat_0[2]),.dinb(w_G92gat_0[0]),.dout(n322),.clk(gclk));
	jor g266(.dina(n322),.dinb(w_n254_0[0]),.dout(n323),.clk(gclk));
	jand g267(.dina(n323),.dinb(w_n313_0[0]),.dout(n324),.clk(gclk));
	jand g268(.dina(w_n303_0[0]),.dinb(w_n317_0[1]),.dout(n325),.clk(gclk));
	jand g269(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jand g270(.dina(w_n317_0[0]),.dinb(w_n283_0[0]),.dout(n327),.clk(gclk));
	jor g271(.dina(n327),.dinb(w_n286_0[0]),.dout(n328),.clk(gclk));
	jor g272(.dina(n328),.dinb(w_n319_0[0]),.dout(n329),.clk(gclk));
	jor g273(.dina(n329),.dinb(w_dff_B_Cy7OM6LL8_1),.dout(G432gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_G4gat_0[0]),.doutb(w_G4gat_0[1]),.doutc(w_G4gat_0[2]),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G11gat_0(.douta(w_G11gat_0[0]),.doutb(w_G11gat_0[1]),.doutc(w_G11gat_0[2]),.din(G11gat));
	jspl3 jspl3_w_G14gat_0(.douta(w_G14gat_0[0]),.doutb(w_G14gat_0[1]),.doutc(w_G14gat_0[2]),.din(G14gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_G21gat_0[0]),.doutb(w_G21gat_0[1]),.doutc(w_G21gat_0[2]),.din(G21gat));
	jspl jspl_w_G21gat_1(.douta(w_G21gat_1[0]),.doutb(w_G21gat_1[1]),.din(w_G21gat_0[0]));
	jspl jspl_w_G24gat_0(.douta(w_G24gat_0[0]),.doutb(w_G24gat_0[1]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_G27gat_0[0]),.doutb(w_G27gat_0[1]),.din(G27gat));
	jspl jspl_w_G30gat_0(.douta(w_G30gat_0[0]),.doutb(w_G30gat_0[1]),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_G34gat_0[0]),.doutb(w_G34gat_0[1]),.doutc(w_G34gat_0[2]),.din(G34gat));
	jspl3 jspl3_w_G37gat_0(.douta(w_G37gat_0[0]),.doutb(w_G37gat_0[1]),.doutc(w_G37gat_0[2]),.din(G37gat));
	jspl jspl_w_G40gat_0(.douta(w_G40gat_0[0]),.doutb(w_G40gat_0[1]),.din(G40gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_G43gat_0[0]),.doutb(w_G43gat_0[1]),.doutc(w_G43gat_0[2]),.din(G43gat));
	jspl jspl_w_G43gat_1(.douta(w_G43gat_1[0]),.doutb(w_G43gat_1[1]),.din(w_G43gat_0[0]));
	jspl jspl_w_G47gat_0(.douta(w_G47gat_0[0]),.doutb(w_G47gat_0[1]),.din(G47gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_G50gat_0[0]),.doutb(w_G50gat_0[1]),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_G53gat_0[0]),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_G56gat_0[0]),.doutb(w_G56gat_0[1]),.doutc(w_G56gat_0[2]),.din(G56gat));
	jspl3 jspl3_w_G60gat_0(.douta(w_G60gat_0[0]),.doutb(w_G60gat_0[1]),.doutc(w_G60gat_0[2]),.din(G60gat));
	jspl3 jspl3_w_G63gat_0(.douta(w_G63gat_0[0]),.doutb(w_G63gat_0[1]),.doutc(w_G63gat_0[2]),.din(G63gat));
	jspl jspl_w_G66gat_0(.douta(w_G66gat_0[0]),.doutb(w_G66gat_0[1]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G73gat_0(.douta(w_G73gat_0[0]),.doutb(w_G73gat_0[1]),.doutc(w_G73gat_0[2]),.din(G73gat));
	jspl jspl_w_G76gat_0(.douta(w_G76gat_0[0]),.doutb(w_G76gat_0[1]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_G79gat_0[0]),.doutb(w_G79gat_0[1]),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_G82gat_0[0]),.doutb(w_G82gat_0[1]),.doutc(w_G82gat_0[2]),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl jspl_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G89gat_0(.douta(w_G89gat_0[0]),.doutb(w_G89gat_0[1]),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_G92gat_0[0]),.doutb(w_G92gat_0[1]),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_G95gat_0[0]),.doutb(w_G95gat_0[1]),.doutc(w_G95gat_0[2]),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_G99gat_0[0]),.doutb(w_G99gat_0[1]),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl3 jspl3_w_G102gat_0(.douta(w_G102gat_0[0]),.doutb(w_G102gat_0[1]),.doutc(w_G102gat_0[2]),.din(G102gat));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_G105gat_0[1]),.din(G105gat));
	jspl3 jspl3_w_G108gat_0(.douta(w_G108gat_0[0]),.doutb(w_G108gat_0[1]),.doutc(w_G108gat_0[2]),.din(G108gat));
	jspl3 jspl3_w_G112gat_0(.douta(w_G112gat_0[0]),.doutb(w_G112gat_0[1]),.doutc(w_G112gat_0[2]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_G115gat_0[0]),.doutb(w_G115gat_0[1]),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(w_dff_A_U2myqVlw1_2),.din(w_G223gat_0[2]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl3 jspl3_w_G329gat_4(.douta(w_G329gat_4[0]),.doutb(w_G329gat_4[1]),.doutc(w_G329gat_4[2]),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G329gat_5(.douta(w_G329gat_5[0]),.doutb(w_G329gat_5[1]),.doutc(w_G329gat_5[2]),.din(w_G329gat_1[1]));
	jspl jspl_w_G329gat_6(.douta(w_G329gat_6),.doutb(w_dff_A_6BlOj4PO6_1),.din(w_G329gat_1[2]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_G370gat_1[2]),.din(w_G370gat_0[0]));
	jspl jspl_w_G370gat_2(.douta(w_G370gat_2),.doutb(w_dff_A_iURVVgb10_1),.din(w_G370gat_0[1]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(w_dff_A_C8M0FakO9_1),.din(G430gat_fa_));
	jspl jspl_w_n43_0(.douta(w_n43_0[0]),.doutb(w_n43_0[1]),.din(n43));
	jspl jspl_w_n44_0(.douta(w_n44_0[0]),.doutb(w_n44_0[1]),.din(n44));
	jspl jspl_w_n47_0(.douta(w_n47_0[0]),.doutb(w_n47_0[1]),.din(n47));
	jspl jspl_w_n52_0(.douta(w_n52_0[0]),.doutb(w_n52_0[1]),.din(n52));
	jspl jspl_w_n53_0(.douta(w_n53_0[0]),.doutb(w_n53_0[1]),.din(n53));
	jspl jspl_w_n56_0(.douta(w_n56_0[0]),.doutb(w_n56_0[1]),.din(n56));
	jspl jspl_w_n58_0(.douta(w_n58_0[0]),.doutb(w_n58_0[1]),.din(n58));
	jspl jspl_w_n61_0(.douta(w_n61_0[0]),.doutb(w_n61_0[1]),.din(n61));
	jspl jspl_w_n63_0(.douta(w_n63_0[0]),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n69_0(.douta(w_n69_0[0]),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n72_0(.douta(w_n72_0[0]),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.din(n79));
	jspl jspl_w_n82_0(.douta(w_n82_0[0]),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n87_0(.douta(w_n87_0[0]),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_n89_0[0]),.doutb(w_n89_0[1]),.din(n89));
	jspl3 jspl3_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl3 jspl3_w_n94_1(.douta(w_n94_1[0]),.doutb(w_n94_1[1]),.doutc(w_n94_1[2]),.din(w_n94_0[0]));
	jspl3 jspl3_w_n94_2(.douta(w_n94_2[0]),.doutb(w_n94_2[1]),.doutc(w_n94_2[2]),.din(w_n94_0[1]));
	jspl3 jspl3_w_n94_3(.douta(w_n94_3[0]),.doutb(w_n94_3[1]),.doutc(w_n94_3[2]),.din(w_n94_0[2]));
	jspl jspl_w_n94_4(.douta(w_n94_4[0]),.doutb(w_n94_4[1]),.din(w_n94_1[0]));
	jspl jspl_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n100_0(.douta(w_n100_0[0]),.doutb(w_n100_0[1]),.din(n100));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n114_0(.douta(w_n114_0[0]),.doutb(w_n114_0[1]),.doutc(w_n114_0[2]),.din(n114));
	jspl jspl_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.din(n115));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.din(n123));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(n128));
	jspl3 jspl3_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.doutc(w_n130_0[2]),.din(n130));
	jspl jspl_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.din(n132));
	jspl jspl_w_n139_0(.douta(w_n139_0[0]),.doutb(w_dff_A_4wpWuhcS5_1),.din(n139));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_dff_A_HeeEoTy64_0),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n145_0(.douta(w_dff_A_HK2fndwt2_0),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_iDTa47vb4_1),.din(n146));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl jspl_w_n150_0(.douta(w_n150_0[0]),.doutb(w_n150_0[1]),.din(n150));
	jspl jspl_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.din(n151));
	jspl jspl_w_n154_0(.douta(w_dff_A_KANBbx909_0),.doutb(w_n154_0[1]),.din(w_dff_B_R2JwCoqq6_2));
	jspl jspl_w_n156_0(.douta(w_dff_A_CZVKhSoJ6_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n159_0(.douta(w_dff_A_SXewAdwv0_0),.doutb(w_n159_0[1]),.din(n159));
	jspl jspl_w_n164_0(.douta(w_dff_A_H9jgYljp9_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n170_0(.douta(w_dff_A_y5ZGbqtw9_0),.doutb(w_n170_0[1]),.din(w_dff_B_5Z31j0s29_2));
	jspl jspl_w_n174_0(.douta(w_dff_A_RISmnG7W4_0),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n177_0(.douta(w_dff_A_GeqVoK4M6_0),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n182_2(.douta(w_n182_2[0]),.doutb(w_n182_2[1]),.doutc(w_n182_2[2]),.din(w_n182_0[1]));
	jspl jspl_w_n182_3(.douta(w_n182_3[0]),.doutb(w_n182_3[1]),.din(w_n182_0[2]));
	jspl jspl_w_n184_0(.douta(w_dff_A_0jaXmlQm8_0),.doutb(w_n184_0[1]),.din(n184));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.din(n191));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.din(n193));
	jspl jspl_w_n197_0(.douta(w_dff_A_FVGC99NZ8_0),.doutb(w_n197_0[1]),.din(n197));
	jspl jspl_w_n198_0(.douta(w_dff_A_r64e4DY39_0),.doutb(w_n198_0[1]),.din(w_dff_B_dCAN8GhJ7_2));
	jspl jspl_w_n204_0(.douta(w_dff_A_0CZK0CXH3_0),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n205_0(.douta(w_dff_A_aR5lBUSR9_0),.doutb(w_n205_0[1]),.din(w_dff_B_4HksJLIe0_2));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n222_0(.douta(w_dff_A_CYPpKWXV4_0),.doutb(w_n222_0[1]),.din(w_dff_B_tiu2edyZ9_2));
	jspl jspl_w_n224_0(.douta(w_dff_A_HQnMQAMg9_0),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_dff_A_401m6pOU5_1),.din(n231));
	jspl jspl_w_n254_0(.douta(w_dff_A_RDuB9J604_0),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_n271_1[0]),.doutb(w_n271_1[1]),.doutc(w_n271_1[2]),.din(w_n271_0[0]));
	jspl3 jspl3_w_n271_2(.douta(w_n271_2[0]),.doutb(w_n271_2[1]),.doutc(w_n271_2[2]),.din(w_n271_0[1]));
	jspl jspl_w_n271_3(.douta(w_n271_3[0]),.doutb(w_n271_3[1]),.din(w_n271_0[2]));
	jspl jspl_w_n274_0(.douta(w_dff_A_w4LmiAQl5_0),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n281_0(.douta(w_dff_A_elp8uBYG5_0),.doutb(w_n281_0[1]),.din(n281));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.din(n283));
	jspl jspl_w_n286_0(.douta(w_dff_A_ZCGVbZ6j3_0),.doutb(w_n286_0[1]),.din(n286));
	jspl jspl_w_n290_0(.douta(w_dff_A_Io8wu6CR0_0),.doutb(w_n290_0[1]),.din(n290));
	jspl jspl_w_n293_0(.douta(w_dff_A_WEGfJ7D77_0),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n296_0(.douta(w_dff_A_CPVisDct8_0),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(n305));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.din(n314));
	jspl3 jspl3_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.doutc(w_n317_0[2]),.din(n317));
	jspl jspl_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.din(n319));
	jdff dff_B_XtHeAfHt3_1(.din(n233),.dout(w_dff_B_XtHeAfHt3_1),.clk(gclk));
	jdff dff_B_mU4a1R0G9_1(.din(w_dff_B_XtHeAfHt3_1),.dout(w_dff_B_mU4a1R0G9_1),.clk(gclk));
	jdff dff_B_rtAp55pV5_1(.din(w_dff_B_mU4a1R0G9_1),.dout(w_dff_B_rtAp55pV5_1),.clk(gclk));
	jdff dff_B_zXWR4QiJ6_0(.din(n275),.dout(w_dff_B_zXWR4QiJ6_0),.clk(gclk));
	jdff dff_B_nHXfgPoY1_0(.din(w_dff_B_zXWR4QiJ6_0),.dout(w_dff_B_nHXfgPoY1_0),.clk(gclk));
	jdff dff_B_bNEI4rL86_0(.din(w_dff_B_nHXfgPoY1_0),.dout(w_dff_B_bNEI4rL86_0),.clk(gclk));
	jdff dff_B_IMDGVjcC1_0(.din(w_dff_B_bNEI4rL86_0),.dout(w_dff_B_IMDGVjcC1_0),.clk(gclk));
	jdff dff_B_aRJZPg1J1_0(.din(w_dff_B_IMDGVjcC1_0),.dout(w_dff_B_aRJZPg1J1_0),.clk(gclk));
	jdff dff_B_iDU98mng5_1(.din(n315),.dout(w_dff_B_iDU98mng5_1),.clk(gclk));
	jdff dff_A_WEGfJ7D77_0(.dout(w_n293_0[0]),.din(w_dff_A_WEGfJ7D77_0),.clk(gclk));
	jdff dff_B_2fu6BJoY9_0(.din(n291),.dout(w_dff_B_2fu6BJoY9_0),.clk(gclk));
	jdff dff_B_yGPvgfJt3_0(.din(w_dff_B_2fu6BJoY9_0),.dout(w_dff_B_yGPvgfJt3_0),.clk(gclk));
	jdff dff_B_9Xu2oV544_0(.din(w_dff_B_yGPvgfJt3_0),.dout(w_dff_B_9Xu2oV544_0),.clk(gclk));
	jdff dff_B_nTjcGx367_0(.din(w_dff_B_9Xu2oV544_0),.dout(w_dff_B_nTjcGx367_0),.clk(gclk));
	jdff dff_B_XsdkV8eb0_0(.din(w_dff_B_nTjcGx367_0),.dout(w_dff_B_XsdkV8eb0_0),.clk(gclk));
	jdff dff_A_CPVisDct8_0(.dout(w_n296_0[0]),.din(w_dff_A_CPVisDct8_0),.clk(gclk));
	jdff dff_B_Cy7OM6LL8_1(.din(n326),.dout(w_dff_B_Cy7OM6LL8_1),.clk(gclk));
	jdff dff_B_Tz57h5cV9_0(.din(n282),.dout(w_dff_B_Tz57h5cV9_0),.clk(gclk));
	jdff dff_B_vvFGQoVh3_0(.din(w_dff_B_Tz57h5cV9_0),.dout(w_dff_B_vvFGQoVh3_0),.clk(gclk));
	jdff dff_B_LZ0A1fIT9_0(.din(w_dff_B_vvFGQoVh3_0),.dout(w_dff_B_LZ0A1fIT9_0),.clk(gclk));
	jdff dff_B_Fgsm36Nb6_0(.din(w_dff_B_LZ0A1fIT9_0),.dout(w_dff_B_Fgsm36Nb6_0),.clk(gclk));
	jdff dff_B_dr6xUBbA2_0(.din(w_dff_B_Fgsm36Nb6_0),.dout(w_dff_B_dr6xUBbA2_0),.clk(gclk));
	jdff dff_A_ZCGVbZ6j3_0(.dout(w_n286_0[0]),.din(w_dff_A_ZCGVbZ6j3_0),.clk(gclk));
	jdff dff_A_hPDd8nNh7_0(.dout(w_n274_0[0]),.din(w_dff_A_hPDd8nNh7_0),.clk(gclk));
	jdff dff_A_62pZ9gad9_0(.dout(w_dff_A_hPDd8nNh7_0),.din(w_dff_A_62pZ9gad9_0),.clk(gclk));
	jdff dff_A_LP1iDE6J0_0(.dout(w_dff_A_62pZ9gad9_0),.din(w_dff_A_LP1iDE6J0_0),.clk(gclk));
	jdff dff_A_lX0tC26d5_0(.dout(w_dff_A_LP1iDE6J0_0),.din(w_dff_A_lX0tC26d5_0),.clk(gclk));
	jdff dff_A_6NAHzLAd6_0(.dout(w_dff_A_lX0tC26d5_0),.din(w_dff_A_6NAHzLAd6_0),.clk(gclk));
	jdff dff_A_w4LmiAQl5_0(.dout(w_dff_A_6NAHzLAd6_0),.din(w_dff_A_w4LmiAQl5_0),.clk(gclk));
	jdff dff_B_5YqJoV4e2_1(.din(n300),.dout(w_dff_B_5YqJoV4e2_1),.clk(gclk));
	jdff dff_B_k5ymrU9g7_1(.din(w_dff_B_5YqJoV4e2_1),.dout(w_dff_B_k5ymrU9g7_1),.clk(gclk));
	jdff dff_B_MXFl03cr1_1(.din(w_dff_B_k5ymrU9g7_1),.dout(w_dff_B_MXFl03cr1_1),.clk(gclk));
	jdff dff_B_6vj4xBQp7_1(.din(w_dff_B_MXFl03cr1_1),.dout(w_dff_B_6vj4xBQp7_1),.clk(gclk));
	jdff dff_B_VsfiNflG8_1(.din(w_dff_B_6vj4xBQp7_1),.dout(w_dff_B_VsfiNflG8_1),.clk(gclk));
	jdff dff_B_SLaXVEXg4_1(.din(n301),.dout(w_dff_B_SLaXVEXg4_1),.clk(gclk));
	jdff dff_B_a73vCTRQ3_1(.din(w_dff_B_SLaXVEXg4_1),.dout(w_dff_B_a73vCTRQ3_1),.clk(gclk));
	jdff dff_B_H0wA1PPA9_1(.din(w_dff_B_a73vCTRQ3_1),.dout(w_dff_B_H0wA1PPA9_1),.clk(gclk));
	jdff dff_B_y6aSXzkD7_1(.din(w_dff_B_H0wA1PPA9_1),.dout(w_dff_B_y6aSXzkD7_1),.clk(gclk));
	jdff dff_B_CH96FsCJ4_1(.din(w_dff_B_y6aSXzkD7_1),.dout(w_dff_B_CH96FsCJ4_1),.clk(gclk));
	jdff dff_B_VbQXb5dF0_1(.din(w_dff_B_CH96FsCJ4_1),.dout(w_dff_B_VbQXb5dF0_1),.clk(gclk));
	jdff dff_B_AVqRZJd08_1(.din(w_dff_B_VbQXb5dF0_1),.dout(w_dff_B_AVqRZJd08_1),.clk(gclk));
	jdff dff_B_CHTtVXaK8_1(.din(w_dff_B_AVqRZJd08_1),.dout(w_dff_B_CHTtVXaK8_1),.clk(gclk));
	jdff dff_B_Vvdh6JPd3_1(.din(w_dff_B_CHTtVXaK8_1),.dout(w_dff_B_Vvdh6JPd3_1),.clk(gclk));
	jdff dff_B_9t1Ri9rA7_1(.din(w_dff_B_Vvdh6JPd3_1),.dout(w_dff_B_9t1Ri9rA7_1),.clk(gclk));
	jdff dff_B_29msO7Ij6_1(.din(w_dff_B_9t1Ri9rA7_1),.dout(w_dff_B_29msO7Ij6_1),.clk(gclk));
	jdff dff_B_TP2ysv185_1(.din(w_dff_B_29msO7Ij6_1),.dout(w_dff_B_TP2ysv185_1),.clk(gclk));
	jdff dff_B_kOZLYA213_1(.din(w_dff_B_TP2ysv185_1),.dout(w_dff_B_kOZLYA213_1),.clk(gclk));
	jdff dff_B_4CizjBJQ7_1(.din(w_dff_B_kOZLYA213_1),.dout(w_dff_B_4CizjBJQ7_1),.clk(gclk));
	jdff dff_B_7d2hg9nE5_1(.din(w_dff_B_4CizjBJQ7_1),.dout(w_dff_B_7d2hg9nE5_1),.clk(gclk));
	jdff dff_B_t64QZ5Sx5_1(.din(w_dff_B_7d2hg9nE5_1),.dout(w_dff_B_t64QZ5Sx5_1),.clk(gclk));
	jdff dff_B_stNHmWmI6_1(.din(w_dff_B_t64QZ5Sx5_1),.dout(w_dff_B_stNHmWmI6_1),.clk(gclk));
	jdff dff_B_ElDv60aw7_1(.din(w_dff_B_stNHmWmI6_1),.dout(w_dff_B_ElDv60aw7_1),.clk(gclk));
	jdff dff_B_1fsV7m6g8_1(.din(w_dff_B_ElDv60aw7_1),.dout(w_dff_B_1fsV7m6g8_1),.clk(gclk));
	jdff dff_B_dXfHzVvI2_1(.din(n242),.dout(w_dff_B_dXfHzVvI2_1),.clk(gclk));
	jdff dff_B_YuoYgjBp9_1(.din(n252),.dout(w_dff_B_YuoYgjBp9_1),.clk(gclk));
	jdff dff_B_Le00bwyL1_1(.din(n264),.dout(w_dff_B_Le00bwyL1_1),.clk(gclk));
	jdff dff_B_FissYN5J5_0(.din(n262),.dout(w_dff_B_FissYN5J5_0),.clk(gclk));
	jdff dff_B_9gYMrj778_0(.din(w_dff_B_FissYN5J5_0),.dout(w_dff_B_9gYMrj778_0),.clk(gclk));
	jdff dff_B_cwhqTbIK1_0(.din(w_dff_B_9gYMrj778_0),.dout(w_dff_B_cwhqTbIK1_0),.clk(gclk));
	jdff dff_A_uSygbgaG4_1(.dout(w_n231_0[1]),.din(w_dff_A_uSygbgaG4_1),.clk(gclk));
	jdff dff_A_lX7HOrsH8_1(.dout(w_dff_A_uSygbgaG4_1),.din(w_dff_A_lX7HOrsH8_1),.clk(gclk));
	jdff dff_A_UIBVQYQS0_1(.dout(w_dff_A_lX7HOrsH8_1),.din(w_dff_A_UIBVQYQS0_1),.clk(gclk));
	jdff dff_A_QGG2jtbD0_1(.dout(w_dff_A_UIBVQYQS0_1),.din(w_dff_A_QGG2jtbD0_1),.clk(gclk));
	jdff dff_A_PSVXGahE5_1(.dout(w_dff_A_QGG2jtbD0_1),.din(w_dff_A_PSVXGahE5_1),.clk(gclk));
	jdff dff_A_401m6pOU5_1(.dout(w_dff_A_PSVXGahE5_1),.din(w_dff_A_401m6pOU5_1),.clk(gclk));
	jdff dff_B_JYpo5TJY7_1(.din(n246),.dout(w_dff_B_JYpo5TJY7_1),.clk(gclk));
	jdff dff_B_WNoS3vJn2_0(.din(n244),.dout(w_dff_B_WNoS3vJn2_0),.clk(gclk));
	jdff dff_B_xXpzcbdI5_0(.din(w_dff_B_WNoS3vJn2_0),.dout(w_dff_B_xXpzcbdI5_0),.clk(gclk));
	jdff dff_B_5pVV6fYM3_0(.din(w_dff_B_xXpzcbdI5_0),.dout(w_dff_B_5pVV6fYM3_0),.clk(gclk));
	jdff dff_B_nwK4xXoc8_0(.din(w_dff_B_5pVV6fYM3_0),.dout(w_dff_B_nwK4xXoc8_0),.clk(gclk));
	jdff dff_B_LU7xsRHL2_0(.din(w_dff_B_nwK4xXoc8_0),.dout(w_dff_B_LU7xsRHL2_0),.clk(gclk));
	jdff dff_B_PJdAhUWv3_1(.din(n237),.dout(w_dff_B_PJdAhUWv3_1),.clk(gclk));
	jdff dff_B_N0MoOT9q2_0(.din(n235),.dout(w_dff_B_N0MoOT9q2_0),.clk(gclk));
	jdff dff_B_Wmb5Vblx7_0(.din(w_dff_B_N0MoOT9q2_0),.dout(w_dff_B_Wmb5Vblx7_0),.clk(gclk));
	jdff dff_B_1tvf18FW4_0(.din(w_dff_B_Wmb5Vblx7_0),.dout(w_dff_B_1tvf18FW4_0),.clk(gclk));
	jdff dff_B_rOrn4pq43_0(.din(w_dff_B_1tvf18FW4_0),.dout(w_dff_B_rOrn4pq43_0),.clk(gclk));
	jdff dff_A_fy0OtTh78_0(.dout(w_n290_0[0]),.din(w_dff_A_fy0OtTh78_0),.clk(gclk));
	jdff dff_A_06P2op1q6_0(.dout(w_dff_A_fy0OtTh78_0),.din(w_dff_A_06P2op1q6_0),.clk(gclk));
	jdff dff_A_Auye3inr6_0(.dout(w_dff_A_06P2op1q6_0),.din(w_dff_A_Auye3inr6_0),.clk(gclk));
	jdff dff_A_VfJ30puZ9_0(.dout(w_dff_A_Auye3inr6_0),.din(w_dff_A_VfJ30puZ9_0),.clk(gclk));
	jdff dff_A_ZtLsp5To9_0(.dout(w_dff_A_VfJ30puZ9_0),.din(w_dff_A_ZtLsp5To9_0),.clk(gclk));
	jdff dff_A_Io8wu6CR0_0(.dout(w_dff_A_ZtLsp5To9_0),.din(w_dff_A_Io8wu6CR0_0),.clk(gclk));
	jdff dff_A_mDAUDbsT8_0(.dout(w_n254_0[0]),.din(w_dff_A_mDAUDbsT8_0),.clk(gclk));
	jdff dff_A_dmfuDBAc4_0(.dout(w_dff_A_mDAUDbsT8_0),.din(w_dff_A_dmfuDBAc4_0),.clk(gclk));
	jdff dff_A_fakqwGEj0_0(.dout(w_dff_A_dmfuDBAc4_0),.din(w_dff_A_fakqwGEj0_0),.clk(gclk));
	jdff dff_A_qMYvcXrW2_0(.dout(w_dff_A_fakqwGEj0_0),.din(w_dff_A_qMYvcXrW2_0),.clk(gclk));
	jdff dff_A_lHtqvvXo0_0(.dout(w_dff_A_qMYvcXrW2_0),.din(w_dff_A_lHtqvvXo0_0),.clk(gclk));
	jdff dff_A_RDuB9J604_0(.dout(w_dff_A_lHtqvvXo0_0),.din(w_dff_A_RDuB9J604_0),.clk(gclk));
	jdff dff_A_KiXnnO0H1_0(.dout(w_n281_0[0]),.din(w_dff_A_KiXnnO0H1_0),.clk(gclk));
	jdff dff_A_rRNuASCT2_0(.dout(w_dff_A_KiXnnO0H1_0),.din(w_dff_A_rRNuASCT2_0),.clk(gclk));
	jdff dff_A_k3ABFhLk2_0(.dout(w_dff_A_rRNuASCT2_0),.din(w_dff_A_k3ABFhLk2_0),.clk(gclk));
	jdff dff_A_TWJ76dEY2_0(.dout(w_dff_A_k3ABFhLk2_0),.din(w_dff_A_TWJ76dEY2_0),.clk(gclk));
	jdff dff_A_EOkWvfXL5_0(.dout(w_dff_A_TWJ76dEY2_0),.din(w_dff_A_EOkWvfXL5_0),.clk(gclk));
	jdff dff_A_elp8uBYG5_0(.dout(w_dff_A_EOkWvfXL5_0),.din(w_dff_A_elp8uBYG5_0),.clk(gclk));
	jdff dff_B_0pQmMgYh3_0(.din(n280),.dout(w_dff_B_0pQmMgYh3_0),.clk(gclk));
	jdff dff_B_Ei3srVPx3_0(.din(w_dff_B_0pQmMgYh3_0),.dout(w_dff_B_Ei3srVPx3_0),.clk(gclk));
	jdff dff_B_FfSBo8dk2_0(.din(w_dff_B_Ei3srVPx3_0),.dout(w_dff_B_FfSBo8dk2_0),.clk(gclk));
	jdff dff_B_3GouIE3F3_0(.din(w_dff_B_FfSBo8dk2_0),.dout(w_dff_B_3GouIE3F3_0),.clk(gclk));
	jdff dff_B_zut9mmyo8_0(.din(w_dff_B_3GouIE3F3_0),.dout(w_dff_B_zut9mmyo8_0),.clk(gclk));
	jdff dff_B_GD1r0xmC1_0(.din(w_dff_B_zut9mmyo8_0),.dout(w_dff_B_GD1r0xmC1_0),.clk(gclk));
	jdff dff_B_8MFLnt5m9_1(.din(n187),.dout(w_dff_B_8MFLnt5m9_1),.clk(gclk));
	jdff dff_B_VWnVZ5F89_1(.din(n202),.dout(w_dff_B_VWnVZ5F89_1),.clk(gclk));
	jdff dff_B_ErEIblJx5_1(.din(n221),.dout(w_dff_B_ErEIblJx5_1),.clk(gclk));
	jdff dff_A_jAzNkW4y0_0(.dout(w_n224_0[0]),.din(w_dff_A_jAzNkW4y0_0),.clk(gclk));
	jdff dff_A_Z94B9Lvk9_0(.dout(w_dff_A_jAzNkW4y0_0),.din(w_dff_A_Z94B9Lvk9_0),.clk(gclk));
	jdff dff_A_hwgTDZLm7_0(.dout(w_dff_A_Z94B9Lvk9_0),.din(w_dff_A_hwgTDZLm7_0),.clk(gclk));
	jdff dff_A_xhCE7X622_0(.dout(w_dff_A_hwgTDZLm7_0),.din(w_dff_A_xhCE7X622_0),.clk(gclk));
	jdff dff_A_nkxJFDy28_0(.dout(w_dff_A_xhCE7X622_0),.din(w_dff_A_nkxJFDy28_0),.clk(gclk));
	jdff dff_A_HQnMQAMg9_0(.dout(w_dff_A_nkxJFDy28_0),.din(w_dff_A_HQnMQAMg9_0),.clk(gclk));
	jdff dff_A_Wh1RiAQx6_0(.dout(w_n222_0[0]),.din(w_dff_A_Wh1RiAQx6_0),.clk(gclk));
	jdff dff_A_UjGwj7CU3_0(.dout(w_dff_A_Wh1RiAQx6_0),.din(w_dff_A_UjGwj7CU3_0),.clk(gclk));
	jdff dff_A_ALys9RFq4_0(.dout(w_dff_A_UjGwj7CU3_0),.din(w_dff_A_ALys9RFq4_0),.clk(gclk));
	jdff dff_A_31UNmNVu2_0(.dout(w_dff_A_ALys9RFq4_0),.din(w_dff_A_31UNmNVu2_0),.clk(gclk));
	jdff dff_A_CYPpKWXV4_0(.dout(w_dff_A_31UNmNVu2_0),.din(w_dff_A_CYPpKWXV4_0),.clk(gclk));
	jdff dff_B_qg7mWGb20_2(.din(n222),.dout(w_dff_B_qg7mWGb20_2),.clk(gclk));
	jdff dff_B_MW5gfkNF4_2(.din(w_dff_B_qg7mWGb20_2),.dout(w_dff_B_MW5gfkNF4_2),.clk(gclk));
	jdff dff_B_rsVgH1GT7_2(.din(w_dff_B_MW5gfkNF4_2),.dout(w_dff_B_rsVgH1GT7_2),.clk(gclk));
	jdff dff_B_o2BQCpRe8_2(.din(w_dff_B_rsVgH1GT7_2),.dout(w_dff_B_o2BQCpRe8_2),.clk(gclk));
	jdff dff_B_Ak0plN7W2_2(.din(w_dff_B_o2BQCpRe8_2),.dout(w_dff_B_Ak0plN7W2_2),.clk(gclk));
	jdff dff_B_2qaQWBAQ4_2(.din(w_dff_B_Ak0plN7W2_2),.dout(w_dff_B_2qaQWBAQ4_2),.clk(gclk));
	jdff dff_B_yjhHwxmA9_2(.din(w_dff_B_2qaQWBAQ4_2),.dout(w_dff_B_yjhHwxmA9_2),.clk(gclk));
	jdff dff_B_fFVjhWS68_2(.din(w_dff_B_yjhHwxmA9_2),.dout(w_dff_B_fFVjhWS68_2),.clk(gclk));
	jdff dff_B_woW1UOno0_2(.din(w_dff_B_fFVjhWS68_2),.dout(w_dff_B_woW1UOno0_2),.clk(gclk));
	jdff dff_B_ivtfX5JB3_2(.din(w_dff_B_woW1UOno0_2),.dout(w_dff_B_ivtfX5JB3_2),.clk(gclk));
	jdff dff_B_Vqrr3Xeq4_2(.din(w_dff_B_ivtfX5JB3_2),.dout(w_dff_B_Vqrr3Xeq4_2),.clk(gclk));
	jdff dff_B_hfXbhLSj7_2(.din(w_dff_B_Vqrr3Xeq4_2),.dout(w_dff_B_hfXbhLSj7_2),.clk(gclk));
	jdff dff_B_TqRYiniu7_2(.din(w_dff_B_hfXbhLSj7_2),.dout(w_dff_B_TqRYiniu7_2),.clk(gclk));
	jdff dff_B_tiu2edyZ9_2(.din(w_dff_B_TqRYiniu7_2),.dout(w_dff_B_tiu2edyZ9_2),.clk(gclk));
	jdff dff_B_FyFM8Ygp2_1(.din(n214),.dout(w_dff_B_FyFM8Ygp2_1),.clk(gclk));
	jdff dff_B_eNrwTtNg3_1(.din(w_dff_B_FyFM8Ygp2_1),.dout(w_dff_B_eNrwTtNg3_1),.clk(gclk));
	jdff dff_B_yggQB6Ys8_1(.din(w_dff_B_eNrwTtNg3_1),.dout(w_dff_B_yggQB6Ys8_1),.clk(gclk));
	jdff dff_B_U0MpGuxn5_1(.din(w_dff_B_yggQB6Ys8_1),.dout(w_dff_B_U0MpGuxn5_1),.clk(gclk));
	jdff dff_B_NYlgNJl09_1(.din(w_dff_B_U0MpGuxn5_1),.dout(w_dff_B_NYlgNJl09_1),.clk(gclk));
	jdff dff_B_x5QkcuRc4_1(.din(w_dff_B_NYlgNJl09_1),.dout(w_dff_B_x5QkcuRc4_1),.clk(gclk));
	jdff dff_B_HcES8P0P0_1(.din(w_dff_B_x5QkcuRc4_1),.dout(w_dff_B_HcES8P0P0_1),.clk(gclk));
	jdff dff_B_ppmixOzB9_1(.din(w_dff_B_HcES8P0P0_1),.dout(w_dff_B_ppmixOzB9_1),.clk(gclk));
	jdff dff_B_vmiTmYiF4_1(.din(w_dff_B_ppmixOzB9_1),.dout(w_dff_B_vmiTmYiF4_1),.clk(gclk));
	jdff dff_B_OYUCZ4l41_1(.din(w_dff_B_vmiTmYiF4_1),.dout(w_dff_B_OYUCZ4l41_1),.clk(gclk));
	jdff dff_B_aHMr6rBz7_1(.din(w_dff_B_OYUCZ4l41_1),.dout(w_dff_B_aHMr6rBz7_1),.clk(gclk));
	jdff dff_B_QLbN3OC24_1(.din(w_dff_B_aHMr6rBz7_1),.dout(w_dff_B_QLbN3OC24_1),.clk(gclk));
	jdff dff_B_AM95yKvk0_1(.din(n209),.dout(w_dff_B_AM95yKvk0_1),.clk(gclk));
	jdff dff_B_CHp7zuqa4_1(.din(w_dff_B_AM95yKvk0_1),.dout(w_dff_B_CHp7zuqa4_1),.clk(gclk));
	jdff dff_B_Y2xHbUVu2_1(.din(w_dff_B_CHp7zuqa4_1),.dout(w_dff_B_Y2xHbUVu2_1),.clk(gclk));
	jdff dff_B_laHDFc1W2_1(.din(w_dff_B_Y2xHbUVu2_1),.dout(w_dff_B_laHDFc1W2_1),.clk(gclk));
	jdff dff_B_kGyIrKsw1_1(.din(w_dff_B_laHDFc1W2_1),.dout(w_dff_B_kGyIrKsw1_1),.clk(gclk));
	jdff dff_B_KgFU634u2_1(.din(w_dff_B_kGyIrKsw1_1),.dout(w_dff_B_KgFU634u2_1),.clk(gclk));
	jdff dff_B_My7Aav3g5_1(.din(w_dff_B_KgFU634u2_1),.dout(w_dff_B_My7Aav3g5_1),.clk(gclk));
	jdff dff_B_ngP0PGs45_1(.din(w_dff_B_My7Aav3g5_1),.dout(w_dff_B_ngP0PGs45_1),.clk(gclk));
	jdff dff_B_I2tvJizq0_1(.din(w_dff_B_ngP0PGs45_1),.dout(w_dff_B_I2tvJizq0_1),.clk(gclk));
	jdff dff_B_moXcOpP59_1(.din(w_dff_B_I2tvJizq0_1),.dout(w_dff_B_moXcOpP59_1),.clk(gclk));
	jdff dff_B_CxDoqWCF9_1(.din(w_dff_B_moXcOpP59_1),.dout(w_dff_B_CxDoqWCF9_1),.clk(gclk));
	jdff dff_B_bQ8DlPv90_1(.din(w_dff_B_CxDoqWCF9_1),.dout(w_dff_B_bQ8DlPv90_1),.clk(gclk));
	jdff dff_B_NKML2GtR0_1(.din(w_dff_B_bQ8DlPv90_1),.dout(w_dff_B_NKML2GtR0_1),.clk(gclk));
	jdff dff_B_9K2odaVq1_1(.din(w_dff_B_NKML2GtR0_1),.dout(w_dff_B_9K2odaVq1_1),.clk(gclk));
	jdff dff_A_zbikquwd1_0(.dout(w_n205_0[0]),.din(w_dff_A_zbikquwd1_0),.clk(gclk));
	jdff dff_A_QVn7yNck3_0(.dout(w_dff_A_zbikquwd1_0),.din(w_dff_A_QVn7yNck3_0),.clk(gclk));
	jdff dff_A_n0TYYcXN6_0(.dout(w_dff_A_QVn7yNck3_0),.din(w_dff_A_n0TYYcXN6_0),.clk(gclk));
	jdff dff_A_ECPX5BkF9_0(.dout(w_dff_A_n0TYYcXN6_0),.din(w_dff_A_ECPX5BkF9_0),.clk(gclk));
	jdff dff_A_A6r9DdmE6_0(.dout(w_dff_A_ECPX5BkF9_0),.din(w_dff_A_A6r9DdmE6_0),.clk(gclk));
	jdff dff_A_aR5lBUSR9_0(.dout(w_dff_A_A6r9DdmE6_0),.din(w_dff_A_aR5lBUSR9_0),.clk(gclk));
	jdff dff_B_EMSPp0NZ0_2(.din(n205),.dout(w_dff_B_EMSPp0NZ0_2),.clk(gclk));
	jdff dff_B_hQvT0f3E4_2(.din(w_dff_B_EMSPp0NZ0_2),.dout(w_dff_B_hQvT0f3E4_2),.clk(gclk));
	jdff dff_B_25WKhGGk9_2(.din(w_dff_B_hQvT0f3E4_2),.dout(w_dff_B_25WKhGGk9_2),.clk(gclk));
	jdff dff_B_mh33z2Yd4_2(.din(w_dff_B_25WKhGGk9_2),.dout(w_dff_B_mh33z2Yd4_2),.clk(gclk));
	jdff dff_B_uQoBKJ9X1_2(.din(w_dff_B_mh33z2Yd4_2),.dout(w_dff_B_uQoBKJ9X1_2),.clk(gclk));
	jdff dff_B_5kEo7zCX8_2(.din(w_dff_B_uQoBKJ9X1_2),.dout(w_dff_B_5kEo7zCX8_2),.clk(gclk));
	jdff dff_B_9kmsZGCh0_2(.din(w_dff_B_5kEo7zCX8_2),.dout(w_dff_B_9kmsZGCh0_2),.clk(gclk));
	jdff dff_B_pXCl8kXn9_2(.din(w_dff_B_9kmsZGCh0_2),.dout(w_dff_B_pXCl8kXn9_2),.clk(gclk));
	jdff dff_B_k24UfNbR5_2(.din(w_dff_B_pXCl8kXn9_2),.dout(w_dff_B_k24UfNbR5_2),.clk(gclk));
	jdff dff_B_izS80gCz9_2(.din(w_dff_B_k24UfNbR5_2),.dout(w_dff_B_izS80gCz9_2),.clk(gclk));
	jdff dff_B_kemnXx8M0_2(.din(w_dff_B_izS80gCz9_2),.dout(w_dff_B_kemnXx8M0_2),.clk(gclk));
	jdff dff_B_R3jnqyQA0_2(.din(w_dff_B_kemnXx8M0_2),.dout(w_dff_B_R3jnqyQA0_2),.clk(gclk));
	jdff dff_B_4HksJLIe0_2(.din(w_dff_B_R3jnqyQA0_2),.dout(w_dff_B_4HksJLIe0_2),.clk(gclk));
	jdff dff_A_uViN6cTm4_0(.dout(w_n204_0[0]),.din(w_dff_A_uViN6cTm4_0),.clk(gclk));
	jdff dff_A_nnKjElT53_0(.dout(w_dff_A_uViN6cTm4_0),.din(w_dff_A_nnKjElT53_0),.clk(gclk));
	jdff dff_A_vbNNgIQg3_0(.dout(w_dff_A_nnKjElT53_0),.din(w_dff_A_vbNNgIQg3_0),.clk(gclk));
	jdff dff_A_Ah0ngBQz4_0(.dout(w_dff_A_vbNNgIQg3_0),.din(w_dff_A_Ah0ngBQz4_0),.clk(gclk));
	jdff dff_A_Qbd9lZ5L1_0(.dout(w_dff_A_Ah0ngBQz4_0),.din(w_dff_A_Qbd9lZ5L1_0),.clk(gclk));
	jdff dff_A_0CZK0CXH3_0(.dout(w_dff_A_Qbd9lZ5L1_0),.din(w_dff_A_0CZK0CXH3_0),.clk(gclk));
	jdff dff_A_r845OfmA6_0(.dout(w_n198_0[0]),.din(w_dff_A_r845OfmA6_0),.clk(gclk));
	jdff dff_A_eCkCE2r60_0(.dout(w_dff_A_r845OfmA6_0),.din(w_dff_A_eCkCE2r60_0),.clk(gclk));
	jdff dff_A_Laa5sYIB7_0(.dout(w_dff_A_eCkCE2r60_0),.din(w_dff_A_Laa5sYIB7_0),.clk(gclk));
	jdff dff_A_360d4E9j8_0(.dout(w_dff_A_Laa5sYIB7_0),.din(w_dff_A_360d4E9j8_0),.clk(gclk));
	jdff dff_A_6lc62de52_0(.dout(w_dff_A_360d4E9j8_0),.din(w_dff_A_6lc62de52_0),.clk(gclk));
	jdff dff_A_r64e4DY39_0(.dout(w_dff_A_6lc62de52_0),.din(w_dff_A_r64e4DY39_0),.clk(gclk));
	jdff dff_B_VBOZ7g2j6_2(.din(n198),.dout(w_dff_B_VBOZ7g2j6_2),.clk(gclk));
	jdff dff_B_eV0S1xYl3_2(.din(w_dff_B_VBOZ7g2j6_2),.dout(w_dff_B_eV0S1xYl3_2),.clk(gclk));
	jdff dff_B_KPEBxuUq7_2(.din(w_dff_B_eV0S1xYl3_2),.dout(w_dff_B_KPEBxuUq7_2),.clk(gclk));
	jdff dff_B_CEDaHPVs2_2(.din(w_dff_B_KPEBxuUq7_2),.dout(w_dff_B_CEDaHPVs2_2),.clk(gclk));
	jdff dff_B_cqlO6qAm3_2(.din(w_dff_B_CEDaHPVs2_2),.dout(w_dff_B_cqlO6qAm3_2),.clk(gclk));
	jdff dff_B_ZBpyvRCx3_2(.din(w_dff_B_cqlO6qAm3_2),.dout(w_dff_B_ZBpyvRCx3_2),.clk(gclk));
	jdff dff_B_bi592kgC7_2(.din(w_dff_B_ZBpyvRCx3_2),.dout(w_dff_B_bi592kgC7_2),.clk(gclk));
	jdff dff_B_l1YZ9jLP0_2(.din(w_dff_B_bi592kgC7_2),.dout(w_dff_B_l1YZ9jLP0_2),.clk(gclk));
	jdff dff_B_uG2bxopE2_2(.din(w_dff_B_l1YZ9jLP0_2),.dout(w_dff_B_uG2bxopE2_2),.clk(gclk));
	jdff dff_B_3BRfc02z0_2(.din(w_dff_B_uG2bxopE2_2),.dout(w_dff_B_3BRfc02z0_2),.clk(gclk));
	jdff dff_B_dh96HMii8_2(.din(w_dff_B_3BRfc02z0_2),.dout(w_dff_B_dh96HMii8_2),.clk(gclk));
	jdff dff_B_yLoxZPxV0_2(.din(w_dff_B_dh96HMii8_2),.dout(w_dff_B_yLoxZPxV0_2),.clk(gclk));
	jdff dff_B_dCAN8GhJ7_2(.din(w_dff_B_yLoxZPxV0_2),.dout(w_dff_B_dCAN8GhJ7_2),.clk(gclk));
	jdff dff_A_6tWAUU271_0(.dout(w_n197_0[0]),.din(w_dff_A_6tWAUU271_0),.clk(gclk));
	jdff dff_A_6WZoJxMl3_0(.dout(w_dff_A_6tWAUU271_0),.din(w_dff_A_6WZoJxMl3_0),.clk(gclk));
	jdff dff_A_2Eqx7S8l2_0(.dout(w_dff_A_6WZoJxMl3_0),.din(w_dff_A_2Eqx7S8l2_0),.clk(gclk));
	jdff dff_A_PYtGB0pE4_0(.dout(w_dff_A_2Eqx7S8l2_0),.din(w_dff_A_PYtGB0pE4_0),.clk(gclk));
	jdff dff_A_pVQUDdVA1_0(.dout(w_dff_A_PYtGB0pE4_0),.din(w_dff_A_pVQUDdVA1_0),.clk(gclk));
	jdff dff_A_FVGC99NZ8_0(.dout(w_dff_A_pVQUDdVA1_0),.din(w_dff_A_FVGC99NZ8_0),.clk(gclk));
	jdff dff_A_4TF5M3ij0_0(.dout(w_n184_0[0]),.din(w_dff_A_4TF5M3ij0_0),.clk(gclk));
	jdff dff_A_7kQZIIpO5_0(.dout(w_dff_A_4TF5M3ij0_0),.din(w_dff_A_7kQZIIpO5_0),.clk(gclk));
	jdff dff_A_K3LifHUO9_0(.dout(w_dff_A_7kQZIIpO5_0),.din(w_dff_A_K3LifHUO9_0),.clk(gclk));
	jdff dff_A_1bHFImJt9_0(.dout(w_dff_A_K3LifHUO9_0),.din(w_dff_A_1bHFImJt9_0),.clk(gclk));
	jdff dff_A_JQPDQPyt7_0(.dout(w_dff_A_1bHFImJt9_0),.din(w_dff_A_JQPDQPyt7_0),.clk(gclk));
	jdff dff_A_0jaXmlQm8_0(.dout(w_dff_A_JQPDQPyt7_0),.din(w_dff_A_0jaXmlQm8_0),.clk(gclk));
	jdff dff_B_30JJ7VWd1_1(.din(n167),.dout(w_dff_B_30JJ7VWd1_1),.clk(gclk));
	jdff dff_A_0Kr7sAnf0_0(.dout(w_n177_0[0]),.din(w_dff_A_0Kr7sAnf0_0),.clk(gclk));
	jdff dff_A_3FKVdAia8_0(.dout(w_dff_A_0Kr7sAnf0_0),.din(w_dff_A_3FKVdAia8_0),.clk(gclk));
	jdff dff_A_6dUHppkX9_0(.dout(w_dff_A_3FKVdAia8_0),.din(w_dff_A_6dUHppkX9_0),.clk(gclk));
	jdff dff_A_caFBgMjP5_0(.dout(w_dff_A_6dUHppkX9_0),.din(w_dff_A_caFBgMjP5_0),.clk(gclk));
	jdff dff_A_Cg9vU7Wc4_0(.dout(w_dff_A_caFBgMjP5_0),.din(w_dff_A_Cg9vU7Wc4_0),.clk(gclk));
	jdff dff_A_GeqVoK4M6_0(.dout(w_dff_A_Cg9vU7Wc4_0),.din(w_dff_A_GeqVoK4M6_0),.clk(gclk));
	jdff dff_A_hTuuCm4F8_0(.dout(w_n174_0[0]),.din(w_dff_A_hTuuCm4F8_0),.clk(gclk));
	jdff dff_A_s5PcXhe91_0(.dout(w_dff_A_hTuuCm4F8_0),.din(w_dff_A_s5PcXhe91_0),.clk(gclk));
	jdff dff_A_Zd29BN252_0(.dout(w_dff_A_s5PcXhe91_0),.din(w_dff_A_Zd29BN252_0),.clk(gclk));
	jdff dff_A_2sWQGN515_0(.dout(w_dff_A_Zd29BN252_0),.din(w_dff_A_2sWQGN515_0),.clk(gclk));
	jdff dff_A_OJmXFrQB0_0(.dout(w_dff_A_2sWQGN515_0),.din(w_dff_A_OJmXFrQB0_0),.clk(gclk));
	jdff dff_A_RISmnG7W4_0(.dout(w_dff_A_OJmXFrQB0_0),.din(w_dff_A_RISmnG7W4_0),.clk(gclk));
	jdff dff_B_sda6iCdK6_1(.din(n172),.dout(w_dff_B_sda6iCdK6_1),.clk(gclk));
	jdff dff_B_8UbO43Uq1_1(.din(w_dff_B_sda6iCdK6_1),.dout(w_dff_B_8UbO43Uq1_1),.clk(gclk));
	jdff dff_B_KDKRnPY56_1(.din(w_dff_B_8UbO43Uq1_1),.dout(w_dff_B_KDKRnPY56_1),.clk(gclk));
	jdff dff_B_bLrzaVhU1_1(.din(w_dff_B_KDKRnPY56_1),.dout(w_dff_B_bLrzaVhU1_1),.clk(gclk));
	jdff dff_B_yRRxXC9F0_1(.din(w_dff_B_bLrzaVhU1_1),.dout(w_dff_B_yRRxXC9F0_1),.clk(gclk));
	jdff dff_B_6pAiUECP2_1(.din(w_dff_B_yRRxXC9F0_1),.dout(w_dff_B_6pAiUECP2_1),.clk(gclk));
	jdff dff_A_uOjPQsTM7_0(.dout(w_n170_0[0]),.din(w_dff_A_uOjPQsTM7_0),.clk(gclk));
	jdff dff_A_FhGZDlhD1_0(.dout(w_dff_A_uOjPQsTM7_0),.din(w_dff_A_FhGZDlhD1_0),.clk(gclk));
	jdff dff_A_Sz5H8gib4_0(.dout(w_dff_A_FhGZDlhD1_0),.din(w_dff_A_Sz5H8gib4_0),.clk(gclk));
	jdff dff_A_y5ZGbqtw9_0(.dout(w_dff_A_Sz5H8gib4_0),.din(w_dff_A_y5ZGbqtw9_0),.clk(gclk));
	jdff dff_B_5Z31j0s29_2(.din(n170),.dout(w_dff_B_5Z31j0s29_2),.clk(gclk));
	jdff dff_A_qRBfRAPu7_0(.dout(w_n164_0[0]),.din(w_dff_A_qRBfRAPu7_0),.clk(gclk));
	jdff dff_A_PefwWC5e3_0(.dout(w_dff_A_qRBfRAPu7_0),.din(w_dff_A_PefwWC5e3_0),.clk(gclk));
	jdff dff_A_Py2NcyGQ4_0(.dout(w_dff_A_PefwWC5e3_0),.din(w_dff_A_Py2NcyGQ4_0),.clk(gclk));
	jdff dff_A_g0hdhvdd4_0(.dout(w_dff_A_Py2NcyGQ4_0),.din(w_dff_A_g0hdhvdd4_0),.clk(gclk));
	jdff dff_A_PuumVz3v9_0(.dout(w_dff_A_g0hdhvdd4_0),.din(w_dff_A_PuumVz3v9_0),.clk(gclk));
	jdff dff_A_H9jgYljp9_0(.dout(w_dff_A_PuumVz3v9_0),.din(w_dff_A_H9jgYljp9_0),.clk(gclk));
	jdff dff_A_FbOkL3oh9_0(.dout(w_n159_0[0]),.din(w_dff_A_FbOkL3oh9_0),.clk(gclk));
	jdff dff_A_LB8qNsp02_0(.dout(w_dff_A_FbOkL3oh9_0),.din(w_dff_A_LB8qNsp02_0),.clk(gclk));
	jdff dff_A_N6GA9OXz6_0(.dout(w_dff_A_LB8qNsp02_0),.din(w_dff_A_N6GA9OXz6_0),.clk(gclk));
	jdff dff_A_7jkH8cLA8_0(.dout(w_dff_A_N6GA9OXz6_0),.din(w_dff_A_7jkH8cLA8_0),.clk(gclk));
	jdff dff_A_yDCvhztt5_0(.dout(w_dff_A_7jkH8cLA8_0),.din(w_dff_A_yDCvhztt5_0),.clk(gclk));
	jdff dff_A_SXewAdwv0_0(.dout(w_dff_A_yDCvhztt5_0),.din(w_dff_A_SXewAdwv0_0),.clk(gclk));
	jdff dff_A_tgyV8E6r7_0(.dout(w_n156_0[0]),.din(w_dff_A_tgyV8E6r7_0),.clk(gclk));
	jdff dff_A_1Jq4nkXF1_0(.dout(w_dff_A_tgyV8E6r7_0),.din(w_dff_A_1Jq4nkXF1_0),.clk(gclk));
	jdff dff_A_yJLP9fDB7_0(.dout(w_dff_A_1Jq4nkXF1_0),.din(w_dff_A_yJLP9fDB7_0),.clk(gclk));
	jdff dff_A_bIl8ee3p0_0(.dout(w_dff_A_yJLP9fDB7_0),.din(w_dff_A_bIl8ee3p0_0),.clk(gclk));
	jdff dff_A_WQ2gkHU33_0(.dout(w_dff_A_bIl8ee3p0_0),.din(w_dff_A_WQ2gkHU33_0),.clk(gclk));
	jdff dff_A_CZVKhSoJ6_0(.dout(w_dff_A_WQ2gkHU33_0),.din(w_dff_A_CZVKhSoJ6_0),.clk(gclk));
	jdff dff_A_lPNB9SXU5_0(.dout(w_n154_0[0]),.din(w_dff_A_lPNB9SXU5_0),.clk(gclk));
	jdff dff_A_7Ts3aUSM7_0(.dout(w_dff_A_lPNB9SXU5_0),.din(w_dff_A_7Ts3aUSM7_0),.clk(gclk));
	jdff dff_A_f1iMwhNx3_0(.dout(w_dff_A_7Ts3aUSM7_0),.din(w_dff_A_f1iMwhNx3_0),.clk(gclk));
	jdff dff_A_FZkAdwT63_0(.dout(w_dff_A_f1iMwhNx3_0),.din(w_dff_A_FZkAdwT63_0),.clk(gclk));
	jdff dff_A_KANBbx909_0(.dout(w_dff_A_FZkAdwT63_0),.din(w_dff_A_KANBbx909_0),.clk(gclk));
	jdff dff_B_MIhgDrZp5_2(.din(n154),.dout(w_dff_B_MIhgDrZp5_2),.clk(gclk));
	jdff dff_B_QuZuGzNj1_2(.din(w_dff_B_MIhgDrZp5_2),.dout(w_dff_B_QuZuGzNj1_2),.clk(gclk));
	jdff dff_B_vuG75snK7_2(.din(w_dff_B_QuZuGzNj1_2),.dout(w_dff_B_vuG75snK7_2),.clk(gclk));
	jdff dff_B_AbNuQma71_2(.din(w_dff_B_vuG75snK7_2),.dout(w_dff_B_AbNuQma71_2),.clk(gclk));
	jdff dff_B_Zkvwf1hd9_2(.din(w_dff_B_AbNuQma71_2),.dout(w_dff_B_Zkvwf1hd9_2),.clk(gclk));
	jdff dff_B_1k3jrDMp1_2(.din(w_dff_B_Zkvwf1hd9_2),.dout(w_dff_B_1k3jrDMp1_2),.clk(gclk));
	jdff dff_B_3eMPSOt68_2(.din(w_dff_B_1k3jrDMp1_2),.dout(w_dff_B_3eMPSOt68_2),.clk(gclk));
	jdff dff_B_jGDwblWz6_2(.din(w_dff_B_3eMPSOt68_2),.dout(w_dff_B_jGDwblWz6_2),.clk(gclk));
	jdff dff_B_bcqC3Odf5_2(.din(w_dff_B_jGDwblWz6_2),.dout(w_dff_B_bcqC3Odf5_2),.clk(gclk));
	jdff dff_B_UNxknqTt3_2(.din(w_dff_B_bcqC3Odf5_2),.dout(w_dff_B_UNxknqTt3_2),.clk(gclk));
	jdff dff_B_QNKmPUo10_2(.din(w_dff_B_UNxknqTt3_2),.dout(w_dff_B_QNKmPUo10_2),.clk(gclk));
	jdff dff_B_V9oMdfJU2_2(.din(w_dff_B_QNKmPUo10_2),.dout(w_dff_B_V9oMdfJU2_2),.clk(gclk));
	jdff dff_B_lDNCmbYg3_2(.din(w_dff_B_V9oMdfJU2_2),.dout(w_dff_B_lDNCmbYg3_2),.clk(gclk));
	jdff dff_B_R2JwCoqq6_2(.din(w_dff_B_lDNCmbYg3_2),.dout(w_dff_B_R2JwCoqq6_2),.clk(gclk));
	jdff dff_A_g6hg80xF5_1(.dout(w_n146_0[1]),.din(w_dff_A_g6hg80xF5_1),.clk(gclk));
	jdff dff_A_6uNmkRof2_1(.dout(w_dff_A_g6hg80xF5_1),.din(w_dff_A_6uNmkRof2_1),.clk(gclk));
	jdff dff_A_T4EavMuv3_1(.dout(w_dff_A_6uNmkRof2_1),.din(w_dff_A_T4EavMuv3_1),.clk(gclk));
	jdff dff_A_iDTa47vb4_1(.dout(w_dff_A_T4EavMuv3_1),.din(w_dff_A_iDTa47vb4_1),.clk(gclk));
	jdff dff_A_Sd3vZQAW8_0(.dout(w_n145_0[0]),.din(w_dff_A_Sd3vZQAW8_0),.clk(gclk));
	jdff dff_A_TWd66Ggc0_0(.dout(w_dff_A_Sd3vZQAW8_0),.din(w_dff_A_TWd66Ggc0_0),.clk(gclk));
	jdff dff_A_ZFkON3pV8_0(.dout(w_dff_A_TWd66Ggc0_0),.din(w_dff_A_ZFkON3pV8_0),.clk(gclk));
	jdff dff_A_tC9e8ZTm8_0(.dout(w_dff_A_ZFkON3pV8_0),.din(w_dff_A_tC9e8ZTm8_0),.clk(gclk));
	jdff dff_A_Tv1nYxhP5_0(.dout(w_dff_A_tC9e8ZTm8_0),.din(w_dff_A_Tv1nYxhP5_0),.clk(gclk));
	jdff dff_A_HK2fndwt2_0(.dout(w_dff_A_Tv1nYxhP5_0),.din(w_dff_A_HK2fndwt2_0),.clk(gclk));
	jdff dff_A_HeeEoTy64_0(.dout(w_n142_0[0]),.din(w_dff_A_HeeEoTy64_0),.clk(gclk));
	jdff dff_A_n5GzK4zV6_1(.dout(w_n139_0[1]),.din(w_dff_A_n5GzK4zV6_1),.clk(gclk));
	jdff dff_A_DoLX5AFt6_1(.dout(w_dff_A_n5GzK4zV6_1),.din(w_dff_A_DoLX5AFt6_1),.clk(gclk));
	jdff dff_A_YaurMj0r3_1(.dout(w_dff_A_DoLX5AFt6_1),.din(w_dff_A_YaurMj0r3_1),.clk(gclk));
	jdff dff_A_F6Ecdgn17_1(.dout(w_dff_A_YaurMj0r3_1),.din(w_dff_A_F6Ecdgn17_1),.clk(gclk));
	jdff dff_A_O5uDvHnT1_1(.dout(w_dff_A_F6Ecdgn17_1),.din(w_dff_A_O5uDvHnT1_1),.clk(gclk));
	jdff dff_A_4wpWuhcS5_1(.dout(w_dff_A_O5uDvHnT1_1),.din(w_dff_A_4wpWuhcS5_1),.clk(gclk));
	jdff dff_A_U2myqVlw1_2(.dout(w_dff_A_r1PolYoN8_0),.din(w_dff_A_U2myqVlw1_2),.clk(gclk));
	jdff dff_A_r1PolYoN8_0(.dout(w_dff_A_npYM2eh68_0),.din(w_dff_A_r1PolYoN8_0),.clk(gclk));
	jdff dff_A_npYM2eh68_0(.dout(w_dff_A_vxUEi8dk1_0),.din(w_dff_A_npYM2eh68_0),.clk(gclk));
	jdff dff_A_vxUEi8dk1_0(.dout(w_dff_A_oDi1ha292_0),.din(w_dff_A_vxUEi8dk1_0),.clk(gclk));
	jdff dff_A_oDi1ha292_0(.dout(w_dff_A_LP3ezWcE7_0),.din(w_dff_A_oDi1ha292_0),.clk(gclk));
	jdff dff_A_LP3ezWcE7_0(.dout(w_dff_A_5IA7FVEp8_0),.din(w_dff_A_LP3ezWcE7_0),.clk(gclk));
	jdff dff_A_5IA7FVEp8_0(.dout(w_dff_A_rUXUmbIs5_0),.din(w_dff_A_5IA7FVEp8_0),.clk(gclk));
	jdff dff_A_rUXUmbIs5_0(.dout(w_dff_A_WfCN4ii01_0),.din(w_dff_A_rUXUmbIs5_0),.clk(gclk));
	jdff dff_A_WfCN4ii01_0(.dout(w_dff_A_FEVZJuwM1_0),.din(w_dff_A_WfCN4ii01_0),.clk(gclk));
	jdff dff_A_FEVZJuwM1_0(.dout(w_dff_A_qrQbfMeW7_0),.din(w_dff_A_FEVZJuwM1_0),.clk(gclk));
	jdff dff_A_qrQbfMeW7_0(.dout(w_dff_A_LDgfQkT33_0),.din(w_dff_A_qrQbfMeW7_0),.clk(gclk));
	jdff dff_A_LDgfQkT33_0(.dout(w_dff_A_Rn7gZ7Wo9_0),.din(w_dff_A_LDgfQkT33_0),.clk(gclk));
	jdff dff_A_Rn7gZ7Wo9_0(.dout(w_dff_A_ILLmIjGa0_0),.din(w_dff_A_Rn7gZ7Wo9_0),.clk(gclk));
	jdff dff_A_ILLmIjGa0_0(.dout(w_dff_A_ThmFGEWB0_0),.din(w_dff_A_ILLmIjGa0_0),.clk(gclk));
	jdff dff_A_ThmFGEWB0_0(.dout(w_dff_A_IbJyhUjl3_0),.din(w_dff_A_ThmFGEWB0_0),.clk(gclk));
	jdff dff_A_IbJyhUjl3_0(.dout(w_dff_A_drZFLKzm1_0),.din(w_dff_A_IbJyhUjl3_0),.clk(gclk));
	jdff dff_A_drZFLKzm1_0(.dout(w_dff_A_DHS1iso26_0),.din(w_dff_A_drZFLKzm1_0),.clk(gclk));
	jdff dff_A_DHS1iso26_0(.dout(w_dff_A_BntL2tG77_0),.din(w_dff_A_DHS1iso26_0),.clk(gclk));
	jdff dff_A_BntL2tG77_0(.dout(w_dff_A_PCOFOU9c5_0),.din(w_dff_A_BntL2tG77_0),.clk(gclk));
	jdff dff_A_PCOFOU9c5_0(.dout(G223gat),.din(w_dff_A_PCOFOU9c5_0),.clk(gclk));
	jdff dff_A_6BlOj4PO6_1(.dout(w_dff_A_gJ9QO1IN4_0),.din(w_dff_A_6BlOj4PO6_1),.clk(gclk));
	jdff dff_A_gJ9QO1IN4_0(.dout(w_dff_A_YyOfjQmG0_0),.din(w_dff_A_gJ9QO1IN4_0),.clk(gclk));
	jdff dff_A_YyOfjQmG0_0(.dout(w_dff_A_VNlNLTow8_0),.din(w_dff_A_YyOfjQmG0_0),.clk(gclk));
	jdff dff_A_VNlNLTow8_0(.dout(w_dff_A_ei14NpkH3_0),.din(w_dff_A_VNlNLTow8_0),.clk(gclk));
	jdff dff_A_ei14NpkH3_0(.dout(w_dff_A_nXsGjgZx3_0),.din(w_dff_A_ei14NpkH3_0),.clk(gclk));
	jdff dff_A_nXsGjgZx3_0(.dout(w_dff_A_PEk6LAkq2_0),.din(w_dff_A_nXsGjgZx3_0),.clk(gclk));
	jdff dff_A_PEk6LAkq2_0(.dout(w_dff_A_geYzOqFe7_0),.din(w_dff_A_PEk6LAkq2_0),.clk(gclk));
	jdff dff_A_geYzOqFe7_0(.dout(w_dff_A_OewmXfb11_0),.din(w_dff_A_geYzOqFe7_0),.clk(gclk));
	jdff dff_A_OewmXfb11_0(.dout(w_dff_A_HoXvt9rV9_0),.din(w_dff_A_OewmXfb11_0),.clk(gclk));
	jdff dff_A_HoXvt9rV9_0(.dout(w_dff_A_4pRC4xYS3_0),.din(w_dff_A_HoXvt9rV9_0),.clk(gclk));
	jdff dff_A_4pRC4xYS3_0(.dout(w_dff_A_mWAVF39O0_0),.din(w_dff_A_4pRC4xYS3_0),.clk(gclk));
	jdff dff_A_mWAVF39O0_0(.dout(w_dff_A_zFdNpgDY2_0),.din(w_dff_A_mWAVF39O0_0),.clk(gclk));
	jdff dff_A_zFdNpgDY2_0(.dout(G329gat),.din(w_dff_A_zFdNpgDY2_0),.clk(gclk));
	jdff dff_A_iURVVgb10_1(.dout(w_dff_A_6oMFTJmt9_0),.din(w_dff_A_iURVVgb10_1),.clk(gclk));
	jdff dff_A_6oMFTJmt9_0(.dout(w_dff_A_Z3cxfR5c0_0),.din(w_dff_A_6oMFTJmt9_0),.clk(gclk));
	jdff dff_A_Z3cxfR5c0_0(.dout(w_dff_A_T4u4e5Ml8_0),.din(w_dff_A_Z3cxfR5c0_0),.clk(gclk));
	jdff dff_A_T4u4e5Ml8_0(.dout(w_dff_A_zyEgun1U8_0),.din(w_dff_A_T4u4e5Ml8_0),.clk(gclk));
	jdff dff_A_zyEgun1U8_0(.dout(w_dff_A_l0pFLbh48_0),.din(w_dff_A_zyEgun1U8_0),.clk(gclk));
	jdff dff_A_l0pFLbh48_0(.dout(G370gat),.din(w_dff_A_l0pFLbh48_0),.clk(gclk));
	jdff dff_A_C8M0FakO9_1(.dout(w_dff_A_gmAmFeKr4_0),.din(w_dff_A_C8M0FakO9_1),.clk(gclk));
	jdff dff_A_gmAmFeKr4_0(.dout(G430gat),.din(w_dff_A_gmAmFeKr4_0),.clk(gclk));
endmodule

