/*

top:
	jxor: 603
	jspl: 1591
	jspl3: 1428
	jnot: 630
	jdff: 985
	jor: 1152
	jand: 2691

Summary:
	jxor: 603
	jspl: 1591
	jspl3: 1428
	jnot: 630
	jdff: 985
	jor: 1152
	jand: 2691

The maximum logic level gap of any gate:
	top: 127
*/

module rf_sin(gclk, a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, sin0, sin1, sin2, sin3, sin4, sin5, sin6, sin7, sin8, sin9, sin10, sin11, sin12, sin13, sin14, sin15, sin16, sin17, sin18, sin19, sin20, sin21, sin22, sin23, sin24);
	input gclk;
	input a0;
	input a1;
	input a2;
	input a3;
	input a4;
	input a5;
	input a6;
	input a7;
	input a8;
	input a9;
	input a10;
	input a11;
	input a12;
	input a13;
	input a14;
	input a15;
	input a16;
	input a17;
	input a18;
	input a19;
	input a20;
	input a21;
	input a22;
	input a23;
	output sin0;
	output sin1;
	output sin2;
	output sin3;
	output sin4;
	output sin5;
	output sin6;
	output sin7;
	output sin8;
	output sin9;
	output sin10;
	output sin11;
	output sin12;
	output sin13;
	output sin14;
	output sin15;
	output sin16;
	output sin17;
	output sin18;
	output sin19;
	output sin20;
	output sin21;
	output sin22;
	output sin23;
	output sin24;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n808;
	wire n810;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1063;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1100;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1147;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1704;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1821;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1837;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire n1852;
	wire n1853;
	wire n1854;
	wire n1855;
	wire n1856;
	wire n1857;
	wire n1858;
	wire n1859;
	wire n1860;
	wire n1861;
	wire n1862;
	wire n1863;
	wire n1864;
	wire n1865;
	wire n1866;
	wire n1867;
	wire n1868;
	wire n1869;
	wire n1870;
	wire n1871;
	wire n1872;
	wire n1873;
	wire n1874;
	wire n1875;
	wire n1876;
	wire n1877;
	wire n1878;
	wire n1879;
	wire n1880;
	wire n1881;
	wire n1882;
	wire n1883;
	wire n1884;
	wire n1885;
	wire n1886;
	wire n1887;
	wire n1888;
	wire n1889;
	wire n1890;
	wire n1891;
	wire n1892;
	wire n1893;
	wire n1894;
	wire n1895;
	wire n1896;
	wire n1897;
	wire n1898;
	wire n1899;
	wire n1900;
	wire n1901;
	wire n1902;
	wire n1903;
	wire n1904;
	wire n1905;
	wire n1906;
	wire n1907;
	wire n1908;
	wire n1909;
	wire n1910;
	wire n1911;
	wire n1912;
	wire n1913;
	wire n1914;
	wire n1915;
	wire n1916;
	wire n1917;
	wire n1918;
	wire n1919;
	wire n1920;
	wire n1921;
	wire n1922;
	wire n1923;
	wire n1924;
	wire n1925;
	wire n1926;
	wire n1927;
	wire n1928;
	wire n1929;
	wire n1930;
	wire n1931;
	wire n1932;
	wire n1933;
	wire n1934;
	wire n1935;
	wire n1936;
	wire n1937;
	wire n1938;
	wire n1939;
	wire n1940;
	wire n1941;
	wire n1942;
	wire n1943;
	wire n1944;
	wire n1945;
	wire n1946;
	wire n1947;
	wire n1948;
	wire n1949;
	wire n1950;
	wire n1951;
	wire n1952;
	wire n1953;
	wire n1954;
	wire n1955;
	wire n1956;
	wire n1957;
	wire n1958;
	wire n1959;
	wire n1960;
	wire n1961;
	wire n1962;
	wire n1963;
	wire n1964;
	wire n1965;
	wire n1966;
	wire n1967;
	wire n1968;
	wire n1969;
	wire n1970;
	wire n1971;
	wire n1972;
	wire n1973;
	wire n1974;
	wire n1975;
	wire n1976;
	wire n1977;
	wire n1978;
	wire n1979;
	wire n1980;
	wire n1981;
	wire n1982;
	wire n1983;
	wire n1984;
	wire n1985;
	wire n1986;
	wire n1987;
	wire n1988;
	wire n1989;
	wire n1990;
	wire n1991;
	wire n1992;
	wire n1993;
	wire n1994;
	wire n1995;
	wire n1996;
	wire n1997;
	wire n1998;
	wire n1999;
	wire n2000;
	wire n2001;
	wire n2002;
	wire n2003;
	wire n2004;
	wire n2005;
	wire n2006;
	wire n2007;
	wire n2008;
	wire n2009;
	wire n2010;
	wire n2011;
	wire n2012;
	wire n2013;
	wire n2014;
	wire n2015;
	wire n2016;
	wire n2017;
	wire n2018;
	wire n2019;
	wire n2020;
	wire n2021;
	wire n2022;
	wire n2023;
	wire n2024;
	wire n2025;
	wire n2026;
	wire n2027;
	wire n2028;
	wire n2029;
	wire n2030;
	wire n2031;
	wire n2032;
	wire n2033;
	wire n2034;
	wire n2035;
	wire n2036;
	wire n2037;
	wire n2038;
	wire n2039;
	wire n2040;
	wire n2041;
	wire n2042;
	wire n2043;
	wire n2044;
	wire n2045;
	wire n2046;
	wire n2047;
	wire n2048;
	wire n2049;
	wire n2050;
	wire n2051;
	wire n2052;
	wire n2053;
	wire n2054;
	wire n2055;
	wire n2056;
	wire n2057;
	wire n2058;
	wire n2059;
	wire n2060;
	wire n2061;
	wire n2062;
	wire n2063;
	wire n2064;
	wire n2065;
	wire n2066;
	wire n2067;
	wire n2068;
	wire n2069;
	wire n2070;
	wire n2071;
	wire n2072;
	wire n2073;
	wire n2074;
	wire n2075;
	wire n2076;
	wire n2077;
	wire n2078;
	wire n2079;
	wire n2080;
	wire n2081;
	wire n2082;
	wire n2083;
	wire n2084;
	wire n2085;
	wire n2086;
	wire n2087;
	wire n2088;
	wire n2089;
	wire n2090;
	wire n2091;
	wire n2092;
	wire n2093;
	wire n2094;
	wire n2095;
	wire n2096;
	wire n2097;
	wire n2098;
	wire n2099;
	wire n2100;
	wire n2101;
	wire n2102;
	wire n2103;
	wire n2104;
	wire n2105;
	wire n2106;
	wire n2107;
	wire n2108;
	wire n2109;
	wire n2110;
	wire n2111;
	wire n2112;
	wire n2113;
	wire n2114;
	wire n2115;
	wire n2116;
	wire n2117;
	wire n2118;
	wire n2119;
	wire n2120;
	wire n2121;
	wire n2122;
	wire n2123;
	wire n2124;
	wire n2125;
	wire n2126;
	wire n2127;
	wire n2128;
	wire n2129;
	wire n2130;
	wire n2131;
	wire n2132;
	wire n2133;
	wire n2134;
	wire n2135;
	wire n2136;
	wire n2137;
	wire n2138;
	wire n2139;
	wire n2140;
	wire n2141;
	wire n2142;
	wire n2143;
	wire n2144;
	wire n2145;
	wire n2146;
	wire n2147;
	wire n2148;
	wire n2149;
	wire n2150;
	wire n2151;
	wire n2152;
	wire n2153;
	wire n2154;
	wire n2155;
	wire n2156;
	wire n2157;
	wire n2158;
	wire n2159;
	wire n2160;
	wire n2161;
	wire n2162;
	wire n2163;
	wire n2164;
	wire n2165;
	wire n2166;
	wire n2167;
	wire n2168;
	wire n2169;
	wire n2170;
	wire n2171;
	wire n2172;
	wire n2173;
	wire n2174;
	wire n2175;
	wire n2176;
	wire n2177;
	wire n2178;
	wire n2179;
	wire n2180;
	wire n2181;
	wire n2182;
	wire n2183;
	wire n2184;
	wire n2185;
	wire n2186;
	wire n2187;
	wire n2188;
	wire n2189;
	wire n2190;
	wire n2191;
	wire n2192;
	wire n2193;
	wire n2194;
	wire n2195;
	wire n2196;
	wire n2197;
	wire n2198;
	wire n2199;
	wire n2200;
	wire n2201;
	wire n2202;
	wire n2203;
	wire n2204;
	wire n2205;
	wire n2206;
	wire n2207;
	wire n2208;
	wire n2209;
	wire n2210;
	wire n2211;
	wire n2212;
	wire n2213;
	wire n2214;
	wire n2215;
	wire n2216;
	wire n2217;
	wire n2218;
	wire n2219;
	wire n2220;
	wire n2221;
	wire n2222;
	wire n2223;
	wire n2224;
	wire n2225;
	wire n2226;
	wire n2227;
	wire n2228;
	wire n2229;
	wire n2230;
	wire n2231;
	wire n2232;
	wire n2233;
	wire n2234;
	wire n2235;
	wire n2236;
	wire n2237;
	wire n2238;
	wire n2239;
	wire n2240;
	wire n2241;
	wire n2242;
	wire n2243;
	wire n2244;
	wire n2245;
	wire n2246;
	wire n2247;
	wire n2248;
	wire n2249;
	wire n2250;
	wire n2251;
	wire n2252;
	wire n2253;
	wire n2254;
	wire n2255;
	wire n2256;
	wire n2257;
	wire n2258;
	wire n2259;
	wire n2260;
	wire n2261;
	wire n2262;
	wire n2263;
	wire n2264;
	wire n2265;
	wire n2266;
	wire n2267;
	wire n2268;
	wire n2269;
	wire n2270;
	wire n2272;
	wire n2275;
	wire n2276;
	wire n2277;
	wire n2278;
	wire n2279;
	wire n2280;
	wire n2281;
	wire n2282;
	wire n2283;
	wire n2284;
	wire n2285;
	wire n2286;
	wire n2287;
	wire n2288;
	wire n2289;
	wire n2290;
	wire n2291;
	wire n2292;
	wire n2293;
	wire n2294;
	wire n2295;
	wire n2296;
	wire n2297;
	wire n2298;
	wire n2299;
	wire n2300;
	wire n2301;
	wire n2302;
	wire n2303;
	wire n2304;
	wire n2305;
	wire n2306;
	wire n2307;
	wire n2308;
	wire n2309;
	wire n2310;
	wire n2311;
	wire n2312;
	wire n2313;
	wire n2314;
	wire n2315;
	wire n2316;
	wire n2317;
	wire n2318;
	wire n2319;
	wire n2320;
	wire n2321;
	wire n2322;
	wire n2323;
	wire n2324;
	wire n2325;
	wire n2326;
	wire n2327;
	wire n2328;
	wire n2329;
	wire n2330;
	wire n2331;
	wire n2332;
	wire n2333;
	wire n2334;
	wire n2335;
	wire n2336;
	wire n2337;
	wire n2338;
	wire n2339;
	wire n2340;
	wire n2341;
	wire n2342;
	wire n2343;
	wire n2344;
	wire n2345;
	wire n2346;
	wire n2347;
	wire n2348;
	wire n2349;
	wire n2350;
	wire n2351;
	wire n2352;
	wire n2353;
	wire n2354;
	wire n2355;
	wire n2356;
	wire n2357;
	wire n2358;
	wire n2359;
	wire n2360;
	wire n2361;
	wire n2362;
	wire n2363;
	wire n2364;
	wire n2365;
	wire n2366;
	wire n2367;
	wire n2368;
	wire n2369;
	wire n2370;
	wire n2371;
	wire n2372;
	wire n2373;
	wire n2374;
	wire n2375;
	wire n2376;
	wire n2377;
	wire n2378;
	wire n2379;
	wire n2380;
	wire n2381;
	wire n2382;
	wire n2383;
	wire n2384;
	wire n2385;
	wire n2386;
	wire n2387;
	wire n2388;
	wire n2389;
	wire n2390;
	wire n2391;
	wire n2392;
	wire n2393;
	wire n2394;
	wire n2395;
	wire n2396;
	wire n2397;
	wire n2398;
	wire n2399;
	wire n2400;
	wire n2401;
	wire n2402;
	wire n2403;
	wire n2404;
	wire n2405;
	wire n2406;
	wire n2407;
	wire n2408;
	wire n2409;
	wire n2410;
	wire n2411;
	wire n2412;
	wire n2413;
	wire n2414;
	wire n2415;
	wire n2416;
	wire n2417;
	wire n2418;
	wire n2419;
	wire n2420;
	wire n2421;
	wire n2422;
	wire n2423;
	wire n2424;
	wire n2425;
	wire n2426;
	wire n2427;
	wire n2428;
	wire n2429;
	wire n2430;
	wire n2431;
	wire n2432;
	wire n2433;
	wire n2434;
	wire n2435;
	wire n2436;
	wire n2437;
	wire n2438;
	wire n2439;
	wire n2440;
	wire n2441;
	wire n2442;
	wire n2443;
	wire n2444;
	wire n2445;
	wire n2446;
	wire n2447;
	wire n2448;
	wire n2449;
	wire n2450;
	wire n2451;
	wire n2452;
	wire n2453;
	wire n2454;
	wire n2455;
	wire n2456;
	wire n2457;
	wire n2458;
	wire n2459;
	wire n2460;
	wire n2461;
	wire n2462;
	wire n2463;
	wire n2464;
	wire n2465;
	wire n2466;
	wire n2467;
	wire n2468;
	wire n2469;
	wire n2470;
	wire n2471;
	wire n2472;
	wire n2473;
	wire n2474;
	wire n2475;
	wire n2476;
	wire n2477;
	wire n2478;
	wire n2479;
	wire n2480;
	wire n2481;
	wire n2482;
	wire n2483;
	wire n2484;
	wire n2485;
	wire n2486;
	wire n2487;
	wire n2488;
	wire n2489;
	wire n2490;
	wire n2491;
	wire n2492;
	wire n2493;
	wire n2494;
	wire n2495;
	wire n2496;
	wire n2497;
	wire n2498;
	wire n2499;
	wire n2500;
	wire n2501;
	wire n2502;
	wire n2503;
	wire n2504;
	wire n2505;
	wire n2506;
	wire n2507;
	wire n2508;
	wire n2509;
	wire n2510;
	wire n2511;
	wire n2512;
	wire n2513;
	wire n2514;
	wire n2515;
	wire n2516;
	wire n2517;
	wire n2518;
	wire n2519;
	wire n2520;
	wire n2521;
	wire n2522;
	wire n2523;
	wire n2524;
	wire n2525;
	wire n2526;
	wire n2527;
	wire n2528;
	wire n2529;
	wire n2530;
	wire n2531;
	wire n2532;
	wire n2533;
	wire n2534;
	wire n2535;
	wire n2536;
	wire n2537;
	wire n2538;
	wire n2539;
	wire n2540;
	wire n2541;
	wire n2542;
	wire n2543;
	wire n2544;
	wire n2545;
	wire n2546;
	wire n2547;
	wire n2548;
	wire n2549;
	wire n2550;
	wire n2551;
	wire n2552;
	wire n2553;
	wire n2554;
	wire n2555;
	wire n2556;
	wire n2557;
	wire n2558;
	wire n2559;
	wire n2560;
	wire n2561;
	wire n2562;
	wire n2563;
	wire n2564;
	wire n2565;
	wire n2566;
	wire n2567;
	wire n2568;
	wire n2569;
	wire n2570;
	wire n2571;
	wire n2572;
	wire n2573;
	wire n2574;
	wire n2575;
	wire n2576;
	wire n2577;
	wire n2578;
	wire n2579;
	wire n2580;
	wire n2581;
	wire n2582;
	wire n2583;
	wire n2584;
	wire n2585;
	wire n2586;
	wire n2587;
	wire n2588;
	wire n2589;
	wire n2590;
	wire n2591;
	wire n2592;
	wire n2593;
	wire n2594;
	wire n2595;
	wire n2596;
	wire n2597;
	wire n2598;
	wire n2599;
	wire n2600;
	wire n2601;
	wire n2602;
	wire n2603;
	wire n2604;
	wire n2605;
	wire n2606;
	wire n2607;
	wire n2608;
	wire n2609;
	wire n2610;
	wire n2611;
	wire n2612;
	wire n2613;
	wire n2614;
	wire n2615;
	wire n2616;
	wire n2617;
	wire n2618;
	wire n2619;
	wire n2620;
	wire n2621;
	wire n2622;
	wire n2623;
	wire n2624;
	wire n2625;
	wire n2626;
	wire n2627;
	wire n2628;
	wire n2629;
	wire n2630;
	wire n2632;
	wire n2633;
	wire n2634;
	wire n2635;
	wire n2636;
	wire n2637;
	wire n2638;
	wire n2639;
	wire n2640;
	wire n2641;
	wire n2642;
	wire n2643;
	wire n2644;
	wire n2645;
	wire n2646;
	wire n2647;
	wire n2648;
	wire n2649;
	wire n2650;
	wire n2651;
	wire n2652;
	wire n2653;
	wire n2654;
	wire n2655;
	wire n2656;
	wire n2657;
	wire n2658;
	wire n2659;
	wire n2660;
	wire n2661;
	wire n2662;
	wire n2663;
	wire n2664;
	wire n2665;
	wire n2666;
	wire n2667;
	wire n2668;
	wire n2669;
	wire n2670;
	wire n2671;
	wire n2672;
	wire n2673;
	wire n2674;
	wire n2675;
	wire n2676;
	wire n2677;
	wire n2678;
	wire n2679;
	wire n2680;
	wire n2681;
	wire n2682;
	wire n2683;
	wire n2684;
	wire n2685;
	wire n2686;
	wire n2687;
	wire n2688;
	wire n2689;
	wire n2690;
	wire n2691;
	wire n2692;
	wire n2693;
	wire n2694;
	wire n2695;
	wire n2696;
	wire n2697;
	wire n2698;
	wire n2699;
	wire n2700;
	wire n2701;
	wire n2702;
	wire n2703;
	wire n2704;
	wire n2705;
	wire n2706;
	wire n2707;
	wire n2708;
	wire n2709;
	wire n2710;
	wire n2711;
	wire n2712;
	wire n2713;
	wire n2714;
	wire n2715;
	wire n2716;
	wire n2717;
	wire n2718;
	wire n2719;
	wire n2720;
	wire n2721;
	wire n2722;
	wire n2723;
	wire n2724;
	wire n2725;
	wire n2726;
	wire n2727;
	wire n2728;
	wire n2729;
	wire n2730;
	wire n2731;
	wire n2732;
	wire n2733;
	wire n2734;
	wire n2735;
	wire n2736;
	wire n2737;
	wire n2738;
	wire n2739;
	wire n2740;
	wire n2741;
	wire n2742;
	wire n2743;
	wire n2744;
	wire n2745;
	wire n2746;
	wire n2747;
	wire n2748;
	wire n2749;
	wire n2750;
	wire n2751;
	wire n2752;
	wire n2753;
	wire n2754;
	wire n2757;
	wire n2758;
	wire n2759;
	wire n2760;
	wire n2761;
	wire n2762;
	wire n2763;
	wire n2764;
	wire n2765;
	wire n2766;
	wire n2767;
	wire n2768;
	wire n2769;
	wire n2770;
	wire n2771;
	wire n2772;
	wire n2773;
	wire n2774;
	wire n2775;
	wire n2776;
	wire n2777;
	wire n2778;
	wire n2779;
	wire n2780;
	wire n2781;
	wire n2782;
	wire n2783;
	wire n2784;
	wire n2785;
	wire n2786;
	wire n2787;
	wire n2788;
	wire n2789;
	wire n2790;
	wire n2791;
	wire n2792;
	wire n2793;
	wire n2794;
	wire n2795;
	wire n2796;
	wire n2797;
	wire n2798;
	wire n2799;
	wire n2800;
	wire n2801;
	wire n2802;
	wire n2803;
	wire n2804;
	wire n2805;
	wire n2806;
	wire n2807;
	wire n2808;
	wire n2809;
	wire n2810;
	wire n2811;
	wire n2812;
	wire n2813;
	wire n2814;
	wire n2815;
	wire n2816;
	wire n2817;
	wire n2818;
	wire n2819;
	wire n2820;
	wire n2821;
	wire n2822;
	wire n2823;
	wire n2824;
	wire n2825;
	wire n2826;
	wire n2827;
	wire n2828;
	wire n2829;
	wire n2830;
	wire n2831;
	wire n2832;
	wire n2833;
	wire n2834;
	wire n2835;
	wire n2836;
	wire n2837;
	wire n2838;
	wire n2839;
	wire n2840;
	wire n2841;
	wire n2842;
	wire n2843;
	wire n2844;
	wire n2845;
	wire n2846;
	wire n2847;
	wire n2848;
	wire n2849;
	wire n2850;
	wire n2851;
	wire n2852;
	wire n2853;
	wire n2854;
	wire n2855;
	wire n2856;
	wire n2857;
	wire n2858;
	wire n2859;
	wire n2860;
	wire n2861;
	wire n2862;
	wire n2863;
	wire n2864;
	wire n2865;
	wire n2866;
	wire n2867;
	wire n2868;
	wire n2869;
	wire n2870;
	wire n2871;
	wire n2872;
	wire n2873;
	wire n2874;
	wire n2875;
	wire n2876;
	wire n2877;
	wire n2878;
	wire n2879;
	wire n2880;
	wire n2881;
	wire n2882;
	wire n2883;
	wire n2884;
	wire n2885;
	wire n2886;
	wire n2887;
	wire n2888;
	wire n2889;
	wire n2890;
	wire n2891;
	wire n2892;
	wire n2893;
	wire n2894;
	wire n2895;
	wire n2896;
	wire n2897;
	wire n2898;
	wire n2899;
	wire n2900;
	wire n2901;
	wire n2902;
	wire n2903;
	wire n2904;
	wire n2905;
	wire n2906;
	wire n2907;
	wire n2908;
	wire n2909;
	wire n2910;
	wire n2911;
	wire n2912;
	wire n2913;
	wire n2914;
	wire n2915;
	wire n2916;
	wire n2917;
	wire n2918;
	wire n2919;
	wire n2920;
	wire n2921;
	wire n2922;
	wire n2923;
	wire n2924;
	wire n2925;
	wire n2926;
	wire n2927;
	wire n2928;
	wire n2929;
	wire n2930;
	wire n2931;
	wire n2932;
	wire n2933;
	wire n2934;
	wire n2935;
	wire n2936;
	wire n2937;
	wire n2938;
	wire n2939;
	wire n2940;
	wire n2941;
	wire n2942;
	wire n2943;
	wire n2944;
	wire n2945;
	wire n2946;
	wire n2947;
	wire n2948;
	wire n2949;
	wire n2950;
	wire n2951;
	wire n2952;
	wire n2953;
	wire n2954;
	wire n2955;
	wire n2956;
	wire n2957;
	wire n2958;
	wire n2959;
	wire n2960;
	wire n2961;
	wire n2962;
	wire n2963;
	wire n2964;
	wire n2965;
	wire n2966;
	wire n2967;
	wire n2968;
	wire n2969;
	wire n2970;
	wire n2971;
	wire n2972;
	wire n2973;
	wire n2974;
	wire n2975;
	wire n2976;
	wire n2977;
	wire n2978;
	wire n2979;
	wire n2980;
	wire n2981;
	wire n2982;
	wire n2983;
	wire n2984;
	wire n2985;
	wire n2986;
	wire n2987;
	wire n2988;
	wire n2989;
	wire n2990;
	wire n2991;
	wire n2992;
	wire n2993;
	wire n2994;
	wire n2995;
	wire n2996;
	wire n2997;
	wire n2998;
	wire n2999;
	wire n3000;
	wire n3001;
	wire n3002;
	wire n3003;
	wire n3004;
	wire n3005;
	wire n3006;
	wire n3007;
	wire n3008;
	wire n3009;
	wire n3010;
	wire n3011;
	wire n3012;
	wire n3013;
	wire n3014;
	wire n3015;
	wire n3016;
	wire n3017;
	wire n3018;
	wire n3019;
	wire n3020;
	wire n3021;
	wire n3022;
	wire n3023;
	wire n3024;
	wire n3025;
	wire n3026;
	wire n3027;
	wire n3028;
	wire n3029;
	wire n3030;
	wire n3031;
	wire n3032;
	wire n3033;
	wire n3034;
	wire n3035;
	wire n3036;
	wire n3037;
	wire n3038;
	wire n3039;
	wire n3040;
	wire n3041;
	wire n3042;
	wire n3043;
	wire n3044;
	wire n3045;
	wire n3046;
	wire n3047;
	wire n3048;
	wire n3049;
	wire n3050;
	wire n3051;
	wire n3052;
	wire n3053;
	wire n3054;
	wire n3055;
	wire n3056;
	wire n3057;
	wire n3058;
	wire n3059;
	wire n3060;
	wire n3061;
	wire n3062;
	wire n3063;
	wire n3064;
	wire n3065;
	wire n3066;
	wire n3067;
	wire n3068;
	wire n3069;
	wire n3070;
	wire n3071;
	wire n3072;
	wire n3073;
	wire n3074;
	wire n3075;
	wire n3076;
	wire n3077;
	wire n3078;
	wire n3079;
	wire n3080;
	wire n3081;
	wire n3082;
	wire n3083;
	wire n3084;
	wire n3085;
	wire n3086;
	wire n3087;
	wire n3088;
	wire n3089;
	wire n3090;
	wire n3091;
	wire n3092;
	wire n3093;
	wire n3094;
	wire n3095;
	wire n3096;
	wire n3097;
	wire n3098;
	wire n3099;
	wire n3100;
	wire n3101;
	wire n3102;
	wire n3103;
	wire n3104;
	wire n3105;
	wire n3106;
	wire n3107;
	wire n3108;
	wire n3109;
	wire n3110;
	wire n3111;
	wire n3112;
	wire n3113;
	wire n3114;
	wire n3115;
	wire n3116;
	wire n3117;
	wire n3118;
	wire n3119;
	wire n3120;
	wire n3121;
	wire n3122;
	wire n3123;
	wire n3124;
	wire n3125;
	wire n3126;
	wire n3127;
	wire n3128;
	wire n3129;
	wire n3130;
	wire n3131;
	wire n3132;
	wire n3133;
	wire n3134;
	wire n3135;
	wire n3136;
	wire n3137;
	wire n3138;
	wire n3139;
	wire n3140;
	wire n3141;
	wire n3142;
	wire n3143;
	wire n3144;
	wire n3145;
	wire n3146;
	wire n3147;
	wire n3148;
	wire n3149;
	wire n3150;
	wire n3151;
	wire n3152;
	wire n3153;
	wire n3154;
	wire n3155;
	wire n3156;
	wire n3157;
	wire n3158;
	wire n3159;
	wire n3160;
	wire n3161;
	wire n3162;
	wire n3163;
	wire n3164;
	wire n3165;
	wire n3166;
	wire n3167;
	wire n3168;
	wire n3169;
	wire n3170;
	wire n3171;
	wire n3172;
	wire n3173;
	wire n3174;
	wire n3175;
	wire n3176;
	wire n3177;
	wire n3178;
	wire n3179;
	wire n3180;
	wire n3181;
	wire n3182;
	wire n3183;
	wire n3184;
	wire n3185;
	wire n3186;
	wire n3187;
	wire n3188;
	wire n3189;
	wire n3190;
	wire n3191;
	wire n3192;
	wire n3193;
	wire n3194;
	wire n3195;
	wire n3196;
	wire n3197;
	wire n3198;
	wire n3199;
	wire n3200;
	wire n3201;
	wire n3202;
	wire n3203;
	wire n3204;
	wire n3205;
	wire n3206;
	wire n3207;
	wire n3208;
	wire n3209;
	wire n3210;
	wire n3211;
	wire n3212;
	wire n3213;
	wire n3214;
	wire n3215;
	wire n3216;
	wire n3217;
	wire n3218;
	wire n3219;
	wire n3220;
	wire n3221;
	wire n3222;
	wire n3223;
	wire n3224;
	wire n3225;
	wire n3226;
	wire n3227;
	wire n3228;
	wire n3229;
	wire n3230;
	wire n3231;
	wire n3232;
	wire n3233;
	wire n3234;
	wire n3235;
	wire n3236;
	wire n3237;
	wire n3238;
	wire n3239;
	wire n3240;
	wire n3241;
	wire n3242;
	wire n3243;
	wire n3244;
	wire n3245;
	wire n3246;
	wire n3247;
	wire n3248;
	wire n3249;
	wire n3250;
	wire n3251;
	wire n3252;
	wire n3253;
	wire n3254;
	wire n3255;
	wire n3256;
	wire n3257;
	wire n3258;
	wire n3259;
	wire n3260;
	wire n3261;
	wire n3262;
	wire n3263;
	wire n3264;
	wire n3265;
	wire n3266;
	wire n3267;
	wire n3268;
	wire n3269;
	wire n3270;
	wire n3271;
	wire n3272;
	wire n3273;
	wire n3274;
	wire n3275;
	wire n3276;
	wire n3277;
	wire n3278;
	wire n3279;
	wire n3280;
	wire n3281;
	wire n3282;
	wire n3283;
	wire n3284;
	wire n3285;
	wire n3286;
	wire n3287;
	wire n3288;
	wire n3289;
	wire n3290;
	wire n3291;
	wire n3292;
	wire n3293;
	wire n3294;
	wire n3295;
	wire n3296;
	wire n3297;
	wire n3298;
	wire n3299;
	wire n3300;
	wire n3301;
	wire n3302;
	wire n3303;
	wire n3304;
	wire n3305;
	wire n3306;
	wire n3307;
	wire n3308;
	wire n3309;
	wire n3310;
	wire n3311;
	wire n3312;
	wire n3313;
	wire n3314;
	wire n3315;
	wire n3316;
	wire n3317;
	wire n3318;
	wire n3319;
	wire n3320;
	wire n3321;
	wire n3322;
	wire n3323;
	wire n3324;
	wire n3325;
	wire n3326;
	wire n3327;
	wire n3328;
	wire n3329;
	wire n3330;
	wire n3331;
	wire n3332;
	wire n3333;
	wire n3334;
	wire n3335;
	wire n3336;
	wire n3337;
	wire n3338;
	wire n3339;
	wire n3340;
	wire n3341;
	wire n3342;
	wire n3343;
	wire n3344;
	wire n3345;
	wire n3346;
	wire n3347;
	wire n3348;
	wire n3349;
	wire n3350;
	wire n3351;
	wire n3352;
	wire n3353;
	wire n3354;
	wire n3355;
	wire n3356;
	wire n3357;
	wire n3358;
	wire n3359;
	wire n3360;
	wire n3361;
	wire n3362;
	wire n3363;
	wire n3364;
	wire n3365;
	wire n3366;
	wire n3367;
	wire n3368;
	wire n3369;
	wire n3370;
	wire n3371;
	wire n3372;
	wire n3373;
	wire n3374;
	wire n3375;
	wire n3376;
	wire n3377;
	wire n3378;
	wire n3379;
	wire n3380;
	wire n3381;
	wire n3382;
	wire n3383;
	wire n3384;
	wire n3385;
	wire n3386;
	wire n3387;
	wire n3388;
	wire n3389;
	wire n3390;
	wire n3391;
	wire n3392;
	wire n3393;
	wire n3394;
	wire n3395;
	wire n3396;
	wire n3397;
	wire n3398;
	wire n3399;
	wire n3400;
	wire n3401;
	wire n3402;
	wire n3403;
	wire n3404;
	wire n3405;
	wire n3406;
	wire n3407;
	wire n3408;
	wire n3409;
	wire n3410;
	wire n3411;
	wire n3412;
	wire n3413;
	wire n3414;
	wire n3415;
	wire n3416;
	wire n3417;
	wire n3418;
	wire n3419;
	wire n3420;
	wire n3421;
	wire n3422;
	wire n3423;
	wire n3424;
	wire n3425;
	wire n3426;
	wire n3427;
	wire n3428;
	wire n3429;
	wire n3430;
	wire n3431;
	wire n3432;
	wire n3433;
	wire n3434;
	wire n3435;
	wire n3436;
	wire n3437;
	wire n3438;
	wire n3439;
	wire n3440;
	wire n3441;
	wire n3442;
	wire n3443;
	wire n3444;
	wire n3445;
	wire n3446;
	wire n3447;
	wire n3448;
	wire n3449;
	wire n3450;
	wire n3451;
	wire n3452;
	wire n3453;
	wire n3454;
	wire n3455;
	wire n3456;
	wire n3457;
	wire n3458;
	wire n3459;
	wire n3460;
	wire n3461;
	wire n3462;
	wire n3463;
	wire n3464;
	wire n3465;
	wire n3466;
	wire n3467;
	wire n3468;
	wire n3469;
	wire n3470;
	wire n3471;
	wire n3472;
	wire n3473;
	wire n3474;
	wire n3475;
	wire n3476;
	wire n3477;
	wire n3478;
	wire n3479;
	wire n3480;
	wire n3481;
	wire n3482;
	wire n3483;
	wire n3484;
	wire n3485;
	wire n3486;
	wire n3487;
	wire n3488;
	wire n3489;
	wire n3490;
	wire n3491;
	wire n3492;
	wire n3493;
	wire n3494;
	wire n3495;
	wire n3496;
	wire n3497;
	wire n3498;
	wire n3499;
	wire n3500;
	wire n3501;
	wire n3502;
	wire n3503;
	wire n3504;
	wire n3505;
	wire n3506;
	wire n3507;
	wire n3508;
	wire n3509;
	wire n3510;
	wire n3511;
	wire n3512;
	wire n3513;
	wire n3514;
	wire n3515;
	wire n3516;
	wire n3517;
	wire n3518;
	wire n3519;
	wire n3520;
	wire n3521;
	wire n3522;
	wire n3523;
	wire n3524;
	wire n3525;
	wire n3526;
	wire n3527;
	wire n3528;
	wire n3529;
	wire n3530;
	wire n3531;
	wire n3532;
	wire n3533;
	wire n3534;
	wire n3535;
	wire n3536;
	wire n3537;
	wire n3538;
	wire n3539;
	wire n3540;
	wire n3541;
	wire n3542;
	wire n3543;
	wire n3544;
	wire n3545;
	wire n3546;
	wire n3547;
	wire n3548;
	wire n3549;
	wire n3550;
	wire n3551;
	wire n3552;
	wire n3553;
	wire n3554;
	wire n3555;
	wire n3556;
	wire n3557;
	wire n3558;
	wire n3559;
	wire n3560;
	wire n3561;
	wire n3562;
	wire n3563;
	wire n3564;
	wire n3565;
	wire n3566;
	wire n3567;
	wire n3568;
	wire n3569;
	wire n3570;
	wire n3571;
	wire n3572;
	wire n3573;
	wire n3574;
	wire n3575;
	wire n3576;
	wire n3577;
	wire n3578;
	wire n3579;
	wire n3580;
	wire n3581;
	wire n3582;
	wire n3583;
	wire n3584;
	wire n3585;
	wire n3586;
	wire n3587;
	wire n3588;
	wire n3589;
	wire n3590;
	wire n3591;
	wire n3592;
	wire n3593;
	wire n3594;
	wire n3595;
	wire n3596;
	wire n3597;
	wire n3598;
	wire n3599;
	wire n3600;
	wire n3601;
	wire n3602;
	wire n3603;
	wire n3604;
	wire n3605;
	wire n3606;
	wire n3607;
	wire n3608;
	wire n3609;
	wire n3610;
	wire n3611;
	wire n3612;
	wire n3613;
	wire n3614;
	wire n3615;
	wire n3616;
	wire n3617;
	wire n3618;
	wire n3619;
	wire n3620;
	wire n3621;
	wire n3622;
	wire n3623;
	wire n3624;
	wire n3625;
	wire n3626;
	wire n3627;
	wire n3628;
	wire n3629;
	wire n3630;
	wire n3631;
	wire n3632;
	wire n3633;
	wire n3634;
	wire n3635;
	wire n3636;
	wire n3637;
	wire n3638;
	wire n3639;
	wire n3640;
	wire n3641;
	wire n3642;
	wire n3643;
	wire n3644;
	wire n3645;
	wire n3646;
	wire n3647;
	wire n3648;
	wire n3649;
	wire n3650;
	wire n3651;
	wire n3652;
	wire n3653;
	wire n3654;
	wire n3655;
	wire n3656;
	wire n3657;
	wire n3658;
	wire n3659;
	wire n3660;
	wire n3661;
	wire n3662;
	wire n3663;
	wire n3664;
	wire n3665;
	wire n3666;
	wire n3667;
	wire n3668;
	wire n3669;
	wire n3670;
	wire n3671;
	wire n3672;
	wire n3673;
	wire n3674;
	wire n3675;
	wire n3676;
	wire n3677;
	wire n3678;
	wire n3679;
	wire n3680;
	wire n3681;
	wire n3682;
	wire n3683;
	wire n3684;
	wire n3685;
	wire n3686;
	wire n3687;
	wire n3688;
	wire n3689;
	wire n3690;
	wire n3691;
	wire n3692;
	wire n3693;
	wire n3694;
	wire n3695;
	wire n3696;
	wire n3697;
	wire n3698;
	wire n3699;
	wire n3700;
	wire n3701;
	wire n3702;
	wire n3703;
	wire n3704;
	wire n3705;
	wire n3706;
	wire n3707;
	wire n3708;
	wire n3709;
	wire n3710;
	wire n3711;
	wire n3712;
	wire n3713;
	wire n3714;
	wire n3715;
	wire n3716;
	wire n3717;
	wire n3718;
	wire n3719;
	wire n3720;
	wire n3721;
	wire n3722;
	wire n3723;
	wire n3724;
	wire n3725;
	wire n3726;
	wire n3727;
	wire n3728;
	wire n3729;
	wire n3730;
	wire n3731;
	wire n3732;
	wire n3733;
	wire n3734;
	wire n3735;
	wire n3736;
	wire n3737;
	wire n3738;
	wire n3739;
	wire n3740;
	wire n3741;
	wire n3742;
	wire n3743;
	wire n3744;
	wire n3745;
	wire n3746;
	wire n3747;
	wire n3748;
	wire n3749;
	wire n3750;
	wire n3751;
	wire n3752;
	wire n3753;
	wire n3754;
	wire n3755;
	wire n3756;
	wire n3757;
	wire n3758;
	wire n3759;
	wire n3760;
	wire n3761;
	wire n3762;
	wire n3763;
	wire n3764;
	wire n3765;
	wire n3766;
	wire n3767;
	wire n3768;
	wire n3769;
	wire n3770;
	wire n3771;
	wire n3772;
	wire n3773;
	wire n3774;
	wire n3775;
	wire n3776;
	wire n3777;
	wire n3778;
	wire n3779;
	wire n3780;
	wire n3781;
	wire n3782;
	wire n3783;
	wire n3784;
	wire n3785;
	wire n3786;
	wire n3787;
	wire n3788;
	wire n3789;
	wire n3790;
	wire n3791;
	wire n3792;
	wire n3793;
	wire n3794;
	wire n3795;
	wire n3796;
	wire n3797;
	wire n3798;
	wire n3799;
	wire n3800;
	wire n3801;
	wire n3802;
	wire n3803;
	wire n3804;
	wire n3805;
	wire n3806;
	wire n3807;
	wire n3808;
	wire n3809;
	wire n3810;
	wire n3811;
	wire n3812;
	wire n3813;
	wire n3814;
	wire n3815;
	wire n3816;
	wire n3817;
	wire n3818;
	wire n3819;
	wire n3820;
	wire n3821;
	wire n3822;
	wire n3823;
	wire n3824;
	wire n3825;
	wire n3826;
	wire n3827;
	wire n3828;
	wire n3829;
	wire n3830;
	wire n3831;
	wire n3832;
	wire n3833;
	wire n3834;
	wire n3835;
	wire n3836;
	wire n3837;
	wire n3838;
	wire n3839;
	wire n3840;
	wire n3841;
	wire n3842;
	wire n3843;
	wire n3844;
	wire n3845;
	wire n3846;
	wire n3847;
	wire n3848;
	wire n3849;
	wire n3850;
	wire n3851;
	wire n3852;
	wire n3853;
	wire n3854;
	wire n3855;
	wire n3856;
	wire n3857;
	wire n3858;
	wire n3859;
	wire n3860;
	wire n3861;
	wire n3862;
	wire n3863;
	wire n3864;
	wire n3865;
	wire n3866;
	wire n3867;
	wire n3868;
	wire n3869;
	wire n3870;
	wire n3871;
	wire n3872;
	wire n3873;
	wire n3874;
	wire n3875;
	wire n3876;
	wire n3877;
	wire n3878;
	wire n3879;
	wire n3880;
	wire n3881;
	wire n3882;
	wire n3883;
	wire n3884;
	wire n3885;
	wire n3886;
	wire n3887;
	wire n3888;
	wire n3889;
	wire n3890;
	wire n3891;
	wire n3893;
	wire n3894;
	wire n3895;
	wire n3896;
	wire n3897;
	wire n3898;
	wire n3899;
	wire n3900;
	wire n3901;
	wire n3902;
	wire n3904;
	wire n3905;
	wire n3906;
	wire n3907;
	wire n3908;
	wire n3909;
	wire n3910;
	wire n3911;
	wire n3912;
	wire n3913;
	wire n3914;
	wire n3915;
	wire n3916;
	wire n3917;
	wire n3918;
	wire n3919;
	wire n3920;
	wire n3923;
	wire n3924;
	wire n3925;
	wire n3926;
	wire n3927;
	wire n3928;
	wire n3929;
	wire n3930;
	wire n3931;
	wire n3932;
	wire n3933;
	wire n3934;
	wire n3935;
	wire n3936;
	wire n3937;
	wire n3938;
	wire n3939;
	wire n3940;
	wire n3941;
	wire n3942;
	wire n3943;
	wire n3944;
	wire n3945;
	wire n3946;
	wire n3947;
	wire n3948;
	wire n3949;
	wire n3950;
	wire n3951;
	wire n3952;
	wire n3953;
	wire n3954;
	wire n3955;
	wire n3956;
	wire n3957;
	wire n3958;
	wire n3959;
	wire n3960;
	wire n3961;
	wire n3962;
	wire n3963;
	wire n3964;
	wire n3965;
	wire n3966;
	wire n3967;
	wire n3968;
	wire n3969;
	wire n3970;
	wire n3971;
	wire n3972;
	wire n3973;
	wire n3974;
	wire n3975;
	wire n3976;
	wire n3977;
	wire n3978;
	wire n3979;
	wire n3980;
	wire n3981;
	wire n3982;
	wire n3983;
	wire n3984;
	wire n3985;
	wire n3986;
	wire n3987;
	wire n3988;
	wire n3989;
	wire n3990;
	wire n3991;
	wire n3992;
	wire n3993;
	wire n3994;
	wire n3995;
	wire n3996;
	wire n3997;
	wire n3998;
	wire n3999;
	wire n4000;
	wire n4001;
	wire n4002;
	wire n4003;
	wire n4004;
	wire n4005;
	wire n4006;
	wire n4007;
	wire n4008;
	wire n4009;
	wire n4010;
	wire n4011;
	wire n4012;
	wire n4013;
	wire n4014;
	wire n4015;
	wire n4016;
	wire n4017;
	wire n4018;
	wire n4019;
	wire n4021;
	wire n4022;
	wire n4023;
	wire n4024;
	wire n4025;
	wire n4026;
	wire n4027;
	wire n4028;
	wire n4029;
	wire n4030;
	wire n4031;
	wire n4032;
	wire n4033;
	wire n4034;
	wire n4035;
	wire n4036;
	wire n4037;
	wire n4038;
	wire n4039;
	wire n4040;
	wire n4041;
	wire n4042;
	wire n4043;
	wire n4044;
	wire n4045;
	wire n4046;
	wire n4047;
	wire n4048;
	wire n4049;
	wire n4050;
	wire n4051;
	wire n4052;
	wire n4053;
	wire n4054;
	wire n4055;
	wire n4056;
	wire n4057;
	wire n4058;
	wire n4059;
	wire n4060;
	wire n4061;
	wire n4062;
	wire n4063;
	wire n4064;
	wire n4065;
	wire n4066;
	wire n4067;
	wire n4068;
	wire n4069;
	wire n4070;
	wire n4071;
	wire n4072;
	wire n4073;
	wire n4074;
	wire n4075;
	wire n4076;
	wire n4077;
	wire n4078;
	wire n4079;
	wire n4080;
	wire n4081;
	wire n4082;
	wire n4083;
	wire n4084;
	wire n4085;
	wire n4086;
	wire n4087;
	wire n4088;
	wire n4089;
	wire n4090;
	wire n4091;
	wire n4092;
	wire n4093;
	wire n4094;
	wire n4095;
	wire n4096;
	wire n4097;
	wire n4098;
	wire n4099;
	wire n4100;
	wire n4101;
	wire n4102;
	wire n4103;
	wire n4104;
	wire n4105;
	wire n4106;
	wire n4107;
	wire n4108;
	wire n4109;
	wire n4110;
	wire n4111;
	wire n4112;
	wire n4113;
	wire n4114;
	wire n4115;
	wire n4116;
	wire n4117;
	wire n4118;
	wire n4119;
	wire n4120;
	wire n4121;
	wire n4123;
	wire n4124;
	wire n4125;
	wire n4126;
	wire n4127;
	wire n4128;
	wire n4129;
	wire n4130;
	wire n4131;
	wire n4132;
	wire n4133;
	wire n4134;
	wire n4135;
	wire n4136;
	wire n4137;
	wire n4138;
	wire n4139;
	wire n4140;
	wire n4141;
	wire n4142;
	wire n4143;
	wire n4144;
	wire n4145;
	wire n4146;
	wire n4147;
	wire n4148;
	wire n4149;
	wire n4150;
	wire n4151;
	wire n4152;
	wire n4153;
	wire n4154;
	wire n4155;
	wire n4156;
	wire n4157;
	wire n4158;
	wire n4159;
	wire n4160;
	wire n4161;
	wire n4162;
	wire n4163;
	wire n4164;
	wire n4165;
	wire n4166;
	wire n4167;
	wire n4168;
	wire n4169;
	wire n4170;
	wire n4171;
	wire n4172;
	wire n4173;
	wire n4174;
	wire n4175;
	wire n4176;
	wire n4177;
	wire n4178;
	wire n4179;
	wire n4180;
	wire n4181;
	wire n4182;
	wire n4183;
	wire n4184;
	wire n4185;
	wire n4186;
	wire n4187;
	wire n4188;
	wire n4189;
	wire n4190;
	wire n4191;
	wire n4192;
	wire n4193;
	wire n4194;
	wire n4195;
	wire n4196;
	wire n4197;
	wire n4198;
	wire n4199;
	wire n4200;
	wire n4201;
	wire n4202;
	wire n4203;
	wire n4204;
	wire n4205;
	wire n4206;
	wire n4207;
	wire n4208;
	wire n4209;
	wire n4211;
	wire n4212;
	wire n4213;
	wire n4214;
	wire n4215;
	wire n4216;
	wire n4217;
	wire n4218;
	wire n4219;
	wire n4220;
	wire n4221;
	wire n4222;
	wire n4223;
	wire n4224;
	wire n4225;
	wire n4226;
	wire n4227;
	wire n4228;
	wire n4229;
	wire n4230;
	wire n4231;
	wire n4232;
	wire n4233;
	wire n4234;
	wire n4235;
	wire n4236;
	wire n4237;
	wire n4238;
	wire n4239;
	wire n4240;
	wire n4241;
	wire n4242;
	wire n4243;
	wire n4244;
	wire n4245;
	wire n4246;
	wire n4247;
	wire n4248;
	wire n4249;
	wire n4250;
	wire n4251;
	wire n4252;
	wire n4253;
	wire n4254;
	wire n4255;
	wire n4256;
	wire n4257;
	wire n4258;
	wire n4259;
	wire n4260;
	wire n4261;
	wire n4262;
	wire n4263;
	wire n4264;
	wire n4265;
	wire n4266;
	wire n4267;
	wire n4268;
	wire n4269;
	wire n4270;
	wire n4271;
	wire n4272;
	wire n4273;
	wire n4274;
	wire n4275;
	wire n4276;
	wire n4277;
	wire n4278;
	wire n4279;
	wire n4280;
	wire n4281;
	wire n4282;
	wire n4283;
	wire n4284;
	wire n4285;
	wire n4286;
	wire n4287;
	wire n4288;
	wire n4289;
	wire n4290;
	wire n4291;
	wire n4293;
	wire n4294;
	wire n4295;
	wire n4296;
	wire n4297;
	wire n4298;
	wire n4299;
	wire n4300;
	wire n4301;
	wire n4302;
	wire n4303;
	wire n4304;
	wire n4305;
	wire n4306;
	wire n4307;
	wire n4308;
	wire n4309;
	wire n4310;
	wire n4311;
	wire n4312;
	wire n4313;
	wire n4314;
	wire n4315;
	wire n4316;
	wire n4317;
	wire n4318;
	wire n4319;
	wire n4320;
	wire n4321;
	wire n4322;
	wire n4323;
	wire n4324;
	wire n4325;
	wire n4326;
	wire n4327;
	wire n4328;
	wire n4329;
	wire n4330;
	wire n4331;
	wire n4332;
	wire n4333;
	wire n4334;
	wire n4335;
	wire n4336;
	wire n4337;
	wire n4338;
	wire n4339;
	wire n4340;
	wire n4341;
	wire n4342;
	wire n4343;
	wire n4344;
	wire n4345;
	wire n4346;
	wire n4347;
	wire n4348;
	wire n4349;
	wire n4350;
	wire n4351;
	wire n4352;
	wire n4353;
	wire n4354;
	wire n4355;
	wire n4356;
	wire n4357;
	wire n4358;
	wire n4359;
	wire n4360;
	wire n4361;
	wire n4362;
	wire n4363;
	wire n4364;
	wire n4365;
	wire n4366;
	wire n4367;
	wire n4368;
	wire n4369;
	wire n4370;
	wire n4371;
	wire n4372;
	wire n4373;
	wire n4375;
	wire n4376;
	wire n4377;
	wire n4378;
	wire n4379;
	wire n4380;
	wire n4381;
	wire n4382;
	wire n4383;
	wire n4384;
	wire n4385;
	wire n4386;
	wire n4387;
	wire n4388;
	wire n4389;
	wire n4390;
	wire n4391;
	wire n4392;
	wire n4393;
	wire n4394;
	wire n4395;
	wire n4396;
	wire n4397;
	wire n4398;
	wire n4399;
	wire n4400;
	wire n4401;
	wire n4402;
	wire n4403;
	wire n4404;
	wire n4405;
	wire n4406;
	wire n4407;
	wire n4408;
	wire n4409;
	wire n4410;
	wire n4411;
	wire n4412;
	wire n4413;
	wire n4414;
	wire n4415;
	wire n4416;
	wire n4417;
	wire n4418;
	wire n4419;
	wire n4420;
	wire n4421;
	wire n4422;
	wire n4423;
	wire n4424;
	wire n4425;
	wire n4426;
	wire n4427;
	wire n4428;
	wire n4429;
	wire n4430;
	wire n4431;
	wire n4432;
	wire n4433;
	wire n4434;
	wire n4435;
	wire n4436;
	wire n4437;
	wire n4438;
	wire n4439;
	wire n4440;
	wire n4441;
	wire n4442;
	wire n4443;
	wire n4444;
	wire n4445;
	wire n4446;
	wire n4447;
	wire n4448;
	wire n4449;
	wire n4450;
	wire n4451;
	wire n4452;
	wire n4453;
	wire n4454;
	wire n4455;
	wire n4457;
	wire n4458;
	wire n4459;
	wire n4460;
	wire n4461;
	wire n4462;
	wire n4463;
	wire n4464;
	wire n4465;
	wire n4466;
	wire n4467;
	wire n4468;
	wire n4469;
	wire n4470;
	wire n4471;
	wire n4472;
	wire n4473;
	wire n4474;
	wire n4475;
	wire n4476;
	wire n4477;
	wire n4478;
	wire n4479;
	wire n4480;
	wire n4481;
	wire n4482;
	wire n4483;
	wire n4484;
	wire n4485;
	wire n4486;
	wire n4487;
	wire n4488;
	wire n4489;
	wire n4490;
	wire n4491;
	wire n4492;
	wire n4493;
	wire n4494;
	wire n4495;
	wire n4496;
	wire n4497;
	wire n4498;
	wire n4499;
	wire n4500;
	wire n4501;
	wire n4502;
	wire n4503;
	wire n4504;
	wire n4505;
	wire n4506;
	wire n4507;
	wire n4508;
	wire n4509;
	wire n4510;
	wire n4511;
	wire n4512;
	wire n4513;
	wire n4514;
	wire n4515;
	wire n4516;
	wire n4517;
	wire n4518;
	wire n4519;
	wire n4520;
	wire n4521;
	wire n4522;
	wire n4523;
	wire n4524;
	wire n4525;
	wire n4526;
	wire n4527;
	wire n4528;
	wire n4530;
	wire n4531;
	wire n4532;
	wire n4533;
	wire n4534;
	wire n4535;
	wire n4536;
	wire n4537;
	wire n4538;
	wire n4539;
	wire n4540;
	wire n4541;
	wire n4542;
	wire n4543;
	wire n4544;
	wire n4545;
	wire n4546;
	wire n4547;
	wire n4548;
	wire n4549;
	wire n4550;
	wire n4551;
	wire n4552;
	wire n4553;
	wire n4554;
	wire n4555;
	wire n4556;
	wire n4557;
	wire n4558;
	wire n4559;
	wire n4560;
	wire n4561;
	wire n4562;
	wire n4563;
	wire n4564;
	wire n4565;
	wire n4566;
	wire n4567;
	wire n4568;
	wire n4569;
	wire n4570;
	wire n4571;
	wire n4572;
	wire n4573;
	wire n4574;
	wire n4575;
	wire n4576;
	wire n4577;
	wire n4578;
	wire n4579;
	wire n4580;
	wire n4581;
	wire n4582;
	wire n4583;
	wire n4584;
	wire n4585;
	wire n4586;
	wire n4587;
	wire n4588;
	wire n4589;
	wire n4590;
	wire n4591;
	wire n4592;
	wire n4593;
	wire n4594;
	wire n4595;
	wire n4596;
	wire n4597;
	wire n4598;
	wire n4599;
	wire n4600;
	wire n4601;
	wire n4602;
	wire n4603;
	wire n4604;
	wire n4606;
	wire n4607;
	wire n4608;
	wire n4609;
	wire n4610;
	wire n4611;
	wire n4612;
	wire n4613;
	wire n4614;
	wire n4615;
	wire n4616;
	wire n4617;
	wire n4618;
	wire n4619;
	wire n4620;
	wire n4621;
	wire n4622;
	wire n4623;
	wire n4624;
	wire n4625;
	wire n4626;
	wire n4627;
	wire n4628;
	wire n4629;
	wire n4630;
	wire n4631;
	wire n4632;
	wire n4633;
	wire n4634;
	wire n4635;
	wire n4636;
	wire n4637;
	wire n4638;
	wire n4639;
	wire n4640;
	wire n4641;
	wire n4642;
	wire n4643;
	wire n4644;
	wire n4645;
	wire n4646;
	wire n4647;
	wire n4648;
	wire n4649;
	wire n4650;
	wire n4651;
	wire n4652;
	wire n4653;
	wire n4654;
	wire n4655;
	wire n4656;
	wire n4657;
	wire n4658;
	wire n4659;
	wire n4660;
	wire n4661;
	wire n4662;
	wire n4663;
	wire n4664;
	wire n4665;
	wire n4666;
	wire n4667;
	wire n4668;
	wire n4670;
	wire n4671;
	wire n4672;
	wire n4673;
	wire n4674;
	wire n4675;
	wire n4676;
	wire n4677;
	wire n4678;
	wire n4679;
	wire n4680;
	wire n4681;
	wire n4682;
	wire n4683;
	wire n4684;
	wire n4685;
	wire n4686;
	wire n4687;
	wire n4688;
	wire n4689;
	wire n4690;
	wire n4691;
	wire n4692;
	wire n4693;
	wire n4694;
	wire n4695;
	wire n4696;
	wire n4697;
	wire n4698;
	wire n4699;
	wire n4700;
	wire n4701;
	wire n4702;
	wire n4703;
	wire n4704;
	wire n4705;
	wire n4706;
	wire n4707;
	wire n4708;
	wire n4709;
	wire n4710;
	wire n4711;
	wire n4712;
	wire n4713;
	wire n4714;
	wire n4715;
	wire n4716;
	wire n4717;
	wire n4718;
	wire n4719;
	wire n4720;
	wire n4721;
	wire n4722;
	wire n4723;
	wire n4724;
	wire n4725;
	wire n4726;
	wire n4727;
	wire n4728;
	wire n4729;
	wire n4730;
	wire n4731;
	wire n4732;
	wire n4733;
	wire n4735;
	wire n4736;
	wire n4737;
	wire n4738;
	wire n4739;
	wire n4740;
	wire n4741;
	wire n4742;
	wire n4743;
	wire n4744;
	wire n4745;
	wire n4746;
	wire n4747;
	wire n4748;
	wire n4749;
	wire n4750;
	wire n4751;
	wire n4752;
	wire n4753;
	wire n4754;
	wire n4755;
	wire n4756;
	wire n4757;
	wire n4758;
	wire n4759;
	wire n4760;
	wire n4761;
	wire n4762;
	wire n4763;
	wire n4764;
	wire n4765;
	wire n4766;
	wire n4767;
	wire n4768;
	wire n4769;
	wire n4770;
	wire n4771;
	wire n4772;
	wire n4773;
	wire n4774;
	wire n4775;
	wire n4776;
	wire n4777;
	wire n4778;
	wire n4779;
	wire n4780;
	wire n4781;
	wire n4782;
	wire n4783;
	wire n4784;
	wire n4785;
	wire n4786;
	wire n4787;
	wire n4788;
	wire n4789;
	wire n4790;
	wire n4792;
	wire n4793;
	wire n4794;
	wire n4795;
	wire n4796;
	wire n4797;
	wire n4798;
	wire n4799;
	wire n4800;
	wire n4801;
	wire n4802;
	wire n4803;
	wire n4804;
	wire n4805;
	wire n4806;
	wire n4807;
	wire n4808;
	wire n4809;
	wire n4810;
	wire n4811;
	wire n4812;
	wire n4813;
	wire n4814;
	wire n4815;
	wire n4816;
	wire n4817;
	wire n4818;
	wire n4819;
	wire n4820;
	wire n4821;
	wire n4822;
	wire n4823;
	wire n4824;
	wire n4825;
	wire n4826;
	wire n4827;
	wire n4828;
	wire n4829;
	wire n4830;
	wire n4831;
	wire n4832;
	wire n4833;
	wire n4834;
	wire n4835;
	wire n4836;
	wire n4837;
	wire n4838;
	wire n4839;
	wire n4840;
	wire n4841;
	wire n4843;
	wire n4844;
	wire n4845;
	wire n4846;
	wire n4847;
	wire n4848;
	wire n4849;
	wire n4850;
	wire n4851;
	wire n4852;
	wire n4853;
	wire n4854;
	wire n4855;
	wire n4856;
	wire n4857;
	wire n4858;
	wire n4859;
	wire n4860;
	wire n4861;
	wire n4862;
	wire n4863;
	wire n4864;
	wire n4865;
	wire n4866;
	wire n4867;
	wire n4868;
	wire n4869;
	wire n4870;
	wire n4871;
	wire n4872;
	wire n4873;
	wire n4874;
	wire n4875;
	wire n4876;
	wire n4877;
	wire n4878;
	wire n4879;
	wire n4880;
	wire n4881;
	wire n4882;
	wire n4883;
	wire n4884;
	wire n4885;
	wire n4886;
	wire n4887;
	wire n4888;
	wire n4889;
	wire n4890;
	wire n4891;
	wire n4892;
	wire n4893;
	wire n4894;
	wire n4895;
	wire n4896;
	wire n4897;
	wire n4899;
	wire n4900;
	wire n4901;
	wire n4902;
	wire n4903;
	wire n4904;
	wire n4905;
	wire n4906;
	wire n4907;
	wire n4908;
	wire n4909;
	wire n4910;
	wire n4911;
	wire n4912;
	wire n4913;
	wire n4914;
	wire n4915;
	wire n4916;
	wire n4917;
	wire n4918;
	wire n4919;
	wire n4920;
	wire n4921;
	wire n4922;
	wire n4923;
	wire n4924;
	wire n4925;
	wire n4926;
	wire n4927;
	wire n4928;
	wire n4929;
	wire n4930;
	wire n4931;
	wire n4932;
	wire n4933;
	wire n4934;
	wire n4935;
	wire n4936;
	wire n4937;
	wire n4938;
	wire n4939;
	wire n4940;
	wire n4941;
	wire n4942;
	wire n4943;
	wire n4944;
	wire n4946;
	wire n4947;
	wire n4948;
	wire n4949;
	wire n4950;
	wire n4951;
	wire n4952;
	wire n4953;
	wire n4954;
	wire n4955;
	wire n4956;
	wire n4957;
	wire n4958;
	wire n4959;
	wire n4960;
	wire n4961;
	wire n4962;
	wire n4963;
	wire n4964;
	wire n4965;
	wire n4966;
	wire n4967;
	wire n4968;
	wire n4969;
	wire n4970;
	wire n4971;
	wire n4972;
	wire n4973;
	wire n4974;
	wire n4975;
	wire n4976;
	wire n4977;
	wire n4978;
	wire n4979;
	wire n4980;
	wire n4981;
	wire n4982;
	wire n4983;
	wire n4984;
	wire n4985;
	wire n4986;
	wire n4987;
	wire n4989;
	wire n4990;
	wire n4991;
	wire n4992;
	wire n4993;
	wire n4994;
	wire n4995;
	wire n4996;
	wire n4997;
	wire n4998;
	wire n4999;
	wire n5000;
	wire n5001;
	wire n5002;
	wire n5003;
	wire n5004;
	wire n5005;
	wire n5006;
	wire n5007;
	wire n5008;
	wire n5009;
	wire n5010;
	wire n5011;
	wire n5012;
	wire n5013;
	wire n5014;
	wire n5015;
	wire n5016;
	wire n5017;
	wire n5018;
	wire n5019;
	wire n5020;
	wire n5021;
	wire n5022;
	wire n5024;
	wire n5025;
	wire n5026;
	wire n5027;
	wire n5028;
	wire n5029;
	wire n5030;
	wire n5031;
	wire n5032;
	wire n5033;
	wire n5034;
	wire n5035;
	wire n5036;
	wire n5037;
	wire n5038;
	wire n5039;
	wire n5040;
	wire n5041;
	wire n5042;
	wire n5043;
	wire n5044;
	wire n5046;
	wire n5047;
	wire n5048;
	wire n5049;
	wire n5050;
	wire n5051;
	wire n5052;
	wire n5053;
	wire n5054;
	wire n5055;
	wire n5056;
	wire n5057;
	wire n5058;
	wire n5059;
	wire n5060;
	wire n5061;
	wire n5062;
	wire n5063;
	wire n5064;
	wire n5065;
	wire n5066;
	wire n5067;
	wire n5068;
	wire n5069;
	wire n5071;
	wire n5072;
	wire n5073;
	wire n5074;
	wire n5075;
	wire n5076;
	wire n5077;
	wire n5078;
	wire n5079;
	wire n5080;
	wire n5081;
	wire n5082;
	wire n5083;
	wire n5084;
	wire n5085;
	wire n5086;
	wire n5087;
	wire n5088;
	wire n5089;
	wire n5091;
	wire n5092;
	wire n5093;
	wire n5094;
	wire n5095;
	wire n5096;
	wire n5097;
	wire n5098;
	wire n5099;
	wire n5100;
	wire n5101;
	wire n5102;
	wire n5103;
	wire n5104;
	wire n5105;
	wire n5106;
	wire n5107;
	wire n5108;
	wire n5109;
	wire n5110;
	wire n5112;
	wire n5113;
	wire n5114;
	wire n5115;
	wire n5116;
	wire n5117;
	wire n5118;
	wire n5119;
	wire n5120;
	wire n5121;
	wire n5122;
	wire n5123;
	wire n5124;
	wire n5126;
	wire n5127;
	wire n5128;
	wire n5129;
	wire n5130;
	wire n5131;
	wire n5132;
	wire n5133;
	wire n5135;
	wire n5136;
	wire n5137;
	wire n5138;
	wire n5139;
	wire n5140;
	wire n5141;
	wire n5142;
	wire n5143;
	wire n5144;
	wire n5145;
	wire n5146;
	wire n5147;
	wire n5148;
	wire n5149;
	wire n5151;
	wire n5153;
	wire n5154;
	wire n5155;
	wire n5156;
	wire n5157;
	wire n5158;
	wire n5159;
	wire n5160;
	wire[2:0] w_a0_0;
	wire[1:0] w_a0_1;
	wire[2:0] w_a1_0;
	wire[2:0] w_a2_0;
	wire[2:0] w_a2_1;
	wire[2:0] w_a3_0;
	wire[2:0] w_a4_0;
	wire[1:0] w_a4_1;
	wire[2:0] w_a5_0;
	wire[2:0] w_a6_0;
	wire[1:0] w_a6_1;
	wire[2:0] w_a7_0;
	wire[2:0] w_a8_0;
	wire[1:0] w_a8_1;
	wire[2:0] w_a9_0;
	wire[2:0] w_a10_0;
	wire[1:0] w_a10_1;
	wire[2:0] w_a11_0;
	wire[2:0] w_a12_0;
	wire[1:0] w_a12_1;
	wire[2:0] w_a13_0;
	wire[2:0] w_a14_0;
	wire[1:0] w_a14_1;
	wire[2:0] w_a15_0;
	wire[1:0] w_a15_1;
	wire[2:0] w_a16_0;
	wire[1:0] w_a17_0;
	wire[2:0] w_a18_0;
	wire[1:0] w_a18_1;
	wire[2:0] w_a19_0;
	wire[2:0] w_a20_0;
	wire[1:0] w_a20_1;
	wire[1:0] w_a21_0;
	wire[2:0] w_a22_0;
	wire[2:0] w_a22_1;
	wire[2:0] w_a22_2;
	wire[2:0] w_a22_3;
	wire[2:0] w_a22_4;
	wire[2:0] w_a22_5;
	wire[1:0] w_a22_6;
	wire[1:0] w_sin0_0;
	wire sin0_fa_;
	wire[2:0] w_n49_0;
	wire[2:0] w_n49_1;
	wire[2:0] w_n49_2;
	wire[2:0] w_n49_3;
	wire[2:0] w_n49_4;
	wire[1:0] w_n49_5;
	wire[1:0] w_n51_0;
	wire[1:0] w_n52_0;
	wire[1:0] w_n53_0;
	wire[1:0] w_n54_0;
	wire[2:0] w_n55_0;
	wire[2:0] w_n55_1;
	wire[2:0] w_n55_2;
	wire[2:0] w_n55_3;
	wire[2:0] w_n55_4;
	wire[2:0] w_n55_5;
	wire[2:0] w_n55_6;
	wire[2:0] w_n55_7;
	wire[2:0] w_n55_8;
	wire[2:0] w_n55_9;
	wire[2:0] w_n56_0;
	wire[2:0] w_n56_1;
	wire[2:0] w_n56_2;
	wire[2:0] w_n56_3;
	wire[2:0] w_n56_4;
	wire[2:0] w_n56_5;
	wire[2:0] w_n56_6;
	wire[2:0] w_n56_7;
	wire[2:0] w_n56_8;
	wire[2:0] w_n56_9;
	wire[2:0] w_n56_10;
	wire[2:0] w_n56_11;
	wire[2:0] w_n56_12;
	wire[1:0] w_n57_0;
	wire[2:0] w_n58_0;
	wire[2:0] w_n58_1;
	wire[2:0] w_n58_2;
	wire[2:0] w_n58_3;
	wire[2:0] w_n58_4;
	wire[2:0] w_n59_0;
	wire[2:0] w_n59_1;
	wire[2:0] w_n59_2;
	wire[1:0] w_n59_3;
	wire[2:0] w_n61_0;
	wire[2:0] w_n61_1;
	wire[2:0] w_n62_0;
	wire[2:0] w_n63_0;
	wire[2:0] w_n63_1;
	wire[2:0] w_n63_2;
	wire[1:0] w_n64_0;
	wire[2:0] w_n68_0;
	wire[2:0] w_n68_1;
	wire[2:0] w_n68_2;
	wire[2:0] w_n68_3;
	wire[2:0] w_n68_4;
	wire[2:0] w_n68_5;
	wire[2:0] w_n68_6;
	wire[2:0] w_n69_0;
	wire[2:0] w_n70_0;
	wire[2:0] w_n75_0;
	wire[2:0] w_n75_1;
	wire[2:0] w_n75_2;
	wire[2:0] w_n75_3;
	wire[2:0] w_n75_4;
	wire[2:0] w_n75_5;
	wire[1:0] w_n76_0;
	wire[1:0] w_n77_0;
	wire[2:0] w_n78_0;
	wire[2:0] w_n78_1;
	wire[2:0] w_n78_2;
	wire[2:0] w_n79_0;
	wire[2:0] w_n79_1;
	wire[2:0] w_n79_2;
	wire[2:0] w_n79_3;
	wire[2:0] w_n79_4;
	wire[2:0] w_n79_5;
	wire[1:0] w_n79_6;
	wire[1:0] w_n81_0;
	wire[1:0] w_n82_0;
	wire[1:0] w_n83_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n85_0;
	wire[1:0] w_n86_0;
	wire[1:0] w_n87_0;
	wire[1:0] w_n88_0;
	wire[1:0] w_n89_0;
	wire[1:0] w_n90_0;
	wire[1:0] w_n91_0;
	wire[1:0] w_n92_0;
	wire[2:0] w_n96_0;
	wire[2:0] w_n96_1;
	wire[2:0] w_n96_2;
	wire[2:0] w_n96_3;
	wire[2:0] w_n96_4;
	wire[2:0] w_n96_5;
	wire[1:0] w_n97_0;
	wire[1:0] w_n98_0;
	wire[1:0] w_n99_0;
	wire[1:0] w_n100_0;
	wire[1:0] w_n102_0;
	wire[2:0] w_n103_0;
	wire[1:0] w_n103_1;
	wire[1:0] w_n104_0;
	wire[1:0] w_n105_0;
	wire[2:0] w_n108_0;
	wire[1:0] w_n108_1;
	wire[2:0] w_n109_0;
	wire[2:0] w_n109_1;
	wire[1:0] w_n109_2;
	wire[2:0] w_n110_0;
	wire[2:0] w_n110_1;
	wire[2:0] w_n110_2;
	wire[2:0] w_n110_3;
	wire[2:0] w_n110_4;
	wire[2:0] w_n110_5;
	wire[1:0] w_n110_6;
	wire[1:0] w_n112_0;
	wire[2:0] w_n116_0;
	wire[1:0] w_n116_1;
	wire[1:0] w_n117_0;
	wire[2:0] w_n118_0;
	wire[1:0] w_n119_0;
	wire[2:0] w_n120_0;
	wire[1:0] w_n121_0;
	wire[2:0] w_n123_0;
	wire[1:0] w_n123_1;
	wire[1:0] w_n125_0;
	wire[2:0] w_n126_0;
	wire[2:0] w_n127_0;
	wire[1:0] w_n127_1;
	wire[2:0] w_n128_0;
	wire[2:0] w_n128_1;
	wire[2:0] w_n128_2;
	wire[2:0] w_n130_0;
	wire[2:0] w_n130_1;
	wire[2:0] w_n130_2;
	wire[1:0] w_n131_0;
	wire[2:0] w_n132_0;
	wire[2:0] w_n134_0;
	wire[1:0] w_n134_1;
	wire[2:0] w_n135_0;
	wire[2:0] w_n135_1;
	wire[2:0] w_n135_2;
	wire[2:0] w_n136_0;
	wire[1:0] w_n137_0;
	wire[2:0] w_n138_0;
	wire[2:0] w_n138_1;
	wire[2:0] w_n138_2;
	wire[2:0] w_n138_3;
	wire[1:0] w_n138_4;
	wire[2:0] w_n139_0;
	wire[1:0] w_n139_1;
	wire[2:0] w_n140_0;
	wire[1:0] w_n140_1;
	wire[2:0] w_n141_0;
	wire[2:0] w_n141_1;
	wire[1:0] w_n141_2;
	wire[2:0] w_n142_0;
	wire[1:0] w_n142_1;
	wire[2:0] w_n143_0;
	wire[2:0] w_n143_1;
	wire[2:0] w_n143_2;
	wire[2:0] w_n143_3;
	wire[2:0] w_n143_4;
	wire[2:0] w_n143_5;
	wire[1:0] w_n143_6;
	wire[2:0] w_n144_0;
	wire[2:0] w_n145_0;
	wire[1:0] w_n145_1;
	wire[2:0] w_n146_0;
	wire[2:0] w_n146_1;
	wire[2:0] w_n146_2;
	wire[2:0] w_n146_3;
	wire[2:0] w_n146_4;
	wire[2:0] w_n147_0;
	wire[2:0] w_n147_1;
	wire[2:0] w_n147_2;
	wire[2:0] w_n147_3;
	wire[1:0] w_n147_4;
	wire[2:0] w_n151_0;
	wire[2:0] w_n151_1;
	wire[2:0] w_n151_2;
	wire[2:0] w_n151_3;
	wire[2:0] w_n151_4;
	wire[2:0] w_n151_5;
	wire[1:0] w_n151_6;
	wire[1:0] w_n152_0;
	wire[2:0] w_n153_0;
	wire[1:0] w_n153_1;
	wire[2:0] w_n154_0;
	wire[1:0] w_n154_1;
	wire[2:0] w_n155_0;
	wire[1:0] w_n155_1;
	wire[1:0] w_n156_0;
	wire[2:0] w_n157_0;
	wire[2:0] w_n157_1;
	wire[2:0] w_n158_0;
	wire[1:0] w_n158_1;
	wire[2:0] w_n160_0;
	wire[2:0] w_n161_0;
	wire[2:0] w_n162_0;
	wire[1:0] w_n162_1;
	wire[2:0] w_n163_0;
	wire[2:0] w_n163_1;
	wire[2:0] w_n163_2;
	wire[2:0] w_n164_0;
	wire[1:0] w_n165_0;
	wire[1:0] w_n167_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n207_0;
	wire[1:0] w_n210_0;
	wire[2:0] w_n211_0;
	wire[1:0] w_n211_1;
	wire[2:0] w_n212_0;
	wire[2:0] w_n212_1;
	wire[2:0] w_n212_2;
	wire[1:0] w_n212_3;
	wire[2:0] w_n213_0;
	wire[1:0] w_n213_1;
	wire[2:0] w_n214_0;
	wire[2:0] w_n214_1;
	wire[2:0] w_n214_2;
	wire[2:0] w_n215_0;
	wire[2:0] w_n215_1;
	wire[1:0] w_n215_2;
	wire[2:0] w_n216_0;
	wire[2:0] w_n216_1;
	wire[2:0] w_n216_2;
	wire[2:0] w_n216_3;
	wire[1:0] w_n216_4;
	wire[1:0] w_n218_0;
	wire[2:0] w_n219_0;
	wire[1:0] w_n219_1;
	wire[2:0] w_n220_0;
	wire[2:0] w_n220_1;
	wire[2:0] w_n220_2;
	wire[1:0] w_n220_3;
	wire[2:0] w_n222_0;
	wire[2:0] w_n222_1;
	wire[1:0] w_n222_2;
	wire[2:0] w_n223_0;
	wire[2:0] w_n223_1;
	wire[2:0] w_n223_2;
	wire[2:0] w_n224_0;
	wire[2:0] w_n225_0;
	wire[2:0] w_n225_1;
	wire[2:0] w_n225_2;
	wire[2:0] w_n227_0;
	wire[2:0] w_n227_1;
	wire[1:0] w_n227_2;
	wire[1:0] w_n228_0;
	wire[2:0] w_n229_0;
	wire[2:0] w_n229_1;
	wire[2:0] w_n229_2;
	wire[2:0] w_n230_0;
	wire[2:0] w_n230_1;
	wire[1:0] w_n230_2;
	wire[1:0] w_n231_0;
	wire[2:0] w_n232_0;
	wire[2:0] w_n232_1;
	wire[2:0] w_n232_2;
	wire[1:0] w_n234_0;
	wire[2:0] w_n235_0;
	wire[2:0] w_n236_0;
	wire[2:0] w_n236_1;
	wire[2:0] w_n236_2;
	wire[1:0] w_n236_3;
	wire[1:0] w_n239_0;
	wire[2:0] w_n240_0;
	wire[2:0] w_n241_0;
	wire[1:0] w_n241_1;
	wire[1:0] w_n242_0;
	wire[2:0] w_n243_0;
	wire[2:0] w_n243_1;
	wire[2:0] w_n243_2;
	wire[2:0] w_n243_3;
	wire[2:0] w_n243_4;
	wire[1:0] w_n246_0;
	wire[2:0] w_n247_0;
	wire[2:0] w_n247_1;
	wire[2:0] w_n247_2;
	wire[2:0] w_n249_0;
	wire[2:0] w_n249_1;
	wire[1:0] w_n249_2;
	wire[1:0] w_n250_0;
	wire[2:0] w_n251_0;
	wire[2:0] w_n251_1;
	wire[2:0] w_n251_2;
	wire[1:0] w_n251_3;
	wire[2:0] w_n254_0;
	wire[2:0] w_n254_1;
	wire[2:0] w_n254_2;
	wire[1:0] w_n254_3;
	wire[2:0] w_n256_0;
	wire[2:0] w_n256_1;
	wire[1:0] w_n256_2;
	wire[2:0] w_n259_0;
	wire[2:0] w_n259_1;
	wire[2:0] w_n259_2;
	wire[1:0] w_n259_3;
	wire[1:0] w_n260_0;
	wire[2:0] w_n261_0;
	wire[2:0] w_n261_1;
	wire[2:0] w_n262_0;
	wire[2:0] w_n262_1;
	wire[2:0] w_n262_2;
	wire[2:0] w_n262_3;
	wire[1:0] w_n263_0;
	wire[2:0] w_n264_0;
	wire[2:0] w_n264_1;
	wire[2:0] w_n264_2;
	wire[2:0] w_n265_0;
	wire[2:0] w_n266_0;
	wire[1:0] w_n266_1;
	wire[2:0] w_n267_0;
	wire[2:0] w_n267_1;
	wire[2:0] w_n268_0;
	wire[2:0] w_n268_1;
	wire[2:0] w_n268_2;
	wire[2:0] w_n269_0;
	wire[2:0] w_n270_0;
	wire[2:0] w_n270_1;
	wire[2:0] w_n270_2;
	wire[1:0] w_n275_0;
	wire[2:0] w_n276_0;
	wire[2:0] w_n277_0;
	wire[2:0] w_n277_1;
	wire[2:0] w_n277_2;
	wire[1:0] w_n277_3;
	wire[1:0] w_n278_0;
	wire[2:0] w_n279_0;
	wire[2:0] w_n279_1;
	wire[1:0] w_n279_2;
	wire[2:0] w_n280_0;
	wire[1:0] w_n280_1;
	wire[1:0] w_n281_0;
	wire[2:0] w_n282_0;
	wire[2:0] w_n282_1;
	wire[2:0] w_n282_2;
	wire[1:0] w_n282_3;
	wire[2:0] w_n283_0;
	wire[2:0] w_n283_1;
	wire[2:0] w_n283_2;
	wire[1:0] w_n283_3;
	wire[1:0] w_n284_0;
	wire[2:0] w_n285_0;
	wire[2:0] w_n285_1;
	wire[1:0] w_n285_2;
	wire[2:0] w_n286_0;
	wire[2:0] w_n286_1;
	wire[1:0] w_n287_0;
	wire[2:0] w_n288_0;
	wire[1:0] w_n288_1;
	wire[1:0] w_n290_0;
	wire[2:0] w_n291_0;
	wire[2:0] w_n291_1;
	wire[1:0] w_n291_2;
	wire[2:0] w_n294_0;
	wire[2:0] w_n294_1;
	wire[2:0] w_n294_2;
	wire[1:0] w_n294_3;
	wire[2:0] w_n295_0;
	wire[2:0] w_n295_1;
	wire[2:0] w_n295_2;
	wire[2:0] w_n295_3;
	wire[2:0] w_n298_0;
	wire[2:0] w_n299_0;
	wire[1:0] w_n300_0;
	wire[2:0] w_n301_0;
	wire[2:0] w_n301_1;
	wire[2:0] w_n301_2;
	wire[2:0] w_n303_0;
	wire[2:0] w_n303_1;
	wire[2:0] w_n303_2;
	wire[2:0] w_n303_3;
	wire[1:0] w_n303_4;
	wire[2:0] w_n304_0;
	wire[2:0] w_n304_1;
	wire[2:0] w_n304_2;
	wire[1:0] w_n304_3;
	wire[2:0] w_n305_0;
	wire[1:0] w_n308_0;
	wire[1:0] w_n309_0;
	wire[2:0] w_n310_0;
	wire[2:0] w_n310_1;
	wire[2:0] w_n312_0;
	wire[2:0] w_n312_1;
	wire[2:0] w_n312_2;
	wire[2:0] w_n312_3;
	wire[2:0] w_n314_0;
	wire[1:0] w_n314_1;
	wire[2:0] w_n315_0;
	wire[1:0] w_n319_0;
	wire[2:0] w_n320_0;
	wire[2:0] w_n321_0;
	wire[1:0] w_n321_1;
	wire[1:0] w_n322_0;
	wire[2:0] w_n323_0;
	wire[2:0] w_n323_1;
	wire[2:0] w_n323_2;
	wire[1:0] w_n323_3;
	wire[2:0] w_n324_0;
	wire[1:0] w_n324_1;
	wire[1:0] w_n325_0;
	wire[1:0] w_n326_0;
	wire[2:0] w_n327_0;
	wire[2:0] w_n327_1;
	wire[2:0] w_n327_2;
	wire[2:0] w_n328_0;
	wire[2:0] w_n334_0;
	wire[2:0] w_n334_1;
	wire[2:0] w_n335_0;
	wire[2:0] w_n335_1;
	wire[2:0] w_n335_2;
	wire[2:0] w_n335_3;
	wire[2:0] w_n335_4;
	wire[2:0] w_n335_5;
	wire[2:0] w_n335_6;
	wire[1:0] w_n336_0;
	wire[2:0] w_n337_0;
	wire[2:0] w_n337_1;
	wire[2:0] w_n337_2;
	wire[2:0] w_n337_3;
	wire[2:0] w_n337_4;
	wire[1:0] w_n337_5;
	wire[2:0] w_n338_0;
	wire[1:0] w_n338_1;
	wire[2:0] w_n339_0;
	wire[2:0] w_n340_0;
	wire[2:0] w_n340_1;
	wire[1:0] w_n340_2;
	wire[2:0] w_n341_0;
	wire[2:0] w_n341_1;
	wire[2:0] w_n341_2;
	wire[2:0] w_n341_3;
	wire[1:0] w_n341_4;
	wire[1:0] w_n342_0;
	wire[2:0] w_n343_0;
	wire[2:0] w_n343_1;
	wire[1:0] w_n343_2;
	wire[2:0] w_n345_0;
	wire[2:0] w_n346_0;
	wire[2:0] w_n346_1;
	wire[2:0] w_n346_2;
	wire[2:0] w_n346_3;
	wire[2:0] w_n346_4;
	wire[2:0] w_n346_5;
	wire[2:0] w_n346_6;
	wire[1:0] w_n346_7;
	wire[2:0] w_n348_0;
	wire[2:0] w_n348_1;
	wire[2:0] w_n348_2;
	wire[2:0] w_n349_0;
	wire[2:0] w_n349_1;
	wire[2:0] w_n349_2;
	wire[2:0] w_n349_3;
	wire[2:0] w_n349_4;
	wire[2:0] w_n349_5;
	wire[2:0] w_n349_6;
	wire[2:0] w_n351_0;
	wire[2:0] w_n351_1;
	wire[1:0] w_n351_2;
	wire[2:0] w_n353_0;
	wire[2:0] w_n354_0;
	wire[2:0] w_n354_1;
	wire[2:0] w_n354_2;
	wire[2:0] w_n354_3;
	wire[1:0] w_n354_4;
	wire[1:0] w_n355_0;
	wire[2:0] w_n356_0;
	wire[2:0] w_n356_1;
	wire[2:0] w_n358_0;
	wire[2:0] w_n358_1;
	wire[1:0] w_n358_2;
	wire[1:0] w_n361_0;
	wire[1:0] w_n362_0;
	wire[2:0] w_n363_0;
	wire[2:0] w_n363_1;
	wire[1:0] w_n363_2;
	wire[1:0] w_n364_0;
	wire[2:0] w_n365_0;
	wire[2:0] w_n365_1;
	wire[1:0] w_n366_0;
	wire[2:0] w_n367_0;
	wire[2:0] w_n367_1;
	wire[2:0] w_n367_2;
	wire[2:0] w_n368_0;
	wire[2:0] w_n368_1;
	wire[2:0] w_n368_2;
	wire[1:0] w_n369_0;
	wire[2:0] w_n370_0;
	wire[2:0] w_n370_1;
	wire[1:0] w_n370_2;
	wire[1:0] w_n371_0;
	wire[2:0] w_n372_0;
	wire[2:0] w_n372_1;
	wire[1:0] w_n373_0;
	wire[2:0] w_n374_0;
	wire[2:0] w_n374_1;
	wire[2:0] w_n374_2;
	wire[1:0] w_n378_0;
	wire[2:0] w_n379_0;
	wire[2:0] w_n379_1;
	wire[2:0] w_n380_0;
	wire[1:0] w_n380_1;
	wire[2:0] w_n381_0;
	wire[2:0] w_n381_1;
	wire[2:0] w_n381_2;
	wire[1:0] w_n382_0;
	wire[2:0] w_n383_0;
	wire[2:0] w_n383_1;
	wire[2:0] w_n383_2;
	wire[2:0] w_n384_0;
	wire[1:0] w_n384_1;
	wire[2:0] w_n385_0;
	wire[1:0] w_n385_1;
	wire[2:0] w_n386_0;
	wire[2:0] w_n387_0;
	wire[2:0] w_n387_1;
	wire[1:0] w_n388_0;
	wire[1:0] w_n389_0;
	wire[2:0] w_n390_0;
	wire[2:0] w_n390_1;
	wire[2:0] w_n392_0;
	wire[2:0] w_n395_0;
	wire[2:0] w_n397_0;
	wire[2:0] w_n397_1;
	wire[1:0] w_n398_0;
	wire[1:0] w_n399_0;
	wire[1:0] w_n400_0;
	wire[2:0] w_n401_0;
	wire[2:0] w_n401_1;
	wire[2:0] w_n401_2;
	wire[2:0] w_n402_0;
	wire[2:0] w_n402_1;
	wire[2:0] w_n402_2;
	wire[1:0] w_n402_3;
	wire[1:0] w_n403_0;
	wire[1:0] w_n405_0;
	wire[2:0] w_n406_0;
	wire[1:0] w_n406_1;
	wire[1:0] w_n407_0;
	wire[1:0] w_n408_0;
	wire[1:0] w_n409_0;
	wire[2:0] w_n410_0;
	wire[2:0] w_n410_1;
	wire[1:0] w_n411_0;
	wire[2:0] w_n412_0;
	wire[2:0] w_n412_1;
	wire[1:0] w_n412_2;
	wire[1:0] w_n413_0;
	wire[1:0] w_n414_0;
	wire[2:0] w_n415_0;
	wire[2:0] w_n417_0;
	wire[2:0] w_n417_1;
	wire[2:0] w_n420_0;
	wire[2:0] w_n420_1;
	wire[1:0] w_n420_2;
	wire[2:0] w_n421_0;
	wire[2:0] w_n421_1;
	wire[2:0] w_n421_2;
	wire[1:0] w_n421_3;
	wire[2:0] w_n422_0;
	wire[2:0] w_n422_1;
	wire[2:0] w_n422_2;
	wire[1:0] w_n424_0;
	wire[1:0] w_n425_0;
	wire[2:0] w_n426_0;
	wire[2:0] w_n426_1;
	wire[2:0] w_n426_2;
	wire[2:0] w_n426_3;
	wire[2:0] w_n427_0;
	wire[2:0] w_n427_1;
	wire[2:0] w_n427_2;
	wire[1:0] w_n427_3;
	wire[2:0] w_n428_0;
	wire[1:0] w_n429_0;
	wire[2:0] w_n430_0;
	wire[2:0] w_n430_1;
	wire[2:0] w_n430_2;
	wire[1:0] w_n434_0;
	wire[1:0] w_n435_0;
	wire[2:0] w_n436_0;
	wire[2:0] w_n436_1;
	wire[2:0] w_n436_2;
	wire[2:0] w_n437_0;
	wire[2:0] w_n437_1;
	wire[1:0] w_n437_2;
	wire[1:0] w_n439_0;
	wire[2:0] w_n440_0;
	wire[2:0] w_n441_0;
	wire[2:0] w_n441_1;
	wire[1:0] w_n443_0;
	wire[1:0] w_n444_0;
	wire[2:0] w_n445_0;
	wire[2:0] w_n445_1;
	wire[2:0] w_n445_2;
	wire[2:0] w_n451_0;
	wire[2:0] w_n451_1;
	wire[2:0] w_n451_2;
	wire[1:0] w_n451_3;
	wire[1:0] w_n453_0;
	wire[2:0] w_n454_0;
	wire[2:0] w_n454_1;
	wire[2:0] w_n454_2;
	wire[1:0] w_n457_0;
	wire[2:0] w_n458_0;
	wire[2:0] w_n458_1;
	wire[1:0] w_n459_0;
	wire[1:0] w_n460_0;
	wire[2:0] w_n461_0;
	wire[2:0] w_n461_1;
	wire[2:0] w_n461_2;
	wire[2:0] w_n463_0;
	wire[2:0] w_n463_1;
	wire[2:0] w_n463_2;
	wire[1:0] w_n463_3;
	wire[1:0] w_n466_0;
	wire[2:0] w_n467_0;
	wire[1:0] w_n467_1;
	wire[1:0] w_n468_0;
	wire[1:0] w_n469_0;
	wire[2:0] w_n470_0;
	wire[2:0] w_n470_1;
	wire[1:0] w_n471_0;
	wire[1:0] w_n472_0;
	wire[2:0] w_n473_0;
	wire[2:0] w_n473_1;
	wire[1:0] w_n473_2;
	wire[2:0] w_n475_0;
	wire[1:0] w_n475_1;
	wire[2:0] w_n477_0;
	wire[2:0] w_n477_1;
	wire[2:0] w_n477_2;
	wire[1:0] w_n478_0;
	wire[2:0] w_n479_0;
	wire[2:0] w_n479_1;
	wire[1:0] w_n479_2;
	wire[1:0] w_n482_0;
	wire[2:0] w_n486_0;
	wire[1:0] w_n486_1;
	wire[1:0] w_n487_0;
	wire[2:0] w_n488_0;
	wire[2:0] w_n488_1;
	wire[1:0] w_n490_0;
	wire[1:0] w_n491_0;
	wire[1:0] w_n493_0;
	wire[1:0] w_n494_0;
	wire[2:0] w_n497_0;
	wire[1:0] w_n497_1;
	wire[2:0] w_n499_0;
	wire[2:0] w_n499_1;
	wire[1:0] w_n500_0;
	wire[2:0] w_n501_0;
	wire[2:0] w_n501_1;
	wire[2:0] w_n501_2;
	wire[2:0] w_n504_0;
	wire[1:0] w_n505_0;
	wire[2:0] w_n506_0;
	wire[2:0] w_n506_1;
	wire[1:0] w_n506_2;
	wire[2:0] w_n507_0;
	wire[1:0] w_n507_1;
	wire[2:0] w_n509_0;
	wire[2:0] w_n511_0;
	wire[1:0] w_n511_1;
	wire[2:0] w_n513_0;
	wire[2:0] w_n515_0;
	wire[2:0] w_n515_1;
	wire[2:0] w_n515_2;
	wire[1:0] w_n516_0;
	wire[2:0] w_n518_0;
	wire[1:0] w_n519_0;
	wire[2:0] w_n521_0;
	wire[1:0] w_n522_0;
	wire[2:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n525_0;
	wire[1:0] w_n531_0;
	wire[2:0] w_n532_0;
	wire[2:0] w_n532_1;
	wire[2:0] w_n532_2;
	wire[1:0] w_n534_0;
	wire[2:0] w_n535_0;
	wire[1:0] w_n535_1;
	wire[2:0] w_n538_0;
	wire[1:0] w_n541_0;
	wire[2:0] w_n543_0;
	wire[1:0] w_n543_1;
	wire[1:0] w_n545_0;
	wire[1:0] w_n548_0;
	wire[1:0] w_n550_0;
	wire[2:0] w_n551_0;
	wire[2:0] w_n552_0;
	wire[2:0] w_n554_0;
	wire[1:0] w_n556_0;
	wire[1:0] w_n557_0;
	wire[1:0] w_n560_0;
	wire[2:0] w_n561_0;
	wire[2:0] w_n561_1;
	wire[1:0] w_n561_2;
	wire[1:0] w_n562_0;
	wire[2:0] w_n563_0;
	wire[1:0] w_n564_0;
	wire[2:0] w_n565_0;
	wire[1:0] w_n565_1;
	wire[2:0] w_n568_0;
	wire[2:0] w_n571_0;
	wire[2:0] w_n574_0;
	wire[1:0] w_n577_0;
	wire[1:0] w_n578_0;
	wire[2:0] w_n579_0;
	wire[2:0] w_n579_1;
	wire[2:0] w_n579_2;
	wire[1:0] w_n580_0;
	wire[1:0] w_n581_0;
	wire[1:0] w_n584_0;
	wire[1:0] w_n586_0;
	wire[1:0] w_n587_0;
	wire[2:0] w_n588_0;
	wire[1:0] w_n588_1;
	wire[1:0] w_n590_0;
	wire[1:0] w_n591_0;
	wire[2:0] w_n592_0;
	wire[2:0] w_n592_1;
	wire[2:0] w_n592_2;
	wire[1:0] w_n592_3;
	wire[1:0] w_n593_0;
	wire[2:0] w_n594_0;
	wire[2:0] w_n594_1;
	wire[2:0] w_n594_2;
	wire[2:0] w_n595_0;
	wire[2:0] w_n596_0;
	wire[2:0] w_n597_0;
	wire[2:0] w_n597_1;
	wire[1:0] w_n597_2;
	wire[1:0] w_n598_0;
	wire[2:0] w_n604_0;
	wire[1:0] w_n605_0;
	wire[2:0] w_n606_0;
	wire[2:0] w_n608_0;
	wire[2:0] w_n611_0;
	wire[1:0] w_n611_1;
	wire[2:0] w_n612_0;
	wire[2:0] w_n612_1;
	wire[2:0] w_n612_2;
	wire[2:0] w_n612_3;
	wire[2:0] w_n614_0;
	wire[2:0] w_n614_1;
	wire[2:0] w_n614_2;
	wire[2:0] w_n619_0;
	wire[2:0] w_n619_1;
	wire[2:0] w_n622_0;
	wire[2:0] w_n622_1;
	wire[1:0] w_n623_0;
	wire[2:0] w_n624_0;
	wire[2:0] w_n624_1;
	wire[2:0] w_n624_2;
	wire[1:0] w_n625_0;
	wire[2:0] w_n626_0;
	wire[1:0] w_n626_1;
	wire[1:0] w_n630_0;
	wire[2:0] w_n631_0;
	wire[2:0] w_n632_0;
	wire[2:0] w_n632_1;
	wire[1:0] w_n632_2;
	wire[1:0] w_n633_0;
	wire[1:0] w_n636_0;
	wire[1:0] w_n637_0;
	wire[2:0] w_n638_0;
	wire[1:0] w_n641_0;
	wire[2:0] w_n642_0;
	wire[2:0] w_n642_1;
	wire[1:0] w_n643_0;
	wire[1:0] w_n644_0;
	wire[2:0] w_n645_0;
	wire[2:0] w_n645_1;
	wire[1:0] w_n645_2;
	wire[2:0] w_n646_0;
	wire[1:0] w_n648_0;
	wire[1:0] w_n650_0;
	wire[1:0] w_n651_0;
	wire[1:0] w_n655_0;
	wire[1:0] w_n661_0;
	wire[2:0] w_n662_0;
	wire[2:0] w_n662_1;
	wire[2:0] w_n662_2;
	wire[2:0] w_n664_0;
	wire[2:0] w_n665_0;
	wire[2:0] w_n665_1;
	wire[2:0] w_n665_2;
	wire[1:0] w_n667_0;
	wire[2:0] w_n668_0;
	wire[2:0] w_n668_1;
	wire[2:0] w_n668_2;
	wire[1:0] w_n669_0;
	wire[2:0] w_n670_0;
	wire[2:0] w_n675_0;
	wire[2:0] w_n676_0;
	wire[1:0] w_n676_1;
	wire[2:0] w_n677_0;
	wire[1:0] w_n678_0;
	wire[2:0] w_n679_0;
	wire[2:0] w_n679_1;
	wire[1:0] w_n679_2;
	wire[2:0] w_n680_0;
	wire[1:0] w_n680_1;
	wire[1:0] w_n681_0;
	wire[1:0] w_n685_0;
	wire[2:0] w_n688_0;
	wire[1:0] w_n690_0;
	wire[2:0] w_n691_0;
	wire[2:0] w_n691_1;
	wire[1:0] w_n693_0;
	wire[1:0] w_n695_0;
	wire[2:0] w_n699_0;
	wire[2:0] w_n699_1;
	wire[2:0] w_n699_2;
	wire[2:0] w_n699_3;
	wire[2:0] w_n699_4;
	wire[2:0] w_n699_5;
	wire[2:0] w_n699_6;
	wire[2:0] w_n699_7;
	wire[2:0] w_n699_8;
	wire[2:0] w_n699_9;
	wire[2:0] w_n699_10;
	wire[2:0] w_n699_11;
	wire[2:0] w_n699_12;
	wire[2:0] w_n699_13;
	wire[1:0] w_n700_0;
	wire[1:0] w_n702_0;
	wire[1:0] w_n704_0;
	wire[2:0] w_n708_0;
	wire[2:0] w_n708_1;
	wire[2:0] w_n708_2;
	wire[2:0] w_n708_3;
	wire[2:0] w_n708_4;
	wire[2:0] w_n708_5;
	wire[1:0] w_n708_6;
	wire[2:0] w_n709_0;
	wire[1:0] w_n709_1;
	wire[2:0] w_n710_0;
	wire[2:0] w_n710_1;
	wire[2:0] w_n710_2;
	wire[1:0] w_n710_3;
	wire[1:0] w_n711_0;
	wire[2:0] w_n712_0;
	wire[1:0] w_n713_0;
	wire[2:0] w_n719_0;
	wire[1:0] w_n719_1;
	wire[1:0] w_n722_0;
	wire[2:0] w_n724_0;
	wire[2:0] w_n724_1;
	wire[2:0] w_n724_2;
	wire[1:0] w_n725_0;
	wire[1:0] w_n726_0;
	wire[1:0] w_n727_0;
	wire[1:0] w_n728_0;
	wire[2:0] w_n730_0;
	wire[1:0] w_n730_1;
	wire[2:0] w_n731_0;
	wire[2:0] w_n732_0;
	wire[2:0] w_n732_1;
	wire[2:0] w_n732_2;
	wire[1:0] w_n732_3;
	wire[2:0] w_n733_0;
	wire[1:0] w_n733_1;
	wire[2:0] w_n734_0;
	wire[2:0] w_n734_1;
	wire[1:0] w_n735_0;
	wire[2:0] w_n739_0;
	wire[1:0] w_n740_0;
	wire[2:0] w_n741_0;
	wire[1:0] w_n741_1;
	wire[1:0] w_n742_0;
	wire[2:0] w_n744_0;
	wire[2:0] w_n744_1;
	wire[2:0] w_n744_2;
	wire[2:0] w_n746_0;
	wire[2:0] w_n748_0;
	wire[1:0] w_n748_1;
	wire[2:0] w_n749_0;
	wire[1:0] w_n749_1;
	wire[1:0] w_n750_0;
	wire[2:0] w_n751_0;
	wire[2:0] w_n751_1;
	wire[1:0] w_n751_2;
	wire[1:0] w_n754_0;
	wire[1:0] w_n756_0;
	wire[1:0] w_n757_0;
	wire[1:0] w_n758_0;
	wire[2:0] w_n762_0;
	wire[2:0] w_n762_1;
	wire[1:0] w_n762_2;
	wire[2:0] w_n763_0;
	wire[2:0] w_n763_1;
	wire[1:0] w_n763_2;
	wire[2:0] w_n764_0;
	wire[2:0] w_n765_0;
	wire[2:0] w_n765_1;
	wire[1:0] w_n767_0;
	wire[2:0] w_n768_0;
	wire[2:0] w_n768_1;
	wire[2:0] w_n768_2;
	wire[2:0] w_n771_0;
	wire[2:0] w_n771_1;
	wire[1:0] w_n771_2;
	wire[2:0] w_n772_0;
	wire[2:0] w_n772_1;
	wire[2:0] w_n772_2;
	wire[1:0] w_n773_0;
	wire[1:0] w_n776_0;
	wire[1:0] w_n779_0;
	wire[1:0] w_n780_0;
	wire[2:0] w_n781_0;
	wire[2:0] w_n781_1;
	wire[1:0] w_n781_2;
	wire[1:0] w_n784_0;
	wire[2:0] w_n786_0;
	wire[1:0] w_n786_1;
	wire[2:0] w_n788_0;
	wire[2:0] w_n789_0;
	wire[2:0] w_n789_1;
	wire[2:0] w_n789_2;
	wire[2:0] w_n789_3;
	wire[2:0] w_n789_4;
	wire[1:0] w_n789_5;
	wire[2:0] w_n790_0;
	wire[2:0] w_n792_0;
	wire[2:0] w_n794_0;
	wire[2:0] w_n794_1;
	wire[2:0] w_n794_2;
	wire[2:0] w_n794_3;
	wire[2:0] w_n794_4;
	wire[2:0] w_n795_0;
	wire[1:0] w_n795_1;
	wire[2:0] w_n799_0;
	wire[2:0] w_n799_1;
	wire[2:0] w_n799_2;
	wire[2:0] w_n799_3;
	wire[2:0] w_n800_0;
	wire[2:0] w_n803_0;
	wire[2:0] w_n803_1;
	wire[2:0] w_n803_2;
	wire[2:0] w_n803_3;
	wire[2:0] w_n803_4;
	wire[2:0] w_n803_5;
	wire[2:0] w_n803_6;
	wire[2:0] w_n803_7;
	wire[2:0] w_n803_8;
	wire[2:0] w_n804_0;
	wire[2:0] w_n804_1;
	wire[2:0] w_n804_2;
	wire[2:0] w_n804_3;
	wire[2:0] w_n808_0;
	wire[2:0] w_n808_1;
	wire[2:0] w_n808_2;
	wire[2:0] w_n808_3;
	wire[2:0] w_n808_4;
	wire[2:0] w_n808_5;
	wire[2:0] w_n808_6;
	wire[2:0] w_n808_7;
	wire[2:0] w_n808_8;
	wire[2:0] w_n808_9;
	wire[2:0] w_n808_10;
	wire[2:0] w_n808_11;
	wire[2:0] w_n808_12;
	wire[2:0] w_n808_13;
	wire[1:0] w_n813_0;
	wire[2:0] w_n820_0;
	wire[2:0] w_n820_1;
	wire[2:0] w_n820_2;
	wire[2:0] w_n820_3;
	wire[2:0] w_n820_4;
	wire[2:0] w_n820_5;
	wire[2:0] w_n821_0;
	wire[1:0] w_n821_1;
	wire[2:0] w_n822_0;
	wire[2:0] w_n822_1;
	wire[1:0] w_n822_2;
	wire[1:0] w_n824_0;
	wire[2:0] w_n825_0;
	wire[2:0] w_n825_1;
	wire[2:0] w_n832_0;
	wire[1:0] w_n832_1;
	wire[1:0] w_n834_0;
	wire[1:0] w_n836_0;
	wire[2:0] w_n837_0;
	wire[2:0] w_n837_1;
	wire[1:0] w_n837_2;
	wire[1:0] w_n843_0;
	wire[1:0] w_n846_0;
	wire[2:0] w_n849_0;
	wire[2:0] w_n849_1;
	wire[1:0] w_n849_2;
	wire[1:0] w_n850_0;
	wire[1:0] w_n852_0;
	wire[2:0] w_n853_0;
	wire[2:0] w_n853_1;
	wire[2:0] w_n853_2;
	wire[2:0] w_n854_0;
	wire[1:0] w_n855_0;
	wire[1:0] w_n856_0;
	wire[1:0] w_n858_0;
	wire[1:0] w_n860_0;
	wire[1:0] w_n863_0;
	wire[1:0] w_n865_0;
	wire[1:0] w_n866_0;
	wire[2:0] w_n868_0;
	wire[1:0] w_n868_1;
	wire[2:0] w_n869_0;
	wire[1:0] w_n876_0;
	wire[1:0] w_n877_0;
	wire[2:0] w_n878_0;
	wire[1:0] w_n878_1;
	wire[1:0] w_n880_0;
	wire[2:0] w_n881_0;
	wire[1:0] w_n881_1;
	wire[2:0] w_n882_0;
	wire[2:0] w_n882_1;
	wire[1:0] w_n882_2;
	wire[1:0] w_n883_0;
	wire[1:0] w_n885_0;
	wire[2:0] w_n890_0;
	wire[2:0] w_n890_1;
	wire[1:0] w_n893_0;
	wire[1:0] w_n894_0;
	wire[1:0] w_n895_0;
	wire[2:0] w_n897_0;
	wire[1:0] w_n898_0;
	wire[1:0] w_n902_0;
	wire[1:0] w_n904_0;
	wire[1:0] w_n905_0;
	wire[1:0] w_n906_0;
	wire[1:0] w_n912_0;
	wire[1:0] w_n914_0;
	wire[1:0] w_n917_0;
	wire[2:0] w_n918_0;
	wire[2:0] w_n918_1;
	wire[1:0] w_n918_2;
	wire[1:0] w_n920_0;
	wire[1:0] w_n923_0;
	wire[2:0] w_n924_0;
	wire[2:0] w_n924_1;
	wire[2:0] w_n925_0;
	wire[1:0] w_n925_1;
	wire[1:0] w_n929_0;
	wire[2:0] w_n930_0;
	wire[1:0] w_n930_1;
	wire[1:0] w_n932_0;
	wire[1:0] w_n933_0;
	wire[2:0] w_n934_0;
	wire[2:0] w_n935_0;
	wire[2:0] w_n935_1;
	wire[2:0] w_n935_2;
	wire[1:0] w_n935_3;
	wire[2:0] w_n936_0;
	wire[2:0] w_n938_0;
	wire[2:0] w_n942_0;
	wire[1:0] w_n943_0;
	wire[1:0] w_n950_0;
	wire[2:0] w_n951_0;
	wire[2:0] w_n951_1;
	wire[2:0] w_n952_0;
	wire[2:0] w_n952_1;
	wire[2:0] w_n952_2;
	wire[2:0] w_n952_3;
	wire[1:0] w_n952_4;
	wire[2:0] w_n954_0;
	wire[2:0] w_n954_1;
	wire[2:0] w_n954_2;
	wire[2:0] w_n954_3;
	wire[2:0] w_n954_4;
	wire[2:0] w_n954_5;
	wire[2:0] w_n954_6;
	wire[2:0] w_n954_7;
	wire[2:0] w_n954_8;
	wire[2:0] w_n954_9;
	wire[2:0] w_n954_10;
	wire[2:0] w_n954_11;
	wire[2:0] w_n954_12;
	wire[2:0] w_n954_13;
	wire[2:0] w_n954_14;
	wire[2:0] w_n954_15;
	wire[2:0] w_n954_16;
	wire[2:0] w_n954_17;
	wire[2:0] w_n954_18;
	wire[2:0] w_n954_19;
	wire[2:0] w_n954_20;
	wire[2:0] w_n954_21;
	wire[2:0] w_n954_22;
	wire[2:0] w_n954_23;
	wire[1:0] w_n954_24;
	wire[2:0] w_n955_0;
	wire[2:0] w_n956_0;
	wire[2:0] w_n956_1;
	wire[2:0] w_n956_2;
	wire[2:0] w_n956_3;
	wire[1:0] w_n956_4;
	wire[1:0] w_n959_0;
	wire[2:0] w_n960_0;
	wire[2:0] w_n960_1;
	wire[2:0] w_n960_2;
	wire[2:0] w_n960_3;
	wire[2:0] w_n960_4;
	wire[2:0] w_n960_5;
	wire[2:0] w_n961_0;
	wire[2:0] w_n961_1;
	wire[2:0] w_n961_2;
	wire[2:0] w_n961_3;
	wire[2:0] w_n961_4;
	wire[1:0] w_n961_5;
	wire[1:0] w_n962_0;
	wire[2:0] w_n964_0;
	wire[1:0] w_n964_1;
	wire[1:0] w_n965_0;
	wire[2:0] w_n966_0;
	wire[2:0] w_n966_1;
	wire[2:0] w_n966_2;
	wire[2:0] w_n966_3;
	wire[1:0] w_n966_4;
	wire[1:0] w_n968_0;
	wire[2:0] w_n970_0;
	wire[2:0] w_n971_0;
	wire[2:0] w_n971_1;
	wire[2:0] w_n971_2;
	wire[2:0] w_n971_3;
	wire[1:0] w_n971_4;
	wire[1:0] w_n975_0;
	wire[2:0] w_n980_0;
	wire[2:0] w_n980_1;
	wire[2:0] w_n980_2;
	wire[2:0] w_n980_3;
	wire[2:0] w_n980_4;
	wire[2:0] w_n980_5;
	wire[1:0] w_n980_6;
	wire[2:0] w_n981_0;
	wire[2:0] w_n981_1;
	wire[2:0] w_n981_2;
	wire[2:0] w_n981_3;
	wire[2:0] w_n981_4;
	wire[1:0] w_n985_0;
	wire[1:0] w_n986_0;
	wire[2:0] w_n987_0;
	wire[2:0] w_n987_1;
	wire[1:0] w_n988_0;
	wire[1:0] w_n991_0;
	wire[2:0] w_n992_0;
	wire[2:0] w_n992_1;
	wire[2:0] w_n993_0;
	wire[2:0] w_n993_1;
	wire[1:0] w_n994_0;
	wire[2:0] w_n999_0;
	wire[1:0] w_n1000_0;
	wire[1:0] w_n1002_0;
	wire[1:0] w_n1006_0;
	wire[1:0] w_n1011_0;
	wire[1:0] w_n1013_0;
	wire[1:0] w_n1017_0;
	wire[2:0] w_n1018_0;
	wire[1:0] w_n1018_1;
	wire[1:0] w_n1020_0;
	wire[1:0] w_n1021_0;
	wire[2:0] w_n1022_0;
	wire[2:0] w_n1025_0;
	wire[1:0] w_n1026_0;
	wire[2:0] w_n1027_0;
	wire[1:0] w_n1032_0;
	wire[2:0] w_n1033_0;
	wire[2:0] w_n1033_1;
	wire[2:0] w_n1034_0;
	wire[2:0] w_n1034_1;
	wire[2:0] w_n1034_2;
	wire[2:0] w_n1034_3;
	wire[2:0] w_n1035_0;
	wire[2:0] w_n1037_0;
	wire[2:0] w_n1037_1;
	wire[2:0] w_n1037_2;
	wire[2:0] w_n1037_3;
	wire[2:0] w_n1038_0;
	wire[2:0] w_n1042_0;
	wire[2:0] w_n1043_0;
	wire[2:0] w_n1043_1;
	wire[2:0] w_n1043_2;
	wire[2:0] w_n1043_3;
	wire[1:0] w_n1043_4;
	wire[1:0] w_n1045_0;
	wire[2:0] w_n1047_0;
	wire[1:0] w_n1047_1;
	wire[2:0] w_n1049_0;
	wire[2:0] w_n1049_1;
	wire[2:0] w_n1049_2;
	wire[2:0] w_n1049_3;
	wire[1:0] w_n1049_4;
	wire[1:0] w_n1053_0;
	wire[1:0] w_n1055_0;
	wire[2:0] w_n1057_0;
	wire[2:0] w_n1057_1;
	wire[2:0] w_n1057_2;
	wire[2:0] w_n1057_3;
	wire[2:0] w_n1057_4;
	wire[1:0] w_n1057_5;
	wire[2:0] w_n1059_0;
	wire[2:0] w_n1059_1;
	wire[2:0] w_n1059_2;
	wire[2:0] w_n1059_3;
	wire[2:0] w_n1059_4;
	wire[2:0] w_n1059_5;
	wire[1:0] w_n1066_0;
	wire[1:0] w_n1068_0;
	wire[1:0] w_n1069_0;
	wire[1:0] w_n1071_0;
	wire[1:0] w_n1072_0;
	wire[2:0] w_n1073_0;
	wire[1:0] w_n1074_0;
	wire[1:0] w_n1075_0;
	wire[1:0] w_n1076_0;
	wire[1:0] w_n1078_0;
	wire[1:0] w_n1083_0;
	wire[1:0] w_n1085_0;
	wire[1:0] w_n1093_0;
	wire[1:0] w_n1095_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1109_0;
	wire[1:0] w_n1110_0;
	wire[1:0] w_n1111_0;
	wire[1:0] w_n1113_0;
	wire[1:0] w_n1114_0;
	wire[2:0] w_n1115_0;
	wire[1:0] w_n1120_0;
	wire[1:0] w_n1121_0;
	wire[1:0] w_n1129_0;
	wire[1:0] w_n1130_0;
	wire[1:0] w_n1133_0;
	wire[1:0] w_n1138_0;
	wire[1:0] w_n1139_0;
	wire[1:0] w_n1140_0;
	wire[2:0] w_n1143_0;
	wire[2:0] w_n1143_1;
	wire[2:0] w_n1143_2;
	wire[2:0] w_n1143_3;
	wire[2:0] w_n1143_4;
	wire[2:0] w_n1143_5;
	wire[2:0] w_n1143_6;
	wire[2:0] w_n1143_7;
	wire[2:0] w_n1143_8;
	wire[1:0] w_n1143_9;
	wire[1:0] w_n1150_0;
	wire[1:0] w_n1152_0;
	wire[1:0] w_n1159_0;
	wire[1:0] w_n1163_0;
	wire[1:0] w_n1169_0;
	wire[2:0] w_n1170_0;
	wire[1:0] w_n1175_0;
	wire[1:0] w_n1176_0;
	wire[1:0] w_n1179_0;
	wire[2:0] w_n1185_0;
	wire[2:0] w_n1185_1;
	wire[2:0] w_n1187_0;
	wire[1:0] w_n1188_0;
	wire[2:0] w_n1189_0;
	wire[1:0] w_n1189_1;
	wire[1:0] w_n1190_0;
	wire[1:0] w_n1192_0;
	wire[1:0] w_n1193_0;
	wire[2:0] w_n1196_0;
	wire[1:0] w_n1197_0;
	wire[1:0] w_n1198_0;
	wire[2:0] w_n1203_0;
	wire[2:0] w_n1204_0;
	wire[1:0] w_n1204_1;
	wire[2:0] w_n1209_0;
	wire[2:0] w_n1209_1;
	wire[1:0] w_n1210_0;
	wire[1:0] w_n1214_0;
	wire[1:0] w_n1215_0;
	wire[2:0] w_n1217_0;
	wire[2:0] w_n1218_0;
	wire[1:0] w_n1224_0;
	wire[1:0] w_n1227_0;
	wire[1:0] w_n1228_0;
	wire[2:0] w_n1231_0;
	wire[1:0] w_n1232_0;
	wire[1:0] w_n1239_0;
	wire[1:0] w_n1240_0;
	wire[2:0] w_n1243_0;
	wire[2:0] w_n1243_1;
	wire[1:0] w_n1243_2;
	wire[1:0] w_n1245_0;
	wire[1:0] w_n1259_0;
	wire[2:0] w_n1283_0;
	wire[2:0] w_n1283_1;
	wire[2:0] w_n1283_2;
	wire[2:0] w_n1283_3;
	wire[2:0] w_n1283_4;
	wire[2:0] w_n1283_5;
	wire[2:0] w_n1283_6;
	wire[2:0] w_n1283_7;
	wire[2:0] w_n1283_8;
	wire[2:0] w_n1283_9;
	wire[2:0] w_n1283_10;
	wire[2:0] w_n1283_11;
	wire[2:0] w_n1283_12;
	wire[1:0] w_n1285_0;
	wire[1:0] w_n1288_0;
	wire[1:0] w_n1292_0;
	wire[1:0] w_n1293_0;
	wire[1:0] w_n1294_0;
	wire[1:0] w_n1299_0;
	wire[1:0] w_n1302_0;
	wire[1:0] w_n1307_0;
	wire[1:0] w_n1309_0;
	wire[1:0] w_n1310_0;
	wire[1:0] w_n1312_0;
	wire[1:0] w_n1319_0;
	wire[1:0] w_n1322_0;
	wire[1:0] w_n1325_0;
	wire[2:0] w_n1328_0;
	wire[1:0] w_n1329_0;
	wire[1:0] w_n1332_0;
	wire[2:0] w_n1338_0;
	wire[2:0] w_n1339_0;
	wire[2:0] w_n1340_0;
	wire[1:0] w_n1342_0;
	wire[2:0] w_n1347_0;
	wire[2:0] w_n1347_1;
	wire[2:0] w_n1347_2;
	wire[2:0] w_n1347_3;
	wire[2:0] w_n1347_4;
	wire[2:0] w_n1347_5;
	wire[1:0] w_n1347_6;
	wire[1:0] w_n1348_0;
	wire[1:0] w_n1350_0;
	wire[1:0] w_n1351_0;
	wire[1:0] w_n1354_0;
	wire[2:0] w_n1356_0;
	wire[1:0] w_n1356_1;
	wire[1:0] w_n1358_0;
	wire[1:0] w_n1361_0;
	wire[2:0] w_n1362_0;
	wire[1:0] w_n1364_0;
	wire[1:0] w_n1367_0;
	wire[1:0] w_n1375_0;
	wire[1:0] w_n1377_0;
	wire[1:0] w_n1379_0;
	wire[1:0] w_n1380_0;
	wire[1:0] w_n1382_0;
	wire[1:0] w_n1383_0;
	wire[1:0] w_n1385_0;
	wire[1:0] w_n1386_0;
	wire[1:0] w_n1388_0;
	wire[1:0] w_n1389_0;
	wire[2:0] w_n1391_0;
	wire[2:0] w_n1391_1;
	wire[2:0] w_n1391_2;
	wire[2:0] w_n1391_3;
	wire[2:0] w_n1391_4;
	wire[2:0] w_n1391_5;
	wire[1:0] w_n1399_0;
	wire[1:0] w_n1407_0;
	wire[1:0] w_n1409_0;
	wire[2:0] w_n1411_0;
	wire[2:0] w_n1411_1;
	wire[2:0] w_n1411_2;
	wire[1:0] w_n1413_0;
	wire[2:0] w_n1414_0;
	wire[2:0] w_n1414_1;
	wire[2:0] w_n1414_2;
	wire[1:0] w_n1417_0;
	wire[2:0] w_n1418_0;
	wire[2:0] w_n1418_1;
	wire[2:0] w_n1418_2;
	wire[2:0] w_n1418_3;
	wire[1:0] w_n1418_4;
	wire[1:0] w_n1420_0;
	wire[2:0] w_n1421_0;
	wire[2:0] w_n1421_1;
	wire[2:0] w_n1421_2;
	wire[2:0] w_n1421_3;
	wire[1:0] w_n1421_4;
	wire[1:0] w_n1425_0;
	wire[1:0] w_n1427_0;
	wire[1:0] w_n1428_0;
	wire[1:0] w_n1430_0;
	wire[1:0] w_n1431_0;
	wire[1:0] w_n1433_0;
	wire[1:0] w_n1434_0;
	wire[1:0] w_n1436_0;
	wire[1:0] w_n1437_0;
	wire[1:0] w_n1439_0;
	wire[1:0] w_n1440_0;
	wire[1:0] w_n1442_0;
	wire[1:0] w_n1446_0;
	wire[1:0] w_n1454_0;
	wire[1:0] w_n1456_0;
	wire[1:0] w_n1458_0;
	wire[1:0] w_n1513_0;
	wire[1:0] w_n1514_0;
	wire[1:0] w_n1515_0;
	wire[1:0] w_n1517_0;
	wire[2:0] w_n1520_0;
	wire[1:0] w_n1521_0;
	wire[1:0] w_n1524_0;
	wire[1:0] w_n1526_0;
	wire[1:0] w_n1527_0;
	wire[1:0] w_n1529_0;
	wire[2:0] w_n1533_0;
	wire[2:0] w_n1533_1;
	wire[2:0] w_n1535_0;
	wire[2:0] w_n1535_1;
	wire[1:0] w_n1539_0;
	wire[1:0] w_n1541_0;
	wire[1:0] w_n1548_0;
	wire[1:0] w_n1550_0;
	wire[1:0] w_n1558_0;
	wire[1:0] w_n1560_0;
	wire[1:0] w_n1561_0;
	wire[1:0] w_n1563_0;
	wire[1:0] w_n1565_0;
	wire[2:0] w_n1566_0;
	wire[2:0] w_n1566_1;
	wire[2:0] w_n1566_2;
	wire[1:0] w_n1566_3;
	wire[2:0] w_n1568_0;
	wire[2:0] w_n1568_1;
	wire[2:0] w_n1568_2;
	wire[1:0] w_n1568_3;
	wire[2:0] w_n1571_0;
	wire[1:0] w_n1571_1;
	wire[2:0] w_n1572_0;
	wire[2:0] w_n1572_1;
	wire[2:0] w_n1572_2;
	wire[1:0] w_n1572_3;
	wire[1:0] w_n1574_0;
	wire[1:0] w_n1575_0;
	wire[2:0] w_n1576_0;
	wire[2:0] w_n1577_0;
	wire[2:0] w_n1577_1;
	wire[2:0] w_n1577_2;
	wire[1:0] w_n1577_3;
	wire[1:0] w_n1581_0;
	wire[1:0] w_n1583_0;
	wire[2:0] w_n1584_0;
	wire[2:0] w_n1584_1;
	wire[2:0] w_n1584_2;
	wire[2:0] w_n1584_3;
	wire[2:0] w_n1584_4;
	wire[1:0] w_n1592_0;
	wire[1:0] w_n1594_0;
	wire[1:0] w_n1595_0;
	wire[1:0] w_n1597_0;
	wire[1:0] w_n1604_0;
	wire[1:0] w_n1612_0;
	wire[1:0] w_n1614_0;
	wire[1:0] w_n1622_0;
	wire[1:0] w_n1624_0;
	wire[1:0] w_n1626_0;
	wire[1:0] w_n1627_0;
	wire[1:0] w_n1629_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1632_0;
	wire[1:0] w_n1634_0;
	wire[1:0] w_n1635_0;
	wire[1:0] w_n1637_0;
	wire[1:0] w_n1638_0;
	wire[1:0] w_n1640_0;
	wire[1:0] w_n1641_0;
	wire[2:0] w_n1646_0;
	wire[1:0] w_n1653_0;
	wire[1:0] w_n1658_0;
	wire[1:0] w_n1669_0;
	wire[1:0] w_n1673_0;
	wire[1:0] w_n1675_0;
	wire[1:0] w_n1676_0;
	wire[1:0] w_n1679_0;
	wire[2:0] w_n1682_0;
	wire[2:0] w_n1682_1;
	wire[2:0] w_n1682_2;
	wire[2:0] w_n1682_3;
	wire[2:0] w_n1682_4;
	wire[1:0] w_n1682_5;
	wire[2:0] w_n1683_0;
	wire[2:0] w_n1683_1;
	wire[2:0] w_n1683_2;
	wire[2:0] w_n1683_3;
	wire[2:0] w_n1683_4;
	wire[1:0] w_n1685_0;
	wire[1:0] w_n1687_0;
	wire[2:0] w_n1688_0;
	wire[1:0] w_n1688_1;
	wire[2:0] w_n1690_0;
	wire[1:0] w_n1690_1;
	wire[1:0] w_n1697_0;
	wire[1:0] w_n1699_0;
	wire[1:0] w_n1707_0;
	wire[1:0] w_n1709_0;
	wire[1:0] w_n1717_0;
	wire[1:0] w_n1725_0;
	wire[1:0] w_n1727_0;
	wire[1:0] w_n1735_0;
	wire[1:0] w_n1737_0;
	wire[1:0] w_n1739_0;
	wire[1:0] w_n1740_0;
	wire[1:0] w_n1742_0;
	wire[1:0] w_n1743_0;
	wire[1:0] w_n1745_0;
	wire[1:0] w_n1746_0;
	wire[1:0] w_n1748_0;
	wire[1:0] w_n1749_0;
	wire[1:0] w_n1751_0;
	wire[1:0] w_n1754_0;
	wire[1:0] w_n1760_0;
	wire[1:0] w_n1761_0;
	wire[2:0] w_n1762_0;
	wire[2:0] w_n1762_1;
	wire[2:0] w_n1762_2;
	wire[2:0] w_n1762_3;
	wire[2:0] w_n1762_4;
	wire[1:0] w_n1762_5;
	wire[1:0] w_n1770_0;
	wire[1:0] w_n1779_0;
	wire[1:0] w_n1787_0;
	wire[1:0] w_n1789_0;
	wire[1:0] w_n1797_0;
	wire[1:0] w_n1799_0;
	wire[1:0] w_n1800_0;
	wire[1:0] w_n1802_0;
	wire[1:0] w_n1803_0;
	wire[1:0] w_n1805_0;
	wire[1:0] w_n1806_0;
	wire[1:0] w_n1808_0;
	wire[1:0] w_n1809_0;
	wire[1:0] w_n1811_0;
	wire[1:0] w_n1812_0;
	wire[1:0] w_n1814_0;
	wire[1:0] w_n1815_0;
	wire[1:0] w_n1824_0;
	wire[1:0] w_n1832_0;
	wire[1:0] w_n1834_0;
	wire[1:0] w_n1835_0;
	wire[1:0] w_n1837_0;
	wire[1:0] w_n1838_0;
	wire[1:0] w_n1840_0;
	wire[1:0] w_n1841_0;
	wire[1:0] w_n1843_0;
	wire[1:0] w_n1844_0;
	wire[1:0] w_n1846_0;
	wire[1:0] w_n1847_0;
	wire[1:0] w_n1849_0;
	wire[1:0] w_n1850_0;
	wire[1:0] w_n1858_0;
	wire[1:0] w_n1866_0;
	wire[2:0] w_n1869_0;
	wire[1:0] w_n1871_0;
	wire[1:0] w_n1872_0;
	wire[1:0] w_n1878_0;
	wire[1:0] w_n1879_0;
	wire[1:0] w_n1880_0;
	wire[1:0] w_n1882_0;
	wire[1:0] w_n1883_0;
	wire[1:0] w_n1889_0;
	wire[1:0] w_n1897_0;
	wire[1:0] w_n1899_0;
	wire[1:0] w_n1907_0;
	wire[1:0] w_n1909_0;
	wire[1:0] w_n1911_0;
	wire[1:0] w_n1912_0;
	wire[1:0] w_n1914_0;
	wire[1:0] w_n1915_0;
	wire[1:0] w_n1917_0;
	wire[1:0] w_n1918_0;
	wire[1:0] w_n1920_0;
	wire[1:0] w_n1921_0;
	wire[1:0] w_n1930_0;
	wire[1:0] w_n1938_0;
	wire[1:0] w_n1940_0;
	wire[1:0] w_n1948_0;
	wire[1:0] w_n1950_0;
	wire[1:0] w_n1952_0;
	wire[1:0] w_n1953_0;
	wire[1:0] w_n1955_0;
	wire[1:0] w_n1956_0;
	wire[1:0] w_n1958_0;
	wire[1:0] w_n1959_0;
	wire[1:0] w_n1961_0;
	wire[1:0] w_n1962_0;
	wire[1:0] w_n1964_0;
	wire[1:0] w_n1965_0;
	wire[1:0] w_n1973_0;
	wire[1:0] w_n1975_0;
	wire[1:0] w_n1981_0;
	wire[1:0] w_n1989_0;
	wire[1:0] w_n1991_0;
	wire[1:0] w_n1999_0;
	wire[1:0] w_n2001_0;
	wire[1:0] w_n2002_0;
	wire[1:0] w_n2004_0;
	wire[1:0] w_n2005_0;
	wire[1:0] w_n2007_0;
	wire[1:0] w_n2008_0;
	wire[1:0] w_n2010_0;
	wire[2:0] w_n2011_0;
	wire[1:0] w_n2013_0;
	wire[1:0] w_n2014_0;
	wire[1:0] w_n2020_0;
	wire[1:0] w_n2021_0;
	wire[1:0] w_n2029_0;
	wire[1:0] w_n2031_0;
	wire[1:0] w_n2033_0;
	wire[1:0] w_n2034_0;
	wire[1:0] w_n2036_0;
	wire[1:0] w_n2037_0;
	wire[1:0] w_n2039_0;
	wire[1:0] w_n2047_0;
	wire[1:0] w_n2055_0;
	wire[1:0] w_n2057_0;
	wire[1:0] w_n2065_0;
	wire[1:0] w_n2067_0;
	wire[1:0] w_n2068_0;
	wire[1:0] w_n2070_0;
	wire[1:0] w_n2071_0;
	wire[1:0] w_n2073_0;
	wire[1:0] w_n2074_0;
	wire[1:0] w_n2075_0;
	wire[1:0] w_n2081_0;
	wire[1:0] w_n2089_0;
	wire[1:0] w_n2091_0;
	wire[1:0] w_n2099_0;
	wire[1:0] w_n2101_0;
	wire[1:0] w_n2103_0;
	wire[1:0] w_n2104_0;
	wire[1:0] w_n2106_0;
	wire[2:0] w_n2107_0;
	wire[1:0] w_n2109_0;
	wire[1:0] w_n2110_0;
	wire[1:0] w_n2116_0;
	wire[1:0] w_n2117_0;
	wire[1:0] w_n2125_0;
	wire[1:0] w_n2132_0;
	wire[1:0] w_n2134_0;
	wire[1:0] w_n2135_0;
	wire[1:0] w_n2137_0;
	wire[1:0] w_n2138_0;
	wire[1:0] w_n2140_0;
	wire[1:0] w_n2141_0;
	wire[1:0] w_n2142_0;
	wire[1:0] w_n2148_0;
	wire[1:0] w_n2155_0;
	wire[1:0] w_n2157_0;
	wire[1:0] w_n2159_0;
	wire[1:0] w_n2160_0;
	wire[1:0] w_n2166_0;
	wire[1:0] w_n2167_0;
	wire[1:0] w_n2168_0;
	wire[1:0] w_n2170_0;
	wire[1:0] w_n2171_0;
	wire[1:0] w_n2174_0;
	wire[1:0] w_n2180_0;
	wire[1:0] w_n2184_0;
	wire[1:0] w_n2187_0;
	wire[1:0] w_n2191_0;
	wire[1:0] w_n2197_0;
	wire[1:0] w_n2201_0;
	wire[1:0] w_n2208_0;
	wire[1:0] w_n2213_0;
	wire[1:0] w_n2218_0;
	wire[1:0] w_n2223_0;
	wire[1:0] w_n2228_0;
	wire[1:0] w_n2233_0;
	wire[1:0] w_n2238_0;
	wire[1:0] w_n2240_0;
	wire[1:0] w_n2241_0;
	wire[1:0] w_n2243_0;
	wire[1:0] w_n2244_0;
	wire[1:0] w_n2246_0;
	wire[1:0] w_n2247_0;
	wire[1:0] w_n2249_0;
	wire[1:0] w_n2250_0;
	wire[1:0] w_n2252_0;
	wire[1:0] w_n2253_0;
	wire[1:0] w_n2255_0;
	wire[1:0] w_n2256_0;
	wire[1:0] w_n2258_0;
	wire[1:0] w_n2259_0;
	wire[1:0] w_n2261_0;
	wire[1:0] w_n2262_0;
	wire[1:0] w_n2264_0;
	wire[1:0] w_n2267_0;
	wire[1:0] w_n2270_0;
	wire[1:0] w_n2278_0;
	wire[1:0] w_n2279_0;
	wire[1:0] w_n2280_0;
	wire[1:0] w_n2281_0;
	wire[1:0] w_n2282_0;
	wire[1:0] w_n2283_0;
	wire[1:0] w_n2284_0;
	wire[1:0] w_n2285_0;
	wire[1:0] w_n2286_0;
	wire[1:0] w_n2287_0;
	wire[1:0] w_n2289_0;
	wire[1:0] w_n2300_0;
	wire[1:0] w_n2302_0;
	wire[1:0] w_n2305_0;
	wire[1:0] w_n2307_0;
	wire[1:0] w_n2313_0;
	wire[1:0] w_n2315_0;
	wire[2:0] w_n2321_0;
	wire[1:0] w_n2323_0;
	wire[2:0] w_n2326_0;
	wire[1:0] w_n2330_0;
	wire[1:0] w_n2331_0;
	wire[1:0] w_n2332_0;
	wire[2:0] w_n2334_0;
	wire[1:0] w_n2335_0;
	wire[1:0] w_n2339_0;
	wire[1:0] w_n2345_0;
	wire[1:0] w_n2347_0;
	wire[1:0] w_n2350_0;
	wire[1:0] w_n2351_0;
	wire[1:0] w_n2359_0;
	wire[1:0] w_n2360_0;
	wire[2:0] w_n2365_0;
	wire[2:0] w_n2372_0;
	wire[1:0] w_n2377_0;
	wire[1:0] w_n2379_0;
	wire[2:0] w_n2380_0;
	wire[2:0] w_n2380_1;
	wire[2:0] w_n2380_2;
	wire[1:0] w_n2380_3;
	wire[1:0] w_n2382_0;
	wire[2:0] w_n2385_0;
	wire[1:0] w_n2385_1;
	wire[1:0] w_n2387_0;
	wire[1:0] w_n2391_0;
	wire[1:0] w_n2396_0;
	wire[1:0] w_n2398_0;
	wire[1:0] w_n2402_0;
	wire[1:0] w_n2406_0;
	wire[1:0] w_n2412_0;
	wire[1:0] w_n2414_0;
	wire[2:0] w_n2417_0;
	wire[1:0] w_n2424_0;
	wire[2:0] w_n2427_0;
	wire[1:0] w_n2428_0;
	wire[2:0] w_n2429_0;
	wire[1:0] w_n2429_1;
	wire[1:0] w_n2438_0;
	wire[1:0] w_n2440_0;
	wire[1:0] w_n2442_0;
	wire[1:0] w_n2449_0;
	wire[1:0] w_n2451_0;
	wire[1:0] w_n2453_0;
	wire[2:0] w_n2456_0;
	wire[1:0] w_n2457_0;
	wire[1:0] w_n2461_0;
	wire[1:0] w_n2466_0;
	wire[1:0] w_n2477_0;
	wire[2:0] w_n2479_0;
	wire[1:0] w_n2486_0;
	wire[1:0] w_n2490_0;
	wire[1:0] w_n2498_0;
	wire[2:0] w_n2504_0;
	wire[1:0] w_n2506_0;
	wire[2:0] w_n2511_0;
	wire[1:0] w_n2511_1;
	wire[1:0] w_n2514_0;
	wire[2:0] w_n2515_0;
	wire[2:0] w_n2520_0;
	wire[2:0] w_n2521_0;
	wire[1:0] w_n2521_1;
	wire[1:0] w_n2534_0;
	wire[1:0] w_n2536_0;
	wire[1:0] w_n2538_0;
	wire[1:0] w_n2540_0;
	wire[1:0] w_n2541_0;
	wire[1:0] w_n2542_0;
	wire[1:0] w_n2544_0;
	wire[1:0] w_n2551_0;
	wire[1:0] w_n2552_0;
	wire[1:0] w_n2564_0;
	wire[1:0] w_n2566_0;
	wire[1:0] w_n2571_0;
	wire[2:0] w_n2575_0;
	wire[1:0] w_n2580_0;
	wire[1:0] w_n2586_0;
	wire[1:0] w_n2587_0;
	wire[2:0] w_n2589_0;
	wire[1:0] w_n2591_0;
	wire[1:0] w_n2593_0;
	wire[1:0] w_n2595_0;
	wire[1:0] w_n2599_0;
	wire[1:0] w_n2600_0;
	wire[2:0] w_n2603_0;
	wire[1:0] w_n2604_0;
	wire[1:0] w_n2605_0;
	wire[1:0] w_n2607_0;
	wire[1:0] w_n2608_0;
	wire[1:0] w_n2611_0;
	wire[1:0] w_n2612_0;
	wire[1:0] w_n2615_0;
	wire[1:0] w_n2617_0;
	wire[1:0] w_n2620_0;
	wire[1:0] w_n2621_0;
	wire[1:0] w_n2624_0;
	wire[1:0] w_n2627_0;
	wire[1:0] w_n2630_0;
	wire[1:0] w_n2633_0;
	wire[1:0] w_n2634_0;
	wire[1:0] w_n2640_0;
	wire[1:0] w_n2641_0;
	wire[1:0] w_n2642_0;
	wire[1:0] w_n2643_0;
	wire[1:0] w_n2644_0;
	wire[1:0] w_n2655_0;
	wire[1:0] w_n2658_0;
	wire[1:0] w_n2665_0;
	wire[1:0] w_n2667_0;
	wire[1:0] w_n2668_0;
	wire[2:0] w_n2669_0;
	wire[2:0] w_n2669_1;
	wire[2:0] w_n2669_2;
	wire[2:0] w_n2669_3;
	wire[2:0] w_n2670_0;
	wire[2:0] w_n2670_1;
	wire[2:0] w_n2670_2;
	wire[2:0] w_n2670_3;
	wire[2:0] w_n2670_4;
	wire[2:0] w_n2670_5;
	wire[2:0] w_n2671_0;
	wire[2:0] w_n2671_1;
	wire[2:0] w_n2671_2;
	wire[2:0] w_n2671_3;
	wire[2:0] w_n2671_4;
	wire[2:0] w_n2671_5;
	wire[1:0] w_n2671_6;
	wire[2:0] w_n2672_0;
	wire[2:0] w_n2672_1;
	wire[2:0] w_n2672_2;
	wire[2:0] w_n2674_0;
	wire[2:0] w_n2674_1;
	wire[2:0] w_n2674_2;
	wire[2:0] w_n2674_3;
	wire[1:0] w_n2674_4;
	wire[2:0] w_n2677_0;
	wire[2:0] w_n2677_1;
	wire[2:0] w_n2677_2;
	wire[2:0] w_n2677_3;
	wire[2:0] w_n2677_4;
	wire[2:0] w_n2678_0;
	wire[2:0] w_n2678_1;
	wire[2:0] w_n2678_2;
	wire[2:0] w_n2678_3;
	wire[2:0] w_n2678_4;
	wire[2:0] w_n2678_5;
	wire[1:0] w_n2678_6;
	wire[2:0] w_n2679_0;
	wire[2:0] w_n2679_1;
	wire[2:0] w_n2679_2;
	wire[1:0] w_n2679_3;
	wire[2:0] w_n2681_0;
	wire[2:0] w_n2681_1;
	wire[2:0] w_n2681_2;
	wire[2:0] w_n2681_3;
	wire[2:0] w_n2681_4;
	wire[1:0] w_n2681_5;
	wire[2:0] w_n2684_0;
	wire[2:0] w_n2684_1;
	wire[2:0] w_n2684_2;
	wire[2:0] w_n2684_3;
	wire[1:0] w_n2684_4;
	wire[2:0] w_n2685_0;
	wire[2:0] w_n2685_1;
	wire[1:0] w_n2685_2;
	wire[2:0] w_n2687_0;
	wire[2:0] w_n2687_1;
	wire[2:0] w_n2687_2;
	wire[2:0] w_n2687_3;
	wire[2:0] w_n2687_4;
	wire[2:0] w_n2687_5;
	wire[2:0] w_n2687_6;
	wire[1:0] w_n2687_7;
	wire[2:0] w_n2688_0;
	wire[2:0] w_n2688_1;
	wire[2:0] w_n2688_2;
	wire[2:0] w_n2688_3;
	wire[2:0] w_n2688_4;
	wire[2:0] w_n2688_5;
	wire[2:0] w_n2688_6;
	wire[2:0] w_n2688_7;
	wire[2:0] w_n2688_8;
	wire[2:0] w_n2691_0;
	wire[2:0] w_n2691_1;
	wire[2:0] w_n2691_2;
	wire[2:0] w_n2691_3;
	wire[2:0] w_n2691_4;
	wire[2:0] w_n2691_5;
	wire[2:0] w_n2691_6;
	wire[2:0] w_n2691_7;
	wire[2:0] w_n2691_8;
	wire[2:0] w_n2693_0;
	wire[2:0] w_n2693_1;
	wire[2:0] w_n2693_2;
	wire[2:0] w_n2693_3;
	wire[2:0] w_n2693_4;
	wire[2:0] w_n2694_0;
	wire[2:0] w_n2694_1;
	wire[2:0] w_n2694_2;
	wire[2:0] w_n2694_3;
	wire[2:0] w_n2694_4;
	wire[2:0] w_n2696_0;
	wire[2:0] w_n2697_0;
	wire[1:0] w_n2697_1;
	wire[2:0] w_n2698_0;
	wire[2:0] w_n2698_1;
	wire[2:0] w_n2698_2;
	wire[2:0] w_n2698_3;
	wire[2:0] w_n2698_4;
	wire[2:0] w_n2698_5;
	wire[1:0] w_n2698_6;
	wire[2:0] w_n2700_0;
	wire[2:0] w_n2700_1;
	wire[2:0] w_n2700_2;
	wire[2:0] w_n2700_3;
	wire[2:0] w_n2700_4;
	wire[2:0] w_n2700_5;
	wire[1:0] w_n2701_0;
	wire[1:0] w_n2702_0;
	wire[1:0] w_n2704_0;
	wire[1:0] w_n2705_0;
	wire[1:0] w_n2708_0;
	wire[1:0] w_n2711_0;
	wire[1:0] w_n2713_0;
	wire[1:0] w_n2715_0;
	wire[1:0] w_n2718_0;
	wire[1:0] w_n2719_0;
	wire[1:0] w_n2721_0;
	wire[1:0] w_n2722_0;
	wire[1:0] w_n2724_0;
	wire[1:0] w_n2725_0;
	wire[1:0] w_n2727_0;
	wire[1:0] w_n2733_0;
	wire[2:0] w_n2734_0;
	wire[2:0] w_n2736_0;
	wire[1:0] w_n2736_1;
	wire[1:0] w_n2743_0;
	wire[1:0] w_n2745_0;
	wire[2:0] w_n2750_0;
	wire[1:0] w_n2751_0;
	wire[2:0] w_n2752_0;
	wire[2:0] w_n2767_0;
	wire[2:0] w_n2769_0;
	wire[2:0] w_n2769_1;
	wire[2:0] w_n2769_2;
	wire[2:0] w_n2769_3;
	wire[1:0] w_n2769_4;
	wire[2:0] w_n2770_0;
	wire[2:0] w_n2771_0;
	wire[2:0] w_n2771_1;
	wire[2:0] w_n2773_0;
	wire[2:0] w_n2773_1;
	wire[2:0] w_n2773_2;
	wire[2:0] w_n2773_3;
	wire[2:0] w_n2773_4;
	wire[2:0] w_n2774_0;
	wire[2:0] w_n2774_1;
	wire[1:0] w_n2774_2;
	wire[2:0] w_n2775_0;
	wire[2:0] w_n2775_1;
	wire[2:0] w_n2775_2;
	wire[2:0] w_n2775_3;
	wire[2:0] w_n2775_4;
	wire[2:0] w_n2775_5;
	wire[1:0] w_n2777_0;
	wire[2:0] w_n2779_0;
	wire[2:0] w_n2779_1;
	wire[2:0] w_n2779_2;
	wire[2:0] w_n2780_0;
	wire[2:0] w_n2780_1;
	wire[2:0] w_n2780_2;
	wire[2:0] w_n2780_3;
	wire[2:0] w_n2780_4;
	wire[2:0] w_n2780_5;
	wire[2:0] w_n2783_0;
	wire[2:0] w_n2783_1;
	wire[1:0] w_n2783_2;
	wire[2:0] w_n2784_0;
	wire[2:0] w_n2784_1;
	wire[2:0] w_n2784_2;
	wire[2:0] w_n2784_3;
	wire[2:0] w_n2784_4;
	wire[2:0] w_n2784_5;
	wire[1:0] w_n2784_6;
	wire[1:0] w_n2789_0;
	wire[2:0] w_n2790_0;
	wire[2:0] w_n2791_0;
	wire[1:0] w_n2792_0;
	wire[1:0] w_n2793_0;
	wire[2:0] w_n2794_0;
	wire[2:0] w_n2794_1;
	wire[2:0] w_n2794_2;
	wire[2:0] w_n2795_0;
	wire[2:0] w_n2795_1;
	wire[2:0] w_n2795_2;
	wire[2:0] w_n2795_3;
	wire[2:0] w_n2795_4;
	wire[2:0] w_n2795_5;
	wire[1:0] w_n2795_6;
	wire[2:0] w_n2797_0;
	wire[2:0] w_n2797_1;
	wire[2:0] w_n2799_0;
	wire[2:0] w_n2799_1;
	wire[1:0] w_n2799_2;
	wire[2:0] w_n2800_0;
	wire[2:0] w_n2800_1;
	wire[2:0] w_n2800_2;
	wire[2:0] w_n2800_3;
	wire[2:0] w_n2800_4;
	wire[2:0] w_n2800_5;
	wire[1:0] w_n2802_0;
	wire[2:0] w_n2804_0;
	wire[2:0] w_n2804_1;
	wire[2:0] w_n2804_2;
	wire[2:0] w_n2805_0;
	wire[2:0] w_n2805_1;
	wire[2:0] w_n2805_2;
	wire[2:0] w_n2805_3;
	wire[2:0] w_n2805_4;
	wire[2:0] w_n2805_5;
	wire[2:0] w_n2808_0;
	wire[2:0] w_n2808_1;
	wire[1:0] w_n2808_2;
	wire[2:0] w_n2809_0;
	wire[2:0] w_n2809_1;
	wire[2:0] w_n2809_2;
	wire[2:0] w_n2809_3;
	wire[2:0] w_n2809_4;
	wire[2:0] w_n2809_5;
	wire[1:0] w_n2809_6;
	wire[1:0] w_n2815_0;
	wire[2:0] w_n2816_0;
	wire[2:0] w_n2817_0;
	wire[1:0] w_n2817_1;
	wire[2:0] w_n2818_0;
	wire[1:0] w_n2821_0;
	wire[1:0] w_n2822_0;
	wire[2:0] w_n2823_0;
	wire[1:0] w_n2823_1;
	wire[2:0] w_n2824_0;
	wire[2:0] w_n2825_0;
	wire[1:0] w_n2826_0;
	wire[1:0] w_n2827_0;
	wire[2:0] w_n2828_0;
	wire[2:0] w_n2828_1;
	wire[2:0] w_n2828_2;
	wire[1:0] w_n2830_0;
	wire[2:0] w_n2832_0;
	wire[2:0] w_n2832_1;
	wire[2:0] w_n2832_2;
	wire[2:0] w_n2834_0;
	wire[2:0] w_n2834_1;
	wire[1:0] w_n2834_2;
	wire[1:0] w_n2837_0;
	wire[2:0] w_n2839_0;
	wire[1:0] w_n2839_1;
	wire[1:0] w_n2842_0;
	wire[2:0] w_n2844_0;
	wire[1:0] w_n2844_1;
	wire[2:0] w_n2848_0;
	wire[2:0] w_n2848_1;
	wire[1:0] w_n2848_2;
	wire[1:0] w_n2854_0;
	wire[1:0] w_n2855_0;
	wire[2:0] w_n2857_0;
	wire[2:0] w_n2857_1;
	wire[2:0] w_n2857_2;
	wire[2:0] w_n2857_3;
	wire[2:0] w_n2857_4;
	wire[2:0] w_n2857_5;
	wire[1:0] w_n2857_6;
	wire[2:0] w_n2858_0;
	wire[2:0] w_n2858_1;
	wire[2:0] w_n2860_0;
	wire[2:0] w_n2860_1;
	wire[2:0] w_n2860_2;
	wire[2:0] w_n2860_3;
	wire[2:0] w_n2860_4;
	wire[2:0] w_n2860_5;
	wire[2:0] w_n2862_0;
	wire[2:0] w_n2862_1;
	wire[2:0] w_n2862_2;
	wire[2:0] w_n2863_0;
	wire[2:0] w_n2863_1;
	wire[2:0] w_n2863_2;
	wire[2:0] w_n2863_3;
	wire[2:0] w_n2863_4;
	wire[2:0] w_n2863_5;
	wire[1:0] w_n2863_6;
	wire[2:0] w_n2865_0;
	wire[2:0] w_n2865_1;
	wire[2:0] w_n2865_2;
	wire[2:0] w_n2865_3;
	wire[2:0] w_n2865_4;
	wire[2:0] w_n2865_5;
	wire[1:0] w_n2870_0;
	wire[1:0] w_n2871_0;
	wire[1:0] w_n2873_0;
	wire[2:0] w_n2874_0;
	wire[2:0] w_n2874_1;
	wire[1:0] w_n2882_0;
	wire[2:0] w_n2883_0;
	wire[2:0] w_n2883_1;
	wire[2:0] w_n2883_2;
	wire[1:0] w_n2883_3;
	wire[1:0] w_n2885_0;
	wire[2:0] w_n2887_0;
	wire[2:0] w_n2887_1;
	wire[2:0] w_n2887_2;
	wire[2:0] w_n2887_3;
	wire[2:0] w_n2887_4;
	wire[2:0] w_n2889_0;
	wire[2:0] w_n2889_1;
	wire[2:0] w_n2889_2;
	wire[2:0] w_n2889_3;
	wire[1:0] w_n2889_4;
	wire[1:0] w_n2892_0;
	wire[2:0] w_n2893_0;
	wire[1:0] w_n2895_0;
	wire[1:0] w_n2896_0;
	wire[1:0] w_n2897_0;
	wire[2:0] w_n2899_0;
	wire[2:0] w_n2899_1;
	wire[1:0] w_n2907_0;
	wire[1:0] w_n2908_0;
	wire[2:0] w_n2911_0;
	wire[2:0] w_n2911_1;
	wire[1:0] w_n2920_0;
	wire[1:0] w_n2922_0;
	wire[1:0] w_n2931_0;
	wire[1:0] w_n2933_0;
	wire[1:0] w_n2939_0;
	wire[2:0] w_n2941_0;
	wire[1:0] w_n2941_1;
	wire[1:0] w_n2944_0;
	wire[1:0] w_n2952_0;
	wire[1:0] w_n2953_0;
	wire[1:0] w_n2963_0;
	wire[1:0] w_n2964_0;
	wire[1:0] w_n2966_0;
	wire[1:0] w_n2967_0;
	wire[1:0] w_n2969_0;
	wire[1:0] w_n2970_0;
	wire[1:0] w_n2972_0;
	wire[1:0] w_n2973_0;
	wire[1:0] w_n2975_0;
	wire[1:0] w_n2976_0;
	wire[1:0] w_n2978_0;
	wire[1:0] w_n2981_0;
	wire[1:0] w_n2989_0;
	wire[1:0] w_n2990_0;
	wire[2:0] w_n2995_0;
	wire[2:0] w_n2995_1;
	wire[2:0] w_n2995_2;
	wire[2:0] w_n2995_3;
	wire[2:0] w_n2995_4;
	wire[1:0] w_n3000_0;
	wire[1:0] w_n3001_0;
	wire[1:0] w_n3002_0;
	wire[1:0] w_n3003_0;
	wire[2:0] w_n3004_0;
	wire[2:0] w_n3004_1;
	wire[1:0] w_n3012_0;
	wire[1:0] w_n3013_0;
	wire[1:0] w_n3014_0;
	wire[2:0] w_n3016_0;
	wire[2:0] w_n3016_1;
	wire[1:0] w_n3024_0;
	wire[1:0] w_n3025_0;
	wire[2:0] w_n3028_0;
	wire[2:0] w_n3028_1;
	wire[1:0] w_n3036_0;
	wire[1:0] w_n3037_0;
	wire[1:0] w_n3046_0;
	wire[1:0] w_n3047_0;
	wire[1:0] w_n3056_0;
	wire[1:0] w_n3057_0;
	wire[1:0] w_n3066_0;
	wire[1:0] w_n3067_0;
	wire[1:0] w_n3076_0;
	wire[1:0] w_n3078_0;
	wire[1:0] w_n3087_0;
	wire[1:0] w_n3089_0;
	wire[1:0] w_n3095_0;
	wire[2:0] w_n3097_0;
	wire[1:0] w_n3100_0;
	wire[1:0] w_n3107_0;
	wire[1:0] w_n3109_0;
	wire[1:0] w_n3118_0;
	wire[1:0] w_n3119_0;
	wire[1:0] w_n3121_0;
	wire[1:0] w_n3122_0;
	wire[1:0] w_n3124_0;
	wire[1:0] w_n3125_0;
	wire[1:0] w_n3127_0;
	wire[1:0] w_n3128_0;
	wire[1:0] w_n3130_0;
	wire[1:0] w_n3131_0;
	wire[1:0] w_n3133_0;
	wire[1:0] w_n3134_0;
	wire[1:0] w_n3136_0;
	wire[1:0] w_n3137_0;
	wire[1:0] w_n3139_0;
	wire[1:0] w_n3140_0;
	wire[1:0] w_n3142_0;
	wire[1:0] w_n3143_0;
	wire[1:0] w_n3145_0;
	wire[1:0] w_n3148_0;
	wire[1:0] w_n3154_0;
	wire[1:0] w_n3155_0;
	wire[1:0] w_n3159_0;
	wire[1:0] w_n3171_0;
	wire[2:0] w_n3172_0;
	wire[2:0] w_n3172_1;
	wire[2:0] w_n3172_2;
	wire[2:0] w_n3172_3;
	wire[2:0] w_n3172_4;
	wire[2:0] w_n3172_5;
	wire[1:0] w_n3172_6;
	wire[1:0] w_n3173_0;
	wire[2:0] w_n3174_0;
	wire[2:0] w_n3174_1;
	wire[2:0] w_n3176_0;
	wire[2:0] w_n3176_1;
	wire[2:0] w_n3176_2;
	wire[1:0] w_n3183_0;
	wire[1:0] w_n3186_0;
	wire[1:0] w_n3189_0;
	wire[1:0] w_n3197_0;
	wire[2:0] w_n3198_0;
	wire[2:0] w_n3198_1;
	wire[2:0] w_n3198_2;
	wire[2:0] w_n3198_3;
	wire[2:0] w_n3198_4;
	wire[2:0] w_n3198_5;
	wire[2:0] w_n3200_0;
	wire[2:0] w_n3200_1;
	wire[2:0] w_n3200_2;
	wire[2:0] w_n3200_3;
	wire[2:0] w_n3202_0;
	wire[2:0] w_n3202_1;
	wire[2:0] w_n3202_2;
	wire[2:0] w_n3202_3;
	wire[2:0] w_n3204_0;
	wire[2:0] w_n3204_1;
	wire[2:0] w_n3204_2;
	wire[2:0] w_n3204_3;
	wire[1:0] w_n3210_0;
	wire[1:0] w_n3212_0;
	wire[1:0] w_n3215_0;
	wire[1:0] w_n3217_0;
	wire[1:0] w_n3218_0;
	wire[1:0] w_n3219_0;
	wire[1:0] w_n3220_0;
	wire[1:0] w_n3228_0;
	wire[1:0] w_n3229_0;
	wire[1:0] w_n3230_0;
	wire[1:0] w_n3231_0;
	wire[1:0] w_n3232_0;
	wire[2:0] w_n3233_0;
	wire[2:0] w_n3233_1;
	wire[2:0] w_n3233_2;
	wire[2:0] w_n3233_3;
	wire[2:0] w_n3233_4;
	wire[2:0] w_n3233_5;
	wire[2:0] w_n3233_6;
	wire[2:0] w_n3233_7;
	wire[2:0] w_n3233_8;
	wire[2:0] w_n3233_9;
	wire[1:0] w_n3235_0;
	wire[1:0] w_n3236_0;
	wire[2:0] w_n3237_0;
	wire[2:0] w_n3237_1;
	wire[1:0] w_n3237_2;
	wire[2:0] w_n3238_0;
	wire[2:0] w_n3238_1;
	wire[2:0] w_n3238_2;
	wire[2:0] w_n3238_3;
	wire[2:0] w_n3238_4;
	wire[2:0] w_n3238_5;
	wire[2:0] w_n3238_6;
	wire[1:0] w_n3238_7;
	wire[1:0] w_n3240_0;
	wire[2:0] w_n3242_0;
	wire[1:0] w_n3250_0;
	wire[2:0] w_n3256_0;
	wire[1:0] w_n3257_0;
	wire[2:0] w_n3258_0;
	wire[2:0] w_n3258_1;
	wire[1:0] w_n3263_0;
	wire[2:0] w_n3270_0;
	wire[1:0] w_n3271_0;
	wire[1:0] w_n3274_0;
	wire[2:0] w_n3282_0;
	wire[2:0] w_n3283_0;
	wire[2:0] w_n3283_1;
	wire[2:0] w_n3283_2;
	wire[2:0] w_n3283_3;
	wire[2:0] w_n3283_4;
	wire[2:0] w_n3283_5;
	wire[2:0] w_n3283_6;
	wire[2:0] w_n3283_7;
	wire[1:0] w_n3283_8;
	wire[2:0] w_n3284_0;
	wire[2:0] w_n3284_1;
	wire[2:0] w_n3284_2;
	wire[2:0] w_n3284_3;
	wire[2:0] w_n3284_4;
	wire[2:0] w_n3284_5;
	wire[2:0] w_n3284_6;
	wire[2:0] w_n3284_7;
	wire[2:0] w_n3284_8;
	wire[1:0] w_n3285_0;
	wire[1:0] w_n3287_0;
	wire[1:0] w_n3291_0;
	wire[1:0] w_n3294_0;
	wire[1:0] w_n3296_0;
	wire[2:0] w_n3299_0;
	wire[1:0] w_n3301_0;
	wire[2:0] w_n3302_0;
	wire[1:0] w_n3303_0;
	wire[2:0] w_n3307_0;
	wire[2:0] w_n3307_1;
	wire[2:0] w_n3314_0;
	wire[2:0] w_n3315_0;
	wire[2:0] w_n3315_1;
	wire[2:0] w_n3315_2;
	wire[2:0] w_n3315_3;
	wire[2:0] w_n3315_4;
	wire[2:0] w_n3315_5;
	wire[2:0] w_n3315_6;
	wire[2:0] w_n3315_7;
	wire[2:0] w_n3316_0;
	wire[1:0] w_n3317_0;
	wire[1:0] w_n3319_0;
	wire[2:0] w_n3320_0;
	wire[2:0] w_n3320_1;
	wire[2:0] w_n3322_0;
	wire[2:0] w_n3322_1;
	wire[2:0] w_n3322_2;
	wire[2:0] w_n3322_3;
	wire[2:0] w_n3322_4;
	wire[2:0] w_n3322_5;
	wire[2:0] w_n3322_6;
	wire[1:0] w_n3322_7;
	wire[2:0] w_n3324_0;
	wire[2:0] w_n3324_1;
	wire[1:0] w_n3324_2;
	wire[2:0] w_n3325_0;
	wire[2:0] w_n3325_1;
	wire[2:0] w_n3325_2;
	wire[2:0] w_n3325_3;
	wire[2:0] w_n3325_4;
	wire[1:0] w_n3325_5;
	wire[2:0] w_n3328_0;
	wire[2:0] w_n3328_1;
	wire[2:0] w_n3328_2;
	wire[2:0] w_n3328_3;
	wire[2:0] w_n3328_4;
	wire[2:0] w_n3328_5;
	wire[1:0] w_n3333_0;
	wire[1:0] w_n3335_0;
	wire[2:0] w_n3337_0;
	wire[2:0] w_n3337_1;
	wire[1:0] w_n3345_0;
	wire[1:0] w_n3347_0;
	wire[2:0] w_n3348_0;
	wire[2:0] w_n3349_0;
	wire[2:0] w_n3350_0;
	wire[2:0] w_n3351_0;
	wire[2:0] w_n3352_0;
	wire[2:0] w_n3353_0;
	wire[2:0] w_n3354_0;
	wire[2:0] w_n3362_0;
	wire[2:0] w_n3365_0;
	wire[2:0] w_n3367_0;
	wire[1:0] w_n3373_0;
	wire[1:0] w_n3375_0;
	wire[1:0] w_n3379_0;
	wire[1:0] w_n3394_0;
	wire[1:0] w_n3396_0;
	wire[1:0] w_n3397_0;
	wire[1:0] w_n3406_0;
	wire[1:0] w_n3408_0;
	wire[1:0] w_n3409_0;
	wire[1:0] w_n3418_0;
	wire[1:0] w_n3420_0;
	wire[1:0] w_n3421_0;
	wire[1:0] w_n3423_0;
	wire[1:0] w_n3425_0;
	wire[1:0] w_n3426_0;
	wire[1:0] w_n3435_0;
	wire[1:0] w_n3437_0;
	wire[1:0] w_n3438_0;
	wire[1:0] w_n3446_0;
	wire[1:0] w_n3452_0;
	wire[1:0] w_n3454_0;
	wire[1:0] w_n3455_0;
	wire[1:0] w_n3464_0;
	wire[1:0] w_n3466_0;
	wire[1:0] w_n3467_0;
	wire[1:0] w_n3475_0;
	wire[1:0] w_n3482_0;
	wire[1:0] w_n3484_0;
	wire[1:0] w_n3485_0;
	wire[1:0] w_n3494_0;
	wire[1:0] w_n3496_0;
	wire[1:0] w_n3497_0;
	wire[1:0] w_n3504_0;
	wire[1:0] w_n3510_0;
	wire[1:0] w_n3512_0;
	wire[1:0] w_n3513_0;
	wire[2:0] w_n3516_0;
	wire[2:0] w_n3516_1;
	wire[1:0] w_n3524_0;
	wire[1:0] w_n3528_0;
	wire[1:0] w_n3529_0;
	wire[1:0] w_n3530_0;
	wire[1:0] w_n3532_0;
	wire[1:0] w_n3535_0;
	wire[1:0] w_n3543_0;
	wire[1:0] w_n3546_0;
	wire[1:0] w_n3554_0;
	wire[1:0] w_n3557_0;
	wire[1:0] w_n3565_0;
	wire[1:0] w_n3567_0;
	wire[2:0] w_n3571_0;
	wire[1:0] w_n3571_1;
	wire[2:0] w_n3573_0;
	wire[1:0] w_n3579_0;
	wire[1:0] w_n3580_0;
	wire[1:0] w_n3581_0;
	wire[1:0] w_n3582_0;
	wire[1:0] w_n3583_0;
	wire[1:0] w_n3584_0;
	wire[1:0] w_n3585_0;
	wire[1:0] w_n3586_0;
	wire[1:0] w_n3587_0;
	wire[1:0] w_n3590_0;
	wire[1:0] w_n3591_0;
	wire[1:0] w_n3592_0;
	wire[2:0] w_n3599_0;
	wire[2:0] w_n3600_0;
	wire[2:0] w_n3600_1;
	wire[2:0] w_n3600_2;
	wire[2:0] w_n3600_3;
	wire[2:0] w_n3600_4;
	wire[2:0] w_n3600_5;
	wire[2:0] w_n3600_6;
	wire[2:0] w_n3600_7;
	wire[2:0] w_n3600_8;
	wire[2:0] w_n3601_0;
	wire[1:0] w_n3601_1;
	wire[1:0] w_n3602_0;
	wire[1:0] w_n3604_0;
	wire[2:0] w_n3605_0;
	wire[2:0] w_n3605_1;
	wire[1:0] w_n3613_0;
	wire[1:0] w_n3614_0;
	wire[1:0] w_n3615_0;
	wire[1:0] w_n3620_0;
	wire[2:0] w_n3624_0;
	wire[1:0] w_n3626_0;
	wire[1:0] w_n3630_0;
	wire[1:0] w_n3633_0;
	wire[1:0] w_n3634_0;
	wire[1:0] w_n3638_0;
	wire[1:0] w_n3650_0;
	wire[1:0] w_n3652_0;
	wire[1:0] w_n3654_0;
	wire[1:0] w_n3663_0;
	wire[1:0] w_n3666_0;
	wire[1:0] w_n3669_0;
	wire[1:0] w_n3676_0;
	wire[1:0] w_n3686_0;
	wire[2:0] w_n3693_0;
	wire[1:0] w_n3696_0;
	wire[1:0] w_n3779_0;
	wire[1:0] w_n3781_0;
	wire[1:0] w_n3784_0;
	wire[1:0] w_n3787_0;
	wire[1:0] w_n3794_0;
	wire[1:0] w_n3805_0;
	wire[2:0] w_n3806_0;
	wire[2:0] w_n3806_1;
	wire[2:0] w_n3806_2;
	wire[2:0] w_n3806_3;
	wire[2:0] w_n3806_4;
	wire[2:0] w_n3806_5;
	wire[2:0] w_n3807_0;
	wire[2:0] w_n3807_1;
	wire[2:0] w_n3807_2;
	wire[1:0] w_n3807_3;
	wire[1:0] w_n3808_0;
	wire[1:0] w_n3810_0;
	wire[2:0] w_n3811_0;
	wire[2:0] w_n3811_1;
	wire[1:0] w_n3820_0;
	wire[1:0] w_n3823_0;
	wire[1:0] w_n3826_0;
	wire[1:0] w_n3835_0;
	wire[1:0] w_n3838_0;
	wire[1:0] w_n3848_0;
	wire[1:0] w_n3849_0;
	wire[1:0] w_n3853_0;
	wire[1:0] w_n3854_0;
	wire[1:0] w_n3862_0;
	wire[1:0] w_n3863_0;
	wire[1:0] w_n3864_0;
	wire[1:0] w_n3865_0;
	wire[1:0] w_n3866_0;
	wire[1:0] w_n3874_0;
	wire[1:0] w_n3875_0;
	wire[1:0] w_n3876_0;
	wire[1:0] w_n3877_0;
	wire[1:0] w_n3878_0;
	wire[1:0] w_n3888_0;
	wire[1:0] w_n3889_0;
	wire[1:0] w_n3890_0;
	wire[1:0] w_n3891_0;
	wire[1:0] w_n3896_0;
	wire[1:0] w_n3899_0;
	wire[1:0] w_n3900_0;
	wire[1:0] w_n3902_0;
	wire[1:0] w_n3909_0;
	wire[1:0] w_n3911_0;
	wire[2:0] w_n3919_0;
	wire[2:0] w_n3919_1;
	wire[2:0] w_n3919_2;
	wire[2:0] w_n3919_3;
	wire[2:0] w_n3919_4;
	wire[2:0] w_n3919_5;
	wire[2:0] w_n3920_0;
	wire[2:0] w_n3920_1;
	wire[2:0] w_n3920_2;
	wire[1:0] w_n3920_3;
	wire[1:0] w_n3924_0;
	wire[1:0] w_n3925_0;
	wire[2:0] w_n3927_0;
	wire[2:0] w_n3927_1;
	wire[1:0] w_n3936_0;
	wire[1:0] w_n3939_0;
	wire[1:0] w_n3942_0;
	wire[1:0] w_n3951_0;
	wire[1:0] w_n3954_0;
	wire[1:0] w_n3962_0;
	wire[1:0] w_n3972_0;
	wire[1:0] w_n3973_0;
	wire[1:0] w_n3977_0;
	wire[1:0] w_n3978_0;
	wire[1:0] w_n3979_0;
	wire[1:0] w_n3980_0;
	wire[1:0] w_n3981_0;
	wire[1:0] w_n3982_0;
	wire[1:0] w_n3990_0;
	wire[1:0] w_n3991_0;
	wire[1:0] w_n3992_0;
	wire[1:0] w_n3993_0;
	wire[1:0] w_n3994_0;
	wire[2:0] w_n4000_0;
	wire[1:0] w_n4009_0;
	wire[1:0] w_n4010_0;
	wire[2:0] w_n4011_0;
	wire[2:0] w_n4013_0;
	wire[2:0] w_n4013_1;
	wire[2:0] w_n4013_2;
	wire[2:0] w_n4013_3;
	wire[2:0] w_n4013_4;
	wire[2:0] w_n4013_5;
	wire[2:0] w_n4013_6;
	wire[2:0] w_n4013_7;
	wire[2:0] w_n4013_8;
	wire[2:0] w_n4013_9;
	wire[2:0] w_n4013_10;
	wire[1:0] w_n4014_0;
	wire[1:0] w_n4017_0;
	wire[1:0] w_n4018_0;
	wire[1:0] w_n4021_0;
	wire[1:0] w_n4025_0;
	wire[1:0] w_n4028_0;
	wire[1:0] w_n4031_0;
	wire[1:0] w_n4034_0;
	wire[1:0] w_n4043_0;
	wire[1:0] w_n4046_0;
	wire[1:0] w_n4054_0;
	wire[1:0] w_n4064_0;
	wire[1:0] w_n4065_0;
	wire[1:0] w_n4069_0;
	wire[1:0] w_n4070_0;
	wire[1:0] w_n4071_0;
	wire[1:0] w_n4072_0;
	wire[1:0] w_n4073_0;
	wire[1:0] w_n4074_0;
	wire[1:0] w_n4082_0;
	wire[1:0] w_n4083_0;
	wire[1:0] w_n4084_0;
	wire[1:0] w_n4086_0;
	wire[1:0] w_n4088_0;
	wire[2:0] w_n4090_0;
	wire[2:0] w_n4090_1;
	wire[1:0] w_n4092_0;
	wire[1:0] w_n4099_0;
	wire[1:0] w_n4100_0;
	wire[1:0] w_n4101_0;
	wire[1:0] w_n4106_0;
	wire[1:0] w_n4116_0;
	wire[1:0] w_n4117_0;
	wire[1:0] w_n4118_0;
	wire[1:0] w_n4119_0;
	wire[1:0] w_n4120_0;
	wire[1:0] w_n4123_0;
	wire[1:0] w_n4125_0;
	wire[1:0] w_n4129_0;
	wire[1:0] w_n4132_0;
	wire[1:0] w_n4135_0;
	wire[2:0] w_n4136_0;
	wire[2:0] w_n4136_1;
	wire[1:0] w_n4141_0;
	wire[1:0] w_n4144_0;
	wire[1:0] w_n4153_0;
	wire[1:0] w_n4156_0;
	wire[1:0] w_n4164_0;
	wire[1:0] w_n4172_0;
	wire[1:0] w_n4173_0;
	wire[1:0] w_n4177_0;
	wire[1:0] w_n4178_0;
	wire[1:0] w_n4179_0;
	wire[1:0] w_n4180_0;
	wire[1:0] w_n4181_0;
	wire[1:0] w_n4182_0;
	wire[1:0] w_n4190_0;
	wire[1:0] w_n4191_0;
	wire[1:0] w_n4192_0;
	wire[1:0] w_n4193_0;
	wire[1:0] w_n4194_0;
	wire[1:0] w_n4206_0;
	wire[1:0] w_n4207_0;
	wire[1:0] w_n4208_0;
	wire[1:0] w_n4209_0;
	wire[1:0] w_n4211_0;
	wire[1:0] w_n4215_0;
	wire[1:0] w_n4218_0;
	wire[1:0] w_n4221_0;
	wire[1:0] w_n4224_0;
	wire[1:0] w_n4233_0;
	wire[1:0] w_n4236_0;
	wire[1:0] w_n4245_0;
	wire[1:0] w_n4246_0;
	wire[1:0] w_n4247_0;
	wire[1:0] w_n4248_0;
	wire[1:0] w_n4253_0;
	wire[1:0] w_n4254_0;
	wire[1:0] w_n4262_0;
	wire[1:0] w_n4263_0;
	wire[1:0] w_n4264_0;
	wire[1:0] w_n4265_0;
	wire[1:0] w_n4266_0;
	wire[1:0] w_n4274_0;
	wire[1:0] w_n4275_0;
	wire[1:0] w_n4276_0;
	wire[1:0] w_n4277_0;
	wire[1:0] w_n4286_0;
	wire[1:0] w_n4287_0;
	wire[1:0] w_n4288_0;
	wire[1:0] w_n4289_0;
	wire[1:0] w_n4290_0;
	wire[1:0] w_n4293_0;
	wire[1:0] w_n4297_0;
	wire[1:0] w_n4300_0;
	wire[1:0] w_n4303_0;
	wire[1:0] w_n4309_0;
	wire[1:0] w_n4312_0;
	wire[1:0] w_n4321_0;
	wire[1:0] w_n4324_0;
	wire[1:0] w_n4332_0;
	wire[1:0] w_n4340_0;
	wire[1:0] w_n4343_0;
	wire[1:0] w_n4344_0;
	wire[1:0] w_n4345_0;
	wire[1:0] w_n4346_0;
	wire[1:0] w_n4347_0;
	wire[1:0] w_n4348_0;
	wire[1:0] w_n4349_0;
	wire[1:0] w_n4350_0;
	wire[1:0] w_n4351_0;
	wire[1:0] w_n4352_0;
	wire[1:0] w_n4353_0;
	wire[1:0] w_n4354_0;
	wire[1:0] w_n4355_0;
	wire[2:0] w_n4357_0;
	wire[1:0] w_n4368_0;
	wire[1:0] w_n4369_0;
	wire[1:0] w_n4370_0;
	wire[1:0] w_n4371_0;
	wire[1:0] w_n4372_0;
	wire[1:0] w_n4375_0;
	wire[1:0] w_n4379_0;
	wire[1:0] w_n4382_0;
	wire[1:0] w_n4385_0;
	wire[1:0] w_n4389_0;
	wire[1:0] w_n4393_0;
	wire[1:0] w_n4394_0;
	wire[1:0] w_n4403_0;
	wire[1:0] w_n4406_0;
	wire[1:0] w_n4414_0;
	wire[1:0] w_n4422_0;
	wire[1:0] w_n4425_0;
	wire[1:0] w_n4426_0;
	wire[1:0] w_n4427_0;
	wire[1:0] w_n4428_0;
	wire[1:0] w_n4429_0;
	wire[1:0] w_n4430_0;
	wire[1:0] w_n4431_0;
	wire[1:0] w_n4432_0;
	wire[1:0] w_n4433_0;
	wire[1:0] w_n4434_0;
	wire[1:0] w_n4435_0;
	wire[1:0] w_n4442_0;
	wire[1:0] w_n4450_0;
	wire[1:0] w_n4451_0;
	wire[1:0] w_n4452_0;
	wire[1:0] w_n4453_0;
	wire[1:0] w_n4454_0;
	wire[1:0] w_n4457_0;
	wire[1:0] w_n4461_0;
	wire[1:0] w_n4464_0;
	wire[1:0] w_n4469_0;
	wire[1:0] w_n4472_0;
	wire[1:0] w_n4480_0;
	wire[1:0] w_n4481_0;
	wire[1:0] w_n4484_0;
	wire[1:0] w_n4487_0;
	wire[1:0] w_n4496_0;
	wire[1:0] w_n4497_0;
	wire[1:0] w_n4498_0;
	wire[1:0] w_n4499_0;
	wire[1:0] w_n4500_0;
	wire[1:0] w_n4501_0;
	wire[1:0] w_n4509_0;
	wire[1:0] w_n4510_0;
	wire[1:0] w_n4511_0;
	wire[1:0] w_n4512_0;
	wire[1:0] w_n4513_0;
	wire[1:0] w_n4514_0;
	wire[1:0] w_n4523_0;
	wire[1:0] w_n4524_0;
	wire[1:0] w_n4525_0;
	wire[1:0] w_n4526_0;
	wire[1:0] w_n4527_0;
	wire[1:0] w_n4530_0;
	wire[1:0] w_n4534_0;
	wire[1:0] w_n4537_0;
	wire[1:0] w_n4540_0;
	wire[1:0] w_n4547_0;
	wire[1:0] w_n4550_0;
	wire[1:0] w_n4558_0;
	wire[1:0] w_n4561_0;
	wire[1:0] w_n4569_0;
	wire[1:0] w_n4570_0;
	wire[2:0] w_n4571_0;
	wire[1:0] w_n4574_0;
	wire[1:0] w_n4575_0;
	wire[1:0] w_n4576_0;
	wire[1:0] w_n4577_0;
	wire[1:0] w_n4578_0;
	wire[1:0] w_n4579_0;
	wire[1:0] w_n4580_0;
	wire[1:0] w_n4581_0;
	wire[1:0] w_n4582_0;
	wire[1:0] w_n4589_0;
	wire[1:0] w_n4599_0;
	wire[1:0] w_n4600_0;
	wire[1:0] w_n4601_0;
	wire[1:0] w_n4602_0;
	wire[1:0] w_n4603_0;
	wire[1:0] w_n4606_0;
	wire[1:0] w_n4610_0;
	wire[1:0] w_n4613_0;
	wire[1:0] w_n4616_0;
	wire[1:0] w_n4620_0;
	wire[1:0] w_n4624_0;
	wire[1:0] w_n4625_0;
	wire[1:0] w_n4628_0;
	wire[1:0] w_n4636_0;
	wire[1:0] w_n4637_0;
	wire[1:0] w_n4638_0;
	wire[1:0] w_n4639_0;
	wire[1:0] w_n4647_0;
	wire[1:0] w_n4648_0;
	wire[1:0] w_n4649_0;
	wire[1:0] w_n4650_0;
	wire[1:0] w_n4651_0;
	wire[1:0] w_n4663_0;
	wire[1:0] w_n4664_0;
	wire[1:0] w_n4665_0;
	wire[1:0] w_n4666_0;
	wire[1:0] w_n4667_0;
	wire[1:0] w_n4670_0;
	wire[1:0] w_n4674_0;
	wire[1:0] w_n4677_0;
	wire[1:0] w_n4682_0;
	wire[1:0] w_n4685_0;
	wire[1:0] w_n4693_0;
	wire[1:0] w_n4694_0;
	wire[1:0] w_n4703_0;
	wire[2:0] w_n4704_0;
	wire[2:0] w_n4706_0;
	wire[2:0] w_n4711_0;
	wire[1:0] w_n4713_0;
	wire[1:0] w_n4714_0;
	wire[1:0] w_n4715_0;
	wire[1:0] w_n4716_0;
	wire[1:0] w_n4728_0;
	wire[1:0] w_n4729_0;
	wire[1:0] w_n4730_0;
	wire[1:0] w_n4731_0;
	wire[1:0] w_n4732_0;
	wire[1:0] w_n4735_0;
	wire[1:0] w_n4739_0;
	wire[1:0] w_n4742_0;
	wire[1:0] w_n4745_0;
	wire[1:0] w_n4751_0;
	wire[1:0] w_n4759_0;
	wire[2:0] w_n4760_0;
	wire[1:0] w_n4766_0;
	wire[1:0] w_n4767_0;
	wire[1:0] w_n4768_0;
	wire[1:0] w_n4775_0;
	wire[1:0] w_n4776_0;
	wire[1:0] w_n4777_0;
	wire[1:0] w_n4778_0;
	wire[1:0] w_n4779_0;
	wire[1:0] w_n4785_0;
	wire[1:0] w_n4786_0;
	wire[1:0] w_n4787_0;
	wire[1:0] w_n4788_0;
	wire[1:0] w_n4789_0;
	wire[1:0] w_n4792_0;
	wire[1:0] w_n4796_0;
	wire[1:0] w_n4799_0;
	wire[1:0] w_n4802_0;
	wire[1:0] w_n4806_0;
	wire[1:0] w_n4807_0;
	wire[1:0] w_n4808_0;
	wire[1:0] w_n4816_0;
	wire[1:0] w_n4820_0;
	wire[1:0] w_n4821_0;
	wire[1:0] w_n4822_0;
	wire[1:0] w_n4823_0;
	wire[1:0] w_n4824_0;
	wire[1:0] w_n4832_0;
	wire[1:0] w_n4836_0;
	wire[1:0] w_n4837_0;
	wire[1:0] w_n4838_0;
	wire[1:0] w_n4839_0;
	wire[1:0] w_n4840_0;
	wire[1:0] w_n4843_0;
	wire[1:0] w_n4847_0;
	wire[1:0] w_n4850_0;
	wire[1:0] w_n4855_0;
	wire[1:0] w_n4859_0;
	wire[1:0] w_n4868_0;
	wire[1:0] w_n4869_0;
	wire[1:0] w_n4870_0;
	wire[1:0] w_n4871_0;
	wire[1:0] w_n4872_0;
	wire[1:0] w_n4873_0;
	wire[1:0] w_n4874_0;
	wire[1:0] w_n4875_0;
	wire[1:0] w_n4876_0;
	wire[1:0] w_n4880_0;
	wire[1:0] w_n4892_0;
	wire[1:0] w_n4893_0;
	wire[1:0] w_n4894_0;
	wire[1:0] w_n4895_0;
	wire[1:0] w_n4896_0;
	wire[1:0] w_n4899_0;
	wire[1:0] w_n4903_0;
	wire[1:0] w_n4906_0;
	wire[1:0] w_n4909_0;
	wire[1:0] w_n4915_0;
	wire[1:0] w_n4917_0;
	wire[1:0] w_n4920_0;
	wire[1:0] w_n4921_0;
	wire[1:0] w_n4922_0;
	wire[1:0] w_n4923_0;
	wire[1:0] w_n4924_0;
	wire[1:0] w_n4931_0;
	wire[1:0] w_n4939_0;
	wire[1:0] w_n4940_0;
	wire[1:0] w_n4941_0;
	wire[1:0] w_n4942_0;
	wire[1:0] w_n4943_0;
	wire[1:0] w_n4946_0;
	wire[1:0] w_n4950_0;
	wire[1:0] w_n4953_0;
	wire[1:0] w_n4957_0;
	wire[1:0] w_n4959_0;
	wire[1:0] w_n4960_0;
	wire[1:0] w_n4964_0;
	wire[1:0] w_n4965_0;
	wire[1:0] w_n4968_0;
	wire[1:0] w_n4969_0;
	wire[1:0] w_n4972_0;
	wire[1:0] w_n4982_0;
	wire[1:0] w_n4983_0;
	wire[1:0] w_n4984_0;
	wire[1:0] w_n4985_0;
	wire[1:0] w_n4986_0;
	wire[1:0] w_n4989_0;
	wire[1:0] w_n4993_0;
	wire[1:0] w_n4994_0;
	wire[2:0] w_n5003_0;
	wire[1:0] w_n5007_0;
	wire[1:0] w_n5016_0;
	wire[1:0] w_n5017_0;
	wire[1:0] w_n5018_0;
	wire[1:0] w_n5019_0;
	wire[1:0] w_n5020_0;
	wire[1:0] w_n5021_0;
	wire[2:0] w_n5024_0;
	wire[2:0] w_n5026_0;
	wire[1:0] w_n5027_0;
	wire[1:0] w_n5031_0;
	wire[2:0] w_n5042_0;
	wire[1:0] w_n5042_1;
	wire[2:0] w_n5043_0;
	wire[1:0] w_n5044_0;
	wire[1:0] w_n5046_0;
	wire[1:0] w_n5048_0;
	wire[1:0] w_n5050_0;
	wire[1:0] w_n5054_0;
	wire[1:0] w_n5056_0;
	wire[1:0] w_n5057_0;
	wire[1:0] w_n5058_0;
	wire[2:0] w_n5068_0;
	wire[1:0] w_n5068_1;
	wire[1:0] w_n5069_0;
	wire[2:0] w_n5081_0;
	wire[1:0] w_n5082_0;
	wire[2:0] w_n5083_0;
	wire[2:0] w_n5084_0;
	wire[1:0] w_n5085_0;
	wire[1:0] w_n5088_0;
	wire[1:0] w_n5091_0;
	wire[1:0] w_n5092_0;
	wire[1:0] w_n5095_0;
	wire[1:0] w_n5098_0;
	wire[1:0] w_n5099_0;
	wire[1:0] w_n5100_0;
	wire[2:0] w_n5109_0;
	wire[1:0] w_n5110_0;
	wire[2:0] w_n5112_0;
	wire[2:0] w_n5113_0;
	wire[1:0] w_n5116_0;
	wire[1:0] w_n5117_0;
	wire[1:0] w_n5118_0;
	wire[2:0] w_n5119_0;
	wire[1:0] w_n5120_0;
	wire[1:0] w_n5123_0;
	wire[1:0] w_n5126_0;
	wire[1:0] w_n5128_0;
	wire[1:0] w_n5129_0;
	wire[1:0] w_n5130_0;
	wire[1:0] w_n5132_0;
	wire[1:0] w_n5133_0;
	wire[1:0] w_n5137_0;
	wire[1:0] w_n5138_0;
	wire[1:0] w_n5140_0;
	wire[1:0] w_n5142_0;
	wire w_dff_A_RiPtSZDk9_1;
	wire w_dff_A_NGXHeKO55_0;
	wire w_dff_A_37IA4n3O4_0;
	wire w_dff_A_4OtQlOja2_0;
	wire w_dff_A_TpbVPwI53_0;
	wire w_dff_A_kpphw58F3_0;
	wire w_dff_A_vlPZ0Ent8_1;
	wire w_dff_A_UoKBhK4Y5_1;
	wire w_dff_A_Hx1Ouz7H2_1;
	wire w_dff_A_MZ7mXmkf2_0;
	wire w_dff_A_sF759xAa4_0;
	wire w_dff_A_gKWP81xO2_0;
	wire w_dff_A_s4kVgoWW2_0;
	wire w_dff_A_71ea6gqc1_1;
	wire w_dff_A_ucqtqfZU9_1;
	wire w_dff_A_z1uSxqiA1_0;
	wire w_dff_A_5FLG8NpT4_0;
	wire w_dff_A_PyH5QJbQ1_0;
	wire w_dff_A_VEC9hgaD8_0;
	wire w_dff_A_VBobKaBi6_1;
	wire w_dff_A_TV7kAWfk8_1;
	wire w_dff_A_GJdWBh692_0;
	wire w_dff_A_kVOWvjKY5_0;
	wire w_dff_A_aOryP3WK4_0;
	wire w_dff_A_GJdM5i5M9_0;
	wire w_dff_A_wQjDLugB6_1;
	wire w_dff_A_hKKpVgtY8_1;
	wire w_dff_A_GbhPl4H60_0;
	wire w_dff_A_HxOgasBy2_0;
	wire w_dff_A_B0Y8cdCP8_0;
	wire w_dff_A_pLKYVyp88_0;
	wire w_dff_A_EkEHmc8d2_0;
	wire w_dff_A_LkUnTVjy1_0;
	wire w_dff_A_a1aj6vRM7_0;
	wire w_dff_A_pZnZyIvF9_0;
	wire w_dff_A_9hCSOo2w9_0;
	wire w_dff_A_ZsQ6Rmqk2_0;
	wire w_dff_A_IUPVafqv2_0;
	wire w_dff_A_zFz06Ms96_0;
	wire w_dff_A_c1FXsuoM0_1;
	wire w_dff_A_s4A9eYcR0_1;
	wire w_dff_A_QopHYMRW9_1;
	wire w_dff_A_h7oPp7wq6_1;
	wire w_dff_A_ApGqMT1D4_1;
	wire w_dff_A_bJB9Q22H3_1;
	wire w_dff_A_rbEHx83I3_0;
	wire w_dff_A_DgJBwDXc8_0;
	wire w_dff_A_EtaMr0GE0_0;
	wire w_dff_A_wMefoSvl1_0;
	wire w_dff_A_uAUH7fgJ9_1;
	wire w_dff_A_dBDyGrTJ0_1;
	wire w_dff_B_eZEzychJ4_0;
	wire w_dff_A_RBDOLeeS2_0;
	wire w_dff_A_m2X92ovI5_0;
	wire w_dff_A_bZ09vicW3_0;
	wire w_dff_B_5RI4xp2g0_2;
	wire w_dff_B_dhiVQU502_2;
	wire w_dff_B_jcaxrZF74_2;
	wire w_dff_B_w3sdJIzj0_2;
	wire w_dff_B_BAThx7lY3_2;
	wire w_dff_B_riTWdShy8_2;
	wire w_dff_B_ULl67ORI8_2;
	wire w_dff_B_MXVV6Kuo8_2;
	wire w_dff_B_yGx9f0w05_2;
	wire w_dff_B_Qr16cTJg6_2;
	wire w_dff_B_mCu6o7Is6_2;
	wire w_dff_B_YLo8Csg21_2;
	wire w_dff_B_VK4p86qM3_2;
	wire w_dff_B_sWi4cVC18_2;
	wire w_dff_B_XwE082Vg1_2;
	wire w_dff_B_Eu7QGMNU6_2;
	wire w_dff_B_icLouTRe3_2;
	wire w_dff_B_JCU59h5a4_2;
	wire w_dff_B_jlC6hA1j8_2;
	wire w_dff_B_cBNuyFzy2_2;
	wire w_dff_B_Y9FVxNhB9_2;
	wire w_dff_B_o6QWkKQA0_2;
	wire w_dff_B_EydgXy3w4_2;
	wire w_dff_B_m3IjCvmS5_2;
	wire w_dff_B_jup1g00q9_2;
	wire w_dff_B_PUkG8ZRw4_2;
	wire w_dff_B_wgMSX9l29_2;
	wire w_dff_B_A71ehwnI3_2;
	wire w_dff_B_XZV6JPhW1_2;
	wire w_dff_B_qlKAxEia2_2;
	wire w_dff_B_gvL5aKzK1_2;
	wire w_dff_B_CsliOohJ7_2;
	wire w_dff_B_G6YBppBM0_2;
	wire w_dff_B_ZzJf2LJC4_2;
	wire w_dff_B_WEHirB0f9_2;
	wire w_dff_B_OzwR54au9_2;
	wire w_dff_B_Exl1FNYz6_2;
	wire w_dff_B_9k2eQFIa7_2;
	wire w_dff_B_2VstCvap2_2;
	wire w_dff_B_uBVkdo3C0_2;
	wire w_dff_B_s1VBUl6w1_2;
	wire w_dff_B_Qa9YHEfh9_2;
	wire w_dff_B_MgMvnRTs0_2;
	wire w_dff_B_Vg5ZcwMW4_2;
	wire w_dff_B_GK3MlLa02_2;
	wire w_dff_B_3J0Az0Tj9_2;
	wire w_dff_B_iJMDOdGD0_2;
	wire w_dff_B_3Y6m6eYG7_2;
	wire w_dff_B_5kGmypLt0_2;
	wire w_dff_B_bmvoXJ8M9_2;
	wire w_dff_B_NQNAA8pr0_2;
	wire w_dff_B_vxJaR31t8_2;
	wire w_dff_B_Wxo4ZPjh9_2;
	wire w_dff_B_rj1wjVlq7_2;
	wire w_dff_B_ZR1DnZ4i9_2;
	wire w_dff_B_OCgBxrtb4_2;
	wire w_dff_B_X9TYsqmO2_2;
	wire w_dff_B_ottB5zyD7_2;
	wire w_dff_B_eWTgTqtM5_2;
	wire w_dff_B_pTRErxPb5_2;
	wire w_dff_B_Milp0czy0_2;
	wire w_dff_B_7yseujS22_2;
	wire w_dff_B_sw3dxI9g4_2;
	wire w_dff_B_fz22z2qR1_2;
	wire w_dff_B_Gt05YMW87_2;
	wire w_dff_B_HEL5L0zz2_2;
	wire w_dff_B_TMjOVxqT5_2;
	wire w_dff_B_KcW4lYA00_2;
	wire w_dff_B_fuyAr6Pq3_2;
	wire w_dff_B_44woTVgy3_2;
	wire w_dff_B_KDKBNM6v0_2;
	wire w_dff_B_1E3aRSXX0_2;
	wire w_dff_B_TISKl5955_2;
	wire w_dff_B_Jyxz7DFM1_2;
	wire w_dff_B_3sRop2Ie6_2;
	wire w_dff_B_y7ccUvVH1_2;
	wire w_dff_B_UFNe7O7N9_2;
	wire w_dff_B_NJFkvd9n3_2;
	wire w_dff_B_O9A2viQI7_2;
	wire w_dff_B_OhJT1iyq9_2;
	wire w_dff_B_FaBiW03U2_2;
	wire w_dff_B_5j6zucTg2_2;
	wire w_dff_B_i20OsPjB8_2;
	wire w_dff_B_Rs7NWEAE4_2;
	wire w_dff_B_QP4PSIAd5_2;
	wire w_dff_B_AftEnVhu8_2;
	wire w_dff_B_AM5Bs5ur0_2;
	wire w_dff_B_TmSKnfvk0_2;
	wire w_dff_B_Le8JZY4E5_2;
	wire w_dff_B_PLHNxj171_2;
	wire w_dff_B_fkiWHb5z7_2;
	wire w_dff_B_wsJydkto0_2;
	wire w_dff_B_9cKC052I7_2;
	wire w_dff_B_KOsJ800c0_2;
	wire w_dff_B_SufTqADf2_2;
	wire w_dff_B_ETFt5nf87_2;
	wire w_dff_B_q5szTSDk8_2;
	wire w_dff_B_awuJZjRy1_2;
	wire w_dff_B_NaRMWG1q4_2;
	wire w_dff_B_houcbZNh6_2;
	wire w_dff_B_pcKV86BE1_2;
	wire w_dff_B_AzKsezPA4_2;
	wire w_dff_B_vxaNRlZp0_2;
	wire w_dff_B_yiPpV30k0_2;
	wire w_dff_B_8qirCfdf9_2;
	wire w_dff_B_vQ1IGsp82_2;
	wire w_dff_B_LAmnM0vh0_2;
	wire w_dff_B_FUdmWInD1_2;
	wire w_dff_B_Ryt8C1hJ5_2;
	wire w_dff_B_VYJQqXnf0_2;
	wire w_dff_B_LxKP9G961_2;
	wire w_dff_B_PigctOHU8_2;
	wire w_dff_B_MH55XeHM6_2;
	wire w_dff_B_yHPASRXz5_2;
	wire w_dff_B_0LaGRlav8_2;
	wire w_dff_B_6mfeIp3z0_2;
	wire w_dff_B_yD7dkkhi9_2;
	wire w_dff_B_LQiHz9fy5_2;
	wire w_dff_B_uEyTSu8O3_2;
	wire w_dff_B_cHfGK3wW5_2;
	wire w_dff_B_KjLceTJ15_2;
	wire w_dff_B_Fx4HYKGK9_2;
	wire w_dff_B_QcR9J9D45_2;
	wire w_dff_B_CWSG3c6X3_2;
	wire w_dff_B_FYi19mux6_2;
	wire w_dff_B_UGfytwYE5_2;
	wire w_dff_B_fTmfuLci5_2;
	wire w_dff_B_wgwNlq0s6_2;
	wire w_dff_B_B9hxklVT5_2;
	wire w_dff_B_H1CEOAzK2_2;
	wire w_dff_B_yQCmSbu72_2;
	wire w_dff_B_xkNf9owQ5_2;
	wire w_dff_B_PNEGI4yT5_2;
	wire w_dff_B_fJ7zhDrm9_2;
	wire w_dff_B_46lDhABu1_2;
	wire w_dff_B_qgr76Lbj5_2;
	wire w_dff_B_1a890rbd8_2;
	wire w_dff_B_YkOE5CkR1_2;
	wire w_dff_B_qL6rScVZ8_2;
	wire w_dff_B_4CHZKSur9_2;
	wire w_dff_B_BeYRFeNT9_2;
	wire w_dff_B_FEK6rsfi1_2;
	wire w_dff_B_0bWCEVVm3_2;
	wire w_dff_B_gd2Mccjr1_2;
	wire w_dff_B_vnp5ZE708_2;
	wire w_dff_B_yCAK8FC23_2;
	wire w_dff_B_nPPCaf1Q4_2;
	wire w_dff_B_Gw348KKn2_2;
	wire w_dff_B_ysrD9GaZ8_2;
	wire w_dff_B_Zm7EjNgg7_2;
	wire w_dff_B_YYcRPf0b8_2;
	wire w_dff_B_CtoyzuH37_2;
	wire w_dff_B_1Q9Go4ez0_2;
	wire w_dff_B_iL8QFOMo9_2;
	wire w_dff_B_5eDBnhxR4_2;
	wire w_dff_B_mIQBAR6E9_2;
	wire w_dff_B_wcw2K1gk7_2;
	wire w_dff_A_mEdyEIrL5_0;
	wire w_dff_A_Bw0aCnDm9_0;
	wire w_dff_A_b6PhEX3p8_0;
	wire w_dff_A_ypy0WxOY7_1;
	wire w_dff_A_QWOvLrxd2_1;
	wire w_dff_A_GY2RnPJc4_1;
	wire w_dff_A_WhFlsVOj3_1;
	wire w_dff_B_2rz4dWGZ7_1;
	wire w_dff_A_B735v1Ea2_1;
	wire w_dff_B_OP6iqswc4_1;
	wire w_dff_A_h2PYpQyn7_0;
	wire w_dff_A_EohMCOr02_1;
	wire w_dff_A_N6sxVGld7_1;
	wire w_dff_B_kKOZmqN48_2;
	wire w_dff_B_7rDoO9sx7_2;
	wire w_dff_B_CeDtLGO62_2;
	wire w_dff_B_DzGFTP3B4_2;
	wire w_dff_B_g2D3wdph1_2;
	wire w_dff_B_zcOhCS2a8_2;
	wire w_dff_B_B8QSZ5Zm7_2;
	wire w_dff_B_yDTR2Y3x7_2;
	wire w_dff_B_nlmpukMG7_2;
	wire w_dff_B_ANgszXzq4_2;
	wire w_dff_B_lKfhn1IJ8_2;
	wire w_dff_B_0TJPPYYb2_2;
	wire w_dff_B_4uDgwDES3_2;
	wire w_dff_B_KCex5Kn38_2;
	wire w_dff_B_8QGrpRFt9_2;
	wire w_dff_B_PDW74LMp1_2;
	wire w_dff_B_AJj62i627_2;
	wire w_dff_B_BIBiy4dV7_2;
	wire w_dff_B_oRiamI7y5_2;
	wire w_dff_B_Fudaf5rG0_2;
	wire w_dff_B_7uJfallg2_2;
	wire w_dff_B_6RnCNS9P7_2;
	wire w_dff_B_HyMnj4nP1_2;
	wire w_dff_B_3XFrlSPU0_2;
	wire w_dff_B_r5j9ZkxA8_2;
	wire w_dff_B_73cJfVwZ1_2;
	wire w_dff_B_tyBm301x7_2;
	wire w_dff_B_xBaAXZT70_2;
	wire w_dff_B_AuhgSYuF1_2;
	wire w_dff_B_i6hB622j1_2;
	wire w_dff_B_o0qEQHwN2_2;
	wire w_dff_B_qpojBUg34_2;
	wire w_dff_B_v3nsYcVk8_2;
	wire w_dff_B_IL6YDOLP7_2;
	wire w_dff_B_W9idEL0R0_2;
	wire w_dff_B_rwQv5M8l5_2;
	wire w_dff_B_039ssV2g5_2;
	wire w_dff_B_2tKs1Km07_2;
	wire w_dff_B_KjNMdo2c6_2;
	wire w_dff_B_2JwdyTnF4_2;
	wire w_dff_B_83U5kNYX4_2;
	wire w_dff_B_eRRRpXIp0_2;
	wire w_dff_B_IVmAjTV78_2;
	wire w_dff_B_gwNpEnUi9_2;
	wire w_dff_B_qQtLCcZW8_2;
	wire w_dff_B_US5NXbHh4_2;
	wire w_dff_B_stTWBR3N5_2;
	wire w_dff_B_G3VAygMi9_2;
	wire w_dff_B_iK4WsCJd2_2;
	wire w_dff_B_ROPJrve65_2;
	wire w_dff_B_9niJIMgr0_2;
	wire w_dff_B_EdPmcdeZ2_2;
	wire w_dff_B_rFZjnwEp4_2;
	wire w_dff_B_BIhyteCr6_2;
	wire w_dff_B_WIVEVmRH9_2;
	wire w_dff_B_sM6oXN572_2;
	wire w_dff_B_rNzDtf1p1_2;
	wire w_dff_B_wYEHWQGJ7_2;
	wire w_dff_B_R32K0NNh2_2;
	wire w_dff_B_aqMaFA1e4_2;
	wire w_dff_B_fwWN6pFr6_2;
	wire w_dff_B_5LmGhSp79_2;
	wire w_dff_B_8vziuG1U6_2;
	wire w_dff_B_lTvL2yLB7_2;
	wire w_dff_B_bLrpStSI8_2;
	wire w_dff_B_e2mE2qLA2_2;
	wire w_dff_B_f3mcrV686_2;
	wire w_dff_B_nqXoUMTE8_2;
	wire w_dff_B_KjwFphHi1_2;
	wire w_dff_B_wz9CJPBy5_2;
	wire w_dff_B_FidPeKuk3_2;
	wire w_dff_B_dt1fWUPw1_2;
	wire w_dff_B_NIFoP6fq5_2;
	wire w_dff_B_9Pn1QdBa0_2;
	wire w_dff_B_Mwdr0ex54_2;
	wire w_dff_B_kehcM6Nf6_2;
	wire w_dff_B_5VJFioyt2_2;
	wire w_dff_B_nVuxINDG6_2;
	wire w_dff_B_0dhcWmTo6_2;
	wire w_dff_B_9KcLHECc0_2;
	wire w_dff_B_USHaZjdi7_2;
	wire w_dff_B_G5BEgudb6_2;
	wire w_dff_B_KgmKOHcP4_2;
	wire w_dff_B_arB0yoaU3_2;
	wire w_dff_B_60rVC1rb0_2;
	wire w_dff_B_pu4gjLdZ1_2;
	wire w_dff_B_P27OR78m7_2;
	wire w_dff_B_IN61Kn5F7_2;
	wire w_dff_B_x2hBgIs82_2;
	wire w_dff_B_5H9dfX1j9_2;
	wire w_dff_B_nnpwLxU44_2;
	wire w_dff_B_sCNFtcAp6_2;
	wire w_dff_B_l6vTRmli8_2;
	wire w_dff_B_eztTHDde1_2;
	wire w_dff_B_3OrDKUJj0_2;
	wire w_dff_B_CsiPZSAa2_2;
	wire w_dff_B_A3V6HJoQ5_2;
	wire w_dff_B_ZfCni8gI2_2;
	wire w_dff_B_RXClBM164_2;
	wire w_dff_B_des7wfFf4_2;
	wire w_dff_B_wZOj33dQ6_2;
	wire w_dff_B_IZsVzRmh2_2;
	wire w_dff_B_Q1a9kF4g0_2;
	wire w_dff_B_2dB8pYrl2_2;
	wire w_dff_B_5VfWGz4r1_2;
	wire w_dff_B_jekYDuP48_2;
	wire w_dff_B_DPSlNoRU3_2;
	wire w_dff_B_UaVO9muF5_2;
	wire w_dff_B_XY4keW9r7_2;
	wire w_dff_B_PMzv3sup1_2;
	wire w_dff_B_MZZPo2KJ3_2;
	wire w_dff_B_ZcgGVSla1_2;
	wire w_dff_B_CSnHakR16_2;
	wire w_dff_B_WopNUl880_2;
	wire w_dff_B_kpt5IzMd0_2;
	wire w_dff_B_qTnEM4Pf4_2;
	wire w_dff_B_29I4CNV09_2;
	wire w_dff_B_uO0oUmgB6_2;
	wire w_dff_B_tDJHiKPo9_2;
	wire w_dff_B_4qVYnJ1F4_2;
	wire w_dff_B_xXAtKyuR3_2;
	wire w_dff_B_uISo6LVc5_2;
	wire w_dff_B_IoTRuWhs9_2;
	wire w_dff_B_fouTRMzq4_2;
	wire w_dff_B_upVwaqff9_2;
	wire w_dff_B_9K6zKB0w6_2;
	wire w_dff_B_RdJkpfpH4_2;
	wire w_dff_B_zUuRNuqY6_2;
	wire w_dff_B_TemKBV990_2;
	wire w_dff_B_TeEVRnbd9_2;
	wire w_dff_B_8hC2alfW9_2;
	wire w_dff_B_G9uczfGb9_2;
	wire w_dff_B_IPG6jWwi7_2;
	wire w_dff_B_RTxZitcs4_2;
	wire w_dff_B_7ujJIy5n9_2;
	wire w_dff_B_9RaeZEvG0_2;
	wire w_dff_B_xRMqeGPe7_2;
	wire w_dff_B_stWHUBP12_2;
	wire w_dff_B_OWlWKqxz0_2;
	wire w_dff_B_5SXokDAm3_2;
	wire w_dff_B_9U6RuGSZ9_2;
	wire w_dff_B_J653GGjn7_2;
	wire w_dff_B_389mS7mG7_2;
	wire w_dff_B_d9hBrptt6_0;
	wire w_dff_A_OaMuw6Hb9_1;
	wire w_dff_B_4LMWvph54_1;
	wire w_dff_A_Xhuy3IJF7_0;
	wire w_dff_A_awo5l0ir3_0;
	wire w_dff_A_HPuTasns0_0;
	wire w_dff_A_wxzz2WBi3_0;
	wire w_dff_A_e94k11f77_0;
	wire w_dff_A_yIbGSoVr3_0;
	wire w_dff_A_sOErIqr07_0;
	wire w_dff_A_fGY52gbv0_0;
	wire w_dff_A_72JVXFet2_0;
	wire w_dff_A_J0qwBfzZ9_0;
	wire w_dff_A_h9g6HZkd4_0;
	wire w_dff_A_SMxcsPby6_0;
	wire w_dff_A_gjRzRkwI1_0;
	wire w_dff_A_t9pi2k7w5_0;
	wire w_dff_A_uVwNu9Rb1_0;
	wire w_dff_A_vDPcnB1Q5_0;
	wire w_dff_A_l5ALSQ9k4_0;
	wire w_dff_A_UK3GPCLL0_0;
	wire w_dff_A_Op0hX5fq0_0;
	wire w_dff_A_W48FiSy24_1;
	wire w_dff_B_elMsNUXc0_2;
	wire w_dff_A_lr3QEvLc2_1;
	wire w_dff_B_QvlyzZXy5_2;
	wire w_dff_A_UKMe566N2_1;
	wire w_dff_A_fx7a37RG8_1;
	wire w_dff_A_FN0f6bzQ8_1;
	wire w_dff_A_o1vAK5iq7_1;
	wire w_dff_A_nBj4kGVC4_1;
	wire w_dff_A_jzz1ksPd0_1;
	wire w_dff_A_2BWMdtY83_1;
	wire w_dff_A_xcEohffX4_1;
	wire w_dff_A_C2jk7L929_1;
	wire w_dff_A_jFPvwqMJ4_1;
	wire w_dff_A_dWFmD96g4_1;
	wire w_dff_A_itrUM3iV6_1;
	wire w_dff_A_ECp7BdkB5_1;
	wire w_dff_A_YkCbqYno9_1;
	wire w_dff_A_onfvbgBw3_1;
	wire w_dff_A_hngeokM71_1;
	wire w_dff_A_s9ntx8NO3_1;
	wire w_dff_A_qzWxn6461_1;
	wire w_dff_A_ut645Deh1_1;
	wire w_dff_A_V7hMOjCO9_1;
	wire w_dff_A_YIRDUDk07_1;
	wire w_dff_A_gVYHnMqv1_1;
	wire w_dff_A_fTytwo4O6_1;
	wire w_dff_A_z38fvWZc0_1;
	wire w_dff_A_Vzxv9Uwi8_1;
	wire w_dff_A_rmUArDBM2_1;
	wire w_dff_A_p1UN0wUm4_1;
	wire w_dff_A_RyfUTes05_1;
	wire w_dff_A_SZhjyTSy6_1;
	wire w_dff_A_aj04g3bj4_1;
	wire w_dff_A_gY7FIhkc5_1;
	wire w_dff_A_wCli2Gti0_1;
	wire w_dff_A_5vjv4XYO9_1;
	wire w_dff_A_b9mZ2KQB0_1;
	wire w_dff_A_ivunJrwH4_1;
	wire w_dff_A_lGfZrXAS9_1;
	wire w_dff_A_7IGeBWFh0_1;
	wire w_dff_A_1coDZ5kC2_1;
	wire w_dff_A_sEhaFDJJ0_1;
	wire w_dff_A_y5jKn7ty6_1;
	wire w_dff_A_TPHP4biu1_1;
	wire w_dff_A_pxaZNlSl4_1;
	wire w_dff_A_RAC8Yl7x7_1;
	wire w_dff_A_0eyV9lEz2_1;
	wire w_dff_A_mNgCQiig8_2;
	wire w_dff_A_y1nXRSnK5_2;
	wire w_dff_A_B5Ac0O8K5_2;
	wire w_dff_A_swxcqNDD5_2;
	wire w_dff_A_T8Lxu1iO5_2;
	wire w_dff_A_73Tdf7ol7_2;
	wire w_dff_A_4SoxahjL2_2;
	wire w_dff_A_WFxcwB9S2_2;
	wire w_dff_A_9sVERyzN7_2;
	wire w_dff_A_3CfDnksh3_2;
	wire w_dff_A_5pjEuW558_2;
	wire w_dff_A_f6tYevuC1_2;
	wire w_dff_A_AhKoH0QZ0_2;
	wire w_dff_A_HjELsC5A1_2;
	wire w_dff_A_8q8Q82ie9_2;
	wire w_dff_A_3QogiG4a1_2;
	wire w_dff_A_7fIuVTFi8_2;
	wire w_dff_A_udxvaf216_2;
	wire w_dff_A_vY1EVIxP6_2;
	wire w_dff_A_wWyWsqDQ0_2;
	wire w_dff_A_RjO5YV3n9_2;
	wire w_dff_A_Vdt1oG7S1_2;
	wire w_dff_A_8zMVLYsD9_2;
	wire w_dff_A_ibcF77I59_2;
	wire w_dff_A_7ubQB2Fm9_2;
	wire w_dff_A_AcWnmXhW1_2;
	wire w_dff_A_p7j1aMtU4_2;
	wire w_dff_A_UNRhocXR4_2;
	wire w_dff_A_Gdxe3ZOr8_2;
	wire w_dff_A_fzySm9kS8_2;
	wire w_dff_A_31Yp8lUP4_2;
	wire w_dff_A_YLtUBQWC8_2;
	wire w_dff_A_ctpukIw40_2;
	wire w_dff_A_MG8GSihc2_2;
	wire w_dff_A_WvCZHVW40_2;
	wire w_dff_A_bg1MJ6p33_2;
	wire w_dff_A_A8d9CICa0_2;
	wire w_dff_A_6lPvK0jv6_2;
	wire w_dff_A_uotJZMkN8_2;
	wire w_dff_A_z8MM6RZQ8_2;
	wire w_dff_A_aRGfLVlE1_2;
	wire w_dff_A_OxUIVHDa5_2;
	wire w_dff_A_D1xwlsPT1_2;
	wire w_dff_A_YXCB7zUl6_0;
	wire w_dff_A_70lp1gHR9_0;
	wire w_dff_A_M3Z5D07K8_0;
	wire w_dff_A_tEixc4cS7_0;
	wire w_dff_A_4kdarGqW1_0;
	wire w_dff_A_r4dvnVmN5_0;
	wire w_dff_A_iJdPwCoZ2_0;
	wire w_dff_A_hWB0jgn51_0;
	wire w_dff_A_AbMz5S2W1_0;
	wire w_dff_A_pVHLXphT4_0;
	wire w_dff_A_zgCEQf6q4_0;
	wire w_dff_A_xYlQIh4F1_0;
	wire w_dff_A_jUJfMBc59_0;
	wire w_dff_A_j28GR6Ov8_0;
	wire w_dff_A_61HnOdxT1_0;
	wire w_dff_A_zkxOXXab0_0;
	wire w_dff_A_JcGOeZhc4_0;
	wire w_dff_A_wJDD0g888_0;
	wire w_dff_A_kpW8vJ3c7_0;
	wire w_dff_A_J0azdLdr1_0;
	wire w_dff_A_bXsos5Wl2_0;
	wire w_dff_A_enFVIsB98_0;
	wire w_dff_A_OWD1bF6y3_0;
	wire w_dff_A_m8hIAkfz1_0;
	wire w_dff_A_uCWGAXRX0_0;
	wire w_dff_A_iBSl5plc3_0;
	wire w_dff_A_zuskG7SG9_0;
	wire w_dff_A_HhPqdd4l1_0;
	wire w_dff_A_jIrz6R3B2_0;
	wire w_dff_A_q483wXra7_0;
	wire w_dff_A_6nVV6T3c0_0;
	wire w_dff_A_Sd21q1ia2_0;
	wire w_dff_A_NBkdc1KW1_0;
	wire w_dff_A_YBOdL1Ul3_0;
	wire w_dff_A_JKNGIHdO0_0;
	wire w_dff_A_D7N8Y8dP1_0;
	wire w_dff_A_9WzGAwzG9_0;
	wire w_dff_A_NeaAda4q1_0;
	wire w_dff_A_OPaaCXiF3_0;
	wire w_dff_A_Jdw2fPxG9_0;
	wire w_dff_A_MNJYD7c20_0;
	wire w_dff_A_Qwv3AjZl5_0;
	wire w_dff_A_X6vwduPr4_0;
	wire w_dff_A_cV0ii5IC2_0;
	wire w_dff_A_lIGy9qnK1_2;
	wire w_dff_A_Yms946IM2_0;
	wire w_dff_A_3O9aB6np8_0;
	wire w_dff_A_PAMpttRC2_0;
	wire w_dff_A_zrqntBIf8_0;
	wire w_dff_A_145wPxLy7_0;
	wire w_dff_A_9KthTZRE2_0;
	wire w_dff_A_Hs8fM28S0_0;
	wire w_dff_A_19YwcVEl1_0;
	wire w_dff_A_kJTNWExQ8_0;
	wire w_dff_A_lsY5VVDK4_0;
	wire w_dff_A_VFXng7rv1_0;
	wire w_dff_A_QKhzTLtn4_0;
	wire w_dff_A_6yBjoo4p9_0;
	wire w_dff_A_Naqlk2Mc8_0;
	wire w_dff_A_qk9xSDyE9_0;
	wire w_dff_A_IbWlIuzf6_0;
	wire w_dff_A_IUL2BnbZ9_0;
	wire w_dff_A_CwQY95RY8_0;
	wire w_dff_A_jmmDeEed0_0;
	wire w_dff_A_8TPblaNh9_0;
	wire w_dff_A_f7gjjkT66_0;
	wire w_dff_A_fokDOBqX0_0;
	wire w_dff_A_EOkUnT3Y9_0;
	wire w_dff_A_TU7oweEo5_0;
	wire w_dff_A_aEPT9noN2_0;
	wire w_dff_A_aXfgFULw2_0;
	wire w_dff_A_hgtTWBIc1_0;
	wire w_dff_A_YNVxmON74_0;
	wire w_dff_A_YGRqTFNp7_0;
	wire w_dff_A_QprqWveD2_0;
	wire w_dff_A_v4vjErgD4_0;
	wire w_dff_A_tOf1XTz83_0;
	wire w_dff_A_Juh47g114_0;
	wire w_dff_A_0VznXvK52_0;
	wire w_dff_A_sVyrxLrU4_0;
	wire w_dff_A_BJ9tlNVC8_0;
	wire w_dff_A_bY5QyAMS3_0;
	wire w_dff_A_2EigPglX2_0;
	wire w_dff_A_oo1LMv3F4_0;
	wire w_dff_A_baA821cv6_0;
	wire w_dff_A_QWIijunn1_2;
	wire w_dff_A_qNegFRs30_0;
	wire w_dff_A_avbzxA8K5_0;
	wire w_dff_A_XFhLLati8_0;
	wire w_dff_A_2M6rdHWa8_0;
	wire w_dff_A_gaQyrKER4_0;
	wire w_dff_A_evMP8BRa7_0;
	wire w_dff_A_Odanodd16_0;
	wire w_dff_A_FHhu5GBy0_0;
	wire w_dff_A_knwUz8vb8_0;
	wire w_dff_A_PPjjr6Ek2_0;
	wire w_dff_A_9yiZoM3N6_0;
	wire w_dff_A_cLiY4Yhy8_0;
	wire w_dff_A_aMxejYF88_0;
	wire w_dff_A_Co6zi4pN5_0;
	wire w_dff_A_JQmPX4R77_0;
	wire w_dff_A_dzK2YkCF7_0;
	wire w_dff_A_GyJafjJW1_0;
	wire w_dff_A_yr4ym27S8_0;
	wire w_dff_A_baeF2ZlL2_0;
	wire w_dff_A_kDNFZZ2I5_0;
	wire w_dff_A_Ld6cAEeq4_0;
	wire w_dff_A_tMFe6DGo4_0;
	wire w_dff_A_Jp9QMmEh5_0;
	wire w_dff_A_ummB57JS2_0;
	wire w_dff_A_kwixWjqq2_0;
	wire w_dff_A_Lga8gxrU1_0;
	wire w_dff_A_HmNCNAau6_0;
	wire w_dff_A_DoGQ16Dh2_0;
	wire w_dff_A_I7ubIESY7_0;
	wire w_dff_A_NQW85L9I3_0;
	wire w_dff_A_V0xTlsNd1_0;
	wire w_dff_A_Z1bnETvS7_0;
	wire w_dff_A_7ZGjbFEt9_0;
	wire w_dff_A_TK6DAxyF5_0;
	wire w_dff_A_b7vkck2R3_0;
	wire w_dff_A_QfGEX16i3_0;
	wire w_dff_A_RLCHDuhN6_0;
	wire w_dff_A_5YaOfvIe5_0;
	wire w_dff_A_WcfqmgfR5_0;
	wire w_dff_A_oRAz1Nyn2_2;
	wire w_dff_A_ZIdj2CVd0_0;
	wire w_dff_A_YrCGUe8g1_0;
	wire w_dff_A_qezTTKHw5_0;
	wire w_dff_A_HMjCTgyV9_0;
	wire w_dff_A_9LHthM2C0_0;
	wire w_dff_A_pyry5Pkw5_0;
	wire w_dff_A_yDgyKOuz4_0;
	wire w_dff_A_eXPvLlUl4_0;
	wire w_dff_A_KvjIEHiq3_0;
	wire w_dff_A_BPaUnHmN9_0;
	wire w_dff_A_Cw7Z87zf2_0;
	wire w_dff_A_O8sqpJQt9_0;
	wire w_dff_A_uyKQpU0Y5_0;
	wire w_dff_A_phWk8JiG6_0;
	wire w_dff_A_rqHnH6dV9_0;
	wire w_dff_A_45NN33Gw6_0;
	wire w_dff_A_HfbiPsJi3_0;
	wire w_dff_A_UOM9hux63_0;
	wire w_dff_A_cmqib9Zr2_0;
	wire w_dff_A_xWbaMkqZ0_0;
	wire w_dff_A_a4sGhVbG8_0;
	wire w_dff_A_w9uwQoXl7_0;
	wire w_dff_A_D9xK50206_0;
	wire w_dff_A_507e3veY6_0;
	wire w_dff_A_sU5wOAP63_0;
	wire w_dff_A_M7uRXGEH2_0;
	wire w_dff_A_7JZim46d9_0;
	wire w_dff_A_YeLKkgj59_0;
	wire w_dff_A_czoAlkgL1_0;
	wire w_dff_A_SvsvTzZc5_0;
	wire w_dff_A_nQWmn73N5_0;
	wire w_dff_A_gtEukHTK3_0;
	wire w_dff_A_774uUGHS4_0;
	wire w_dff_A_rk9oiF4S5_0;
	wire w_dff_A_Wc8Xy8Bm5_0;
	wire w_dff_A_ljXuj8UG9_0;
	wire w_dff_A_th4yLU1a9_0;
	wire w_dff_A_fQgYMzmB5_2;
	wire w_dff_A_Vm4r6kSA9_0;
	wire w_dff_A_cKM4hrn19_0;
	wire w_dff_A_VQLF6I0m4_0;
	wire w_dff_A_lzWt3GkF0_0;
	wire w_dff_A_JB4e1KLY0_0;
	wire w_dff_A_38sI1FJt2_0;
	wire w_dff_A_MSoVkhbI7_0;
	wire w_dff_A_61DNhxX66_0;
	wire w_dff_A_Ww5t9rKI9_0;
	wire w_dff_A_iiJwCTWB2_0;
	wire w_dff_A_hhVg1E5R5_0;
	wire w_dff_A_I46BmDXm9_0;
	wire w_dff_A_UIdOnfCi7_0;
	wire w_dff_A_ZnWYDBmG7_0;
	wire w_dff_A_5QpdIZtF9_0;
	wire w_dff_A_gLvrGR2Y3_0;
	wire w_dff_A_2j5wV0QH8_0;
	wire w_dff_A_hoEDNDer6_0;
	wire w_dff_A_cPOyXQ3M7_0;
	wire w_dff_A_rjbXorsZ3_0;
	wire w_dff_A_igl3qT3p1_0;
	wire w_dff_A_be6Owouh8_0;
	wire w_dff_A_X4ZsCPTt0_0;
	wire w_dff_A_dcgbj7sH3_0;
	wire w_dff_A_znBA6ZiU0_0;
	wire w_dff_A_WvlBKI9K8_0;
	wire w_dff_A_lSRhZmJy2_0;
	wire w_dff_A_6Mim457e3_0;
	wire w_dff_A_SElGqOG34_0;
	wire w_dff_A_ARUYfesm0_0;
	wire w_dff_A_EODH7g842_0;
	wire w_dff_A_296RwDxi7_0;
	wire w_dff_A_eCqOjRHE4_0;
	wire w_dff_A_fUDJXR8i0_0;
	wire w_dff_A_4U5OUJGW4_0;
	wire w_dff_A_Zdk0dlCk2_2;
	wire w_dff_A_9yFvthSH3_0;
	wire w_dff_A_6JejdKBu5_0;
	wire w_dff_A_SszONaO97_0;
	wire w_dff_A_DC1s2nnq2_0;
	wire w_dff_A_CJmFnuZt5_0;
	wire w_dff_A_O5pdFJEe5_0;
	wire w_dff_A_ft8TwJPZ9_0;
	wire w_dff_A_HxNumhOn6_0;
	wire w_dff_A_jIooTm9d3_0;
	wire w_dff_A_i9vGzzLv4_0;
	wire w_dff_A_3lJLA2Yt9_0;
	wire w_dff_A_9VrcpKBu3_0;
	wire w_dff_A_XYftsUyd9_0;
	wire w_dff_A_ocGg1ky89_0;
	wire w_dff_A_vi0nIyCM3_0;
	wire w_dff_A_RnnA6yeb6_0;
	wire w_dff_A_6OnaoYbA1_0;
	wire w_dff_A_3b6lSHj47_0;
	wire w_dff_A_qzTRnjzg0_0;
	wire w_dff_A_3ViHq50n9_0;
	wire w_dff_A_eNBB4EP73_0;
	wire w_dff_A_5oXrXCIH3_0;
	wire w_dff_A_TOVy9fie3_0;
	wire w_dff_A_f6Dq06jn3_0;
	wire w_dff_A_4ZkwPbzT3_0;
	wire w_dff_A_S1q3s3Fz0_0;
	wire w_dff_A_eLE1IRuJ8_0;
	wire w_dff_A_bGLybw8o0_0;
	wire w_dff_A_DbqWJFSd7_0;
	wire w_dff_A_vfZVeqtS2_0;
	wire w_dff_A_gO82Gl7T1_0;
	wire w_dff_A_2Aa8zRq84_0;
	wire w_dff_A_Qta0xbLt4_0;
	wire w_dff_A_y6UHYdvt4_2;
	wire w_dff_A_VSczgI9a5_0;
	wire w_dff_A_Cd928ia36_0;
	wire w_dff_A_V4ucMXfr3_0;
	wire w_dff_A_PghwdNzX0_0;
	wire w_dff_A_CZT15yUT9_0;
	wire w_dff_A_XWStr6gT2_0;
	wire w_dff_A_njAZfeca5_0;
	wire w_dff_A_nGr7frN61_0;
	wire w_dff_A_BX1N2P5a4_0;
	wire w_dff_A_vLHec2pN9_0;
	wire w_dff_A_fiV0BgNN1_0;
	wire w_dff_A_yuT1EXrx2_0;
	wire w_dff_A_2xevLxyK6_0;
	wire w_dff_A_lFASKJbU0_0;
	wire w_dff_A_GKPY07cg4_0;
	wire w_dff_A_jAOyFJTn7_0;
	wire w_dff_A_d8IGNN0A8_0;
	wire w_dff_A_MYDDFt994_0;
	wire w_dff_A_TJnfdsga9_0;
	wire w_dff_A_UVY9Iozz4_0;
	wire w_dff_A_9FAIB4Ar5_0;
	wire w_dff_A_0p8MIe4W5_0;
	wire w_dff_A_Gx0IniJa7_0;
	wire w_dff_A_0CRCesfm7_0;
	wire w_dff_A_A3uCyWZb8_0;
	wire w_dff_A_tULTtL3L6_0;
	wire w_dff_A_TSzkUqFK7_0;
	wire w_dff_A_6XgM8n5L3_0;
	wire w_dff_A_Bka5OWbA6_0;
	wire w_dff_A_Ybo2tHbZ1_0;
	wire w_dff_A_Wg5zbNkE5_0;
	wire w_dff_A_RryB5Bx36_2;
	wire w_dff_A_2q2xAQeC6_0;
	wire w_dff_A_ZPXUbUTb3_0;
	wire w_dff_A_nxCr2dCa0_0;
	wire w_dff_A_WVoKf6jI4_0;
	wire w_dff_A_yeK30YaD2_0;
	wire w_dff_A_k6gT5kZQ2_0;
	wire w_dff_A_5oEVdd244_0;
	wire w_dff_A_smd1EMQt4_0;
	wire w_dff_A_NxAkp4N11_0;
	wire w_dff_A_7xEYWvSz5_0;
	wire w_dff_A_A5UiPDDN7_0;
	wire w_dff_A_gAbQAD9q5_0;
	wire w_dff_A_1OxsGPe50_0;
	wire w_dff_A_jh7oYIIn3_0;
	wire w_dff_A_axZCnYeL3_0;
	wire w_dff_A_jeRq0WL24_0;
	wire w_dff_A_hp2rcP6N9_0;
	wire w_dff_A_GhLQdO0E4_0;
	wire w_dff_A_BRkMEQ5r8_0;
	wire w_dff_A_JxBDSVW62_0;
	wire w_dff_A_4mf4bNWe1_0;
	wire w_dff_A_HTcJQbg33_0;
	wire w_dff_A_IZfYf7nS2_0;
	wire w_dff_A_LjAx4rqT4_0;
	wire w_dff_A_chrLxxQm0_0;
	wire w_dff_A_6DcrJCLa9_0;
	wire w_dff_A_09szml5I4_0;
	wire w_dff_A_vFVYQM431_0;
	wire w_dff_A_jfDZfkmv1_0;
	wire w_dff_A_bZHWsZ3E8_2;
	wire w_dff_A_SA1CQeSI7_0;
	wire w_dff_A_vFywo5td6_0;
	wire w_dff_A_7q9XyUWj2_0;
	wire w_dff_A_4hASwI6f9_0;
	wire w_dff_A_Ydyk6nff2_0;
	wire w_dff_A_azSuLj7Q9_0;
	wire w_dff_A_Sz0SlQX26_0;
	wire w_dff_A_YkPWNupc7_0;
	wire w_dff_A_I3sfRKQf6_0;
	wire w_dff_A_DksUjKGx6_0;
	wire w_dff_A_zgn3vwlh0_0;
	wire w_dff_A_wxl2hvhu1_0;
	wire w_dff_A_j0UnreYl0_0;
	wire w_dff_A_v7jindob5_0;
	wire w_dff_A_NCarShOt9_0;
	wire w_dff_A_TMW7sxXM8_0;
	wire w_dff_A_h6szTUnb4_0;
	wire w_dff_A_y4WB1Hpz1_0;
	wire w_dff_A_hblJQGDh8_0;
	wire w_dff_A_sIfycOJl3_0;
	wire w_dff_A_UoyzXXtz8_0;
	wire w_dff_A_B20mjgdN9_0;
	wire w_dff_A_7Mrz7gZ40_0;
	wire w_dff_A_1qMKwhEQ7_0;
	wire w_dff_A_I4JQ4Did4_0;
	wire w_dff_A_7NuQY5cf0_0;
	wire w_dff_A_wIweRCIZ6_0;
	wire w_dff_A_u8ZD7jxR4_2;
	wire w_dff_A_xIjmN53W8_0;
	wire w_dff_A_VvJfRlVy1_0;
	wire w_dff_A_rpnuCX2m3_0;
	wire w_dff_A_en97lUwR2_0;
	wire w_dff_A_lTJkpVQQ7_0;
	wire w_dff_A_TPzfFAbM5_0;
	wire w_dff_A_WY9GZPqX7_0;
	wire w_dff_A_J19n05Kp8_0;
	wire w_dff_A_uY42FFpW9_0;
	wire w_dff_A_EorRc6GK5_0;
	wire w_dff_A_UTAfM9Ld6_0;
	wire w_dff_A_WoguPPsq8_0;
	wire w_dff_A_wTXLXwnW0_0;
	wire w_dff_A_eIlvoaGs8_0;
	wire w_dff_A_W7ALtZPI5_0;
	wire w_dff_A_zHaN7Vux1_0;
	wire w_dff_A_TbGOdZon0_0;
	wire w_dff_A_4lwN3GCC4_0;
	wire w_dff_A_LDf80yb75_0;
	wire w_dff_A_w5dAdQPn1_0;
	wire w_dff_A_toEoJcX35_0;
	wire w_dff_A_TzyBSbEB7_0;
	wire w_dff_A_hkJdPfo42_0;
	wire w_dff_A_SzG6izqJ5_0;
	wire w_dff_A_Wh7Nsh6u6_0;
	wire w_dff_A_SP0xCeW41_2;
	wire w_dff_A_zCw8m8dq0_0;
	wire w_dff_A_wcuoHtPZ2_0;
	wire w_dff_A_cBxi1A4y6_0;
	wire w_dff_A_zNCMFdRD3_0;
	wire w_dff_A_6w1qM55O1_0;
	wire w_dff_A_j4gC81zA6_0;
	wire w_dff_A_jAlXBA9k3_0;
	wire w_dff_A_mboHtXUS9_0;
	wire w_dff_A_kx82cDBm4_0;
	wire w_dff_A_5NLq3L9W2_0;
	wire w_dff_A_N3M452Qp5_0;
	wire w_dff_A_20zhR8K87_0;
	wire w_dff_A_nIeJ6drv6_0;
	wire w_dff_A_fFimfUza6_0;
	wire w_dff_A_Agh7AKyL0_0;
	wire w_dff_A_oH248Y4P4_0;
	wire w_dff_A_81AFO8ut4_0;
	wire w_dff_A_xE382PUD8_0;
	wire w_dff_A_WiLblRlj2_0;
	wire w_dff_A_mXqmIs4H4_0;
	wire w_dff_A_Dg6kfu2O1_0;
	wire w_dff_A_rziDBC9L5_0;
	wire w_dff_A_S10WfadL7_0;
	wire w_dff_A_gP8OwZoN2_2;
	wire w_dff_A_vYEU9rof4_0;
	wire w_dff_A_cmBoHTo26_0;
	wire w_dff_A_xZ2zrSHd7_0;
	wire w_dff_A_6YawxdGv6_0;
	wire w_dff_A_xWOYFBbj2_0;
	wire w_dff_A_ezdOWVDX2_0;
	wire w_dff_A_Oy0RtZ3C6_0;
	wire w_dff_A_EkJtWrnA6_0;
	wire w_dff_A_R873z4GN2_0;
	wire w_dff_A_dKfo5FFq8_0;
	wire w_dff_A_euFG9zf55_0;
	wire w_dff_A_x39Ff9zt8_0;
	wire w_dff_A_meAbKCtT8_0;
	wire w_dff_A_iZJ3QSDR9_0;
	wire w_dff_A_GYdczOMX1_0;
	wire w_dff_A_zaOeb0f63_0;
	wire w_dff_A_pwtacHqE4_0;
	wire w_dff_A_XuWS0maq8_0;
	wire w_dff_A_PYTOf91n7_0;
	wire w_dff_A_m7Rav7Rh8_0;
	wire w_dff_A_xyIOOBwo1_0;
	wire w_dff_A_5LHruE6g9_2;
	wire w_dff_A_XraBX9ax8_0;
	wire w_dff_A_36XP6H9o3_0;
	wire w_dff_A_oMdRGqlV4_0;
	wire w_dff_A_jRegBd9L2_0;
	wire w_dff_A_gQxxtX7L3_0;
	wire w_dff_A_2G8L8kIx3_0;
	wire w_dff_A_0LDLR0aL2_0;
	wire w_dff_A_V8hz3nfq6_0;
	wire w_dff_A_KKZotsfK4_0;
	wire w_dff_A_QETzy8Qf0_0;
	wire w_dff_A_tC1zSLKx6_0;
	wire w_dff_A_kPOlxqHF4_0;
	wire w_dff_A_FiwSAyo31_0;
	wire w_dff_A_eOmUKcvu1_0;
	wire w_dff_A_FgYbu4IE2_0;
	wire w_dff_A_CX4aF0us2_0;
	wire w_dff_A_Hfxu5oWq8_0;
	wire w_dff_A_btSXAvG23_0;
	wire w_dff_A_QWZuBYSD7_0;
	wire w_dff_A_oxEVAVgt4_2;
	wire w_dff_A_FPVKDFJ45_0;
	wire w_dff_A_ToSWAq2x5_0;
	wire w_dff_A_wM0OhjKk0_0;
	wire w_dff_A_V9Yf3nlK6_0;
	wire w_dff_A_bHPpDfnj2_0;
	wire w_dff_A_J67J2Nt24_0;
	wire w_dff_A_Y5IUSRh22_0;
	wire w_dff_A_WUHuYyqG9_0;
	wire w_dff_A_9w0Xae3d8_0;
	wire w_dff_A_PoAdZYf43_0;
	wire w_dff_A_NfoXnuL88_0;
	wire w_dff_A_o6vZFeEC2_0;
	wire w_dff_A_wAH8io2v1_0;
	wire w_dff_A_ywLq8MK66_0;
	wire w_dff_A_u4gMFVF98_0;
	wire w_dff_A_Ge9anYdW7_0;
	wire w_dff_A_OOy7QXUP8_0;
	wire w_dff_A_CHdzBFmi0_2;
	wire w_dff_A_UnU6ipts8_0;
	wire w_dff_A_URYwyff68_0;
	wire w_dff_A_DJO6BGWh1_0;
	wire w_dff_A_XK0V8Yav0_0;
	wire w_dff_A_lrIuidol1_0;
	wire w_dff_A_8k3b3W493_0;
	wire w_dff_A_scJTSTg71_0;
	wire w_dff_A_X5d0iTYj7_0;
	wire w_dff_A_yaIwIwEV5_0;
	wire w_dff_A_mp6WrrJI0_0;
	wire w_dff_A_wFhcnsMx3_0;
	wire w_dff_A_xzfUSp979_0;
	wire w_dff_A_sdbpSfTh9_0;
	wire w_dff_A_8pzOy3UG5_0;
	wire w_dff_A_hEgTE9hf0_0;
	wire w_dff_A_rLUmXsuL3_2;
	wire w_dff_A_otiGIucp1_0;
	wire w_dff_A_QCIAlclO5_0;
	wire w_dff_A_PKNUWaTc8_0;
	wire w_dff_A_tnvxfwEx6_0;
	wire w_dff_A_bI7eZstP8_0;
	wire w_dff_A_LfD11Ul04_0;
	wire w_dff_A_uCEdhaHI9_0;
	wire w_dff_A_VSNBlYSA8_0;
	wire w_dff_A_DunAigsW4_0;
	wire w_dff_A_ws1ZNx7D7_0;
	wire w_dff_A_eQ2uXRjN7_0;
	wire w_dff_A_qkbQYpJS9_0;
	wire w_dff_A_6w7bUJw38_0;
	wire w_dff_A_J2WpamXl7_2;
	wire w_dff_A_SSc9x9V91_0;
	wire w_dff_A_RoJR0kUy8_0;
	wire w_dff_A_VFhQUbqC4_0;
	wire w_dff_A_gKxJifTD3_0;
	wire w_dff_A_zK6tjDpz5_0;
	wire w_dff_A_2EczkCpu2_0;
	wire w_dff_A_7dlymOGj7_0;
	wire w_dff_A_KcxQcDa58_0;
	wire w_dff_A_6qiLiz9K4_0;
	wire w_dff_A_QV6JNCbe6_0;
	wire w_dff_A_k0YYIuNo5_2;
	wire w_dff_A_7bgQ0bRC0_0;
	wire w_dff_A_wxlMlu5M2_0;
	wire w_dff_A_SCmN7kIq5_0;
	wire w_dff_A_GBCejgwR2_0;
	wire w_dff_A_rLusq6RD4_0;
	wire w_dff_A_wOGxBmPA5_0;
	wire w_dff_A_rqlcZPUQ3_0;
	wire w_dff_A_wzXcXi204_0;
	wire w_dff_A_0nVz4h2P4_2;
	wire w_dff_A_7ztwvdHZ5_0;
	wire w_dff_A_HxzPE9Ro9_0;
	wire w_dff_A_6itk3QDR1_0;
	wire w_dff_A_J1zHO9iV7_0;
	wire w_dff_A_PHDW0HQK8_0;
	wire w_dff_A_cGXW2PwO3_0;
	wire w_dff_A_Cw7elsfJ2_2;
	wire w_dff_A_SQqGAZ728_0;
	wire w_dff_A_ieToSDME3_0;
	wire w_dff_A_r1o6n5ps1_0;
	wire w_dff_A_GC1Xlu628_0;
	wire w_dff_A_gS2lI5Ue9_2;
	wire w_dff_A_G2ckHM4a8_0;
	wire w_dff_A_xrK6u3Nq1_0;
	wire w_dff_A_UG9OPTVc9_0;
	wire w_dff_A_TNSINLGv9_2;
	wire w_dff_A_mEOc6pxz8_0;
	wire w_dff_A_S7Y49kXp0_0;
	wire w_dff_A_HR8wY1806_2;
	wire w_dff_A_b1AKM4qo9_0;
	jnot g0000(.din(w_a22_6[1]),.dout(n49),.clk(gclk));
	jor g0001(.dina(w_a2_1[2]),.dinb(w_a1_0[2]),.dout(n50),.clk(gclk));
	jor g0002(.dina(n50),.dinb(w_a0_1[1]),.dout(n51),.clk(gclk));
	jor g0003(.dina(w_n51_0[1]),.dinb(w_a3_0[2]),.dout(n52),.clk(gclk));
	jor g0004(.dina(w_n52_0[1]),.dinb(w_a4_1[1]),.dout(n53),.clk(gclk));
	jand g0005(.dina(w_n53_0[1]),.dinb(w_n49_5[1]),.dout(n54),.clk(gclk));
	jxor g0006(.dina(w_n54_0[1]),.dinb(w_a5_0[2]),.dout(n55),.clk(gclk));
	jnot g0007(.din(w_n55_9[2]),.dout(n56),.clk(gclk));
	jand g0008(.dina(w_n51_0[0]),.dinb(w_n49_5[0]),.dout(n57),.clk(gclk));
	jxor g0009(.dina(w_n57_0[1]),.dinb(w_a3_0[1]),.dout(n58),.clk(gclk));
	jnot g0010(.din(w_n58_4[2]),.dout(n59),.clk(gclk));
	jand g0011(.dina(w_a22_6[0]),.dinb(w_a2_1[1]),.dout(n60),.clk(gclk));
	jnot g0012(.din(w_a0_1[0]),.dout(n61),.clk(gclk));
	jnot g0013(.din(w_a1_0[1]),.dout(n62),.clk(gclk));
	jand g0014(.dina(w_n62_0[2]),.dinb(w_n61_1[2]),.dout(n63),.clk(gclk));
	jnot g0015(.din(w_n63_2[2]),.dout(n64),.clk(gclk));
	jand g0016(.dina(w_n64_0[1]),.dinb(w_a2_1[0]),.dout(n65),.clk(gclk));
	jnot g0017(.din(n65),.dout(n66),.clk(gclk));
	jand g0018(.dina(n66),.dinb(w_n57_0[0]),.dout(n67),.clk(gclk));
	jor g0019(.dina(n67),.dinb(n60),.dout(n68),.clk(gclk));
	jxor g0020(.dina(w_n68_6[2]),.dinb(w_n59_3[1]),.dout(n69),.clk(gclk));
	jnot g0021(.din(w_n69_0[2]),.dout(n70),.clk(gclk));
	jand g0022(.dina(w_a22_5[2]),.dinb(w_a4_1[0]),.dout(n71),.clk(gclk));
	jand g0023(.dina(w_n52_0[0]),.dinb(w_a4_0[2]),.dout(n72),.clk(gclk));
	jnot g0024(.din(n72),.dout(n73),.clk(gclk));
	jand g0025(.dina(n73),.dinb(w_n54_0[0]),.dout(n74),.clk(gclk));
	jor g0026(.dina(n74),.dinb(n71),.dout(n75),.clk(gclk));
	jxor g0027(.dina(w_n75_5[2]),.dinb(w_n56_12[2]),.dout(n76),.clk(gclk));
	jnot g0028(.din(w_n76_0[1]),.dout(n77),.clk(gclk));
	jand g0029(.dina(w_n77_0[1]),.dinb(w_n70_0[2]),.dout(n78),.clk(gclk));
	jnot g0030(.din(w_n78_2[2]),.dout(n79),.clk(gclk));
	jand g0031(.dina(w_a22_5[1]),.dinb(w_a15_1[1]),.dout(n80),.clk(gclk));
	jor g0032(.dina(w_n53_0[0]),.dinb(w_a5_0[1]),.dout(n81),.clk(gclk));
	jor g0033(.dina(w_n81_0[1]),.dinb(w_a6_1[1]),.dout(n82),.clk(gclk));
	jor g0034(.dina(w_n82_0[1]),.dinb(w_a7_0[2]),.dout(n83),.clk(gclk));
	jor g0035(.dina(w_n83_0[1]),.dinb(w_a8_1[1]),.dout(n84),.clk(gclk));
	jor g0036(.dina(w_n84_0[1]),.dinb(w_a9_0[2]),.dout(n85),.clk(gclk));
	jor g0037(.dina(w_n85_0[1]),.dinb(w_a10_1[1]),.dout(n86),.clk(gclk));
	jor g0038(.dina(w_n86_0[1]),.dinb(w_a11_0[2]),.dout(n87),.clk(gclk));
	jor g0039(.dina(w_n87_0[1]),.dinb(w_a12_1[1]),.dout(n88),.clk(gclk));
	jor g0040(.dina(w_n88_0[1]),.dinb(w_a13_0[2]),.dout(n89),.clk(gclk));
	jor g0041(.dina(w_n89_0[1]),.dinb(w_a14_1[1]),.dout(n90),.clk(gclk));
	jor g0042(.dina(w_n90_0[1]),.dinb(w_a15_1[0]),.dout(n91),.clk(gclk));
	jand g0043(.dina(w_n91_0[1]),.dinb(w_n49_4[2]),.dout(n92),.clk(gclk));
	jand g0044(.dina(w_n90_0[0]),.dinb(w_a15_0[2]),.dout(n93),.clk(gclk));
	jnot g0045(.din(n93),.dout(n94),.clk(gclk));
	jand g0046(.dina(n94),.dinb(w_n92_0[1]),.dout(n95),.clk(gclk));
	jor g0047(.dina(n95),.dinb(n80),.dout(n96),.clk(gclk));
	jor g0048(.dina(w_n91_0[0]),.dinb(w_a16_0[2]),.dout(n97),.clk(gclk));
	jor g0049(.dina(w_n97_0[1]),.dinb(w_a17_0[1]),.dout(n98),.clk(gclk));
	jor g0050(.dina(w_n98_0[1]),.dinb(w_a18_1[1]),.dout(n99),.clk(gclk));
	jor g0051(.dina(w_n99_0[1]),.dinb(w_a19_0[2]),.dout(n100),.clk(gclk));
	jor g0052(.dina(w_n100_0[1]),.dinb(w_a20_1[1]),.dout(n101),.clk(gclk));
	jand g0053(.dina(n101),.dinb(w_n49_4[1]),.dout(n102),.clk(gclk));
	jxor g0054(.dina(w_n102_0[1]),.dinb(w_a21_0[1]),.dout(n103),.clk(gclk));
	jand g0055(.dina(w_a22_5[0]),.dinb(w_a20_1[0]),.dout(n104),.clk(gclk));
	jand g0056(.dina(w_n100_0[0]),.dinb(w_a20_0[2]),.dout(n105),.clk(gclk));
	jnot g0057(.din(w_n105_0[1]),.dout(n106),.clk(gclk));
	jand g0058(.dina(n106),.dinb(w_n102_0[0]),.dout(n107),.clk(gclk));
	jor g0059(.dina(n107),.dinb(w_n104_0[1]),.dout(n108),.clk(gclk));
	jand g0060(.dina(w_n108_1[1]),.dinb(w_n103_1[1]),.dout(n109),.clk(gclk));
	jand g0061(.dina(w_n109_2[1]),.dinb(w_n96_5[2]),.dout(n110),.clk(gclk));
	jand g0062(.dina(w_a22_4[2]),.dinb(w_a18_1[0]),.dout(n111),.clk(gclk));
	jand g0063(.dina(w_n99_0[0]),.dinb(w_n49_4[0]),.dout(n112),.clk(gclk));
	jand g0064(.dina(w_n98_0[0]),.dinb(w_a18_0[2]),.dout(n113),.clk(gclk));
	jnot g0065(.din(n113),.dout(n114),.clk(gclk));
	jand g0066(.dina(n114),.dinb(w_n112_0[1]),.dout(n115),.clk(gclk));
	jor g0067(.dina(n115),.dinb(n111),.dout(n116),.clk(gclk));
	jxor g0068(.dina(w_n112_0[0]),.dinb(w_a19_0[1]),.dout(n117),.clk(gclk));
	jnot g0069(.din(w_n117_0[1]),.dout(n118),.clk(gclk));
	jor g0070(.dina(w_n118_0[2]),.dinb(w_n116_1[1]),.dout(n119),.clk(gclk));
	jnot g0071(.din(w_n119_0[1]),.dout(n120),.clk(gclk));
	jnot g0072(.din(w_a17_0[0]),.dout(n121),.clk(gclk));
	jand g0073(.dina(w_n97_0[0]),.dinb(w_n49_3[2]),.dout(n122),.clk(gclk));
	jxor g0074(.dina(n122),.dinb(w_n121_0[1]),.dout(n123),.clk(gclk));
	jnot g0075(.din(w_n123_1[1]),.dout(n124),.clk(gclk));
	jxor g0076(.dina(w_n92_0[0]),.dinb(w_a16_0[1]),.dout(n125),.clk(gclk));
	jnot g0077(.din(w_n125_0[1]),.dout(n126),.clk(gclk));
	jand g0078(.dina(w_n126_0[2]),.dinb(n124),.dout(n127),.clk(gclk));
	jand g0079(.dina(w_n127_1[1]),.dinb(w_n120_0[2]),.dout(n128),.clk(gclk));
	jand g0080(.dina(w_n128_2[2]),.dinb(w_n110_6[1]),.dout(n129),.clk(gclk));
	jnot g0081(.din(n129),.dout(n130),.clk(gclk));
	jor g0082(.dina(w_n126_0[1]),.dinb(w_n123_1[0]),.dout(n131),.clk(gclk));
	jnot g0083(.din(w_n131_0[1]),.dout(n132),.clk(gclk));
	jnot g0084(.din(w_n116_1[0]),.dout(n133),.clk(gclk));
	jand g0085(.dina(w_n118_0[1]),.dinb(n133),.dout(n134),.clk(gclk));
	jand g0086(.dina(w_n134_1[1]),.dinb(w_n132_0[2]),.dout(n135),.clk(gclk));
	jand g0087(.dina(w_n135_2[2]),.dinb(w_n109_2[0]),.dout(n136),.clk(gclk));
	jand g0088(.dina(w_n136_0[2]),.dinb(w_n96_5[1]),.dout(n137),.clk(gclk));
	jnot g0089(.din(w_n137_0[1]),.dout(n138),.clk(gclk));
	jand g0090(.dina(w_n117_0[0]),.dinb(w_n116_0[2]),.dout(n139),.clk(gclk));
	jand g0091(.dina(w_n125_0[0]),.dinb(w_n123_0[2]),.dout(n140),.clk(gclk));
	jand g0092(.dina(w_n140_1[1]),.dinb(w_n139_1[1]),.dout(n141),.clk(gclk));
	jnot g0093(.din(w_n141_2[1]),.dout(n142),.clk(gclk));
	jnot g0094(.din(w_n96_5[0]),.dout(n143),.clk(gclk));
	jnot g0095(.din(w_n103_1[0]),.dout(n144),.clk(gclk));
	jor g0096(.dina(w_n108_1[0]),.dinb(w_n144_0[2]),.dout(n145),.clk(gclk));
	jor g0097(.dina(w_n145_1[1]),.dinb(w_n143_6[1]),.dout(n146),.clk(gclk));
	jor g0098(.dina(w_n146_4[2]),.dinb(w_n142_1[1]),.dout(n147),.clk(gclk));
	jand g0099(.dina(w_n147_4[1]),.dinb(w_n138_4[1]),.dout(n148),.clk(gclk));
	jand g0100(.dina(n148),.dinb(w_n130_2[2]),.dout(n149),.clk(gclk));
	jnot g0101(.din(n149),.dout(n150),.clk(gclk));
	jand g0102(.dina(w_n109_1[2]),.dinb(w_n143_6[0]),.dout(n151),.clk(gclk));
	jand g0103(.dina(w_n151_6[1]),.dinb(w_n128_2[1]),.dout(n152),.clk(gclk));
	jnot g0104(.din(w_n152_0[1]),.dout(n153),.clk(gclk));
	jor g0105(.dina(w_n131_0[0]),.dinb(w_n119_0[0]),.dout(n154),.clk(gclk));
	jnot g0106(.din(w_n154_1[1]),.dout(n155),.clk(gclk));
	jand g0107(.dina(w_n155_1[1]),.dinb(w_n151_6[0]),.dout(n156),.clk(gclk));
	jnot g0108(.din(w_n156_0[1]),.dout(n157),.clk(gclk));
	jand g0109(.dina(w_n157_1[2]),.dinb(w_n153_1[1]),.dout(n158),.clk(gclk));
	jnot g0110(.din(w_n158_1[1]),.dout(n159),.clk(gclk));
	jand g0111(.dina(w_n136_0[1]),.dinb(w_n143_5[2]),.dout(n160),.clk(gclk));
	jnot g0112(.din(w_n146_4[1]),.dout(n161),.clk(gclk));
	jand g0113(.dina(w_n126_0[0]),.dinb(w_n123_0[1]),.dout(n162),.clk(gclk));
	jand g0114(.dina(w_n162_1[1]),.dinb(w_n139_1[0]),.dout(n163),.clk(gclk));
	jand g0115(.dina(w_n163_2[2]),.dinb(w_n161_0[2]),.dout(n164),.clk(gclk));
	jor g0116(.dina(w_n164_0[2]),.dinb(w_n160_0[2]),.dout(n165),.clk(gclk));
	jor g0117(.dina(w_n165_0[1]),.dinb(n159),.dout(n166),.clk(gclk));
	jor g0118(.dina(n166),.dinb(n150),.dout(n167),.clk(gclk));
	jnot g0119(.din(w_n167_0[1]),.dout(n168),.clk(gclk));
	jnot g0120(.din(w_n104_0[0]),.dout(n169),.clk(gclk));
	jnot g0121(.din(w_a20_0[1]),.dout(n170),.clk(gclk));
	jnot g0122(.din(w_a19_0[0]),.dout(n171),.clk(gclk));
	jnot g0123(.din(w_a18_0[1]),.dout(n172),.clk(gclk));
	jnot g0124(.din(w_a16_0[0]),.dout(n173),.clk(gclk));
	jnot g0125(.din(w_a15_0[1]),.dout(n174),.clk(gclk));
	jnot g0126(.din(w_a14_1[0]),.dout(n175),.clk(gclk));
	jnot g0127(.din(w_a13_0[1]),.dout(n176),.clk(gclk));
	jnot g0128(.din(w_a12_1[0]),.dout(n177),.clk(gclk));
	jnot g0129(.din(w_a11_0[1]),.dout(n178),.clk(gclk));
	jnot g0130(.din(w_a10_1[0]),.dout(n179),.clk(gclk));
	jnot g0131(.din(w_a9_0[1]),.dout(n180),.clk(gclk));
	jnot g0132(.din(w_a8_1[0]),.dout(n181),.clk(gclk));
	jnot g0133(.din(w_a7_0[1]),.dout(n182),.clk(gclk));
	jnot g0134(.din(w_a6_1[0]),.dout(n183),.clk(gclk));
	jnot g0135(.din(w_a5_0[0]),.dout(n184),.clk(gclk));
	jnot g0136(.din(w_a4_0[1]),.dout(n185),.clk(gclk));
	jnot g0137(.din(w_a3_0[0]),.dout(n186),.clk(gclk));
	jnot g0138(.din(w_a2_0[2]),.dout(n187),.clk(gclk));
	jand g0139(.dina(n187),.dinb(w_n62_0[1]),.dout(n188),.clk(gclk));
	jand g0140(.dina(n188),.dinb(w_n61_1[1]),.dout(n189),.clk(gclk));
	jand g0141(.dina(n189),.dinb(n186),.dout(n190),.clk(gclk));
	jand g0142(.dina(n190),.dinb(n185),.dout(n191),.clk(gclk));
	jand g0143(.dina(n191),.dinb(n184),.dout(n192),.clk(gclk));
	jand g0144(.dina(n192),.dinb(n183),.dout(n193),.clk(gclk));
	jand g0145(.dina(n193),.dinb(n182),.dout(n194),.clk(gclk));
	jand g0146(.dina(n194),.dinb(n181),.dout(n195),.clk(gclk));
	jand g0147(.dina(n195),.dinb(n180),.dout(n196),.clk(gclk));
	jand g0148(.dina(n196),.dinb(n179),.dout(n197),.clk(gclk));
	jand g0149(.dina(n197),.dinb(n178),.dout(n198),.clk(gclk));
	jand g0150(.dina(n198),.dinb(n177),.dout(n199),.clk(gclk));
	jand g0151(.dina(n199),.dinb(n176),.dout(n200),.clk(gclk));
	jand g0152(.dina(n200),.dinb(n175),.dout(n201),.clk(gclk));
	jand g0153(.dina(w_n201_0[1]),.dinb(n174),.dout(n202),.clk(gclk));
	jand g0154(.dina(n202),.dinb(n173),.dout(n203),.clk(gclk));
	jand g0155(.dina(n203),.dinb(w_n121_0[0]),.dout(n204),.clk(gclk));
	jand g0156(.dina(n204),.dinb(n172),.dout(n205),.clk(gclk));
	jand g0157(.dina(n205),.dinb(n171),.dout(n206),.clk(gclk));
	jand g0158(.dina(n206),.dinb(n170),.dout(n207),.clk(gclk));
	jor g0159(.dina(w_n207_0[1]),.dinb(w_a22_4[1]),.dout(n208),.clk(gclk));
	jor g0160(.dina(w_n105_0[0]),.dinb(n208),.dout(n209),.clk(gclk));
	jand g0161(.dina(n209),.dinb(n169),.dout(n210),.clk(gclk));
	jand g0162(.dina(w_n210_0[1]),.dinb(w_n103_0[2]),.dout(n211),.clk(gclk));
	jand g0163(.dina(w_n211_1[1]),.dinb(w_n143_5[1]),.dout(n212),.clk(gclk));
	jand g0164(.dina(w_n212_3[1]),.dinb(w_n163_2[1]),.dout(n213),.clk(gclk));
	jnot g0165(.din(w_n213_1[1]),.dout(n214),.clk(gclk));
	jor g0166(.dina(w_n145_1[0]),.dinb(w_n96_4[2]),.dout(n215),.clk(gclk));
	jor g0167(.dina(w_n215_2[1]),.dinb(w_n142_1[0]),.dout(n216),.clk(gclk));
	jand g0168(.dina(w_n216_4[1]),.dinb(w_n214_2[2]),.dout(n217),.clk(gclk));
	jand g0169(.dina(n217),.dinb(n168),.dout(n218),.clk(gclk));
	jand g0170(.dina(w_n118_0[0]),.dinb(w_n116_0[1]),.dout(n219),.clk(gclk));
	jand g0171(.dina(w_n219_1[1]),.dinb(w_n132_0[1]),.dout(n220),.clk(gclk));
	jand g0172(.dina(w_n220_3[1]),.dinb(w_n151_5[2]),.dout(n221),.clk(gclk));
	jnot g0173(.din(n221),.dout(n222),.clk(gclk));
	jand g0174(.dina(w_n140_1[0]),.dinb(w_n120_0[1]),.dout(n223),.clk(gclk));
	jand g0175(.dina(w_n223_2[2]),.dinb(w_n212_3[0]),.dout(n224),.clk(gclk));
	jnot g0176(.din(w_n224_0[2]),.dout(n225),.clk(gclk));
	jand g0177(.dina(w_n225_2[2]),.dinb(w_n222_2[1]),.dout(n226),.clk(gclk));
	jand g0178(.dina(w_n219_1[0]),.dinb(w_n162_1[0]),.dout(n227),.clk(gclk));
	jand g0179(.dina(w_n227_2[1]),.dinb(w_n151_5[1]),.dout(n228),.clk(gclk));
	jnot g0180(.din(w_n228_0[1]),.dout(n229),.clk(gclk));
	jand g0181(.dina(w_n219_0[2]),.dinb(w_n127_1[0]),.dout(n230),.clk(gclk));
	jand g0182(.dina(w_n230_2[1]),.dinb(w_n110_6[0]),.dout(n231),.clk(gclk));
	jnot g0183(.din(w_n231_0[1]),.dout(n232),.clk(gclk));
	jand g0184(.dina(w_n232_2[2]),.dinb(w_n229_2[2]),.dout(n233),.clk(gclk));
	jand g0185(.dina(n233),.dinb(n226),.dout(n234),.clk(gclk));
	jand g0186(.dina(w_n220_3[0]),.dinb(w_n110_5[2]),.dout(n235),.clk(gclk));
	jand g0187(.dina(w_n162_0[2]),.dinb(w_n120_0[0]),.dout(n236),.clk(gclk));
	jand g0188(.dina(w_n236_3[1]),.dinb(w_n211_1[0]),.dout(n237),.clk(gclk));
	jor g0189(.dina(n237),.dinb(w_n235_0[2]),.dout(n238),.clk(gclk));
	jnot g0190(.din(n238),.dout(n239),.clk(gclk));
	jand g0191(.dina(w_n227_2[0]),.dinb(w_n110_5[1]),.dout(n240),.clk(gclk));
	jnot g0192(.din(w_n240_0[2]),.dout(n241),.clk(gclk));
	jnot g0193(.din(w_n223_2[1]),.dout(n242),.clk(gclk));
	jor g0194(.dina(w_n242_0[1]),.dinb(w_n146_4[0]),.dout(n243),.clk(gclk));
	jand g0195(.dina(w_n243_4[2]),.dinb(w_n241_1[1]),.dout(n244),.clk(gclk));
	jand g0196(.dina(n244),.dinb(w_n239_0[1]),.dout(n245),.clk(gclk));
	jand g0197(.dina(n245),.dinb(w_n234_0[1]),.dout(n246),.clk(gclk));
	jand g0198(.dina(w_n140_0[2]),.dinb(w_n134_1[0]),.dout(n247),.clk(gclk));
	jand g0199(.dina(w_n247_2[2]),.dinb(w_n151_5[0]),.dout(n248),.clk(gclk));
	jnot g0200(.din(n248),.dout(n249),.clk(gclk));
	jand g0201(.dina(w_n141_2[0]),.dinb(w_n110_5[0]),.dout(n250),.clk(gclk));
	jnot g0202(.din(w_n250_0[1]),.dout(n251),.clk(gclk));
	jand g0203(.dina(w_n251_3[1]),.dinb(w_n249_2[1]),.dout(n252),.clk(gclk));
	jand g0204(.dina(w_n223_2[0]),.dinb(w_n110_4[2]),.dout(n253),.clk(gclk));
	jnot g0205(.din(n253),.dout(n254),.clk(gclk));
	jand g0206(.dina(w_n151_4[2]),.dinb(w_n141_1[2]),.dout(n255),.clk(gclk));
	jnot g0207(.din(n255),.dout(n256),.clk(gclk));
	jand g0208(.dina(w_n256_2[1]),.dinb(w_n254_3[1]),.dout(n257),.clk(gclk));
	jand g0209(.dina(n257),.dinb(n252),.dout(n258),.clk(gclk));
	jand g0210(.dina(w_n162_0[1]),.dinb(w_n134_0[2]),.dout(n259),.clk(gclk));
	jand g0211(.dina(w_n259_3[1]),.dinb(w_n151_4[1]),.dout(n260),.clk(gclk));
	jnot g0212(.din(w_n260_0[1]),.dout(n261),.clk(gclk));
	jand g0213(.dina(w_n139_0[2]),.dinb(w_n132_0[0]),.dout(n262),.clk(gclk));
	jand g0214(.dina(w_n262_3[2]),.dinb(w_n161_0[1]),.dout(n263),.clk(gclk));
	jnot g0215(.din(w_n263_0[1]),.dout(n264),.clk(gclk));
	jand g0216(.dina(w_n264_2[2]),.dinb(w_n261_1[2]),.dout(n265),.clk(gclk));
	jand g0217(.dina(w_n259_3[0]),.dinb(w_n110_4[1]),.dout(n266),.clk(gclk));
	jnot g0218(.din(w_n266_1[1]),.dout(n267),.clk(gclk));
	jand g0219(.dina(w_n139_0[1]),.dinb(w_n127_0[2]),.dout(n268),.clk(gclk));
	jand g0220(.dina(w_n268_2[2]),.dinb(w_n151_4[0]),.dout(n269),.clk(gclk));
	jnot g0221(.din(w_n269_0[2]),.dout(n270),.clk(gclk));
	jand g0222(.dina(w_n270_2[2]),.dinb(w_n267_1[2]),.dout(n271),.clk(gclk));
	jand g0223(.dina(n271),.dinb(w_n265_0[2]),.dout(n272),.clk(gclk));
	jand g0224(.dina(n272),.dinb(n258),.dout(n273),.clk(gclk));
	jand g0225(.dina(n273),.dinb(w_n246_0[1]),.dout(n274),.clk(gclk));
	jand g0226(.dina(n274),.dinb(w_n218_0[1]),.dout(n275),.clk(gclk));
	jnot g0227(.din(w_n230_2[0]),.dout(n276),.clk(gclk));
	jor g0228(.dina(w_n276_0[2]),.dinb(w_n146_3[2]),.dout(n277),.clk(gclk));
	jand g0229(.dina(w_n220_2[2]),.dinb(w_n212_2[2]),.dout(n278),.clk(gclk));
	jnot g0230(.din(w_n278_0[1]),.dout(n279),.clk(gclk));
	jand g0231(.dina(w_n279_2[1]),.dinb(w_n277_3[1]),.dout(n280),.clk(gclk));
	jnot g0232(.din(w_n220_2[1]),.dout(n281),.clk(gclk));
	jor g0233(.dina(w_n281_0[1]),.dinb(w_n146_3[1]),.dout(n282),.clk(gclk));
	jand g0234(.dina(w_n219_0[1]),.dinb(w_n140_0[1]),.dout(n283),.clk(gclk));
	jand g0235(.dina(w_n283_3[1]),.dinb(w_n110_4[0]),.dout(n284),.clk(gclk));
	jnot g0236(.din(w_n284_0[1]),.dout(n285),.clk(gclk));
	jand g0237(.dina(w_n285_2[1]),.dinb(w_n282_3[1]),.dout(n286),.clk(gclk));
	jand g0238(.dina(w_n286_1[2]),.dinb(w_n280_1[1]),.dout(n287),.clk(gclk));
	jand g0239(.dina(w_n211_0[2]),.dinb(w_n128_2[0]),.dout(n288),.clk(gclk));
	jnot g0240(.din(w_n288_1[1]),.dout(n289),.clk(gclk));
	jand g0241(.dina(w_n283_3[0]),.dinb(w_n151_3[2]),.dout(n290),.clk(gclk));
	jnot g0242(.din(w_n290_0[1]),.dout(n291),.clk(gclk));
	jand g0243(.dina(w_n291_2[1]),.dinb(n289),.dout(n292),.clk(gclk));
	jand g0244(.dina(w_n236_3[0]),.dinb(w_n110_3[2]),.dout(n293),.clk(gclk));
	jnot g0245(.din(n293),.dout(n294),.clk(gclk));
	jor g0246(.dina(w_n154_1[0]),.dinb(w_n146_3[0]),.dout(n295),.clk(gclk));
	jand g0247(.dina(w_n295_3[2]),.dinb(w_n294_3[1]),.dout(n296),.clk(gclk));
	jand g0248(.dina(n296),.dinb(n292),.dout(n297),.clk(gclk));
	jand g0249(.dina(w_n223_1[2]),.dinb(w_n151_3[1]),.dout(n298),.clk(gclk));
	jand g0250(.dina(w_n230_1[2]),.dinb(w_n151_3[0]),.dout(n299),.clk(gclk));
	jor g0251(.dina(w_n299_0[2]),.dinb(w_n298_0[2]),.dout(n300),.clk(gclk));
	jnot g0252(.din(w_n300_0[1]),.dout(n301),.clk(gclk));
	jand g0253(.dina(w_n236_2[2]),.dinb(w_n151_2[2]),.dout(n302),.clk(gclk));
	jnot g0254(.din(n302),.dout(n303),.clk(gclk));
	jor g0255(.dina(w_n215_2[0]),.dinb(w_n154_0[2]),.dout(n304),.clk(gclk));
	jand g0256(.dina(w_n304_3[1]),.dinb(w_n303_4[1]),.dout(n305),.clk(gclk));
	jand g0257(.dina(w_n305_0[2]),.dinb(w_n301_2[2]),.dout(n306),.clk(gclk));
	jand g0258(.dina(n306),.dinb(n297),.dout(n307),.clk(gclk));
	jand g0259(.dina(n307),.dinb(w_n287_0[1]),.dout(n308),.clk(gclk));
	jand g0260(.dina(w_n262_3[1]),.dinb(w_n212_2[1]),.dout(n309),.clk(gclk));
	jnot g0261(.din(w_n309_0[1]),.dout(n310),.clk(gclk));
	jand g0262(.dina(w_n155_1[0]),.dinb(w_n110_3[1]),.dout(n311),.clk(gclk));
	jnot g0263(.din(n311),.dout(n312),.clk(gclk));
	jnot g0264(.din(w_n268_2[1]),.dout(n313),.clk(gclk));
	jor g0265(.dina(n313),.dinb(w_n145_0[2]),.dout(n314),.clk(gclk));
	jand g0266(.dina(w_n163_2[0]),.dinb(w_n109_1[1]),.dout(n315),.clk(gclk));
	jnot g0267(.din(w_n315_0[2]),.dout(n316),.clk(gclk));
	jand g0268(.dina(n316),.dinb(w_n314_1[1]),.dout(n317),.clk(gclk));
	jand g0269(.dina(n317),.dinb(w_n312_3[2]),.dout(n318),.clk(gclk));
	jand g0270(.dina(n318),.dinb(w_n310_1[2]),.dout(n319),.clk(gclk));
	jand g0271(.dina(w_n268_2[0]),.dinb(w_n110_3[0]),.dout(n320),.clk(gclk));
	jnot g0272(.din(w_n320_0[2]),.dout(n321),.clk(gclk));
	jand g0273(.dina(w_n247_2[1]),.dinb(w_n110_2[2]),.dout(n322),.clk(gclk));
	jnot g0274(.din(w_n322_0[1]),.dout(n323),.clk(gclk));
	jand g0275(.dina(w_n323_3[1]),.dinb(w_n321_1[1]),.dout(n324),.clk(gclk));
	jnot g0276(.din(w_n109_1[0]),.dout(n325),.clk(gclk));
	jnot g0277(.din(w_n262_3[0]),.dout(n326),.clk(gclk));
	jand g0278(.dina(w_n134_0[1]),.dinb(w_n127_0[1]),.dout(n327),.clk(gclk));
	jnot g0279(.din(w_n327_2[2]),.dout(n328),.clk(gclk));
	jand g0280(.dina(w_n328_0[2]),.dinb(w_n326_0[1]),.dout(n329),.clk(gclk));
	jor g0281(.dina(n329),.dinb(w_n325_0[1]),.dout(n330),.clk(gclk));
	jand g0282(.dina(n330),.dinb(w_n324_1[1]),.dout(n331),.clk(gclk));
	jand g0283(.dina(n331),.dinb(w_n319_0[1]),.dout(n332),.clk(gclk));
	jand g0284(.dina(n332),.dinb(w_n308_0[1]),.dout(n333),.clk(gclk));
	jand g0285(.dina(n333),.dinb(w_n275_0[1]),.dout(n334),.clk(gclk));
	jnot g0286(.din(w_n334_1[2]),.dout(n335),.clk(gclk));
	jand g0287(.dina(w_n82_0[0]),.dinb(w_n49_3[1]),.dout(n336),.clk(gclk));
	jxor g0288(.dina(w_n336_0[1]),.dinb(w_a7_0[0]),.dout(n337),.clk(gclk));
	jand g0289(.dina(w_n337_5[1]),.dinb(w_n335_6[2]),.dout(n338),.clk(gclk));
	jor g0290(.dina(w_n108_0[2]),.dinb(w_n103_0[1]),.dout(n339),.clk(gclk));
	jor g0291(.dina(w_n339_0[2]),.dinb(w_n96_4[1]),.dout(n340),.clk(gclk));
	jnot g0292(.din(w_n340_2[1]),.dout(n341),.clk(gclk));
	jand g0293(.dina(w_n341_4[1]),.dinb(w_n236_2[1]),.dout(n342),.clk(gclk));
	jnot g0294(.din(w_n342_0[1]),.dout(n343),.clk(gclk));
	jand g0295(.dina(w_n343_2[1]),.dinb(w_n303_4[0]),.dout(n344),.clk(gclk));
	jand g0296(.dina(w_n108_0[1]),.dinb(w_n144_0[1]),.dout(n345),.clk(gclk));
	jand g0297(.dina(w_n345_0[2]),.dinb(w_n143_5[0]),.dout(n346),.clk(gclk));
	jand g0298(.dina(w_n346_7[1]),.dinb(w_n223_1[1]),.dout(n347),.clk(gclk));
	jnot g0299(.din(n347),.dout(n348),.clk(gclk));
	jand g0300(.dina(w_n345_0[1]),.dinb(w_n96_4[0]),.dout(n349),.clk(gclk));
	jand g0301(.dina(w_n349_6[2]),.dinb(w_n247_2[0]),.dout(n350),.clk(gclk));
	jnot g0302(.din(n350),.dout(n351),.clk(gclk));
	jand g0303(.dina(w_n351_2[1]),.dinb(w_n348_2[2]),.dout(n352),.clk(gclk));
	jand g0304(.dina(w_n210_0[0]),.dinb(w_n144_0[0]),.dout(n353),.clk(gclk));
	jand g0305(.dina(w_n353_0[2]),.dinb(w_n96_3[2]),.dout(n354),.clk(gclk));
	jand g0306(.dina(w_n354_4[1]),.dinb(w_n268_1[2]),.dout(n355),.clk(gclk));
	jnot g0307(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jand g0308(.dina(w_n346_7[0]),.dinb(w_n230_1[1]),.dout(n357),.clk(gclk));
	jnot g0309(.din(n357),.dout(n358),.clk(gclk));
	jand g0310(.dina(w_n358_2[1]),.dinb(w_n356_1[2]),.dout(n359),.clk(gclk));
	jand g0311(.dina(n359),.dinb(n352),.dout(n360),.clk(gclk));
	jand g0312(.dina(n360),.dinb(n344),.dout(n361),.clk(gclk));
	jand g0313(.dina(w_n349_6[1]),.dinb(w_n327_2[1]),.dout(n362),.clk(gclk));
	jnot g0314(.din(w_n362_0[1]),.dout(n363),.clk(gclk));
	jand g0315(.dina(w_n349_6[0]),.dinb(w_n163_1[2]),.dout(n364),.clk(gclk));
	jnot g0316(.din(w_n364_0[1]),.dout(n365),.clk(gclk));
	jand g0317(.dina(w_n365_1[2]),.dinb(w_n363_2[1]),.dout(n366),.clk(gclk));
	jor g0318(.dina(w_n339_0[1]),.dinb(w_n143_4[2]),.dout(n367),.clk(gclk));
	jor g0319(.dina(w_n367_2[2]),.dinb(w_n328_0[1]),.dout(n368),.clk(gclk));
	jand g0320(.dina(w_n341_4[0]),.dinb(w_n268_1[1]),.dout(n369),.clk(gclk));
	jnot g0321(.din(w_n369_0[1]),.dout(n370),.clk(gclk));
	jand g0322(.dina(w_n370_2[1]),.dinb(w_n368_2[2]),.dout(n371),.clk(gclk));
	jnot g0323(.din(w_n298_0[1]),.dout(n372),.clk(gclk));
	jand g0324(.dina(w_n349_5[2]),.dinb(w_n220_2[0]),.dout(n373),.clk(gclk));
	jnot g0325(.din(w_n373_0[1]),.dout(n374),.clk(gclk));
	jand g0326(.dina(w_n374_2[2]),.dinb(w_n372_1[2]),.dout(n375),.clk(gclk));
	jand g0327(.dina(n375),.dinb(w_n371_0[1]),.dout(n376),.clk(gclk));
	jand g0328(.dina(n376),.dinb(w_n366_0[1]),.dout(n377),.clk(gclk));
	jand g0329(.dina(w_n349_5[1]),.dinb(w_n259_2[2]),.dout(n378),.clk(gclk));
	jnot g0330(.din(w_n378_0[1]),.dout(n379),.clk(gclk));
	jnot g0331(.din(w_n227_1[2]),.dout(n380),.clk(gclk));
	jor g0332(.dina(w_n380_1[1]),.dinb(w_n146_2[2]),.dout(n381),.clk(gclk));
	jnot g0333(.din(w_n283_2[2]),.dout(n382),.clk(gclk));
	jor g0334(.dina(w_n382_0[1]),.dinb(w_n146_2[1]),.dout(n383),.clk(gclk));
	jand g0335(.dina(w_n383_2[2]),.dinb(w_n381_2[2]),.dout(n384),.clk(gclk));
	jand g0336(.dina(w_n384_1[1]),.dinb(w_n379_1[2]),.dout(n385),.clk(gclk));
	jand g0337(.dina(w_n354_4[0]),.dinb(w_n247_1[2]),.dout(n386),.clk(gclk));
	jnot g0338(.din(w_n386_0[2]),.dout(n387),.clk(gclk));
	jand g0339(.dina(w_n387_1[2]),.dinb(w_n295_3[1]),.dout(n388),.clk(gclk));
	jand g0340(.dina(w_n346_6[2]),.dinb(w_n128_1[2]),.dout(n389),.clk(gclk));
	jnot g0341(.din(w_n389_0[1]),.dout(n390),.clk(gclk));
	jand g0342(.dina(w_n390_1[2]),.dinb(w_n243_4[1]),.dout(n391),.clk(gclk));
	jand g0343(.dina(n391),.dinb(w_n388_0[1]),.dout(n392),.clk(gclk));
	jand g0344(.dina(w_n392_0[2]),.dinb(w_n385_1[1]),.dout(n393),.clk(gclk));
	jand g0345(.dina(n393),.dinb(n377),.dout(n394),.clk(gclk));
	jand g0346(.dina(n394),.dinb(w_n361_0[1]),.dout(n395),.clk(gclk));
	jand g0347(.dina(w_n288_1[0]),.dinb(w_n143_4[1]),.dout(n396),.clk(gclk));
	jnot g0348(.din(n396),.dout(n397),.clk(gclk));
	jand g0349(.dina(w_n397_1[2]),.dinb(w_n214_2[1]),.dout(n398),.clk(gclk));
	jand g0350(.dina(w_n294_3[0]),.dinb(w_n222_2[0]),.dout(n399),.clk(gclk));
	jand g0351(.dina(w_n346_6[1]),.dinb(w_n283_2[1]),.dout(n400),.clk(gclk));
	jnot g0352(.din(w_n400_0[1]),.dout(n401),.clk(gclk));
	jor g0353(.dina(w_n276_0[1]),.dinb(w_n215_1[2]),.dout(n402),.clk(gclk));
	jand g0354(.dina(w_n402_3[1]),.dinb(w_n401_2[2]),.dout(n403),.clk(gclk));
	jand g0355(.dina(w_n403_0[1]),.dinb(w_n399_0[1]),.dout(n404),.clk(gclk));
	jand g0356(.dina(n404),.dinb(w_n398_0[1]),.dout(n405),.clk(gclk));
	jand g0357(.dina(w_n341_3[2]),.dinb(w_n220_1[2]),.dout(n406),.clk(gclk));
	jor g0358(.dina(w_n406_1[1]),.dinb(w_n160_0[1]),.dout(n407),.clk(gclk));
	jnot g0359(.din(w_n407_0[1]),.dout(n408),.clk(gclk));
	jnot g0360(.din(w_n236_2[0]),.dout(n409),.clk(gclk));
	jor g0361(.dina(w_n409_0[1]),.dinb(w_n215_1[1]),.dout(n410),.clk(gclk));
	jand g0362(.dina(w_n346_6[0]),.dinb(w_n268_1[0]),.dout(n411),.clk(gclk));
	jnot g0363(.din(w_n411_0[1]),.dout(n412),.clk(gclk));
	jand g0364(.dina(w_n412_2[1]),.dinb(w_n410_1[2]),.dout(n413),.clk(gclk));
	jand g0365(.dina(w_n354_3[2]),.dinb(w_n230_1[0]),.dout(n414),.clk(gclk));
	jand g0366(.dina(w_n349_5[0]),.dinb(w_n236_1[2]),.dout(n415),.clk(gclk));
	jor g0367(.dina(w_n415_0[2]),.dinb(w_n414_0[1]),.dout(n416),.clk(gclk));
	jnot g0368(.din(n416),.dout(n417),.clk(gclk));
	jand g0369(.dina(w_n417_1[2]),.dinb(w_n413_0[1]),.dout(n418),.clk(gclk));
	jand g0370(.dina(n418),.dinb(w_n408_0[1]),.dout(n419),.clk(gclk));
	jor g0371(.dina(w_n380_1[0]),.dinb(w_n215_1[0]),.dout(n420),.clk(gclk));
	jor g0372(.dina(w_n367_2[1]),.dinb(w_n382_0[0]),.dout(n421),.clk(gclk));
	jor g0373(.dina(w_n367_2[0]),.dinb(w_n380_0[2]),.dout(n422),.clk(gclk));
	jand g0374(.dina(w_n422_2[2]),.dinb(w_n421_3[1]),.dout(n423),.clk(gclk));
	jand g0375(.dina(n423),.dinb(w_n420_2[1]),.dout(n424),.clk(gclk));
	jand g0376(.dina(w_n349_4[2]),.dinb(w_n262_2[2]),.dout(n425),.clk(gclk));
	jnot g0377(.din(w_n425_0[1]),.dout(n426),.clk(gclk));
	jor g0378(.dina(w_n340_2[0]),.dinb(w_n142_0[2]),.dout(n427),.clk(gclk));
	jand g0379(.dina(w_n427_3[1]),.dinb(w_n426_3[2]),.dout(n428),.clk(gclk));
	jand g0380(.dina(w_n341_3[1]),.dinb(w_n223_1[0]),.dout(n429),.clk(gclk));
	jnot g0381(.din(w_n429_0[1]),.dout(n430),.clk(gclk));
	jand g0382(.dina(w_n430_2[2]),.dinb(w_n428_0[2]),.dout(n431),.clk(gclk));
	jand g0383(.dina(n431),.dinb(w_n424_0[1]),.dout(n432),.clk(gclk));
	jand g0384(.dina(n432),.dinb(n419),.dout(n433),.clk(gclk));
	jand g0385(.dina(n433),.dinb(w_n405_0[1]),.dout(n434),.clk(gclk));
	jnot g0386(.din(w_n247_1[1]),.dout(n435),.clk(gclk));
	jor g0387(.dina(w_n435_0[1]),.dinb(w_n215_0[2]),.dout(n436),.clk(gclk));
	jor g0388(.dina(w_n328_0[0]),.dinb(w_n146_2[0]),.dout(n437),.clk(gclk));
	jand g0389(.dina(w_n437_2[1]),.dinb(w_n436_2[2]),.dout(n438),.clk(gclk));
	jand g0390(.dina(n438),.dinb(w_n147_4[0]),.dout(n439),.clk(gclk));
	jand g0391(.dina(w_n349_4[1]),.dinb(w_n230_0[2]),.dout(n440),.clk(gclk));
	jnot g0392(.din(w_n440_0[2]),.dout(n441),.clk(gclk));
	jand g0393(.dina(w_n441_1[2]),.dinb(w_n267_1[1]),.dout(n442),.clk(gclk));
	jand g0394(.dina(n442),.dinb(w_n241_1[0]),.dout(n443),.clk(gclk));
	jand g0395(.dina(w_n354_3[1]),.dinb(w_n135_2[1]),.dout(n444),.clk(gclk));
	jnot g0396(.din(w_n444_0[1]),.dout(n445),.clk(gclk));
	jand g0397(.dina(w_n314_1[0]),.dinb(w_n229_2[1]),.dout(n446),.clk(gclk));
	jand g0398(.dina(n446),.dinb(w_n445_2[2]),.dout(n447),.clk(gclk));
	jand g0399(.dina(n447),.dinb(w_n443_0[1]),.dout(n448),.clk(gclk));
	jand g0400(.dina(n448),.dinb(w_n439_0[1]),.dout(n449),.clk(gclk));
	jand g0401(.dina(w_n346_5[2]),.dinb(w_n227_1[1]),.dout(n450),.clk(gclk));
	jnot g0402(.din(n450),.dout(n451),.clk(gclk));
	jand g0403(.dina(w_n451_3[1]),.dinb(w_n261_1[1]),.dout(n452),.clk(gclk));
	jand g0404(.dina(w_n346_5[1]),.dinb(w_n141_1[1]),.dout(n453),.clk(gclk));
	jnot g0405(.din(w_n453_0[1]),.dout(n454),.clk(gclk));
	jand g0406(.dina(w_n454_2[2]),.dinb(w_n138_4[0]),.dout(n455),.clk(gclk));
	jand g0407(.dina(n455),.dinb(n452),.dout(n456),.clk(gclk));
	jnot g0408(.din(w_n259_2[1]),.dout(n457),.clk(gclk));
	jor g0409(.dina(w_n367_1[2]),.dinb(w_n457_0[1]),.dout(n458),.clk(gclk));
	jand g0410(.dina(w_n458_1[2]),.dinb(w_n249_2[0]),.dout(n459),.clk(gclk));
	jand g0411(.dina(w_n341_3[0]),.dinb(w_n128_1[1]),.dout(n460),.clk(gclk));
	jnot g0412(.din(w_n460_0[1]),.dout(n461),.clk(gclk));
	jnot g0413(.din(w_n163_1[1]),.dout(n462),.clk(gclk));
	jor g0414(.dina(w_n340_1[2]),.dinb(n462),.dout(n463),.clk(gclk));
	jand g0415(.dina(w_n463_3[1]),.dinb(w_n461_2[2]),.dout(n464),.clk(gclk));
	jand g0416(.dina(n464),.dinb(w_n459_0[1]),.dout(n465),.clk(gclk));
	jand g0417(.dina(n465),.dinb(n456),.dout(n466),.clk(gclk));
	jnot g0418(.din(w_n235_0[1]),.dout(n467),.clk(gclk));
	jand g0419(.dina(w_n353_0[1]),.dinb(w_n155_0[2]),.dout(n468),.clk(gclk));
	jand g0420(.dina(w_n468_0[1]),.dinb(w_n143_4[0]),.dout(n469),.clk(gclk));
	jnot g0421(.din(w_n469_0[1]),.dout(n470),.clk(gclk));
	jand g0422(.dina(w_n470_1[2]),.dinb(w_n467_1[1]),.dout(n471),.clk(gclk));
	jand g0423(.dina(w_n354_3[0]),.dinb(w_n262_2[1]),.dout(n472),.clk(gclk));
	jnot g0424(.din(w_n472_0[1]),.dout(n473),.clk(gclk));
	jand g0425(.dina(w_n473_2[1]),.dinb(w_n282_3[0]),.dout(n474),.clk(gclk));
	jand g0426(.dina(w_n345_0[0]),.dinb(w_n155_0[1]),.dout(n475),.clk(gclk));
	jand g0427(.dina(w_n475_1[1]),.dinb(w_n96_3[1]),.dout(n476),.clk(gclk));
	jnot g0428(.din(n476),.dout(n477),.clk(gclk));
	jand g0429(.dina(w_n346_5[0]),.dinb(w_n135_2[0]),.dout(n478),.clk(gclk));
	jnot g0430(.din(w_n478_0[1]),.dout(n479),.clk(gclk));
	jand g0431(.dina(w_n479_2[1]),.dinb(w_n477_2[2]),.dout(n480),.clk(gclk));
	jand g0432(.dina(n480),.dinb(n474),.dout(n481),.clk(gclk));
	jand g0433(.dina(n481),.dinb(w_n471_0[1]),.dout(n482),.clk(gclk));
	jand g0434(.dina(w_n482_0[1]),.dinb(w_n466_0[1]),.dout(n483),.clk(gclk));
	jand g0435(.dina(n483),.dinb(n449),.dout(n484),.clk(gclk));
	jand g0436(.dina(n484),.dinb(w_n434_0[1]),.dout(n485),.clk(gclk));
	jand g0437(.dina(n485),.dinb(w_n395_0[2]),.dout(n486),.clk(gclk));
	jand g0438(.dina(w_n327_2[0]),.dinb(w_n110_2[1]),.dout(n487),.clk(gclk));
	jnot g0439(.din(w_n487_0[1]),.dout(n488),.clk(gclk));
	jand g0440(.dina(w_n488_1[2]),.dinb(w_n277_3[0]),.dout(n489),.clk(gclk));
	jand g0441(.dina(n489),.dinb(w_n270_2[1]),.dout(n490),.clk(gclk));
	jand g0442(.dina(w_n346_4[2]),.dinb(w_n236_1[1]),.dout(n491),.clk(gclk));
	jor g0443(.dina(w_n491_0[1]),.dinb(w_n478_0[0]),.dout(n492),.clk(gclk));
	jnot g0444(.din(n492),.dout(n493),.clk(gclk));
	jand g0445(.dina(w_n426_3[1]),.dinb(w_n310_1[1]),.dout(n494),.clk(gclk));
	jand g0446(.dina(w_n494_0[1]),.dinb(w_n286_1[1]),.dout(n495),.clk(gclk));
	jand g0447(.dina(n495),.dinb(w_n493_0[1]),.dout(n496),.clk(gclk));
	jand g0448(.dina(n496),.dinb(w_n490_0[1]),.dout(n497),.clk(gclk));
	jnot g0449(.din(w_n497_1[1]),.dout(n498),.clk(gclk));
	jnot g0450(.din(w_n406_1[0]),.dout(n499),.clk(gclk));
	jor g0451(.dina(w_n339_0[0]),.dinb(w_n154_0[1]),.dout(n500),.clk(gclk));
	jor g0452(.dina(w_n500_0[1]),.dinb(w_n143_3[2]),.dout(n501),.clk(gclk));
	jand g0453(.dina(w_n501_2[2]),.dinb(w_n368_2[1]),.dout(n502),.clk(gclk));
	jand g0454(.dina(n502),.dinb(w_n499_1[2]),.dout(n503),.clk(gclk));
	jand g0455(.dina(w_n412_2[0]),.dinb(w_n256_2[0]),.dout(n504),.clk(gclk));
	jand g0456(.dina(w_n259_2[0]),.dinb(w_n161_0[0]),.dout(n505),.clk(gclk));
	jnot g0457(.din(w_n505_0[1]),.dout(n506),.clk(gclk));
	jand g0458(.dina(w_n506_2[1]),.dinb(w_n454_2[1]),.dout(n507),.clk(gclk));
	jand g0459(.dina(w_n507_1[1]),.dinb(w_n504_0[2]),.dout(n508),.clk(gclk));
	jand g0460(.dina(n508),.dinb(n503),.dout(n509),.clk(gclk));
	jnot g0461(.din(w_n509_0[2]),.dout(n510),.clk(gclk));
	jand g0462(.dina(w_n463_3[0]),.dinb(w_n304_3[0]),.dout(n511),.clk(gclk));
	jand g0463(.dina(w_n511_1[1]),.dinb(w_n397_1[1]),.dout(n512),.clk(gclk));
	jand g0464(.dina(n512),.dinb(w_n459_0[0]),.dout(n513),.clk(gclk));
	jnot g0465(.din(w_n513_0[2]),.dout(n514),.clk(gclk));
	jor g0466(.dina(w_n367_1[1]),.dinb(w_n281_0[0]),.dout(n515),.clk(gclk));
	jand g0467(.dina(w_n515_2[2]),.dinb(w_n374_2[1]),.dout(n516),.clk(gclk));
	jnot g0468(.din(w_n516_0[1]),.dout(n517),.clk(gclk));
	jand g0469(.dina(w_n262_2[0]),.dinb(w_n151_2[1]),.dout(n518),.clk(gclk));
	jor g0470(.dina(w_n518_0[2]),.dinb(w_n164_0[1]),.dout(n519),.clk(gclk));
	jor g0471(.dina(w_n519_0[1]),.dinb(n517),.dout(n520),.clk(gclk));
	jand g0472(.dina(w_n346_4[1]),.dinb(w_n163_1[0]),.dout(n521),.clk(gclk));
	jor g0473(.dina(w_n521_0[2]),.dinb(w_n440_0[1]),.dout(n522),.clk(gclk));
	jnot g0474(.din(w_n522_0[1]),.dout(n523),.clk(gclk));
	jand g0475(.dina(w_n351_2[0]),.dinb(w_n157_1[1]),.dout(n524),.clk(gclk));
	jand g0476(.dina(w_n524_0[1]),.dinb(w_n523_0[2]),.dout(n525),.clk(gclk));
	jnot g0477(.din(w_n525_0[1]),.dout(n526),.clk(gclk));
	jor g0478(.dina(n526),.dinb(n520),.dout(n527),.clk(gclk));
	jor g0479(.dina(n527),.dinb(n514),.dout(n528),.clk(gclk));
	jor g0480(.dina(n528),.dinb(n510),.dout(n529),.clk(gclk));
	jor g0481(.dina(n529),.dinb(n498),.dout(n530),.clk(gclk));
	jand g0482(.dina(w_n341_2[2]),.dinb(w_n262_1[2]),.dout(n531),.clk(gclk));
	jnot g0483(.din(w_n531_0[1]),.dout(n532),.clk(gclk));
	jand g0484(.dina(w_n532_2[2]),.dinb(w_n390_1[1]),.dout(n533),.clk(gclk));
	jand g0485(.dina(w_n341_2[1]),.dinb(w_n135_1[2]),.dout(n534),.clk(gclk));
	jnot g0486(.din(w_n534_0[1]),.dout(n535),.clk(gclk));
	jand g0487(.dina(w_n535_1[1]),.dinb(w_n130_2[1]),.dout(n536),.clk(gclk));
	jand g0488(.dina(n536),.dinb(n533),.dout(n537),.clk(gclk));
	jand g0489(.dina(n537),.dinb(w_n239_0[0]),.dout(n538),.clk(gclk));
	jnot g0490(.din(w_n538_0[2]),.dout(n539),.clk(gclk));
	jand g0491(.dina(w_n401_2[1]),.dinb(w_n138_3[2]),.dout(n540),.clk(gclk));
	jand g0492(.dina(n540),.dinb(w_n225_2[1]),.dout(n541),.clk(gclk));
	jnot g0493(.din(w_n541_0[1]),.dout(n542),.clk(gclk));
	jand g0494(.dina(w_n348_2[1]),.dinb(w_n251_3[0]),.dout(n543),.clk(gclk));
	jnot g0495(.din(w_n543_1[1]),.dout(n544),.clk(gclk));
	jor g0496(.dina(w_n298_0[0]),.dinb(w_n278_0[0]),.dout(n545),.clk(gclk));
	jor g0497(.dina(w_n545_0[1]),.dinb(n544),.dout(n546),.clk(gclk));
	jor g0498(.dina(n546),.dinb(n542),.dout(n547),.clk(gclk));
	jand g0499(.dina(w_n349_4[0]),.dinb(w_n135_1[1]),.dout(n548),.clk(gclk));
	jor g0500(.dina(w_n548_0[1]),.dinb(w_n444_0[0]),.dout(n549),.clk(gclk));
	jor g0501(.dina(n549),.dinb(w_n472_0[0]),.dout(n550),.clk(gclk));
	jand g0502(.dina(w_n327_1[2]),.dinb(w_n212_2[0]),.dout(n551),.clk(gclk));
	jand g0503(.dina(w_n354_2[2]),.dinb(w_n236_1[0]),.dout(n552),.clk(gclk));
	jor g0504(.dina(w_n552_0[2]),.dinb(w_n551_0[2]),.dout(n553),.clk(gclk));
	jand g0505(.dina(w_n346_4[0]),.dinb(w_n262_1[1]),.dout(n554),.clk(gclk));
	jor g0506(.dina(w_n554_0[2]),.dinb(w_n429_0[0]),.dout(n555),.clk(gclk));
	jor g0507(.dina(n555),.dinb(n553),.dout(n556),.clk(gclk));
	jor g0508(.dina(w_n556_0[1]),.dinb(w_n550_0[1]),.dout(n557),.clk(gclk));
	jor g0509(.dina(w_n557_0[1]),.dinb(n547),.dout(n558),.clk(gclk));
	jor g0510(.dina(n558),.dinb(n539),.dout(n559),.clk(gclk));
	jand g0511(.dina(w_n262_1[0]),.dinb(w_n110_2[0]),.dout(n560),.clk(gclk));
	jnot g0512(.din(w_n560_0[1]),.dout(n561),.clk(gclk));
	jand g0513(.dina(w_n475_1[0]),.dinb(w_n143_3[1]),.dout(n562),.clk(gclk));
	jnot g0514(.din(w_n562_0[1]),.dout(n563),.clk(gclk));
	jand g0515(.dina(w_n563_0[2]),.dinb(w_n561_2[1]),.dout(n564),.clk(gclk));
	jand g0516(.dina(w_n564_0[1]),.dinb(w_n356_1[1]),.dout(n565),.clk(gclk));
	jnot g0517(.din(w_n565_1[1]),.dout(n566),.clk(gclk));
	jand g0518(.dina(w_n381_2[1]),.dinb(w_n232_2[1]),.dout(n567),.clk(gclk));
	jand g0519(.dina(n567),.dinb(w_n295_3[0]),.dout(n568),.clk(gclk));
	jnot g0520(.din(w_n568_0[2]),.dout(n569),.clk(gclk));
	jor g0521(.dina(w_n342_0[0]),.dinb(w_n320_0[1]),.dout(n570),.clk(gclk));
	jor g0522(.dina(n570),.dinb(w_n240_0[1]),.dout(n571),.clk(gclk));
	jor g0523(.dina(w_n571_0[2]),.dinb(n569),.dout(n572),.clk(gclk));
	jor g0524(.dina(n572),.dinb(n566),.dout(n573),.clk(gclk));
	jand g0525(.dina(w_n354_2[1]),.dinb(w_n163_0[2]),.dout(n574),.clk(gclk));
	jor g0526(.dina(w_n574_0[2]),.dinb(w_n266_1[0]),.dout(n575),.clk(gclk));
	jor g0527(.dina(n575),.dinb(w_n386_0[1]),.dout(n576),.clk(gclk));
	jnot g0528(.din(w_n420_2[0]),.dout(n577),.clk(gclk));
	jor g0529(.dina(w_n577_0[1]),.dinb(w_n213_1[0]),.dout(n578),.clk(gclk));
	jor g0530(.dina(w_n314_0[2]),.dinb(w_n143_3[0]),.dout(n579),.clk(gclk));
	jnot g0531(.din(w_n579_2[2]),.dout(n580),.clk(gclk));
	jand g0532(.dina(w_n288_0[2]),.dinb(w_n96_3[0]),.dout(n581),.clk(gclk));
	jor g0533(.dina(w_n581_0[1]),.dinb(w_n580_0[1]),.dout(n582),.clk(gclk));
	jor g0534(.dina(n582),.dinb(w_n578_0[1]),.dout(n583),.clk(gclk));
	jor g0535(.dina(n583),.dinb(n576),.dout(n584),.clk(gclk));
	jnot g0536(.din(w_n437_2[0]),.dout(n585),.clk(gclk));
	jand g0537(.dina(w_n341_2[0]),.dinb(w_n327_1[1]),.dout(n586),.clk(gclk));
	jor g0538(.dina(w_n586_0[1]),.dinb(n585),.dout(n587),.clk(gclk));
	jand g0539(.dina(w_n341_1[2]),.dinb(w_n247_1[0]),.dout(n588),.clk(gclk));
	jor g0540(.dina(w_n588_1[1]),.dinb(w_n263_0[0]),.dout(n589),.clk(gclk));
	jor g0541(.dina(n589),.dinb(w_n587_0[1]),.dout(n590),.clk(gclk));
	jand g0542(.dina(w_n349_3[2]),.dinb(w_n227_1[0]),.dout(n591),.clk(gclk));
	jnot g0543(.din(w_n591_0[1]),.dout(n592),.clk(gclk));
	jand g0544(.dina(w_n346_3[2]),.dinb(w_n247_0[2]),.dout(n593),.clk(gclk));
	jnot g0545(.din(w_n593_0[1]),.dout(n594),.clk(gclk));
	jand g0546(.dina(w_n594_2[2]),.dinb(w_n592_3[1]),.dout(n595),.clk(gclk));
	jor g0547(.dina(w_n340_1[1]),.dinb(w_n457_0[0]),.dout(n596),.clk(gclk));
	jand g0548(.dina(w_n596_0[2]),.dinb(w_n243_4[0]),.dout(n597),.clk(gclk));
	jand g0549(.dina(w_n597_2[1]),.dinb(w_n595_0[2]),.dout(n598),.clk(gclk));
	jnot g0550(.din(w_n598_0[1]),.dout(n599),.clk(gclk));
	jor g0551(.dina(n599),.dinb(w_n590_0[1]),.dout(n600),.clk(gclk));
	jor g0552(.dina(n600),.dinb(w_n584_0[1]),.dout(n601),.clk(gclk));
	jor g0553(.dina(n601),.dinb(n573),.dout(n602),.clk(gclk));
	jor g0554(.dina(n602),.dinb(n559),.dout(n603),.clk(gclk));
	jor g0555(.dina(n603),.dinb(n530),.dout(n604),.clk(gclk));
	jnot g0556(.din(w_n556_0[0]),.dout(n605),.clk(gclk));
	jand g0557(.dina(w_n349_3[1]),.dinb(w_n141_1[0]),.dout(n606),.clk(gclk));
	jor g0558(.dina(w_n606_0[2]),.dinb(w_n518_0[1]),.dout(n607),.clk(gclk));
	jand g0559(.dina(w_n315_0[1]),.dinb(w_n143_2[2]),.dout(n608),.clk(gclk));
	jor g0560(.dina(w_n608_0[2]),.dinb(w_n269_0[1]),.dout(n609),.clk(gclk));
	jor g0561(.dina(n609),.dinb(n607),.dout(n610),.clk(gclk));
	jnot g0562(.din(n610),.dout(n611),.clk(gclk));
	jor g0563(.dina(w_n367_1[0]),.dinb(w_n242_0[0]),.dout(n612),.clk(gclk));
	jand g0564(.dina(w_n327_1[0]),.dinb(w_n151_2[0]),.dout(n613),.clk(gclk));
	jnot g0565(.din(n613),.dout(n614),.clk(gclk));
	jand g0566(.dina(w_n614_2[2]),.dinb(w_n612_3[2]),.dout(n615),.clk(gclk));
	jand g0567(.dina(n615),.dinb(w_n232_2[0]),.dout(n616),.clk(gclk));
	jand g0568(.dina(n616),.dinb(w_n611_1[1]),.dout(n617),.clk(gclk));
	jand g0569(.dina(n617),.dinb(w_n605_0[1]),.dout(n618),.clk(gclk));
	jand g0570(.dina(w_n249_1[2]),.dinb(w_n229_2[0]),.dout(n619),.clk(gclk));
	jand g0571(.dina(w_n561_2[0]),.dinb(w_n216_4[0]),.dout(n620),.clk(gclk));
	jand g0572(.dina(n620),.dinb(w_n294_2[2]),.dout(n621),.clk(gclk));
	jand g0573(.dina(n621),.dinb(w_n619_1[2]),.dout(n622),.clk(gclk));
	jand g0574(.dina(w_n379_1[1]),.dinb(w_n251_2[2]),.dout(n623),.clk(gclk));
	jor g0575(.dina(w_n314_0[1]),.dinb(w_n96_2[2]),.dout(n624),.clk(gclk));
	jand g0576(.dina(w_n624_2[2]),.dinb(w_n454_2[0]),.dout(n625),.clk(gclk));
	jand g0577(.dina(w_n436_2[1]),.dinb(w_n264_2[1]),.dout(n626),.clk(gclk));
	jand g0578(.dina(w_n626_1[1]),.dinb(w_n625_0[1]),.dout(n627),.clk(gclk));
	jand g0579(.dina(n627),.dinb(w_n623_0[1]),.dout(n628),.clk(gclk));
	jand g0580(.dina(n628),.dinb(w_n622_1[2]),.dout(n629),.clk(gclk));
	jand g0581(.dina(n629),.dinb(n618),.dout(n630),.clk(gclk));
	jand g0582(.dina(w_n315_0[0]),.dinb(w_n96_2[1]),.dout(n631),.clk(gclk));
	jnot g0583(.din(w_n631_0[2]),.dout(n632),.clk(gclk));
	jand g0584(.dina(w_n632_2[1]),.dinb(w_n303_3[2]),.dout(n633),.clk(gclk));
	jand g0585(.dina(w_n499_1[1]),.dinb(w_n343_2[0]),.dout(n634),.clk(gclk));
	jand g0586(.dina(n634),.dinb(w_n633_0[1]),.dout(n635),.clk(gclk));
	jand g0587(.dina(n635),.dinb(w_n630_0[1]),.dout(n636),.clk(gclk));
	jor g0588(.dina(w_n487_0[0]),.dinb(w_n240_0[0]),.dout(n637),.clk(gclk));
	jnot g0589(.din(w_n637_0[1]),.dout(n638),.clk(gclk));
	jand g0590(.dina(w_n515_2[1]),.dinb(w_n312_3[1]),.dout(n639),.clk(gclk));
	jand g0591(.dina(n639),.dinb(w_n638_0[2]),.dout(n640),.clk(gclk));
	jand g0592(.dina(w_n283_2[0]),.dinb(w_n212_1[2]),.dout(n641),.clk(gclk));
	jnot g0593(.din(w_n641_0[1]),.dout(n642),.clk(gclk));
	jand g0594(.dina(w_n642_1[2]),.dinb(w_n402_3[0]),.dout(n643),.clk(gclk));
	jand g0595(.dina(w_n346_3[1]),.dinb(w_n259_1[2]),.dout(n644),.clk(gclk));
	jnot g0596(.din(w_n644_0[1]),.dout(n645),.clk(gclk));
	jand g0597(.dina(w_n645_2[1]),.dinb(w_n356_1[0]),.dout(n646),.clk(gclk));
	jand g0598(.dina(w_n646_0[2]),.dinb(w_n643_0[1]),.dout(n647),.clk(gclk));
	jand g0599(.dina(n647),.dinb(n640),.dout(n648),.clk(gclk));
	jnot g0600(.din(w_n304_2[2]),.dout(n649),.clk(gclk));
	jor g0601(.dina(w_n562_0[0]),.dinb(w_n440_0[0]),.dout(n650),.clk(gclk));
	jor g0602(.dina(w_n650_0[1]),.dinb(n649),.dout(n651),.clk(gclk));
	jnot g0603(.din(w_n381_2[0]),.dout(n652),.clk(gclk));
	jor g0604(.dina(w_n469_0[0]),.dinb(n652),.dout(n653),.clk(gclk));
	jor g0605(.dina(n653),.dinb(w_n651_0[1]),.dout(n654),.clk(gclk));
	jnot g0606(.din(n654),.dout(n655),.clk(gclk));
	jand g0607(.dina(w_n532_2[1]),.dinb(w_n348_2[0]),.dout(n656),.clk(gclk));
	jand g0608(.dina(n656),.dinb(w_n225_2[0]),.dout(n657),.clk(gclk));
	jand g0609(.dina(n657),.dinb(w_n301_2[1]),.dout(n658),.clk(gclk));
	jand g0610(.dina(n658),.dinb(w_n655_0[1]),.dout(n659),.clk(gclk));
	jand g0611(.dina(n659),.dinb(w_n648_0[1]),.dout(n660),.clk(gclk));
	jand g0612(.dina(w_n349_3[0]),.dinb(w_n223_0[2]),.dout(n661),.clk(gclk));
	jnot g0613(.din(w_n661_0[1]),.dout(n662),.clk(gclk));
	jnot g0614(.din(w_n135_1[0]),.dout(n663),.clk(gclk));
	jor g0615(.dina(w_n145_0[1]),.dinb(n663),.dout(n664),.clk(gclk));
	jor g0616(.dina(w_n664_0[2]),.dinb(w_n143_2[1]),.dout(n665),.clk(gclk));
	jand g0617(.dina(w_n665_2[2]),.dinb(w_n662_2[2]),.dout(n666),.clk(gclk));
	jand g0618(.dina(n666),.dinb(w_n477_2[1]),.dout(n667),.clk(gclk));
	jnot g0619(.din(w_n548_0[0]),.dout(n668),.clk(gclk));
	jand g0620(.dina(w_n668_2[2]),.dinb(w_n451_3[0]),.dout(n669),.clk(gclk));
	jand g0621(.dina(w_n346_3[0]),.dinb(w_n220_1[1]),.dout(n670),.clk(gclk));
	jor g0622(.dina(w_n670_0[2]),.dinb(w_n320_0[0]),.dout(n671),.clk(gclk));
	jnot g0623(.din(n671),.dout(n672),.clk(gclk));
	jand g0624(.dina(n672),.dinb(w_n398_0[0]),.dout(n673),.clk(gclk));
	jand g0625(.dina(n673),.dinb(w_n669_0[1]),.dout(n674),.clk(gclk));
	jand g0626(.dina(n674),.dinb(w_n667_0[1]),.dout(n675),.clk(gclk));
	jand g0627(.dina(w_n579_2[1]),.dinb(w_n410_1[1]),.dout(n676),.clk(gclk));
	jand g0628(.dina(w_n676_1[1]),.dinb(w_n461_2[1]),.dout(n677),.clk(gclk));
	jand g0629(.dina(w_n354_2[0]),.dinb(w_n128_1[0]),.dout(n678),.clk(gclk));
	jnot g0630(.din(w_n678_0[1]),.dout(n679),.clk(gclk));
	jand g0631(.dina(w_n679_2[1]),.dinb(w_n473_2[0]),.dout(n680),.clk(gclk));
	jand g0632(.dina(w_n506_2[0]),.dinb(w_n256_1[2]),.dout(n681),.clk(gclk));
	jand g0633(.dina(w_n479_2[0]),.dinb(w_n279_2[0]),.dout(n682),.clk(gclk));
	jand g0634(.dina(n682),.dinb(w_n681_0[1]),.dout(n683),.clk(gclk));
	jand g0635(.dina(n683),.dinb(w_n680_1[1]),.dout(n684),.clk(gclk));
	jand g0636(.dina(n684),.dinb(w_n677_0[2]),.dout(n685),.clk(gclk));
	jand g0637(.dina(w_n685_0[1]),.dinb(w_n675_0[2]),.dout(n686),.clk(gclk));
	jand g0638(.dina(n686),.dinb(n660),.dout(n687),.clk(gclk));
	jand g0639(.dina(n687),.dinb(w_n636_0[1]),.dout(n688),.clk(gclk));
	jnot g0640(.din(w_n688_0[2]),.dout(n689),.clk(gclk));
	jand g0641(.dina(n689),.dinb(w_n604_0[2]),.dout(n690),.clk(gclk));
	jor g0642(.dina(w_n690_0[1]),.dinb(w_n486_1[1]),.dout(n691),.clk(gclk));
	jand g0643(.dina(w_n691_1[2]),.dinb(w_n338_1[1]),.dout(n692),.clk(gclk));
	jxor g0644(.dina(w_n691_1[1]),.dinb(w_n338_1[0]),.dout(n693),.clk(gclk));
	jand g0645(.dina(w_a22_4[0]),.dinb(w_a8_0[2]),.dout(n694),.clk(gclk));
	jand g0646(.dina(w_n84_0[0]),.dinb(w_n49_3[0]),.dout(n695),.clk(gclk));
	jand g0647(.dina(w_n83_0[0]),.dinb(w_a8_0[1]),.dout(n696),.clk(gclk));
	jnot g0648(.din(n696),.dout(n697),.clk(gclk));
	jand g0649(.dina(n697),.dinb(w_n695_0[1]),.dout(n698),.clk(gclk));
	jor g0650(.dina(n698),.dinb(n694),.dout(n699),.clk(gclk));
	jand g0651(.dina(w_n699_13[2]),.dinb(w_n335_6[1]),.dout(n700),.clk(gclk));
	jand g0652(.dina(w_n700_0[1]),.dinb(w_n693_0[1]),.dout(n701),.clk(gclk));
	jor g0653(.dina(n701),.dinb(n692),.dout(n702),.clk(gclk));
	jand g0654(.dina(w_a22_3[2]),.dinb(w_a10_0[2]),.dout(n703),.clk(gclk));
	jand g0655(.dina(w_n86_0[0]),.dinb(w_n49_2[2]),.dout(n704),.clk(gclk));
	jand g0656(.dina(w_n85_0[0]),.dinb(w_a10_0[1]),.dout(n705),.clk(gclk));
	jnot g0657(.din(n705),.dout(n706),.clk(gclk));
	jand g0658(.dina(n706),.dinb(w_n704_0[1]),.dout(n707),.clk(gclk));
	jor g0659(.dina(n707),.dinb(n703),.dout(n708),.clk(gclk));
	jnot g0660(.din(w_n574_0[1]),.dout(n709),.clk(gclk));
	jor g0661(.dina(w_n367_0[2]),.dinb(w_n142_0[1]),.dout(n710),.clk(gclk));
	jand g0662(.dina(w_n710_3[1]),.dinb(w_n709_1[1]),.dout(n711),.clk(gclk));
	jand g0663(.dina(w_n642_1[1]),.dinb(w_n420_1[2]),.dout(n712),.clk(gclk));
	jand g0664(.dina(w_n532_2[0]),.dinb(w_n427_3[0]),.dout(n713),.clk(gclk));
	jand g0665(.dina(w_n713_0[1]),.dinb(w_n712_0[2]),.dout(n714),.clk(gclk));
	jand g0666(.dina(n714),.dinb(w_n711_0[1]),.dout(n715),.clk(gclk));
	jand g0667(.dina(w_n473_1[2]),.dinb(w_n370_2[0]),.dout(n716),.clk(gclk));
	jand g0668(.dina(n716),.dinb(w_n646_0[1]),.dout(n717),.clk(gclk));
	jand g0669(.dina(n717),.dinb(w_n385_1[0]),.dout(n718),.clk(gclk));
	jand g0670(.dina(n718),.dinb(n715),.dout(n719),.clk(gclk));
	jand g0671(.dina(w_n500_0[0]),.dinb(w_n463_2[2]),.dout(n720),.clk(gclk));
	jand g0672(.dina(n720),.dinb(w_n679_2[0]),.dout(n721),.clk(gclk));
	jand g0673(.dina(n721),.dinb(w_n719_1[1]),.dout(n722),.clk(gclk));
	jand g0674(.dina(w_n259_1[1]),.dinb(w_n212_1[1]),.dout(n723),.clk(gclk));
	jnot g0675(.din(n723),.dout(n724),.clk(gclk));
	jand g0676(.dina(w_n211_0[1]),.dinb(w_n135_0[2]),.dout(n725),.clk(gclk));
	jand g0677(.dina(w_n725_0[1]),.dinb(w_n96_2[0]),.dout(n726),.clk(gclk));
	jor g0678(.dina(w_n726_0[1]),.dinb(w_n551_0[1]),.dout(n727),.clk(gclk));
	jnot g0679(.din(w_n727_0[1]),.dout(n728),.clk(gclk));
	jand g0680(.dina(w_n728_0[1]),.dinb(w_n724_2[2]),.dout(n729),.clk(gclk));
	jnot g0681(.din(w_n554_0[1]),.dout(n730),.clk(gclk));
	jand g0682(.dina(w_n730_1[1]),.dinb(w_n402_2[2]),.dout(n731),.clk(gclk));
	jor g0683(.dina(w_n435_0[0]),.dinb(w_n146_1[2]),.dout(n732),.clk(gclk));
	jand g0684(.dina(w_n732_3[1]),.dinb(w_n437_1[2]),.dout(n733),.clk(gclk));
	jnot g0685(.din(w_n521_0[1]),.dout(n734),.clk(gclk));
	jand g0686(.dina(w_n734_1[2]),.dinb(w_n506_1[2]),.dout(n735),.clk(gclk));
	jand g0687(.dina(w_n735_0[1]),.dinb(w_n733_1[1]),.dout(n736),.clk(gclk));
	jand g0688(.dina(n736),.dinb(w_n731_0[2]),.dout(n737),.clk(gclk));
	jand g0689(.dina(n737),.dinb(n729),.dout(n738),.clk(gclk));
	jnot g0690(.din(w_n606_0[1]),.dout(n739),.clk(gclk));
	jand g0691(.dina(w_n739_0[2]),.dinb(w_n365_1[1]),.dout(n740),.clk(gclk));
	jand g0692(.dina(w_n740_0[1]),.dinb(w_n454_1[2]),.dout(n741),.clk(gclk));
	jnot g0693(.din(w_n475_0[2]),.dout(n742),.clk(gclk));
	jand g0694(.dina(w_n349_2[2]),.dinb(w_n268_0[2]),.dout(n743),.clk(gclk));
	jnot g0695(.din(n743),.dout(n744),.clk(gclk));
	jand g0696(.dina(w_n744_2[2]),.dinb(w_n742_0[1]),.dout(n745),.clk(gclk));
	jand g0697(.dina(n745),.dinb(w_n741_1[1]),.dout(n746),.clk(gclk));
	jand g0698(.dina(w_n436_2[0]),.dinb(w_n412_1[2]),.dout(n747),.clk(gclk));
	jand g0699(.dina(w_n725_0[0]),.dinb(w_n143_2[0]),.dout(n748),.clk(gclk));
	jnot g0700(.din(w_n748_1[1]),.dout(n749),.clk(gclk));
	jand g0701(.dina(w_n349_2[1]),.dinb(w_n128_0[2]),.dout(n750),.clk(gclk));
	jnot g0702(.din(w_n750_0[1]),.dout(n751),.clk(gclk));
	jand g0703(.dina(w_n751_2[1]),.dinb(w_n426_3[0]),.dout(n752),.clk(gclk));
	jand g0704(.dina(n752),.dinb(w_n749_1[1]),.dout(n753),.clk(gclk));
	jand g0705(.dina(n753),.dinb(n747),.dout(n754),.clk(gclk));
	jand g0706(.dina(w_n754_0[1]),.dinb(w_n746_0[2]),.dout(n755),.clk(gclk));
	jand g0707(.dina(n755),.dinb(n738),.dout(n756),.clk(gclk));
	jnot g0708(.din(w_n552_0[1]),.dout(n757),.clk(gclk));
	jand g0709(.dina(w_n612_3[1]),.dinb(w_n757_0[1]),.dout(n758),.clk(gclk));
	jand g0710(.dina(w_n461_2[0]),.dinb(w_n430_2[1]),.dout(n759),.clk(gclk));
	jand g0711(.dina(n759),.dinb(w_n758_0[1]),.dout(n760),.clk(gclk));
	jand g0712(.dina(n760),.dinb(w_n756_0[1]),.dout(n761),.clk(gclk));
	jand g0713(.dina(n761),.dinb(w_n722_0[1]),.dout(n762),.clk(gclk));
	jnot g0714(.din(w_n670_0[1]),.dout(n763),.clk(gclk));
	jand g0715(.dina(w_n349_2[0]),.dinb(w_n283_1[2]),.dout(n764),.clk(gclk));
	jnot g0716(.din(w_n764_0[2]),.dout(n765),.clk(gclk));
	jand g0717(.dina(w_n765_1[2]),.dinb(w_n763_2[1]),.dout(n766),.clk(gclk));
	jand g0718(.dina(n766),.dinb(w_n358_2[0]),.dout(n767),.clk(gclk));
	jnot g0719(.din(w_n415_0[1]),.dout(n768),.clk(gclk));
	jand g0720(.dina(w_n662_2[1]),.dinb(w_n441_1[1]),.dout(n769),.clk(gclk));
	jand g0721(.dina(n769),.dinb(w_n768_2[2]),.dout(n770),.clk(gclk));
	jand g0722(.dina(w_n390_1[0]),.dinb(w_n374_2[0]),.dout(n771),.clk(gclk));
	jnot g0723(.din(w_n491_0[0]),.dout(n772),.clk(gclk));
	jand g0724(.dina(w_n772_2[2]),.dinb(w_n348_1[2]),.dout(n773),.clk(gclk));
	jand g0725(.dina(w_n773_0[1]),.dinb(w_n771_2[1]),.dout(n774),.clk(gclk));
	jand g0726(.dina(n774),.dinb(n770),.dout(n775),.clk(gclk));
	jand g0727(.dina(n775),.dinb(w_n767_0[1]),.dout(n776),.clk(gclk));
	jand g0728(.dina(w_n712_0[1]),.dinb(w_n384_1[0]),.dout(n777),.clk(gclk));
	jand g0729(.dina(n777),.dinb(w_n776_0[1]),.dout(n778),.clk(gclk));
	jand g0730(.dina(n778),.dinb(w_n756_0[0]),.dout(n779),.clk(gclk));
	jand g0731(.dina(w_n346_2[2]),.dinb(w_n327_0[2]),.dout(n780),.clk(gclk));
	jnot g0732(.din(w_n780_0[1]),.dout(n781),.clk(gclk));
	jand g0733(.dina(w_n781_2[1]),.dinb(w_n479_1[2]),.dout(n782),.clk(gclk));
	jand g0734(.dina(n782),.dinb(w_n351_1[2]),.dout(n783),.clk(gclk));
	jand g0735(.dina(n783),.dinb(w_n595_0[1]),.dout(n784),.clk(gclk));
	jand g0736(.dina(w_n669_0[0]),.dinb(w_n363_2[0]),.dout(n785),.clk(gclk));
	jand g0737(.dina(n785),.dinb(w_n784_0[1]),.dout(n786),.clk(gclk));
	jand g0738(.dina(w_n786_1[1]),.dinb(w_n401_2[0]),.dout(n787),.clk(gclk));
	jand g0739(.dina(n787),.dinb(w_n779_0[1]),.dout(n788),.clk(gclk));
	jxor g0740(.dina(w_n788_0[2]),.dinb(w_n762_2[1]),.dout(n789),.clk(gclk));
	jnot g0741(.din(w_n762_2[0]),.dout(n790),.clk(gclk));
	jor g0742(.dina(w_n790_0[2]),.dinb(w_n789_5[1]),.dout(n792),.clk(gclk));
	jand g0743(.dina(w_n792_0[2]),.dinb(w_n708_6[1]),.dout(n793),.clk(gclk));
	jnot g0744(.din(w_n708_6[0]),.dout(n794),.clk(gclk));
	jnot g0745(.din(w_n789_5[0]),.dout(n795),.clk(gclk));
	jor g0746(.dina(w_n788_0[1]),.dinb(w_n762_1[2]),.dout(n796),.clk(gclk));
	jand g0747(.dina(w_n334_1[1]),.dinb(w_n795_1[1]),.dout(n799),.clk(gclk));
	jnot g0748(.din(w_n799_3[2]),.dout(n800),.clk(gclk));
	jand g0749(.dina(w_n800_0[2]),.dinb(w_n794_4[2]),.dout(n801),.clk(gclk));
	jor g0750(.dina(n801),.dinb(n793),.dout(n802),.clk(gclk));
	jxor g0751(.dina(w_n704_0[0]),.dinb(w_a11_0[0]),.dout(n803),.clk(gclk));
	jand g0752(.dina(w_n788_0[0]),.dinb(w_n762_1[1]),.dout(n804),.clk(gclk));
	jnot g0753(.din(w_n803_8[2]),.dout(n808),.clk(gclk));
	jand g0754(.dina(w_n789_4[2]),.dinb(w_n808_13[2]),.dout(n810),.clk(gclk));
	jnot g0755(.din(n810),.dout(n812),.clk(gclk));
	jand g0756(.dina(n812),.dinb(n802),.dout(n813),.clk(gclk));
	jand g0757(.dina(w_n813_0[1]),.dinb(w_n702_0[1]),.dout(n814),.clk(gclk));
	jand g0758(.dina(w_a22_3[1]),.dinb(w_a14_0[2]),.dout(n815),.clk(gclk));
	jnot g0759(.din(n815),.dout(n816),.clk(gclk));
	jand g0760(.dina(w_n89_0[0]),.dinb(w_a14_0[1]),.dout(n817),.clk(gclk));
	jor g0761(.dina(n817),.dinb(w_a22_3[0]),.dout(n818),.clk(gclk));
	jor g0762(.dina(n818),.dinb(w_n201_0[0]),.dout(n819),.clk(gclk));
	jand g0763(.dina(n819),.dinb(n816),.dout(n820),.clk(gclk));
	jand g0764(.dina(w_n744_2[1]),.dinb(w_n401_1[2]),.dout(n821),.clk(gclk));
	jand g0765(.dina(w_n515_2[0]),.dinb(w_n321_1[0]),.dout(n822),.clk(gclk));
	jand g0766(.dina(w_n822_2[1]),.dinb(w_n821_1[1]),.dout(n823),.clk(gclk));
	jand g0767(.dina(n823),.dinb(w_n158_1[0]),.dout(n824),.clk(gclk));
	jnot g0768(.din(w_n414_0[0]),.dout(n825),.clk(gclk));
	jand g0769(.dina(w_n825_1[2]),.dinb(w_n467_1[0]),.dout(n826),.clk(gclk));
	jand g0770(.dina(n826),.dinb(w_n579_2[0]),.dout(n827),.clk(gclk));
	jand g0771(.dina(w_n254_3[0]),.dinb(w_n222_1[2]),.dout(n828),.clk(gclk));
	jand g0772(.dina(n828),.dinb(w_n301_2[0]),.dout(n829),.clk(gclk));
	jand g0773(.dina(n829),.dinb(w_n504_0[1]),.dout(n830),.clk(gclk));
	jand g0774(.dina(n830),.dinb(n827),.dout(n831),.clk(gclk));
	jand g0775(.dina(n831),.dinb(w_n824_0[1]),.dout(n832),.clk(gclk));
	jand g0776(.dina(w_n451_2[2]),.dinb(w_n294_2[1]),.dout(n833),.clk(gclk));
	jand g0777(.dina(n833),.dinb(w_n832_1[1]),.dout(n834),.clk(gclk));
	jand g0778(.dina(w_n561_1[2]),.dinb(w_n312_3[0]),.dout(n835),.clk(gclk));
	jand g0779(.dina(n835),.dinb(w_n130_2[0]),.dout(n836),.clk(gclk));
	jnot g0780(.din(w_n586_0[0]),.dout(n837),.clk(gclk));
	jand g0781(.dina(w_n402_2[1]),.dinb(w_n270_2[0]),.dout(n838),.clk(gclk));
	jand g0782(.dina(n838),.dinb(w_n837_2[1]),.dout(n839),.clk(gclk));
	jand g0783(.dina(n839),.dinb(w_n836_0[1]),.dout(n840),.clk(gclk));
	jnot g0784(.din(w_n550_0[0]),.dout(n841),.clk(gclk));
	jand g0785(.dina(w_n501_2[1]),.dinb(w_n216_3[2]),.dout(n842),.clk(gclk));
	jand g0786(.dina(n842),.dinb(w_n147_3[2]),.dout(n843),.clk(gclk));
	jand g0787(.dina(w_n843_0[1]),.dinb(n841),.dout(n844),.clk(gclk));
	jand g0788(.dina(n844),.dinb(n840),.dout(n845),.clk(gclk));
	jand g0789(.dina(w_n662_2[0]),.dinb(w_n470_1[1]),.dout(n846),.clk(gclk));
	jand g0790(.dina(w_n632_2[0]),.dinb(w_n304_2[1]),.dout(n847),.clk(gclk));
	jand g0791(.dina(n847),.dinb(w_n846_0[1]),.dout(n848),.clk(gclk));
	jnot g0792(.din(w_n608_0[1]),.dout(n849),.clk(gclk));
	jand g0793(.dina(w_n849_2[1]),.dinb(w_n420_1[1]),.dout(n850),.clk(gclk));
	jand g0794(.dina(w_n850_0[1]),.dinb(w_n623_0[0]),.dout(n851),.clk(gclk));
	jand g0795(.dina(n851),.dinb(n848),.dout(n852),.clk(gclk));
	jor g0796(.dina(w_n340_1[0]),.dinb(w_n276_0[0]),.dout(n853),.clk(gclk));
	jand g0797(.dina(w_n853_2[2]),.dinb(w_n368_2[0]),.dout(n854),.clk(gclk));
	jand g0798(.dina(w_n854_0[2]),.dinb(w_n532_1[2]),.dout(n855),.clk(gclk));
	jand g0799(.dina(w_n283_1[1]),.dinb(w_n109_0[2]),.dout(n856),.clk(gclk));
	jnot g0800(.din(w_n856_0[1]),.dout(n857),.clk(gclk));
	jand g0801(.dina(n857),.dinb(w_n855_0[1]),.dout(n858),.clk(gclk));
	jand g0802(.dina(w_n858_0[1]),.dinb(w_n852_0[1]),.dout(n859),.clk(gclk));
	jand g0803(.dina(n859),.dinb(n845),.dout(n860),.clk(gclk));
	jor g0804(.dina(w_n748_1[0]),.dinb(w_n641_0[0]),.dout(n861),.clk(gclk));
	jor g0805(.dina(w_n606_0[0]),.dinb(w_n213_0[2]),.dout(n862),.clk(gclk));
	jor g0806(.dina(n862),.dinb(n861),.dout(n863),.clk(gclk));
	jnot g0807(.din(w_n863_0[1]),.dout(n864),.clk(gclk));
	jand g0808(.dina(w_n645_2[0]),.dinb(w_n768_2[1]),.dout(n865),.clk(gclk));
	jor g0809(.dina(w_n554_0[0]),.dinb(w_n406_0[2]),.dout(n866),.clk(gclk));
	jnot g0810(.din(w_n866_0[1]),.dout(n867),.clk(gclk));
	jnot g0811(.din(w_n164_0[0]),.dout(n868),.clk(gclk));
	jand g0812(.dina(w_n535_1[0]),.dinb(w_n868_1[1]),.dout(n869),.clk(gclk));
	jand g0813(.dina(w_n869_0[2]),.dinb(n867),.dout(n870),.clk(gclk));
	jand g0814(.dina(n870),.dinb(w_n865_0[1]),.dout(n871),.clk(gclk));
	jand g0815(.dina(n871),.dinb(n864),.dout(n872),.clk(gclk));
	jand g0816(.dina(w_n463_2[1]),.dinb(w_n303_3[1]),.dout(n873),.clk(gclk));
	jand g0817(.dina(w_n665_2[1]),.dinb(w_n426_2[2]),.dout(n874),.clk(gclk));
	jand g0818(.dina(n874),.dinb(n873),.dout(n875),.clk(gclk));
	jand g0819(.dina(n875),.dinb(w_n568_0[1]),.dout(n876),.clk(gclk));
	jand g0820(.dina(w_n390_0[2]),.dinb(w_n383_2[1]),.dout(n877),.clk(gclk));
	jnot g0821(.din(w_n581_0[0]),.dout(n878),.clk(gclk));
	jand g0822(.dina(w_n624_2[1]),.dinb(w_n878_1[1]),.dout(n879),.clk(gclk));
	jand g0823(.dina(n879),.dinb(w_n343_1[2]),.dout(n880),.clk(gclk));
	jand g0824(.dina(w_n880_0[1]),.dinb(w_n877_0[1]),.dout(n881),.clk(gclk));
	jnot g0825(.din(w_n518_0[0]),.dout(n882),.clk(gclk));
	jand g0826(.dina(w_n592_3[0]),.dinb(w_n882_2[1]),.dout(n883),.clk(gclk));
	jand g0827(.dina(w_n883_0[1]),.dinb(w_n679_1[2]),.dout(n884),.clk(gclk));
	jand g0828(.dina(n884),.dinb(w_n773_0[0]),.dout(n885),.clk(gclk));
	jand g0829(.dina(w_n885_0[1]),.dinb(w_n881_1[1]),.dout(n886),.clk(gclk));
	jand g0830(.dina(n886),.dinb(w_n876_0[1]),.dout(n887),.clk(gclk));
	jand g0831(.dina(n887),.dinb(n872),.dout(n888),.clk(gclk));
	jand g0832(.dina(n888),.dinb(w_n860_0[1]),.dout(n889),.clk(gclk));
	jand g0833(.dina(n889),.dinb(w_n834_0[1]),.dout(n890),.clk(gclk));
	jand g0834(.dina(w_n763_2[0]),.dinb(w_n383_2[0]),.dout(n891),.clk(gclk));
	jand g0835(.dina(n891),.dinb(w_n158_0[2]),.dout(n892),.clk(gclk));
	jand g0836(.dina(w_n341_1[1]),.dinb(w_n283_1[0]),.dout(n893),.clk(gclk));
	jor g0837(.dina(w_n893_0[1]),.dinb(w_n269_0[0]),.dout(n894),.clk(gclk));
	jnot g0838(.din(w_n894_0[1]),.dout(n895),.clk(gclk));
	jand g0839(.dina(w_n895_0[1]),.dinb(w_n324_1[0]),.dout(n896),.clk(gclk));
	jnot g0840(.din(w_n160_0[0]),.dout(n897),.clk(gclk));
	jand g0841(.dina(w_n229_1[2]),.dinb(w_n897_0[2]),.dout(n898),.clk(gclk));
	jand g0842(.dina(w_n898_0[1]),.dinb(w_n771_2[0]),.dout(n899),.clk(gclk));
	jand g0843(.dina(n899),.dinb(n896),.dout(n900),.clk(gclk));
	jand g0844(.dina(n900),.dinb(n892),.dout(n901),.clk(gclk));
	jand g0845(.dina(n901),.dinb(w_n648_0[0]),.dout(n902),.clk(gclk));
	jand g0846(.dina(w_n561_1[1]),.dinb(w_n343_1[1]),.dout(n903),.clk(gclk));
	jand g0847(.dina(n903),.dinb(w_n902_0[1]),.dout(n904),.clk(gclk));
	jand g0848(.dina(w_n479_1[1]),.dinb(w_n397_1[0]),.dout(n905),.clk(gclk));
	jand g0849(.dina(w_n579_1[2]),.dinb(w_n370_1[2]),.dout(n906),.clk(gclk));
	jand g0850(.dina(w_n216_3[1]),.dinb(w_n138_3[1]),.dout(n907),.clk(gclk));
	jand g0851(.dina(n907),.dinb(w_n906_0[1]),.dout(n908),.clk(gclk));
	jand g0852(.dina(n908),.dinb(w_n905_0[1]),.dout(n909),.clk(gclk));
	jand g0853(.dina(w_n662_1[2]),.dinb(w_n612_3[0]),.dout(n910),.clk(gclk));
	jand g0854(.dina(w_n730_1[0]),.dinb(w_n868_1[0]),.dout(n911),.clk(gclk));
	jand g0855(.dina(n911),.dinb(n910),.dout(n912),.clk(gclk));
	jand g0856(.dina(w_n849_2[0]),.dinb(w_n254_2[2]),.dout(n913),.clk(gclk));
	jand g0857(.dina(n913),.dinb(w_n426_2[1]),.dout(n914),.clk(gclk));
	jand g0858(.dina(w_n914_0[1]),.dinb(w_n912_0[1]),.dout(n915),.clk(gclk));
	jand g0859(.dina(w_n734_1[1]),.dinb(w_n251_2[1]),.dout(n916),.clk(gclk));
	jand g0860(.dina(n916),.dinb(w_n463_2[0]),.dout(n917),.clk(gclk));
	jnot g0861(.din(w_n551_0[0]),.dout(n918),.clk(gclk));
	jand g0862(.dina(w_n614_2[1]),.dinb(w_n918_2[1]),.dout(n919),.clk(gclk));
	jand g0863(.dina(n919),.dinb(w_n130_1[2]),.dout(n920),.clk(gclk));
	jand g0864(.dina(w_n920_0[1]),.dinb(w_n917_0[1]),.dout(n921),.clk(gclk));
	jand g0865(.dina(n921),.dinb(n915),.dout(n922),.clk(gclk));
	jand g0866(.dina(n922),.dinb(n909),.dout(n923),.clk(gclk));
	jand g0867(.dina(w_n437_1[1]),.dinb(w_n421_3[0]),.dout(n924),.clk(gclk));
	jnot g0868(.din(w_n588_1[0]),.dout(n925),.clk(gclk));
	jand g0869(.dina(w_n925_1[1]),.dinb(w_n461_1[2]),.dout(n926),.clk(gclk));
	jand g0870(.dina(n926),.dinb(w_n924_1[2]),.dout(n927),.clk(gclk));
	jnot g0871(.din(w_n732_3[0]),.dout(n928),.clk(gclk));
	jor g0872(.dina(n928),.dinb(w_n534_0[0]),.dout(n929),.clk(gclk));
	jnot g0873(.din(w_n929_0[1]),.dout(n930),.clk(gclk));
	jand g0874(.dina(w_n930_1[1]),.dinb(w_n821_1[0]),.dout(n931),.clk(gclk));
	jand g0875(.dina(n931),.dinb(n927),.dout(n932),.clk(gclk));
	jand g0876(.dina(w_n932_0[1]),.dinb(w_n366_0[0]),.dout(n933),.clk(gclk));
	jand g0877(.dina(w_n632_1[2]),.dinb(w_n243_3[2]),.dout(n934),.clk(gclk));
	jor g0878(.dina(w_n409_0[0]),.dinb(w_n146_1[1]),.dout(n935),.clk(gclk));
	jand g0879(.dina(w_n935_3[1]),.dinb(w_n256_1[1]),.dout(n936),.clk(gclk));
	jand g0880(.dina(w_n936_0[2]),.dinb(w_n934_0[2]),.dout(n937),.clk(gclk));
	jand g0881(.dina(w_n225_1[2]),.dinb(w_n147_3[1]),.dout(n938),.clk(gclk));
	jand g0882(.dina(w_n938_0[2]),.dinb(w_n883_0[0]),.dout(n939),.clk(gclk));
	jand g0883(.dina(n939),.dinb(n937),.dout(n940),.clk(gclk));
	jand g0884(.dina(w_n710_3[0]),.dinb(w_n445_2[1]),.dout(n941),.clk(gclk));
	jand g0885(.dina(n941),.dinb(w_n625_0[0]),.dout(n942),.clk(gclk));
	jand g0886(.dina(w_n501_2[0]),.dinb(w_n387_1[1]),.dout(n943),.clk(gclk));
	jand g0887(.dina(w_n781_2[0]),.dinb(w_n379_1[0]),.dout(n944),.clk(gclk));
	jand g0888(.dina(n944),.dinb(w_n943_0[1]),.dout(n945),.clk(gclk));
	jand g0889(.dina(n945),.dinb(w_n942_0[2]),.dout(n946),.clk(gclk));
	jand g0890(.dina(n946),.dinb(n940),.dout(n947),.clk(gclk));
	jand g0891(.dina(n947),.dinb(w_n933_0[1]),.dout(n948),.clk(gclk));
	jand g0892(.dina(n948),.dinb(w_n923_0[1]),.dout(n949),.clk(gclk));
	jand g0893(.dina(n949),.dinb(w_n904_0[1]),.dout(n950),.clk(gclk));
	jxor g0894(.dina(w_n950_0[1]),.dinb(w_n486_1[0]),.dout(n951),.clk(gclk));
	jand g0895(.dina(w_n951_1[2]),.dinb(w_n890_1[2]),.dout(n952),.clk(gclk));
	jand g0896(.dina(w_n952_4[1]),.dinb(w_n820_5[2]),.dout(n953),.clk(gclk));
	jnot g0897(.din(w_n820_5[1]),.dout(n954),.clk(gclk));
	jnot g0898(.din(w_n890_1[1]),.dout(n955),.clk(gclk));
	jand g0899(.dina(w_n951_1[1]),.dinb(w_n955_0[2]),.dout(n956),.clk(gclk));
	jand g0900(.dina(w_n956_4[1]),.dinb(w_n954_24[1]),.dout(n957),.clk(gclk));
	jor g0901(.dina(n957),.dinb(n953),.dout(n958),.clk(gclk));
	jand g0902(.dina(w_n88_0[0]),.dinb(w_n49_2[1]),.dout(n959),.clk(gclk));
	jxor g0903(.dina(w_n959_0[1]),.dinb(w_a13_0[0]),.dout(n960),.clk(gclk));
	jnot g0904(.din(w_n960_5[2]),.dout(n961),.clk(gclk));
	jnot g0905(.din(w_n951_1[0]),.dout(n962),.clk(gclk));
	jor g0906(.dina(w_n950_0[0]),.dinb(w_n486_0[2]),.dout(n963),.clk(gclk));
	jand g0907(.dina(n963),.dinb(w_n955_0[1]),.dout(n964),.clk(gclk));
	jnot g0908(.din(w_n964_1[1]),.dout(n965),.clk(gclk));
	jand g0909(.dina(w_n965_0[1]),.dinb(w_n962_0[1]),.dout(n966),.clk(gclk));
	jand g0910(.dina(w_n966_4[1]),.dinb(w_n961_5[1]),.dout(n967),.clk(gclk));
	jnot g0911(.din(w_n486_0[1]),.dout(n968),.clk(gclk));
	jand g0912(.dina(w_n890_1[0]),.dinb(w_n968_0[1]),.dout(n969),.clk(gclk));
	jor g0913(.dina(n969),.dinb(w_n951_0[2]),.dout(n970),.clk(gclk));
	jnot g0914(.din(w_n970_0[2]),.dout(n971),.clk(gclk));
	jand g0915(.dina(w_n971_4[1]),.dinb(w_n960_5[1]),.dout(n972),.clk(gclk));
	jor g0916(.dina(n972),.dinb(n967),.dout(n973),.clk(gclk));
	jor g0917(.dina(n973),.dinb(n958),.dout(n974),.clk(gclk));
	jnot g0918(.din(n974),.dout(n975),.clk(gclk));
	jand g0919(.dina(w_a22_2[2]),.dinb(w_a12_0[2]),.dout(n976),.clk(gclk));
	jand g0920(.dina(w_n87_0[0]),.dinb(w_a12_0[1]),.dout(n977),.clk(gclk));
	jnot g0921(.din(n977),.dout(n978),.clk(gclk));
	jand g0922(.dina(n978),.dinb(w_n959_0[0]),.dout(n979),.clk(gclk));
	jor g0923(.dina(n979),.dinb(n976),.dout(n980),.clk(gclk));
	jnot g0924(.din(w_n980_6[1]),.dout(n981),.clk(gclk));
	jand g0925(.dina(w_n379_0[2]),.dinb(w_n254_2[1]),.dout(n982),.clk(gclk));
	jand g0926(.dina(w_n853_2[1]),.dinb(w_n232_1[2]),.dout(n983),.clk(gclk));
	jand g0927(.dina(n983),.dinb(n982),.dout(n984),.clk(gclk));
	jand g0928(.dina(w_n354_1[2]),.dinb(w_n227_0[2]),.dout(n985),.clk(gclk));
	jor g0929(.dina(w_n985_0[1]),.dinb(w_n369_0[0]),.dout(n986),.clk(gclk));
	jnot g0930(.din(w_n986_0[1]),.dout(n987),.clk(gclk));
	jand g0931(.dina(w_n768_2[0]),.dinb(w_n358_1[2]),.dout(n988),.clk(gclk));
	jand g0932(.dina(w_n988_0[1]),.dinb(w_n301_1[2]),.dout(n989),.clk(gclk));
	jand g0933(.dina(n989),.dinb(w_n987_1[2]),.dout(n990),.clk(gclk));
	jand g0934(.dina(n990),.dinb(n984),.dout(n991),.clk(gclk));
	jand g0935(.dina(w_n749_1[0]),.dinb(w_n709_1[0]),.dout(n992),.clk(gclk));
	jor g0936(.dina(w_n340_0[2]),.dinb(w_n380_0[1]),.dout(n993),.clk(gclk));
	jand g0937(.dina(w_n993_1[2]),.dinb(w_n421_2[2]),.dout(n994),.clk(gclk));
	jand g0938(.dina(w_n506_1[1]),.dinb(w_n381_1[2]),.dout(n995),.clk(gclk));
	jand g0939(.dina(n995),.dinb(w_n994_0[1]),.dout(n996),.clk(gclk));
	jand g0940(.dina(n996),.dinb(w_n992_1[2]),.dout(n997),.clk(gclk));
	jand g0941(.dina(w_n772_2[1]),.dinb(w_n249_1[1]),.dout(n998),.clk(gclk));
	jand g0942(.dina(n998),.dinb(w_n303_3[0]),.dout(n999),.clk(gclk));
	jand g0943(.dina(w_n291_2[0]),.dinb(w_n267_1[0]),.dout(n1000),.clk(gclk));
	jand g0944(.dina(w_n662_1[1]),.dinb(w_n467_0[2]),.dout(n1001),.clk(gclk));
	jand g0945(.dina(n1001),.dinb(w_n1000_0[1]),.dout(n1002),.clk(gclk));
	jand g0946(.dina(w_n1002_0[1]),.dinb(w_n999_0[2]),.dout(n1003),.clk(gclk));
	jand g0947(.dina(n1003),.dinb(n997),.dout(n1004),.clk(gclk));
	jand g0948(.dina(n1004),.dinb(w_n991_0[1]),.dout(n1005),.clk(gclk));
	jand g0949(.dina(n1005),.dinb(w_n904_0[0]),.dout(n1006),.clk(gclk));
	jand g0950(.dina(w_n473_1[1]),.dinb(w_n825_1[1]),.dout(n1007),.clk(gclk));
	jand g0951(.dina(w_n285_2[0]),.dinb(w_n256_1[0]),.dout(n1008),.clk(gclk));
	jand g0952(.dina(n1008),.dinb(n1007),.dout(n1009),.clk(gclk));
	jand g0953(.dina(n1009),.dinb(w_n626_1[0]),.dout(n1010),.clk(gclk));
	jand g0954(.dina(n1010),.dinb(w_n920_0[0]),.dout(n1011),.clk(gclk));
	jand g0955(.dina(w_n732_2[2]),.dinb(w_n138_3[0]),.dout(n1012),.clk(gclk));
	jand g0956(.dina(n1012),.dinb(w_n1011_0[1]),.dout(n1013),.clk(gclk));
	jand g0957(.dina(w_n632_1[1]),.dinb(w_n882_2[0]),.dout(n1014),.clk(gclk));
	jand g0958(.dina(w_n441_1[0]),.dinb(w_n437_1[0]),.dout(n1015),.clk(gclk));
	jand g0959(.dina(n1015),.dinb(n1014),.dout(n1016),.clk(gclk));
	jor g0960(.dina(w_n309_0[0]),.dinb(w_n260_0[0]),.dout(n1017),.clk(gclk));
	jnot g0961(.din(w_n1017_0[1]),.dout(n1018),.clk(gclk));
	jand g0962(.dina(w_n1018_1[1]),.dinb(w_n543_1[0]),.dout(n1019),.clk(gclk));
	jand g0963(.dina(n1019),.dinb(n1016),.dout(n1020),.clk(gclk));
	jand g0964(.dina(w_n765_1[1]),.dinb(w_n665_2[0]),.dout(n1021),.clk(gclk));
	jand g0965(.dina(w_n532_1[1]),.dinb(w_n420_1[0]),.dout(n1022),.clk(gclk));
	jand g0966(.dina(w_n1022_0[2]),.dinb(w_n499_1[0]),.dout(n1023),.clk(gclk));
	jand g0967(.dina(n1023),.dinb(w_n1021_0[1]),.dout(n1024),.clk(gclk));
	jand g0968(.dina(w_n724_2[1]),.dinb(w_n427_2[2]),.dout(n1025),.clk(gclk));
	jand g0969(.dina(w_n1025_0[2]),.dinb(w_n849_1[2]),.dout(n1026),.clk(gclk));
	jand g0970(.dina(w_n710_2[2]),.dinb(w_n399_0[0]),.dout(n1027),.clk(gclk));
	jand g0971(.dina(w_n1027_0[2]),.dinb(w_n1026_0[1]),.dout(n1028),.clk(gclk));
	jand g0972(.dina(n1028),.dinb(n1024),.dout(n1029),.clk(gclk));
	jand g0973(.dina(n1029),.dinb(w_n1020_0[1]),.dout(n1030),.clk(gclk));
	jand g0974(.dina(n1030),.dinb(w_n1013_0[1]),.dout(n1031),.clk(gclk));
	jand g0975(.dina(n1031),.dinb(w_n1006_0[1]),.dout(n1032),.clk(gclk));
	jxor g0976(.dina(w_n1032_0[1]),.dinb(w_n890_0[2]),.dout(n1033),.clk(gclk));
	jand g0977(.dina(w_n1033_1[2]),.dinb(w_n762_1[0]),.dout(n1034),.clk(gclk));
	jnot g0978(.din(w_n1034_3[2]),.dout(n1035),.clk(gclk));
	jand g0979(.dina(w_n1035_0[2]),.dinb(w_n981_4[2]),.dout(n1036),.clk(gclk));
	jand g0980(.dina(w_n1033_1[1]),.dinb(w_n790_0[1]),.dout(n1037),.clk(gclk));
	jnot g0981(.din(w_n1037_3[2]),.dout(n1038),.clk(gclk));
	jand g0982(.dina(w_n1038_0[2]),.dinb(w_n980_6[0]),.dout(n1039),.clk(gclk));
	jor g0983(.dina(n1039),.dinb(n1036),.dout(n1040),.clk(gclk));
	jand g0984(.dina(w_n955_0[0]),.dinb(w_n762_0[2]),.dout(n1041),.clk(gclk));
	jor g0985(.dina(n1041),.dinb(w_n1033_1[0]),.dout(n1042),.clk(gclk));
	jnot g0986(.din(w_n1042_0[2]),.dout(n1043),.clk(gclk));
	jand g0987(.dina(w_n1043_4[1]),.dinb(w_n803_8[1]),.dout(n1044),.clk(gclk));
	jnot g0988(.din(w_n1033_0[2]),.dout(n1045),.clk(gclk));
	jor g0989(.dina(w_n1032_0[0]),.dinb(w_n890_0[1]),.dout(n1046),.clk(gclk));
	jand g0990(.dina(n1046),.dinb(w_n790_0[0]),.dout(n1047),.clk(gclk));
	jnot g0991(.din(w_n1047_1[1]),.dout(n1048),.clk(gclk));
	jand g0992(.dina(n1048),.dinb(w_n1045_0[1]),.dout(n1049),.clk(gclk));
	jand g0993(.dina(w_n1049_4[1]),.dinb(w_n808_13[1]),.dout(n1050),.clk(gclk));
	jor g0994(.dina(n1050),.dinb(n1044),.dout(n1051),.clk(gclk));
	jnot g0995(.din(n1051),.dout(n1052),.clk(gclk));
	jand g0996(.dina(n1052),.dinb(n1040),.dout(n1053),.clk(gclk));
	jand g0997(.dina(w_n1053_0[1]),.dinb(w_n975_0[1]),.dout(n1054),.clk(gclk));
	jxor g0998(.dina(w_n1053_0[0]),.dinb(w_n975_0[0]),.dout(n1055),.clk(gclk));
	jxor g0999(.dina(w_n695_0[0]),.dinb(w_a9_0[0]),.dout(n1057),.clk(gclk));
	jand g1000(.dina(w_n1057_5[1]),.dinb(w_n804_3[2]),.dout(n1058),.clk(gclk));
	jnot g1001(.din(w_n1057_5[0]),.dout(n1059),.clk(gclk));
	jand g1002(.dina(w_n1059_5[2]),.dinb(w_n799_3[1]),.dout(n1060),.clk(gclk));
	jor g1003(.dina(n1060),.dinb(n1058),.dout(n1061),.clk(gclk));
	jand g1004(.dina(w_n789_4[1]),.dinb(w_n794_4[1]),.dout(n1063),.clk(gclk));
	jor g1005(.dina(n1063),.dinb(n1061),.dout(n1065),.clk(gclk));
	jnot g1006(.din(n1065),.dout(n1066),.clk(gclk));
	jand g1007(.dina(w_n1066_0[1]),.dinb(w_n1055_0[1]),.dout(n1067),.clk(gclk));
	jor g1008(.dina(n1067),.dinb(n1054),.dout(n1068),.clk(gclk));
	jxor g1009(.dina(w_n813_0[0]),.dinb(w_n702_0[0]),.dout(n1069),.clk(gclk));
	jand g1010(.dina(w_n1069_0[1]),.dinb(w_n1068_0[1]),.dout(n1070),.clk(gclk));
	jor g1011(.dina(n1070),.dinb(n814),.dout(n1071),.clk(gclk));
	jand g1012(.dina(w_n1057_4[2]),.dinb(w_n335_6[0]),.dout(n1072),.clk(gclk));
	jnot g1013(.din(w_n1072_0[1]),.dout(n1073),.clk(gclk));
	jxor g1014(.dina(w_n1073_0[2]),.dinb(w_n964_1[0]),.dout(n1074),.clk(gclk));
	jand g1015(.dina(w_n708_5[2]),.dinb(w_n335_5[2]),.dout(n1075),.clk(gclk));
	jxor g1016(.dina(w_n1075_0[1]),.dinb(w_n1074_0[1]),.dout(n1076),.clk(gclk));
	jand g1017(.dina(w_n1076_0[1]),.dinb(w_n1071_0[1]),.dout(n1077),.clk(gclk));
	jxor g1018(.dina(w_n1076_0[0]),.dinb(w_n1071_0[0]),.dout(n1078),.clk(gclk));
	jand g1019(.dina(w_n962_0[0]),.dinb(w_n954_24[0]),.dout(n1079),.clk(gclk));
	jor g1020(.dina(n1079),.dinb(w_n964_0[2]),.dout(n1080),.clk(gclk));
	jand g1021(.dina(w_n971_4[0]),.dinb(w_n954_23[2]),.dout(n1081),.clk(gclk));
	jnot g1022(.din(n1081),.dout(n1082),.clk(gclk));
	jand g1023(.dina(n1082),.dinb(n1080),.dout(n1083),.clk(gclk));
	jand g1024(.dina(w_n1083_0[1]),.dinb(w_n1073_0[1]),.dout(n1084),.clk(gclk));
	jxor g1025(.dina(w_n1083_0[0]),.dinb(w_n1073_0[0]),.dout(n1085),.clk(gclk));
	jand g1026(.dina(w_n1037_3[1]),.dinb(w_n960_5[0]),.dout(n1086),.clk(gclk));
	jand g1027(.dina(w_n1034_3[1]),.dinb(w_n961_5[0]),.dout(n1087),.clk(gclk));
	jor g1028(.dina(n1087),.dinb(n1086),.dout(n1088),.clk(gclk));
	jand g1029(.dina(w_n1043_4[0]),.dinb(w_n980_5[2]),.dout(n1089),.clk(gclk));
	jand g1030(.dina(w_n1049_4[0]),.dinb(w_n981_4[1]),.dout(n1090),.clk(gclk));
	jor g1031(.dina(n1090),.dinb(n1089),.dout(n1091),.clk(gclk));
	jor g1032(.dina(n1091),.dinb(n1088),.dout(n1092),.clk(gclk));
	jnot g1033(.din(n1092),.dout(n1093),.clk(gclk));
	jand g1034(.dina(w_n1093_0[1]),.dinb(w_n1085_0[1]),.dout(n1094),.clk(gclk));
	jor g1035(.dina(n1094),.dinb(n1084),.dout(n1095),.clk(gclk));
	jand g1036(.dina(w_n803_8[0]),.dinb(w_n804_3[1]),.dout(n1096),.clk(gclk));
	jand g1037(.dina(w_n808_13[0]),.dinb(w_n799_3[0]),.dout(n1097),.clk(gclk));
	jor g1038(.dina(n1097),.dinb(n1096),.dout(n1098),.clk(gclk));
	jand g1039(.dina(w_n981_4[0]),.dinb(w_n789_4[0]),.dout(n1100),.clk(gclk));
	jor g1040(.dina(n1100),.dinb(n1098),.dout(n1102),.clk(gclk));
	jand g1041(.dina(w_n1034_3[0]),.dinb(w_n820_5[0]),.dout(n1103),.clk(gclk));
	jand g1042(.dina(w_n1037_3[0]),.dinb(w_n954_23[1]),.dout(n1104),.clk(gclk));
	jor g1043(.dina(n1104),.dinb(n1103),.dout(n1105),.clk(gclk));
	jand g1044(.dina(w_n1049_3[2]),.dinb(w_n961_4[2]),.dout(n1106),.clk(gclk));
	jand g1045(.dina(w_n1043_3[2]),.dinb(w_n960_4[2]),.dout(n1107),.clk(gclk));
	jor g1046(.dina(n1107),.dinb(n1106),.dout(n1108),.clk(gclk));
	jor g1047(.dina(n1108),.dinb(n1105),.dout(n1109),.clk(gclk));
	jxor g1048(.dina(w_n1109_0[1]),.dinb(w_n1102_0[1]),.dout(n1110),.clk(gclk));
	jxor g1049(.dina(w_n1110_0[1]),.dinb(w_n1095_0[1]),.dout(n1111),.clk(gclk));
	jand g1050(.dina(w_n1111_0[1]),.dinb(w_n1078_0[1]),.dout(n1112),.clk(gclk));
	jor g1051(.dina(n1112),.dinb(n1077),.dout(n1113),.clk(gclk));
	jand g1052(.dina(w_n803_7[2]),.dinb(w_n335_5[1]),.dout(n1114),.clk(gclk));
	jnot g1053(.din(w_n1114_0[1]),.dout(n1115),.clk(gclk));
	jand g1054(.dina(w_n1045_0[0]),.dinb(w_n954_23[0]),.dout(n1116),.clk(gclk));
	jor g1055(.dina(n1116),.dinb(w_n1047_1[0]),.dout(n1117),.clk(gclk));
	jand g1056(.dina(w_n1043_3[1]),.dinb(w_n954_22[2]),.dout(n1118),.clk(gclk));
	jnot g1057(.din(n1118),.dout(n1119),.clk(gclk));
	jand g1058(.dina(n1119),.dinb(n1117),.dout(n1120),.clk(gclk));
	jxor g1059(.dina(w_n1120_0[1]),.dinb(w_n1115_0[2]),.dout(n1121),.clk(gclk));
	jand g1060(.dina(w_n981_3[2]),.dinb(w_n799_2[2]),.dout(n1122),.clk(gclk));
	jand g1061(.dina(w_n980_5[1]),.dinb(w_n804_3[0]),.dout(n1123),.clk(gclk));
	jor g1062(.dina(n1123),.dinb(n1122),.dout(n1124),.clk(gclk));
	jand g1063(.dina(w_n961_4[1]),.dinb(w_n789_3[2]),.dout(n1125),.clk(gclk));
	jor g1064(.dina(n1125),.dinb(n1124),.dout(n1128),.clk(gclk));
	jnot g1065(.din(n1128),.dout(n1129),.clk(gclk));
	jxor g1066(.dina(w_n1129_0[1]),.dinb(w_n1121_0[1]),.dout(n1130),.clk(gclk));
	jand g1067(.dina(w_n1072_0[0]),.dinb(w_n965_0[0]),.dout(n1131),.clk(gclk));
	jand g1068(.dina(w_n1075_0[0]),.dinb(w_n1074_0[0]),.dout(n1132),.clk(gclk));
	jor g1069(.dina(n1132),.dinb(n1131),.dout(n1133),.clk(gclk));
	jnot g1070(.din(w_n1102_0[0]),.dout(n1134),.clk(gclk));
	jnot g1071(.din(w_n1109_0[0]),.dout(n1135),.clk(gclk));
	jand g1072(.dina(n1135),.dinb(n1134),.dout(n1136),.clk(gclk));
	jand g1073(.dina(w_n1110_0[0]),.dinb(w_n1095_0[0]),.dout(n1137),.clk(gclk));
	jor g1074(.dina(n1137),.dinb(n1136),.dout(n1138),.clk(gclk));
	jxor g1075(.dina(w_n1138_0[1]),.dinb(w_n1133_0[1]),.dout(n1139),.clk(gclk));
	jxor g1076(.dina(w_n1139_0[1]),.dinb(w_n1130_0[1]),.dout(n1140),.clk(gclk));
	jand g1077(.dina(w_n1140_0[1]),.dinb(w_n1113_0[1]),.dout(n1141),.clk(gclk));
	jand g1078(.dina(w_n792_0[1]),.dinb(w_n699_13[1]),.dout(n1142),.clk(gclk));
	jnot g1079(.din(w_n699_13[0]),.dout(n1143),.clk(gclk));
	jand g1080(.dina(w_n800_0[1]),.dinb(w_n1143_9[1]),.dout(n1144),.clk(gclk));
	jor g1081(.dina(n1144),.dinb(n1142),.dout(n1145),.clk(gclk));
	jand g1082(.dina(w_n1059_5[1]),.dinb(w_n789_3[1]),.dout(n1147),.clk(gclk));
	jnot g1083(.din(n1147),.dout(n1149),.clk(gclk));
	jand g1084(.dina(n1149),.dinb(n1145),.dout(n1150),.clk(gclk));
	jand g1085(.dina(w_n1042_0[1]),.dinb(w_n708_5[1]),.dout(n1151),.clk(gclk));
	jnot g1086(.din(w_n1049_3[1]),.dout(n1152),.clk(gclk));
	jand g1087(.dina(w_n1152_0[1]),.dinb(w_n794_4[0]),.dout(n1153),.clk(gclk));
	jor g1088(.dina(n1153),.dinb(n1151),.dout(n1154),.clk(gclk));
	jand g1089(.dina(w_n1037_2[2]),.dinb(w_n803_7[1]),.dout(n1155),.clk(gclk));
	jand g1090(.dina(w_n1034_2[2]),.dinb(w_n808_12[2]),.dout(n1156),.clk(gclk));
	jor g1091(.dina(n1156),.dinb(n1155),.dout(n1157),.clk(gclk));
	jnot g1092(.din(n1157),.dout(n1158),.clk(gclk));
	jand g1093(.dina(n1158),.dinb(n1154),.dout(n1159),.clk(gclk));
	jand g1094(.dina(w_n1159_0[1]),.dinb(w_n1150_0[1]),.dout(n1160),.clk(gclk));
	jnot g1095(.din(n1160),.dout(n1161),.clk(gclk));
	jxor g1096(.dina(w_n1159_0[0]),.dinb(w_n1150_0[0]),.dout(n1162),.clk(gclk));
	jnot g1097(.din(n1162),.dout(n1163),.clk(gclk));
	jnot g1098(.din(w_n519_0[0]),.dout(n1164),.clk(gclk));
	jand g1099(.dina(n1164),.dinb(w_n516_0[0]),.dout(n1165),.clk(gclk));
	jand g1100(.dina(w_n525_0[0]),.dinb(n1165),.dout(n1166),.clk(gclk));
	jand g1101(.dina(n1166),.dinb(w_n513_0[1]),.dout(n1167),.clk(gclk));
	jand g1102(.dina(n1167),.dinb(w_n509_0[1]),.dout(n1168),.clk(gclk));
	jand g1103(.dina(n1168),.dinb(w_n497_1[0]),.dout(n1169),.clk(gclk));
	jnot g1104(.din(w_n545_0[0]),.dout(n1170),.clk(gclk));
	jand g1105(.dina(w_n1170_0[2]),.dinb(w_n543_0[2]),.dout(n1171),.clk(gclk));
	jand g1106(.dina(n1171),.dinb(w_n541_0[0]),.dout(n1172),.clk(gclk));
	jnot g1107(.din(w_n557_0[0]),.dout(n1173),.clk(gclk));
	jand g1108(.dina(n1173),.dinb(n1172),.dout(n1174),.clk(gclk));
	jand g1109(.dina(n1174),.dinb(w_n538_0[1]),.dout(n1175),.clk(gclk));
	jnot g1110(.din(w_n571_0[1]),.dout(n1176),.clk(gclk));
	jand g1111(.dina(w_n1176_0[1]),.dinb(w_n568_0[0]),.dout(n1177),.clk(gclk));
	jand g1112(.dina(n1177),.dinb(w_n565_1[0]),.dout(n1178),.clk(gclk));
	jnot g1113(.din(w_n584_0[0]),.dout(n1179),.clk(gclk));
	jnot g1114(.din(w_n590_0[0]),.dout(n1180),.clk(gclk));
	jand g1115(.dina(w_n598_0[0]),.dinb(n1180),.dout(n1181),.clk(gclk));
	jand g1116(.dina(n1181),.dinb(w_n1179_0[1]),.dout(n1182),.clk(gclk));
	jand g1117(.dina(n1182),.dinb(n1178),.dout(n1183),.clk(gclk));
	jand g1118(.dina(n1183),.dinb(w_n1175_0[1]),.dout(n1184),.clk(gclk));
	jand g1119(.dina(n1184),.dinb(w_n1169_0[1]),.dout(n1185),.clk(gclk));
	jand g1120(.dina(w_n624_2[0]),.dinb(w_n506_1[0]),.dout(n1186),.clk(gclk));
	jand g1121(.dina(n1186),.dinb(w_n837_2[0]),.dout(n1187),.clk(gclk));
	jand g1122(.dina(w_n402_2[0]),.dinb(w_n351_1[1]),.dout(n1188),.clk(gclk));
	jand g1123(.dina(w_n1188_0[1]),.dinb(w_n594_2[1]),.dout(n1189),.clk(gclk));
	jor g1124(.dina(w_n748_0[2]),.dinb(w_n631_0[1]),.dout(n1190),.clk(gclk));
	jnot g1125(.din(w_n1190_0[1]),.dout(n1191),.clk(gclk));
	jand g1126(.dina(w_n427_2[1]),.dinb(w_n348_1[1]),.dout(n1192),.clk(gclk));
	jand g1127(.dina(w_n1192_0[1]),.dinb(n1191),.dout(n1193),.clk(gclk));
	jand g1128(.dina(w_n1193_0[1]),.dinb(w_n1189_1[1]),.dout(n1194),.clk(gclk));
	jand g1129(.dina(n1194),.dinb(w_n1187_0[2]),.dout(n1195),.clk(gclk));
	jand g1130(.dina(w_n744_2[0]),.dinb(w_n279_1[2]),.dout(n1196),.clk(gclk));
	jand g1131(.dina(w_n882_1[2]),.dinb(w_n426_2[0]),.dout(n1197),.clk(gclk));
	jor g1132(.dina(w_n678_0[0]),.dinb(w_n400_0[0]),.dout(n1198),.clk(gclk));
	jnot g1133(.din(w_n1198_0[1]),.dout(n1199),.clk(gclk));
	jand g1134(.dina(n1199),.dinb(w_n1197_0[1]),.dout(n1200),.clk(gclk));
	jand g1135(.dina(n1200),.dinb(w_n1196_0[2]),.dout(n1201),.clk(gclk));
	jand g1136(.dina(n1201),.dinb(w_n622_1[1]),.dout(n1202),.clk(gclk));
	jand g1137(.dina(n1202),.dinb(n1195),.dout(n1203),.clk(gclk));
	jand g1138(.dina(w_n993_1[1]),.dinb(w_n612_2[2]),.dout(n1204),.clk(gclk));
	jand g1139(.dina(w_n1204_1[1]),.dinb(w_n638_0[1]),.dout(n1205),.clk(gclk));
	jand g1140(.dina(n1205),.dinb(w_n408_0[0]),.dout(n1206),.clk(gclk));
	jand g1141(.dina(w_n579_1[1]),.dinb(w_n363_1[2]),.dout(n1207),.clk(gclk));
	jand g1142(.dina(n1207),.dinb(w_n454_1[1]),.dout(n1208),.clk(gclk));
	jnot g1143(.din(w_n299_0[1]),.dout(n1209),.clk(gclk));
	jand g1144(.dina(w_n935_3[0]),.dinb(w_n1209_1[2]),.dout(n1210),.clk(gclk));
	jand g1145(.dina(w_n1210_0[1]),.dinb(w_n597_2[0]),.dout(n1211),.clk(gclk));
	jand g1146(.dina(n1211),.dinb(n1208),.dout(n1212),.clk(gclk));
	jand g1147(.dina(n1212),.dinb(n1206),.dout(n1213),.clk(gclk));
	jor g1148(.dina(w_n355_0[0]),.dinb(w_n288_0[1]),.dout(n1214),.clk(gclk));
	jor g1149(.dina(w_n750_0[0]),.dinb(w_n591_0[0]),.dout(n1215),.clk(gclk));
	jor g1150(.dina(w_n1215_0[1]),.dinb(w_n475_0[1]),.dout(n1216),.clk(gclk));
	jor g1151(.dina(n1216),.dinb(w_n1214_0[1]),.dout(n1217),.clk(gclk));
	jnot g1152(.din(w_n1217_0[2]),.dout(n1218),.clk(gclk));
	jand g1153(.dina(w_n1218_0[2]),.dinb(w_n858_0[0]),.dout(n1219),.clk(gclk));
	jand g1154(.dina(n1219),.dinb(n1213),.dout(n1220),.clk(gclk));
	jor g1155(.dina(w_n415_0[0]),.dinb(w_n224_0[1]),.dout(n1221),.clk(gclk));
	jand g1156(.dina(w_n501_1[2]),.dinb(w_n381_1[1]),.dout(n1222),.clk(gclk));
	jnot g1157(.din(n1222),.dout(n1223),.clk(gclk));
	jor g1158(.dina(n1223),.dinb(n1221),.dout(n1224),.clk(gclk));
	jnot g1159(.din(w_n1224_0[1]),.dout(n1225),.clk(gclk));
	jand g1160(.dina(w_n924_1[1]),.dinb(w_n523_0[1]),.dout(n1226),.clk(gclk));
	jor g1161(.dina(w_n364_0[0]),.dinb(w_n235_0[0]),.dout(n1227),.clk(gclk));
	jnot g1162(.din(w_n1227_0[1]),.dout(n1228),.clk(gclk));
	jand g1163(.dina(w_n1228_0[1]),.dinb(w_n850_0[0]),.dout(n1229),.clk(gclk));
	jand g1164(.dina(n1229),.dinb(n1226),.dout(n1230),.clk(gclk));
	jand g1165(.dina(n1230),.dinb(n1225),.dout(n1231),.clk(gclk));
	jand g1166(.dina(w_n354_1[1]),.dinb(w_n259_1[0]),.dout(n1232),.clk(gclk));
	jor g1167(.dina(w_n1232_0[1]),.dinb(w_n213_0[1]),.dout(n1233),.clk(gclk));
	jor g1168(.dina(n1233),.dinb(w_n552_0[0]),.dout(n1234),.clk(gclk));
	jor g1169(.dina(w_n780_0[0]),.dinb(w_n250_0[0]),.dout(n1235),.clk(gclk));
	jor g1170(.dina(w_n373_0[0]),.dinb(w_n266_0[2]),.dout(n1236),.clk(gclk));
	jor g1171(.dina(n1236),.dinb(n1235),.dout(n1237),.clk(gclk));
	jor g1172(.dina(n1237),.dinb(w_n727_0[0]),.dout(n1238),.clk(gclk));
	jor g1173(.dina(n1238),.dinb(n1234),.dout(n1239),.clk(gclk));
	jnot g1174(.din(w_n1239_0[1]),.dout(n1240),.clk(gclk));
	jand g1175(.dina(w_n1240_0[1]),.dinb(w_n1231_0[2]),.dout(n1241),.clk(gclk));
	jand g1176(.dina(n1241),.dinb(n1220),.dout(n1242),.clk(gclk));
	jand g1177(.dina(n1242),.dinb(w_n1203_0[2]),.dout(n1243),.clk(gclk));
	jand g1178(.dina(w_n1243_2[1]),.dinb(w_n1185_1[2]),.dout(n1244),.clk(gclk));
	jnot g1179(.din(n1244),.dout(n1245),.clk(gclk));
	jnot g1180(.din(w_n1187_0[1]),.dout(n1246),.clk(gclk));
	jnot g1181(.din(w_n1189_1[0]),.dout(n1247),.clk(gclk));
	jnot g1182(.din(w_n1192_0[0]),.dout(n1248),.clk(gclk));
	jor g1183(.dina(n1248),.dinb(w_n1190_0[0]),.dout(n1249),.clk(gclk));
	jor g1184(.dina(n1249),.dinb(n1247),.dout(n1250),.clk(gclk));
	jor g1185(.dina(n1250),.dinb(n1246),.dout(n1251),.clk(gclk));
	jnot g1186(.din(w_n622_1[0]),.dout(n1252),.clk(gclk));
	jnot g1187(.din(w_n1196_0[1]),.dout(n1253),.clk(gclk));
	jnot g1188(.din(w_n1197_0[0]),.dout(n1254),.clk(gclk));
	jor g1189(.dina(w_n1198_0[0]),.dinb(n1254),.dout(n1255),.clk(gclk));
	jor g1190(.dina(n1255),.dinb(n1253),.dout(n1256),.clk(gclk));
	jor g1191(.dina(n1256),.dinb(n1252),.dout(n1257),.clk(gclk));
	jor g1192(.dina(n1257),.dinb(n1251),.dout(n1258),.clk(gclk));
	jnot g1193(.din(w_n1204_1[0]),.dout(n1259),.clk(gclk));
	jor g1194(.dina(w_n1259_0[1]),.dinb(w_n637_0[0]),.dout(n1260),.clk(gclk));
	jor g1195(.dina(n1260),.dinb(w_n407_0[0]),.dout(n1261),.clk(gclk));
	jor g1196(.dina(w_n580_0[0]),.dinb(w_n362_0[0]),.dout(n1262),.clk(gclk));
	jor g1197(.dina(n1262),.dinb(w_n453_0[0]),.dout(n1263),.clk(gclk));
	jnot g1198(.din(w_n597_1[2]),.dout(n1264),.clk(gclk));
	jnot g1199(.din(w_n935_2[2]),.dout(n1265),.clk(gclk));
	jor g1200(.dina(n1265),.dinb(w_n299_0[0]),.dout(n1266),.clk(gclk));
	jor g1201(.dina(n1266),.dinb(n1264),.dout(n1267),.clk(gclk));
	jor g1202(.dina(n1267),.dinb(n1263),.dout(n1268),.clk(gclk));
	jor g1203(.dina(n1268),.dinb(n1261),.dout(n1269),.clk(gclk));
	jnot g1204(.din(w_n854_0[1]),.dout(n1270),.clk(gclk));
	jor g1205(.dina(n1270),.dinb(w_n531_0[0]),.dout(n1271),.clk(gclk));
	jor g1206(.dina(w_n856_0[0]),.dinb(n1271),.dout(n1272),.clk(gclk));
	jor g1207(.dina(w_n1217_0[1]),.dinb(n1272),.dout(n1273),.clk(gclk));
	jor g1208(.dina(n1273),.dinb(n1269),.dout(n1274),.clk(gclk));
	jnot g1209(.din(w_n924_1[0]),.dout(n1275),.clk(gclk));
	jor g1210(.dina(n1275),.dinb(w_n522_0[0]),.dout(n1276),.clk(gclk));
	jor g1211(.dina(w_n608_0[0]),.dinb(w_n577_0[0]),.dout(n1277),.clk(gclk));
	jor g1212(.dina(w_n1227_0[0]),.dinb(n1277),.dout(n1278),.clk(gclk));
	jor g1213(.dina(n1278),.dinb(n1276),.dout(n1279),.clk(gclk));
	jor g1214(.dina(n1279),.dinb(w_n1224_0[0]),.dout(n1280),.clk(gclk));
	jor g1215(.dina(w_n1239_0[0]),.dinb(n1280),.dout(n1281),.clk(gclk));
	jor g1216(.dina(n1281),.dinb(n1274),.dout(n1282),.clk(gclk));
	jor g1217(.dina(n1282),.dinb(n1258),.dout(n1283),.clk(gclk));
	jand g1218(.dina(w_n882_1[1]),.dinb(w_n479_1[0]),.dout(n1284),.clk(gclk));
	jand g1219(.dina(n1284),.dinb(w_n724_2[0]),.dout(n1285),.clk(gclk));
	jand g1220(.dina(w_n1285_0[1]),.dinb(w_n1176_0[0]),.dout(n1286),.clk(gclk));
	jand g1221(.dina(n1286),.dinb(w_n1027_0[1]),.dout(n1287),.clk(gclk));
	jor g1222(.dina(w_n560_0[0]),.dinb(w_n231_0[0]),.dout(n1288),.clk(gclk));
	jnot g1223(.din(w_n1288_0[1]),.dout(n1289),.clk(gclk));
	jand g1224(.dina(n1289),.dinb(w_n733_1[0]),.dout(n1290),.clk(gclk));
	jand g1225(.dina(w_n1204_0[2]),.dinb(w_n934_0[1]),.dout(n1291),.clk(gclk));
	jand g1226(.dina(n1291),.dinb(n1290),.dout(n1292),.clk(gclk));
	jor g1227(.dina(w_n661_0[0]),.dinb(w_n152_0[0]),.dout(n1293),.clk(gclk));
	jnot g1228(.din(w_n1293_0[1]),.dout(n1294),.clk(gclk));
	jand g1229(.dina(w_n1294_0[1]),.dinb(w_n286_1[0]),.dout(n1295),.clk(gclk));
	jand g1230(.dina(n1295),.dinb(w_n895_0[0]),.dout(n1296),.clk(gclk));
	jand g1231(.dina(n1296),.dinb(w_n1292_0[1]),.dout(n1297),.clk(gclk));
	jand g1232(.dina(n1297),.dinb(w_n1218_0[1]),.dout(n1298),.clk(gclk));
	jand g1233(.dina(n1298),.dinb(n1287),.dout(n1299),.clk(gclk));
	jor g1234(.dina(w_n406_0[1]),.dinb(w_n386_0[0]),.dout(n1300),.clk(gclk));
	jor g1235(.dina(w_n266_0[1]),.dinb(w_n224_0[0]),.dout(n1301),.clk(gclk));
	jor g1236(.dina(n1301),.dinb(n1300),.dout(n1302),.clk(gclk));
	jnot g1237(.din(w_n1302_0[1]),.dout(n1303),.clk(gclk));
	jand g1238(.dina(w_n402_1[2]),.dinb(w_n323_3[0]),.dout(n1304),.clk(gclk));
	jand g1239(.dina(n1304),.dinb(w_n511_1[0]),.dout(n1305),.clk(gclk));
	jand g1240(.dina(n1305),.dinb(w_n1018_1[0]),.dout(n1306),.clk(gclk));
	jand g1241(.dina(n1306),.dinb(n1303),.dout(n1307),.clk(gclk));
	jnot g1242(.din(w_n596_0[1]),.dout(n1308),.clk(gclk));
	jor g1243(.dina(n1308),.dinb(w_n588_0[2]),.dout(n1309),.clk(gclk));
	jnot g1244(.din(w_n1309_0[1]),.dout(n1310),.clk(gclk));
	jand g1245(.dina(w_n935_2[1]),.dinb(w_n515_1[2]),.dout(n1311),.clk(gclk));
	jand g1246(.dina(n1311),.dinb(w_n384_0[2]),.dout(n1312),.clk(gclk));
	jand g1247(.dina(w_n1312_0[1]),.dinb(w_n1310_0[1]),.dout(n1313),.clk(gclk));
	jand g1248(.dina(w_n458_1[1]),.dinb(w_n422_2[1]),.dout(n1314),.clk(gclk));
	jand g1249(.dina(n1314),.dinb(w_n295_2[2]),.dout(n1315),.clk(gclk));
	jand g1250(.dina(n1315),.dinb(w_n843_0[0]),.dout(n1316),.clk(gclk));
	jand g1251(.dina(n1316),.dinb(w_n677_0[1]),.dout(n1317),.clk(gclk));
	jand g1252(.dina(n1317),.dinb(n1313),.dout(n1318),.clk(gclk));
	jand g1253(.dina(n1318),.dinb(w_n1307_0[1]),.dout(n1319),.clk(gclk));
	jor g1254(.dina(w_n521_0[0]),.dinb(w_n411_0[0]),.dout(n1320),.clk(gclk));
	jor g1255(.dina(w_n290_0[0]),.dinb(w_n228_0[0]),.dout(n1321),.clk(gclk));
	jor g1256(.dina(n1321),.dinb(n1320),.dout(n1322),.clk(gclk));
	jor g1257(.dina(w_n593_0[0]),.dinb(w_n137_0[0]),.dout(n1323),.clk(gclk));
	jor g1258(.dina(n1323),.dinb(w_n156_0[0]),.dout(n1324),.clk(gclk));
	jor g1259(.dina(n1324),.dinb(w_n1322_0[1]),.dout(n1325),.clk(gclk));
	jnot g1260(.din(w_n1325_0[1]),.dout(n1326),.clk(gclk));
	jand g1261(.dina(n1326),.dinb(w_n741_1[0]),.dout(n1327),.clk(gclk));
	jand g1262(.dina(w_n781_1[2]),.dinb(w_n451_2[1]),.dout(n1328),.clk(gclk));
	jor g1263(.dina(w_n670_0[0]),.dinb(w_n644_0[0]),.dout(n1329),.clk(gclk));
	jnot g1264(.din(w_n1329_0[1]),.dout(n1330),.clk(gclk));
	jand g1265(.dina(n1330),.dinb(w_n1021_0[0]),.dout(n1331),.clk(gclk));
	jand g1266(.dina(n1331),.dinb(w_n1328_0[2]),.dout(n1332),.clk(gclk));
	jand g1267(.dina(w_n428_0[1]),.dinb(w_n301_1[1]),.dout(n1333),.clk(gclk));
	jand g1268(.dina(n1333),.dinb(w_n771_1[2]),.dout(n1334),.clk(gclk));
	jand g1269(.dina(n1334),.dinb(w_n1332_0[1]),.dout(n1335),.clk(gclk));
	jand g1270(.dina(n1335),.dinb(n1327),.dout(n1336),.clk(gclk));
	jand g1271(.dina(n1336),.dinb(w_n1319_0[1]),.dout(n1337),.clk(gclk));
	jand g1272(.dina(n1337),.dinb(w_n1299_0[1]),.dout(n1338),.clk(gclk));
	jor g1273(.dina(w_n1338_0[2]),.dinb(w_n1243_2[0]),.dout(n1339),.clk(gclk));
	jand g1274(.dina(w_n1339_0[2]),.dinb(w_n604_0[1]),.dout(n1340),.clk(gclk));
	jand g1275(.dina(w_n1340_0[2]),.dinb(w_n1283_12[2]),.dout(n1341),.clk(gclk));
	jnot g1276(.din(n1341),.dout(n1342),.clk(gclk));
	jand g1277(.dina(w_a22_2[1]),.dinb(w_a6_0[2]),.dout(n1343),.clk(gclk));
	jand g1278(.dina(w_n81_0[0]),.dinb(w_a6_0[1]),.dout(n1344),.clk(gclk));
	jnot g1279(.din(n1344),.dout(n1345),.clk(gclk));
	jand g1280(.dina(n1345),.dinb(w_n336_0[0]),.dout(n1346),.clk(gclk));
	jor g1281(.dina(n1346),.dinb(n1343),.dout(n1347),.clk(gclk));
	jand g1282(.dina(w_n1347_6[1]),.dinb(w_n335_5[0]),.dout(n1348),.clk(gclk));
	jand g1283(.dina(w_n1348_0[1]),.dinb(w_n1342_0[1]),.dout(n1349),.clk(gclk));
	jnot g1284(.din(n1349),.dout(n1350),.clk(gclk));
	jand g1285(.dina(w_n1350_0[1]),.dinb(w_n1245_0[1]),.dout(n1351),.clk(gclk));
	jor g1286(.dina(w_n1351_0[1]),.dinb(w_n1163_0[1]),.dout(n1352),.clk(gclk));
	jand g1287(.dina(n1352),.dinb(n1161),.dout(n1353),.clk(gclk));
	jnot g1288(.din(n1353),.dout(n1354),.clk(gclk));
	jnot g1289(.din(w_n338_0[2]),.dout(n1355),.clk(gclk));
	jxor g1290(.dina(w_n688_0[1]),.dinb(w_n1185_1[1]),.dout(n1356),.clk(gclk));
	jnot g1291(.din(w_n1356_1[1]),.dout(n1357),.clk(gclk));
	jand g1292(.dina(n1357),.dinb(w_n954_22[1]),.dout(n1358),.clk(gclk));
	jnot g1293(.din(w_n1358_0[1]),.dout(n1359),.clk(gclk));
	jand g1294(.dina(n1359),.dinb(w_n691_1[0]),.dout(n1360),.clk(gclk));
	jand g1295(.dina(w_n688_0[0]),.dinb(w_n1185_1[0]),.dout(n1361),.clk(gclk));
	jor g1296(.dina(w_n1361_0[1]),.dinb(w_n968_0[0]),.dout(n1362),.clk(gclk));
	jand g1297(.dina(w_n1362_0[2]),.dinb(w_n1358_0[0]),.dout(n1363),.clk(gclk));
	jor g1298(.dina(n1363),.dinb(n1360),.dout(n1364),.clk(gclk));
	jnot g1299(.din(w_n1364_0[1]),.dout(n1365),.clk(gclk));
	jand g1300(.dina(n1365),.dinb(n1355),.dout(n1366),.clk(gclk));
	jxor g1301(.dina(w_n1364_0[0]),.dinb(w_n338_0[1]),.dout(n1367),.clk(gclk));
	jand g1302(.dina(w_n960_4[1]),.dinb(w_n956_4[0]),.dout(n1368),.clk(gclk));
	jand g1303(.dina(w_n961_4[0]),.dinb(w_n952_4[0]),.dout(n1369),.clk(gclk));
	jor g1304(.dina(n1369),.dinb(n1368),.dout(n1370),.clk(gclk));
	jand g1305(.dina(w_n980_5[0]),.dinb(w_n971_3[2]),.dout(n1371),.clk(gclk));
	jand g1306(.dina(w_n981_3[1]),.dinb(w_n966_4[0]),.dout(n1372),.clk(gclk));
	jor g1307(.dina(n1372),.dinb(n1371),.dout(n1373),.clk(gclk));
	jor g1308(.dina(n1373),.dinb(n1370),.dout(n1374),.clk(gclk));
	jnot g1309(.din(n1374),.dout(n1375),.clk(gclk));
	jand g1310(.dina(w_n1375_0[1]),.dinb(w_n1367_0[1]),.dout(n1376),.clk(gclk));
	jor g1311(.dina(n1376),.dinb(n1366),.dout(n1377),.clk(gclk));
	jand g1312(.dina(w_n1377_0[1]),.dinb(w_n1354_0[1]),.dout(n1378),.clk(gclk));
	jxor g1313(.dina(w_n700_0[0]),.dinb(w_n693_0[0]),.dout(n1379),.clk(gclk));
	jxor g1314(.dina(w_n1377_0[0]),.dinb(w_n1354_0[0]),.dout(n1380),.clk(gclk));
	jand g1315(.dina(w_n1380_0[1]),.dinb(w_n1379_0[1]),.dout(n1381),.clk(gclk));
	jor g1316(.dina(n1381),.dinb(n1378),.dout(n1382),.clk(gclk));
	jxor g1317(.dina(w_n1093_0[0]),.dinb(w_n1085_0[0]),.dout(n1383),.clk(gclk));
	jand g1318(.dina(w_n1383_0[1]),.dinb(w_n1382_0[1]),.dout(n1384),.clk(gclk));
	jxor g1319(.dina(w_n1383_0[0]),.dinb(w_n1382_0[0]),.dout(n1385),.clk(gclk));
	jxor g1320(.dina(w_n1069_0[0]),.dinb(w_n1068_0[0]),.dout(n1386),.clk(gclk));
	jand g1321(.dina(w_n1386_0[1]),.dinb(w_n1385_0[1]),.dout(n1387),.clk(gclk));
	jor g1322(.dina(n1387),.dinb(n1384),.dout(n1388),.clk(gclk));
	jxor g1323(.dina(w_n1111_0[0]),.dinb(w_n1078_0[0]),.dout(n1389),.clk(gclk));
	jand g1324(.dina(w_n1389_0[1]),.dinb(w_n1388_0[1]),.dout(n1390),.clk(gclk));
	jnot g1325(.din(w_n337_5[0]),.dout(n1391),.clk(gclk));
	jand g1326(.dina(w_n799_2[1]),.dinb(w_n1391_5[2]),.dout(n1392),.clk(gclk));
	jnot g1327(.din(n1392),.dout(n1393),.clk(gclk));
	jand g1328(.dina(w_n804_2[2]),.dinb(w_n337_4[2]),.dout(n1394),.clk(gclk));
	jnot g1329(.din(n1394),.dout(n1395),.clk(gclk));
	jxor g1330(.dina(w_n1143_9[0]),.dinb(w_n334_1[0]),.dout(n1396),.clk(gclk));
	jor g1331(.dina(n1396),.dinb(w_n795_1[0]),.dout(n1397),.clk(gclk));
	jand g1332(.dina(n1397),.dinb(n1395),.dout(n1398),.clk(gclk));
	jand g1333(.dina(n1398),.dinb(n1393),.dout(n1399),.clk(gclk));
	jand g1334(.dina(w_n1035_0[1]),.dinb(w_n794_3[2]),.dout(n1400),.clk(gclk));
	jand g1335(.dina(w_n1038_0[1]),.dinb(w_n708_5[0]),.dout(n1401),.clk(gclk));
	jor g1336(.dina(n1401),.dinb(n1400),.dout(n1402),.clk(gclk));
	jand g1337(.dina(w_n1057_4[1]),.dinb(w_n1043_3[0]),.dout(n1403),.clk(gclk));
	jand g1338(.dina(w_n1059_5[0]),.dinb(w_n1049_3[0]),.dout(n1404),.clk(gclk));
	jor g1339(.dina(n1404),.dinb(n1403),.dout(n1405),.clk(gclk));
	jnot g1340(.din(n1405),.dout(n1406),.clk(gclk));
	jand g1341(.dina(n1406),.dinb(n1402),.dout(n1407),.clk(gclk));
	jand g1342(.dina(w_n1407_0[1]),.dinb(w_n1399_0[1]),.dout(n1408),.clk(gclk));
	jxor g1343(.dina(w_n1407_0[0]),.dinb(w_n1399_0[0]),.dout(n1409),.clk(gclk));
	jnot g1344(.din(w_n1362_0[1]),.dout(n1410),.clk(gclk));
	jor g1345(.dina(n1410),.dinb(w_n1356_1[0]),.dout(n1411),.clk(gclk));
	jand g1346(.dina(w_n1411_2[2]),.dinb(w_n960_4[0]),.dout(n1412),.clk(gclk));
	jnot g1347(.din(w_n691_0[2]),.dout(n1413),.clk(gclk));
	jor g1348(.dina(w_n1356_0[2]),.dinb(w_n1413_0[1]),.dout(n1414),.clk(gclk));
	jand g1349(.dina(w_n1414_2[2]),.dinb(w_n961_3[2]),.dout(n1415),.clk(gclk));
	jor g1350(.dina(n1415),.dinb(n1412),.dout(n1416),.clk(gclk));
	jor g1351(.dina(w_n1361_0[0]),.dinb(w_n691_0[1]),.dout(n1417),.clk(gclk));
	jnot g1352(.din(w_n1417_0[1]),.dout(n1418),.clk(gclk));
	jand g1353(.dina(w_n1418_4[1]),.dinb(w_n954_22[0]),.dout(n1419),.clk(gclk));
	jor g1354(.dina(w_n1362_0[0]),.dinb(w_n690_0[0]),.dout(n1420),.clk(gclk));
	jnot g1355(.din(w_n1420_0[1]),.dout(n1421),.clk(gclk));
	jand g1356(.dina(w_n1421_4[1]),.dinb(w_n820_4[2]),.dout(n1422),.clk(gclk));
	jor g1357(.dina(n1422),.dinb(n1419),.dout(n1423),.clk(gclk));
	jnot g1358(.din(n1423),.dout(n1424),.clk(gclk));
	jand g1359(.dina(n1424),.dinb(n1416),.dout(n1425),.clk(gclk));
	jand g1360(.dina(w_n1425_0[1]),.dinb(w_n1409_0[1]),.dout(n1426),.clk(gclk));
	jor g1361(.dina(n1426),.dinb(n1408),.dout(n1427),.clk(gclk));
	jxor g1362(.dina(w_n1375_0[0]),.dinb(w_n1367_0[0]),.dout(n1428),.clk(gclk));
	jand g1363(.dina(w_n1428_0[1]),.dinb(w_n1427_0[1]),.dout(n1429),.clk(gclk));
	jxor g1364(.dina(w_n1351_0[0]),.dinb(w_n1163_0[0]),.dout(n1430),.clk(gclk));
	jxor g1365(.dina(w_n1428_0[0]),.dinb(w_n1427_0[0]),.dout(n1431),.clk(gclk));
	jand g1366(.dina(w_n1431_0[1]),.dinb(w_n1430_0[1]),.dout(n1432),.clk(gclk));
	jor g1367(.dina(n1432),.dinb(n1429),.dout(n1433),.clk(gclk));
	jxor g1368(.dina(w_n1066_0[0]),.dinb(w_n1055_0[0]),.dout(n1434),.clk(gclk));
	jand g1369(.dina(w_n1434_0[1]),.dinb(w_n1433_0[1]),.dout(n1435),.clk(gclk));
	jxor g1370(.dina(w_n1434_0[0]),.dinb(w_n1433_0[0]),.dout(n1436),.clk(gclk));
	jxor g1371(.dina(w_n1380_0[0]),.dinb(w_n1379_0[0]),.dout(n1437),.clk(gclk));
	jand g1372(.dina(w_n1437_0[1]),.dinb(w_n1436_0[1]),.dout(n1438),.clk(gclk));
	jor g1373(.dina(n1438),.dinb(n1435),.dout(n1439),.clk(gclk));
	jxor g1374(.dina(w_n1386_0[0]),.dinb(w_n1385_0[0]),.dout(n1440),.clk(gclk));
	jand g1375(.dina(w_n1440_0[1]),.dinb(w_n1439_0[1]),.dout(n1441),.clk(gclk));
	jand g1376(.dina(w_n1342_0[0]),.dinb(w_n1245_0[0]),.dout(n1442),.clk(gclk));
	jnot g1377(.din(w_n1442_0[1]),.dout(n1443),.clk(gclk));
	jand g1378(.dina(n1443),.dinb(w_n1348_0[0]),.dout(n1444),.clk(gclk));
	jand g1379(.dina(w_n1442_0[0]),.dinb(w_n1350_0[0]),.dout(n1445),.clk(gclk));
	jor g1380(.dina(n1445),.dinb(n1444),.dout(n1446),.clk(gclk));
	jand g1381(.dina(w_n981_3[0]),.dinb(w_n952_3[2]),.dout(n1447),.clk(gclk));
	jand g1382(.dina(w_n980_4[2]),.dinb(w_n956_3[2]),.dout(n1448),.clk(gclk));
	jor g1383(.dina(n1448),.dinb(n1447),.dout(n1449),.clk(gclk));
	jand g1384(.dina(w_n966_3[2]),.dinb(w_n808_12[1]),.dout(n1450),.clk(gclk));
	jand g1385(.dina(w_n971_3[1]),.dinb(w_n803_7[0]),.dout(n1451),.clk(gclk));
	jor g1386(.dina(n1451),.dinb(n1450),.dout(n1452),.clk(gclk));
	jor g1387(.dina(n1452),.dinb(n1449),.dout(n1453),.clk(gclk));
	jnot g1388(.din(n1453),.dout(n1454),.clk(gclk));
	jand g1389(.dina(w_n1454_0[1]),.dinb(w_n1446_0[1]),.dout(n1455),.clk(gclk));
	jand g1390(.dina(w_n335_4[2]),.dinb(w_n55_9[1]),.dout(n1456),.clk(gclk));
	jand g1391(.dina(w_n1456_0[1]),.dinb(w_n1283_12[1]),.dout(n1457),.clk(gclk));
	jxor g1392(.dina(w_n1456_0[0]),.dinb(w_n1283_12[0]),.dout(n1458),.clk(gclk));
	jnot g1393(.din(w_n1027_0[0]),.dout(n1459),.clk(gclk));
	jnot g1394(.din(w_n1285_0[0]),.dout(n1460),.clk(gclk));
	jor g1395(.dina(n1460),.dinb(w_n571_0[0]),.dout(n1461),.clk(gclk));
	jor g1396(.dina(n1461),.dinb(n1459),.dout(n1462),.clk(gclk));
	jnot g1397(.din(w_n733_0[2]),.dout(n1463),.clk(gclk));
	jor g1398(.dina(w_n1288_0[0]),.dinb(n1463),.dout(n1464),.clk(gclk));
	jnot g1399(.din(w_n243_3[1]),.dout(n1465),.clk(gclk));
	jor g1400(.dina(w_n631_0[0]),.dinb(n1465),.dout(n1466),.clk(gclk));
	jor g1401(.dina(w_n1259_0[0]),.dinb(n1466),.dout(n1467),.clk(gclk));
	jor g1402(.dina(n1467),.dinb(n1464),.dout(n1468),.clk(gclk));
	jnot g1403(.din(w_n282_2[2]),.dout(n1469),.clk(gclk));
	jor g1404(.dina(w_n284_0[0]),.dinb(n1469),.dout(n1470),.clk(gclk));
	jor g1405(.dina(w_n1293_0[0]),.dinb(n1470),.dout(n1471),.clk(gclk));
	jor g1406(.dina(n1471),.dinb(w_n894_0[0]),.dout(n1472),.clk(gclk));
	jor g1407(.dina(n1472),.dinb(n1468),.dout(n1473),.clk(gclk));
	jor g1408(.dina(n1473),.dinb(w_n1217_0[0]),.dout(n1474),.clk(gclk));
	jor g1409(.dina(n1474),.dinb(n1462),.dout(n1475),.clk(gclk));
	jnot g1410(.din(w_n511_0[2]),.dout(n1476),.clk(gclk));
	jnot g1411(.din(w_n402_1[1]),.dout(n1477),.clk(gclk));
	jor g1412(.dina(n1477),.dinb(w_n322_0[0]),.dout(n1478),.clk(gclk));
	jor g1413(.dina(n1478),.dinb(n1476),.dout(n1479),.clk(gclk));
	jor g1414(.dina(n1479),.dinb(w_n1017_0[0]),.dout(n1480),.clk(gclk));
	jor g1415(.dina(n1480),.dinb(w_n1302_0[0]),.dout(n1481),.clk(gclk));
	jnot g1416(.din(w_n1312_0[0]),.dout(n1482),.clk(gclk));
	jor g1417(.dina(n1482),.dinb(w_n1309_0[0]),.dout(n1483),.clk(gclk));
	jnot g1418(.din(w_n676_1[0]),.dout(n1484),.clk(gclk));
	jor g1419(.dina(n1484),.dinb(w_n460_0[0]),.dout(n1485),.clk(gclk));
	jnot g1420(.din(w_n147_3[0]),.dout(n1486),.clk(gclk));
	jand g1421(.dina(w_n212_1[0]),.dinb(w_n141_0[2]),.dout(n1487),.clk(gclk));
	jand g1422(.dina(w_n468_0[0]),.dinb(w_n96_1[2]),.dout(n1488),.clk(gclk));
	jor g1423(.dina(n1488),.dinb(n1487),.dout(n1489),.clk(gclk));
	jor g1424(.dina(n1489),.dinb(n1486),.dout(n1490),.clk(gclk));
	jnot g1425(.din(w_n295_2[1]),.dout(n1491),.clk(gclk));
	jor g1426(.dina(w_n1232_0[0]),.dinb(w_n985_0[0]),.dout(n1492),.clk(gclk));
	jor g1427(.dina(n1492),.dinb(n1491),.dout(n1493),.clk(gclk));
	jor g1428(.dina(n1493),.dinb(n1490),.dout(n1494),.clk(gclk));
	jor g1429(.dina(n1494),.dinb(n1485),.dout(n1495),.clk(gclk));
	jor g1430(.dina(n1495),.dinb(n1483),.dout(n1496),.clk(gclk));
	jor g1431(.dina(n1496),.dinb(n1481),.dout(n1497),.clk(gclk));
	jnot g1432(.din(w_n741_0[2]),.dout(n1498),.clk(gclk));
	jor g1433(.dina(w_n1325_0[0]),.dinb(n1498),.dout(n1499),.clk(gclk));
	jnot g1434(.din(w_n1328_0[1]),.dout(n1500),.clk(gclk));
	jor g1435(.dina(w_n764_0[1]),.dinb(w_n726_0[0]),.dout(n1501),.clk(gclk));
	jor g1436(.dina(w_n1329_0[0]),.dinb(n1501),.dout(n1502),.clk(gclk));
	jor g1437(.dina(n1502),.dinb(n1500),.dout(n1503),.clk(gclk));
	jnot g1438(.din(w_n771_1[1]),.dout(n1504),.clk(gclk));
	jnot g1439(.din(w_n427_2[0]),.dout(n1505),.clk(gclk));
	jor g1440(.dina(n1505),.dinb(w_n425_0[0]),.dout(n1506),.clk(gclk));
	jor g1441(.dina(n1506),.dinb(w_n300_0[0]),.dout(n1507),.clk(gclk));
	jor g1442(.dina(n1507),.dinb(n1504),.dout(n1508),.clk(gclk));
	jor g1443(.dina(n1508),.dinb(n1503),.dout(n1509),.clk(gclk));
	jor g1444(.dina(n1509),.dinb(n1499),.dout(n1510),.clk(gclk));
	jor g1445(.dina(n1510),.dinb(n1497),.dout(n1511),.clk(gclk));
	jor g1446(.dina(n1511),.dinb(n1475),.dout(n1512),.clk(gclk));
	jand g1447(.dina(n1512),.dinb(w_n1283_11[2]),.dout(n1513),.clk(gclk));
	jor g1448(.dina(w_n1513_0[1]),.dinb(w_n1185_0[2]),.dout(n1514),.clk(gclk));
	jxor g1449(.dina(w_n1338_0[1]),.dinb(w_n1243_1[2]),.dout(n1515),.clk(gclk));
	jnot g1450(.din(w_n1515_0[1]),.dout(n1516),.clk(gclk));
	jand g1451(.dina(n1516),.dinb(w_n954_21[2]),.dout(n1517),.clk(gclk));
	jnot g1452(.din(w_n1517_0[1]),.dout(n1518),.clk(gclk));
	jand g1453(.dina(n1518),.dinb(w_n1514_0[1]),.dout(n1519),.clk(gclk));
	jand g1454(.dina(w_n1338_0[0]),.dinb(w_n1243_1[1]),.dout(n1520),.clk(gclk));
	jor g1455(.dina(w_n1520_0[2]),.dinb(w_n604_0[0]),.dout(n1521),.clk(gclk));
	jand g1456(.dina(w_n1521_0[1]),.dinb(w_n1517_0[0]),.dout(n1522),.clk(gclk));
	jor g1457(.dina(n1522),.dinb(n1519),.dout(n1523),.clk(gclk));
	jnot g1458(.din(n1523),.dout(n1524),.clk(gclk));
	jand g1459(.dina(w_n1524_0[1]),.dinb(w_n1458_0[1]),.dout(n1525),.clk(gclk));
	jor g1460(.dina(n1525),.dinb(n1457),.dout(n1526),.clk(gclk));
	jxor g1461(.dina(w_n1454_0[0]),.dinb(w_n1446_0[0]),.dout(n1527),.clk(gclk));
	jand g1462(.dina(w_n1527_0[1]),.dinb(w_n1526_0[1]),.dout(n1528),.clk(gclk));
	jor g1463(.dina(n1528),.dinb(n1455),.dout(n1529),.clk(gclk));
	jand g1464(.dina(w_n1418_4[0]),.dinb(w_n960_3[2]),.dout(n1530),.clk(gclk));
	jand g1465(.dina(w_n1421_4[0]),.dinb(w_n961_3[1]),.dout(n1531),.clk(gclk));
	jor g1466(.dina(n1531),.dinb(n1530),.dout(n1532),.clk(gclk));
	jnot g1467(.din(w_n1411_2[1]),.dout(n1533),.clk(gclk));
	jand g1468(.dina(w_n1533_1[2]),.dinb(w_n980_4[1]),.dout(n1534),.clk(gclk));
	jnot g1469(.din(w_n1414_2[1]),.dout(n1535),.clk(gclk));
	jand g1470(.dina(w_n1535_1[2]),.dinb(w_n981_2[2]),.dout(n1536),.clk(gclk));
	jor g1471(.dina(n1536),.dinb(n1534),.dout(n1537),.clk(gclk));
	jor g1472(.dina(n1537),.dinb(n1532),.dout(n1538),.clk(gclk));
	jnot g1473(.din(n1538),.dout(n1539),.clk(gclk));
	jand g1474(.dina(w_n970_0[1]),.dinb(w_n708_4[2]),.dout(n1540),.clk(gclk));
	jnot g1475(.din(w_n966_3[1]),.dout(n1541),.clk(gclk));
	jand g1476(.dina(w_n1541_0[1]),.dinb(w_n794_3[1]),.dout(n1542),.clk(gclk));
	jor g1477(.dina(n1542),.dinb(n1540),.dout(n1543),.clk(gclk));
	jand g1478(.dina(w_n956_3[1]),.dinb(w_n803_6[2]),.dout(n1544),.clk(gclk));
	jand g1479(.dina(w_n952_3[1]),.dinb(w_n808_12[0]),.dout(n1545),.clk(gclk));
	jor g1480(.dina(n1545),.dinb(n1544),.dout(n1546),.clk(gclk));
	jnot g1481(.din(n1546),.dout(n1547),.clk(gclk));
	jand g1482(.dina(n1547),.dinb(n1543),.dout(n1548),.clk(gclk));
	jand g1483(.dina(w_n1548_0[1]),.dinb(w_n1539_0[1]),.dout(n1549),.clk(gclk));
	jxor g1484(.dina(w_n1548_0[0]),.dinb(w_n1539_0[0]),.dout(n1550),.clk(gclk));
	jand g1485(.dina(w_n1042_0[0]),.dinb(w_n699_12[2]),.dout(n1551),.clk(gclk));
	jand g1486(.dina(w_n1152_0[0]),.dinb(w_n1143_8[2]),.dout(n1552),.clk(gclk));
	jor g1487(.dina(n1552),.dinb(n1551),.dout(n1553),.clk(gclk));
	jand g1488(.dina(w_n1057_4[0]),.dinb(w_n1037_2[1]),.dout(n1554),.clk(gclk));
	jand g1489(.dina(w_n1059_4[2]),.dinb(w_n1034_2[1]),.dout(n1555),.clk(gclk));
	jor g1490(.dina(n1555),.dinb(n1554),.dout(n1556),.clk(gclk));
	jnot g1491(.din(n1556),.dout(n1557),.clk(gclk));
	jand g1492(.dina(n1557),.dinb(n1553),.dout(n1558),.clk(gclk));
	jand g1493(.dina(w_n1558_0[1]),.dinb(w_n1550_0[1]),.dout(n1559),.clk(gclk));
	jor g1494(.dina(n1559),.dinb(n1549),.dout(n1560),.clk(gclk));
	jxor g1495(.dina(w_n1425_0[0]),.dinb(w_n1409_0[0]),.dout(n1561),.clk(gclk));
	jand g1496(.dina(w_n1561_0[1]),.dinb(w_n1560_0[1]),.dout(n1562),.clk(gclk));
	jand g1497(.dina(w_n335_4[1]),.dinb(w_n75_5[1]),.dout(n1563),.clk(gclk));
	jand g1498(.dina(w_n1563_0[1]),.dinb(w_n1283_11[1]),.dout(n1564),.clk(gclk));
	jxor g1499(.dina(w_n1563_0[0]),.dinb(w_n1283_11[0]),.dout(n1565),.clk(gclk));
	jor g1500(.dina(w_n1521_0[0]),.dinb(w_n1513_0[0]),.dout(n1566),.clk(gclk));
	jand g1501(.dina(w_n1566_3[1]),.dinb(w_n820_4[1]),.dout(n1567),.clk(gclk));
	jor g1502(.dina(w_n1520_0[1]),.dinb(w_n1514_0[0]),.dout(n1568),.clk(gclk));
	jand g1503(.dina(w_n1568_3[1]),.dinb(w_n954_21[1]),.dout(n1569),.clk(gclk));
	jor g1504(.dina(n1569),.dinb(n1567),.dout(n1570),.clk(gclk));
	jor g1505(.dina(w_n1515_0[0]),.dinb(w_n1340_0[1]),.dout(n1571),.clk(gclk));
	jnot g1506(.din(w_n1571_1[1]),.dout(n1572),.clk(gclk));
	jand g1507(.dina(w_n1572_3[1]),.dinb(w_n961_3[0]),.dout(n1573),.clk(gclk));
	jnot g1508(.din(w_n1520_0[0]),.dout(n1574),.clk(gclk));
	jor g1509(.dina(w_n1339_0[1]),.dinb(w_n1185_0[1]),.dout(n1575),.clk(gclk));
	jand g1510(.dina(w_n1575_0[1]),.dinb(w_n1574_0[1]),.dout(n1576),.clk(gclk));
	jnot g1511(.din(w_n1576_0[2]),.dout(n1577),.clk(gclk));
	jand g1512(.dina(w_n1577_3[1]),.dinb(w_n960_3[1]),.dout(n1578),.clk(gclk));
	jor g1513(.dina(n1578),.dinb(n1573),.dout(n1579),.clk(gclk));
	jnot g1514(.din(n1579),.dout(n1580),.clk(gclk));
	jand g1515(.dina(n1580),.dinb(n1570),.dout(n1581),.clk(gclk));
	jand g1516(.dina(w_n1581_0[1]),.dinb(w_n1565_0[1]),.dout(n1582),.clk(gclk));
	jor g1517(.dina(n1582),.dinb(n1564),.dout(n1583),.clk(gclk));
	jnot g1518(.din(w_n1347_6[0]),.dout(n1584),.clk(gclk));
	jand g1519(.dina(w_n1584_4[2]),.dinb(w_n799_2[0]),.dout(n1585),.clk(gclk));
	jand g1520(.dina(w_n1347_5[2]),.dinb(w_n804_2[1]),.dout(n1586),.clk(gclk));
	jor g1521(.dina(n1586),.dinb(n1585),.dout(n1587),.clk(gclk));
	jand g1522(.dina(w_n789_3[0]),.dinb(w_n1391_5[1]),.dout(n1588),.clk(gclk));
	jor g1523(.dina(n1588),.dinb(n1587),.dout(n1591),.clk(gclk));
	jnot g1524(.din(n1591),.dout(n1592),.clk(gclk));
	jand g1525(.dina(w_n1592_0[1]),.dinb(w_n1583_0[1]),.dout(n1593),.clk(gclk));
	jxor g1526(.dina(w_n1592_0[0]),.dinb(w_n1583_0[0]),.dout(n1594),.clk(gclk));
	jnot g1527(.din(w_n952_3[0]),.dout(n1595),.clk(gclk));
	jand g1528(.dina(w_n1595_0[1]),.dinb(w_n794_3[0]),.dout(n1596),.clk(gclk));
	jnot g1529(.din(w_n956_3[0]),.dout(n1597),.clk(gclk));
	jand g1530(.dina(w_n1597_0[1]),.dinb(w_n708_4[1]),.dout(n1598),.clk(gclk));
	jor g1531(.dina(n1598),.dinb(n1596),.dout(n1599),.clk(gclk));
	jand g1532(.dina(w_n1057_3[2]),.dinb(w_n971_3[0]),.dout(n1600),.clk(gclk));
	jand g1533(.dina(w_n1059_4[1]),.dinb(w_n966_3[0]),.dout(n1601),.clk(gclk));
	jor g1534(.dina(n1601),.dinb(n1600),.dout(n1602),.clk(gclk));
	jnot g1535(.din(n1602),.dout(n1603),.clk(gclk));
	jand g1536(.dina(n1603),.dinb(n1599),.dout(n1604),.clk(gclk));
	jand g1537(.dina(w_n1411_2[0]),.dinb(w_n803_6[1]),.dout(n1605),.clk(gclk));
	jand g1538(.dina(w_n1414_2[0]),.dinb(w_n808_11[2]),.dout(n1606),.clk(gclk));
	jor g1539(.dina(n1606),.dinb(n1605),.dout(n1607),.clk(gclk));
	jand g1540(.dina(w_n1418_3[2]),.dinb(w_n980_4[0]),.dout(n1608),.clk(gclk));
	jand g1541(.dina(w_n1421_3[2]),.dinb(w_n981_2[1]),.dout(n1609),.clk(gclk));
	jor g1542(.dina(n1609),.dinb(n1608),.dout(n1610),.clk(gclk));
	jnot g1543(.din(n1610),.dout(n1611),.clk(gclk));
	jand g1544(.dina(n1611),.dinb(n1607),.dout(n1612),.clk(gclk));
	jand g1545(.dina(w_n1612_0[1]),.dinb(w_n1604_0[1]),.dout(n1613),.clk(gclk));
	jxor g1546(.dina(w_n1612_0[0]),.dinb(w_n1604_0[0]),.dout(n1614),.clk(gclk));
	jand g1547(.dina(w_n1035_0[0]),.dinb(w_n1143_8[1]),.dout(n1615),.clk(gclk));
	jand g1548(.dina(w_n1038_0[0]),.dinb(w_n699_12[1]),.dout(n1616),.clk(gclk));
	jor g1549(.dina(n1616),.dinb(n1615),.dout(n1617),.clk(gclk));
	jand g1550(.dina(w_n1043_2[2]),.dinb(w_n337_4[1]),.dout(n1618),.clk(gclk));
	jand g1551(.dina(w_n1049_2[2]),.dinb(w_n1391_5[0]),.dout(n1619),.clk(gclk));
	jor g1552(.dina(n1619),.dinb(n1618),.dout(n1620),.clk(gclk));
	jnot g1553(.din(n1620),.dout(n1621),.clk(gclk));
	jand g1554(.dina(n1621),.dinb(n1617),.dout(n1622),.clk(gclk));
	jand g1555(.dina(w_n1622_0[1]),.dinb(w_n1614_0[1]),.dout(n1623),.clk(gclk));
	jor g1556(.dina(n1623),.dinb(n1613),.dout(n1624),.clk(gclk));
	jand g1557(.dina(w_n1624_0[1]),.dinb(w_n1594_0[1]),.dout(n1625),.clk(gclk));
	jor g1558(.dina(n1625),.dinb(n1593),.dout(n1626),.clk(gclk));
	jxor g1559(.dina(w_n1561_0[0]),.dinb(w_n1560_0[0]),.dout(n1627),.clk(gclk));
	jand g1560(.dina(w_n1627_0[1]),.dinb(w_n1626_0[1]),.dout(n1628),.clk(gclk));
	jor g1561(.dina(n1628),.dinb(n1562),.dout(n1629),.clk(gclk));
	jand g1562(.dina(w_n1629_0[1]),.dinb(w_n1529_0[1]),.dout(n1630),.clk(gclk));
	jxor g1563(.dina(w_n1431_0[0]),.dinb(w_n1430_0[0]),.dout(n1631),.clk(gclk));
	jxor g1564(.dina(w_n1629_0[0]),.dinb(w_n1529_0[0]),.dout(n1632),.clk(gclk));
	jand g1565(.dina(w_n1632_0[1]),.dinb(w_n1631_0[1]),.dout(n1633),.clk(gclk));
	jor g1566(.dina(n1633),.dinb(n1630),.dout(n1634),.clk(gclk));
	jxor g1567(.dina(w_n1437_0[0]),.dinb(w_n1436_0[0]),.dout(n1635),.clk(gclk));
	jand g1568(.dina(w_n1635_0[1]),.dinb(w_n1634_0[1]),.dout(n1636),.clk(gclk));
	jxor g1569(.dina(w_n1524_0[0]),.dinb(w_n1458_0[0]),.dout(n1637),.clk(gclk));
	jxor g1570(.dina(w_n1558_0[0]),.dinb(w_n1550_0[0]),.dout(n1638),.clk(gclk));
	jand g1571(.dina(w_n1638_0[1]),.dinb(w_n1637_0[1]),.dout(n1639),.clk(gclk));
	jand g1572(.dina(w_n335_4[0]),.dinb(w_n58_4[1]),.dout(n1640),.clk(gclk));
	jand g1573(.dina(w_n724_1[2]),.dinb(w_n267_0[2]),.dout(n1641),.clk(gclk));
	jand g1574(.dina(w_n1641_0[1]),.dinb(w_n324_0[2]),.dout(n1642),.clk(gclk));
	jand g1575(.dina(w_n713_0[0]),.dinb(w_n676_0[2]),.dout(n1643),.clk(gclk));
	jand g1576(.dina(n1643),.dinb(n1642),.dout(n1644),.clk(gclk));
	jnot g1577(.din(n1644),.dout(n1645),.clk(gclk));
	jand g1578(.dina(w_n905_0[0]),.dinb(w_n232_1[1]),.dout(n1646),.clk(gclk));
	jnot g1579(.din(w_n1646_0[2]),.dout(n1647),.clk(gclk));
	jand g1580(.dina(w_n668_2[1]),.dinb(w_n303_2[2]),.dout(n1648),.clk(gclk));
	jand g1581(.dina(n1648),.dinb(w_n216_3[0]),.dout(n1649),.clk(gclk));
	jnot g1582(.din(n1649),.dout(n1650),.clk(gclk));
	jor g1583(.dina(n1650),.dinb(w_n863_0[0]),.dout(n1651),.clk(gclk));
	jor g1584(.dina(n1651),.dinb(n1647),.dout(n1652),.clk(gclk));
	jor g1585(.dina(n1652),.dinb(n1645),.dout(n1653),.clk(gclk));
	jand g1586(.dina(w_n592_2[2]),.dinb(w_n291_1[2]),.dout(n1654),.clk(gclk));
	jand g1587(.dina(n1654),.dinb(w_n849_1[1]),.dout(n1655),.clk(gclk));
	jnot g1588(.din(n1655),.dout(n1656),.clk(gclk));
	jnot g1589(.din(w_n994_0[0]),.dout(n1657),.clk(gclk));
	jor g1590(.dina(w_n764_0[0]),.dinb(w_n588_0[1]),.dout(n1658),.clk(gclk));
	jor g1591(.dina(w_n1658_0[1]),.dinb(n1657),.dout(n1659),.clk(gclk));
	jor g1592(.dina(n1659),.dinb(w_n986_0[0]),.dout(n1660),.clk(gclk));
	jor g1593(.dina(n1660),.dinb(n1656),.dout(n1661),.clk(gclk));
	jor g1594(.dina(n1661),.dinb(w_n167_0[0]),.dout(n1662),.clk(gclk));
	jand g1595(.dina(w_n285_1[2]),.dinb(w_n243_3[0]),.dout(n1663),.clk(gclk));
	jand g1596(.dina(w_n426_1[2]),.dinb(w_n304_2[0]),.dout(n1664),.clk(gclk));
	jand g1597(.dina(n1664),.dinb(n1663),.dout(n1665),.clk(gclk));
	jnot g1598(.din(n1665),.dout(n1666),.clk(gclk));
	jor g1599(.dina(w_n929_0[0]),.dinb(w_n587_0[0]),.dout(n1667),.clk(gclk));
	jor g1600(.dina(n1667),.dinb(w_n866_0[0]),.dout(n1668),.clk(gclk));
	jor g1601(.dina(n1668),.dinb(n1666),.dout(n1669),.clk(gclk));
	jand g1602(.dina(w_n596_0[0]),.dinb(w_n515_1[1]),.dout(n1670),.clk(gclk));
	jand g1603(.dina(n1670),.dinb(w_n665_1[2]),.dout(n1671),.clk(gclk));
	jnot g1604(.din(n1671),.dout(n1672),.clk(gclk));
	jand g1605(.dina(w_n645_1[2]),.dinb(w_n348_1[0]),.dout(n1673),.clk(gclk));
	jnot g1606(.din(w_n1673_0[1]),.dout(n1674),.clk(gclk));
	jor g1607(.dina(w_n389_0[0]),.dinb(w_n378_0[0]),.dout(n1675),.clk(gclk));
	jor g1608(.dina(w_n574_0[0]),.dinb(w_n505_0[0]),.dout(n1676),.clk(gclk));
	jor g1609(.dina(w_n1676_0[1]),.dinb(w_n1675_0[1]),.dout(n1677),.clk(gclk));
	jor g1610(.dina(n1677),.dinb(n1674),.dout(n1678),.clk(gclk));
	jor g1611(.dina(n1678),.dinb(n1672),.dout(n1679),.clk(gclk));
	jor g1612(.dina(w_n1679_0[1]),.dinb(w_n1669_0[1]),.dout(n1680),.clk(gclk));
	jor g1613(.dina(n1680),.dinb(n1662),.dout(n1681),.clk(gclk));
	jor g1614(.dina(n1681),.dinb(w_n1653_0[1]),.dout(n1682),.clk(gclk));
	jand g1615(.dina(w_n1682_5[1]),.dinb(w_n1283_10[2]),.dout(n1683),.clk(gclk));
	jand g1616(.dina(w_n1283_10[1]),.dinb(w_n820_4[0]),.dout(n1684),.clk(gclk));
	jor g1617(.dina(n1684),.dinb(w_n1683_4[2]),.dout(n1685),.clk(gclk));
	jand g1618(.dina(w_n1685_0[1]),.dinb(w_n1640_0[1]),.dout(n1686),.clk(gclk));
	jxor g1619(.dina(w_n1685_0[0]),.dinb(w_n1640_0[0]),.dout(n1687),.clk(gclk));
	jnot g1620(.din(w_n1568_3[0]),.dout(n1688),.clk(gclk));
	jand g1621(.dina(w_n1688_1[1]),.dinb(w_n960_3[0]),.dout(n1689),.clk(gclk));
	jnot g1622(.din(w_n1566_3[0]),.dout(n1690),.clk(gclk));
	jand g1623(.dina(w_n1690_1[1]),.dinb(w_n961_2[2]),.dout(n1691),.clk(gclk));
	jor g1624(.dina(n1691),.dinb(n1689),.dout(n1692),.clk(gclk));
	jand g1625(.dina(w_n1577_3[0]),.dinb(w_n980_3[2]),.dout(n1693),.clk(gclk));
	jand g1626(.dina(w_n1572_3[0]),.dinb(w_n981_2[0]),.dout(n1694),.clk(gclk));
	jor g1627(.dina(n1694),.dinb(n1693),.dout(n1695),.clk(gclk));
	jor g1628(.dina(n1695),.dinb(n1692),.dout(n1696),.clk(gclk));
	jnot g1629(.din(n1696),.dout(n1697),.clk(gclk));
	jand g1630(.dina(w_n1697_0[1]),.dinb(w_n1687_0[1]),.dout(n1698),.clk(gclk));
	jor g1631(.dina(n1698),.dinb(n1686),.dout(n1699),.clk(gclk));
	jand g1632(.dina(w_n804_2[0]),.dinb(w_n55_9[0]),.dout(n1700),.clk(gclk));
	jand g1633(.dina(w_n799_1[2]),.dinb(w_n56_12[1]),.dout(n1701),.clk(gclk));
	jor g1634(.dina(n1701),.dinb(n1700),.dout(n1702),.clk(gclk));
	jand g1635(.dina(w_n1584_4[1]),.dinb(w_n789_2[2]),.dout(n1704),.clk(gclk));
	jor g1636(.dina(n1704),.dinb(n1702),.dout(n1706),.clk(gclk));
	jnot g1637(.din(n1706),.dout(n1707),.clk(gclk));
	jand g1638(.dina(w_n1707_0[1]),.dinb(w_n1699_0[1]),.dout(n1708),.clk(gclk));
	jxor g1639(.dina(w_n1707_0[0]),.dinb(w_n1699_0[0]),.dout(n1709),.clk(gclk));
	jand g1640(.dina(w_n970_0[0]),.dinb(w_n699_12[0]),.dout(n1710),.clk(gclk));
	jand g1641(.dina(w_n1541_0[0]),.dinb(w_n1143_8[0]),.dout(n1711),.clk(gclk));
	jor g1642(.dina(n1711),.dinb(n1710),.dout(n1712),.clk(gclk));
	jand g1643(.dina(w_n1057_3[1]),.dinb(w_n956_2[2]),.dout(n1713),.clk(gclk));
	jand g1644(.dina(w_n1059_4[0]),.dinb(w_n952_2[2]),.dout(n1714),.clk(gclk));
	jor g1645(.dina(n1714),.dinb(n1713),.dout(n1715),.clk(gclk));
	jnot g1646(.din(n1715),.dout(n1716),.clk(gclk));
	jand g1647(.dina(n1716),.dinb(n1712),.dout(n1717),.clk(gclk));
	jand g1648(.dina(w_n1418_3[1]),.dinb(w_n803_6[0]),.dout(n1718),.clk(gclk));
	jand g1649(.dina(w_n1421_3[1]),.dinb(w_n808_11[1]),.dout(n1719),.clk(gclk));
	jor g1650(.dina(n1719),.dinb(n1718),.dout(n1720),.clk(gclk));
	jand g1651(.dina(w_n1533_1[1]),.dinb(w_n708_4[0]),.dout(n1721),.clk(gclk));
	jand g1652(.dina(w_n1535_1[1]),.dinb(w_n794_2[2]),.dout(n1722),.clk(gclk));
	jor g1653(.dina(n1722),.dinb(n1721),.dout(n1723),.clk(gclk));
	jor g1654(.dina(n1723),.dinb(n1720),.dout(n1724),.clk(gclk));
	jnot g1655(.din(n1724),.dout(n1725),.clk(gclk));
	jand g1656(.dina(w_n1725_0[1]),.dinb(w_n1717_0[1]),.dout(n1726),.clk(gclk));
	jxor g1657(.dina(w_n1725_0[0]),.dinb(w_n1717_0[0]),.dout(n1727),.clk(gclk));
	jand g1658(.dina(w_n1037_2[0]),.dinb(w_n337_4[0]),.dout(n1728),.clk(gclk));
	jand g1659(.dina(w_n1034_2[0]),.dinb(w_n1391_4[2]),.dout(n1729),.clk(gclk));
	jor g1660(.dina(n1729),.dinb(n1728),.dout(n1730),.clk(gclk));
	jand g1661(.dina(w_n1347_5[1]),.dinb(w_n1043_2[1]),.dout(n1731),.clk(gclk));
	jand g1662(.dina(w_n1584_4[0]),.dinb(w_n1049_2[1]),.dout(n1732),.clk(gclk));
	jor g1663(.dina(n1732),.dinb(n1731),.dout(n1733),.clk(gclk));
	jor g1664(.dina(n1733),.dinb(n1730),.dout(n1734),.clk(gclk));
	jnot g1665(.din(n1734),.dout(n1735),.clk(gclk));
	jand g1666(.dina(w_n1735_0[1]),.dinb(w_n1727_0[1]),.dout(n1736),.clk(gclk));
	jor g1667(.dina(n1736),.dinb(n1726),.dout(n1737),.clk(gclk));
	jand g1668(.dina(w_n1737_0[1]),.dinb(w_n1709_0[1]),.dout(n1738),.clk(gclk));
	jor g1669(.dina(n1738),.dinb(n1708),.dout(n1739),.clk(gclk));
	jxor g1670(.dina(w_n1638_0[0]),.dinb(w_n1637_0[0]),.dout(n1740),.clk(gclk));
	jand g1671(.dina(w_n1740_0[1]),.dinb(w_n1739_0[1]),.dout(n1741),.clk(gclk));
	jor g1672(.dina(n1741),.dinb(n1639),.dout(n1742),.clk(gclk));
	jxor g1673(.dina(w_n1527_0[0]),.dinb(w_n1526_0[0]),.dout(n1743),.clk(gclk));
	jand g1674(.dina(w_n1743_0[1]),.dinb(w_n1742_0[1]),.dout(n1744),.clk(gclk));
	jxor g1675(.dina(w_n1743_0[0]),.dinb(w_n1742_0[0]),.dout(n1745),.clk(gclk));
	jxor g1676(.dina(w_n1627_0[0]),.dinb(w_n1626_0[0]),.dout(n1746),.clk(gclk));
	jand g1677(.dina(w_n1746_0[1]),.dinb(w_n1745_0[1]),.dout(n1747),.clk(gclk));
	jor g1678(.dina(n1747),.dinb(n1744),.dout(n1748),.clk(gclk));
	jxor g1679(.dina(w_n1632_0[0]),.dinb(w_n1631_0[0]),.dout(n1749),.clk(gclk));
	jand g1680(.dina(w_n1749_0[1]),.dinb(w_n1748_0[1]),.dout(n1750),.clk(gclk));
	jand g1681(.dina(w_n789_2[1]),.dinb(w_n58_4[0]),.dout(n1751),.clk(gclk));
	jand g1682(.dina(w_n1682_5[0]),.dinb(w_n954_21[0]),.dout(n1754),.clk(gclk));
	jand g1683(.dina(w_n1754_0[1]),.dinb(w_n1283_10[0]),.dout(n1755),.clk(gclk));
	jnot g1684(.din(n1755),.dout(n1756),.clk(gclk));
	jand g1685(.dina(w_n1283_9[2]),.dinb(w_n961_2[1]),.dout(n1757),.clk(gclk));
	jor g1686(.dina(n1757),.dinb(w_n1754_0[0]),.dout(n1758),.clk(gclk));
	jor g1687(.dina(n1758),.dinb(w_n1683_4[1]),.dout(n1759),.clk(gclk));
	jand g1688(.dina(n1759),.dinb(n1756),.dout(n1760),.clk(gclk));
	jand g1689(.dina(w_n1760_0[1]),.dinb(w_n335_3[2]),.dout(n1761),.clk(gclk));
	jnot g1690(.din(w_n75_5[0]),.dout(n1762),.clk(gclk));
	jand g1691(.dina(w_n799_1[1]),.dinb(w_n1762_5[1]),.dout(n1763),.clk(gclk));
	jand g1692(.dina(w_n804_1[2]),.dinb(w_n75_4[2]),.dout(n1764),.clk(gclk));
	jor g1693(.dina(n1764),.dinb(n1763),.dout(n1765),.clk(gclk));
	jand g1694(.dina(w_n789_2[0]),.dinb(w_n56_12[0]),.dout(n1766),.clk(gclk));
	jor g1695(.dina(n1766),.dinb(n1765),.dout(n1769),.clk(gclk));
	jnot g1696(.din(n1769),.dout(n1770),.clk(gclk));
	jand g1697(.dina(w_n1770_0[1]),.dinb(w_n1761_0[1]),.dout(n1771),.clk(gclk));
	jand g1698(.dina(w_n1595_0[0]),.dinb(w_n1143_7[2]),.dout(n1772),.clk(gclk));
	jand g1699(.dina(w_n1597_0[0]),.dinb(w_n699_11[2]),.dout(n1773),.clk(gclk));
	jor g1700(.dina(n1773),.dinb(n1772),.dout(n1774),.clk(gclk));
	jand g1701(.dina(w_n971_2[2]),.dinb(w_n337_3[2]),.dout(n1775),.clk(gclk));
	jand g1702(.dina(w_n966_2[2]),.dinb(w_n1391_4[1]),.dout(n1776),.clk(gclk));
	jor g1703(.dina(n1776),.dinb(n1775),.dout(n1777),.clk(gclk));
	jnot g1704(.din(n1777),.dout(n1778),.clk(gclk));
	jand g1705(.dina(n1778),.dinb(n1774),.dout(n1779),.clk(gclk));
	jand g1706(.dina(w_n1584_3[2]),.dinb(w_n1034_1[2]),.dout(n1780),.clk(gclk));
	jand g1707(.dina(w_n1347_5[0]),.dinb(w_n1037_1[2]),.dout(n1781),.clk(gclk));
	jor g1708(.dina(n1781),.dinb(n1780),.dout(n1782),.clk(gclk));
	jand g1709(.dina(w_n1049_2[0]),.dinb(w_n56_11[2]),.dout(n1783),.clk(gclk));
	jand g1710(.dina(w_n1043_2[0]),.dinb(w_n55_8[2]),.dout(n1784),.clk(gclk));
	jor g1711(.dina(n1784),.dinb(n1783),.dout(n1785),.clk(gclk));
	jor g1712(.dina(n1785),.dinb(n1782),.dout(n1786),.clk(gclk));
	jnot g1713(.din(n1786),.dout(n1787),.clk(gclk));
	jand g1714(.dina(w_n1787_0[1]),.dinb(w_n1779_0[1]),.dout(n1788),.clk(gclk));
	jxor g1715(.dina(w_n1787_0[0]),.dinb(w_n1779_0[0]),.dout(n1789),.clk(gclk));
	jand g1716(.dina(w_n1411_1[2]),.dinb(w_n1057_3[0]),.dout(n1790),.clk(gclk));
	jand g1717(.dina(w_n1414_1[2]),.dinb(w_n1059_3[2]),.dout(n1791),.clk(gclk));
	jor g1718(.dina(n1791),.dinb(n1790),.dout(n1792),.clk(gclk));
	jand g1719(.dina(w_n1418_3[0]),.dinb(w_n708_3[2]),.dout(n1793),.clk(gclk));
	jand g1720(.dina(w_n1421_3[0]),.dinb(w_n794_2[1]),.dout(n1794),.clk(gclk));
	jor g1721(.dina(n1794),.dinb(n1793),.dout(n1795),.clk(gclk));
	jnot g1722(.din(n1795),.dout(n1796),.clk(gclk));
	jand g1723(.dina(n1796),.dinb(n1792),.dout(n1797),.clk(gclk));
	jand g1724(.dina(w_n1797_0[1]),.dinb(w_n1789_0[1]),.dout(n1798),.clk(gclk));
	jor g1725(.dina(n1798),.dinb(n1788),.dout(n1799),.clk(gclk));
	jxor g1726(.dina(w_n1770_0[0]),.dinb(w_n1761_0[0]),.dout(n1800),.clk(gclk));
	jand g1727(.dina(w_n1800_0[1]),.dinb(w_n1799_0[1]),.dout(n1801),.clk(gclk));
	jor g1728(.dina(n1801),.dinb(n1771),.dout(n1802),.clk(gclk));
	jxor g1729(.dina(w_n1581_0[0]),.dinb(w_n1565_0[0]),.dout(n1803),.clk(gclk));
	jand g1730(.dina(w_n1803_0[1]),.dinb(w_n1802_0[1]),.dout(n1804),.clk(gclk));
	jxor g1731(.dina(w_n1803_0[0]),.dinb(w_n1802_0[0]),.dout(n1805),.clk(gclk));
	jxor g1732(.dina(w_n1622_0[0]),.dinb(w_n1614_0[0]),.dout(n1806),.clk(gclk));
	jand g1733(.dina(w_n1806_0[1]),.dinb(w_n1805_0[1]),.dout(n1807),.clk(gclk));
	jor g1734(.dina(n1807),.dinb(n1804),.dout(n1808),.clk(gclk));
	jxor g1735(.dina(w_n1624_0[0]),.dinb(w_n1594_0[0]),.dout(n1809),.clk(gclk));
	jand g1736(.dina(w_n1809_0[1]),.dinb(w_n1808_0[1]),.dout(n1810),.clk(gclk));
	jxor g1737(.dina(w_n1809_0[0]),.dinb(w_n1808_0[0]),.dout(n1811),.clk(gclk));
	jxor g1738(.dina(w_n1740_0[0]),.dinb(w_n1739_0[0]),.dout(n1812),.clk(gclk));
	jand g1739(.dina(w_n1812_0[1]),.dinb(w_n1811_0[1]),.dout(n1813),.clk(gclk));
	jor g1740(.dina(n1813),.dinb(n1810),.dout(n1814),.clk(gclk));
	jxor g1741(.dina(w_n1746_0[0]),.dinb(w_n1745_0[0]),.dout(n1815),.clk(gclk));
	jand g1742(.dina(w_n1815_0[1]),.dinb(w_n1814_0[1]),.dout(n1816),.clk(gclk));
	jand g1743(.dina(w_n804_1[1]),.dinb(w_n58_3[2]),.dout(n1817),.clk(gclk));
	jand g1744(.dina(w_n799_1[0]),.dinb(w_n59_3[0]),.dout(n1818),.clk(gclk));
	jor g1745(.dina(n1818),.dinb(n1817),.dout(n1819),.clk(gclk));
	jand g1746(.dina(w_n789_1[2]),.dinb(w_n1762_5[0]),.dout(n1821),.clk(gclk));
	jor g1747(.dina(n1821),.dinb(n1819),.dout(n1823),.clk(gclk));
	jnot g1748(.din(n1823),.dout(n1824),.clk(gclk));
	jand g1749(.dina(w_n1566_2[2]),.dinb(w_n981_1[2]),.dout(n1825),.clk(gclk));
	jand g1750(.dina(w_n1568_2[2]),.dinb(w_n980_3[1]),.dout(n1826),.clk(gclk));
	jor g1751(.dina(n1826),.dinb(n1825),.dout(n1827),.clk(gclk));
	jand g1752(.dina(w_n1572_2[2]),.dinb(w_n808_11[0]),.dout(n1828),.clk(gclk));
	jand g1753(.dina(w_n1577_2[2]),.dinb(w_n803_5[2]),.dout(n1829),.clk(gclk));
	jor g1754(.dina(n1829),.dinb(n1828),.dout(n1830),.clk(gclk));
	jnot g1755(.din(n1830),.dout(n1831),.clk(gclk));
	jand g1756(.dina(n1831),.dinb(n1827),.dout(n1832),.clk(gclk));
	jand g1757(.dina(w_n1832_0[1]),.dinb(w_n1824_0[1]),.dout(n1833),.clk(gclk));
	jxor g1758(.dina(w_n1760_0[0]),.dinb(w_n335_3[1]),.dout(n1834),.clk(gclk));
	jxor g1759(.dina(w_n1832_0[0]),.dinb(w_n1824_0[0]),.dout(n1835),.clk(gclk));
	jand g1760(.dina(w_n1835_0[1]),.dinb(w_n1834_0[1]),.dout(n1836),.clk(gclk));
	jor g1761(.dina(n1836),.dinb(n1833),.dout(n1837),.clk(gclk));
	jxor g1762(.dina(w_n1697_0[0]),.dinb(w_n1687_0[0]),.dout(n1838),.clk(gclk));
	jand g1763(.dina(w_n1838_0[1]),.dinb(w_n1837_0[1]),.dout(n1839),.clk(gclk));
	jxor g1764(.dina(w_n1838_0[0]),.dinb(w_n1837_0[0]),.dout(n1840),.clk(gclk));
	jxor g1765(.dina(w_n1735_0[0]),.dinb(w_n1727_0[0]),.dout(n1841),.clk(gclk));
	jand g1766(.dina(w_n1841_0[1]),.dinb(w_n1840_0[1]),.dout(n1842),.clk(gclk));
	jor g1767(.dina(n1842),.dinb(n1839),.dout(n1843),.clk(gclk));
	jxor g1768(.dina(w_n1737_0[0]),.dinb(w_n1709_0[0]),.dout(n1844),.clk(gclk));
	jand g1769(.dina(w_n1844_0[1]),.dinb(w_n1843_0[1]),.dout(n1845),.clk(gclk));
	jxor g1770(.dina(w_n1844_0[0]),.dinb(w_n1843_0[0]),.dout(n1846),.clk(gclk));
	jxor g1771(.dina(w_n1806_0[0]),.dinb(w_n1805_0[0]),.dout(n1847),.clk(gclk));
	jand g1772(.dina(w_n1847_0[1]),.dinb(w_n1846_0[1]),.dout(n1848),.clk(gclk));
	jor g1773(.dina(n1848),.dinb(n1845),.dout(n1849),.clk(gclk));
	jxor g1774(.dina(w_n1812_0[0]),.dinb(w_n1811_0[0]),.dout(n1850),.clk(gclk));
	jand g1775(.dina(w_n1850_0[1]),.dinb(w_n1849_0[1]),.dout(n1851),.clk(gclk));
	jand g1776(.dina(w_n1418_2[2]),.dinb(w_n1057_2[2]),.dout(n1852),.clk(gclk));
	jand g1777(.dina(w_n1421_2[2]),.dinb(w_n1059_3[1]),.dout(n1853),.clk(gclk));
	jor g1778(.dina(n1853),.dinb(n1852),.dout(n1854),.clk(gclk));
	jand g1779(.dina(w_n1533_1[0]),.dinb(w_n699_11[1]),.dout(n1855),.clk(gclk));
	jand g1780(.dina(w_n1535_1[0]),.dinb(w_n1143_7[1]),.dout(n1856),.clk(gclk));
	jor g1781(.dina(n1856),.dinb(n1855),.dout(n1857),.clk(gclk));
	jor g1782(.dina(n1857),.dinb(n1854),.dout(n1858),.clk(gclk));
	jnot g1783(.din(w_n1858_0[1]),.dout(n1859),.clk(gclk));
	jand g1784(.dina(w_n956_2[1]),.dinb(w_n337_3[1]),.dout(n1860),.clk(gclk));
	jand g1785(.dina(w_n952_2[1]),.dinb(w_n1391_4[0]),.dout(n1861),.clk(gclk));
	jor g1786(.dina(n1861),.dinb(n1860),.dout(n1862),.clk(gclk));
	jand g1787(.dina(w_n1347_4[2]),.dinb(w_n971_2[1]),.dout(n1863),.clk(gclk));
	jand g1788(.dina(w_n1584_3[1]),.dinb(w_n966_2[1]),.dout(n1864),.clk(gclk));
	jor g1789(.dina(n1864),.dinb(n1863),.dout(n1865),.clk(gclk));
	jor g1790(.dina(n1865),.dinb(n1862),.dout(n1866),.clk(gclk));
	jnot g1791(.din(w_n1866_0[1]),.dout(n1867),.clk(gclk));
	jand g1792(.dina(n1867),.dinb(n1859),.dout(n1868),.clk(gclk));
	jand g1793(.dina(w_n1033_0[1]),.dinb(w_n58_3[1]),.dout(n1869),.clk(gclk));
	jnot g1794(.din(w_n1869_0[2]),.dout(n1870),.clk(gclk));
	jand g1795(.dina(n1870),.dinb(w_n1047_0[2]),.dout(n1871),.clk(gclk));
	jand g1796(.dina(w_n1682_4[2]),.dinb(w_n980_3[0]),.dout(n1872),.clk(gclk));
	jand g1797(.dina(w_n1872_0[1]),.dinb(w_n1283_9[1]),.dout(n1873),.clk(gclk));
	jnot g1798(.din(n1873),.dout(n1874),.clk(gclk));
	jand g1799(.dina(w_n1283_9[0]),.dinb(w_n808_10[2]),.dout(n1875),.clk(gclk));
	jor g1800(.dina(n1875),.dinb(w_n1872_0[0]),.dout(n1876),.clk(gclk));
	jor g1801(.dina(n1876),.dinb(w_n1683_4[0]),.dout(n1877),.clk(gclk));
	jand g1802(.dina(n1877),.dinb(n1874),.dout(n1878),.clk(gclk));
	jand g1803(.dina(w_n1878_0[1]),.dinb(w_n1871_0[1]),.dout(n1879),.clk(gclk));
	jxor g1804(.dina(w_n1866_0[0]),.dinb(w_n1858_0[0]),.dout(n1880),.clk(gclk));
	jand g1805(.dina(w_n1880_0[1]),.dinb(w_n1879_0[1]),.dout(n1881),.clk(gclk));
	jor g1806(.dina(n1881),.dinb(n1868),.dout(n1882),.clk(gclk));
	jand g1807(.dina(w_n1682_4[1]),.dinb(w_n960_2[2]),.dout(n1883),.clk(gclk));
	jand g1808(.dina(w_n1883_0[1]),.dinb(w_n1283_8[2]),.dout(n1884),.clk(gclk));
	jnot g1809(.din(n1884),.dout(n1885),.clk(gclk));
	jand g1810(.dina(w_n1283_8[1]),.dinb(w_n981_1[1]),.dout(n1886),.clk(gclk));
	jor g1811(.dina(n1886),.dinb(w_n1883_0[0]),.dout(n1887),.clk(gclk));
	jor g1812(.dina(n1887),.dinb(w_n1683_3[2]),.dout(n1888),.clk(gclk));
	jand g1813(.dina(n1888),.dinb(n1885),.dout(n1889),.clk(gclk));
	jand g1814(.dina(w_n1688_1[0]),.dinb(w_n803_5[1]),.dout(n1890),.clk(gclk));
	jand g1815(.dina(w_n1690_1[0]),.dinb(w_n808_10[1]),.dout(n1891),.clk(gclk));
	jor g1816(.dina(n1891),.dinb(n1890),.dout(n1892),.clk(gclk));
	jand g1817(.dina(w_n1577_2[1]),.dinb(w_n708_3[1]),.dout(n1893),.clk(gclk));
	jand g1818(.dina(w_n1572_2[1]),.dinb(w_n794_2[0]),.dout(n1894),.clk(gclk));
	jor g1819(.dina(n1894),.dinb(n1893),.dout(n1895),.clk(gclk));
	jor g1820(.dina(n1895),.dinb(n1892),.dout(n1896),.clk(gclk));
	jnot g1821(.din(n1896),.dout(n1897),.clk(gclk));
	jand g1822(.dina(w_n1897_0[1]),.dinb(w_n1889_0[1]),.dout(n1898),.clk(gclk));
	jxor g1823(.dina(w_n1897_0[0]),.dinb(w_n1889_0[0]),.dout(n1899),.clk(gclk));
	jand g1824(.dina(w_n1037_1[1]),.dinb(w_n55_8[1]),.dout(n1900),.clk(gclk));
	jand g1825(.dina(w_n1034_1[1]),.dinb(w_n56_11[1]),.dout(n1901),.clk(gclk));
	jor g1826(.dina(n1901),.dinb(n1900),.dout(n1902),.clk(gclk));
	jand g1827(.dina(w_n1043_1[2]),.dinb(w_n75_4[1]),.dout(n1903),.clk(gclk));
	jand g1828(.dina(w_n1049_1[2]),.dinb(w_n1762_4[2]),.dout(n1904),.clk(gclk));
	jor g1829(.dina(n1904),.dinb(n1903),.dout(n1905),.clk(gclk));
	jor g1830(.dina(n1905),.dinb(n1902),.dout(n1906),.clk(gclk));
	jnot g1831(.din(n1906),.dout(n1907),.clk(gclk));
	jand g1832(.dina(w_n1907_0[1]),.dinb(w_n1899_0[1]),.dout(n1908),.clk(gclk));
	jor g1833(.dina(n1908),.dinb(n1898),.dout(n1909),.clk(gclk));
	jand g1834(.dina(w_n1909_0[1]),.dinb(w_n1882_0[1]),.dout(n1910),.clk(gclk));
	jxor g1835(.dina(w_n1909_0[0]),.dinb(w_n1882_0[0]),.dout(n1911),.clk(gclk));
	jxor g1836(.dina(w_n1797_0[0]),.dinb(w_n1789_0[0]),.dout(n1912),.clk(gclk));
	jand g1837(.dina(w_n1912_0[1]),.dinb(w_n1911_0[1]),.dout(n1913),.clk(gclk));
	jor g1838(.dina(n1913),.dinb(n1910),.dout(n1914),.clk(gclk));
	jxor g1839(.dina(w_n1800_0[0]),.dinb(w_n1799_0[0]),.dout(n1915),.clk(gclk));
	jand g1840(.dina(w_n1915_0[1]),.dinb(w_n1914_0[1]),.dout(n1916),.clk(gclk));
	jxor g1841(.dina(w_n1915_0[0]),.dinb(w_n1914_0[0]),.dout(n1917),.clk(gclk));
	jxor g1842(.dina(w_n1841_0[0]),.dinb(w_n1840_0[0]),.dout(n1918),.clk(gclk));
	jand g1843(.dina(w_n1918_0[1]),.dinb(w_n1917_0[1]),.dout(n1919),.clk(gclk));
	jor g1844(.dina(n1919),.dinb(n1916),.dout(n1920),.clk(gclk));
	jxor g1845(.dina(w_n1847_0[0]),.dinb(w_n1846_0[0]),.dout(n1921),.clk(gclk));
	jand g1846(.dina(w_n1921_0[1]),.dinb(w_n1920_0[1]),.dout(n1922),.clk(gclk));
	jand g1847(.dina(w_n1566_2[1]),.dinb(w_n794_1[2]),.dout(n1923),.clk(gclk));
	jand g1848(.dina(w_n1568_2[1]),.dinb(w_n708_3[0]),.dout(n1924),.clk(gclk));
	jor g1849(.dina(n1924),.dinb(n1923),.dout(n1925),.clk(gclk));
	jand g1850(.dina(w_n1572_2[0]),.dinb(w_n1059_3[0]),.dout(n1926),.clk(gclk));
	jand g1851(.dina(w_n1577_2[0]),.dinb(w_n1057_2[1]),.dout(n1927),.clk(gclk));
	jor g1852(.dina(n1927),.dinb(n1926),.dout(n1928),.clk(gclk));
	jnot g1853(.din(n1928),.dout(n1929),.clk(gclk));
	jand g1854(.dina(n1929),.dinb(n1925),.dout(n1930),.clk(gclk));
	jand g1855(.dina(w_n1584_3[0]),.dinb(w_n952_2[0]),.dout(n1931),.clk(gclk));
	jand g1856(.dina(w_n1347_4[1]),.dinb(w_n956_2[0]),.dout(n1932),.clk(gclk));
	jor g1857(.dina(n1932),.dinb(n1931),.dout(n1933),.clk(gclk));
	jand g1858(.dina(w_n966_2[0]),.dinb(w_n56_11[0]),.dout(n1934),.clk(gclk));
	jand g1859(.dina(w_n971_2[0]),.dinb(w_n55_8[0]),.dout(n1935),.clk(gclk));
	jor g1860(.dina(n1935),.dinb(n1934),.dout(n1936),.clk(gclk));
	jor g1861(.dina(n1936),.dinb(n1933),.dout(n1937),.clk(gclk));
	jnot g1862(.din(n1937),.dout(n1938),.clk(gclk));
	jand g1863(.dina(w_n1938_0[1]),.dinb(w_n1930_0[1]),.dout(n1939),.clk(gclk));
	jxor g1864(.dina(w_n1938_0[0]),.dinb(w_n1930_0[0]),.dout(n1940),.clk(gclk));
	jand g1865(.dina(w_n1411_1[1]),.dinb(w_n337_3[0]),.dout(n1941),.clk(gclk));
	jand g1866(.dina(w_n1414_1[1]),.dinb(w_n1391_3[2]),.dout(n1942),.clk(gclk));
	jor g1867(.dina(n1942),.dinb(n1941),.dout(n1943),.clk(gclk));
	jand g1868(.dina(w_n1418_2[1]),.dinb(w_n699_11[0]),.dout(n1944),.clk(gclk));
	jand g1869(.dina(w_n1421_2[1]),.dinb(w_n1143_7[0]),.dout(n1945),.clk(gclk));
	jor g1870(.dina(n1945),.dinb(n1944),.dout(n1946),.clk(gclk));
	jnot g1871(.din(n1946),.dout(n1947),.clk(gclk));
	jand g1872(.dina(n1947),.dinb(n1943),.dout(n1948),.clk(gclk));
	jand g1873(.dina(w_n1948_0[1]),.dinb(w_n1940_0[1]),.dout(n1949),.clk(gclk));
	jor g1874(.dina(n1949),.dinb(n1939),.dout(n1950),.clk(gclk));
	jand g1875(.dina(w_n1950_0[1]),.dinb(w_n1751_0[1]),.dout(n1951),.clk(gclk));
	jxor g1876(.dina(w_n1880_0[0]),.dinb(w_n1879_0[0]),.dout(n1952),.clk(gclk));
	jxor g1877(.dina(w_n1950_0[0]),.dinb(w_n1751_0[0]),.dout(n1953),.clk(gclk));
	jand g1878(.dina(w_n1953_0[1]),.dinb(w_n1952_0[1]),.dout(n1954),.clk(gclk));
	jor g1879(.dina(n1954),.dinb(n1951),.dout(n1955),.clk(gclk));
	jxor g1880(.dina(w_n1835_0[0]),.dinb(w_n1834_0[0]),.dout(n1956),.clk(gclk));
	jand g1881(.dina(w_n1956_0[1]),.dinb(w_n1955_0[1]),.dout(n1957),.clk(gclk));
	jxor g1882(.dina(w_n1956_0[0]),.dinb(w_n1955_0[0]),.dout(n1958),.clk(gclk));
	jxor g1883(.dina(w_n1912_0[0]),.dinb(w_n1911_0[0]),.dout(n1959),.clk(gclk));
	jand g1884(.dina(w_n1959_0[1]),.dinb(w_n1958_0[1]),.dout(n1960),.clk(gclk));
	jor g1885(.dina(n1960),.dinb(n1957),.dout(n1961),.clk(gclk));
	jxor g1886(.dina(w_n1918_0[0]),.dinb(w_n1917_0[0]),.dout(n1962),.clk(gclk));
	jand g1887(.dina(w_n1962_0[1]),.dinb(w_n1961_0[1]),.dout(n1963),.clk(gclk));
	jxor g1888(.dina(w_n1962_0[0]),.dinb(w_n1961_0[0]),.dout(n1964),.clk(gclk));
	jxor g1889(.dina(w_n1878_0[0]),.dinb(w_n1871_0[0]),.dout(n1965),.clk(gclk));
	jand g1890(.dina(w_n1034_1[0]),.dinb(w_n1762_4[1]),.dout(n1966),.clk(gclk));
	jand g1891(.dina(w_n1037_1[0]),.dinb(w_n75_4[0]),.dout(n1967),.clk(gclk));
	jor g1892(.dina(n1967),.dinb(n1966),.dout(n1968),.clk(gclk));
	jand g1893(.dina(w_n1049_1[1]),.dinb(w_n59_2[2]),.dout(n1969),.clk(gclk));
	jand g1894(.dina(w_n1043_1[1]),.dinb(w_n58_3[0]),.dout(n1970),.clk(gclk));
	jor g1895(.dina(n1970),.dinb(n1969),.dout(n1971),.clk(gclk));
	jor g1896(.dina(n1971),.dinb(n1968),.dout(n1972),.clk(gclk));
	jnot g1897(.din(n1972),.dout(n1973),.clk(gclk));
	jand g1898(.dina(w_n1973_0[1]),.dinb(w_n1965_0[1]),.dout(n1974),.clk(gclk));
	jand g1899(.dina(w_n1682_4[0]),.dinb(w_n803_5[0]),.dout(n1975),.clk(gclk));
	jand g1900(.dina(w_n1975_0[1]),.dinb(w_n1283_8[0]),.dout(n1976),.clk(gclk));
	jnot g1901(.din(n1976),.dout(n1977),.clk(gclk));
	jand g1902(.dina(w_n1283_7[2]),.dinb(w_n794_1[1]),.dout(n1978),.clk(gclk));
	jor g1903(.dina(n1978),.dinb(w_n1975_0[0]),.dout(n1979),.clk(gclk));
	jor g1904(.dina(n1979),.dinb(w_n1683_3[1]),.dout(n1980),.clk(gclk));
	jand g1905(.dina(n1980),.dinb(n1977),.dout(n1981),.clk(gclk));
	jand g1906(.dina(w_n1688_0[2]),.dinb(w_n1057_2[0]),.dout(n1982),.clk(gclk));
	jand g1907(.dina(w_n1690_0[2]),.dinb(w_n1059_2[2]),.dout(n1983),.clk(gclk));
	jor g1908(.dina(n1983),.dinb(n1982),.dout(n1984),.clk(gclk));
	jand g1909(.dina(w_n1577_1[2]),.dinb(w_n699_10[2]),.dout(n1985),.clk(gclk));
	jand g1910(.dina(w_n1572_1[2]),.dinb(w_n1143_6[2]),.dout(n1986),.clk(gclk));
	jor g1911(.dina(n1986),.dinb(n1985),.dout(n1987),.clk(gclk));
	jor g1912(.dina(n1987),.dinb(n1984),.dout(n1988),.clk(gclk));
	jnot g1913(.din(n1988),.dout(n1989),.clk(gclk));
	jand g1914(.dina(w_n1989_0[1]),.dinb(w_n1981_0[1]),.dout(n1990),.clk(gclk));
	jxor g1915(.dina(w_n1989_0[0]),.dinb(w_n1981_0[0]),.dout(n1991),.clk(gclk));
	jand g1916(.dina(w_n1418_2[0]),.dinb(w_n337_2[2]),.dout(n1992),.clk(gclk));
	jand g1917(.dina(w_n1421_2[0]),.dinb(w_n1391_3[1]),.dout(n1993),.clk(gclk));
	jor g1918(.dina(n1993),.dinb(n1992),.dout(n1994),.clk(gclk));
	jand g1919(.dina(w_n1533_0[2]),.dinb(w_n1347_4[0]),.dout(n1995),.clk(gclk));
	jand g1920(.dina(w_n1535_0[2]),.dinb(w_n1584_2[2]),.dout(n1996),.clk(gclk));
	jor g1921(.dina(n1996),.dinb(n1995),.dout(n1997),.clk(gclk));
	jor g1922(.dina(n1997),.dinb(n1994),.dout(n1998),.clk(gclk));
	jnot g1923(.din(n1998),.dout(n1999),.clk(gclk));
	jand g1924(.dina(w_n1999_0[1]),.dinb(w_n1991_0[1]),.dout(n2000),.clk(gclk));
	jor g1925(.dina(n2000),.dinb(n1990),.dout(n2001),.clk(gclk));
	jxor g1926(.dina(w_n1973_0[0]),.dinb(w_n1965_0[0]),.dout(n2002),.clk(gclk));
	jand g1927(.dina(w_n2002_0[1]),.dinb(w_n2001_0[1]),.dout(n2003),.clk(gclk));
	jor g1928(.dina(n2003),.dinb(n1974),.dout(n2004),.clk(gclk));
	jxor g1929(.dina(w_n1907_0[0]),.dinb(w_n1899_0[0]),.dout(n2005),.clk(gclk));
	jand g1930(.dina(w_n2005_0[1]),.dinb(w_n2004_0[1]),.dout(n2006),.clk(gclk));
	jxor g1931(.dina(w_n1953_0[0]),.dinb(w_n1952_0[0]),.dout(n2007),.clk(gclk));
	jxor g1932(.dina(w_n2005_0[0]),.dinb(w_n2004_0[0]),.dout(n2008),.clk(gclk));
	jand g1933(.dina(w_n2008_0[1]),.dinb(w_n2007_0[1]),.dout(n2009),.clk(gclk));
	jor g1934(.dina(n2009),.dinb(n2006),.dout(n2010),.clk(gclk));
	jand g1935(.dina(w_n951_0[1]),.dinb(w_n58_2[2]),.dout(n2011),.clk(gclk));
	jnot g1936(.din(w_n2011_0[2]),.dout(n2012),.clk(gclk));
	jand g1937(.dina(n2012),.dinb(w_n964_0[1]),.dout(n2013),.clk(gclk));
	jand g1938(.dina(w_n1682_3[2]),.dinb(w_n708_2[2]),.dout(n2014),.clk(gclk));
	jand g1939(.dina(w_n2014_0[1]),.dinb(w_n1283_7[1]),.dout(n2015),.clk(gclk));
	jnot g1940(.din(n2015),.dout(n2016),.clk(gclk));
	jand g1941(.dina(w_n1283_7[0]),.dinb(w_n1059_2[1]),.dout(n2017),.clk(gclk));
	jor g1942(.dina(n2017),.dinb(w_n2014_0[0]),.dout(n2018),.clk(gclk));
	jor g1943(.dina(n2018),.dinb(w_n1683_3[0]),.dout(n2019),.clk(gclk));
	jand g1944(.dina(n2019),.dinb(n2016),.dout(n2020),.clk(gclk));
	jand g1945(.dina(w_n2020_0[1]),.dinb(w_n2013_0[1]),.dout(n2021),.clk(gclk));
	jand g1946(.dina(w_n956_1[2]),.dinb(w_n55_7[2]),.dout(n2022),.clk(gclk));
	jand g1947(.dina(w_n952_1[2]),.dinb(w_n56_10[2]),.dout(n2023),.clk(gclk));
	jor g1948(.dina(n2023),.dinb(n2022),.dout(n2024),.clk(gclk));
	jand g1949(.dina(w_n971_1[2]),.dinb(w_n75_3[2]),.dout(n2025),.clk(gclk));
	jand g1950(.dina(w_n966_1[2]),.dinb(w_n1762_4[0]),.dout(n2026),.clk(gclk));
	jor g1951(.dina(n2026),.dinb(n2025),.dout(n2027),.clk(gclk));
	jor g1952(.dina(n2027),.dinb(n2024),.dout(n2028),.clk(gclk));
	jnot g1953(.din(n2028),.dout(n2029),.clk(gclk));
	jand g1954(.dina(w_n2029_0[1]),.dinb(w_n2021_0[1]),.dout(n2030),.clk(gclk));
	jxor g1955(.dina(w_n2029_0[0]),.dinb(w_n2021_0[0]),.dout(n2031),.clk(gclk));
	jand g1956(.dina(w_n2031_0[1]),.dinb(w_n1869_0[1]),.dout(n2032),.clk(gclk));
	jor g1957(.dina(n2032),.dinb(n2030),.dout(n2033),.clk(gclk));
	jxor g1958(.dina(w_n1948_0[0]),.dinb(w_n1940_0[0]),.dout(n2034),.clk(gclk));
	jand g1959(.dina(w_n2034_0[1]),.dinb(w_n2033_0[1]),.dout(n2035),.clk(gclk));
	jxor g1960(.dina(w_n2034_0[0]),.dinb(w_n2033_0[0]),.dout(n2036),.clk(gclk));
	jxor g1961(.dina(w_n2002_0[0]),.dinb(w_n2001_0[0]),.dout(n2037),.clk(gclk));
	jand g1962(.dina(w_n2037_0[1]),.dinb(w_n2036_0[1]),.dout(n2038),.clk(gclk));
	jor g1963(.dina(n2038),.dinb(n2035),.dout(n2039),.clk(gclk));
	jand g1964(.dina(w_n1566_2[0]),.dinb(w_n1143_6[1]),.dout(n2040),.clk(gclk));
	jand g1965(.dina(w_n1568_2[0]),.dinb(w_n699_10[1]),.dout(n2041),.clk(gclk));
	jor g1966(.dina(n2041),.dinb(n2040),.dout(n2042),.clk(gclk));
	jand g1967(.dina(w_n1572_1[1]),.dinb(w_n1391_3[0]),.dout(n2043),.clk(gclk));
	jand g1968(.dina(w_n1577_1[1]),.dinb(w_n337_2[1]),.dout(n2044),.clk(gclk));
	jor g1969(.dina(n2044),.dinb(n2043),.dout(n2045),.clk(gclk));
	jnot g1970(.din(n2045),.dout(n2046),.clk(gclk));
	jand g1971(.dina(n2046),.dinb(n2042),.dout(n2047),.clk(gclk));
	jand g1972(.dina(w_n1411_1[0]),.dinb(w_n55_7[1]),.dout(n2048),.clk(gclk));
	jand g1973(.dina(w_n1414_1[0]),.dinb(w_n56_10[1]),.dout(n2049),.clk(gclk));
	jor g1974(.dina(n2049),.dinb(n2048),.dout(n2050),.clk(gclk));
	jand g1975(.dina(w_n1418_1[2]),.dinb(w_n1347_3[2]),.dout(n2051),.clk(gclk));
	jand g1976(.dina(w_n1421_1[2]),.dinb(w_n1584_2[1]),.dout(n2052),.clk(gclk));
	jor g1977(.dina(n2052),.dinb(n2051),.dout(n2053),.clk(gclk));
	jnot g1978(.din(n2053),.dout(n2054),.clk(gclk));
	jand g1979(.dina(n2054),.dinb(n2050),.dout(n2055),.clk(gclk));
	jand g1980(.dina(w_n2055_0[1]),.dinb(w_n2047_0[1]),.dout(n2056),.clk(gclk));
	jxor g1981(.dina(w_n2055_0[0]),.dinb(w_n2047_0[0]),.dout(n2057),.clk(gclk));
	jand g1982(.dina(w_n952_1[1]),.dinb(w_n1762_3[2]),.dout(n2058),.clk(gclk));
	jand g1983(.dina(w_n956_1[1]),.dinb(w_n75_3[1]),.dout(n2059),.clk(gclk));
	jor g1984(.dina(n2059),.dinb(n2058),.dout(n2060),.clk(gclk));
	jand g1985(.dina(w_n966_1[1]),.dinb(w_n59_2[1]),.dout(n2061),.clk(gclk));
	jand g1986(.dina(w_n971_1[1]),.dinb(w_n58_2[1]),.dout(n2062),.clk(gclk));
	jor g1987(.dina(n2062),.dinb(n2061),.dout(n2063),.clk(gclk));
	jor g1988(.dina(n2063),.dinb(n2060),.dout(n2064),.clk(gclk));
	jnot g1989(.din(n2064),.dout(n2065),.clk(gclk));
	jand g1990(.dina(w_n2065_0[1]),.dinb(w_n2057_0[1]),.dout(n2066),.clk(gclk));
	jor g1991(.dina(n2066),.dinb(n2056),.dout(n2067),.clk(gclk));
	jxor g1992(.dina(w_n1999_0[0]),.dinb(w_n1991_0[0]),.dout(n2068),.clk(gclk));
	jand g1993(.dina(w_n2068_0[1]),.dinb(w_n2067_0[1]),.dout(n2069),.clk(gclk));
	jxor g1994(.dina(w_n2031_0[0]),.dinb(w_n1869_0[0]),.dout(n2070),.clk(gclk));
	jxor g1995(.dina(w_n2068_0[0]),.dinb(w_n2067_0[0]),.dout(n2071),.clk(gclk));
	jand g1996(.dina(w_n2071_0[1]),.dinb(w_n2070_0[1]),.dout(n2072),.clk(gclk));
	jor g1997(.dina(n2072),.dinb(n2069),.dout(n2073),.clk(gclk));
	jxor g1998(.dina(w_n2020_0[0]),.dinb(w_n2013_0[0]),.dout(n2074),.clk(gclk));
	jand g1999(.dina(w_n1682_3[1]),.dinb(w_n1057_1[2]),.dout(n2075),.clk(gclk));
	jand g2000(.dina(w_n2075_0[1]),.dinb(w_n1283_6[2]),.dout(n2076),.clk(gclk));
	jnot g2001(.din(n2076),.dout(n2077),.clk(gclk));
	jand g2002(.dina(w_n1283_6[1]),.dinb(w_n1143_6[0]),.dout(n2078),.clk(gclk));
	jor g2003(.dina(n2078),.dinb(w_n2075_0[0]),.dout(n2079),.clk(gclk));
	jor g2004(.dina(n2079),.dinb(w_n1683_2[2]),.dout(n2080),.clk(gclk));
	jand g2005(.dina(n2080),.dinb(n2077),.dout(n2081),.clk(gclk));
	jand g2006(.dina(w_n1688_0[1]),.dinb(w_n337_2[0]),.dout(n2082),.clk(gclk));
	jand g2007(.dina(w_n1690_0[1]),.dinb(w_n1391_2[2]),.dout(n2083),.clk(gclk));
	jor g2008(.dina(n2083),.dinb(n2082),.dout(n2084),.clk(gclk));
	jand g2009(.dina(w_n1577_1[0]),.dinb(w_n1347_3[1]),.dout(n2085),.clk(gclk));
	jand g2010(.dina(w_n1572_1[0]),.dinb(w_n1584_2[0]),.dout(n2086),.clk(gclk));
	jor g2011(.dina(n2086),.dinb(n2085),.dout(n2087),.clk(gclk));
	jor g2012(.dina(n2087),.dinb(n2084),.dout(n2088),.clk(gclk));
	jnot g2013(.din(n2088),.dout(n2089),.clk(gclk));
	jand g2014(.dina(w_n2089_0[1]),.dinb(w_n2081_0[1]),.dout(n2090),.clk(gclk));
	jxor g2015(.dina(w_n2089_0[0]),.dinb(w_n2081_0[0]),.dout(n2091),.clk(gclk));
	jand g2016(.dina(w_n1418_1[1]),.dinb(w_n55_7[0]),.dout(n2092),.clk(gclk));
	jand g2017(.dina(w_n1421_1[1]),.dinb(w_n56_10[0]),.dout(n2093),.clk(gclk));
	jor g2018(.dina(n2093),.dinb(n2092),.dout(n2094),.clk(gclk));
	jand g2019(.dina(w_n1533_0[1]),.dinb(w_n75_3[0]),.dout(n2095),.clk(gclk));
	jand g2020(.dina(w_n1535_0[1]),.dinb(w_n1762_3[1]),.dout(n2096),.clk(gclk));
	jor g2021(.dina(n2096),.dinb(n2095),.dout(n2097),.clk(gclk));
	jor g2022(.dina(n2097),.dinb(n2094),.dout(n2098),.clk(gclk));
	jnot g2023(.din(n2098),.dout(n2099),.clk(gclk));
	jand g2024(.dina(w_n2099_0[1]),.dinb(w_n2091_0[1]),.dout(n2100),.clk(gclk));
	jor g2025(.dina(n2100),.dinb(n2090),.dout(n2101),.clk(gclk));
	jand g2026(.dina(w_n2101_0[1]),.dinb(w_n2074_0[1]),.dout(n2102),.clk(gclk));
	jxor g2027(.dina(w_n2101_0[0]),.dinb(w_n2074_0[0]),.dout(n2103),.clk(gclk));
	jxor g2028(.dina(w_n2065_0[0]),.dinb(w_n2057_0[0]),.dout(n2104),.clk(gclk));
	jand g2029(.dina(w_n2104_0[1]),.dinb(w_n2103_0[1]),.dout(n2105),.clk(gclk));
	jor g2030(.dina(n2105),.dinb(n2102),.dout(n2106),.clk(gclk));
	jand g2031(.dina(w_n1356_0[1]),.dinb(w_n58_2[0]),.dout(n2107),.clk(gclk));
	jnot g2032(.din(w_n2107_0[2]),.dout(n2108),.clk(gclk));
	jand g2033(.dina(n2108),.dinb(w_n1413_0[0]),.dout(n2109),.clk(gclk));
	jand g2034(.dina(w_n1682_3[0]),.dinb(w_n699_10[0]),.dout(n2110),.clk(gclk));
	jand g2035(.dina(w_n2110_0[1]),.dinb(w_n1283_6[0]),.dout(n2111),.clk(gclk));
	jnot g2036(.din(n2111),.dout(n2112),.clk(gclk));
	jand g2037(.dina(w_n1283_5[2]),.dinb(w_n1391_2[1]),.dout(n2113),.clk(gclk));
	jor g2038(.dina(n2113),.dinb(w_n2110_0[0]),.dout(n2114),.clk(gclk));
	jor g2039(.dina(n2114),.dinb(w_n1683_2[1]),.dout(n2115),.clk(gclk));
	jand g2040(.dina(n2115),.dinb(n2112),.dout(n2116),.clk(gclk));
	jand g2041(.dina(w_n2116_0[1]),.dinb(w_n2109_0[1]),.dout(n2117),.clk(gclk));
	jand g2042(.dina(w_n2117_0[1]),.dinb(w_n2011_0[1]),.dout(n2118),.clk(gclk));
	jand g2043(.dina(w_n1420_0[0]),.dinb(w_n1762_3[0]),.dout(n2119),.clk(gclk));
	jand g2044(.dina(w_n1417_0[0]),.dinb(w_n75_2[2]),.dout(n2120),.clk(gclk));
	jor g2045(.dina(n2120),.dinb(n2119),.dout(n2121),.clk(gclk));
	jand g2046(.dina(w_n1411_0[2]),.dinb(w_n58_1[2]),.dout(n2122),.clk(gclk));
	jand g2047(.dina(w_n1414_0[2]),.dinb(w_n59_2[0]),.dout(n2123),.clk(gclk));
	jor g2048(.dina(n2123),.dinb(n2122),.dout(n2124),.clk(gclk));
	jand g2049(.dina(n2124),.dinb(n2121),.dout(n2125),.clk(gclk));
	jand g2050(.dina(w_n1566_1[2]),.dinb(w_n1584_1[2]),.dout(n2126),.clk(gclk));
	jand g2051(.dina(w_n1568_1[2]),.dinb(w_n1347_3[0]),.dout(n2127),.clk(gclk));
	jor g2052(.dina(n2127),.dinb(n2126),.dout(n2128),.clk(gclk));
	jor g2053(.dina(w_n1571_1[0]),.dinb(w_n55_6[2]),.dout(n2129),.clk(gclk));
	jor g2054(.dina(w_n1576_0[1]),.dinb(w_n56_9[2]),.dout(n2130),.clk(gclk));
	jand g2055(.dina(n2130),.dinb(n2129),.dout(n2131),.clk(gclk));
	jand g2056(.dina(n2131),.dinb(n2128),.dout(n2132),.clk(gclk));
	jand g2057(.dina(w_n2132_0[1]),.dinb(w_n2125_0[1]),.dout(n2133),.clk(gclk));
	jxor g2058(.dina(w_n2116_0[0]),.dinb(w_n2109_0[0]),.dout(n2134),.clk(gclk));
	jxor g2059(.dina(w_n2132_0[0]),.dinb(w_n2125_0[0]),.dout(n2135),.clk(gclk));
	jand g2060(.dina(w_n2135_0[1]),.dinb(w_n2134_0[1]),.dout(n2136),.clk(gclk));
	jor g2061(.dina(n2136),.dinb(n2133),.dout(n2137),.clk(gclk));
	jxor g2062(.dina(w_n2117_0[0]),.dinb(w_n2011_0[0]),.dout(n2138),.clk(gclk));
	jand g2063(.dina(w_n2138_0[1]),.dinb(w_n2137_0[1]),.dout(n2139),.clk(gclk));
	jor g2064(.dina(n2139),.dinb(n2118),.dout(n2140),.clk(gclk));
	jxor g2065(.dina(w_n2138_0[0]),.dinb(w_n2137_0[0]),.dout(n2141),.clk(gclk));
	jand g2066(.dina(w_n1682_2[2]),.dinb(w_n337_1[2]),.dout(n2142),.clk(gclk));
	jand g2067(.dina(w_n2142_0[1]),.dinb(w_n1283_5[1]),.dout(n2143),.clk(gclk));
	jnot g2068(.din(n2143),.dout(n2144),.clk(gclk));
	jand g2069(.dina(w_n1584_1[1]),.dinb(w_n1283_5[0]),.dout(n2145),.clk(gclk));
	jor g2070(.dina(n2145),.dinb(w_n2142_0[0]),.dout(n2146),.clk(gclk));
	jor g2071(.dina(n2146),.dinb(w_n1683_2[0]),.dout(n2147),.clk(gclk));
	jand g2072(.dina(n2147),.dinb(n2144),.dout(n2148),.clk(gclk));
	jor g2073(.dina(w_n1568_1[1]),.dinb(w_n56_9[1]),.dout(n2149),.clk(gclk));
	jor g2074(.dina(w_n1566_1[1]),.dinb(w_n55_6[1]),.dout(n2150),.clk(gclk));
	jand g2075(.dina(n2150),.dinb(n2149),.dout(n2151),.clk(gclk));
	jor g2076(.dina(w_n1576_0[0]),.dinb(w_n1762_2[2]),.dout(n2152),.clk(gclk));
	jor g2077(.dina(w_n1571_0[2]),.dinb(w_n75_2[1]),.dout(n2153),.clk(gclk));
	jand g2078(.dina(n2153),.dinb(n2152),.dout(n2154),.clk(gclk));
	jand g2079(.dina(n2154),.dinb(n2151),.dout(n2155),.clk(gclk));
	jand g2080(.dina(w_n2155_0[1]),.dinb(w_n2148_0[1]),.dout(n2156),.clk(gclk));
	jand g2081(.dina(w_n1574_0[0]),.dinb(w_n58_1[1]),.dout(n2157),.clk(gclk));
	jnot g2082(.din(w_n2157_0[1]),.dout(n2158),.clk(gclk));
	jand g2083(.dina(n2158),.dinb(w_n1340_0[0]),.dout(n2159),.clk(gclk));
	jand g2084(.dina(w_n1682_2[1]),.dinb(w_n1347_2[2]),.dout(n2160),.clk(gclk));
	jnot g2085(.din(w_n2160_0[1]),.dout(n2161),.clk(gclk));
	jor g2086(.dina(n2161),.dinb(w_n1243_1[0]),.dout(n2162),.clk(gclk));
	jand g2087(.dina(w_n1283_4[2]),.dinb(w_n56_9[0]),.dout(n2163),.clk(gclk));
	jor g2088(.dina(n2163),.dinb(w_n2160_0[0]),.dout(n2164),.clk(gclk));
	jor g2089(.dina(n2164),.dinb(w_n1683_1[2]),.dout(n2165),.clk(gclk));
	jand g2090(.dina(n2165),.dinb(n2162),.dout(n2166),.clk(gclk));
	jand g2091(.dina(w_n2166_0[1]),.dinb(w_n2159_0[1]),.dout(n2167),.clk(gclk));
	jxor g2092(.dina(w_n2155_0[0]),.dinb(w_n2148_0[0]),.dout(n2168),.clk(gclk));
	jand g2093(.dina(w_n2168_0[1]),.dinb(w_n2167_0[1]),.dout(n2169),.clk(gclk));
	jor g2094(.dina(n2169),.dinb(n2156),.dout(n2170),.clk(gclk));
	jxor g2095(.dina(w_n2135_0[0]),.dinb(w_n2134_0[0]),.dout(n2171),.clk(gclk));
	jor g2096(.dina(w_n2171_0[1]),.dinb(w_n2170_0[1]),.dout(n2172),.clk(gclk));
	jand g2097(.dina(w_n2171_0[0]),.dinb(w_n2170_0[0]),.dout(n2173),.clk(gclk));
	jand g2098(.dina(w_n1682_2[0]),.dinb(w_n55_6[0]),.dout(n2174),.clk(gclk));
	jnot g2099(.din(w_n2174_0[1]),.dout(n2175),.clk(gclk));
	jor g2100(.dina(n2175),.dinb(w_n1243_0[2]),.dout(n2176),.clk(gclk));
	jand g2101(.dina(w_n1283_4[1]),.dinb(w_n1762_2[1]),.dout(n2177),.clk(gclk));
	jor g2102(.dina(n2177),.dinb(w_n2174_0[0]),.dout(n2178),.clk(gclk));
	jor g2103(.dina(n2178),.dinb(w_n1683_1[1]),.dout(n2179),.clk(gclk));
	jand g2104(.dina(n2179),.dinb(n2176),.dout(n2180),.clk(gclk));
	jnot g2105(.din(w_n1682_1[2]),.dout(n2181),.clk(gclk));
	jor g2106(.dina(n2181),.dinb(w_n1762_2[0]),.dout(n2182),.clk(gclk));
	jand g2107(.dina(w_n1283_4[0]),.dinb(w_n59_1[2]),.dout(n2183),.clk(gclk));
	jand g2108(.dina(n2183),.dinb(n2182),.dout(n2184),.clk(gclk));
	jor g2109(.dina(w_n2184_0[1]),.dinb(w_n2180_0[1]),.dout(n2185),.clk(gclk));
	jand g2110(.dina(w_n2184_0[0]),.dinb(w_n2180_0[0]),.dout(n2186),.clk(gclk));
	jand g2111(.dina(w_n2157_0[0]),.dinb(w_n1575_0[0]),.dout(n2187),.clk(gclk));
	jand g2112(.dina(w_n2187_0[1]),.dinb(w_n1339_0[0]),.dout(n2188),.clk(gclk));
	jor g2113(.dina(n2188),.dinb(n2186),.dout(n2189),.clk(gclk));
	jand g2114(.dina(n2189),.dinb(n2185),.dout(n2190),.clk(gclk));
	jxor g2115(.dina(w_n2166_0[0]),.dinb(w_n2159_0[0]),.dout(n2191),.clk(gclk));
	jand g2116(.dina(w_n1571_0[1]),.dinb(w_n59_1[1]),.dout(n2192),.clk(gclk));
	jor g2117(.dina(n2192),.dinb(w_n2187_0[0]),.dout(n2193),.clk(gclk));
	jor g2118(.dina(w_n1568_1[0]),.dinb(w_n1762_1[2]),.dout(n2194),.clk(gclk));
	jor g2119(.dina(w_n1566_1[0]),.dinb(w_n75_2[0]),.dout(n2195),.clk(gclk));
	jand g2120(.dina(n2195),.dinb(n2194),.dout(n2196),.clk(gclk));
	jand g2121(.dina(n2196),.dinb(n2193),.dout(n2197),.clk(gclk));
	jand g2122(.dina(w_n2197_0[1]),.dinb(w_n2191_0[1]),.dout(n2198),.clk(gclk));
	jor g2123(.dina(n2198),.dinb(n2190),.dout(n2199),.clk(gclk));
	jor g2124(.dina(w_n2197_0[0]),.dinb(w_n2191_0[0]),.dout(n2200),.clk(gclk));
	jand g2125(.dina(n2200),.dinb(n2199),.dout(n2201),.clk(gclk));
	jor g2126(.dina(w_n2201_0[1]),.dinb(w_n2107_0[1]),.dout(n2202),.clk(gclk));
	jand g2127(.dina(w_n2201_0[0]),.dinb(w_n2107_0[0]),.dout(n2203),.clk(gclk));
	jxor g2128(.dina(w_n2168_0[0]),.dinb(w_n2167_0[0]),.dout(n2204),.clk(gclk));
	jor g2129(.dina(n2204),.dinb(n2203),.dout(n2205),.clk(gclk));
	jand g2130(.dina(n2205),.dinb(n2202),.dout(n2206),.clk(gclk));
	jor g2131(.dina(n2206),.dinb(n2173),.dout(n2207),.clk(gclk));
	jand g2132(.dina(n2207),.dinb(n2172),.dout(n2208),.clk(gclk));
	jor g2133(.dina(w_n2208_0[1]),.dinb(w_n2141_0[1]),.dout(n2209),.clk(gclk));
	jand g2134(.dina(w_n2208_0[0]),.dinb(w_n2141_0[0]),.dout(n2210),.clk(gclk));
	jxor g2135(.dina(w_n2099_0[0]),.dinb(w_n2091_0[0]),.dout(n2211),.clk(gclk));
	jor g2136(.dina(n2211),.dinb(n2210),.dout(n2212),.clk(gclk));
	jand g2137(.dina(n2212),.dinb(n2209),.dout(n2213),.clk(gclk));
	jor g2138(.dina(w_n2213_0[1]),.dinb(w_n2140_0[1]),.dout(n2214),.clk(gclk));
	jand g2139(.dina(w_n2213_0[0]),.dinb(w_n2140_0[0]),.dout(n2215),.clk(gclk));
	jxor g2140(.dina(w_n2104_0[0]),.dinb(w_n2103_0[0]),.dout(n2216),.clk(gclk));
	jor g2141(.dina(n2216),.dinb(n2215),.dout(n2217),.clk(gclk));
	jand g2142(.dina(n2217),.dinb(n2214),.dout(n2218),.clk(gclk));
	jor g2143(.dina(w_n2218_0[1]),.dinb(w_n2106_0[1]),.dout(n2219),.clk(gclk));
	jand g2144(.dina(w_n2218_0[0]),.dinb(w_n2106_0[0]),.dout(n2220),.clk(gclk));
	jxor g2145(.dina(w_n2071_0[0]),.dinb(w_n2070_0[0]),.dout(n2221),.clk(gclk));
	jor g2146(.dina(n2221),.dinb(n2220),.dout(n2222),.clk(gclk));
	jand g2147(.dina(n2222),.dinb(n2219),.dout(n2223),.clk(gclk));
	jor g2148(.dina(w_n2223_0[1]),.dinb(w_n2073_0[1]),.dout(n2224),.clk(gclk));
	jand g2149(.dina(w_n2223_0[0]),.dinb(w_n2073_0[0]),.dout(n2225),.clk(gclk));
	jxor g2150(.dina(w_n2037_0[0]),.dinb(w_n2036_0[0]),.dout(n2226),.clk(gclk));
	jor g2151(.dina(n2226),.dinb(n2225),.dout(n2227),.clk(gclk));
	jand g2152(.dina(n2227),.dinb(n2224),.dout(n2228),.clk(gclk));
	jor g2153(.dina(w_n2228_0[1]),.dinb(w_n2039_0[1]),.dout(n2229),.clk(gclk));
	jand g2154(.dina(w_n2228_0[0]),.dinb(w_n2039_0[0]),.dout(n2230),.clk(gclk));
	jxor g2155(.dina(w_n2008_0[0]),.dinb(w_n2007_0[0]),.dout(n2231),.clk(gclk));
	jor g2156(.dina(n2231),.dinb(n2230),.dout(n2232),.clk(gclk));
	jand g2157(.dina(n2232),.dinb(n2229),.dout(n2233),.clk(gclk));
	jor g2158(.dina(w_n2233_0[1]),.dinb(w_n2010_0[1]),.dout(n2234),.clk(gclk));
	jand g2159(.dina(w_n2233_0[0]),.dinb(w_n2010_0[0]),.dout(n2235),.clk(gclk));
	jxor g2160(.dina(w_n1959_0[0]),.dinb(w_n1958_0[0]),.dout(n2236),.clk(gclk));
	jor g2161(.dina(n2236),.dinb(n2235),.dout(n2237),.clk(gclk));
	jand g2162(.dina(n2237),.dinb(n2234),.dout(n2238),.clk(gclk));
	jand g2163(.dina(w_n2238_0[1]),.dinb(w_n1964_0[1]),.dout(n2239),.clk(gclk));
	jor g2164(.dina(n2239),.dinb(n1963),.dout(n2240),.clk(gclk));
	jxor g2165(.dina(w_n1921_0[0]),.dinb(w_n1920_0[0]),.dout(n2241),.clk(gclk));
	jand g2166(.dina(w_n2241_0[1]),.dinb(w_n2240_0[1]),.dout(n2242),.clk(gclk));
	jor g2167(.dina(n2242),.dinb(n1922),.dout(n2243),.clk(gclk));
	jxor g2168(.dina(w_n1850_0[0]),.dinb(w_n1849_0[0]),.dout(n2244),.clk(gclk));
	jand g2169(.dina(w_n2244_0[1]),.dinb(w_n2243_0[1]),.dout(n2245),.clk(gclk));
	jor g2170(.dina(n2245),.dinb(n1851),.dout(n2246),.clk(gclk));
	jxor g2171(.dina(w_n1815_0[0]),.dinb(w_n1814_0[0]),.dout(n2247),.clk(gclk));
	jand g2172(.dina(w_n2247_0[1]),.dinb(w_n2246_0[1]),.dout(n2248),.clk(gclk));
	jor g2173(.dina(n2248),.dinb(n1816),.dout(n2249),.clk(gclk));
	jxor g2174(.dina(w_n1749_0[0]),.dinb(w_n1748_0[0]),.dout(n2250),.clk(gclk));
	jand g2175(.dina(w_n2250_0[1]),.dinb(w_n2249_0[1]),.dout(n2251),.clk(gclk));
	jor g2176(.dina(n2251),.dinb(n1750),.dout(n2252),.clk(gclk));
	jxor g2177(.dina(w_n1635_0[0]),.dinb(w_n1634_0[0]),.dout(n2253),.clk(gclk));
	jand g2178(.dina(w_n2253_0[1]),.dinb(w_n2252_0[1]),.dout(n2254),.clk(gclk));
	jor g2179(.dina(n2254),.dinb(n1636),.dout(n2255),.clk(gclk));
	jxor g2180(.dina(w_n1440_0[0]),.dinb(w_n1439_0[0]),.dout(n2256),.clk(gclk));
	jand g2181(.dina(w_n2256_0[1]),.dinb(w_n2255_0[1]),.dout(n2257),.clk(gclk));
	jor g2182(.dina(n2257),.dinb(n1441),.dout(n2258),.clk(gclk));
	jxor g2183(.dina(w_n1389_0[0]),.dinb(w_n1388_0[0]),.dout(n2259),.clk(gclk));
	jand g2184(.dina(w_n2259_0[1]),.dinb(w_n2258_0[1]),.dout(n2260),.clk(gclk));
	jor g2185(.dina(n2260),.dinb(n1390),.dout(n2261),.clk(gclk));
	jxor g2186(.dina(w_n1140_0[0]),.dinb(w_n1113_0[0]),.dout(n2262),.clk(gclk));
	jand g2187(.dina(w_n2262_0[1]),.dinb(w_n2261_0[1]),.dout(n2263),.clk(gclk));
	jor g2188(.dina(n2263),.dinb(n1141),.dout(n2264),.clk(gclk));
	jand g2189(.dina(w_n1138_0[0]),.dinb(w_n1133_0[0]),.dout(n2265),.clk(gclk));
	jand g2190(.dina(w_n1139_0[0]),.dinb(w_n1130_0[0]),.dout(n2266),.clk(gclk));
	jor g2191(.dina(n2266),.dinb(n2265),.dout(n2267),.clk(gclk));
	jand g2192(.dina(w_n1120_0[0]),.dinb(w_n1115_0[1]),.dout(n2268),.clk(gclk));
	jand g2193(.dina(w_n1129_0[0]),.dinb(w_n1121_0[0]),.dout(n2269),.clk(gclk));
	jor g2194(.dina(n2269),.dinb(n2268),.dout(n2270),.clk(gclk));
	jor g2195(.dina(w_n954_20[2]),.dinb(w_n795_0[2]),.dout(n2272),.clk(gclk));
	jor g2196(.dina(w_n960_2[1]),.dinb(w_n800_0[0]),.dout(n2275),.clk(gclk));
	jor g2197(.dina(w_n961_2[0]),.dinb(w_n792_0[0]),.dout(n2276),.clk(gclk));
	jand g2198(.dina(n2276),.dinb(n2275),.dout(n2277),.clk(gclk));
	jand g2199(.dina(n2277),.dinb(n2272),.dout(n2278),.clk(gclk));
	jxor g2200(.dina(w_n2278_0[1]),.dinb(w_n2270_0[1]),.dout(n2279),.clk(gclk));
	jxor g2201(.dina(w_n1115_0[0]),.dinb(w_n1047_0[1]),.dout(n2280),.clk(gclk));
	jand g2202(.dina(w_n980_2[2]),.dinb(w_n335_3[0]),.dout(n2281),.clk(gclk));
	jxor g2203(.dina(w_n2281_0[1]),.dinb(w_n2280_0[1]),.dout(n2282),.clk(gclk));
	jxor g2204(.dina(w_n2282_0[1]),.dinb(w_n2279_0[1]),.dout(n2283),.clk(gclk));
	jxor g2205(.dina(w_n2283_0[1]),.dinb(w_n2267_0[1]),.dout(n2284),.clk(gclk));
	jxor g2206(.dina(w_n2284_0[1]),.dinb(w_n2264_0[1]),.dout(n2285),.clk(gclk));
	jand g2207(.dina(w_n645_1[1]),.dinb(w_n261_1[0]),.dout(n2286),.clk(gclk));
	jand g2208(.dina(w_n356_0[2]),.dinb(w_n310_1[0]),.dout(n2287),.clk(gclk));
	jand g2209(.dina(w_n2287_0[1]),.dinb(w_n2286_0[1]),.dout(n2288),.clk(gclk));
	jand g2210(.dina(w_n445_2[0]),.dinb(w_n365_1[0]),.dout(n2289),.clk(gclk));
	jand g2211(.dina(w_n2289_0[1]),.dinb(w_n504_0[0]),.dout(n2290),.clk(gclk));
	jand g2212(.dina(n2290),.dinb(n2288),.dout(n2291),.clk(gclk));
	jand g2213(.dina(w_n781_1[1]),.dinb(w_n732_2[1]),.dout(n2292),.clk(gclk));
	jand g2214(.dina(n2292),.dinb(w_n470_1[0]),.dout(n2293),.clk(gclk));
	jand g2215(.dina(n2293),.dinb(w_n917_0[0]),.dout(n2294),.clk(gclk));
	jand g2216(.dina(w_n490_0[0]),.dinb(w_n392_0[1]),.dout(n2295),.clk(gclk));
	jand g2217(.dina(n2295),.dinb(n2294),.dout(n2296),.clk(gclk));
	jand g2218(.dina(n2296),.dinb(n2291),.dout(n2297),.clk(gclk));
	jand g2219(.dina(w_n991_0[0]),.dinb(w_n675_0[1]),.dout(n2298),.clk(gclk));
	jand g2220(.dina(n2298),.dinb(n2297),.dout(n2299),.clk(gclk));
	jand g2221(.dina(n2299),.dinb(w_n1203_0[1]),.dout(n2300),.clk(gclk));
	jor g2222(.dina(w_n2300_0[1]),.dinb(w_n2285_0[1]),.dout(n2301),.clk(gclk));
	jxor g2223(.dina(w_n2262_0[0]),.dinb(w_n2261_0[0]),.dout(n2302),.clk(gclk));
	jand g2224(.dina(w_n477_2[0]),.dinb(w_n401_1[1]),.dout(n2303),.clk(gclk));
	jand g2225(.dina(n2303),.dinb(w_n436_1[2]),.dout(n2304),.clk(gclk));
	jand g2226(.dina(w_n734_1[0]),.dinb(w_n368_1[2]),.dout(n2305),.clk(gclk));
	jand g2227(.dina(w_n2305_0[1]),.dinb(w_n507_1[0]),.dout(n2306),.clk(gclk));
	jand g2228(.dina(n2306),.dinb(n2304),.dout(n2307),.clk(gclk));
	jand g2229(.dina(w_n312_2[2]),.dinb(w_n216_2[2]),.dout(n2308),.clk(gclk));
	jand g2230(.dina(w_n387_1[0]),.dinb(w_n243_2[2]),.dout(n2309),.clk(gclk));
	jand g2231(.dina(n2309),.dinb(n2308),.dout(n2310),.clk(gclk));
	jand g2232(.dina(n2310),.dinb(w_n1002_0[0]),.dout(n2311),.clk(gclk));
	jand g2233(.dina(n2311),.dinb(w_n885_0[0]),.dout(n2312),.clk(gclk));
	jand g2234(.dina(n2312),.dinb(w_n2307_0[1]),.dout(n2313),.clk(gclk));
	jand g2235(.dina(w_n765_1[0]),.dinb(w_n412_1[1]),.dout(n2314),.clk(gclk));
	jand g2236(.dina(n2314),.dinb(w_n676_0[1]),.dout(n2315),.clk(gclk));
	jand g2237(.dina(w_n561_1[0]),.dinb(w_n363_1[1]),.dout(n2316),.clk(gclk));
	jand g2238(.dina(w_n285_1[1]),.dinb(w_n147_2[2]),.dout(n2317),.clk(gclk));
	jand g2239(.dina(n2317),.dinb(n2316),.dout(n2318),.clk(gclk));
	jand g2240(.dina(n2318),.dinb(w_n2315_0[1]),.dout(n2319),.clk(gclk));
	jand g2241(.dina(w_n757_0[0]),.dinb(w_n254_2[0]),.dout(n2320),.clk(gclk));
	jand g2242(.dina(n2320),.dinb(w_n138_2[2]),.dout(n2321),.clk(gclk));
	jand g2243(.dina(w_n642_1[0]),.dinb(w_n264_2[0]),.dout(n2322),.clk(gclk));
	jand g2244(.dina(n2322),.dinb(w_n614_2[0]),.dout(n2323),.clk(gclk));
	jand g2245(.dina(w_n2323_0[1]),.dinb(w_n2321_0[2]),.dout(n2324),.clk(gclk));
	jand g2246(.dina(n2324),.dinb(n2319),.dout(n2325),.clk(gclk));
	jand g2247(.dina(w_n668_2[0]),.dinb(w_n356_0[1]),.dout(n2326),.clk(gclk));
	jand g2248(.dina(w_n2326_0[2]),.dinb(w_n1018_0[2]),.dout(n2327),.clk(gclk));
	jand g2249(.dina(n2327),.dinb(w_n924_0[2]),.dout(n2328),.clk(gclk));
	jand g2250(.dina(n2328),.dinb(w_n881_1[0]),.dout(n2329),.clk(gclk));
	jand g2251(.dina(n2329),.dinb(n2325),.dout(n2330),.clk(gclk));
	jand g2252(.dina(w_n430_2[0]),.dinb(w_n282_2[1]),.dout(n2331),.clk(gclk));
	jand g2253(.dina(w_n2331_0[1]),.dinb(w_n441_0[2]),.dout(n2332),.clk(gclk));
	jand g2254(.dina(w_n849_1[0]),.dinb(w_n358_1[1]),.dout(n2333),.clk(gclk));
	jand g2255(.dina(n2333),.dinb(w_n473_1[0]),.dout(n2334),.clk(gclk));
	jand g2256(.dina(w_n935_2[0]),.dinb(w_n709_0[2]),.dout(n2335),.clk(gclk));
	jand g2257(.dina(w_n2335_0[1]),.dinb(w_n710_2[1]),.dout(n2336),.clk(gclk));
	jand g2258(.dina(n2336),.dinb(w_n2334_0[2]),.dout(n2337),.clk(gclk));
	jand g2259(.dina(n2337),.dinb(w_n2332_0[1]),.dout(n2338),.clk(gclk));
	jand g2260(.dina(w_n853_2[0]),.dinb(w_n488_1[1]),.dout(n2339),.clk(gclk));
	jand g2261(.dina(w_n1025_0[1]),.dinb(w_n822_2[0]),.dout(n2340),.clk(gclk));
	jand g2262(.dina(n2340),.dinb(w_n2339_0[1]),.dout(n2341),.clk(gclk));
	jand g2263(.dina(n2341),.dinb(w_n876_0[0]),.dout(n2342),.clk(gclk));
	jand g2264(.dina(n2342),.dinb(n2338),.dout(n2343),.clk(gclk));
	jand g2265(.dina(n2343),.dinb(w_n2330_0[1]),.dout(n2344),.clk(gclk));
	jand g2266(.dina(n2344),.dinb(w_n2313_0[1]),.dout(n2345),.clk(gclk));
	jor g2267(.dina(w_n2345_0[1]),.dinb(w_n2302_0[1]),.dout(n2346),.clk(gclk));
	jxor g2268(.dina(w_n2259_0[0]),.dinb(w_n2258_0[0]),.dout(n2347),.clk(gclk));
	jand g2269(.dina(w_n501_1[1]),.dinb(w_n157_1[0]),.dout(n2348),.clk(gclk));
	jand g2270(.dina(n2348),.dinb(w_n422_2[0]),.dout(n2349),.clk(gclk));
	jand g2271(.dina(n2349),.dinb(w_n2330_0[0]),.dout(n2350),.clk(gclk));
	jand g2272(.dina(w_n594_2[0]),.dinb(w_n897_0[1]),.dout(n2351),.clk(gclk));
	jand g2273(.dina(w_n532_1[0]),.dinb(w_n270_1[2]),.dout(n2352),.clk(gclk));
	jand g2274(.dina(n2352),.dinb(w_n2351_0[1]),.dout(n2353),.clk(gclk));
	jand g2275(.dina(n2353),.dinb(w_n305_0[1]),.dout(n2354),.clk(gclk));
	jand g2276(.dina(w_n993_1[0]),.dinb(w_n451_2[0]),.dout(n2355),.clk(gclk));
	jand g2277(.dina(n2355),.dinb(w_n372_1[1]),.dout(n2356),.clk(gclk));
	jand g2278(.dina(n2356),.dinb(w_n741_0[1]),.dout(n2357),.clk(gclk));
	jand g2279(.dina(n2357),.dinb(w_n2334_0[1]),.dout(n2358),.clk(gclk));
	jand g2280(.dina(n2358),.dinb(n2354),.dout(n2359),.clk(gclk));
	jand g2281(.dina(w_n401_1[0]),.dinb(w_n225_1[1]),.dout(n2360),.clk(gclk));
	jand g2282(.dina(w_n732_2[0]),.dinb(w_n1209_1[1]),.dout(n2361),.clk(gclk));
	jand g2283(.dina(w_n763_1[2]),.dinb(w_n837_1[2]),.dout(n2362),.clk(gclk));
	jand g2284(.dina(n2362),.dinb(n2361),.dout(n2363),.clk(gclk));
	jand g2285(.dina(n2363),.dinb(w_n2360_0[1]),.dout(n2364),.clk(gclk));
	jand g2286(.dina(n2364),.dinb(w_n912_0[0]),.dout(n2365),.clk(gclk));
	jand g2287(.dina(w_n664_0[1]),.dinb(w_n295_2[0]),.dout(n2366),.clk(gclk));
	jand g2288(.dina(w_n282_2[0]),.dinb(w_n251_2[0]),.dout(n2367),.clk(gclk));
	jand g2289(.dina(n2367),.dinb(n2366),.dout(n2368),.clk(gclk));
	jand g2290(.dina(w_n619_1[1]),.dinb(w_n597_1[1]),.dout(n2369),.clk(gclk));
	jand g2291(.dina(n2369),.dinb(n2368),.dout(n2370),.clk(gclk));
	jand g2292(.dina(w_n477_1[2]),.dinb(w_n445_1[2]),.dout(n2371),.clk(gclk));
	jand g2293(.dina(n2371),.dinb(w_n499_0[2]),.dout(n2372),.clk(gclk));
	jand g2294(.dina(w_n2372_0[2]),.dinb(w_n1646_0[1]),.dout(n2373),.clk(gclk));
	jand g2295(.dina(n2373),.dinb(n2370),.dout(n2374),.clk(gclk));
	jand g2296(.dina(n2374),.dinb(w_n2365_0[2]),.dout(n2375),.clk(gclk));
	jand g2297(.dina(n2375),.dinb(w_n2359_0[1]),.dout(n2376),.clk(gclk));
	jand g2298(.dina(n2376),.dinb(w_n2350_0[1]),.dout(n2377),.clk(gclk));
	jor g2299(.dina(w_n2377_0[1]),.dinb(w_n2347_0[1]),.dout(n2378),.clk(gclk));
	jxor g2300(.dina(w_n2256_0[0]),.dinb(w_n2255_0[0]),.dout(n2379),.clk(gclk));
	jnot g2301(.din(w_n893_0[0]),.dout(n2380),.clk(gclk));
	jand g2302(.dina(w_n2380_3[1]),.dinb(w_n370_1[1]),.dout(n2381),.clk(gclk));
	jand g2303(.dina(n2381),.dinb(w_n1169_0[0]),.dout(n2382),.clk(gclk));
	jand g2304(.dina(w_n732_1[2]),.dinb(w_n730_0[2]),.dout(n2383),.clk(gclk));
	jand g2305(.dina(n2383),.dinb(w_n1204_0[1]),.dout(n2384),.clk(gclk));
	jand g2306(.dina(w_n461_1[1]),.dinb(w_n130_1[1]),.dout(n2385),.clk(gclk));
	jand g2307(.dina(w_n2385_1[1]),.dinb(w_n1025_0[0]),.dout(n2386),.clk(gclk));
	jand g2308(.dina(w_n477_1[1]),.dinb(w_n303_2[1]),.dout(n2387),.clk(gclk));
	jand g2309(.dina(w_n2387_0[1]),.dinb(w_n301_1[0]),.dout(n2388),.clk(gclk));
	jand g2310(.dina(n2388),.dinb(n2386),.dout(n2389),.clk(gclk));
	jand g2311(.dina(n2389),.dinb(n2384),.dout(n2390),.clk(gclk));
	jand g2312(.dina(n2390),.dinb(w_n1179_0[0]),.dout(n2391),.clk(gclk));
	jand g2313(.dina(w_n470_0[2]),.dinb(w_n243_2[1]),.dout(n2392),.clk(gclk));
	jand g2314(.dina(w_n668_1[2]),.dinb(w_n222_1[1]),.dout(n2393),.clk(gclk));
	jand g2315(.dina(n2393),.dinb(n2392),.dout(n2394),.clk(gclk));
	jnot g2316(.din(w_n1675_0[0]),.dout(n2395),.clk(gclk));
	jand g2317(.dina(w_n763_1[1]),.dinb(w_n312_2[1]),.dout(n2396),.clk(gclk));
	jand g2318(.dina(w_n2396_0[1]),.dinb(n2395),.dout(n2397),.clk(gclk));
	jand g2319(.dina(n2397),.dinb(n2394),.dout(n2398),.clk(gclk));
	jand g2320(.dina(w_n679_1[1]),.dinb(w_n421_2[1]),.dout(n2399),.clk(gclk));
	jand g2321(.dina(w_n744_1[2]),.dinb(w_n294_2[0]),.dout(n2400),.clk(gclk));
	jand g2322(.dina(n2400),.dinb(w_n383_1[2]),.dout(n2401),.clk(gclk));
	jand g2323(.dina(n2401),.dinb(n2399),.dout(n2402),.clk(gclk));
	jand g2324(.dina(w_n614_1[2]),.dinb(w_n138_2[1]),.dout(n2403),.clk(gclk));
	jand g2325(.dina(w_n768_1[2]),.dinb(w_n229_1[1]),.dout(n2404),.clk(gclk));
	jand g2326(.dina(n2404),.dinb(n2403),.dout(n2405),.clk(gclk));
	jand g2327(.dina(w_n430_1[2]),.dinb(w_n323_2[2]),.dout(n2406),.clk(gclk));
	jand g2328(.dina(w_n2406_0[1]),.dinb(w_n740_0[0]),.dout(n2407),.clk(gclk));
	jand g2329(.dina(n2407),.dinb(n2405),.dout(n2408),.clk(gclk));
	jand g2330(.dina(n2408),.dinb(w_n2402_0[1]),.dout(n2409),.clk(gclk));
	jand g2331(.dina(n2409),.dinb(w_n2398_0[1]),.dout(n2410),.clk(gclk));
	jand g2332(.dina(n2410),.dinb(w_n2391_0[1]),.dout(n2411),.clk(gclk));
	jand g2333(.dina(n2411),.dinb(w_n2382_0[1]),.dout(n2412),.clk(gclk));
	jor g2334(.dina(w_n2412_0[1]),.dinb(w_n2379_0[1]),.dout(n2413),.clk(gclk));
	jxor g2335(.dina(w_n2253_0[0]),.dinb(w_n2252_0[0]),.dout(n2414),.clk(gclk));
	jand g2336(.dina(w_n458_1[0]),.dinb(w_n387_0[2]),.dout(n2415),.clk(gclk));
	jand g2337(.dina(n2415),.dinb(w_n724_1[1]),.dout(n2416),.clk(gclk));
	jand g2338(.dina(n2416),.dinb(w_n767_0[0]),.dout(n2417),.clk(gclk));
	jand g2339(.dina(w_n992_1[1]),.dinb(w_n524_0[0]),.dout(n2418),.clk(gclk));
	jand g2340(.dina(n2418),.dinb(w_n286_0[2]),.dout(n2419),.clk(gclk));
	jand g2341(.dina(n2419),.dinb(w_n2417_0[2]),.dout(n2420),.clk(gclk));
	jand g2342(.dina(n2420),.dinb(w_n538_0[0]),.dout(n2421),.clk(gclk));
	jand g2343(.dina(w_n662_1[0]),.dinb(w_n772_2[0]),.dout(n2422),.clk(gclk));
	jand g2344(.dina(n2422),.dinb(w_n523_0[0]),.dout(n2423),.clk(gclk));
	jand g2345(.dina(w_n2380_3[0]),.dinb(w_n679_1[0]),.dout(n2424),.clk(gclk));
	jand g2346(.dina(w_n2424_0[1]),.dinb(w_n1170_0[1]),.dout(n2425),.clk(gclk));
	jand g2347(.dina(n2425),.dinb(n2423),.dout(n2426),.clk(gclk));
	jand g2348(.dina(n2426),.dinb(w_n424_0[0]),.dout(n2427),.clk(gclk));
	jand g2349(.dina(w_n402_1[0]),.dinb(w_n371_0[0]),.dout(n2428),.clk(gclk));
	jand g2350(.dina(w_n744_1[1]),.dinb(w_n222_1[0]),.dout(n2429),.clk(gclk));
	jand g2351(.dina(w_n592_2[1]),.dinb(w_n383_1[1]),.dout(n2430),.clk(gclk));
	jand g2352(.dina(n2430),.dinb(w_n2429_1[1]),.dout(n2431),.clk(gclk));
	jnot g2353(.din(w_n1214_0[0]),.dout(n2432),.clk(gclk));
	jand g2354(.dina(n2432),.dinb(w_n324_0[1]),.dout(n2433),.clk(gclk));
	jand g2355(.dina(n2433),.dinb(n2431),.dout(n2434),.clk(gclk));
	jand g2356(.dina(n2434),.dinb(w_n2428_0[1]),.dout(n2435),.clk(gclk));
	jand g2357(.dina(n2435),.dinb(w_n2427_0[2]),.dout(n2436),.clk(gclk));
	jand g2358(.dina(n2436),.dinb(n2421),.dout(n2437),.clk(gclk));
	jand g2359(.dina(n2437),.dinb(w_n630_0[0]),.dout(n2438),.clk(gclk));
	jor g2360(.dina(w_n2438_0[1]),.dinb(w_n2414_0[1]),.dout(n2439),.clk(gclk));
	jxor g2361(.dina(w_n2250_0[0]),.dinb(w_n2249_0[0]),.dout(n2440),.clk(gclk));
	jand g2362(.dina(w_n918_2[0]),.dinb(w_n532_0[2]),.dout(n2441),.clk(gclk));
	jand g2363(.dina(n2441),.dinb(w_n2385_1[0]),.dout(n2442),.clk(gclk));
	jand g2364(.dina(w_n744_1[0]),.dinb(w_n612_2[1]),.dout(n2443),.clk(gclk));
	jand g2365(.dina(w_n579_1[0]),.dinb(w_n304_1[2]),.dout(n2444),.clk(gclk));
	jand g2366(.dina(n2444),.dinb(n2443),.dout(n2445),.clk(gclk));
	jand g2367(.dina(n2445),.dinb(w_n987_1[1]),.dout(n2446),.clk(gclk));
	jand g2368(.dina(n2446),.dinb(w_n2442_0[1]),.dout(n2447),.clk(gclk));
	jand g2369(.dina(w_n1332_0[0]),.dinb(w_n881_0[2]),.dout(n2448),.clk(gclk));
	jand g2370(.dina(n2448),.dinb(n2447),.dout(n2449),.clk(gclk));
	jand g2371(.dina(w_n822_1[2]),.dinb(w_n397_0[2]),.dout(n2450),.clk(gclk));
	jand g2372(.dina(n2450),.dinb(w_n2449_0[1]),.dout(n2451),.clk(gclk));
	jand g2373(.dina(w_n853_1[2]),.dinb(w_n264_1[2]),.dout(n2452),.clk(gclk));
	jand g2374(.dina(n2452),.dinb(w_n739_0[1]),.dout(n2453),.clk(gclk));
	jand g2375(.dina(w_n348_0[2]),.dinb(w_n897_0[0]),.dout(n2454),.clk(gclk));
	jand g2376(.dina(n2454),.dinb(w_n643_0[0]),.dout(n2455),.clk(gclk));
	jand g2377(.dina(w_n445_1[1]),.dinb(w_n323_2[1]),.dout(n2456),.clk(gclk));
	jand g2378(.dina(w_n381_1[0]),.dinb(w_n279_1[1]),.dout(n2457),.clk(gclk));
	jand g2379(.dina(w_n2457_0[1]),.dinb(w_n2456_0[2]),.dout(n2458),.clk(gclk));
	jand g2380(.dina(n2458),.dinb(n2455),.dout(n2459),.clk(gclk));
	jand g2381(.dina(n2459),.dinb(w_n2453_0[1]),.dout(n2460),.clk(gclk));
	jand g2382(.dina(n2460),.dinb(w_n509_0[0]),.dout(n2461),.clk(gclk));
	jand g2383(.dina(w_n837_1[1]),.dinb(w_n282_1[2]),.dout(n2462),.clk(gclk));
	jand g2384(.dina(w_n751_2[0]),.dinb(w_n216_2[1]),.dout(n2463),.clk(gclk));
	jand g2385(.dina(n2463),.dinb(n2462),.dout(n2464),.clk(gclk));
	jand g2386(.dina(w_n2287_0[0]),.dinb(w_n301_0[2]),.dout(n2465),.clk(gclk));
	jand g2387(.dina(n2465),.dinb(n2464),.dout(n2466),.clk(gclk));
	jand g2388(.dina(w_n742_0[0]),.dinb(w_n427_1[2]),.dout(n2467),.clk(gclk));
	jand g2389(.dina(w_n295_1[2]),.dinb(w_n285_1[0]),.dout(n2468),.clk(gclk));
	jand g2390(.dina(n2468),.dinb(n2467),.dout(n2469),.clk(gclk));
	jnot g2391(.din(w_n346_2[1]),.dout(n2470),.clk(gclk));
	jand g2392(.dina(n2470),.dinb(w_n325_0[0]),.dout(n2471),.clk(gclk));
	jor g2393(.dina(n2471),.dinb(w_n326_0[0]),.dout(n2472),.clk(gclk));
	jand g2394(.dina(n2472),.dinb(w_n417_1[1]),.dout(n2473),.clk(gclk));
	jand g2395(.dina(n2473),.dinb(n2469),.dout(n2474),.clk(gclk));
	jand g2396(.dina(n2474),.dinb(w_n2466_0[1]),.dout(n2475),.clk(gclk));
	jand g2397(.dina(n2475),.dinb(w_n2461_0[1]),.dout(n2476),.clk(gclk));
	jand g2398(.dina(n2476),.dinb(w_n2451_0[1]),.dout(n2477),.clk(gclk));
	jor g2399(.dina(w_n2477_0[1]),.dinb(w_n2440_0[1]),.dout(n2478),.clk(gclk));
	jxor g2400(.dina(w_n2247_0[0]),.dinb(w_n2246_0[0]),.dout(n2479),.clk(gclk));
	jand g2401(.dina(w_n2380_2[2]),.dinb(w_n612_2[0]),.dout(n2480),.clk(gclk));
	jand g2402(.dina(w_n665_1[1]),.dinb(w_n772_1[2]),.dout(n2481),.clk(gclk));
	jand g2403(.dina(n2481),.dinb(n2480),.dout(n2482),.clk(gclk));
	jand g2404(.dina(n2482),.dinb(w_n507_0[2]),.dout(n2483),.clk(gclk));
	jand g2405(.dina(w_n2332_0[0]),.dinb(w_n836_0[0]),.dout(n2484),.clk(gclk));
	jand g2406(.dina(n2484),.dinb(w_n234_0[0]),.dout(n2485),.clk(gclk));
	jand g2407(.dina(n2485),.dinb(n2483),.dout(n2486),.clk(gclk));
	jand g2408(.dina(w_n853_1[1]),.dinb(w_n925_1[0]),.dout(n2487),.clk(gclk));
	jand g2409(.dina(n2487),.dinb(w_n501_1[0]),.dout(n2488),.clk(gclk));
	jand g2410(.dina(w_n668_1[1]),.dinb(w_n138_2[0]),.dout(n2489),.clk(gclk));
	jand g2411(.dina(w_n624_1[2]),.dinb(w_n294_1[2]),.dout(n2490),.clk(gclk));
	jand g2412(.dina(w_n2490_0[1]),.dinb(n2489),.dout(n2491),.clk(gclk));
	jand g2413(.dina(n2491),.dinb(n2488),.dout(n2492),.clk(gclk));
	jand g2414(.dina(n2492),.dinb(w_n611_1[0]),.dout(n2493),.clk(gclk));
	jnot g2415(.din(w_n1215_0[0]),.dout(n2494),.clk(gclk));
	jand g2416(.dina(w_n642_0[2]),.dinb(w_n768_1[1]),.dout(n2495),.clk(gclk));
	jand g2417(.dina(n2495),.dinb(n2494),.dout(n2496),.clk(gclk));
	jand g2418(.dina(w_n1022_0[1]),.dinb(w_n265_0[1]),.dout(n2497),.clk(gclk));
	jand g2419(.dina(n2497),.dinb(n2496),.dout(n2498),.clk(gclk));
	jand g2420(.dina(w_n2335_0[0]),.dinb(w_n821_0[2]),.dout(n2499),.clk(gclk));
	jand g2421(.dina(n2499),.dinb(w_n869_0[1]),.dout(n2500),.clk(gclk));
	jand g2422(.dina(n2500),.dinb(w_n2498_0[1]),.dout(n2501),.clk(gclk));
	jand g2423(.dina(n2501),.dinb(n2493),.dout(n2502),.clk(gclk));
	jand g2424(.dina(n2502),.dinb(w_n2486_0[1]),.dout(n2503),.clk(gclk));
	jand g2425(.dina(n2503),.dinb(w_n395_0[1]),.dout(n2504),.clk(gclk));
	jor g2426(.dina(w_n2504_0[2]),.dinb(w_n2479_0[2]),.dout(n2505),.clk(gclk));
	jxor g2427(.dina(w_n2244_0[0]),.dinb(w_n2243_0[0]),.dout(n2506),.clk(gclk));
	jand g2428(.dina(w_n612_1[2]),.dinb(w_n427_1[1]),.dout(n2507),.clk(gclk));
	jand g2429(.dina(n2507),.dinb(w_n987_1[0]),.dout(n2508),.clk(gclk));
	jand g2430(.dina(n2508),.dinb(w_n605_0[0]),.dout(n2509),.clk(gclk));
	jand g2431(.dina(n2509),.dinb(w_n2372_0[1]),.dout(n2510),.clk(gclk));
	jand g2432(.dina(w_n993_0[2]),.dinb(w_n837_1[0]),.dout(n2511),.clk(gclk));
	jand g2433(.dina(w_n710_2[0]),.dinb(w_n594_1[2]),.dout(n2512),.clk(gclk));
	jand g2434(.dina(n2512),.dinb(w_n734_0[2]),.dout(n2513),.clk(gclk));
	jand g2435(.dina(n2513),.dinb(w_n2511_1[1]),.dout(n2514),.clk(gclk));
	jand g2436(.dina(w_n739_0[0]),.dinb(w_n501_0[2]),.dout(n2515),.clk(gclk));
	jand g2437(.dina(w_n2515_0[2]),.dinb(w_n680_1[0]),.dout(n2516),.clk(gclk));
	jand g2438(.dina(n2516),.dinb(w_n1328_0[0]),.dout(n2517),.clk(gclk));
	jand g2439(.dina(n2517),.dinb(w_n2417_0[1]),.dout(n2518),.clk(gclk));
	jand g2440(.dina(n2518),.dinb(w_n2514_0[1]),.dout(n2519),.clk(gclk));
	jand g2441(.dina(n2519),.dinb(n2510),.dout(n2520),.clk(gclk));
	jand g2442(.dina(w_n374_1[2]),.dinb(w_n343_1[0]),.dout(n2521),.clk(gclk));
	jand g2443(.dina(w_n2521_1[1]),.dinb(w_n597_1[0]),.dout(n2522),.clk(gclk));
	jand g2444(.dina(n2522),.dinb(w_n938_0[1]),.dout(n2523),.clk(gclk));
	jand g2445(.dina(w_n368_1[1]),.dinb(w_n267_0[1]),.dout(n2524),.clk(gclk));
	jand g2446(.dina(n2524),.dinb(w_n410_1[0]),.dout(n2525),.clk(gclk));
	jand g2447(.dina(w_n665_1[0]),.dinb(w_n614_1[1]),.dout(n2526),.clk(gclk));
	jand g2448(.dina(n2526),.dinb(w_n305_0[0]),.dout(n2527),.clk(gclk));
	jand g2449(.dina(n2527),.dinb(n2525),.dout(n2528),.clk(gclk));
	jand g2450(.dina(n2528),.dinb(n2523),.dout(n2529),.clk(gclk));
	jand g2451(.dina(w_n2498_0[0]),.dinb(w_n622_0[2]),.dout(n2530),.clk(gclk));
	jand g2452(.dina(n2530),.dinb(n2529),.dout(n2531),.clk(gclk));
	jand g2453(.dina(n2531),.dinb(w_n497_0[2]),.dout(n2532),.clk(gclk));
	jand g2454(.dina(n2532),.dinb(w_n832_1[0]),.dout(n2533),.clk(gclk));
	jand g2455(.dina(n2533),.dinb(w_n2520_0[2]),.dout(n2534),.clk(gclk));
	jor g2456(.dina(w_n2534_0[1]),.dinb(w_n2506_0[1]),.dout(n2535),.clk(gclk));
	jxor g2457(.dina(w_n2241_0[0]),.dinb(w_n2240_0[0]),.dout(n2536),.clk(gclk));
	jand g2458(.dina(w_n825_1[0]),.dinb(w_n310_0[2]),.dout(n2537),.clk(gclk));
	jand g2459(.dina(w_n765_0[2]),.dinb(w_n251_1[2]),.dout(n2538),.clk(gclk));
	jand g2460(.dina(w_n2538_0[1]),.dinb(w_n918_1[2]),.dout(n2539),.clk(gclk));
	jand g2461(.dina(n2539),.dinb(n2537),.dout(n2540),.clk(gclk));
	jand g2462(.dina(w_n1210_0[0]),.dinb(w_n730_0[1]),.dout(n2541),.clk(gclk));
	jand g2463(.dina(w_n853_1[0]),.dinb(w_n312_2[0]),.dout(n2542),.clk(gclk));
	jand g2464(.dina(w_n2542_0[1]),.dinb(w_n157_0[2]),.dout(n2543),.clk(gclk));
	jand g2465(.dina(n2543),.dinb(w_n2541_0[1]),.dout(n2544),.clk(gclk));
	jand g2466(.dina(w_n353_0[0]),.dinb(w_n220_1[0]),.dout(n2545),.clk(gclk));
	jor g2467(.dina(n2545),.dinb(w_n748_0[1]),.dout(n2546),.clk(gclk));
	jnot g2468(.din(n2546),.dout(n2547),.clk(gclk));
	jand g2469(.dina(w_n732_1[1]),.dinb(w_n451_1[2]),.dout(n2548),.clk(gclk));
	jand g2470(.dina(n2548),.dinb(n2547),.dout(n2549),.clk(gclk));
	jand g2471(.dina(n2549),.dinb(w_n2544_0[1]),.dout(n2550),.clk(gclk));
	jand g2472(.dina(n2550),.dinb(w_n2540_0[1]),.dout(n2551),.clk(gclk));
	jand g2473(.dina(w_n291_1[1]),.dinb(w_n254_1[2]),.dout(n2552),.clk(gclk));
	jand g2474(.dina(w_n2552_0[1]),.dinb(w_n2515_0[1]),.dout(n2553),.clk(gclk));
	jand g2475(.dina(n2553),.dinb(w_n646_0[0]),.dout(n2554),.clk(gclk));
	jand g2476(.dina(w_n878_1[0]),.dinb(w_n243_2[0]),.dout(n2555),.clk(gclk));
	jand g2477(.dina(w_n430_1[1]),.dinb(w_n303_2[0]),.dout(n2556),.clk(gclk));
	jand g2478(.dina(n2556),.dinb(n2555),.dout(n2557),.clk(gclk));
	jand g2479(.dina(w_n751_1[2]),.dinb(w_n763_1[0]),.dout(n2558),.clk(gclk));
	jand g2480(.dina(n2558),.dinb(w_n626_0[2]),.dout(n2559),.clk(gclk));
	jand g2481(.dina(n2559),.dinb(n2557),.dout(n2560),.clk(gclk));
	jand g2482(.dina(n2560),.dinb(w_n942_0[1]),.dout(n2561),.clk(gclk));
	jand g2483(.dina(n2561),.dinb(n2554),.dout(n2562),.clk(gclk));
	jand g2484(.dina(n2562),.dinb(w_n2427_0[1]),.dout(n2563),.clk(gclk));
	jand g2485(.dina(n2563),.dinb(w_n2551_0[1]),.dout(n2564),.clk(gclk));
	jor g2486(.dina(w_n2564_0[1]),.dinb(w_n2536_0[1]),.dout(n2565),.clk(gclk));
	jxor g2487(.dina(w_n2238_0[0]),.dinb(w_n1964_0[0]),.dout(n2566),.clk(gclk));
	jand g2488(.dina(w_n1189_0[2]),.dinb(w_n385_0[2]),.dout(n2567),.clk(gclk));
	jand g2489(.dina(w_n2315_0[0]),.dinb(w_n611_0[2]),.dout(n2568),.clk(gclk));
	jand g2490(.dina(n2568),.dinb(n2567),.dout(n2569),.clk(gclk));
	jand g2491(.dina(w_n2286_0[0]),.dinb(w_n365_0[2]),.dout(n2570),.clk(gclk));
	jand g2492(.dina(n2570),.dinb(w_n1000_0[0]),.dout(n2571),.clk(gclk));
	jand g2493(.dina(w_n854_0[0]),.dinb(w_n515_1[0]),.dout(n2572),.clk(gclk));
	jand g2494(.dina(n2572),.dinb(w_n417_1[0]),.dout(n2573),.clk(gclk));
	jand g2495(.dina(n2573),.dinb(w_n2571_0[1]),.dout(n2574),.clk(gclk));
	jand g2496(.dina(n2574),.dinb(n2569),.dout(n2575),.clk(gclk));
	jand g2497(.dina(w_n1193_0[0]),.dinb(w_n439_0[0]),.dout(n2576),.clk(gclk));
	jand g2498(.dina(n2576),.dinb(w_n392_0[0]),.dout(n2577),.clk(gclk));
	jand g2499(.dina(w_n993_0[1]),.dinb(w_n216_2[0]),.dout(n2578),.clk(gclk));
	jand g2500(.dina(n2578),.dinb(w_n781_1[0]),.dout(n2579),.clk(gclk));
	jand g2501(.dina(w_n878_0[2]),.dinb(w_n563_0[1]),.dout(n2580),.clk(gclk));
	jand g2502(.dina(w_n2580_0[1]),.dinb(w_n987_0[2]),.dout(n2581),.clk(gclk));
	jand g2503(.dina(n2581),.dinb(n2579),.dout(n2582),.clk(gclk));
	jand g2504(.dina(n2582),.dinb(w_n513_0[0]),.dout(n2583),.clk(gclk));
	jand g2505(.dina(n2583),.dinb(n2577),.dout(n2584),.clk(gclk));
	jand g2506(.dina(n2584),.dinb(w_n2575_0[2]),.dout(n2585),.clk(gclk));
	jand g2507(.dina(n2585),.dinb(w_n2486_0[0]),.dout(n2586),.clk(gclk));
	jand g2508(.dina(w_n2586_0[1]),.dinb(w_n2566_0[1]),.dout(n2587),.clk(gclk));
	jnot g2509(.din(w_n2564_0[0]),.dout(n2588),.clk(gclk));
	jxor g2510(.dina(n2588),.dinb(w_n2536_0[0]),.dout(n2589),.clk(gclk));
	jor g2511(.dina(w_n2589_0[2]),.dinb(w_n2587_0[1]),.dout(n2590),.clk(gclk));
	jand g2512(.dina(n2590),.dinb(n2565),.dout(n2591),.clk(gclk));
	jnot g2513(.din(w_n2534_0[0]),.dout(n2592),.clk(gclk));
	jxor g2514(.dina(n2592),.dinb(w_n2506_0[0]),.dout(n2593),.clk(gclk));
	jor g2515(.dina(w_n2593_0[1]),.dinb(w_n2591_0[1]),.dout(n2594),.clk(gclk));
	jand g2516(.dina(n2594),.dinb(n2535),.dout(n2595),.clk(gclk));
	jnot g2517(.din(w_n2504_0[1]),.dout(n2596),.clk(gclk));
	jxor g2518(.dina(n2596),.dinb(w_n2479_0[1]),.dout(n2597),.clk(gclk));
	jor g2519(.dina(n2597),.dinb(w_n2595_0[1]),.dout(n2598),.clk(gclk));
	jand g2520(.dina(n2598),.dinb(n2505),.dout(n2599),.clk(gclk));
	jxor g2521(.dina(w_n2477_0[0]),.dinb(w_n2440_0[0]),.dout(n2600),.clk(gclk));
	jnot g2522(.din(w_n2600_0[1]),.dout(n2601),.clk(gclk));
	jor g2523(.dina(n2601),.dinb(w_n2599_0[1]),.dout(n2602),.clk(gclk));
	jand g2524(.dina(n2602),.dinb(n2478),.dout(n2603),.clk(gclk));
	jxor g2525(.dina(w_n2438_0[0]),.dinb(w_n2414_0[0]),.dout(n2604),.clk(gclk));
	jnot g2526(.din(w_n2604_0[1]),.dout(n2605),.clk(gclk));
	jor g2527(.dina(w_n2605_0[1]),.dinb(w_n2603_0[2]),.dout(n2606),.clk(gclk));
	jand g2528(.dina(n2606),.dinb(n2439),.dout(n2607),.clk(gclk));
	jxor g2529(.dina(w_n2412_0[0]),.dinb(w_n2379_0[0]),.dout(n2608),.clk(gclk));
	jnot g2530(.din(w_n2608_0[1]),.dout(n2609),.clk(gclk));
	jor g2531(.dina(n2609),.dinb(w_n2607_0[1]),.dout(n2610),.clk(gclk));
	jand g2532(.dina(n2610),.dinb(n2413),.dout(n2611),.clk(gclk));
	jxor g2533(.dina(w_n2377_0[0]),.dinb(w_n2347_0[0]),.dout(n2612),.clk(gclk));
	jnot g2534(.din(w_n2612_0[1]),.dout(n2613),.clk(gclk));
	jor g2535(.dina(n2613),.dinb(w_n2611_0[1]),.dout(n2614),.clk(gclk));
	jand g2536(.dina(n2614),.dinb(n2378),.dout(n2615),.clk(gclk));
	jnot g2537(.din(w_n2615_0[1]),.dout(n2616),.clk(gclk));
	jxor g2538(.dina(w_n2345_0[0]),.dinb(w_n2302_0[0]),.dout(n2617),.clk(gclk));
	jand g2539(.dina(w_n2617_0[1]),.dinb(n2616),.dout(n2618),.clk(gclk));
	jnot g2540(.din(n2618),.dout(n2619),.clk(gclk));
	jand g2541(.dina(n2619),.dinb(n2346),.dout(n2620),.clk(gclk));
	jxor g2542(.dina(w_n2300_0[0]),.dinb(w_n2285_0[0]),.dout(n2621),.clk(gclk));
	jnot g2543(.din(w_n2621_0[1]),.dout(n2622),.clk(gclk));
	jor g2544(.dina(n2622),.dinb(w_n2620_0[1]),.dout(n2623),.clk(gclk));
	jand g2545(.dina(n2623),.dinb(n2301),.dout(n2624),.clk(gclk));
	jand g2546(.dina(w_n2283_0[0]),.dinb(w_n2267_0[0]),.dout(n2625),.clk(gclk));
	jand g2547(.dina(w_n2284_0[0]),.dinb(w_n2264_0[0]),.dout(n2626),.clk(gclk));
	jor g2548(.dina(n2626),.dinb(n2625),.dout(n2627),.clk(gclk));
	jand g2549(.dina(w_n2278_0[0]),.dinb(w_n2270_0[0]),.dout(n2628),.clk(gclk));
	jand g2550(.dina(w_n2282_0[0]),.dinb(w_n2279_0[0]),.dout(n2629),.clk(gclk));
	jor g2551(.dina(n2629),.dinb(n2628),.dout(n2630),.clk(gclk));
	jand g2552(.dina(w_n2281_0[0]),.dinb(w_n2280_0[0]),.dout(n2632),.clk(gclk));
	jor g2553(.dina(n2632),.dinb(w_n1114_0[0]),.dout(n2633),.clk(gclk));
	jand g2554(.dina(w_n960_2[0]),.dinb(w_n335_2[2]),.dout(n2634),.clk(gclk));
	jand g2555(.dina(w_n954_20[1]),.dinb(w_n795_0[1]),.dout(n2635),.clk(gclk));
	jor g2556(.dina(n2635),.dinb(w_n335_2[1]),.dout(n2636),.clk(gclk));
	jand g2557(.dina(w_n954_20[0]),.dinb(w_n804_1[0]),.dout(n2637),.clk(gclk));
	jnot g2558(.din(n2637),.dout(n2638),.clk(gclk));
	jand g2559(.dina(n2638),.dinb(n2636),.dout(n2639),.clk(gclk));
	jnot g2560(.din(n2639),.dout(n2640),.clk(gclk));
	jxor g2561(.dina(w_n2640_0[1]),.dinb(w_n2634_0[1]),.dout(n2641),.clk(gclk));
	jxor g2562(.dina(w_n2641_0[1]),.dinb(w_n2633_0[1]),.dout(n2642),.clk(gclk));
	jxor g2563(.dina(w_n2642_0[1]),.dinb(w_n2630_0[1]),.dout(n2643),.clk(gclk));
	jxor g2564(.dina(w_n2643_0[1]),.dinb(w_n2627_0[1]),.dout(n2644),.clk(gclk));
	jand g2565(.dina(w_n936_0[1]),.dinb(w_n158_0[1]),.dout(n2645),.clk(gclk));
	jand g2566(.dina(w_n1022_0[0]),.dinb(w_n280_1[0]),.dout(n2646),.clk(gclk));
	jand g2567(.dina(n2646),.dinb(n2645),.dout(n2647),.clk(gclk));
	jand g2568(.dina(w_n614_1[0]),.dinb(w_n422_1[2]),.dout(n2648),.clk(gclk));
	jand g2569(.dina(w_n374_1[1]),.dinb(w_n294_1[1]),.dout(n2649),.clk(gclk));
	jand g2570(.dina(n2649),.dinb(n2648),.dout(n2650),.clk(gclk));
	jand g2571(.dina(n2650),.dinb(w_n2321_0[1]),.dout(n2651),.clk(gclk));
	jand g2572(.dina(n2651),.dinb(n2647),.dout(n2652),.clk(gclk));
	jand g2573(.dina(n2652),.dinb(w_n482_0[0]),.dout(n2653),.clk(gclk));
	jand g2574(.dina(n2653),.dinb(w_n2365_0[1]),.dout(n2654),.clk(gclk));
	jand g2575(.dina(w_n781_0[2]),.dinb(w_n709_0[1]),.dout(n2655),.clk(gclk));
	jand g2576(.dina(w_n642_0[1]),.dinb(w_n436_1[1]),.dout(n2656),.clk(gclk));
	jand g2577(.dina(n2656),.dinb(w_n2380_2[1]),.dout(n2657),.clk(gclk));
	jand g2578(.dina(n2657),.dinb(w_n2655_0[1]),.dout(n2658),.clk(gclk));
	jand g2579(.dina(w_n624_1[1]),.dinb(w_n535_0[2]),.dout(n2659),.clk(gclk));
	jand g2580(.dina(n2659),.dinb(w_n563_0[0]),.dout(n2660),.clk(gclk));
	jand g2581(.dina(w_n363_1[0]),.dinb(w_n214_2[0]),.dout(n2661),.clk(gclk));
	jand g2582(.dina(n2661),.dinb(w_n388_0[0]),.dout(n2662),.clk(gclk));
	jand g2583(.dina(n2662),.dinb(w_n428_0[0]),.dout(n2663),.clk(gclk));
	jand g2584(.dina(n2663),.dinb(n2660),.dout(n2664),.clk(gclk));
	jand g2585(.dina(n2664),.dinb(w_n2658_0[1]),.dout(n2665),.clk(gclk));
	jand g2586(.dina(w_n2665_0[1]),.dinb(w_n2575_0[1]),.dout(n2666),.clk(gclk));
	jand g2587(.dina(n2666),.dinb(n2654),.dout(n2667),.clk(gclk));
	jxor g2588(.dina(w_n2667_0[1]),.dinb(w_n2644_0[1]),.dout(n2668),.clk(gclk));
	jxor g2589(.dina(w_n2668_0[1]),.dinb(w_n2624_0[1]),.dout(n2669),.clk(gclk));
	jnot g2590(.din(w_n2669_3[2]),.dout(n2670),.clk(gclk));
	jxor g2591(.dina(w_n2621_0[0]),.dinb(w_n2620_0[0]),.dout(n2671),.clk(gclk));
	jnot g2592(.din(w_n2671_6[1]),.dout(n2672),.clk(gclk));
	jand g2593(.dina(w_n2672_2[2]),.dinb(w_n2670_5[2]),.dout(n2673),.clk(gclk));
	jxor g2594(.dina(w_n2617_0[0]),.dinb(w_n2615_0[0]),.dout(n2674),.clk(gclk));
	jor g2595(.dina(w_n2674_4[1]),.dinb(w_n2671_6[0]),.dout(n2675),.clk(gclk));
	jnot g2596(.din(n2675),.dout(n2676),.clk(gclk));
	jnot g2597(.din(w_n2674_4[0]),.dout(n2677),.clk(gclk));
	jxor g2598(.dina(w_n2612_0[0]),.dinb(w_n2611_0[0]),.dout(n2678),.clk(gclk));
	jnot g2599(.din(w_n2678_6[1]),.dout(n2679),.clk(gclk));
	jand g2600(.dina(w_n2679_3[1]),.dinb(w_n2677_4[2]),.dout(n2680),.clk(gclk));
	jxor g2601(.dina(w_n2608_0[0]),.dinb(w_n2607_0[0]),.dout(n2681),.clk(gclk));
	jor g2602(.dina(w_n2681_5[1]),.dinb(w_n2678_6[0]),.dout(n2682),.clk(gclk));
	jnot g2603(.din(n2682),.dout(n2683),.clk(gclk));
	jnot g2604(.din(w_n2681_5[0]),.dout(n2684),.clk(gclk));
	jxor g2605(.dina(w_n2605_0[0]),.dinb(w_n2603_0[1]),.dout(n2685),.clk(gclk));
	jand g2606(.dina(w_n2685_2[1]),.dinb(w_n2684_4[1]),.dout(n2686),.clk(gclk));
	jxor g2607(.dina(w_n2604_0[0]),.dinb(w_n2603_0[0]),.dout(n2687),.clk(gclk));
	jxor g2608(.dina(w_n2600_0[0]),.dinb(w_n2599_0[0]),.dout(n2688),.clk(gclk));
	jor g2609(.dina(w_n2688_8[2]),.dinb(w_n2687_7[1]),.dout(n2689),.clk(gclk));
	jxor g2610(.dina(w_n2504_0[0]),.dinb(w_n2479_0[0]),.dout(n2690),.clk(gclk));
	jxor g2611(.dina(n2690),.dinb(w_n2595_0[0]),.dout(n2691),.clk(gclk));
	jor g2612(.dina(w_n2691_8[2]),.dinb(w_n2688_8[1]),.dout(n2692),.clk(gclk));
	jxor g2613(.dina(w_n2593_0[0]),.dinb(w_n2591_0[0]),.dout(n2693),.clk(gclk));
	jnot g2614(.din(w_n2693_4[2]),.dout(n2694),.clk(gclk));
	jor g2615(.dina(w_n2694_4[2]),.dinb(w_n2691_8[1]),.dout(n2695),.clk(gclk));
	jxor g2616(.dina(w_n2693_4[1]),.dinb(w_n2691_8[0]),.dout(n2696),.clk(gclk));
	jxor g2617(.dina(w_n2586_0[0]),.dinb(w_n2566_0[0]),.dout(n2697),.clk(gclk));
	jnot g2618(.din(w_n2697_1[1]),.dout(n2698),.clk(gclk));
	jor g2619(.dina(w_n2698_6[1]),.dinb(w_n2693_4[0]),.dout(n2699),.clk(gclk));
	jxor g2620(.dina(w_n2589_0[1]),.dinb(w_n2587_0[0]),.dout(n2700),.clk(gclk));
	jand g2621(.dina(w_n2700_5[2]),.dinb(n2699),.dout(n2701),.clk(gclk));
	jnot g2622(.din(w_n2701_0[1]),.dout(n2702),.clk(gclk));
	jor g2623(.dina(w_n2702_0[1]),.dinb(w_n2696_0[2]),.dout(n2703),.clk(gclk));
	jand g2624(.dina(n2703),.dinb(n2695),.dout(n2704),.clk(gclk));
	jxor g2625(.dina(w_n2691_7[2]),.dinb(w_n2688_8[0]),.dout(n2705),.clk(gclk));
	jnot g2626(.din(w_n2705_0[1]),.dout(n2706),.clk(gclk));
	jor g2627(.dina(n2706),.dinb(w_n2704_0[1]),.dout(n2707),.clk(gclk));
	jand g2628(.dina(n2707),.dinb(n2692),.dout(n2708),.clk(gclk));
	jxor g2629(.dina(w_n2688_7[2]),.dinb(w_n2685_2[0]),.dout(n2709),.clk(gclk));
	jor g2630(.dina(n2709),.dinb(w_n2708_0[1]),.dout(n2710),.clk(gclk));
	jand g2631(.dina(n2710),.dinb(n2689),.dout(n2711),.clk(gclk));
	jnot g2632(.din(w_n2711_0[1]),.dout(n2712),.clk(gclk));
	jxor g2633(.dina(w_n2687_7[0]),.dinb(w_n2681_4[2]),.dout(n2713),.clk(gclk));
	jand g2634(.dina(w_n2713_0[1]),.dinb(n2712),.dout(n2714),.clk(gclk));
	jor g2635(.dina(n2714),.dinb(n2686),.dout(n2715),.clk(gclk));
	jxor g2636(.dina(w_n2681_4[1]),.dinb(w_n2678_5[2]),.dout(n2716),.clk(gclk));
	jand g2637(.dina(n2716),.dinb(w_n2715_0[1]),.dout(n2717),.clk(gclk));
	jor g2638(.dina(n2717),.dinb(n2683),.dout(n2718),.clk(gclk));
	jxor g2639(.dina(w_n2678_5[1]),.dinb(w_n2674_3[2]),.dout(n2719),.clk(gclk));
	jand g2640(.dina(w_n2719_0[1]),.dinb(w_n2718_0[1]),.dout(n2720),.clk(gclk));
	jor g2641(.dina(n2720),.dinb(n2680),.dout(n2721),.clk(gclk));
	jxor g2642(.dina(w_n2674_3[1]),.dinb(w_n2671_5[2]),.dout(n2722),.clk(gclk));
	jand g2643(.dina(w_n2722_0[1]),.dinb(w_n2721_0[1]),.dout(n2723),.clk(gclk));
	jor g2644(.dina(n2723),.dinb(n2676),.dout(n2724),.clk(gclk));
	jxor g2645(.dina(w_n2671_5[1]),.dinb(w_n2669_3[1]),.dout(n2725),.clk(gclk));
	jand g2646(.dina(w_n2725_0[1]),.dinb(w_n2724_0[1]),.dout(n2726),.clk(gclk));
	jor g2647(.dina(n2726),.dinb(n2673),.dout(n2727),.clk(gclk));
	jnot g2648(.din(w_n2727_0[1]),.dout(n2728),.clk(gclk));
	jor g2649(.dina(w_n2667_0[0]),.dinb(w_n2644_0[0]),.dout(n2729),.clk(gclk));
	jnot g2650(.din(n2729),.dout(n2730),.clk(gclk));
	jnot g2651(.din(w_n2624_0[0]),.dout(n2731),.clk(gclk));
	jand g2652(.dina(w_n2668_0[0]),.dinb(n2731),.dout(n2732),.clk(gclk));
	jor g2653(.dina(n2732),.dinb(n2730),.dout(n2733),.clk(gclk));
	jand g2654(.dina(w_n458_0[2]),.dinb(w_n153_1[0]),.dout(n2734),.clk(gclk));
	jand g2655(.dina(w_n2734_0[2]),.dinb(w_n597_0[2]),.dout(n2735),.clk(gclk));
	jand g2656(.dina(w_n925_0[2]),.dinb(w_n410_0[2]),.dout(n2736),.clk(gclk));
	jand g2657(.dina(w_n2736_1[1]),.dinb(w_n731_0[1]),.dout(n2737),.clk(gclk));
	jand g2658(.dina(w_n2552_0[0]),.dinb(w_n992_1[0]),.dout(n2738),.clk(gclk));
	jand g2659(.dina(n2738),.dinb(n2737),.dout(n2739),.clk(gclk));
	jand g2660(.dina(n2739),.dinb(n2735),.dout(n2740),.clk(gclk));
	jand g2661(.dina(w_n2380_2[0]),.dinb(w_n279_1[0]),.dout(n2741),.clk(gclk));
	jand g2662(.dina(n2741),.dinb(w_n470_0[1]),.dout(n2742),.clk(gclk));
	jand g2663(.dina(n2742),.dinb(w_n2323_0[0]),.dout(n2743),.clk(gclk));
	jand g2664(.dina(w_n935_1[2]),.dinb(w_n633_0[0]),.dout(n2744),.clk(gclk));
	jand g2665(.dina(n2744),.dinb(w_n2351_0[0]),.dout(n2745),.clk(gclk));
	jand g2666(.dina(w_n2745_0[1]),.dinb(w_n2743_0[1]),.dout(n2746),.clk(gclk));
	jand g2667(.dina(n2746),.dinb(n2740),.dout(n2747),.clk(gclk));
	jand g2668(.dina(w_n1231_0[1]),.dinb(w_n497_0[1]),.dout(n2748),.clk(gclk));
	jand g2669(.dina(n2748),.dinb(n2747),.dout(n2749),.clk(gclk));
	jand g2670(.dina(n2749),.dinb(w_n2451_0[0]),.dout(n2750),.clk(gclk));
	jxor g2671(.dina(w_n960_1[2]),.dinb(w_n820_3[2]),.dout(n2751),.clk(gclk));
	jnot g2672(.din(w_n2751_0[1]),.dout(n2752),.clk(gclk));
	jand g2673(.dina(w_n2752_0[2]),.dinb(n796),.dout(n2753),.clk(gclk));
	jnot g2674(.din(n2753),.dout(n2754),.clk(gclk));
	jand g2675(.dina(w_n335_2[0]),.dinb(n2754),.dout(n2757),.clk(gclk));
	jand g2676(.dina(w_n2642_0[0]),.dinb(w_n2630_0[0]),.dout(n2758),.clk(gclk));
	jand g2677(.dina(w_n2643_0[0]),.dinb(w_n2627_0[0]),.dout(n2759),.clk(gclk));
	jor g2678(.dina(n2759),.dinb(n2758),.dout(n2760),.clk(gclk));
	jor g2679(.dina(w_n2640_0[0]),.dinb(w_n2634_0[0]),.dout(n2761),.clk(gclk));
	jnot g2680(.din(w_n2633_0[0]),.dout(n2762),.clk(gclk));
	jnot g2681(.din(w_n2641_0[0]),.dout(n2763),.clk(gclk));
	jor g2682(.dina(n2763),.dinb(n2762),.dout(n2764),.clk(gclk));
	jand g2683(.dina(n2764),.dinb(n2761),.dout(n2765),.clk(gclk));
	jxor g2684(.dina(n2765),.dinb(n2760),.dout(n2766),.clk(gclk));
	jxor g2685(.dina(n2766),.dinb(n2757),.dout(n2767),.clk(gclk));
	jxor g2686(.dina(w_n2767_0[2]),.dinb(w_n2750_0[2]),.dout(n2768),.clk(gclk));
	jxor g2687(.dina(n2768),.dinb(w_n2733_0[1]),.dout(n2769),.clk(gclk));
	jxor g2688(.dina(w_n2769_4[1]),.dinb(w_n2670_5[1]),.dout(n2770),.clk(gclk));
	jxor g2689(.dina(w_n2770_0[2]),.dinb(n2728),.dout(n2771),.clk(gclk));
	jor g2690(.dina(w_n2771_1[2]),.dinb(w_n79_6[1]),.dout(n2772),.clk(gclk));
	jnot g2691(.din(w_n2769_4[0]),.dout(n2773),.clk(gclk));
	jand g2692(.dina(w_n76_0[0]),.dinb(w_n70_0[1]),.dout(n2774),.clk(gclk));
	jnot g2693(.din(w_n2774_2[1]),.dout(n2775),.clk(gclk));
	jor g2694(.dina(w_n2775_5[2]),.dinb(w_n2773_4[2]),.dout(n2776),.clk(gclk));
	jxor g2695(.dina(w_n75_1[2]),.dinb(w_n59_1[0]),.dout(n2777),.clk(gclk));
	jnot g2696(.din(w_n2777_0[1]),.dout(n2778),.clk(gclk));
	jand g2697(.dina(n2778),.dinb(w_n69_0[1]),.dout(n2779),.clk(gclk));
	jnot g2698(.din(w_n2779_2[2]),.dout(n2780),.clk(gclk));
	jor g2699(.dina(w_n2780_5[2]),.dinb(w_n2669_3[0]),.dout(n2781),.clk(gclk));
	jand g2700(.dina(w_n77_0[0]),.dinb(w_n69_0[0]),.dout(n2782),.clk(gclk));
	jand g2701(.dina(n2782),.dinb(w_n2777_0[0]),.dout(n2783),.clk(gclk));
	jnot g2702(.din(w_n2783_2[1]),.dout(n2784),.clk(gclk));
	jor g2703(.dina(w_n2784_6[1]),.dinb(w_n2671_5[0]),.dout(n2785),.clk(gclk));
	jand g2704(.dina(n2785),.dinb(n2781),.dout(n2786),.clk(gclk));
	jand g2705(.dina(n2786),.dinb(n2776),.dout(n2787),.clk(gclk));
	jand g2706(.dina(n2787),.dinb(n2772),.dout(n2788),.clk(gclk));
	jxor g2707(.dina(n2788),.dinb(w_n56_8[2]),.dout(n2789),.clk(gclk));
	jxor g2708(.dina(w_n1347_2[1]),.dinb(w_n56_8[1]),.dout(n2790),.clk(gclk));
	jnot g2709(.din(w_n2790_0[2]),.dout(n2791),.clk(gclk));
	jxor g2710(.dina(w_n699_9[2]),.dinb(w_n1391_2[0]),.dout(n2792),.clk(gclk));
	jnot g2711(.din(w_n2792_0[1]),.dout(n2793),.clk(gclk));
	jand g2712(.dina(w_n2793_0[1]),.dinb(w_n2791_0[2]),.dout(n2794),.clk(gclk));
	jnot g2713(.din(w_n2794_2[2]),.dout(n2795),.clk(gclk));
	jxor g2714(.dina(w_n2684_4[0]),.dinb(w_n2678_5[0]),.dout(n2796),.clk(gclk));
	jxor g2715(.dina(n2796),.dinb(w_n2715_0[0]),.dout(n2797),.clk(gclk));
	jor g2716(.dina(w_n2797_1[2]),.dinb(w_n2795_6[1]),.dout(n2798),.clk(gclk));
	jand g2717(.dina(w_n2792_0[0]),.dinb(w_n2791_0[1]),.dout(n2799),.clk(gclk));
	jnot g2718(.din(w_n2799_2[1]),.dout(n2800),.clk(gclk));
	jor g2719(.dina(w_n2800_5[2]),.dinb(w_n2678_4[2]),.dout(n2801),.clk(gclk));
	jxor g2720(.dina(w_n1347_2[0]),.dinb(w_n1391_1[2]),.dout(n2802),.clk(gclk));
	jnot g2721(.din(w_n2802_0[1]),.dout(n2803),.clk(gclk));
	jand g2722(.dina(n2803),.dinb(w_n2790_0[1]),.dout(n2804),.clk(gclk));
	jnot g2723(.din(w_n2804_2[2]),.dout(n2805),.clk(gclk));
	jor g2724(.dina(w_n2805_5[2]),.dinb(w_n2681_4[0]),.dout(n2806),.clk(gclk));
	jand g2725(.dina(w_n2802_0[0]),.dinb(w_n2790_0[0]),.dout(n2807),.clk(gclk));
	jand g2726(.dina(n2807),.dinb(w_n2793_0[0]),.dout(n2808),.clk(gclk));
	jnot g2727(.din(w_n2808_2[1]),.dout(n2809),.clk(gclk));
	jor g2728(.dina(w_n2809_6[1]),.dinb(w_n2687_6[2]),.dout(n2810),.clk(gclk));
	jand g2729(.dina(n2810),.dinb(n2806),.dout(n2811),.clk(gclk));
	jand g2730(.dina(n2811),.dinb(n2801),.dout(n2812),.clk(gclk));
	jand g2731(.dina(n2812),.dinb(n2798),.dout(n2813),.clk(gclk));
	jxor g2732(.dina(n2813),.dinb(w_n699_9[1]),.dout(n2814),.clk(gclk));
	jnot g2733(.din(n2814),.dout(n2815),.clk(gclk));
	jxor g2734(.dina(w_n980_2[1]),.dinb(w_n808_10[0]),.dout(n2816),.clk(gclk));
	jnot g2735(.din(w_n2816_0[2]),.dout(n2817),.clk(gclk));
	jand g2736(.dina(w_n2817_1[1]),.dinb(w_n2698_6[0]),.dout(n2818),.clk(gclk));
	jor g2737(.dina(w_n2700_5[1]),.dinb(w_n2697_1[0]),.dout(n2819),.clk(gclk));
	jand g2738(.dina(w_n2697_0[2]),.dinb(w_n2589_0[0]),.dout(n2820),.clk(gclk));
	jnot g2739(.din(n2820),.dout(n2821),.clk(gclk));
	jand g2740(.dina(w_n2821_0[1]),.dinb(n2819),.dout(n2822),.clk(gclk));
	jnot g2741(.din(w_n2822_0[1]),.dout(n2823),.clk(gclk));
	jxor g2742(.dina(w_n1059_2[0]),.dinb(w_n699_9[0]),.dout(n2824),.clk(gclk));
	jnot g2743(.din(w_n2824_0[2]),.dout(n2825),.clk(gclk));
	jxor g2744(.dina(w_n808_9[2]),.dinb(w_n708_2[1]),.dout(n2826),.clk(gclk));
	jnot g2745(.din(w_n2826_0[1]),.dout(n2827),.clk(gclk));
	jand g2746(.dina(w_n2827_0[1]),.dinb(w_n2825_0[2]),.dout(n2828),.clk(gclk));
	jand g2747(.dina(w_n2828_2[2]),.dinb(w_n2823_1[1]),.dout(n2829),.clk(gclk));
	jxor g2748(.dina(w_n1059_1[2]),.dinb(w_n708_2[0]),.dout(n2830),.clk(gclk));
	jnot g2749(.din(w_n2830_0[1]),.dout(n2831),.clk(gclk));
	jand g2750(.dina(n2831),.dinb(w_n2824_0[1]),.dout(n2832),.clk(gclk));
	jand g2751(.dina(w_n2832_2[2]),.dinb(w_n2698_5[2]),.dout(n2833),.clk(gclk));
	jand g2752(.dina(w_n2826_0[0]),.dinb(w_n2825_0[1]),.dout(n2834),.clk(gclk));
	jand g2753(.dina(w_n2834_2[1]),.dinb(w_n2700_5[0]),.dout(n2835),.clk(gclk));
	jor g2754(.dina(n2835),.dinb(n2833),.dout(n2836),.clk(gclk));
	jor g2755(.dina(n2836),.dinb(n2829),.dout(n2837),.clk(gclk));
	jnot g2756(.din(w_n2837_0[1]),.dout(n2838),.clk(gclk));
	jand g2757(.dina(w_n2825_0[0]),.dinb(w_n2698_5[1]),.dout(n2839),.clk(gclk));
	jnot g2758(.din(w_n2839_1[1]),.dout(n2840),.clk(gclk));
	jand g2759(.dina(n2840),.dinb(w_n803_4[2]),.dout(n2841),.clk(gclk));
	jand g2760(.dina(n2841),.dinb(n2838),.dout(n2842),.clk(gclk));
	jxor g2761(.dina(w_n2821_0[0]),.dinb(w_n2693_3[2]),.dout(n2843),.clk(gclk));
	jnot g2762(.din(n2843),.dout(n2844),.clk(gclk));
	jand g2763(.dina(w_n2844_1[1]),.dinb(w_n2828_2[1]),.dout(n2845),.clk(gclk));
	jand g2764(.dina(w_n2834_2[0]),.dinb(w_n2693_3[1]),.dout(n2846),.clk(gclk));
	jand g2765(.dina(w_n2830_0[0]),.dinb(w_n2824_0[0]),.dout(n2847),.clk(gclk));
	jand g2766(.dina(n2847),.dinb(w_n2827_0[0]),.dout(n2848),.clk(gclk));
	jand g2767(.dina(w_n2848_2[1]),.dinb(w_n2698_5[0]),.dout(n2849),.clk(gclk));
	jand g2768(.dina(w_n2832_2[1]),.dinb(w_n2700_4[2]),.dout(n2850),.clk(gclk));
	jor g2769(.dina(n2850),.dinb(n2849),.dout(n2851),.clk(gclk));
	jor g2770(.dina(n2851),.dinb(n2846),.dout(n2852),.clk(gclk));
	jor g2771(.dina(n2852),.dinb(n2845),.dout(n2853),.clk(gclk));
	jnot g2772(.din(n2853),.dout(n2854),.clk(gclk));
	jand g2773(.dina(w_n2854_0[1]),.dinb(w_n2842_0[1]),.dout(n2855),.clk(gclk));
	jand g2774(.dina(w_n2855_0[1]),.dinb(w_n2818_0[2]),.dout(n2856),.clk(gclk));
	jnot g2775(.din(w_n2828_2[0]),.dout(n2857),.clk(gclk));
	jxor g2776(.dina(w_n2701_0[0]),.dinb(w_n2696_0[1]),.dout(n2858),.clk(gclk));
	jor g2777(.dina(w_n2858_1[2]),.dinb(w_n2857_6[1]),.dout(n2859),.clk(gclk));
	jnot g2778(.din(w_n2834_1[2]),.dout(n2860),.clk(gclk));
	jor g2779(.dina(w_n2860_5[2]),.dinb(w_n2691_7[1]),.dout(n2861),.clk(gclk));
	jnot g2780(.din(w_n2700_4[1]),.dout(n2862),.clk(gclk));
	jnot g2781(.din(w_n2848_2[0]),.dout(n2863),.clk(gclk));
	jor g2782(.dina(w_n2863_6[1]),.dinb(w_n2862_2[2]),.dout(n2864),.clk(gclk));
	jnot g2783(.din(w_n2832_2[0]),.dout(n2865),.clk(gclk));
	jor g2784(.dina(w_n2865_5[2]),.dinb(w_n2694_4[1]),.dout(n2866),.clk(gclk));
	jand g2785(.dina(n2866),.dinb(n2864),.dout(n2867),.clk(gclk));
	jand g2786(.dina(n2867),.dinb(n2861),.dout(n2868),.clk(gclk));
	jand g2787(.dina(n2868),.dinb(n2859),.dout(n2869),.clk(gclk));
	jxor g2788(.dina(n2869),.dinb(w_n808_9[1]),.dout(n2870),.clk(gclk));
	jxor g2789(.dina(w_n2855_0[0]),.dinb(w_n2818_0[1]),.dout(n2871),.clk(gclk));
	jand g2790(.dina(w_n2871_0[1]),.dinb(w_n2870_0[1]),.dout(n2872),.clk(gclk));
	jor g2791(.dina(n2872),.dinb(n2856),.dout(n2873),.clk(gclk));
	jxor g2792(.dina(w_n2705_0[0]),.dinb(w_n2704_0[0]),.dout(n2874),.clk(gclk));
	jor g2793(.dina(w_n2874_1[2]),.dinb(w_n2857_6[0]),.dout(n2875),.clk(gclk));
	jor g2794(.dina(w_n2860_5[1]),.dinb(w_n2688_7[1]),.dout(n2876),.clk(gclk));
	jor g2795(.dina(w_n2865_5[1]),.dinb(w_n2691_7[0]),.dout(n2877),.clk(gclk));
	jor g2796(.dina(w_n2863_6[0]),.dinb(w_n2694_4[0]),.dout(n2878),.clk(gclk));
	jand g2797(.dina(n2878),.dinb(n2877),.dout(n2879),.clk(gclk));
	jand g2798(.dina(n2879),.dinb(n2876),.dout(n2880),.clk(gclk));
	jand g2799(.dina(n2880),.dinb(n2875),.dout(n2881),.clk(gclk));
	jxor g2800(.dina(n2881),.dinb(w_n808_9[0]),.dout(n2882),.clk(gclk));
	jand g2801(.dina(w_n2817_1[0]),.dinb(w_n2752_0[1]),.dout(n2883),.clk(gclk));
	jand g2802(.dina(w_n2883_3[1]),.dinb(w_n2823_1[0]),.dout(n2884),.clk(gclk));
	jxor g2803(.dina(w_n980_2[0]),.dinb(w_n961_1[2]),.dout(n2885),.clk(gclk));
	jnot g2804(.din(w_n2885_0[1]),.dout(n2886),.clk(gclk));
	jand g2805(.dina(n2886),.dinb(w_n2816_0[1]),.dout(n2887),.clk(gclk));
	jand g2806(.dina(w_n2887_4[2]),.dinb(w_n2698_4[2]),.dout(n2888),.clk(gclk));
	jand g2807(.dina(w_n2817_0[2]),.dinb(w_n2751_0[0]),.dout(n2889),.clk(gclk));
	jand g2808(.dina(w_n2889_4[1]),.dinb(w_n2700_4[0]),.dout(n2890),.clk(gclk));
	jor g2809(.dina(n2890),.dinb(n2888),.dout(n2891),.clk(gclk));
	jor g2810(.dina(n2891),.dinb(n2884),.dout(n2892),.clk(gclk));
	jand g2811(.dina(w_n2698_4[1]),.dinb(w_n954_19[2]),.dout(n2893),.clk(gclk));
	jand g2812(.dina(w_n2893_0[2]),.dinb(w_n2817_0[1]),.dout(n2894),.clk(gclk));
	jxor g2813(.dina(n2894),.dinb(w_n2892_0[1]),.dout(n2895),.clk(gclk));
	jxor g2814(.dina(w_n2895_0[1]),.dinb(w_n2882_0[1]),.dout(n2896),.clk(gclk));
	jxor g2815(.dina(w_n2896_0[1]),.dinb(w_n2873_0[1]),.dout(n2897),.clk(gclk));
	jand g2816(.dina(w_n2897_0[1]),.dinb(w_n2815_0[1]),.dout(n2898),.clk(gclk));
	jxor g2817(.dina(w_n2713_0[0]),.dinb(w_n2711_0[0]),.dout(n2899),.clk(gclk));
	jor g2818(.dina(w_n2899_1[2]),.dinb(w_n2795_6[0]),.dout(n2900),.clk(gclk));
	jor g2819(.dina(w_n2800_5[1]),.dinb(w_n2681_3[2]),.dout(n2901),.clk(gclk));
	jor g2820(.dina(w_n2805_5[1]),.dinb(w_n2687_6[1]),.dout(n2902),.clk(gclk));
	jor g2821(.dina(w_n2809_6[0]),.dinb(w_n2688_7[0]),.dout(n2903),.clk(gclk));
	jand g2822(.dina(n2903),.dinb(n2902),.dout(n2904),.clk(gclk));
	jand g2823(.dina(n2904),.dinb(n2901),.dout(n2905),.clk(gclk));
	jand g2824(.dina(n2905),.dinb(n2900),.dout(n2906),.clk(gclk));
	jxor g2825(.dina(n2906),.dinb(w_n1143_5[2]),.dout(n2907),.clk(gclk));
	jxor g2826(.dina(w_n2871_0[0]),.dinb(w_n2870_0[0]),.dout(n2908),.clk(gclk));
	jand g2827(.dina(w_n2908_0[1]),.dinb(w_n2907_0[1]),.dout(n2909),.clk(gclk));
	jxor g2828(.dina(w_n2688_6[2]),.dinb(w_n2687_6[0]),.dout(n2910),.clk(gclk));
	jxor g2829(.dina(n2910),.dinb(w_n2708_0[0]),.dout(n2911),.clk(gclk));
	jor g2830(.dina(w_n2911_1[2]),.dinb(w_n2795_5[2]),.dout(n2912),.clk(gclk));
	jor g2831(.dina(w_n2800_5[0]),.dinb(w_n2687_5[2]),.dout(n2913),.clk(gclk));
	jor g2832(.dina(w_n2805_5[0]),.dinb(w_n2688_6[1]),.dout(n2914),.clk(gclk));
	jor g2833(.dina(w_n2809_5[2]),.dinb(w_n2691_6[2]),.dout(n2915),.clk(gclk));
	jand g2834(.dina(n2915),.dinb(n2914),.dout(n2916),.clk(gclk));
	jand g2835(.dina(n2916),.dinb(n2913),.dout(n2917),.clk(gclk));
	jand g2836(.dina(n2917),.dinb(n2912),.dout(n2918),.clk(gclk));
	jxor g2837(.dina(n2918),.dinb(w_n699_8[2]),.dout(n2919),.clk(gclk));
	jnot g2838(.din(n2919),.dout(n2920),.clk(gclk));
	jor g2839(.dina(w_n2842_0[0]),.dinb(w_n808_8[2]),.dout(n2921),.clk(gclk));
	jxor g2840(.dina(n2921),.dinb(w_n2854_0[0]),.dout(n2922),.clk(gclk));
	jand g2841(.dina(w_n2922_0[1]),.dinb(w_n2920_0[1]),.dout(n2923),.clk(gclk));
	jor g2842(.dina(w_n2874_1[1]),.dinb(w_n2795_5[1]),.dout(n2924),.clk(gclk));
	jor g2843(.dina(w_n2800_4[2]),.dinb(w_n2688_6[0]),.dout(n2925),.clk(gclk));
	jor g2844(.dina(w_n2805_4[2]),.dinb(w_n2691_6[1]),.dout(n2926),.clk(gclk));
	jor g2845(.dina(w_n2809_5[1]),.dinb(w_n2694_3[2]),.dout(n2927),.clk(gclk));
	jand g2846(.dina(n2927),.dinb(n2926),.dout(n2928),.clk(gclk));
	jand g2847(.dina(n2928),.dinb(n2925),.dout(n2929),.clk(gclk));
	jand g2848(.dina(n2929),.dinb(n2924),.dout(n2930),.clk(gclk));
	jxor g2849(.dina(n2930),.dinb(w_n1143_5[1]),.dout(n2931),.clk(gclk));
	jand g2850(.dina(w_n2839_1[0]),.dinb(w_n803_4[1]),.dout(n2932),.clk(gclk));
	jxor g2851(.dina(n2932),.dinb(w_n2837_0[0]),.dout(n2933),.clk(gclk));
	jand g2852(.dina(w_n2933_0[1]),.dinb(w_n2931_0[1]),.dout(n2934),.clk(gclk));
	jand g2853(.dina(w_n2823_0[2]),.dinb(w_n2794_2[1]),.dout(n2935),.clk(gclk));
	jand g2854(.dina(w_n2804_2[1]),.dinb(w_n2698_4[0]),.dout(n2936),.clk(gclk));
	jand g2855(.dina(w_n2799_2[0]),.dinb(w_n2700_3[2]),.dout(n2937),.clk(gclk));
	jor g2856(.dina(n2937),.dinb(n2936),.dout(n2938),.clk(gclk));
	jor g2857(.dina(n2938),.dinb(n2935),.dout(n2939),.clk(gclk));
	jnot g2858(.din(w_n2939_0[1]),.dout(n2940),.clk(gclk));
	jand g2859(.dina(w_n2791_0[0]),.dinb(w_n2698_3[2]),.dout(n2941),.clk(gclk));
	jnot g2860(.din(w_n2941_1[1]),.dout(n2942),.clk(gclk));
	jand g2861(.dina(n2942),.dinb(w_n699_8[1]),.dout(n2943),.clk(gclk));
	jand g2862(.dina(n2943),.dinb(n2940),.dout(n2944),.clk(gclk));
	jand g2863(.dina(w_n2844_1[0]),.dinb(w_n2794_2[0]),.dout(n2945),.clk(gclk));
	jand g2864(.dina(w_n2799_1[2]),.dinb(w_n2693_3[0]),.dout(n2946),.clk(gclk));
	jand g2865(.dina(w_n2808_2[0]),.dinb(w_n2698_3[1]),.dout(n2947),.clk(gclk));
	jand g2866(.dina(w_n2804_2[0]),.dinb(w_n2700_3[1]),.dout(n2948),.clk(gclk));
	jor g2867(.dina(n2948),.dinb(n2947),.dout(n2949),.clk(gclk));
	jor g2868(.dina(n2949),.dinb(n2946),.dout(n2950),.clk(gclk));
	jor g2869(.dina(n2950),.dinb(n2945),.dout(n2951),.clk(gclk));
	jnot g2870(.din(n2951),.dout(n2952),.clk(gclk));
	jand g2871(.dina(w_n2952_0[1]),.dinb(w_n2944_0[1]),.dout(n2953),.clk(gclk));
	jand g2872(.dina(w_n2953_0[1]),.dinb(w_n2839_0[2]),.dout(n2954),.clk(gclk));
	jor g2873(.dina(w_n2858_1[1]),.dinb(w_n2795_5[0]),.dout(n2955),.clk(gclk));
	jor g2874(.dina(w_n2800_4[1]),.dinb(w_n2691_6[0]),.dout(n2956),.clk(gclk));
	jor g2875(.dina(w_n2809_5[0]),.dinb(w_n2862_2[1]),.dout(n2957),.clk(gclk));
	jor g2876(.dina(w_n2805_4[1]),.dinb(w_n2694_3[1]),.dout(n2958),.clk(gclk));
	jand g2877(.dina(n2958),.dinb(n2957),.dout(n2959),.clk(gclk));
	jand g2878(.dina(n2959),.dinb(n2956),.dout(n2960),.clk(gclk));
	jand g2879(.dina(n2960),.dinb(n2955),.dout(n2961),.clk(gclk));
	jxor g2880(.dina(n2961),.dinb(w_n699_8[0]),.dout(n2962),.clk(gclk));
	jnot g2881(.din(n2962),.dout(n2963),.clk(gclk));
	jxor g2882(.dina(w_n2953_0[0]),.dinb(w_n2839_0[1]),.dout(n2964),.clk(gclk));
	jand g2883(.dina(w_n2964_0[1]),.dinb(w_n2963_0[1]),.dout(n2965),.clk(gclk));
	jor g2884(.dina(n2965),.dinb(n2954),.dout(n2966),.clk(gclk));
	jxor g2885(.dina(w_n2933_0[0]),.dinb(w_n2931_0[0]),.dout(n2967),.clk(gclk));
	jand g2886(.dina(w_n2967_0[1]),.dinb(w_n2966_0[1]),.dout(n2968),.clk(gclk));
	jor g2887(.dina(n2968),.dinb(n2934),.dout(n2969),.clk(gclk));
	jxor g2888(.dina(w_n2922_0[0]),.dinb(w_n2920_0[0]),.dout(n2970),.clk(gclk));
	jand g2889(.dina(w_n2970_0[1]),.dinb(w_n2969_0[1]),.dout(n2971),.clk(gclk));
	jor g2890(.dina(n2971),.dinb(n2923),.dout(n2972),.clk(gclk));
	jxor g2891(.dina(w_n2908_0[0]),.dinb(w_n2907_0[0]),.dout(n2973),.clk(gclk));
	jand g2892(.dina(w_n2973_0[1]),.dinb(w_n2972_0[1]),.dout(n2974),.clk(gclk));
	jor g2893(.dina(n2974),.dinb(n2909),.dout(n2975),.clk(gclk));
	jxor g2894(.dina(w_n2897_0[0]),.dinb(w_n2815_0[0]),.dout(n2976),.clk(gclk));
	jand g2895(.dina(w_n2976_0[1]),.dinb(w_n2975_0[1]),.dout(n2977),.clk(gclk));
	jor g2896(.dina(n2977),.dinb(n2898),.dout(n2978),.clk(gclk));
	jand g2897(.dina(w_n2895_0[0]),.dinb(w_n2882_0[0]),.dout(n2979),.clk(gclk));
	jand g2898(.dina(w_n2896_0[0]),.dinb(w_n2873_0[0]),.dout(n2980),.clk(gclk));
	jor g2899(.dina(n2980),.dinb(n2979),.dout(n2981),.clk(gclk));
	jor g2900(.dina(w_n2911_1[1]),.dinb(w_n2857_5[2]),.dout(n2982),.clk(gclk));
	jor g2901(.dina(w_n2860_5[0]),.dinb(w_n2687_5[1]),.dout(n2983),.clk(gclk));
	jor g2902(.dina(w_n2865_5[0]),.dinb(w_n2688_5[2]),.dout(n2984),.clk(gclk));
	jor g2903(.dina(w_n2863_5[2]),.dinb(w_n2691_5[2]),.dout(n2985),.clk(gclk));
	jand g2904(.dina(n2985),.dinb(n2984),.dout(n2986),.clk(gclk));
	jand g2905(.dina(n2986),.dinb(n2983),.dout(n2987),.clk(gclk));
	jand g2906(.dina(n2987),.dinb(n2982),.dout(n2988),.clk(gclk));
	jxor g2907(.dina(n2988),.dinb(w_n808_8[1]),.dout(n2989),.clk(gclk));
	jor g2908(.dina(w_n2892_0[0]),.dinb(w_n2818_0[0]),.dout(n2990),.clk(gclk));
	jand g2909(.dina(w_n2990_0[1]),.dinb(w_n954_19[1]),.dout(n2991),.clk(gclk));
	jand g2910(.dina(w_n2883_3[0]),.dinb(w_n2844_0[2]),.dout(n2992),.clk(gclk));
	jand g2911(.dina(w_n2889_4[0]),.dinb(w_n2693_2[2]),.dout(n2993),.clk(gclk));
	jand g2912(.dina(w_n2885_0[0]),.dinb(w_n2816_0[0]),.dout(n2994),.clk(gclk));
	jand g2913(.dina(n2994),.dinb(w_n2752_0[0]),.dout(n2995),.clk(gclk));
	jand g2914(.dina(w_n2995_4[2]),.dinb(w_n2698_3[0]),.dout(n2996),.clk(gclk));
	jand g2915(.dina(w_n2887_4[1]),.dinb(w_n2700_3[0]),.dout(n2997),.clk(gclk));
	jor g2916(.dina(n2997),.dinb(n2996),.dout(n2998),.clk(gclk));
	jor g2917(.dina(n2998),.dinb(n2993),.dout(n2999),.clk(gclk));
	jor g2918(.dina(n2999),.dinb(n2992),.dout(n3000),.clk(gclk));
	jxor g2919(.dina(w_n3000_0[1]),.dinb(n2991),.dout(n3001),.clk(gclk));
	jxor g2920(.dina(w_n3001_0[1]),.dinb(w_n2989_0[1]),.dout(n3002),.clk(gclk));
	jxor g2921(.dina(w_n3002_0[1]),.dinb(w_n2981_0[1]),.dout(n3003),.clk(gclk));
	jxor g2922(.dina(w_n2719_0[0]),.dinb(w_n2718_0[0]),.dout(n3004),.clk(gclk));
	jand g2923(.dina(w_n3004_1[2]),.dinb(w_n2794_1[2]),.dout(n3005),.clk(gclk));
	jand g2924(.dina(w_n2799_1[1]),.dinb(w_n2677_4[1]),.dout(n3006),.clk(gclk));
	jand g2925(.dina(w_n2808_1[2]),.dinb(w_n2684_3[2]),.dout(n3007),.clk(gclk));
	jand g2926(.dina(w_n2804_1[2]),.dinb(w_n2679_3[0]),.dout(n3008),.clk(gclk));
	jor g2927(.dina(n3008),.dinb(n3007),.dout(n3009),.clk(gclk));
	jor g2928(.dina(n3009),.dinb(n3006),.dout(n3010),.clk(gclk));
	jor g2929(.dina(n3010),.dinb(n3005),.dout(n3011),.clk(gclk));
	jxor g2930(.dina(n3011),.dinb(w_n699_7[2]),.dout(n3012),.clk(gclk));
	jxor g2931(.dina(w_n3012_0[1]),.dinb(w_n3003_0[1]),.dout(n3013),.clk(gclk));
	jxor g2932(.dina(w_n3013_0[1]),.dinb(w_n2978_0[1]),.dout(n3014),.clk(gclk));
	jand g2933(.dina(w_n3014_0[1]),.dinb(w_n2789_0[1]),.dout(n3015),.clk(gclk));
	jxor g2934(.dina(w_n2725_0[0]),.dinb(w_n2724_0[0]),.dout(n3016),.clk(gclk));
	jand g2935(.dina(w_n3016_1[2]),.dinb(w_n78_2[1]),.dout(n3017),.clk(gclk));
	jand g2936(.dina(w_n2774_2[0]),.dinb(w_n2670_5[0]),.dout(n3018),.clk(gclk));
	jand g2937(.dina(w_n2783_2[0]),.dinb(w_n2677_4[0]),.dout(n3019),.clk(gclk));
	jand g2938(.dina(w_n2779_2[1]),.dinb(w_n2672_2[1]),.dout(n3020),.clk(gclk));
	jor g2939(.dina(n3020),.dinb(n3019),.dout(n3021),.clk(gclk));
	jor g2940(.dina(n3021),.dinb(n3018),.dout(n3022),.clk(gclk));
	jor g2941(.dina(n3022),.dinb(n3017),.dout(n3023),.clk(gclk));
	jxor g2942(.dina(n3023),.dinb(w_n55_5[2]),.dout(n3024),.clk(gclk));
	jxor g2943(.dina(w_n2976_0[0]),.dinb(w_n2975_0[0]),.dout(n3025),.clk(gclk));
	jand g2944(.dina(w_n3025_0[1]),.dinb(w_n3024_0[1]),.dout(n3026),.clk(gclk));
	jnot g2945(.din(w_n2721_0[0]),.dout(n3027),.clk(gclk));
	jxor g2946(.dina(w_n2722_0[0]),.dinb(n3027),.dout(n3028),.clk(gclk));
	jor g2947(.dina(w_n3028_1[2]),.dinb(w_n79_6[0]),.dout(n3029),.clk(gclk));
	jor g2948(.dina(w_n2775_5[1]),.dinb(w_n2671_4[2]),.dout(n3030),.clk(gclk));
	jor g2949(.dina(w_n2780_5[1]),.dinb(w_n2674_3[0]),.dout(n3031),.clk(gclk));
	jor g2950(.dina(w_n2784_6[0]),.dinb(w_n2678_4[1]),.dout(n3032),.clk(gclk));
	jand g2951(.dina(n3032),.dinb(n3031),.dout(n3033),.clk(gclk));
	jand g2952(.dina(n3033),.dinb(n3030),.dout(n3034),.clk(gclk));
	jand g2953(.dina(n3034),.dinb(n3029),.dout(n3035),.clk(gclk));
	jxor g2954(.dina(n3035),.dinb(w_n56_8[0]),.dout(n3036),.clk(gclk));
	jxor g2955(.dina(w_n2973_0[0]),.dinb(w_n2972_0[0]),.dout(n3037),.clk(gclk));
	jand g2956(.dina(w_n3037_0[1]),.dinb(w_n3036_0[1]),.dout(n3038),.clk(gclk));
	jand g2957(.dina(w_n3004_1[1]),.dinb(w_n78_2[0]),.dout(n3039),.clk(gclk));
	jand g2958(.dina(w_n2774_1[2]),.dinb(w_n2677_3[2]),.dout(n3040),.clk(gclk));
	jand g2959(.dina(w_n2783_1[2]),.dinb(w_n2684_3[1]),.dout(n3041),.clk(gclk));
	jand g2960(.dina(w_n2779_2[0]),.dinb(w_n2679_2[2]),.dout(n3042),.clk(gclk));
	jor g2961(.dina(n3042),.dinb(n3041),.dout(n3043),.clk(gclk));
	jor g2962(.dina(n3043),.dinb(n3040),.dout(n3044),.clk(gclk));
	jor g2963(.dina(n3044),.dinb(n3039),.dout(n3045),.clk(gclk));
	jxor g2964(.dina(n3045),.dinb(w_n55_5[1]),.dout(n3046),.clk(gclk));
	jxor g2965(.dina(w_n2970_0[0]),.dinb(w_n2969_0[0]),.dout(n3047),.clk(gclk));
	jand g2966(.dina(w_n3047_0[1]),.dinb(w_n3046_0[1]),.dout(n3048),.clk(gclk));
	jor g2967(.dina(w_n2797_1[1]),.dinb(w_n79_5[2]),.dout(n3049),.clk(gclk));
	jor g2968(.dina(w_n2775_5[0]),.dinb(w_n2678_4[0]),.dout(n3050),.clk(gclk));
	jor g2969(.dina(w_n2780_5[0]),.dinb(w_n2681_3[1]),.dout(n3051),.clk(gclk));
	jor g2970(.dina(w_n2784_5[2]),.dinb(w_n2687_5[0]),.dout(n3052),.clk(gclk));
	jand g2971(.dina(n3052),.dinb(n3051),.dout(n3053),.clk(gclk));
	jand g2972(.dina(n3053),.dinb(n3050),.dout(n3054),.clk(gclk));
	jand g2973(.dina(n3054),.dinb(n3049),.dout(n3055),.clk(gclk));
	jxor g2974(.dina(n3055),.dinb(w_n56_7[2]),.dout(n3056),.clk(gclk));
	jxor g2975(.dina(w_n2967_0[0]),.dinb(w_n2966_0[0]),.dout(n3057),.clk(gclk));
	jand g2976(.dina(w_n3057_0[1]),.dinb(w_n3056_0[1]),.dout(n3058),.clk(gclk));
	jor g2977(.dina(w_n2899_1[1]),.dinb(w_n79_5[1]),.dout(n3059),.clk(gclk));
	jor g2978(.dina(w_n2775_4[2]),.dinb(w_n2681_3[0]),.dout(n3060),.clk(gclk));
	jor g2979(.dina(w_n2780_4[2]),.dinb(w_n2687_4[2]),.dout(n3061),.clk(gclk));
	jor g2980(.dina(w_n2784_5[1]),.dinb(w_n2688_5[1]),.dout(n3062),.clk(gclk));
	jand g2981(.dina(n3062),.dinb(n3061),.dout(n3063),.clk(gclk));
	jand g2982(.dina(n3063),.dinb(n3060),.dout(n3064),.clk(gclk));
	jand g2983(.dina(n3064),.dinb(n3059),.dout(n3065),.clk(gclk));
	jxor g2984(.dina(n3065),.dinb(w_n56_7[1]),.dout(n3066),.clk(gclk));
	jxor g2985(.dina(w_n2964_0[0]),.dinb(w_n2963_0[0]),.dout(n3067),.clk(gclk));
	jand g2986(.dina(w_n3067_0[1]),.dinb(w_n3066_0[1]),.dout(n3068),.clk(gclk));
	jor g2987(.dina(w_n2911_1[0]),.dinb(w_n79_5[0]),.dout(n3069),.clk(gclk));
	jor g2988(.dina(w_n2775_4[1]),.dinb(w_n2687_4[1]),.dout(n3070),.clk(gclk));
	jor g2989(.dina(w_n2780_4[1]),.dinb(w_n2688_5[0]),.dout(n3071),.clk(gclk));
	jor g2990(.dina(w_n2784_5[0]),.dinb(w_n2691_5[1]),.dout(n3072),.clk(gclk));
	jand g2991(.dina(n3072),.dinb(n3071),.dout(n3073),.clk(gclk));
	jand g2992(.dina(n3073),.dinb(n3070),.dout(n3074),.clk(gclk));
	jand g2993(.dina(n3074),.dinb(n3069),.dout(n3075),.clk(gclk));
	jxor g2994(.dina(n3075),.dinb(w_n56_7[0]),.dout(n3076),.clk(gclk));
	jor g2995(.dina(w_n2944_0[0]),.dinb(w_n1143_5[0]),.dout(n3077),.clk(gclk));
	jxor g2996(.dina(n3077),.dinb(w_n2952_0[0]),.dout(n3078),.clk(gclk));
	jand g2997(.dina(w_n3078_0[1]),.dinb(w_n3076_0[1]),.dout(n3079),.clk(gclk));
	jor g2998(.dina(w_n2874_1[0]),.dinb(w_n79_4[2]),.dout(n3080),.clk(gclk));
	jor g2999(.dina(w_n2775_4[0]),.dinb(w_n2688_4[2]),.dout(n3081),.clk(gclk));
	jor g3000(.dina(w_n2780_4[0]),.dinb(w_n2691_5[0]),.dout(n3082),.clk(gclk));
	jor g3001(.dina(w_n2784_4[2]),.dinb(w_n2694_3[0]),.dout(n3083),.clk(gclk));
	jand g3002(.dina(n3083),.dinb(n3082),.dout(n3084),.clk(gclk));
	jand g3003(.dina(n3084),.dinb(n3081),.dout(n3085),.clk(gclk));
	jand g3004(.dina(n3085),.dinb(n3080),.dout(n3086),.clk(gclk));
	jxor g3005(.dina(n3086),.dinb(w_n56_6[2]),.dout(n3087),.clk(gclk));
	jand g3006(.dina(w_n2941_1[0]),.dinb(w_n699_7[1]),.dout(n3088),.clk(gclk));
	jxor g3007(.dina(n3088),.dinb(w_n2939_0[0]),.dout(n3089),.clk(gclk));
	jand g3008(.dina(w_n3089_0[1]),.dinb(w_n3087_0[1]),.dout(n3090),.clk(gclk));
	jand g3009(.dina(w_n2823_0[1]),.dinb(w_n78_1[2]),.dout(n3091),.clk(gclk));
	jand g3010(.dina(w_n2779_1[2]),.dinb(w_n2698_2[2]),.dout(n3092),.clk(gclk));
	jand g3011(.dina(w_n2774_1[1]),.dinb(w_n2700_2[2]),.dout(n3093),.clk(gclk));
	jor g3012(.dina(n3093),.dinb(n3092),.dout(n3094),.clk(gclk));
	jor g3013(.dina(n3094),.dinb(n3091),.dout(n3095),.clk(gclk));
	jnot g3014(.din(w_n3095_0[1]),.dout(n3096),.clk(gclk));
	jand g3015(.dina(w_n2698_2[1]),.dinb(w_n70_0[0]),.dout(n3097),.clk(gclk));
	jnot g3016(.din(w_n3097_0[2]),.dout(n3098),.clk(gclk));
	jand g3017(.dina(n3098),.dinb(w_n55_5[0]),.dout(n3099),.clk(gclk));
	jand g3018(.dina(n3099),.dinb(n3096),.dout(n3100),.clk(gclk));
	jand g3019(.dina(w_n2844_0[1]),.dinb(w_n78_1[1]),.dout(n3101),.clk(gclk));
	jand g3020(.dina(w_n2774_1[0]),.dinb(w_n2693_2[1]),.dout(n3102),.clk(gclk));
	jand g3021(.dina(w_n2783_1[1]),.dinb(w_n2698_2[0]),.dout(n3103),.clk(gclk));
	jand g3022(.dina(w_n2779_1[1]),.dinb(w_n2700_2[1]),.dout(n3104),.clk(gclk));
	jor g3023(.dina(n3104),.dinb(n3103),.dout(n3105),.clk(gclk));
	jor g3024(.dina(n3105),.dinb(n3102),.dout(n3106),.clk(gclk));
	jor g3025(.dina(n3106),.dinb(n3101),.dout(n3107),.clk(gclk));
	jnot g3026(.din(w_n3107_0[1]),.dout(n3108),.clk(gclk));
	jand g3027(.dina(n3108),.dinb(w_n3100_0[1]),.dout(n3109),.clk(gclk));
	jand g3028(.dina(w_n3109_0[1]),.dinb(w_n2941_0[2]),.dout(n3110),.clk(gclk));
	jor g3029(.dina(w_n2858_1[0]),.dinb(w_n79_4[1]),.dout(n3111),.clk(gclk));
	jor g3030(.dina(w_n2775_3[2]),.dinb(w_n2691_4[2]),.dout(n3112),.clk(gclk));
	jor g3031(.dina(w_n2784_4[1]),.dinb(w_n2862_2[0]),.dout(n3113),.clk(gclk));
	jor g3032(.dina(w_n2780_3[2]),.dinb(w_n2694_2[2]),.dout(n3114),.clk(gclk));
	jand g3033(.dina(n3114),.dinb(n3113),.dout(n3115),.clk(gclk));
	jand g3034(.dina(n3115),.dinb(n3112),.dout(n3116),.clk(gclk));
	jand g3035(.dina(n3116),.dinb(n3111),.dout(n3117),.clk(gclk));
	jxor g3036(.dina(n3117),.dinb(w_n56_6[1]),.dout(n3118),.clk(gclk));
	jxor g3037(.dina(w_n3109_0[0]),.dinb(w_n2941_0[1]),.dout(n3119),.clk(gclk));
	jand g3038(.dina(w_n3119_0[1]),.dinb(w_n3118_0[1]),.dout(n3120),.clk(gclk));
	jor g3039(.dina(n3120),.dinb(n3110),.dout(n3121),.clk(gclk));
	jxor g3040(.dina(w_n3089_0[0]),.dinb(w_n3087_0[0]),.dout(n3122),.clk(gclk));
	jand g3041(.dina(w_n3122_0[1]),.dinb(w_n3121_0[1]),.dout(n3123),.clk(gclk));
	jor g3042(.dina(n3123),.dinb(n3090),.dout(n3124),.clk(gclk));
	jxor g3043(.dina(w_n3078_0[0]),.dinb(w_n3076_0[0]),.dout(n3125),.clk(gclk));
	jand g3044(.dina(w_n3125_0[1]),.dinb(w_n3124_0[1]),.dout(n3126),.clk(gclk));
	jor g3045(.dina(n3126),.dinb(n3079),.dout(n3127),.clk(gclk));
	jxor g3046(.dina(w_n3067_0[0]),.dinb(w_n3066_0[0]),.dout(n3128),.clk(gclk));
	jand g3047(.dina(w_n3128_0[1]),.dinb(w_n3127_0[1]),.dout(n3129),.clk(gclk));
	jor g3048(.dina(n3129),.dinb(n3068),.dout(n3130),.clk(gclk));
	jxor g3049(.dina(w_n3057_0[0]),.dinb(w_n3056_0[0]),.dout(n3131),.clk(gclk));
	jand g3050(.dina(w_n3131_0[1]),.dinb(w_n3130_0[1]),.dout(n3132),.clk(gclk));
	jor g3051(.dina(n3132),.dinb(n3058),.dout(n3133),.clk(gclk));
	jxor g3052(.dina(w_n3047_0[0]),.dinb(w_n3046_0[0]),.dout(n3134),.clk(gclk));
	jand g3053(.dina(w_n3134_0[1]),.dinb(w_n3133_0[1]),.dout(n3135),.clk(gclk));
	jor g3054(.dina(n3135),.dinb(n3048),.dout(n3136),.clk(gclk));
	jxor g3055(.dina(w_n3037_0[0]),.dinb(w_n3036_0[0]),.dout(n3137),.clk(gclk));
	jand g3056(.dina(w_n3137_0[1]),.dinb(w_n3136_0[1]),.dout(n3138),.clk(gclk));
	jor g3057(.dina(n3138),.dinb(n3038),.dout(n3139),.clk(gclk));
	jxor g3058(.dina(w_n3025_0[0]),.dinb(w_n3024_0[0]),.dout(n3140),.clk(gclk));
	jand g3059(.dina(w_n3140_0[1]),.dinb(w_n3139_0[1]),.dout(n3141),.clk(gclk));
	jor g3060(.dina(n3141),.dinb(n3026),.dout(n3142),.clk(gclk));
	jxor g3061(.dina(w_n3014_0[0]),.dinb(w_n2789_0[0]),.dout(n3143),.clk(gclk));
	jand g3062(.dina(w_n3143_0[1]),.dinb(w_n3142_0[1]),.dout(n3144),.clk(gclk));
	jor g3063(.dina(n3144),.dinb(n3015),.dout(n3145),.clk(gclk));
	jand g3064(.dina(w_n2769_3[2]),.dinb(w_n2670_4[2]),.dout(n3146),.clk(gclk));
	jand g3065(.dina(w_n2770_0[1]),.dinb(w_n2727_0[0]),.dout(n3147),.clk(gclk));
	jor g3066(.dina(n3147),.dinb(n3146),.dout(n3148),.clk(gclk));
	jor g3067(.dina(w_n2767_0[1]),.dinb(w_n2750_0[1]),.dout(n3149),.clk(gclk));
	jnot g3068(.din(n3149),.dout(n3150),.clk(gclk));
	jand g3069(.dina(w_n2767_0[0]),.dinb(w_n2750_0[0]),.dout(n3151),.clk(gclk));
	jnot g3070(.din(n3151),.dout(n3152),.clk(gclk));
	jand g3071(.dina(n3152),.dinb(w_n2733_0[0]),.dout(n3153),.clk(gclk));
	jor g3072(.dina(n3153),.dinb(n3150),.dout(n3154),.clk(gclk));
	jnot g3073(.din(w_n1653_0[0]),.dout(n3155),.clk(gclk));
	jand g3074(.dina(w_n461_1[0]),.dinb(w_n312_1[2]),.dout(n3156),.clk(gclk));
	jand g3075(.dina(n3156),.dinb(w_n304_1[1]),.dout(n3157),.clk(gclk));
	jand g3076(.dina(n3157),.dinb(w_n898_0[0]),.dout(n3158),.clk(gclk));
	jand g3077(.dina(n3158),.dinb(w_n914_0[0]),.dout(n3159),.clk(gclk));
	jand g3078(.dina(w_n711_0[0]),.dinb(w_n564_0[0]),.dout(n3160),.clk(gclk));
	jand g3079(.dina(n3160),.dinb(w_n821_0[1]),.dout(n3161),.clk(gclk));
	jand g3080(.dina(w_n612_1[1]),.dinb(w_n499_0[1]),.dout(n3162),.clk(gclk));
	jand g3081(.dina(w_n853_0[2]),.dinb(w_n225_1[0]),.dout(n3163),.clk(gclk));
	jand g3082(.dina(n3163),.dinb(n3162),.dout(n3164),.clk(gclk));
	jand g3083(.dina(n3164),.dinb(w_n1189_0[1]),.dout(n3165),.clk(gclk));
	jand g3084(.dina(n3165),.dinb(n3161),.dout(n3166),.clk(gclk));
	jand g3085(.dina(n3166),.dinb(w_n3159_0[1]),.dout(n3167),.clk(gclk));
	jand g3086(.dina(w_n2427_0[0]),.dinb(w_n1011_0[0]),.dout(n3168),.clk(gclk));
	jand g3087(.dina(n3168),.dinb(n3167),.dout(n3169),.clk(gclk));
	jand g3088(.dina(n3169),.dinb(w_n3155_0[1]),.dout(n3170),.clk(gclk));
	jnot g3089(.din(n3170),.dout(n3171),.clk(gclk));
	jxor g3090(.dina(w_n3171_0[1]),.dinb(w_n3154_0[1]),.dout(n3172),.clk(gclk));
	jxor g3091(.dina(w_n3172_6[1]),.dinb(w_n2773_4[1]),.dout(n3173),.clk(gclk));
	jxor g3092(.dina(w_n3173_0[1]),.dinb(w_n3148_0[1]),.dout(n3174),.clk(gclk));
	jand g3093(.dina(w_n3174_1[2]),.dinb(w_n78_1[0]),.dout(n3175),.clk(gclk));
	jnot g3094(.din(w_n3172_6[0]),.dout(n3176),.clk(gclk));
	jand g3095(.dina(w_n3176_2[2]),.dinb(w_n2774_0[2]),.dout(n3177),.clk(gclk));
	jand g3096(.dina(w_n2783_1[0]),.dinb(w_n2670_4[1]),.dout(n3178),.clk(gclk));
	jand g3097(.dina(w_n2779_1[0]),.dinb(w_n2769_3[1]),.dout(n3179),.clk(gclk));
	jor g3098(.dina(n3179),.dinb(n3178),.dout(n3180),.clk(gclk));
	jor g3099(.dina(n3180),.dinb(n3177),.dout(n3181),.clk(gclk));
	jor g3100(.dina(n3181),.dinb(n3175),.dout(n3182),.clk(gclk));
	jxor g3101(.dina(n3182),.dinb(w_n55_4[2]),.dout(n3183),.clk(gclk));
	jand g3102(.dina(w_n3012_0[0]),.dinb(w_n3003_0[0]),.dout(n3184),.clk(gclk));
	jand g3103(.dina(w_n3013_0[0]),.dinb(w_n2978_0[0]),.dout(n3185),.clk(gclk));
	jor g3104(.dina(n3185),.dinb(n3184),.dout(n3186),.clk(gclk));
	jand g3105(.dina(w_n3001_0[0]),.dinb(w_n2989_0[0]),.dout(n3187),.clk(gclk));
	jand g3106(.dina(w_n3002_0[0]),.dinb(w_n2981_0[0]),.dout(n3188),.clk(gclk));
	jor g3107(.dina(n3188),.dinb(n3187),.dout(n3189),.clk(gclk));
	jor g3108(.dina(w_n2899_1[0]),.dinb(w_n2857_5[1]),.dout(n3190),.clk(gclk));
	jor g3109(.dina(w_n2860_4[2]),.dinb(w_n2681_2[2]),.dout(n3191),.clk(gclk));
	jor g3110(.dina(w_n2865_4[2]),.dinb(w_n2687_4[0]),.dout(n3192),.clk(gclk));
	jor g3111(.dina(w_n2863_5[1]),.dinb(w_n2688_4[1]),.dout(n3193),.clk(gclk));
	jand g3112(.dina(n3193),.dinb(n3192),.dout(n3194),.clk(gclk));
	jand g3113(.dina(n3194),.dinb(n3191),.dout(n3195),.clk(gclk));
	jand g3114(.dina(n3195),.dinb(n3190),.dout(n3196),.clk(gclk));
	jxor g3115(.dina(n3196),.dinb(w_n808_8[0]),.dout(n3197),.clk(gclk));
	jnot g3116(.din(w_n2883_2[2]),.dout(n3198),.clk(gclk));
	jor g3117(.dina(w_n3198_5[2]),.dinb(w_n2858_0[2]),.dout(n3199),.clk(gclk));
	jnot g3118(.din(w_n2889_3[2]),.dout(n3200),.clk(gclk));
	jor g3119(.dina(w_n3200_3[2]),.dinb(w_n2691_4[1]),.dout(n3201),.clk(gclk));
	jnot g3120(.din(w_n2995_4[1]),.dout(n3202),.clk(gclk));
	jor g3121(.dina(w_n3202_3[2]),.dinb(w_n2862_1[2]),.dout(n3203),.clk(gclk));
	jnot g3122(.din(w_n2887_4[0]),.dout(n3204),.clk(gclk));
	jor g3123(.dina(w_n3204_3[2]),.dinb(w_n2694_2[1]),.dout(n3205),.clk(gclk));
	jand g3124(.dina(n3205),.dinb(n3203),.dout(n3206),.clk(gclk));
	jand g3125(.dina(n3206),.dinb(n3201),.dout(n3207),.clk(gclk));
	jand g3126(.dina(n3207),.dinb(n3199),.dout(n3208),.clk(gclk));
	jxor g3127(.dina(n3208),.dinb(w_n954_19[0]),.dout(n3209),.clk(gclk));
	jnot g3128(.din(n3209),.dout(n3210),.clk(gclk));
	jor g3129(.dina(w_n3000_0[0]),.dinb(w_n2990_0[0]),.dout(n3211),.clk(gclk));
	jnot g3130(.din(n3211),.dout(n3212),.clk(gclk));
	jand g3131(.dina(w_n3212_0[1]),.dinb(w_n954_18[2]),.dout(n3213),.clk(gclk));
	jor g3132(.dina(n3213),.dinb(w_n2893_0[1]),.dout(n3214),.clk(gclk));
	jand g3133(.dina(w_n3212_0[0]),.dinb(w_n2893_0[0]),.dout(n3215),.clk(gclk));
	jnot g3134(.din(w_n3215_0[1]),.dout(n3216),.clk(gclk));
	jand g3135(.dina(n3216),.dinb(n3214),.dout(n3217),.clk(gclk));
	jxor g3136(.dina(w_n3217_0[1]),.dinb(w_n3210_0[1]),.dout(n3218),.clk(gclk));
	jxor g3137(.dina(w_n3218_0[1]),.dinb(w_n3197_0[1]),.dout(n3219),.clk(gclk));
	jxor g3138(.dina(w_n3219_0[1]),.dinb(w_n3189_0[1]),.dout(n3220),.clk(gclk));
	jor g3139(.dina(w_n3028_1[1]),.dinb(w_n2795_4[2]),.dout(n3221),.clk(gclk));
	jor g3140(.dina(w_n2800_4[0]),.dinb(w_n2671_4[1]),.dout(n3222),.clk(gclk));
	jor g3141(.dina(w_n2805_4[0]),.dinb(w_n2674_2[2]),.dout(n3223),.clk(gclk));
	jor g3142(.dina(w_n2809_4[2]),.dinb(w_n2678_3[2]),.dout(n3224),.clk(gclk));
	jand g3143(.dina(n3224),.dinb(n3223),.dout(n3225),.clk(gclk));
	jand g3144(.dina(n3225),.dinb(n3222),.dout(n3226),.clk(gclk));
	jand g3145(.dina(n3226),.dinb(n3221),.dout(n3227),.clk(gclk));
	jxor g3146(.dina(n3227),.dinb(w_n1143_4[2]),.dout(n3228),.clk(gclk));
	jxor g3147(.dina(w_n3228_0[1]),.dinb(w_n3220_0[1]),.dout(n3229),.clk(gclk));
	jxor g3148(.dina(w_n3229_0[1]),.dinb(w_n3186_0[1]),.dout(n3230),.clk(gclk));
	jxor g3149(.dina(w_n3230_0[1]),.dinb(w_n3183_0[1]),.dout(n3231),.clk(gclk));
	jxor g3150(.dina(w_n3231_0[1]),.dinb(w_n3145_0[1]),.dout(n3232),.clk(gclk));
	jnot g3151(.din(w_n68_6[1]),.dout(n3233),.clk(gclk));
	jand g3152(.dina(w_n49_2[0]),.dinb(w_a0_0[2]),.dout(n3234),.clk(gclk));
	jxor g3153(.dina(n3234),.dinb(w_n62_0[0]),.dout(n3235),.clk(gclk));
	jxor g3154(.dina(w_n3235_0[1]),.dinb(w_n3233_9[2]),.dout(n3236),.clk(gclk));
	jand g3155(.dina(w_n3236_0[1]),.dinb(w_a0_0[1]),.dout(n3237),.clk(gclk));
	jnot g3156(.din(w_n3237_2[1]),.dout(n3238),.clk(gclk));
	jor g3157(.dina(w_n3171_0[0]),.dinb(w_n3154_0[0]),.dout(n3239),.clk(gclk));
	jnot g3158(.din(n3239),.dout(n3240),.clk(gclk));
	jand g3159(.dina(w_n2380_1[2]),.dinb(w_n437_0[2]),.dout(n3241),.clk(gclk));
	jand g3160(.dina(n3241),.dinb(w_n936_0[0]),.dout(n3242),.clk(gclk));
	jand g3161(.dina(w_n772_1[1]),.dinb(w_n477_1[0]),.dout(n3243),.clk(gclk));
	jand g3162(.dina(w_n624_1[0]),.dinb(w_n261_0[2]),.dout(n3244),.clk(gclk));
	jand g3163(.dina(n3244),.dinb(n3243),.dout(n3245),.clk(gclk));
	jand g3164(.dina(n3245),.dinb(w_n3242_0[2]),.dout(n3246),.clk(gclk));
	jand g3165(.dina(n3246),.dinb(w_n2321_0[0]),.dout(n3247),.clk(gclk));
	jand g3166(.dina(w_n882_1[0]),.dinb(w_n323_2[0]),.dout(n3248),.clk(gclk));
	jand g3167(.dina(n3248),.dinb(w_n381_0[2]),.dout(n3249),.clk(gclk));
	jand g3168(.dina(n3249),.dinb(w_n2580_0[0]),.dout(n3250),.clk(gclk));
	jand g3169(.dina(w_n724_1[0]),.dinb(w_n918_1[1]),.dout(n3251),.clk(gclk));
	jand g3170(.dina(w_n594_1[1]),.dinb(w_n370_1[0]),.dout(n3252),.clk(gclk));
	jand g3171(.dina(n3252),.dinb(n3251),.dout(n3253),.clk(gclk));
	jand g3172(.dina(n3253),.dinb(w_n2655_0[0]),.dout(n3254),.clk(gclk));
	jand g3173(.dina(n3254),.dinb(w_n3250_0[1]),.dout(n3255),.clk(gclk));
	jand g3174(.dina(n3255),.dinb(n3247),.dout(n3256),.clk(gclk));
	jand g3175(.dina(w_n363_0[2]),.dinb(w_n291_1[0]),.dout(n3257),.clk(gclk));
	jand g3176(.dina(w_n3257_0[1]),.dinb(w_n277_2[2]),.dout(n3258),.clk(gclk));
	jand g3177(.dina(w_n710_1[2]),.dinb(w_n232_1[0]),.dout(n3259),.clk(gclk));
	jand g3178(.dina(n3259),.dinb(w_n2538_0[0]),.dout(n3260),.clk(gclk));
	jand g3179(.dina(n3260),.dinb(w_n3258_1[2]),.dout(n3261),.clk(gclk));
	jand g3180(.dina(n3261),.dinb(w_n2453_0[0]),.dout(n3262),.clk(gclk));
	jand g3181(.dina(w_n868_0[2]),.dinb(w_n153_0[2]),.dout(n3263),.clk(gclk));
	jand g3182(.dina(w_n506_0[2]),.dinb(w_n312_1[1]),.dout(n3264),.clk(gclk));
	jand g3183(.dina(n3264),.dinb(w_n3263_0[1]),.dout(n3265),.clk(gclk));
	jand g3184(.dina(n3265),.dinb(w_n822_1[1]),.dout(n3266),.clk(gclk));
	jand g3185(.dina(n3266),.dinb(w_n361_0[0]),.dout(n3267),.clk(gclk));
	jand g3186(.dina(n3267),.dinb(n3262),.dout(n3268),.clk(gclk));
	jand g3187(.dina(n3268),.dinb(w_n3256_0[2]),.dout(n3269),.clk(gclk));
	jand g3188(.dina(n3269),.dinb(w_n434_0[0]),.dout(n3270),.clk(gclk));
	jand g3189(.dina(w_n3270_0[2]),.dinb(w_n3240_0[1]),.dout(n3271),.clk(gclk));
	jand g3190(.dina(w_n426_1[1]),.dinb(w_n374_1[0]),.dout(n3272),.clk(gclk));
	jand g3191(.dina(n3272),.dinb(w_n2289_0[0]),.dout(n3273),.clk(gclk));
	jnot g3192(.din(w_n650_0[0]),.dout(n3274),.clk(gclk));
	jand g3193(.dina(w_n1310_0[0]),.dinb(w_n3274_0[1]),.dout(n3275),.clk(gclk));
	jand g3194(.dina(w_n2511_1[0]),.dinb(w_n930_1[0]),.dout(n3276),.clk(gclk));
	jand g3195(.dina(n3276),.dinb(n3275),.dout(n3277),.clk(gclk));
	jand g3196(.dina(n3277),.dinb(n3273),.dout(n3278),.clk(gclk));
	jand g3197(.dina(w_n2417_0[0]),.dinb(w_n2307_0[0]),.dout(n3279),.clk(gclk));
	jand g3198(.dina(n3279),.dinb(n3278),.dout(n3280),.clk(gclk));
	jand g3199(.dina(n3280),.dinb(w_n719_1[0]),.dout(n3281),.clk(gclk));
	jand g3200(.dina(n3281),.dinb(w_n275_0[0]),.dout(n3282),.clk(gclk));
	jxor g3201(.dina(w_n3282_0[2]),.dinb(w_n3271_0[1]),.dout(n3283),.clk(gclk));
	jxor g3202(.dina(w_n3270_0[1]),.dinb(w_n3240_0[0]),.dout(n3284),.clk(gclk));
	jor g3203(.dina(w_n3284_8[2]),.dinb(w_n3283_8[1]),.dout(n3285),.clk(gclk));
	jnot g3204(.din(w_n3285_0[1]),.dout(n3286),.clk(gclk));
	jor g3205(.dina(w_n3284_8[1]),.dinb(w_n3172_5[2]),.dout(n3287),.clk(gclk));
	jnot g3206(.din(w_n3287_0[1]),.dout(n3288),.clk(gclk));
	jand g3207(.dina(w_n3176_2[1]),.dinb(w_n2769_3[0]),.dout(n3289),.clk(gclk));
	jand g3208(.dina(w_n3173_0[0]),.dinb(w_n3148_0[0]),.dout(n3290),.clk(gclk));
	jor g3209(.dina(n3290),.dinb(n3289),.dout(n3291),.clk(gclk));
	jand g3210(.dina(w_n3270_0[0]),.dinb(w_n3172_5[1]),.dout(n3292),.clk(gclk));
	jnot g3211(.din(n3292),.dout(n3293),.clk(gclk));
	jand g3212(.dina(n3293),.dinb(w_n3287_0[0]),.dout(n3294),.clk(gclk));
	jand g3213(.dina(w_n3294_0[1]),.dinb(w_n3291_0[1]),.dout(n3295),.clk(gclk));
	jor g3214(.dina(n3295),.dinb(n3288),.dout(n3296),.clk(gclk));
	jand g3215(.dina(w_n3284_8[0]),.dinb(w_n3282_0[1]),.dout(n3297),.clk(gclk));
	jnot g3216(.din(n3297),.dout(n3298),.clk(gclk));
	jand g3217(.dina(n3298),.dinb(w_n3285_0[0]),.dout(n3299),.clk(gclk));
	jand g3218(.dina(w_n3299_0[2]),.dinb(w_n3296_0[1]),.dout(n3300),.clk(gclk));
	jor g3219(.dina(n3300),.dinb(n3286),.dout(n3301),.clk(gclk));
	jnot g3220(.din(w_n3283_8[0]),.dout(n3302),.clk(gclk));
	jand g3221(.dina(w_n3282_0[0]),.dinb(w_n3271_0[0]),.dout(n3303),.clk(gclk));
	jnot g3222(.din(w_n1322_0[0]),.dout(n3304),.clk(gclk));
	jand g3223(.dina(n3304),.dinb(w_n319_0[0]),.dout(n3305),.clk(gclk));
	jand g3224(.dina(n3305),.dinb(w_n287_0[0]),.dout(n3306),.clk(gclk));
	jand g3225(.dina(w_n254_1[1]),.dinb(w_n241_0[2]),.dout(n3307),.clk(gclk));
	jand g3226(.dina(w_n3307_1[2]),.dinb(w_n1209_1[0]),.dout(n3308),.clk(gclk));
	jand g3227(.dina(n3308),.dinb(w_n731_0[0]),.dout(n3309),.clk(gclk));
	jand g3228(.dina(n3309),.dinb(w_n746_0[1]),.dout(n3310),.clk(gclk));
	jand g3229(.dina(n3310),.dinb(n3306),.dout(n3311),.clk(gclk));
	jand g3230(.dina(w_n786_1[0]),.dinb(w_n719_0[2]),.dout(n3312),.clk(gclk));
	jand g3231(.dina(n3312),.dinb(w_n218_0[0]),.dout(n3313),.clk(gclk));
	jand g3232(.dina(n3313),.dinb(n3311),.dout(n3314),.clk(gclk));
	jxor g3233(.dina(w_n3314_0[2]),.dinb(w_n3303_0[1]),.dout(n3315),.clk(gclk));
	jnot g3234(.din(w_n3315_7[2]),.dout(n3316),.clk(gclk));
	jand g3235(.dina(w_n3316_0[2]),.dinb(w_n3302_0[2]),.dout(n3317),.clk(gclk));
	jand g3236(.dina(w_n3314_0[1]),.dinb(w_n3283_7[2]),.dout(n3318),.clk(gclk));
	jor g3237(.dina(n3318),.dinb(w_n3317_0[1]),.dout(n3319),.clk(gclk));
	jxor g3238(.dina(w_n3319_0[1]),.dinb(w_n3301_0[1]),.dout(n3320),.clk(gclk));
	jor g3239(.dina(w_n3320_1[2]),.dinb(w_n3238_7[1]),.dout(n3321),.clk(gclk));
	jor g3240(.dina(w_n3236_0[0]),.dinb(w_n61_1[0]),.dout(n3322),.clk(gclk));
	jor g3241(.dina(w_n3322_7[1]),.dinb(w_n3315_7[1]),.dout(n3323),.clk(gclk));
	jand g3242(.dina(w_a1_0[0]),.dinb(w_n61_0[2]),.dout(n3324),.clk(gclk));
	jnot g3243(.din(w_n3324_2[1]),.dout(n3325),.clk(gclk));
	jor g3244(.dina(w_n3325_5[1]),.dinb(w_n3283_7[1]),.dout(n3326),.clk(gclk));
	jand g3245(.dina(w_n63_2[1]),.dinb(w_a2_0[1]),.dout(n3327),.clk(gclk));
	jnot g3246(.din(n3327),.dout(n3328),.clk(gclk));
	jor g3247(.dina(w_n3328_5[2]),.dinb(w_n3284_7[2]),.dout(n3329),.clk(gclk));
	jand g3248(.dina(n3329),.dinb(n3326),.dout(n3330),.clk(gclk));
	jand g3249(.dina(n3330),.dinb(n3323),.dout(n3331),.clk(gclk));
	jand g3250(.dina(n3331),.dinb(n3321),.dout(n3332),.clk(gclk));
	jxor g3251(.dina(n3332),.dinb(w_n3233_9[1]),.dout(n3333),.clk(gclk));
	jand g3252(.dina(w_n3333_0[1]),.dinb(w_n3232_0[1]),.dout(n3334),.clk(gclk));
	jxor g3253(.dina(w_n3143_0[0]),.dinb(w_n3142_0[0]),.dout(n3335),.clk(gclk));
	jnot g3254(.din(w_n3299_0[1]),.dout(n3336),.clk(gclk));
	jxor g3255(.dina(n3336),.dinb(w_n3296_0[0]),.dout(n3337),.clk(gclk));
	jor g3256(.dina(w_n3337_1[2]),.dinb(w_n3238_7[0]),.dout(n3338),.clk(gclk));
	jor g3257(.dina(w_n3322_7[0]),.dinb(w_n3283_7[0]),.dout(n3339),.clk(gclk));
	jor g3258(.dina(w_n3325_5[0]),.dinb(w_n3284_7[1]),.dout(n3340),.clk(gclk));
	jor g3259(.dina(w_n3328_5[1]),.dinb(w_n3172_5[0]),.dout(n3341),.clk(gclk));
	jand g3260(.dina(n3341),.dinb(n3340),.dout(n3342),.clk(gclk));
	jand g3261(.dina(n3342),.dinb(n3339),.dout(n3343),.clk(gclk));
	jand g3262(.dina(n3343),.dinb(n3338),.dout(n3344),.clk(gclk));
	jxor g3263(.dina(n3344),.dinb(w_n3233_9[0]),.dout(n3345),.clk(gclk));
	jand g3264(.dina(w_n3345_0[1]),.dinb(w_n3335_0[1]),.dout(n3346),.clk(gclk));
	jxor g3265(.dina(w_n3345_0[0]),.dinb(w_n3335_0[0]),.dout(n3347),.clk(gclk));
	jxor g3266(.dina(w_n3140_0[0]),.dinb(w_n3139_0[0]),.dout(n3348),.clk(gclk));
	jxor g3267(.dina(w_n3137_0[0]),.dinb(w_n3136_0[0]),.dout(n3349),.clk(gclk));
	jxor g3268(.dina(w_n3134_0[0]),.dinb(w_n3133_0[0]),.dout(n3350),.clk(gclk));
	jxor g3269(.dina(w_n3131_0[0]),.dinb(w_n3130_0[0]),.dout(n3351),.clk(gclk));
	jxor g3270(.dina(w_n3128_0[0]),.dinb(w_n3127_0[0]),.dout(n3352),.clk(gclk));
	jxor g3271(.dina(w_n3125_0[0]),.dinb(w_n3124_0[0]),.dout(n3353),.clk(gclk));
	jxor g3272(.dina(w_n3122_0[0]),.dinb(w_n3121_0[0]),.dout(n3354),.clk(gclk));
	jor g3273(.dina(w_n3238_6[2]),.dinb(w_n2899_0[2]),.dout(n3355),.clk(gclk));
	jor g3274(.dina(w_n3322_6[2]),.dinb(w_n2681_2[1]),.dout(n3356),.clk(gclk));
	jor g3275(.dina(w_n3325_4[2]),.dinb(w_n2687_3[2]),.dout(n3357),.clk(gclk));
	jor g3276(.dina(w_n3328_5[0]),.dinb(w_n2688_4[0]),.dout(n3358),.clk(gclk));
	jand g3277(.dina(n3358),.dinb(n3357),.dout(n3359),.clk(gclk));
	jand g3278(.dina(n3359),.dinb(n3356),.dout(n3360),.clk(gclk));
	jand g3279(.dina(n3360),.dinb(n3355),.dout(n3361),.clk(gclk));
	jxor g3280(.dina(n3361),.dinb(w_n3233_8[2]),.dout(n3362),.clk(gclk));
	jnot g3281(.din(w_n3100_0[0]),.dout(n3363),.clk(gclk));
	jand g3282(.dina(n3363),.dinb(w_n55_4[1]),.dout(n3364),.clk(gclk));
	jxor g3283(.dina(n3364),.dinb(w_n3107_0[0]),.dout(n3365),.clk(gclk));
	jand g3284(.dina(w_n3097_0[1]),.dinb(w_n55_4[0]),.dout(n3366),.clk(gclk));
	jxor g3285(.dina(n3366),.dinb(w_n3095_0[0]),.dout(n3367),.clk(gclk));
	jxor g3286(.dina(w_n2702_0[0]),.dinb(w_n2696_0[0]),.dout(n3368),.clk(gclk));
	jand g3287(.dina(w_n3237_2[0]),.dinb(n3368),.dout(n3369),.clk(gclk));
	jor g3288(.dina(w_n3322_6[1]),.dinb(w_n2691_4[0]),.dout(n3370),.clk(gclk));
	jand g3289(.dina(w_n3324_2[0]),.dinb(w_n2693_2[0]),.dout(n3371),.clk(gclk));
	jnot g3290(.din(n3371),.dout(n3372),.clk(gclk));
	jand g3291(.dina(n3372),.dinb(n3370),.dout(n3373),.clk(gclk));
	jnot g3292(.din(w_n3373_0[1]),.dout(n3374),.clk(gclk));
	jor g3293(.dina(n3374),.dinb(n3369),.dout(n3375),.clk(gclk));
	jand g3294(.dina(w_n2700_2[0]),.dinb(w_n63_2[0]),.dout(n3376),.clk(gclk));
	jor g3295(.dina(n3376),.dinb(w_n3233_8[1]),.dout(n3377),.clk(gclk));
	jnot g3296(.din(n3377),.dout(n3378),.clk(gclk));
	jor g3297(.dina(n3378),.dinb(w_n3375_0[1]),.dout(n3379),.clk(gclk));
	jor g3298(.dina(w_n3238_6[1]),.dinb(w_n2858_0[1]),.dout(n3380),.clk(gclk));
	jand g3299(.dina(w_n3373_0[0]),.dinb(n3380),.dout(n3381),.clk(gclk));
	jor g3300(.dina(n3381),.dinb(w_n3233_8[0]),.dout(n3382),.clk(gclk));
	jand g3301(.dina(w_n3238_6[0]),.dinb(w_n2862_1[1]),.dout(n3383),.clk(gclk));
	jand g3302(.dina(w_n3238_5[2]),.dinb(w_n64_0[0]),.dout(n3384),.clk(gclk));
	jnot g3303(.din(n3384),.dout(n3385),.clk(gclk));
	jand g3304(.dina(n3385),.dinb(w_n2822_0[0]),.dout(n3386),.clk(gclk));
	jor g3305(.dina(n3386),.dinb(n3383),.dout(n3387),.clk(gclk));
	jand g3306(.dina(n3387),.dinb(w_n2694_2[0]),.dout(n3388),.clk(gclk));
	jor g3307(.dina(w_n3235_0[0]),.dinb(w_n2862_1[0]),.dout(n3389),.clk(gclk));
	jand g3308(.dina(n3389),.dinb(w_n61_0[1]),.dout(n3390),.clk(gclk));
	jor g3309(.dina(n3390),.dinb(n3388),.dout(n3391),.clk(gclk));
	jand g3310(.dina(w_n2697_0[1]),.dinb(w_n68_6[0]),.dout(n3392),.clk(gclk));
	jand g3311(.dina(n3392),.dinb(n3391),.dout(n3393),.clk(gclk));
	jor g3312(.dina(n3393),.dinb(w_n3097_0[0]),.dout(n3394),.clk(gclk));
	jand g3313(.dina(w_n3394_0[1]),.dinb(n3382),.dout(n3395),.clk(gclk));
	jand g3314(.dina(n3395),.dinb(w_n3379_0[1]),.dout(n3396),.clk(gclk));
	jand g3315(.dina(w_n3396_0[1]),.dinb(w_n3367_0[2]),.dout(n3397),.clk(gclk));
	jor g3316(.dina(w_n3396_0[0]),.dinb(w_n3367_0[1]),.dout(n3398),.clk(gclk));
	jor g3317(.dina(w_n3238_5[1]),.dinb(w_n2874_0[2]),.dout(n3399),.clk(gclk));
	jor g3318(.dina(w_n3322_6[0]),.dinb(w_n2688_3[2]),.dout(n3400),.clk(gclk));
	jor g3319(.dina(w_n3325_4[1]),.dinb(w_n2691_3[2]),.dout(n3401),.clk(gclk));
	jor g3320(.dina(w_n3328_4[2]),.dinb(w_n2694_1[2]),.dout(n3402),.clk(gclk));
	jand g3321(.dina(n3402),.dinb(n3401),.dout(n3403),.clk(gclk));
	jand g3322(.dina(n3403),.dinb(n3400),.dout(n3404),.clk(gclk));
	jand g3323(.dina(n3404),.dinb(n3399),.dout(n3405),.clk(gclk));
	jxor g3324(.dina(n3405),.dinb(w_n3233_7[2]),.dout(n3406),.clk(gclk));
	jand g3325(.dina(w_n3406_0[1]),.dinb(n3398),.dout(n3407),.clk(gclk));
	jor g3326(.dina(n3407),.dinb(w_n3397_0[1]),.dout(n3408),.clk(gclk));
	jor g3327(.dina(w_n3408_0[1]),.dinb(w_n3365_0[2]),.dout(n3409),.clk(gclk));
	jand g3328(.dina(w_n3408_0[0]),.dinb(w_n3365_0[1]),.dout(n3410),.clk(gclk));
	jor g3329(.dina(w_n3238_5[0]),.dinb(w_n2911_0[2]),.dout(n3411),.clk(gclk));
	jor g3330(.dina(w_n3322_5[2]),.dinb(w_n2687_3[1]),.dout(n3412),.clk(gclk));
	jor g3331(.dina(w_n3325_4[0]),.dinb(w_n2688_3[1]),.dout(n3413),.clk(gclk));
	jor g3332(.dina(w_n3328_4[1]),.dinb(w_n2691_3[1]),.dout(n3414),.clk(gclk));
	jand g3333(.dina(n3414),.dinb(n3413),.dout(n3415),.clk(gclk));
	jand g3334(.dina(n3415),.dinb(n3412),.dout(n3416),.clk(gclk));
	jand g3335(.dina(n3416),.dinb(n3411),.dout(n3417),.clk(gclk));
	jxor g3336(.dina(n3417),.dinb(w_n3233_7[1]),.dout(n3418),.clk(gclk));
	jor g3337(.dina(w_n3418_0[1]),.dinb(n3410),.dout(n3419),.clk(gclk));
	jand g3338(.dina(n3419),.dinb(w_n3409_0[1]),.dout(n3420),.clk(gclk));
	jand g3339(.dina(w_n3420_0[1]),.dinb(w_n3362_0[2]),.dout(n3421),.clk(gclk));
	jor g3340(.dina(w_n3420_0[0]),.dinb(w_n3362_0[1]),.dout(n3422),.clk(gclk));
	jxor g3341(.dina(w_n3119_0[0]),.dinb(w_n3118_0[0]),.dout(n3423),.clk(gclk));
	jand g3342(.dina(w_n3423_0[1]),.dinb(n3422),.dout(n3424),.clk(gclk));
	jor g3343(.dina(n3424),.dinb(w_n3421_0[1]),.dout(n3425),.clk(gclk));
	jor g3344(.dina(w_n3425_0[1]),.dinb(w_n3354_0[2]),.dout(n3426),.clk(gclk));
	jand g3345(.dina(w_n3425_0[0]),.dinb(w_n3354_0[1]),.dout(n3427),.clk(gclk));
	jor g3346(.dina(w_n3238_4[2]),.dinb(w_n2797_1[0]),.dout(n3428),.clk(gclk));
	jor g3347(.dina(w_n3322_5[1]),.dinb(w_n2678_3[1]),.dout(n3429),.clk(gclk));
	jor g3348(.dina(w_n3325_3[2]),.dinb(w_n2681_2[0]),.dout(n3430),.clk(gclk));
	jor g3349(.dina(w_n3328_4[0]),.dinb(w_n2687_3[0]),.dout(n3431),.clk(gclk));
	jand g3350(.dina(n3431),.dinb(n3430),.dout(n3432),.clk(gclk));
	jand g3351(.dina(n3432),.dinb(n3429),.dout(n3433),.clk(gclk));
	jand g3352(.dina(n3433),.dinb(n3428),.dout(n3434),.clk(gclk));
	jxor g3353(.dina(n3434),.dinb(w_n3233_7[0]),.dout(n3435),.clk(gclk));
	jor g3354(.dina(w_n3435_0[1]),.dinb(n3427),.dout(n3436),.clk(gclk));
	jand g3355(.dina(n3436),.dinb(w_n3426_0[1]),.dout(n3437),.clk(gclk));
	jand g3356(.dina(w_n3437_0[1]),.dinb(w_n3353_0[2]),.dout(n3438),.clk(gclk));
	jor g3357(.dina(w_n3437_0[0]),.dinb(w_n3353_0[1]),.dout(n3439),.clk(gclk));
	jand g3358(.dina(w_n3237_1[2]),.dinb(w_n3004_1[0]),.dout(n3440),.clk(gclk));
	jor g3359(.dina(w_n3322_5[0]),.dinb(w_n2674_2[1]),.dout(n3441),.clk(gclk));
	jand g3360(.dina(w_n3324_1[2]),.dinb(w_n2679_2[1]),.dout(n3442),.clk(gclk));
	jnot g3361(.din(n3442),.dout(n3443),.clk(gclk));
	jand g3362(.dina(n3443),.dinb(n3441),.dout(n3444),.clk(gclk));
	jnot g3363(.din(n3444),.dout(n3445),.clk(gclk));
	jor g3364(.dina(n3445),.dinb(n3440),.dout(n3446),.clk(gclk));
	jand g3365(.dina(w_n3446_0[1]),.dinb(w_n3233_6[2]),.dout(n3447),.clk(gclk));
	jand g3366(.dina(w_n2684_3[0]),.dinb(w_n63_1[2]),.dout(n3448),.clk(gclk));
	jor g3367(.dina(n3448),.dinb(w_n3233_6[1]),.dout(n3449),.clk(gclk));
	jor g3368(.dina(n3449),.dinb(w_n3446_0[0]),.dout(n3450),.clk(gclk));
	jnot g3369(.din(n3450),.dout(n3451),.clk(gclk));
	jor g3370(.dina(n3451),.dinb(n3447),.dout(n3452),.clk(gclk));
	jand g3371(.dina(w_n3452_0[1]),.dinb(n3439),.dout(n3453),.clk(gclk));
	jor g3372(.dina(n3453),.dinb(w_n3438_0[1]),.dout(n3454),.clk(gclk));
	jand g3373(.dina(w_n3454_0[1]),.dinb(w_n3352_0[2]),.dout(n3455),.clk(gclk));
	jor g3374(.dina(w_n3454_0[0]),.dinb(w_n3352_0[1]),.dout(n3456),.clk(gclk));
	jor g3375(.dina(w_n3238_4[1]),.dinb(w_n3028_1[0]),.dout(n3457),.clk(gclk));
	jor g3376(.dina(w_n3322_4[2]),.dinb(w_n2671_4[0]),.dout(n3458),.clk(gclk));
	jor g3377(.dina(w_n3325_3[1]),.dinb(w_n2674_2[0]),.dout(n3459),.clk(gclk));
	jor g3378(.dina(w_n3328_3[2]),.dinb(w_n2678_3[0]),.dout(n3460),.clk(gclk));
	jand g3379(.dina(n3460),.dinb(n3459),.dout(n3461),.clk(gclk));
	jand g3380(.dina(n3461),.dinb(n3458),.dout(n3462),.clk(gclk));
	jand g3381(.dina(n3462),.dinb(n3457),.dout(n3463),.clk(gclk));
	jxor g3382(.dina(n3463),.dinb(w_n3233_6[0]),.dout(n3464),.clk(gclk));
	jand g3383(.dina(w_n3464_0[1]),.dinb(n3456),.dout(n3465),.clk(gclk));
	jor g3384(.dina(n3465),.dinb(w_n3455_0[1]),.dout(n3466),.clk(gclk));
	jand g3385(.dina(w_n3466_0[1]),.dinb(w_n3351_0[2]),.dout(n3467),.clk(gclk));
	jor g3386(.dina(w_n3466_0[0]),.dinb(w_n3351_0[1]),.dout(n3468),.clk(gclk));
	jand g3387(.dina(w_n3237_1[1]),.dinb(w_n3016_1[1]),.dout(n3469),.clk(gclk));
	jnot g3388(.din(n3469),.dout(n3470),.clk(gclk));
	jor g3389(.dina(w_n3322_4[1]),.dinb(w_n2669_2[2]),.dout(n3471),.clk(gclk));
	jand g3390(.dina(w_n3324_1[1]),.dinb(w_n2672_2[0]),.dout(n3472),.clk(gclk));
	jnot g3391(.din(n3472),.dout(n3473),.clk(gclk));
	jand g3392(.dina(n3473),.dinb(n3471),.dout(n3474),.clk(gclk));
	jand g3393(.dina(n3474),.dinb(n3470),.dout(n3475),.clk(gclk));
	jnot g3394(.din(w_n3475_0[1]),.dout(n3476),.clk(gclk));
	jand g3395(.dina(n3476),.dinb(w_n3233_5[2]),.dout(n3477),.clk(gclk));
	jand g3396(.dina(w_n2677_3[1]),.dinb(w_n63_1[1]),.dout(n3478),.clk(gclk));
	jor g3397(.dina(n3478),.dinb(w_n3233_5[1]),.dout(n3479),.clk(gclk));
	jnot g3398(.din(n3479),.dout(n3480),.clk(gclk));
	jand g3399(.dina(n3480),.dinb(w_n3475_0[0]),.dout(n3481),.clk(gclk));
	jor g3400(.dina(n3481),.dinb(n3477),.dout(n3482),.clk(gclk));
	jand g3401(.dina(w_n3482_0[1]),.dinb(n3468),.dout(n3483),.clk(gclk));
	jor g3402(.dina(n3483),.dinb(w_n3467_0[1]),.dout(n3484),.clk(gclk));
	jor g3403(.dina(w_n3484_0[1]),.dinb(w_n3350_0[2]),.dout(n3485),.clk(gclk));
	jand g3404(.dina(w_n3484_0[0]),.dinb(w_n3350_0[1]),.dout(n3486),.clk(gclk));
	jor g3405(.dina(w_n3238_4[0]),.dinb(w_n2771_1[1]),.dout(n3487),.clk(gclk));
	jor g3406(.dina(w_n3322_4[0]),.dinb(w_n2773_4[0]),.dout(n3488),.clk(gclk));
	jor g3407(.dina(w_n3325_3[0]),.dinb(w_n2669_2[1]),.dout(n3489),.clk(gclk));
	jor g3408(.dina(w_n3328_3[1]),.dinb(w_n2671_3[2]),.dout(n3490),.clk(gclk));
	jand g3409(.dina(n3490),.dinb(n3489),.dout(n3491),.clk(gclk));
	jand g3410(.dina(n3491),.dinb(n3488),.dout(n3492),.clk(gclk));
	jand g3411(.dina(n3492),.dinb(n3487),.dout(n3493),.clk(gclk));
	jxor g3412(.dina(n3493),.dinb(w_n3233_5[0]),.dout(n3494),.clk(gclk));
	jor g3413(.dina(w_n3494_0[1]),.dinb(n3486),.dout(n3495),.clk(gclk));
	jand g3414(.dina(n3495),.dinb(w_n3485_0[1]),.dout(n3496),.clk(gclk));
	jand g3415(.dina(w_n3496_0[1]),.dinb(w_n3349_0[2]),.dout(n3497),.clk(gclk));
	jor g3416(.dina(w_n3496_0[0]),.dinb(w_n3349_0[1]),.dout(n3498),.clk(gclk));
	jand g3417(.dina(w_n3237_1[0]),.dinb(w_n3174_1[1]),.dout(n3499),.clk(gclk));
	jnot g3418(.din(w_n3322_3[2]),.dout(n3500),.clk(gclk));
	jand g3419(.dina(n3500),.dinb(w_n3176_2[0]),.dout(n3501),.clk(gclk));
	jand g3420(.dina(w_n3324_1[0]),.dinb(w_n2769_2[2]),.dout(n3502),.clk(gclk));
	jor g3421(.dina(n3502),.dinb(n3501),.dout(n3503),.clk(gclk));
	jor g3422(.dina(n3503),.dinb(n3499),.dout(n3504),.clk(gclk));
	jand g3423(.dina(w_n3504_0[1]),.dinb(w_n3233_4[2]),.dout(n3505),.clk(gclk));
	jand g3424(.dina(w_n2670_4[0]),.dinb(w_n63_1[0]),.dout(n3506),.clk(gclk));
	jor g3425(.dina(n3506),.dinb(w_n3233_4[1]),.dout(n3507),.clk(gclk));
	jor g3426(.dina(n3507),.dinb(w_n3504_0[0]),.dout(n3508),.clk(gclk));
	jnot g3427(.din(n3508),.dout(n3509),.clk(gclk));
	jor g3428(.dina(n3509),.dinb(n3505),.dout(n3510),.clk(gclk));
	jand g3429(.dina(w_n3510_0[1]),.dinb(n3498),.dout(n3511),.clk(gclk));
	jor g3430(.dina(n3511),.dinb(w_n3497_0[1]),.dout(n3512),.clk(gclk));
	jor g3431(.dina(w_n3512_0[1]),.dinb(w_n3348_0[2]),.dout(n3513),.clk(gclk));
	jand g3432(.dina(w_n3512_0[0]),.dinb(w_n3348_0[1]),.dout(n3514),.clk(gclk));
	jnot g3433(.din(w_n3291_0[0]),.dout(n3515),.clk(gclk));
	jxor g3434(.dina(w_n3294_0[0]),.dinb(n3515),.dout(n3516),.clk(gclk));
	jor g3435(.dina(w_n3516_1[2]),.dinb(w_n3238_3[2]),.dout(n3517),.clk(gclk));
	jor g3436(.dina(w_n3322_3[1]),.dinb(w_n3284_7[0]),.dout(n3518),.clk(gclk));
	jor g3437(.dina(w_n3325_2[2]),.dinb(w_n3172_4[2]),.dout(n3519),.clk(gclk));
	jor g3438(.dina(w_n3328_3[0]),.dinb(w_n2773_3[2]),.dout(n3520),.clk(gclk));
	jand g3439(.dina(n3520),.dinb(n3519),.dout(n3521),.clk(gclk));
	jand g3440(.dina(n3521),.dinb(n3518),.dout(n3522),.clk(gclk));
	jand g3441(.dina(n3522),.dinb(n3517),.dout(n3523),.clk(gclk));
	jxor g3442(.dina(n3523),.dinb(w_n68_5[2]),.dout(n3524),.clk(gclk));
	jnot g3443(.din(w_n3524_0[1]),.dout(n3525),.clk(gclk));
	jor g3444(.dina(n3525),.dinb(n3514),.dout(n3526),.clk(gclk));
	jand g3445(.dina(n3526),.dinb(w_n3513_0[1]),.dout(n3527),.clk(gclk));
	jand g3446(.dina(n3527),.dinb(w_n3347_0[1]),.dout(n3528),.clk(gclk));
	jor g3447(.dina(w_n3528_0[1]),.dinb(n3346),.dout(n3529),.clk(gclk));
	jxor g3448(.dina(w_n3333_0[0]),.dinb(w_n3232_0[0]),.dout(n3530),.clk(gclk));
	jand g3449(.dina(w_n3530_0[1]),.dinb(w_n3529_0[1]),.dout(n3531),.clk(gclk));
	jor g3450(.dina(n3531),.dinb(n3334),.dout(n3532),.clk(gclk));
	jand g3451(.dina(w_n3230_0[0]),.dinb(w_n3183_0[0]),.dout(n3533),.clk(gclk));
	jand g3452(.dina(w_n3231_0[0]),.dinb(w_n3145_0[0]),.dout(n3534),.clk(gclk));
	jor g3453(.dina(n3534),.dinb(n3533),.dout(n3535),.clk(gclk));
	jor g3454(.dina(w_n3516_1[1]),.dinb(w_n79_4[0]),.dout(n3536),.clk(gclk));
	jor g3455(.dina(w_n3284_6[2]),.dinb(w_n2775_3[1]),.dout(n3537),.clk(gclk));
	jor g3456(.dina(w_n3172_4[1]),.dinb(w_n2780_3[1]),.dout(n3538),.clk(gclk));
	jor g3457(.dina(w_n2784_4[0]),.dinb(w_n2773_3[1]),.dout(n3539),.clk(gclk));
	jand g3458(.dina(n3539),.dinb(n3538),.dout(n3540),.clk(gclk));
	jand g3459(.dina(n3540),.dinb(n3537),.dout(n3541),.clk(gclk));
	jand g3460(.dina(n3541),.dinb(n3536),.dout(n3542),.clk(gclk));
	jxor g3461(.dina(n3542),.dinb(w_n56_6[0]),.dout(n3543),.clk(gclk));
	jand g3462(.dina(w_n3228_0[0]),.dinb(w_n3220_0[0]),.dout(n3544),.clk(gclk));
	jand g3463(.dina(w_n3229_0[0]),.dinb(w_n3186_0[0]),.dout(n3545),.clk(gclk));
	jor g3464(.dina(n3545),.dinb(n3544),.dout(n3546),.clk(gclk));
	jand g3465(.dina(w_n3016_1[0]),.dinb(w_n2794_1[1]),.dout(n3547),.clk(gclk));
	jand g3466(.dina(w_n2799_1[0]),.dinb(w_n2670_3[2]),.dout(n3548),.clk(gclk));
	jand g3467(.dina(w_n2808_1[1]),.dinb(w_n2677_3[0]),.dout(n3549),.clk(gclk));
	jand g3468(.dina(w_n2804_1[1]),.dinb(w_n2672_1[2]),.dout(n3550),.clk(gclk));
	jor g3469(.dina(n3550),.dinb(n3549),.dout(n3551),.clk(gclk));
	jor g3470(.dina(n3551),.dinb(n3548),.dout(n3552),.clk(gclk));
	jor g3471(.dina(n3552),.dinb(n3547),.dout(n3553),.clk(gclk));
	jxor g3472(.dina(n3553),.dinb(w_n699_7[0]),.dout(n3554),.clk(gclk));
	jand g3473(.dina(w_n3218_0[0]),.dinb(w_n3197_0[0]),.dout(n3555),.clk(gclk));
	jand g3474(.dina(w_n3219_0[0]),.dinb(w_n3189_0[0]),.dout(n3556),.clk(gclk));
	jor g3475(.dina(n3556),.dinb(n3555),.dout(n3557),.clk(gclk));
	jor g3476(.dina(w_n2857_5[0]),.dinb(w_n2797_0[2]),.dout(n3558),.clk(gclk));
	jor g3477(.dina(w_n2860_4[1]),.dinb(w_n2678_2[2]),.dout(n3559),.clk(gclk));
	jor g3478(.dina(w_n2865_4[1]),.dinb(w_n2681_1[2]),.dout(n3560),.clk(gclk));
	jor g3479(.dina(w_n2863_5[0]),.dinb(w_n2687_2[2]),.dout(n3561),.clk(gclk));
	jand g3480(.dina(n3561),.dinb(n3560),.dout(n3562),.clk(gclk));
	jand g3481(.dina(n3562),.dinb(n3559),.dout(n3563),.clk(gclk));
	jand g3482(.dina(n3563),.dinb(n3558),.dout(n3564),.clk(gclk));
	jxor g3483(.dina(n3564),.dinb(w_n808_7[2]),.dout(n3565),.clk(gclk));
	jand g3484(.dina(w_n3217_0[0]),.dinb(w_n3210_0[0]),.dout(n3566),.clk(gclk));
	jor g3485(.dina(n3566),.dinb(w_n3215_0[0]),.dout(n3567),.clk(gclk));
	jand g3486(.dina(w_n2862_0[2]),.dinb(w_n954_18[1]),.dout(n3568),.clk(gclk));
	jnot g3487(.din(n3568),.dout(n3569),.clk(gclk));
	jor g3488(.dina(w_n3198_5[1]),.dinb(w_n2874_0[1]),.dout(n3570),.clk(gclk));
	jnot g3489(.din(w_n2688_3[0]),.dout(n3571),.clk(gclk));
	jand g3490(.dina(w_n2889_3[1]),.dinb(w_n3571_1[1]),.dout(n3572),.clk(gclk));
	jnot g3491(.din(w_n2691_3[0]),.dout(n3573),.clk(gclk));
	jand g3492(.dina(w_n2887_3[2]),.dinb(w_n3573_0[2]),.dout(n3574),.clk(gclk));
	jand g3493(.dina(w_n2995_4[0]),.dinb(w_n2693_1[2]),.dout(n3575),.clk(gclk));
	jor g3494(.dina(n3575),.dinb(n3574),.dout(n3576),.clk(gclk));
	jor g3495(.dina(n3576),.dinb(n3572),.dout(n3577),.clk(gclk));
	jnot g3496(.din(n3577),.dout(n3578),.clk(gclk));
	jand g3497(.dina(n3578),.dinb(n3570),.dout(n3579),.clk(gclk));
	jxor g3498(.dina(w_n3579_0[1]),.dinb(n3569),.dout(n3580),.clk(gclk));
	jxor g3499(.dina(w_n3580_0[1]),.dinb(w_n3567_0[1]),.dout(n3581),.clk(gclk));
	jxor g3500(.dina(w_n3581_0[1]),.dinb(w_n3565_0[1]),.dout(n3582),.clk(gclk));
	jxor g3501(.dina(w_n3582_0[1]),.dinb(w_n3557_0[1]),.dout(n3583),.clk(gclk));
	jxor g3502(.dina(w_n3583_0[1]),.dinb(w_n3554_0[1]),.dout(n3584),.clk(gclk));
	jxor g3503(.dina(w_n3584_0[1]),.dinb(w_n3546_0[1]),.dout(n3585),.clk(gclk));
	jxor g3504(.dina(w_n3585_0[1]),.dinb(w_n3543_0[1]),.dout(n3586),.clk(gclk));
	jxor g3505(.dina(w_n3586_0[1]),.dinb(w_n3535_0[1]),.dout(n3587),.clk(gclk));
	jnot g3506(.din(w_n3319_0[0]),.dout(n3588),.clk(gclk));
	jand g3507(.dina(n3588),.dinb(w_n3301_0[0]),.dout(n3589),.clk(gclk));
	jor g3508(.dina(n3589),.dinb(w_n3317_0[0]),.dout(n3590),.clk(gclk));
	jand g3509(.dina(w_n3314_0[0]),.dinb(w_n3303_0[0]),.dout(n3591),.clk(gclk));
	jand g3510(.dina(w_n786_0[2]),.dinb(w_n403_0[0]),.dout(n3592),.clk(gclk));
	jnot g3511(.din(w_n136_0[0]),.dout(n3593),.clk(gclk));
	jand g3512(.dina(w_n751_1[1]),.dinb(n3593),.dout(n3594),.clk(gclk));
	jand g3513(.dina(n3594),.dinb(w_n246_0[0]),.dout(n3595),.clk(gclk));
	jand g3514(.dina(n3595),.dinb(w_n776_0[0]),.dout(n3596),.clk(gclk));
	jand g3515(.dina(w_n719_0[1]),.dinb(w_n308_0[0]),.dout(n3597),.clk(gclk));
	jand g3516(.dina(n3597),.dinb(n3596),.dout(n3598),.clk(gclk));
	jand g3517(.dina(n3598),.dinb(w_n3592_0[1]),.dout(n3599),.clk(gclk));
	jxor g3518(.dina(w_n3599_0[2]),.dinb(w_n3591_0[1]),.dout(n3600),.clk(gclk));
	jnot g3519(.din(w_n3600_8[2]),.dout(n3601),.clk(gclk));
	jand g3520(.dina(w_n3601_1[1]),.dinb(w_n3316_0[1]),.dout(n3602),.clk(gclk));
	jand g3521(.dina(w_n3599_0[1]),.dinb(w_n3315_7[0]),.dout(n3603),.clk(gclk));
	jor g3522(.dina(n3603),.dinb(w_n3602_0[1]),.dout(n3604),.clk(gclk));
	jxor g3523(.dina(w_n3604_0[1]),.dinb(w_n3590_0[1]),.dout(n3605),.clk(gclk));
	jor g3524(.dina(w_n3605_1[2]),.dinb(w_n3238_3[1]),.dout(n3606),.clk(gclk));
	jor g3525(.dina(w_n3600_8[1]),.dinb(w_n3322_3[0]),.dout(n3607),.clk(gclk));
	jor g3526(.dina(w_n3325_2[1]),.dinb(w_n3315_6[2]),.dout(n3608),.clk(gclk));
	jor g3527(.dina(w_n3328_2[2]),.dinb(w_n3283_6[2]),.dout(n3609),.clk(gclk));
	jand g3528(.dina(n3609),.dinb(n3608),.dout(n3610),.clk(gclk));
	jand g3529(.dina(n3610),.dinb(n3607),.dout(n3611),.clk(gclk));
	jand g3530(.dina(n3611),.dinb(n3606),.dout(n3612),.clk(gclk));
	jxor g3531(.dina(n3612),.dinb(w_n3233_4[0]),.dout(n3613),.clk(gclk));
	jxor g3532(.dina(w_n3613_0[1]),.dinb(w_n3587_0[1]),.dout(n3614),.clk(gclk));
	jxor g3533(.dina(w_n3614_0[1]),.dinb(w_n3532_0[1]),.dout(n3615),.clk(gclk));
	jnot g3534(.din(w_n3615_0[1]),.dout(n3616),.clk(gclk));
	jand g3535(.dina(w_n312_1[0]),.dinb(w_n147_2[1]),.dout(n3617),.clk(gclk));
	jand g3536(.dina(w_n751_1[0]),.dinb(w_n612_1[0]),.dout(n3618),.clk(gclk));
	jand g3537(.dina(n3618),.dinb(n3617),.dout(n3619),.clk(gclk));
	jand g3538(.dina(n3619),.dinb(w_n2490_0[0]),.dout(n3620),.clk(gclk));
	jand g3539(.dina(w_n249_1[0]),.dinb(w_n214_1[2]),.dout(n3621),.clk(gclk));
	jand g3540(.dina(w_n422_1[1]),.dinb(w_n232_0[2]),.dout(n3622),.clk(gclk));
	jand g3541(.dina(n3622),.dinb(n3621),.dout(n3623),.clk(gclk));
	jand g3542(.dina(w_n445_1[0]),.dinb(w_n368_1[0]),.dout(n3624),.clk(gclk));
	jand g3543(.dina(w_n3624_0[2]),.dinb(w_n877_0[0]),.dout(n3625),.clk(gclk));
	jand g3544(.dina(w_n285_0[2]),.dinb(w_n138_1[2]),.dout(n3626),.clk(gclk));
	jand g3545(.dina(w_n3626_0[1]),.dinb(w_n2326_0[1]),.dout(n3627),.clk(gclk));
	jand g3546(.dina(n3627),.dinb(n3625),.dout(n3628),.clk(gclk));
	jand g3547(.dina(n3628),.dinb(n3623),.dout(n3629),.clk(gclk));
	jand g3548(.dina(n3629),.dinb(w_n3620_0[1]),.dout(n3630),.clk(gclk));
	jand g3549(.dina(w_n426_1[0]),.dinb(w_n421_2[0]),.dout(n3631),.clk(gclk));
	jand g3550(.dina(n3631),.dinb(w_n1641_0[0]),.dout(n3632),.clk(gclk));
	jand g3551(.dina(n3632),.dinb(w_n3630_0[1]),.dout(n3633),.clk(gclk));
	jnot g3552(.din(w_n165_0[0]),.dout(n3634),.clk(gclk));
	jand g3553(.dina(w_n454_1[0]),.dinb(w_n295_1[1]),.dout(n3635),.clk(gclk));
	jand g3554(.dina(n3635),.dinb(w_n3634_0[1]),.dout(n3636),.clk(gclk));
	jand g3555(.dina(n3636),.dinb(w_n3250_0[0]),.dout(n3637),.clk(gclk));
	jand g3556(.dina(n3637),.dinb(w_n852_0[0]),.dout(n3638),.clk(gclk));
	jand g3557(.dina(w_n243_1[2]),.dinb(w_n130_1[0]),.dout(n3639),.clk(gclk));
	jand g3558(.dina(w_n592_2[0]),.dinb(w_n270_1[1]),.dout(n3640),.clk(gclk));
	jand g3559(.dina(n3640),.dinb(n3639),.dout(n3641),.clk(gclk));
	jand g3560(.dina(w_n2736_1[0]),.dinb(w_n626_0[1]),.dout(n3642),.clk(gclk));
	jand g3561(.dina(n3642),.dinb(n3641),.dout(n3643),.clk(gclk));
	jand g3562(.dina(w_n734_0[1]),.dinb(w_n370_0[2]),.dout(n3644),.clk(gclk));
	jand g3563(.dina(n3644),.dinb(w_n772_1[0]),.dout(n3645),.clk(gclk));
	jand g3564(.dina(n3645),.dinb(w_n3258_1[1]),.dout(n3646),.clk(gclk));
	jand g3565(.dina(n3646),.dinb(n3643),.dout(n3647),.clk(gclk));
	jand g3566(.dina(n3647),.dinb(w_n832_0[2]),.dout(n3648),.clk(gclk));
	jand g3567(.dina(n3648),.dinb(w_n3638_0[1]),.dout(n3649),.clk(gclk));
	jand g3568(.dina(n3649),.dinb(w_n3633_0[1]),.dout(n3650),.clk(gclk));
	jor g3569(.dina(w_n3650_0[1]),.dinb(n3616),.dout(n3651),.clk(gclk));
	jxor g3570(.dina(w_n3650_0[0]),.dinb(w_n3615_0[0]),.dout(n3652),.clk(gclk));
	jnot g3571(.din(w_n3530_0[0]),.dout(n3653),.clk(gclk));
	jxor g3572(.dina(n3653),.dinb(w_n3529_0[0]),.dout(n3654),.clk(gclk));
	jand g3573(.dina(w_n837_0[2]),.dinb(w_n264_1[1]),.dout(n3655),.clk(gclk));
	jand g3574(.dina(w_n422_1[0]),.dinb(w_n383_1[0]),.dout(n3656),.clk(gclk));
	jand g3575(.dina(n3656),.dinb(n3655),.dout(n3657),.clk(gclk));
	jand g3576(.dina(n3657),.dinb(w_n771_1[0]),.dout(n3658),.clk(gclk));
	jand g3577(.dina(w_n473_0[2]),.dinb(w_n351_1[0]),.dout(n3659),.clk(gclk));
	jand g3578(.dina(n3659),.dinb(w_n430_1[0]),.dout(n3660),.clk(gclk));
	jand g3579(.dina(n3660),.dinb(w_n2442_0[0]),.dout(n3661),.clk(gclk));
	jand g3580(.dina(n3661),.dinb(n3658),.dout(n3662),.clk(gclk));
	jand g3581(.dina(n3662),.dinb(w_n1292_0[0]),.dout(n3663),.clk(gclk));
	jand g3582(.dina(w_n768_1[0]),.dinb(w_n216_1[2]),.dout(n3664),.clk(gclk));
	jand g3583(.dina(n3664),.dinb(w_n942_0[0]),.dout(n3665),.clk(gclk));
	jand g3584(.dina(n3665),.dinb(w_n3663_0[1]),.dout(n3666),.clk(gclk));
	jand g3585(.dina(w_n772_0[2]),.dinb(w_n358_1[0]),.dout(n3667),.clk(gclk));
	jand g3586(.dina(n3667),.dinb(w_n515_0[2]),.dout(n3668),.clk(gclk));
	jand g3587(.dina(n3668),.dinb(w_n943_0[0]),.dout(n3669),.clk(gclk));
	jand g3588(.dina(w_n412_1[0]),.dinb(w_n372_1[0]),.dout(n3670),.clk(gclk));
	jand g3589(.dina(w_n451_1[1]),.dinb(w_n282_1[1]),.dout(n3671),.clk(gclk));
	jand g3590(.dina(n3671),.dinb(n3670),.dout(n3672),.clk(gclk));
	jand g3591(.dina(w_n3263_0[0]),.dinb(w_n906_0[0]),.dout(n3673),.clk(gclk));
	jand g3592(.dina(n3673),.dinb(w_n938_0[0]),.dout(n3674),.clk(gclk));
	jand g3593(.dina(n3674),.dinb(n3672),.dout(n3675),.clk(gclk));
	jand g3594(.dina(n3675),.dinb(w_n3669_0[1]),.dout(n3676),.clk(gclk));
	jnot g3595(.din(w_n1676_0[0]),.dout(n3677),.clk(gclk));
	jand g3596(.dina(n3677),.dinb(w_n463_1[2]),.dout(n3678),.clk(gclk));
	jand g3597(.dina(w_n594_1[0]),.dinb(w_n436_1[0]),.dout(n3679),.clk(gclk));
	jand g3598(.dina(n3679),.dinb(w_n1228_0[0]),.dout(n3680),.clk(gclk));
	jand g3599(.dina(w_n1196_0[0]),.dinb(w_n619_1[0]),.dout(n3681),.clk(gclk));
	jand g3600(.dina(n3681),.dinb(n3680),.dout(n3682),.clk(gclk));
	jand g3601(.dina(n3682),.dinb(n3678),.dout(n3683),.clk(gclk));
	jand g3602(.dina(n3683),.dinb(w_n2544_0[0]),.dout(n3684),.clk(gclk));
	jand g3603(.dina(n3684),.dinb(w_n3676_0[1]),.dout(n3685),.clk(gclk));
	jand g3604(.dina(n3685),.dinb(w_n3666_0[1]),.dout(n3686),.clk(gclk));
	jand g3605(.dina(w_n3686_0[1]),.dinb(w_n3654_0[1]),.dout(n3687),.clk(gclk));
	jor g3606(.dina(w_n3686_0[0]),.dinb(w_n3654_0[0]),.dout(n3688),.clk(gclk));
	jand g3607(.dina(w_n710_1[1]),.dinb(w_n256_0[2]),.dout(n3689),.clk(gclk));
	jand g3608(.dina(n3689),.dinb(w_n280_0[2]),.dout(n3690),.clk(gclk));
	jand g3609(.dina(n3690),.dinb(w_n1673_0[0]),.dout(n3691),.clk(gclk));
	jand g3610(.dina(n3691),.dinb(w_n2372_0[0]),.dout(n3692),.clk(gclk));
	jand g3611(.dina(n3692),.dinb(w_n2398_0[0]),.dout(n3693),.clk(gclk));
	jand g3612(.dina(w_n321_0[2]),.dinb(w_n467_0[1]),.dout(n3694),.clk(gclk));
	jand g3613(.dina(n3694),.dinb(w_n2745_0[0]),.dout(n3695),.clk(gclk));
	jand g3614(.dina(n3695),.dinb(w_n932_0[0]),.dout(n3696),.clk(gclk));
	jand g3615(.dina(w_n2515_0[0]),.dinb(w_n992_0[2]),.dout(n3697),.clk(gclk));
	jand g3616(.dina(w_n2521_1[0]),.dinb(w_n728_0[0]),.dout(n3698),.clk(gclk));
	jand g3617(.dina(n3698),.dinb(n3697),.dout(n3699),.clk(gclk));
	jand g3618(.dina(w_n214_1[1]),.dinb(w_n138_1[1]),.dout(n3700),.clk(gclk));
	jand g3619(.dina(n3700),.dinb(w_n153_0[1]),.dout(n3701),.clk(gclk));
	jand g3620(.dina(w_n441_0[1]),.dinb(w_n304_1[0]),.dout(n3702),.clk(gclk));
	jand g3621(.dina(w_n488_1[0]),.dinb(w_n261_0[1]),.dout(n3703),.clk(gclk));
	jand g3622(.dina(n3703),.dinb(n3702),.dout(n3704),.clk(gclk));
	jand g3623(.dina(n3704),.dinb(n3701),.dout(n3705),.clk(gclk));
	jand g3624(.dina(n3705),.dinb(n3699),.dout(n3706),.clk(gclk));
	jand g3625(.dina(n3706),.dinb(w_n2466_0[0]),.dout(n3707),.clk(gclk));
	jand g3626(.dina(n3707),.dinb(w_n3696_0[1]),.dout(n3708),.clk(gclk));
	jand g3627(.dina(n3708),.dinb(w_n3693_0[2]),.dout(n3709),.clk(gclk));
	jnot g3628(.din(w_n3347_0[0]),.dout(n3710),.clk(gclk));
	jnot g3629(.din(w_n3513_0[0]),.dout(n3711),.clk(gclk));
	jnot g3630(.din(w_n3348_0[0]),.dout(n3712),.clk(gclk));
	jnot g3631(.din(w_n3497_0[0]),.dout(n3713),.clk(gclk));
	jnot g3632(.din(w_n3349_0[0]),.dout(n3714),.clk(gclk));
	jnot g3633(.din(w_n3485_0[0]),.dout(n3715),.clk(gclk));
	jnot g3634(.din(w_n3350_0[0]),.dout(n3716),.clk(gclk));
	jnot g3635(.din(w_n3467_0[0]),.dout(n3717),.clk(gclk));
	jnot g3636(.din(w_n3351_0[0]),.dout(n3718),.clk(gclk));
	jnot g3637(.din(w_n3455_0[0]),.dout(n3719),.clk(gclk));
	jnot g3638(.din(w_n3352_0[0]),.dout(n3720),.clk(gclk));
	jnot g3639(.din(w_n3438_0[0]),.dout(n3721),.clk(gclk));
	jnot g3640(.din(w_n3353_0[0]),.dout(n3722),.clk(gclk));
	jnot g3641(.din(w_n3426_0[0]),.dout(n3723),.clk(gclk));
	jnot g3642(.din(w_n3354_0[0]),.dout(n3724),.clk(gclk));
	jnot g3643(.din(w_n3421_0[0]),.dout(n3725),.clk(gclk));
	jnot g3644(.din(w_n3362_0[0]),.dout(n3726),.clk(gclk));
	jnot g3645(.din(w_n3409_0[0]),.dout(n3727),.clk(gclk));
	jnot g3646(.din(w_n3365_0[0]),.dout(n3728),.clk(gclk));
	jnot g3647(.din(w_n3397_0[0]),.dout(n3729),.clk(gclk));
	jnot g3648(.din(w_n3367_0[0]),.dout(n3730),.clk(gclk));
	jnot g3649(.din(w_n3379_0[0]),.dout(n3731),.clk(gclk));
	jand g3650(.dina(w_n3375_0[0]),.dinb(w_n68_5[1]),.dout(n3732),.clk(gclk));
	jnot g3651(.din(w_n3394_0[0]),.dout(n3733),.clk(gclk));
	jor g3652(.dina(n3733),.dinb(n3732),.dout(n3734),.clk(gclk));
	jor g3653(.dina(n3734),.dinb(n3731),.dout(n3735),.clk(gclk));
	jand g3654(.dina(n3735),.dinb(n3730),.dout(n3736),.clk(gclk));
	jnot g3655(.din(w_n3406_0[0]),.dout(n3737),.clk(gclk));
	jor g3656(.dina(n3737),.dinb(n3736),.dout(n3738),.clk(gclk));
	jand g3657(.dina(n3738),.dinb(n3729),.dout(n3739),.clk(gclk));
	jor g3658(.dina(n3739),.dinb(n3728),.dout(n3740),.clk(gclk));
	jnot g3659(.din(w_n3418_0[0]),.dout(n3741),.clk(gclk));
	jand g3660(.dina(n3741),.dinb(n3740),.dout(n3742),.clk(gclk));
	jor g3661(.dina(n3742),.dinb(n3727),.dout(n3743),.clk(gclk));
	jand g3662(.dina(n3743),.dinb(n3726),.dout(n3744),.clk(gclk));
	jnot g3663(.din(w_n3423_0[0]),.dout(n3745),.clk(gclk));
	jor g3664(.dina(n3745),.dinb(n3744),.dout(n3746),.clk(gclk));
	jand g3665(.dina(n3746),.dinb(n3725),.dout(n3747),.clk(gclk));
	jor g3666(.dina(n3747),.dinb(n3724),.dout(n3748),.clk(gclk));
	jnot g3667(.din(w_n3435_0[0]),.dout(n3749),.clk(gclk));
	jand g3668(.dina(n3749),.dinb(n3748),.dout(n3750),.clk(gclk));
	jor g3669(.dina(n3750),.dinb(n3723),.dout(n3751),.clk(gclk));
	jand g3670(.dina(n3751),.dinb(n3722),.dout(n3752),.clk(gclk));
	jnot g3671(.din(w_n3452_0[0]),.dout(n3753),.clk(gclk));
	jor g3672(.dina(n3753),.dinb(n3752),.dout(n3754),.clk(gclk));
	jand g3673(.dina(n3754),.dinb(n3721),.dout(n3755),.clk(gclk));
	jand g3674(.dina(n3755),.dinb(n3720),.dout(n3756),.clk(gclk));
	jnot g3675(.din(w_n3464_0[0]),.dout(n3757),.clk(gclk));
	jor g3676(.dina(n3757),.dinb(n3756),.dout(n3758),.clk(gclk));
	jand g3677(.dina(n3758),.dinb(n3719),.dout(n3759),.clk(gclk));
	jand g3678(.dina(n3759),.dinb(n3718),.dout(n3760),.clk(gclk));
	jnot g3679(.din(w_n3482_0[0]),.dout(n3761),.clk(gclk));
	jor g3680(.dina(n3761),.dinb(n3760),.dout(n3762),.clk(gclk));
	jand g3681(.dina(n3762),.dinb(n3717),.dout(n3763),.clk(gclk));
	jor g3682(.dina(n3763),.dinb(n3716),.dout(n3764),.clk(gclk));
	jnot g3683(.din(w_n3494_0[0]),.dout(n3765),.clk(gclk));
	jand g3684(.dina(n3765),.dinb(n3764),.dout(n3766),.clk(gclk));
	jor g3685(.dina(n3766),.dinb(n3715),.dout(n3767),.clk(gclk));
	jand g3686(.dina(n3767),.dinb(n3714),.dout(n3768),.clk(gclk));
	jnot g3687(.din(w_n3510_0[0]),.dout(n3769),.clk(gclk));
	jor g3688(.dina(n3769),.dinb(n3768),.dout(n3770),.clk(gclk));
	jand g3689(.dina(n3770),.dinb(n3713),.dout(n3771),.clk(gclk));
	jor g3690(.dina(n3771),.dinb(n3712),.dout(n3772),.clk(gclk));
	jand g3691(.dina(w_n3524_0[0]),.dinb(n3772),.dout(n3773),.clk(gclk));
	jor g3692(.dina(n3773),.dinb(n3711),.dout(n3774),.clk(gclk));
	jand g3693(.dina(n3774),.dinb(n3710),.dout(n3775),.clk(gclk));
	jor g3694(.dina(n3775),.dinb(n3709),.dout(n3776),.clk(gclk));
	jor g3695(.dina(n3776),.dinb(w_n3528_0[0]),.dout(n3777),.clk(gclk));
	jand g3696(.dina(n3777),.dinb(n3688),.dout(n3778),.clk(gclk));
	jor g3697(.dina(n3778),.dinb(n3687),.dout(n3779),.clk(gclk));
	jor g3698(.dina(w_n3779_0[1]),.dinb(w_n3652_0[1]),.dout(n3780),.clk(gclk));
	jand g3699(.dina(n3780),.dinb(n3651),.dout(n3781),.clk(gclk));
	jand g3700(.dina(w_n3613_0[0]),.dinb(w_n3587_0[0]),.dout(n3782),.clk(gclk));
	jand g3701(.dina(w_n3614_0[0]),.dinb(w_n3532_0[0]),.dout(n3783),.clk(gclk));
	jor g3702(.dina(n3783),.dinb(n3782),.dout(n3784),.clk(gclk));
	jnot g3703(.din(w_n3604_0[0]),.dout(n3785),.clk(gclk));
	jand g3704(.dina(n3785),.dinb(w_n3590_0[0]),.dout(n3786),.clk(gclk));
	jor g3705(.dina(n3786),.dinb(w_n3602_0[0]),.dout(n3787),.clk(gclk));
	jand g3706(.dina(w_n3599_0[0]),.dinb(w_n3591_0[0]),.dout(n3788),.clk(gclk));
	jand g3707(.dina(w_n397_0[1]),.dinb(w_n243_1[1]),.dout(n3789),.clk(gclk));
	jand g3708(.dina(w_n679_0[2]),.dinb(w_n277_2[1]),.dout(n3790),.clk(gclk));
	jand g3709(.dina(n3790),.dinb(n3789),.dout(n3791),.clk(gclk));
	jand g3710(.dina(w_n2331_0[0]),.dinb(w_n869_0[0]),.dout(n3792),.clk(gclk));
	jand g3711(.dina(n3792),.dinb(w_n3624_0[1]),.dout(n3793),.clk(gclk));
	jand g3712(.dina(n3793),.dinb(n3791),.dout(n3794),.clk(gclk));
	jand g3713(.dina(w_n2511_0[2]),.dinb(w_n758_0[0]),.dout(n3795),.clk(gclk));
	jnot g3714(.din(w_n578_0[0]),.dout(n3796),.clk(gclk));
	jand g3715(.dina(w_n2339_0[0]),.dinb(n3796),.dout(n3797),.clk(gclk));
	jand g3716(.dina(n3797),.dinb(n3795),.dout(n3798),.clk(gclk));
	jand g3717(.dina(w_n825_0[2]),.dinb(w_n249_0[2]),.dout(n3799),.clk(gclk));
	jand g3718(.dina(n3799),.dinb(w_n421_1[2]),.dout(n3800),.clk(gclk));
	jand g3719(.dina(n3800),.dinb(w_n880_0[0]),.dout(n3801),.clk(gclk));
	jand g3720(.dina(n3801),.dinb(n3798),.dout(n3802),.clk(gclk));
	jand g3721(.dina(n3802),.dinb(w_n2743_0[0]),.dout(n3803),.clk(gclk));
	jand g3722(.dina(n3803),.dinb(w_n3794_0[1]),.dout(n3804),.clk(gclk));
	jand g3723(.dina(n3804),.dinb(w_n1319_0[0]),.dout(n3805),.clk(gclk));
	jxor g3724(.dina(w_n3805_0[1]),.dinb(n3788),.dout(n3806),.clk(gclk));
	jnot g3725(.din(w_n3806_5[2]),.dout(n3807),.clk(gclk));
	jand g3726(.dina(w_n3807_3[1]),.dinb(w_n3601_1[0]),.dout(n3808),.clk(gclk));
	jand g3727(.dina(w_n3805_0[0]),.dinb(w_n3600_8[0]),.dout(n3809),.clk(gclk));
	jor g3728(.dina(n3809),.dinb(w_n3808_0[1]),.dout(n3810),.clk(gclk));
	jxor g3729(.dina(w_n3810_0[1]),.dinb(w_n3787_0[1]),.dout(n3811),.clk(gclk));
	jor g3730(.dina(w_n3811_1[2]),.dinb(w_n3238_3[0]),.dout(n3812),.clk(gclk));
	jor g3731(.dina(w_n3806_5[1]),.dinb(w_n3322_2[2]),.dout(n3813),.clk(gclk));
	jor g3732(.dina(w_n3600_7[2]),.dinb(w_n3325_2[0]),.dout(n3814),.clk(gclk));
	jor g3733(.dina(w_n3328_2[1]),.dinb(w_n3315_6[1]),.dout(n3815),.clk(gclk));
	jand g3734(.dina(n3815),.dinb(n3814),.dout(n3816),.clk(gclk));
	jand g3735(.dina(n3816),.dinb(n3813),.dout(n3817),.clk(gclk));
	jand g3736(.dina(n3817),.dinb(n3812),.dout(n3818),.clk(gclk));
	jxor g3737(.dina(n3818),.dinb(w_n68_5[0]),.dout(n3819),.clk(gclk));
	jnot g3738(.din(n3819),.dout(n3820),.clk(gclk));
	jand g3739(.dina(w_n3585_0[0]),.dinb(w_n3543_0[0]),.dout(n3821),.clk(gclk));
	jand g3740(.dina(w_n3586_0[0]),.dinb(w_n3535_0[0]),.dout(n3822),.clk(gclk));
	jor g3741(.dina(n3822),.dinb(n3821),.dout(n3823),.clk(gclk));
	jand g3742(.dina(w_n3583_0[0]),.dinb(w_n3554_0[0]),.dout(n3824),.clk(gclk));
	jand g3743(.dina(w_n3584_0[0]),.dinb(w_n3546_0[0]),.dout(n3825),.clk(gclk));
	jor g3744(.dina(n3825),.dinb(n3824),.dout(n3826),.clk(gclk));
	jor g3745(.dina(w_n2795_4[1]),.dinb(w_n2771_1[0]),.dout(n3827),.clk(gclk));
	jor g3746(.dina(w_n2800_3[2]),.dinb(w_n2773_3[0]),.dout(n3828),.clk(gclk));
	jor g3747(.dina(w_n2805_3[2]),.dinb(w_n2669_2[0]),.dout(n3829),.clk(gclk));
	jor g3748(.dina(w_n2809_4[1]),.dinb(w_n2671_3[1]),.dout(n3830),.clk(gclk));
	jand g3749(.dina(n3830),.dinb(n3829),.dout(n3831),.clk(gclk));
	jand g3750(.dina(n3831),.dinb(n3828),.dout(n3832),.clk(gclk));
	jand g3751(.dina(n3832),.dinb(n3827),.dout(n3833),.clk(gclk));
	jxor g3752(.dina(n3833),.dinb(w_n699_6[2]),.dout(n3834),.clk(gclk));
	jnot g3753(.din(n3834),.dout(n3835),.clk(gclk));
	jand g3754(.dina(w_n3581_0[0]),.dinb(w_n3565_0[0]),.dout(n3836),.clk(gclk));
	jand g3755(.dina(w_n3582_0[0]),.dinb(w_n3557_0[0]),.dout(n3837),.clk(gclk));
	jor g3756(.dina(n3837),.dinb(n3836),.dout(n3838),.clk(gclk));
	jand g3757(.dina(w_n2694_1[1]),.dinb(w_n954_18[0]),.dout(n3839),.clk(gclk));
	jnot g3758(.din(n3839),.dout(n3840),.clk(gclk));
	jor g3759(.dina(w_n2911_0[1]),.dinb(w_n3198_5[0]),.dout(n3841),.clk(gclk));
	jand g3760(.dina(w_n2889_3[0]),.dinb(w_n2685_1[2]),.dout(n3842),.clk(gclk));
	jand g3761(.dina(w_n2887_3[1]),.dinb(w_n3571_1[0]),.dout(n3843),.clk(gclk));
	jand g3762(.dina(w_n2995_3[2]),.dinb(w_n3573_0[1]),.dout(n3844),.clk(gclk));
	jor g3763(.dina(n3844),.dinb(n3843),.dout(n3845),.clk(gclk));
	jor g3764(.dina(n3845),.dinb(n3842),.dout(n3846),.clk(gclk));
	jnot g3765(.din(n3846),.dout(n3847),.clk(gclk));
	jand g3766(.dina(n3847),.dinb(n3841),.dout(n3848),.clk(gclk));
	jxor g3767(.dina(w_n3848_0[1]),.dinb(n3840),.dout(n3849),.clk(gclk));
	jand g3768(.dina(w_n3580_0[0]),.dinb(w_n3567_0[0]),.dout(n3850),.clk(gclk));
	jand g3769(.dina(w_n2700_1[2]),.dinb(w_n954_17[2]),.dout(n3851),.clk(gclk));
	jand g3770(.dina(n3851),.dinb(w_n3579_0[0]),.dout(n3852),.clk(gclk));
	jor g3771(.dina(n3852),.dinb(n3850),.dout(n3853),.clk(gclk));
	jxor g3772(.dina(w_n3853_0[1]),.dinb(w_n3849_0[1]),.dout(n3854),.clk(gclk));
	jand g3773(.dina(w_n3004_0[2]),.dinb(w_n2828_1[2]),.dout(n3855),.clk(gclk));
	jand g3774(.dina(w_n2834_1[1]),.dinb(w_n2677_2[2]),.dout(n3856),.clk(gclk));
	jand g3775(.dina(w_n2848_1[2]),.dinb(w_n2684_2[2]),.dout(n3857),.clk(gclk));
	jand g3776(.dina(w_n2832_1[2]),.dinb(w_n2679_2[0]),.dout(n3858),.clk(gclk));
	jor g3777(.dina(n3858),.dinb(n3857),.dout(n3859),.clk(gclk));
	jor g3778(.dina(n3859),.dinb(n3856),.dout(n3860),.clk(gclk));
	jor g3779(.dina(n3860),.dinb(n3855),.dout(n3861),.clk(gclk));
	jxor g3780(.dina(n3861),.dinb(w_n803_4[0]),.dout(n3862),.clk(gclk));
	jxor g3781(.dina(w_n3862_0[1]),.dinb(w_n3854_0[1]),.dout(n3863),.clk(gclk));
	jxor g3782(.dina(w_n3863_0[1]),.dinb(w_n3838_0[1]),.dout(n3864),.clk(gclk));
	jxor g3783(.dina(w_n3864_0[1]),.dinb(w_n3835_0[1]),.dout(n3865),.clk(gclk));
	jxor g3784(.dina(w_n3865_0[1]),.dinb(w_n3826_0[1]),.dout(n3866),.clk(gclk));
	jor g3785(.dina(w_n3337_1[1]),.dinb(w_n79_3[2]),.dout(n3867),.clk(gclk));
	jor g3786(.dina(w_n3283_6[1]),.dinb(w_n2775_3[0]),.dout(n3868),.clk(gclk));
	jor g3787(.dina(w_n3284_6[1]),.dinb(w_n2780_3[0]),.dout(n3869),.clk(gclk));
	jor g3788(.dina(w_n3172_4[0]),.dinb(w_n2784_3[2]),.dout(n3870),.clk(gclk));
	jand g3789(.dina(n3870),.dinb(n3869),.dout(n3871),.clk(gclk));
	jand g3790(.dina(n3871),.dinb(n3868),.dout(n3872),.clk(gclk));
	jand g3791(.dina(n3872),.dinb(n3867),.dout(n3873),.clk(gclk));
	jxor g3792(.dina(n3873),.dinb(w_n56_5[2]),.dout(n3874),.clk(gclk));
	jxor g3793(.dina(w_n3874_0[1]),.dinb(w_n3866_0[1]),.dout(n3875),.clk(gclk));
	jxor g3794(.dina(w_n3875_0[1]),.dinb(w_n3823_0[1]),.dout(n3876),.clk(gclk));
	jxor g3795(.dina(w_n3876_0[1]),.dinb(w_n3820_0[1]),.dout(n3877),.clk(gclk));
	jxor g3796(.dina(w_n3877_0[1]),.dinb(w_n3784_0[1]),.dout(n3878),.clk(gclk));
	jand g3797(.dina(w_n3258_1[0]),.dinb(w_n1187_0[0]),.dout(n3879),.clk(gclk));
	jand g3798(.dina(n3879),.dinb(w_n1646_0[0]),.dout(n3880),.clk(gclk));
	jand g3799(.dina(w_n458_0[1]),.dinb(w_n264_1[0]),.dout(n3881),.clk(gclk));
	jand g3800(.dina(n3881),.dinb(w_n147_2[0]),.dout(n3882),.clk(gclk));
	jand g3801(.dina(w_n3624_0[0]),.dinb(w_n2360_0[0]),.dout(n3883),.clk(gclk));
	jand g3802(.dina(n3883),.dinb(n3882),.dout(n3884),.clk(gclk));
	jand g3803(.dina(n3884),.dinb(w_n1020_0[0]),.dout(n3885),.clk(gclk));
	jand g3804(.dina(n3885),.dinb(n3880),.dout(n3886),.clk(gclk));
	jand g3805(.dina(n3886),.dinb(w_n902_0[0]),.dout(n3887),.clk(gclk));
	jand g3806(.dina(n3887),.dinb(w_n2391_0[0]),.dout(n3888),.clk(gclk));
	jxor g3807(.dina(w_n3888_0[1]),.dinb(w_n3878_0[1]),.dout(n3889),.clk(gclk));
	jxor g3808(.dina(w_n3889_0[1]),.dinb(w_n3781_0[1]),.dout(n3890),.clk(gclk));
	jxor g3809(.dina(w_n3779_0[0]),.dinb(w_n3652_0[0]),.dout(n3891),.clk(gclk));
	jxor g3810(.dina(w_n3891_0[1]),.dinb(w_n3890_0[1]),.dout(sin0_fa_),.clk(gclk));
	jnot g3811(.din(w_n3878_0[0]),.dout(n3893),.clk(gclk));
	jor g3812(.dina(w_n3888_0[0]),.dinb(n3893),.dout(n3894),.clk(gclk));
	jor g3813(.dina(w_n3889_0[0]),.dinb(w_n3781_0[0]),.dout(n3895),.clk(gclk));
	jand g3814(.dina(n3895),.dinb(n3894),.dout(n3896),.clk(gclk));
	jand g3815(.dina(w_n3876_0[0]),.dinb(w_n3820_0[0]),.dout(n3897),.clk(gclk));
	jand g3816(.dina(w_n3877_0[0]),.dinb(w_n3784_0[0]),.dout(n3898),.clk(gclk));
	jor g3817(.dina(n3898),.dinb(n3897),.dout(n3899),.clk(gclk));
	jnot g3818(.din(w_n3810_0[0]),.dout(n3900),.clk(gclk));
	jand g3819(.dina(w_n3900_0[1]),.dinb(w_n3787_0[0]),.dout(n3901),.clk(gclk));
	jor g3820(.dina(n3901),.dinb(w_n3808_0[0]),.dout(n3902),.clk(gclk));
	jand g3821(.dina(w_n592_1[2]),.dinb(w_n454_0[2]),.dout(n3904),.clk(gclk));
	jand g3822(.dina(n3904),.dinb(w_n2326_0[0]),.dout(n3905),.clk(gclk));
	jand g3823(.dina(w_n2521_0[2]),.dinb(w_n417_0[2]),.dout(n3906),.clk(gclk));
	jand g3824(.dina(n3906),.dinb(w_n846_0[0]),.dout(n3907),.clk(gclk));
	jand g3825(.dina(n3907),.dinb(n3905),.dout(n3908),.clk(gclk));
	jand g3826(.dina(n3908),.dinb(w_n754_0[0]),.dout(n3909),.clk(gclk));
	jnot g3827(.din(w_n1679_0[0]),.dout(n3910),.clk(gclk));
	jand g3828(.dina(w_n3274_0[0]),.dinb(w_n493_0[0]),.dout(n3911),.clk(gclk));
	jand g3829(.dina(w_n463_1[1]),.dinb(w_n351_0[2]),.dout(n3912),.clk(gclk));
	jand g3830(.dina(n3912),.dinb(w_n2380_1[1]),.dout(n3913),.clk(gclk));
	jand g3831(.dina(n3913),.dinb(w_n855_0[0]),.dout(n3914),.clk(gclk));
	jand g3832(.dina(n3914),.dinb(w_n3911_0[1]),.dout(n3915),.clk(gclk));
	jand g3833(.dina(n3915),.dinb(n3910),.dout(n3916),.clk(gclk));
	jand g3834(.dina(n3916),.dinb(w_n933_0[0]),.dout(n3917),.clk(gclk));
	jand g3835(.dina(n3917),.dinb(w_n3909_0[1]),.dout(n3918),.clk(gclk));
	jand g3836(.dina(n3918),.dinb(w_n2520_0[1]),.dout(n3919),.clk(gclk));
	jnot g3837(.din(w_n3919_5[2]),.dout(n3920),.clk(gclk));
	jand g3838(.dina(w_n3919_5[1]),.dinb(w_n3807_3[0]),.dout(n3923),.clk(gclk));
	jand g3839(.dina(w_n3920_3[1]),.dinb(w_n3806_5[0]),.dout(n3924),.clk(gclk));
	jor g3840(.dina(w_n3924_0[1]),.dinb(n3923),.dout(n3925),.clk(gclk));
	jnot g3841(.din(w_n3925_0[1]),.dout(n3926),.clk(gclk));
	jxor g3842(.dina(n3926),.dinb(w_n3902_0[1]),.dout(n3927),.clk(gclk));
	jor g3843(.dina(w_n3927_1[2]),.dinb(w_n3238_2[2]),.dout(n3928),.clk(gclk));
	jor g3844(.dina(w_n3919_5[0]),.dinb(w_n3322_2[1]),.dout(n3929),.clk(gclk));
	jor g3845(.dina(w_n3806_4[2]),.dinb(w_n3325_1[2]),.dout(n3930),.clk(gclk));
	jor g3846(.dina(w_n3600_7[1]),.dinb(w_n3328_2[0]),.dout(n3931),.clk(gclk));
	jand g3847(.dina(n3931),.dinb(n3930),.dout(n3932),.clk(gclk));
	jand g3848(.dina(n3932),.dinb(n3929),.dout(n3933),.clk(gclk));
	jand g3849(.dina(n3933),.dinb(n3928),.dout(n3934),.clk(gclk));
	jxor g3850(.dina(n3934),.dinb(w_n68_4[2]),.dout(n3935),.clk(gclk));
	jnot g3851(.din(n3935),.dout(n3936),.clk(gclk));
	jand g3852(.dina(w_n3874_0[0]),.dinb(w_n3866_0[0]),.dout(n3937),.clk(gclk));
	jand g3853(.dina(w_n3875_0[0]),.dinb(w_n3823_0[0]),.dout(n3938),.clk(gclk));
	jor g3854(.dina(n3938),.dinb(n3937),.dout(n3939),.clk(gclk));
	jand g3855(.dina(w_n3864_0[0]),.dinb(w_n3835_0[0]),.dout(n3940),.clk(gclk));
	jand g3856(.dina(w_n3865_0[0]),.dinb(w_n3826_0[0]),.dout(n3941),.clk(gclk));
	jor g3857(.dina(n3941),.dinb(n3940),.dout(n3942),.clk(gclk));
	jand g3858(.dina(w_n3174_1[0]),.dinb(w_n2794_1[0]),.dout(n3943),.clk(gclk));
	jand g3859(.dina(w_n3176_1[2]),.dinb(w_n2799_0[2]),.dout(n3944),.clk(gclk));
	jand g3860(.dina(w_n2808_1[0]),.dinb(w_n2670_3[1]),.dout(n3945),.clk(gclk));
	jand g3861(.dina(w_n2804_1[0]),.dinb(w_n2769_2[1]),.dout(n3946),.clk(gclk));
	jor g3862(.dina(n3946),.dinb(n3945),.dout(n3947),.clk(gclk));
	jor g3863(.dina(n3947),.dinb(n3944),.dout(n3948),.clk(gclk));
	jor g3864(.dina(n3948),.dinb(n3943),.dout(n3949),.clk(gclk));
	jxor g3865(.dina(n3949),.dinb(w_n1143_4[1]),.dout(n3950),.clk(gclk));
	jnot g3866(.din(n3950),.dout(n3951),.clk(gclk));
	jand g3867(.dina(w_n3862_0[0]),.dinb(w_n3854_0[0]),.dout(n3952),.clk(gclk));
	jand g3868(.dina(w_n3863_0[0]),.dinb(w_n3838_0[0]),.dout(n3953),.clk(gclk));
	jor g3869(.dina(n3953),.dinb(n3952),.dout(n3954),.clk(gclk));
	jor g3870(.dina(w_n3028_0[2]),.dinb(w_n2857_4[2]),.dout(n3955),.clk(gclk));
	jor g3871(.dina(w_n2860_4[0]),.dinb(w_n2671_3[0]),.dout(n3956),.clk(gclk));
	jor g3872(.dina(w_n2865_4[0]),.dinb(w_n2674_1[2]),.dout(n3957),.clk(gclk));
	jor g3873(.dina(w_n2863_4[2]),.dinb(w_n2678_2[1]),.dout(n3958),.clk(gclk));
	jand g3874(.dina(n3958),.dinb(n3957),.dout(n3959),.clk(gclk));
	jand g3875(.dina(n3959),.dinb(n3956),.dout(n3960),.clk(gclk));
	jand g3876(.dina(n3960),.dinb(n3955),.dout(n3961),.clk(gclk));
	jxor g3877(.dina(n3961),.dinb(w_n808_7[1]),.dout(n3962),.clk(gclk));
	jand g3878(.dina(w_n2691_2[2]),.dinb(w_n954_17[1]),.dout(n3963),.clk(gclk));
	jnot g3879(.din(n3963),.dout(n3964),.clk(gclk));
	jor g3880(.dina(w_n2899_0[1]),.dinb(w_n3198_4[2]),.dout(n3965),.clk(gclk));
	jand g3881(.dina(w_n2889_2[2]),.dinb(w_n2684_2[1]),.dout(n3966),.clk(gclk));
	jand g3882(.dina(w_n2887_3[0]),.dinb(w_n2685_1[1]),.dout(n3967),.clk(gclk));
	jand g3883(.dina(w_n2995_3[1]),.dinb(w_n3571_0[2]),.dout(n3968),.clk(gclk));
	jor g3884(.dina(n3968),.dinb(n3967),.dout(n3969),.clk(gclk));
	jor g3885(.dina(n3969),.dinb(n3966),.dout(n3970),.clk(gclk));
	jnot g3886(.din(n3970),.dout(n3971),.clk(gclk));
	jand g3887(.dina(n3971),.dinb(n3965),.dout(n3972),.clk(gclk));
	jxor g3888(.dina(w_n3972_0[1]),.dinb(n3964),.dout(n3973),.clk(gclk));
	jand g3889(.dina(w_n3853_0[0]),.dinb(w_n3849_0[0]),.dout(n3974),.clk(gclk));
	jand g3890(.dina(w_n2693_1[1]),.dinb(w_n954_17[0]),.dout(n3975),.clk(gclk));
	jand g3891(.dina(n3975),.dinb(w_n3848_0[0]),.dout(n3976),.clk(gclk));
	jor g3892(.dina(n3976),.dinb(n3974),.dout(n3977),.clk(gclk));
	jxor g3893(.dina(w_n3977_0[1]),.dinb(w_n3973_0[1]),.dout(n3978),.clk(gclk));
	jxor g3894(.dina(w_n3978_0[1]),.dinb(w_n3962_0[1]),.dout(n3979),.clk(gclk));
	jxor g3895(.dina(w_n3979_0[1]),.dinb(w_n3954_0[1]),.dout(n3980),.clk(gclk));
	jxor g3896(.dina(w_n3980_0[1]),.dinb(w_n3951_0[1]),.dout(n3981),.clk(gclk));
	jxor g3897(.dina(w_n3981_0[1]),.dinb(w_n3942_0[1]),.dout(n3982),.clk(gclk));
	jor g3898(.dina(w_n3320_1[1]),.dinb(w_n79_3[1]),.dout(n3983),.clk(gclk));
	jor g3899(.dina(w_n3315_6[0]),.dinb(w_n2775_2[2]),.dout(n3984),.clk(gclk));
	jor g3900(.dina(w_n3283_6[0]),.dinb(w_n2780_2[2]),.dout(n3985),.clk(gclk));
	jor g3901(.dina(w_n3284_6[0]),.dinb(w_n2784_3[1]),.dout(n3986),.clk(gclk));
	jand g3902(.dina(n3986),.dinb(n3985),.dout(n3987),.clk(gclk));
	jand g3903(.dina(n3987),.dinb(n3984),.dout(n3988),.clk(gclk));
	jand g3904(.dina(n3988),.dinb(n3983),.dout(n3989),.clk(gclk));
	jxor g3905(.dina(n3989),.dinb(w_n56_5[1]),.dout(n3990),.clk(gclk));
	jxor g3906(.dina(w_n3990_0[1]),.dinb(w_n3982_0[1]),.dout(n3991),.clk(gclk));
	jxor g3907(.dina(w_n3991_0[1]),.dinb(w_n3939_0[1]),.dout(n3992),.clk(gclk));
	jxor g3908(.dina(w_n3992_0[1]),.dinb(w_n3936_0[1]),.dout(n3993),.clk(gclk));
	jxor g3909(.dina(w_n3993_0[1]),.dinb(w_n3899_0[1]),.dout(n3994),.clk(gclk));
	jand g3910(.dina(w_n1018_0[1]),.dinb(w_n417_0[1]),.dout(n3995),.clk(gclk));
	jand g3911(.dina(w_n2457_0[0]),.dinb(w_n2429_1[0]),.dout(n3996),.clk(gclk));
	jand g3912(.dina(n3996),.dinb(n3995),.dout(n3997),.clk(gclk));
	jnot g3913(.din(w_n1658_0[0]),.dout(n3998),.clk(gclk));
	jand g3914(.dina(w_n1209_0[2]),.dinb(w_n241_0[1]),.dout(n3999),.clk(gclk));
	jand g3915(.dina(n3999),.dinb(n3998),.dout(n4000),.clk(gclk));
	jand g3916(.dina(w_n592_1[1]),.dinb(w_n430_0[2]),.dout(n4001),.clk(gclk));
	jand g3917(.dina(w_n632_1[0]),.dinb(w_n321_0[1]),.dout(n4002),.clk(gclk));
	jand g3918(.dina(n4002),.dinb(n4001),.dout(n4003),.clk(gclk));
	jand g3919(.dina(n4003),.dinb(w_n4000_0[2]),.dout(n4004),.clk(gclk));
	jand g3920(.dina(w_n3258_0[2]),.dinb(w_n3242_0[1]),.dout(n4005),.clk(gclk));
	jand g3921(.dina(n4005),.dinb(n4004),.dout(n4006),.clk(gclk));
	jand g3922(.dina(n4006),.dinb(n3997),.dout(n4007),.clk(gclk));
	jand g3923(.dina(n4007),.dinb(w_n3630_0[0]),.dout(n4008),.clk(gclk));
	jand g3924(.dina(n4008),.dinb(w_n2359_0[0]),.dout(n4009),.clk(gclk));
	jxor g3925(.dina(w_n4009_0[1]),.dinb(w_n3994_0[1]),.dout(n4010),.clk(gclk));
	jxor g3926(.dina(w_n4010_0[1]),.dinb(w_n3896_0[1]),.dout(n4011),.clk(gclk));
	jnot g3927(.din(w_n4011_0[2]),.dout(n4012),.clk(gclk));
	jxor g3928(.dina(a23),.dinb(w_a22_2[0]),.dout(n4013),.clk(gclk));
	jand g3929(.dina(w_n4013_10[2]),.dinb(w_sin0_0[1]),.dout(n4014),.clk(gclk));
	jand g3930(.dina(w_n4014_0[1]),.dinb(n4012),.dout(n4015),.clk(gclk));
	jnot g3931(.din(w_n4014_0[0]),.dout(n4016),.clk(gclk));
	jand g3932(.dina(w_n3891_0[0]),.dinb(w_n3890_0[0]),.dout(n4017),.clk(gclk));
	jxor g3933(.dina(w_n4011_0[1]),.dinb(w_n4017_0[1]),.dout(n4018),.clk(gclk));
	jand g3934(.dina(w_n4018_0[1]),.dinb(n4016),.dout(n4019),.clk(gclk));
	jor g3935(.dina(n4019),.dinb(n4015),.dout(w_dff_A_lIGy9qnK1_2),.clk(gclk));
	jand g3936(.dina(w_n4011_0[0]),.dinb(w_n4017_0[0]),.dout(n4021),.clk(gclk));
	jnot g3937(.din(w_n3994_0[0]),.dout(n4022),.clk(gclk));
	jor g3938(.dina(w_n4009_0[0]),.dinb(n4022),.dout(n4023),.clk(gclk));
	jor g3939(.dina(w_n4010_0[0]),.dinb(w_n3896_0[0]),.dout(n4024),.clk(gclk));
	jand g3940(.dina(n4024),.dinb(n4023),.dout(n4025),.clk(gclk));
	jand g3941(.dina(w_n3992_0[0]),.dinb(w_n3936_0[0]),.dout(n4026),.clk(gclk));
	jand g3942(.dina(w_n3993_0[0]),.dinb(w_n3899_0[0]),.dout(n4027),.clk(gclk));
	jor g3943(.dina(n4027),.dinb(n4026),.dout(n4028),.clk(gclk));
	jand g3944(.dina(w_n3990_0[0]),.dinb(w_n3982_0[0]),.dout(n4029),.clk(gclk));
	jand g3945(.dina(w_n3991_0[0]),.dinb(w_n3939_0[0]),.dout(n4030),.clk(gclk));
	jor g3946(.dina(n4030),.dinb(n4029),.dout(n4031),.clk(gclk));
	jand g3947(.dina(w_n3980_0[0]),.dinb(w_n3951_0[0]),.dout(n4032),.clk(gclk));
	jand g3948(.dina(w_n3981_0[0]),.dinb(w_n3942_0[0]),.dout(n4033),.clk(gclk));
	jor g3949(.dina(n4033),.dinb(n4032),.dout(n4034),.clk(gclk));
	jor g3950(.dina(w_n3516_1[0]),.dinb(w_n2795_4[0]),.dout(n4035),.clk(gclk));
	jor g3951(.dina(w_n3284_5[2]),.dinb(w_n2800_3[1]),.dout(n4036),.clk(gclk));
	jor g3952(.dina(w_n3172_3[2]),.dinb(w_n2805_3[1]),.dout(n4037),.clk(gclk));
	jor g3953(.dina(w_n2809_4[0]),.dinb(w_n2773_2[2]),.dout(n4038),.clk(gclk));
	jand g3954(.dina(n4038),.dinb(n4037),.dout(n4039),.clk(gclk));
	jand g3955(.dina(n4039),.dinb(n4036),.dout(n4040),.clk(gclk));
	jand g3956(.dina(n4040),.dinb(n4035),.dout(n4041),.clk(gclk));
	jxor g3957(.dina(n4041),.dinb(w_n699_6[1]),.dout(n4042),.clk(gclk));
	jnot g3958(.din(n4042),.dout(n4043),.clk(gclk));
	jand g3959(.dina(w_n3978_0[0]),.dinb(w_n3962_0[0]),.dout(n4044),.clk(gclk));
	jand g3960(.dina(w_n3979_0[0]),.dinb(w_n3954_0[0]),.dout(n4045),.clk(gclk));
	jor g3961(.dina(n4045),.dinb(n4044),.dout(n4046),.clk(gclk));
	jand g3962(.dina(w_n3016_0[2]),.dinb(w_n2828_1[1]),.dout(n4047),.clk(gclk));
	jand g3963(.dina(w_n2834_1[0]),.dinb(w_n2670_3[0]),.dout(n4048),.clk(gclk));
	jand g3964(.dina(w_n2848_1[1]),.dinb(w_n2677_2[1]),.dout(n4049),.clk(gclk));
	jand g3965(.dina(w_n2832_1[1]),.dinb(w_n2672_1[1]),.dout(n4050),.clk(gclk));
	jor g3966(.dina(n4050),.dinb(n4049),.dout(n4051),.clk(gclk));
	jor g3967(.dina(n4051),.dinb(n4048),.dout(n4052),.clk(gclk));
	jor g3968(.dina(n4052),.dinb(n4047),.dout(n4053),.clk(gclk));
	jxor g3969(.dina(n4053),.dinb(w_n803_3[2]),.dout(n4054),.clk(gclk));
	jand g3970(.dina(w_n2688_2[2]),.dinb(w_n954_16[2]),.dout(n4055),.clk(gclk));
	jnot g3971(.din(n4055),.dout(n4056),.clk(gclk));
	jor g3972(.dina(w_n3198_4[1]),.dinb(w_n2797_0[1]),.dout(n4057),.clk(gclk));
	jand g3973(.dina(w_n2889_2[1]),.dinb(w_n2679_1[2]),.dout(n4058),.clk(gclk));
	jand g3974(.dina(w_n2887_2[2]),.dinb(w_n2684_2[0]),.dout(n4059),.clk(gclk));
	jand g3975(.dina(w_n2995_3[0]),.dinb(w_n2685_1[0]),.dout(n4060),.clk(gclk));
	jor g3976(.dina(n4060),.dinb(n4059),.dout(n4061),.clk(gclk));
	jor g3977(.dina(n4061),.dinb(n4058),.dout(n4062),.clk(gclk));
	jnot g3978(.din(n4062),.dout(n4063),.clk(gclk));
	jand g3979(.dina(n4063),.dinb(n4057),.dout(n4064),.clk(gclk));
	jxor g3980(.dina(w_n4064_0[1]),.dinb(n4056),.dout(n4065),.clk(gclk));
	jand g3981(.dina(w_n3977_0[0]),.dinb(w_n3973_0[0]),.dout(n4066),.clk(gclk));
	jand g3982(.dina(w_n3573_0[0]),.dinb(w_n954_16[1]),.dout(n4067),.clk(gclk));
	jand g3983(.dina(n4067),.dinb(w_n3972_0[0]),.dout(n4068),.clk(gclk));
	jor g3984(.dina(n4068),.dinb(n4066),.dout(n4069),.clk(gclk));
	jxor g3985(.dina(w_n4069_0[1]),.dinb(w_n4065_0[1]),.dout(n4070),.clk(gclk));
	jxor g3986(.dina(w_n4070_0[1]),.dinb(w_n4054_0[1]),.dout(n4071),.clk(gclk));
	jxor g3987(.dina(w_n4071_0[1]),.dinb(w_n4046_0[1]),.dout(n4072),.clk(gclk));
	jxor g3988(.dina(w_n4072_0[1]),.dinb(w_n4043_0[1]),.dout(n4073),.clk(gclk));
	jxor g3989(.dina(w_n4073_0[1]),.dinb(w_n4034_0[1]),.dout(n4074),.clk(gclk));
	jor g3990(.dina(w_n3605_1[1]),.dinb(w_n79_3[0]),.dout(n4075),.clk(gclk));
	jor g3991(.dina(w_n3600_7[0]),.dinb(w_n2775_2[1]),.dout(n4076),.clk(gclk));
	jor g3992(.dina(w_n3315_5[2]),.dinb(w_n2780_2[1]),.dout(n4077),.clk(gclk));
	jor g3993(.dina(w_n3283_5[2]),.dinb(w_n2784_3[0]),.dout(n4078),.clk(gclk));
	jand g3994(.dina(n4078),.dinb(n4077),.dout(n4079),.clk(gclk));
	jand g3995(.dina(n4079),.dinb(n4076),.dout(n4080),.clk(gclk));
	jand g3996(.dina(n4080),.dinb(n4075),.dout(n4081),.clk(gclk));
	jxor g3997(.dina(n4081),.dinb(w_n56_5[0]),.dout(n4082),.clk(gclk));
	jxor g3998(.dina(w_n4082_0[1]),.dinb(w_n4074_0[1]),.dout(n4083),.clk(gclk));
	jxor g3999(.dina(w_n4083_0[1]),.dinb(w_n4031_0[1]),.dout(n4084),.clk(gclk));
	jand g4000(.dina(w_n3920_3[0]),.dinb(w_n3324_0[2]),.dout(n4085),.clk(gclk));
	jand g4001(.dina(w_n3925_0[0]),.dinb(w_n3902_0[0]),.dout(n4086),.clk(gclk));
	jand g4002(.dina(w_n4086_0[1]),.dinb(w_n3919_4[2]),.dout(n4087),.clk(gclk));
	jnot g4003(.din(w_n4086_0[0]),.dout(n4088),.clk(gclk));
	jand g4004(.dina(w_n4088_0[1]),.dinb(w_n3924_0[0]),.dout(n4089),.clk(gclk));
	jor g4005(.dina(n4089),.dinb(n4087),.dout(n4090),.clk(gclk));
	jand g4006(.dina(w_n4090_1[2]),.dinb(w_n3237_0[2]),.dout(n4091),.clk(gclk));
	jor g4007(.dina(n4091),.dinb(n4085),.dout(n4092),.clk(gclk));
	jand g4008(.dina(w_n3807_2[2]),.dinb(w_n63_0[2]),.dout(n4093),.clk(gclk));
	jor g4009(.dina(n4093),.dinb(w_n3233_3[2]),.dout(n4094),.clk(gclk));
	jnot g4010(.din(n4094),.dout(n4095),.clk(gclk));
	jor g4011(.dina(n4095),.dinb(w_n4092_0[1]),.dout(n4096),.clk(gclk));
	jnot g4012(.din(w_n4092_0[0]),.dout(n4097),.clk(gclk));
	jor g4013(.dina(n4097),.dinb(w_n3233_3[1]),.dout(n4098),.clk(gclk));
	jand g4014(.dina(n4098),.dinb(n4096),.dout(n4099),.clk(gclk));
	jxor g4015(.dina(w_n4099_0[1]),.dinb(w_n4084_0[1]),.dout(n4100),.clk(gclk));
	jxor g4016(.dina(w_n4100_0[1]),.dinb(w_n4028_0[1]),.dout(n4101),.clk(gclk));
	jand g4017(.dina(w_n294_1[0]),.dinb(w_n229_1[0]),.dout(n4102),.clk(gclk));
	jand g4018(.dina(n4102),.dinb(w_n825_0[1]),.dout(n4103),.clk(gclk));
	jand g4019(.dina(w_n412_0[2]),.dinb(w_n270_1[0]),.dout(n4104),.clk(gclk));
	jand g4020(.dina(n4104),.dinb(w_n2734_0[1]),.dout(n4105),.clk(gclk));
	jand g4021(.dina(n4105),.dinb(n4103),.dout(n4106),.clk(gclk));
	jand g4022(.dina(w_n744_0[2]),.dinb(w_n282_1[0]),.dout(n4107),.clk(gclk));
	jand g4023(.dina(n4107),.dinb(w_n265_0[0]),.dout(n4108),.clk(gclk));
	jand g4024(.dina(n4108),.dinb(w_n988_0[0]),.dout(n4109),.clk(gclk));
	jand g4025(.dina(w_n2380_1[0]),.dinb(w_n732_1[0]),.dout(n4110),.clk(gclk));
	jand g4026(.dina(n4110),.dinb(w_n374_0[2]),.dout(n4111),.clk(gclk));
	jand g4027(.dina(n4111),.dinb(w_n999_0[1]),.dout(n4112),.clk(gclk));
	jand g4028(.dina(n4112),.dinb(n4109),.dout(n4113),.clk(gclk));
	jand g4029(.dina(n4113),.dinb(w_n4106_0[1]),.dout(n4114),.clk(gclk));
	jand g4030(.dina(n4114),.dinb(w_n923_0[0]),.dout(n4115),.clk(gclk));
	jand g4031(.dina(n4115),.dinb(w_n3693_0[1]),.dout(n4116),.clk(gclk));
	jxor g4032(.dina(w_n4116_0[1]),.dinb(w_n4101_0[1]),.dout(n4117),.clk(gclk));
	jxor g4033(.dina(w_n4117_0[1]),.dinb(w_n4025_0[1]),.dout(n4118),.clk(gclk));
	jxor g4034(.dina(w_n4118_0[1]),.dinb(w_n4021_0[1]),.dout(n4119),.clk(gclk));
	jor g4035(.dina(w_n4018_0[0]),.dinb(w_sin0_0[0]),.dout(n4120),.clk(gclk));
	jand g4036(.dina(w_n4120_0[1]),.dinb(w_n4013_10[1]),.dout(n4121),.clk(gclk));
	jxor g4037(.dina(n4121),.dinb(w_n4119_0[1]),.dout(w_dff_A_QWIijunn1_2),.clk(gclk));
	jor g4038(.dina(w_n4120_0[0]),.dinb(w_n4119_0[0]),.dout(n4123),.clk(gclk));
	jand g4039(.dina(w_n4123_0[1]),.dinb(w_n4013_10[0]),.dout(n4124),.clk(gclk));
	jand g4040(.dina(w_n4118_0[0]),.dinb(w_n4021_0[0]),.dout(n4125),.clk(gclk));
	jnot g4041(.din(w_n4101_0[0]),.dout(n4126),.clk(gclk));
	jor g4042(.dina(w_n4116_0[0]),.dinb(n4126),.dout(n4127),.clk(gclk));
	jor g4043(.dina(w_n4117_0[0]),.dinb(w_n4025_0[0]),.dout(n4128),.clk(gclk));
	jand g4044(.dina(n4128),.dinb(n4127),.dout(n4129),.clk(gclk));
	jand g4045(.dina(w_n4099_0[0]),.dinb(w_n4084_0[0]),.dout(n4130),.clk(gclk));
	jand g4046(.dina(w_n4100_0[0]),.dinb(w_n4028_0[0]),.dout(n4131),.clk(gclk));
	jor g4047(.dina(n4131),.dinb(n4130),.dout(n4132),.clk(gclk));
	jand g4048(.dina(w_n4082_0[0]),.dinb(w_n4074_0[0]),.dout(n4133),.clk(gclk));
	jand g4049(.dina(w_n4083_0[0]),.dinb(w_n4031_0[0]),.dout(n4134),.clk(gclk));
	jor g4050(.dina(n4134),.dinb(n4133),.dout(n4135),.clk(gclk));
	jand g4051(.dina(w_n4088_0[0]),.dinb(w_n3806_4[1]),.dout(n4136),.clk(gclk));
	jor g4052(.dina(w_n4136_1[2]),.dinb(w_n3238_2[1]),.dout(n4137),.clk(gclk));
	jand g4053(.dina(n4137),.dinb(w_n3328_1[2]),.dout(n4138),.clk(gclk));
	jor g4054(.dina(n4138),.dinb(w_n3919_4[1]),.dout(n4139),.clk(gclk));
	jxor g4055(.dina(n4139),.dinb(w_n68_4[1]),.dout(n4140),.clk(gclk));
	jnot g4056(.din(n4140),.dout(n4141),.clk(gclk));
	jand g4057(.dina(w_n4072_0[0]),.dinb(w_n4043_0[0]),.dout(n4142),.clk(gclk));
	jand g4058(.dina(w_n4073_0[0]),.dinb(w_n4034_0[0]),.dout(n4143),.clk(gclk));
	jor g4059(.dina(n4143),.dinb(n4142),.dout(n4144),.clk(gclk));
	jor g4060(.dina(w_n3337_1[0]),.dinb(w_n2795_3[2]),.dout(n4145),.clk(gclk));
	jor g4061(.dina(w_n3283_5[1]),.dinb(w_n2800_3[0]),.dout(n4146),.clk(gclk));
	jor g4062(.dina(w_n3284_5[1]),.dinb(w_n2805_3[0]),.dout(n4147),.clk(gclk));
	jor g4063(.dina(w_n3172_3[1]),.dinb(w_n2809_3[2]),.dout(n4148),.clk(gclk));
	jand g4064(.dina(n4148),.dinb(n4147),.dout(n4149),.clk(gclk));
	jand g4065(.dina(n4149),.dinb(n4146),.dout(n4150),.clk(gclk));
	jand g4066(.dina(n4150),.dinb(n4145),.dout(n4151),.clk(gclk));
	jxor g4067(.dina(n4151),.dinb(w_n699_6[0]),.dout(n4152),.clk(gclk));
	jnot g4068(.din(n4152),.dout(n4153),.clk(gclk));
	jand g4069(.dina(w_n4070_0[0]),.dinb(w_n4054_0[0]),.dout(n4154),.clk(gclk));
	jand g4070(.dina(w_n4071_0[0]),.dinb(w_n4046_0[0]),.dout(n4155),.clk(gclk));
	jor g4071(.dina(n4155),.dinb(n4154),.dout(n4156),.clk(gclk));
	jor g4072(.dina(w_n2857_4[1]),.dinb(w_n2771_0[2]),.dout(n4157),.clk(gclk));
	jor g4073(.dina(w_n2860_3[2]),.dinb(w_n2773_2[1]),.dout(n4158),.clk(gclk));
	jor g4074(.dina(w_n2865_3[2]),.dinb(w_n2669_1[2]),.dout(n4159),.clk(gclk));
	jor g4075(.dina(w_n2863_4[1]),.dinb(w_n2671_2[2]),.dout(n4160),.clk(gclk));
	jand g4076(.dina(n4160),.dinb(n4159),.dout(n4161),.clk(gclk));
	jand g4077(.dina(n4161),.dinb(n4158),.dout(n4162),.clk(gclk));
	jand g4078(.dina(n4162),.dinb(n4157),.dout(n4163),.clk(gclk));
	jxor g4079(.dina(n4163),.dinb(w_n808_7[0]),.dout(n4164),.clk(gclk));
	jand g4080(.dina(w_n2687_2[1]),.dinb(w_n954_16[0]),.dout(n4165),.clk(gclk));
	jand g4081(.dina(w_n3004_0[1]),.dinb(w_n2883_2[1]),.dout(n4166),.clk(gclk));
	jand g4082(.dina(w_n2889_2[0]),.dinb(w_n2677_2[0]),.dout(n4167),.clk(gclk));
	jand g4083(.dina(w_n2995_2[2]),.dinb(w_n2684_1[2]),.dout(n4168),.clk(gclk));
	jand g4084(.dina(w_n2887_2[1]),.dinb(w_n2679_1[1]),.dout(n4169),.clk(gclk));
	jor g4085(.dina(n4169),.dinb(n4168),.dout(n4170),.clk(gclk));
	jor g4086(.dina(n4170),.dinb(n4167),.dout(n4171),.clk(gclk));
	jor g4087(.dina(n4171),.dinb(n4166),.dout(n4172),.clk(gclk));
	jxor g4088(.dina(w_n4172_0[1]),.dinb(n4165),.dout(n4173),.clk(gclk));
	jand g4089(.dina(w_n4069_0[0]),.dinb(w_n4065_0[0]),.dout(n4174),.clk(gclk));
	jand g4090(.dina(w_n3571_0[1]),.dinb(w_n954_15[2]),.dout(n4175),.clk(gclk));
	jand g4091(.dina(n4175),.dinb(w_n4064_0[0]),.dout(n4176),.clk(gclk));
	jor g4092(.dina(n4176),.dinb(n4174),.dout(n4177),.clk(gclk));
	jxor g4093(.dina(w_n4177_0[1]),.dinb(w_n4173_0[1]),.dout(n4178),.clk(gclk));
	jxor g4094(.dina(w_n4178_0[1]),.dinb(w_n4164_0[1]),.dout(n4179),.clk(gclk));
	jxor g4095(.dina(w_n4179_0[1]),.dinb(w_n4156_0[1]),.dout(n4180),.clk(gclk));
	jxor g4096(.dina(w_n4180_0[1]),.dinb(w_n4153_0[1]),.dout(n4181),.clk(gclk));
	jxor g4097(.dina(w_n4181_0[1]),.dinb(w_n4144_0[1]),.dout(n4182),.clk(gclk));
	jor g4098(.dina(w_n3811_1[1]),.dinb(w_n79_2[2]),.dout(n4183),.clk(gclk));
	jor g4099(.dina(w_n3806_4[0]),.dinb(w_n2775_2[0]),.dout(n4184),.clk(gclk));
	jor g4100(.dina(w_n3600_6[2]),.dinb(w_n2780_2[0]),.dout(n4185),.clk(gclk));
	jor g4101(.dina(w_n3315_5[1]),.dinb(w_n2784_2[2]),.dout(n4186),.clk(gclk));
	jand g4102(.dina(n4186),.dinb(n4185),.dout(n4187),.clk(gclk));
	jand g4103(.dina(n4187),.dinb(n4184),.dout(n4188),.clk(gclk));
	jand g4104(.dina(n4188),.dinb(n4183),.dout(n4189),.clk(gclk));
	jxor g4105(.dina(n4189),.dinb(w_n56_4[2]),.dout(n4190),.clk(gclk));
	jxor g4106(.dina(w_n4190_0[1]),.dinb(w_n4182_0[1]),.dout(n4191),.clk(gclk));
	jxor g4107(.dina(w_n4191_0[1]),.dinb(w_n4141_0[1]),.dout(n4192),.clk(gclk));
	jxor g4108(.dina(w_n4192_0[1]),.dinb(w_n4135_0[1]),.dout(n4193),.clk(gclk));
	jxor g4109(.dina(w_n4193_0[1]),.dinb(w_n4132_0[1]),.dout(n4194),.clk(gclk));
	jand g4110(.dina(w_n3669_0[0]),.dinb(w_n466_0[0]),.dout(n4195),.clk(gclk));
	jand g4111(.dina(n4195),.dinb(w_n881_0[1]),.dout(n4196),.clk(gclk));
	jand g4112(.dina(w_n2429_0[2]),.dinb(w_n2305_0[0]),.dout(n4197),.clk(gclk));
	jand g4113(.dina(n4197),.dinb(w_n280_0[1]),.dout(n4198),.clk(gclk));
	jand g4114(.dina(w_n925_0[1]),.dinb(w_n918_1[0]),.dout(n4199),.clk(gclk));
	jand g4115(.dina(w_n632_0[2]),.dinb(w_n488_0[2]),.dout(n4200),.clk(gclk));
	jand g4116(.dina(n4200),.dinb(n4199),.dout(n4201),.clk(gclk));
	jand g4117(.dina(n4201),.dinb(w_n565_0[2]),.dout(n4202),.clk(gclk));
	jand g4118(.dina(n4202),.dinb(n4198),.dout(n4203),.clk(gclk));
	jand g4119(.dina(n4203),.dinb(w_n2365_0[0]),.dout(n4204),.clk(gclk));
	jand g4120(.dina(n4204),.dinb(n4196),.dout(n4205),.clk(gclk));
	jand g4121(.dina(n4205),.dinb(w_n3155_0[0]),.dout(n4206),.clk(gclk));
	jxor g4122(.dina(w_n4206_0[1]),.dinb(w_n4194_0[1]),.dout(n4207),.clk(gclk));
	jxor g4123(.dina(w_n4207_0[1]),.dinb(w_n4129_0[1]),.dout(n4208),.clk(gclk));
	jxor g4124(.dina(w_n4208_0[1]),.dinb(w_n4125_0[1]),.dout(n4209),.clk(gclk));
	jxor g4125(.dina(w_n4209_0[1]),.dinb(n4124),.dout(w_dff_A_oRAz1Nyn2_2),.clk(gclk));
	jand g4126(.dina(w_n4208_0[0]),.dinb(w_n4125_0[0]),.dout(n4211),.clk(gclk));
	jnot g4127(.din(w_n4194_0[0]),.dout(n4212),.clk(gclk));
	jor g4128(.dina(w_n4206_0[0]),.dinb(n4212),.dout(n4213),.clk(gclk));
	jor g4129(.dina(w_n4207_0[0]),.dinb(w_n4129_0[0]),.dout(n4214),.clk(gclk));
	jand g4130(.dina(n4214),.dinb(n4213),.dout(n4215),.clk(gclk));
	jand g4131(.dina(w_n4192_0[0]),.dinb(w_n4135_0[0]),.dout(n4216),.clk(gclk));
	jand g4132(.dina(w_n4193_0[0]),.dinb(w_n4132_0[0]),.dout(n4217),.clk(gclk));
	jor g4133(.dina(n4217),.dinb(n4216),.dout(n4218),.clk(gclk));
	jand g4134(.dina(w_n4190_0[0]),.dinb(w_n4182_0[0]),.dout(n4219),.clk(gclk));
	jand g4135(.dina(w_n4191_0[0]),.dinb(w_n4141_0[0]),.dout(n4220),.clk(gclk));
	jor g4136(.dina(n4220),.dinb(n4219),.dout(n4221),.clk(gclk));
	jand g4137(.dina(w_n4180_0[0]),.dinb(w_n4153_0[0]),.dout(n4222),.clk(gclk));
	jand g4138(.dina(w_n4181_0[0]),.dinb(w_n4144_0[0]),.dout(n4223),.clk(gclk));
	jor g4139(.dina(n4223),.dinb(n4222),.dout(n4224),.clk(gclk));
	jor g4140(.dina(w_n3320_1[0]),.dinb(w_n2795_3[1]),.dout(n4225),.clk(gclk));
	jor g4141(.dina(w_n3315_5[0]),.dinb(w_n2800_2[2]),.dout(n4226),.clk(gclk));
	jor g4142(.dina(w_n3283_5[0]),.dinb(w_n2805_2[2]),.dout(n4227),.clk(gclk));
	jor g4143(.dina(w_n3284_5[0]),.dinb(w_n2809_3[1]),.dout(n4228),.clk(gclk));
	jand g4144(.dina(n4228),.dinb(n4227),.dout(n4229),.clk(gclk));
	jand g4145(.dina(n4229),.dinb(n4226),.dout(n4230),.clk(gclk));
	jand g4146(.dina(n4230),.dinb(n4225),.dout(n4231),.clk(gclk));
	jxor g4147(.dina(n4231),.dinb(w_n699_5[2]),.dout(n4232),.clk(gclk));
	jnot g4148(.din(n4232),.dout(n4233),.clk(gclk));
	jand g4149(.dina(w_n4178_0[0]),.dinb(w_n4164_0[0]),.dout(n4234),.clk(gclk));
	jand g4150(.dina(w_n4179_0[0]),.dinb(w_n4156_0[0]),.dout(n4235),.clk(gclk));
	jor g4151(.dina(n4235),.dinb(n4234),.dout(n4236),.clk(gclk));
	jor g4152(.dina(w_n3028_0[1]),.dinb(w_n3198_4[0]),.dout(n4237),.clk(gclk));
	jor g4153(.dina(w_n3200_3[1]),.dinb(w_n2671_2[1]),.dout(n4238),.clk(gclk));
	jor g4154(.dina(w_n3204_3[1]),.dinb(w_n2674_1[1]),.dout(n4239),.clk(gclk));
	jor g4155(.dina(w_n3202_3[1]),.dinb(w_n2678_2[0]),.dout(n4240),.clk(gclk));
	jand g4156(.dina(n4240),.dinb(n4239),.dout(n4241),.clk(gclk));
	jand g4157(.dina(n4241),.dinb(n4238),.dout(n4242),.clk(gclk));
	jand g4158(.dina(n4242),.dinb(n4237),.dout(n4243),.clk(gclk));
	jxor g4159(.dina(n4243),.dinb(w_n954_15[1]),.dout(n4244),.clk(gclk));
	jnot g4160(.din(n4244),.dout(n4245),.clk(gclk));
	jand g4161(.dina(w_n2684_1[1]),.dinb(w_n954_15[0]),.dout(n4246),.clk(gclk));
	jxor g4162(.dina(w_n4246_0[1]),.dinb(w_n68_4[0]),.dout(n4247),.clk(gclk));
	jxor g4163(.dina(w_n4247_0[1]),.dinb(w_n4245_0[1]),.dout(n4248),.clk(gclk));
	jand g4164(.dina(w_n4177_0[0]),.dinb(w_n4173_0[0]),.dout(n4249),.clk(gclk));
	jnot g4165(.din(w_n4172_0[0]),.dout(n4250),.clk(gclk));
	jand g4166(.dina(w_n2685_0[2]),.dinb(w_n954_14[2]),.dout(n4251),.clk(gclk));
	jand g4167(.dina(n4251),.dinb(n4250),.dout(n4252),.clk(gclk));
	jor g4168(.dina(n4252),.dinb(n4249),.dout(n4253),.clk(gclk));
	jxor g4169(.dina(w_n4253_0[1]),.dinb(w_n4248_0[1]),.dout(n4254),.clk(gclk));
	jand g4170(.dina(w_n3174_0[2]),.dinb(w_n2828_1[0]),.dout(n4255),.clk(gclk));
	jand g4171(.dina(w_n3176_1[1]),.dinb(w_n2834_0[2]),.dout(n4256),.clk(gclk));
	jand g4172(.dina(w_n2848_1[0]),.dinb(w_n2670_2[2]),.dout(n4257),.clk(gclk));
	jand g4173(.dina(w_n2832_1[0]),.dinb(w_n2769_2[0]),.dout(n4258),.clk(gclk));
	jor g4174(.dina(n4258),.dinb(n4257),.dout(n4259),.clk(gclk));
	jor g4175(.dina(n4259),.dinb(n4256),.dout(n4260),.clk(gclk));
	jor g4176(.dina(n4260),.dinb(n4255),.dout(n4261),.clk(gclk));
	jxor g4177(.dina(n4261),.dinb(w_n803_3[1]),.dout(n4262),.clk(gclk));
	jxor g4178(.dina(w_n4262_0[1]),.dinb(w_n4254_0[1]),.dout(n4263),.clk(gclk));
	jxor g4179(.dina(w_n4263_0[1]),.dinb(w_n4236_0[1]),.dout(n4264),.clk(gclk));
	jxor g4180(.dina(w_n4264_0[1]),.dinb(w_n4233_0[1]),.dout(n4265),.clk(gclk));
	jxor g4181(.dina(w_n4265_0[1]),.dinb(w_n4224_0[1]),.dout(n4266),.clk(gclk));
	jor g4182(.dina(w_n3927_1[1]),.dinb(w_n79_2[1]),.dout(n4267),.clk(gclk));
	jor g4183(.dina(w_n3919_4[0]),.dinb(w_n2775_1[2]),.dout(n4268),.clk(gclk));
	jor g4184(.dina(w_n3806_3[2]),.dinb(w_n2780_1[2]),.dout(n4269),.clk(gclk));
	jor g4185(.dina(w_n3600_6[1]),.dinb(w_n2784_2[1]),.dout(n4270),.clk(gclk));
	jand g4186(.dina(n4270),.dinb(n4269),.dout(n4271),.clk(gclk));
	jand g4187(.dina(n4271),.dinb(n4268),.dout(n4272),.clk(gclk));
	jand g4188(.dina(n4272),.dinb(n4267),.dout(n4273),.clk(gclk));
	jxor g4189(.dina(n4273),.dinb(w_n56_4[1]),.dout(n4274),.clk(gclk));
	jxor g4190(.dina(w_n4274_0[1]),.dinb(w_n4266_0[1]),.dout(n4275),.clk(gclk));
	jxor g4191(.dina(w_n4275_0[1]),.dinb(w_n4221_0[1]),.dout(n4276),.clk(gclk));
	jxor g4192(.dina(w_n4276_0[1]),.dinb(w_n4218_0[1]),.dout(n4277),.clk(gclk));
	jand g4193(.dina(w_n2511_0[1]),.dinb(w_n595_0[0]),.dout(n4278),.clk(gclk));
	jand g4194(.dina(n4278),.dinb(w_n924_0[1]),.dout(n4279),.clk(gclk));
	jand g4195(.dina(w_n535_0[1]),.dinb(w_n323_1[2]),.dout(n4280),.clk(gclk));
	jand g4196(.dina(n4280),.dinb(w_n2734_0[0]),.dout(n4281),.clk(gclk));
	jand g4197(.dina(n4281),.dinb(w_n1026_0[0]),.dout(n4282),.clk(gclk));
	jand g4198(.dina(n4282),.dinb(n4279),.dout(n4283),.clk(gclk));
	jand g4199(.dina(n4283),.dinb(w_n685_0[0]),.dout(n4284),.clk(gclk));
	jand g4200(.dina(n4284),.dinb(w_n2551_0[0]),.dout(n4285),.clk(gclk));
	jand g4201(.dina(n4285),.dinb(w_n395_0[0]),.dout(n4286),.clk(gclk));
	jxor g4202(.dina(w_n4286_0[1]),.dinb(w_n4277_0[1]),.dout(n4287),.clk(gclk));
	jxor g4203(.dina(w_n4287_0[1]),.dinb(w_n4215_0[1]),.dout(n4288),.clk(gclk));
	jxor g4204(.dina(w_n4288_0[1]),.dinb(w_n4211_0[1]),.dout(n4289),.clk(gclk));
	jor g4205(.dina(w_n4209_0[0]),.dinb(w_n4123_0[0]),.dout(n4290),.clk(gclk));
	jand g4206(.dina(w_n4290_0[1]),.dinb(w_n4013_9[2]),.dout(n4291),.clk(gclk));
	jxor g4207(.dina(n4291),.dinb(w_n4289_0[1]),.dout(w_dff_A_fQgYMzmB5_2),.clk(gclk));
	jand g4208(.dina(w_n4288_0[0]),.dinb(w_n4211_0[0]),.dout(n4293),.clk(gclk));
	jnot g4209(.din(w_n4277_0[0]),.dout(n4294),.clk(gclk));
	jor g4210(.dina(w_n4286_0[0]),.dinb(n4294),.dout(n4295),.clk(gclk));
	jor g4211(.dina(w_n4287_0[0]),.dinb(w_n4215_0[0]),.dout(n4296),.clk(gclk));
	jand g4212(.dina(n4296),.dinb(n4295),.dout(n4297),.clk(gclk));
	jand g4213(.dina(w_n4275_0[0]),.dinb(w_n4221_0[0]),.dout(n4298),.clk(gclk));
	jand g4214(.dina(w_n4276_0[0]),.dinb(w_n4218_0[0]),.dout(n4299),.clk(gclk));
	jor g4215(.dina(n4299),.dinb(n4298),.dout(n4300),.clk(gclk));
	jand g4216(.dina(w_n4265_0[0]),.dinb(w_n4224_0[0]),.dout(n4301),.clk(gclk));
	jand g4217(.dina(w_n4274_0[0]),.dinb(w_n4266_0[0]),.dout(n4302),.clk(gclk));
	jor g4218(.dina(n4302),.dinb(n4301),.dout(n4303),.clk(gclk));
	jand g4219(.dina(w_n4090_1[1]),.dinb(w_n78_0[2]),.dout(n4304),.clk(gclk));
	jand g4220(.dina(w_n3807_2[1]),.dinb(w_n2783_0[2]),.dout(n4305),.clk(gclk));
	jand g4221(.dina(w_n3920_2[2]),.dinb(w_n2779_0[2]),.dout(n4306),.clk(gclk));
	jor g4222(.dina(n4306),.dinb(n4305),.dout(n4307),.clk(gclk));
	jor g4223(.dina(n4307),.dinb(n4304),.dout(n4308),.clk(gclk));
	jxor g4224(.dina(n4308),.dinb(w_n55_3[2]),.dout(n4309),.clk(gclk));
	jand g4225(.dina(w_n4263_0[0]),.dinb(w_n4236_0[0]),.dout(n4310),.clk(gclk));
	jand g4226(.dina(w_n4264_0[0]),.dinb(w_n4233_0[0]),.dout(n4311),.clk(gclk));
	jor g4227(.dina(n4311),.dinb(n4310),.dout(n4312),.clk(gclk));
	jor g4228(.dina(w_n3605_1[0]),.dinb(w_n2795_3[0]),.dout(n4313),.clk(gclk));
	jor g4229(.dina(w_n3600_6[0]),.dinb(w_n2800_2[1]),.dout(n4314),.clk(gclk));
	jor g4230(.dina(w_n3315_4[2]),.dinb(w_n2805_2[1]),.dout(n4315),.clk(gclk));
	jor g4231(.dina(w_n3283_4[2]),.dinb(w_n2809_3[0]),.dout(n4316),.clk(gclk));
	jand g4232(.dina(n4316),.dinb(n4315),.dout(n4317),.clk(gclk));
	jand g4233(.dina(n4317),.dinb(n4314),.dout(n4318),.clk(gclk));
	jand g4234(.dina(n4318),.dinb(n4313),.dout(n4319),.clk(gclk));
	jxor g4235(.dina(n4319),.dinb(w_n699_5[1]),.dout(n4320),.clk(gclk));
	jnot g4236(.din(n4320),.dout(n4321),.clk(gclk));
	jand g4237(.dina(w_n4253_0[0]),.dinb(w_n4248_0[0]),.dout(n4322),.clk(gclk));
	jand g4238(.dina(w_n4262_0[0]),.dinb(w_n4254_0[0]),.dout(n4323),.clk(gclk));
	jor g4239(.dina(n4323),.dinb(n4322),.dout(n4324),.clk(gclk));
	jor g4240(.dina(w_n3516_0[2]),.dinb(w_n2857_4[0]),.dout(n4325),.clk(gclk));
	jor g4241(.dina(w_n3284_4[2]),.dinb(w_n2860_3[1]),.dout(n4326),.clk(gclk));
	jor g4242(.dina(w_n3172_3[0]),.dinb(w_n2865_3[1]),.dout(n4327),.clk(gclk));
	jor g4243(.dina(w_n2863_4[0]),.dinb(w_n2773_2[0]),.dout(n4328),.clk(gclk));
	jand g4244(.dina(n4328),.dinb(n4327),.dout(n4329),.clk(gclk));
	jand g4245(.dina(n4329),.dinb(n4326),.dout(n4330),.clk(gclk));
	jand g4246(.dina(n4330),.dinb(n4325),.dout(n4331),.clk(gclk));
	jxor g4247(.dina(n4331),.dinb(w_n808_6[2]),.dout(n4332),.clk(gclk));
	jand g4248(.dina(w_n3016_0[1]),.dinb(w_n2883_2[0]),.dout(n4333),.clk(gclk));
	jand g4249(.dina(w_n2889_1[2]),.dinb(w_n2670_2[1]),.dout(n4334),.clk(gclk));
	jand g4250(.dina(w_n2995_2[1]),.dinb(w_n2677_1[2]),.dout(n4335),.clk(gclk));
	jand g4251(.dina(w_n2887_2[0]),.dinb(w_n2672_1[0]),.dout(n4336),.clk(gclk));
	jor g4252(.dina(n4336),.dinb(n4335),.dout(n4337),.clk(gclk));
	jor g4253(.dina(n4337),.dinb(n4334),.dout(n4338),.clk(gclk));
	jor g4254(.dina(n4338),.dinb(n4333),.dout(n4339),.clk(gclk));
	jxor g4255(.dina(n4339),.dinb(w_n954_14[1]),.dout(n4340),.clk(gclk));
	jand g4256(.dina(w_n4246_0[0]),.dinb(w_n68_3[2]),.dout(n4341),.clk(gclk));
	jand g4257(.dina(w_n4247_0[0]),.dinb(w_n4245_0[0]),.dout(n4342),.clk(gclk));
	jor g4258(.dina(n4342),.dinb(n4341),.dout(n4343),.clk(gclk));
	jand g4259(.dina(w_n2679_1[0]),.dinb(w_n954_14[0]),.dout(n4344),.clk(gclk));
	jxor g4260(.dina(w_n4344_0[1]),.dinb(w_n68_3[1]),.dout(n4345),.clk(gclk));
	jxor g4261(.dina(w_n4345_0[1]),.dinb(w_n4343_0[1]),.dout(n4346),.clk(gclk));
	jxor g4262(.dina(w_n4346_0[1]),.dinb(w_n4340_0[1]),.dout(n4347),.clk(gclk));
	jxor g4263(.dina(w_n4347_0[1]),.dinb(w_n4332_0[1]),.dout(n4348),.clk(gclk));
	jxor g4264(.dina(w_n4348_0[1]),.dinb(w_n4324_0[1]),.dout(n4349),.clk(gclk));
	jxor g4265(.dina(w_n4349_0[1]),.dinb(w_n4321_0[1]),.dout(n4350),.clk(gclk));
	jxor g4266(.dina(w_n4350_0[1]),.dinb(w_n4312_0[1]),.dout(n4351),.clk(gclk));
	jxor g4267(.dina(w_n4351_0[1]),.dinb(w_n4309_0[1]),.dout(n4352),.clk(gclk));
	jxor g4268(.dina(w_n4352_0[1]),.dinb(w_n4303_0[1]),.dout(n4353),.clk(gclk));
	jxor g4269(.dina(w_n4353_0[1]),.dinb(w_n4300_0[1]),.dout(n4354),.clk(gclk));
	jand g4270(.dina(w_n2385_0[2]),.dinb(w_n3634_0[0]),.dout(n4355),.clk(gclk));
	jand g4271(.dina(w_n488_0[1]),.dinb(w_n427_1[0]),.dout(n4356),.clk(gclk));
	jand g4272(.dina(n4356),.dinb(w_n451_1[0]),.dout(n4357),.clk(gclk));
	jand g4273(.dina(w_n4357_0[2]),.dinb(w_n4355_0[1]),.dout(n4358),.clk(gclk));
	jand g4274(.dina(n4358),.dinb(w_n4000_0[1]),.dout(n4359),.clk(gclk));
	jand g4275(.dina(w_n849_0[2]),.dinb(w_n216_1[1]),.dout(n4360),.clk(gclk));
	jand g4276(.dina(w_n445_0[2]),.dinb(w_n225_0[2]),.dout(n4361),.clk(gclk));
	jand g4277(.dina(n4361),.dinb(n4360),.dout(n4362),.clk(gclk));
	jand g4278(.dina(w_n934_0[0]),.dinb(w_n286_0[1]),.dout(n4363),.clk(gclk));
	jand g4279(.dina(n4363),.dinb(n4362),.dout(n4364),.clk(gclk));
	jand g4280(.dina(n4364),.dinb(w_n2402_0[0]),.dout(n4365),.clk(gclk));
	jand g4281(.dina(n4365),.dinb(n4359),.dout(n4366),.clk(gclk));
	jand g4282(.dina(n4366),.dinb(w_n3909_0[0]),.dout(n4367),.clk(gclk));
	jand g4283(.dina(n4367),.dinb(w_n3256_0[1]),.dout(n4368),.clk(gclk));
	jxor g4284(.dina(w_n4368_0[1]),.dinb(w_n4354_0[1]),.dout(n4369),.clk(gclk));
	jxor g4285(.dina(w_n4369_0[1]),.dinb(w_n4297_0[1]),.dout(n4370),.clk(gclk));
	jxor g4286(.dina(w_n4370_0[1]),.dinb(w_n4293_0[1]),.dout(n4371),.clk(gclk));
	jor g4287(.dina(w_n4290_0[0]),.dinb(w_n4289_0[0]),.dout(n4372),.clk(gclk));
	jand g4288(.dina(w_n4372_0[1]),.dinb(w_n4013_9[1]),.dout(n4373),.clk(gclk));
	jxor g4289(.dina(n4373),.dinb(w_n4371_0[1]),.dout(w_dff_A_Zdk0dlCk2_2),.clk(gclk));
	jand g4290(.dina(w_n4370_0[0]),.dinb(w_n4293_0[0]),.dout(n4375),.clk(gclk));
	jnot g4291(.din(w_n4354_0[0]),.dout(n4376),.clk(gclk));
	jor g4292(.dina(w_n4368_0[0]),.dinb(n4376),.dout(n4377),.clk(gclk));
	jor g4293(.dina(w_n4369_0[0]),.dinb(w_n4297_0[0]),.dout(n4378),.clk(gclk));
	jand g4294(.dina(n4378),.dinb(n4377),.dout(n4379),.clk(gclk));
	jand g4295(.dina(w_n4352_0[0]),.dinb(w_n4303_0[0]),.dout(n4380),.clk(gclk));
	jand g4296(.dina(w_n4353_0[0]),.dinb(w_n4300_0[0]),.dout(n4381),.clk(gclk));
	jor g4297(.dina(n4381),.dinb(n4380),.dout(n4382),.clk(gclk));
	jand g4298(.dina(w_n4350_0[0]),.dinb(w_n4312_0[0]),.dout(n4383),.clk(gclk));
	jand g4299(.dina(w_n4351_0[0]),.dinb(w_n4309_0[0]),.dout(n4384),.clk(gclk));
	jor g4300(.dina(n4384),.dinb(n4383),.dout(n4385),.clk(gclk));
	jand g4301(.dina(w_n4348_0[0]),.dinb(w_n4324_0[0]),.dout(n4386),.clk(gclk));
	jand g4302(.dina(w_n4349_0[0]),.dinb(w_n4321_0[0]),.dout(n4387),.clk(gclk));
	jor g4303(.dina(n4387),.dinb(n4386),.dout(n4388),.clk(gclk));
	jnot g4304(.din(n4388),.dout(n4389),.clk(gclk));
	jor g4305(.dina(w_n4136_1[1]),.dinb(w_n79_2[0]),.dout(n4390),.clk(gclk));
	jand g4306(.dina(n4390),.dinb(w_n2784_2[0]),.dout(n4391),.clk(gclk));
	jor g4307(.dina(n4391),.dinb(w_n3919_3[2]),.dout(n4392),.clk(gclk));
	jxor g4308(.dina(n4392),.dinb(w_n55_3[1]),.dout(n4393),.clk(gclk));
	jxor g4309(.dina(w_n4393_0[1]),.dinb(w_n4389_0[1]),.dout(n4394),.clk(gclk));
	jor g4310(.dina(w_n3811_1[0]),.dinb(w_n2795_2[2]),.dout(n4395),.clk(gclk));
	jor g4311(.dina(w_n3806_3[1]),.dinb(w_n2800_2[0]),.dout(n4396),.clk(gclk));
	jor g4312(.dina(w_n3600_5[2]),.dinb(w_n2805_2[0]),.dout(n4397),.clk(gclk));
	jor g4313(.dina(w_n3315_4[1]),.dinb(w_n2809_2[2]),.dout(n4398),.clk(gclk));
	jand g4314(.dina(n4398),.dinb(n4397),.dout(n4399),.clk(gclk));
	jand g4315(.dina(n4399),.dinb(n4396),.dout(n4400),.clk(gclk));
	jand g4316(.dina(n4400),.dinb(n4395),.dout(n4401),.clk(gclk));
	jxor g4317(.dina(n4401),.dinb(w_n699_5[0]),.dout(n4402),.clk(gclk));
	jnot g4318(.din(n4402),.dout(n4403),.clk(gclk));
	jand g4319(.dina(w_n4346_0[0]),.dinb(w_n4340_0[0]),.dout(n4404),.clk(gclk));
	jand g4320(.dina(w_n4347_0[0]),.dinb(w_n4332_0[0]),.dout(n4405),.clk(gclk));
	jor g4321(.dina(n4405),.dinb(n4404),.dout(n4406),.clk(gclk));
	jor g4322(.dina(w_n3337_0[2]),.dinb(w_n2857_3[2]),.dout(n4407),.clk(gclk));
	jor g4323(.dina(w_n3283_4[1]),.dinb(w_n2860_3[0]),.dout(n4408),.clk(gclk));
	jor g4324(.dina(w_n3284_4[1]),.dinb(w_n2865_3[0]),.dout(n4409),.clk(gclk));
	jor g4325(.dina(w_n3172_2[2]),.dinb(w_n2863_3[2]),.dout(n4410),.clk(gclk));
	jand g4326(.dina(n4410),.dinb(n4409),.dout(n4411),.clk(gclk));
	jand g4327(.dina(n4411),.dinb(n4408),.dout(n4412),.clk(gclk));
	jand g4328(.dina(n4412),.dinb(n4407),.dout(n4413),.clk(gclk));
	jxor g4329(.dina(n4413),.dinb(w_n808_6[1]),.dout(n4414),.clk(gclk));
	jor g4330(.dina(w_n3198_3[2]),.dinb(w_n2771_0[1]),.dout(n4415),.clk(gclk));
	jor g4331(.dina(w_n3200_3[0]),.dinb(w_n2773_1[2]),.dout(n4416),.clk(gclk));
	jor g4332(.dina(w_n3204_3[0]),.dinb(w_n2669_1[1]),.dout(n4417),.clk(gclk));
	jor g4333(.dina(w_n3202_3[0]),.dinb(w_n2671_2[0]),.dout(n4418),.clk(gclk));
	jand g4334(.dina(n4418),.dinb(n4417),.dout(n4419),.clk(gclk));
	jand g4335(.dina(n4419),.dinb(n4416),.dout(n4420),.clk(gclk));
	jand g4336(.dina(n4420),.dinb(n4415),.dout(n4421),.clk(gclk));
	jxor g4337(.dina(n4421),.dinb(w_n820_3[1]),.dout(n4422),.clk(gclk));
	jand g4338(.dina(w_n4344_0[0]),.dinb(w_n68_3[0]),.dout(n4423),.clk(gclk));
	jand g4339(.dina(w_n4345_0[0]),.dinb(w_n4343_0[0]),.dout(n4424),.clk(gclk));
	jor g4340(.dina(n4424),.dinb(n4423),.dout(n4425),.clk(gclk));
	jand g4341(.dina(w_n2677_1[1]),.dinb(w_n954_13[2]),.dout(n4426),.clk(gclk));
	jxor g4342(.dina(w_n4426_0[1]),.dinb(w_n68_2[2]),.dout(n4427),.clk(gclk));
	jxor g4343(.dina(w_n4427_0[1]),.dinb(w_n4425_0[1]),.dout(n4428),.clk(gclk));
	jxor g4344(.dina(w_n4428_0[1]),.dinb(w_n4422_0[1]),.dout(n4429),.clk(gclk));
	jxor g4345(.dina(w_n4429_0[1]),.dinb(w_n4414_0[1]),.dout(n4430),.clk(gclk));
	jxor g4346(.dina(w_n4430_0[1]),.dinb(w_n4406_0[1]),.dout(n4431),.clk(gclk));
	jxor g4347(.dina(w_n4431_0[1]),.dinb(w_n4403_0[1]),.dout(n4432),.clk(gclk));
	jxor g4348(.dina(w_n4432_0[1]),.dinb(w_n4394_0[1]),.dout(n4433),.clk(gclk));
	jxor g4349(.dina(w_n4433_0[1]),.dinb(w_n4385_0[1]),.dout(n4434),.clk(gclk));
	jxor g4350(.dina(w_n4434_0[1]),.dinb(w_n4382_0[1]),.dout(n4435),.clk(gclk));
	jand g4351(.dina(w_n2429_0[1]),.dinb(w_n763_0[2]),.dout(n4436),.clk(gclk));
	jand g4352(.dina(n4436),.dinb(w_n3911_0[0]),.dout(n4437),.clk(gclk));
	jand g4353(.dina(n4437),.dinb(w_n2541_0[0]),.dout(n4438),.clk(gclk));
	jand g4354(.dina(w_n865_0[0]),.dinb(w_n822_1[0]),.dout(n4439),.clk(gclk));
	jand g4355(.dina(n4439),.dinb(w_n2385_0[1]),.dout(n4440),.clk(gclk));
	jand g4356(.dina(n4440),.dinb(w_n2514_0[0]),.dout(n4441),.clk(gclk));
	jand g4357(.dina(n4441),.dinb(n4438),.dout(n4442),.clk(gclk));
	jand g4358(.dina(w_n401_0[2]),.dinb(w_n379_0[1]),.dout(n4443),.clk(gclk));
	jand g4359(.dina(n4443),.dinb(w_n680_0[2]),.dout(n4444),.clk(gclk));
	jand g4360(.dina(w_n3307_1[1]),.dinb(w_n1294_0[0]),.dout(n4445),.clk(gclk));
	jand g4361(.dina(n4445),.dinb(w_n2387_0[0]),.dout(n4446),.clk(gclk));
	jand g4362(.dina(n4446),.dinb(n4444),.dout(n4447),.clk(gclk));
	jand g4363(.dina(n4447),.dinb(w_n2540_0[0]),.dout(n4448),.clk(gclk));
	jand g4364(.dina(n4448),.dinb(w_n4442_0[1]),.dout(n4449),.clk(gclk));
	jand g4365(.dina(n4449),.dinb(w_n3633_0[0]),.dout(n4450),.clk(gclk));
	jxor g4366(.dina(w_n4450_0[1]),.dinb(w_n4435_0[1]),.dout(n4451),.clk(gclk));
	jxor g4367(.dina(w_n4451_0[1]),.dinb(w_n4379_0[1]),.dout(n4452),.clk(gclk));
	jxor g4368(.dina(w_n4452_0[1]),.dinb(w_n4375_0[1]),.dout(n4453),.clk(gclk));
	jor g4369(.dina(w_n4372_0[0]),.dinb(w_n4371_0[0]),.dout(n4454),.clk(gclk));
	jand g4370(.dina(w_n4454_0[1]),.dinb(w_n4013_9[0]),.dout(n4455),.clk(gclk));
	jxor g4371(.dina(n4455),.dinb(w_n4453_0[1]),.dout(w_dff_A_y6UHYdvt4_2),.clk(gclk));
	jand g4372(.dina(w_n4452_0[0]),.dinb(w_n4375_0[0]),.dout(n4457),.clk(gclk));
	jnot g4373(.din(w_n4435_0[0]),.dout(n4458),.clk(gclk));
	jor g4374(.dina(w_n4450_0[0]),.dinb(n4458),.dout(n4459),.clk(gclk));
	jor g4375(.dina(w_n4451_0[0]),.dinb(w_n4379_0[0]),.dout(n4460),.clk(gclk));
	jand g4376(.dina(n4460),.dinb(n4459),.dout(n4461),.clk(gclk));
	jand g4377(.dina(w_n4433_0[0]),.dinb(w_n4385_0[0]),.dout(n4462),.clk(gclk));
	jand g4378(.dina(w_n4434_0[0]),.dinb(w_n4382_0[0]),.dout(n4463),.clk(gclk));
	jor g4379(.dina(n4463),.dinb(n4462),.dout(n4464),.clk(gclk));
	jor g4380(.dina(w_n4393_0[0]),.dinb(w_n4389_0[0]),.dout(n4465),.clk(gclk));
	jand g4381(.dina(w_n4432_0[0]),.dinb(w_n4394_0[0]),.dout(n4466),.clk(gclk));
	jnot g4382(.din(n4466),.dout(n4467),.clk(gclk));
	jand g4383(.dina(n4467),.dinb(n4465),.dout(n4468),.clk(gclk));
	jnot g4384(.din(n4468),.dout(n4469),.clk(gclk));
	jand g4385(.dina(w_n4430_0[0]),.dinb(w_n4406_0[0]),.dout(n4470),.clk(gclk));
	jand g4386(.dina(w_n4431_0[0]),.dinb(w_n4403_0[0]),.dout(n4471),.clk(gclk));
	jor g4387(.dina(n4471),.dinb(n4470),.dout(n4472),.clk(gclk));
	jor g4388(.dina(w_n3927_1[0]),.dinb(w_n2795_2[1]),.dout(n4473),.clk(gclk));
	jor g4389(.dina(w_n3919_3[1]),.dinb(w_n2800_1[2]),.dout(n4474),.clk(gclk));
	jor g4390(.dina(w_n3806_3[0]),.dinb(w_n2805_1[2]),.dout(n4475),.clk(gclk));
	jor g4391(.dina(w_n3600_5[1]),.dinb(w_n2809_2[1]),.dout(n4476),.clk(gclk));
	jand g4392(.dina(n4476),.dinb(n4475),.dout(n4477),.clk(gclk));
	jand g4393(.dina(n4477),.dinb(n4474),.dout(n4478),.clk(gclk));
	jand g4394(.dina(n4478),.dinb(n4473),.dout(n4479),.clk(gclk));
	jxor g4395(.dina(n4479),.dinb(w_n1143_4[0]),.dout(n4480),.clk(gclk));
	jxor g4396(.dina(w_n4480_0[1]),.dinb(w_n4472_0[1]),.dout(n4481),.clk(gclk));
	jand g4397(.dina(w_n4428_0[0]),.dinb(w_n4422_0[0]),.dout(n4482),.clk(gclk));
	jand g4398(.dina(w_n4429_0[0]),.dinb(w_n4414_0[0]),.dout(n4483),.clk(gclk));
	jor g4399(.dina(n4483),.dinb(n4482),.dout(n4484),.clk(gclk));
	jand g4400(.dina(w_n4426_0[0]),.dinb(w_n68_2[1]),.dout(n4485),.clk(gclk));
	jand g4401(.dina(w_n4427_0[0]),.dinb(w_n4425_0[0]),.dout(n4486),.clk(gclk));
	jor g4402(.dina(n4486),.dinb(n4485),.dout(n4487),.clk(gclk));
	jand g4403(.dina(w_n3174_0[1]),.dinb(w_n2883_1[2]),.dout(n4488),.clk(gclk));
	jand g4404(.dina(w_n3176_1[0]),.dinb(w_n2889_1[1]),.dout(n4489),.clk(gclk));
	jand g4405(.dina(w_n2995_2[0]),.dinb(w_n2670_2[0]),.dout(n4490),.clk(gclk));
	jand g4406(.dina(w_n2887_1[2]),.dinb(w_n2769_1[2]),.dout(n4491),.clk(gclk));
	jor g4407(.dina(n4491),.dinb(n4490),.dout(n4492),.clk(gclk));
	jor g4408(.dina(n4492),.dinb(n4489),.dout(n4493),.clk(gclk));
	jor g4409(.dina(n4493),.dinb(n4488),.dout(n4494),.clk(gclk));
	jxor g4410(.dina(n4494),.dinb(w_n820_3[0]),.dout(n4495),.clk(gclk));
	jnot g4411(.din(n4495),.dout(n4496),.clk(gclk));
	jand g4412(.dina(w_n2672_0[2]),.dinb(w_n954_13[1]),.dout(n4497),.clk(gclk));
	jxor g4413(.dina(w_n68_2[0]),.dinb(w_n55_3[0]),.dout(n4498),.clk(gclk));
	jxor g4414(.dina(w_n4498_0[1]),.dinb(w_n4497_0[1]),.dout(n4499),.clk(gclk));
	jxor g4415(.dina(w_n4499_0[1]),.dinb(w_n4496_0[1]),.dout(n4500),.clk(gclk));
	jxor g4416(.dina(w_n4500_0[1]),.dinb(w_n4487_0[1]),.dout(n4501),.clk(gclk));
	jor g4417(.dina(w_n3320_0[2]),.dinb(w_n2857_3[1]),.dout(n4502),.clk(gclk));
	jor g4418(.dina(w_n3315_4[0]),.dinb(w_n2860_2[2]),.dout(n4503),.clk(gclk));
	jor g4419(.dina(w_n3283_4[0]),.dinb(w_n2865_2[2]),.dout(n4504),.clk(gclk));
	jor g4420(.dina(w_n3284_4[0]),.dinb(w_n2863_3[1]),.dout(n4505),.clk(gclk));
	jand g4421(.dina(n4505),.dinb(n4504),.dout(n4506),.clk(gclk));
	jand g4422(.dina(n4506),.dinb(n4503),.dout(n4507),.clk(gclk));
	jand g4423(.dina(n4507),.dinb(n4502),.dout(n4508),.clk(gclk));
	jxor g4424(.dina(n4508),.dinb(w_n808_6[0]),.dout(n4509),.clk(gclk));
	jxor g4425(.dina(w_n4509_0[1]),.dinb(w_n4501_0[1]),.dout(n4510),.clk(gclk));
	jxor g4426(.dina(w_n4510_0[1]),.dinb(w_n4484_0[1]),.dout(n4511),.clk(gclk));
	jxor g4427(.dina(w_n4511_0[1]),.dinb(w_n4481_0[1]),.dout(n4512),.clk(gclk));
	jxor g4428(.dina(w_n4512_0[1]),.dinb(w_n4469_0[1]),.dout(n4513),.clk(gclk));
	jxor g4429(.dina(w_n4513_0[1]),.dinb(w_n4464_0[1]),.dout(n4514),.clk(gclk));
	jand g4430(.dina(w_n1188_0[0]),.dinb(w_n471_0[0]),.dout(n4515),.clk(gclk));
	jand g4431(.dina(w_n2406_0[0]),.dinb(w_n1170_0[0]),.dout(n4516),.clk(gclk));
	jand g4432(.dina(n4516),.dinb(n4515),.dout(n4517),.clk(gclk));
	jand g4433(.dina(w_n270_0[2]),.dinb(w_n214_1[0]),.dout(n4518),.clk(gclk));
	jand g4434(.dina(n4518),.dinb(w_n930_0[2]),.dout(n4519),.clk(gclk));
	jand g4435(.dina(n4519),.dinb(w_n4357_0[1]),.dout(n4520),.clk(gclk));
	jand g4436(.dina(n4520),.dinb(n4517),.dout(n4521),.clk(gclk));
	jand g4437(.dina(n4521),.dinb(w_n4442_0[0]),.dout(n4522),.clk(gclk));
	jand g4438(.dina(n4522),.dinb(w_n2350_0[0]),.dout(n4523),.clk(gclk));
	jxor g4439(.dina(w_n4523_0[1]),.dinb(w_n4514_0[1]),.dout(n4524),.clk(gclk));
	jxor g4440(.dina(w_n4524_0[1]),.dinb(w_n4461_0[1]),.dout(n4525),.clk(gclk));
	jxor g4441(.dina(w_n4525_0[1]),.dinb(w_n4457_0[1]),.dout(n4526),.clk(gclk));
	jor g4442(.dina(w_n4454_0[0]),.dinb(w_n4453_0[0]),.dout(n4527),.clk(gclk));
	jand g4443(.dina(w_n4527_0[1]),.dinb(w_n4013_8[2]),.dout(n4528),.clk(gclk));
	jxor g4444(.dina(n4528),.dinb(w_n4526_0[1]),.dout(w_dff_A_RryB5Bx36_2),.clk(gclk));
	jand g4445(.dina(w_n4525_0[0]),.dinb(w_n4457_0[0]),.dout(n4530),.clk(gclk));
	jnot g4446(.din(w_n4514_0[0]),.dout(n4531),.clk(gclk));
	jor g4447(.dina(w_n4523_0[0]),.dinb(n4531),.dout(n4532),.clk(gclk));
	jor g4448(.dina(w_n4524_0[0]),.dinb(w_n4461_0[0]),.dout(n4533),.clk(gclk));
	jand g4449(.dina(n4533),.dinb(n4532),.dout(n4534),.clk(gclk));
	jand g4450(.dina(w_n4512_0[0]),.dinb(w_n4469_0[0]),.dout(n4535),.clk(gclk));
	jand g4451(.dina(w_n4513_0[0]),.dinb(w_n4464_0[0]),.dout(n4536),.clk(gclk));
	jor g4452(.dina(n4536),.dinb(n4535),.dout(n4537),.clk(gclk));
	jand g4453(.dina(w_n4480_0[0]),.dinb(w_n4472_0[0]),.dout(n4538),.clk(gclk));
	jand g4454(.dina(w_n4511_0[0]),.dinb(w_n4481_0[0]),.dout(n4539),.clk(gclk));
	jor g4455(.dina(n4539),.dinb(n4538),.dout(n4540),.clk(gclk));
	jand g4456(.dina(w_n4090_1[0]),.dinb(w_n2794_0[2]),.dout(n4541),.clk(gclk));
	jand g4457(.dina(w_n3807_2[0]),.dinb(w_n2808_0[2]),.dout(n4542),.clk(gclk));
	jand g4458(.dina(w_n3920_2[1]),.dinb(w_n2804_0[2]),.dout(n4543),.clk(gclk));
	jor g4459(.dina(n4543),.dinb(n4542),.dout(n4544),.clk(gclk));
	jor g4460(.dina(n4544),.dinb(n4541),.dout(n4545),.clk(gclk));
	jxor g4461(.dina(n4545),.dinb(w_n1143_3[2]),.dout(n4546),.clk(gclk));
	jnot g4462(.din(n4546),.dout(n4547),.clk(gclk));
	jand g4463(.dina(w_n4509_0[0]),.dinb(w_n4501_0[0]),.dout(n4548),.clk(gclk));
	jand g4464(.dina(w_n4510_0[0]),.dinb(w_n4484_0[0]),.dout(n4549),.clk(gclk));
	jor g4465(.dina(n4549),.dinb(n4548),.dout(n4550),.clk(gclk));
	jor g4466(.dina(w_n3605_0[2]),.dinb(w_n2857_3[0]),.dout(n4551),.clk(gclk));
	jor g4467(.dina(w_n3600_5[0]),.dinb(w_n2860_2[1]),.dout(n4552),.clk(gclk));
	jor g4468(.dina(w_n3315_3[2]),.dinb(w_n2865_2[1]),.dout(n4553),.clk(gclk));
	jor g4469(.dina(w_n3283_3[2]),.dinb(w_n2863_3[0]),.dout(n4554),.clk(gclk));
	jand g4470(.dina(n4554),.dinb(n4553),.dout(n4555),.clk(gclk));
	jand g4471(.dina(n4555),.dinb(n4552),.dout(n4556),.clk(gclk));
	jand g4472(.dina(n4556),.dinb(n4551),.dout(n4557),.clk(gclk));
	jxor g4473(.dina(n4557),.dinb(w_n808_5[2]),.dout(n4558),.clk(gclk));
	jand g4474(.dina(w_n4499_0[0]),.dinb(w_n4496_0[0]),.dout(n4559),.clk(gclk));
	jand g4475(.dina(w_n4500_0[0]),.dinb(w_n4487_0[0]),.dout(n4560),.clk(gclk));
	jor g4476(.dina(n4560),.dinb(n4559),.dout(n4561),.clk(gclk));
	jor g4477(.dina(w_n3516_0[1]),.dinb(w_n3198_3[1]),.dout(n4562),.clk(gclk));
	jor g4478(.dina(w_n3284_3[2]),.dinb(w_n3200_2[2]),.dout(n4563),.clk(gclk));
	jor g4479(.dina(w_n3172_2[1]),.dinb(w_n3204_2[2]),.dout(n4564),.clk(gclk));
	jor g4480(.dina(w_n3202_2[2]),.dinb(w_n2773_1[1]),.dout(n4565),.clk(gclk));
	jand g4481(.dina(n4565),.dinb(n4564),.dout(n4566),.clk(gclk));
	jand g4482(.dina(n4566),.dinb(n4563),.dout(n4567),.clk(gclk));
	jand g4483(.dina(n4567),.dinb(n4562),.dout(n4568),.clk(gclk));
	jxor g4484(.dina(n4568),.dinb(w_n820_2[2]),.dout(n4569),.clk(gclk));
	jand g4485(.dina(w_n2670_1[2]),.dinb(w_n954_13[0]),.dout(n4570),.clk(gclk));
	jnot g4486(.din(w_n4570_0[1]),.dout(n4571),.clk(gclk));
	jand g4487(.dina(w_n3233_3[0]),.dinb(w_n56_4[0]),.dout(n4572),.clk(gclk));
	jand g4488(.dina(w_n4498_0[0]),.dinb(w_n4497_0[0]),.dout(n4573),.clk(gclk));
	jor g4489(.dina(n4573),.dinb(n4572),.dout(n4574),.clk(gclk));
	jxor g4490(.dina(w_n4574_0[1]),.dinb(w_n4571_0[2]),.dout(n4575),.clk(gclk));
	jxor g4491(.dina(w_n4575_0[1]),.dinb(w_n4569_0[1]),.dout(n4576),.clk(gclk));
	jxor g4492(.dina(w_n4576_0[1]),.dinb(w_n4561_0[1]),.dout(n4577),.clk(gclk));
	jxor g4493(.dina(w_n4577_0[1]),.dinb(w_n4558_0[1]),.dout(n4578),.clk(gclk));
	jxor g4494(.dina(w_n4578_0[1]),.dinb(w_n4550_0[1]),.dout(n4579),.clk(gclk));
	jxor g4495(.dina(w_n4579_0[1]),.dinb(w_n4547_0[1]),.dout(n4580),.clk(gclk));
	jxor g4496(.dina(w_n4580_0[1]),.dinb(w_n4540_0[1]),.dout(n4581),.clk(gclk));
	jxor g4497(.dina(w_n4581_0[1]),.dinb(w_n4537_0[1]),.dout(n4582),.clk(gclk));
	jand g4498(.dina(w_n421_1[1]),.dinb(w_n147_1[2]),.dout(n4583),.clk(gclk));
	jand g4499(.dina(n4583),.dinb(w_n295_1[0]),.dout(n4584),.clk(gclk));
	jand g4500(.dina(w_n735_0[0]),.dinb(w_n638_0[0]),.dout(n4585),.clk(gclk));
	jand g4501(.dina(n4585),.dinb(w_n3626_0[0]),.dout(n4586),.clk(gclk));
	jand g4502(.dina(n4586),.dinb(n4584),.dout(n4587),.clk(gclk));
	jand g4503(.dina(n4587),.dinb(w_n2571_0[0]),.dout(n4588),.clk(gclk));
	jand g4504(.dina(n4588),.dinb(w_n832_0[1]),.dout(n4589),.clk(gclk));
	jand g4505(.dina(w_n277_2[0]),.dinb(w_n229_0[2]),.dout(n4590),.clk(gclk));
	jand g4506(.dina(n4590),.dinb(w_n410_0[1]),.dout(n4591),.clk(gclk));
	jand g4507(.dina(w_n765_0[1]),.dinb(w_n751_0[2]),.dout(n4592),.clk(gclk));
	jand g4508(.dina(n4592),.dinb(w_n2424_0[0]),.dout(n4593),.clk(gclk));
	jand g4509(.dina(n4593),.dinb(n4591),.dout(n4594),.clk(gclk));
	jand g4510(.dina(w_n2428_0[0]),.dinb(w_n667_0[0]),.dout(n4595),.clk(gclk));
	jand g4511(.dina(n4595),.dinb(n4594),.dout(n4596),.clk(gclk));
	jand g4512(.dina(n4596),.dinb(w_n655_0[0]),.dout(n4597),.clk(gclk));
	jand g4513(.dina(n4597),.dinb(w_n4589_0[1]),.dout(n4598),.clk(gclk));
	jand g4514(.dina(n4598),.dinb(w_n3666_0[0]),.dout(n4599),.clk(gclk));
	jxor g4515(.dina(w_n4599_0[1]),.dinb(w_n4582_0[1]),.dout(n4600),.clk(gclk));
	jxor g4516(.dina(w_n4600_0[1]),.dinb(w_n4534_0[1]),.dout(n4601),.clk(gclk));
	jxor g4517(.dina(w_n4601_0[1]),.dinb(w_n4530_0[1]),.dout(n4602),.clk(gclk));
	jor g4518(.dina(w_n4527_0[0]),.dinb(w_n4526_0[0]),.dout(n4603),.clk(gclk));
	jand g4519(.dina(w_n4603_0[1]),.dinb(w_n4013_8[1]),.dout(n4604),.clk(gclk));
	jxor g4520(.dina(n4604),.dinb(w_n4602_0[1]),.dout(w_dff_A_bZHWsZ3E8_2),.clk(gclk));
	jand g4521(.dina(w_n4601_0[0]),.dinb(w_n4530_0[0]),.dout(n4606),.clk(gclk));
	jnot g4522(.din(w_n4582_0[0]),.dout(n4607),.clk(gclk));
	jor g4523(.dina(w_n4599_0[0]),.dinb(n4607),.dout(n4608),.clk(gclk));
	jor g4524(.dina(w_n4600_0[0]),.dinb(w_n4534_0[0]),.dout(n4609),.clk(gclk));
	jand g4525(.dina(n4609),.dinb(n4608),.dout(n4610),.clk(gclk));
	jand g4526(.dina(w_n4580_0[0]),.dinb(w_n4540_0[0]),.dout(n4611),.clk(gclk));
	jand g4527(.dina(w_n4581_0[0]),.dinb(w_n4537_0[0]),.dout(n4612),.clk(gclk));
	jor g4528(.dina(n4612),.dinb(n4611),.dout(n4613),.clk(gclk));
	jand g4529(.dina(w_n4578_0[0]),.dinb(w_n4550_0[0]),.dout(n4614),.clk(gclk));
	jand g4530(.dina(w_n4579_0[0]),.dinb(w_n4547_0[0]),.dout(n4615),.clk(gclk));
	jor g4531(.dina(n4615),.dinb(n4614),.dout(n4616),.clk(gclk));
	jand g4532(.dina(w_n4576_0[0]),.dinb(w_n4561_0[0]),.dout(n4617),.clk(gclk));
	jand g4533(.dina(w_n4577_0[0]),.dinb(w_n4558_0[0]),.dout(n4618),.clk(gclk));
	jor g4534(.dina(n4618),.dinb(n4617),.dout(n4619),.clk(gclk));
	jnot g4535(.din(n4619),.dout(n4620),.clk(gclk));
	jor g4536(.dina(w_n4136_1[0]),.dinb(w_n2795_2[0]),.dout(n4621),.clk(gclk));
	jand g4537(.dina(n4621),.dinb(w_n2809_2[0]),.dout(n4622),.clk(gclk));
	jor g4538(.dina(n4622),.dinb(w_n3919_3[0]),.dout(n4623),.clk(gclk));
	jxor g4539(.dina(n4623),.dinb(w_n699_4[2]),.dout(n4624),.clk(gclk));
	jxor g4540(.dina(w_n4624_0[1]),.dinb(w_n4620_0[1]),.dout(n4625),.clk(gclk));
	jand g4541(.dina(w_n4574_0[0]),.dinb(w_n4571_0[1]),.dout(n4626),.clk(gclk));
	jand g4542(.dina(w_n4575_0[0]),.dinb(w_n4569_0[0]),.dout(n4627),.clk(gclk));
	jor g4543(.dina(n4627),.dinb(n4626),.dout(n4628),.clk(gclk));
	jor g4544(.dina(w_n3337_0[1]),.dinb(w_n3198_3[0]),.dout(n4629),.clk(gclk));
	jor g4545(.dina(w_n3283_3[1]),.dinb(w_n3200_2[1]),.dout(n4630),.clk(gclk));
	jor g4546(.dina(w_n3284_3[1]),.dinb(w_n3204_2[1]),.dout(n4631),.clk(gclk));
	jor g4547(.dina(w_n3172_2[0]),.dinb(w_n3202_2[1]),.dout(n4632),.clk(gclk));
	jand g4548(.dina(n4632),.dinb(n4631),.dout(n4633),.clk(gclk));
	jand g4549(.dina(n4633),.dinb(n4630),.dout(n4634),.clk(gclk));
	jand g4550(.dina(n4634),.dinb(n4629),.dout(n4635),.clk(gclk));
	jxor g4551(.dina(n4635),.dinb(w_n954_12[2]),.dout(n4636),.clk(gclk));
	jand g4552(.dina(w_n2770_0[0]),.dinb(w_n954_12[1]),.dout(n4637),.clk(gclk));
	jxor g4553(.dina(w_n4637_0[1]),.dinb(w_n4636_0[1]),.dout(n4638),.clk(gclk));
	jxor g4554(.dina(w_n4638_0[1]),.dinb(w_n4628_0[1]),.dout(n4639),.clk(gclk));
	jor g4555(.dina(w_n3811_0[2]),.dinb(w_n2857_2[2]),.dout(n4640),.clk(gclk));
	jor g4556(.dina(w_n3806_2[2]),.dinb(w_n2860_2[0]),.dout(n4641),.clk(gclk));
	jor g4557(.dina(w_n3600_4[2]),.dinb(w_n2865_2[0]),.dout(n4642),.clk(gclk));
	jor g4558(.dina(w_n3315_3[1]),.dinb(w_n2863_2[2]),.dout(n4643),.clk(gclk));
	jand g4559(.dina(n4643),.dinb(n4642),.dout(n4644),.clk(gclk));
	jand g4560(.dina(n4644),.dinb(n4641),.dout(n4645),.clk(gclk));
	jand g4561(.dina(n4645),.dinb(n4640),.dout(n4646),.clk(gclk));
	jxor g4562(.dina(n4646),.dinb(w_n808_5[1]),.dout(n4647),.clk(gclk));
	jxor g4563(.dina(w_n4647_0[1]),.dinb(w_n4639_0[1]),.dout(n4648),.clk(gclk));
	jxor g4564(.dina(w_n4648_0[1]),.dinb(w_n4625_0[1]),.dout(n4649),.clk(gclk));
	jxor g4565(.dina(w_n4649_0[1]),.dinb(w_n4616_0[1]),.dout(n4650),.clk(gclk));
	jxor g4566(.dina(w_n4650_0[1]),.dinb(w_n4613_0[1]),.dout(n4651),.clk(gclk));
	jand g4567(.dina(w_n668_1[0]),.dinb(w_n279_0[2]),.dout(n4652),.clk(gclk));
	jand g4568(.dina(w_n645_1[0]),.dinb(w_n147_1[1]),.dout(n4653),.clk(gclk));
	jand g4569(.dina(n4653),.dinb(n4652),.dout(n4654),.clk(gclk));
	jand g4570(.dina(w_n3307_1[0]),.dinb(w_n930_0[1]),.dout(n4655),.clk(gclk));
	jand g4571(.dina(n4655),.dinb(n4654),.dout(n4656),.clk(gclk));
	jand g4572(.dina(w_n579_0[2]),.dinb(w_n390_0[1]),.dout(n4657),.clk(gclk));
	jand g4573(.dina(n4657),.dinb(w_n303_1[2]),.dout(n4658),.clk(gclk));
	jand g4574(.dina(n4658),.dinb(w_n3242_0[0]),.dout(n4659),.clk(gclk));
	jand g4575(.dina(n4659),.dinb(n4656),.dout(n4660),.clk(gclk));
	jand g4576(.dina(n4660),.dinb(w_n405_0[0]),.dout(n4661),.clk(gclk));
	jand g4577(.dina(n4661),.dinb(w_n3638_0[0]),.dout(n4662),.clk(gclk));
	jand g4578(.dina(n4662),.dinb(w_n2520_0[0]),.dout(n4663),.clk(gclk));
	jxor g4579(.dina(w_n4663_0[1]),.dinb(w_n4651_0[1]),.dout(n4664),.clk(gclk));
	jxor g4580(.dina(w_n4664_0[1]),.dinb(w_n4610_0[1]),.dout(n4665),.clk(gclk));
	jxor g4581(.dina(w_n4665_0[1]),.dinb(w_n4606_0[1]),.dout(n4666),.clk(gclk));
	jor g4582(.dina(w_n4603_0[0]),.dinb(w_n4602_0[0]),.dout(n4667),.clk(gclk));
	jand g4583(.dina(w_n4667_0[1]),.dinb(w_n4013_8[0]),.dout(n4668),.clk(gclk));
	jxor g4584(.dina(n4668),.dinb(w_n4666_0[1]),.dout(w_dff_A_u8ZD7jxR4_2),.clk(gclk));
	jand g4585(.dina(w_n4665_0[0]),.dinb(w_n4606_0[0]),.dout(n4670),.clk(gclk));
	jnot g4586(.din(w_n4651_0[0]),.dout(n4671),.clk(gclk));
	jor g4587(.dina(w_n4663_0[0]),.dinb(n4671),.dout(n4672),.clk(gclk));
	jor g4588(.dina(w_n4664_0[0]),.dinb(w_n4610_0[0]),.dout(n4673),.clk(gclk));
	jand g4589(.dina(n4673),.dinb(n4672),.dout(n4674),.clk(gclk));
	jand g4590(.dina(w_n4649_0[0]),.dinb(w_n4616_0[0]),.dout(n4675),.clk(gclk));
	jand g4591(.dina(w_n4650_0[0]),.dinb(w_n4613_0[0]),.dout(n4676),.clk(gclk));
	jor g4592(.dina(n4676),.dinb(n4675),.dout(n4677),.clk(gclk));
	jor g4593(.dina(w_n4624_0[0]),.dinb(w_n4620_0[0]),.dout(n4678),.clk(gclk));
	jand g4594(.dina(w_n4648_0[0]),.dinb(w_n4625_0[0]),.dout(n4679),.clk(gclk));
	jnot g4595(.din(n4679),.dout(n4680),.clk(gclk));
	jand g4596(.dina(n4680),.dinb(n4678),.dout(n4681),.clk(gclk));
	jnot g4597(.din(n4681),.dout(n4682),.clk(gclk));
	jand g4598(.dina(w_n4638_0[0]),.dinb(w_n4628_0[0]),.dout(n4683),.clk(gclk));
	jand g4599(.dina(w_n4647_0[0]),.dinb(w_n4639_0[0]),.dout(n4684),.clk(gclk));
	jor g4600(.dina(n4684),.dinb(n4683),.dout(n4685),.clk(gclk));
	jor g4601(.dina(w_n3927_0[2]),.dinb(w_n2857_2[1]),.dout(n4686),.clk(gclk));
	jor g4602(.dina(w_n3919_2[2]),.dinb(w_n2860_1[2]),.dout(n4687),.clk(gclk));
	jor g4603(.dina(w_n3806_2[1]),.dinb(w_n2865_1[2]),.dout(n4688),.clk(gclk));
	jor g4604(.dina(w_n3600_4[1]),.dinb(w_n2863_2[1]),.dout(n4689),.clk(gclk));
	jand g4605(.dina(n4689),.dinb(n4688),.dout(n4690),.clk(gclk));
	jand g4606(.dina(n4690),.dinb(n4687),.dout(n4691),.clk(gclk));
	jand g4607(.dina(n4691),.dinb(n4686),.dout(n4692),.clk(gclk));
	jxor g4608(.dina(n4692),.dinb(w_n808_5[0]),.dout(n4693),.clk(gclk));
	jxor g4609(.dina(w_n4693_0[1]),.dinb(w_n4685_0[1]),.dout(n4694),.clk(gclk));
	jor g4610(.dina(w_n3320_0[1]),.dinb(w_n3198_2[2]),.dout(n4695),.clk(gclk));
	jor g4611(.dina(w_n3315_3[0]),.dinb(w_n3200_2[0]),.dout(n4696),.clk(gclk));
	jor g4612(.dina(w_n3283_3[0]),.dinb(w_n3204_2[0]),.dout(n4697),.clk(gclk));
	jor g4613(.dina(w_n3284_3[0]),.dinb(w_n3202_2[0]),.dout(n4698),.clk(gclk));
	jand g4614(.dina(n4698),.dinb(n4697),.dout(n4699),.clk(gclk));
	jand g4615(.dina(n4699),.dinb(n4696),.dout(n4700),.clk(gclk));
	jand g4616(.dina(n4700),.dinb(n4695),.dout(n4701),.clk(gclk));
	jxor g4617(.dina(n4701),.dinb(w_n954_12[0]),.dout(n4702),.clk(gclk));
	jnot g4618(.din(n4702),.dout(n4703),.clk(gclk));
	jand g4619(.dina(w_n3176_0[2]),.dinb(w_n954_11[2]),.dout(n4704),.clk(gclk));
	jxor g4620(.dina(w_n4704_0[2]),.dinb(w_n1143_3[1]),.dout(n4705),.clk(gclk));
	jxor g4621(.dina(n4705),.dinb(w_n4571_0[0]),.dout(n4706),.clk(gclk));
	jor g4622(.dina(w_n4637_0[0]),.dinb(w_n4636_0[0]),.dout(n4707),.clk(gclk));
	jand g4623(.dina(w_n2669_1[0]),.dinb(w_n954_11[1]),.dout(n4708),.clk(gclk));
	jand g4624(.dina(n4708),.dinb(w_n2769_1[1]),.dout(n4709),.clk(gclk));
	jnot g4625(.din(n4709),.dout(n4710),.clk(gclk));
	jand g4626(.dina(n4710),.dinb(n4707),.dout(n4711),.clk(gclk));
	jxor g4627(.dina(w_n4711_0[2]),.dinb(w_n4706_0[2]),.dout(n4712),.clk(gclk));
	jxor g4628(.dina(n4712),.dinb(w_n4703_0[1]),.dout(n4713),.clk(gclk));
	jxor g4629(.dina(w_n4713_0[1]),.dinb(w_n4694_0[1]),.dout(n4714),.clk(gclk));
	jxor g4630(.dina(w_n4714_0[1]),.dinb(w_n4682_0[1]),.dout(n4715),.clk(gclk));
	jxor g4631(.dina(w_n4715_0[1]),.dinb(w_n4677_0[1]),.dout(n4716),.clk(gclk));
	jand g4632(.dina(w_n3307_0[2]),.dinb(w_n2736_0[2]),.dout(n4717),.clk(gclk));
	jand g4633(.dina(n4717),.dinb(w_n771_0[2]),.dout(n4718),.clk(gclk));
	jand g4634(.dina(w_n878_0[1]),.dinb(w_n310_0[1]),.dout(n4719),.clk(gclk));
	jand g4635(.dina(n4719),.dinb(w_n479_0[2]),.dout(n4720),.clk(gclk));
	jand g4636(.dina(n4720),.dinb(w_n385_0[1]),.dout(n4721),.clk(gclk));
	jnot g4637(.din(w_n651_0[0]),.dout(n4722),.clk(gclk));
	jand g4638(.dina(w_n3258_0[1]),.dinb(n4722),.dout(n4723),.clk(gclk));
	jand g4639(.dina(n4723),.dinb(n4721),.dout(n4724),.clk(gclk));
	jand g4640(.dina(n4724),.dinb(n4718),.dout(n4725),.clk(gclk));
	jand g4641(.dina(n4725),.dinb(w_n1203_0[0]),.dout(n4726),.clk(gclk));
	jand g4642(.dina(w_n3676_0[0]),.dinb(w_n1013_0[0]),.dout(n4727),.clk(gclk));
	jand g4643(.dina(n4727),.dinb(n4726),.dout(n4728),.clk(gclk));
	jxor g4644(.dina(w_n4728_0[1]),.dinb(w_n4716_0[1]),.dout(n4729),.clk(gclk));
	jxor g4645(.dina(w_n4729_0[1]),.dinb(w_n4674_0[1]),.dout(n4730),.clk(gclk));
	jxor g4646(.dina(w_n4730_0[1]),.dinb(w_n4670_0[1]),.dout(n4731),.clk(gclk));
	jor g4647(.dina(w_n4667_0[0]),.dinb(w_n4666_0[0]),.dout(n4732),.clk(gclk));
	jand g4648(.dina(w_n4732_0[1]),.dinb(w_n4013_7[2]),.dout(n4733),.clk(gclk));
	jxor g4649(.dina(n4733),.dinb(w_n4731_0[1]),.dout(w_dff_A_SP0xCeW41_2),.clk(gclk));
	jand g4650(.dina(w_n4730_0[0]),.dinb(w_n4670_0[0]),.dout(n4735),.clk(gclk));
	jnot g4651(.din(w_n4716_0[0]),.dout(n4736),.clk(gclk));
	jor g4652(.dina(w_n4728_0[0]),.dinb(n4736),.dout(n4737),.clk(gclk));
	jor g4653(.dina(w_n4729_0[0]),.dinb(w_n4674_0[0]),.dout(n4738),.clk(gclk));
	jand g4654(.dina(n4738),.dinb(n4737),.dout(n4739),.clk(gclk));
	jand g4655(.dina(w_n4714_0[0]),.dinb(w_n4682_0[0]),.dout(n4740),.clk(gclk));
	jand g4656(.dina(w_n4715_0[0]),.dinb(w_n4677_0[0]),.dout(n4741),.clk(gclk));
	jor g4657(.dina(n4741),.dinb(n4740),.dout(n4742),.clk(gclk));
	jand g4658(.dina(w_n4693_0[0]),.dinb(w_n4685_0[0]),.dout(n4743),.clk(gclk));
	jand g4659(.dina(w_n4713_0[0]),.dinb(w_n4694_0[0]),.dout(n4744),.clk(gclk));
	jor g4660(.dina(n4744),.dinb(n4743),.dout(n4745),.clk(gclk));
	jand g4661(.dina(w_n4090_0[2]),.dinb(w_n2828_0[2]),.dout(n4746),.clk(gclk));
	jand g4662(.dina(w_n3807_1[2]),.dinb(w_n2848_0[2]),.dout(n4747),.clk(gclk));
	jand g4663(.dina(w_n3920_2[0]),.dinb(w_n2832_0[2]),.dout(n4748),.clk(gclk));
	jor g4664(.dina(n4748),.dinb(n4747),.dout(n4749),.clk(gclk));
	jor g4665(.dina(n4749),.dinb(n4746),.dout(n4750),.clk(gclk));
	jxor g4666(.dina(n4750),.dinb(w_n803_3[0]),.dout(n4751),.clk(gclk));
	jor g4667(.dina(w_n3605_0[1]),.dinb(w_n3198_2[1]),.dout(n4752),.clk(gclk));
	jor g4668(.dina(w_n3600_4[0]),.dinb(w_n3200_1[2]),.dout(n4753),.clk(gclk));
	jor g4669(.dina(w_n3315_2[2]),.dinb(w_n3204_1[2]),.dout(n4754),.clk(gclk));
	jor g4670(.dina(w_n3283_2[2]),.dinb(w_n3202_1[2]),.dout(n4755),.clk(gclk));
	jand g4671(.dina(n4755),.dinb(n4754),.dout(n4756),.clk(gclk));
	jand g4672(.dina(n4756),.dinb(n4753),.dout(n4757),.clk(gclk));
	jand g4673(.dina(n4757),.dinb(n4752),.dout(n4758),.clk(gclk));
	jxor g4674(.dina(n4758),.dinb(w_n820_2[1]),.dout(n4759),.clk(gclk));
	jor g4675(.dina(w_n3284_2[2]),.dinb(w_n820_2[0]),.dout(n4760),.clk(gclk));
	jnot g4676(.din(w_n4704_0[1]),.dout(n4761),.clk(gclk));
	jand g4677(.dina(n4761),.dinb(w_n699_4[1]),.dout(n4762),.clk(gclk));
	jnot g4678(.din(n4762),.dout(n4763),.clk(gclk));
	jand g4679(.dina(w_n4704_0[0]),.dinb(w_n1143_3[0]),.dout(n4764),.clk(gclk));
	jor g4680(.dina(n4764),.dinb(w_n4570_0[0]),.dout(n4765),.clk(gclk));
	jand g4681(.dina(n4765),.dinb(n4763),.dout(n4766),.clk(gclk));
	jxor g4682(.dina(w_n4766_0[1]),.dinb(w_n4760_0[2]),.dout(n4767),.clk(gclk));
	jxor g4683(.dina(w_n4767_0[1]),.dinb(w_n4759_0[1]),.dout(n4768),.clk(gclk));
	jand g4684(.dina(w_n4711_0[1]),.dinb(w_n4706_0[1]),.dout(n4769),.clk(gclk));
	jnot g4685(.din(n4769),.dout(n4770),.clk(gclk));
	jnot g4686(.din(w_n4706_0[0]),.dout(n4771),.clk(gclk));
	jnot g4687(.din(w_n4711_0[0]),.dout(n4772),.clk(gclk));
	jand g4688(.dina(n4772),.dinb(n4771),.dout(n4773),.clk(gclk));
	jor g4689(.dina(n4773),.dinb(w_n4703_0[0]),.dout(n4774),.clk(gclk));
	jand g4690(.dina(n4774),.dinb(n4770),.dout(n4775),.clk(gclk));
	jxor g4691(.dina(w_n4775_0[1]),.dinb(w_n4768_0[1]),.dout(n4776),.clk(gclk));
	jxor g4692(.dina(w_n4776_0[1]),.dinb(w_n4751_0[1]),.dout(n4777),.clk(gclk));
	jxor g4693(.dina(w_n4777_0[1]),.dinb(w_n4745_0[1]),.dout(n4778),.clk(gclk));
	jxor g4694(.dina(w_n4778_0[1]),.dinb(w_n4742_0[1]),.dout(n4779),.clk(gclk));
	jand g4695(.dina(w_n935_1[1]),.dinb(w_n511_0[1]),.dout(n4780),.clk(gclk));
	jand g4696(.dina(n4780),.dinb(w_n677_0[0]),.dout(n4781),.clk(gclk));
	jand g4697(.dina(n4781),.dinb(w_n746_0[0]),.dout(n4782),.clk(gclk));
	jand g4698(.dina(n4782),.dinb(w_n784_0[0]),.dout(n4783),.clk(gclk));
	jand g4699(.dina(n4783),.dinb(w_n3794_0[0]),.dout(n4784),.clk(gclk));
	jand g4700(.dina(n4784),.dinb(w_n1006_0[0]),.dout(n4785),.clk(gclk));
	jxor g4701(.dina(w_n4785_0[1]),.dinb(w_n4779_0[1]),.dout(n4786),.clk(gclk));
	jxor g4702(.dina(w_n4786_0[1]),.dinb(w_n4739_0[1]),.dout(n4787),.clk(gclk));
	jxor g4703(.dina(w_n4787_0[1]),.dinb(w_n4735_0[1]),.dout(n4788),.clk(gclk));
	jor g4704(.dina(w_n4732_0[0]),.dinb(w_n4731_0[0]),.dout(n4789),.clk(gclk));
	jand g4705(.dina(w_n4789_0[1]),.dinb(w_n4013_7[1]),.dout(n4790),.clk(gclk));
	jxor g4706(.dina(n4790),.dinb(w_n4788_0[1]),.dout(w_dff_A_gP8OwZoN2_2),.clk(gclk));
	jand g4707(.dina(w_n4787_0[0]),.dinb(w_n4735_0[0]),.dout(n4792),.clk(gclk));
	jnot g4708(.din(w_n4779_0[0]),.dout(n4793),.clk(gclk));
	jor g4709(.dina(w_n4785_0[0]),.dinb(n4793),.dout(n4794),.clk(gclk));
	jor g4710(.dina(w_n4786_0[0]),.dinb(w_n4739_0[0]),.dout(n4795),.clk(gclk));
	jand g4711(.dina(n4795),.dinb(n4794),.dout(n4796),.clk(gclk));
	jand g4712(.dina(w_n4777_0[0]),.dinb(w_n4745_0[0]),.dout(n4797),.clk(gclk));
	jand g4713(.dina(w_n4778_0[0]),.dinb(w_n4742_0[0]),.dout(n4798),.clk(gclk));
	jor g4714(.dina(n4798),.dinb(n4797),.dout(n4799),.clk(gclk));
	jand g4715(.dina(w_n4775_0[0]),.dinb(w_n4768_0[0]),.dout(n4800),.clk(gclk));
	jand g4716(.dina(w_n4776_0[0]),.dinb(w_n4751_0[0]),.dout(n4801),.clk(gclk));
	jor g4717(.dina(n4801),.dinb(n4800),.dout(n4802),.clk(gclk));
	jand g4718(.dina(w_n4766_0[0]),.dinb(w_n4760_0[1]),.dout(n4803),.clk(gclk));
	jand g4719(.dina(w_n4767_0[0]),.dinb(w_n4759_0[0]),.dout(n4804),.clk(gclk));
	jor g4720(.dina(n4804),.dinb(n4803),.dout(n4805),.clk(gclk));
	jnot g4721(.din(n4805),.dout(n4806),.clk(gclk));
	jand g4722(.dina(w_n3299_0[0]),.dinb(w_n954_11[0]),.dout(n4807),.clk(gclk));
	jxor g4723(.dina(w_n4807_0[1]),.dinb(w_n4806_0[1]),.dout(n4808),.clk(gclk));
	jor g4724(.dina(w_n3811_0[1]),.dinb(w_n3198_2[0]),.dout(n4809),.clk(gclk));
	jor g4725(.dina(w_n3806_2[0]),.dinb(w_n3200_1[1]),.dout(n4810),.clk(gclk));
	jor g4726(.dina(w_n3600_3[2]),.dinb(w_n3204_1[1]),.dout(n4811),.clk(gclk));
	jor g4727(.dina(w_n3315_2[1]),.dinb(w_n3202_1[1]),.dout(n4812),.clk(gclk));
	jand g4728(.dina(n4812),.dinb(n4811),.dout(n4813),.clk(gclk));
	jand g4729(.dina(n4813),.dinb(n4810),.dout(n4814),.clk(gclk));
	jand g4730(.dina(n4814),.dinb(n4809),.dout(n4815),.clk(gclk));
	jxor g4731(.dina(n4815),.dinb(w_n954_10[2]),.dout(n4816),.clk(gclk));
	jor g4732(.dina(w_n4136_0[2]),.dinb(w_n2857_2[0]),.dout(n4817),.clk(gclk));
	jand g4733(.dina(n4817),.dinb(w_n2863_2[0]),.dout(n4818),.clk(gclk));
	jor g4734(.dina(n4818),.dinb(w_n3919_2[1]),.dout(n4819),.clk(gclk));
	jxor g4735(.dina(n4819),.dinb(w_n803_2[2]),.dout(n4820),.clk(gclk));
	jxor g4736(.dina(w_n4820_0[1]),.dinb(w_n4816_0[1]),.dout(n4821),.clk(gclk));
	jxor g4737(.dina(w_n4821_0[1]),.dinb(w_n4808_0[1]),.dout(n4822),.clk(gclk));
	jxor g4738(.dina(w_n4822_0[1]),.dinb(w_n4802_0[1]),.dout(n4823),.clk(gclk));
	jxor g4739(.dina(w_n4823_0[1]),.dinb(w_n4799_0[1]),.dout(n4824),.clk(gclk));
	jand g4740(.dina(w_n421_1[0]),.dinb(w_n254_1[0]),.dout(n4825),.clk(gclk));
	jand g4741(.dina(n4825),.dinb(w_n372_0[2]),.dout(n4826),.clk(gclk));
	jand g4742(.dina(n4826),.dinb(w_n2456_0[1]),.dout(n4827),.clk(gclk));
	jand g4743(.dina(n4827),.dinb(w_n565_0[1]),.dout(n4828),.clk(gclk));
	jand g4744(.dina(w_n668_0[2]),.dinb(w_n420_0[2]),.dout(n4829),.clk(gclk));
	jand g4745(.dina(w_n594_0[2]),.dinb(w_n868_0[1]),.dout(n4830),.clk(gclk));
	jand g4746(.dina(n4830),.dinb(w_n277_1[2]),.dout(n4831),.clk(gclk));
	jand g4747(.dina(n4831),.dinb(n4829),.dout(n4832),.clk(gclk));
	jand g4748(.dina(w_n4832_0[1]),.dinb(w_n4106_0[0]),.dout(n4833),.clk(gclk));
	jand g4749(.dina(n4833),.dinb(n4828),.dout(n4834),.clk(gclk));
	jand g4750(.dina(n4834),.dinb(w_n2449_0[0]),.dout(n4835),.clk(gclk));
	jand g4751(.dina(n4835),.dinb(w_n2313_0[0]),.dout(n4836),.clk(gclk));
	jxor g4752(.dina(w_n4836_0[1]),.dinb(w_n4824_0[1]),.dout(n4837),.clk(gclk));
	jxor g4753(.dina(w_n4837_0[1]),.dinb(w_n4796_0[1]),.dout(n4838),.clk(gclk));
	jxor g4754(.dina(w_n4838_0[1]),.dinb(w_n4792_0[1]),.dout(n4839),.clk(gclk));
	jor g4755(.dina(w_n4789_0[0]),.dinb(w_n4788_0[0]),.dout(n4840),.clk(gclk));
	jand g4756(.dina(w_n4840_0[1]),.dinb(w_n4013_7[0]),.dout(n4841),.clk(gclk));
	jxor g4757(.dina(n4841),.dinb(w_n4839_0[1]),.dout(w_dff_A_5LHruE6g9_2),.clk(gclk));
	jand g4758(.dina(w_n4838_0[0]),.dinb(w_n4792_0[0]),.dout(n4843),.clk(gclk));
	jnot g4759(.din(w_n4824_0[0]),.dout(n4844),.clk(gclk));
	jor g4760(.dina(w_n4836_0[0]),.dinb(n4844),.dout(n4845),.clk(gclk));
	jor g4761(.dina(w_n4837_0[0]),.dinb(w_n4796_0[0]),.dout(n4846),.clk(gclk));
	jand g4762(.dina(n4846),.dinb(n4845),.dout(n4847),.clk(gclk));
	jand g4763(.dina(w_n4822_0[0]),.dinb(w_n4802_0[0]),.dout(n4848),.clk(gclk));
	jand g4764(.dina(w_n4823_0[0]),.dinb(w_n4799_0[0]),.dout(n4849),.clk(gclk));
	jor g4765(.dina(n4849),.dinb(n4848),.dout(n4850),.clk(gclk));
	jor g4766(.dina(w_n4820_0[0]),.dinb(w_n4816_0[0]),.dout(n4851),.clk(gclk));
	jand g4767(.dina(w_n4821_0[0]),.dinb(w_n4808_0[0]),.dout(n4852),.clk(gclk));
	jnot g4768(.din(n4852),.dout(n4853),.clk(gclk));
	jand g4769(.dina(n4853),.dinb(n4851),.dout(n4854),.clk(gclk));
	jnot g4770(.din(n4854),.dout(n4855),.clk(gclk));
	jor g4771(.dina(w_n4807_0[0]),.dinb(w_n4806_0[0]),.dout(n4856),.clk(gclk));
	jor g4772(.dina(w_n4760_0[0]),.dinb(w_n3302_0[1]),.dout(n4857),.clk(gclk));
	jand g4773(.dina(n4857),.dinb(n4856),.dout(n4858),.clk(gclk));
	jnot g4774(.din(n4858),.dout(n4859),.clk(gclk));
	jor g4775(.dina(w_n3927_0[1]),.dinb(w_n3198_1[2]),.dout(n4860),.clk(gclk));
	jor g4776(.dina(w_n3919_2[0]),.dinb(w_n3200_1[0]),.dout(n4861),.clk(gclk));
	jor g4777(.dina(w_n3806_1[2]),.dinb(w_n3204_1[0]),.dout(n4862),.clk(gclk));
	jor g4778(.dina(w_n3600_3[1]),.dinb(w_n3202_1[0]),.dout(n4863),.clk(gclk));
	jand g4779(.dina(n4863),.dinb(n4862),.dout(n4864),.clk(gclk));
	jand g4780(.dina(n4864),.dinb(n4861),.dout(n4865),.clk(gclk));
	jand g4781(.dina(n4865),.dinb(n4860),.dout(n4866),.clk(gclk));
	jxor g4782(.dina(n4866),.dinb(w_n954_10[1]),.dout(n4867),.clk(gclk));
	jnot g4783(.din(n4867),.dout(n4868),.clk(gclk));
	jand g4784(.dina(w_n3302_0[0]),.dinb(w_n954_10[0]),.dout(n4869),.clk(gclk));
	jxor g4785(.dina(w_n4869_0[1]),.dinb(w_n808_4[2]),.dout(n4870),.clk(gclk));
	jand g4786(.dina(w_n3316_0[0]),.dinb(w_n954_9[2]),.dout(n4871),.clk(gclk));
	jxor g4787(.dina(w_n4871_0[1]),.dinb(w_n4870_0[1]),.dout(n4872),.clk(gclk));
	jxor g4788(.dina(w_n4872_0[1]),.dinb(w_n4868_0[1]),.dout(n4873),.clk(gclk));
	jxor g4789(.dina(w_n4873_0[1]),.dinb(w_n4859_0[1]),.dout(n4874),.clk(gclk));
	jxor g4790(.dina(w_n4874_0[1]),.dinb(w_n4855_0[1]),.dout(n4875),.clk(gclk));
	jxor g4791(.dina(w_n4875_0[1]),.dinb(w_n4850_0[1]),.dout(n4876),.clk(gclk));
	jand g4792(.dina(w_n592_1[0]),.dinb(w_n323_1[1]),.dout(n4877),.clk(gclk));
	jand g4793(.dina(w_n665_0[2]),.dinb(w_n561_0[2]),.dout(n4878),.clk(gclk));
	jand g4794(.dina(n4878),.dinb(w_n264_0[2]),.dout(n4879),.clk(gclk));
	jand g4795(.dina(n4879),.dinb(n4877),.dout(n4880),.clk(gclk));
	jand g4796(.dina(w_n662_0[2]),.dinb(w_n463_1[0]),.dout(n4881),.clk(gclk));
	jand g4797(.dina(n4881),.dinb(w_n619_0[2]),.dout(n4882),.clk(gclk));
	jand g4798(.dina(w_n822_0[2]),.dinb(w_n413_0[0]),.dout(n4883),.clk(gclk));
	jand g4799(.dina(n4883),.dinb(n4882),.dout(n4884),.clk(gclk));
	jand g4800(.dina(w_n749_0[2]),.dinb(w_n343_0[2]),.dout(n4885),.clk(gclk));
	jand g4801(.dina(n4885),.dinb(w_n882_0[2]),.dout(n4886),.clk(gclk));
	jand g4802(.dina(n4886),.dinb(w_n4000_0[0]),.dout(n4887),.clk(gclk));
	jand g4803(.dina(n4887),.dinb(n4884),.dout(n4888),.clk(gclk));
	jand g4804(.dina(n4888),.dinb(w_n4880_0[1]),.dout(n4889),.clk(gclk));
	jand g4805(.dina(n4889),.dinb(w_n1231_0[0]),.dout(n4890),.clk(gclk));
	jand g4806(.dina(w_n3693_0[0]),.dinb(w_n2665_0[0]),.dout(n4891),.clk(gclk));
	jand g4807(.dina(n4891),.dinb(n4890),.dout(n4892),.clk(gclk));
	jxor g4808(.dina(w_n4892_0[1]),.dinb(w_n4876_0[1]),.dout(n4893),.clk(gclk));
	jxor g4809(.dina(w_n4893_0[1]),.dinb(w_n4847_0[1]),.dout(n4894),.clk(gclk));
	jxor g4810(.dina(w_n4894_0[1]),.dinb(w_n4843_0[1]),.dout(n4895),.clk(gclk));
	jor g4811(.dina(w_n4840_0[0]),.dinb(w_n4839_0[0]),.dout(n4896),.clk(gclk));
	jand g4812(.dina(w_n4896_0[1]),.dinb(w_n4013_6[2]),.dout(n4897),.clk(gclk));
	jxor g4813(.dina(n4897),.dinb(w_n4895_0[1]),.dout(w_dff_A_oxEVAVgt4_2),.clk(gclk));
	jand g4814(.dina(w_n4894_0[0]),.dinb(w_n4843_0[0]),.dout(n4899),.clk(gclk));
	jnot g4815(.din(w_n4876_0[0]),.dout(n4900),.clk(gclk));
	jor g4816(.dina(w_n4892_0[0]),.dinb(n4900),.dout(n4901),.clk(gclk));
	jor g4817(.dina(w_n4893_0[0]),.dinb(w_n4847_0[0]),.dout(n4902),.clk(gclk));
	jand g4818(.dina(n4902),.dinb(n4901),.dout(n4903),.clk(gclk));
	jand g4819(.dina(w_n4874_0[0]),.dinb(w_n4855_0[0]),.dout(n4904),.clk(gclk));
	jand g4820(.dina(w_n4875_0[0]),.dinb(w_n4850_0[0]),.dout(n4905),.clk(gclk));
	jor g4821(.dina(n4905),.dinb(n4904),.dout(n4906),.clk(gclk));
	jand g4822(.dina(w_n4872_0[0]),.dinb(w_n4868_0[0]),.dout(n4907),.clk(gclk));
	jand g4823(.dina(w_n4873_0[0]),.dinb(w_n4859_0[0]),.dout(n4908),.clk(gclk));
	jor g4824(.dina(n4908),.dinb(n4907),.dout(n4909),.clk(gclk));
	jand g4825(.dina(w_n4090_0[1]),.dinb(w_n2883_1[1]),.dout(n4910),.clk(gclk));
	jand g4826(.dina(w_n3807_1[1]),.dinb(w_n2995_1[2]),.dout(n4911),.clk(gclk));
	jand g4827(.dina(w_n3920_1[2]),.dinb(w_n2887_1[1]),.dout(n4912),.clk(gclk));
	jor g4828(.dina(n4912),.dinb(n4911),.dout(n4913),.clk(gclk));
	jor g4829(.dina(n4913),.dinb(n4910),.dout(n4914),.clk(gclk));
	jxor g4830(.dina(n4914),.dinb(w_n954_9[1]),.dout(n4915),.clk(gclk));
	jand g4831(.dina(w_n3601_0[2]),.dinb(w_n954_9[0]),.dout(n4916),.clk(gclk));
	jnot g4832(.din(n4916),.dout(n4917),.clk(gclk));
	jand g4833(.dina(w_n4869_0[0]),.dinb(w_n808_4[1]),.dout(n4918),.clk(gclk));
	jand g4834(.dina(w_n4871_0[0]),.dinb(w_n4870_0[0]),.dout(n4919),.clk(gclk));
	jor g4835(.dina(n4919),.dinb(n4918),.dout(n4920),.clk(gclk));
	jxor g4836(.dina(w_n4920_0[1]),.dinb(w_n4917_0[1]),.dout(n4921),.clk(gclk));
	jxor g4837(.dina(w_n4921_0[1]),.dinb(w_n4915_0[1]),.dout(n4922),.clk(gclk));
	jxor g4838(.dina(w_n4922_0[1]),.dinb(w_n4909_0[1]),.dout(n4923),.clk(gclk));
	jxor g4839(.dina(w_n4923_0[1]),.dinb(w_n4906_0[1]),.dout(n4924),.clk(gclk));
	jand g4840(.dina(w_n2456_0[0]),.dinb(w_n712_0[0]),.dout(n4925),.clk(gclk));
	jand g4841(.dina(w_n3307_0[1]),.dinb(w_n2521_0[1]),.dout(n4926),.clk(gclk));
	jand g4842(.dina(n4926),.dinb(n4925),.dout(n4927),.clk(gclk));
	jand g4843(.dina(w_n749_0[1]),.dinb(w_n222_0[2]),.dout(n4928),.clk(gclk));
	jand g4844(.dina(n4928),.dinb(w_n918_0[2]),.dout(n4929),.clk(gclk));
	jand g4845(.dina(w_n935_1[0]),.dinb(w_n251_1[1]),.dout(n4930),.clk(gclk));
	jand g4846(.dina(w_n358_0[2]),.dinb(w_n130_0[2]),.dout(n4931),.clk(gclk));
	jand g4847(.dina(w_n4931_0[1]),.dinb(n4930),.dout(n4932),.clk(gclk));
	jand g4848(.dina(n4932),.dinb(n4929),.dout(n4933),.clk(gclk));
	jand g4849(.dina(n4933),.dinb(n4927),.dout(n4934),.clk(gclk));
	jand g4850(.dina(n4934),.dinb(w_n622_0[1]),.dout(n4935),.clk(gclk));
	jnot g4851(.din(w_n1669_0[0]),.dout(n4936),.clk(gclk));
	jand g4852(.dina(n4936),.dinb(w_n675_0[0]),.dout(n4937),.clk(gclk));
	jand g4853(.dina(n4937),.dinb(n4935),.dout(n4938),.clk(gclk));
	jand g4854(.dina(n4938),.dinb(w_n2575_0[0]),.dout(n4939),.clk(gclk));
	jxor g4855(.dina(w_n4939_0[1]),.dinb(w_n4924_0[1]),.dout(n4940),.clk(gclk));
	jxor g4856(.dina(w_n4940_0[1]),.dinb(w_n4903_0[1]),.dout(n4941),.clk(gclk));
	jxor g4857(.dina(w_n4941_0[1]),.dinb(w_n4899_0[1]),.dout(n4942),.clk(gclk));
	jor g4858(.dina(w_n4896_0[0]),.dinb(w_n4895_0[0]),.dout(n4943),.clk(gclk));
	jand g4859(.dina(w_n4943_0[1]),.dinb(w_n4013_6[1]),.dout(n4944),.clk(gclk));
	jxor g4860(.dina(n4944),.dinb(w_n4942_0[1]),.dout(w_dff_A_CHdzBFmi0_2),.clk(gclk));
	jand g4861(.dina(w_n4941_0[0]),.dinb(w_n4899_0[0]),.dout(n4946),.clk(gclk));
	jnot g4862(.din(w_n4924_0[0]),.dout(n4947),.clk(gclk));
	jor g4863(.dina(w_n4939_0[0]),.dinb(n4947),.dout(n4948),.clk(gclk));
	jor g4864(.dina(w_n4940_0[0]),.dinb(w_n4903_0[0]),.dout(n4949),.clk(gclk));
	jand g4865(.dina(n4949),.dinb(n4948),.dout(n4950),.clk(gclk));
	jand g4866(.dina(w_n4920_0[0]),.dinb(w_n4917_0[0]),.dout(n4951),.clk(gclk));
	jand g4867(.dina(w_n4921_0[0]),.dinb(w_n4915_0[0]),.dout(n4952),.clk(gclk));
	jor g4868(.dina(n4952),.dinb(n4951),.dout(n4953),.clk(gclk));
	jnot g4869(.din(w_n4136_0[1]),.dout(n4954),.clk(gclk));
	jand g4870(.dina(n4954),.dinb(w_n2883_1[0]),.dout(n4955),.clk(gclk));
	jor g4871(.dina(n4955),.dinb(w_n2995_1[1]),.dout(n4956),.clk(gclk));
	jand g4872(.dina(n4956),.dinb(w_n3920_1[1]),.dout(n4957),.clk(gclk));
	jxor g4873(.dina(w_n4957_0[1]),.dinb(w_n820_1[2]),.dout(n4958),.clk(gclk));
	jand g4874(.dina(w_n3900_0[0]),.dinb(w_n954_8[2]),.dout(n4959),.clk(gclk));
	jor g4875(.dina(w_n4959_0[1]),.dinb(n4958),.dout(n4960),.clk(gclk));
	jnot g4876(.din(w_n4957_0[0]),.dout(n4961),.clk(gclk));
	jnot g4877(.din(w_n4959_0[0]),.dout(n4962),.clk(gclk));
	jor g4878(.dina(n4962),.dinb(n4961),.dout(n4963),.clk(gclk));
	jand g4879(.dina(n4963),.dinb(w_n4960_0[1]),.dout(n4964),.clk(gclk));
	jxor g4880(.dina(w_n4964_0[1]),.dinb(w_n4953_0[1]),.dout(n4965),.clk(gclk));
	jand g4881(.dina(w_n4922_0[0]),.dinb(w_n4909_0[0]),.dout(n4966),.clk(gclk));
	jand g4882(.dina(w_n4923_0[0]),.dinb(w_n4906_0[0]),.dout(n4967),.clk(gclk));
	jor g4883(.dina(n4967),.dinb(n4966),.dout(n4968),.clk(gclk));
	jxor g4884(.dina(w_n4968_0[1]),.dinb(w_n4965_0[1]),.dout(n4969),.clk(gclk));
	jand g4885(.dina(w_n614_0[2]),.dinb(w_n436_0[2]),.dout(n4970),.clk(gclk));
	jand g4886(.dina(n4970),.dinb(w_n303_1[1]),.dout(n4971),.clk(gclk));
	jand g4887(.dina(n4971),.dinb(w_n1299_0[0]),.dout(n4972),.clk(gclk));
	jand g4888(.dina(w_n387_0[1]),.dinb(w_n383_0[2]),.dout(n4973),.clk(gclk));
	jand g4889(.dina(n4973),.dinb(w_n4931_0[0]),.dout(n4974),.clk(gclk));
	jand g4890(.dina(w_n645_0[2]),.dinb(w_n624_0[2]),.dout(n4975),.clk(gclk));
	jand g4891(.dina(n4975),.dinb(w_n992_0[1]),.dout(n4976),.clk(gclk));
	jand g4892(.dina(n4976),.dinb(w_n680_0[1]),.dout(n4977),.clk(gclk));
	jand g4893(.dina(n4977),.dinb(n4974),.dout(n4978),.clk(gclk));
	jand g4894(.dina(n4978),.dinb(w_n4832_0[0]),.dout(n4979),.clk(gclk));
	jand g4895(.dina(n4979),.dinb(w_n1240_0[0]),.dout(n4980),.clk(gclk));
	jand g4896(.dina(n4980),.dinb(w_n2461_0[0]),.dout(n4981),.clk(gclk));
	jand g4897(.dina(n4981),.dinb(w_n4972_0[1]),.dout(n4982),.clk(gclk));
	jxor g4898(.dina(w_n4982_0[1]),.dinb(w_n4969_0[1]),.dout(n4983),.clk(gclk));
	jxor g4899(.dina(w_n4983_0[1]),.dinb(w_n4950_0[1]),.dout(n4984),.clk(gclk));
	jxor g4900(.dina(w_n4984_0[1]),.dinb(w_n4946_0[1]),.dout(n4985),.clk(gclk));
	jor g4901(.dina(w_n4943_0[0]),.dinb(w_n4942_0[0]),.dout(n4986),.clk(gclk));
	jand g4902(.dina(w_n4986_0[1]),.dinb(w_n4013_6[0]),.dout(n4987),.clk(gclk));
	jxor g4903(.dina(n4987),.dinb(w_n4985_0[1]),.dout(w_dff_A_rLUmXsuL3_2),.clk(gclk));
	jand g4904(.dina(w_n4984_0[0]),.dinb(w_n4946_0[0]),.dout(n4989),.clk(gclk));
	jnot g4905(.din(w_n4969_0[0]),.dout(n4990),.clk(gclk));
	jor g4906(.dina(w_n4982_0[0]),.dinb(n4990),.dout(n4991),.clk(gclk));
	jor g4907(.dina(w_n4983_0[0]),.dinb(w_n4950_0[0]),.dout(n4992),.clk(gclk));
	jand g4908(.dina(n4992),.dinb(n4991),.dout(n4993),.clk(gclk));
	jnot g4909(.din(w_n4993_0[1]),.dout(n4994),.clk(gclk));
	jand g4910(.dina(w_n477_0[2]),.dinb(w_n291_0[2]),.dout(n4995),.clk(gclk));
	jand g4911(.dina(n4995),.dinb(w_n710_1[0]),.dout(n4996),.clk(gclk));
	jand g4912(.dina(w_n543_0[1]),.dinb(w_n384_0[1]),.dout(n4997),.clk(gclk));
	jand g4913(.dina(n4997),.dinb(n4996),.dout(n4998),.clk(gclk));
	jand g4914(.dina(n4998),.dinb(w_n2334_0[0]),.dout(n4999),.clk(gclk));
	jand g4915(.dina(w_n4880_0[0]),.dinb(w_n3620_0[0]),.dout(n5000),.clk(gclk));
	jand g4916(.dina(n5000),.dinb(n4999),.dout(n5001),.clk(gclk));
	jand g4917(.dina(n5001),.dinb(w_n3696_0[0]),.dout(n5002),.clk(gclk));
	jand g4918(.dina(n5002),.dinb(w_n2382_0[0]),.dout(n5003),.clk(gclk));
	jand g4919(.dina(w_n3600_3[0]),.dinb(w_n954_8[1]),.dout(n5004),.clk(gclk));
	jand g4920(.dina(n5004),.dinb(w_n3807_1[0]),.dout(n5005),.clk(gclk));
	jnot g4921(.din(n5005),.dout(n5006),.clk(gclk));
	jand g4922(.dina(n5006),.dinb(w_n4960_0[0]),.dout(n5007),.clk(gclk));
	jnot g4923(.din(w_n5007_0[1]),.dout(n5008),.clk(gclk));
	jand g4924(.dina(w_n4964_0[0]),.dinb(w_n4953_0[0]),.dout(n5009),.clk(gclk));
	jand g4925(.dina(w_n4968_0[0]),.dinb(w_n4965_0[0]),.dout(n5010),.clk(gclk));
	jor g4926(.dina(n5010),.dinb(n5009),.dout(n5011),.clk(gclk));
	jor g4927(.dina(w_n3920_1[0]),.dinb(w_n3600_2[2]),.dout(n5012),.clk(gclk));
	jor g4928(.dina(w_n3919_1[2]),.dinb(w_n3601_0[1]),.dout(n5013),.clk(gclk));
	jand g4929(.dina(n5013),.dinb(w_n954_8[0]),.dout(n5014),.clk(gclk));
	jand g4930(.dina(n5014),.dinb(n5012),.dout(n5015),.clk(gclk));
	jxor g4931(.dina(n5015),.dinb(n5011),.dout(n5016),.clk(gclk));
	jxor g4932(.dina(w_n5016_0[1]),.dinb(n5008),.dout(n5017),.clk(gclk));
	jxor g4933(.dina(w_n5017_0[1]),.dinb(w_n5003_0[2]),.dout(n5018),.clk(gclk));
	jxor g4934(.dina(w_n5018_0[1]),.dinb(w_n4994_0[1]),.dout(n5019),.clk(gclk));
	jxor g4935(.dina(w_n5019_0[1]),.dinb(w_n4989_0[1]),.dout(n5020),.clk(gclk));
	jor g4936(.dina(w_n4986_0[0]),.dinb(w_n4985_0[0]),.dout(n5021),.clk(gclk));
	jand g4937(.dina(w_n5021_0[1]),.dinb(w_n4013_5[2]),.dout(n5022),.clk(gclk));
	jxor g4938(.dina(w_dff_B_eZEzychJ4_0),.dinb(w_n5020_0[1]),.dout(w_dff_A_J2WpamXl7_2),.clk(gclk));
	jor g4939(.dina(w_n5021_0[0]),.dinb(w_n5020_0[0]),.dout(n5024),.clk(gclk));
	jand g4940(.dina(w_n5024_0[2]),.dinb(w_n4013_5[1]),.dout(n5025),.clk(gclk));
	jand g4941(.dina(w_n5019_0[0]),.dinb(w_n4989_0[0]),.dout(n5026),.clk(gclk));
	jor g4942(.dina(w_n5017_0[0]),.dinb(w_n5003_0[1]),.dout(n5027),.clk(gclk));
	jxor g4943(.dina(w_n5016_0[0]),.dinb(w_n5007_0[0]),.dout(n5028),.clk(gclk));
	jxor g4944(.dina(n5028),.dinb(w_n5003_0[0]),.dout(n5029),.clk(gclk));
	jor g4945(.dina(n5029),.dinb(w_n4993_0[0]),.dout(n5030),.clk(gclk));
	jand g4946(.dina(n5030),.dinb(w_n5027_0[1]),.dout(n5031),.clk(gclk));
	jand g4947(.dina(w_n461_0[2]),.dinb(w_n372_0[1]),.dout(n5032),.clk(gclk));
	jand g4948(.dina(n5032),.dinb(w_n619_0[1]),.dout(n5033),.clk(gclk));
	jand g4949(.dina(w_n2736_0[1]),.dinb(w_n507_0[1]),.dout(n5034),.clk(gclk));
	jand g4950(.dina(n5034),.dinb(n5033),.dout(n5035),.clk(gclk));
	jand g4951(.dina(w_n365_0[1]),.dinb(w_n277_1[1]),.dout(n5036),.clk(gclk));
	jand g4952(.dina(n5036),.dinb(w_n422_0[2]),.dout(n5037),.clk(gclk));
	jand g4953(.dina(n5037),.dinb(w_n443_0[0]),.dout(n5038),.clk(gclk));
	jand g4954(.dina(n5038),.dinb(n5035),.dout(n5039),.clk(gclk));
	jand g4955(.dina(n5039),.dinb(w_n824_0[0]),.dout(n5040),.clk(gclk));
	jand g4956(.dina(n5040),.dinb(w_n3256_0[0]),.dout(n5041),.clk(gclk));
	jand g4957(.dina(n5041),.dinb(w_n860_0[0]),.dout(n5042),.clk(gclk));
	jxor g4958(.dina(w_n5042_1[1]),.dinb(w_n5031_0[1]),.dout(n5043),.clk(gclk));
	jxor g4959(.dina(w_n5043_0[2]),.dinb(w_n5026_0[2]),.dout(n5044),.clk(gclk));
	jxor g4960(.dina(w_n5044_0[1]),.dinb(n5025),.dout(w_dff_A_k0YYIuNo5_2),.clk(gclk));
	jnot g4961(.din(w_n4013_5[0]),.dout(n5046),.clk(gclk));
	jnot g4962(.din(w_n5024_0[1]),.dout(n5047),.clk(gclk));
	jnot g4963(.din(w_n5026_0[1]),.dout(n5048),.clk(gclk));
	jxor g4964(.dina(w_n5043_0[1]),.dinb(w_n5048_0[1]),.dout(n5049),.clk(gclk));
	jand g4965(.dina(n5049),.dinb(n5047),.dout(n5050),.clk(gclk));
	jor g4966(.dina(w_n5050_0[1]),.dinb(w_n5046_0[1]),.dout(n5051),.clk(gclk));
	jnot g4967(.din(w_n5027_0[0]),.dout(n5052),.clk(gclk));
	jand g4968(.dina(w_n5018_0[0]),.dinb(w_n4994_0[0]),.dout(n5053),.clk(gclk));
	jor g4969(.dina(n5053),.dinb(n5052),.dout(n5054),.clk(gclk));
	jnot g4970(.din(w_n5042_1[0]),.dout(n5055),.clk(gclk));
	jand g4971(.dina(n5055),.dinb(w_n5054_0[1]),.dout(n5056),.clk(gclk));
	jand g4972(.dina(w_n5043_0[0]),.dinb(w_n5026_0[0]),.dout(n5057),.clk(gclk));
	jor g4973(.dina(w_n5057_0[1]),.dinb(w_n5056_0[1]),.dout(n5058),.clk(gclk));
	jand g4974(.dina(w_n277_1[0]),.dinb(w_n251_1[0]),.dout(n5059),.clk(gclk));
	jand g4975(.dina(n5059),.dinb(w_n368_0[2]),.dout(n5060),.clk(gclk));
	jand g4976(.dina(n5060),.dinb(w_n2396_0[0]),.dout(n5061),.clk(gclk));
	jand g4977(.dina(w_n999_0[0]),.dinb(w_n611_0[1]),.dout(n5062),.clk(gclk));
	jand g4978(.dina(n5062),.dinb(n5061),.dout(n5063),.clk(gclk));
	jand g4979(.dina(w_n2658_0[0]),.dinb(w_n1218_0[0]),.dout(n5064),.clk(gclk));
	jand g4980(.dina(n5064),.dinb(n5063),.dout(n5065),.clk(gclk));
	jand g4981(.dina(n5065),.dinb(w_n1307_0[0]),.dout(n5066),.clk(gclk));
	jand g4982(.dina(n5066),.dinb(w_n3663_0[0]),.dout(n5067),.clk(gclk));
	jand g4983(.dina(n5067),.dinb(w_n834_0[0]),.dout(n5068),.clk(gclk));
	jxor g4984(.dina(w_n5068_1[1]),.dinb(w_n5058_0[1]),.dout(n5069),.clk(gclk));
	jxor g4985(.dina(w_n5069_0[1]),.dinb(n5051),.dout(w_dff_A_0nVz4h2P4_2),.clk(gclk));
	jor g4986(.dina(w_n5042_0[2]),.dinb(w_n5031_0[0]),.dout(n5071),.clk(gclk));
	jor g4987(.dina(w_n5068_1[0]),.dinb(n5071),.dout(n5072),.clk(gclk));
	jand g4988(.dina(w_n3257_0[0]),.dinb(w_n681_0[0]),.dout(n5073),.clk(gclk));
	jand g4989(.dina(n5073),.dinb(w_n987_0[1]),.dout(n5074),.clk(gclk));
	jand g4990(.dina(w_n768_0[2]),.dinb(w_n157_0[1]),.dout(n5075),.clk(gclk));
	jand g4991(.dina(n5075),.dinb(w_n1209_0[1]),.dout(n5076),.clk(gclk));
	jand g4992(.dina(n5076),.dinb(w_n4357_0[0]),.dout(n5077),.clk(gclk));
	jand g4993(.dina(n5077),.dinb(n5074),.dout(n5078),.clk(gclk));
	jand g4994(.dina(n5078),.dinb(w_n3159_0[0]),.dout(n5079),.clk(gclk));
	jand g4995(.dina(n5079),.dinb(w_n1175_0[0]),.dout(n5080),.clk(gclk));
	jand g4996(.dina(n5080),.dinb(w_n4972_0[0]),.dout(n5081),.clk(gclk));
	jxor g4997(.dina(w_n5081_0[2]),.dinb(n5072),.dout(n5082),.clk(gclk));
	jnot g4998(.din(w_n5068_0[2]),.dout(n5083),.clk(gclk));
	jand g4999(.dina(w_n5083_0[2]),.dinb(w_n5057_0[0]),.dout(n5084),.clk(gclk));
	jxor g5000(.dina(w_n5084_0[2]),.dinb(w_n5082_0[1]),.dout(n5085),.clk(gclk));
	jor g5001(.dina(w_n5044_0[0]),.dinb(w_n5024_0[0]),.dout(n5086),.clk(gclk));
	jxor g5002(.dina(w_n5083_0[1]),.dinb(w_n5058_0[0]),.dout(n5087),.clk(gclk));
	jor g5003(.dina(n5087),.dinb(w_dff_B_4LMWvph54_1),.dout(n5088),.clk(gclk));
	jand g5004(.dina(w_n5088_0[1]),.dinb(w_n4013_4[2]),.dout(n5089),.clk(gclk));
	jxor g5005(.dina(n5089),.dinb(w_n5085_0[1]),.dout(w_dff_A_Cw7elsfJ2_2),.clk(gclk));
	jand g5006(.dina(w_n5083_0[0]),.dinb(w_n5056_0[0]),.dout(n5091),.clk(gclk));
	jxor g5007(.dina(w_n5081_0[1]),.dinb(w_n5091_0[1]),.dout(n5092),.clk(gclk));
	jxor g5008(.dina(w_n5084_0[1]),.dinb(w_n5092_0[1]),.dout(n5093),.clk(gclk));
	jand g5009(.dina(w_n5069_0[0]),.dinb(w_n5050_0[0]),.dout(n5094),.clk(gclk));
	jand g5010(.dina(n5094),.dinb(w_dff_B_OP6iqswc4_1),.dout(n5095),.clk(gclk));
	jor g5011(.dina(w_n5095_0[1]),.dinb(w_n5046_0[0]),.dout(n5096),.clk(gclk));
	jnot g5012(.din(w_n5081_0[0]),.dout(n5097),.clk(gclk));
	jand g5013(.dina(n5097),.dinb(w_n5091_0[0]),.dout(n5098),.clk(gclk));
	jand g5014(.dina(w_n5084_0[0]),.dinb(w_n5082_0[0]),.dout(n5099),.clk(gclk));
	jor g5015(.dina(w_n5099_0[1]),.dinb(w_n5098_0[1]),.dout(n5100),.clk(gclk));
	jand g5016(.dina(w_n733_0[1]),.dinb(w_n494_0[0]),.dout(n5101),.clk(gclk));
	jand g5017(.dina(n5101),.dinb(w_n2542_0[0]),.dout(n5102),.clk(gclk));
	jand g5018(.dina(w_n724_0[2]),.dinb(w_n323_1[0]),.dout(n5103),.clk(gclk));
	jand g5019(.dina(n5103),.dinb(w_n214_0[2]),.dout(n5104),.clk(gclk));
	jand g5020(.dina(n5104),.dinb(w_n4355_0[0]),.dout(n5105),.clk(gclk));
	jand g5021(.dina(n5105),.dinb(n5102),.dout(n5106),.clk(gclk));
	jand g5022(.dina(n5106),.dinb(w_n786_0[1]),.dout(n5107),.clk(gclk));
	jand g5023(.dina(n5107),.dinb(w_n4589_0[0]),.dout(n5108),.clk(gclk));
	jand g5024(.dina(n5108),.dinb(w_n636_0[0]),.dout(n5109),.clk(gclk));
	jxor g5025(.dina(w_n5109_0[2]),.dinb(w_n5100_0[1]),.dout(n5110),.clk(gclk));
	jxor g5026(.dina(w_n5110_0[1]),.dinb(n5096),.dout(w_dff_A_gS2lI5Ue9_2),.clk(gclk));
	jnot g5027(.din(w_n5109_0[1]),.dout(n5112),.clk(gclk));
	jand g5028(.dina(w_n5112_0[2]),.dinb(w_n5098_0[0]),.dout(n5113),.clk(gclk));
	jand g5029(.dina(w_n3592_0[0]),.dinb(w_n664_0[0]),.dout(n5114),.clk(gclk));
	jand g5030(.dina(n5114),.dinb(w_n722_0[0]),.dout(n5115),.clk(gclk));
	jand g5031(.dina(n5115),.dinb(w_n334_0[2]),.dout(n5116),.clk(gclk));
	jnot g5032(.din(w_n5116_0[1]),.dout(n5117),.clk(gclk));
	jxor g5033(.dina(w_n5117_0[1]),.dinb(w_n5113_0[2]),.dout(n5118),.clk(gclk));
	jand g5034(.dina(w_n5112_0[1]),.dinb(w_n5099_0[0]),.dout(n5119),.clk(gclk));
	jxor g5035(.dina(w_n5119_0[2]),.dinb(w_n5118_0[1]),.dout(n5120),.clk(gclk));
	jor g5036(.dina(w_n5088_0[0]),.dinb(w_n5085_0[0]),.dout(n5121),.clk(gclk));
	jxor g5037(.dina(w_n5112_0[0]),.dinb(w_n5100_0[0]),.dout(n5122),.clk(gclk));
	jor g5038(.dina(n5122),.dinb(n5121),.dout(n5123),.clk(gclk));
	jand g5039(.dina(w_n5123_0[1]),.dinb(w_n4013_4[1]),.dout(n5124),.clk(gclk));
	jxor g5040(.dina(n5124),.dinb(w_n5120_0[1]),.dout(w_dff_A_TNSINLGv9_2),.clk(gclk));
	jor g5041(.dina(w_n5123_0[0]),.dinb(w_n5120_0[0]),.dout(n5126),.clk(gclk));
	jand g5042(.dina(w_n5126_0[1]),.dinb(w_n4013_4[0]),.dout(n5127),.clk(gclk));
	jand g5043(.dina(w_n779_0[0]),.dinb(w_n334_0[1]),.dout(n5128),.clk(gclk));
	jnot g5044(.din(w_n5128_0[1]),.dout(n5129),.clk(gclk));
	jand g5045(.dina(w_n5117_0[0]),.dinb(w_n5113_0[1]),.dout(n5130),.clk(gclk));
	jand g5046(.dina(w_n5119_0[1]),.dinb(w_n5118_0[0]),.dout(n5131),.clk(gclk));
	jor g5047(.dina(n5131),.dinb(w_n5130_0[1]),.dout(n5132),.clk(gclk));
	jxor g5048(.dina(w_n5132_0[1]),.dinb(w_n5129_0[1]),.dout(n5133),.clk(gclk));
	jxor g5049(.dina(w_n5133_0[1]),.dinb(n5127),.dout(w_dff_A_HR8wY1806_2),.clk(gclk));
	jnot g5050(.din(w_a21_0[0]),.dout(n5135),.clk(gclk));
	jand g5051(.dina(w_n49_1[2]),.dinb(n5135),.dout(n5136),.clk(gclk));
	jand g5052(.dina(n5136),.dinb(w_n207_0[0]),.dout(n5137),.clk(gclk));
	jor g5053(.dina(w_n5133_0[0]),.dinb(w_n5126_0[0]),.dout(n5138),.clk(gclk));
	jand g5054(.dina(w_n5138_0[1]),.dinb(w_n4013_3[2]),.dout(n5139),.clk(gclk));
	jand g5055(.dina(w_n5132_0[0]),.dinb(w_n5129_0[0]),.dout(n5140),.clk(gclk));
	jnot g5056(.din(w_n5130_0[0]),.dout(n5141),.clk(gclk));
	jxor g5057(.dina(w_n5116_0[0]),.dinb(w_n5113_0[0]),.dout(n5142),.clk(gclk));
	jxor g5058(.dina(w_n5042_0[1]),.dinb(w_n5054_0[0]),.dout(n5143),.clk(gclk));
	jor g5059(.dina(n5143),.dinb(w_n5048_0[0]),.dout(n5144),.clk(gclk));
	jor g5060(.dina(w_n5068_0[1]),.dinb(n5144),.dout(n5145),.clk(gclk));
	jor g5061(.dina(n5145),.dinb(w_n5092_0[0]),.dout(n5146),.clk(gclk));
	jor g5062(.dina(w_n5109_0[0]),.dinb(n5146),.dout(n5147),.clk(gclk));
	jor g5063(.dina(n5147),.dinb(w_n5142_0[1]),.dout(n5148),.clk(gclk));
	jor g5064(.dina(n5148),.dinb(n5141),.dout(n5149),.clk(gclk));
	jxor g5065(.dina(w_n5140_0[1]),.dinb(n5139),.dout(n5151),.clk(gclk));
	jor g5066(.dina(n5151),.dinb(w_n5137_0[1]),.dout(sin23),.clk(gclk));
	jor g5067(.dina(n5149),.dinb(w_n5128_0[0]),.dout(n5153),.clk(gclk));
	jand g5068(.dina(w_dff_B_d9hBrptt6_0),.dinb(w_n5138_0[0]),.dout(n5154),.clk(gclk));
	jxor g5069(.dina(w_n5119_0[0]),.dinb(w_n5142_0[0]),.dout(n5155),.clk(gclk));
	jand g5070(.dina(w_n5110_0[0]),.dinb(w_n5095_0[0]),.dout(n5156),.clk(gclk));
	jand g5071(.dina(n5156),.dinb(w_dff_B_2rz4dWGZ7_1),.dout(n5157),.clk(gclk));
	jand g5072(.dina(w_n5140_0[0]),.dinb(n5157),.dout(n5158),.clk(gclk));
	jor g5073(.dina(n5158),.dinb(w_n5137_0[0]),.dout(n5159),.clk(gclk));
	jor g5074(.dina(n5159),.dinb(n5154),.dout(n5160),.clk(gclk));
	jand g5075(.dina(n5160),.dinb(w_n4013_3[1]),.dout(sin24),.clk(gclk));
	jspl3 jspl3_w_a0_0(.douta(w_a0_0[0]),.doutb(w_a0_0[1]),.doutc(w_a0_0[2]),.din(a0));
	jspl jspl_w_a0_1(.douta(w_a0_1[0]),.doutb(w_a0_1[1]),.din(w_a0_0[0]));
	jspl3 jspl3_w_a1_0(.douta(w_a1_0[0]),.doutb(w_a1_0[1]),.doutc(w_a1_0[2]),.din(a1));
	jspl3 jspl3_w_a2_0(.douta(w_a2_0[0]),.doutb(w_a2_0[1]),.doutc(w_a2_0[2]),.din(a2));
	jspl3 jspl3_w_a2_1(.douta(w_a2_1[0]),.doutb(w_a2_1[1]),.doutc(w_a2_1[2]),.din(w_a2_0[0]));
	jspl3 jspl3_w_a3_0(.douta(w_a3_0[0]),.doutb(w_a3_0[1]),.doutc(w_a3_0[2]),.din(a3));
	jspl3 jspl3_w_a4_0(.douta(w_a4_0[0]),.doutb(w_a4_0[1]),.doutc(w_a4_0[2]),.din(a4));
	jspl jspl_w_a4_1(.douta(w_a4_1[0]),.doutb(w_a4_1[1]),.din(w_a4_0[0]));
	jspl3 jspl3_w_a5_0(.douta(w_a5_0[0]),.doutb(w_a5_0[1]),.doutc(w_a5_0[2]),.din(a5));
	jspl3 jspl3_w_a6_0(.douta(w_a6_0[0]),.doutb(w_a6_0[1]),.doutc(w_a6_0[2]),.din(a6));
	jspl jspl_w_a6_1(.douta(w_a6_1[0]),.doutb(w_a6_1[1]),.din(w_a6_0[0]));
	jspl3 jspl3_w_a7_0(.douta(w_a7_0[0]),.doutb(w_a7_0[1]),.doutc(w_a7_0[2]),.din(a7));
	jspl3 jspl3_w_a8_0(.douta(w_a8_0[0]),.doutb(w_a8_0[1]),.doutc(w_a8_0[2]),.din(a8));
	jspl jspl_w_a8_1(.douta(w_a8_1[0]),.doutb(w_a8_1[1]),.din(w_a8_0[0]));
	jspl3 jspl3_w_a9_0(.douta(w_a9_0[0]),.doutb(w_a9_0[1]),.doutc(w_a9_0[2]),.din(a9));
	jspl3 jspl3_w_a10_0(.douta(w_a10_0[0]),.doutb(w_a10_0[1]),.doutc(w_a10_0[2]),.din(a10));
	jspl jspl_w_a10_1(.douta(w_a10_1[0]),.doutb(w_a10_1[1]),.din(w_a10_0[0]));
	jspl3 jspl3_w_a11_0(.douta(w_a11_0[0]),.doutb(w_a11_0[1]),.doutc(w_a11_0[2]),.din(a11));
	jspl3 jspl3_w_a12_0(.douta(w_a12_0[0]),.doutb(w_a12_0[1]),.doutc(w_a12_0[2]),.din(a12));
	jspl jspl_w_a12_1(.douta(w_a12_1[0]),.doutb(w_a12_1[1]),.din(w_a12_0[0]));
	jspl3 jspl3_w_a13_0(.douta(w_a13_0[0]),.doutb(w_a13_0[1]),.doutc(w_a13_0[2]),.din(a13));
	jspl3 jspl3_w_a14_0(.douta(w_a14_0[0]),.doutb(w_a14_0[1]),.doutc(w_a14_0[2]),.din(a14));
	jspl jspl_w_a14_1(.douta(w_a14_1[0]),.doutb(w_a14_1[1]),.din(w_a14_0[0]));
	jspl3 jspl3_w_a15_0(.douta(w_a15_0[0]),.doutb(w_a15_0[1]),.doutc(w_a15_0[2]),.din(a15));
	jspl jspl_w_a15_1(.douta(w_a15_1[0]),.doutb(w_a15_1[1]),.din(w_a15_0[0]));
	jspl3 jspl3_w_a16_0(.douta(w_a16_0[0]),.doutb(w_a16_0[1]),.doutc(w_a16_0[2]),.din(a16));
	jspl jspl_w_a17_0(.douta(w_a17_0[0]),.doutb(w_a17_0[1]),.din(a17));
	jspl3 jspl3_w_a18_0(.douta(w_a18_0[0]),.doutb(w_a18_0[1]),.doutc(w_a18_0[2]),.din(a18));
	jspl jspl_w_a18_1(.douta(w_a18_1[0]),.doutb(w_a18_1[1]),.din(w_a18_0[0]));
	jspl3 jspl3_w_a19_0(.douta(w_a19_0[0]),.doutb(w_a19_0[1]),.doutc(w_a19_0[2]),.din(a19));
	jspl3 jspl3_w_a20_0(.douta(w_a20_0[0]),.doutb(w_a20_0[1]),.doutc(w_a20_0[2]),.din(a20));
	jspl jspl_w_a20_1(.douta(w_a20_1[0]),.doutb(w_a20_1[1]),.din(w_a20_0[0]));
	jspl jspl_w_a21_0(.douta(w_a21_0[0]),.doutb(w_a21_0[1]),.din(a21));
	jspl3 jspl3_w_a22_0(.douta(w_a22_0[0]),.doutb(w_a22_0[1]),.doutc(w_a22_0[2]),.din(a22));
	jspl3 jspl3_w_a22_1(.douta(w_a22_1[0]),.doutb(w_a22_1[1]),.doutc(w_a22_1[2]),.din(w_a22_0[0]));
	jspl3 jspl3_w_a22_2(.douta(w_a22_2[0]),.doutb(w_a22_2[1]),.doutc(w_a22_2[2]),.din(w_a22_0[1]));
	jspl3 jspl3_w_a22_3(.douta(w_a22_3[0]),.doutb(w_a22_3[1]),.doutc(w_a22_3[2]),.din(w_a22_0[2]));
	jspl3 jspl3_w_a22_4(.douta(w_a22_4[0]),.doutb(w_a22_4[1]),.doutc(w_a22_4[2]),.din(w_a22_1[0]));
	jspl3 jspl3_w_a22_5(.douta(w_a22_5[0]),.doutb(w_a22_5[1]),.doutc(w_a22_5[2]),.din(w_a22_1[1]));
	jspl jspl_w_a22_6(.douta(w_a22_6[0]),.doutb(w_a22_6[1]),.din(w_a22_1[2]));
	jspl3 jspl3_w_sin0_0(.douta(w_dff_A_Op0hX5fq0_0),.doutb(w_sin0_0[1]),.doutc(w_dff_A_D1xwlsPT1_2),.din(sin0_fa_));
	jspl3 jspl3_w_n49_0(.douta(w_n49_0[0]),.doutb(w_n49_0[1]),.doutc(w_n49_0[2]),.din(n49));
	jspl3 jspl3_w_n49_1(.douta(w_n49_1[0]),.doutb(w_n49_1[1]),.doutc(w_n49_1[2]),.din(w_n49_0[0]));
	jspl3 jspl3_w_n49_2(.douta(w_n49_2[0]),.doutb(w_n49_2[1]),.doutc(w_n49_2[2]),.din(w_n49_0[1]));
	jspl3 jspl3_w_n49_3(.douta(w_n49_3[0]),.doutb(w_n49_3[1]),.doutc(w_n49_3[2]),.din(w_n49_0[2]));
	jspl3 jspl3_w_n49_4(.douta(w_n49_4[0]),.doutb(w_n49_4[1]),.doutc(w_n49_4[2]),.din(w_n49_1[0]));
	jspl jspl_w_n49_5(.douta(w_n49_5[0]),.doutb(w_n49_5[1]),.din(w_n49_1[1]));
	jspl jspl_w_n51_0(.douta(w_n51_0[0]),.doutb(w_n51_0[1]),.din(n51));
	jspl jspl_w_n52_0(.douta(w_n52_0[0]),.doutb(w_n52_0[1]),.din(n52));
	jspl jspl_w_n53_0(.douta(w_n53_0[0]),.doutb(w_n53_0[1]),.din(n53));
	jspl jspl_w_n54_0(.douta(w_n54_0[0]),.doutb(w_n54_0[1]),.din(n54));
	jspl3 jspl3_w_n55_0(.douta(w_n55_0[0]),.doutb(w_n55_0[1]),.doutc(w_n55_0[2]),.din(n55));
	jspl3 jspl3_w_n55_1(.douta(w_n55_1[0]),.doutb(w_n55_1[1]),.doutc(w_n55_1[2]),.din(w_n55_0[0]));
	jspl3 jspl3_w_n55_2(.douta(w_n55_2[0]),.doutb(w_n55_2[1]),.doutc(w_n55_2[2]),.din(w_n55_0[1]));
	jspl3 jspl3_w_n55_3(.douta(w_n55_3[0]),.doutb(w_n55_3[1]),.doutc(w_n55_3[2]),.din(w_n55_0[2]));
	jspl3 jspl3_w_n55_4(.douta(w_n55_4[0]),.doutb(w_n55_4[1]),.doutc(w_n55_4[2]),.din(w_n55_1[0]));
	jspl3 jspl3_w_n55_5(.douta(w_n55_5[0]),.doutb(w_n55_5[1]),.doutc(w_n55_5[2]),.din(w_n55_1[1]));
	jspl3 jspl3_w_n55_6(.douta(w_n55_6[0]),.doutb(w_n55_6[1]),.doutc(w_n55_6[2]),.din(w_n55_1[2]));
	jspl3 jspl3_w_n55_7(.douta(w_n55_7[0]),.doutb(w_n55_7[1]),.doutc(w_n55_7[2]),.din(w_n55_2[0]));
	jspl3 jspl3_w_n55_8(.douta(w_n55_8[0]),.doutb(w_n55_8[1]),.doutc(w_n55_8[2]),.din(w_n55_2[1]));
	jspl3 jspl3_w_n55_9(.douta(w_n55_9[0]),.doutb(w_n55_9[1]),.doutc(w_n55_9[2]),.din(w_n55_2[2]));
	jspl3 jspl3_w_n56_0(.douta(w_n56_0[0]),.doutb(w_n56_0[1]),.doutc(w_n56_0[2]),.din(n56));
	jspl3 jspl3_w_n56_1(.douta(w_n56_1[0]),.doutb(w_n56_1[1]),.doutc(w_n56_1[2]),.din(w_n56_0[0]));
	jspl3 jspl3_w_n56_2(.douta(w_n56_2[0]),.doutb(w_n56_2[1]),.doutc(w_n56_2[2]),.din(w_n56_0[1]));
	jspl3 jspl3_w_n56_3(.douta(w_n56_3[0]),.doutb(w_n56_3[1]),.doutc(w_n56_3[2]),.din(w_n56_0[2]));
	jspl3 jspl3_w_n56_4(.douta(w_n56_4[0]),.doutb(w_n56_4[1]),.doutc(w_n56_4[2]),.din(w_n56_1[0]));
	jspl3 jspl3_w_n56_5(.douta(w_n56_5[0]),.doutb(w_n56_5[1]),.doutc(w_n56_5[2]),.din(w_n56_1[1]));
	jspl3 jspl3_w_n56_6(.douta(w_n56_6[0]),.doutb(w_n56_6[1]),.doutc(w_n56_6[2]),.din(w_n56_1[2]));
	jspl3 jspl3_w_n56_7(.douta(w_n56_7[0]),.doutb(w_n56_7[1]),.doutc(w_n56_7[2]),.din(w_n56_2[0]));
	jspl3 jspl3_w_n56_8(.douta(w_n56_8[0]),.doutb(w_n56_8[1]),.doutc(w_n56_8[2]),.din(w_n56_2[1]));
	jspl3 jspl3_w_n56_9(.douta(w_n56_9[0]),.doutb(w_n56_9[1]),.doutc(w_n56_9[2]),.din(w_n56_2[2]));
	jspl3 jspl3_w_n56_10(.douta(w_n56_10[0]),.doutb(w_n56_10[1]),.doutc(w_n56_10[2]),.din(w_n56_3[0]));
	jspl3 jspl3_w_n56_11(.douta(w_n56_11[0]),.doutb(w_n56_11[1]),.doutc(w_n56_11[2]),.din(w_n56_3[1]));
	jspl3 jspl3_w_n56_12(.douta(w_n56_12[0]),.doutb(w_n56_12[1]),.doutc(w_n56_12[2]),.din(w_n56_3[2]));
	jspl jspl_w_n57_0(.douta(w_n57_0[0]),.doutb(w_n57_0[1]),.din(n57));
	jspl3 jspl3_w_n58_0(.douta(w_n58_0[0]),.doutb(w_n58_0[1]),.doutc(w_n58_0[2]),.din(n58));
	jspl3 jspl3_w_n58_1(.douta(w_n58_1[0]),.doutb(w_n58_1[1]),.doutc(w_n58_1[2]),.din(w_n58_0[0]));
	jspl3 jspl3_w_n58_2(.douta(w_n58_2[0]),.doutb(w_n58_2[1]),.doutc(w_n58_2[2]),.din(w_n58_0[1]));
	jspl3 jspl3_w_n58_3(.douta(w_n58_3[0]),.doutb(w_n58_3[1]),.doutc(w_n58_3[2]),.din(w_n58_0[2]));
	jspl3 jspl3_w_n58_4(.douta(w_n58_4[0]),.doutb(w_n58_4[1]),.doutc(w_n58_4[2]),.din(w_n58_1[0]));
	jspl3 jspl3_w_n59_0(.douta(w_n59_0[0]),.doutb(w_n59_0[1]),.doutc(w_n59_0[2]),.din(n59));
	jspl3 jspl3_w_n59_1(.douta(w_n59_1[0]),.doutb(w_n59_1[1]),.doutc(w_n59_1[2]),.din(w_n59_0[0]));
	jspl3 jspl3_w_n59_2(.douta(w_n59_2[0]),.doutb(w_n59_2[1]),.doutc(w_n59_2[2]),.din(w_n59_0[1]));
	jspl jspl_w_n59_3(.douta(w_n59_3[0]),.doutb(w_n59_3[1]),.din(w_n59_0[2]));
	jspl3 jspl3_w_n61_0(.douta(w_n61_0[0]),.doutb(w_n61_0[1]),.doutc(w_n61_0[2]),.din(n61));
	jspl3 jspl3_w_n61_1(.douta(w_n61_1[0]),.doutb(w_n61_1[1]),.doutc(w_n61_1[2]),.din(w_n61_0[0]));
	jspl3 jspl3_w_n62_0(.douta(w_n62_0[0]),.doutb(w_n62_0[1]),.doutc(w_n62_0[2]),.din(n62));
	jspl3 jspl3_w_n63_0(.douta(w_n63_0[0]),.doutb(w_n63_0[1]),.doutc(w_n63_0[2]),.din(n63));
	jspl3 jspl3_w_n63_1(.douta(w_n63_1[0]),.doutb(w_n63_1[1]),.doutc(w_n63_1[2]),.din(w_n63_0[0]));
	jspl3 jspl3_w_n63_2(.douta(w_n63_2[0]),.doutb(w_n63_2[1]),.doutc(w_n63_2[2]),.din(w_n63_0[1]));
	jspl jspl_w_n64_0(.douta(w_n64_0[0]),.doutb(w_n64_0[1]),.din(n64));
	jspl3 jspl3_w_n68_0(.douta(w_n68_0[0]),.doutb(w_n68_0[1]),.doutc(w_n68_0[2]),.din(n68));
	jspl3 jspl3_w_n68_1(.douta(w_n68_1[0]),.doutb(w_n68_1[1]),.doutc(w_n68_1[2]),.din(w_n68_0[0]));
	jspl3 jspl3_w_n68_2(.douta(w_n68_2[0]),.doutb(w_n68_2[1]),.doutc(w_n68_2[2]),.din(w_n68_0[1]));
	jspl3 jspl3_w_n68_3(.douta(w_n68_3[0]),.doutb(w_n68_3[1]),.doutc(w_n68_3[2]),.din(w_n68_0[2]));
	jspl3 jspl3_w_n68_4(.douta(w_n68_4[0]),.doutb(w_n68_4[1]),.doutc(w_n68_4[2]),.din(w_n68_1[0]));
	jspl3 jspl3_w_n68_5(.douta(w_n68_5[0]),.doutb(w_n68_5[1]),.doutc(w_n68_5[2]),.din(w_n68_1[1]));
	jspl3 jspl3_w_n68_6(.douta(w_n68_6[0]),.doutb(w_n68_6[1]),.doutc(w_n68_6[2]),.din(w_n68_1[2]));
	jspl3 jspl3_w_n69_0(.douta(w_n69_0[0]),.doutb(w_n69_0[1]),.doutc(w_n69_0[2]),.din(n69));
	jspl3 jspl3_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.doutc(w_n70_0[2]),.din(n70));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.doutc(w_n75_0[2]),.din(n75));
	jspl3 jspl3_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.doutc(w_n75_1[2]),.din(w_n75_0[0]));
	jspl3 jspl3_w_n75_2(.douta(w_n75_2[0]),.doutb(w_n75_2[1]),.doutc(w_n75_2[2]),.din(w_n75_0[1]));
	jspl3 jspl3_w_n75_3(.douta(w_n75_3[0]),.doutb(w_n75_3[1]),.doutc(w_n75_3[2]),.din(w_n75_0[2]));
	jspl3 jspl3_w_n75_4(.douta(w_n75_4[0]),.doutb(w_n75_4[1]),.doutc(w_n75_4[2]),.din(w_n75_1[0]));
	jspl3 jspl3_w_n75_5(.douta(w_n75_5[0]),.doutb(w_n75_5[1]),.doutc(w_n75_5[2]),.din(w_n75_1[1]));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.din(n76));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl3 jspl3_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.doutc(w_n78_0[2]),.din(n78));
	jspl3 jspl3_w_n78_1(.douta(w_n78_1[0]),.doutb(w_n78_1[1]),.doutc(w_n78_1[2]),.din(w_n78_0[0]));
	jspl3 jspl3_w_n78_2(.douta(w_n78_2[0]),.doutb(w_n78_2[1]),.doutc(w_n78_2[2]),.din(w_n78_0[1]));
	jspl3 jspl3_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.doutc(w_n79_0[2]),.din(n79));
	jspl3 jspl3_w_n79_1(.douta(w_n79_1[0]),.doutb(w_n79_1[1]),.doutc(w_n79_1[2]),.din(w_n79_0[0]));
	jspl3 jspl3_w_n79_2(.douta(w_n79_2[0]),.doutb(w_n79_2[1]),.doutc(w_n79_2[2]),.din(w_n79_0[1]));
	jspl3 jspl3_w_n79_3(.douta(w_n79_3[0]),.doutb(w_n79_3[1]),.doutc(w_n79_3[2]),.din(w_n79_0[2]));
	jspl3 jspl3_w_n79_4(.douta(w_n79_4[0]),.doutb(w_n79_4[1]),.doutc(w_n79_4[2]),.din(w_n79_1[0]));
	jspl3 jspl3_w_n79_5(.douta(w_n79_5[0]),.doutb(w_n79_5[1]),.doutc(w_n79_5[2]),.din(w_n79_1[1]));
	jspl jspl_w_n79_6(.douta(w_n79_6[0]),.doutb(w_n79_6[1]),.din(w_n79_1[2]));
	jspl jspl_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.din(n81));
	jspl jspl_w_n82_0(.douta(w_n82_0[0]),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n87_0(.douta(w_n87_0[0]),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n89_0(.douta(w_n89_0[0]),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.din(n91));
	jspl jspl_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.din(n92));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.doutc(w_n96_0[2]),.din(n96));
	jspl3 jspl3_w_n96_1(.douta(w_n96_1[0]),.doutb(w_n96_1[1]),.doutc(w_n96_1[2]),.din(w_n96_0[0]));
	jspl3 jspl3_w_n96_2(.douta(w_n96_2[0]),.doutb(w_n96_2[1]),.doutc(w_n96_2[2]),.din(w_n96_0[1]));
	jspl3 jspl3_w_n96_3(.douta(w_n96_3[0]),.doutb(w_n96_3[1]),.doutc(w_n96_3[2]),.din(w_n96_0[2]));
	jspl3 jspl3_w_n96_4(.douta(w_n96_4[0]),.doutb(w_n96_4[1]),.doutc(w_n96_4[2]),.din(w_n96_1[0]));
	jspl3 jspl3_w_n96_5(.douta(w_n96_5[0]),.doutb(w_n96_5[1]),.doutc(w_n96_5[2]),.din(w_n96_1[1]));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n100_0(.douta(w_n100_0[0]),.doutb(w_n100_0[1]),.din(n100));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.doutc(w_n103_0[2]),.din(n103));
	jspl jspl_w_n103_1(.douta(w_n103_1[0]),.doutb(w_n103_1[1]),.din(w_n103_0[0]));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n105_0(.douta(w_n105_0[0]),.doutb(w_n105_0[1]),.din(n105));
	jspl3 jspl3_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.doutc(w_n108_0[2]),.din(n108));
	jspl jspl_w_n108_1(.douta(w_n108_1[0]),.doutb(w_n108_1[1]),.din(w_n108_0[0]));
	jspl3 jspl3_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.doutc(w_n109_0[2]),.din(n109));
	jspl3 jspl3_w_n109_1(.douta(w_n109_1[0]),.doutb(w_n109_1[1]),.doutc(w_n109_1[2]),.din(w_n109_0[0]));
	jspl jspl_w_n109_2(.douta(w_n109_2[0]),.doutb(w_n109_2[1]),.din(w_n109_0[1]));
	jspl3 jspl3_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.doutc(w_n110_0[2]),.din(n110));
	jspl3 jspl3_w_n110_1(.douta(w_n110_1[0]),.doutb(w_n110_1[1]),.doutc(w_n110_1[2]),.din(w_n110_0[0]));
	jspl3 jspl3_w_n110_2(.douta(w_n110_2[0]),.doutb(w_n110_2[1]),.doutc(w_n110_2[2]),.din(w_n110_0[1]));
	jspl3 jspl3_w_n110_3(.douta(w_n110_3[0]),.doutb(w_n110_3[1]),.doutc(w_n110_3[2]),.din(w_n110_0[2]));
	jspl3 jspl3_w_n110_4(.douta(w_n110_4[0]),.doutb(w_n110_4[1]),.doutc(w_n110_4[2]),.din(w_n110_1[0]));
	jspl3 jspl3_w_n110_5(.douta(w_n110_5[0]),.doutb(w_n110_5[1]),.doutc(w_n110_5[2]),.din(w_n110_1[1]));
	jspl jspl_w_n110_6(.douta(w_n110_6[0]),.doutb(w_n110_6[1]),.din(w_n110_1[2]));
	jspl jspl_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.doutc(w_n116_0[2]),.din(n116));
	jspl jspl_w_n116_1(.douta(w_n116_1[0]),.doutb(w_n116_1[1]),.din(w_n116_0[0]));
	jspl jspl_w_n117_0(.douta(w_n117_0[0]),.doutb(w_n117_0[1]),.din(n117));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl3 jspl3_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.doutc(w_n120_0[2]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl3 jspl3_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.doutc(w_n123_0[2]),.din(n123));
	jspl jspl_w_n123_1(.douta(w_n123_1[0]),.doutb(w_n123_1[1]),.din(w_n123_0[0]));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl3 jspl3_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.doutc(w_n127_0[2]),.din(n127));
	jspl jspl_w_n127_1(.douta(w_n127_1[0]),.doutb(w_n127_1[1]),.din(w_n127_0[0]));
	jspl3 jspl3_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.doutc(w_n128_0[2]),.din(n128));
	jspl3 jspl3_w_n128_1(.douta(w_n128_1[0]),.doutb(w_n128_1[1]),.doutc(w_n128_1[2]),.din(w_n128_0[0]));
	jspl3 jspl3_w_n128_2(.douta(w_n128_2[0]),.doutb(w_n128_2[1]),.doutc(w_n128_2[2]),.din(w_n128_0[1]));
	jspl3 jspl3_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.doutc(w_n130_0[2]),.din(n130));
	jspl3 jspl3_w_n130_1(.douta(w_n130_1[0]),.doutb(w_n130_1[1]),.doutc(w_n130_1[2]),.din(w_n130_0[0]));
	jspl3 jspl3_w_n130_2(.douta(w_n130_2[0]),.doutb(w_n130_2[1]),.doutc(w_n130_2[2]),.din(w_n130_0[1]));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n134_0(.douta(w_n134_0[0]),.doutb(w_n134_0[1]),.doutc(w_n134_0[2]),.din(n134));
	jspl jspl_w_n134_1(.douta(w_n134_1[0]),.doutb(w_n134_1[1]),.din(w_n134_0[0]));
	jspl3 jspl3_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.doutc(w_n135_0[2]),.din(n135));
	jspl3 jspl3_w_n135_1(.douta(w_n135_1[0]),.doutb(w_n135_1[1]),.doutc(w_n135_1[2]),.din(w_n135_0[0]));
	jspl3 jspl3_w_n135_2(.douta(w_n135_2[0]),.doutb(w_n135_2[1]),.doutc(w_n135_2[2]),.din(w_n135_0[1]));
	jspl3 jspl3_w_n136_0(.douta(w_n136_0[0]),.doutb(w_n136_0[1]),.doutc(w_n136_0[2]),.din(n136));
	jspl jspl_w_n137_0(.douta(w_n137_0[0]),.doutb(w_n137_0[1]),.din(n137));
	jspl3 jspl3_w_n138_0(.douta(w_n138_0[0]),.doutb(w_n138_0[1]),.doutc(w_n138_0[2]),.din(n138));
	jspl3 jspl3_w_n138_1(.douta(w_n138_1[0]),.doutb(w_n138_1[1]),.doutc(w_n138_1[2]),.din(w_n138_0[0]));
	jspl3 jspl3_w_n138_2(.douta(w_n138_2[0]),.doutb(w_n138_2[1]),.doutc(w_n138_2[2]),.din(w_n138_0[1]));
	jspl3 jspl3_w_n138_3(.douta(w_n138_3[0]),.doutb(w_n138_3[1]),.doutc(w_n138_3[2]),.din(w_n138_0[2]));
	jspl jspl_w_n138_4(.douta(w_n138_4[0]),.doutb(w_n138_4[1]),.din(w_n138_1[0]));
	jspl3 jspl3_w_n139_0(.douta(w_n139_0[0]),.doutb(w_n139_0[1]),.doutc(w_n139_0[2]),.din(n139));
	jspl jspl_w_n139_1(.douta(w_n139_1[0]),.doutb(w_n139_1[1]),.din(w_n139_0[0]));
	jspl3 jspl3_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.doutc(w_n140_0[2]),.din(n140));
	jspl jspl_w_n140_1(.douta(w_n140_1[0]),.doutb(w_n140_1[1]),.din(w_n140_0[0]));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl3 jspl3_w_n141_1(.douta(w_n141_1[0]),.doutb(w_n141_1[1]),.doutc(w_n141_1[2]),.din(w_n141_0[0]));
	jspl jspl_w_n141_2(.douta(w_n141_2[0]),.doutb(w_n141_2[1]),.din(w_n141_0[1]));
	jspl3 jspl3_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.doutc(w_n142_0[2]),.din(n142));
	jspl jspl_w_n142_1(.douta(w_n142_1[0]),.doutb(w_n142_1[1]),.din(w_n142_0[0]));
	jspl3 jspl3_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.doutc(w_n143_0[2]),.din(n143));
	jspl3 jspl3_w_n143_1(.douta(w_n143_1[0]),.doutb(w_n143_1[1]),.doutc(w_n143_1[2]),.din(w_n143_0[0]));
	jspl3 jspl3_w_n143_2(.douta(w_n143_2[0]),.doutb(w_n143_2[1]),.doutc(w_n143_2[2]),.din(w_n143_0[1]));
	jspl3 jspl3_w_n143_3(.douta(w_n143_3[0]),.doutb(w_n143_3[1]),.doutc(w_n143_3[2]),.din(w_n143_0[2]));
	jspl3 jspl3_w_n143_4(.douta(w_n143_4[0]),.doutb(w_n143_4[1]),.doutc(w_n143_4[2]),.din(w_n143_1[0]));
	jspl3 jspl3_w_n143_5(.douta(w_n143_5[0]),.doutb(w_n143_5[1]),.doutc(w_n143_5[2]),.din(w_n143_1[1]));
	jspl jspl_w_n143_6(.douta(w_n143_6[0]),.doutb(w_n143_6[1]),.din(w_n143_1[2]));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.doutc(w_n145_0[2]),.din(n145));
	jspl jspl_w_n145_1(.douta(w_n145_1[0]),.doutb(w_n145_1[1]),.din(w_n145_0[0]));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.doutc(w_n146_0[2]),.din(n146));
	jspl3 jspl3_w_n146_1(.douta(w_n146_1[0]),.doutb(w_n146_1[1]),.doutc(w_n146_1[2]),.din(w_n146_0[0]));
	jspl3 jspl3_w_n146_2(.douta(w_n146_2[0]),.doutb(w_n146_2[1]),.doutc(w_n146_2[2]),.din(w_n146_0[1]));
	jspl3 jspl3_w_n146_3(.douta(w_n146_3[0]),.doutb(w_n146_3[1]),.doutc(w_n146_3[2]),.din(w_n146_0[2]));
	jspl3 jspl3_w_n146_4(.douta(w_n146_4[0]),.doutb(w_n146_4[1]),.doutc(w_n146_4[2]),.din(w_n146_1[0]));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl3 jspl3_w_n147_1(.douta(w_n147_1[0]),.doutb(w_n147_1[1]),.doutc(w_n147_1[2]),.din(w_n147_0[0]));
	jspl3 jspl3_w_n147_2(.douta(w_n147_2[0]),.doutb(w_n147_2[1]),.doutc(w_n147_2[2]),.din(w_n147_0[1]));
	jspl3 jspl3_w_n147_3(.douta(w_n147_3[0]),.doutb(w_n147_3[1]),.doutc(w_n147_3[2]),.din(w_n147_0[2]));
	jspl jspl_w_n147_4(.douta(w_n147_4[0]),.doutb(w_n147_4[1]),.din(w_n147_1[0]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_n151_1[1]),.doutc(w_n151_1[2]),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_n151_2[0]),.doutb(w_n151_2[1]),.doutc(w_n151_2[2]),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_n151_3[0]),.doutb(w_n151_3[1]),.doutc(w_n151_3[2]),.din(w_n151_0[2]));
	jspl3 jspl3_w_n151_4(.douta(w_n151_4[0]),.doutb(w_n151_4[1]),.doutc(w_n151_4[2]),.din(w_n151_1[0]));
	jspl3 jspl3_w_n151_5(.douta(w_n151_5[0]),.doutb(w_n151_5[1]),.doutc(w_n151_5[2]),.din(w_n151_1[1]));
	jspl jspl_w_n151_6(.douta(w_n151_6[0]),.doutb(w_n151_6[1]),.din(w_n151_1[2]));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl jspl_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_n154_0[2]),.din(n154));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl jspl_w_n155_1(.douta(w_n155_1[0]),.doutb(w_n155_1[1]),.din(w_n155_0[0]));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.doutc(w_n157_0[2]),.din(n157));
	jspl3 jspl3_w_n157_1(.douta(w_n157_1[0]),.doutb(w_n157_1[1]),.doutc(w_n157_1[2]),.din(w_n157_0[0]));
	jspl3 jspl3_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.doutc(w_n158_0[2]),.din(n158));
	jspl jspl_w_n158_1(.douta(w_n158_1[0]),.doutb(w_n158_1[1]),.din(w_n158_0[0]));
	jspl3 jspl3_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.doutc(w_n160_0[2]),.din(n160));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl3 jspl3_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.doutc(w_n162_0[2]),.din(n162));
	jspl jspl_w_n162_1(.douta(w_n162_1[0]),.doutb(w_n162_1[1]),.din(w_n162_0[0]));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_n163_0[2]),.din(n163));
	jspl3 jspl3_w_n163_1(.douta(w_n163_1[0]),.doutb(w_n163_1[1]),.doutc(w_n163_1[2]),.din(w_n163_0[0]));
	jspl3 jspl3_w_n163_2(.douta(w_n163_2[0]),.doutb(w_n163_2[1]),.doutc(w_n163_2[2]),.din(w_n163_0[1]));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_n164_0[2]),.din(n164));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(n165));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl3 jspl3_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.doutc(w_n211_0[2]),.din(n211));
	jspl jspl_w_n211_1(.douta(w_n211_1[0]),.doutb(w_n211_1[1]),.din(w_n211_0[0]));
	jspl3 jspl3_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.doutc(w_n212_0[2]),.din(n212));
	jspl3 jspl3_w_n212_1(.douta(w_n212_1[0]),.doutb(w_n212_1[1]),.doutc(w_n212_1[2]),.din(w_n212_0[0]));
	jspl3 jspl3_w_n212_2(.douta(w_n212_2[0]),.doutb(w_n212_2[1]),.doutc(w_n212_2[2]),.din(w_n212_0[1]));
	jspl jspl_w_n212_3(.douta(w_n212_3[0]),.doutb(w_n212_3[1]),.din(w_n212_0[2]));
	jspl3 jspl3_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.doutc(w_n213_0[2]),.din(n213));
	jspl jspl_w_n213_1(.douta(w_n213_1[0]),.doutb(w_n213_1[1]),.din(w_n213_0[0]));
	jspl3 jspl3_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.doutc(w_n214_0[2]),.din(n214));
	jspl3 jspl3_w_n214_1(.douta(w_n214_1[0]),.doutb(w_n214_1[1]),.doutc(w_n214_1[2]),.din(w_n214_0[0]));
	jspl3 jspl3_w_n214_2(.douta(w_n214_2[0]),.doutb(w_n214_2[1]),.doutc(w_n214_2[2]),.din(w_n214_0[1]));
	jspl3 jspl3_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.doutc(w_n215_0[2]),.din(n215));
	jspl3 jspl3_w_n215_1(.douta(w_n215_1[0]),.doutb(w_n215_1[1]),.doutc(w_n215_1[2]),.din(w_n215_0[0]));
	jspl jspl_w_n215_2(.douta(w_n215_2[0]),.doutb(w_n215_2[1]),.din(w_n215_0[1]));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.doutc(w_n216_0[2]),.din(n216));
	jspl3 jspl3_w_n216_1(.douta(w_n216_1[0]),.doutb(w_n216_1[1]),.doutc(w_n216_1[2]),.din(w_n216_0[0]));
	jspl3 jspl3_w_n216_2(.douta(w_n216_2[0]),.doutb(w_n216_2[1]),.doutc(w_n216_2[2]),.din(w_n216_0[1]));
	jspl3 jspl3_w_n216_3(.douta(w_n216_3[0]),.doutb(w_n216_3[1]),.doutc(w_n216_3[2]),.din(w_n216_0[2]));
	jspl jspl_w_n216_4(.douta(w_n216_4[0]),.doutb(w_n216_4[1]),.din(w_n216_1[0]));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.doutc(w_n219_0[2]),.din(n219));
	jspl jspl_w_n219_1(.douta(w_n219_1[0]),.doutb(w_n219_1[1]),.din(w_n219_0[0]));
	jspl3 jspl3_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.doutc(w_n220_0[2]),.din(n220));
	jspl3 jspl3_w_n220_1(.douta(w_n220_1[0]),.doutb(w_n220_1[1]),.doutc(w_n220_1[2]),.din(w_n220_0[0]));
	jspl3 jspl3_w_n220_2(.douta(w_n220_2[0]),.doutb(w_n220_2[1]),.doutc(w_n220_2[2]),.din(w_n220_0[1]));
	jspl jspl_w_n220_3(.douta(w_n220_3[0]),.doutb(w_n220_3[1]),.din(w_n220_0[2]));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.doutc(w_n222_0[2]),.din(n222));
	jspl3 jspl3_w_n222_1(.douta(w_n222_1[0]),.doutb(w_n222_1[1]),.doutc(w_n222_1[2]),.din(w_n222_0[0]));
	jspl jspl_w_n222_2(.douta(w_n222_2[0]),.doutb(w_n222_2[1]),.din(w_n222_0[1]));
	jspl3 jspl3_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.doutc(w_n223_0[2]),.din(n223));
	jspl3 jspl3_w_n223_1(.douta(w_n223_1[0]),.doutb(w_n223_1[1]),.doutc(w_n223_1[2]),.din(w_n223_0[0]));
	jspl3 jspl3_w_n223_2(.douta(w_n223_2[0]),.doutb(w_n223_2[1]),.doutc(w_n223_2[2]),.din(w_n223_0[1]));
	jspl3 jspl3_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.doutc(w_n224_0[2]),.din(n224));
	jspl3 jspl3_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.doutc(w_n225_0[2]),.din(n225));
	jspl3 jspl3_w_n225_1(.douta(w_n225_1[0]),.doutb(w_n225_1[1]),.doutc(w_n225_1[2]),.din(w_n225_0[0]));
	jspl3 jspl3_w_n225_2(.douta(w_n225_2[0]),.doutb(w_n225_2[1]),.doutc(w_n225_2[2]),.din(w_n225_0[1]));
	jspl3 jspl3_w_n227_0(.douta(w_n227_0[0]),.doutb(w_n227_0[1]),.doutc(w_n227_0[2]),.din(n227));
	jspl3 jspl3_w_n227_1(.douta(w_n227_1[0]),.doutb(w_n227_1[1]),.doutc(w_n227_1[2]),.din(w_n227_0[0]));
	jspl jspl_w_n227_2(.douta(w_n227_2[0]),.doutb(w_n227_2[1]),.din(w_n227_0[1]));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl3 jspl3_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.doutc(w_n229_0[2]),.din(n229));
	jspl3 jspl3_w_n229_1(.douta(w_n229_1[0]),.doutb(w_n229_1[1]),.doutc(w_n229_1[2]),.din(w_n229_0[0]));
	jspl3 jspl3_w_n229_2(.douta(w_n229_2[0]),.doutb(w_n229_2[1]),.doutc(w_n229_2[2]),.din(w_n229_0[1]));
	jspl3 jspl3_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.doutc(w_n230_0[2]),.din(n230));
	jspl3 jspl3_w_n230_1(.douta(w_n230_1[0]),.doutb(w_n230_1[1]),.doutc(w_n230_1[2]),.din(w_n230_0[0]));
	jspl jspl_w_n230_2(.douta(w_n230_2[0]),.doutb(w_n230_2[1]),.din(w_n230_0[1]));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.din(n231));
	jspl3 jspl3_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.doutc(w_n232_0[2]),.din(n232));
	jspl3 jspl3_w_n232_1(.douta(w_n232_1[0]),.doutb(w_n232_1[1]),.doutc(w_n232_1[2]),.din(w_n232_0[0]));
	jspl3 jspl3_w_n232_2(.douta(w_n232_2[0]),.doutb(w_n232_2[1]),.doutc(w_n232_2[2]),.din(w_n232_0[1]));
	jspl jspl_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.din(n234));
	jspl3 jspl3_w_n235_0(.douta(w_n235_0[0]),.doutb(w_n235_0[1]),.doutc(w_n235_0[2]),.din(n235));
	jspl3 jspl3_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.doutc(w_n236_0[2]),.din(n236));
	jspl3 jspl3_w_n236_1(.douta(w_n236_1[0]),.doutb(w_n236_1[1]),.doutc(w_n236_1[2]),.din(w_n236_0[0]));
	jspl3 jspl3_w_n236_2(.douta(w_n236_2[0]),.doutb(w_n236_2[1]),.doutc(w_n236_2[2]),.din(w_n236_0[1]));
	jspl jspl_w_n236_3(.douta(w_n236_3[0]),.doutb(w_n236_3[1]),.din(w_n236_0[2]));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(n239));
	jspl3 jspl3_w_n240_0(.douta(w_n240_0[0]),.doutb(w_n240_0[1]),.doutc(w_n240_0[2]),.din(n240));
	jspl3 jspl3_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.doutc(w_n241_0[2]),.din(n241));
	jspl jspl_w_n241_1(.douta(w_n241_1[0]),.doutb(w_n241_1[1]),.din(w_n241_0[0]));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl3 jspl3_w_n243_1(.douta(w_n243_1[0]),.doutb(w_n243_1[1]),.doutc(w_n243_1[2]),.din(w_n243_0[0]));
	jspl3 jspl3_w_n243_2(.douta(w_n243_2[0]),.doutb(w_n243_2[1]),.doutc(w_n243_2[2]),.din(w_n243_0[1]));
	jspl3 jspl3_w_n243_3(.douta(w_n243_3[0]),.doutb(w_n243_3[1]),.doutc(w_n243_3[2]),.din(w_n243_0[2]));
	jspl3 jspl3_w_n243_4(.douta(w_n243_4[0]),.doutb(w_n243_4[1]),.doutc(w_n243_4[2]),.din(w_n243_1[0]));
	jspl jspl_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.din(n246));
	jspl3 jspl3_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.doutc(w_n247_0[2]),.din(n247));
	jspl3 jspl3_w_n247_1(.douta(w_n247_1[0]),.doutb(w_n247_1[1]),.doutc(w_n247_1[2]),.din(w_n247_0[0]));
	jspl3 jspl3_w_n247_2(.douta(w_n247_2[0]),.doutb(w_n247_2[1]),.doutc(w_n247_2[2]),.din(w_n247_0[1]));
	jspl3 jspl3_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.doutc(w_n249_0[2]),.din(n249));
	jspl3 jspl3_w_n249_1(.douta(w_n249_1[0]),.doutb(w_n249_1[1]),.doutc(w_n249_1[2]),.din(w_n249_0[0]));
	jspl jspl_w_n249_2(.douta(w_n249_2[0]),.doutb(w_n249_2[1]),.din(w_n249_0[1]));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl3 jspl3_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.doutc(w_n251_0[2]),.din(n251));
	jspl3 jspl3_w_n251_1(.douta(w_n251_1[0]),.doutb(w_n251_1[1]),.doutc(w_n251_1[2]),.din(w_n251_0[0]));
	jspl3 jspl3_w_n251_2(.douta(w_n251_2[0]),.doutb(w_n251_2[1]),.doutc(w_n251_2[2]),.din(w_n251_0[1]));
	jspl jspl_w_n251_3(.douta(w_n251_3[0]),.doutb(w_n251_3[1]),.din(w_n251_0[2]));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl3 jspl3_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.doutc(w_n254_1[2]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n254_2(.douta(w_n254_2[0]),.doutb(w_n254_2[1]),.doutc(w_n254_2[2]),.din(w_n254_0[1]));
	jspl jspl_w_n254_3(.douta(w_n254_3[0]),.doutb(w_n254_3[1]),.din(w_n254_0[2]));
	jspl3 jspl3_w_n256_0(.douta(w_n256_0[0]),.doutb(w_n256_0[1]),.doutc(w_n256_0[2]),.din(n256));
	jspl3 jspl3_w_n256_1(.douta(w_n256_1[0]),.doutb(w_n256_1[1]),.doutc(w_n256_1[2]),.din(w_n256_0[0]));
	jspl jspl_w_n256_2(.douta(w_n256_2[0]),.doutb(w_n256_2[1]),.din(w_n256_0[1]));
	jspl3 jspl3_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.doutc(w_n259_0[2]),.din(n259));
	jspl3 jspl3_w_n259_1(.douta(w_n259_1[0]),.doutb(w_n259_1[1]),.doutc(w_n259_1[2]),.din(w_n259_0[0]));
	jspl3 jspl3_w_n259_2(.douta(w_n259_2[0]),.doutb(w_n259_2[1]),.doutc(w_n259_2[2]),.din(w_n259_0[1]));
	jspl jspl_w_n259_3(.douta(w_n259_3[0]),.doutb(w_n259_3[1]),.din(w_n259_0[2]));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl3 jspl3_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.doutc(w_n261_0[2]),.din(n261));
	jspl3 jspl3_w_n261_1(.douta(w_n261_1[0]),.doutb(w_n261_1[1]),.doutc(w_n261_1[2]),.din(w_n261_0[0]));
	jspl3 jspl3_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.doutc(w_n262_0[2]),.din(n262));
	jspl3 jspl3_w_n262_1(.douta(w_n262_1[0]),.doutb(w_n262_1[1]),.doutc(w_n262_1[2]),.din(w_n262_0[0]));
	jspl3 jspl3_w_n262_2(.douta(w_n262_2[0]),.doutb(w_n262_2[1]),.doutc(w_n262_2[2]),.din(w_n262_0[1]));
	jspl3 jspl3_w_n262_3(.douta(w_n262_3[0]),.doutb(w_n262_3[1]),.doutc(w_n262_3[2]),.din(w_n262_0[2]));
	jspl jspl_w_n263_0(.douta(w_n263_0[0]),.doutb(w_n263_0[1]),.din(n263));
	jspl3 jspl3_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.doutc(w_n264_0[2]),.din(n264));
	jspl3 jspl3_w_n264_1(.douta(w_n264_1[0]),.doutb(w_n264_1[1]),.doutc(w_n264_1[2]),.din(w_n264_0[0]));
	jspl3 jspl3_w_n264_2(.douta(w_n264_2[0]),.doutb(w_n264_2[1]),.doutc(w_n264_2[2]),.din(w_n264_0[1]));
	jspl3 jspl3_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.doutc(w_n265_0[2]),.din(n265));
	jspl3 jspl3_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.doutc(w_n266_0[2]),.din(n266));
	jspl jspl_w_n266_1(.douta(w_n266_1[0]),.doutb(w_n266_1[1]),.din(w_n266_0[0]));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.doutc(w_n267_0[2]),.din(n267));
	jspl3 jspl3_w_n267_1(.douta(w_n267_1[0]),.doutb(w_n267_1[1]),.doutc(w_n267_1[2]),.din(w_n267_0[0]));
	jspl3 jspl3_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.doutc(w_n268_0[2]),.din(n268));
	jspl3 jspl3_w_n268_1(.douta(w_n268_1[0]),.doutb(w_n268_1[1]),.doutc(w_n268_1[2]),.din(w_n268_0[0]));
	jspl3 jspl3_w_n268_2(.douta(w_n268_2[0]),.doutb(w_n268_2[1]),.doutc(w_n268_2[2]),.din(w_n268_0[1]));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.doutc(w_n270_0[2]),.din(n270));
	jspl3 jspl3_w_n270_1(.douta(w_n270_1[0]),.doutb(w_n270_1[1]),.doutc(w_n270_1[2]),.din(w_n270_0[0]));
	jspl3 jspl3_w_n270_2(.douta(w_n270_2[0]),.doutb(w_n270_2[1]),.doutc(w_n270_2[2]),.din(w_n270_0[1]));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl3 jspl3_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.doutc(w_n276_0[2]),.din(n276));
	jspl3 jspl3_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.doutc(w_n277_0[2]),.din(n277));
	jspl3 jspl3_w_n277_1(.douta(w_n277_1[0]),.doutb(w_n277_1[1]),.doutc(w_n277_1[2]),.din(w_n277_0[0]));
	jspl3 jspl3_w_n277_2(.douta(w_n277_2[0]),.doutb(w_n277_2[1]),.doutc(w_n277_2[2]),.din(w_n277_0[1]));
	jspl jspl_w_n277_3(.douta(w_n277_3[0]),.doutb(w_n277_3[1]),.din(w_n277_0[2]));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(n278));
	jspl3 jspl3_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.doutc(w_n279_0[2]),.din(n279));
	jspl3 jspl3_w_n279_1(.douta(w_n279_1[0]),.doutb(w_n279_1[1]),.doutc(w_n279_1[2]),.din(w_n279_0[0]));
	jspl jspl_w_n279_2(.douta(w_n279_2[0]),.doutb(w_n279_2[1]),.din(w_n279_0[1]));
	jspl3 jspl3_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.doutc(w_n280_0[2]),.din(n280));
	jspl jspl_w_n280_1(.douta(w_n280_1[0]),.doutb(w_n280_1[1]),.din(w_n280_0[0]));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.din(n281));
	jspl3 jspl3_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.doutc(w_n282_0[2]),.din(n282));
	jspl3 jspl3_w_n282_1(.douta(w_n282_1[0]),.doutb(w_n282_1[1]),.doutc(w_n282_1[2]),.din(w_n282_0[0]));
	jspl3 jspl3_w_n282_2(.douta(w_n282_2[0]),.doutb(w_n282_2[1]),.doutc(w_n282_2[2]),.din(w_n282_0[1]));
	jspl jspl_w_n282_3(.douta(w_n282_3[0]),.doutb(w_n282_3[1]),.din(w_n282_0[2]));
	jspl3 jspl3_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.doutc(w_n283_0[2]),.din(n283));
	jspl3 jspl3_w_n283_1(.douta(w_n283_1[0]),.doutb(w_n283_1[1]),.doutc(w_n283_1[2]),.din(w_n283_0[0]));
	jspl3 jspl3_w_n283_2(.douta(w_n283_2[0]),.doutb(w_n283_2[1]),.doutc(w_n283_2[2]),.din(w_n283_0[1]));
	jspl jspl_w_n283_3(.douta(w_n283_3[0]),.doutb(w_n283_3[1]),.din(w_n283_0[2]));
	jspl jspl_w_n284_0(.douta(w_n284_0[0]),.doutb(w_n284_0[1]),.din(n284));
	jspl3 jspl3_w_n285_0(.douta(w_n285_0[0]),.doutb(w_n285_0[1]),.doutc(w_n285_0[2]),.din(n285));
	jspl3 jspl3_w_n285_1(.douta(w_n285_1[0]),.doutb(w_n285_1[1]),.doutc(w_n285_1[2]),.din(w_n285_0[0]));
	jspl jspl_w_n285_2(.douta(w_n285_2[0]),.doutb(w_n285_2[1]),.din(w_n285_0[1]));
	jspl3 jspl3_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.doutc(w_n286_0[2]),.din(n286));
	jspl3 jspl3_w_n286_1(.douta(w_n286_1[0]),.doutb(w_n286_1[1]),.doutc(w_n286_1[2]),.din(w_n286_0[0]));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n288_1(.douta(w_n288_1[0]),.doutb(w_n288_1[1]),.din(w_n288_0[0]));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(n290));
	jspl3 jspl3_w_n291_0(.douta(w_n291_0[0]),.doutb(w_n291_0[1]),.doutc(w_n291_0[2]),.din(n291));
	jspl3 jspl3_w_n291_1(.douta(w_n291_1[0]),.doutb(w_n291_1[1]),.doutc(w_n291_1[2]),.din(w_n291_0[0]));
	jspl jspl_w_n291_2(.douta(w_n291_2[0]),.doutb(w_n291_2[1]),.din(w_n291_0[1]));
	jspl3 jspl3_w_n294_0(.douta(w_n294_0[0]),.doutb(w_n294_0[1]),.doutc(w_n294_0[2]),.din(n294));
	jspl3 jspl3_w_n294_1(.douta(w_n294_1[0]),.doutb(w_n294_1[1]),.doutc(w_n294_1[2]),.din(w_n294_0[0]));
	jspl3 jspl3_w_n294_2(.douta(w_n294_2[0]),.doutb(w_n294_2[1]),.doutc(w_n294_2[2]),.din(w_n294_0[1]));
	jspl jspl_w_n294_3(.douta(w_n294_3[0]),.doutb(w_n294_3[1]),.din(w_n294_0[2]));
	jspl3 jspl3_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.doutc(w_n295_0[2]),.din(n295));
	jspl3 jspl3_w_n295_1(.douta(w_n295_1[0]),.doutb(w_n295_1[1]),.doutc(w_n295_1[2]),.din(w_n295_0[0]));
	jspl3 jspl3_w_n295_2(.douta(w_n295_2[0]),.doutb(w_n295_2[1]),.doutc(w_n295_2[2]),.din(w_n295_0[1]));
	jspl3 jspl3_w_n295_3(.douta(w_n295_3[0]),.doutb(w_n295_3[1]),.doutc(w_n295_3[2]),.din(w_n295_0[2]));
	jspl3 jspl3_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.doutc(w_n298_0[2]),.din(n298));
	jspl3 jspl3_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.doutc(w_n299_0[2]),.din(n299));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_n300_0[1]),.din(n300));
	jspl3 jspl3_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.doutc(w_n301_0[2]),.din(n301));
	jspl3 jspl3_w_n301_1(.douta(w_n301_1[0]),.doutb(w_n301_1[1]),.doutc(w_n301_1[2]),.din(w_n301_0[0]));
	jspl3 jspl3_w_n301_2(.douta(w_n301_2[0]),.doutb(w_n301_2[1]),.doutc(w_n301_2[2]),.din(w_n301_0[1]));
	jspl3 jspl3_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.doutc(w_n303_0[2]),.din(n303));
	jspl3 jspl3_w_n303_1(.douta(w_n303_1[0]),.doutb(w_n303_1[1]),.doutc(w_n303_1[2]),.din(w_n303_0[0]));
	jspl3 jspl3_w_n303_2(.douta(w_n303_2[0]),.doutb(w_n303_2[1]),.doutc(w_n303_2[2]),.din(w_n303_0[1]));
	jspl3 jspl3_w_n303_3(.douta(w_n303_3[0]),.doutb(w_n303_3[1]),.doutc(w_n303_3[2]),.din(w_n303_0[2]));
	jspl jspl_w_n303_4(.douta(w_n303_4[0]),.doutb(w_n303_4[1]),.din(w_n303_1[0]));
	jspl3 jspl3_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.doutc(w_n304_0[2]),.din(n304));
	jspl3 jspl3_w_n304_1(.douta(w_n304_1[0]),.doutb(w_n304_1[1]),.doutc(w_n304_1[2]),.din(w_n304_0[0]));
	jspl3 jspl3_w_n304_2(.douta(w_n304_2[0]),.doutb(w_n304_2[1]),.doutc(w_n304_2[2]),.din(w_n304_0[1]));
	jspl jspl_w_n304_3(.douta(w_n304_3[0]),.doutb(w_n304_3[1]),.din(w_n304_0[2]));
	jspl3 jspl3_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.doutc(w_n305_0[2]),.din(n305));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(n309));
	jspl3 jspl3_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.doutc(w_n310_0[2]),.din(n310));
	jspl3 jspl3_w_n310_1(.douta(w_n310_1[0]),.doutb(w_n310_1[1]),.doutc(w_n310_1[2]),.din(w_n310_0[0]));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.doutc(w_n312_0[2]),.din(n312));
	jspl3 jspl3_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.doutc(w_n312_1[2]),.din(w_n312_0[0]));
	jspl3 jspl3_w_n312_2(.douta(w_n312_2[0]),.doutb(w_n312_2[1]),.doutc(w_n312_2[2]),.din(w_n312_0[1]));
	jspl3 jspl3_w_n312_3(.douta(w_n312_3[0]),.doutb(w_n312_3[1]),.doutc(w_n312_3[2]),.din(w_n312_0[2]));
	jspl3 jspl3_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.doutc(w_n314_0[2]),.din(n314));
	jspl jspl_w_n314_1(.douta(w_n314_1[0]),.doutb(w_n314_1[1]),.din(w_n314_0[0]));
	jspl3 jspl3_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.doutc(w_n315_0[2]),.din(n315));
	jspl jspl_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.din(n319));
	jspl3 jspl3_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.doutc(w_n320_0[2]),.din(n320));
	jspl3 jspl3_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.doutc(w_n321_0[2]),.din(n321));
	jspl jspl_w_n321_1(.douta(w_n321_1[0]),.doutb(w_n321_1[1]),.din(w_n321_0[0]));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl3 jspl3_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.doutc(w_n323_0[2]),.din(n323));
	jspl3 jspl3_w_n323_1(.douta(w_n323_1[0]),.doutb(w_n323_1[1]),.doutc(w_n323_1[2]),.din(w_n323_0[0]));
	jspl3 jspl3_w_n323_2(.douta(w_n323_2[0]),.doutb(w_n323_2[1]),.doutc(w_n323_2[2]),.din(w_n323_0[1]));
	jspl jspl_w_n323_3(.douta(w_n323_3[0]),.doutb(w_n323_3[1]),.din(w_n323_0[2]));
	jspl3 jspl3_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.doutc(w_n324_0[2]),.din(n324));
	jspl jspl_w_n324_1(.douta(w_n324_1[0]),.doutb(w_n324_1[1]),.din(w_n324_0[0]));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.din(n326));
	jspl3 jspl3_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.doutc(w_n327_0[2]),.din(n327));
	jspl3 jspl3_w_n327_1(.douta(w_n327_1[0]),.doutb(w_n327_1[1]),.doutc(w_n327_1[2]),.din(w_n327_0[0]));
	jspl3 jspl3_w_n327_2(.douta(w_n327_2[0]),.doutb(w_n327_2[1]),.doutc(w_n327_2[2]),.din(w_n327_0[1]));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl3 jspl3_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.doutc(w_n334_0[2]),.din(n334));
	jspl3 jspl3_w_n334_1(.douta(w_n334_1[0]),.doutb(w_n334_1[1]),.doutc(w_n334_1[2]),.din(w_n334_0[0]));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.doutc(w_n335_1[2]),.din(w_n335_0[0]));
	jspl3 jspl3_w_n335_2(.douta(w_n335_2[0]),.doutb(w_n335_2[1]),.doutc(w_n335_2[2]),.din(w_n335_0[1]));
	jspl3 jspl3_w_n335_3(.douta(w_n335_3[0]),.doutb(w_n335_3[1]),.doutc(w_n335_3[2]),.din(w_n335_0[2]));
	jspl3 jspl3_w_n335_4(.douta(w_n335_4[0]),.doutb(w_n335_4[1]),.doutc(w_n335_4[2]),.din(w_n335_1[0]));
	jspl3 jspl3_w_n335_5(.douta(w_n335_5[0]),.doutb(w_n335_5[1]),.doutc(w_n335_5[2]),.din(w_n335_1[1]));
	jspl3 jspl3_w_n335_6(.douta(w_n335_6[0]),.doutb(w_n335_6[1]),.doutc(w_n335_6[2]),.din(w_n335_1[2]));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl3 jspl3_w_n337_0(.douta(w_n337_0[0]),.doutb(w_n337_0[1]),.doutc(w_n337_0[2]),.din(n337));
	jspl3 jspl3_w_n337_1(.douta(w_n337_1[0]),.doutb(w_n337_1[1]),.doutc(w_n337_1[2]),.din(w_n337_0[0]));
	jspl3 jspl3_w_n337_2(.douta(w_n337_2[0]),.doutb(w_n337_2[1]),.doutc(w_n337_2[2]),.din(w_n337_0[1]));
	jspl3 jspl3_w_n337_3(.douta(w_n337_3[0]),.doutb(w_n337_3[1]),.doutc(w_n337_3[2]),.din(w_n337_0[2]));
	jspl3 jspl3_w_n337_4(.douta(w_n337_4[0]),.doutb(w_n337_4[1]),.doutc(w_n337_4[2]),.din(w_n337_1[0]));
	jspl jspl_w_n337_5(.douta(w_n337_5[0]),.doutb(w_n337_5[1]),.din(w_n337_1[1]));
	jspl3 jspl3_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.doutc(w_n338_0[2]),.din(n338));
	jspl jspl_w_n338_1(.douta(w_n338_1[0]),.doutb(w_n338_1[1]),.din(w_n338_0[0]));
	jspl3 jspl3_w_n339_0(.douta(w_n339_0[0]),.doutb(w_n339_0[1]),.doutc(w_n339_0[2]),.din(n339));
	jspl3 jspl3_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.doutc(w_n340_0[2]),.din(n340));
	jspl3 jspl3_w_n340_1(.douta(w_n340_1[0]),.doutb(w_n340_1[1]),.doutc(w_n340_1[2]),.din(w_n340_0[0]));
	jspl jspl_w_n340_2(.douta(w_n340_2[0]),.doutb(w_n340_2[1]),.din(w_n340_0[1]));
	jspl3 jspl3_w_n341_0(.douta(w_n341_0[0]),.doutb(w_n341_0[1]),.doutc(w_n341_0[2]),.din(n341));
	jspl3 jspl3_w_n341_1(.douta(w_n341_1[0]),.doutb(w_n341_1[1]),.doutc(w_n341_1[2]),.din(w_n341_0[0]));
	jspl3 jspl3_w_n341_2(.douta(w_n341_2[0]),.doutb(w_n341_2[1]),.doutc(w_n341_2[2]),.din(w_n341_0[1]));
	jspl3 jspl3_w_n341_3(.douta(w_n341_3[0]),.doutb(w_n341_3[1]),.doutc(w_n341_3[2]),.din(w_n341_0[2]));
	jspl jspl_w_n341_4(.douta(w_n341_4[0]),.doutb(w_n341_4[1]),.din(w_n341_1[0]));
	jspl jspl_w_n342_0(.douta(w_n342_0[0]),.doutb(w_n342_0[1]),.din(n342));
	jspl3 jspl3_w_n343_0(.douta(w_n343_0[0]),.doutb(w_n343_0[1]),.doutc(w_n343_0[2]),.din(n343));
	jspl3 jspl3_w_n343_1(.douta(w_n343_1[0]),.doutb(w_n343_1[1]),.doutc(w_n343_1[2]),.din(w_n343_0[0]));
	jspl jspl_w_n343_2(.douta(w_n343_2[0]),.doutb(w_n343_2[1]),.din(w_n343_0[1]));
	jspl3 jspl3_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.doutc(w_n345_0[2]),.din(n345));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl3 jspl3_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.doutc(w_n346_1[2]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n346_2(.douta(w_n346_2[0]),.doutb(w_n346_2[1]),.doutc(w_n346_2[2]),.din(w_n346_0[1]));
	jspl3 jspl3_w_n346_3(.douta(w_n346_3[0]),.doutb(w_n346_3[1]),.doutc(w_n346_3[2]),.din(w_n346_0[2]));
	jspl3 jspl3_w_n346_4(.douta(w_n346_4[0]),.doutb(w_n346_4[1]),.doutc(w_n346_4[2]),.din(w_n346_1[0]));
	jspl3 jspl3_w_n346_5(.douta(w_n346_5[0]),.doutb(w_n346_5[1]),.doutc(w_n346_5[2]),.din(w_n346_1[1]));
	jspl3 jspl3_w_n346_6(.douta(w_n346_6[0]),.doutb(w_n346_6[1]),.doutc(w_n346_6[2]),.din(w_n346_1[2]));
	jspl jspl_w_n346_7(.douta(w_n346_7[0]),.doutb(w_n346_7[1]),.din(w_n346_2[0]));
	jspl3 jspl3_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.doutc(w_n348_0[2]),.din(n348));
	jspl3 jspl3_w_n348_1(.douta(w_n348_1[0]),.doutb(w_n348_1[1]),.doutc(w_n348_1[2]),.din(w_n348_0[0]));
	jspl3 jspl3_w_n348_2(.douta(w_n348_2[0]),.doutb(w_n348_2[1]),.doutc(w_n348_2[2]),.din(w_n348_0[1]));
	jspl3 jspl3_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.doutc(w_n349_0[2]),.din(n349));
	jspl3 jspl3_w_n349_1(.douta(w_n349_1[0]),.doutb(w_n349_1[1]),.doutc(w_n349_1[2]),.din(w_n349_0[0]));
	jspl3 jspl3_w_n349_2(.douta(w_n349_2[0]),.doutb(w_n349_2[1]),.doutc(w_n349_2[2]),.din(w_n349_0[1]));
	jspl3 jspl3_w_n349_3(.douta(w_n349_3[0]),.doutb(w_n349_3[1]),.doutc(w_n349_3[2]),.din(w_n349_0[2]));
	jspl3 jspl3_w_n349_4(.douta(w_n349_4[0]),.doutb(w_n349_4[1]),.doutc(w_n349_4[2]),.din(w_n349_1[0]));
	jspl3 jspl3_w_n349_5(.douta(w_n349_5[0]),.doutb(w_n349_5[1]),.doutc(w_n349_5[2]),.din(w_n349_1[1]));
	jspl3 jspl3_w_n349_6(.douta(w_n349_6[0]),.doutb(w_n349_6[1]),.doutc(w_n349_6[2]),.din(w_n349_1[2]));
	jspl3 jspl3_w_n351_0(.douta(w_n351_0[0]),.doutb(w_n351_0[1]),.doutc(w_n351_0[2]),.din(n351));
	jspl3 jspl3_w_n351_1(.douta(w_n351_1[0]),.doutb(w_n351_1[1]),.doutc(w_n351_1[2]),.din(w_n351_0[0]));
	jspl jspl_w_n351_2(.douta(w_n351_2[0]),.doutb(w_n351_2[1]),.din(w_n351_0[1]));
	jspl3 jspl3_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.doutc(w_n353_0[2]),.din(n353));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_n354_0[2]),.din(n354));
	jspl3 jspl3_w_n354_1(.douta(w_n354_1[0]),.doutb(w_n354_1[1]),.doutc(w_n354_1[2]),.din(w_n354_0[0]));
	jspl3 jspl3_w_n354_2(.douta(w_n354_2[0]),.doutb(w_n354_2[1]),.doutc(w_n354_2[2]),.din(w_n354_0[1]));
	jspl3 jspl3_w_n354_3(.douta(w_n354_3[0]),.doutb(w_n354_3[1]),.doutc(w_n354_3[2]),.din(w_n354_0[2]));
	jspl jspl_w_n354_4(.douta(w_n354_4[0]),.doutb(w_n354_4[1]),.din(w_n354_1[0]));
	jspl jspl_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.din(n355));
	jspl3 jspl3_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.doutc(w_n356_0[2]),.din(n356));
	jspl3 jspl3_w_n356_1(.douta(w_n356_1[0]),.doutb(w_n356_1[1]),.doutc(w_n356_1[2]),.din(w_n356_0[0]));
	jspl3 jspl3_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.doutc(w_n358_0[2]),.din(n358));
	jspl3 jspl3_w_n358_1(.douta(w_n358_1[0]),.doutb(w_n358_1[1]),.doutc(w_n358_1[2]),.din(w_n358_0[0]));
	jspl jspl_w_n358_2(.douta(w_n358_2[0]),.doutb(w_n358_2[1]),.din(w_n358_0[1]));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.doutc(w_n363_0[2]),.din(n363));
	jspl3 jspl3_w_n363_1(.douta(w_n363_1[0]),.doutb(w_n363_1[1]),.doutc(w_n363_1[2]),.din(w_n363_0[0]));
	jspl jspl_w_n363_2(.douta(w_n363_2[0]),.doutb(w_n363_2[1]),.din(w_n363_0[1]));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl3 jspl3_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.doutc(w_n365_0[2]),.din(n365));
	jspl3 jspl3_w_n365_1(.douta(w_n365_1[0]),.doutb(w_n365_1[1]),.doutc(w_n365_1[2]),.din(w_n365_0[0]));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(n366));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl3 jspl3_w_n367_1(.douta(w_n367_1[0]),.doutb(w_n367_1[1]),.doutc(w_n367_1[2]),.din(w_n367_0[0]));
	jspl3 jspl3_w_n367_2(.douta(w_n367_2[0]),.doutb(w_n367_2[1]),.doutc(w_n367_2[2]),.din(w_n367_0[1]));
	jspl3 jspl3_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.doutc(w_n368_0[2]),.din(n368));
	jspl3 jspl3_w_n368_1(.douta(w_n368_1[0]),.doutb(w_n368_1[1]),.doutc(w_n368_1[2]),.din(w_n368_0[0]));
	jspl3 jspl3_w_n368_2(.douta(w_n368_2[0]),.doutb(w_n368_2[1]),.doutc(w_n368_2[2]),.din(w_n368_0[1]));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl3 jspl3_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.doutc(w_n370_0[2]),.din(n370));
	jspl3 jspl3_w_n370_1(.douta(w_n370_1[0]),.doutb(w_n370_1[1]),.doutc(w_n370_1[2]),.din(w_n370_0[0]));
	jspl jspl_w_n370_2(.douta(w_n370_2[0]),.doutb(w_n370_2[1]),.din(w_n370_0[1]));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.doutc(w_n372_0[2]),.din(n372));
	jspl3 jspl3_w_n372_1(.douta(w_n372_1[0]),.doutb(w_n372_1[1]),.doutc(w_n372_1[2]),.din(w_n372_0[0]));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl3 jspl3_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.doutc(w_n374_0[2]),.din(n374));
	jspl3 jspl3_w_n374_1(.douta(w_n374_1[0]),.doutb(w_n374_1[1]),.doutc(w_n374_1[2]),.din(w_n374_0[0]));
	jspl3 jspl3_w_n374_2(.douta(w_n374_2[0]),.doutb(w_n374_2[1]),.doutc(w_n374_2[2]),.din(w_n374_0[1]));
	jspl jspl_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.din(n378));
	jspl3 jspl3_w_n379_0(.douta(w_n379_0[0]),.doutb(w_n379_0[1]),.doutc(w_n379_0[2]),.din(n379));
	jspl3 jspl3_w_n379_1(.douta(w_n379_1[0]),.doutb(w_n379_1[1]),.doutc(w_n379_1[2]),.din(w_n379_0[0]));
	jspl3 jspl3_w_n380_0(.douta(w_n380_0[0]),.doutb(w_n380_0[1]),.doutc(w_n380_0[2]),.din(n380));
	jspl jspl_w_n380_1(.douta(w_n380_1[0]),.doutb(w_n380_1[1]),.din(w_n380_0[0]));
	jspl3 jspl3_w_n381_0(.douta(w_n381_0[0]),.doutb(w_n381_0[1]),.doutc(w_n381_0[2]),.din(n381));
	jspl3 jspl3_w_n381_1(.douta(w_n381_1[0]),.doutb(w_n381_1[1]),.doutc(w_n381_1[2]),.din(w_n381_0[0]));
	jspl3 jspl3_w_n381_2(.douta(w_n381_2[0]),.doutb(w_n381_2[1]),.doutc(w_n381_2[2]),.din(w_n381_0[1]));
	jspl jspl_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.din(n382));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n383_1(.douta(w_n383_1[0]),.doutb(w_n383_1[1]),.doutc(w_n383_1[2]),.din(w_n383_0[0]));
	jspl3 jspl3_w_n383_2(.douta(w_n383_2[0]),.doutb(w_n383_2[1]),.doutc(w_n383_2[2]),.din(w_n383_0[1]));
	jspl3 jspl3_w_n384_0(.douta(w_n384_0[0]),.doutb(w_n384_0[1]),.doutc(w_n384_0[2]),.din(n384));
	jspl jspl_w_n384_1(.douta(w_n384_1[0]),.doutb(w_n384_1[1]),.din(w_n384_0[0]));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl jspl_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl3 jspl3_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.doutc(w_n387_1[2]),.din(w_n387_0[0]));
	jspl jspl_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.din(n388));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.din(n389));
	jspl3 jspl3_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.doutc(w_n390_0[2]),.din(n390));
	jspl3 jspl3_w_n390_1(.douta(w_n390_1[0]),.doutb(w_n390_1[1]),.doutc(w_n390_1[2]),.din(w_n390_0[0]));
	jspl3 jspl3_w_n392_0(.douta(w_n392_0[0]),.doutb(w_n392_0[1]),.doutc(w_n392_0[2]),.din(n392));
	jspl3 jspl3_w_n395_0(.douta(w_n395_0[0]),.doutb(w_n395_0[1]),.doutc(w_n395_0[2]),.din(n395));
	jspl3 jspl3_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.doutc(w_n397_0[2]),.din(n397));
	jspl3 jspl3_w_n397_1(.douta(w_n397_1[0]),.doutb(w_n397_1[1]),.doutc(w_n397_1[2]),.din(w_n397_0[0]));
	jspl jspl_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.din(n398));
	jspl jspl_w_n399_0(.douta(w_n399_0[0]),.doutb(w_n399_0[1]),.din(n399));
	jspl jspl_w_n400_0(.douta(w_n400_0[0]),.doutb(w_n400_0[1]),.din(n400));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n401_1(.douta(w_n401_1[0]),.doutb(w_n401_1[1]),.doutc(w_n401_1[2]),.din(w_n401_0[0]));
	jspl3 jspl3_w_n401_2(.douta(w_n401_2[0]),.doutb(w_n401_2[1]),.doutc(w_n401_2[2]),.din(w_n401_0[1]));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n402_1(.douta(w_n402_1[0]),.doutb(w_n402_1[1]),.doutc(w_n402_1[2]),.din(w_n402_0[0]));
	jspl3 jspl3_w_n402_2(.douta(w_n402_2[0]),.doutb(w_n402_2[1]),.doutc(w_n402_2[2]),.din(w_n402_0[1]));
	jspl jspl_w_n402_3(.douta(w_n402_3[0]),.doutb(w_n402_3[1]),.din(w_n402_0[2]));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.doutc(w_n406_0[2]),.din(n406));
	jspl jspl_w_n406_1(.douta(w_n406_1[0]),.doutb(w_n406_1[1]),.din(w_n406_0[0]));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl jspl_w_n409_0(.douta(w_n409_0[0]),.doutb(w_n409_0[1]),.din(n409));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_n410_0[2]),.din(n410));
	jspl3 jspl3_w_n410_1(.douta(w_n410_1[0]),.doutb(w_n410_1[1]),.doutc(w_n410_1[2]),.din(w_n410_0[0]));
	jspl jspl_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.din(n411));
	jspl3 jspl3_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.doutc(w_n412_0[2]),.din(n412));
	jspl3 jspl3_w_n412_1(.douta(w_n412_1[0]),.doutb(w_n412_1[1]),.doutc(w_n412_1[2]),.din(w_n412_0[0]));
	jspl jspl_w_n412_2(.douta(w_n412_2[0]),.doutb(w_n412_2[1]),.din(w_n412_0[1]));
	jspl jspl_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.din(n413));
	jspl jspl_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.din(n414));
	jspl3 jspl3_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.doutc(w_n415_0[2]),.din(n415));
	jspl3 jspl3_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.doutc(w_n417_0[2]),.din(n417));
	jspl3 jspl3_w_n417_1(.douta(w_n417_1[0]),.doutb(w_n417_1[1]),.doutc(w_n417_1[2]),.din(w_n417_0[0]));
	jspl3 jspl3_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jspl3 jspl3_w_n420_1(.douta(w_n420_1[0]),.doutb(w_n420_1[1]),.doutc(w_n420_1[2]),.din(w_n420_0[0]));
	jspl jspl_w_n420_2(.douta(w_n420_2[0]),.doutb(w_n420_2[1]),.din(w_n420_0[1]));
	jspl3 jspl3_w_n421_0(.douta(w_n421_0[0]),.doutb(w_n421_0[1]),.doutc(w_n421_0[2]),.din(n421));
	jspl3 jspl3_w_n421_1(.douta(w_n421_1[0]),.doutb(w_n421_1[1]),.doutc(w_n421_1[2]),.din(w_n421_0[0]));
	jspl3 jspl3_w_n421_2(.douta(w_n421_2[0]),.doutb(w_n421_2[1]),.doutc(w_n421_2[2]),.din(w_n421_0[1]));
	jspl jspl_w_n421_3(.douta(w_n421_3[0]),.doutb(w_n421_3[1]),.din(w_n421_0[2]));
	jspl3 jspl3_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.doutc(w_n422_0[2]),.din(n422));
	jspl3 jspl3_w_n422_1(.douta(w_n422_1[0]),.doutb(w_n422_1[1]),.doutc(w_n422_1[2]),.din(w_n422_0[0]));
	jspl3 jspl3_w_n422_2(.douta(w_n422_2[0]),.doutb(w_n422_2[1]),.doutc(w_n422_2[2]),.din(w_n422_0[1]));
	jspl jspl_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.din(n424));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl3 jspl3_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.doutc(w_n426_0[2]),.din(n426));
	jspl3 jspl3_w_n426_1(.douta(w_n426_1[0]),.doutb(w_n426_1[1]),.doutc(w_n426_1[2]),.din(w_n426_0[0]));
	jspl3 jspl3_w_n426_2(.douta(w_n426_2[0]),.doutb(w_n426_2[1]),.doutc(w_n426_2[2]),.din(w_n426_0[1]));
	jspl3 jspl3_w_n426_3(.douta(w_n426_3[0]),.doutb(w_n426_3[1]),.doutc(w_n426_3[2]),.din(w_n426_0[2]));
	jspl3 jspl3_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.doutc(w_n427_0[2]),.din(n427));
	jspl3 jspl3_w_n427_1(.douta(w_n427_1[0]),.doutb(w_n427_1[1]),.doutc(w_n427_1[2]),.din(w_n427_0[0]));
	jspl3 jspl3_w_n427_2(.douta(w_n427_2[0]),.doutb(w_n427_2[1]),.doutc(w_n427_2[2]),.din(w_n427_0[1]));
	jspl jspl_w_n427_3(.douta(w_n427_3[0]),.doutb(w_n427_3[1]),.din(w_n427_0[2]));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.doutc(w_n428_0[2]),.din(n428));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl3 jspl3_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.doutc(w_n430_0[2]),.din(n430));
	jspl3 jspl3_w_n430_1(.douta(w_n430_1[0]),.doutb(w_n430_1[1]),.doutc(w_n430_1[2]),.din(w_n430_0[0]));
	jspl3 jspl3_w_n430_2(.douta(w_n430_2[0]),.doutb(w_n430_2[1]),.doutc(w_n430_2[2]),.din(w_n430_0[1]));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n436_1(.douta(w_n436_1[0]),.doutb(w_n436_1[1]),.doutc(w_n436_1[2]),.din(w_n436_0[0]));
	jspl3 jspl3_w_n436_2(.douta(w_n436_2[0]),.doutb(w_n436_2[1]),.doutc(w_n436_2[2]),.din(w_n436_0[1]));
	jspl3 jspl3_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.doutc(w_n437_0[2]),.din(n437));
	jspl3 jspl3_w_n437_1(.douta(w_n437_1[0]),.doutb(w_n437_1[1]),.doutc(w_n437_1[2]),.din(w_n437_0[0]));
	jspl jspl_w_n437_2(.douta(w_n437_2[0]),.doutb(w_n437_2[1]),.din(w_n437_0[1]));
	jspl jspl_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.din(n439));
	jspl3 jspl3_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.doutc(w_n440_0[2]),.din(n440));
	jspl3 jspl3_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.doutc(w_n441_0[2]),.din(n441));
	jspl3 jspl3_w_n441_1(.douta(w_n441_1[0]),.doutb(w_n441_1[1]),.doutc(w_n441_1[2]),.din(w_n441_0[0]));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n444_0(.douta(w_n444_0[0]),.doutb(w_n444_0[1]),.din(n444));
	jspl3 jspl3_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.doutc(w_n445_0[2]),.din(n445));
	jspl3 jspl3_w_n445_1(.douta(w_n445_1[0]),.doutb(w_n445_1[1]),.doutc(w_n445_1[2]),.din(w_n445_0[0]));
	jspl3 jspl3_w_n445_2(.douta(w_n445_2[0]),.doutb(w_n445_2[1]),.doutc(w_n445_2[2]),.din(w_n445_0[1]));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_n451_0[1]),.doutc(w_n451_0[2]),.din(n451));
	jspl3 jspl3_w_n451_1(.douta(w_n451_1[0]),.doutb(w_n451_1[1]),.doutc(w_n451_1[2]),.din(w_n451_0[0]));
	jspl3 jspl3_w_n451_2(.douta(w_n451_2[0]),.doutb(w_n451_2[1]),.doutc(w_n451_2[2]),.din(w_n451_0[1]));
	jspl jspl_w_n451_3(.douta(w_n451_3[0]),.doutb(w_n451_3[1]),.din(w_n451_0[2]));
	jspl jspl_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.din(n453));
	jspl3 jspl3_w_n454_0(.douta(w_n454_0[0]),.doutb(w_n454_0[1]),.doutc(w_n454_0[2]),.din(n454));
	jspl3 jspl3_w_n454_1(.douta(w_n454_1[0]),.doutb(w_n454_1[1]),.doutc(w_n454_1[2]),.din(w_n454_0[0]));
	jspl3 jspl3_w_n454_2(.douta(w_n454_2[0]),.doutb(w_n454_2[1]),.doutc(w_n454_2[2]),.din(w_n454_0[1]));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n458_0(.douta(w_n458_0[0]),.doutb(w_n458_0[1]),.doutc(w_n458_0[2]),.din(n458));
	jspl3 jspl3_w_n458_1(.douta(w_n458_1[0]),.doutb(w_n458_1[1]),.doutc(w_n458_1[2]),.din(w_n458_0[0]));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(n459));
	jspl jspl_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.din(n460));
	jspl3 jspl3_w_n461_0(.douta(w_n461_0[0]),.doutb(w_n461_0[1]),.doutc(w_n461_0[2]),.din(n461));
	jspl3 jspl3_w_n461_1(.douta(w_n461_1[0]),.doutb(w_n461_1[1]),.doutc(w_n461_1[2]),.din(w_n461_0[0]));
	jspl3 jspl3_w_n461_2(.douta(w_n461_2[0]),.doutb(w_n461_2[1]),.doutc(w_n461_2[2]),.din(w_n461_0[1]));
	jspl3 jspl3_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.doutc(w_n463_0[2]),.din(n463));
	jspl3 jspl3_w_n463_1(.douta(w_n463_1[0]),.doutb(w_n463_1[1]),.doutc(w_n463_1[2]),.din(w_n463_0[0]));
	jspl3 jspl3_w_n463_2(.douta(w_n463_2[0]),.doutb(w_n463_2[1]),.doutc(w_n463_2[2]),.din(w_n463_0[1]));
	jspl jspl_w_n463_3(.douta(w_n463_3[0]),.doutb(w_n463_3[1]),.din(w_n463_0[2]));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(n466));
	jspl3 jspl3_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.doutc(w_n467_0[2]),.din(n467));
	jspl jspl_w_n467_1(.douta(w_n467_1[0]),.doutb(w_n467_1[1]),.din(w_n467_0[0]));
	jspl jspl_w_n468_0(.douta(w_n468_0[0]),.doutb(w_n468_0[1]),.din(n468));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(n469));
	jspl3 jspl3_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.doutc(w_n470_0[2]),.din(n470));
	jspl3 jspl3_w_n470_1(.douta(w_n470_1[0]),.doutb(w_n470_1[1]),.doutc(w_n470_1[2]),.din(w_n470_0[0]));
	jspl jspl_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.din(n471));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.doutc(w_n473_0[2]),.din(n473));
	jspl3 jspl3_w_n473_1(.douta(w_n473_1[0]),.doutb(w_n473_1[1]),.doutc(w_n473_1[2]),.din(w_n473_0[0]));
	jspl jspl_w_n473_2(.douta(w_n473_2[0]),.doutb(w_n473_2[1]),.din(w_n473_0[1]));
	jspl3 jspl3_w_n475_0(.douta(w_n475_0[0]),.doutb(w_n475_0[1]),.doutc(w_n475_0[2]),.din(n475));
	jspl jspl_w_n475_1(.douta(w_n475_1[0]),.doutb(w_n475_1[1]),.din(w_n475_0[0]));
	jspl3 jspl3_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.doutc(w_n477_0[2]),.din(n477));
	jspl3 jspl3_w_n477_1(.douta(w_n477_1[0]),.doutb(w_n477_1[1]),.doutc(w_n477_1[2]),.din(w_n477_0[0]));
	jspl3 jspl3_w_n477_2(.douta(w_n477_2[0]),.doutb(w_n477_2[1]),.doutc(w_n477_2[2]),.din(w_n477_0[1]));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl3 jspl3_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.doutc(w_n479_0[2]),.din(n479));
	jspl3 jspl3_w_n479_1(.douta(w_n479_1[0]),.doutb(w_n479_1[1]),.doutc(w_n479_1[2]),.din(w_n479_0[0]));
	jspl jspl_w_n479_2(.douta(w_n479_2[0]),.doutb(w_n479_2[1]),.din(w_n479_0[1]));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(n482));
	jspl3 jspl3_w_n486_0(.douta(w_n486_0[0]),.doutb(w_n486_0[1]),.doutc(w_n486_0[2]),.din(n486));
	jspl jspl_w_n486_1(.douta(w_n486_1[0]),.doutb(w_n486_1[1]),.din(w_n486_0[0]));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl3 jspl3_w_n488_0(.douta(w_n488_0[0]),.doutb(w_n488_0[1]),.doutc(w_n488_0[2]),.din(n488));
	jspl3 jspl3_w_n488_1(.douta(w_n488_1[0]),.doutb(w_n488_1[1]),.doutc(w_n488_1[2]),.din(w_n488_0[0]));
	jspl jspl_w_n490_0(.douta(w_n490_0[0]),.doutb(w_n490_0[1]),.din(n490));
	jspl jspl_w_n491_0(.douta(w_n491_0[0]),.doutb(w_n491_0[1]),.din(n491));
	jspl jspl_w_n493_0(.douta(w_n493_0[0]),.doutb(w_n493_0[1]),.din(n493));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl3 jspl3_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.doutc(w_n497_0[2]),.din(n497));
	jspl jspl_w_n497_1(.douta(w_n497_1[0]),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl3 jspl3_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.doutc(w_n499_0[2]),.din(n499));
	jspl3 jspl3_w_n499_1(.douta(w_n499_1[0]),.doutb(w_n499_1[1]),.doutc(w_n499_1[2]),.din(w_n499_0[0]));
	jspl jspl_w_n500_0(.douta(w_n500_0[0]),.doutb(w_n500_0[1]),.din(n500));
	jspl3 jspl3_w_n501_0(.douta(w_n501_0[0]),.doutb(w_n501_0[1]),.doutc(w_n501_0[2]),.din(n501));
	jspl3 jspl3_w_n501_1(.douta(w_n501_1[0]),.doutb(w_n501_1[1]),.doutc(w_n501_1[2]),.din(w_n501_0[0]));
	jspl3 jspl3_w_n501_2(.douta(w_n501_2[0]),.doutb(w_n501_2[1]),.doutc(w_n501_2[2]),.din(w_n501_0[1]));
	jspl3 jspl3_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.doutc(w_n504_0[2]),.din(n504));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl3 jspl3_w_n506_0(.douta(w_n506_0[0]),.doutb(w_n506_0[1]),.doutc(w_n506_0[2]),.din(n506));
	jspl3 jspl3_w_n506_1(.douta(w_n506_1[0]),.doutb(w_n506_1[1]),.doutc(w_n506_1[2]),.din(w_n506_0[0]));
	jspl jspl_w_n506_2(.douta(w_n506_2[0]),.doutb(w_n506_2[1]),.din(w_n506_0[1]));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl jspl_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.din(w_n507_0[0]));
	jspl3 jspl3_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.doutc(w_n509_0[2]),.din(n509));
	jspl3 jspl3_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.doutc(w_n511_0[2]),.din(n511));
	jspl jspl_w_n511_1(.douta(w_n511_1[0]),.doutb(w_n511_1[1]),.din(w_n511_0[0]));
	jspl3 jspl3_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.doutc(w_n513_0[2]),.din(n513));
	jspl3 jspl3_w_n515_0(.douta(w_n515_0[0]),.doutb(w_n515_0[1]),.doutc(w_n515_0[2]),.din(n515));
	jspl3 jspl3_w_n515_1(.douta(w_n515_1[0]),.doutb(w_n515_1[1]),.doutc(w_n515_1[2]),.din(w_n515_0[0]));
	jspl3 jspl3_w_n515_2(.douta(w_n515_2[0]),.doutb(w_n515_2[1]),.doutc(w_n515_2[2]),.din(w_n515_0[1]));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(n519));
	jspl3 jspl3_w_n521_0(.douta(w_n521_0[0]),.doutb(w_n521_0[1]),.doutc(w_n521_0[2]),.din(n521));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.doutc(w_n523_0[2]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n525_0(.douta(w_n525_0[0]),.doutb(w_n525_0[1]),.din(n525));
	jspl jspl_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.din(n531));
	jspl3 jspl3_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.doutc(w_n532_0[2]),.din(n532));
	jspl3 jspl3_w_n532_1(.douta(w_n532_1[0]),.doutb(w_n532_1[1]),.doutc(w_n532_1[2]),.din(w_n532_0[0]));
	jspl3 jspl3_w_n532_2(.douta(w_n532_2[0]),.doutb(w_n532_2[1]),.doutc(w_n532_2[2]),.din(w_n532_0[1]));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl3 jspl3_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.doutc(w_n535_0[2]),.din(n535));
	jspl jspl_w_n535_1(.douta(w_n535_1[0]),.doutb(w_n535_1[1]),.din(w_n535_0[0]));
	jspl3 jspl3_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.doutc(w_n538_0[2]),.din(n538));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl3 jspl3_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.doutc(w_n543_0[2]),.din(n543));
	jspl jspl_w_n543_1(.douta(w_n543_1[0]),.doutb(w_n543_1[1]),.din(w_n543_0[0]));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl3 jspl3_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.doutc(w_n551_0[2]),.din(n551));
	jspl3 jspl3_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.doutc(w_n552_0[2]),.din(n552));
	jspl3 jspl3_w_n554_0(.douta(w_n554_0[0]),.doutb(w_n554_0[1]),.doutc(w_n554_0[2]),.din(n554));
	jspl jspl_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.din(n556));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl3 jspl3_w_n561_1(.douta(w_n561_1[0]),.doutb(w_n561_1[1]),.doutc(w_n561_1[2]),.din(w_n561_0[0]));
	jspl jspl_w_n561_2(.douta(w_n561_2[0]),.doutb(w_n561_2[1]),.din(w_n561_0[1]));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.doutc(w_n563_0[2]),.din(n563));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_n564_0[1]),.din(n564));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl jspl_w_n565_1(.douta(w_n565_1[0]),.doutb(w_n565_1[1]),.din(w_n565_0[0]));
	jspl3 jspl3_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.doutc(w_n568_0[2]),.din(n568));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_n571_0[2]),.din(n571));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(n577));
	jspl jspl_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.din(n578));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.doutc(w_n579_0[2]),.din(n579));
	jspl3 jspl3_w_n579_1(.douta(w_n579_1[0]),.doutb(w_n579_1[1]),.doutc(w_n579_1[2]),.din(w_n579_0[0]));
	jspl3 jspl3_w_n579_2(.douta(w_n579_2[0]),.doutb(w_n579_2[1]),.doutc(w_n579_2[2]),.din(w_n579_0[1]));
	jspl jspl_w_n580_0(.douta(w_n580_0[0]),.doutb(w_n580_0[1]),.din(n580));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl jspl_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.din(n586));
	jspl jspl_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.din(n587));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl jspl_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.din(n590));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl3 jspl3_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.doutc(w_n592_0[2]),.din(n592));
	jspl3 jspl3_w_n592_1(.douta(w_n592_1[0]),.doutb(w_n592_1[1]),.doutc(w_n592_1[2]),.din(w_n592_0[0]));
	jspl3 jspl3_w_n592_2(.douta(w_n592_2[0]),.doutb(w_n592_2[1]),.doutc(w_n592_2[2]),.din(w_n592_0[1]));
	jspl jspl_w_n592_3(.douta(w_n592_3[0]),.doutb(w_n592_3[1]),.din(w_n592_0[2]));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl3 jspl3_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.doutc(w_n594_0[2]),.din(n594));
	jspl3 jspl3_w_n594_1(.douta(w_n594_1[0]),.doutb(w_n594_1[1]),.doutc(w_n594_1[2]),.din(w_n594_0[0]));
	jspl3 jspl3_w_n594_2(.douta(w_n594_2[0]),.doutb(w_n594_2[1]),.doutc(w_n594_2[2]),.din(w_n594_0[1]));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.doutc(w_n595_0[2]),.din(n595));
	jspl3 jspl3_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl3 jspl3_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.doutc(w_n597_0[2]),.din(n597));
	jspl3 jspl3_w_n597_1(.douta(w_n597_1[0]),.doutb(w_n597_1[1]),.doutc(w_n597_1[2]),.din(w_n597_0[0]));
	jspl jspl_w_n597_2(.douta(w_n597_2[0]),.doutb(w_n597_2[1]),.din(w_n597_0[1]));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl3 jspl3_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.doutc(w_n604_0[2]),.din(n604));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl3 jspl3_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.doutc(w_n606_0[2]),.din(n606));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.doutc(w_n608_0[2]),.din(n608));
	jspl3 jspl3_w_n611_0(.douta(w_n611_0[0]),.doutb(w_n611_0[1]),.doutc(w_n611_0[2]),.din(n611));
	jspl jspl_w_n611_1(.douta(w_n611_1[0]),.doutb(w_n611_1[1]),.din(w_n611_0[0]));
	jspl3 jspl3_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.doutc(w_n612_0[2]),.din(n612));
	jspl3 jspl3_w_n612_1(.douta(w_n612_1[0]),.doutb(w_n612_1[1]),.doutc(w_n612_1[2]),.din(w_n612_0[0]));
	jspl3 jspl3_w_n612_2(.douta(w_n612_2[0]),.doutb(w_n612_2[1]),.doutc(w_n612_2[2]),.din(w_n612_0[1]));
	jspl3 jspl3_w_n612_3(.douta(w_n612_3[0]),.doutb(w_n612_3[1]),.doutc(w_n612_3[2]),.din(w_n612_0[2]));
	jspl3 jspl3_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.doutc(w_n614_0[2]),.din(n614));
	jspl3 jspl3_w_n614_1(.douta(w_n614_1[0]),.doutb(w_n614_1[1]),.doutc(w_n614_1[2]),.din(w_n614_0[0]));
	jspl3 jspl3_w_n614_2(.douta(w_n614_2[0]),.doutb(w_n614_2[1]),.doutc(w_n614_2[2]),.din(w_n614_0[1]));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n619_1(.douta(w_n619_1[0]),.doutb(w_n619_1[1]),.doutc(w_n619_1[2]),.din(w_n619_0[0]));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_n622_0[2]),.din(n622));
	jspl3 jspl3_w_n622_1(.douta(w_n622_1[0]),.doutb(w_n622_1[1]),.doutc(w_n622_1[2]),.din(w_n622_0[0]));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.doutc(w_n624_0[2]),.din(n624));
	jspl3 jspl3_w_n624_1(.douta(w_n624_1[0]),.doutb(w_n624_1[1]),.doutc(w_n624_1[2]),.din(w_n624_0[0]));
	jspl3 jspl3_w_n624_2(.douta(w_n624_2[0]),.doutb(w_n624_2[1]),.doutc(w_n624_2[2]),.din(w_n624_0[1]));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.din(n625));
	jspl3 jspl3_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.doutc(w_n626_0[2]),.din(n626));
	jspl jspl_w_n626_1(.douta(w_n626_1[0]),.doutb(w_n626_1[1]),.din(w_n626_0[0]));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl3 jspl3_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.doutc(w_n631_0[2]),.din(n631));
	jspl3 jspl3_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.doutc(w_n632_0[2]),.din(n632));
	jspl3 jspl3_w_n632_1(.douta(w_n632_1[0]),.doutb(w_n632_1[1]),.doutc(w_n632_1[2]),.din(w_n632_0[0]));
	jspl jspl_w_n632_2(.douta(w_n632_2[0]),.doutb(w_n632_2[1]),.din(w_n632_0[1]));
	jspl jspl_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.din(n633));
	jspl jspl_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.din(n636));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(n637));
	jspl3 jspl3_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.doutc(w_n638_0[2]),.din(n638));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl3 jspl3_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.doutc(w_n642_0[2]),.din(n642));
	jspl3 jspl3_w_n642_1(.douta(w_n642_1[0]),.doutb(w_n642_1[1]),.doutc(w_n642_1[2]),.din(w_n642_0[0]));
	jspl jspl_w_n643_0(.douta(w_n643_0[0]),.doutb(w_n643_0[1]),.din(n643));
	jspl jspl_w_n644_0(.douta(w_n644_0[0]),.doutb(w_n644_0[1]),.din(n644));
	jspl3 jspl3_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.doutc(w_n645_0[2]),.din(n645));
	jspl3 jspl3_w_n645_1(.douta(w_n645_1[0]),.doutb(w_n645_1[1]),.doutc(w_n645_1[2]),.din(w_n645_0[0]));
	jspl jspl_w_n645_2(.douta(w_n645_2[0]),.doutb(w_n645_2[1]),.din(w_n645_0[1]));
	jspl3 jspl3_w_n646_0(.douta(w_n646_0[0]),.doutb(w_n646_0[1]),.doutc(w_n646_0[2]),.din(n646));
	jspl jspl_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.din(n648));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.din(n651));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl3 jspl3_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.doutc(w_n662_0[2]),.din(n662));
	jspl3 jspl3_w_n662_1(.douta(w_n662_1[0]),.doutb(w_n662_1[1]),.doutc(w_n662_1[2]),.din(w_n662_0[0]));
	jspl3 jspl3_w_n662_2(.douta(w_n662_2[0]),.doutb(w_n662_2[1]),.doutc(w_n662_2[2]),.din(w_n662_0[1]));
	jspl3 jspl3_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.doutc(w_n664_0[2]),.din(n664));
	jspl3 jspl3_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.doutc(w_n665_0[2]),.din(n665));
	jspl3 jspl3_w_n665_1(.douta(w_n665_1[0]),.doutb(w_n665_1[1]),.doutc(w_n665_1[2]),.din(w_n665_0[0]));
	jspl3 jspl3_w_n665_2(.douta(w_n665_2[0]),.doutb(w_n665_2[1]),.doutc(w_n665_2[2]),.din(w_n665_0[1]));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(n667));
	jspl3 jspl3_w_n668_0(.douta(w_n668_0[0]),.doutb(w_n668_0[1]),.doutc(w_n668_0[2]),.din(n668));
	jspl3 jspl3_w_n668_1(.douta(w_n668_1[0]),.doutb(w_n668_1[1]),.doutc(w_n668_1[2]),.din(w_n668_0[0]));
	jspl3 jspl3_w_n668_2(.douta(w_n668_2[0]),.doutb(w_n668_2[1]),.doutc(w_n668_2[2]),.din(w_n668_0[1]));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(n669));
	jspl3 jspl3_w_n670_0(.douta(w_n670_0[0]),.doutb(w_n670_0[1]),.doutc(w_n670_0[2]),.din(n670));
	jspl3 jspl3_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.doutc(w_n675_0[2]),.din(n675));
	jspl3 jspl3_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.doutc(w_n676_0[2]),.din(n676));
	jspl jspl_w_n676_1(.douta(w_n676_1[0]),.doutb(w_n676_1[1]),.din(w_n676_0[0]));
	jspl3 jspl3_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.doutc(w_n677_0[2]),.din(n677));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl3 jspl3_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.doutc(w_n679_0[2]),.din(n679));
	jspl3 jspl3_w_n679_1(.douta(w_n679_1[0]),.doutb(w_n679_1[1]),.doutc(w_n679_1[2]),.din(w_n679_0[0]));
	jspl jspl_w_n679_2(.douta(w_n679_2[0]),.doutb(w_n679_2[1]),.din(w_n679_0[1]));
	jspl3 jspl3_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.doutc(w_n680_0[2]),.din(n680));
	jspl jspl_w_n680_1(.douta(w_n680_1[0]),.doutb(w_n680_1[1]),.din(w_n680_0[0]));
	jspl jspl_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.din(n681));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl3 jspl3_w_n688_0(.douta(w_n688_0[0]),.doutb(w_n688_0[1]),.doutc(w_n688_0[2]),.din(n688));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl3 jspl3_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.doutc(w_n691_0[2]),.din(n691));
	jspl3 jspl3_w_n691_1(.douta(w_n691_1[0]),.doutb(w_n691_1[1]),.doutc(w_n691_1[2]),.din(w_n691_0[0]));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl3 jspl3_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.doutc(w_n699_0[2]),.din(n699));
	jspl3 jspl3_w_n699_1(.douta(w_n699_1[0]),.doutb(w_n699_1[1]),.doutc(w_n699_1[2]),.din(w_n699_0[0]));
	jspl3 jspl3_w_n699_2(.douta(w_n699_2[0]),.doutb(w_n699_2[1]),.doutc(w_n699_2[2]),.din(w_n699_0[1]));
	jspl3 jspl3_w_n699_3(.douta(w_n699_3[0]),.doutb(w_n699_3[1]),.doutc(w_n699_3[2]),.din(w_n699_0[2]));
	jspl3 jspl3_w_n699_4(.douta(w_n699_4[0]),.doutb(w_n699_4[1]),.doutc(w_n699_4[2]),.din(w_n699_1[0]));
	jspl3 jspl3_w_n699_5(.douta(w_n699_5[0]),.doutb(w_n699_5[1]),.doutc(w_n699_5[2]),.din(w_n699_1[1]));
	jspl3 jspl3_w_n699_6(.douta(w_n699_6[0]),.doutb(w_n699_6[1]),.doutc(w_n699_6[2]),.din(w_n699_1[2]));
	jspl3 jspl3_w_n699_7(.douta(w_n699_7[0]),.doutb(w_n699_7[1]),.doutc(w_n699_7[2]),.din(w_n699_2[0]));
	jspl3 jspl3_w_n699_8(.douta(w_n699_8[0]),.doutb(w_n699_8[1]),.doutc(w_n699_8[2]),.din(w_n699_2[1]));
	jspl3 jspl3_w_n699_9(.douta(w_n699_9[0]),.doutb(w_n699_9[1]),.doutc(w_n699_9[2]),.din(w_n699_2[2]));
	jspl3 jspl3_w_n699_10(.douta(w_n699_10[0]),.doutb(w_n699_10[1]),.doutc(w_n699_10[2]),.din(w_n699_3[0]));
	jspl3 jspl3_w_n699_11(.douta(w_n699_11[0]),.doutb(w_n699_11[1]),.doutc(w_n699_11[2]),.din(w_n699_3[1]));
	jspl3 jspl3_w_n699_12(.douta(w_n699_12[0]),.doutb(w_n699_12[1]),.doutc(w_n699_12[2]),.din(w_n699_3[2]));
	jspl3 jspl3_w_n699_13(.douta(w_n699_13[0]),.doutb(w_n699_13[1]),.doutc(w_n699_13[2]),.din(w_n699_4[0]));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_n700_0[1]),.din(n700));
	jspl jspl_w_n702_0(.douta(w_n702_0[0]),.doutb(w_n702_0[1]),.din(n702));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl3 jspl3_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.doutc(w_n708_0[2]),.din(n708));
	jspl3 jspl3_w_n708_1(.douta(w_n708_1[0]),.doutb(w_n708_1[1]),.doutc(w_n708_1[2]),.din(w_n708_0[0]));
	jspl3 jspl3_w_n708_2(.douta(w_n708_2[0]),.doutb(w_n708_2[1]),.doutc(w_n708_2[2]),.din(w_n708_0[1]));
	jspl3 jspl3_w_n708_3(.douta(w_n708_3[0]),.doutb(w_n708_3[1]),.doutc(w_n708_3[2]),.din(w_n708_0[2]));
	jspl3 jspl3_w_n708_4(.douta(w_n708_4[0]),.doutb(w_n708_4[1]),.doutc(w_n708_4[2]),.din(w_n708_1[0]));
	jspl3 jspl3_w_n708_5(.douta(w_n708_5[0]),.doutb(w_n708_5[1]),.doutc(w_n708_5[2]),.din(w_n708_1[1]));
	jspl jspl_w_n708_6(.douta(w_n708_6[0]),.doutb(w_n708_6[1]),.din(w_n708_1[2]));
	jspl3 jspl3_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.doutc(w_n709_0[2]),.din(n709));
	jspl jspl_w_n709_1(.douta(w_n709_1[0]),.doutb(w_n709_1[1]),.din(w_n709_0[0]));
	jspl3 jspl3_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.doutc(w_n710_0[2]),.din(n710));
	jspl3 jspl3_w_n710_1(.douta(w_n710_1[0]),.doutb(w_n710_1[1]),.doutc(w_n710_1[2]),.din(w_n710_0[0]));
	jspl3 jspl3_w_n710_2(.douta(w_n710_2[0]),.doutb(w_n710_2[1]),.doutc(w_n710_2[2]),.din(w_n710_0[1]));
	jspl jspl_w_n710_3(.douta(w_n710_3[0]),.doutb(w_n710_3[1]),.din(w_n710_0[2]));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl3 jspl3_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.doutc(w_n712_0[2]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl3 jspl3_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.doutc(w_n719_0[2]),.din(n719));
	jspl jspl_w_n719_1(.douta(w_n719_1[0]),.doutb(w_n719_1[1]),.din(w_n719_0[0]));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl3 jspl3_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.doutc(w_n724_0[2]),.din(n724));
	jspl3 jspl3_w_n724_1(.douta(w_n724_1[0]),.doutb(w_n724_1[1]),.doutc(w_n724_1[2]),.din(w_n724_0[0]));
	jspl3 jspl3_w_n724_2(.douta(w_n724_2[0]),.doutb(w_n724_2[1]),.doutc(w_n724_2[2]),.din(w_n724_0[1]));
	jspl jspl_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.din(n725));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n730_0(.douta(w_n730_0[0]),.doutb(w_n730_0[1]),.doutc(w_n730_0[2]),.din(n730));
	jspl jspl_w_n730_1(.douta(w_n730_1[0]),.doutb(w_n730_1[1]),.din(w_n730_0[0]));
	jspl3 jspl3_w_n731_0(.douta(w_n731_0[0]),.doutb(w_n731_0[1]),.doutc(w_n731_0[2]),.din(n731));
	jspl3 jspl3_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.doutc(w_n732_0[2]),.din(n732));
	jspl3 jspl3_w_n732_1(.douta(w_n732_1[0]),.doutb(w_n732_1[1]),.doutc(w_n732_1[2]),.din(w_n732_0[0]));
	jspl3 jspl3_w_n732_2(.douta(w_n732_2[0]),.doutb(w_n732_2[1]),.doutc(w_n732_2[2]),.din(w_n732_0[1]));
	jspl jspl_w_n732_3(.douta(w_n732_3[0]),.doutb(w_n732_3[1]),.din(w_n732_0[2]));
	jspl3 jspl3_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.doutc(w_n733_0[2]),.din(n733));
	jspl jspl_w_n733_1(.douta(w_n733_1[0]),.doutb(w_n733_1[1]),.din(w_n733_0[0]));
	jspl3 jspl3_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.doutc(w_n734_0[2]),.din(n734));
	jspl3 jspl3_w_n734_1(.douta(w_n734_1[0]),.doutb(w_n734_1[1]),.doutc(w_n734_1[2]),.din(w_n734_0[0]));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.din(n735));
	jspl3 jspl3_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.doutc(w_n739_0[2]),.din(n739));
	jspl jspl_w_n740_0(.douta(w_n740_0[0]),.doutb(w_n740_0[1]),.din(n740));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n741_1(.douta(w_n741_1[0]),.doutb(w_n741_1[1]),.din(w_n741_0[0]));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_n744_0[2]),.din(n744));
	jspl3 jspl3_w_n744_1(.douta(w_n744_1[0]),.doutb(w_n744_1[1]),.doutc(w_n744_1[2]),.din(w_n744_0[0]));
	jspl3 jspl3_w_n744_2(.douta(w_n744_2[0]),.doutb(w_n744_2[1]),.doutc(w_n744_2[2]),.din(w_n744_0[1]));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.doutc(w_n746_0[2]),.din(n746));
	jspl3 jspl3_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.doutc(w_n748_0[2]),.din(n748));
	jspl jspl_w_n748_1(.douta(w_n748_1[0]),.doutb(w_n748_1[1]),.din(w_n748_0[0]));
	jspl3 jspl3_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.doutc(w_n749_0[2]),.din(n749));
	jspl jspl_w_n749_1(.douta(w_n749_1[0]),.doutb(w_n749_1[1]),.din(w_n749_0[0]));
	jspl jspl_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.din(n750));
	jspl3 jspl3_w_n751_0(.douta(w_n751_0[0]),.doutb(w_n751_0[1]),.doutc(w_n751_0[2]),.din(n751));
	jspl3 jspl3_w_n751_1(.douta(w_n751_1[0]),.doutb(w_n751_1[1]),.doutc(w_n751_1[2]),.din(w_n751_0[0]));
	jspl jspl_w_n751_2(.douta(w_n751_2[0]),.doutb(w_n751_2[1]),.din(w_n751_0[1]));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl jspl_w_n756_0(.douta(w_n756_0[0]),.doutb(w_n756_0[1]),.din(n756));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n758_0(.douta(w_n758_0[0]),.doutb(w_n758_0[1]),.din(n758));
	jspl3 jspl3_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.doutc(w_n762_0[2]),.din(n762));
	jspl3 jspl3_w_n762_1(.douta(w_n762_1[0]),.doutb(w_n762_1[1]),.doutc(w_n762_1[2]),.din(w_n762_0[0]));
	jspl jspl_w_n762_2(.douta(w_n762_2[0]),.doutb(w_n762_2[1]),.din(w_n762_0[1]));
	jspl3 jspl3_w_n763_0(.douta(w_n763_0[0]),.doutb(w_n763_0[1]),.doutc(w_n763_0[2]),.din(n763));
	jspl3 jspl3_w_n763_1(.douta(w_n763_1[0]),.doutb(w_n763_1[1]),.doutc(w_n763_1[2]),.din(w_n763_0[0]));
	jspl jspl_w_n763_2(.douta(w_n763_2[0]),.doutb(w_n763_2[1]),.din(w_n763_0[1]));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_n764_0[2]),.din(n764));
	jspl3 jspl3_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.doutc(w_n765_0[2]),.din(n765));
	jspl3 jspl3_w_n765_1(.douta(w_n765_1[0]),.doutb(w_n765_1[1]),.doutc(w_n765_1[2]),.din(w_n765_0[0]));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl3 jspl3_w_n768_0(.douta(w_n768_0[0]),.doutb(w_n768_0[1]),.doutc(w_n768_0[2]),.din(n768));
	jspl3 jspl3_w_n768_1(.douta(w_n768_1[0]),.doutb(w_n768_1[1]),.doutc(w_n768_1[2]),.din(w_n768_0[0]));
	jspl3 jspl3_w_n768_2(.douta(w_n768_2[0]),.doutb(w_n768_2[1]),.doutc(w_n768_2[2]),.din(w_n768_0[1]));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_n771_0[2]),.din(n771));
	jspl3 jspl3_w_n771_1(.douta(w_n771_1[0]),.doutb(w_n771_1[1]),.doutc(w_n771_1[2]),.din(w_n771_0[0]));
	jspl jspl_w_n771_2(.douta(w_n771_2[0]),.doutb(w_n771_2[1]),.din(w_n771_0[1]));
	jspl3 jspl3_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.doutc(w_n772_0[2]),.din(n772));
	jspl3 jspl3_w_n772_1(.douta(w_n772_1[0]),.doutb(w_n772_1[1]),.doutc(w_n772_1[2]),.din(w_n772_0[0]));
	jspl3 jspl3_w_n772_2(.douta(w_n772_2[0]),.doutb(w_n772_2[1]),.doutc(w_n772_2[2]),.din(w_n772_0[1]));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n776_0(.douta(w_n776_0[0]),.doutb(w_n776_0[1]),.din(n776));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.din(n779));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl3 jspl3_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.doutc(w_n781_0[2]),.din(n781));
	jspl3 jspl3_w_n781_1(.douta(w_n781_1[0]),.doutb(w_n781_1[1]),.doutc(w_n781_1[2]),.din(w_n781_0[0]));
	jspl jspl_w_n781_2(.douta(w_n781_2[0]),.doutb(w_n781_2[1]),.din(w_n781_0[1]));
	jspl jspl_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.din(n784));
	jspl3 jspl3_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.doutc(w_n786_0[2]),.din(n786));
	jspl jspl_w_n786_1(.douta(w_n786_1[0]),.doutb(w_n786_1[1]),.din(w_n786_0[0]));
	jspl3 jspl3_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.doutc(w_n788_0[2]),.din(n788));
	jspl3 jspl3_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.doutc(w_n789_0[2]),.din(n789));
	jspl3 jspl3_w_n789_1(.douta(w_n789_1[0]),.doutb(w_n789_1[1]),.doutc(w_n789_1[2]),.din(w_n789_0[0]));
	jspl3 jspl3_w_n789_2(.douta(w_n789_2[0]),.doutb(w_n789_2[1]),.doutc(w_n789_2[2]),.din(w_n789_0[1]));
	jspl3 jspl3_w_n789_3(.douta(w_n789_3[0]),.doutb(w_n789_3[1]),.doutc(w_n789_3[2]),.din(w_n789_0[2]));
	jspl3 jspl3_w_n789_4(.douta(w_n789_4[0]),.doutb(w_n789_4[1]),.doutc(w_n789_4[2]),.din(w_n789_1[0]));
	jspl jspl_w_n789_5(.douta(w_n789_5[0]),.doutb(w_n789_5[1]),.din(w_n789_1[1]));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.doutc(w_n790_0[2]),.din(n790));
	jspl3 jspl3_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.doutc(w_n792_0[2]),.din(n792));
	jspl3 jspl3_w_n794_0(.douta(w_n794_0[0]),.doutb(w_n794_0[1]),.doutc(w_n794_0[2]),.din(n794));
	jspl3 jspl3_w_n794_1(.douta(w_n794_1[0]),.doutb(w_n794_1[1]),.doutc(w_n794_1[2]),.din(w_n794_0[0]));
	jspl3 jspl3_w_n794_2(.douta(w_n794_2[0]),.doutb(w_n794_2[1]),.doutc(w_n794_2[2]),.din(w_n794_0[1]));
	jspl3 jspl3_w_n794_3(.douta(w_n794_3[0]),.doutb(w_n794_3[1]),.doutc(w_n794_3[2]),.din(w_n794_0[2]));
	jspl3 jspl3_w_n794_4(.douta(w_n794_4[0]),.doutb(w_n794_4[1]),.doutc(w_n794_4[2]),.din(w_n794_1[0]));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl3 jspl3_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.doutc(w_n799_0[2]),.din(n799));
	jspl3 jspl3_w_n799_1(.douta(w_n799_1[0]),.doutb(w_n799_1[1]),.doutc(w_n799_1[2]),.din(w_n799_0[0]));
	jspl3 jspl3_w_n799_2(.douta(w_n799_2[0]),.doutb(w_n799_2[1]),.doutc(w_n799_2[2]),.din(w_n799_0[1]));
	jspl3 jspl3_w_n799_3(.douta(w_n799_3[0]),.doutb(w_n799_3[1]),.doutc(w_n799_3[2]),.din(w_n799_0[2]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.doutc(w_n800_0[2]),.din(n800));
	jspl3 jspl3_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.doutc(w_n803_0[2]),.din(n803));
	jspl3 jspl3_w_n803_1(.douta(w_n803_1[0]),.doutb(w_n803_1[1]),.doutc(w_n803_1[2]),.din(w_n803_0[0]));
	jspl3 jspl3_w_n803_2(.douta(w_n803_2[0]),.doutb(w_n803_2[1]),.doutc(w_n803_2[2]),.din(w_n803_0[1]));
	jspl3 jspl3_w_n803_3(.douta(w_n803_3[0]),.doutb(w_n803_3[1]),.doutc(w_n803_3[2]),.din(w_n803_0[2]));
	jspl3 jspl3_w_n803_4(.douta(w_n803_4[0]),.doutb(w_n803_4[1]),.doutc(w_n803_4[2]),.din(w_n803_1[0]));
	jspl3 jspl3_w_n803_5(.douta(w_n803_5[0]),.doutb(w_n803_5[1]),.doutc(w_n803_5[2]),.din(w_n803_1[1]));
	jspl3 jspl3_w_n803_6(.douta(w_n803_6[0]),.doutb(w_n803_6[1]),.doutc(w_n803_6[2]),.din(w_n803_1[2]));
	jspl3 jspl3_w_n803_7(.douta(w_n803_7[0]),.doutb(w_n803_7[1]),.doutc(w_n803_7[2]),.din(w_n803_2[0]));
	jspl3 jspl3_w_n803_8(.douta(w_n803_8[0]),.doutb(w_n803_8[1]),.doutc(w_n803_8[2]),.din(w_n803_2[1]));
	jspl3 jspl3_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.doutc(w_n804_0[2]),.din(n804));
	jspl3 jspl3_w_n804_1(.douta(w_n804_1[0]),.doutb(w_n804_1[1]),.doutc(w_n804_1[2]),.din(w_n804_0[0]));
	jspl3 jspl3_w_n804_2(.douta(w_n804_2[0]),.doutb(w_n804_2[1]),.doutc(w_n804_2[2]),.din(w_n804_0[1]));
	jspl3 jspl3_w_n804_3(.douta(w_n804_3[0]),.doutb(w_n804_3[1]),.doutc(w_n804_3[2]),.din(w_n804_0[2]));
	jspl3 jspl3_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.doutc(w_n808_0[2]),.din(n808));
	jspl3 jspl3_w_n808_1(.douta(w_n808_1[0]),.doutb(w_n808_1[1]),.doutc(w_n808_1[2]),.din(w_n808_0[0]));
	jspl3 jspl3_w_n808_2(.douta(w_n808_2[0]),.doutb(w_n808_2[1]),.doutc(w_n808_2[2]),.din(w_n808_0[1]));
	jspl3 jspl3_w_n808_3(.douta(w_n808_3[0]),.doutb(w_n808_3[1]),.doutc(w_n808_3[2]),.din(w_n808_0[2]));
	jspl3 jspl3_w_n808_4(.douta(w_n808_4[0]),.doutb(w_n808_4[1]),.doutc(w_n808_4[2]),.din(w_n808_1[0]));
	jspl3 jspl3_w_n808_5(.douta(w_n808_5[0]),.doutb(w_n808_5[1]),.doutc(w_n808_5[2]),.din(w_n808_1[1]));
	jspl3 jspl3_w_n808_6(.douta(w_n808_6[0]),.doutb(w_n808_6[1]),.doutc(w_n808_6[2]),.din(w_n808_1[2]));
	jspl3 jspl3_w_n808_7(.douta(w_n808_7[0]),.doutb(w_n808_7[1]),.doutc(w_n808_7[2]),.din(w_n808_2[0]));
	jspl3 jspl3_w_n808_8(.douta(w_n808_8[0]),.doutb(w_n808_8[1]),.doutc(w_n808_8[2]),.din(w_n808_2[1]));
	jspl3 jspl3_w_n808_9(.douta(w_n808_9[0]),.doutb(w_n808_9[1]),.doutc(w_n808_9[2]),.din(w_n808_2[2]));
	jspl3 jspl3_w_n808_10(.douta(w_n808_10[0]),.doutb(w_n808_10[1]),.doutc(w_n808_10[2]),.din(w_n808_3[0]));
	jspl3 jspl3_w_n808_11(.douta(w_n808_11[0]),.doutb(w_n808_11[1]),.doutc(w_n808_11[2]),.din(w_n808_3[1]));
	jspl3 jspl3_w_n808_12(.douta(w_n808_12[0]),.doutb(w_n808_12[1]),.doutc(w_n808_12[2]),.din(w_n808_3[2]));
	jspl3 jspl3_w_n808_13(.douta(w_n808_13[0]),.doutb(w_n808_13[1]),.doutc(w_n808_13[2]),.din(w_n808_4[0]));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl3 jspl3_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.doutc(w_n820_0[2]),.din(n820));
	jspl3 jspl3_w_n820_1(.douta(w_n820_1[0]),.doutb(w_n820_1[1]),.doutc(w_n820_1[2]),.din(w_n820_0[0]));
	jspl3 jspl3_w_n820_2(.douta(w_n820_2[0]),.doutb(w_n820_2[1]),.doutc(w_n820_2[2]),.din(w_n820_0[1]));
	jspl3 jspl3_w_n820_3(.douta(w_n820_3[0]),.doutb(w_n820_3[1]),.doutc(w_n820_3[2]),.din(w_n820_0[2]));
	jspl3 jspl3_w_n820_4(.douta(w_n820_4[0]),.doutb(w_n820_4[1]),.doutc(w_n820_4[2]),.din(w_n820_1[0]));
	jspl3 jspl3_w_n820_5(.douta(w_n820_5[0]),.doutb(w_n820_5[1]),.doutc(w_n820_5[2]),.din(w_n820_1[1]));
	jspl3 jspl3_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.doutc(w_n821_0[2]),.din(n821));
	jspl jspl_w_n821_1(.douta(w_n821_1[0]),.doutb(w_n821_1[1]),.din(w_n821_0[0]));
	jspl3 jspl3_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.doutc(w_n822_0[2]),.din(n822));
	jspl3 jspl3_w_n822_1(.douta(w_n822_1[0]),.doutb(w_n822_1[1]),.doutc(w_n822_1[2]),.din(w_n822_0[0]));
	jspl jspl_w_n822_2(.douta(w_n822_2[0]),.doutb(w_n822_2[1]),.din(w_n822_0[1]));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl3 jspl3_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.doutc(w_n825_0[2]),.din(n825));
	jspl3 jspl3_w_n825_1(.douta(w_n825_1[0]),.doutb(w_n825_1[1]),.doutc(w_n825_1[2]),.din(w_n825_0[0]));
	jspl3 jspl3_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.doutc(w_n832_0[2]),.din(n832));
	jspl jspl_w_n832_1(.douta(w_n832_1[0]),.doutb(w_n832_1[1]),.din(w_n832_0[0]));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n836_0(.douta(w_n836_0[0]),.doutb(w_n836_0[1]),.din(n836));
	jspl3 jspl3_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.doutc(w_n837_0[2]),.din(n837));
	jspl3 jspl3_w_n837_1(.douta(w_n837_1[0]),.doutb(w_n837_1[1]),.doutc(w_n837_1[2]),.din(w_n837_0[0]));
	jspl jspl_w_n837_2(.douta(w_n837_2[0]),.doutb(w_n837_2[1]),.din(w_n837_0[1]));
	jspl jspl_w_n843_0(.douta(w_n843_0[0]),.doutb(w_n843_0[1]),.din(n843));
	jspl jspl_w_n846_0(.douta(w_n846_0[0]),.doutb(w_n846_0[1]),.din(n846));
	jspl3 jspl3_w_n849_0(.douta(w_n849_0[0]),.doutb(w_n849_0[1]),.doutc(w_n849_0[2]),.din(n849));
	jspl3 jspl3_w_n849_1(.douta(w_n849_1[0]),.doutb(w_n849_1[1]),.doutc(w_n849_1[2]),.din(w_n849_0[0]));
	jspl jspl_w_n849_2(.douta(w_n849_2[0]),.doutb(w_n849_2[1]),.din(w_n849_0[1]));
	jspl jspl_w_n850_0(.douta(w_n850_0[0]),.doutb(w_n850_0[1]),.din(n850));
	jspl jspl_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.din(n852));
	jspl3 jspl3_w_n853_0(.douta(w_n853_0[0]),.doutb(w_n853_0[1]),.doutc(w_n853_0[2]),.din(n853));
	jspl3 jspl3_w_n853_1(.douta(w_n853_1[0]),.doutb(w_n853_1[1]),.doutc(w_n853_1[2]),.din(w_n853_0[0]));
	jspl3 jspl3_w_n853_2(.douta(w_n853_2[0]),.doutb(w_n853_2[1]),.doutc(w_n853_2[2]),.din(w_n853_0[1]));
	jspl3 jspl3_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.doutc(w_n854_0[2]),.din(n854));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl jspl_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.din(n858));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.din(n863));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.din(n865));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(n866));
	jspl3 jspl3_w_n868_0(.douta(w_n868_0[0]),.doutb(w_n868_0[1]),.doutc(w_n868_0[2]),.din(n868));
	jspl jspl_w_n868_1(.douta(w_n868_1[0]),.doutb(w_n868_1[1]),.din(w_n868_0[0]));
	jspl3 jspl3_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.doutc(w_n869_0[2]),.din(n869));
	jspl jspl_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.din(n876));
	jspl jspl_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.din(n877));
	jspl3 jspl3_w_n878_0(.douta(w_n878_0[0]),.doutb(w_n878_0[1]),.doutc(w_n878_0[2]),.din(n878));
	jspl jspl_w_n878_1(.douta(w_n878_1[0]),.doutb(w_n878_1[1]),.din(w_n878_0[0]));
	jspl jspl_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.din(n880));
	jspl3 jspl3_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.doutc(w_n881_0[2]),.din(n881));
	jspl jspl_w_n881_1(.douta(w_n881_1[0]),.doutb(w_n881_1[1]),.din(w_n881_0[0]));
	jspl3 jspl3_w_n882_0(.douta(w_n882_0[0]),.doutb(w_n882_0[1]),.doutc(w_n882_0[2]),.din(n882));
	jspl3 jspl3_w_n882_1(.douta(w_n882_1[0]),.doutb(w_n882_1[1]),.doutc(w_n882_1[2]),.din(w_n882_0[0]));
	jspl jspl_w_n882_2(.douta(w_n882_2[0]),.doutb(w_n882_2[1]),.din(w_n882_0[1]));
	jspl jspl_w_n883_0(.douta(w_n883_0[0]),.doutb(w_n883_0[1]),.din(n883));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl3 jspl3_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.doutc(w_n890_0[2]),.din(n890));
	jspl3 jspl3_w_n890_1(.douta(w_n890_1[0]),.doutb(w_n890_1[1]),.doutc(w_n890_1[2]),.din(w_n890_0[0]));
	jspl jspl_w_n893_0(.douta(w_n893_0[0]),.doutb(w_n893_0[1]),.din(n893));
	jspl jspl_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl3 jspl3_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.doutc(w_n897_0[2]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(n898));
	jspl jspl_w_n902_0(.douta(w_n902_0[0]),.doutb(w_n902_0[1]),.din(n902));
	jspl jspl_w_n904_0(.douta(w_n904_0[0]),.doutb(w_n904_0[1]),.din(n904));
	jspl jspl_w_n905_0(.douta(w_n905_0[0]),.doutb(w_n905_0[1]),.din(n905));
	jspl jspl_w_n906_0(.douta(w_n906_0[0]),.doutb(w_n906_0[1]),.din(n906));
	jspl jspl_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.din(n912));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n917_0(.douta(w_n917_0[0]),.doutb(w_n917_0[1]),.din(n917));
	jspl3 jspl3_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.doutc(w_n918_0[2]),.din(n918));
	jspl3 jspl3_w_n918_1(.douta(w_n918_1[0]),.doutb(w_n918_1[1]),.doutc(w_n918_1[2]),.din(w_n918_0[0]));
	jspl jspl_w_n918_2(.douta(w_n918_2[0]),.doutb(w_n918_2[1]),.din(w_n918_0[1]));
	jspl jspl_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.din(n920));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(n923));
	jspl3 jspl3_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.doutc(w_n924_0[2]),.din(n924));
	jspl3 jspl3_w_n924_1(.douta(w_n924_1[0]),.doutb(w_n924_1[1]),.doutc(w_n924_1[2]),.din(w_n924_0[0]));
	jspl3 jspl3_w_n925_0(.douta(w_n925_0[0]),.doutb(w_n925_0[1]),.doutc(w_n925_0[2]),.din(n925));
	jspl jspl_w_n925_1(.douta(w_n925_1[0]),.doutb(w_n925_1[1]),.din(w_n925_0[0]));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(n929));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_n930_0[2]),.din(n930));
	jspl jspl_w_n930_1(.douta(w_n930_1[0]),.doutb(w_n930_1[1]),.din(w_n930_0[0]));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n933_0(.douta(w_n933_0[0]),.doutb(w_n933_0[1]),.din(n933));
	jspl3 jspl3_w_n934_0(.douta(w_n934_0[0]),.doutb(w_n934_0[1]),.doutc(w_n934_0[2]),.din(n934));
	jspl3 jspl3_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.doutc(w_n935_0[2]),.din(n935));
	jspl3 jspl3_w_n935_1(.douta(w_n935_1[0]),.doutb(w_n935_1[1]),.doutc(w_n935_1[2]),.din(w_n935_0[0]));
	jspl3 jspl3_w_n935_2(.douta(w_n935_2[0]),.doutb(w_n935_2[1]),.doutc(w_n935_2[2]),.din(w_n935_0[1]));
	jspl jspl_w_n935_3(.douta(w_n935_3[0]),.doutb(w_n935_3[1]),.din(w_n935_0[2]));
	jspl3 jspl3_w_n936_0(.douta(w_n936_0[0]),.doutb(w_n936_0[1]),.doutc(w_n936_0[2]),.din(n936));
	jspl3 jspl3_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.doutc(w_n938_0[2]),.din(n938));
	jspl3 jspl3_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.doutc(w_n942_0[2]),.din(n942));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_n943_0[1]),.din(n943));
	jspl jspl_w_n950_0(.douta(w_n950_0[0]),.doutb(w_n950_0[1]),.din(n950));
	jspl3 jspl3_w_n951_0(.douta(w_n951_0[0]),.doutb(w_n951_0[1]),.doutc(w_n951_0[2]),.din(n951));
	jspl3 jspl3_w_n951_1(.douta(w_n951_1[0]),.doutb(w_n951_1[1]),.doutc(w_n951_1[2]),.din(w_n951_0[0]));
	jspl3 jspl3_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.doutc(w_n952_0[2]),.din(n952));
	jspl3 jspl3_w_n952_1(.douta(w_n952_1[0]),.doutb(w_n952_1[1]),.doutc(w_n952_1[2]),.din(w_n952_0[0]));
	jspl3 jspl3_w_n952_2(.douta(w_n952_2[0]),.doutb(w_n952_2[1]),.doutc(w_n952_2[2]),.din(w_n952_0[1]));
	jspl3 jspl3_w_n952_3(.douta(w_n952_3[0]),.doutb(w_n952_3[1]),.doutc(w_n952_3[2]),.din(w_n952_0[2]));
	jspl jspl_w_n952_4(.douta(w_n952_4[0]),.doutb(w_n952_4[1]),.din(w_n952_1[0]));
	jspl3 jspl3_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.doutc(w_n954_0[2]),.din(n954));
	jspl3 jspl3_w_n954_1(.douta(w_n954_1[0]),.doutb(w_n954_1[1]),.doutc(w_n954_1[2]),.din(w_n954_0[0]));
	jspl3 jspl3_w_n954_2(.douta(w_n954_2[0]),.doutb(w_n954_2[1]),.doutc(w_n954_2[2]),.din(w_n954_0[1]));
	jspl3 jspl3_w_n954_3(.douta(w_n954_3[0]),.doutb(w_n954_3[1]),.doutc(w_n954_3[2]),.din(w_n954_0[2]));
	jspl3 jspl3_w_n954_4(.douta(w_n954_4[0]),.doutb(w_n954_4[1]),.doutc(w_n954_4[2]),.din(w_n954_1[0]));
	jspl3 jspl3_w_n954_5(.douta(w_n954_5[0]),.doutb(w_n954_5[1]),.doutc(w_n954_5[2]),.din(w_n954_1[1]));
	jspl3 jspl3_w_n954_6(.douta(w_n954_6[0]),.doutb(w_n954_6[1]),.doutc(w_n954_6[2]),.din(w_n954_1[2]));
	jspl3 jspl3_w_n954_7(.douta(w_n954_7[0]),.doutb(w_n954_7[1]),.doutc(w_n954_7[2]),.din(w_n954_2[0]));
	jspl3 jspl3_w_n954_8(.douta(w_n954_8[0]),.doutb(w_n954_8[1]),.doutc(w_n954_8[2]),.din(w_n954_2[1]));
	jspl3 jspl3_w_n954_9(.douta(w_n954_9[0]),.doutb(w_n954_9[1]),.doutc(w_n954_9[2]),.din(w_n954_2[2]));
	jspl3 jspl3_w_n954_10(.douta(w_n954_10[0]),.doutb(w_n954_10[1]),.doutc(w_n954_10[2]),.din(w_n954_3[0]));
	jspl3 jspl3_w_n954_11(.douta(w_n954_11[0]),.doutb(w_n954_11[1]),.doutc(w_n954_11[2]),.din(w_n954_3[1]));
	jspl3 jspl3_w_n954_12(.douta(w_n954_12[0]),.doutb(w_n954_12[1]),.doutc(w_n954_12[2]),.din(w_n954_3[2]));
	jspl3 jspl3_w_n954_13(.douta(w_n954_13[0]),.doutb(w_n954_13[1]),.doutc(w_n954_13[2]),.din(w_n954_4[0]));
	jspl3 jspl3_w_n954_14(.douta(w_n954_14[0]),.doutb(w_n954_14[1]),.doutc(w_n954_14[2]),.din(w_n954_4[1]));
	jspl3 jspl3_w_n954_15(.douta(w_n954_15[0]),.doutb(w_n954_15[1]),.doutc(w_n954_15[2]),.din(w_n954_4[2]));
	jspl3 jspl3_w_n954_16(.douta(w_n954_16[0]),.doutb(w_n954_16[1]),.doutc(w_n954_16[2]),.din(w_n954_5[0]));
	jspl3 jspl3_w_n954_17(.douta(w_n954_17[0]),.doutb(w_n954_17[1]),.doutc(w_n954_17[2]),.din(w_n954_5[1]));
	jspl3 jspl3_w_n954_18(.douta(w_n954_18[0]),.doutb(w_n954_18[1]),.doutc(w_n954_18[2]),.din(w_n954_5[2]));
	jspl3 jspl3_w_n954_19(.douta(w_n954_19[0]),.doutb(w_n954_19[1]),.doutc(w_n954_19[2]),.din(w_n954_6[0]));
	jspl3 jspl3_w_n954_20(.douta(w_n954_20[0]),.doutb(w_n954_20[1]),.doutc(w_n954_20[2]),.din(w_n954_6[1]));
	jspl3 jspl3_w_n954_21(.douta(w_n954_21[0]),.doutb(w_n954_21[1]),.doutc(w_n954_21[2]),.din(w_n954_6[2]));
	jspl3 jspl3_w_n954_22(.douta(w_n954_22[0]),.doutb(w_n954_22[1]),.doutc(w_n954_22[2]),.din(w_n954_7[0]));
	jspl3 jspl3_w_n954_23(.douta(w_n954_23[0]),.doutb(w_n954_23[1]),.doutc(w_n954_23[2]),.din(w_n954_7[1]));
	jspl jspl_w_n954_24(.douta(w_n954_24[0]),.doutb(w_n954_24[1]),.din(w_n954_7[2]));
	jspl3 jspl3_w_n955_0(.douta(w_n955_0[0]),.doutb(w_n955_0[1]),.doutc(w_n955_0[2]),.din(n955));
	jspl3 jspl3_w_n956_0(.douta(w_n956_0[0]),.doutb(w_n956_0[1]),.doutc(w_n956_0[2]),.din(n956));
	jspl3 jspl3_w_n956_1(.douta(w_n956_1[0]),.doutb(w_n956_1[1]),.doutc(w_n956_1[2]),.din(w_n956_0[0]));
	jspl3 jspl3_w_n956_2(.douta(w_n956_2[0]),.doutb(w_n956_2[1]),.doutc(w_n956_2[2]),.din(w_n956_0[1]));
	jspl3 jspl3_w_n956_3(.douta(w_n956_3[0]),.doutb(w_n956_3[1]),.doutc(w_n956_3[2]),.din(w_n956_0[2]));
	jspl jspl_w_n956_4(.douta(w_n956_4[0]),.doutb(w_n956_4[1]),.din(w_n956_1[0]));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(n959));
	jspl3 jspl3_w_n960_0(.douta(w_n960_0[0]),.doutb(w_n960_0[1]),.doutc(w_n960_0[2]),.din(n960));
	jspl3 jspl3_w_n960_1(.douta(w_n960_1[0]),.doutb(w_n960_1[1]),.doutc(w_n960_1[2]),.din(w_n960_0[0]));
	jspl3 jspl3_w_n960_2(.douta(w_n960_2[0]),.doutb(w_n960_2[1]),.doutc(w_n960_2[2]),.din(w_n960_0[1]));
	jspl3 jspl3_w_n960_3(.douta(w_n960_3[0]),.doutb(w_n960_3[1]),.doutc(w_n960_3[2]),.din(w_n960_0[2]));
	jspl3 jspl3_w_n960_4(.douta(w_n960_4[0]),.doutb(w_n960_4[1]),.doutc(w_n960_4[2]),.din(w_n960_1[0]));
	jspl3 jspl3_w_n960_5(.douta(w_n960_5[0]),.doutb(w_n960_5[1]),.doutc(w_n960_5[2]),.din(w_n960_1[1]));
	jspl3 jspl3_w_n961_0(.douta(w_n961_0[0]),.doutb(w_n961_0[1]),.doutc(w_n961_0[2]),.din(n961));
	jspl3 jspl3_w_n961_1(.douta(w_n961_1[0]),.doutb(w_n961_1[1]),.doutc(w_n961_1[2]),.din(w_n961_0[0]));
	jspl3 jspl3_w_n961_2(.douta(w_n961_2[0]),.doutb(w_n961_2[1]),.doutc(w_n961_2[2]),.din(w_n961_0[1]));
	jspl3 jspl3_w_n961_3(.douta(w_n961_3[0]),.doutb(w_n961_3[1]),.doutc(w_n961_3[2]),.din(w_n961_0[2]));
	jspl3 jspl3_w_n961_4(.douta(w_n961_4[0]),.doutb(w_n961_4[1]),.doutc(w_n961_4[2]),.din(w_n961_1[0]));
	jspl jspl_w_n961_5(.douta(w_n961_5[0]),.doutb(w_n961_5[1]),.din(w_n961_1[1]));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl3 jspl3_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.doutc(w_n964_0[2]),.din(n964));
	jspl jspl_w_n964_1(.douta(w_n964_1[0]),.doutb(w_n964_1[1]),.din(w_n964_0[0]));
	jspl jspl_w_n965_0(.douta(w_n965_0[0]),.doutb(w_n965_0[1]),.din(n965));
	jspl3 jspl3_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.doutc(w_n966_0[2]),.din(n966));
	jspl3 jspl3_w_n966_1(.douta(w_n966_1[0]),.doutb(w_n966_1[1]),.doutc(w_n966_1[2]),.din(w_n966_0[0]));
	jspl3 jspl3_w_n966_2(.douta(w_n966_2[0]),.doutb(w_n966_2[1]),.doutc(w_n966_2[2]),.din(w_n966_0[1]));
	jspl3 jspl3_w_n966_3(.douta(w_n966_3[0]),.doutb(w_n966_3[1]),.doutc(w_n966_3[2]),.din(w_n966_0[2]));
	jspl jspl_w_n966_4(.douta(w_n966_4[0]),.doutb(w_n966_4[1]),.din(w_n966_1[0]));
	jspl jspl_w_n968_0(.douta(w_n968_0[0]),.doutb(w_n968_0[1]),.din(n968));
	jspl3 jspl3_w_n970_0(.douta(w_n970_0[0]),.doutb(w_n970_0[1]),.doutc(w_n970_0[2]),.din(n970));
	jspl3 jspl3_w_n971_0(.douta(w_n971_0[0]),.doutb(w_n971_0[1]),.doutc(w_n971_0[2]),.din(n971));
	jspl3 jspl3_w_n971_1(.douta(w_n971_1[0]),.doutb(w_n971_1[1]),.doutc(w_n971_1[2]),.din(w_n971_0[0]));
	jspl3 jspl3_w_n971_2(.douta(w_n971_2[0]),.doutb(w_n971_2[1]),.doutc(w_n971_2[2]),.din(w_n971_0[1]));
	jspl3 jspl3_w_n971_3(.douta(w_n971_3[0]),.doutb(w_n971_3[1]),.doutc(w_n971_3[2]),.din(w_n971_0[2]));
	jspl jspl_w_n971_4(.douta(w_n971_4[0]),.doutb(w_n971_4[1]),.din(w_n971_1[0]));
	jspl jspl_w_n975_0(.douta(w_n975_0[0]),.doutb(w_n975_0[1]),.din(n975));
	jspl3 jspl3_w_n980_0(.douta(w_n980_0[0]),.doutb(w_n980_0[1]),.doutc(w_n980_0[2]),.din(n980));
	jspl3 jspl3_w_n980_1(.douta(w_n980_1[0]),.doutb(w_n980_1[1]),.doutc(w_n980_1[2]),.din(w_n980_0[0]));
	jspl3 jspl3_w_n980_2(.douta(w_n980_2[0]),.doutb(w_n980_2[1]),.doutc(w_n980_2[2]),.din(w_n980_0[1]));
	jspl3 jspl3_w_n980_3(.douta(w_n980_3[0]),.doutb(w_n980_3[1]),.doutc(w_n980_3[2]),.din(w_n980_0[2]));
	jspl3 jspl3_w_n980_4(.douta(w_n980_4[0]),.doutb(w_n980_4[1]),.doutc(w_n980_4[2]),.din(w_n980_1[0]));
	jspl3 jspl3_w_n980_5(.douta(w_n980_5[0]),.doutb(w_n980_5[1]),.doutc(w_n980_5[2]),.din(w_n980_1[1]));
	jspl jspl_w_n980_6(.douta(w_n980_6[0]),.doutb(w_n980_6[1]),.din(w_n980_1[2]));
	jspl3 jspl3_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.doutc(w_n981_0[2]),.din(n981));
	jspl3 jspl3_w_n981_1(.douta(w_n981_1[0]),.doutb(w_n981_1[1]),.doutc(w_n981_1[2]),.din(w_n981_0[0]));
	jspl3 jspl3_w_n981_2(.douta(w_n981_2[0]),.doutb(w_n981_2[1]),.doutc(w_n981_2[2]),.din(w_n981_0[1]));
	jspl3 jspl3_w_n981_3(.douta(w_n981_3[0]),.doutb(w_n981_3[1]),.doutc(w_n981_3[2]),.din(w_n981_0[2]));
	jspl3 jspl3_w_n981_4(.douta(w_n981_4[0]),.doutb(w_n981_4[1]),.doutc(w_n981_4[2]),.din(w_n981_1[0]));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl3 jspl3_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.doutc(w_n987_0[2]),.din(n987));
	jspl3 jspl3_w_n987_1(.douta(w_n987_1[0]),.doutb(w_n987_1[1]),.doutc(w_n987_1[2]),.din(w_n987_0[0]));
	jspl jspl_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.din(n988));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(n991));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl3 jspl3_w_n992_1(.douta(w_n992_1[0]),.doutb(w_n992_1[1]),.doutc(w_n992_1[2]),.din(w_n992_0[0]));
	jspl3 jspl3_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.doutc(w_n993_0[2]),.din(n993));
	jspl3 jspl3_w_n993_1(.douta(w_n993_1[0]),.doutb(w_n993_1[1]),.doutc(w_n993_1[2]),.din(w_n993_0[0]));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.doutc(w_n999_0[2]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.din(n1002));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.din(n1006));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl3 jspl3_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.doutc(w_n1018_0[2]),.din(n1018));
	jspl jspl_w_n1018_1(.douta(w_n1018_1[0]),.doutb(w_n1018_1[1]),.din(w_n1018_0[0]));
	jspl jspl_w_n1020_0(.douta(w_n1020_0[0]),.doutb(w_n1020_0[1]),.din(n1020));
	jspl jspl_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.din(n1021));
	jspl3 jspl3_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.doutc(w_n1022_0[2]),.din(n1022));
	jspl3 jspl3_w_n1025_0(.douta(w_n1025_0[0]),.doutb(w_n1025_0[1]),.doutc(w_n1025_0[2]),.din(n1025));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl3 jspl3_w_n1027_0(.douta(w_n1027_0[0]),.doutb(w_n1027_0[1]),.doutc(w_n1027_0[2]),.din(n1027));
	jspl jspl_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.din(n1032));
	jspl3 jspl3_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.doutc(w_n1033_0[2]),.din(n1033));
	jspl3 jspl3_w_n1033_1(.douta(w_n1033_1[0]),.doutb(w_n1033_1[1]),.doutc(w_n1033_1[2]),.din(w_n1033_0[0]));
	jspl3 jspl3_w_n1034_0(.douta(w_n1034_0[0]),.doutb(w_n1034_0[1]),.doutc(w_n1034_0[2]),.din(n1034));
	jspl3 jspl3_w_n1034_1(.douta(w_n1034_1[0]),.doutb(w_n1034_1[1]),.doutc(w_n1034_1[2]),.din(w_n1034_0[0]));
	jspl3 jspl3_w_n1034_2(.douta(w_n1034_2[0]),.doutb(w_n1034_2[1]),.doutc(w_n1034_2[2]),.din(w_n1034_0[1]));
	jspl3 jspl3_w_n1034_3(.douta(w_n1034_3[0]),.doutb(w_n1034_3[1]),.doutc(w_n1034_3[2]),.din(w_n1034_0[2]));
	jspl3 jspl3_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.doutc(w_n1035_0[2]),.din(n1035));
	jspl3 jspl3_w_n1037_0(.douta(w_n1037_0[0]),.doutb(w_n1037_0[1]),.doutc(w_n1037_0[2]),.din(n1037));
	jspl3 jspl3_w_n1037_1(.douta(w_n1037_1[0]),.doutb(w_n1037_1[1]),.doutc(w_n1037_1[2]),.din(w_n1037_0[0]));
	jspl3 jspl3_w_n1037_2(.douta(w_n1037_2[0]),.doutb(w_n1037_2[1]),.doutc(w_n1037_2[2]),.din(w_n1037_0[1]));
	jspl3 jspl3_w_n1037_3(.douta(w_n1037_3[0]),.doutb(w_n1037_3[1]),.doutc(w_n1037_3[2]),.din(w_n1037_0[2]));
	jspl3 jspl3_w_n1038_0(.douta(w_n1038_0[0]),.doutb(w_n1038_0[1]),.doutc(w_n1038_0[2]),.din(n1038));
	jspl3 jspl3_w_n1042_0(.douta(w_n1042_0[0]),.doutb(w_n1042_0[1]),.doutc(w_n1042_0[2]),.din(n1042));
	jspl3 jspl3_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.doutc(w_n1043_0[2]),.din(n1043));
	jspl3 jspl3_w_n1043_1(.douta(w_n1043_1[0]),.doutb(w_n1043_1[1]),.doutc(w_n1043_1[2]),.din(w_n1043_0[0]));
	jspl3 jspl3_w_n1043_2(.douta(w_n1043_2[0]),.doutb(w_n1043_2[1]),.doutc(w_n1043_2[2]),.din(w_n1043_0[1]));
	jspl3 jspl3_w_n1043_3(.douta(w_n1043_3[0]),.doutb(w_n1043_3[1]),.doutc(w_n1043_3[2]),.din(w_n1043_0[2]));
	jspl jspl_w_n1043_4(.douta(w_n1043_4[0]),.doutb(w_n1043_4[1]),.din(w_n1043_1[0]));
	jspl jspl_w_n1045_0(.douta(w_n1045_0[0]),.doutb(w_n1045_0[1]),.din(n1045));
	jspl3 jspl3_w_n1047_0(.douta(w_n1047_0[0]),.doutb(w_n1047_0[1]),.doutc(w_n1047_0[2]),.din(n1047));
	jspl jspl_w_n1047_1(.douta(w_n1047_1[0]),.doutb(w_n1047_1[1]),.din(w_n1047_0[0]));
	jspl3 jspl3_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.doutc(w_n1049_0[2]),.din(n1049));
	jspl3 jspl3_w_n1049_1(.douta(w_n1049_1[0]),.doutb(w_n1049_1[1]),.doutc(w_n1049_1[2]),.din(w_n1049_0[0]));
	jspl3 jspl3_w_n1049_2(.douta(w_n1049_2[0]),.doutb(w_n1049_2[1]),.doutc(w_n1049_2[2]),.din(w_n1049_0[1]));
	jspl3 jspl3_w_n1049_3(.douta(w_n1049_3[0]),.doutb(w_n1049_3[1]),.doutc(w_n1049_3[2]),.din(w_n1049_0[2]));
	jspl jspl_w_n1049_4(.douta(w_n1049_4[0]),.doutb(w_n1049_4[1]),.din(w_n1049_1[0]));
	jspl jspl_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.din(n1053));
	jspl jspl_w_n1055_0(.douta(w_n1055_0[0]),.doutb(w_n1055_0[1]),.din(n1055));
	jspl3 jspl3_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.doutc(w_n1057_0[2]),.din(n1057));
	jspl3 jspl3_w_n1057_1(.douta(w_n1057_1[0]),.doutb(w_n1057_1[1]),.doutc(w_n1057_1[2]),.din(w_n1057_0[0]));
	jspl3 jspl3_w_n1057_2(.douta(w_n1057_2[0]),.doutb(w_n1057_2[1]),.doutc(w_n1057_2[2]),.din(w_n1057_0[1]));
	jspl3 jspl3_w_n1057_3(.douta(w_n1057_3[0]),.doutb(w_n1057_3[1]),.doutc(w_n1057_3[2]),.din(w_n1057_0[2]));
	jspl3 jspl3_w_n1057_4(.douta(w_n1057_4[0]),.doutb(w_n1057_4[1]),.doutc(w_n1057_4[2]),.din(w_n1057_1[0]));
	jspl jspl_w_n1057_5(.douta(w_n1057_5[0]),.doutb(w_n1057_5[1]),.din(w_n1057_1[1]));
	jspl3 jspl3_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.doutc(w_n1059_0[2]),.din(n1059));
	jspl3 jspl3_w_n1059_1(.douta(w_n1059_1[0]),.doutb(w_n1059_1[1]),.doutc(w_n1059_1[2]),.din(w_n1059_0[0]));
	jspl3 jspl3_w_n1059_2(.douta(w_n1059_2[0]),.doutb(w_n1059_2[1]),.doutc(w_n1059_2[2]),.din(w_n1059_0[1]));
	jspl3 jspl3_w_n1059_3(.douta(w_n1059_3[0]),.doutb(w_n1059_3[1]),.doutc(w_n1059_3[2]),.din(w_n1059_0[2]));
	jspl3 jspl3_w_n1059_4(.douta(w_n1059_4[0]),.doutb(w_n1059_4[1]),.doutc(w_n1059_4[2]),.din(w_n1059_1[0]));
	jspl3 jspl3_w_n1059_5(.douta(w_n1059_5[0]),.doutb(w_n1059_5[1]),.doutc(w_n1059_5[2]),.din(w_n1059_1[1]));
	jspl jspl_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.din(n1066));
	jspl jspl_w_n1068_0(.douta(w_n1068_0[0]),.doutb(w_n1068_0[1]),.din(n1068));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(n1069));
	jspl jspl_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.din(n1071));
	jspl jspl_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.din(n1072));
	jspl3 jspl3_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.doutc(w_n1073_0[2]),.din(n1073));
	jspl jspl_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.din(n1074));
	jspl jspl_w_n1075_0(.douta(w_n1075_0[0]),.doutb(w_n1075_0[1]),.din(n1075));
	jspl jspl_w_n1076_0(.douta(w_n1076_0[0]),.doutb(w_n1076_0[1]),.din(n1076));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(n1078));
	jspl jspl_w_n1083_0(.douta(w_n1083_0[0]),.doutb(w_n1083_0[1]),.din(n1083));
	jspl jspl_w_n1085_0(.douta(w_n1085_0[0]),.doutb(w_n1085_0[1]),.din(n1085));
	jspl jspl_w_n1093_0(.douta(w_n1093_0[0]),.doutb(w_n1093_0[1]),.din(n1093));
	jspl jspl_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.din(n1095));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1110_0(.douta(w_n1110_0[0]),.doutb(w_n1110_0[1]),.din(n1110));
	jspl jspl_w_n1111_0(.douta(w_n1111_0[0]),.doutb(w_n1111_0[1]),.din(n1111));
	jspl jspl_w_n1113_0(.douta(w_n1113_0[0]),.doutb(w_n1113_0[1]),.din(n1113));
	jspl jspl_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.din(n1114));
	jspl3 jspl3_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.doutc(w_n1115_0[2]),.din(n1115));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl jspl_w_n1121_0(.douta(w_n1121_0[0]),.doutb(w_n1121_0[1]),.din(n1121));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.din(n1133));
	jspl jspl_w_n1138_0(.douta(w_n1138_0[0]),.doutb(w_n1138_0[1]),.din(n1138));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1140_0(.douta(w_n1140_0[0]),.doutb(w_n1140_0[1]),.din(n1140));
	jspl3 jspl3_w_n1143_0(.douta(w_n1143_0[0]),.doutb(w_n1143_0[1]),.doutc(w_n1143_0[2]),.din(n1143));
	jspl3 jspl3_w_n1143_1(.douta(w_n1143_1[0]),.doutb(w_n1143_1[1]),.doutc(w_n1143_1[2]),.din(w_n1143_0[0]));
	jspl3 jspl3_w_n1143_2(.douta(w_n1143_2[0]),.doutb(w_n1143_2[1]),.doutc(w_n1143_2[2]),.din(w_n1143_0[1]));
	jspl3 jspl3_w_n1143_3(.douta(w_n1143_3[0]),.doutb(w_n1143_3[1]),.doutc(w_n1143_3[2]),.din(w_n1143_0[2]));
	jspl3 jspl3_w_n1143_4(.douta(w_n1143_4[0]),.doutb(w_n1143_4[1]),.doutc(w_n1143_4[2]),.din(w_n1143_1[0]));
	jspl3 jspl3_w_n1143_5(.douta(w_n1143_5[0]),.doutb(w_n1143_5[1]),.doutc(w_n1143_5[2]),.din(w_n1143_1[1]));
	jspl3 jspl3_w_n1143_6(.douta(w_n1143_6[0]),.doutb(w_n1143_6[1]),.doutc(w_n1143_6[2]),.din(w_n1143_1[2]));
	jspl3 jspl3_w_n1143_7(.douta(w_n1143_7[0]),.doutb(w_n1143_7[1]),.doutc(w_n1143_7[2]),.din(w_n1143_2[0]));
	jspl3 jspl3_w_n1143_8(.douta(w_n1143_8[0]),.doutb(w_n1143_8[1]),.doutc(w_n1143_8[2]),.din(w_n1143_2[1]));
	jspl jspl_w_n1143_9(.douta(w_n1143_9[0]),.doutb(w_n1143_9[1]),.din(w_n1143_2[2]));
	jspl jspl_w_n1150_0(.douta(w_n1150_0[0]),.doutb(w_n1150_0[1]),.din(n1150));
	jspl jspl_w_n1152_0(.douta(w_n1152_0[0]),.doutb(w_n1152_0[1]),.din(n1152));
	jspl jspl_w_n1159_0(.douta(w_n1159_0[0]),.doutb(w_n1159_0[1]),.din(n1159));
	jspl jspl_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.din(n1163));
	jspl jspl_w_n1169_0(.douta(w_n1169_0[0]),.doutb(w_n1169_0[1]),.din(n1169));
	jspl3 jspl3_w_n1170_0(.douta(w_n1170_0[0]),.doutb(w_n1170_0[1]),.doutc(w_n1170_0[2]),.din(n1170));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_n1175_0[1]),.din(n1175));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(n1176));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl3 jspl3_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.doutc(w_n1185_0[2]),.din(n1185));
	jspl3 jspl3_w_n1185_1(.douta(w_n1185_1[0]),.doutb(w_n1185_1[1]),.doutc(w_n1185_1[2]),.din(w_n1185_0[0]));
	jspl3 jspl3_w_n1187_0(.douta(w_n1187_0[0]),.doutb(w_n1187_0[1]),.doutc(w_n1187_0[2]),.din(n1187));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(n1188));
	jspl3 jspl3_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.doutc(w_n1189_0[2]),.din(n1189));
	jspl jspl_w_n1189_1(.douta(w_n1189_1[0]),.doutb(w_n1189_1[1]),.din(w_n1189_0[0]));
	jspl jspl_w_n1190_0(.douta(w_n1190_0[0]),.doutb(w_n1190_0[1]),.din(n1190));
	jspl jspl_w_n1192_0(.douta(w_n1192_0[0]),.doutb(w_n1192_0[1]),.din(n1192));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(n1193));
	jspl3 jspl3_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.doutc(w_n1196_0[2]),.din(n1196));
	jspl jspl_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.din(n1197));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(n1198));
	jspl3 jspl3_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.doutc(w_n1203_0[2]),.din(n1203));
	jspl3 jspl3_w_n1204_0(.douta(w_n1204_0[0]),.doutb(w_n1204_0[1]),.doutc(w_n1204_0[2]),.din(n1204));
	jspl jspl_w_n1204_1(.douta(w_n1204_1[0]),.doutb(w_n1204_1[1]),.din(w_n1204_0[0]));
	jspl3 jspl3_w_n1209_0(.douta(w_n1209_0[0]),.doutb(w_n1209_0[1]),.doutc(w_n1209_0[2]),.din(n1209));
	jspl3 jspl3_w_n1209_1(.douta(w_n1209_1[0]),.doutb(w_n1209_1[1]),.doutc(w_n1209_1[2]),.din(w_n1209_0[0]));
	jspl jspl_w_n1210_0(.douta(w_n1210_0[0]),.doutb(w_n1210_0[1]),.din(n1210));
	jspl jspl_w_n1214_0(.douta(w_n1214_0[0]),.doutb(w_n1214_0[1]),.din(n1214));
	jspl jspl_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.din(n1215));
	jspl3 jspl3_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.doutc(w_n1217_0[2]),.din(n1217));
	jspl3 jspl3_w_n1218_0(.douta(w_n1218_0[0]),.doutb(w_n1218_0[1]),.doutc(w_n1218_0[2]),.din(n1218));
	jspl jspl_w_n1224_0(.douta(w_n1224_0[0]),.doutb(w_n1224_0[1]),.din(n1224));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(n1227));
	jspl jspl_w_n1228_0(.douta(w_n1228_0[0]),.doutb(w_n1228_0[1]),.din(n1228));
	jspl3 jspl3_w_n1231_0(.douta(w_n1231_0[0]),.doutb(w_n1231_0[1]),.doutc(w_n1231_0[2]),.din(n1231));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(n1232));
	jspl jspl_w_n1239_0(.douta(w_n1239_0[0]),.doutb(w_n1239_0[1]),.din(n1239));
	jspl jspl_w_n1240_0(.douta(w_n1240_0[0]),.doutb(w_n1240_0[1]),.din(n1240));
	jspl3 jspl3_w_n1243_0(.douta(w_n1243_0[0]),.doutb(w_n1243_0[1]),.doutc(w_n1243_0[2]),.din(n1243));
	jspl3 jspl3_w_n1243_1(.douta(w_n1243_1[0]),.doutb(w_n1243_1[1]),.doutc(w_n1243_1[2]),.din(w_n1243_0[0]));
	jspl jspl_w_n1243_2(.douta(w_n1243_2[0]),.doutb(w_n1243_2[1]),.din(w_n1243_0[1]));
	jspl jspl_w_n1245_0(.douta(w_n1245_0[0]),.doutb(w_n1245_0[1]),.din(n1245));
	jspl jspl_w_n1259_0(.douta(w_n1259_0[0]),.doutb(w_n1259_0[1]),.din(n1259));
	jspl3 jspl3_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.doutc(w_n1283_0[2]),.din(n1283));
	jspl3 jspl3_w_n1283_1(.douta(w_n1283_1[0]),.doutb(w_n1283_1[1]),.doutc(w_n1283_1[2]),.din(w_n1283_0[0]));
	jspl3 jspl3_w_n1283_2(.douta(w_n1283_2[0]),.doutb(w_n1283_2[1]),.doutc(w_n1283_2[2]),.din(w_n1283_0[1]));
	jspl3 jspl3_w_n1283_3(.douta(w_n1283_3[0]),.doutb(w_n1283_3[1]),.doutc(w_n1283_3[2]),.din(w_n1283_0[2]));
	jspl3 jspl3_w_n1283_4(.douta(w_n1283_4[0]),.doutb(w_n1283_4[1]),.doutc(w_n1283_4[2]),.din(w_n1283_1[0]));
	jspl3 jspl3_w_n1283_5(.douta(w_n1283_5[0]),.doutb(w_n1283_5[1]),.doutc(w_n1283_5[2]),.din(w_n1283_1[1]));
	jspl3 jspl3_w_n1283_6(.douta(w_n1283_6[0]),.doutb(w_n1283_6[1]),.doutc(w_n1283_6[2]),.din(w_n1283_1[2]));
	jspl3 jspl3_w_n1283_7(.douta(w_n1283_7[0]),.doutb(w_n1283_7[1]),.doutc(w_n1283_7[2]),.din(w_n1283_2[0]));
	jspl3 jspl3_w_n1283_8(.douta(w_n1283_8[0]),.doutb(w_n1283_8[1]),.doutc(w_n1283_8[2]),.din(w_n1283_2[1]));
	jspl3 jspl3_w_n1283_9(.douta(w_n1283_9[0]),.doutb(w_n1283_9[1]),.doutc(w_n1283_9[2]),.din(w_n1283_2[2]));
	jspl3 jspl3_w_n1283_10(.douta(w_n1283_10[0]),.doutb(w_n1283_10[1]),.doutc(w_n1283_10[2]),.din(w_n1283_3[0]));
	jspl3 jspl3_w_n1283_11(.douta(w_n1283_11[0]),.doutb(w_n1283_11[1]),.doutc(w_n1283_11[2]),.din(w_n1283_3[1]));
	jspl3 jspl3_w_n1283_12(.douta(w_n1283_12[0]),.doutb(w_n1283_12[1]),.doutc(w_n1283_12[2]),.din(w_n1283_3[2]));
	jspl jspl_w_n1285_0(.douta(w_n1285_0[0]),.doutb(w_n1285_0[1]),.din(n1285));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(n1288));
	jspl jspl_w_n1292_0(.douta(w_n1292_0[0]),.doutb(w_n1292_0[1]),.din(n1292));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(n1293));
	jspl jspl_w_n1294_0(.douta(w_n1294_0[0]),.doutb(w_n1294_0[1]),.din(n1294));
	jspl jspl_w_n1299_0(.douta(w_n1299_0[0]),.doutb(w_n1299_0[1]),.din(n1299));
	jspl jspl_w_n1302_0(.douta(w_n1302_0[0]),.doutb(w_n1302_0[1]),.din(n1302));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(n1307));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(n1312));
	jspl jspl_w_n1319_0(.douta(w_n1319_0[0]),.doutb(w_n1319_0[1]),.din(n1319));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.din(n1322));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl3 jspl3_w_n1328_0(.douta(w_n1328_0[0]),.doutb(w_n1328_0[1]),.doutc(w_n1328_0[2]),.din(n1328));
	jspl jspl_w_n1329_0(.douta(w_n1329_0[0]),.doutb(w_n1329_0[1]),.din(n1329));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(n1332));
	jspl3 jspl3_w_n1338_0(.douta(w_n1338_0[0]),.doutb(w_n1338_0[1]),.doutc(w_n1338_0[2]),.din(n1338));
	jspl3 jspl3_w_n1339_0(.douta(w_n1339_0[0]),.doutb(w_n1339_0[1]),.doutc(w_n1339_0[2]),.din(n1339));
	jspl3 jspl3_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_n1340_0[1]),.doutc(w_n1340_0[2]),.din(n1340));
	jspl jspl_w_n1342_0(.douta(w_n1342_0[0]),.doutb(w_n1342_0[1]),.din(n1342));
	jspl3 jspl3_w_n1347_0(.douta(w_n1347_0[0]),.doutb(w_n1347_0[1]),.doutc(w_n1347_0[2]),.din(n1347));
	jspl3 jspl3_w_n1347_1(.douta(w_n1347_1[0]),.doutb(w_n1347_1[1]),.doutc(w_n1347_1[2]),.din(w_n1347_0[0]));
	jspl3 jspl3_w_n1347_2(.douta(w_n1347_2[0]),.doutb(w_n1347_2[1]),.doutc(w_n1347_2[2]),.din(w_n1347_0[1]));
	jspl3 jspl3_w_n1347_3(.douta(w_n1347_3[0]),.doutb(w_n1347_3[1]),.doutc(w_n1347_3[2]),.din(w_n1347_0[2]));
	jspl3 jspl3_w_n1347_4(.douta(w_n1347_4[0]),.doutb(w_n1347_4[1]),.doutc(w_n1347_4[2]),.din(w_n1347_1[0]));
	jspl3 jspl3_w_n1347_5(.douta(w_n1347_5[0]),.doutb(w_n1347_5[1]),.doutc(w_n1347_5[2]),.din(w_n1347_1[1]));
	jspl jspl_w_n1347_6(.douta(w_n1347_6[0]),.doutb(w_n1347_6[1]),.din(w_n1347_1[2]));
	jspl jspl_w_n1348_0(.douta(w_n1348_0[0]),.doutb(w_n1348_0[1]),.din(n1348));
	jspl jspl_w_n1350_0(.douta(w_n1350_0[0]),.doutb(w_n1350_0[1]),.din(n1350));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(n1351));
	jspl jspl_w_n1354_0(.douta(w_n1354_0[0]),.doutb(w_n1354_0[1]),.din(n1354));
	jspl3 jspl3_w_n1356_0(.douta(w_n1356_0[0]),.doutb(w_n1356_0[1]),.doutc(w_n1356_0[2]),.din(n1356));
	jspl jspl_w_n1356_1(.douta(w_n1356_1[0]),.doutb(w_n1356_1[1]),.din(w_n1356_0[0]));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl3 jspl3_w_n1362_0(.douta(w_n1362_0[0]),.doutb(w_n1362_0[1]),.doutc(w_n1362_0[2]),.din(n1362));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_n1364_0[1]),.din(n1364));
	jspl jspl_w_n1367_0(.douta(w_n1367_0[0]),.doutb(w_n1367_0[1]),.din(n1367));
	jspl jspl_w_n1375_0(.douta(w_n1375_0[0]),.doutb(w_n1375_0[1]),.din(n1375));
	jspl jspl_w_n1377_0(.douta(w_n1377_0[0]),.doutb(w_n1377_0[1]),.din(n1377));
	jspl jspl_w_n1379_0(.douta(w_n1379_0[0]),.doutb(w_n1379_0[1]),.din(n1379));
	jspl jspl_w_n1380_0(.douta(w_n1380_0[0]),.doutb(w_n1380_0[1]),.din(n1380));
	jspl jspl_w_n1382_0(.douta(w_n1382_0[0]),.doutb(w_n1382_0[1]),.din(n1382));
	jspl jspl_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.din(n1383));
	jspl jspl_w_n1385_0(.douta(w_n1385_0[0]),.doutb(w_n1385_0[1]),.din(n1385));
	jspl jspl_w_n1386_0(.douta(w_n1386_0[0]),.doutb(w_n1386_0[1]),.din(n1386));
	jspl jspl_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_n1388_0[1]),.din(n1388));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(n1389));
	jspl3 jspl3_w_n1391_0(.douta(w_n1391_0[0]),.doutb(w_n1391_0[1]),.doutc(w_n1391_0[2]),.din(n1391));
	jspl3 jspl3_w_n1391_1(.douta(w_n1391_1[0]),.doutb(w_n1391_1[1]),.doutc(w_n1391_1[2]),.din(w_n1391_0[0]));
	jspl3 jspl3_w_n1391_2(.douta(w_n1391_2[0]),.doutb(w_n1391_2[1]),.doutc(w_n1391_2[2]),.din(w_n1391_0[1]));
	jspl3 jspl3_w_n1391_3(.douta(w_n1391_3[0]),.doutb(w_n1391_3[1]),.doutc(w_n1391_3[2]),.din(w_n1391_0[2]));
	jspl3 jspl3_w_n1391_4(.douta(w_n1391_4[0]),.doutb(w_n1391_4[1]),.doutc(w_n1391_4[2]),.din(w_n1391_1[0]));
	jspl3 jspl3_w_n1391_5(.douta(w_n1391_5[0]),.doutb(w_n1391_5[1]),.doutc(w_n1391_5[2]),.din(w_n1391_1[1]));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(n1399));
	jspl jspl_w_n1407_0(.douta(w_n1407_0[0]),.doutb(w_n1407_0[1]),.din(n1407));
	jspl jspl_w_n1409_0(.douta(w_n1409_0[0]),.doutb(w_n1409_0[1]),.din(n1409));
	jspl3 jspl3_w_n1411_0(.douta(w_n1411_0[0]),.doutb(w_n1411_0[1]),.doutc(w_n1411_0[2]),.din(n1411));
	jspl3 jspl3_w_n1411_1(.douta(w_n1411_1[0]),.doutb(w_n1411_1[1]),.doutc(w_n1411_1[2]),.din(w_n1411_0[0]));
	jspl3 jspl3_w_n1411_2(.douta(w_n1411_2[0]),.doutb(w_n1411_2[1]),.doutc(w_n1411_2[2]),.din(w_n1411_0[1]));
	jspl jspl_w_n1413_0(.douta(w_n1413_0[0]),.doutb(w_n1413_0[1]),.din(n1413));
	jspl3 jspl3_w_n1414_0(.douta(w_n1414_0[0]),.doutb(w_n1414_0[1]),.doutc(w_n1414_0[2]),.din(n1414));
	jspl3 jspl3_w_n1414_1(.douta(w_n1414_1[0]),.doutb(w_n1414_1[1]),.doutc(w_n1414_1[2]),.din(w_n1414_0[0]));
	jspl3 jspl3_w_n1414_2(.douta(w_n1414_2[0]),.doutb(w_n1414_2[1]),.doutc(w_n1414_2[2]),.din(w_n1414_0[1]));
	jspl jspl_w_n1417_0(.douta(w_n1417_0[0]),.doutb(w_n1417_0[1]),.din(n1417));
	jspl3 jspl3_w_n1418_0(.douta(w_n1418_0[0]),.doutb(w_n1418_0[1]),.doutc(w_n1418_0[2]),.din(n1418));
	jspl3 jspl3_w_n1418_1(.douta(w_n1418_1[0]),.doutb(w_n1418_1[1]),.doutc(w_n1418_1[2]),.din(w_n1418_0[0]));
	jspl3 jspl3_w_n1418_2(.douta(w_n1418_2[0]),.doutb(w_n1418_2[1]),.doutc(w_n1418_2[2]),.din(w_n1418_0[1]));
	jspl3 jspl3_w_n1418_3(.douta(w_n1418_3[0]),.doutb(w_n1418_3[1]),.doutc(w_n1418_3[2]),.din(w_n1418_0[2]));
	jspl jspl_w_n1418_4(.douta(w_n1418_4[0]),.doutb(w_n1418_4[1]),.din(w_n1418_1[0]));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(n1420));
	jspl3 jspl3_w_n1421_0(.douta(w_n1421_0[0]),.doutb(w_n1421_0[1]),.doutc(w_n1421_0[2]),.din(n1421));
	jspl3 jspl3_w_n1421_1(.douta(w_n1421_1[0]),.doutb(w_n1421_1[1]),.doutc(w_n1421_1[2]),.din(w_n1421_0[0]));
	jspl3 jspl3_w_n1421_2(.douta(w_n1421_2[0]),.doutb(w_n1421_2[1]),.doutc(w_n1421_2[2]),.din(w_n1421_0[1]));
	jspl3 jspl3_w_n1421_3(.douta(w_n1421_3[0]),.doutb(w_n1421_3[1]),.doutc(w_n1421_3[2]),.din(w_n1421_0[2]));
	jspl jspl_w_n1421_4(.douta(w_n1421_4[0]),.doutb(w_n1421_4[1]),.din(w_n1421_1[0]));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1427_0(.douta(w_n1427_0[0]),.doutb(w_n1427_0[1]),.din(n1427));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(n1428));
	jspl jspl_w_n1430_0(.douta(w_n1430_0[0]),.doutb(w_n1430_0[1]),.din(n1430));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(n1431));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(n1436));
	jspl jspl_w_n1437_0(.douta(w_n1437_0[0]),.doutb(w_n1437_0[1]),.din(n1437));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.din(n1440));
	jspl jspl_w_n1442_0(.douta(w_n1442_0[0]),.doutb(w_n1442_0[1]),.din(n1442));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(n1454));
	jspl jspl_w_n1456_0(.douta(w_n1456_0[0]),.doutb(w_n1456_0[1]),.din(n1456));
	jspl jspl_w_n1458_0(.douta(w_n1458_0[0]),.doutb(w_n1458_0[1]),.din(n1458));
	jspl jspl_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.din(n1513));
	jspl jspl_w_n1514_0(.douta(w_n1514_0[0]),.doutb(w_n1514_0[1]),.din(n1514));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(n1515));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(n1517));
	jspl3 jspl3_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.doutc(w_n1520_0[2]),.din(n1520));
	jspl jspl_w_n1521_0(.douta(w_n1521_0[0]),.doutb(w_n1521_0[1]),.din(n1521));
	jspl jspl_w_n1524_0(.douta(w_n1524_0[0]),.doutb(w_n1524_0[1]),.din(n1524));
	jspl jspl_w_n1526_0(.douta(w_n1526_0[0]),.doutb(w_n1526_0[1]),.din(n1526));
	jspl jspl_w_n1527_0(.douta(w_n1527_0[0]),.doutb(w_n1527_0[1]),.din(n1527));
	jspl jspl_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.din(n1529));
	jspl3 jspl3_w_n1533_0(.douta(w_n1533_0[0]),.doutb(w_n1533_0[1]),.doutc(w_n1533_0[2]),.din(n1533));
	jspl3 jspl3_w_n1533_1(.douta(w_n1533_1[0]),.doutb(w_n1533_1[1]),.doutc(w_n1533_1[2]),.din(w_n1533_0[0]));
	jspl3 jspl3_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.doutc(w_n1535_0[2]),.din(n1535));
	jspl3 jspl3_w_n1535_1(.douta(w_n1535_1[0]),.doutb(w_n1535_1[1]),.doutc(w_n1535_1[2]),.din(w_n1535_0[0]));
	jspl jspl_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.din(n1539));
	jspl jspl_w_n1541_0(.douta(w_n1541_0[0]),.doutb(w_n1541_0[1]),.din(n1541));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(n1548));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_n1550_0[1]),.din(n1550));
	jspl jspl_w_n1558_0(.douta(w_n1558_0[0]),.doutb(w_n1558_0[1]),.din(n1558));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1561_0(.douta(w_n1561_0[0]),.doutb(w_n1561_0[1]),.din(n1561));
	jspl jspl_w_n1563_0(.douta(w_n1563_0[0]),.doutb(w_n1563_0[1]),.din(n1563));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(n1565));
	jspl3 jspl3_w_n1566_0(.douta(w_n1566_0[0]),.doutb(w_n1566_0[1]),.doutc(w_n1566_0[2]),.din(n1566));
	jspl3 jspl3_w_n1566_1(.douta(w_n1566_1[0]),.doutb(w_n1566_1[1]),.doutc(w_n1566_1[2]),.din(w_n1566_0[0]));
	jspl3 jspl3_w_n1566_2(.douta(w_n1566_2[0]),.doutb(w_n1566_2[1]),.doutc(w_n1566_2[2]),.din(w_n1566_0[1]));
	jspl jspl_w_n1566_3(.douta(w_n1566_3[0]),.doutb(w_n1566_3[1]),.din(w_n1566_0[2]));
	jspl3 jspl3_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_n1568_0[1]),.doutc(w_n1568_0[2]),.din(n1568));
	jspl3 jspl3_w_n1568_1(.douta(w_n1568_1[0]),.doutb(w_n1568_1[1]),.doutc(w_n1568_1[2]),.din(w_n1568_0[0]));
	jspl3 jspl3_w_n1568_2(.douta(w_n1568_2[0]),.doutb(w_n1568_2[1]),.doutc(w_n1568_2[2]),.din(w_n1568_0[1]));
	jspl jspl_w_n1568_3(.douta(w_n1568_3[0]),.doutb(w_n1568_3[1]),.din(w_n1568_0[2]));
	jspl3 jspl3_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.doutc(w_n1571_0[2]),.din(n1571));
	jspl jspl_w_n1571_1(.douta(w_n1571_1[0]),.doutb(w_n1571_1[1]),.din(w_n1571_0[0]));
	jspl3 jspl3_w_n1572_0(.douta(w_n1572_0[0]),.doutb(w_n1572_0[1]),.doutc(w_n1572_0[2]),.din(n1572));
	jspl3 jspl3_w_n1572_1(.douta(w_n1572_1[0]),.doutb(w_n1572_1[1]),.doutc(w_n1572_1[2]),.din(w_n1572_0[0]));
	jspl3 jspl3_w_n1572_2(.douta(w_n1572_2[0]),.doutb(w_n1572_2[1]),.doutc(w_n1572_2[2]),.din(w_n1572_0[1]));
	jspl jspl_w_n1572_3(.douta(w_n1572_3[0]),.doutb(w_n1572_3[1]),.din(w_n1572_0[2]));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(n1574));
	jspl jspl_w_n1575_0(.douta(w_n1575_0[0]),.doutb(w_n1575_0[1]),.din(n1575));
	jspl3 jspl3_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.doutc(w_n1576_0[2]),.din(n1576));
	jspl3 jspl3_w_n1577_0(.douta(w_n1577_0[0]),.doutb(w_n1577_0[1]),.doutc(w_n1577_0[2]),.din(n1577));
	jspl3 jspl3_w_n1577_1(.douta(w_n1577_1[0]),.doutb(w_n1577_1[1]),.doutc(w_n1577_1[2]),.din(w_n1577_0[0]));
	jspl3 jspl3_w_n1577_2(.douta(w_n1577_2[0]),.doutb(w_n1577_2[1]),.doutc(w_n1577_2[2]),.din(w_n1577_0[1]));
	jspl jspl_w_n1577_3(.douta(w_n1577_3[0]),.doutb(w_n1577_3[1]),.din(w_n1577_0[2]));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_n1581_0[1]),.din(n1581));
	jspl jspl_w_n1583_0(.douta(w_n1583_0[0]),.doutb(w_n1583_0[1]),.din(n1583));
	jspl3 jspl3_w_n1584_0(.douta(w_n1584_0[0]),.doutb(w_n1584_0[1]),.doutc(w_n1584_0[2]),.din(n1584));
	jspl3 jspl3_w_n1584_1(.douta(w_n1584_1[0]),.doutb(w_n1584_1[1]),.doutc(w_n1584_1[2]),.din(w_n1584_0[0]));
	jspl3 jspl3_w_n1584_2(.douta(w_n1584_2[0]),.doutb(w_n1584_2[1]),.doutc(w_n1584_2[2]),.din(w_n1584_0[1]));
	jspl3 jspl3_w_n1584_3(.douta(w_n1584_3[0]),.doutb(w_n1584_3[1]),.doutc(w_n1584_3[2]),.din(w_n1584_0[2]));
	jspl3 jspl3_w_n1584_4(.douta(w_n1584_4[0]),.doutb(w_n1584_4[1]),.doutc(w_n1584_4[2]),.din(w_n1584_1[0]));
	jspl jspl_w_n1592_0(.douta(w_n1592_0[0]),.doutb(w_n1592_0[1]),.din(n1592));
	jspl jspl_w_n1594_0(.douta(w_n1594_0[0]),.doutb(w_n1594_0[1]),.din(n1594));
	jspl jspl_w_n1595_0(.douta(w_n1595_0[0]),.doutb(w_n1595_0[1]),.din(n1595));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(n1597));
	jspl jspl_w_n1604_0(.douta(w_n1604_0[0]),.doutb(w_n1604_0[1]),.din(n1604));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(n1612));
	jspl jspl_w_n1614_0(.douta(w_n1614_0[0]),.doutb(w_n1614_0[1]),.din(n1614));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(n1622));
	jspl jspl_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.din(n1624));
	jspl jspl_w_n1626_0(.douta(w_n1626_0[0]),.doutb(w_n1626_0[1]),.din(n1626));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(n1631));
	jspl jspl_w_n1632_0(.douta(w_n1632_0[0]),.doutb(w_n1632_0[1]),.din(n1632));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(n1634));
	jspl jspl_w_n1635_0(.douta(w_n1635_0[0]),.doutb(w_n1635_0[1]),.din(n1635));
	jspl jspl_w_n1637_0(.douta(w_n1637_0[0]),.doutb(w_n1637_0[1]),.din(n1637));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(n1638));
	jspl jspl_w_n1640_0(.douta(w_n1640_0[0]),.doutb(w_n1640_0[1]),.din(n1640));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_n1641_0[1]),.din(n1641));
	jspl3 jspl3_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.doutc(w_n1646_0[2]),.din(n1646));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(n1653));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(n1658));
	jspl jspl_w_n1669_0(.douta(w_n1669_0[0]),.doutb(w_n1669_0[1]),.din(n1669));
	jspl jspl_w_n1673_0(.douta(w_n1673_0[0]),.doutb(w_n1673_0[1]),.din(n1673));
	jspl jspl_w_n1675_0(.douta(w_n1675_0[0]),.doutb(w_n1675_0[1]),.din(n1675));
	jspl jspl_w_n1676_0(.douta(w_n1676_0[0]),.doutb(w_n1676_0[1]),.din(n1676));
	jspl jspl_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.din(n1679));
	jspl3 jspl3_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.doutc(w_n1682_0[2]),.din(n1682));
	jspl3 jspl3_w_n1682_1(.douta(w_n1682_1[0]),.doutb(w_n1682_1[1]),.doutc(w_n1682_1[2]),.din(w_n1682_0[0]));
	jspl3 jspl3_w_n1682_2(.douta(w_n1682_2[0]),.doutb(w_n1682_2[1]),.doutc(w_n1682_2[2]),.din(w_n1682_0[1]));
	jspl3 jspl3_w_n1682_3(.douta(w_n1682_3[0]),.doutb(w_n1682_3[1]),.doutc(w_n1682_3[2]),.din(w_n1682_0[2]));
	jspl3 jspl3_w_n1682_4(.douta(w_n1682_4[0]),.doutb(w_n1682_4[1]),.doutc(w_n1682_4[2]),.din(w_n1682_1[0]));
	jspl jspl_w_n1682_5(.douta(w_n1682_5[0]),.doutb(w_n1682_5[1]),.din(w_n1682_1[1]));
	jspl3 jspl3_w_n1683_0(.douta(w_n1683_0[0]),.doutb(w_n1683_0[1]),.doutc(w_n1683_0[2]),.din(n1683));
	jspl3 jspl3_w_n1683_1(.douta(w_n1683_1[0]),.doutb(w_n1683_1[1]),.doutc(w_n1683_1[2]),.din(w_n1683_0[0]));
	jspl3 jspl3_w_n1683_2(.douta(w_n1683_2[0]),.doutb(w_n1683_2[1]),.doutc(w_n1683_2[2]),.din(w_n1683_0[1]));
	jspl3 jspl3_w_n1683_3(.douta(w_n1683_3[0]),.doutb(w_n1683_3[1]),.doutc(w_n1683_3[2]),.din(w_n1683_0[2]));
	jspl3 jspl3_w_n1683_4(.douta(w_n1683_4[0]),.doutb(w_n1683_4[1]),.doutc(w_n1683_4[2]),.din(w_n1683_1[0]));
	jspl jspl_w_n1685_0(.douta(w_n1685_0[0]),.doutb(w_n1685_0[1]),.din(n1685));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_n1687_0[1]),.din(n1687));
	jspl3 jspl3_w_n1688_0(.douta(w_n1688_0[0]),.doutb(w_n1688_0[1]),.doutc(w_n1688_0[2]),.din(n1688));
	jspl jspl_w_n1688_1(.douta(w_n1688_1[0]),.doutb(w_n1688_1[1]),.din(w_n1688_0[0]));
	jspl3 jspl3_w_n1690_0(.douta(w_n1690_0[0]),.doutb(w_n1690_0[1]),.doutc(w_n1690_0[2]),.din(n1690));
	jspl jspl_w_n1690_1(.douta(w_n1690_1[0]),.doutb(w_n1690_1[1]),.din(w_n1690_0[0]));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_n1697_0[1]),.din(n1697));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(n1699));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(n1707));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(n1709));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1727_0(.douta(w_n1727_0[0]),.doutb(w_n1727_0[1]),.din(n1727));
	jspl jspl_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.din(n1735));
	jspl jspl_w_n1737_0(.douta(w_n1737_0[0]),.doutb(w_n1737_0[1]),.din(n1737));
	jspl jspl_w_n1739_0(.douta(w_n1739_0[0]),.doutb(w_n1739_0[1]),.din(n1739));
	jspl jspl_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.din(n1740));
	jspl jspl_w_n1742_0(.douta(w_n1742_0[0]),.doutb(w_n1742_0[1]),.din(n1742));
	jspl jspl_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.din(n1743));
	jspl jspl_w_n1745_0(.douta(w_n1745_0[0]),.doutb(w_n1745_0[1]),.din(n1745));
	jspl jspl_w_n1746_0(.douta(w_n1746_0[0]),.doutb(w_n1746_0[1]),.din(n1746));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(n1748));
	jspl jspl_w_n1749_0(.douta(w_n1749_0[0]),.doutb(w_n1749_0[1]),.din(n1749));
	jspl jspl_w_n1751_0(.douta(w_n1751_0[0]),.doutb(w_n1751_0[1]),.din(n1751));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1760_0(.douta(w_n1760_0[0]),.doutb(w_n1760_0[1]),.din(n1760));
	jspl jspl_w_n1761_0(.douta(w_n1761_0[0]),.doutb(w_n1761_0[1]),.din(n1761));
	jspl3 jspl3_w_n1762_0(.douta(w_n1762_0[0]),.doutb(w_n1762_0[1]),.doutc(w_n1762_0[2]),.din(n1762));
	jspl3 jspl3_w_n1762_1(.douta(w_n1762_1[0]),.doutb(w_n1762_1[1]),.doutc(w_n1762_1[2]),.din(w_n1762_0[0]));
	jspl3 jspl3_w_n1762_2(.douta(w_n1762_2[0]),.doutb(w_n1762_2[1]),.doutc(w_n1762_2[2]),.din(w_n1762_0[1]));
	jspl3 jspl3_w_n1762_3(.douta(w_n1762_3[0]),.doutb(w_n1762_3[1]),.doutc(w_n1762_3[2]),.din(w_n1762_0[2]));
	jspl3 jspl3_w_n1762_4(.douta(w_n1762_4[0]),.doutb(w_n1762_4[1]),.doutc(w_n1762_4[2]),.din(w_n1762_1[0]));
	jspl jspl_w_n1762_5(.douta(w_n1762_5[0]),.doutb(w_n1762_5[1]),.din(w_n1762_1[1]));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(n1770));
	jspl jspl_w_n1779_0(.douta(w_n1779_0[0]),.doutb(w_n1779_0[1]),.din(n1779));
	jspl jspl_w_n1787_0(.douta(w_n1787_0[0]),.doutb(w_n1787_0[1]),.din(n1787));
	jspl jspl_w_n1789_0(.douta(w_n1789_0[0]),.doutb(w_n1789_0[1]),.din(n1789));
	jspl jspl_w_n1797_0(.douta(w_n1797_0[0]),.doutb(w_n1797_0[1]),.din(n1797));
	jspl jspl_w_n1799_0(.douta(w_n1799_0[0]),.doutb(w_n1799_0[1]),.din(n1799));
	jspl jspl_w_n1800_0(.douta(w_n1800_0[0]),.doutb(w_n1800_0[1]),.din(n1800));
	jspl jspl_w_n1802_0(.douta(w_n1802_0[0]),.doutb(w_n1802_0[1]),.din(n1802));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(n1803));
	jspl jspl_w_n1805_0(.douta(w_n1805_0[0]),.doutb(w_n1805_0[1]),.din(n1805));
	jspl jspl_w_n1806_0(.douta(w_n1806_0[0]),.doutb(w_n1806_0[1]),.din(n1806));
	jspl jspl_w_n1808_0(.douta(w_n1808_0[0]),.doutb(w_n1808_0[1]),.din(n1808));
	jspl jspl_w_n1809_0(.douta(w_n1809_0[0]),.doutb(w_n1809_0[1]),.din(n1809));
	jspl jspl_w_n1811_0(.douta(w_n1811_0[0]),.doutb(w_n1811_0[1]),.din(n1811));
	jspl jspl_w_n1812_0(.douta(w_n1812_0[0]),.doutb(w_n1812_0[1]),.din(n1812));
	jspl jspl_w_n1814_0(.douta(w_n1814_0[0]),.doutb(w_n1814_0[1]),.din(n1814));
	jspl jspl_w_n1815_0(.douta(w_n1815_0[0]),.doutb(w_n1815_0[1]),.din(n1815));
	jspl jspl_w_n1824_0(.douta(w_n1824_0[0]),.doutb(w_n1824_0[1]),.din(n1824));
	jspl jspl_w_n1832_0(.douta(w_n1832_0[0]),.doutb(w_n1832_0[1]),.din(n1832));
	jspl jspl_w_n1834_0(.douta(w_n1834_0[0]),.doutb(w_n1834_0[1]),.din(n1834));
	jspl jspl_w_n1835_0(.douta(w_n1835_0[0]),.doutb(w_n1835_0[1]),.din(n1835));
	jspl jspl_w_n1837_0(.douta(w_n1837_0[0]),.doutb(w_n1837_0[1]),.din(n1837));
	jspl jspl_w_n1838_0(.douta(w_n1838_0[0]),.doutb(w_n1838_0[1]),.din(n1838));
	jspl jspl_w_n1840_0(.douta(w_n1840_0[0]),.doutb(w_n1840_0[1]),.din(n1840));
	jspl jspl_w_n1841_0(.douta(w_n1841_0[0]),.doutb(w_n1841_0[1]),.din(n1841));
	jspl jspl_w_n1843_0(.douta(w_n1843_0[0]),.doutb(w_n1843_0[1]),.din(n1843));
	jspl jspl_w_n1844_0(.douta(w_n1844_0[0]),.doutb(w_n1844_0[1]),.din(n1844));
	jspl jspl_w_n1846_0(.douta(w_n1846_0[0]),.doutb(w_n1846_0[1]),.din(n1846));
	jspl jspl_w_n1847_0(.douta(w_n1847_0[0]),.doutb(w_n1847_0[1]),.din(n1847));
	jspl jspl_w_n1849_0(.douta(w_n1849_0[0]),.doutb(w_n1849_0[1]),.din(n1849));
	jspl jspl_w_n1850_0(.douta(w_n1850_0[0]),.doutb(w_n1850_0[1]),.din(n1850));
	jspl jspl_w_n1858_0(.douta(w_n1858_0[0]),.doutb(w_n1858_0[1]),.din(n1858));
	jspl jspl_w_n1866_0(.douta(w_n1866_0[0]),.doutb(w_n1866_0[1]),.din(n1866));
	jspl3 jspl3_w_n1869_0(.douta(w_n1869_0[0]),.doutb(w_n1869_0[1]),.doutc(w_n1869_0[2]),.din(n1869));
	jspl jspl_w_n1871_0(.douta(w_n1871_0[0]),.doutb(w_n1871_0[1]),.din(n1871));
	jspl jspl_w_n1872_0(.douta(w_n1872_0[0]),.doutb(w_n1872_0[1]),.din(n1872));
	jspl jspl_w_n1878_0(.douta(w_n1878_0[0]),.doutb(w_n1878_0[1]),.din(n1878));
	jspl jspl_w_n1879_0(.douta(w_n1879_0[0]),.doutb(w_n1879_0[1]),.din(n1879));
	jspl jspl_w_n1880_0(.douta(w_n1880_0[0]),.doutb(w_n1880_0[1]),.din(n1880));
	jspl jspl_w_n1882_0(.douta(w_n1882_0[0]),.doutb(w_n1882_0[1]),.din(n1882));
	jspl jspl_w_n1883_0(.douta(w_n1883_0[0]),.doutb(w_n1883_0[1]),.din(n1883));
	jspl jspl_w_n1889_0(.douta(w_n1889_0[0]),.doutb(w_n1889_0[1]),.din(n1889));
	jspl jspl_w_n1897_0(.douta(w_n1897_0[0]),.doutb(w_n1897_0[1]),.din(n1897));
	jspl jspl_w_n1899_0(.douta(w_n1899_0[0]),.doutb(w_n1899_0[1]),.din(n1899));
	jspl jspl_w_n1907_0(.douta(w_n1907_0[0]),.doutb(w_n1907_0[1]),.din(n1907));
	jspl jspl_w_n1909_0(.douta(w_n1909_0[0]),.doutb(w_n1909_0[1]),.din(n1909));
	jspl jspl_w_n1911_0(.douta(w_n1911_0[0]),.doutb(w_n1911_0[1]),.din(n1911));
	jspl jspl_w_n1912_0(.douta(w_n1912_0[0]),.doutb(w_n1912_0[1]),.din(n1912));
	jspl jspl_w_n1914_0(.douta(w_n1914_0[0]),.doutb(w_n1914_0[1]),.din(n1914));
	jspl jspl_w_n1915_0(.douta(w_n1915_0[0]),.doutb(w_n1915_0[1]),.din(n1915));
	jspl jspl_w_n1917_0(.douta(w_n1917_0[0]),.doutb(w_n1917_0[1]),.din(n1917));
	jspl jspl_w_n1918_0(.douta(w_n1918_0[0]),.doutb(w_n1918_0[1]),.din(n1918));
	jspl jspl_w_n1920_0(.douta(w_n1920_0[0]),.doutb(w_n1920_0[1]),.din(n1920));
	jspl jspl_w_n1921_0(.douta(w_n1921_0[0]),.doutb(w_n1921_0[1]),.din(n1921));
	jspl jspl_w_n1930_0(.douta(w_n1930_0[0]),.doutb(w_n1930_0[1]),.din(n1930));
	jspl jspl_w_n1938_0(.douta(w_n1938_0[0]),.doutb(w_n1938_0[1]),.din(n1938));
	jspl jspl_w_n1940_0(.douta(w_n1940_0[0]),.doutb(w_n1940_0[1]),.din(n1940));
	jspl jspl_w_n1948_0(.douta(w_n1948_0[0]),.doutb(w_n1948_0[1]),.din(n1948));
	jspl jspl_w_n1950_0(.douta(w_n1950_0[0]),.doutb(w_n1950_0[1]),.din(n1950));
	jspl jspl_w_n1952_0(.douta(w_n1952_0[0]),.doutb(w_n1952_0[1]),.din(n1952));
	jspl jspl_w_n1953_0(.douta(w_n1953_0[0]),.doutb(w_n1953_0[1]),.din(n1953));
	jspl jspl_w_n1955_0(.douta(w_n1955_0[0]),.doutb(w_n1955_0[1]),.din(n1955));
	jspl jspl_w_n1956_0(.douta(w_n1956_0[0]),.doutb(w_n1956_0[1]),.din(n1956));
	jspl jspl_w_n1958_0(.douta(w_n1958_0[0]),.doutb(w_n1958_0[1]),.din(n1958));
	jspl jspl_w_n1959_0(.douta(w_n1959_0[0]),.doutb(w_n1959_0[1]),.din(n1959));
	jspl jspl_w_n1961_0(.douta(w_n1961_0[0]),.doutb(w_n1961_0[1]),.din(n1961));
	jspl jspl_w_n1962_0(.douta(w_n1962_0[0]),.doutb(w_n1962_0[1]),.din(n1962));
	jspl jspl_w_n1964_0(.douta(w_n1964_0[0]),.doutb(w_n1964_0[1]),.din(n1964));
	jspl jspl_w_n1965_0(.douta(w_n1965_0[0]),.doutb(w_n1965_0[1]),.din(n1965));
	jspl jspl_w_n1973_0(.douta(w_n1973_0[0]),.doutb(w_n1973_0[1]),.din(n1973));
	jspl jspl_w_n1975_0(.douta(w_n1975_0[0]),.doutb(w_n1975_0[1]),.din(n1975));
	jspl jspl_w_n1981_0(.douta(w_n1981_0[0]),.doutb(w_n1981_0[1]),.din(n1981));
	jspl jspl_w_n1989_0(.douta(w_n1989_0[0]),.doutb(w_n1989_0[1]),.din(n1989));
	jspl jspl_w_n1991_0(.douta(w_n1991_0[0]),.doutb(w_n1991_0[1]),.din(n1991));
	jspl jspl_w_n1999_0(.douta(w_n1999_0[0]),.doutb(w_n1999_0[1]),.din(n1999));
	jspl jspl_w_n2001_0(.douta(w_n2001_0[0]),.doutb(w_n2001_0[1]),.din(n2001));
	jspl jspl_w_n2002_0(.douta(w_n2002_0[0]),.doutb(w_n2002_0[1]),.din(n2002));
	jspl jspl_w_n2004_0(.douta(w_n2004_0[0]),.doutb(w_n2004_0[1]),.din(n2004));
	jspl jspl_w_n2005_0(.douta(w_n2005_0[0]),.doutb(w_n2005_0[1]),.din(n2005));
	jspl jspl_w_n2007_0(.douta(w_n2007_0[0]),.doutb(w_n2007_0[1]),.din(n2007));
	jspl jspl_w_n2008_0(.douta(w_n2008_0[0]),.doutb(w_n2008_0[1]),.din(n2008));
	jspl jspl_w_n2010_0(.douta(w_n2010_0[0]),.doutb(w_n2010_0[1]),.din(n2010));
	jspl3 jspl3_w_n2011_0(.douta(w_n2011_0[0]),.doutb(w_n2011_0[1]),.doutc(w_n2011_0[2]),.din(n2011));
	jspl jspl_w_n2013_0(.douta(w_n2013_0[0]),.doutb(w_n2013_0[1]),.din(n2013));
	jspl jspl_w_n2014_0(.douta(w_n2014_0[0]),.doutb(w_n2014_0[1]),.din(n2014));
	jspl jspl_w_n2020_0(.douta(w_n2020_0[0]),.doutb(w_n2020_0[1]),.din(n2020));
	jspl jspl_w_n2021_0(.douta(w_n2021_0[0]),.doutb(w_n2021_0[1]),.din(n2021));
	jspl jspl_w_n2029_0(.douta(w_n2029_0[0]),.doutb(w_n2029_0[1]),.din(n2029));
	jspl jspl_w_n2031_0(.douta(w_n2031_0[0]),.doutb(w_n2031_0[1]),.din(n2031));
	jspl jspl_w_n2033_0(.douta(w_n2033_0[0]),.doutb(w_n2033_0[1]),.din(n2033));
	jspl jspl_w_n2034_0(.douta(w_n2034_0[0]),.doutb(w_n2034_0[1]),.din(n2034));
	jspl jspl_w_n2036_0(.douta(w_n2036_0[0]),.doutb(w_n2036_0[1]),.din(n2036));
	jspl jspl_w_n2037_0(.douta(w_n2037_0[0]),.doutb(w_n2037_0[1]),.din(n2037));
	jspl jspl_w_n2039_0(.douta(w_n2039_0[0]),.doutb(w_n2039_0[1]),.din(n2039));
	jspl jspl_w_n2047_0(.douta(w_n2047_0[0]),.doutb(w_n2047_0[1]),.din(n2047));
	jspl jspl_w_n2055_0(.douta(w_n2055_0[0]),.doutb(w_n2055_0[1]),.din(n2055));
	jspl jspl_w_n2057_0(.douta(w_n2057_0[0]),.doutb(w_n2057_0[1]),.din(n2057));
	jspl jspl_w_n2065_0(.douta(w_n2065_0[0]),.doutb(w_n2065_0[1]),.din(n2065));
	jspl jspl_w_n2067_0(.douta(w_n2067_0[0]),.doutb(w_n2067_0[1]),.din(n2067));
	jspl jspl_w_n2068_0(.douta(w_n2068_0[0]),.doutb(w_n2068_0[1]),.din(n2068));
	jspl jspl_w_n2070_0(.douta(w_n2070_0[0]),.doutb(w_n2070_0[1]),.din(n2070));
	jspl jspl_w_n2071_0(.douta(w_n2071_0[0]),.doutb(w_n2071_0[1]),.din(n2071));
	jspl jspl_w_n2073_0(.douta(w_n2073_0[0]),.doutb(w_n2073_0[1]),.din(n2073));
	jspl jspl_w_n2074_0(.douta(w_n2074_0[0]),.doutb(w_n2074_0[1]),.din(n2074));
	jspl jspl_w_n2075_0(.douta(w_n2075_0[0]),.doutb(w_n2075_0[1]),.din(n2075));
	jspl jspl_w_n2081_0(.douta(w_n2081_0[0]),.doutb(w_n2081_0[1]),.din(n2081));
	jspl jspl_w_n2089_0(.douta(w_n2089_0[0]),.doutb(w_n2089_0[1]),.din(n2089));
	jspl jspl_w_n2091_0(.douta(w_n2091_0[0]),.doutb(w_n2091_0[1]),.din(n2091));
	jspl jspl_w_n2099_0(.douta(w_n2099_0[0]),.doutb(w_n2099_0[1]),.din(n2099));
	jspl jspl_w_n2101_0(.douta(w_n2101_0[0]),.doutb(w_n2101_0[1]),.din(n2101));
	jspl jspl_w_n2103_0(.douta(w_n2103_0[0]),.doutb(w_n2103_0[1]),.din(n2103));
	jspl jspl_w_n2104_0(.douta(w_n2104_0[0]),.doutb(w_n2104_0[1]),.din(n2104));
	jspl jspl_w_n2106_0(.douta(w_n2106_0[0]),.doutb(w_n2106_0[1]),.din(n2106));
	jspl3 jspl3_w_n2107_0(.douta(w_n2107_0[0]),.doutb(w_n2107_0[1]),.doutc(w_n2107_0[2]),.din(n2107));
	jspl jspl_w_n2109_0(.douta(w_n2109_0[0]),.doutb(w_n2109_0[1]),.din(n2109));
	jspl jspl_w_n2110_0(.douta(w_n2110_0[0]),.doutb(w_n2110_0[1]),.din(n2110));
	jspl jspl_w_n2116_0(.douta(w_n2116_0[0]),.doutb(w_n2116_0[1]),.din(n2116));
	jspl jspl_w_n2117_0(.douta(w_n2117_0[0]),.doutb(w_n2117_0[1]),.din(n2117));
	jspl jspl_w_n2125_0(.douta(w_n2125_0[0]),.doutb(w_n2125_0[1]),.din(n2125));
	jspl jspl_w_n2132_0(.douta(w_n2132_0[0]),.doutb(w_n2132_0[1]),.din(n2132));
	jspl jspl_w_n2134_0(.douta(w_n2134_0[0]),.doutb(w_n2134_0[1]),.din(n2134));
	jspl jspl_w_n2135_0(.douta(w_n2135_0[0]),.doutb(w_n2135_0[1]),.din(n2135));
	jspl jspl_w_n2137_0(.douta(w_n2137_0[0]),.doutb(w_n2137_0[1]),.din(n2137));
	jspl jspl_w_n2138_0(.douta(w_n2138_0[0]),.doutb(w_n2138_0[1]),.din(n2138));
	jspl jspl_w_n2140_0(.douta(w_n2140_0[0]),.doutb(w_n2140_0[1]),.din(n2140));
	jspl jspl_w_n2141_0(.douta(w_n2141_0[0]),.doutb(w_n2141_0[1]),.din(n2141));
	jspl jspl_w_n2142_0(.douta(w_n2142_0[0]),.doutb(w_n2142_0[1]),.din(n2142));
	jspl jspl_w_n2148_0(.douta(w_n2148_0[0]),.doutb(w_n2148_0[1]),.din(n2148));
	jspl jspl_w_n2155_0(.douta(w_n2155_0[0]),.doutb(w_n2155_0[1]),.din(n2155));
	jspl jspl_w_n2157_0(.douta(w_n2157_0[0]),.doutb(w_n2157_0[1]),.din(n2157));
	jspl jspl_w_n2159_0(.douta(w_n2159_0[0]),.doutb(w_n2159_0[1]),.din(n2159));
	jspl jspl_w_n2160_0(.douta(w_n2160_0[0]),.doutb(w_n2160_0[1]),.din(n2160));
	jspl jspl_w_n2166_0(.douta(w_n2166_0[0]),.doutb(w_n2166_0[1]),.din(n2166));
	jspl jspl_w_n2167_0(.douta(w_n2167_0[0]),.doutb(w_n2167_0[1]),.din(n2167));
	jspl jspl_w_n2168_0(.douta(w_n2168_0[0]),.doutb(w_n2168_0[1]),.din(n2168));
	jspl jspl_w_n2170_0(.douta(w_n2170_0[0]),.doutb(w_n2170_0[1]),.din(n2170));
	jspl jspl_w_n2171_0(.douta(w_n2171_0[0]),.doutb(w_n2171_0[1]),.din(n2171));
	jspl jspl_w_n2174_0(.douta(w_n2174_0[0]),.doutb(w_n2174_0[1]),.din(n2174));
	jspl jspl_w_n2180_0(.douta(w_n2180_0[0]),.doutb(w_n2180_0[1]),.din(n2180));
	jspl jspl_w_n2184_0(.douta(w_n2184_0[0]),.doutb(w_n2184_0[1]),.din(n2184));
	jspl jspl_w_n2187_0(.douta(w_n2187_0[0]),.doutb(w_n2187_0[1]),.din(n2187));
	jspl jspl_w_n2191_0(.douta(w_n2191_0[0]),.doutb(w_n2191_0[1]),.din(n2191));
	jspl jspl_w_n2197_0(.douta(w_n2197_0[0]),.doutb(w_n2197_0[1]),.din(n2197));
	jspl jspl_w_n2201_0(.douta(w_n2201_0[0]),.doutb(w_n2201_0[1]),.din(n2201));
	jspl jspl_w_n2208_0(.douta(w_n2208_0[0]),.doutb(w_n2208_0[1]),.din(n2208));
	jspl jspl_w_n2213_0(.douta(w_n2213_0[0]),.doutb(w_n2213_0[1]),.din(n2213));
	jspl jspl_w_n2218_0(.douta(w_n2218_0[0]),.doutb(w_n2218_0[1]),.din(n2218));
	jspl jspl_w_n2223_0(.douta(w_n2223_0[0]),.doutb(w_n2223_0[1]),.din(n2223));
	jspl jspl_w_n2228_0(.douta(w_n2228_0[0]),.doutb(w_n2228_0[1]),.din(n2228));
	jspl jspl_w_n2233_0(.douta(w_n2233_0[0]),.doutb(w_n2233_0[1]),.din(n2233));
	jspl jspl_w_n2238_0(.douta(w_n2238_0[0]),.doutb(w_n2238_0[1]),.din(n2238));
	jspl jspl_w_n2240_0(.douta(w_n2240_0[0]),.doutb(w_n2240_0[1]),.din(n2240));
	jspl jspl_w_n2241_0(.douta(w_n2241_0[0]),.doutb(w_n2241_0[1]),.din(n2241));
	jspl jspl_w_n2243_0(.douta(w_n2243_0[0]),.doutb(w_n2243_0[1]),.din(n2243));
	jspl jspl_w_n2244_0(.douta(w_n2244_0[0]),.doutb(w_n2244_0[1]),.din(n2244));
	jspl jspl_w_n2246_0(.douta(w_n2246_0[0]),.doutb(w_n2246_0[1]),.din(n2246));
	jspl jspl_w_n2247_0(.douta(w_n2247_0[0]),.doutb(w_n2247_0[1]),.din(n2247));
	jspl jspl_w_n2249_0(.douta(w_n2249_0[0]),.doutb(w_n2249_0[1]),.din(n2249));
	jspl jspl_w_n2250_0(.douta(w_n2250_0[0]),.doutb(w_n2250_0[1]),.din(n2250));
	jspl jspl_w_n2252_0(.douta(w_n2252_0[0]),.doutb(w_n2252_0[1]),.din(n2252));
	jspl jspl_w_n2253_0(.douta(w_n2253_0[0]),.doutb(w_n2253_0[1]),.din(n2253));
	jspl jspl_w_n2255_0(.douta(w_n2255_0[0]),.doutb(w_n2255_0[1]),.din(n2255));
	jspl jspl_w_n2256_0(.douta(w_n2256_0[0]),.doutb(w_n2256_0[1]),.din(n2256));
	jspl jspl_w_n2258_0(.douta(w_n2258_0[0]),.doutb(w_n2258_0[1]),.din(n2258));
	jspl jspl_w_n2259_0(.douta(w_n2259_0[0]),.doutb(w_n2259_0[1]),.din(n2259));
	jspl jspl_w_n2261_0(.douta(w_n2261_0[0]),.doutb(w_n2261_0[1]),.din(n2261));
	jspl jspl_w_n2262_0(.douta(w_n2262_0[0]),.doutb(w_n2262_0[1]),.din(n2262));
	jspl jspl_w_n2264_0(.douta(w_n2264_0[0]),.doutb(w_n2264_0[1]),.din(n2264));
	jspl jspl_w_n2267_0(.douta(w_n2267_0[0]),.doutb(w_n2267_0[1]),.din(n2267));
	jspl jspl_w_n2270_0(.douta(w_n2270_0[0]),.doutb(w_n2270_0[1]),.din(n2270));
	jspl jspl_w_n2278_0(.douta(w_n2278_0[0]),.doutb(w_n2278_0[1]),.din(n2278));
	jspl jspl_w_n2279_0(.douta(w_n2279_0[0]),.doutb(w_n2279_0[1]),.din(n2279));
	jspl jspl_w_n2280_0(.douta(w_n2280_0[0]),.doutb(w_n2280_0[1]),.din(n2280));
	jspl jspl_w_n2281_0(.douta(w_n2281_0[0]),.doutb(w_n2281_0[1]),.din(n2281));
	jspl jspl_w_n2282_0(.douta(w_n2282_0[0]),.doutb(w_n2282_0[1]),.din(n2282));
	jspl jspl_w_n2283_0(.douta(w_n2283_0[0]),.doutb(w_n2283_0[1]),.din(n2283));
	jspl jspl_w_n2284_0(.douta(w_n2284_0[0]),.doutb(w_n2284_0[1]),.din(n2284));
	jspl jspl_w_n2285_0(.douta(w_n2285_0[0]),.doutb(w_n2285_0[1]),.din(n2285));
	jspl jspl_w_n2286_0(.douta(w_n2286_0[0]),.doutb(w_n2286_0[1]),.din(n2286));
	jspl jspl_w_n2287_0(.douta(w_n2287_0[0]),.doutb(w_n2287_0[1]),.din(n2287));
	jspl jspl_w_n2289_0(.douta(w_n2289_0[0]),.doutb(w_n2289_0[1]),.din(n2289));
	jspl jspl_w_n2300_0(.douta(w_n2300_0[0]),.doutb(w_n2300_0[1]),.din(n2300));
	jspl jspl_w_n2302_0(.douta(w_n2302_0[0]),.doutb(w_n2302_0[1]),.din(n2302));
	jspl jspl_w_n2305_0(.douta(w_n2305_0[0]),.doutb(w_n2305_0[1]),.din(n2305));
	jspl jspl_w_n2307_0(.douta(w_n2307_0[0]),.doutb(w_n2307_0[1]),.din(n2307));
	jspl jspl_w_n2313_0(.douta(w_n2313_0[0]),.doutb(w_n2313_0[1]),.din(n2313));
	jspl jspl_w_n2315_0(.douta(w_n2315_0[0]),.doutb(w_n2315_0[1]),.din(n2315));
	jspl3 jspl3_w_n2321_0(.douta(w_n2321_0[0]),.doutb(w_n2321_0[1]),.doutc(w_n2321_0[2]),.din(n2321));
	jspl jspl_w_n2323_0(.douta(w_n2323_0[0]),.doutb(w_n2323_0[1]),.din(n2323));
	jspl3 jspl3_w_n2326_0(.douta(w_n2326_0[0]),.doutb(w_n2326_0[1]),.doutc(w_n2326_0[2]),.din(n2326));
	jspl jspl_w_n2330_0(.douta(w_n2330_0[0]),.doutb(w_n2330_0[1]),.din(n2330));
	jspl jspl_w_n2331_0(.douta(w_n2331_0[0]),.doutb(w_n2331_0[1]),.din(n2331));
	jspl jspl_w_n2332_0(.douta(w_n2332_0[0]),.doutb(w_n2332_0[1]),.din(n2332));
	jspl3 jspl3_w_n2334_0(.douta(w_n2334_0[0]),.doutb(w_n2334_0[1]),.doutc(w_n2334_0[2]),.din(n2334));
	jspl jspl_w_n2335_0(.douta(w_n2335_0[0]),.doutb(w_n2335_0[1]),.din(n2335));
	jspl jspl_w_n2339_0(.douta(w_n2339_0[0]),.doutb(w_n2339_0[1]),.din(n2339));
	jspl jspl_w_n2345_0(.douta(w_n2345_0[0]),.doutb(w_n2345_0[1]),.din(n2345));
	jspl jspl_w_n2347_0(.douta(w_n2347_0[0]),.doutb(w_n2347_0[1]),.din(n2347));
	jspl jspl_w_n2350_0(.douta(w_n2350_0[0]),.doutb(w_n2350_0[1]),.din(n2350));
	jspl jspl_w_n2351_0(.douta(w_n2351_0[0]),.doutb(w_n2351_0[1]),.din(n2351));
	jspl jspl_w_n2359_0(.douta(w_n2359_0[0]),.doutb(w_n2359_0[1]),.din(n2359));
	jspl jspl_w_n2360_0(.douta(w_n2360_0[0]),.doutb(w_n2360_0[1]),.din(n2360));
	jspl3 jspl3_w_n2365_0(.douta(w_n2365_0[0]),.doutb(w_n2365_0[1]),.doutc(w_n2365_0[2]),.din(n2365));
	jspl3 jspl3_w_n2372_0(.douta(w_n2372_0[0]),.doutb(w_n2372_0[1]),.doutc(w_n2372_0[2]),.din(n2372));
	jspl jspl_w_n2377_0(.douta(w_n2377_0[0]),.doutb(w_n2377_0[1]),.din(n2377));
	jspl jspl_w_n2379_0(.douta(w_n2379_0[0]),.doutb(w_n2379_0[1]),.din(n2379));
	jspl3 jspl3_w_n2380_0(.douta(w_n2380_0[0]),.doutb(w_n2380_0[1]),.doutc(w_n2380_0[2]),.din(n2380));
	jspl3 jspl3_w_n2380_1(.douta(w_n2380_1[0]),.doutb(w_n2380_1[1]),.doutc(w_n2380_1[2]),.din(w_n2380_0[0]));
	jspl3 jspl3_w_n2380_2(.douta(w_n2380_2[0]),.doutb(w_n2380_2[1]),.doutc(w_n2380_2[2]),.din(w_n2380_0[1]));
	jspl jspl_w_n2380_3(.douta(w_n2380_3[0]),.doutb(w_n2380_3[1]),.din(w_n2380_0[2]));
	jspl jspl_w_n2382_0(.douta(w_n2382_0[0]),.doutb(w_n2382_0[1]),.din(n2382));
	jspl3 jspl3_w_n2385_0(.douta(w_n2385_0[0]),.doutb(w_n2385_0[1]),.doutc(w_n2385_0[2]),.din(n2385));
	jspl jspl_w_n2385_1(.douta(w_n2385_1[0]),.doutb(w_n2385_1[1]),.din(w_n2385_0[0]));
	jspl jspl_w_n2387_0(.douta(w_n2387_0[0]),.doutb(w_n2387_0[1]),.din(n2387));
	jspl jspl_w_n2391_0(.douta(w_n2391_0[0]),.doutb(w_n2391_0[1]),.din(n2391));
	jspl jspl_w_n2396_0(.douta(w_n2396_0[0]),.doutb(w_n2396_0[1]),.din(n2396));
	jspl jspl_w_n2398_0(.douta(w_n2398_0[0]),.doutb(w_n2398_0[1]),.din(n2398));
	jspl jspl_w_n2402_0(.douta(w_n2402_0[0]),.doutb(w_n2402_0[1]),.din(n2402));
	jspl jspl_w_n2406_0(.douta(w_n2406_0[0]),.doutb(w_n2406_0[1]),.din(n2406));
	jspl jspl_w_n2412_0(.douta(w_n2412_0[0]),.doutb(w_n2412_0[1]),.din(n2412));
	jspl jspl_w_n2414_0(.douta(w_n2414_0[0]),.doutb(w_n2414_0[1]),.din(n2414));
	jspl3 jspl3_w_n2417_0(.douta(w_n2417_0[0]),.doutb(w_n2417_0[1]),.doutc(w_n2417_0[2]),.din(n2417));
	jspl jspl_w_n2424_0(.douta(w_n2424_0[0]),.doutb(w_n2424_0[1]),.din(n2424));
	jspl3 jspl3_w_n2427_0(.douta(w_n2427_0[0]),.doutb(w_n2427_0[1]),.doutc(w_n2427_0[2]),.din(n2427));
	jspl jspl_w_n2428_0(.douta(w_n2428_0[0]),.doutb(w_n2428_0[1]),.din(n2428));
	jspl3 jspl3_w_n2429_0(.douta(w_n2429_0[0]),.doutb(w_n2429_0[1]),.doutc(w_n2429_0[2]),.din(n2429));
	jspl jspl_w_n2429_1(.douta(w_n2429_1[0]),.doutb(w_n2429_1[1]),.din(w_n2429_0[0]));
	jspl jspl_w_n2438_0(.douta(w_n2438_0[0]),.doutb(w_n2438_0[1]),.din(n2438));
	jspl jspl_w_n2440_0(.douta(w_n2440_0[0]),.doutb(w_n2440_0[1]),.din(n2440));
	jspl jspl_w_n2442_0(.douta(w_n2442_0[0]),.doutb(w_n2442_0[1]),.din(n2442));
	jspl jspl_w_n2449_0(.douta(w_n2449_0[0]),.doutb(w_n2449_0[1]),.din(n2449));
	jspl jspl_w_n2451_0(.douta(w_n2451_0[0]),.doutb(w_n2451_0[1]),.din(n2451));
	jspl jspl_w_n2453_0(.douta(w_n2453_0[0]),.doutb(w_n2453_0[1]),.din(n2453));
	jspl3 jspl3_w_n2456_0(.douta(w_n2456_0[0]),.doutb(w_n2456_0[1]),.doutc(w_n2456_0[2]),.din(n2456));
	jspl jspl_w_n2457_0(.douta(w_n2457_0[0]),.doutb(w_n2457_0[1]),.din(n2457));
	jspl jspl_w_n2461_0(.douta(w_n2461_0[0]),.doutb(w_n2461_0[1]),.din(n2461));
	jspl jspl_w_n2466_0(.douta(w_n2466_0[0]),.doutb(w_n2466_0[1]),.din(n2466));
	jspl jspl_w_n2477_0(.douta(w_n2477_0[0]),.doutb(w_n2477_0[1]),.din(n2477));
	jspl3 jspl3_w_n2479_0(.douta(w_n2479_0[0]),.doutb(w_n2479_0[1]),.doutc(w_n2479_0[2]),.din(n2479));
	jspl jspl_w_n2486_0(.douta(w_n2486_0[0]),.doutb(w_n2486_0[1]),.din(n2486));
	jspl jspl_w_n2490_0(.douta(w_n2490_0[0]),.doutb(w_n2490_0[1]),.din(n2490));
	jspl jspl_w_n2498_0(.douta(w_n2498_0[0]),.doutb(w_n2498_0[1]),.din(n2498));
	jspl3 jspl3_w_n2504_0(.douta(w_n2504_0[0]),.doutb(w_n2504_0[1]),.doutc(w_n2504_0[2]),.din(n2504));
	jspl jspl_w_n2506_0(.douta(w_n2506_0[0]),.doutb(w_n2506_0[1]),.din(n2506));
	jspl3 jspl3_w_n2511_0(.douta(w_n2511_0[0]),.doutb(w_n2511_0[1]),.doutc(w_n2511_0[2]),.din(n2511));
	jspl jspl_w_n2511_1(.douta(w_n2511_1[0]),.doutb(w_n2511_1[1]),.din(w_n2511_0[0]));
	jspl jspl_w_n2514_0(.douta(w_n2514_0[0]),.doutb(w_n2514_0[1]),.din(n2514));
	jspl3 jspl3_w_n2515_0(.douta(w_n2515_0[0]),.doutb(w_n2515_0[1]),.doutc(w_n2515_0[2]),.din(n2515));
	jspl3 jspl3_w_n2520_0(.douta(w_n2520_0[0]),.doutb(w_n2520_0[1]),.doutc(w_n2520_0[2]),.din(n2520));
	jspl3 jspl3_w_n2521_0(.douta(w_n2521_0[0]),.doutb(w_n2521_0[1]),.doutc(w_n2521_0[2]),.din(n2521));
	jspl jspl_w_n2521_1(.douta(w_n2521_1[0]),.doutb(w_n2521_1[1]),.din(w_n2521_0[0]));
	jspl jspl_w_n2534_0(.douta(w_n2534_0[0]),.doutb(w_n2534_0[1]),.din(n2534));
	jspl jspl_w_n2536_0(.douta(w_n2536_0[0]),.doutb(w_n2536_0[1]),.din(n2536));
	jspl jspl_w_n2538_0(.douta(w_n2538_0[0]),.doutb(w_n2538_0[1]),.din(n2538));
	jspl jspl_w_n2540_0(.douta(w_n2540_0[0]),.doutb(w_n2540_0[1]),.din(n2540));
	jspl jspl_w_n2541_0(.douta(w_n2541_0[0]),.doutb(w_n2541_0[1]),.din(n2541));
	jspl jspl_w_n2542_0(.douta(w_n2542_0[0]),.doutb(w_n2542_0[1]),.din(n2542));
	jspl jspl_w_n2544_0(.douta(w_n2544_0[0]),.doutb(w_n2544_0[1]),.din(n2544));
	jspl jspl_w_n2551_0(.douta(w_n2551_0[0]),.doutb(w_n2551_0[1]),.din(n2551));
	jspl jspl_w_n2552_0(.douta(w_n2552_0[0]),.doutb(w_n2552_0[1]),.din(n2552));
	jspl jspl_w_n2564_0(.douta(w_n2564_0[0]),.doutb(w_n2564_0[1]),.din(n2564));
	jspl jspl_w_n2566_0(.douta(w_n2566_0[0]),.doutb(w_n2566_0[1]),.din(n2566));
	jspl jspl_w_n2571_0(.douta(w_n2571_0[0]),.doutb(w_n2571_0[1]),.din(n2571));
	jspl3 jspl3_w_n2575_0(.douta(w_n2575_0[0]),.doutb(w_n2575_0[1]),.doutc(w_n2575_0[2]),.din(n2575));
	jspl jspl_w_n2580_0(.douta(w_n2580_0[0]),.doutb(w_n2580_0[1]),.din(n2580));
	jspl jspl_w_n2586_0(.douta(w_n2586_0[0]),.doutb(w_n2586_0[1]),.din(n2586));
	jspl jspl_w_n2587_0(.douta(w_n2587_0[0]),.doutb(w_n2587_0[1]),.din(n2587));
	jspl3 jspl3_w_n2589_0(.douta(w_n2589_0[0]),.doutb(w_n2589_0[1]),.doutc(w_n2589_0[2]),.din(n2589));
	jspl jspl_w_n2591_0(.douta(w_n2591_0[0]),.doutb(w_n2591_0[1]),.din(n2591));
	jspl jspl_w_n2593_0(.douta(w_n2593_0[0]),.doutb(w_n2593_0[1]),.din(n2593));
	jspl jspl_w_n2595_0(.douta(w_n2595_0[0]),.doutb(w_n2595_0[1]),.din(n2595));
	jspl jspl_w_n2599_0(.douta(w_n2599_0[0]),.doutb(w_n2599_0[1]),.din(n2599));
	jspl jspl_w_n2600_0(.douta(w_n2600_0[0]),.doutb(w_n2600_0[1]),.din(n2600));
	jspl3 jspl3_w_n2603_0(.douta(w_n2603_0[0]),.doutb(w_n2603_0[1]),.doutc(w_n2603_0[2]),.din(n2603));
	jspl jspl_w_n2604_0(.douta(w_n2604_0[0]),.doutb(w_n2604_0[1]),.din(n2604));
	jspl jspl_w_n2605_0(.douta(w_n2605_0[0]),.doutb(w_n2605_0[1]),.din(n2605));
	jspl jspl_w_n2607_0(.douta(w_n2607_0[0]),.doutb(w_n2607_0[1]),.din(n2607));
	jspl jspl_w_n2608_0(.douta(w_n2608_0[0]),.doutb(w_n2608_0[1]),.din(n2608));
	jspl jspl_w_n2611_0(.douta(w_n2611_0[0]),.doutb(w_n2611_0[1]),.din(n2611));
	jspl jspl_w_n2612_0(.douta(w_n2612_0[0]),.doutb(w_n2612_0[1]),.din(n2612));
	jspl jspl_w_n2615_0(.douta(w_n2615_0[0]),.doutb(w_n2615_0[1]),.din(n2615));
	jspl jspl_w_n2617_0(.douta(w_n2617_0[0]),.doutb(w_n2617_0[1]),.din(n2617));
	jspl jspl_w_n2620_0(.douta(w_n2620_0[0]),.doutb(w_n2620_0[1]),.din(n2620));
	jspl jspl_w_n2621_0(.douta(w_n2621_0[0]),.doutb(w_n2621_0[1]),.din(n2621));
	jspl jspl_w_n2624_0(.douta(w_n2624_0[0]),.doutb(w_n2624_0[1]),.din(n2624));
	jspl jspl_w_n2627_0(.douta(w_n2627_0[0]),.doutb(w_n2627_0[1]),.din(n2627));
	jspl jspl_w_n2630_0(.douta(w_n2630_0[0]),.doutb(w_n2630_0[1]),.din(n2630));
	jspl jspl_w_n2633_0(.douta(w_n2633_0[0]),.doutb(w_n2633_0[1]),.din(n2633));
	jspl jspl_w_n2634_0(.douta(w_n2634_0[0]),.doutb(w_n2634_0[1]),.din(n2634));
	jspl jspl_w_n2640_0(.douta(w_n2640_0[0]),.doutb(w_n2640_0[1]),.din(n2640));
	jspl jspl_w_n2641_0(.douta(w_n2641_0[0]),.doutb(w_n2641_0[1]),.din(n2641));
	jspl jspl_w_n2642_0(.douta(w_n2642_0[0]),.doutb(w_n2642_0[1]),.din(n2642));
	jspl jspl_w_n2643_0(.douta(w_n2643_0[0]),.doutb(w_n2643_0[1]),.din(n2643));
	jspl jspl_w_n2644_0(.douta(w_n2644_0[0]),.doutb(w_n2644_0[1]),.din(n2644));
	jspl jspl_w_n2655_0(.douta(w_n2655_0[0]),.doutb(w_n2655_0[1]),.din(n2655));
	jspl jspl_w_n2658_0(.douta(w_n2658_0[0]),.doutb(w_n2658_0[1]),.din(n2658));
	jspl jspl_w_n2665_0(.douta(w_n2665_0[0]),.doutb(w_n2665_0[1]),.din(n2665));
	jspl jspl_w_n2667_0(.douta(w_n2667_0[0]),.doutb(w_n2667_0[1]),.din(n2667));
	jspl jspl_w_n2668_0(.douta(w_n2668_0[0]),.doutb(w_n2668_0[1]),.din(n2668));
	jspl3 jspl3_w_n2669_0(.douta(w_n2669_0[0]),.doutb(w_n2669_0[1]),.doutc(w_n2669_0[2]),.din(n2669));
	jspl3 jspl3_w_n2669_1(.douta(w_n2669_1[0]),.doutb(w_n2669_1[1]),.doutc(w_n2669_1[2]),.din(w_n2669_0[0]));
	jspl3 jspl3_w_n2669_2(.douta(w_n2669_2[0]),.doutb(w_n2669_2[1]),.doutc(w_n2669_2[2]),.din(w_n2669_0[1]));
	jspl3 jspl3_w_n2669_3(.douta(w_n2669_3[0]),.doutb(w_n2669_3[1]),.doutc(w_n2669_3[2]),.din(w_n2669_0[2]));
	jspl3 jspl3_w_n2670_0(.douta(w_n2670_0[0]),.doutb(w_n2670_0[1]),.doutc(w_n2670_0[2]),.din(n2670));
	jspl3 jspl3_w_n2670_1(.douta(w_n2670_1[0]),.doutb(w_n2670_1[1]),.doutc(w_n2670_1[2]),.din(w_n2670_0[0]));
	jspl3 jspl3_w_n2670_2(.douta(w_n2670_2[0]),.doutb(w_n2670_2[1]),.doutc(w_n2670_2[2]),.din(w_n2670_0[1]));
	jspl3 jspl3_w_n2670_3(.douta(w_n2670_3[0]),.doutb(w_n2670_3[1]),.doutc(w_n2670_3[2]),.din(w_n2670_0[2]));
	jspl3 jspl3_w_n2670_4(.douta(w_n2670_4[0]),.doutb(w_n2670_4[1]),.doutc(w_n2670_4[2]),.din(w_n2670_1[0]));
	jspl3 jspl3_w_n2670_5(.douta(w_n2670_5[0]),.doutb(w_n2670_5[1]),.doutc(w_n2670_5[2]),.din(w_n2670_1[1]));
	jspl3 jspl3_w_n2671_0(.douta(w_n2671_0[0]),.doutb(w_n2671_0[1]),.doutc(w_n2671_0[2]),.din(n2671));
	jspl3 jspl3_w_n2671_1(.douta(w_n2671_1[0]),.doutb(w_n2671_1[1]),.doutc(w_n2671_1[2]),.din(w_n2671_0[0]));
	jspl3 jspl3_w_n2671_2(.douta(w_n2671_2[0]),.doutb(w_n2671_2[1]),.doutc(w_n2671_2[2]),.din(w_n2671_0[1]));
	jspl3 jspl3_w_n2671_3(.douta(w_n2671_3[0]),.doutb(w_n2671_3[1]),.doutc(w_n2671_3[2]),.din(w_n2671_0[2]));
	jspl3 jspl3_w_n2671_4(.douta(w_n2671_4[0]),.doutb(w_n2671_4[1]),.doutc(w_n2671_4[2]),.din(w_n2671_1[0]));
	jspl3 jspl3_w_n2671_5(.douta(w_n2671_5[0]),.doutb(w_n2671_5[1]),.doutc(w_n2671_5[2]),.din(w_n2671_1[1]));
	jspl jspl_w_n2671_6(.douta(w_n2671_6[0]),.doutb(w_n2671_6[1]),.din(w_n2671_1[2]));
	jspl3 jspl3_w_n2672_0(.douta(w_n2672_0[0]),.doutb(w_n2672_0[1]),.doutc(w_n2672_0[2]),.din(n2672));
	jspl3 jspl3_w_n2672_1(.douta(w_n2672_1[0]),.doutb(w_n2672_1[1]),.doutc(w_n2672_1[2]),.din(w_n2672_0[0]));
	jspl3 jspl3_w_n2672_2(.douta(w_n2672_2[0]),.doutb(w_n2672_2[1]),.doutc(w_n2672_2[2]),.din(w_n2672_0[1]));
	jspl3 jspl3_w_n2674_0(.douta(w_n2674_0[0]),.doutb(w_n2674_0[1]),.doutc(w_n2674_0[2]),.din(n2674));
	jspl3 jspl3_w_n2674_1(.douta(w_n2674_1[0]),.doutb(w_n2674_1[1]),.doutc(w_n2674_1[2]),.din(w_n2674_0[0]));
	jspl3 jspl3_w_n2674_2(.douta(w_n2674_2[0]),.doutb(w_n2674_2[1]),.doutc(w_n2674_2[2]),.din(w_n2674_0[1]));
	jspl3 jspl3_w_n2674_3(.douta(w_n2674_3[0]),.doutb(w_n2674_3[1]),.doutc(w_n2674_3[2]),.din(w_n2674_0[2]));
	jspl jspl_w_n2674_4(.douta(w_n2674_4[0]),.doutb(w_n2674_4[1]),.din(w_n2674_1[0]));
	jspl3 jspl3_w_n2677_0(.douta(w_n2677_0[0]),.doutb(w_n2677_0[1]),.doutc(w_n2677_0[2]),.din(n2677));
	jspl3 jspl3_w_n2677_1(.douta(w_n2677_1[0]),.doutb(w_n2677_1[1]),.doutc(w_n2677_1[2]),.din(w_n2677_0[0]));
	jspl3 jspl3_w_n2677_2(.douta(w_n2677_2[0]),.doutb(w_n2677_2[1]),.doutc(w_n2677_2[2]),.din(w_n2677_0[1]));
	jspl3 jspl3_w_n2677_3(.douta(w_n2677_3[0]),.doutb(w_n2677_3[1]),.doutc(w_n2677_3[2]),.din(w_n2677_0[2]));
	jspl3 jspl3_w_n2677_4(.douta(w_n2677_4[0]),.doutb(w_n2677_4[1]),.doutc(w_n2677_4[2]),.din(w_n2677_1[0]));
	jspl3 jspl3_w_n2678_0(.douta(w_n2678_0[0]),.doutb(w_n2678_0[1]),.doutc(w_n2678_0[2]),.din(n2678));
	jspl3 jspl3_w_n2678_1(.douta(w_n2678_1[0]),.doutb(w_n2678_1[1]),.doutc(w_n2678_1[2]),.din(w_n2678_0[0]));
	jspl3 jspl3_w_n2678_2(.douta(w_n2678_2[0]),.doutb(w_n2678_2[1]),.doutc(w_n2678_2[2]),.din(w_n2678_0[1]));
	jspl3 jspl3_w_n2678_3(.douta(w_n2678_3[0]),.doutb(w_n2678_3[1]),.doutc(w_n2678_3[2]),.din(w_n2678_0[2]));
	jspl3 jspl3_w_n2678_4(.douta(w_n2678_4[0]),.doutb(w_n2678_4[1]),.doutc(w_n2678_4[2]),.din(w_n2678_1[0]));
	jspl3 jspl3_w_n2678_5(.douta(w_n2678_5[0]),.doutb(w_n2678_5[1]),.doutc(w_n2678_5[2]),.din(w_n2678_1[1]));
	jspl jspl_w_n2678_6(.douta(w_n2678_6[0]),.doutb(w_n2678_6[1]),.din(w_n2678_1[2]));
	jspl3 jspl3_w_n2679_0(.douta(w_n2679_0[0]),.doutb(w_n2679_0[1]),.doutc(w_n2679_0[2]),.din(n2679));
	jspl3 jspl3_w_n2679_1(.douta(w_n2679_1[0]),.doutb(w_n2679_1[1]),.doutc(w_n2679_1[2]),.din(w_n2679_0[0]));
	jspl3 jspl3_w_n2679_2(.douta(w_n2679_2[0]),.doutb(w_n2679_2[1]),.doutc(w_n2679_2[2]),.din(w_n2679_0[1]));
	jspl jspl_w_n2679_3(.douta(w_n2679_3[0]),.doutb(w_n2679_3[1]),.din(w_n2679_0[2]));
	jspl3 jspl3_w_n2681_0(.douta(w_n2681_0[0]),.doutb(w_n2681_0[1]),.doutc(w_n2681_0[2]),.din(n2681));
	jspl3 jspl3_w_n2681_1(.douta(w_n2681_1[0]),.doutb(w_n2681_1[1]),.doutc(w_n2681_1[2]),.din(w_n2681_0[0]));
	jspl3 jspl3_w_n2681_2(.douta(w_n2681_2[0]),.doutb(w_n2681_2[1]),.doutc(w_n2681_2[2]),.din(w_n2681_0[1]));
	jspl3 jspl3_w_n2681_3(.douta(w_n2681_3[0]),.doutb(w_n2681_3[1]),.doutc(w_n2681_3[2]),.din(w_n2681_0[2]));
	jspl3 jspl3_w_n2681_4(.douta(w_n2681_4[0]),.doutb(w_n2681_4[1]),.doutc(w_n2681_4[2]),.din(w_n2681_1[0]));
	jspl jspl_w_n2681_5(.douta(w_n2681_5[0]),.doutb(w_n2681_5[1]),.din(w_n2681_1[1]));
	jspl3 jspl3_w_n2684_0(.douta(w_n2684_0[0]),.doutb(w_n2684_0[1]),.doutc(w_n2684_0[2]),.din(n2684));
	jspl3 jspl3_w_n2684_1(.douta(w_n2684_1[0]),.doutb(w_n2684_1[1]),.doutc(w_n2684_1[2]),.din(w_n2684_0[0]));
	jspl3 jspl3_w_n2684_2(.douta(w_n2684_2[0]),.doutb(w_n2684_2[1]),.doutc(w_n2684_2[2]),.din(w_n2684_0[1]));
	jspl3 jspl3_w_n2684_3(.douta(w_n2684_3[0]),.doutb(w_n2684_3[1]),.doutc(w_n2684_3[2]),.din(w_n2684_0[2]));
	jspl jspl_w_n2684_4(.douta(w_n2684_4[0]),.doutb(w_n2684_4[1]),.din(w_n2684_1[0]));
	jspl3 jspl3_w_n2685_0(.douta(w_n2685_0[0]),.doutb(w_n2685_0[1]),.doutc(w_n2685_0[2]),.din(n2685));
	jspl3 jspl3_w_n2685_1(.douta(w_n2685_1[0]),.doutb(w_n2685_1[1]),.doutc(w_n2685_1[2]),.din(w_n2685_0[0]));
	jspl jspl_w_n2685_2(.douta(w_n2685_2[0]),.doutb(w_n2685_2[1]),.din(w_n2685_0[1]));
	jspl3 jspl3_w_n2687_0(.douta(w_n2687_0[0]),.doutb(w_n2687_0[1]),.doutc(w_n2687_0[2]),.din(n2687));
	jspl3 jspl3_w_n2687_1(.douta(w_n2687_1[0]),.doutb(w_n2687_1[1]),.doutc(w_n2687_1[2]),.din(w_n2687_0[0]));
	jspl3 jspl3_w_n2687_2(.douta(w_n2687_2[0]),.doutb(w_n2687_2[1]),.doutc(w_n2687_2[2]),.din(w_n2687_0[1]));
	jspl3 jspl3_w_n2687_3(.douta(w_n2687_3[0]),.doutb(w_n2687_3[1]),.doutc(w_n2687_3[2]),.din(w_n2687_0[2]));
	jspl3 jspl3_w_n2687_4(.douta(w_n2687_4[0]),.doutb(w_n2687_4[1]),.doutc(w_n2687_4[2]),.din(w_n2687_1[0]));
	jspl3 jspl3_w_n2687_5(.douta(w_n2687_5[0]),.doutb(w_n2687_5[1]),.doutc(w_n2687_5[2]),.din(w_n2687_1[1]));
	jspl3 jspl3_w_n2687_6(.douta(w_n2687_6[0]),.doutb(w_n2687_6[1]),.doutc(w_n2687_6[2]),.din(w_n2687_1[2]));
	jspl jspl_w_n2687_7(.douta(w_n2687_7[0]),.doutb(w_n2687_7[1]),.din(w_n2687_2[0]));
	jspl3 jspl3_w_n2688_0(.douta(w_n2688_0[0]),.doutb(w_n2688_0[1]),.doutc(w_n2688_0[2]),.din(n2688));
	jspl3 jspl3_w_n2688_1(.douta(w_n2688_1[0]),.doutb(w_n2688_1[1]),.doutc(w_n2688_1[2]),.din(w_n2688_0[0]));
	jspl3 jspl3_w_n2688_2(.douta(w_n2688_2[0]),.doutb(w_n2688_2[1]),.doutc(w_n2688_2[2]),.din(w_n2688_0[1]));
	jspl3 jspl3_w_n2688_3(.douta(w_n2688_3[0]),.doutb(w_n2688_3[1]),.doutc(w_n2688_3[2]),.din(w_n2688_0[2]));
	jspl3 jspl3_w_n2688_4(.douta(w_n2688_4[0]),.doutb(w_n2688_4[1]),.doutc(w_n2688_4[2]),.din(w_n2688_1[0]));
	jspl3 jspl3_w_n2688_5(.douta(w_n2688_5[0]),.doutb(w_n2688_5[1]),.doutc(w_n2688_5[2]),.din(w_n2688_1[1]));
	jspl3 jspl3_w_n2688_6(.douta(w_n2688_6[0]),.doutb(w_n2688_6[1]),.doutc(w_n2688_6[2]),.din(w_n2688_1[2]));
	jspl3 jspl3_w_n2688_7(.douta(w_n2688_7[0]),.doutb(w_n2688_7[1]),.doutc(w_n2688_7[2]),.din(w_n2688_2[0]));
	jspl3 jspl3_w_n2688_8(.douta(w_n2688_8[0]),.doutb(w_n2688_8[1]),.doutc(w_n2688_8[2]),.din(w_n2688_2[1]));
	jspl3 jspl3_w_n2691_0(.douta(w_n2691_0[0]),.doutb(w_n2691_0[1]),.doutc(w_n2691_0[2]),.din(n2691));
	jspl3 jspl3_w_n2691_1(.douta(w_n2691_1[0]),.doutb(w_n2691_1[1]),.doutc(w_n2691_1[2]),.din(w_n2691_0[0]));
	jspl3 jspl3_w_n2691_2(.douta(w_n2691_2[0]),.doutb(w_n2691_2[1]),.doutc(w_n2691_2[2]),.din(w_n2691_0[1]));
	jspl3 jspl3_w_n2691_3(.douta(w_n2691_3[0]),.doutb(w_n2691_3[1]),.doutc(w_n2691_3[2]),.din(w_n2691_0[2]));
	jspl3 jspl3_w_n2691_4(.douta(w_n2691_4[0]),.doutb(w_n2691_4[1]),.doutc(w_n2691_4[2]),.din(w_n2691_1[0]));
	jspl3 jspl3_w_n2691_5(.douta(w_n2691_5[0]),.doutb(w_n2691_5[1]),.doutc(w_n2691_5[2]),.din(w_n2691_1[1]));
	jspl3 jspl3_w_n2691_6(.douta(w_n2691_6[0]),.doutb(w_n2691_6[1]),.doutc(w_n2691_6[2]),.din(w_n2691_1[2]));
	jspl3 jspl3_w_n2691_7(.douta(w_n2691_7[0]),.doutb(w_n2691_7[1]),.doutc(w_n2691_7[2]),.din(w_n2691_2[0]));
	jspl3 jspl3_w_n2691_8(.douta(w_n2691_8[0]),.doutb(w_n2691_8[1]),.doutc(w_n2691_8[2]),.din(w_n2691_2[1]));
	jspl3 jspl3_w_n2693_0(.douta(w_n2693_0[0]),.doutb(w_n2693_0[1]),.doutc(w_n2693_0[2]),.din(n2693));
	jspl3 jspl3_w_n2693_1(.douta(w_n2693_1[0]),.doutb(w_n2693_1[1]),.doutc(w_n2693_1[2]),.din(w_n2693_0[0]));
	jspl3 jspl3_w_n2693_2(.douta(w_n2693_2[0]),.doutb(w_n2693_2[1]),.doutc(w_n2693_2[2]),.din(w_n2693_0[1]));
	jspl3 jspl3_w_n2693_3(.douta(w_n2693_3[0]),.doutb(w_n2693_3[1]),.doutc(w_n2693_3[2]),.din(w_n2693_0[2]));
	jspl3 jspl3_w_n2693_4(.douta(w_n2693_4[0]),.doutb(w_n2693_4[1]),.doutc(w_n2693_4[2]),.din(w_n2693_1[0]));
	jspl3 jspl3_w_n2694_0(.douta(w_n2694_0[0]),.doutb(w_n2694_0[1]),.doutc(w_n2694_0[2]),.din(n2694));
	jspl3 jspl3_w_n2694_1(.douta(w_n2694_1[0]),.doutb(w_n2694_1[1]),.doutc(w_n2694_1[2]),.din(w_n2694_0[0]));
	jspl3 jspl3_w_n2694_2(.douta(w_n2694_2[0]),.doutb(w_n2694_2[1]),.doutc(w_n2694_2[2]),.din(w_n2694_0[1]));
	jspl3 jspl3_w_n2694_3(.douta(w_n2694_3[0]),.doutb(w_n2694_3[1]),.doutc(w_n2694_3[2]),.din(w_n2694_0[2]));
	jspl3 jspl3_w_n2694_4(.douta(w_n2694_4[0]),.doutb(w_n2694_4[1]),.doutc(w_n2694_4[2]),.din(w_n2694_1[0]));
	jspl3 jspl3_w_n2696_0(.douta(w_n2696_0[0]),.doutb(w_n2696_0[1]),.doutc(w_n2696_0[2]),.din(n2696));
	jspl3 jspl3_w_n2697_0(.douta(w_n2697_0[0]),.doutb(w_n2697_0[1]),.doutc(w_n2697_0[2]),.din(n2697));
	jspl jspl_w_n2697_1(.douta(w_n2697_1[0]),.doutb(w_n2697_1[1]),.din(w_n2697_0[0]));
	jspl3 jspl3_w_n2698_0(.douta(w_n2698_0[0]),.doutb(w_n2698_0[1]),.doutc(w_n2698_0[2]),.din(n2698));
	jspl3 jspl3_w_n2698_1(.douta(w_n2698_1[0]),.doutb(w_n2698_1[1]),.doutc(w_n2698_1[2]),.din(w_n2698_0[0]));
	jspl3 jspl3_w_n2698_2(.douta(w_n2698_2[0]),.doutb(w_n2698_2[1]),.doutc(w_n2698_2[2]),.din(w_n2698_0[1]));
	jspl3 jspl3_w_n2698_3(.douta(w_n2698_3[0]),.doutb(w_n2698_3[1]),.doutc(w_n2698_3[2]),.din(w_n2698_0[2]));
	jspl3 jspl3_w_n2698_4(.douta(w_n2698_4[0]),.doutb(w_n2698_4[1]),.doutc(w_n2698_4[2]),.din(w_n2698_1[0]));
	jspl3 jspl3_w_n2698_5(.douta(w_n2698_5[0]),.doutb(w_n2698_5[1]),.doutc(w_n2698_5[2]),.din(w_n2698_1[1]));
	jspl jspl_w_n2698_6(.douta(w_n2698_6[0]),.doutb(w_n2698_6[1]),.din(w_n2698_1[2]));
	jspl3 jspl3_w_n2700_0(.douta(w_n2700_0[0]),.doutb(w_n2700_0[1]),.doutc(w_n2700_0[2]),.din(n2700));
	jspl3 jspl3_w_n2700_1(.douta(w_n2700_1[0]),.doutb(w_n2700_1[1]),.doutc(w_n2700_1[2]),.din(w_n2700_0[0]));
	jspl3 jspl3_w_n2700_2(.douta(w_n2700_2[0]),.doutb(w_n2700_2[1]),.doutc(w_n2700_2[2]),.din(w_n2700_0[1]));
	jspl3 jspl3_w_n2700_3(.douta(w_n2700_3[0]),.doutb(w_n2700_3[1]),.doutc(w_n2700_3[2]),.din(w_n2700_0[2]));
	jspl3 jspl3_w_n2700_4(.douta(w_n2700_4[0]),.doutb(w_n2700_4[1]),.doutc(w_n2700_4[2]),.din(w_n2700_1[0]));
	jspl3 jspl3_w_n2700_5(.douta(w_n2700_5[0]),.doutb(w_n2700_5[1]),.doutc(w_n2700_5[2]),.din(w_n2700_1[1]));
	jspl jspl_w_n2701_0(.douta(w_n2701_0[0]),.doutb(w_n2701_0[1]),.din(n2701));
	jspl jspl_w_n2702_0(.douta(w_n2702_0[0]),.doutb(w_n2702_0[1]),.din(n2702));
	jspl jspl_w_n2704_0(.douta(w_n2704_0[0]),.doutb(w_n2704_0[1]),.din(n2704));
	jspl jspl_w_n2705_0(.douta(w_n2705_0[0]),.doutb(w_n2705_0[1]),.din(n2705));
	jspl jspl_w_n2708_0(.douta(w_n2708_0[0]),.doutb(w_n2708_0[1]),.din(n2708));
	jspl jspl_w_n2711_0(.douta(w_n2711_0[0]),.doutb(w_n2711_0[1]),.din(n2711));
	jspl jspl_w_n2713_0(.douta(w_n2713_0[0]),.doutb(w_n2713_0[1]),.din(n2713));
	jspl jspl_w_n2715_0(.douta(w_n2715_0[0]),.doutb(w_n2715_0[1]),.din(n2715));
	jspl jspl_w_n2718_0(.douta(w_n2718_0[0]),.doutb(w_n2718_0[1]),.din(n2718));
	jspl jspl_w_n2719_0(.douta(w_n2719_0[0]),.doutb(w_n2719_0[1]),.din(n2719));
	jspl jspl_w_n2721_0(.douta(w_n2721_0[0]),.doutb(w_n2721_0[1]),.din(n2721));
	jspl jspl_w_n2722_0(.douta(w_n2722_0[0]),.doutb(w_n2722_0[1]),.din(n2722));
	jspl jspl_w_n2724_0(.douta(w_n2724_0[0]),.doutb(w_n2724_0[1]),.din(n2724));
	jspl jspl_w_n2725_0(.douta(w_n2725_0[0]),.doutb(w_n2725_0[1]),.din(n2725));
	jspl jspl_w_n2727_0(.douta(w_n2727_0[0]),.doutb(w_n2727_0[1]),.din(n2727));
	jspl jspl_w_n2733_0(.douta(w_n2733_0[0]),.doutb(w_n2733_0[1]),.din(n2733));
	jspl3 jspl3_w_n2734_0(.douta(w_n2734_0[0]),.doutb(w_n2734_0[1]),.doutc(w_n2734_0[2]),.din(n2734));
	jspl3 jspl3_w_n2736_0(.douta(w_n2736_0[0]),.doutb(w_n2736_0[1]),.doutc(w_n2736_0[2]),.din(n2736));
	jspl jspl_w_n2736_1(.douta(w_n2736_1[0]),.doutb(w_n2736_1[1]),.din(w_n2736_0[0]));
	jspl jspl_w_n2743_0(.douta(w_n2743_0[0]),.doutb(w_n2743_0[1]),.din(n2743));
	jspl jspl_w_n2745_0(.douta(w_n2745_0[0]),.doutb(w_n2745_0[1]),.din(n2745));
	jspl3 jspl3_w_n2750_0(.douta(w_n2750_0[0]),.doutb(w_n2750_0[1]),.doutc(w_n2750_0[2]),.din(n2750));
	jspl jspl_w_n2751_0(.douta(w_n2751_0[0]),.doutb(w_n2751_0[1]),.din(n2751));
	jspl3 jspl3_w_n2752_0(.douta(w_n2752_0[0]),.doutb(w_n2752_0[1]),.doutc(w_n2752_0[2]),.din(n2752));
	jspl3 jspl3_w_n2767_0(.douta(w_n2767_0[0]),.doutb(w_n2767_0[1]),.doutc(w_n2767_0[2]),.din(n2767));
	jspl3 jspl3_w_n2769_0(.douta(w_n2769_0[0]),.doutb(w_n2769_0[1]),.doutc(w_n2769_0[2]),.din(n2769));
	jspl3 jspl3_w_n2769_1(.douta(w_n2769_1[0]),.doutb(w_n2769_1[1]),.doutc(w_n2769_1[2]),.din(w_n2769_0[0]));
	jspl3 jspl3_w_n2769_2(.douta(w_n2769_2[0]),.doutb(w_n2769_2[1]),.doutc(w_n2769_2[2]),.din(w_n2769_0[1]));
	jspl3 jspl3_w_n2769_3(.douta(w_n2769_3[0]),.doutb(w_n2769_3[1]),.doutc(w_n2769_3[2]),.din(w_n2769_0[2]));
	jspl jspl_w_n2769_4(.douta(w_n2769_4[0]),.doutb(w_n2769_4[1]),.din(w_n2769_1[0]));
	jspl3 jspl3_w_n2770_0(.douta(w_n2770_0[0]),.doutb(w_n2770_0[1]),.doutc(w_n2770_0[2]),.din(n2770));
	jspl3 jspl3_w_n2771_0(.douta(w_n2771_0[0]),.doutb(w_n2771_0[1]),.doutc(w_n2771_0[2]),.din(n2771));
	jspl3 jspl3_w_n2771_1(.douta(w_n2771_1[0]),.doutb(w_n2771_1[1]),.doutc(w_n2771_1[2]),.din(w_n2771_0[0]));
	jspl3 jspl3_w_n2773_0(.douta(w_n2773_0[0]),.doutb(w_n2773_0[1]),.doutc(w_n2773_0[2]),.din(n2773));
	jspl3 jspl3_w_n2773_1(.douta(w_n2773_1[0]),.doutb(w_n2773_1[1]),.doutc(w_n2773_1[2]),.din(w_n2773_0[0]));
	jspl3 jspl3_w_n2773_2(.douta(w_n2773_2[0]),.doutb(w_n2773_2[1]),.doutc(w_n2773_2[2]),.din(w_n2773_0[1]));
	jspl3 jspl3_w_n2773_3(.douta(w_n2773_3[0]),.doutb(w_n2773_3[1]),.doutc(w_n2773_3[2]),.din(w_n2773_0[2]));
	jspl3 jspl3_w_n2773_4(.douta(w_n2773_4[0]),.doutb(w_n2773_4[1]),.doutc(w_n2773_4[2]),.din(w_n2773_1[0]));
	jspl3 jspl3_w_n2774_0(.douta(w_n2774_0[0]),.doutb(w_n2774_0[1]),.doutc(w_n2774_0[2]),.din(n2774));
	jspl3 jspl3_w_n2774_1(.douta(w_n2774_1[0]),.doutb(w_n2774_1[1]),.doutc(w_n2774_1[2]),.din(w_n2774_0[0]));
	jspl jspl_w_n2774_2(.douta(w_n2774_2[0]),.doutb(w_n2774_2[1]),.din(w_n2774_0[1]));
	jspl3 jspl3_w_n2775_0(.douta(w_n2775_0[0]),.doutb(w_n2775_0[1]),.doutc(w_n2775_0[2]),.din(n2775));
	jspl3 jspl3_w_n2775_1(.douta(w_n2775_1[0]),.doutb(w_n2775_1[1]),.doutc(w_n2775_1[2]),.din(w_n2775_0[0]));
	jspl3 jspl3_w_n2775_2(.douta(w_n2775_2[0]),.doutb(w_n2775_2[1]),.doutc(w_n2775_2[2]),.din(w_n2775_0[1]));
	jspl3 jspl3_w_n2775_3(.douta(w_n2775_3[0]),.doutb(w_n2775_3[1]),.doutc(w_n2775_3[2]),.din(w_n2775_0[2]));
	jspl3 jspl3_w_n2775_4(.douta(w_n2775_4[0]),.doutb(w_n2775_4[1]),.doutc(w_n2775_4[2]),.din(w_n2775_1[0]));
	jspl3 jspl3_w_n2775_5(.douta(w_n2775_5[0]),.doutb(w_n2775_5[1]),.doutc(w_n2775_5[2]),.din(w_n2775_1[1]));
	jspl jspl_w_n2777_0(.douta(w_n2777_0[0]),.doutb(w_n2777_0[1]),.din(n2777));
	jspl3 jspl3_w_n2779_0(.douta(w_n2779_0[0]),.doutb(w_n2779_0[1]),.doutc(w_n2779_0[2]),.din(n2779));
	jspl3 jspl3_w_n2779_1(.douta(w_n2779_1[0]),.doutb(w_n2779_1[1]),.doutc(w_n2779_1[2]),.din(w_n2779_0[0]));
	jspl3 jspl3_w_n2779_2(.douta(w_n2779_2[0]),.doutb(w_n2779_2[1]),.doutc(w_n2779_2[2]),.din(w_n2779_0[1]));
	jspl3 jspl3_w_n2780_0(.douta(w_n2780_0[0]),.doutb(w_n2780_0[1]),.doutc(w_n2780_0[2]),.din(n2780));
	jspl3 jspl3_w_n2780_1(.douta(w_n2780_1[0]),.doutb(w_n2780_1[1]),.doutc(w_n2780_1[2]),.din(w_n2780_0[0]));
	jspl3 jspl3_w_n2780_2(.douta(w_n2780_2[0]),.doutb(w_n2780_2[1]),.doutc(w_n2780_2[2]),.din(w_n2780_0[1]));
	jspl3 jspl3_w_n2780_3(.douta(w_n2780_3[0]),.doutb(w_n2780_3[1]),.doutc(w_n2780_3[2]),.din(w_n2780_0[2]));
	jspl3 jspl3_w_n2780_4(.douta(w_n2780_4[0]),.doutb(w_n2780_4[1]),.doutc(w_n2780_4[2]),.din(w_n2780_1[0]));
	jspl3 jspl3_w_n2780_5(.douta(w_n2780_5[0]),.doutb(w_n2780_5[1]),.doutc(w_n2780_5[2]),.din(w_n2780_1[1]));
	jspl3 jspl3_w_n2783_0(.douta(w_n2783_0[0]),.doutb(w_n2783_0[1]),.doutc(w_n2783_0[2]),.din(n2783));
	jspl3 jspl3_w_n2783_1(.douta(w_n2783_1[0]),.doutb(w_n2783_1[1]),.doutc(w_n2783_1[2]),.din(w_n2783_0[0]));
	jspl jspl_w_n2783_2(.douta(w_n2783_2[0]),.doutb(w_n2783_2[1]),.din(w_n2783_0[1]));
	jspl3 jspl3_w_n2784_0(.douta(w_n2784_0[0]),.doutb(w_n2784_0[1]),.doutc(w_n2784_0[2]),.din(n2784));
	jspl3 jspl3_w_n2784_1(.douta(w_n2784_1[0]),.doutb(w_n2784_1[1]),.doutc(w_n2784_1[2]),.din(w_n2784_0[0]));
	jspl3 jspl3_w_n2784_2(.douta(w_n2784_2[0]),.doutb(w_n2784_2[1]),.doutc(w_n2784_2[2]),.din(w_n2784_0[1]));
	jspl3 jspl3_w_n2784_3(.douta(w_n2784_3[0]),.doutb(w_n2784_3[1]),.doutc(w_n2784_3[2]),.din(w_n2784_0[2]));
	jspl3 jspl3_w_n2784_4(.douta(w_n2784_4[0]),.doutb(w_n2784_4[1]),.doutc(w_n2784_4[2]),.din(w_n2784_1[0]));
	jspl3 jspl3_w_n2784_5(.douta(w_n2784_5[0]),.doutb(w_n2784_5[1]),.doutc(w_n2784_5[2]),.din(w_n2784_1[1]));
	jspl jspl_w_n2784_6(.douta(w_n2784_6[0]),.doutb(w_n2784_6[1]),.din(w_n2784_1[2]));
	jspl jspl_w_n2789_0(.douta(w_n2789_0[0]),.doutb(w_n2789_0[1]),.din(n2789));
	jspl3 jspl3_w_n2790_0(.douta(w_n2790_0[0]),.doutb(w_n2790_0[1]),.doutc(w_n2790_0[2]),.din(n2790));
	jspl3 jspl3_w_n2791_0(.douta(w_n2791_0[0]),.doutb(w_n2791_0[1]),.doutc(w_n2791_0[2]),.din(n2791));
	jspl jspl_w_n2792_0(.douta(w_n2792_0[0]),.doutb(w_n2792_0[1]),.din(n2792));
	jspl jspl_w_n2793_0(.douta(w_n2793_0[0]),.doutb(w_n2793_0[1]),.din(n2793));
	jspl3 jspl3_w_n2794_0(.douta(w_n2794_0[0]),.doutb(w_n2794_0[1]),.doutc(w_n2794_0[2]),.din(n2794));
	jspl3 jspl3_w_n2794_1(.douta(w_n2794_1[0]),.doutb(w_n2794_1[1]),.doutc(w_n2794_1[2]),.din(w_n2794_0[0]));
	jspl3 jspl3_w_n2794_2(.douta(w_n2794_2[0]),.doutb(w_n2794_2[1]),.doutc(w_n2794_2[2]),.din(w_n2794_0[1]));
	jspl3 jspl3_w_n2795_0(.douta(w_n2795_0[0]),.doutb(w_n2795_0[1]),.doutc(w_n2795_0[2]),.din(n2795));
	jspl3 jspl3_w_n2795_1(.douta(w_n2795_1[0]),.doutb(w_n2795_1[1]),.doutc(w_n2795_1[2]),.din(w_n2795_0[0]));
	jspl3 jspl3_w_n2795_2(.douta(w_n2795_2[0]),.doutb(w_n2795_2[1]),.doutc(w_n2795_2[2]),.din(w_n2795_0[1]));
	jspl3 jspl3_w_n2795_3(.douta(w_n2795_3[0]),.doutb(w_n2795_3[1]),.doutc(w_n2795_3[2]),.din(w_n2795_0[2]));
	jspl3 jspl3_w_n2795_4(.douta(w_n2795_4[0]),.doutb(w_n2795_4[1]),.doutc(w_n2795_4[2]),.din(w_n2795_1[0]));
	jspl3 jspl3_w_n2795_5(.douta(w_n2795_5[0]),.doutb(w_n2795_5[1]),.doutc(w_n2795_5[2]),.din(w_n2795_1[1]));
	jspl jspl_w_n2795_6(.douta(w_n2795_6[0]),.doutb(w_n2795_6[1]),.din(w_n2795_1[2]));
	jspl3 jspl3_w_n2797_0(.douta(w_n2797_0[0]),.doutb(w_n2797_0[1]),.doutc(w_n2797_0[2]),.din(n2797));
	jspl3 jspl3_w_n2797_1(.douta(w_n2797_1[0]),.doutb(w_n2797_1[1]),.doutc(w_n2797_1[2]),.din(w_n2797_0[0]));
	jspl3 jspl3_w_n2799_0(.douta(w_n2799_0[0]),.doutb(w_n2799_0[1]),.doutc(w_n2799_0[2]),.din(n2799));
	jspl3 jspl3_w_n2799_1(.douta(w_n2799_1[0]),.doutb(w_n2799_1[1]),.doutc(w_n2799_1[2]),.din(w_n2799_0[0]));
	jspl jspl_w_n2799_2(.douta(w_n2799_2[0]),.doutb(w_n2799_2[1]),.din(w_n2799_0[1]));
	jspl3 jspl3_w_n2800_0(.douta(w_n2800_0[0]),.doutb(w_n2800_0[1]),.doutc(w_n2800_0[2]),.din(n2800));
	jspl3 jspl3_w_n2800_1(.douta(w_n2800_1[0]),.doutb(w_n2800_1[1]),.doutc(w_n2800_1[2]),.din(w_n2800_0[0]));
	jspl3 jspl3_w_n2800_2(.douta(w_n2800_2[0]),.doutb(w_n2800_2[1]),.doutc(w_n2800_2[2]),.din(w_n2800_0[1]));
	jspl3 jspl3_w_n2800_3(.douta(w_n2800_3[0]),.doutb(w_n2800_3[1]),.doutc(w_n2800_3[2]),.din(w_n2800_0[2]));
	jspl3 jspl3_w_n2800_4(.douta(w_n2800_4[0]),.doutb(w_n2800_4[1]),.doutc(w_n2800_4[2]),.din(w_n2800_1[0]));
	jspl3 jspl3_w_n2800_5(.douta(w_n2800_5[0]),.doutb(w_n2800_5[1]),.doutc(w_n2800_5[2]),.din(w_n2800_1[1]));
	jspl jspl_w_n2802_0(.douta(w_n2802_0[0]),.doutb(w_n2802_0[1]),.din(n2802));
	jspl3 jspl3_w_n2804_0(.douta(w_n2804_0[0]),.doutb(w_n2804_0[1]),.doutc(w_n2804_0[2]),.din(n2804));
	jspl3 jspl3_w_n2804_1(.douta(w_n2804_1[0]),.doutb(w_n2804_1[1]),.doutc(w_n2804_1[2]),.din(w_n2804_0[0]));
	jspl3 jspl3_w_n2804_2(.douta(w_n2804_2[0]),.doutb(w_n2804_2[1]),.doutc(w_n2804_2[2]),.din(w_n2804_0[1]));
	jspl3 jspl3_w_n2805_0(.douta(w_n2805_0[0]),.doutb(w_n2805_0[1]),.doutc(w_n2805_0[2]),.din(n2805));
	jspl3 jspl3_w_n2805_1(.douta(w_n2805_1[0]),.doutb(w_n2805_1[1]),.doutc(w_n2805_1[2]),.din(w_n2805_0[0]));
	jspl3 jspl3_w_n2805_2(.douta(w_n2805_2[0]),.doutb(w_n2805_2[1]),.doutc(w_n2805_2[2]),.din(w_n2805_0[1]));
	jspl3 jspl3_w_n2805_3(.douta(w_n2805_3[0]),.doutb(w_n2805_3[1]),.doutc(w_n2805_3[2]),.din(w_n2805_0[2]));
	jspl3 jspl3_w_n2805_4(.douta(w_n2805_4[0]),.doutb(w_n2805_4[1]),.doutc(w_n2805_4[2]),.din(w_n2805_1[0]));
	jspl3 jspl3_w_n2805_5(.douta(w_n2805_5[0]),.doutb(w_n2805_5[1]),.doutc(w_n2805_5[2]),.din(w_n2805_1[1]));
	jspl3 jspl3_w_n2808_0(.douta(w_n2808_0[0]),.doutb(w_n2808_0[1]),.doutc(w_n2808_0[2]),.din(n2808));
	jspl3 jspl3_w_n2808_1(.douta(w_n2808_1[0]),.doutb(w_n2808_1[1]),.doutc(w_n2808_1[2]),.din(w_n2808_0[0]));
	jspl jspl_w_n2808_2(.douta(w_n2808_2[0]),.doutb(w_n2808_2[1]),.din(w_n2808_0[1]));
	jspl3 jspl3_w_n2809_0(.douta(w_n2809_0[0]),.doutb(w_n2809_0[1]),.doutc(w_n2809_0[2]),.din(n2809));
	jspl3 jspl3_w_n2809_1(.douta(w_n2809_1[0]),.doutb(w_n2809_1[1]),.doutc(w_n2809_1[2]),.din(w_n2809_0[0]));
	jspl3 jspl3_w_n2809_2(.douta(w_n2809_2[0]),.doutb(w_n2809_2[1]),.doutc(w_n2809_2[2]),.din(w_n2809_0[1]));
	jspl3 jspl3_w_n2809_3(.douta(w_n2809_3[0]),.doutb(w_n2809_3[1]),.doutc(w_n2809_3[2]),.din(w_n2809_0[2]));
	jspl3 jspl3_w_n2809_4(.douta(w_n2809_4[0]),.doutb(w_n2809_4[1]),.doutc(w_n2809_4[2]),.din(w_n2809_1[0]));
	jspl3 jspl3_w_n2809_5(.douta(w_n2809_5[0]),.doutb(w_n2809_5[1]),.doutc(w_n2809_5[2]),.din(w_n2809_1[1]));
	jspl jspl_w_n2809_6(.douta(w_n2809_6[0]),.doutb(w_n2809_6[1]),.din(w_n2809_1[2]));
	jspl jspl_w_n2815_0(.douta(w_n2815_0[0]),.doutb(w_n2815_0[1]),.din(n2815));
	jspl3 jspl3_w_n2816_0(.douta(w_n2816_0[0]),.doutb(w_n2816_0[1]),.doutc(w_n2816_0[2]),.din(n2816));
	jspl3 jspl3_w_n2817_0(.douta(w_n2817_0[0]),.doutb(w_n2817_0[1]),.doutc(w_n2817_0[2]),.din(n2817));
	jspl jspl_w_n2817_1(.douta(w_n2817_1[0]),.doutb(w_n2817_1[1]),.din(w_n2817_0[0]));
	jspl3 jspl3_w_n2818_0(.douta(w_n2818_0[0]),.doutb(w_n2818_0[1]),.doutc(w_n2818_0[2]),.din(n2818));
	jspl jspl_w_n2821_0(.douta(w_n2821_0[0]),.doutb(w_n2821_0[1]),.din(n2821));
	jspl jspl_w_n2822_0(.douta(w_n2822_0[0]),.doutb(w_n2822_0[1]),.din(n2822));
	jspl3 jspl3_w_n2823_0(.douta(w_n2823_0[0]),.doutb(w_n2823_0[1]),.doutc(w_n2823_0[2]),.din(n2823));
	jspl jspl_w_n2823_1(.douta(w_n2823_1[0]),.doutb(w_n2823_1[1]),.din(w_n2823_0[0]));
	jspl3 jspl3_w_n2824_0(.douta(w_n2824_0[0]),.doutb(w_n2824_0[1]),.doutc(w_n2824_0[2]),.din(n2824));
	jspl3 jspl3_w_n2825_0(.douta(w_n2825_0[0]),.doutb(w_n2825_0[1]),.doutc(w_n2825_0[2]),.din(n2825));
	jspl jspl_w_n2826_0(.douta(w_n2826_0[0]),.doutb(w_n2826_0[1]),.din(n2826));
	jspl jspl_w_n2827_0(.douta(w_n2827_0[0]),.doutb(w_n2827_0[1]),.din(n2827));
	jspl3 jspl3_w_n2828_0(.douta(w_n2828_0[0]),.doutb(w_n2828_0[1]),.doutc(w_n2828_0[2]),.din(n2828));
	jspl3 jspl3_w_n2828_1(.douta(w_n2828_1[0]),.doutb(w_n2828_1[1]),.doutc(w_n2828_1[2]),.din(w_n2828_0[0]));
	jspl3 jspl3_w_n2828_2(.douta(w_n2828_2[0]),.doutb(w_n2828_2[1]),.doutc(w_n2828_2[2]),.din(w_n2828_0[1]));
	jspl jspl_w_n2830_0(.douta(w_n2830_0[0]),.doutb(w_n2830_0[1]),.din(n2830));
	jspl3 jspl3_w_n2832_0(.douta(w_n2832_0[0]),.doutb(w_n2832_0[1]),.doutc(w_n2832_0[2]),.din(n2832));
	jspl3 jspl3_w_n2832_1(.douta(w_n2832_1[0]),.doutb(w_n2832_1[1]),.doutc(w_n2832_1[2]),.din(w_n2832_0[0]));
	jspl3 jspl3_w_n2832_2(.douta(w_n2832_2[0]),.doutb(w_n2832_2[1]),.doutc(w_n2832_2[2]),.din(w_n2832_0[1]));
	jspl3 jspl3_w_n2834_0(.douta(w_n2834_0[0]),.doutb(w_n2834_0[1]),.doutc(w_n2834_0[2]),.din(n2834));
	jspl3 jspl3_w_n2834_1(.douta(w_n2834_1[0]),.doutb(w_n2834_1[1]),.doutc(w_n2834_1[2]),.din(w_n2834_0[0]));
	jspl jspl_w_n2834_2(.douta(w_n2834_2[0]),.doutb(w_n2834_2[1]),.din(w_n2834_0[1]));
	jspl jspl_w_n2837_0(.douta(w_n2837_0[0]),.doutb(w_n2837_0[1]),.din(n2837));
	jspl3 jspl3_w_n2839_0(.douta(w_n2839_0[0]),.doutb(w_n2839_0[1]),.doutc(w_n2839_0[2]),.din(n2839));
	jspl jspl_w_n2839_1(.douta(w_n2839_1[0]),.doutb(w_n2839_1[1]),.din(w_n2839_0[0]));
	jspl jspl_w_n2842_0(.douta(w_n2842_0[0]),.doutb(w_n2842_0[1]),.din(n2842));
	jspl3 jspl3_w_n2844_0(.douta(w_n2844_0[0]),.doutb(w_n2844_0[1]),.doutc(w_n2844_0[2]),.din(n2844));
	jspl jspl_w_n2844_1(.douta(w_n2844_1[0]),.doutb(w_n2844_1[1]),.din(w_n2844_0[0]));
	jspl3 jspl3_w_n2848_0(.douta(w_n2848_0[0]),.doutb(w_n2848_0[1]),.doutc(w_n2848_0[2]),.din(n2848));
	jspl3 jspl3_w_n2848_1(.douta(w_n2848_1[0]),.doutb(w_n2848_1[1]),.doutc(w_n2848_1[2]),.din(w_n2848_0[0]));
	jspl jspl_w_n2848_2(.douta(w_n2848_2[0]),.doutb(w_n2848_2[1]),.din(w_n2848_0[1]));
	jspl jspl_w_n2854_0(.douta(w_n2854_0[0]),.doutb(w_n2854_0[1]),.din(n2854));
	jspl jspl_w_n2855_0(.douta(w_n2855_0[0]),.doutb(w_n2855_0[1]),.din(n2855));
	jspl3 jspl3_w_n2857_0(.douta(w_n2857_0[0]),.doutb(w_n2857_0[1]),.doutc(w_n2857_0[2]),.din(n2857));
	jspl3 jspl3_w_n2857_1(.douta(w_n2857_1[0]),.doutb(w_n2857_1[1]),.doutc(w_n2857_1[2]),.din(w_n2857_0[0]));
	jspl3 jspl3_w_n2857_2(.douta(w_n2857_2[0]),.doutb(w_n2857_2[1]),.doutc(w_n2857_2[2]),.din(w_n2857_0[1]));
	jspl3 jspl3_w_n2857_3(.douta(w_n2857_3[0]),.doutb(w_n2857_3[1]),.doutc(w_n2857_3[2]),.din(w_n2857_0[2]));
	jspl3 jspl3_w_n2857_4(.douta(w_n2857_4[0]),.doutb(w_n2857_4[1]),.doutc(w_n2857_4[2]),.din(w_n2857_1[0]));
	jspl3 jspl3_w_n2857_5(.douta(w_n2857_5[0]),.doutb(w_n2857_5[1]),.doutc(w_n2857_5[2]),.din(w_n2857_1[1]));
	jspl jspl_w_n2857_6(.douta(w_n2857_6[0]),.doutb(w_n2857_6[1]),.din(w_n2857_1[2]));
	jspl3 jspl3_w_n2858_0(.douta(w_n2858_0[0]),.doutb(w_n2858_0[1]),.doutc(w_n2858_0[2]),.din(n2858));
	jspl3 jspl3_w_n2858_1(.douta(w_n2858_1[0]),.doutb(w_n2858_1[1]),.doutc(w_n2858_1[2]),.din(w_n2858_0[0]));
	jspl3 jspl3_w_n2860_0(.douta(w_n2860_0[0]),.doutb(w_n2860_0[1]),.doutc(w_n2860_0[2]),.din(n2860));
	jspl3 jspl3_w_n2860_1(.douta(w_n2860_1[0]),.doutb(w_n2860_1[1]),.doutc(w_n2860_1[2]),.din(w_n2860_0[0]));
	jspl3 jspl3_w_n2860_2(.douta(w_n2860_2[0]),.doutb(w_n2860_2[1]),.doutc(w_n2860_2[2]),.din(w_n2860_0[1]));
	jspl3 jspl3_w_n2860_3(.douta(w_n2860_3[0]),.doutb(w_n2860_3[1]),.doutc(w_n2860_3[2]),.din(w_n2860_0[2]));
	jspl3 jspl3_w_n2860_4(.douta(w_n2860_4[0]),.doutb(w_n2860_4[1]),.doutc(w_n2860_4[2]),.din(w_n2860_1[0]));
	jspl3 jspl3_w_n2860_5(.douta(w_n2860_5[0]),.doutb(w_n2860_5[1]),.doutc(w_n2860_5[2]),.din(w_n2860_1[1]));
	jspl3 jspl3_w_n2862_0(.douta(w_n2862_0[0]),.doutb(w_n2862_0[1]),.doutc(w_n2862_0[2]),.din(n2862));
	jspl3 jspl3_w_n2862_1(.douta(w_n2862_1[0]),.doutb(w_n2862_1[1]),.doutc(w_n2862_1[2]),.din(w_n2862_0[0]));
	jspl3 jspl3_w_n2862_2(.douta(w_n2862_2[0]),.doutb(w_n2862_2[1]),.doutc(w_n2862_2[2]),.din(w_n2862_0[1]));
	jspl3 jspl3_w_n2863_0(.douta(w_n2863_0[0]),.doutb(w_n2863_0[1]),.doutc(w_n2863_0[2]),.din(n2863));
	jspl3 jspl3_w_n2863_1(.douta(w_n2863_1[0]),.doutb(w_n2863_1[1]),.doutc(w_n2863_1[2]),.din(w_n2863_0[0]));
	jspl3 jspl3_w_n2863_2(.douta(w_n2863_2[0]),.doutb(w_n2863_2[1]),.doutc(w_n2863_2[2]),.din(w_n2863_0[1]));
	jspl3 jspl3_w_n2863_3(.douta(w_n2863_3[0]),.doutb(w_n2863_3[1]),.doutc(w_n2863_3[2]),.din(w_n2863_0[2]));
	jspl3 jspl3_w_n2863_4(.douta(w_n2863_4[0]),.doutb(w_n2863_4[1]),.doutc(w_n2863_4[2]),.din(w_n2863_1[0]));
	jspl3 jspl3_w_n2863_5(.douta(w_n2863_5[0]),.doutb(w_n2863_5[1]),.doutc(w_n2863_5[2]),.din(w_n2863_1[1]));
	jspl jspl_w_n2863_6(.douta(w_n2863_6[0]),.doutb(w_n2863_6[1]),.din(w_n2863_1[2]));
	jspl3 jspl3_w_n2865_0(.douta(w_n2865_0[0]),.doutb(w_n2865_0[1]),.doutc(w_n2865_0[2]),.din(n2865));
	jspl3 jspl3_w_n2865_1(.douta(w_n2865_1[0]),.doutb(w_n2865_1[1]),.doutc(w_n2865_1[2]),.din(w_n2865_0[0]));
	jspl3 jspl3_w_n2865_2(.douta(w_n2865_2[0]),.doutb(w_n2865_2[1]),.doutc(w_n2865_2[2]),.din(w_n2865_0[1]));
	jspl3 jspl3_w_n2865_3(.douta(w_n2865_3[0]),.doutb(w_n2865_3[1]),.doutc(w_n2865_3[2]),.din(w_n2865_0[2]));
	jspl3 jspl3_w_n2865_4(.douta(w_n2865_4[0]),.doutb(w_n2865_4[1]),.doutc(w_n2865_4[2]),.din(w_n2865_1[0]));
	jspl3 jspl3_w_n2865_5(.douta(w_n2865_5[0]),.doutb(w_n2865_5[1]),.doutc(w_n2865_5[2]),.din(w_n2865_1[1]));
	jspl jspl_w_n2870_0(.douta(w_n2870_0[0]),.doutb(w_n2870_0[1]),.din(n2870));
	jspl jspl_w_n2871_0(.douta(w_n2871_0[0]),.doutb(w_n2871_0[1]),.din(n2871));
	jspl jspl_w_n2873_0(.douta(w_n2873_0[0]),.doutb(w_n2873_0[1]),.din(n2873));
	jspl3 jspl3_w_n2874_0(.douta(w_n2874_0[0]),.doutb(w_n2874_0[1]),.doutc(w_n2874_0[2]),.din(n2874));
	jspl3 jspl3_w_n2874_1(.douta(w_n2874_1[0]),.doutb(w_n2874_1[1]),.doutc(w_n2874_1[2]),.din(w_n2874_0[0]));
	jspl jspl_w_n2882_0(.douta(w_n2882_0[0]),.doutb(w_n2882_0[1]),.din(n2882));
	jspl3 jspl3_w_n2883_0(.douta(w_n2883_0[0]),.doutb(w_n2883_0[1]),.doutc(w_n2883_0[2]),.din(n2883));
	jspl3 jspl3_w_n2883_1(.douta(w_n2883_1[0]),.doutb(w_n2883_1[1]),.doutc(w_n2883_1[2]),.din(w_n2883_0[0]));
	jspl3 jspl3_w_n2883_2(.douta(w_n2883_2[0]),.doutb(w_n2883_2[1]),.doutc(w_n2883_2[2]),.din(w_n2883_0[1]));
	jspl jspl_w_n2883_3(.douta(w_n2883_3[0]),.doutb(w_n2883_3[1]),.din(w_n2883_0[2]));
	jspl jspl_w_n2885_0(.douta(w_n2885_0[0]),.doutb(w_n2885_0[1]),.din(n2885));
	jspl3 jspl3_w_n2887_0(.douta(w_n2887_0[0]),.doutb(w_n2887_0[1]),.doutc(w_n2887_0[2]),.din(n2887));
	jspl3 jspl3_w_n2887_1(.douta(w_n2887_1[0]),.doutb(w_n2887_1[1]),.doutc(w_n2887_1[2]),.din(w_n2887_0[0]));
	jspl3 jspl3_w_n2887_2(.douta(w_n2887_2[0]),.doutb(w_n2887_2[1]),.doutc(w_n2887_2[2]),.din(w_n2887_0[1]));
	jspl3 jspl3_w_n2887_3(.douta(w_n2887_3[0]),.doutb(w_n2887_3[1]),.doutc(w_n2887_3[2]),.din(w_n2887_0[2]));
	jspl3 jspl3_w_n2887_4(.douta(w_n2887_4[0]),.doutb(w_n2887_4[1]),.doutc(w_n2887_4[2]),.din(w_n2887_1[0]));
	jspl3 jspl3_w_n2889_0(.douta(w_n2889_0[0]),.doutb(w_n2889_0[1]),.doutc(w_n2889_0[2]),.din(n2889));
	jspl3 jspl3_w_n2889_1(.douta(w_n2889_1[0]),.doutb(w_n2889_1[1]),.doutc(w_n2889_1[2]),.din(w_n2889_0[0]));
	jspl3 jspl3_w_n2889_2(.douta(w_n2889_2[0]),.doutb(w_n2889_2[1]),.doutc(w_n2889_2[2]),.din(w_n2889_0[1]));
	jspl3 jspl3_w_n2889_3(.douta(w_n2889_3[0]),.doutb(w_n2889_3[1]),.doutc(w_n2889_3[2]),.din(w_n2889_0[2]));
	jspl jspl_w_n2889_4(.douta(w_n2889_4[0]),.doutb(w_n2889_4[1]),.din(w_n2889_1[0]));
	jspl jspl_w_n2892_0(.douta(w_n2892_0[0]),.doutb(w_n2892_0[1]),.din(n2892));
	jspl3 jspl3_w_n2893_0(.douta(w_n2893_0[0]),.doutb(w_n2893_0[1]),.doutc(w_n2893_0[2]),.din(n2893));
	jspl jspl_w_n2895_0(.douta(w_n2895_0[0]),.doutb(w_n2895_0[1]),.din(n2895));
	jspl jspl_w_n2896_0(.douta(w_n2896_0[0]),.doutb(w_n2896_0[1]),.din(n2896));
	jspl jspl_w_n2897_0(.douta(w_n2897_0[0]),.doutb(w_n2897_0[1]),.din(n2897));
	jspl3 jspl3_w_n2899_0(.douta(w_n2899_0[0]),.doutb(w_n2899_0[1]),.doutc(w_n2899_0[2]),.din(n2899));
	jspl3 jspl3_w_n2899_1(.douta(w_n2899_1[0]),.doutb(w_n2899_1[1]),.doutc(w_n2899_1[2]),.din(w_n2899_0[0]));
	jspl jspl_w_n2907_0(.douta(w_n2907_0[0]),.doutb(w_n2907_0[1]),.din(n2907));
	jspl jspl_w_n2908_0(.douta(w_n2908_0[0]),.doutb(w_n2908_0[1]),.din(n2908));
	jspl3 jspl3_w_n2911_0(.douta(w_n2911_0[0]),.doutb(w_n2911_0[1]),.doutc(w_n2911_0[2]),.din(n2911));
	jspl3 jspl3_w_n2911_1(.douta(w_n2911_1[0]),.doutb(w_n2911_1[1]),.doutc(w_n2911_1[2]),.din(w_n2911_0[0]));
	jspl jspl_w_n2920_0(.douta(w_n2920_0[0]),.doutb(w_n2920_0[1]),.din(n2920));
	jspl jspl_w_n2922_0(.douta(w_n2922_0[0]),.doutb(w_n2922_0[1]),.din(n2922));
	jspl jspl_w_n2931_0(.douta(w_n2931_0[0]),.doutb(w_n2931_0[1]),.din(n2931));
	jspl jspl_w_n2933_0(.douta(w_n2933_0[0]),.doutb(w_n2933_0[1]),.din(n2933));
	jspl jspl_w_n2939_0(.douta(w_n2939_0[0]),.doutb(w_n2939_0[1]),.din(n2939));
	jspl3 jspl3_w_n2941_0(.douta(w_n2941_0[0]),.doutb(w_n2941_0[1]),.doutc(w_n2941_0[2]),.din(n2941));
	jspl jspl_w_n2941_1(.douta(w_n2941_1[0]),.doutb(w_n2941_1[1]),.din(w_n2941_0[0]));
	jspl jspl_w_n2944_0(.douta(w_n2944_0[0]),.doutb(w_n2944_0[1]),.din(n2944));
	jspl jspl_w_n2952_0(.douta(w_n2952_0[0]),.doutb(w_n2952_0[1]),.din(n2952));
	jspl jspl_w_n2953_0(.douta(w_n2953_0[0]),.doutb(w_n2953_0[1]),.din(n2953));
	jspl jspl_w_n2963_0(.douta(w_n2963_0[0]),.doutb(w_n2963_0[1]),.din(n2963));
	jspl jspl_w_n2964_0(.douta(w_n2964_0[0]),.doutb(w_n2964_0[1]),.din(n2964));
	jspl jspl_w_n2966_0(.douta(w_n2966_0[0]),.doutb(w_n2966_0[1]),.din(n2966));
	jspl jspl_w_n2967_0(.douta(w_n2967_0[0]),.doutb(w_n2967_0[1]),.din(n2967));
	jspl jspl_w_n2969_0(.douta(w_n2969_0[0]),.doutb(w_n2969_0[1]),.din(n2969));
	jspl jspl_w_n2970_0(.douta(w_n2970_0[0]),.doutb(w_n2970_0[1]),.din(n2970));
	jspl jspl_w_n2972_0(.douta(w_n2972_0[0]),.doutb(w_n2972_0[1]),.din(n2972));
	jspl jspl_w_n2973_0(.douta(w_n2973_0[0]),.doutb(w_n2973_0[1]),.din(n2973));
	jspl jspl_w_n2975_0(.douta(w_n2975_0[0]),.doutb(w_n2975_0[1]),.din(n2975));
	jspl jspl_w_n2976_0(.douta(w_n2976_0[0]),.doutb(w_n2976_0[1]),.din(n2976));
	jspl jspl_w_n2978_0(.douta(w_n2978_0[0]),.doutb(w_n2978_0[1]),.din(n2978));
	jspl jspl_w_n2981_0(.douta(w_n2981_0[0]),.doutb(w_n2981_0[1]),.din(n2981));
	jspl jspl_w_n2989_0(.douta(w_n2989_0[0]),.doutb(w_n2989_0[1]),.din(n2989));
	jspl jspl_w_n2990_0(.douta(w_n2990_0[0]),.doutb(w_n2990_0[1]),.din(n2990));
	jspl3 jspl3_w_n2995_0(.douta(w_n2995_0[0]),.doutb(w_n2995_0[1]),.doutc(w_n2995_0[2]),.din(n2995));
	jspl3 jspl3_w_n2995_1(.douta(w_n2995_1[0]),.doutb(w_n2995_1[1]),.doutc(w_n2995_1[2]),.din(w_n2995_0[0]));
	jspl3 jspl3_w_n2995_2(.douta(w_n2995_2[0]),.doutb(w_n2995_2[1]),.doutc(w_n2995_2[2]),.din(w_n2995_0[1]));
	jspl3 jspl3_w_n2995_3(.douta(w_n2995_3[0]),.doutb(w_n2995_3[1]),.doutc(w_n2995_3[2]),.din(w_n2995_0[2]));
	jspl3 jspl3_w_n2995_4(.douta(w_n2995_4[0]),.doutb(w_n2995_4[1]),.doutc(w_n2995_4[2]),.din(w_n2995_1[0]));
	jspl jspl_w_n3000_0(.douta(w_n3000_0[0]),.doutb(w_n3000_0[1]),.din(n3000));
	jspl jspl_w_n3001_0(.douta(w_n3001_0[0]),.doutb(w_n3001_0[1]),.din(n3001));
	jspl jspl_w_n3002_0(.douta(w_n3002_0[0]),.doutb(w_n3002_0[1]),.din(n3002));
	jspl jspl_w_n3003_0(.douta(w_n3003_0[0]),.doutb(w_n3003_0[1]),.din(n3003));
	jspl3 jspl3_w_n3004_0(.douta(w_n3004_0[0]),.doutb(w_n3004_0[1]),.doutc(w_n3004_0[2]),.din(n3004));
	jspl3 jspl3_w_n3004_1(.douta(w_n3004_1[0]),.doutb(w_n3004_1[1]),.doutc(w_n3004_1[2]),.din(w_n3004_0[0]));
	jspl jspl_w_n3012_0(.douta(w_n3012_0[0]),.doutb(w_n3012_0[1]),.din(n3012));
	jspl jspl_w_n3013_0(.douta(w_n3013_0[0]),.doutb(w_n3013_0[1]),.din(n3013));
	jspl jspl_w_n3014_0(.douta(w_n3014_0[0]),.doutb(w_n3014_0[1]),.din(n3014));
	jspl3 jspl3_w_n3016_0(.douta(w_n3016_0[0]),.doutb(w_n3016_0[1]),.doutc(w_n3016_0[2]),.din(n3016));
	jspl3 jspl3_w_n3016_1(.douta(w_n3016_1[0]),.doutb(w_n3016_1[1]),.doutc(w_n3016_1[2]),.din(w_n3016_0[0]));
	jspl jspl_w_n3024_0(.douta(w_n3024_0[0]),.doutb(w_n3024_0[1]),.din(n3024));
	jspl jspl_w_n3025_0(.douta(w_n3025_0[0]),.doutb(w_n3025_0[1]),.din(n3025));
	jspl3 jspl3_w_n3028_0(.douta(w_n3028_0[0]),.doutb(w_n3028_0[1]),.doutc(w_n3028_0[2]),.din(n3028));
	jspl3 jspl3_w_n3028_1(.douta(w_n3028_1[0]),.doutb(w_n3028_1[1]),.doutc(w_n3028_1[2]),.din(w_n3028_0[0]));
	jspl jspl_w_n3036_0(.douta(w_n3036_0[0]),.doutb(w_n3036_0[1]),.din(n3036));
	jspl jspl_w_n3037_0(.douta(w_n3037_0[0]),.doutb(w_n3037_0[1]),.din(n3037));
	jspl jspl_w_n3046_0(.douta(w_n3046_0[0]),.doutb(w_n3046_0[1]),.din(n3046));
	jspl jspl_w_n3047_0(.douta(w_n3047_0[0]),.doutb(w_n3047_0[1]),.din(n3047));
	jspl jspl_w_n3056_0(.douta(w_n3056_0[0]),.doutb(w_n3056_0[1]),.din(n3056));
	jspl jspl_w_n3057_0(.douta(w_n3057_0[0]),.doutb(w_n3057_0[1]),.din(n3057));
	jspl jspl_w_n3066_0(.douta(w_n3066_0[0]),.doutb(w_n3066_0[1]),.din(n3066));
	jspl jspl_w_n3067_0(.douta(w_n3067_0[0]),.doutb(w_n3067_0[1]),.din(n3067));
	jspl jspl_w_n3076_0(.douta(w_n3076_0[0]),.doutb(w_n3076_0[1]),.din(n3076));
	jspl jspl_w_n3078_0(.douta(w_n3078_0[0]),.doutb(w_n3078_0[1]),.din(n3078));
	jspl jspl_w_n3087_0(.douta(w_n3087_0[0]),.doutb(w_n3087_0[1]),.din(n3087));
	jspl jspl_w_n3089_0(.douta(w_n3089_0[0]),.doutb(w_n3089_0[1]),.din(n3089));
	jspl jspl_w_n3095_0(.douta(w_n3095_0[0]),.doutb(w_n3095_0[1]),.din(n3095));
	jspl3 jspl3_w_n3097_0(.douta(w_n3097_0[0]),.doutb(w_n3097_0[1]),.doutc(w_n3097_0[2]),.din(n3097));
	jspl jspl_w_n3100_0(.douta(w_n3100_0[0]),.doutb(w_n3100_0[1]),.din(n3100));
	jspl jspl_w_n3107_0(.douta(w_n3107_0[0]),.doutb(w_n3107_0[1]),.din(n3107));
	jspl jspl_w_n3109_0(.douta(w_n3109_0[0]),.doutb(w_n3109_0[1]),.din(n3109));
	jspl jspl_w_n3118_0(.douta(w_n3118_0[0]),.doutb(w_n3118_0[1]),.din(n3118));
	jspl jspl_w_n3119_0(.douta(w_n3119_0[0]),.doutb(w_n3119_0[1]),.din(n3119));
	jspl jspl_w_n3121_0(.douta(w_n3121_0[0]),.doutb(w_n3121_0[1]),.din(n3121));
	jspl jspl_w_n3122_0(.douta(w_n3122_0[0]),.doutb(w_n3122_0[1]),.din(n3122));
	jspl jspl_w_n3124_0(.douta(w_n3124_0[0]),.doutb(w_n3124_0[1]),.din(n3124));
	jspl jspl_w_n3125_0(.douta(w_n3125_0[0]),.doutb(w_n3125_0[1]),.din(n3125));
	jspl jspl_w_n3127_0(.douta(w_n3127_0[0]),.doutb(w_n3127_0[1]),.din(n3127));
	jspl jspl_w_n3128_0(.douta(w_n3128_0[0]),.doutb(w_n3128_0[1]),.din(n3128));
	jspl jspl_w_n3130_0(.douta(w_n3130_0[0]),.doutb(w_n3130_0[1]),.din(n3130));
	jspl jspl_w_n3131_0(.douta(w_n3131_0[0]),.doutb(w_n3131_0[1]),.din(n3131));
	jspl jspl_w_n3133_0(.douta(w_n3133_0[0]),.doutb(w_n3133_0[1]),.din(n3133));
	jspl jspl_w_n3134_0(.douta(w_n3134_0[0]),.doutb(w_n3134_0[1]),.din(n3134));
	jspl jspl_w_n3136_0(.douta(w_n3136_0[0]),.doutb(w_n3136_0[1]),.din(n3136));
	jspl jspl_w_n3137_0(.douta(w_n3137_0[0]),.doutb(w_n3137_0[1]),.din(n3137));
	jspl jspl_w_n3139_0(.douta(w_n3139_0[0]),.doutb(w_n3139_0[1]),.din(n3139));
	jspl jspl_w_n3140_0(.douta(w_n3140_0[0]),.doutb(w_n3140_0[1]),.din(n3140));
	jspl jspl_w_n3142_0(.douta(w_n3142_0[0]),.doutb(w_n3142_0[1]),.din(n3142));
	jspl jspl_w_n3143_0(.douta(w_n3143_0[0]),.doutb(w_n3143_0[1]),.din(n3143));
	jspl jspl_w_n3145_0(.douta(w_n3145_0[0]),.doutb(w_n3145_0[1]),.din(n3145));
	jspl jspl_w_n3148_0(.douta(w_n3148_0[0]),.doutb(w_n3148_0[1]),.din(n3148));
	jspl jspl_w_n3154_0(.douta(w_n3154_0[0]),.doutb(w_n3154_0[1]),.din(n3154));
	jspl jspl_w_n3155_0(.douta(w_n3155_0[0]),.doutb(w_n3155_0[1]),.din(n3155));
	jspl jspl_w_n3159_0(.douta(w_n3159_0[0]),.doutb(w_n3159_0[1]),.din(n3159));
	jspl jspl_w_n3171_0(.douta(w_n3171_0[0]),.doutb(w_n3171_0[1]),.din(n3171));
	jspl3 jspl3_w_n3172_0(.douta(w_n3172_0[0]),.doutb(w_n3172_0[1]),.doutc(w_n3172_0[2]),.din(n3172));
	jspl3 jspl3_w_n3172_1(.douta(w_n3172_1[0]),.doutb(w_n3172_1[1]),.doutc(w_n3172_1[2]),.din(w_n3172_0[0]));
	jspl3 jspl3_w_n3172_2(.douta(w_n3172_2[0]),.doutb(w_n3172_2[1]),.doutc(w_n3172_2[2]),.din(w_n3172_0[1]));
	jspl3 jspl3_w_n3172_3(.douta(w_n3172_3[0]),.doutb(w_n3172_3[1]),.doutc(w_n3172_3[2]),.din(w_n3172_0[2]));
	jspl3 jspl3_w_n3172_4(.douta(w_n3172_4[0]),.doutb(w_n3172_4[1]),.doutc(w_n3172_4[2]),.din(w_n3172_1[0]));
	jspl3 jspl3_w_n3172_5(.douta(w_n3172_5[0]),.doutb(w_n3172_5[1]),.doutc(w_n3172_5[2]),.din(w_n3172_1[1]));
	jspl jspl_w_n3172_6(.douta(w_n3172_6[0]),.doutb(w_n3172_6[1]),.din(w_n3172_1[2]));
	jspl jspl_w_n3173_0(.douta(w_n3173_0[0]),.doutb(w_n3173_0[1]),.din(n3173));
	jspl3 jspl3_w_n3174_0(.douta(w_n3174_0[0]),.doutb(w_n3174_0[1]),.doutc(w_n3174_0[2]),.din(n3174));
	jspl3 jspl3_w_n3174_1(.douta(w_n3174_1[0]),.doutb(w_n3174_1[1]),.doutc(w_n3174_1[2]),.din(w_n3174_0[0]));
	jspl3 jspl3_w_n3176_0(.douta(w_n3176_0[0]),.doutb(w_n3176_0[1]),.doutc(w_n3176_0[2]),.din(n3176));
	jspl3 jspl3_w_n3176_1(.douta(w_n3176_1[0]),.doutb(w_n3176_1[1]),.doutc(w_n3176_1[2]),.din(w_n3176_0[0]));
	jspl3 jspl3_w_n3176_2(.douta(w_n3176_2[0]),.doutb(w_n3176_2[1]),.doutc(w_n3176_2[2]),.din(w_n3176_0[1]));
	jspl jspl_w_n3183_0(.douta(w_n3183_0[0]),.doutb(w_n3183_0[1]),.din(n3183));
	jspl jspl_w_n3186_0(.douta(w_n3186_0[0]),.doutb(w_n3186_0[1]),.din(n3186));
	jspl jspl_w_n3189_0(.douta(w_n3189_0[0]),.doutb(w_n3189_0[1]),.din(n3189));
	jspl jspl_w_n3197_0(.douta(w_n3197_0[0]),.doutb(w_n3197_0[1]),.din(n3197));
	jspl3 jspl3_w_n3198_0(.douta(w_n3198_0[0]),.doutb(w_n3198_0[1]),.doutc(w_n3198_0[2]),.din(n3198));
	jspl3 jspl3_w_n3198_1(.douta(w_n3198_1[0]),.doutb(w_n3198_1[1]),.doutc(w_n3198_1[2]),.din(w_n3198_0[0]));
	jspl3 jspl3_w_n3198_2(.douta(w_n3198_2[0]),.doutb(w_n3198_2[1]),.doutc(w_n3198_2[2]),.din(w_n3198_0[1]));
	jspl3 jspl3_w_n3198_3(.douta(w_n3198_3[0]),.doutb(w_n3198_3[1]),.doutc(w_n3198_3[2]),.din(w_n3198_0[2]));
	jspl3 jspl3_w_n3198_4(.douta(w_n3198_4[0]),.doutb(w_n3198_4[1]),.doutc(w_n3198_4[2]),.din(w_n3198_1[0]));
	jspl3 jspl3_w_n3198_5(.douta(w_n3198_5[0]),.doutb(w_n3198_5[1]),.doutc(w_n3198_5[2]),.din(w_n3198_1[1]));
	jspl3 jspl3_w_n3200_0(.douta(w_n3200_0[0]),.doutb(w_n3200_0[1]),.doutc(w_n3200_0[2]),.din(n3200));
	jspl3 jspl3_w_n3200_1(.douta(w_n3200_1[0]),.doutb(w_n3200_1[1]),.doutc(w_n3200_1[2]),.din(w_n3200_0[0]));
	jspl3 jspl3_w_n3200_2(.douta(w_n3200_2[0]),.doutb(w_n3200_2[1]),.doutc(w_n3200_2[2]),.din(w_n3200_0[1]));
	jspl3 jspl3_w_n3200_3(.douta(w_n3200_3[0]),.doutb(w_n3200_3[1]),.doutc(w_n3200_3[2]),.din(w_n3200_0[2]));
	jspl3 jspl3_w_n3202_0(.douta(w_n3202_0[0]),.doutb(w_n3202_0[1]),.doutc(w_n3202_0[2]),.din(n3202));
	jspl3 jspl3_w_n3202_1(.douta(w_n3202_1[0]),.doutb(w_n3202_1[1]),.doutc(w_n3202_1[2]),.din(w_n3202_0[0]));
	jspl3 jspl3_w_n3202_2(.douta(w_n3202_2[0]),.doutb(w_n3202_2[1]),.doutc(w_n3202_2[2]),.din(w_n3202_0[1]));
	jspl3 jspl3_w_n3202_3(.douta(w_n3202_3[0]),.doutb(w_n3202_3[1]),.doutc(w_n3202_3[2]),.din(w_n3202_0[2]));
	jspl3 jspl3_w_n3204_0(.douta(w_n3204_0[0]),.doutb(w_n3204_0[1]),.doutc(w_n3204_0[2]),.din(n3204));
	jspl3 jspl3_w_n3204_1(.douta(w_n3204_1[0]),.doutb(w_n3204_1[1]),.doutc(w_n3204_1[2]),.din(w_n3204_0[0]));
	jspl3 jspl3_w_n3204_2(.douta(w_n3204_2[0]),.doutb(w_n3204_2[1]),.doutc(w_n3204_2[2]),.din(w_n3204_0[1]));
	jspl3 jspl3_w_n3204_3(.douta(w_n3204_3[0]),.doutb(w_n3204_3[1]),.doutc(w_n3204_3[2]),.din(w_n3204_0[2]));
	jspl jspl_w_n3210_0(.douta(w_n3210_0[0]),.doutb(w_n3210_0[1]),.din(n3210));
	jspl jspl_w_n3212_0(.douta(w_n3212_0[0]),.doutb(w_n3212_0[1]),.din(n3212));
	jspl jspl_w_n3215_0(.douta(w_n3215_0[0]),.doutb(w_n3215_0[1]),.din(n3215));
	jspl jspl_w_n3217_0(.douta(w_n3217_0[0]),.doutb(w_n3217_0[1]),.din(n3217));
	jspl jspl_w_n3218_0(.douta(w_n3218_0[0]),.doutb(w_n3218_0[1]),.din(n3218));
	jspl jspl_w_n3219_0(.douta(w_n3219_0[0]),.doutb(w_n3219_0[1]),.din(n3219));
	jspl jspl_w_n3220_0(.douta(w_n3220_0[0]),.doutb(w_n3220_0[1]),.din(n3220));
	jspl jspl_w_n3228_0(.douta(w_n3228_0[0]),.doutb(w_n3228_0[1]),.din(n3228));
	jspl jspl_w_n3229_0(.douta(w_n3229_0[0]),.doutb(w_n3229_0[1]),.din(n3229));
	jspl jspl_w_n3230_0(.douta(w_n3230_0[0]),.doutb(w_n3230_0[1]),.din(n3230));
	jspl jspl_w_n3231_0(.douta(w_n3231_0[0]),.doutb(w_n3231_0[1]),.din(n3231));
	jspl jspl_w_n3232_0(.douta(w_n3232_0[0]),.doutb(w_n3232_0[1]),.din(n3232));
	jspl3 jspl3_w_n3233_0(.douta(w_n3233_0[0]),.doutb(w_n3233_0[1]),.doutc(w_n3233_0[2]),.din(n3233));
	jspl3 jspl3_w_n3233_1(.douta(w_n3233_1[0]),.doutb(w_n3233_1[1]),.doutc(w_n3233_1[2]),.din(w_n3233_0[0]));
	jspl3 jspl3_w_n3233_2(.douta(w_n3233_2[0]),.doutb(w_n3233_2[1]),.doutc(w_n3233_2[2]),.din(w_n3233_0[1]));
	jspl3 jspl3_w_n3233_3(.douta(w_n3233_3[0]),.doutb(w_n3233_3[1]),.doutc(w_n3233_3[2]),.din(w_n3233_0[2]));
	jspl3 jspl3_w_n3233_4(.douta(w_n3233_4[0]),.doutb(w_n3233_4[1]),.doutc(w_n3233_4[2]),.din(w_n3233_1[0]));
	jspl3 jspl3_w_n3233_5(.douta(w_n3233_5[0]),.doutb(w_n3233_5[1]),.doutc(w_n3233_5[2]),.din(w_n3233_1[1]));
	jspl3 jspl3_w_n3233_6(.douta(w_n3233_6[0]),.doutb(w_n3233_6[1]),.doutc(w_n3233_6[2]),.din(w_n3233_1[2]));
	jspl3 jspl3_w_n3233_7(.douta(w_n3233_7[0]),.doutb(w_n3233_7[1]),.doutc(w_n3233_7[2]),.din(w_n3233_2[0]));
	jspl3 jspl3_w_n3233_8(.douta(w_n3233_8[0]),.doutb(w_n3233_8[1]),.doutc(w_n3233_8[2]),.din(w_n3233_2[1]));
	jspl3 jspl3_w_n3233_9(.douta(w_n3233_9[0]),.doutb(w_n3233_9[1]),.doutc(w_n3233_9[2]),.din(w_n3233_2[2]));
	jspl jspl_w_n3235_0(.douta(w_n3235_0[0]),.doutb(w_n3235_0[1]),.din(n3235));
	jspl jspl_w_n3236_0(.douta(w_n3236_0[0]),.doutb(w_n3236_0[1]),.din(n3236));
	jspl3 jspl3_w_n3237_0(.douta(w_n3237_0[0]),.doutb(w_n3237_0[1]),.doutc(w_n3237_0[2]),.din(n3237));
	jspl3 jspl3_w_n3237_1(.douta(w_n3237_1[0]),.doutb(w_n3237_1[1]),.doutc(w_n3237_1[2]),.din(w_n3237_0[0]));
	jspl jspl_w_n3237_2(.douta(w_n3237_2[0]),.doutb(w_n3237_2[1]),.din(w_n3237_0[1]));
	jspl3 jspl3_w_n3238_0(.douta(w_n3238_0[0]),.doutb(w_n3238_0[1]),.doutc(w_n3238_0[2]),.din(n3238));
	jspl3 jspl3_w_n3238_1(.douta(w_n3238_1[0]),.doutb(w_n3238_1[1]),.doutc(w_n3238_1[2]),.din(w_n3238_0[0]));
	jspl3 jspl3_w_n3238_2(.douta(w_n3238_2[0]),.doutb(w_n3238_2[1]),.doutc(w_n3238_2[2]),.din(w_n3238_0[1]));
	jspl3 jspl3_w_n3238_3(.douta(w_n3238_3[0]),.doutb(w_n3238_3[1]),.doutc(w_n3238_3[2]),.din(w_n3238_0[2]));
	jspl3 jspl3_w_n3238_4(.douta(w_n3238_4[0]),.doutb(w_n3238_4[1]),.doutc(w_n3238_4[2]),.din(w_n3238_1[0]));
	jspl3 jspl3_w_n3238_5(.douta(w_n3238_5[0]),.doutb(w_n3238_5[1]),.doutc(w_n3238_5[2]),.din(w_n3238_1[1]));
	jspl3 jspl3_w_n3238_6(.douta(w_n3238_6[0]),.doutb(w_n3238_6[1]),.doutc(w_n3238_6[2]),.din(w_n3238_1[2]));
	jspl jspl_w_n3238_7(.douta(w_n3238_7[0]),.doutb(w_n3238_7[1]),.din(w_n3238_2[0]));
	jspl jspl_w_n3240_0(.douta(w_n3240_0[0]),.doutb(w_n3240_0[1]),.din(n3240));
	jspl3 jspl3_w_n3242_0(.douta(w_n3242_0[0]),.doutb(w_n3242_0[1]),.doutc(w_n3242_0[2]),.din(n3242));
	jspl jspl_w_n3250_0(.douta(w_n3250_0[0]),.doutb(w_n3250_0[1]),.din(n3250));
	jspl3 jspl3_w_n3256_0(.douta(w_n3256_0[0]),.doutb(w_n3256_0[1]),.doutc(w_n3256_0[2]),.din(n3256));
	jspl jspl_w_n3257_0(.douta(w_n3257_0[0]),.doutb(w_n3257_0[1]),.din(n3257));
	jspl3 jspl3_w_n3258_0(.douta(w_n3258_0[0]),.doutb(w_n3258_0[1]),.doutc(w_n3258_0[2]),.din(n3258));
	jspl3 jspl3_w_n3258_1(.douta(w_n3258_1[0]),.doutb(w_n3258_1[1]),.doutc(w_n3258_1[2]),.din(w_n3258_0[0]));
	jspl jspl_w_n3263_0(.douta(w_n3263_0[0]),.doutb(w_n3263_0[1]),.din(n3263));
	jspl3 jspl3_w_n3270_0(.douta(w_n3270_0[0]),.doutb(w_n3270_0[1]),.doutc(w_n3270_0[2]),.din(n3270));
	jspl jspl_w_n3271_0(.douta(w_n3271_0[0]),.doutb(w_n3271_0[1]),.din(n3271));
	jspl jspl_w_n3274_0(.douta(w_n3274_0[0]),.doutb(w_n3274_0[1]),.din(n3274));
	jspl3 jspl3_w_n3282_0(.douta(w_n3282_0[0]),.doutb(w_n3282_0[1]),.doutc(w_n3282_0[2]),.din(n3282));
	jspl3 jspl3_w_n3283_0(.douta(w_n3283_0[0]),.doutb(w_n3283_0[1]),.doutc(w_n3283_0[2]),.din(n3283));
	jspl3 jspl3_w_n3283_1(.douta(w_n3283_1[0]),.doutb(w_n3283_1[1]),.doutc(w_n3283_1[2]),.din(w_n3283_0[0]));
	jspl3 jspl3_w_n3283_2(.douta(w_n3283_2[0]),.doutb(w_n3283_2[1]),.doutc(w_n3283_2[2]),.din(w_n3283_0[1]));
	jspl3 jspl3_w_n3283_3(.douta(w_n3283_3[0]),.doutb(w_n3283_3[1]),.doutc(w_n3283_3[2]),.din(w_n3283_0[2]));
	jspl3 jspl3_w_n3283_4(.douta(w_n3283_4[0]),.doutb(w_n3283_4[1]),.doutc(w_n3283_4[2]),.din(w_n3283_1[0]));
	jspl3 jspl3_w_n3283_5(.douta(w_n3283_5[0]),.doutb(w_n3283_5[1]),.doutc(w_n3283_5[2]),.din(w_n3283_1[1]));
	jspl3 jspl3_w_n3283_6(.douta(w_n3283_6[0]),.doutb(w_n3283_6[1]),.doutc(w_n3283_6[2]),.din(w_n3283_1[2]));
	jspl3 jspl3_w_n3283_7(.douta(w_n3283_7[0]),.doutb(w_n3283_7[1]),.doutc(w_n3283_7[2]),.din(w_n3283_2[0]));
	jspl jspl_w_n3283_8(.douta(w_n3283_8[0]),.doutb(w_n3283_8[1]),.din(w_n3283_2[1]));
	jspl3 jspl3_w_n3284_0(.douta(w_n3284_0[0]),.doutb(w_n3284_0[1]),.doutc(w_n3284_0[2]),.din(n3284));
	jspl3 jspl3_w_n3284_1(.douta(w_n3284_1[0]),.doutb(w_n3284_1[1]),.doutc(w_n3284_1[2]),.din(w_n3284_0[0]));
	jspl3 jspl3_w_n3284_2(.douta(w_n3284_2[0]),.doutb(w_n3284_2[1]),.doutc(w_n3284_2[2]),.din(w_n3284_0[1]));
	jspl3 jspl3_w_n3284_3(.douta(w_n3284_3[0]),.doutb(w_n3284_3[1]),.doutc(w_n3284_3[2]),.din(w_n3284_0[2]));
	jspl3 jspl3_w_n3284_4(.douta(w_n3284_4[0]),.doutb(w_n3284_4[1]),.doutc(w_n3284_4[2]),.din(w_n3284_1[0]));
	jspl3 jspl3_w_n3284_5(.douta(w_n3284_5[0]),.doutb(w_n3284_5[1]),.doutc(w_n3284_5[2]),.din(w_n3284_1[1]));
	jspl3 jspl3_w_n3284_6(.douta(w_n3284_6[0]),.doutb(w_n3284_6[1]),.doutc(w_n3284_6[2]),.din(w_n3284_1[2]));
	jspl3 jspl3_w_n3284_7(.douta(w_n3284_7[0]),.doutb(w_n3284_7[1]),.doutc(w_n3284_7[2]),.din(w_n3284_2[0]));
	jspl3 jspl3_w_n3284_8(.douta(w_n3284_8[0]),.doutb(w_n3284_8[1]),.doutc(w_n3284_8[2]),.din(w_n3284_2[1]));
	jspl jspl_w_n3285_0(.douta(w_n3285_0[0]),.doutb(w_n3285_0[1]),.din(n3285));
	jspl jspl_w_n3287_0(.douta(w_n3287_0[0]),.doutb(w_n3287_0[1]),.din(n3287));
	jspl jspl_w_n3291_0(.douta(w_n3291_0[0]),.doutb(w_n3291_0[1]),.din(n3291));
	jspl jspl_w_n3294_0(.douta(w_n3294_0[0]),.doutb(w_n3294_0[1]),.din(n3294));
	jspl jspl_w_n3296_0(.douta(w_n3296_0[0]),.doutb(w_n3296_0[1]),.din(n3296));
	jspl3 jspl3_w_n3299_0(.douta(w_n3299_0[0]),.doutb(w_n3299_0[1]),.doutc(w_n3299_0[2]),.din(n3299));
	jspl jspl_w_n3301_0(.douta(w_n3301_0[0]),.doutb(w_n3301_0[1]),.din(n3301));
	jspl3 jspl3_w_n3302_0(.douta(w_n3302_0[0]),.doutb(w_n3302_0[1]),.doutc(w_n3302_0[2]),.din(n3302));
	jspl jspl_w_n3303_0(.douta(w_n3303_0[0]),.doutb(w_n3303_0[1]),.din(n3303));
	jspl3 jspl3_w_n3307_0(.douta(w_n3307_0[0]),.doutb(w_n3307_0[1]),.doutc(w_n3307_0[2]),.din(n3307));
	jspl3 jspl3_w_n3307_1(.douta(w_n3307_1[0]),.doutb(w_n3307_1[1]),.doutc(w_n3307_1[2]),.din(w_n3307_0[0]));
	jspl3 jspl3_w_n3314_0(.douta(w_n3314_0[0]),.doutb(w_n3314_0[1]),.doutc(w_n3314_0[2]),.din(n3314));
	jspl3 jspl3_w_n3315_0(.douta(w_n3315_0[0]),.doutb(w_n3315_0[1]),.doutc(w_n3315_0[2]),.din(n3315));
	jspl3 jspl3_w_n3315_1(.douta(w_n3315_1[0]),.doutb(w_n3315_1[1]),.doutc(w_n3315_1[2]),.din(w_n3315_0[0]));
	jspl3 jspl3_w_n3315_2(.douta(w_n3315_2[0]),.doutb(w_n3315_2[1]),.doutc(w_n3315_2[2]),.din(w_n3315_0[1]));
	jspl3 jspl3_w_n3315_3(.douta(w_n3315_3[0]),.doutb(w_n3315_3[1]),.doutc(w_n3315_3[2]),.din(w_n3315_0[2]));
	jspl3 jspl3_w_n3315_4(.douta(w_n3315_4[0]),.doutb(w_n3315_4[1]),.doutc(w_n3315_4[2]),.din(w_n3315_1[0]));
	jspl3 jspl3_w_n3315_5(.douta(w_n3315_5[0]),.doutb(w_n3315_5[1]),.doutc(w_n3315_5[2]),.din(w_n3315_1[1]));
	jspl3 jspl3_w_n3315_6(.douta(w_n3315_6[0]),.doutb(w_n3315_6[1]),.doutc(w_n3315_6[2]),.din(w_n3315_1[2]));
	jspl3 jspl3_w_n3315_7(.douta(w_n3315_7[0]),.doutb(w_n3315_7[1]),.doutc(w_n3315_7[2]),.din(w_n3315_2[0]));
	jspl3 jspl3_w_n3316_0(.douta(w_n3316_0[0]),.doutb(w_n3316_0[1]),.doutc(w_n3316_0[2]),.din(n3316));
	jspl jspl_w_n3317_0(.douta(w_n3317_0[0]),.doutb(w_n3317_0[1]),.din(n3317));
	jspl jspl_w_n3319_0(.douta(w_n3319_0[0]),.doutb(w_n3319_0[1]),.din(n3319));
	jspl3 jspl3_w_n3320_0(.douta(w_n3320_0[0]),.doutb(w_n3320_0[1]),.doutc(w_n3320_0[2]),.din(n3320));
	jspl3 jspl3_w_n3320_1(.douta(w_n3320_1[0]),.doutb(w_n3320_1[1]),.doutc(w_n3320_1[2]),.din(w_n3320_0[0]));
	jspl3 jspl3_w_n3322_0(.douta(w_n3322_0[0]),.doutb(w_n3322_0[1]),.doutc(w_n3322_0[2]),.din(n3322));
	jspl3 jspl3_w_n3322_1(.douta(w_n3322_1[0]),.doutb(w_n3322_1[1]),.doutc(w_n3322_1[2]),.din(w_n3322_0[0]));
	jspl3 jspl3_w_n3322_2(.douta(w_n3322_2[0]),.doutb(w_n3322_2[1]),.doutc(w_n3322_2[2]),.din(w_n3322_0[1]));
	jspl3 jspl3_w_n3322_3(.douta(w_n3322_3[0]),.doutb(w_n3322_3[1]),.doutc(w_n3322_3[2]),.din(w_n3322_0[2]));
	jspl3 jspl3_w_n3322_4(.douta(w_n3322_4[0]),.doutb(w_n3322_4[1]),.doutc(w_n3322_4[2]),.din(w_n3322_1[0]));
	jspl3 jspl3_w_n3322_5(.douta(w_n3322_5[0]),.doutb(w_n3322_5[1]),.doutc(w_n3322_5[2]),.din(w_n3322_1[1]));
	jspl3 jspl3_w_n3322_6(.douta(w_n3322_6[0]),.doutb(w_n3322_6[1]),.doutc(w_n3322_6[2]),.din(w_n3322_1[2]));
	jspl jspl_w_n3322_7(.douta(w_n3322_7[0]),.doutb(w_n3322_7[1]),.din(w_n3322_2[0]));
	jspl3 jspl3_w_n3324_0(.douta(w_n3324_0[0]),.doutb(w_n3324_0[1]),.doutc(w_n3324_0[2]),.din(n3324));
	jspl3 jspl3_w_n3324_1(.douta(w_n3324_1[0]),.doutb(w_n3324_1[1]),.doutc(w_n3324_1[2]),.din(w_n3324_0[0]));
	jspl jspl_w_n3324_2(.douta(w_n3324_2[0]),.doutb(w_n3324_2[1]),.din(w_n3324_0[1]));
	jspl3 jspl3_w_n3325_0(.douta(w_n3325_0[0]),.doutb(w_n3325_0[1]),.doutc(w_n3325_0[2]),.din(n3325));
	jspl3 jspl3_w_n3325_1(.douta(w_n3325_1[0]),.doutb(w_n3325_1[1]),.doutc(w_n3325_1[2]),.din(w_n3325_0[0]));
	jspl3 jspl3_w_n3325_2(.douta(w_n3325_2[0]),.doutb(w_n3325_2[1]),.doutc(w_n3325_2[2]),.din(w_n3325_0[1]));
	jspl3 jspl3_w_n3325_3(.douta(w_n3325_3[0]),.doutb(w_n3325_3[1]),.doutc(w_n3325_3[2]),.din(w_n3325_0[2]));
	jspl3 jspl3_w_n3325_4(.douta(w_n3325_4[0]),.doutb(w_n3325_4[1]),.doutc(w_n3325_4[2]),.din(w_n3325_1[0]));
	jspl jspl_w_n3325_5(.douta(w_n3325_5[0]),.doutb(w_n3325_5[1]),.din(w_n3325_1[1]));
	jspl3 jspl3_w_n3328_0(.douta(w_n3328_0[0]),.doutb(w_n3328_0[1]),.doutc(w_n3328_0[2]),.din(n3328));
	jspl3 jspl3_w_n3328_1(.douta(w_n3328_1[0]),.doutb(w_n3328_1[1]),.doutc(w_n3328_1[2]),.din(w_n3328_0[0]));
	jspl3 jspl3_w_n3328_2(.douta(w_n3328_2[0]),.doutb(w_n3328_2[1]),.doutc(w_n3328_2[2]),.din(w_n3328_0[1]));
	jspl3 jspl3_w_n3328_3(.douta(w_n3328_3[0]),.doutb(w_n3328_3[1]),.doutc(w_n3328_3[2]),.din(w_n3328_0[2]));
	jspl3 jspl3_w_n3328_4(.douta(w_n3328_4[0]),.doutb(w_n3328_4[1]),.doutc(w_n3328_4[2]),.din(w_n3328_1[0]));
	jspl3 jspl3_w_n3328_5(.douta(w_n3328_5[0]),.doutb(w_n3328_5[1]),.doutc(w_n3328_5[2]),.din(w_n3328_1[1]));
	jspl jspl_w_n3333_0(.douta(w_n3333_0[0]),.doutb(w_n3333_0[1]),.din(n3333));
	jspl jspl_w_n3335_0(.douta(w_n3335_0[0]),.doutb(w_n3335_0[1]),.din(n3335));
	jspl3 jspl3_w_n3337_0(.douta(w_n3337_0[0]),.doutb(w_n3337_0[1]),.doutc(w_n3337_0[2]),.din(n3337));
	jspl3 jspl3_w_n3337_1(.douta(w_n3337_1[0]),.doutb(w_n3337_1[1]),.doutc(w_n3337_1[2]),.din(w_n3337_0[0]));
	jspl jspl_w_n3345_0(.douta(w_n3345_0[0]),.doutb(w_n3345_0[1]),.din(n3345));
	jspl jspl_w_n3347_0(.douta(w_n3347_0[0]),.doutb(w_n3347_0[1]),.din(n3347));
	jspl3 jspl3_w_n3348_0(.douta(w_n3348_0[0]),.doutb(w_n3348_0[1]),.doutc(w_n3348_0[2]),.din(n3348));
	jspl3 jspl3_w_n3349_0(.douta(w_n3349_0[0]),.doutb(w_n3349_0[1]),.doutc(w_n3349_0[2]),.din(n3349));
	jspl3 jspl3_w_n3350_0(.douta(w_n3350_0[0]),.doutb(w_n3350_0[1]),.doutc(w_n3350_0[2]),.din(n3350));
	jspl3 jspl3_w_n3351_0(.douta(w_n3351_0[0]),.doutb(w_n3351_0[1]),.doutc(w_n3351_0[2]),.din(n3351));
	jspl3 jspl3_w_n3352_0(.douta(w_n3352_0[0]),.doutb(w_n3352_0[1]),.doutc(w_n3352_0[2]),.din(n3352));
	jspl3 jspl3_w_n3353_0(.douta(w_n3353_0[0]),.doutb(w_n3353_0[1]),.doutc(w_n3353_0[2]),.din(n3353));
	jspl3 jspl3_w_n3354_0(.douta(w_n3354_0[0]),.doutb(w_n3354_0[1]),.doutc(w_n3354_0[2]),.din(n3354));
	jspl3 jspl3_w_n3362_0(.douta(w_n3362_0[0]),.doutb(w_n3362_0[1]),.doutc(w_n3362_0[2]),.din(n3362));
	jspl3 jspl3_w_n3365_0(.douta(w_n3365_0[0]),.doutb(w_n3365_0[1]),.doutc(w_n3365_0[2]),.din(n3365));
	jspl3 jspl3_w_n3367_0(.douta(w_n3367_0[0]),.doutb(w_n3367_0[1]),.doutc(w_n3367_0[2]),.din(n3367));
	jspl jspl_w_n3373_0(.douta(w_n3373_0[0]),.doutb(w_n3373_0[1]),.din(n3373));
	jspl jspl_w_n3375_0(.douta(w_n3375_0[0]),.doutb(w_n3375_0[1]),.din(n3375));
	jspl jspl_w_n3379_0(.douta(w_n3379_0[0]),.doutb(w_n3379_0[1]),.din(n3379));
	jspl jspl_w_n3394_0(.douta(w_n3394_0[0]),.doutb(w_n3394_0[1]),.din(n3394));
	jspl jspl_w_n3396_0(.douta(w_n3396_0[0]),.doutb(w_n3396_0[1]),.din(n3396));
	jspl jspl_w_n3397_0(.douta(w_n3397_0[0]),.doutb(w_n3397_0[1]),.din(n3397));
	jspl jspl_w_n3406_0(.douta(w_n3406_0[0]),.doutb(w_n3406_0[1]),.din(n3406));
	jspl jspl_w_n3408_0(.douta(w_n3408_0[0]),.doutb(w_n3408_0[1]),.din(n3408));
	jspl jspl_w_n3409_0(.douta(w_n3409_0[0]),.doutb(w_n3409_0[1]),.din(n3409));
	jspl jspl_w_n3418_0(.douta(w_n3418_0[0]),.doutb(w_n3418_0[1]),.din(n3418));
	jspl jspl_w_n3420_0(.douta(w_n3420_0[0]),.doutb(w_n3420_0[1]),.din(n3420));
	jspl jspl_w_n3421_0(.douta(w_n3421_0[0]),.doutb(w_n3421_0[1]),.din(n3421));
	jspl jspl_w_n3423_0(.douta(w_n3423_0[0]),.doutb(w_n3423_0[1]),.din(n3423));
	jspl jspl_w_n3425_0(.douta(w_n3425_0[0]),.doutb(w_n3425_0[1]),.din(n3425));
	jspl jspl_w_n3426_0(.douta(w_n3426_0[0]),.doutb(w_n3426_0[1]),.din(n3426));
	jspl jspl_w_n3435_0(.douta(w_n3435_0[0]),.doutb(w_n3435_0[1]),.din(n3435));
	jspl jspl_w_n3437_0(.douta(w_n3437_0[0]),.doutb(w_n3437_0[1]),.din(n3437));
	jspl jspl_w_n3438_0(.douta(w_n3438_0[0]),.doutb(w_n3438_0[1]),.din(n3438));
	jspl jspl_w_n3446_0(.douta(w_n3446_0[0]),.doutb(w_n3446_0[1]),.din(n3446));
	jspl jspl_w_n3452_0(.douta(w_n3452_0[0]),.doutb(w_n3452_0[1]),.din(n3452));
	jspl jspl_w_n3454_0(.douta(w_n3454_0[0]),.doutb(w_n3454_0[1]),.din(n3454));
	jspl jspl_w_n3455_0(.douta(w_n3455_0[0]),.doutb(w_n3455_0[1]),.din(n3455));
	jspl jspl_w_n3464_0(.douta(w_n3464_0[0]),.doutb(w_n3464_0[1]),.din(n3464));
	jspl jspl_w_n3466_0(.douta(w_n3466_0[0]),.doutb(w_n3466_0[1]),.din(n3466));
	jspl jspl_w_n3467_0(.douta(w_n3467_0[0]),.doutb(w_n3467_0[1]),.din(n3467));
	jspl jspl_w_n3475_0(.douta(w_n3475_0[0]),.doutb(w_n3475_0[1]),.din(n3475));
	jspl jspl_w_n3482_0(.douta(w_n3482_0[0]),.doutb(w_n3482_0[1]),.din(n3482));
	jspl jspl_w_n3484_0(.douta(w_n3484_0[0]),.doutb(w_n3484_0[1]),.din(n3484));
	jspl jspl_w_n3485_0(.douta(w_n3485_0[0]),.doutb(w_n3485_0[1]),.din(n3485));
	jspl jspl_w_n3494_0(.douta(w_n3494_0[0]),.doutb(w_n3494_0[1]),.din(n3494));
	jspl jspl_w_n3496_0(.douta(w_n3496_0[0]),.doutb(w_n3496_0[1]),.din(n3496));
	jspl jspl_w_n3497_0(.douta(w_n3497_0[0]),.doutb(w_n3497_0[1]),.din(n3497));
	jspl jspl_w_n3504_0(.douta(w_n3504_0[0]),.doutb(w_n3504_0[1]),.din(n3504));
	jspl jspl_w_n3510_0(.douta(w_n3510_0[0]),.doutb(w_n3510_0[1]),.din(n3510));
	jspl jspl_w_n3512_0(.douta(w_n3512_0[0]),.doutb(w_n3512_0[1]),.din(n3512));
	jspl jspl_w_n3513_0(.douta(w_n3513_0[0]),.doutb(w_n3513_0[1]),.din(n3513));
	jspl3 jspl3_w_n3516_0(.douta(w_n3516_0[0]),.doutb(w_n3516_0[1]),.doutc(w_n3516_0[2]),.din(n3516));
	jspl3 jspl3_w_n3516_1(.douta(w_n3516_1[0]),.doutb(w_n3516_1[1]),.doutc(w_n3516_1[2]),.din(w_n3516_0[0]));
	jspl jspl_w_n3524_0(.douta(w_n3524_0[0]),.doutb(w_n3524_0[1]),.din(n3524));
	jspl jspl_w_n3528_0(.douta(w_n3528_0[0]),.doutb(w_n3528_0[1]),.din(n3528));
	jspl jspl_w_n3529_0(.douta(w_n3529_0[0]),.doutb(w_n3529_0[1]),.din(n3529));
	jspl jspl_w_n3530_0(.douta(w_n3530_0[0]),.doutb(w_n3530_0[1]),.din(n3530));
	jspl jspl_w_n3532_0(.douta(w_n3532_0[0]),.doutb(w_n3532_0[1]),.din(n3532));
	jspl jspl_w_n3535_0(.douta(w_n3535_0[0]),.doutb(w_n3535_0[1]),.din(n3535));
	jspl jspl_w_n3543_0(.douta(w_n3543_0[0]),.doutb(w_n3543_0[1]),.din(n3543));
	jspl jspl_w_n3546_0(.douta(w_n3546_0[0]),.doutb(w_n3546_0[1]),.din(n3546));
	jspl jspl_w_n3554_0(.douta(w_n3554_0[0]),.doutb(w_n3554_0[1]),.din(n3554));
	jspl jspl_w_n3557_0(.douta(w_n3557_0[0]),.doutb(w_n3557_0[1]),.din(n3557));
	jspl jspl_w_n3565_0(.douta(w_n3565_0[0]),.doutb(w_n3565_0[1]),.din(n3565));
	jspl jspl_w_n3567_0(.douta(w_n3567_0[0]),.doutb(w_n3567_0[1]),.din(n3567));
	jspl3 jspl3_w_n3571_0(.douta(w_n3571_0[0]),.doutb(w_n3571_0[1]),.doutc(w_n3571_0[2]),.din(n3571));
	jspl jspl_w_n3571_1(.douta(w_n3571_1[0]),.doutb(w_n3571_1[1]),.din(w_n3571_0[0]));
	jspl3 jspl3_w_n3573_0(.douta(w_n3573_0[0]),.doutb(w_n3573_0[1]),.doutc(w_n3573_0[2]),.din(n3573));
	jspl jspl_w_n3579_0(.douta(w_n3579_0[0]),.doutb(w_n3579_0[1]),.din(n3579));
	jspl jspl_w_n3580_0(.douta(w_n3580_0[0]),.doutb(w_n3580_0[1]),.din(n3580));
	jspl jspl_w_n3581_0(.douta(w_n3581_0[0]),.doutb(w_n3581_0[1]),.din(n3581));
	jspl jspl_w_n3582_0(.douta(w_n3582_0[0]),.doutb(w_n3582_0[1]),.din(n3582));
	jspl jspl_w_n3583_0(.douta(w_n3583_0[0]),.doutb(w_n3583_0[1]),.din(n3583));
	jspl jspl_w_n3584_0(.douta(w_n3584_0[0]),.doutb(w_n3584_0[1]),.din(n3584));
	jspl jspl_w_n3585_0(.douta(w_n3585_0[0]),.doutb(w_n3585_0[1]),.din(n3585));
	jspl jspl_w_n3586_0(.douta(w_n3586_0[0]),.doutb(w_n3586_0[1]),.din(n3586));
	jspl jspl_w_n3587_0(.douta(w_n3587_0[0]),.doutb(w_n3587_0[1]),.din(n3587));
	jspl jspl_w_n3590_0(.douta(w_n3590_0[0]),.doutb(w_n3590_0[1]),.din(n3590));
	jspl jspl_w_n3591_0(.douta(w_n3591_0[0]),.doutb(w_n3591_0[1]),.din(n3591));
	jspl jspl_w_n3592_0(.douta(w_n3592_0[0]),.doutb(w_n3592_0[1]),.din(n3592));
	jspl3 jspl3_w_n3599_0(.douta(w_n3599_0[0]),.doutb(w_n3599_0[1]),.doutc(w_n3599_0[2]),.din(n3599));
	jspl3 jspl3_w_n3600_0(.douta(w_n3600_0[0]),.doutb(w_n3600_0[1]),.doutc(w_n3600_0[2]),.din(n3600));
	jspl3 jspl3_w_n3600_1(.douta(w_n3600_1[0]),.doutb(w_n3600_1[1]),.doutc(w_n3600_1[2]),.din(w_n3600_0[0]));
	jspl3 jspl3_w_n3600_2(.douta(w_n3600_2[0]),.doutb(w_n3600_2[1]),.doutc(w_n3600_2[2]),.din(w_n3600_0[1]));
	jspl3 jspl3_w_n3600_3(.douta(w_n3600_3[0]),.doutb(w_n3600_3[1]),.doutc(w_n3600_3[2]),.din(w_n3600_0[2]));
	jspl3 jspl3_w_n3600_4(.douta(w_n3600_4[0]),.doutb(w_n3600_4[1]),.doutc(w_n3600_4[2]),.din(w_n3600_1[0]));
	jspl3 jspl3_w_n3600_5(.douta(w_n3600_5[0]),.doutb(w_n3600_5[1]),.doutc(w_n3600_5[2]),.din(w_n3600_1[1]));
	jspl3 jspl3_w_n3600_6(.douta(w_n3600_6[0]),.doutb(w_n3600_6[1]),.doutc(w_n3600_6[2]),.din(w_n3600_1[2]));
	jspl3 jspl3_w_n3600_7(.douta(w_n3600_7[0]),.doutb(w_n3600_7[1]),.doutc(w_n3600_7[2]),.din(w_n3600_2[0]));
	jspl3 jspl3_w_n3600_8(.douta(w_n3600_8[0]),.doutb(w_n3600_8[1]),.doutc(w_n3600_8[2]),.din(w_n3600_2[1]));
	jspl3 jspl3_w_n3601_0(.douta(w_n3601_0[0]),.doutb(w_n3601_0[1]),.doutc(w_n3601_0[2]),.din(n3601));
	jspl jspl_w_n3601_1(.douta(w_n3601_1[0]),.doutb(w_n3601_1[1]),.din(w_n3601_0[0]));
	jspl jspl_w_n3602_0(.douta(w_n3602_0[0]),.doutb(w_n3602_0[1]),.din(n3602));
	jspl jspl_w_n3604_0(.douta(w_n3604_0[0]),.doutb(w_n3604_0[1]),.din(n3604));
	jspl3 jspl3_w_n3605_0(.douta(w_n3605_0[0]),.doutb(w_n3605_0[1]),.doutc(w_n3605_0[2]),.din(n3605));
	jspl3 jspl3_w_n3605_1(.douta(w_n3605_1[0]),.doutb(w_n3605_1[1]),.doutc(w_n3605_1[2]),.din(w_n3605_0[0]));
	jspl jspl_w_n3613_0(.douta(w_n3613_0[0]),.doutb(w_n3613_0[1]),.din(n3613));
	jspl jspl_w_n3614_0(.douta(w_n3614_0[0]),.doutb(w_n3614_0[1]),.din(n3614));
	jspl jspl_w_n3615_0(.douta(w_n3615_0[0]),.doutb(w_n3615_0[1]),.din(n3615));
	jspl jspl_w_n3620_0(.douta(w_n3620_0[0]),.doutb(w_n3620_0[1]),.din(n3620));
	jspl3 jspl3_w_n3624_0(.douta(w_n3624_0[0]),.doutb(w_n3624_0[1]),.doutc(w_n3624_0[2]),.din(n3624));
	jspl jspl_w_n3626_0(.douta(w_n3626_0[0]),.doutb(w_n3626_0[1]),.din(n3626));
	jspl jspl_w_n3630_0(.douta(w_n3630_0[0]),.doutb(w_n3630_0[1]),.din(n3630));
	jspl jspl_w_n3633_0(.douta(w_n3633_0[0]),.doutb(w_n3633_0[1]),.din(n3633));
	jspl jspl_w_n3634_0(.douta(w_n3634_0[0]),.doutb(w_n3634_0[1]),.din(n3634));
	jspl jspl_w_n3638_0(.douta(w_n3638_0[0]),.doutb(w_n3638_0[1]),.din(n3638));
	jspl jspl_w_n3650_0(.douta(w_n3650_0[0]),.doutb(w_n3650_0[1]),.din(n3650));
	jspl jspl_w_n3652_0(.douta(w_n3652_0[0]),.doutb(w_n3652_0[1]),.din(n3652));
	jspl jspl_w_n3654_0(.douta(w_n3654_0[0]),.doutb(w_n3654_0[1]),.din(n3654));
	jspl jspl_w_n3663_0(.douta(w_n3663_0[0]),.doutb(w_n3663_0[1]),.din(n3663));
	jspl jspl_w_n3666_0(.douta(w_n3666_0[0]),.doutb(w_n3666_0[1]),.din(n3666));
	jspl jspl_w_n3669_0(.douta(w_n3669_0[0]),.doutb(w_n3669_0[1]),.din(n3669));
	jspl jspl_w_n3676_0(.douta(w_n3676_0[0]),.doutb(w_n3676_0[1]),.din(n3676));
	jspl jspl_w_n3686_0(.douta(w_n3686_0[0]),.doutb(w_n3686_0[1]),.din(n3686));
	jspl3 jspl3_w_n3693_0(.douta(w_n3693_0[0]),.doutb(w_n3693_0[1]),.doutc(w_n3693_0[2]),.din(n3693));
	jspl jspl_w_n3696_0(.douta(w_n3696_0[0]),.doutb(w_n3696_0[1]),.din(n3696));
	jspl jspl_w_n3779_0(.douta(w_n3779_0[0]),.doutb(w_n3779_0[1]),.din(n3779));
	jspl jspl_w_n3781_0(.douta(w_n3781_0[0]),.doutb(w_n3781_0[1]),.din(n3781));
	jspl jspl_w_n3784_0(.douta(w_n3784_0[0]),.doutb(w_n3784_0[1]),.din(n3784));
	jspl jspl_w_n3787_0(.douta(w_n3787_0[0]),.doutb(w_n3787_0[1]),.din(n3787));
	jspl jspl_w_n3794_0(.douta(w_n3794_0[0]),.doutb(w_n3794_0[1]),.din(n3794));
	jspl jspl_w_n3805_0(.douta(w_n3805_0[0]),.doutb(w_n3805_0[1]),.din(n3805));
	jspl3 jspl3_w_n3806_0(.douta(w_n3806_0[0]),.doutb(w_n3806_0[1]),.doutc(w_n3806_0[2]),.din(n3806));
	jspl3 jspl3_w_n3806_1(.douta(w_n3806_1[0]),.doutb(w_n3806_1[1]),.doutc(w_n3806_1[2]),.din(w_n3806_0[0]));
	jspl3 jspl3_w_n3806_2(.douta(w_n3806_2[0]),.doutb(w_n3806_2[1]),.doutc(w_n3806_2[2]),.din(w_n3806_0[1]));
	jspl3 jspl3_w_n3806_3(.douta(w_n3806_3[0]),.doutb(w_n3806_3[1]),.doutc(w_n3806_3[2]),.din(w_n3806_0[2]));
	jspl3 jspl3_w_n3806_4(.douta(w_n3806_4[0]),.doutb(w_n3806_4[1]),.doutc(w_n3806_4[2]),.din(w_n3806_1[0]));
	jspl3 jspl3_w_n3806_5(.douta(w_n3806_5[0]),.doutb(w_n3806_5[1]),.doutc(w_n3806_5[2]),.din(w_n3806_1[1]));
	jspl3 jspl3_w_n3807_0(.douta(w_n3807_0[0]),.doutb(w_n3807_0[1]),.doutc(w_n3807_0[2]),.din(n3807));
	jspl3 jspl3_w_n3807_1(.douta(w_n3807_1[0]),.doutb(w_n3807_1[1]),.doutc(w_n3807_1[2]),.din(w_n3807_0[0]));
	jspl3 jspl3_w_n3807_2(.douta(w_n3807_2[0]),.doutb(w_n3807_2[1]),.doutc(w_n3807_2[2]),.din(w_n3807_0[1]));
	jspl jspl_w_n3807_3(.douta(w_n3807_3[0]),.doutb(w_n3807_3[1]),.din(w_n3807_0[2]));
	jspl jspl_w_n3808_0(.douta(w_n3808_0[0]),.doutb(w_n3808_0[1]),.din(n3808));
	jspl jspl_w_n3810_0(.douta(w_n3810_0[0]),.doutb(w_n3810_0[1]),.din(n3810));
	jspl3 jspl3_w_n3811_0(.douta(w_n3811_0[0]),.doutb(w_n3811_0[1]),.doutc(w_n3811_0[2]),.din(n3811));
	jspl3 jspl3_w_n3811_1(.douta(w_n3811_1[0]),.doutb(w_n3811_1[1]),.doutc(w_n3811_1[2]),.din(w_n3811_0[0]));
	jspl jspl_w_n3820_0(.douta(w_n3820_0[0]),.doutb(w_n3820_0[1]),.din(n3820));
	jspl jspl_w_n3823_0(.douta(w_n3823_0[0]),.doutb(w_n3823_0[1]),.din(n3823));
	jspl jspl_w_n3826_0(.douta(w_n3826_0[0]),.doutb(w_n3826_0[1]),.din(n3826));
	jspl jspl_w_n3835_0(.douta(w_n3835_0[0]),.doutb(w_n3835_0[1]),.din(n3835));
	jspl jspl_w_n3838_0(.douta(w_n3838_0[0]),.doutb(w_n3838_0[1]),.din(n3838));
	jspl jspl_w_n3848_0(.douta(w_n3848_0[0]),.doutb(w_n3848_0[1]),.din(n3848));
	jspl jspl_w_n3849_0(.douta(w_n3849_0[0]),.doutb(w_n3849_0[1]),.din(n3849));
	jspl jspl_w_n3853_0(.douta(w_n3853_0[0]),.doutb(w_n3853_0[1]),.din(n3853));
	jspl jspl_w_n3854_0(.douta(w_n3854_0[0]),.doutb(w_n3854_0[1]),.din(n3854));
	jspl jspl_w_n3862_0(.douta(w_n3862_0[0]),.doutb(w_n3862_0[1]),.din(n3862));
	jspl jspl_w_n3863_0(.douta(w_n3863_0[0]),.doutb(w_n3863_0[1]),.din(n3863));
	jspl jspl_w_n3864_0(.douta(w_n3864_0[0]),.doutb(w_n3864_0[1]),.din(n3864));
	jspl jspl_w_n3865_0(.douta(w_n3865_0[0]),.doutb(w_n3865_0[1]),.din(n3865));
	jspl jspl_w_n3866_0(.douta(w_n3866_0[0]),.doutb(w_n3866_0[1]),.din(n3866));
	jspl jspl_w_n3874_0(.douta(w_n3874_0[0]),.doutb(w_n3874_0[1]),.din(n3874));
	jspl jspl_w_n3875_0(.douta(w_n3875_0[0]),.doutb(w_n3875_0[1]),.din(n3875));
	jspl jspl_w_n3876_0(.douta(w_n3876_0[0]),.doutb(w_n3876_0[1]),.din(n3876));
	jspl jspl_w_n3877_0(.douta(w_n3877_0[0]),.doutb(w_n3877_0[1]),.din(n3877));
	jspl jspl_w_n3878_0(.douta(w_n3878_0[0]),.doutb(w_n3878_0[1]),.din(n3878));
	jspl jspl_w_n3888_0(.douta(w_n3888_0[0]),.doutb(w_n3888_0[1]),.din(n3888));
	jspl jspl_w_n3889_0(.douta(w_n3889_0[0]),.doutb(w_n3889_0[1]),.din(n3889));
	jspl jspl_w_n3890_0(.douta(w_n3890_0[0]),.doutb(w_n3890_0[1]),.din(n3890));
	jspl jspl_w_n3891_0(.douta(w_n3891_0[0]),.doutb(w_n3891_0[1]),.din(n3891));
	jspl jspl_w_n3896_0(.douta(w_n3896_0[0]),.doutb(w_n3896_0[1]),.din(n3896));
	jspl jspl_w_n3899_0(.douta(w_n3899_0[0]),.doutb(w_n3899_0[1]),.din(n3899));
	jspl jspl_w_n3900_0(.douta(w_n3900_0[0]),.doutb(w_n3900_0[1]),.din(n3900));
	jspl jspl_w_n3902_0(.douta(w_n3902_0[0]),.doutb(w_n3902_0[1]),.din(n3902));
	jspl jspl_w_n3909_0(.douta(w_n3909_0[0]),.doutb(w_n3909_0[1]),.din(n3909));
	jspl jspl_w_n3911_0(.douta(w_n3911_0[0]),.doutb(w_n3911_0[1]),.din(n3911));
	jspl3 jspl3_w_n3919_0(.douta(w_n3919_0[0]),.doutb(w_n3919_0[1]),.doutc(w_n3919_0[2]),.din(n3919));
	jspl3 jspl3_w_n3919_1(.douta(w_n3919_1[0]),.doutb(w_n3919_1[1]),.doutc(w_n3919_1[2]),.din(w_n3919_0[0]));
	jspl3 jspl3_w_n3919_2(.douta(w_n3919_2[0]),.doutb(w_n3919_2[1]),.doutc(w_n3919_2[2]),.din(w_n3919_0[1]));
	jspl3 jspl3_w_n3919_3(.douta(w_n3919_3[0]),.doutb(w_n3919_3[1]),.doutc(w_n3919_3[2]),.din(w_n3919_0[2]));
	jspl3 jspl3_w_n3919_4(.douta(w_n3919_4[0]),.doutb(w_n3919_4[1]),.doutc(w_n3919_4[2]),.din(w_n3919_1[0]));
	jspl3 jspl3_w_n3919_5(.douta(w_n3919_5[0]),.doutb(w_n3919_5[1]),.doutc(w_n3919_5[2]),.din(w_n3919_1[1]));
	jspl3 jspl3_w_n3920_0(.douta(w_n3920_0[0]),.doutb(w_n3920_0[1]),.doutc(w_n3920_0[2]),.din(n3920));
	jspl3 jspl3_w_n3920_1(.douta(w_n3920_1[0]),.doutb(w_n3920_1[1]),.doutc(w_n3920_1[2]),.din(w_n3920_0[0]));
	jspl3 jspl3_w_n3920_2(.douta(w_n3920_2[0]),.doutb(w_n3920_2[1]),.doutc(w_n3920_2[2]),.din(w_n3920_0[1]));
	jspl jspl_w_n3920_3(.douta(w_n3920_3[0]),.doutb(w_n3920_3[1]),.din(w_n3920_0[2]));
	jspl jspl_w_n3924_0(.douta(w_n3924_0[0]),.doutb(w_n3924_0[1]),.din(n3924));
	jspl jspl_w_n3925_0(.douta(w_n3925_0[0]),.doutb(w_n3925_0[1]),.din(n3925));
	jspl3 jspl3_w_n3927_0(.douta(w_n3927_0[0]),.doutb(w_n3927_0[1]),.doutc(w_n3927_0[2]),.din(n3927));
	jspl3 jspl3_w_n3927_1(.douta(w_n3927_1[0]),.doutb(w_n3927_1[1]),.doutc(w_n3927_1[2]),.din(w_n3927_0[0]));
	jspl jspl_w_n3936_0(.douta(w_n3936_0[0]),.doutb(w_n3936_0[1]),.din(n3936));
	jspl jspl_w_n3939_0(.douta(w_n3939_0[0]),.doutb(w_n3939_0[1]),.din(n3939));
	jspl jspl_w_n3942_0(.douta(w_n3942_0[0]),.doutb(w_n3942_0[1]),.din(n3942));
	jspl jspl_w_n3951_0(.douta(w_n3951_0[0]),.doutb(w_n3951_0[1]),.din(n3951));
	jspl jspl_w_n3954_0(.douta(w_n3954_0[0]),.doutb(w_n3954_0[1]),.din(n3954));
	jspl jspl_w_n3962_0(.douta(w_n3962_0[0]),.doutb(w_n3962_0[1]),.din(n3962));
	jspl jspl_w_n3972_0(.douta(w_n3972_0[0]),.doutb(w_n3972_0[1]),.din(n3972));
	jspl jspl_w_n3973_0(.douta(w_n3973_0[0]),.doutb(w_n3973_0[1]),.din(n3973));
	jspl jspl_w_n3977_0(.douta(w_n3977_0[0]),.doutb(w_n3977_0[1]),.din(n3977));
	jspl jspl_w_n3978_0(.douta(w_n3978_0[0]),.doutb(w_n3978_0[1]),.din(n3978));
	jspl jspl_w_n3979_0(.douta(w_n3979_0[0]),.doutb(w_n3979_0[1]),.din(n3979));
	jspl jspl_w_n3980_0(.douta(w_n3980_0[0]),.doutb(w_n3980_0[1]),.din(n3980));
	jspl jspl_w_n3981_0(.douta(w_n3981_0[0]),.doutb(w_n3981_0[1]),.din(n3981));
	jspl jspl_w_n3982_0(.douta(w_n3982_0[0]),.doutb(w_n3982_0[1]),.din(n3982));
	jspl jspl_w_n3990_0(.douta(w_n3990_0[0]),.doutb(w_n3990_0[1]),.din(n3990));
	jspl jspl_w_n3991_0(.douta(w_n3991_0[0]),.doutb(w_n3991_0[1]),.din(n3991));
	jspl jspl_w_n3992_0(.douta(w_n3992_0[0]),.doutb(w_n3992_0[1]),.din(n3992));
	jspl jspl_w_n3993_0(.douta(w_n3993_0[0]),.doutb(w_n3993_0[1]),.din(n3993));
	jspl jspl_w_n3994_0(.douta(w_n3994_0[0]),.doutb(w_n3994_0[1]),.din(n3994));
	jspl3 jspl3_w_n4000_0(.douta(w_n4000_0[0]),.doutb(w_n4000_0[1]),.doutc(w_n4000_0[2]),.din(n4000));
	jspl jspl_w_n4009_0(.douta(w_n4009_0[0]),.doutb(w_n4009_0[1]),.din(n4009));
	jspl jspl_w_n4010_0(.douta(w_n4010_0[0]),.doutb(w_n4010_0[1]),.din(n4010));
	jspl3 jspl3_w_n4011_0(.douta(w_n4011_0[0]),.doutb(w_n4011_0[1]),.doutc(w_n4011_0[2]),.din(n4011));
	jspl3 jspl3_w_n4013_0(.douta(w_n4013_0[0]),.doutb(w_n4013_0[1]),.doutc(w_n4013_0[2]),.din(n4013));
	jspl3 jspl3_w_n4013_1(.douta(w_n4013_1[0]),.doutb(w_n4013_1[1]),.doutc(w_n4013_1[2]),.din(w_n4013_0[0]));
	jspl3 jspl3_w_n4013_2(.douta(w_dff_A_zFz06Ms96_0),.doutb(w_dff_A_bJB9Q22H3_1),.doutc(w_n4013_2[2]),.din(w_n4013_0[1]));
	jspl3 jspl3_w_n4013_3(.douta(w_n4013_3[0]),.doutb(w_dff_A_0eyV9lEz2_1),.doutc(w_dff_A_OxUIVHDa5_2),.din(w_n4013_0[2]));
	jspl3 jspl3_w_n4013_4(.douta(w_dff_A_b6PhEX3p8_0),.doutb(w_dff_A_QWOvLrxd2_1),.doutc(w_n4013_4[2]),.din(w_n4013_1[0]));
	jspl3 jspl3_w_n4013_5(.douta(w_n4013_5[0]),.doutb(w_n4013_5[1]),.doutc(w_n4013_5[2]),.din(w_n4013_1[1]));
	jspl3 jspl3_w_n4013_6(.douta(w_dff_A_wMefoSvl1_0),.doutb(w_dff_A_dBDyGrTJ0_1),.doutc(w_n4013_6[2]),.din(w_n4013_1[2]));
	jspl3 jspl3_w_n4013_7(.douta(w_dff_A_GJdM5i5M9_0),.doutb(w_dff_A_hKKpVgtY8_1),.doutc(w_n4013_7[2]),.din(w_n4013_2[0]));
	jspl3 jspl3_w_n4013_8(.douta(w_dff_A_VEC9hgaD8_0),.doutb(w_dff_A_TV7kAWfk8_1),.doutc(w_n4013_8[2]),.din(w_n4013_2[1]));
	jspl3 jspl3_w_n4013_9(.douta(w_dff_A_s4kVgoWW2_0),.doutb(w_dff_A_ucqtqfZU9_1),.doutc(w_n4013_9[2]),.din(w_n4013_2[2]));
	jspl3 jspl3_w_n4013_10(.douta(w_dff_A_kpphw58F3_0),.doutb(w_dff_A_Hx1Ouz7H2_1),.doutc(w_n4013_10[2]),.din(w_n4013_3[0]));
	jspl jspl_w_n4014_0(.douta(w_n4014_0[0]),.doutb(w_dff_A_RiPtSZDk9_1),.din(n4014));
	jspl jspl_w_n4017_0(.douta(w_n4017_0[0]),.doutb(w_n4017_0[1]),.din(n4017));
	jspl jspl_w_n4018_0(.douta(w_n4018_0[0]),.doutb(w_n4018_0[1]),.din(n4018));
	jspl jspl_w_n4021_0(.douta(w_n4021_0[0]),.doutb(w_n4021_0[1]),.din(n4021));
	jspl jspl_w_n4025_0(.douta(w_n4025_0[0]),.doutb(w_n4025_0[1]),.din(n4025));
	jspl jspl_w_n4028_0(.douta(w_n4028_0[0]),.doutb(w_n4028_0[1]),.din(n4028));
	jspl jspl_w_n4031_0(.douta(w_n4031_0[0]),.doutb(w_n4031_0[1]),.din(n4031));
	jspl jspl_w_n4034_0(.douta(w_n4034_0[0]),.doutb(w_n4034_0[1]),.din(n4034));
	jspl jspl_w_n4043_0(.douta(w_n4043_0[0]),.doutb(w_n4043_0[1]),.din(n4043));
	jspl jspl_w_n4046_0(.douta(w_n4046_0[0]),.doutb(w_n4046_0[1]),.din(n4046));
	jspl jspl_w_n4054_0(.douta(w_n4054_0[0]),.doutb(w_n4054_0[1]),.din(n4054));
	jspl jspl_w_n4064_0(.douta(w_n4064_0[0]),.doutb(w_n4064_0[1]),.din(n4064));
	jspl jspl_w_n4065_0(.douta(w_n4065_0[0]),.doutb(w_n4065_0[1]),.din(n4065));
	jspl jspl_w_n4069_0(.douta(w_n4069_0[0]),.doutb(w_n4069_0[1]),.din(n4069));
	jspl jspl_w_n4070_0(.douta(w_n4070_0[0]),.doutb(w_n4070_0[1]),.din(n4070));
	jspl jspl_w_n4071_0(.douta(w_n4071_0[0]),.doutb(w_n4071_0[1]),.din(n4071));
	jspl jspl_w_n4072_0(.douta(w_n4072_0[0]),.doutb(w_n4072_0[1]),.din(n4072));
	jspl jspl_w_n4073_0(.douta(w_n4073_0[0]),.doutb(w_n4073_0[1]),.din(n4073));
	jspl jspl_w_n4074_0(.douta(w_n4074_0[0]),.doutb(w_n4074_0[1]),.din(n4074));
	jspl jspl_w_n4082_0(.douta(w_n4082_0[0]),.doutb(w_n4082_0[1]),.din(n4082));
	jspl jspl_w_n4083_0(.douta(w_n4083_0[0]),.doutb(w_n4083_0[1]),.din(n4083));
	jspl jspl_w_n4084_0(.douta(w_n4084_0[0]),.doutb(w_n4084_0[1]),.din(n4084));
	jspl jspl_w_n4086_0(.douta(w_n4086_0[0]),.doutb(w_n4086_0[1]),.din(n4086));
	jspl jspl_w_n4088_0(.douta(w_n4088_0[0]),.doutb(w_n4088_0[1]),.din(n4088));
	jspl3 jspl3_w_n4090_0(.douta(w_n4090_0[0]),.doutb(w_n4090_0[1]),.doutc(w_n4090_0[2]),.din(n4090));
	jspl3 jspl3_w_n4090_1(.douta(w_n4090_1[0]),.doutb(w_n4090_1[1]),.doutc(w_n4090_1[2]),.din(w_n4090_0[0]));
	jspl jspl_w_n4092_0(.douta(w_n4092_0[0]),.doutb(w_n4092_0[1]),.din(n4092));
	jspl jspl_w_n4099_0(.douta(w_n4099_0[0]),.doutb(w_n4099_0[1]),.din(n4099));
	jspl jspl_w_n4100_0(.douta(w_n4100_0[0]),.doutb(w_n4100_0[1]),.din(n4100));
	jspl jspl_w_n4101_0(.douta(w_n4101_0[0]),.doutb(w_n4101_0[1]),.din(n4101));
	jspl jspl_w_n4106_0(.douta(w_n4106_0[0]),.doutb(w_n4106_0[1]),.din(n4106));
	jspl jspl_w_n4116_0(.douta(w_n4116_0[0]),.doutb(w_n4116_0[1]),.din(n4116));
	jspl jspl_w_n4117_0(.douta(w_n4117_0[0]),.doutb(w_n4117_0[1]),.din(n4117));
	jspl jspl_w_n4118_0(.douta(w_n4118_0[0]),.doutb(w_n4118_0[1]),.din(n4118));
	jspl jspl_w_n4119_0(.douta(w_n4119_0[0]),.doutb(w_n4119_0[1]),.din(n4119));
	jspl jspl_w_n4120_0(.douta(w_dff_A_l5ALSQ9k4_0),.doutb(w_n4120_0[1]),.din(n4120));
	jspl jspl_w_n4123_0(.douta(w_dff_A_vDPcnB1Q5_0),.doutb(w_n4123_0[1]),.din(n4123));
	jspl jspl_w_n4125_0(.douta(w_n4125_0[0]),.doutb(w_n4125_0[1]),.din(n4125));
	jspl jspl_w_n4129_0(.douta(w_n4129_0[0]),.doutb(w_n4129_0[1]),.din(n4129));
	jspl jspl_w_n4132_0(.douta(w_n4132_0[0]),.doutb(w_n4132_0[1]),.din(n4132));
	jspl jspl_w_n4135_0(.douta(w_n4135_0[0]),.doutb(w_n4135_0[1]),.din(n4135));
	jspl3 jspl3_w_n4136_0(.douta(w_n4136_0[0]),.doutb(w_n4136_0[1]),.doutc(w_n4136_0[2]),.din(n4136));
	jspl3 jspl3_w_n4136_1(.douta(w_n4136_1[0]),.doutb(w_n4136_1[1]),.doutc(w_n4136_1[2]),.din(w_n4136_0[0]));
	jspl jspl_w_n4141_0(.douta(w_n4141_0[0]),.doutb(w_n4141_0[1]),.din(n4141));
	jspl jspl_w_n4144_0(.douta(w_n4144_0[0]),.doutb(w_n4144_0[1]),.din(n4144));
	jspl jspl_w_n4153_0(.douta(w_n4153_0[0]),.doutb(w_n4153_0[1]),.din(n4153));
	jspl jspl_w_n4156_0(.douta(w_n4156_0[0]),.doutb(w_n4156_0[1]),.din(n4156));
	jspl jspl_w_n4164_0(.douta(w_n4164_0[0]),.doutb(w_n4164_0[1]),.din(n4164));
	jspl jspl_w_n4172_0(.douta(w_n4172_0[0]),.doutb(w_n4172_0[1]),.din(n4172));
	jspl jspl_w_n4173_0(.douta(w_n4173_0[0]),.doutb(w_n4173_0[1]),.din(n4173));
	jspl jspl_w_n4177_0(.douta(w_n4177_0[0]),.doutb(w_n4177_0[1]),.din(n4177));
	jspl jspl_w_n4178_0(.douta(w_n4178_0[0]),.doutb(w_n4178_0[1]),.din(n4178));
	jspl jspl_w_n4179_0(.douta(w_n4179_0[0]),.doutb(w_n4179_0[1]),.din(n4179));
	jspl jspl_w_n4180_0(.douta(w_n4180_0[0]),.doutb(w_n4180_0[1]),.din(n4180));
	jspl jspl_w_n4181_0(.douta(w_n4181_0[0]),.doutb(w_n4181_0[1]),.din(n4181));
	jspl jspl_w_n4182_0(.douta(w_n4182_0[0]),.doutb(w_n4182_0[1]),.din(n4182));
	jspl jspl_w_n4190_0(.douta(w_n4190_0[0]),.doutb(w_n4190_0[1]),.din(n4190));
	jspl jspl_w_n4191_0(.douta(w_n4191_0[0]),.doutb(w_n4191_0[1]),.din(n4191));
	jspl jspl_w_n4192_0(.douta(w_n4192_0[0]),.doutb(w_n4192_0[1]),.din(n4192));
	jspl jspl_w_n4193_0(.douta(w_n4193_0[0]),.doutb(w_n4193_0[1]),.din(n4193));
	jspl jspl_w_n4194_0(.douta(w_n4194_0[0]),.doutb(w_n4194_0[1]),.din(n4194));
	jspl jspl_w_n4206_0(.douta(w_n4206_0[0]),.doutb(w_n4206_0[1]),.din(n4206));
	jspl jspl_w_n4207_0(.douta(w_n4207_0[0]),.doutb(w_n4207_0[1]),.din(n4207));
	jspl jspl_w_n4208_0(.douta(w_n4208_0[0]),.doutb(w_n4208_0[1]),.din(n4208));
	jspl jspl_w_n4209_0(.douta(w_n4209_0[0]),.doutb(w_n4209_0[1]),.din(n4209));
	jspl jspl_w_n4211_0(.douta(w_n4211_0[0]),.doutb(w_n4211_0[1]),.din(n4211));
	jspl jspl_w_n4215_0(.douta(w_n4215_0[0]),.doutb(w_n4215_0[1]),.din(n4215));
	jspl jspl_w_n4218_0(.douta(w_n4218_0[0]),.doutb(w_n4218_0[1]),.din(n4218));
	jspl jspl_w_n4221_0(.douta(w_n4221_0[0]),.doutb(w_n4221_0[1]),.din(n4221));
	jspl jspl_w_n4224_0(.douta(w_n4224_0[0]),.doutb(w_n4224_0[1]),.din(n4224));
	jspl jspl_w_n4233_0(.douta(w_n4233_0[0]),.doutb(w_n4233_0[1]),.din(n4233));
	jspl jspl_w_n4236_0(.douta(w_n4236_0[0]),.doutb(w_n4236_0[1]),.din(n4236));
	jspl jspl_w_n4245_0(.douta(w_n4245_0[0]),.doutb(w_n4245_0[1]),.din(n4245));
	jspl jspl_w_n4246_0(.douta(w_n4246_0[0]),.doutb(w_n4246_0[1]),.din(n4246));
	jspl jspl_w_n4247_0(.douta(w_n4247_0[0]),.doutb(w_n4247_0[1]),.din(n4247));
	jspl jspl_w_n4248_0(.douta(w_n4248_0[0]),.doutb(w_n4248_0[1]),.din(n4248));
	jspl jspl_w_n4253_0(.douta(w_n4253_0[0]),.doutb(w_n4253_0[1]),.din(n4253));
	jspl jspl_w_n4254_0(.douta(w_n4254_0[0]),.doutb(w_n4254_0[1]),.din(n4254));
	jspl jspl_w_n4262_0(.douta(w_n4262_0[0]),.doutb(w_n4262_0[1]),.din(n4262));
	jspl jspl_w_n4263_0(.douta(w_n4263_0[0]),.doutb(w_n4263_0[1]),.din(n4263));
	jspl jspl_w_n4264_0(.douta(w_n4264_0[0]),.doutb(w_n4264_0[1]),.din(n4264));
	jspl jspl_w_n4265_0(.douta(w_n4265_0[0]),.doutb(w_n4265_0[1]),.din(n4265));
	jspl jspl_w_n4266_0(.douta(w_n4266_0[0]),.doutb(w_n4266_0[1]),.din(n4266));
	jspl jspl_w_n4274_0(.douta(w_n4274_0[0]),.doutb(w_n4274_0[1]),.din(n4274));
	jspl jspl_w_n4275_0(.douta(w_n4275_0[0]),.doutb(w_n4275_0[1]),.din(n4275));
	jspl jspl_w_n4276_0(.douta(w_n4276_0[0]),.doutb(w_n4276_0[1]),.din(n4276));
	jspl jspl_w_n4277_0(.douta(w_n4277_0[0]),.doutb(w_n4277_0[1]),.din(n4277));
	jspl jspl_w_n4286_0(.douta(w_n4286_0[0]),.doutb(w_n4286_0[1]),.din(n4286));
	jspl jspl_w_n4287_0(.douta(w_n4287_0[0]),.doutb(w_n4287_0[1]),.din(n4287));
	jspl jspl_w_n4288_0(.douta(w_n4288_0[0]),.doutb(w_n4288_0[1]),.din(n4288));
	jspl jspl_w_n4289_0(.douta(w_n4289_0[0]),.doutb(w_n4289_0[1]),.din(n4289));
	jspl jspl_w_n4290_0(.douta(w_dff_A_uVwNu9Rb1_0),.doutb(w_n4290_0[1]),.din(n4290));
	jspl jspl_w_n4293_0(.douta(w_n4293_0[0]),.doutb(w_n4293_0[1]),.din(n4293));
	jspl jspl_w_n4297_0(.douta(w_n4297_0[0]),.doutb(w_n4297_0[1]),.din(n4297));
	jspl jspl_w_n4300_0(.douta(w_n4300_0[0]),.doutb(w_n4300_0[1]),.din(n4300));
	jspl jspl_w_n4303_0(.douta(w_n4303_0[0]),.doutb(w_n4303_0[1]),.din(n4303));
	jspl jspl_w_n4309_0(.douta(w_n4309_0[0]),.doutb(w_n4309_0[1]),.din(n4309));
	jspl jspl_w_n4312_0(.douta(w_n4312_0[0]),.doutb(w_n4312_0[1]),.din(n4312));
	jspl jspl_w_n4321_0(.douta(w_n4321_0[0]),.doutb(w_n4321_0[1]),.din(n4321));
	jspl jspl_w_n4324_0(.douta(w_n4324_0[0]),.doutb(w_n4324_0[1]),.din(n4324));
	jspl jspl_w_n4332_0(.douta(w_n4332_0[0]),.doutb(w_n4332_0[1]),.din(n4332));
	jspl jspl_w_n4340_0(.douta(w_n4340_0[0]),.doutb(w_n4340_0[1]),.din(n4340));
	jspl jspl_w_n4343_0(.douta(w_n4343_0[0]),.doutb(w_n4343_0[1]),.din(n4343));
	jspl jspl_w_n4344_0(.douta(w_n4344_0[0]),.doutb(w_n4344_0[1]),.din(n4344));
	jspl jspl_w_n4345_0(.douta(w_n4345_0[0]),.doutb(w_n4345_0[1]),.din(n4345));
	jspl jspl_w_n4346_0(.douta(w_n4346_0[0]),.doutb(w_n4346_0[1]),.din(n4346));
	jspl jspl_w_n4347_0(.douta(w_n4347_0[0]),.doutb(w_n4347_0[1]),.din(n4347));
	jspl jspl_w_n4348_0(.douta(w_n4348_0[0]),.doutb(w_n4348_0[1]),.din(n4348));
	jspl jspl_w_n4349_0(.douta(w_n4349_0[0]),.doutb(w_n4349_0[1]),.din(n4349));
	jspl jspl_w_n4350_0(.douta(w_n4350_0[0]),.doutb(w_n4350_0[1]),.din(n4350));
	jspl jspl_w_n4351_0(.douta(w_n4351_0[0]),.doutb(w_n4351_0[1]),.din(n4351));
	jspl jspl_w_n4352_0(.douta(w_n4352_0[0]),.doutb(w_n4352_0[1]),.din(n4352));
	jspl jspl_w_n4353_0(.douta(w_n4353_0[0]),.doutb(w_n4353_0[1]),.din(n4353));
	jspl jspl_w_n4354_0(.douta(w_n4354_0[0]),.doutb(w_n4354_0[1]),.din(n4354));
	jspl jspl_w_n4355_0(.douta(w_n4355_0[0]),.doutb(w_n4355_0[1]),.din(n4355));
	jspl3 jspl3_w_n4357_0(.douta(w_n4357_0[0]),.doutb(w_n4357_0[1]),.doutc(w_n4357_0[2]),.din(n4357));
	jspl jspl_w_n4368_0(.douta(w_n4368_0[0]),.doutb(w_n4368_0[1]),.din(n4368));
	jspl jspl_w_n4369_0(.douta(w_n4369_0[0]),.doutb(w_n4369_0[1]),.din(n4369));
	jspl jspl_w_n4370_0(.douta(w_n4370_0[0]),.doutb(w_n4370_0[1]),.din(n4370));
	jspl jspl_w_n4371_0(.douta(w_n4371_0[0]),.doutb(w_n4371_0[1]),.din(n4371));
	jspl jspl_w_n4372_0(.douta(w_dff_A_t9pi2k7w5_0),.doutb(w_n4372_0[1]),.din(n4372));
	jspl jspl_w_n4375_0(.douta(w_n4375_0[0]),.doutb(w_n4375_0[1]),.din(n4375));
	jspl jspl_w_n4379_0(.douta(w_n4379_0[0]),.doutb(w_n4379_0[1]),.din(n4379));
	jspl jspl_w_n4382_0(.douta(w_n4382_0[0]),.doutb(w_n4382_0[1]),.din(n4382));
	jspl jspl_w_n4385_0(.douta(w_n4385_0[0]),.doutb(w_n4385_0[1]),.din(n4385));
	jspl jspl_w_n4389_0(.douta(w_n4389_0[0]),.doutb(w_n4389_0[1]),.din(n4389));
	jspl jspl_w_n4393_0(.douta(w_n4393_0[0]),.doutb(w_n4393_0[1]),.din(n4393));
	jspl jspl_w_n4394_0(.douta(w_n4394_0[0]),.doutb(w_n4394_0[1]),.din(n4394));
	jspl jspl_w_n4403_0(.douta(w_n4403_0[0]),.doutb(w_n4403_0[1]),.din(n4403));
	jspl jspl_w_n4406_0(.douta(w_n4406_0[0]),.doutb(w_n4406_0[1]),.din(n4406));
	jspl jspl_w_n4414_0(.douta(w_n4414_0[0]),.doutb(w_n4414_0[1]),.din(n4414));
	jspl jspl_w_n4422_0(.douta(w_n4422_0[0]),.doutb(w_n4422_0[1]),.din(n4422));
	jspl jspl_w_n4425_0(.douta(w_n4425_0[0]),.doutb(w_n4425_0[1]),.din(n4425));
	jspl jspl_w_n4426_0(.douta(w_n4426_0[0]),.doutb(w_n4426_0[1]),.din(n4426));
	jspl jspl_w_n4427_0(.douta(w_n4427_0[0]),.doutb(w_n4427_0[1]),.din(n4427));
	jspl jspl_w_n4428_0(.douta(w_n4428_0[0]),.doutb(w_n4428_0[1]),.din(n4428));
	jspl jspl_w_n4429_0(.douta(w_n4429_0[0]),.doutb(w_n4429_0[1]),.din(n4429));
	jspl jspl_w_n4430_0(.douta(w_n4430_0[0]),.doutb(w_n4430_0[1]),.din(n4430));
	jspl jspl_w_n4431_0(.douta(w_n4431_0[0]),.doutb(w_n4431_0[1]),.din(n4431));
	jspl jspl_w_n4432_0(.douta(w_n4432_0[0]),.doutb(w_n4432_0[1]),.din(n4432));
	jspl jspl_w_n4433_0(.douta(w_n4433_0[0]),.doutb(w_n4433_0[1]),.din(n4433));
	jspl jspl_w_n4434_0(.douta(w_n4434_0[0]),.doutb(w_n4434_0[1]),.din(n4434));
	jspl jspl_w_n4435_0(.douta(w_n4435_0[0]),.doutb(w_n4435_0[1]),.din(n4435));
	jspl jspl_w_n4442_0(.douta(w_n4442_0[0]),.doutb(w_n4442_0[1]),.din(n4442));
	jspl jspl_w_n4450_0(.douta(w_n4450_0[0]),.doutb(w_n4450_0[1]),.din(n4450));
	jspl jspl_w_n4451_0(.douta(w_n4451_0[0]),.doutb(w_n4451_0[1]),.din(n4451));
	jspl jspl_w_n4452_0(.douta(w_n4452_0[0]),.doutb(w_n4452_0[1]),.din(n4452));
	jspl jspl_w_n4453_0(.douta(w_n4453_0[0]),.doutb(w_n4453_0[1]),.din(n4453));
	jspl jspl_w_n4454_0(.douta(w_dff_A_gjRzRkwI1_0),.doutb(w_n4454_0[1]),.din(n4454));
	jspl jspl_w_n4457_0(.douta(w_n4457_0[0]),.doutb(w_n4457_0[1]),.din(n4457));
	jspl jspl_w_n4461_0(.douta(w_n4461_0[0]),.doutb(w_n4461_0[1]),.din(n4461));
	jspl jspl_w_n4464_0(.douta(w_n4464_0[0]),.doutb(w_n4464_0[1]),.din(n4464));
	jspl jspl_w_n4469_0(.douta(w_n4469_0[0]),.doutb(w_n4469_0[1]),.din(n4469));
	jspl jspl_w_n4472_0(.douta(w_n4472_0[0]),.doutb(w_n4472_0[1]),.din(n4472));
	jspl jspl_w_n4480_0(.douta(w_n4480_0[0]),.doutb(w_n4480_0[1]),.din(n4480));
	jspl jspl_w_n4481_0(.douta(w_n4481_0[0]),.doutb(w_n4481_0[1]),.din(n4481));
	jspl jspl_w_n4484_0(.douta(w_n4484_0[0]),.doutb(w_n4484_0[1]),.din(n4484));
	jspl jspl_w_n4487_0(.douta(w_n4487_0[0]),.doutb(w_n4487_0[1]),.din(n4487));
	jspl jspl_w_n4496_0(.douta(w_n4496_0[0]),.doutb(w_n4496_0[1]),.din(n4496));
	jspl jspl_w_n4497_0(.douta(w_n4497_0[0]),.doutb(w_n4497_0[1]),.din(n4497));
	jspl jspl_w_n4498_0(.douta(w_n4498_0[0]),.doutb(w_n4498_0[1]),.din(n4498));
	jspl jspl_w_n4499_0(.douta(w_n4499_0[0]),.doutb(w_n4499_0[1]),.din(n4499));
	jspl jspl_w_n4500_0(.douta(w_n4500_0[0]),.doutb(w_n4500_0[1]),.din(n4500));
	jspl jspl_w_n4501_0(.douta(w_n4501_0[0]),.doutb(w_n4501_0[1]),.din(n4501));
	jspl jspl_w_n4509_0(.douta(w_n4509_0[0]),.doutb(w_n4509_0[1]),.din(n4509));
	jspl jspl_w_n4510_0(.douta(w_n4510_0[0]),.doutb(w_n4510_0[1]),.din(n4510));
	jspl jspl_w_n4511_0(.douta(w_n4511_0[0]),.doutb(w_n4511_0[1]),.din(n4511));
	jspl jspl_w_n4512_0(.douta(w_n4512_0[0]),.doutb(w_n4512_0[1]),.din(n4512));
	jspl jspl_w_n4513_0(.douta(w_n4513_0[0]),.doutb(w_n4513_0[1]),.din(n4513));
	jspl jspl_w_n4514_0(.douta(w_n4514_0[0]),.doutb(w_n4514_0[1]),.din(n4514));
	jspl jspl_w_n4523_0(.douta(w_n4523_0[0]),.doutb(w_n4523_0[1]),.din(n4523));
	jspl jspl_w_n4524_0(.douta(w_n4524_0[0]),.doutb(w_n4524_0[1]),.din(n4524));
	jspl jspl_w_n4525_0(.douta(w_n4525_0[0]),.doutb(w_n4525_0[1]),.din(n4525));
	jspl jspl_w_n4526_0(.douta(w_n4526_0[0]),.doutb(w_n4526_0[1]),.din(n4526));
	jspl jspl_w_n4527_0(.douta(w_dff_A_SMxcsPby6_0),.doutb(w_n4527_0[1]),.din(n4527));
	jspl jspl_w_n4530_0(.douta(w_n4530_0[0]),.doutb(w_n4530_0[1]),.din(n4530));
	jspl jspl_w_n4534_0(.douta(w_n4534_0[0]),.doutb(w_n4534_0[1]),.din(n4534));
	jspl jspl_w_n4537_0(.douta(w_n4537_0[0]),.doutb(w_n4537_0[1]),.din(n4537));
	jspl jspl_w_n4540_0(.douta(w_n4540_0[0]),.doutb(w_n4540_0[1]),.din(n4540));
	jspl jspl_w_n4547_0(.douta(w_n4547_0[0]),.doutb(w_n4547_0[1]),.din(n4547));
	jspl jspl_w_n4550_0(.douta(w_n4550_0[0]),.doutb(w_n4550_0[1]),.din(n4550));
	jspl jspl_w_n4558_0(.douta(w_n4558_0[0]),.doutb(w_n4558_0[1]),.din(n4558));
	jspl jspl_w_n4561_0(.douta(w_n4561_0[0]),.doutb(w_n4561_0[1]),.din(n4561));
	jspl jspl_w_n4569_0(.douta(w_n4569_0[0]),.doutb(w_n4569_0[1]),.din(n4569));
	jspl jspl_w_n4570_0(.douta(w_n4570_0[0]),.doutb(w_n4570_0[1]),.din(n4570));
	jspl3 jspl3_w_n4571_0(.douta(w_n4571_0[0]),.doutb(w_n4571_0[1]),.doutc(w_n4571_0[2]),.din(n4571));
	jspl jspl_w_n4574_0(.douta(w_n4574_0[0]),.doutb(w_n4574_0[1]),.din(n4574));
	jspl jspl_w_n4575_0(.douta(w_n4575_0[0]),.doutb(w_n4575_0[1]),.din(n4575));
	jspl jspl_w_n4576_0(.douta(w_n4576_0[0]),.doutb(w_n4576_0[1]),.din(n4576));
	jspl jspl_w_n4577_0(.douta(w_n4577_0[0]),.doutb(w_n4577_0[1]),.din(n4577));
	jspl jspl_w_n4578_0(.douta(w_n4578_0[0]),.doutb(w_n4578_0[1]),.din(n4578));
	jspl jspl_w_n4579_0(.douta(w_n4579_0[0]),.doutb(w_n4579_0[1]),.din(n4579));
	jspl jspl_w_n4580_0(.douta(w_n4580_0[0]),.doutb(w_n4580_0[1]),.din(n4580));
	jspl jspl_w_n4581_0(.douta(w_n4581_0[0]),.doutb(w_n4581_0[1]),.din(n4581));
	jspl jspl_w_n4582_0(.douta(w_n4582_0[0]),.doutb(w_n4582_0[1]),.din(n4582));
	jspl jspl_w_n4589_0(.douta(w_n4589_0[0]),.doutb(w_n4589_0[1]),.din(n4589));
	jspl jspl_w_n4599_0(.douta(w_n4599_0[0]),.doutb(w_n4599_0[1]),.din(n4599));
	jspl jspl_w_n4600_0(.douta(w_n4600_0[0]),.doutb(w_n4600_0[1]),.din(n4600));
	jspl jspl_w_n4601_0(.douta(w_n4601_0[0]),.doutb(w_n4601_0[1]),.din(n4601));
	jspl jspl_w_n4602_0(.douta(w_n4602_0[0]),.doutb(w_n4602_0[1]),.din(n4602));
	jspl jspl_w_n4603_0(.douta(w_dff_A_h9g6HZkd4_0),.doutb(w_n4603_0[1]),.din(n4603));
	jspl jspl_w_n4606_0(.douta(w_n4606_0[0]),.doutb(w_n4606_0[1]),.din(n4606));
	jspl jspl_w_n4610_0(.douta(w_n4610_0[0]),.doutb(w_n4610_0[1]),.din(n4610));
	jspl jspl_w_n4613_0(.douta(w_n4613_0[0]),.doutb(w_n4613_0[1]),.din(n4613));
	jspl jspl_w_n4616_0(.douta(w_n4616_0[0]),.doutb(w_n4616_0[1]),.din(n4616));
	jspl jspl_w_n4620_0(.douta(w_n4620_0[0]),.doutb(w_n4620_0[1]),.din(n4620));
	jspl jspl_w_n4624_0(.douta(w_n4624_0[0]),.doutb(w_n4624_0[1]),.din(n4624));
	jspl jspl_w_n4625_0(.douta(w_n4625_0[0]),.doutb(w_n4625_0[1]),.din(n4625));
	jspl jspl_w_n4628_0(.douta(w_n4628_0[0]),.doutb(w_n4628_0[1]),.din(n4628));
	jspl jspl_w_n4636_0(.douta(w_n4636_0[0]),.doutb(w_n4636_0[1]),.din(n4636));
	jspl jspl_w_n4637_0(.douta(w_n4637_0[0]),.doutb(w_n4637_0[1]),.din(n4637));
	jspl jspl_w_n4638_0(.douta(w_n4638_0[0]),.doutb(w_n4638_0[1]),.din(n4638));
	jspl jspl_w_n4639_0(.douta(w_n4639_0[0]),.doutb(w_n4639_0[1]),.din(n4639));
	jspl jspl_w_n4647_0(.douta(w_n4647_0[0]),.doutb(w_n4647_0[1]),.din(n4647));
	jspl jspl_w_n4648_0(.douta(w_n4648_0[0]),.doutb(w_n4648_0[1]),.din(n4648));
	jspl jspl_w_n4649_0(.douta(w_n4649_0[0]),.doutb(w_n4649_0[1]),.din(n4649));
	jspl jspl_w_n4650_0(.douta(w_n4650_0[0]),.doutb(w_n4650_0[1]),.din(n4650));
	jspl jspl_w_n4651_0(.douta(w_n4651_0[0]),.doutb(w_n4651_0[1]),.din(n4651));
	jspl jspl_w_n4663_0(.douta(w_n4663_0[0]),.doutb(w_n4663_0[1]),.din(n4663));
	jspl jspl_w_n4664_0(.douta(w_n4664_0[0]),.doutb(w_n4664_0[1]),.din(n4664));
	jspl jspl_w_n4665_0(.douta(w_n4665_0[0]),.doutb(w_n4665_0[1]),.din(n4665));
	jspl jspl_w_n4666_0(.douta(w_n4666_0[0]),.doutb(w_n4666_0[1]),.din(n4666));
	jspl jspl_w_n4667_0(.douta(w_dff_A_J0qwBfzZ9_0),.doutb(w_n4667_0[1]),.din(n4667));
	jspl jspl_w_n4670_0(.douta(w_n4670_0[0]),.doutb(w_n4670_0[1]),.din(n4670));
	jspl jspl_w_n4674_0(.douta(w_n4674_0[0]),.doutb(w_n4674_0[1]),.din(n4674));
	jspl jspl_w_n4677_0(.douta(w_n4677_0[0]),.doutb(w_n4677_0[1]),.din(n4677));
	jspl jspl_w_n4682_0(.douta(w_n4682_0[0]),.doutb(w_n4682_0[1]),.din(n4682));
	jspl jspl_w_n4685_0(.douta(w_n4685_0[0]),.doutb(w_n4685_0[1]),.din(n4685));
	jspl jspl_w_n4693_0(.douta(w_n4693_0[0]),.doutb(w_n4693_0[1]),.din(n4693));
	jspl jspl_w_n4694_0(.douta(w_n4694_0[0]),.doutb(w_n4694_0[1]),.din(n4694));
	jspl jspl_w_n4703_0(.douta(w_n4703_0[0]),.doutb(w_n4703_0[1]),.din(n4703));
	jspl3 jspl3_w_n4704_0(.douta(w_n4704_0[0]),.doutb(w_n4704_0[1]),.doutc(w_n4704_0[2]),.din(n4704));
	jspl3 jspl3_w_n4706_0(.douta(w_n4706_0[0]),.doutb(w_n4706_0[1]),.doutc(w_n4706_0[2]),.din(n4706));
	jspl3 jspl3_w_n4711_0(.douta(w_n4711_0[0]),.doutb(w_n4711_0[1]),.doutc(w_n4711_0[2]),.din(n4711));
	jspl jspl_w_n4713_0(.douta(w_n4713_0[0]),.doutb(w_n4713_0[1]),.din(n4713));
	jspl jspl_w_n4714_0(.douta(w_n4714_0[0]),.doutb(w_n4714_0[1]),.din(n4714));
	jspl jspl_w_n4715_0(.douta(w_n4715_0[0]),.doutb(w_n4715_0[1]),.din(n4715));
	jspl jspl_w_n4716_0(.douta(w_n4716_0[0]),.doutb(w_n4716_0[1]),.din(n4716));
	jspl jspl_w_n4728_0(.douta(w_n4728_0[0]),.doutb(w_n4728_0[1]),.din(n4728));
	jspl jspl_w_n4729_0(.douta(w_n4729_0[0]),.doutb(w_n4729_0[1]),.din(n4729));
	jspl jspl_w_n4730_0(.douta(w_n4730_0[0]),.doutb(w_n4730_0[1]),.din(n4730));
	jspl jspl_w_n4731_0(.douta(w_n4731_0[0]),.doutb(w_n4731_0[1]),.din(n4731));
	jspl jspl_w_n4732_0(.douta(w_dff_A_72JVXFet2_0),.doutb(w_n4732_0[1]),.din(n4732));
	jspl jspl_w_n4735_0(.douta(w_n4735_0[0]),.doutb(w_n4735_0[1]),.din(n4735));
	jspl jspl_w_n4739_0(.douta(w_n4739_0[0]),.doutb(w_n4739_0[1]),.din(n4739));
	jspl jspl_w_n4742_0(.douta(w_n4742_0[0]),.doutb(w_n4742_0[1]),.din(n4742));
	jspl jspl_w_n4745_0(.douta(w_n4745_0[0]),.doutb(w_n4745_0[1]),.din(n4745));
	jspl jspl_w_n4751_0(.douta(w_n4751_0[0]),.doutb(w_n4751_0[1]),.din(n4751));
	jspl jspl_w_n4759_0(.douta(w_n4759_0[0]),.doutb(w_n4759_0[1]),.din(n4759));
	jspl3 jspl3_w_n4760_0(.douta(w_n4760_0[0]),.doutb(w_n4760_0[1]),.doutc(w_n4760_0[2]),.din(n4760));
	jspl jspl_w_n4766_0(.douta(w_n4766_0[0]),.doutb(w_n4766_0[1]),.din(n4766));
	jspl jspl_w_n4767_0(.douta(w_n4767_0[0]),.doutb(w_n4767_0[1]),.din(n4767));
	jspl jspl_w_n4768_0(.douta(w_n4768_0[0]),.doutb(w_n4768_0[1]),.din(n4768));
	jspl jspl_w_n4775_0(.douta(w_n4775_0[0]),.doutb(w_n4775_0[1]),.din(n4775));
	jspl jspl_w_n4776_0(.douta(w_n4776_0[0]),.doutb(w_n4776_0[1]),.din(n4776));
	jspl jspl_w_n4777_0(.douta(w_n4777_0[0]),.doutb(w_n4777_0[1]),.din(n4777));
	jspl jspl_w_n4778_0(.douta(w_n4778_0[0]),.doutb(w_n4778_0[1]),.din(n4778));
	jspl jspl_w_n4779_0(.douta(w_n4779_0[0]),.doutb(w_n4779_0[1]),.din(n4779));
	jspl jspl_w_n4785_0(.douta(w_n4785_0[0]),.doutb(w_n4785_0[1]),.din(n4785));
	jspl jspl_w_n4786_0(.douta(w_n4786_0[0]),.doutb(w_n4786_0[1]),.din(n4786));
	jspl jspl_w_n4787_0(.douta(w_n4787_0[0]),.doutb(w_n4787_0[1]),.din(n4787));
	jspl jspl_w_n4788_0(.douta(w_n4788_0[0]),.doutb(w_n4788_0[1]),.din(n4788));
	jspl jspl_w_n4789_0(.douta(w_dff_A_fGY52gbv0_0),.doutb(w_n4789_0[1]),.din(n4789));
	jspl jspl_w_n4792_0(.douta(w_n4792_0[0]),.doutb(w_n4792_0[1]),.din(n4792));
	jspl jspl_w_n4796_0(.douta(w_n4796_0[0]),.doutb(w_n4796_0[1]),.din(n4796));
	jspl jspl_w_n4799_0(.douta(w_n4799_0[0]),.doutb(w_n4799_0[1]),.din(n4799));
	jspl jspl_w_n4802_0(.douta(w_n4802_0[0]),.doutb(w_n4802_0[1]),.din(n4802));
	jspl jspl_w_n4806_0(.douta(w_n4806_0[0]),.doutb(w_n4806_0[1]),.din(n4806));
	jspl jspl_w_n4807_0(.douta(w_n4807_0[0]),.doutb(w_n4807_0[1]),.din(n4807));
	jspl jspl_w_n4808_0(.douta(w_n4808_0[0]),.doutb(w_n4808_0[1]),.din(n4808));
	jspl jspl_w_n4816_0(.douta(w_n4816_0[0]),.doutb(w_n4816_0[1]),.din(n4816));
	jspl jspl_w_n4820_0(.douta(w_n4820_0[0]),.doutb(w_n4820_0[1]),.din(n4820));
	jspl jspl_w_n4821_0(.douta(w_n4821_0[0]),.doutb(w_n4821_0[1]),.din(n4821));
	jspl jspl_w_n4822_0(.douta(w_n4822_0[0]),.doutb(w_n4822_0[1]),.din(n4822));
	jspl jspl_w_n4823_0(.douta(w_n4823_0[0]),.doutb(w_n4823_0[1]),.din(n4823));
	jspl jspl_w_n4824_0(.douta(w_n4824_0[0]),.doutb(w_n4824_0[1]),.din(n4824));
	jspl jspl_w_n4832_0(.douta(w_n4832_0[0]),.doutb(w_n4832_0[1]),.din(n4832));
	jspl jspl_w_n4836_0(.douta(w_n4836_0[0]),.doutb(w_n4836_0[1]),.din(n4836));
	jspl jspl_w_n4837_0(.douta(w_n4837_0[0]),.doutb(w_n4837_0[1]),.din(n4837));
	jspl jspl_w_n4838_0(.douta(w_n4838_0[0]),.doutb(w_n4838_0[1]),.din(n4838));
	jspl jspl_w_n4839_0(.douta(w_n4839_0[0]),.doutb(w_n4839_0[1]),.din(n4839));
	jspl jspl_w_n4840_0(.douta(w_dff_A_sOErIqr07_0),.doutb(w_n4840_0[1]),.din(n4840));
	jspl jspl_w_n4843_0(.douta(w_n4843_0[0]),.doutb(w_n4843_0[1]),.din(n4843));
	jspl jspl_w_n4847_0(.douta(w_n4847_0[0]),.doutb(w_n4847_0[1]),.din(n4847));
	jspl jspl_w_n4850_0(.douta(w_n4850_0[0]),.doutb(w_n4850_0[1]),.din(n4850));
	jspl jspl_w_n4855_0(.douta(w_n4855_0[0]),.doutb(w_n4855_0[1]),.din(n4855));
	jspl jspl_w_n4859_0(.douta(w_n4859_0[0]),.doutb(w_n4859_0[1]),.din(n4859));
	jspl jspl_w_n4868_0(.douta(w_n4868_0[0]),.doutb(w_n4868_0[1]),.din(n4868));
	jspl jspl_w_n4869_0(.douta(w_n4869_0[0]),.doutb(w_n4869_0[1]),.din(n4869));
	jspl jspl_w_n4870_0(.douta(w_n4870_0[0]),.doutb(w_n4870_0[1]),.din(n4870));
	jspl jspl_w_n4871_0(.douta(w_n4871_0[0]),.doutb(w_n4871_0[1]),.din(n4871));
	jspl jspl_w_n4872_0(.douta(w_n4872_0[0]),.doutb(w_n4872_0[1]),.din(n4872));
	jspl jspl_w_n4873_0(.douta(w_n4873_0[0]),.doutb(w_n4873_0[1]),.din(n4873));
	jspl jspl_w_n4874_0(.douta(w_n4874_0[0]),.doutb(w_n4874_0[1]),.din(n4874));
	jspl jspl_w_n4875_0(.douta(w_n4875_0[0]),.doutb(w_n4875_0[1]),.din(n4875));
	jspl jspl_w_n4876_0(.douta(w_n4876_0[0]),.doutb(w_n4876_0[1]),.din(n4876));
	jspl jspl_w_n4880_0(.douta(w_n4880_0[0]),.doutb(w_n4880_0[1]),.din(n4880));
	jspl jspl_w_n4892_0(.douta(w_n4892_0[0]),.doutb(w_n4892_0[1]),.din(n4892));
	jspl jspl_w_n4893_0(.douta(w_n4893_0[0]),.doutb(w_n4893_0[1]),.din(n4893));
	jspl jspl_w_n4894_0(.douta(w_n4894_0[0]),.doutb(w_n4894_0[1]),.din(n4894));
	jspl jspl_w_n4895_0(.douta(w_n4895_0[0]),.doutb(w_n4895_0[1]),.din(n4895));
	jspl jspl_w_n4896_0(.douta(w_dff_A_yIbGSoVr3_0),.doutb(w_n4896_0[1]),.din(n4896));
	jspl jspl_w_n4899_0(.douta(w_n4899_0[0]),.doutb(w_n4899_0[1]),.din(n4899));
	jspl jspl_w_n4903_0(.douta(w_n4903_0[0]),.doutb(w_n4903_0[1]),.din(n4903));
	jspl jspl_w_n4906_0(.douta(w_n4906_0[0]),.doutb(w_n4906_0[1]),.din(n4906));
	jspl jspl_w_n4909_0(.douta(w_n4909_0[0]),.doutb(w_n4909_0[1]),.din(n4909));
	jspl jspl_w_n4915_0(.douta(w_n4915_0[0]),.doutb(w_n4915_0[1]),.din(n4915));
	jspl jspl_w_n4917_0(.douta(w_n4917_0[0]),.doutb(w_n4917_0[1]),.din(n4917));
	jspl jspl_w_n4920_0(.douta(w_n4920_0[0]),.doutb(w_n4920_0[1]),.din(n4920));
	jspl jspl_w_n4921_0(.douta(w_n4921_0[0]),.doutb(w_n4921_0[1]),.din(n4921));
	jspl jspl_w_n4922_0(.douta(w_n4922_0[0]),.doutb(w_n4922_0[1]),.din(n4922));
	jspl jspl_w_n4923_0(.douta(w_n4923_0[0]),.doutb(w_n4923_0[1]),.din(n4923));
	jspl jspl_w_n4924_0(.douta(w_n4924_0[0]),.doutb(w_n4924_0[1]),.din(n4924));
	jspl jspl_w_n4931_0(.douta(w_n4931_0[0]),.doutb(w_n4931_0[1]),.din(n4931));
	jspl jspl_w_n4939_0(.douta(w_n4939_0[0]),.doutb(w_n4939_0[1]),.din(n4939));
	jspl jspl_w_n4940_0(.douta(w_n4940_0[0]),.doutb(w_n4940_0[1]),.din(n4940));
	jspl jspl_w_n4941_0(.douta(w_n4941_0[0]),.doutb(w_n4941_0[1]),.din(n4941));
	jspl jspl_w_n4942_0(.douta(w_n4942_0[0]),.doutb(w_n4942_0[1]),.din(n4942));
	jspl jspl_w_n4943_0(.douta(w_dff_A_e94k11f77_0),.doutb(w_n4943_0[1]),.din(n4943));
	jspl jspl_w_n4946_0(.douta(w_n4946_0[0]),.doutb(w_n4946_0[1]),.din(n4946));
	jspl jspl_w_n4950_0(.douta(w_n4950_0[0]),.doutb(w_n4950_0[1]),.din(n4950));
	jspl jspl_w_n4953_0(.douta(w_n4953_0[0]),.doutb(w_n4953_0[1]),.din(n4953));
	jspl jspl_w_n4957_0(.douta(w_n4957_0[0]),.doutb(w_n4957_0[1]),.din(n4957));
	jspl jspl_w_n4959_0(.douta(w_n4959_0[0]),.doutb(w_n4959_0[1]),.din(n4959));
	jspl jspl_w_n4960_0(.douta(w_n4960_0[0]),.doutb(w_n4960_0[1]),.din(n4960));
	jspl jspl_w_n4964_0(.douta(w_n4964_0[0]),.doutb(w_n4964_0[1]),.din(n4964));
	jspl jspl_w_n4965_0(.douta(w_n4965_0[0]),.doutb(w_n4965_0[1]),.din(n4965));
	jspl jspl_w_n4968_0(.douta(w_n4968_0[0]),.doutb(w_n4968_0[1]),.din(n4968));
	jspl jspl_w_n4969_0(.douta(w_n4969_0[0]),.doutb(w_n4969_0[1]),.din(n4969));
	jspl jspl_w_n4972_0(.douta(w_n4972_0[0]),.doutb(w_n4972_0[1]),.din(n4972));
	jspl jspl_w_n4982_0(.douta(w_n4982_0[0]),.doutb(w_n4982_0[1]),.din(n4982));
	jspl jspl_w_n4983_0(.douta(w_n4983_0[0]),.doutb(w_n4983_0[1]),.din(n4983));
	jspl jspl_w_n4984_0(.douta(w_n4984_0[0]),.doutb(w_n4984_0[1]),.din(n4984));
	jspl jspl_w_n4985_0(.douta(w_n4985_0[0]),.doutb(w_n4985_0[1]),.din(n4985));
	jspl jspl_w_n4986_0(.douta(w_dff_A_wxzz2WBi3_0),.doutb(w_n4986_0[1]),.din(n4986));
	jspl jspl_w_n4989_0(.douta(w_n4989_0[0]),.doutb(w_n4989_0[1]),.din(n4989));
	jspl jspl_w_n4993_0(.douta(w_n4993_0[0]),.doutb(w_n4993_0[1]),.din(n4993));
	jspl jspl_w_n4994_0(.douta(w_n4994_0[0]),.doutb(w_n4994_0[1]),.din(n4994));
	jspl3 jspl3_w_n5003_0(.douta(w_n5003_0[0]),.doutb(w_n5003_0[1]),.doutc(w_n5003_0[2]),.din(n5003));
	jspl jspl_w_n5007_0(.douta(w_n5007_0[0]),.doutb(w_n5007_0[1]),.din(n5007));
	jspl jspl_w_n5016_0(.douta(w_n5016_0[0]),.doutb(w_n5016_0[1]),.din(n5016));
	jspl jspl_w_n5017_0(.douta(w_n5017_0[0]),.doutb(w_n5017_0[1]),.din(n5017));
	jspl jspl_w_n5018_0(.douta(w_n5018_0[0]),.doutb(w_n5018_0[1]),.din(n5018));
	jspl jspl_w_n5019_0(.douta(w_n5019_0[0]),.doutb(w_n5019_0[1]),.din(n5019));
	jspl jspl_w_n5020_0(.douta(w_n5020_0[0]),.doutb(w_n5020_0[1]),.din(n5020));
	jspl jspl_w_n5021_0(.douta(w_dff_A_HPuTasns0_0),.doutb(w_n5021_0[1]),.din(n5021));
	jspl3 jspl3_w_n5024_0(.douta(w_dff_A_Xhuy3IJF7_0),.doutb(w_n5024_0[1]),.doutc(w_n5024_0[2]),.din(n5024));
	jspl3 jspl3_w_n5026_0(.douta(w_n5026_0[0]),.doutb(w_n5026_0[1]),.doutc(w_n5026_0[2]),.din(n5026));
	jspl jspl_w_n5027_0(.douta(w_n5027_0[0]),.doutb(w_n5027_0[1]),.din(n5027));
	jspl jspl_w_n5031_0(.douta(w_n5031_0[0]),.doutb(w_n5031_0[1]),.din(n5031));
	jspl3 jspl3_w_n5042_0(.douta(w_n5042_0[0]),.doutb(w_n5042_0[1]),.doutc(w_n5042_0[2]),.din(n5042));
	jspl jspl_w_n5042_1(.douta(w_n5042_1[0]),.doutb(w_n5042_1[1]),.din(w_n5042_0[0]));
	jspl3 jspl3_w_n5043_0(.douta(w_n5043_0[0]),.doutb(w_n5043_0[1]),.doutc(w_n5043_0[2]),.din(n5043));
	jspl jspl_w_n5044_0(.douta(w_n5044_0[0]),.doutb(w_n5044_0[1]),.din(n5044));
	jspl jspl_w_n5046_0(.douta(w_dff_A_bZ09vicW3_0),.doutb(w_n5046_0[1]),.din(w_dff_B_wcw2K1gk7_2));
	jspl jspl_w_n5048_0(.douta(w_n5048_0[0]),.doutb(w_n5048_0[1]),.din(n5048));
	jspl jspl_w_n5050_0(.douta(w_dff_A_h2PYpQyn7_0),.doutb(w_n5050_0[1]),.din(n5050));
	jspl jspl_w_n5054_0(.douta(w_n5054_0[0]),.doutb(w_n5054_0[1]),.din(n5054));
	jspl jspl_w_n5056_0(.douta(w_n5056_0[0]),.doutb(w_n5056_0[1]),.din(n5056));
	jspl jspl_w_n5057_0(.douta(w_n5057_0[0]),.doutb(w_n5057_0[1]),.din(n5057));
	jspl jspl_w_n5058_0(.douta(w_n5058_0[0]),.doutb(w_n5058_0[1]),.din(n5058));
	jspl3 jspl3_w_n5068_0(.douta(w_n5068_0[0]),.doutb(w_n5068_0[1]),.doutc(w_n5068_0[2]),.din(n5068));
	jspl jspl_w_n5068_1(.douta(w_n5068_1[0]),.doutb(w_n5068_1[1]),.din(w_n5068_0[0]));
	jspl jspl_w_n5069_0(.douta(w_n5069_0[0]),.doutb(w_n5069_0[1]),.din(n5069));
	jspl3 jspl3_w_n5081_0(.douta(w_n5081_0[0]),.doutb(w_n5081_0[1]),.doutc(w_n5081_0[2]),.din(n5081));
	jspl jspl_w_n5082_0(.douta(w_n5082_0[0]),.doutb(w_n5082_0[1]),.din(n5082));
	jspl3 jspl3_w_n5083_0(.douta(w_n5083_0[0]),.doutb(w_n5083_0[1]),.doutc(w_n5083_0[2]),.din(n5083));
	jspl3 jspl3_w_n5084_0(.douta(w_n5084_0[0]),.doutb(w_n5084_0[1]),.doutc(w_n5084_0[2]),.din(n5084));
	jspl jspl_w_n5085_0(.douta(w_n5085_0[0]),.doutb(w_dff_A_W48FiSy24_1),.din(w_dff_B_elMsNUXc0_2));
	jspl jspl_w_n5088_0(.douta(w_n5088_0[0]),.doutb(w_n5088_0[1]),.din(n5088));
	jspl jspl_w_n5091_0(.douta(w_n5091_0[0]),.doutb(w_n5091_0[1]),.din(n5091));
	jspl jspl_w_n5092_0(.douta(w_n5092_0[0]),.doutb(w_n5092_0[1]),.din(n5092));
	jspl jspl_w_n5095_0(.douta(w_n5095_0[0]),.doutb(w_n5095_0[1]),.din(n5095));
	jspl jspl_w_n5098_0(.douta(w_n5098_0[0]),.doutb(w_n5098_0[1]),.din(n5098));
	jspl jspl_w_n5099_0(.douta(w_n5099_0[0]),.doutb(w_n5099_0[1]),.din(n5099));
	jspl jspl_w_n5100_0(.douta(w_n5100_0[0]),.doutb(w_n5100_0[1]),.din(n5100));
	jspl3 jspl3_w_n5109_0(.douta(w_n5109_0[0]),.doutb(w_n5109_0[1]),.doutc(w_n5109_0[2]),.din(n5109));
	jspl jspl_w_n5110_0(.douta(w_n5110_0[0]),.doutb(w_dff_A_B735v1Ea2_1),.din(n5110));
	jspl3 jspl3_w_n5112_0(.douta(w_n5112_0[0]),.doutb(w_n5112_0[1]),.doutc(w_n5112_0[2]),.din(n5112));
	jspl3 jspl3_w_n5113_0(.douta(w_n5113_0[0]),.doutb(w_n5113_0[1]),.doutc(w_n5113_0[2]),.din(n5113));
	jspl jspl_w_n5116_0(.douta(w_n5116_0[0]),.doutb(w_n5116_0[1]),.din(n5116));
	jspl jspl_w_n5117_0(.douta(w_n5117_0[0]),.doutb(w_n5117_0[1]),.din(n5117));
	jspl jspl_w_n5118_0(.douta(w_n5118_0[0]),.doutb(w_n5118_0[1]),.din(n5118));
	jspl3 jspl3_w_n5119_0(.douta(w_n5119_0[0]),.doutb(w_n5119_0[1]),.doutc(w_n5119_0[2]),.din(n5119));
	jspl jspl_w_n5120_0(.douta(w_n5120_0[0]),.doutb(w_dff_A_lr3QEvLc2_1),.din(w_dff_B_QvlyzZXy5_2));
	jspl jspl_w_n5123_0(.douta(w_n5123_0[0]),.doutb(w_n5123_0[1]),.din(n5123));
	jspl jspl_w_n5126_0(.douta(w_n5126_0[0]),.doutb(w_n5126_0[1]),.din(n5126));
	jspl jspl_w_n5128_0(.douta(w_n5128_0[0]),.doutb(w_n5128_0[1]),.din(n5128));
	jspl jspl_w_n5129_0(.douta(w_n5129_0[0]),.doutb(w_n5129_0[1]),.din(n5129));
	jspl jspl_w_n5130_0(.douta(w_n5130_0[0]),.doutb(w_n5130_0[1]),.din(n5130));
	jspl jspl_w_n5132_0(.douta(w_n5132_0[0]),.doutb(w_n5132_0[1]),.din(n5132));
	jspl jspl_w_n5133_0(.douta(w_n5133_0[0]),.doutb(w_dff_A_OaMuw6Hb9_1),.din(n5133));
	jspl jspl_w_n5137_0(.douta(w_n5137_0[0]),.doutb(w_dff_A_N6sxVGld7_1),.din(w_dff_B_389mS7mG7_2));
	jspl jspl_w_n5138_0(.douta(w_n5138_0[0]),.doutb(w_n5138_0[1]),.din(n5138));
	jspl jspl_w_n5140_0(.douta(w_n5140_0[0]),.doutb(w_dff_A_WhFlsVOj3_1),.din(n5140));
	jspl jspl_w_n5142_0(.douta(w_n5142_0[0]),.doutb(w_n5142_0[1]),.din(n5142));
	jdff dff_A_RiPtSZDk9_1(.dout(w_n4014_0[1]),.din(w_dff_A_RiPtSZDk9_1),.clk(gclk));
	jdff dff_A_NGXHeKO55_0(.dout(w_n4013_10[0]),.din(w_dff_A_NGXHeKO55_0),.clk(gclk));
	jdff dff_A_37IA4n3O4_0(.dout(w_dff_A_NGXHeKO55_0),.din(w_dff_A_37IA4n3O4_0),.clk(gclk));
	jdff dff_A_4OtQlOja2_0(.dout(w_dff_A_37IA4n3O4_0),.din(w_dff_A_4OtQlOja2_0),.clk(gclk));
	jdff dff_A_TpbVPwI53_0(.dout(w_dff_A_4OtQlOja2_0),.din(w_dff_A_TpbVPwI53_0),.clk(gclk));
	jdff dff_A_kpphw58F3_0(.dout(w_dff_A_TpbVPwI53_0),.din(w_dff_A_kpphw58F3_0),.clk(gclk));
	jdff dff_A_vlPZ0Ent8_1(.dout(w_n4013_10[1]),.din(w_dff_A_vlPZ0Ent8_1),.clk(gclk));
	jdff dff_A_UoKBhK4Y5_1(.dout(w_dff_A_vlPZ0Ent8_1),.din(w_dff_A_UoKBhK4Y5_1),.clk(gclk));
	jdff dff_A_Hx1Ouz7H2_1(.dout(w_dff_A_UoKBhK4Y5_1),.din(w_dff_A_Hx1Ouz7H2_1),.clk(gclk));
	jdff dff_A_MZ7mXmkf2_0(.dout(w_n4013_9[0]),.din(w_dff_A_MZ7mXmkf2_0),.clk(gclk));
	jdff dff_A_sF759xAa4_0(.dout(w_dff_A_MZ7mXmkf2_0),.din(w_dff_A_sF759xAa4_0),.clk(gclk));
	jdff dff_A_gKWP81xO2_0(.dout(w_dff_A_sF759xAa4_0),.din(w_dff_A_gKWP81xO2_0),.clk(gclk));
	jdff dff_A_s4kVgoWW2_0(.dout(w_dff_A_gKWP81xO2_0),.din(w_dff_A_s4kVgoWW2_0),.clk(gclk));
	jdff dff_A_71ea6gqc1_1(.dout(w_n4013_9[1]),.din(w_dff_A_71ea6gqc1_1),.clk(gclk));
	jdff dff_A_ucqtqfZU9_1(.dout(w_dff_A_71ea6gqc1_1),.din(w_dff_A_ucqtqfZU9_1),.clk(gclk));
	jdff dff_A_z1uSxqiA1_0(.dout(w_n4013_8[0]),.din(w_dff_A_z1uSxqiA1_0),.clk(gclk));
	jdff dff_A_5FLG8NpT4_0(.dout(w_dff_A_z1uSxqiA1_0),.din(w_dff_A_5FLG8NpT4_0),.clk(gclk));
	jdff dff_A_PyH5QJbQ1_0(.dout(w_dff_A_5FLG8NpT4_0),.din(w_dff_A_PyH5QJbQ1_0),.clk(gclk));
	jdff dff_A_VEC9hgaD8_0(.dout(w_dff_A_PyH5QJbQ1_0),.din(w_dff_A_VEC9hgaD8_0),.clk(gclk));
	jdff dff_A_VBobKaBi6_1(.dout(w_n4013_8[1]),.din(w_dff_A_VBobKaBi6_1),.clk(gclk));
	jdff dff_A_TV7kAWfk8_1(.dout(w_dff_A_VBobKaBi6_1),.din(w_dff_A_TV7kAWfk8_1),.clk(gclk));
	jdff dff_A_GJdWBh692_0(.dout(w_n4013_7[0]),.din(w_dff_A_GJdWBh692_0),.clk(gclk));
	jdff dff_A_kVOWvjKY5_0(.dout(w_dff_A_GJdWBh692_0),.din(w_dff_A_kVOWvjKY5_0),.clk(gclk));
	jdff dff_A_aOryP3WK4_0(.dout(w_dff_A_kVOWvjKY5_0),.din(w_dff_A_aOryP3WK4_0),.clk(gclk));
	jdff dff_A_GJdM5i5M9_0(.dout(w_dff_A_aOryP3WK4_0),.din(w_dff_A_GJdM5i5M9_0),.clk(gclk));
	jdff dff_A_wQjDLugB6_1(.dout(w_n4013_7[1]),.din(w_dff_A_wQjDLugB6_1),.clk(gclk));
	jdff dff_A_hKKpVgtY8_1(.dout(w_dff_A_wQjDLugB6_1),.din(w_dff_A_hKKpVgtY8_1),.clk(gclk));
	jdff dff_A_GbhPl4H60_0(.dout(w_n4013_2[0]),.din(w_dff_A_GbhPl4H60_0),.clk(gclk));
	jdff dff_A_HxOgasBy2_0(.dout(w_dff_A_GbhPl4H60_0),.din(w_dff_A_HxOgasBy2_0),.clk(gclk));
	jdff dff_A_B0Y8cdCP8_0(.dout(w_dff_A_HxOgasBy2_0),.din(w_dff_A_B0Y8cdCP8_0),.clk(gclk));
	jdff dff_A_pLKYVyp88_0(.dout(w_dff_A_B0Y8cdCP8_0),.din(w_dff_A_pLKYVyp88_0),.clk(gclk));
	jdff dff_A_EkEHmc8d2_0(.dout(w_dff_A_pLKYVyp88_0),.din(w_dff_A_EkEHmc8d2_0),.clk(gclk));
	jdff dff_A_LkUnTVjy1_0(.dout(w_dff_A_EkEHmc8d2_0),.din(w_dff_A_LkUnTVjy1_0),.clk(gclk));
	jdff dff_A_a1aj6vRM7_0(.dout(w_dff_A_LkUnTVjy1_0),.din(w_dff_A_a1aj6vRM7_0),.clk(gclk));
	jdff dff_A_pZnZyIvF9_0(.dout(w_dff_A_a1aj6vRM7_0),.din(w_dff_A_pZnZyIvF9_0),.clk(gclk));
	jdff dff_A_9hCSOo2w9_0(.dout(w_dff_A_pZnZyIvF9_0),.din(w_dff_A_9hCSOo2w9_0),.clk(gclk));
	jdff dff_A_ZsQ6Rmqk2_0(.dout(w_dff_A_9hCSOo2w9_0),.din(w_dff_A_ZsQ6Rmqk2_0),.clk(gclk));
	jdff dff_A_IUPVafqv2_0(.dout(w_dff_A_ZsQ6Rmqk2_0),.din(w_dff_A_IUPVafqv2_0),.clk(gclk));
	jdff dff_A_zFz06Ms96_0(.dout(w_dff_A_IUPVafqv2_0),.din(w_dff_A_zFz06Ms96_0),.clk(gclk));
	jdff dff_A_c1FXsuoM0_1(.dout(w_n4013_2[1]),.din(w_dff_A_c1FXsuoM0_1),.clk(gclk));
	jdff dff_A_s4A9eYcR0_1(.dout(w_dff_A_c1FXsuoM0_1),.din(w_dff_A_s4A9eYcR0_1),.clk(gclk));
	jdff dff_A_QopHYMRW9_1(.dout(w_dff_A_s4A9eYcR0_1),.din(w_dff_A_QopHYMRW9_1),.clk(gclk));
	jdff dff_A_h7oPp7wq6_1(.dout(w_dff_A_QopHYMRW9_1),.din(w_dff_A_h7oPp7wq6_1),.clk(gclk));
	jdff dff_A_ApGqMT1D4_1(.dout(w_dff_A_h7oPp7wq6_1),.din(w_dff_A_ApGqMT1D4_1),.clk(gclk));
	jdff dff_A_bJB9Q22H3_1(.dout(w_dff_A_ApGqMT1D4_1),.din(w_dff_A_bJB9Q22H3_1),.clk(gclk));
	jdff dff_A_rbEHx83I3_0(.dout(w_n4013_6[0]),.din(w_dff_A_rbEHx83I3_0),.clk(gclk));
	jdff dff_A_DgJBwDXc8_0(.dout(w_dff_A_rbEHx83I3_0),.din(w_dff_A_DgJBwDXc8_0),.clk(gclk));
	jdff dff_A_EtaMr0GE0_0(.dout(w_dff_A_DgJBwDXc8_0),.din(w_dff_A_EtaMr0GE0_0),.clk(gclk));
	jdff dff_A_wMefoSvl1_0(.dout(w_dff_A_EtaMr0GE0_0),.din(w_dff_A_wMefoSvl1_0),.clk(gclk));
	jdff dff_A_uAUH7fgJ9_1(.dout(w_n4013_6[1]),.din(w_dff_A_uAUH7fgJ9_1),.clk(gclk));
	jdff dff_A_dBDyGrTJ0_1(.dout(w_dff_A_uAUH7fgJ9_1),.din(w_dff_A_dBDyGrTJ0_1),.clk(gclk));
	jdff dff_B_eZEzychJ4_0(.din(n5022),.dout(w_dff_B_eZEzychJ4_0),.clk(gclk));
	jdff dff_A_RBDOLeeS2_0(.dout(w_n5046_0[0]),.din(w_dff_A_RBDOLeeS2_0),.clk(gclk));
	jdff dff_A_m2X92ovI5_0(.dout(w_dff_A_RBDOLeeS2_0),.din(w_dff_A_m2X92ovI5_0),.clk(gclk));
	jdff dff_A_bZ09vicW3_0(.dout(w_dff_A_m2X92ovI5_0),.din(w_dff_A_bZ09vicW3_0),.clk(gclk));
	jdff dff_B_5RI4xp2g0_2(.din(n5046),.dout(w_dff_B_5RI4xp2g0_2),.clk(gclk));
	jdff dff_B_dhiVQU502_2(.din(w_dff_B_5RI4xp2g0_2),.dout(w_dff_B_dhiVQU502_2),.clk(gclk));
	jdff dff_B_jcaxrZF74_2(.din(w_dff_B_dhiVQU502_2),.dout(w_dff_B_jcaxrZF74_2),.clk(gclk));
	jdff dff_B_w3sdJIzj0_2(.din(w_dff_B_jcaxrZF74_2),.dout(w_dff_B_w3sdJIzj0_2),.clk(gclk));
	jdff dff_B_BAThx7lY3_2(.din(w_dff_B_w3sdJIzj0_2),.dout(w_dff_B_BAThx7lY3_2),.clk(gclk));
	jdff dff_B_riTWdShy8_2(.din(w_dff_B_BAThx7lY3_2),.dout(w_dff_B_riTWdShy8_2),.clk(gclk));
	jdff dff_B_ULl67ORI8_2(.din(w_dff_B_riTWdShy8_2),.dout(w_dff_B_ULl67ORI8_2),.clk(gclk));
	jdff dff_B_MXVV6Kuo8_2(.din(w_dff_B_ULl67ORI8_2),.dout(w_dff_B_MXVV6Kuo8_2),.clk(gclk));
	jdff dff_B_yGx9f0w05_2(.din(w_dff_B_MXVV6Kuo8_2),.dout(w_dff_B_yGx9f0w05_2),.clk(gclk));
	jdff dff_B_Qr16cTJg6_2(.din(w_dff_B_yGx9f0w05_2),.dout(w_dff_B_Qr16cTJg6_2),.clk(gclk));
	jdff dff_B_mCu6o7Is6_2(.din(w_dff_B_Qr16cTJg6_2),.dout(w_dff_B_mCu6o7Is6_2),.clk(gclk));
	jdff dff_B_YLo8Csg21_2(.din(w_dff_B_mCu6o7Is6_2),.dout(w_dff_B_YLo8Csg21_2),.clk(gclk));
	jdff dff_B_VK4p86qM3_2(.din(w_dff_B_YLo8Csg21_2),.dout(w_dff_B_VK4p86qM3_2),.clk(gclk));
	jdff dff_B_sWi4cVC18_2(.din(w_dff_B_VK4p86qM3_2),.dout(w_dff_B_sWi4cVC18_2),.clk(gclk));
	jdff dff_B_XwE082Vg1_2(.din(w_dff_B_sWi4cVC18_2),.dout(w_dff_B_XwE082Vg1_2),.clk(gclk));
	jdff dff_B_Eu7QGMNU6_2(.din(w_dff_B_XwE082Vg1_2),.dout(w_dff_B_Eu7QGMNU6_2),.clk(gclk));
	jdff dff_B_icLouTRe3_2(.din(w_dff_B_Eu7QGMNU6_2),.dout(w_dff_B_icLouTRe3_2),.clk(gclk));
	jdff dff_B_JCU59h5a4_2(.din(w_dff_B_icLouTRe3_2),.dout(w_dff_B_JCU59h5a4_2),.clk(gclk));
	jdff dff_B_jlC6hA1j8_2(.din(w_dff_B_JCU59h5a4_2),.dout(w_dff_B_jlC6hA1j8_2),.clk(gclk));
	jdff dff_B_cBNuyFzy2_2(.din(w_dff_B_jlC6hA1j8_2),.dout(w_dff_B_cBNuyFzy2_2),.clk(gclk));
	jdff dff_B_Y9FVxNhB9_2(.din(w_dff_B_cBNuyFzy2_2),.dout(w_dff_B_Y9FVxNhB9_2),.clk(gclk));
	jdff dff_B_o6QWkKQA0_2(.din(w_dff_B_Y9FVxNhB9_2),.dout(w_dff_B_o6QWkKQA0_2),.clk(gclk));
	jdff dff_B_EydgXy3w4_2(.din(w_dff_B_o6QWkKQA0_2),.dout(w_dff_B_EydgXy3w4_2),.clk(gclk));
	jdff dff_B_m3IjCvmS5_2(.din(w_dff_B_EydgXy3w4_2),.dout(w_dff_B_m3IjCvmS5_2),.clk(gclk));
	jdff dff_B_jup1g00q9_2(.din(w_dff_B_m3IjCvmS5_2),.dout(w_dff_B_jup1g00q9_2),.clk(gclk));
	jdff dff_B_PUkG8ZRw4_2(.din(w_dff_B_jup1g00q9_2),.dout(w_dff_B_PUkG8ZRw4_2),.clk(gclk));
	jdff dff_B_wgMSX9l29_2(.din(w_dff_B_PUkG8ZRw4_2),.dout(w_dff_B_wgMSX9l29_2),.clk(gclk));
	jdff dff_B_A71ehwnI3_2(.din(w_dff_B_wgMSX9l29_2),.dout(w_dff_B_A71ehwnI3_2),.clk(gclk));
	jdff dff_B_XZV6JPhW1_2(.din(w_dff_B_A71ehwnI3_2),.dout(w_dff_B_XZV6JPhW1_2),.clk(gclk));
	jdff dff_B_qlKAxEia2_2(.din(w_dff_B_XZV6JPhW1_2),.dout(w_dff_B_qlKAxEia2_2),.clk(gclk));
	jdff dff_B_gvL5aKzK1_2(.din(w_dff_B_qlKAxEia2_2),.dout(w_dff_B_gvL5aKzK1_2),.clk(gclk));
	jdff dff_B_CsliOohJ7_2(.din(w_dff_B_gvL5aKzK1_2),.dout(w_dff_B_CsliOohJ7_2),.clk(gclk));
	jdff dff_B_G6YBppBM0_2(.din(w_dff_B_CsliOohJ7_2),.dout(w_dff_B_G6YBppBM0_2),.clk(gclk));
	jdff dff_B_ZzJf2LJC4_2(.din(w_dff_B_G6YBppBM0_2),.dout(w_dff_B_ZzJf2LJC4_2),.clk(gclk));
	jdff dff_B_WEHirB0f9_2(.din(w_dff_B_ZzJf2LJC4_2),.dout(w_dff_B_WEHirB0f9_2),.clk(gclk));
	jdff dff_B_OzwR54au9_2(.din(w_dff_B_WEHirB0f9_2),.dout(w_dff_B_OzwR54au9_2),.clk(gclk));
	jdff dff_B_Exl1FNYz6_2(.din(w_dff_B_OzwR54au9_2),.dout(w_dff_B_Exl1FNYz6_2),.clk(gclk));
	jdff dff_B_9k2eQFIa7_2(.din(w_dff_B_Exl1FNYz6_2),.dout(w_dff_B_9k2eQFIa7_2),.clk(gclk));
	jdff dff_B_2VstCvap2_2(.din(w_dff_B_9k2eQFIa7_2),.dout(w_dff_B_2VstCvap2_2),.clk(gclk));
	jdff dff_B_uBVkdo3C0_2(.din(w_dff_B_2VstCvap2_2),.dout(w_dff_B_uBVkdo3C0_2),.clk(gclk));
	jdff dff_B_s1VBUl6w1_2(.din(w_dff_B_uBVkdo3C0_2),.dout(w_dff_B_s1VBUl6w1_2),.clk(gclk));
	jdff dff_B_Qa9YHEfh9_2(.din(w_dff_B_s1VBUl6w1_2),.dout(w_dff_B_Qa9YHEfh9_2),.clk(gclk));
	jdff dff_B_MgMvnRTs0_2(.din(w_dff_B_Qa9YHEfh9_2),.dout(w_dff_B_MgMvnRTs0_2),.clk(gclk));
	jdff dff_B_Vg5ZcwMW4_2(.din(w_dff_B_MgMvnRTs0_2),.dout(w_dff_B_Vg5ZcwMW4_2),.clk(gclk));
	jdff dff_B_GK3MlLa02_2(.din(w_dff_B_Vg5ZcwMW4_2),.dout(w_dff_B_GK3MlLa02_2),.clk(gclk));
	jdff dff_B_3J0Az0Tj9_2(.din(w_dff_B_GK3MlLa02_2),.dout(w_dff_B_3J0Az0Tj9_2),.clk(gclk));
	jdff dff_B_iJMDOdGD0_2(.din(w_dff_B_3J0Az0Tj9_2),.dout(w_dff_B_iJMDOdGD0_2),.clk(gclk));
	jdff dff_B_3Y6m6eYG7_2(.din(w_dff_B_iJMDOdGD0_2),.dout(w_dff_B_3Y6m6eYG7_2),.clk(gclk));
	jdff dff_B_5kGmypLt0_2(.din(w_dff_B_3Y6m6eYG7_2),.dout(w_dff_B_5kGmypLt0_2),.clk(gclk));
	jdff dff_B_bmvoXJ8M9_2(.din(w_dff_B_5kGmypLt0_2),.dout(w_dff_B_bmvoXJ8M9_2),.clk(gclk));
	jdff dff_B_NQNAA8pr0_2(.din(w_dff_B_bmvoXJ8M9_2),.dout(w_dff_B_NQNAA8pr0_2),.clk(gclk));
	jdff dff_B_vxJaR31t8_2(.din(w_dff_B_NQNAA8pr0_2),.dout(w_dff_B_vxJaR31t8_2),.clk(gclk));
	jdff dff_B_Wxo4ZPjh9_2(.din(w_dff_B_vxJaR31t8_2),.dout(w_dff_B_Wxo4ZPjh9_2),.clk(gclk));
	jdff dff_B_rj1wjVlq7_2(.din(w_dff_B_Wxo4ZPjh9_2),.dout(w_dff_B_rj1wjVlq7_2),.clk(gclk));
	jdff dff_B_ZR1DnZ4i9_2(.din(w_dff_B_rj1wjVlq7_2),.dout(w_dff_B_ZR1DnZ4i9_2),.clk(gclk));
	jdff dff_B_OCgBxrtb4_2(.din(w_dff_B_ZR1DnZ4i9_2),.dout(w_dff_B_OCgBxrtb4_2),.clk(gclk));
	jdff dff_B_X9TYsqmO2_2(.din(w_dff_B_OCgBxrtb4_2),.dout(w_dff_B_X9TYsqmO2_2),.clk(gclk));
	jdff dff_B_ottB5zyD7_2(.din(w_dff_B_X9TYsqmO2_2),.dout(w_dff_B_ottB5zyD7_2),.clk(gclk));
	jdff dff_B_eWTgTqtM5_2(.din(w_dff_B_ottB5zyD7_2),.dout(w_dff_B_eWTgTqtM5_2),.clk(gclk));
	jdff dff_B_pTRErxPb5_2(.din(w_dff_B_eWTgTqtM5_2),.dout(w_dff_B_pTRErxPb5_2),.clk(gclk));
	jdff dff_B_Milp0czy0_2(.din(w_dff_B_pTRErxPb5_2),.dout(w_dff_B_Milp0czy0_2),.clk(gclk));
	jdff dff_B_7yseujS22_2(.din(w_dff_B_Milp0czy0_2),.dout(w_dff_B_7yseujS22_2),.clk(gclk));
	jdff dff_B_sw3dxI9g4_2(.din(w_dff_B_7yseujS22_2),.dout(w_dff_B_sw3dxI9g4_2),.clk(gclk));
	jdff dff_B_fz22z2qR1_2(.din(w_dff_B_sw3dxI9g4_2),.dout(w_dff_B_fz22z2qR1_2),.clk(gclk));
	jdff dff_B_Gt05YMW87_2(.din(w_dff_B_fz22z2qR1_2),.dout(w_dff_B_Gt05YMW87_2),.clk(gclk));
	jdff dff_B_HEL5L0zz2_2(.din(w_dff_B_Gt05YMW87_2),.dout(w_dff_B_HEL5L0zz2_2),.clk(gclk));
	jdff dff_B_TMjOVxqT5_2(.din(w_dff_B_HEL5L0zz2_2),.dout(w_dff_B_TMjOVxqT5_2),.clk(gclk));
	jdff dff_B_KcW4lYA00_2(.din(w_dff_B_TMjOVxqT5_2),.dout(w_dff_B_KcW4lYA00_2),.clk(gclk));
	jdff dff_B_fuyAr6Pq3_2(.din(w_dff_B_KcW4lYA00_2),.dout(w_dff_B_fuyAr6Pq3_2),.clk(gclk));
	jdff dff_B_44woTVgy3_2(.din(w_dff_B_fuyAr6Pq3_2),.dout(w_dff_B_44woTVgy3_2),.clk(gclk));
	jdff dff_B_KDKBNM6v0_2(.din(w_dff_B_44woTVgy3_2),.dout(w_dff_B_KDKBNM6v0_2),.clk(gclk));
	jdff dff_B_1E3aRSXX0_2(.din(w_dff_B_KDKBNM6v0_2),.dout(w_dff_B_1E3aRSXX0_2),.clk(gclk));
	jdff dff_B_TISKl5955_2(.din(w_dff_B_1E3aRSXX0_2),.dout(w_dff_B_TISKl5955_2),.clk(gclk));
	jdff dff_B_Jyxz7DFM1_2(.din(w_dff_B_TISKl5955_2),.dout(w_dff_B_Jyxz7DFM1_2),.clk(gclk));
	jdff dff_B_3sRop2Ie6_2(.din(w_dff_B_Jyxz7DFM1_2),.dout(w_dff_B_3sRop2Ie6_2),.clk(gclk));
	jdff dff_B_y7ccUvVH1_2(.din(w_dff_B_3sRop2Ie6_2),.dout(w_dff_B_y7ccUvVH1_2),.clk(gclk));
	jdff dff_B_UFNe7O7N9_2(.din(w_dff_B_y7ccUvVH1_2),.dout(w_dff_B_UFNe7O7N9_2),.clk(gclk));
	jdff dff_B_NJFkvd9n3_2(.din(w_dff_B_UFNe7O7N9_2),.dout(w_dff_B_NJFkvd9n3_2),.clk(gclk));
	jdff dff_B_O9A2viQI7_2(.din(w_dff_B_NJFkvd9n3_2),.dout(w_dff_B_O9A2viQI7_2),.clk(gclk));
	jdff dff_B_OhJT1iyq9_2(.din(w_dff_B_O9A2viQI7_2),.dout(w_dff_B_OhJT1iyq9_2),.clk(gclk));
	jdff dff_B_FaBiW03U2_2(.din(w_dff_B_OhJT1iyq9_2),.dout(w_dff_B_FaBiW03U2_2),.clk(gclk));
	jdff dff_B_5j6zucTg2_2(.din(w_dff_B_FaBiW03U2_2),.dout(w_dff_B_5j6zucTg2_2),.clk(gclk));
	jdff dff_B_i20OsPjB8_2(.din(w_dff_B_5j6zucTg2_2),.dout(w_dff_B_i20OsPjB8_2),.clk(gclk));
	jdff dff_B_Rs7NWEAE4_2(.din(w_dff_B_i20OsPjB8_2),.dout(w_dff_B_Rs7NWEAE4_2),.clk(gclk));
	jdff dff_B_QP4PSIAd5_2(.din(w_dff_B_Rs7NWEAE4_2),.dout(w_dff_B_QP4PSIAd5_2),.clk(gclk));
	jdff dff_B_AftEnVhu8_2(.din(w_dff_B_QP4PSIAd5_2),.dout(w_dff_B_AftEnVhu8_2),.clk(gclk));
	jdff dff_B_AM5Bs5ur0_2(.din(w_dff_B_AftEnVhu8_2),.dout(w_dff_B_AM5Bs5ur0_2),.clk(gclk));
	jdff dff_B_TmSKnfvk0_2(.din(w_dff_B_AM5Bs5ur0_2),.dout(w_dff_B_TmSKnfvk0_2),.clk(gclk));
	jdff dff_B_Le8JZY4E5_2(.din(w_dff_B_TmSKnfvk0_2),.dout(w_dff_B_Le8JZY4E5_2),.clk(gclk));
	jdff dff_B_PLHNxj171_2(.din(w_dff_B_Le8JZY4E5_2),.dout(w_dff_B_PLHNxj171_2),.clk(gclk));
	jdff dff_B_fkiWHb5z7_2(.din(w_dff_B_PLHNxj171_2),.dout(w_dff_B_fkiWHb5z7_2),.clk(gclk));
	jdff dff_B_wsJydkto0_2(.din(w_dff_B_fkiWHb5z7_2),.dout(w_dff_B_wsJydkto0_2),.clk(gclk));
	jdff dff_B_9cKC052I7_2(.din(w_dff_B_wsJydkto0_2),.dout(w_dff_B_9cKC052I7_2),.clk(gclk));
	jdff dff_B_KOsJ800c0_2(.din(w_dff_B_9cKC052I7_2),.dout(w_dff_B_KOsJ800c0_2),.clk(gclk));
	jdff dff_B_SufTqADf2_2(.din(w_dff_B_KOsJ800c0_2),.dout(w_dff_B_SufTqADf2_2),.clk(gclk));
	jdff dff_B_ETFt5nf87_2(.din(w_dff_B_SufTqADf2_2),.dout(w_dff_B_ETFt5nf87_2),.clk(gclk));
	jdff dff_B_q5szTSDk8_2(.din(w_dff_B_ETFt5nf87_2),.dout(w_dff_B_q5szTSDk8_2),.clk(gclk));
	jdff dff_B_awuJZjRy1_2(.din(w_dff_B_q5szTSDk8_2),.dout(w_dff_B_awuJZjRy1_2),.clk(gclk));
	jdff dff_B_NaRMWG1q4_2(.din(w_dff_B_awuJZjRy1_2),.dout(w_dff_B_NaRMWG1q4_2),.clk(gclk));
	jdff dff_B_houcbZNh6_2(.din(w_dff_B_NaRMWG1q4_2),.dout(w_dff_B_houcbZNh6_2),.clk(gclk));
	jdff dff_B_pcKV86BE1_2(.din(w_dff_B_houcbZNh6_2),.dout(w_dff_B_pcKV86BE1_2),.clk(gclk));
	jdff dff_B_AzKsezPA4_2(.din(w_dff_B_pcKV86BE1_2),.dout(w_dff_B_AzKsezPA4_2),.clk(gclk));
	jdff dff_B_vxaNRlZp0_2(.din(w_dff_B_AzKsezPA4_2),.dout(w_dff_B_vxaNRlZp0_2),.clk(gclk));
	jdff dff_B_yiPpV30k0_2(.din(w_dff_B_vxaNRlZp0_2),.dout(w_dff_B_yiPpV30k0_2),.clk(gclk));
	jdff dff_B_8qirCfdf9_2(.din(w_dff_B_yiPpV30k0_2),.dout(w_dff_B_8qirCfdf9_2),.clk(gclk));
	jdff dff_B_vQ1IGsp82_2(.din(w_dff_B_8qirCfdf9_2),.dout(w_dff_B_vQ1IGsp82_2),.clk(gclk));
	jdff dff_B_LAmnM0vh0_2(.din(w_dff_B_vQ1IGsp82_2),.dout(w_dff_B_LAmnM0vh0_2),.clk(gclk));
	jdff dff_B_FUdmWInD1_2(.din(w_dff_B_LAmnM0vh0_2),.dout(w_dff_B_FUdmWInD1_2),.clk(gclk));
	jdff dff_B_Ryt8C1hJ5_2(.din(w_dff_B_FUdmWInD1_2),.dout(w_dff_B_Ryt8C1hJ5_2),.clk(gclk));
	jdff dff_B_VYJQqXnf0_2(.din(w_dff_B_Ryt8C1hJ5_2),.dout(w_dff_B_VYJQqXnf0_2),.clk(gclk));
	jdff dff_B_LxKP9G961_2(.din(w_dff_B_VYJQqXnf0_2),.dout(w_dff_B_LxKP9G961_2),.clk(gclk));
	jdff dff_B_PigctOHU8_2(.din(w_dff_B_LxKP9G961_2),.dout(w_dff_B_PigctOHU8_2),.clk(gclk));
	jdff dff_B_MH55XeHM6_2(.din(w_dff_B_PigctOHU8_2),.dout(w_dff_B_MH55XeHM6_2),.clk(gclk));
	jdff dff_B_yHPASRXz5_2(.din(w_dff_B_MH55XeHM6_2),.dout(w_dff_B_yHPASRXz5_2),.clk(gclk));
	jdff dff_B_0LaGRlav8_2(.din(w_dff_B_yHPASRXz5_2),.dout(w_dff_B_0LaGRlav8_2),.clk(gclk));
	jdff dff_B_6mfeIp3z0_2(.din(w_dff_B_0LaGRlav8_2),.dout(w_dff_B_6mfeIp3z0_2),.clk(gclk));
	jdff dff_B_yD7dkkhi9_2(.din(w_dff_B_6mfeIp3z0_2),.dout(w_dff_B_yD7dkkhi9_2),.clk(gclk));
	jdff dff_B_LQiHz9fy5_2(.din(w_dff_B_yD7dkkhi9_2),.dout(w_dff_B_LQiHz9fy5_2),.clk(gclk));
	jdff dff_B_uEyTSu8O3_2(.din(w_dff_B_LQiHz9fy5_2),.dout(w_dff_B_uEyTSu8O3_2),.clk(gclk));
	jdff dff_B_cHfGK3wW5_2(.din(w_dff_B_uEyTSu8O3_2),.dout(w_dff_B_cHfGK3wW5_2),.clk(gclk));
	jdff dff_B_KjLceTJ15_2(.din(w_dff_B_cHfGK3wW5_2),.dout(w_dff_B_KjLceTJ15_2),.clk(gclk));
	jdff dff_B_Fx4HYKGK9_2(.din(w_dff_B_KjLceTJ15_2),.dout(w_dff_B_Fx4HYKGK9_2),.clk(gclk));
	jdff dff_B_QcR9J9D45_2(.din(w_dff_B_Fx4HYKGK9_2),.dout(w_dff_B_QcR9J9D45_2),.clk(gclk));
	jdff dff_B_CWSG3c6X3_2(.din(w_dff_B_QcR9J9D45_2),.dout(w_dff_B_CWSG3c6X3_2),.clk(gclk));
	jdff dff_B_FYi19mux6_2(.din(w_dff_B_CWSG3c6X3_2),.dout(w_dff_B_FYi19mux6_2),.clk(gclk));
	jdff dff_B_UGfytwYE5_2(.din(w_dff_B_FYi19mux6_2),.dout(w_dff_B_UGfytwYE5_2),.clk(gclk));
	jdff dff_B_fTmfuLci5_2(.din(w_dff_B_UGfytwYE5_2),.dout(w_dff_B_fTmfuLci5_2),.clk(gclk));
	jdff dff_B_wgwNlq0s6_2(.din(w_dff_B_fTmfuLci5_2),.dout(w_dff_B_wgwNlq0s6_2),.clk(gclk));
	jdff dff_B_B9hxklVT5_2(.din(w_dff_B_wgwNlq0s6_2),.dout(w_dff_B_B9hxklVT5_2),.clk(gclk));
	jdff dff_B_H1CEOAzK2_2(.din(w_dff_B_B9hxklVT5_2),.dout(w_dff_B_H1CEOAzK2_2),.clk(gclk));
	jdff dff_B_yQCmSbu72_2(.din(w_dff_B_H1CEOAzK2_2),.dout(w_dff_B_yQCmSbu72_2),.clk(gclk));
	jdff dff_B_xkNf9owQ5_2(.din(w_dff_B_yQCmSbu72_2),.dout(w_dff_B_xkNf9owQ5_2),.clk(gclk));
	jdff dff_B_PNEGI4yT5_2(.din(w_dff_B_xkNf9owQ5_2),.dout(w_dff_B_PNEGI4yT5_2),.clk(gclk));
	jdff dff_B_fJ7zhDrm9_2(.din(w_dff_B_PNEGI4yT5_2),.dout(w_dff_B_fJ7zhDrm9_2),.clk(gclk));
	jdff dff_B_46lDhABu1_2(.din(w_dff_B_fJ7zhDrm9_2),.dout(w_dff_B_46lDhABu1_2),.clk(gclk));
	jdff dff_B_qgr76Lbj5_2(.din(w_dff_B_46lDhABu1_2),.dout(w_dff_B_qgr76Lbj5_2),.clk(gclk));
	jdff dff_B_1a890rbd8_2(.din(w_dff_B_qgr76Lbj5_2),.dout(w_dff_B_1a890rbd8_2),.clk(gclk));
	jdff dff_B_YkOE5CkR1_2(.din(w_dff_B_1a890rbd8_2),.dout(w_dff_B_YkOE5CkR1_2),.clk(gclk));
	jdff dff_B_qL6rScVZ8_2(.din(w_dff_B_YkOE5CkR1_2),.dout(w_dff_B_qL6rScVZ8_2),.clk(gclk));
	jdff dff_B_4CHZKSur9_2(.din(w_dff_B_qL6rScVZ8_2),.dout(w_dff_B_4CHZKSur9_2),.clk(gclk));
	jdff dff_B_BeYRFeNT9_2(.din(w_dff_B_4CHZKSur9_2),.dout(w_dff_B_BeYRFeNT9_2),.clk(gclk));
	jdff dff_B_FEK6rsfi1_2(.din(w_dff_B_BeYRFeNT9_2),.dout(w_dff_B_FEK6rsfi1_2),.clk(gclk));
	jdff dff_B_0bWCEVVm3_2(.din(w_dff_B_FEK6rsfi1_2),.dout(w_dff_B_0bWCEVVm3_2),.clk(gclk));
	jdff dff_B_gd2Mccjr1_2(.din(w_dff_B_0bWCEVVm3_2),.dout(w_dff_B_gd2Mccjr1_2),.clk(gclk));
	jdff dff_B_vnp5ZE708_2(.din(w_dff_B_gd2Mccjr1_2),.dout(w_dff_B_vnp5ZE708_2),.clk(gclk));
	jdff dff_B_yCAK8FC23_2(.din(w_dff_B_vnp5ZE708_2),.dout(w_dff_B_yCAK8FC23_2),.clk(gclk));
	jdff dff_B_nPPCaf1Q4_2(.din(w_dff_B_yCAK8FC23_2),.dout(w_dff_B_nPPCaf1Q4_2),.clk(gclk));
	jdff dff_B_Gw348KKn2_2(.din(w_dff_B_nPPCaf1Q4_2),.dout(w_dff_B_Gw348KKn2_2),.clk(gclk));
	jdff dff_B_ysrD9GaZ8_2(.din(w_dff_B_Gw348KKn2_2),.dout(w_dff_B_ysrD9GaZ8_2),.clk(gclk));
	jdff dff_B_Zm7EjNgg7_2(.din(w_dff_B_ysrD9GaZ8_2),.dout(w_dff_B_Zm7EjNgg7_2),.clk(gclk));
	jdff dff_B_YYcRPf0b8_2(.din(w_dff_B_Zm7EjNgg7_2),.dout(w_dff_B_YYcRPf0b8_2),.clk(gclk));
	jdff dff_B_CtoyzuH37_2(.din(w_dff_B_YYcRPf0b8_2),.dout(w_dff_B_CtoyzuH37_2),.clk(gclk));
	jdff dff_B_1Q9Go4ez0_2(.din(w_dff_B_CtoyzuH37_2),.dout(w_dff_B_1Q9Go4ez0_2),.clk(gclk));
	jdff dff_B_iL8QFOMo9_2(.din(w_dff_B_1Q9Go4ez0_2),.dout(w_dff_B_iL8QFOMo9_2),.clk(gclk));
	jdff dff_B_5eDBnhxR4_2(.din(w_dff_B_iL8QFOMo9_2),.dout(w_dff_B_5eDBnhxR4_2),.clk(gclk));
	jdff dff_B_mIQBAR6E9_2(.din(w_dff_B_5eDBnhxR4_2),.dout(w_dff_B_mIQBAR6E9_2),.clk(gclk));
	jdff dff_B_wcw2K1gk7_2(.din(w_dff_B_mIQBAR6E9_2),.dout(w_dff_B_wcw2K1gk7_2),.clk(gclk));
	jdff dff_A_mEdyEIrL5_0(.dout(w_n4013_4[0]),.din(w_dff_A_mEdyEIrL5_0),.clk(gclk));
	jdff dff_A_Bw0aCnDm9_0(.dout(w_dff_A_mEdyEIrL5_0),.din(w_dff_A_Bw0aCnDm9_0),.clk(gclk));
	jdff dff_A_b6PhEX3p8_0(.dout(w_dff_A_Bw0aCnDm9_0),.din(w_dff_A_b6PhEX3p8_0),.clk(gclk));
	jdff dff_A_ypy0WxOY7_1(.dout(w_n4013_4[1]),.din(w_dff_A_ypy0WxOY7_1),.clk(gclk));
	jdff dff_A_QWOvLrxd2_1(.dout(w_dff_A_ypy0WxOY7_1),.din(w_dff_A_QWOvLrxd2_1),.clk(gclk));
	jdff dff_A_GY2RnPJc4_1(.dout(w_n5140_0[1]),.din(w_dff_A_GY2RnPJc4_1),.clk(gclk));
	jdff dff_A_WhFlsVOj3_1(.dout(w_dff_A_GY2RnPJc4_1),.din(w_dff_A_WhFlsVOj3_1),.clk(gclk));
	jdff dff_B_2rz4dWGZ7_1(.din(n5155),.dout(w_dff_B_2rz4dWGZ7_1),.clk(gclk));
	jdff dff_A_B735v1Ea2_1(.dout(w_n5110_0[1]),.din(w_dff_A_B735v1Ea2_1),.clk(gclk));
	jdff dff_B_OP6iqswc4_1(.din(n5093),.dout(w_dff_B_OP6iqswc4_1),.clk(gclk));
	jdff dff_A_h2PYpQyn7_0(.dout(w_n5050_0[0]),.din(w_dff_A_h2PYpQyn7_0),.clk(gclk));
	jdff dff_A_EohMCOr02_1(.dout(w_n5137_0[1]),.din(w_dff_A_EohMCOr02_1),.clk(gclk));
	jdff dff_A_N6sxVGld7_1(.dout(w_dff_A_EohMCOr02_1),.din(w_dff_A_N6sxVGld7_1),.clk(gclk));
	jdff dff_B_kKOZmqN48_2(.din(n5137),.dout(w_dff_B_kKOZmqN48_2),.clk(gclk));
	jdff dff_B_7rDoO9sx7_2(.din(w_dff_B_kKOZmqN48_2),.dout(w_dff_B_7rDoO9sx7_2),.clk(gclk));
	jdff dff_B_CeDtLGO62_2(.din(w_dff_B_7rDoO9sx7_2),.dout(w_dff_B_CeDtLGO62_2),.clk(gclk));
	jdff dff_B_DzGFTP3B4_2(.din(w_dff_B_CeDtLGO62_2),.dout(w_dff_B_DzGFTP3B4_2),.clk(gclk));
	jdff dff_B_g2D3wdph1_2(.din(w_dff_B_DzGFTP3B4_2),.dout(w_dff_B_g2D3wdph1_2),.clk(gclk));
	jdff dff_B_zcOhCS2a8_2(.din(w_dff_B_g2D3wdph1_2),.dout(w_dff_B_zcOhCS2a8_2),.clk(gclk));
	jdff dff_B_B8QSZ5Zm7_2(.din(w_dff_B_zcOhCS2a8_2),.dout(w_dff_B_B8QSZ5Zm7_2),.clk(gclk));
	jdff dff_B_yDTR2Y3x7_2(.din(w_dff_B_B8QSZ5Zm7_2),.dout(w_dff_B_yDTR2Y3x7_2),.clk(gclk));
	jdff dff_B_nlmpukMG7_2(.din(w_dff_B_yDTR2Y3x7_2),.dout(w_dff_B_nlmpukMG7_2),.clk(gclk));
	jdff dff_B_ANgszXzq4_2(.din(w_dff_B_nlmpukMG7_2),.dout(w_dff_B_ANgszXzq4_2),.clk(gclk));
	jdff dff_B_lKfhn1IJ8_2(.din(w_dff_B_ANgszXzq4_2),.dout(w_dff_B_lKfhn1IJ8_2),.clk(gclk));
	jdff dff_B_0TJPPYYb2_2(.din(w_dff_B_lKfhn1IJ8_2),.dout(w_dff_B_0TJPPYYb2_2),.clk(gclk));
	jdff dff_B_4uDgwDES3_2(.din(w_dff_B_0TJPPYYb2_2),.dout(w_dff_B_4uDgwDES3_2),.clk(gclk));
	jdff dff_B_KCex5Kn38_2(.din(w_dff_B_4uDgwDES3_2),.dout(w_dff_B_KCex5Kn38_2),.clk(gclk));
	jdff dff_B_8QGrpRFt9_2(.din(w_dff_B_KCex5Kn38_2),.dout(w_dff_B_8QGrpRFt9_2),.clk(gclk));
	jdff dff_B_PDW74LMp1_2(.din(w_dff_B_8QGrpRFt9_2),.dout(w_dff_B_PDW74LMp1_2),.clk(gclk));
	jdff dff_B_AJj62i627_2(.din(w_dff_B_PDW74LMp1_2),.dout(w_dff_B_AJj62i627_2),.clk(gclk));
	jdff dff_B_BIBiy4dV7_2(.din(w_dff_B_AJj62i627_2),.dout(w_dff_B_BIBiy4dV7_2),.clk(gclk));
	jdff dff_B_oRiamI7y5_2(.din(w_dff_B_BIBiy4dV7_2),.dout(w_dff_B_oRiamI7y5_2),.clk(gclk));
	jdff dff_B_Fudaf5rG0_2(.din(w_dff_B_oRiamI7y5_2),.dout(w_dff_B_Fudaf5rG0_2),.clk(gclk));
	jdff dff_B_7uJfallg2_2(.din(w_dff_B_Fudaf5rG0_2),.dout(w_dff_B_7uJfallg2_2),.clk(gclk));
	jdff dff_B_6RnCNS9P7_2(.din(w_dff_B_7uJfallg2_2),.dout(w_dff_B_6RnCNS9P7_2),.clk(gclk));
	jdff dff_B_HyMnj4nP1_2(.din(w_dff_B_6RnCNS9P7_2),.dout(w_dff_B_HyMnj4nP1_2),.clk(gclk));
	jdff dff_B_3XFrlSPU0_2(.din(w_dff_B_HyMnj4nP1_2),.dout(w_dff_B_3XFrlSPU0_2),.clk(gclk));
	jdff dff_B_r5j9ZkxA8_2(.din(w_dff_B_3XFrlSPU0_2),.dout(w_dff_B_r5j9ZkxA8_2),.clk(gclk));
	jdff dff_B_73cJfVwZ1_2(.din(w_dff_B_r5j9ZkxA8_2),.dout(w_dff_B_73cJfVwZ1_2),.clk(gclk));
	jdff dff_B_tyBm301x7_2(.din(w_dff_B_73cJfVwZ1_2),.dout(w_dff_B_tyBm301x7_2),.clk(gclk));
	jdff dff_B_xBaAXZT70_2(.din(w_dff_B_tyBm301x7_2),.dout(w_dff_B_xBaAXZT70_2),.clk(gclk));
	jdff dff_B_AuhgSYuF1_2(.din(w_dff_B_xBaAXZT70_2),.dout(w_dff_B_AuhgSYuF1_2),.clk(gclk));
	jdff dff_B_i6hB622j1_2(.din(w_dff_B_AuhgSYuF1_2),.dout(w_dff_B_i6hB622j1_2),.clk(gclk));
	jdff dff_B_o0qEQHwN2_2(.din(w_dff_B_i6hB622j1_2),.dout(w_dff_B_o0qEQHwN2_2),.clk(gclk));
	jdff dff_B_qpojBUg34_2(.din(w_dff_B_o0qEQHwN2_2),.dout(w_dff_B_qpojBUg34_2),.clk(gclk));
	jdff dff_B_v3nsYcVk8_2(.din(w_dff_B_qpojBUg34_2),.dout(w_dff_B_v3nsYcVk8_2),.clk(gclk));
	jdff dff_B_IL6YDOLP7_2(.din(w_dff_B_v3nsYcVk8_2),.dout(w_dff_B_IL6YDOLP7_2),.clk(gclk));
	jdff dff_B_W9idEL0R0_2(.din(w_dff_B_IL6YDOLP7_2),.dout(w_dff_B_W9idEL0R0_2),.clk(gclk));
	jdff dff_B_rwQv5M8l5_2(.din(w_dff_B_W9idEL0R0_2),.dout(w_dff_B_rwQv5M8l5_2),.clk(gclk));
	jdff dff_B_039ssV2g5_2(.din(w_dff_B_rwQv5M8l5_2),.dout(w_dff_B_039ssV2g5_2),.clk(gclk));
	jdff dff_B_2tKs1Km07_2(.din(w_dff_B_039ssV2g5_2),.dout(w_dff_B_2tKs1Km07_2),.clk(gclk));
	jdff dff_B_KjNMdo2c6_2(.din(w_dff_B_2tKs1Km07_2),.dout(w_dff_B_KjNMdo2c6_2),.clk(gclk));
	jdff dff_B_2JwdyTnF4_2(.din(w_dff_B_KjNMdo2c6_2),.dout(w_dff_B_2JwdyTnF4_2),.clk(gclk));
	jdff dff_B_83U5kNYX4_2(.din(w_dff_B_2JwdyTnF4_2),.dout(w_dff_B_83U5kNYX4_2),.clk(gclk));
	jdff dff_B_eRRRpXIp0_2(.din(w_dff_B_83U5kNYX4_2),.dout(w_dff_B_eRRRpXIp0_2),.clk(gclk));
	jdff dff_B_IVmAjTV78_2(.din(w_dff_B_eRRRpXIp0_2),.dout(w_dff_B_IVmAjTV78_2),.clk(gclk));
	jdff dff_B_gwNpEnUi9_2(.din(w_dff_B_IVmAjTV78_2),.dout(w_dff_B_gwNpEnUi9_2),.clk(gclk));
	jdff dff_B_qQtLCcZW8_2(.din(w_dff_B_gwNpEnUi9_2),.dout(w_dff_B_qQtLCcZW8_2),.clk(gclk));
	jdff dff_B_US5NXbHh4_2(.din(w_dff_B_qQtLCcZW8_2),.dout(w_dff_B_US5NXbHh4_2),.clk(gclk));
	jdff dff_B_stTWBR3N5_2(.din(w_dff_B_US5NXbHh4_2),.dout(w_dff_B_stTWBR3N5_2),.clk(gclk));
	jdff dff_B_G3VAygMi9_2(.din(w_dff_B_stTWBR3N5_2),.dout(w_dff_B_G3VAygMi9_2),.clk(gclk));
	jdff dff_B_iK4WsCJd2_2(.din(w_dff_B_G3VAygMi9_2),.dout(w_dff_B_iK4WsCJd2_2),.clk(gclk));
	jdff dff_B_ROPJrve65_2(.din(w_dff_B_iK4WsCJd2_2),.dout(w_dff_B_ROPJrve65_2),.clk(gclk));
	jdff dff_B_9niJIMgr0_2(.din(w_dff_B_ROPJrve65_2),.dout(w_dff_B_9niJIMgr0_2),.clk(gclk));
	jdff dff_B_EdPmcdeZ2_2(.din(w_dff_B_9niJIMgr0_2),.dout(w_dff_B_EdPmcdeZ2_2),.clk(gclk));
	jdff dff_B_rFZjnwEp4_2(.din(w_dff_B_EdPmcdeZ2_2),.dout(w_dff_B_rFZjnwEp4_2),.clk(gclk));
	jdff dff_B_BIhyteCr6_2(.din(w_dff_B_rFZjnwEp4_2),.dout(w_dff_B_BIhyteCr6_2),.clk(gclk));
	jdff dff_B_WIVEVmRH9_2(.din(w_dff_B_BIhyteCr6_2),.dout(w_dff_B_WIVEVmRH9_2),.clk(gclk));
	jdff dff_B_sM6oXN572_2(.din(w_dff_B_WIVEVmRH9_2),.dout(w_dff_B_sM6oXN572_2),.clk(gclk));
	jdff dff_B_rNzDtf1p1_2(.din(w_dff_B_sM6oXN572_2),.dout(w_dff_B_rNzDtf1p1_2),.clk(gclk));
	jdff dff_B_wYEHWQGJ7_2(.din(w_dff_B_rNzDtf1p1_2),.dout(w_dff_B_wYEHWQGJ7_2),.clk(gclk));
	jdff dff_B_R32K0NNh2_2(.din(w_dff_B_wYEHWQGJ7_2),.dout(w_dff_B_R32K0NNh2_2),.clk(gclk));
	jdff dff_B_aqMaFA1e4_2(.din(w_dff_B_R32K0NNh2_2),.dout(w_dff_B_aqMaFA1e4_2),.clk(gclk));
	jdff dff_B_fwWN6pFr6_2(.din(w_dff_B_aqMaFA1e4_2),.dout(w_dff_B_fwWN6pFr6_2),.clk(gclk));
	jdff dff_B_5LmGhSp79_2(.din(w_dff_B_fwWN6pFr6_2),.dout(w_dff_B_5LmGhSp79_2),.clk(gclk));
	jdff dff_B_8vziuG1U6_2(.din(w_dff_B_5LmGhSp79_2),.dout(w_dff_B_8vziuG1U6_2),.clk(gclk));
	jdff dff_B_lTvL2yLB7_2(.din(w_dff_B_8vziuG1U6_2),.dout(w_dff_B_lTvL2yLB7_2),.clk(gclk));
	jdff dff_B_bLrpStSI8_2(.din(w_dff_B_lTvL2yLB7_2),.dout(w_dff_B_bLrpStSI8_2),.clk(gclk));
	jdff dff_B_e2mE2qLA2_2(.din(w_dff_B_bLrpStSI8_2),.dout(w_dff_B_e2mE2qLA2_2),.clk(gclk));
	jdff dff_B_f3mcrV686_2(.din(w_dff_B_e2mE2qLA2_2),.dout(w_dff_B_f3mcrV686_2),.clk(gclk));
	jdff dff_B_nqXoUMTE8_2(.din(w_dff_B_f3mcrV686_2),.dout(w_dff_B_nqXoUMTE8_2),.clk(gclk));
	jdff dff_B_KjwFphHi1_2(.din(w_dff_B_nqXoUMTE8_2),.dout(w_dff_B_KjwFphHi1_2),.clk(gclk));
	jdff dff_B_wz9CJPBy5_2(.din(w_dff_B_KjwFphHi1_2),.dout(w_dff_B_wz9CJPBy5_2),.clk(gclk));
	jdff dff_B_FidPeKuk3_2(.din(w_dff_B_wz9CJPBy5_2),.dout(w_dff_B_FidPeKuk3_2),.clk(gclk));
	jdff dff_B_dt1fWUPw1_2(.din(w_dff_B_FidPeKuk3_2),.dout(w_dff_B_dt1fWUPw1_2),.clk(gclk));
	jdff dff_B_NIFoP6fq5_2(.din(w_dff_B_dt1fWUPw1_2),.dout(w_dff_B_NIFoP6fq5_2),.clk(gclk));
	jdff dff_B_9Pn1QdBa0_2(.din(w_dff_B_NIFoP6fq5_2),.dout(w_dff_B_9Pn1QdBa0_2),.clk(gclk));
	jdff dff_B_Mwdr0ex54_2(.din(w_dff_B_9Pn1QdBa0_2),.dout(w_dff_B_Mwdr0ex54_2),.clk(gclk));
	jdff dff_B_kehcM6Nf6_2(.din(w_dff_B_Mwdr0ex54_2),.dout(w_dff_B_kehcM6Nf6_2),.clk(gclk));
	jdff dff_B_5VJFioyt2_2(.din(w_dff_B_kehcM6Nf6_2),.dout(w_dff_B_5VJFioyt2_2),.clk(gclk));
	jdff dff_B_nVuxINDG6_2(.din(w_dff_B_5VJFioyt2_2),.dout(w_dff_B_nVuxINDG6_2),.clk(gclk));
	jdff dff_B_0dhcWmTo6_2(.din(w_dff_B_nVuxINDG6_2),.dout(w_dff_B_0dhcWmTo6_2),.clk(gclk));
	jdff dff_B_9KcLHECc0_2(.din(w_dff_B_0dhcWmTo6_2),.dout(w_dff_B_9KcLHECc0_2),.clk(gclk));
	jdff dff_B_USHaZjdi7_2(.din(w_dff_B_9KcLHECc0_2),.dout(w_dff_B_USHaZjdi7_2),.clk(gclk));
	jdff dff_B_G5BEgudb6_2(.din(w_dff_B_USHaZjdi7_2),.dout(w_dff_B_G5BEgudb6_2),.clk(gclk));
	jdff dff_B_KgmKOHcP4_2(.din(w_dff_B_G5BEgudb6_2),.dout(w_dff_B_KgmKOHcP4_2),.clk(gclk));
	jdff dff_B_arB0yoaU3_2(.din(w_dff_B_KgmKOHcP4_2),.dout(w_dff_B_arB0yoaU3_2),.clk(gclk));
	jdff dff_B_60rVC1rb0_2(.din(w_dff_B_arB0yoaU3_2),.dout(w_dff_B_60rVC1rb0_2),.clk(gclk));
	jdff dff_B_pu4gjLdZ1_2(.din(w_dff_B_60rVC1rb0_2),.dout(w_dff_B_pu4gjLdZ1_2),.clk(gclk));
	jdff dff_B_P27OR78m7_2(.din(w_dff_B_pu4gjLdZ1_2),.dout(w_dff_B_P27OR78m7_2),.clk(gclk));
	jdff dff_B_IN61Kn5F7_2(.din(w_dff_B_P27OR78m7_2),.dout(w_dff_B_IN61Kn5F7_2),.clk(gclk));
	jdff dff_B_x2hBgIs82_2(.din(w_dff_B_IN61Kn5F7_2),.dout(w_dff_B_x2hBgIs82_2),.clk(gclk));
	jdff dff_B_5H9dfX1j9_2(.din(w_dff_B_x2hBgIs82_2),.dout(w_dff_B_5H9dfX1j9_2),.clk(gclk));
	jdff dff_B_nnpwLxU44_2(.din(w_dff_B_5H9dfX1j9_2),.dout(w_dff_B_nnpwLxU44_2),.clk(gclk));
	jdff dff_B_sCNFtcAp6_2(.din(w_dff_B_nnpwLxU44_2),.dout(w_dff_B_sCNFtcAp6_2),.clk(gclk));
	jdff dff_B_l6vTRmli8_2(.din(w_dff_B_sCNFtcAp6_2),.dout(w_dff_B_l6vTRmli8_2),.clk(gclk));
	jdff dff_B_eztTHDde1_2(.din(w_dff_B_l6vTRmli8_2),.dout(w_dff_B_eztTHDde1_2),.clk(gclk));
	jdff dff_B_3OrDKUJj0_2(.din(w_dff_B_eztTHDde1_2),.dout(w_dff_B_3OrDKUJj0_2),.clk(gclk));
	jdff dff_B_CsiPZSAa2_2(.din(w_dff_B_3OrDKUJj0_2),.dout(w_dff_B_CsiPZSAa2_2),.clk(gclk));
	jdff dff_B_A3V6HJoQ5_2(.din(w_dff_B_CsiPZSAa2_2),.dout(w_dff_B_A3V6HJoQ5_2),.clk(gclk));
	jdff dff_B_ZfCni8gI2_2(.din(w_dff_B_A3V6HJoQ5_2),.dout(w_dff_B_ZfCni8gI2_2),.clk(gclk));
	jdff dff_B_RXClBM164_2(.din(w_dff_B_ZfCni8gI2_2),.dout(w_dff_B_RXClBM164_2),.clk(gclk));
	jdff dff_B_des7wfFf4_2(.din(w_dff_B_RXClBM164_2),.dout(w_dff_B_des7wfFf4_2),.clk(gclk));
	jdff dff_B_wZOj33dQ6_2(.din(w_dff_B_des7wfFf4_2),.dout(w_dff_B_wZOj33dQ6_2),.clk(gclk));
	jdff dff_B_IZsVzRmh2_2(.din(w_dff_B_wZOj33dQ6_2),.dout(w_dff_B_IZsVzRmh2_2),.clk(gclk));
	jdff dff_B_Q1a9kF4g0_2(.din(w_dff_B_IZsVzRmh2_2),.dout(w_dff_B_Q1a9kF4g0_2),.clk(gclk));
	jdff dff_B_2dB8pYrl2_2(.din(w_dff_B_Q1a9kF4g0_2),.dout(w_dff_B_2dB8pYrl2_2),.clk(gclk));
	jdff dff_B_5VfWGz4r1_2(.din(w_dff_B_2dB8pYrl2_2),.dout(w_dff_B_5VfWGz4r1_2),.clk(gclk));
	jdff dff_B_jekYDuP48_2(.din(w_dff_B_5VfWGz4r1_2),.dout(w_dff_B_jekYDuP48_2),.clk(gclk));
	jdff dff_B_DPSlNoRU3_2(.din(w_dff_B_jekYDuP48_2),.dout(w_dff_B_DPSlNoRU3_2),.clk(gclk));
	jdff dff_B_UaVO9muF5_2(.din(w_dff_B_DPSlNoRU3_2),.dout(w_dff_B_UaVO9muF5_2),.clk(gclk));
	jdff dff_B_XY4keW9r7_2(.din(w_dff_B_UaVO9muF5_2),.dout(w_dff_B_XY4keW9r7_2),.clk(gclk));
	jdff dff_B_PMzv3sup1_2(.din(w_dff_B_XY4keW9r7_2),.dout(w_dff_B_PMzv3sup1_2),.clk(gclk));
	jdff dff_B_MZZPo2KJ3_2(.din(w_dff_B_PMzv3sup1_2),.dout(w_dff_B_MZZPo2KJ3_2),.clk(gclk));
	jdff dff_B_ZcgGVSla1_2(.din(w_dff_B_MZZPo2KJ3_2),.dout(w_dff_B_ZcgGVSla1_2),.clk(gclk));
	jdff dff_B_CSnHakR16_2(.din(w_dff_B_ZcgGVSla1_2),.dout(w_dff_B_CSnHakR16_2),.clk(gclk));
	jdff dff_B_WopNUl880_2(.din(w_dff_B_CSnHakR16_2),.dout(w_dff_B_WopNUl880_2),.clk(gclk));
	jdff dff_B_kpt5IzMd0_2(.din(w_dff_B_WopNUl880_2),.dout(w_dff_B_kpt5IzMd0_2),.clk(gclk));
	jdff dff_B_qTnEM4Pf4_2(.din(w_dff_B_kpt5IzMd0_2),.dout(w_dff_B_qTnEM4Pf4_2),.clk(gclk));
	jdff dff_B_29I4CNV09_2(.din(w_dff_B_qTnEM4Pf4_2),.dout(w_dff_B_29I4CNV09_2),.clk(gclk));
	jdff dff_B_uO0oUmgB6_2(.din(w_dff_B_29I4CNV09_2),.dout(w_dff_B_uO0oUmgB6_2),.clk(gclk));
	jdff dff_B_tDJHiKPo9_2(.din(w_dff_B_uO0oUmgB6_2),.dout(w_dff_B_tDJHiKPo9_2),.clk(gclk));
	jdff dff_B_4qVYnJ1F4_2(.din(w_dff_B_tDJHiKPo9_2),.dout(w_dff_B_4qVYnJ1F4_2),.clk(gclk));
	jdff dff_B_xXAtKyuR3_2(.din(w_dff_B_4qVYnJ1F4_2),.dout(w_dff_B_xXAtKyuR3_2),.clk(gclk));
	jdff dff_B_uISo6LVc5_2(.din(w_dff_B_xXAtKyuR3_2),.dout(w_dff_B_uISo6LVc5_2),.clk(gclk));
	jdff dff_B_IoTRuWhs9_2(.din(w_dff_B_uISo6LVc5_2),.dout(w_dff_B_IoTRuWhs9_2),.clk(gclk));
	jdff dff_B_fouTRMzq4_2(.din(w_dff_B_IoTRuWhs9_2),.dout(w_dff_B_fouTRMzq4_2),.clk(gclk));
	jdff dff_B_upVwaqff9_2(.din(w_dff_B_fouTRMzq4_2),.dout(w_dff_B_upVwaqff9_2),.clk(gclk));
	jdff dff_B_9K6zKB0w6_2(.din(w_dff_B_upVwaqff9_2),.dout(w_dff_B_9K6zKB0w6_2),.clk(gclk));
	jdff dff_B_RdJkpfpH4_2(.din(w_dff_B_9K6zKB0w6_2),.dout(w_dff_B_RdJkpfpH4_2),.clk(gclk));
	jdff dff_B_zUuRNuqY6_2(.din(w_dff_B_RdJkpfpH4_2),.dout(w_dff_B_zUuRNuqY6_2),.clk(gclk));
	jdff dff_B_TemKBV990_2(.din(w_dff_B_zUuRNuqY6_2),.dout(w_dff_B_TemKBV990_2),.clk(gclk));
	jdff dff_B_TeEVRnbd9_2(.din(w_dff_B_TemKBV990_2),.dout(w_dff_B_TeEVRnbd9_2),.clk(gclk));
	jdff dff_B_8hC2alfW9_2(.din(w_dff_B_TeEVRnbd9_2),.dout(w_dff_B_8hC2alfW9_2),.clk(gclk));
	jdff dff_B_G9uczfGb9_2(.din(w_dff_B_8hC2alfW9_2),.dout(w_dff_B_G9uczfGb9_2),.clk(gclk));
	jdff dff_B_IPG6jWwi7_2(.din(w_dff_B_G9uczfGb9_2),.dout(w_dff_B_IPG6jWwi7_2),.clk(gclk));
	jdff dff_B_RTxZitcs4_2(.din(w_dff_B_IPG6jWwi7_2),.dout(w_dff_B_RTxZitcs4_2),.clk(gclk));
	jdff dff_B_7ujJIy5n9_2(.din(w_dff_B_RTxZitcs4_2),.dout(w_dff_B_7ujJIy5n9_2),.clk(gclk));
	jdff dff_B_9RaeZEvG0_2(.din(w_dff_B_7ujJIy5n9_2),.dout(w_dff_B_9RaeZEvG0_2),.clk(gclk));
	jdff dff_B_xRMqeGPe7_2(.din(w_dff_B_9RaeZEvG0_2),.dout(w_dff_B_xRMqeGPe7_2),.clk(gclk));
	jdff dff_B_stWHUBP12_2(.din(w_dff_B_xRMqeGPe7_2),.dout(w_dff_B_stWHUBP12_2),.clk(gclk));
	jdff dff_B_OWlWKqxz0_2(.din(w_dff_B_stWHUBP12_2),.dout(w_dff_B_OWlWKqxz0_2),.clk(gclk));
	jdff dff_B_5SXokDAm3_2(.din(w_dff_B_OWlWKqxz0_2),.dout(w_dff_B_5SXokDAm3_2),.clk(gclk));
	jdff dff_B_9U6RuGSZ9_2(.din(w_dff_B_5SXokDAm3_2),.dout(w_dff_B_9U6RuGSZ9_2),.clk(gclk));
	jdff dff_B_J653GGjn7_2(.din(w_dff_B_9U6RuGSZ9_2),.dout(w_dff_B_J653GGjn7_2),.clk(gclk));
	jdff dff_B_389mS7mG7_2(.din(w_dff_B_J653GGjn7_2),.dout(w_dff_B_389mS7mG7_2),.clk(gclk));
	jdff dff_B_d9hBrptt6_0(.din(n5153),.dout(w_dff_B_d9hBrptt6_0),.clk(gclk));
	jdff dff_A_OaMuw6Hb9_1(.dout(w_n5133_0[1]),.din(w_dff_A_OaMuw6Hb9_1),.clk(gclk));
	jdff dff_B_4LMWvph54_1(.din(n5086),.dout(w_dff_B_4LMWvph54_1),.clk(gclk));
	jdff dff_A_Xhuy3IJF7_0(.dout(w_n5024_0[0]),.din(w_dff_A_Xhuy3IJF7_0),.clk(gclk));
	jdff dff_A_awo5l0ir3_0(.dout(w_n5021_0[0]),.din(w_dff_A_awo5l0ir3_0),.clk(gclk));
	jdff dff_A_HPuTasns0_0(.dout(w_dff_A_awo5l0ir3_0),.din(w_dff_A_HPuTasns0_0),.clk(gclk));
	jdff dff_A_wxzz2WBi3_0(.dout(w_n4986_0[0]),.din(w_dff_A_wxzz2WBi3_0),.clk(gclk));
	jdff dff_A_e94k11f77_0(.dout(w_n4943_0[0]),.din(w_dff_A_e94k11f77_0),.clk(gclk));
	jdff dff_A_yIbGSoVr3_0(.dout(w_n4896_0[0]),.din(w_dff_A_yIbGSoVr3_0),.clk(gclk));
	jdff dff_A_sOErIqr07_0(.dout(w_n4840_0[0]),.din(w_dff_A_sOErIqr07_0),.clk(gclk));
	jdff dff_A_fGY52gbv0_0(.dout(w_n4789_0[0]),.din(w_dff_A_fGY52gbv0_0),.clk(gclk));
	jdff dff_A_72JVXFet2_0(.dout(w_n4732_0[0]),.din(w_dff_A_72JVXFet2_0),.clk(gclk));
	jdff dff_A_J0qwBfzZ9_0(.dout(w_n4667_0[0]),.din(w_dff_A_J0qwBfzZ9_0),.clk(gclk));
	jdff dff_A_h9g6HZkd4_0(.dout(w_n4603_0[0]),.din(w_dff_A_h9g6HZkd4_0),.clk(gclk));
	jdff dff_A_SMxcsPby6_0(.dout(w_n4527_0[0]),.din(w_dff_A_SMxcsPby6_0),.clk(gclk));
	jdff dff_A_gjRzRkwI1_0(.dout(w_n4454_0[0]),.din(w_dff_A_gjRzRkwI1_0),.clk(gclk));
	jdff dff_A_t9pi2k7w5_0(.dout(w_n4372_0[0]),.din(w_dff_A_t9pi2k7w5_0),.clk(gclk));
	jdff dff_A_uVwNu9Rb1_0(.dout(w_n4290_0[0]),.din(w_dff_A_uVwNu9Rb1_0),.clk(gclk));
	jdff dff_A_vDPcnB1Q5_0(.dout(w_n4123_0[0]),.din(w_dff_A_vDPcnB1Q5_0),.clk(gclk));
	jdff dff_A_l5ALSQ9k4_0(.dout(w_n4120_0[0]),.din(w_dff_A_l5ALSQ9k4_0),.clk(gclk));
	jdff dff_A_UK3GPCLL0_0(.dout(w_sin0_0[0]),.din(w_dff_A_UK3GPCLL0_0),.clk(gclk));
	jdff dff_A_Op0hX5fq0_0(.dout(w_dff_A_UK3GPCLL0_0),.din(w_dff_A_Op0hX5fq0_0),.clk(gclk));
	jdff dff_A_W48FiSy24_1(.dout(w_n5085_0[1]),.din(w_dff_A_W48FiSy24_1),.clk(gclk));
	jdff dff_B_elMsNUXc0_2(.din(n5085),.dout(w_dff_B_elMsNUXc0_2),.clk(gclk));
	jdff dff_A_lr3QEvLc2_1(.dout(w_n5120_0[1]),.din(w_dff_A_lr3QEvLc2_1),.clk(gclk));
	jdff dff_B_QvlyzZXy5_2(.din(n5120),.dout(w_dff_B_QvlyzZXy5_2),.clk(gclk));
	jdff dff_A_UKMe566N2_1(.dout(w_n4013_3[1]),.din(w_dff_A_UKMe566N2_1),.clk(gclk));
	jdff dff_A_fx7a37RG8_1(.dout(w_dff_A_UKMe566N2_1),.din(w_dff_A_fx7a37RG8_1),.clk(gclk));
	jdff dff_A_FN0f6bzQ8_1(.dout(w_dff_A_fx7a37RG8_1),.din(w_dff_A_FN0f6bzQ8_1),.clk(gclk));
	jdff dff_A_o1vAK5iq7_1(.dout(w_dff_A_FN0f6bzQ8_1),.din(w_dff_A_o1vAK5iq7_1),.clk(gclk));
	jdff dff_A_nBj4kGVC4_1(.dout(w_dff_A_o1vAK5iq7_1),.din(w_dff_A_nBj4kGVC4_1),.clk(gclk));
	jdff dff_A_jzz1ksPd0_1(.dout(w_dff_A_nBj4kGVC4_1),.din(w_dff_A_jzz1ksPd0_1),.clk(gclk));
	jdff dff_A_2BWMdtY83_1(.dout(w_dff_A_jzz1ksPd0_1),.din(w_dff_A_2BWMdtY83_1),.clk(gclk));
	jdff dff_A_xcEohffX4_1(.dout(w_dff_A_2BWMdtY83_1),.din(w_dff_A_xcEohffX4_1),.clk(gclk));
	jdff dff_A_C2jk7L929_1(.dout(w_dff_A_xcEohffX4_1),.din(w_dff_A_C2jk7L929_1),.clk(gclk));
	jdff dff_A_jFPvwqMJ4_1(.dout(w_dff_A_C2jk7L929_1),.din(w_dff_A_jFPvwqMJ4_1),.clk(gclk));
	jdff dff_A_dWFmD96g4_1(.dout(w_dff_A_jFPvwqMJ4_1),.din(w_dff_A_dWFmD96g4_1),.clk(gclk));
	jdff dff_A_itrUM3iV6_1(.dout(w_dff_A_dWFmD96g4_1),.din(w_dff_A_itrUM3iV6_1),.clk(gclk));
	jdff dff_A_ECp7BdkB5_1(.dout(w_dff_A_itrUM3iV6_1),.din(w_dff_A_ECp7BdkB5_1),.clk(gclk));
	jdff dff_A_YkCbqYno9_1(.dout(w_dff_A_ECp7BdkB5_1),.din(w_dff_A_YkCbqYno9_1),.clk(gclk));
	jdff dff_A_onfvbgBw3_1(.dout(w_dff_A_YkCbqYno9_1),.din(w_dff_A_onfvbgBw3_1),.clk(gclk));
	jdff dff_A_hngeokM71_1(.dout(w_dff_A_onfvbgBw3_1),.din(w_dff_A_hngeokM71_1),.clk(gclk));
	jdff dff_A_s9ntx8NO3_1(.dout(w_dff_A_hngeokM71_1),.din(w_dff_A_s9ntx8NO3_1),.clk(gclk));
	jdff dff_A_qzWxn6461_1(.dout(w_dff_A_s9ntx8NO3_1),.din(w_dff_A_qzWxn6461_1),.clk(gclk));
	jdff dff_A_ut645Deh1_1(.dout(w_dff_A_qzWxn6461_1),.din(w_dff_A_ut645Deh1_1),.clk(gclk));
	jdff dff_A_V7hMOjCO9_1(.dout(w_dff_A_ut645Deh1_1),.din(w_dff_A_V7hMOjCO9_1),.clk(gclk));
	jdff dff_A_YIRDUDk07_1(.dout(w_dff_A_V7hMOjCO9_1),.din(w_dff_A_YIRDUDk07_1),.clk(gclk));
	jdff dff_A_gVYHnMqv1_1(.dout(w_dff_A_YIRDUDk07_1),.din(w_dff_A_gVYHnMqv1_1),.clk(gclk));
	jdff dff_A_fTytwo4O6_1(.dout(w_dff_A_gVYHnMqv1_1),.din(w_dff_A_fTytwo4O6_1),.clk(gclk));
	jdff dff_A_z38fvWZc0_1(.dout(w_dff_A_fTytwo4O6_1),.din(w_dff_A_z38fvWZc0_1),.clk(gclk));
	jdff dff_A_Vzxv9Uwi8_1(.dout(w_dff_A_z38fvWZc0_1),.din(w_dff_A_Vzxv9Uwi8_1),.clk(gclk));
	jdff dff_A_rmUArDBM2_1(.dout(w_dff_A_Vzxv9Uwi8_1),.din(w_dff_A_rmUArDBM2_1),.clk(gclk));
	jdff dff_A_p1UN0wUm4_1(.dout(w_dff_A_rmUArDBM2_1),.din(w_dff_A_p1UN0wUm4_1),.clk(gclk));
	jdff dff_A_RyfUTes05_1(.dout(w_dff_A_p1UN0wUm4_1),.din(w_dff_A_RyfUTes05_1),.clk(gclk));
	jdff dff_A_SZhjyTSy6_1(.dout(w_dff_A_RyfUTes05_1),.din(w_dff_A_SZhjyTSy6_1),.clk(gclk));
	jdff dff_A_aj04g3bj4_1(.dout(w_dff_A_SZhjyTSy6_1),.din(w_dff_A_aj04g3bj4_1),.clk(gclk));
	jdff dff_A_gY7FIhkc5_1(.dout(w_dff_A_aj04g3bj4_1),.din(w_dff_A_gY7FIhkc5_1),.clk(gclk));
	jdff dff_A_wCli2Gti0_1(.dout(w_dff_A_gY7FIhkc5_1),.din(w_dff_A_wCli2Gti0_1),.clk(gclk));
	jdff dff_A_5vjv4XYO9_1(.dout(w_dff_A_wCli2Gti0_1),.din(w_dff_A_5vjv4XYO9_1),.clk(gclk));
	jdff dff_A_b9mZ2KQB0_1(.dout(w_dff_A_5vjv4XYO9_1),.din(w_dff_A_b9mZ2KQB0_1),.clk(gclk));
	jdff dff_A_ivunJrwH4_1(.dout(w_dff_A_b9mZ2KQB0_1),.din(w_dff_A_ivunJrwH4_1),.clk(gclk));
	jdff dff_A_lGfZrXAS9_1(.dout(w_dff_A_ivunJrwH4_1),.din(w_dff_A_lGfZrXAS9_1),.clk(gclk));
	jdff dff_A_7IGeBWFh0_1(.dout(w_dff_A_lGfZrXAS9_1),.din(w_dff_A_7IGeBWFh0_1),.clk(gclk));
	jdff dff_A_1coDZ5kC2_1(.dout(w_dff_A_7IGeBWFh0_1),.din(w_dff_A_1coDZ5kC2_1),.clk(gclk));
	jdff dff_A_sEhaFDJJ0_1(.dout(w_dff_A_1coDZ5kC2_1),.din(w_dff_A_sEhaFDJJ0_1),.clk(gclk));
	jdff dff_A_y5jKn7ty6_1(.dout(w_dff_A_sEhaFDJJ0_1),.din(w_dff_A_y5jKn7ty6_1),.clk(gclk));
	jdff dff_A_TPHP4biu1_1(.dout(w_dff_A_y5jKn7ty6_1),.din(w_dff_A_TPHP4biu1_1),.clk(gclk));
	jdff dff_A_pxaZNlSl4_1(.dout(w_dff_A_TPHP4biu1_1),.din(w_dff_A_pxaZNlSl4_1),.clk(gclk));
	jdff dff_A_RAC8Yl7x7_1(.dout(w_dff_A_pxaZNlSl4_1),.din(w_dff_A_RAC8Yl7x7_1),.clk(gclk));
	jdff dff_A_0eyV9lEz2_1(.dout(w_dff_A_RAC8Yl7x7_1),.din(w_dff_A_0eyV9lEz2_1),.clk(gclk));
	jdff dff_A_mNgCQiig8_2(.dout(w_n4013_3[2]),.din(w_dff_A_mNgCQiig8_2),.clk(gclk));
	jdff dff_A_y1nXRSnK5_2(.dout(w_dff_A_mNgCQiig8_2),.din(w_dff_A_y1nXRSnK5_2),.clk(gclk));
	jdff dff_A_B5Ac0O8K5_2(.dout(w_dff_A_y1nXRSnK5_2),.din(w_dff_A_B5Ac0O8K5_2),.clk(gclk));
	jdff dff_A_swxcqNDD5_2(.dout(w_dff_A_B5Ac0O8K5_2),.din(w_dff_A_swxcqNDD5_2),.clk(gclk));
	jdff dff_A_T8Lxu1iO5_2(.dout(w_dff_A_swxcqNDD5_2),.din(w_dff_A_T8Lxu1iO5_2),.clk(gclk));
	jdff dff_A_73Tdf7ol7_2(.dout(w_dff_A_T8Lxu1iO5_2),.din(w_dff_A_73Tdf7ol7_2),.clk(gclk));
	jdff dff_A_4SoxahjL2_2(.dout(w_dff_A_73Tdf7ol7_2),.din(w_dff_A_4SoxahjL2_2),.clk(gclk));
	jdff dff_A_WFxcwB9S2_2(.dout(w_dff_A_4SoxahjL2_2),.din(w_dff_A_WFxcwB9S2_2),.clk(gclk));
	jdff dff_A_9sVERyzN7_2(.dout(w_dff_A_WFxcwB9S2_2),.din(w_dff_A_9sVERyzN7_2),.clk(gclk));
	jdff dff_A_3CfDnksh3_2(.dout(w_dff_A_9sVERyzN7_2),.din(w_dff_A_3CfDnksh3_2),.clk(gclk));
	jdff dff_A_5pjEuW558_2(.dout(w_dff_A_3CfDnksh3_2),.din(w_dff_A_5pjEuW558_2),.clk(gclk));
	jdff dff_A_f6tYevuC1_2(.dout(w_dff_A_5pjEuW558_2),.din(w_dff_A_f6tYevuC1_2),.clk(gclk));
	jdff dff_A_AhKoH0QZ0_2(.dout(w_dff_A_f6tYevuC1_2),.din(w_dff_A_AhKoH0QZ0_2),.clk(gclk));
	jdff dff_A_HjELsC5A1_2(.dout(w_dff_A_AhKoH0QZ0_2),.din(w_dff_A_HjELsC5A1_2),.clk(gclk));
	jdff dff_A_8q8Q82ie9_2(.dout(w_dff_A_HjELsC5A1_2),.din(w_dff_A_8q8Q82ie9_2),.clk(gclk));
	jdff dff_A_3QogiG4a1_2(.dout(w_dff_A_8q8Q82ie9_2),.din(w_dff_A_3QogiG4a1_2),.clk(gclk));
	jdff dff_A_7fIuVTFi8_2(.dout(w_dff_A_3QogiG4a1_2),.din(w_dff_A_7fIuVTFi8_2),.clk(gclk));
	jdff dff_A_udxvaf216_2(.dout(w_dff_A_7fIuVTFi8_2),.din(w_dff_A_udxvaf216_2),.clk(gclk));
	jdff dff_A_vY1EVIxP6_2(.dout(w_dff_A_udxvaf216_2),.din(w_dff_A_vY1EVIxP6_2),.clk(gclk));
	jdff dff_A_wWyWsqDQ0_2(.dout(w_dff_A_vY1EVIxP6_2),.din(w_dff_A_wWyWsqDQ0_2),.clk(gclk));
	jdff dff_A_RjO5YV3n9_2(.dout(w_dff_A_wWyWsqDQ0_2),.din(w_dff_A_RjO5YV3n9_2),.clk(gclk));
	jdff dff_A_Vdt1oG7S1_2(.dout(w_dff_A_RjO5YV3n9_2),.din(w_dff_A_Vdt1oG7S1_2),.clk(gclk));
	jdff dff_A_8zMVLYsD9_2(.dout(w_dff_A_Vdt1oG7S1_2),.din(w_dff_A_8zMVLYsD9_2),.clk(gclk));
	jdff dff_A_ibcF77I59_2(.dout(w_dff_A_8zMVLYsD9_2),.din(w_dff_A_ibcF77I59_2),.clk(gclk));
	jdff dff_A_7ubQB2Fm9_2(.dout(w_dff_A_ibcF77I59_2),.din(w_dff_A_7ubQB2Fm9_2),.clk(gclk));
	jdff dff_A_AcWnmXhW1_2(.dout(w_dff_A_7ubQB2Fm9_2),.din(w_dff_A_AcWnmXhW1_2),.clk(gclk));
	jdff dff_A_p7j1aMtU4_2(.dout(w_dff_A_AcWnmXhW1_2),.din(w_dff_A_p7j1aMtU4_2),.clk(gclk));
	jdff dff_A_UNRhocXR4_2(.dout(w_dff_A_p7j1aMtU4_2),.din(w_dff_A_UNRhocXR4_2),.clk(gclk));
	jdff dff_A_Gdxe3ZOr8_2(.dout(w_dff_A_UNRhocXR4_2),.din(w_dff_A_Gdxe3ZOr8_2),.clk(gclk));
	jdff dff_A_fzySm9kS8_2(.dout(w_dff_A_Gdxe3ZOr8_2),.din(w_dff_A_fzySm9kS8_2),.clk(gclk));
	jdff dff_A_31Yp8lUP4_2(.dout(w_dff_A_fzySm9kS8_2),.din(w_dff_A_31Yp8lUP4_2),.clk(gclk));
	jdff dff_A_YLtUBQWC8_2(.dout(w_dff_A_31Yp8lUP4_2),.din(w_dff_A_YLtUBQWC8_2),.clk(gclk));
	jdff dff_A_ctpukIw40_2(.dout(w_dff_A_YLtUBQWC8_2),.din(w_dff_A_ctpukIw40_2),.clk(gclk));
	jdff dff_A_MG8GSihc2_2(.dout(w_dff_A_ctpukIw40_2),.din(w_dff_A_MG8GSihc2_2),.clk(gclk));
	jdff dff_A_WvCZHVW40_2(.dout(w_dff_A_MG8GSihc2_2),.din(w_dff_A_WvCZHVW40_2),.clk(gclk));
	jdff dff_A_bg1MJ6p33_2(.dout(w_dff_A_WvCZHVW40_2),.din(w_dff_A_bg1MJ6p33_2),.clk(gclk));
	jdff dff_A_A8d9CICa0_2(.dout(w_dff_A_bg1MJ6p33_2),.din(w_dff_A_A8d9CICa0_2),.clk(gclk));
	jdff dff_A_6lPvK0jv6_2(.dout(w_dff_A_A8d9CICa0_2),.din(w_dff_A_6lPvK0jv6_2),.clk(gclk));
	jdff dff_A_uotJZMkN8_2(.dout(w_dff_A_6lPvK0jv6_2),.din(w_dff_A_uotJZMkN8_2),.clk(gclk));
	jdff dff_A_z8MM6RZQ8_2(.dout(w_dff_A_uotJZMkN8_2),.din(w_dff_A_z8MM6RZQ8_2),.clk(gclk));
	jdff dff_A_aRGfLVlE1_2(.dout(w_dff_A_z8MM6RZQ8_2),.din(w_dff_A_aRGfLVlE1_2),.clk(gclk));
	jdff dff_A_OxUIVHDa5_2(.dout(w_dff_A_aRGfLVlE1_2),.din(w_dff_A_OxUIVHDa5_2),.clk(gclk));
	jdff dff_A_D1xwlsPT1_2(.dout(w_dff_A_YXCB7zUl6_0),.din(w_dff_A_D1xwlsPT1_2),.clk(gclk));
	jdff dff_A_YXCB7zUl6_0(.dout(w_dff_A_70lp1gHR9_0),.din(w_dff_A_YXCB7zUl6_0),.clk(gclk));
	jdff dff_A_70lp1gHR9_0(.dout(w_dff_A_M3Z5D07K8_0),.din(w_dff_A_70lp1gHR9_0),.clk(gclk));
	jdff dff_A_M3Z5D07K8_0(.dout(w_dff_A_tEixc4cS7_0),.din(w_dff_A_M3Z5D07K8_0),.clk(gclk));
	jdff dff_A_tEixc4cS7_0(.dout(w_dff_A_4kdarGqW1_0),.din(w_dff_A_tEixc4cS7_0),.clk(gclk));
	jdff dff_A_4kdarGqW1_0(.dout(w_dff_A_r4dvnVmN5_0),.din(w_dff_A_4kdarGqW1_0),.clk(gclk));
	jdff dff_A_r4dvnVmN5_0(.dout(w_dff_A_iJdPwCoZ2_0),.din(w_dff_A_r4dvnVmN5_0),.clk(gclk));
	jdff dff_A_iJdPwCoZ2_0(.dout(w_dff_A_hWB0jgn51_0),.din(w_dff_A_iJdPwCoZ2_0),.clk(gclk));
	jdff dff_A_hWB0jgn51_0(.dout(w_dff_A_AbMz5S2W1_0),.din(w_dff_A_hWB0jgn51_0),.clk(gclk));
	jdff dff_A_AbMz5S2W1_0(.dout(w_dff_A_pVHLXphT4_0),.din(w_dff_A_AbMz5S2W1_0),.clk(gclk));
	jdff dff_A_pVHLXphT4_0(.dout(w_dff_A_zgCEQf6q4_0),.din(w_dff_A_pVHLXphT4_0),.clk(gclk));
	jdff dff_A_zgCEQf6q4_0(.dout(w_dff_A_xYlQIh4F1_0),.din(w_dff_A_zgCEQf6q4_0),.clk(gclk));
	jdff dff_A_xYlQIh4F1_0(.dout(w_dff_A_jUJfMBc59_0),.din(w_dff_A_xYlQIh4F1_0),.clk(gclk));
	jdff dff_A_jUJfMBc59_0(.dout(w_dff_A_j28GR6Ov8_0),.din(w_dff_A_jUJfMBc59_0),.clk(gclk));
	jdff dff_A_j28GR6Ov8_0(.dout(w_dff_A_61HnOdxT1_0),.din(w_dff_A_j28GR6Ov8_0),.clk(gclk));
	jdff dff_A_61HnOdxT1_0(.dout(w_dff_A_zkxOXXab0_0),.din(w_dff_A_61HnOdxT1_0),.clk(gclk));
	jdff dff_A_zkxOXXab0_0(.dout(w_dff_A_JcGOeZhc4_0),.din(w_dff_A_zkxOXXab0_0),.clk(gclk));
	jdff dff_A_JcGOeZhc4_0(.dout(w_dff_A_wJDD0g888_0),.din(w_dff_A_JcGOeZhc4_0),.clk(gclk));
	jdff dff_A_wJDD0g888_0(.dout(w_dff_A_kpW8vJ3c7_0),.din(w_dff_A_wJDD0g888_0),.clk(gclk));
	jdff dff_A_kpW8vJ3c7_0(.dout(w_dff_A_J0azdLdr1_0),.din(w_dff_A_kpW8vJ3c7_0),.clk(gclk));
	jdff dff_A_J0azdLdr1_0(.dout(w_dff_A_bXsos5Wl2_0),.din(w_dff_A_J0azdLdr1_0),.clk(gclk));
	jdff dff_A_bXsos5Wl2_0(.dout(w_dff_A_enFVIsB98_0),.din(w_dff_A_bXsos5Wl2_0),.clk(gclk));
	jdff dff_A_enFVIsB98_0(.dout(w_dff_A_OWD1bF6y3_0),.din(w_dff_A_enFVIsB98_0),.clk(gclk));
	jdff dff_A_OWD1bF6y3_0(.dout(w_dff_A_m8hIAkfz1_0),.din(w_dff_A_OWD1bF6y3_0),.clk(gclk));
	jdff dff_A_m8hIAkfz1_0(.dout(w_dff_A_uCWGAXRX0_0),.din(w_dff_A_m8hIAkfz1_0),.clk(gclk));
	jdff dff_A_uCWGAXRX0_0(.dout(w_dff_A_iBSl5plc3_0),.din(w_dff_A_uCWGAXRX0_0),.clk(gclk));
	jdff dff_A_iBSl5plc3_0(.dout(w_dff_A_zuskG7SG9_0),.din(w_dff_A_iBSl5plc3_0),.clk(gclk));
	jdff dff_A_zuskG7SG9_0(.dout(w_dff_A_HhPqdd4l1_0),.din(w_dff_A_zuskG7SG9_0),.clk(gclk));
	jdff dff_A_HhPqdd4l1_0(.dout(w_dff_A_jIrz6R3B2_0),.din(w_dff_A_HhPqdd4l1_0),.clk(gclk));
	jdff dff_A_jIrz6R3B2_0(.dout(w_dff_A_q483wXra7_0),.din(w_dff_A_jIrz6R3B2_0),.clk(gclk));
	jdff dff_A_q483wXra7_0(.dout(w_dff_A_6nVV6T3c0_0),.din(w_dff_A_q483wXra7_0),.clk(gclk));
	jdff dff_A_6nVV6T3c0_0(.dout(w_dff_A_Sd21q1ia2_0),.din(w_dff_A_6nVV6T3c0_0),.clk(gclk));
	jdff dff_A_Sd21q1ia2_0(.dout(w_dff_A_NBkdc1KW1_0),.din(w_dff_A_Sd21q1ia2_0),.clk(gclk));
	jdff dff_A_NBkdc1KW1_0(.dout(w_dff_A_YBOdL1Ul3_0),.din(w_dff_A_NBkdc1KW1_0),.clk(gclk));
	jdff dff_A_YBOdL1Ul3_0(.dout(w_dff_A_JKNGIHdO0_0),.din(w_dff_A_YBOdL1Ul3_0),.clk(gclk));
	jdff dff_A_JKNGIHdO0_0(.dout(w_dff_A_D7N8Y8dP1_0),.din(w_dff_A_JKNGIHdO0_0),.clk(gclk));
	jdff dff_A_D7N8Y8dP1_0(.dout(w_dff_A_9WzGAwzG9_0),.din(w_dff_A_D7N8Y8dP1_0),.clk(gclk));
	jdff dff_A_9WzGAwzG9_0(.dout(w_dff_A_NeaAda4q1_0),.din(w_dff_A_9WzGAwzG9_0),.clk(gclk));
	jdff dff_A_NeaAda4q1_0(.dout(w_dff_A_OPaaCXiF3_0),.din(w_dff_A_NeaAda4q1_0),.clk(gclk));
	jdff dff_A_OPaaCXiF3_0(.dout(w_dff_A_Jdw2fPxG9_0),.din(w_dff_A_OPaaCXiF3_0),.clk(gclk));
	jdff dff_A_Jdw2fPxG9_0(.dout(w_dff_A_MNJYD7c20_0),.din(w_dff_A_Jdw2fPxG9_0),.clk(gclk));
	jdff dff_A_MNJYD7c20_0(.dout(w_dff_A_Qwv3AjZl5_0),.din(w_dff_A_MNJYD7c20_0),.clk(gclk));
	jdff dff_A_Qwv3AjZl5_0(.dout(w_dff_A_X6vwduPr4_0),.din(w_dff_A_Qwv3AjZl5_0),.clk(gclk));
	jdff dff_A_X6vwduPr4_0(.dout(w_dff_A_cV0ii5IC2_0),.din(w_dff_A_X6vwduPr4_0),.clk(gclk));
	jdff dff_A_cV0ii5IC2_0(.dout(sin0),.din(w_dff_A_cV0ii5IC2_0),.clk(gclk));
	jdff dff_A_lIGy9qnK1_2(.dout(w_dff_A_Yms946IM2_0),.din(w_dff_A_lIGy9qnK1_2),.clk(gclk));
	jdff dff_A_Yms946IM2_0(.dout(w_dff_A_3O9aB6np8_0),.din(w_dff_A_Yms946IM2_0),.clk(gclk));
	jdff dff_A_3O9aB6np8_0(.dout(w_dff_A_PAMpttRC2_0),.din(w_dff_A_3O9aB6np8_0),.clk(gclk));
	jdff dff_A_PAMpttRC2_0(.dout(w_dff_A_zrqntBIf8_0),.din(w_dff_A_PAMpttRC2_0),.clk(gclk));
	jdff dff_A_zrqntBIf8_0(.dout(w_dff_A_145wPxLy7_0),.din(w_dff_A_zrqntBIf8_0),.clk(gclk));
	jdff dff_A_145wPxLy7_0(.dout(w_dff_A_9KthTZRE2_0),.din(w_dff_A_145wPxLy7_0),.clk(gclk));
	jdff dff_A_9KthTZRE2_0(.dout(w_dff_A_Hs8fM28S0_0),.din(w_dff_A_9KthTZRE2_0),.clk(gclk));
	jdff dff_A_Hs8fM28S0_0(.dout(w_dff_A_19YwcVEl1_0),.din(w_dff_A_Hs8fM28S0_0),.clk(gclk));
	jdff dff_A_19YwcVEl1_0(.dout(w_dff_A_kJTNWExQ8_0),.din(w_dff_A_19YwcVEl1_0),.clk(gclk));
	jdff dff_A_kJTNWExQ8_0(.dout(w_dff_A_lsY5VVDK4_0),.din(w_dff_A_kJTNWExQ8_0),.clk(gclk));
	jdff dff_A_lsY5VVDK4_0(.dout(w_dff_A_VFXng7rv1_0),.din(w_dff_A_lsY5VVDK4_0),.clk(gclk));
	jdff dff_A_VFXng7rv1_0(.dout(w_dff_A_QKhzTLtn4_0),.din(w_dff_A_VFXng7rv1_0),.clk(gclk));
	jdff dff_A_QKhzTLtn4_0(.dout(w_dff_A_6yBjoo4p9_0),.din(w_dff_A_QKhzTLtn4_0),.clk(gclk));
	jdff dff_A_6yBjoo4p9_0(.dout(w_dff_A_Naqlk2Mc8_0),.din(w_dff_A_6yBjoo4p9_0),.clk(gclk));
	jdff dff_A_Naqlk2Mc8_0(.dout(w_dff_A_qk9xSDyE9_0),.din(w_dff_A_Naqlk2Mc8_0),.clk(gclk));
	jdff dff_A_qk9xSDyE9_0(.dout(w_dff_A_IbWlIuzf6_0),.din(w_dff_A_qk9xSDyE9_0),.clk(gclk));
	jdff dff_A_IbWlIuzf6_0(.dout(w_dff_A_IUL2BnbZ9_0),.din(w_dff_A_IbWlIuzf6_0),.clk(gclk));
	jdff dff_A_IUL2BnbZ9_0(.dout(w_dff_A_CwQY95RY8_0),.din(w_dff_A_IUL2BnbZ9_0),.clk(gclk));
	jdff dff_A_CwQY95RY8_0(.dout(w_dff_A_jmmDeEed0_0),.din(w_dff_A_CwQY95RY8_0),.clk(gclk));
	jdff dff_A_jmmDeEed0_0(.dout(w_dff_A_8TPblaNh9_0),.din(w_dff_A_jmmDeEed0_0),.clk(gclk));
	jdff dff_A_8TPblaNh9_0(.dout(w_dff_A_f7gjjkT66_0),.din(w_dff_A_8TPblaNh9_0),.clk(gclk));
	jdff dff_A_f7gjjkT66_0(.dout(w_dff_A_fokDOBqX0_0),.din(w_dff_A_f7gjjkT66_0),.clk(gclk));
	jdff dff_A_fokDOBqX0_0(.dout(w_dff_A_EOkUnT3Y9_0),.din(w_dff_A_fokDOBqX0_0),.clk(gclk));
	jdff dff_A_EOkUnT3Y9_0(.dout(w_dff_A_TU7oweEo5_0),.din(w_dff_A_EOkUnT3Y9_0),.clk(gclk));
	jdff dff_A_TU7oweEo5_0(.dout(w_dff_A_aEPT9noN2_0),.din(w_dff_A_TU7oweEo5_0),.clk(gclk));
	jdff dff_A_aEPT9noN2_0(.dout(w_dff_A_aXfgFULw2_0),.din(w_dff_A_aEPT9noN2_0),.clk(gclk));
	jdff dff_A_aXfgFULw2_0(.dout(w_dff_A_hgtTWBIc1_0),.din(w_dff_A_aXfgFULw2_0),.clk(gclk));
	jdff dff_A_hgtTWBIc1_0(.dout(w_dff_A_YNVxmON74_0),.din(w_dff_A_hgtTWBIc1_0),.clk(gclk));
	jdff dff_A_YNVxmON74_0(.dout(w_dff_A_YGRqTFNp7_0),.din(w_dff_A_YNVxmON74_0),.clk(gclk));
	jdff dff_A_YGRqTFNp7_0(.dout(w_dff_A_QprqWveD2_0),.din(w_dff_A_YGRqTFNp7_0),.clk(gclk));
	jdff dff_A_QprqWveD2_0(.dout(w_dff_A_v4vjErgD4_0),.din(w_dff_A_QprqWveD2_0),.clk(gclk));
	jdff dff_A_v4vjErgD4_0(.dout(w_dff_A_tOf1XTz83_0),.din(w_dff_A_v4vjErgD4_0),.clk(gclk));
	jdff dff_A_tOf1XTz83_0(.dout(w_dff_A_Juh47g114_0),.din(w_dff_A_tOf1XTz83_0),.clk(gclk));
	jdff dff_A_Juh47g114_0(.dout(w_dff_A_0VznXvK52_0),.din(w_dff_A_Juh47g114_0),.clk(gclk));
	jdff dff_A_0VznXvK52_0(.dout(w_dff_A_sVyrxLrU4_0),.din(w_dff_A_0VznXvK52_0),.clk(gclk));
	jdff dff_A_sVyrxLrU4_0(.dout(w_dff_A_BJ9tlNVC8_0),.din(w_dff_A_sVyrxLrU4_0),.clk(gclk));
	jdff dff_A_BJ9tlNVC8_0(.dout(w_dff_A_bY5QyAMS3_0),.din(w_dff_A_BJ9tlNVC8_0),.clk(gclk));
	jdff dff_A_bY5QyAMS3_0(.dout(w_dff_A_2EigPglX2_0),.din(w_dff_A_bY5QyAMS3_0),.clk(gclk));
	jdff dff_A_2EigPglX2_0(.dout(w_dff_A_oo1LMv3F4_0),.din(w_dff_A_2EigPglX2_0),.clk(gclk));
	jdff dff_A_oo1LMv3F4_0(.dout(w_dff_A_baA821cv6_0),.din(w_dff_A_oo1LMv3F4_0),.clk(gclk));
	jdff dff_A_baA821cv6_0(.dout(sin1),.din(w_dff_A_baA821cv6_0),.clk(gclk));
	jdff dff_A_QWIijunn1_2(.dout(w_dff_A_qNegFRs30_0),.din(w_dff_A_QWIijunn1_2),.clk(gclk));
	jdff dff_A_qNegFRs30_0(.dout(w_dff_A_avbzxA8K5_0),.din(w_dff_A_qNegFRs30_0),.clk(gclk));
	jdff dff_A_avbzxA8K5_0(.dout(w_dff_A_XFhLLati8_0),.din(w_dff_A_avbzxA8K5_0),.clk(gclk));
	jdff dff_A_XFhLLati8_0(.dout(w_dff_A_2M6rdHWa8_0),.din(w_dff_A_XFhLLati8_0),.clk(gclk));
	jdff dff_A_2M6rdHWa8_0(.dout(w_dff_A_gaQyrKER4_0),.din(w_dff_A_2M6rdHWa8_0),.clk(gclk));
	jdff dff_A_gaQyrKER4_0(.dout(w_dff_A_evMP8BRa7_0),.din(w_dff_A_gaQyrKER4_0),.clk(gclk));
	jdff dff_A_evMP8BRa7_0(.dout(w_dff_A_Odanodd16_0),.din(w_dff_A_evMP8BRa7_0),.clk(gclk));
	jdff dff_A_Odanodd16_0(.dout(w_dff_A_FHhu5GBy0_0),.din(w_dff_A_Odanodd16_0),.clk(gclk));
	jdff dff_A_FHhu5GBy0_0(.dout(w_dff_A_knwUz8vb8_0),.din(w_dff_A_FHhu5GBy0_0),.clk(gclk));
	jdff dff_A_knwUz8vb8_0(.dout(w_dff_A_PPjjr6Ek2_0),.din(w_dff_A_knwUz8vb8_0),.clk(gclk));
	jdff dff_A_PPjjr6Ek2_0(.dout(w_dff_A_9yiZoM3N6_0),.din(w_dff_A_PPjjr6Ek2_0),.clk(gclk));
	jdff dff_A_9yiZoM3N6_0(.dout(w_dff_A_cLiY4Yhy8_0),.din(w_dff_A_9yiZoM3N6_0),.clk(gclk));
	jdff dff_A_cLiY4Yhy8_0(.dout(w_dff_A_aMxejYF88_0),.din(w_dff_A_cLiY4Yhy8_0),.clk(gclk));
	jdff dff_A_aMxejYF88_0(.dout(w_dff_A_Co6zi4pN5_0),.din(w_dff_A_aMxejYF88_0),.clk(gclk));
	jdff dff_A_Co6zi4pN5_0(.dout(w_dff_A_JQmPX4R77_0),.din(w_dff_A_Co6zi4pN5_0),.clk(gclk));
	jdff dff_A_JQmPX4R77_0(.dout(w_dff_A_dzK2YkCF7_0),.din(w_dff_A_JQmPX4R77_0),.clk(gclk));
	jdff dff_A_dzK2YkCF7_0(.dout(w_dff_A_GyJafjJW1_0),.din(w_dff_A_dzK2YkCF7_0),.clk(gclk));
	jdff dff_A_GyJafjJW1_0(.dout(w_dff_A_yr4ym27S8_0),.din(w_dff_A_GyJafjJW1_0),.clk(gclk));
	jdff dff_A_yr4ym27S8_0(.dout(w_dff_A_baeF2ZlL2_0),.din(w_dff_A_yr4ym27S8_0),.clk(gclk));
	jdff dff_A_baeF2ZlL2_0(.dout(w_dff_A_kDNFZZ2I5_0),.din(w_dff_A_baeF2ZlL2_0),.clk(gclk));
	jdff dff_A_kDNFZZ2I5_0(.dout(w_dff_A_Ld6cAEeq4_0),.din(w_dff_A_kDNFZZ2I5_0),.clk(gclk));
	jdff dff_A_Ld6cAEeq4_0(.dout(w_dff_A_tMFe6DGo4_0),.din(w_dff_A_Ld6cAEeq4_0),.clk(gclk));
	jdff dff_A_tMFe6DGo4_0(.dout(w_dff_A_Jp9QMmEh5_0),.din(w_dff_A_tMFe6DGo4_0),.clk(gclk));
	jdff dff_A_Jp9QMmEh5_0(.dout(w_dff_A_ummB57JS2_0),.din(w_dff_A_Jp9QMmEh5_0),.clk(gclk));
	jdff dff_A_ummB57JS2_0(.dout(w_dff_A_kwixWjqq2_0),.din(w_dff_A_ummB57JS2_0),.clk(gclk));
	jdff dff_A_kwixWjqq2_0(.dout(w_dff_A_Lga8gxrU1_0),.din(w_dff_A_kwixWjqq2_0),.clk(gclk));
	jdff dff_A_Lga8gxrU1_0(.dout(w_dff_A_HmNCNAau6_0),.din(w_dff_A_Lga8gxrU1_0),.clk(gclk));
	jdff dff_A_HmNCNAau6_0(.dout(w_dff_A_DoGQ16Dh2_0),.din(w_dff_A_HmNCNAau6_0),.clk(gclk));
	jdff dff_A_DoGQ16Dh2_0(.dout(w_dff_A_I7ubIESY7_0),.din(w_dff_A_DoGQ16Dh2_0),.clk(gclk));
	jdff dff_A_I7ubIESY7_0(.dout(w_dff_A_NQW85L9I3_0),.din(w_dff_A_I7ubIESY7_0),.clk(gclk));
	jdff dff_A_NQW85L9I3_0(.dout(w_dff_A_V0xTlsNd1_0),.din(w_dff_A_NQW85L9I3_0),.clk(gclk));
	jdff dff_A_V0xTlsNd1_0(.dout(w_dff_A_Z1bnETvS7_0),.din(w_dff_A_V0xTlsNd1_0),.clk(gclk));
	jdff dff_A_Z1bnETvS7_0(.dout(w_dff_A_7ZGjbFEt9_0),.din(w_dff_A_Z1bnETvS7_0),.clk(gclk));
	jdff dff_A_7ZGjbFEt9_0(.dout(w_dff_A_TK6DAxyF5_0),.din(w_dff_A_7ZGjbFEt9_0),.clk(gclk));
	jdff dff_A_TK6DAxyF5_0(.dout(w_dff_A_b7vkck2R3_0),.din(w_dff_A_TK6DAxyF5_0),.clk(gclk));
	jdff dff_A_b7vkck2R3_0(.dout(w_dff_A_QfGEX16i3_0),.din(w_dff_A_b7vkck2R3_0),.clk(gclk));
	jdff dff_A_QfGEX16i3_0(.dout(w_dff_A_RLCHDuhN6_0),.din(w_dff_A_QfGEX16i3_0),.clk(gclk));
	jdff dff_A_RLCHDuhN6_0(.dout(w_dff_A_5YaOfvIe5_0),.din(w_dff_A_RLCHDuhN6_0),.clk(gclk));
	jdff dff_A_5YaOfvIe5_0(.dout(w_dff_A_WcfqmgfR5_0),.din(w_dff_A_5YaOfvIe5_0),.clk(gclk));
	jdff dff_A_WcfqmgfR5_0(.dout(sin2),.din(w_dff_A_WcfqmgfR5_0),.clk(gclk));
	jdff dff_A_oRAz1Nyn2_2(.dout(w_dff_A_ZIdj2CVd0_0),.din(w_dff_A_oRAz1Nyn2_2),.clk(gclk));
	jdff dff_A_ZIdj2CVd0_0(.dout(w_dff_A_YrCGUe8g1_0),.din(w_dff_A_ZIdj2CVd0_0),.clk(gclk));
	jdff dff_A_YrCGUe8g1_0(.dout(w_dff_A_qezTTKHw5_0),.din(w_dff_A_YrCGUe8g1_0),.clk(gclk));
	jdff dff_A_qezTTKHw5_0(.dout(w_dff_A_HMjCTgyV9_0),.din(w_dff_A_qezTTKHw5_0),.clk(gclk));
	jdff dff_A_HMjCTgyV9_0(.dout(w_dff_A_9LHthM2C0_0),.din(w_dff_A_HMjCTgyV9_0),.clk(gclk));
	jdff dff_A_9LHthM2C0_0(.dout(w_dff_A_pyry5Pkw5_0),.din(w_dff_A_9LHthM2C0_0),.clk(gclk));
	jdff dff_A_pyry5Pkw5_0(.dout(w_dff_A_yDgyKOuz4_0),.din(w_dff_A_pyry5Pkw5_0),.clk(gclk));
	jdff dff_A_yDgyKOuz4_0(.dout(w_dff_A_eXPvLlUl4_0),.din(w_dff_A_yDgyKOuz4_0),.clk(gclk));
	jdff dff_A_eXPvLlUl4_0(.dout(w_dff_A_KvjIEHiq3_0),.din(w_dff_A_eXPvLlUl4_0),.clk(gclk));
	jdff dff_A_KvjIEHiq3_0(.dout(w_dff_A_BPaUnHmN9_0),.din(w_dff_A_KvjIEHiq3_0),.clk(gclk));
	jdff dff_A_BPaUnHmN9_0(.dout(w_dff_A_Cw7Z87zf2_0),.din(w_dff_A_BPaUnHmN9_0),.clk(gclk));
	jdff dff_A_Cw7Z87zf2_0(.dout(w_dff_A_O8sqpJQt9_0),.din(w_dff_A_Cw7Z87zf2_0),.clk(gclk));
	jdff dff_A_O8sqpJQt9_0(.dout(w_dff_A_uyKQpU0Y5_0),.din(w_dff_A_O8sqpJQt9_0),.clk(gclk));
	jdff dff_A_uyKQpU0Y5_0(.dout(w_dff_A_phWk8JiG6_0),.din(w_dff_A_uyKQpU0Y5_0),.clk(gclk));
	jdff dff_A_phWk8JiG6_0(.dout(w_dff_A_rqHnH6dV9_0),.din(w_dff_A_phWk8JiG6_0),.clk(gclk));
	jdff dff_A_rqHnH6dV9_0(.dout(w_dff_A_45NN33Gw6_0),.din(w_dff_A_rqHnH6dV9_0),.clk(gclk));
	jdff dff_A_45NN33Gw6_0(.dout(w_dff_A_HfbiPsJi3_0),.din(w_dff_A_45NN33Gw6_0),.clk(gclk));
	jdff dff_A_HfbiPsJi3_0(.dout(w_dff_A_UOM9hux63_0),.din(w_dff_A_HfbiPsJi3_0),.clk(gclk));
	jdff dff_A_UOM9hux63_0(.dout(w_dff_A_cmqib9Zr2_0),.din(w_dff_A_UOM9hux63_0),.clk(gclk));
	jdff dff_A_cmqib9Zr2_0(.dout(w_dff_A_xWbaMkqZ0_0),.din(w_dff_A_cmqib9Zr2_0),.clk(gclk));
	jdff dff_A_xWbaMkqZ0_0(.dout(w_dff_A_a4sGhVbG8_0),.din(w_dff_A_xWbaMkqZ0_0),.clk(gclk));
	jdff dff_A_a4sGhVbG8_0(.dout(w_dff_A_w9uwQoXl7_0),.din(w_dff_A_a4sGhVbG8_0),.clk(gclk));
	jdff dff_A_w9uwQoXl7_0(.dout(w_dff_A_D9xK50206_0),.din(w_dff_A_w9uwQoXl7_0),.clk(gclk));
	jdff dff_A_D9xK50206_0(.dout(w_dff_A_507e3veY6_0),.din(w_dff_A_D9xK50206_0),.clk(gclk));
	jdff dff_A_507e3veY6_0(.dout(w_dff_A_sU5wOAP63_0),.din(w_dff_A_507e3veY6_0),.clk(gclk));
	jdff dff_A_sU5wOAP63_0(.dout(w_dff_A_M7uRXGEH2_0),.din(w_dff_A_sU5wOAP63_0),.clk(gclk));
	jdff dff_A_M7uRXGEH2_0(.dout(w_dff_A_7JZim46d9_0),.din(w_dff_A_M7uRXGEH2_0),.clk(gclk));
	jdff dff_A_7JZim46d9_0(.dout(w_dff_A_YeLKkgj59_0),.din(w_dff_A_7JZim46d9_0),.clk(gclk));
	jdff dff_A_YeLKkgj59_0(.dout(w_dff_A_czoAlkgL1_0),.din(w_dff_A_YeLKkgj59_0),.clk(gclk));
	jdff dff_A_czoAlkgL1_0(.dout(w_dff_A_SvsvTzZc5_0),.din(w_dff_A_czoAlkgL1_0),.clk(gclk));
	jdff dff_A_SvsvTzZc5_0(.dout(w_dff_A_nQWmn73N5_0),.din(w_dff_A_SvsvTzZc5_0),.clk(gclk));
	jdff dff_A_nQWmn73N5_0(.dout(w_dff_A_gtEukHTK3_0),.din(w_dff_A_nQWmn73N5_0),.clk(gclk));
	jdff dff_A_gtEukHTK3_0(.dout(w_dff_A_774uUGHS4_0),.din(w_dff_A_gtEukHTK3_0),.clk(gclk));
	jdff dff_A_774uUGHS4_0(.dout(w_dff_A_rk9oiF4S5_0),.din(w_dff_A_774uUGHS4_0),.clk(gclk));
	jdff dff_A_rk9oiF4S5_0(.dout(w_dff_A_Wc8Xy8Bm5_0),.din(w_dff_A_rk9oiF4S5_0),.clk(gclk));
	jdff dff_A_Wc8Xy8Bm5_0(.dout(w_dff_A_ljXuj8UG9_0),.din(w_dff_A_Wc8Xy8Bm5_0),.clk(gclk));
	jdff dff_A_ljXuj8UG9_0(.dout(w_dff_A_th4yLU1a9_0),.din(w_dff_A_ljXuj8UG9_0),.clk(gclk));
	jdff dff_A_th4yLU1a9_0(.dout(sin3),.din(w_dff_A_th4yLU1a9_0),.clk(gclk));
	jdff dff_A_fQgYMzmB5_2(.dout(w_dff_A_Vm4r6kSA9_0),.din(w_dff_A_fQgYMzmB5_2),.clk(gclk));
	jdff dff_A_Vm4r6kSA9_0(.dout(w_dff_A_cKM4hrn19_0),.din(w_dff_A_Vm4r6kSA9_0),.clk(gclk));
	jdff dff_A_cKM4hrn19_0(.dout(w_dff_A_VQLF6I0m4_0),.din(w_dff_A_cKM4hrn19_0),.clk(gclk));
	jdff dff_A_VQLF6I0m4_0(.dout(w_dff_A_lzWt3GkF0_0),.din(w_dff_A_VQLF6I0m4_0),.clk(gclk));
	jdff dff_A_lzWt3GkF0_0(.dout(w_dff_A_JB4e1KLY0_0),.din(w_dff_A_lzWt3GkF0_0),.clk(gclk));
	jdff dff_A_JB4e1KLY0_0(.dout(w_dff_A_38sI1FJt2_0),.din(w_dff_A_JB4e1KLY0_0),.clk(gclk));
	jdff dff_A_38sI1FJt2_0(.dout(w_dff_A_MSoVkhbI7_0),.din(w_dff_A_38sI1FJt2_0),.clk(gclk));
	jdff dff_A_MSoVkhbI7_0(.dout(w_dff_A_61DNhxX66_0),.din(w_dff_A_MSoVkhbI7_0),.clk(gclk));
	jdff dff_A_61DNhxX66_0(.dout(w_dff_A_Ww5t9rKI9_0),.din(w_dff_A_61DNhxX66_0),.clk(gclk));
	jdff dff_A_Ww5t9rKI9_0(.dout(w_dff_A_iiJwCTWB2_0),.din(w_dff_A_Ww5t9rKI9_0),.clk(gclk));
	jdff dff_A_iiJwCTWB2_0(.dout(w_dff_A_hhVg1E5R5_0),.din(w_dff_A_iiJwCTWB2_0),.clk(gclk));
	jdff dff_A_hhVg1E5R5_0(.dout(w_dff_A_I46BmDXm9_0),.din(w_dff_A_hhVg1E5R5_0),.clk(gclk));
	jdff dff_A_I46BmDXm9_0(.dout(w_dff_A_UIdOnfCi7_0),.din(w_dff_A_I46BmDXm9_0),.clk(gclk));
	jdff dff_A_UIdOnfCi7_0(.dout(w_dff_A_ZnWYDBmG7_0),.din(w_dff_A_UIdOnfCi7_0),.clk(gclk));
	jdff dff_A_ZnWYDBmG7_0(.dout(w_dff_A_5QpdIZtF9_0),.din(w_dff_A_ZnWYDBmG7_0),.clk(gclk));
	jdff dff_A_5QpdIZtF9_0(.dout(w_dff_A_gLvrGR2Y3_0),.din(w_dff_A_5QpdIZtF9_0),.clk(gclk));
	jdff dff_A_gLvrGR2Y3_0(.dout(w_dff_A_2j5wV0QH8_0),.din(w_dff_A_gLvrGR2Y3_0),.clk(gclk));
	jdff dff_A_2j5wV0QH8_0(.dout(w_dff_A_hoEDNDer6_0),.din(w_dff_A_2j5wV0QH8_0),.clk(gclk));
	jdff dff_A_hoEDNDer6_0(.dout(w_dff_A_cPOyXQ3M7_0),.din(w_dff_A_hoEDNDer6_0),.clk(gclk));
	jdff dff_A_cPOyXQ3M7_0(.dout(w_dff_A_rjbXorsZ3_0),.din(w_dff_A_cPOyXQ3M7_0),.clk(gclk));
	jdff dff_A_rjbXorsZ3_0(.dout(w_dff_A_igl3qT3p1_0),.din(w_dff_A_rjbXorsZ3_0),.clk(gclk));
	jdff dff_A_igl3qT3p1_0(.dout(w_dff_A_be6Owouh8_0),.din(w_dff_A_igl3qT3p1_0),.clk(gclk));
	jdff dff_A_be6Owouh8_0(.dout(w_dff_A_X4ZsCPTt0_0),.din(w_dff_A_be6Owouh8_0),.clk(gclk));
	jdff dff_A_X4ZsCPTt0_0(.dout(w_dff_A_dcgbj7sH3_0),.din(w_dff_A_X4ZsCPTt0_0),.clk(gclk));
	jdff dff_A_dcgbj7sH3_0(.dout(w_dff_A_znBA6ZiU0_0),.din(w_dff_A_dcgbj7sH3_0),.clk(gclk));
	jdff dff_A_znBA6ZiU0_0(.dout(w_dff_A_WvlBKI9K8_0),.din(w_dff_A_znBA6ZiU0_0),.clk(gclk));
	jdff dff_A_WvlBKI9K8_0(.dout(w_dff_A_lSRhZmJy2_0),.din(w_dff_A_WvlBKI9K8_0),.clk(gclk));
	jdff dff_A_lSRhZmJy2_0(.dout(w_dff_A_6Mim457e3_0),.din(w_dff_A_lSRhZmJy2_0),.clk(gclk));
	jdff dff_A_6Mim457e3_0(.dout(w_dff_A_SElGqOG34_0),.din(w_dff_A_6Mim457e3_0),.clk(gclk));
	jdff dff_A_SElGqOG34_0(.dout(w_dff_A_ARUYfesm0_0),.din(w_dff_A_SElGqOG34_0),.clk(gclk));
	jdff dff_A_ARUYfesm0_0(.dout(w_dff_A_EODH7g842_0),.din(w_dff_A_ARUYfesm0_0),.clk(gclk));
	jdff dff_A_EODH7g842_0(.dout(w_dff_A_296RwDxi7_0),.din(w_dff_A_EODH7g842_0),.clk(gclk));
	jdff dff_A_296RwDxi7_0(.dout(w_dff_A_eCqOjRHE4_0),.din(w_dff_A_296RwDxi7_0),.clk(gclk));
	jdff dff_A_eCqOjRHE4_0(.dout(w_dff_A_fUDJXR8i0_0),.din(w_dff_A_eCqOjRHE4_0),.clk(gclk));
	jdff dff_A_fUDJXR8i0_0(.dout(w_dff_A_4U5OUJGW4_0),.din(w_dff_A_fUDJXR8i0_0),.clk(gclk));
	jdff dff_A_4U5OUJGW4_0(.dout(sin4),.din(w_dff_A_4U5OUJGW4_0),.clk(gclk));
	jdff dff_A_Zdk0dlCk2_2(.dout(w_dff_A_9yFvthSH3_0),.din(w_dff_A_Zdk0dlCk2_2),.clk(gclk));
	jdff dff_A_9yFvthSH3_0(.dout(w_dff_A_6JejdKBu5_0),.din(w_dff_A_9yFvthSH3_0),.clk(gclk));
	jdff dff_A_6JejdKBu5_0(.dout(w_dff_A_SszONaO97_0),.din(w_dff_A_6JejdKBu5_0),.clk(gclk));
	jdff dff_A_SszONaO97_0(.dout(w_dff_A_DC1s2nnq2_0),.din(w_dff_A_SszONaO97_0),.clk(gclk));
	jdff dff_A_DC1s2nnq2_0(.dout(w_dff_A_CJmFnuZt5_0),.din(w_dff_A_DC1s2nnq2_0),.clk(gclk));
	jdff dff_A_CJmFnuZt5_0(.dout(w_dff_A_O5pdFJEe5_0),.din(w_dff_A_CJmFnuZt5_0),.clk(gclk));
	jdff dff_A_O5pdFJEe5_0(.dout(w_dff_A_ft8TwJPZ9_0),.din(w_dff_A_O5pdFJEe5_0),.clk(gclk));
	jdff dff_A_ft8TwJPZ9_0(.dout(w_dff_A_HxNumhOn6_0),.din(w_dff_A_ft8TwJPZ9_0),.clk(gclk));
	jdff dff_A_HxNumhOn6_0(.dout(w_dff_A_jIooTm9d3_0),.din(w_dff_A_HxNumhOn6_0),.clk(gclk));
	jdff dff_A_jIooTm9d3_0(.dout(w_dff_A_i9vGzzLv4_0),.din(w_dff_A_jIooTm9d3_0),.clk(gclk));
	jdff dff_A_i9vGzzLv4_0(.dout(w_dff_A_3lJLA2Yt9_0),.din(w_dff_A_i9vGzzLv4_0),.clk(gclk));
	jdff dff_A_3lJLA2Yt9_0(.dout(w_dff_A_9VrcpKBu3_0),.din(w_dff_A_3lJLA2Yt9_0),.clk(gclk));
	jdff dff_A_9VrcpKBu3_0(.dout(w_dff_A_XYftsUyd9_0),.din(w_dff_A_9VrcpKBu3_0),.clk(gclk));
	jdff dff_A_XYftsUyd9_0(.dout(w_dff_A_ocGg1ky89_0),.din(w_dff_A_XYftsUyd9_0),.clk(gclk));
	jdff dff_A_ocGg1ky89_0(.dout(w_dff_A_vi0nIyCM3_0),.din(w_dff_A_ocGg1ky89_0),.clk(gclk));
	jdff dff_A_vi0nIyCM3_0(.dout(w_dff_A_RnnA6yeb6_0),.din(w_dff_A_vi0nIyCM3_0),.clk(gclk));
	jdff dff_A_RnnA6yeb6_0(.dout(w_dff_A_6OnaoYbA1_0),.din(w_dff_A_RnnA6yeb6_0),.clk(gclk));
	jdff dff_A_6OnaoYbA1_0(.dout(w_dff_A_3b6lSHj47_0),.din(w_dff_A_6OnaoYbA1_0),.clk(gclk));
	jdff dff_A_3b6lSHj47_0(.dout(w_dff_A_qzTRnjzg0_0),.din(w_dff_A_3b6lSHj47_0),.clk(gclk));
	jdff dff_A_qzTRnjzg0_0(.dout(w_dff_A_3ViHq50n9_0),.din(w_dff_A_qzTRnjzg0_0),.clk(gclk));
	jdff dff_A_3ViHq50n9_0(.dout(w_dff_A_eNBB4EP73_0),.din(w_dff_A_3ViHq50n9_0),.clk(gclk));
	jdff dff_A_eNBB4EP73_0(.dout(w_dff_A_5oXrXCIH3_0),.din(w_dff_A_eNBB4EP73_0),.clk(gclk));
	jdff dff_A_5oXrXCIH3_0(.dout(w_dff_A_TOVy9fie3_0),.din(w_dff_A_5oXrXCIH3_0),.clk(gclk));
	jdff dff_A_TOVy9fie3_0(.dout(w_dff_A_f6Dq06jn3_0),.din(w_dff_A_TOVy9fie3_0),.clk(gclk));
	jdff dff_A_f6Dq06jn3_0(.dout(w_dff_A_4ZkwPbzT3_0),.din(w_dff_A_f6Dq06jn3_0),.clk(gclk));
	jdff dff_A_4ZkwPbzT3_0(.dout(w_dff_A_S1q3s3Fz0_0),.din(w_dff_A_4ZkwPbzT3_0),.clk(gclk));
	jdff dff_A_S1q3s3Fz0_0(.dout(w_dff_A_eLE1IRuJ8_0),.din(w_dff_A_S1q3s3Fz0_0),.clk(gclk));
	jdff dff_A_eLE1IRuJ8_0(.dout(w_dff_A_bGLybw8o0_0),.din(w_dff_A_eLE1IRuJ8_0),.clk(gclk));
	jdff dff_A_bGLybw8o0_0(.dout(w_dff_A_DbqWJFSd7_0),.din(w_dff_A_bGLybw8o0_0),.clk(gclk));
	jdff dff_A_DbqWJFSd7_0(.dout(w_dff_A_vfZVeqtS2_0),.din(w_dff_A_DbqWJFSd7_0),.clk(gclk));
	jdff dff_A_vfZVeqtS2_0(.dout(w_dff_A_gO82Gl7T1_0),.din(w_dff_A_vfZVeqtS2_0),.clk(gclk));
	jdff dff_A_gO82Gl7T1_0(.dout(w_dff_A_2Aa8zRq84_0),.din(w_dff_A_gO82Gl7T1_0),.clk(gclk));
	jdff dff_A_2Aa8zRq84_0(.dout(w_dff_A_Qta0xbLt4_0),.din(w_dff_A_2Aa8zRq84_0),.clk(gclk));
	jdff dff_A_Qta0xbLt4_0(.dout(sin5),.din(w_dff_A_Qta0xbLt4_0),.clk(gclk));
	jdff dff_A_y6UHYdvt4_2(.dout(w_dff_A_VSczgI9a5_0),.din(w_dff_A_y6UHYdvt4_2),.clk(gclk));
	jdff dff_A_VSczgI9a5_0(.dout(w_dff_A_Cd928ia36_0),.din(w_dff_A_VSczgI9a5_0),.clk(gclk));
	jdff dff_A_Cd928ia36_0(.dout(w_dff_A_V4ucMXfr3_0),.din(w_dff_A_Cd928ia36_0),.clk(gclk));
	jdff dff_A_V4ucMXfr3_0(.dout(w_dff_A_PghwdNzX0_0),.din(w_dff_A_V4ucMXfr3_0),.clk(gclk));
	jdff dff_A_PghwdNzX0_0(.dout(w_dff_A_CZT15yUT9_0),.din(w_dff_A_PghwdNzX0_0),.clk(gclk));
	jdff dff_A_CZT15yUT9_0(.dout(w_dff_A_XWStr6gT2_0),.din(w_dff_A_CZT15yUT9_0),.clk(gclk));
	jdff dff_A_XWStr6gT2_0(.dout(w_dff_A_njAZfeca5_0),.din(w_dff_A_XWStr6gT2_0),.clk(gclk));
	jdff dff_A_njAZfeca5_0(.dout(w_dff_A_nGr7frN61_0),.din(w_dff_A_njAZfeca5_0),.clk(gclk));
	jdff dff_A_nGr7frN61_0(.dout(w_dff_A_BX1N2P5a4_0),.din(w_dff_A_nGr7frN61_0),.clk(gclk));
	jdff dff_A_BX1N2P5a4_0(.dout(w_dff_A_vLHec2pN9_0),.din(w_dff_A_BX1N2P5a4_0),.clk(gclk));
	jdff dff_A_vLHec2pN9_0(.dout(w_dff_A_fiV0BgNN1_0),.din(w_dff_A_vLHec2pN9_0),.clk(gclk));
	jdff dff_A_fiV0BgNN1_0(.dout(w_dff_A_yuT1EXrx2_0),.din(w_dff_A_fiV0BgNN1_0),.clk(gclk));
	jdff dff_A_yuT1EXrx2_0(.dout(w_dff_A_2xevLxyK6_0),.din(w_dff_A_yuT1EXrx2_0),.clk(gclk));
	jdff dff_A_2xevLxyK6_0(.dout(w_dff_A_lFASKJbU0_0),.din(w_dff_A_2xevLxyK6_0),.clk(gclk));
	jdff dff_A_lFASKJbU0_0(.dout(w_dff_A_GKPY07cg4_0),.din(w_dff_A_lFASKJbU0_0),.clk(gclk));
	jdff dff_A_GKPY07cg4_0(.dout(w_dff_A_jAOyFJTn7_0),.din(w_dff_A_GKPY07cg4_0),.clk(gclk));
	jdff dff_A_jAOyFJTn7_0(.dout(w_dff_A_d8IGNN0A8_0),.din(w_dff_A_jAOyFJTn7_0),.clk(gclk));
	jdff dff_A_d8IGNN0A8_0(.dout(w_dff_A_MYDDFt994_0),.din(w_dff_A_d8IGNN0A8_0),.clk(gclk));
	jdff dff_A_MYDDFt994_0(.dout(w_dff_A_TJnfdsga9_0),.din(w_dff_A_MYDDFt994_0),.clk(gclk));
	jdff dff_A_TJnfdsga9_0(.dout(w_dff_A_UVY9Iozz4_0),.din(w_dff_A_TJnfdsga9_0),.clk(gclk));
	jdff dff_A_UVY9Iozz4_0(.dout(w_dff_A_9FAIB4Ar5_0),.din(w_dff_A_UVY9Iozz4_0),.clk(gclk));
	jdff dff_A_9FAIB4Ar5_0(.dout(w_dff_A_0p8MIe4W5_0),.din(w_dff_A_9FAIB4Ar5_0),.clk(gclk));
	jdff dff_A_0p8MIe4W5_0(.dout(w_dff_A_Gx0IniJa7_0),.din(w_dff_A_0p8MIe4W5_0),.clk(gclk));
	jdff dff_A_Gx0IniJa7_0(.dout(w_dff_A_0CRCesfm7_0),.din(w_dff_A_Gx0IniJa7_0),.clk(gclk));
	jdff dff_A_0CRCesfm7_0(.dout(w_dff_A_A3uCyWZb8_0),.din(w_dff_A_0CRCesfm7_0),.clk(gclk));
	jdff dff_A_A3uCyWZb8_0(.dout(w_dff_A_tULTtL3L6_0),.din(w_dff_A_A3uCyWZb8_0),.clk(gclk));
	jdff dff_A_tULTtL3L6_0(.dout(w_dff_A_TSzkUqFK7_0),.din(w_dff_A_tULTtL3L6_0),.clk(gclk));
	jdff dff_A_TSzkUqFK7_0(.dout(w_dff_A_6XgM8n5L3_0),.din(w_dff_A_TSzkUqFK7_0),.clk(gclk));
	jdff dff_A_6XgM8n5L3_0(.dout(w_dff_A_Bka5OWbA6_0),.din(w_dff_A_6XgM8n5L3_0),.clk(gclk));
	jdff dff_A_Bka5OWbA6_0(.dout(w_dff_A_Ybo2tHbZ1_0),.din(w_dff_A_Bka5OWbA6_0),.clk(gclk));
	jdff dff_A_Ybo2tHbZ1_0(.dout(w_dff_A_Wg5zbNkE5_0),.din(w_dff_A_Ybo2tHbZ1_0),.clk(gclk));
	jdff dff_A_Wg5zbNkE5_0(.dout(sin6),.din(w_dff_A_Wg5zbNkE5_0),.clk(gclk));
	jdff dff_A_RryB5Bx36_2(.dout(w_dff_A_2q2xAQeC6_0),.din(w_dff_A_RryB5Bx36_2),.clk(gclk));
	jdff dff_A_2q2xAQeC6_0(.dout(w_dff_A_ZPXUbUTb3_0),.din(w_dff_A_2q2xAQeC6_0),.clk(gclk));
	jdff dff_A_ZPXUbUTb3_0(.dout(w_dff_A_nxCr2dCa0_0),.din(w_dff_A_ZPXUbUTb3_0),.clk(gclk));
	jdff dff_A_nxCr2dCa0_0(.dout(w_dff_A_WVoKf6jI4_0),.din(w_dff_A_nxCr2dCa0_0),.clk(gclk));
	jdff dff_A_WVoKf6jI4_0(.dout(w_dff_A_yeK30YaD2_0),.din(w_dff_A_WVoKf6jI4_0),.clk(gclk));
	jdff dff_A_yeK30YaD2_0(.dout(w_dff_A_k6gT5kZQ2_0),.din(w_dff_A_yeK30YaD2_0),.clk(gclk));
	jdff dff_A_k6gT5kZQ2_0(.dout(w_dff_A_5oEVdd244_0),.din(w_dff_A_k6gT5kZQ2_0),.clk(gclk));
	jdff dff_A_5oEVdd244_0(.dout(w_dff_A_smd1EMQt4_0),.din(w_dff_A_5oEVdd244_0),.clk(gclk));
	jdff dff_A_smd1EMQt4_0(.dout(w_dff_A_NxAkp4N11_0),.din(w_dff_A_smd1EMQt4_0),.clk(gclk));
	jdff dff_A_NxAkp4N11_0(.dout(w_dff_A_7xEYWvSz5_0),.din(w_dff_A_NxAkp4N11_0),.clk(gclk));
	jdff dff_A_7xEYWvSz5_0(.dout(w_dff_A_A5UiPDDN7_0),.din(w_dff_A_7xEYWvSz5_0),.clk(gclk));
	jdff dff_A_A5UiPDDN7_0(.dout(w_dff_A_gAbQAD9q5_0),.din(w_dff_A_A5UiPDDN7_0),.clk(gclk));
	jdff dff_A_gAbQAD9q5_0(.dout(w_dff_A_1OxsGPe50_0),.din(w_dff_A_gAbQAD9q5_0),.clk(gclk));
	jdff dff_A_1OxsGPe50_0(.dout(w_dff_A_jh7oYIIn3_0),.din(w_dff_A_1OxsGPe50_0),.clk(gclk));
	jdff dff_A_jh7oYIIn3_0(.dout(w_dff_A_axZCnYeL3_0),.din(w_dff_A_jh7oYIIn3_0),.clk(gclk));
	jdff dff_A_axZCnYeL3_0(.dout(w_dff_A_jeRq0WL24_0),.din(w_dff_A_axZCnYeL3_0),.clk(gclk));
	jdff dff_A_jeRq0WL24_0(.dout(w_dff_A_hp2rcP6N9_0),.din(w_dff_A_jeRq0WL24_0),.clk(gclk));
	jdff dff_A_hp2rcP6N9_0(.dout(w_dff_A_GhLQdO0E4_0),.din(w_dff_A_hp2rcP6N9_0),.clk(gclk));
	jdff dff_A_GhLQdO0E4_0(.dout(w_dff_A_BRkMEQ5r8_0),.din(w_dff_A_GhLQdO0E4_0),.clk(gclk));
	jdff dff_A_BRkMEQ5r8_0(.dout(w_dff_A_JxBDSVW62_0),.din(w_dff_A_BRkMEQ5r8_0),.clk(gclk));
	jdff dff_A_JxBDSVW62_0(.dout(w_dff_A_4mf4bNWe1_0),.din(w_dff_A_JxBDSVW62_0),.clk(gclk));
	jdff dff_A_4mf4bNWe1_0(.dout(w_dff_A_HTcJQbg33_0),.din(w_dff_A_4mf4bNWe1_0),.clk(gclk));
	jdff dff_A_HTcJQbg33_0(.dout(w_dff_A_IZfYf7nS2_0),.din(w_dff_A_HTcJQbg33_0),.clk(gclk));
	jdff dff_A_IZfYf7nS2_0(.dout(w_dff_A_LjAx4rqT4_0),.din(w_dff_A_IZfYf7nS2_0),.clk(gclk));
	jdff dff_A_LjAx4rqT4_0(.dout(w_dff_A_chrLxxQm0_0),.din(w_dff_A_LjAx4rqT4_0),.clk(gclk));
	jdff dff_A_chrLxxQm0_0(.dout(w_dff_A_6DcrJCLa9_0),.din(w_dff_A_chrLxxQm0_0),.clk(gclk));
	jdff dff_A_6DcrJCLa9_0(.dout(w_dff_A_09szml5I4_0),.din(w_dff_A_6DcrJCLa9_0),.clk(gclk));
	jdff dff_A_09szml5I4_0(.dout(w_dff_A_vFVYQM431_0),.din(w_dff_A_09szml5I4_0),.clk(gclk));
	jdff dff_A_vFVYQM431_0(.dout(w_dff_A_jfDZfkmv1_0),.din(w_dff_A_vFVYQM431_0),.clk(gclk));
	jdff dff_A_jfDZfkmv1_0(.dout(sin7),.din(w_dff_A_jfDZfkmv1_0),.clk(gclk));
	jdff dff_A_bZHWsZ3E8_2(.dout(w_dff_A_SA1CQeSI7_0),.din(w_dff_A_bZHWsZ3E8_2),.clk(gclk));
	jdff dff_A_SA1CQeSI7_0(.dout(w_dff_A_vFywo5td6_0),.din(w_dff_A_SA1CQeSI7_0),.clk(gclk));
	jdff dff_A_vFywo5td6_0(.dout(w_dff_A_7q9XyUWj2_0),.din(w_dff_A_vFywo5td6_0),.clk(gclk));
	jdff dff_A_7q9XyUWj2_0(.dout(w_dff_A_4hASwI6f9_0),.din(w_dff_A_7q9XyUWj2_0),.clk(gclk));
	jdff dff_A_4hASwI6f9_0(.dout(w_dff_A_Ydyk6nff2_0),.din(w_dff_A_4hASwI6f9_0),.clk(gclk));
	jdff dff_A_Ydyk6nff2_0(.dout(w_dff_A_azSuLj7Q9_0),.din(w_dff_A_Ydyk6nff2_0),.clk(gclk));
	jdff dff_A_azSuLj7Q9_0(.dout(w_dff_A_Sz0SlQX26_0),.din(w_dff_A_azSuLj7Q9_0),.clk(gclk));
	jdff dff_A_Sz0SlQX26_0(.dout(w_dff_A_YkPWNupc7_0),.din(w_dff_A_Sz0SlQX26_0),.clk(gclk));
	jdff dff_A_YkPWNupc7_0(.dout(w_dff_A_I3sfRKQf6_0),.din(w_dff_A_YkPWNupc7_0),.clk(gclk));
	jdff dff_A_I3sfRKQf6_0(.dout(w_dff_A_DksUjKGx6_0),.din(w_dff_A_I3sfRKQf6_0),.clk(gclk));
	jdff dff_A_DksUjKGx6_0(.dout(w_dff_A_zgn3vwlh0_0),.din(w_dff_A_DksUjKGx6_0),.clk(gclk));
	jdff dff_A_zgn3vwlh0_0(.dout(w_dff_A_wxl2hvhu1_0),.din(w_dff_A_zgn3vwlh0_0),.clk(gclk));
	jdff dff_A_wxl2hvhu1_0(.dout(w_dff_A_j0UnreYl0_0),.din(w_dff_A_wxl2hvhu1_0),.clk(gclk));
	jdff dff_A_j0UnreYl0_0(.dout(w_dff_A_v7jindob5_0),.din(w_dff_A_j0UnreYl0_0),.clk(gclk));
	jdff dff_A_v7jindob5_0(.dout(w_dff_A_NCarShOt9_0),.din(w_dff_A_v7jindob5_0),.clk(gclk));
	jdff dff_A_NCarShOt9_0(.dout(w_dff_A_TMW7sxXM8_0),.din(w_dff_A_NCarShOt9_0),.clk(gclk));
	jdff dff_A_TMW7sxXM8_0(.dout(w_dff_A_h6szTUnb4_0),.din(w_dff_A_TMW7sxXM8_0),.clk(gclk));
	jdff dff_A_h6szTUnb4_0(.dout(w_dff_A_y4WB1Hpz1_0),.din(w_dff_A_h6szTUnb4_0),.clk(gclk));
	jdff dff_A_y4WB1Hpz1_0(.dout(w_dff_A_hblJQGDh8_0),.din(w_dff_A_y4WB1Hpz1_0),.clk(gclk));
	jdff dff_A_hblJQGDh8_0(.dout(w_dff_A_sIfycOJl3_0),.din(w_dff_A_hblJQGDh8_0),.clk(gclk));
	jdff dff_A_sIfycOJl3_0(.dout(w_dff_A_UoyzXXtz8_0),.din(w_dff_A_sIfycOJl3_0),.clk(gclk));
	jdff dff_A_UoyzXXtz8_0(.dout(w_dff_A_B20mjgdN9_0),.din(w_dff_A_UoyzXXtz8_0),.clk(gclk));
	jdff dff_A_B20mjgdN9_0(.dout(w_dff_A_7Mrz7gZ40_0),.din(w_dff_A_B20mjgdN9_0),.clk(gclk));
	jdff dff_A_7Mrz7gZ40_0(.dout(w_dff_A_1qMKwhEQ7_0),.din(w_dff_A_7Mrz7gZ40_0),.clk(gclk));
	jdff dff_A_1qMKwhEQ7_0(.dout(w_dff_A_I4JQ4Did4_0),.din(w_dff_A_1qMKwhEQ7_0),.clk(gclk));
	jdff dff_A_I4JQ4Did4_0(.dout(w_dff_A_7NuQY5cf0_0),.din(w_dff_A_I4JQ4Did4_0),.clk(gclk));
	jdff dff_A_7NuQY5cf0_0(.dout(w_dff_A_wIweRCIZ6_0),.din(w_dff_A_7NuQY5cf0_0),.clk(gclk));
	jdff dff_A_wIweRCIZ6_0(.dout(sin8),.din(w_dff_A_wIweRCIZ6_0),.clk(gclk));
	jdff dff_A_u8ZD7jxR4_2(.dout(w_dff_A_xIjmN53W8_0),.din(w_dff_A_u8ZD7jxR4_2),.clk(gclk));
	jdff dff_A_xIjmN53W8_0(.dout(w_dff_A_VvJfRlVy1_0),.din(w_dff_A_xIjmN53W8_0),.clk(gclk));
	jdff dff_A_VvJfRlVy1_0(.dout(w_dff_A_rpnuCX2m3_0),.din(w_dff_A_VvJfRlVy1_0),.clk(gclk));
	jdff dff_A_rpnuCX2m3_0(.dout(w_dff_A_en97lUwR2_0),.din(w_dff_A_rpnuCX2m3_0),.clk(gclk));
	jdff dff_A_en97lUwR2_0(.dout(w_dff_A_lTJkpVQQ7_0),.din(w_dff_A_en97lUwR2_0),.clk(gclk));
	jdff dff_A_lTJkpVQQ7_0(.dout(w_dff_A_TPzfFAbM5_0),.din(w_dff_A_lTJkpVQQ7_0),.clk(gclk));
	jdff dff_A_TPzfFAbM5_0(.dout(w_dff_A_WY9GZPqX7_0),.din(w_dff_A_TPzfFAbM5_0),.clk(gclk));
	jdff dff_A_WY9GZPqX7_0(.dout(w_dff_A_J19n05Kp8_0),.din(w_dff_A_WY9GZPqX7_0),.clk(gclk));
	jdff dff_A_J19n05Kp8_0(.dout(w_dff_A_uY42FFpW9_0),.din(w_dff_A_J19n05Kp8_0),.clk(gclk));
	jdff dff_A_uY42FFpW9_0(.dout(w_dff_A_EorRc6GK5_0),.din(w_dff_A_uY42FFpW9_0),.clk(gclk));
	jdff dff_A_EorRc6GK5_0(.dout(w_dff_A_UTAfM9Ld6_0),.din(w_dff_A_EorRc6GK5_0),.clk(gclk));
	jdff dff_A_UTAfM9Ld6_0(.dout(w_dff_A_WoguPPsq8_0),.din(w_dff_A_UTAfM9Ld6_0),.clk(gclk));
	jdff dff_A_WoguPPsq8_0(.dout(w_dff_A_wTXLXwnW0_0),.din(w_dff_A_WoguPPsq8_0),.clk(gclk));
	jdff dff_A_wTXLXwnW0_0(.dout(w_dff_A_eIlvoaGs8_0),.din(w_dff_A_wTXLXwnW0_0),.clk(gclk));
	jdff dff_A_eIlvoaGs8_0(.dout(w_dff_A_W7ALtZPI5_0),.din(w_dff_A_eIlvoaGs8_0),.clk(gclk));
	jdff dff_A_W7ALtZPI5_0(.dout(w_dff_A_zHaN7Vux1_0),.din(w_dff_A_W7ALtZPI5_0),.clk(gclk));
	jdff dff_A_zHaN7Vux1_0(.dout(w_dff_A_TbGOdZon0_0),.din(w_dff_A_zHaN7Vux1_0),.clk(gclk));
	jdff dff_A_TbGOdZon0_0(.dout(w_dff_A_4lwN3GCC4_0),.din(w_dff_A_TbGOdZon0_0),.clk(gclk));
	jdff dff_A_4lwN3GCC4_0(.dout(w_dff_A_LDf80yb75_0),.din(w_dff_A_4lwN3GCC4_0),.clk(gclk));
	jdff dff_A_LDf80yb75_0(.dout(w_dff_A_w5dAdQPn1_0),.din(w_dff_A_LDf80yb75_0),.clk(gclk));
	jdff dff_A_w5dAdQPn1_0(.dout(w_dff_A_toEoJcX35_0),.din(w_dff_A_w5dAdQPn1_0),.clk(gclk));
	jdff dff_A_toEoJcX35_0(.dout(w_dff_A_TzyBSbEB7_0),.din(w_dff_A_toEoJcX35_0),.clk(gclk));
	jdff dff_A_TzyBSbEB7_0(.dout(w_dff_A_hkJdPfo42_0),.din(w_dff_A_TzyBSbEB7_0),.clk(gclk));
	jdff dff_A_hkJdPfo42_0(.dout(w_dff_A_SzG6izqJ5_0),.din(w_dff_A_hkJdPfo42_0),.clk(gclk));
	jdff dff_A_SzG6izqJ5_0(.dout(w_dff_A_Wh7Nsh6u6_0),.din(w_dff_A_SzG6izqJ5_0),.clk(gclk));
	jdff dff_A_Wh7Nsh6u6_0(.dout(sin9),.din(w_dff_A_Wh7Nsh6u6_0),.clk(gclk));
	jdff dff_A_SP0xCeW41_2(.dout(w_dff_A_zCw8m8dq0_0),.din(w_dff_A_SP0xCeW41_2),.clk(gclk));
	jdff dff_A_zCw8m8dq0_0(.dout(w_dff_A_wcuoHtPZ2_0),.din(w_dff_A_zCw8m8dq0_0),.clk(gclk));
	jdff dff_A_wcuoHtPZ2_0(.dout(w_dff_A_cBxi1A4y6_0),.din(w_dff_A_wcuoHtPZ2_0),.clk(gclk));
	jdff dff_A_cBxi1A4y6_0(.dout(w_dff_A_zNCMFdRD3_0),.din(w_dff_A_cBxi1A4y6_0),.clk(gclk));
	jdff dff_A_zNCMFdRD3_0(.dout(w_dff_A_6w1qM55O1_0),.din(w_dff_A_zNCMFdRD3_0),.clk(gclk));
	jdff dff_A_6w1qM55O1_0(.dout(w_dff_A_j4gC81zA6_0),.din(w_dff_A_6w1qM55O1_0),.clk(gclk));
	jdff dff_A_j4gC81zA6_0(.dout(w_dff_A_jAlXBA9k3_0),.din(w_dff_A_j4gC81zA6_0),.clk(gclk));
	jdff dff_A_jAlXBA9k3_0(.dout(w_dff_A_mboHtXUS9_0),.din(w_dff_A_jAlXBA9k3_0),.clk(gclk));
	jdff dff_A_mboHtXUS9_0(.dout(w_dff_A_kx82cDBm4_0),.din(w_dff_A_mboHtXUS9_0),.clk(gclk));
	jdff dff_A_kx82cDBm4_0(.dout(w_dff_A_5NLq3L9W2_0),.din(w_dff_A_kx82cDBm4_0),.clk(gclk));
	jdff dff_A_5NLq3L9W2_0(.dout(w_dff_A_N3M452Qp5_0),.din(w_dff_A_5NLq3L9W2_0),.clk(gclk));
	jdff dff_A_N3M452Qp5_0(.dout(w_dff_A_20zhR8K87_0),.din(w_dff_A_N3M452Qp5_0),.clk(gclk));
	jdff dff_A_20zhR8K87_0(.dout(w_dff_A_nIeJ6drv6_0),.din(w_dff_A_20zhR8K87_0),.clk(gclk));
	jdff dff_A_nIeJ6drv6_0(.dout(w_dff_A_fFimfUza6_0),.din(w_dff_A_nIeJ6drv6_0),.clk(gclk));
	jdff dff_A_fFimfUza6_0(.dout(w_dff_A_Agh7AKyL0_0),.din(w_dff_A_fFimfUza6_0),.clk(gclk));
	jdff dff_A_Agh7AKyL0_0(.dout(w_dff_A_oH248Y4P4_0),.din(w_dff_A_Agh7AKyL0_0),.clk(gclk));
	jdff dff_A_oH248Y4P4_0(.dout(w_dff_A_81AFO8ut4_0),.din(w_dff_A_oH248Y4P4_0),.clk(gclk));
	jdff dff_A_81AFO8ut4_0(.dout(w_dff_A_xE382PUD8_0),.din(w_dff_A_81AFO8ut4_0),.clk(gclk));
	jdff dff_A_xE382PUD8_0(.dout(w_dff_A_WiLblRlj2_0),.din(w_dff_A_xE382PUD8_0),.clk(gclk));
	jdff dff_A_WiLblRlj2_0(.dout(w_dff_A_mXqmIs4H4_0),.din(w_dff_A_WiLblRlj2_0),.clk(gclk));
	jdff dff_A_mXqmIs4H4_0(.dout(w_dff_A_Dg6kfu2O1_0),.din(w_dff_A_mXqmIs4H4_0),.clk(gclk));
	jdff dff_A_Dg6kfu2O1_0(.dout(w_dff_A_rziDBC9L5_0),.din(w_dff_A_Dg6kfu2O1_0),.clk(gclk));
	jdff dff_A_rziDBC9L5_0(.dout(w_dff_A_S10WfadL7_0),.din(w_dff_A_rziDBC9L5_0),.clk(gclk));
	jdff dff_A_S10WfadL7_0(.dout(sin10),.din(w_dff_A_S10WfadL7_0),.clk(gclk));
	jdff dff_A_gP8OwZoN2_2(.dout(w_dff_A_vYEU9rof4_0),.din(w_dff_A_gP8OwZoN2_2),.clk(gclk));
	jdff dff_A_vYEU9rof4_0(.dout(w_dff_A_cmBoHTo26_0),.din(w_dff_A_vYEU9rof4_0),.clk(gclk));
	jdff dff_A_cmBoHTo26_0(.dout(w_dff_A_xZ2zrSHd7_0),.din(w_dff_A_cmBoHTo26_0),.clk(gclk));
	jdff dff_A_xZ2zrSHd7_0(.dout(w_dff_A_6YawxdGv6_0),.din(w_dff_A_xZ2zrSHd7_0),.clk(gclk));
	jdff dff_A_6YawxdGv6_0(.dout(w_dff_A_xWOYFBbj2_0),.din(w_dff_A_6YawxdGv6_0),.clk(gclk));
	jdff dff_A_xWOYFBbj2_0(.dout(w_dff_A_ezdOWVDX2_0),.din(w_dff_A_xWOYFBbj2_0),.clk(gclk));
	jdff dff_A_ezdOWVDX2_0(.dout(w_dff_A_Oy0RtZ3C6_0),.din(w_dff_A_ezdOWVDX2_0),.clk(gclk));
	jdff dff_A_Oy0RtZ3C6_0(.dout(w_dff_A_EkJtWrnA6_0),.din(w_dff_A_Oy0RtZ3C6_0),.clk(gclk));
	jdff dff_A_EkJtWrnA6_0(.dout(w_dff_A_R873z4GN2_0),.din(w_dff_A_EkJtWrnA6_0),.clk(gclk));
	jdff dff_A_R873z4GN2_0(.dout(w_dff_A_dKfo5FFq8_0),.din(w_dff_A_R873z4GN2_0),.clk(gclk));
	jdff dff_A_dKfo5FFq8_0(.dout(w_dff_A_euFG9zf55_0),.din(w_dff_A_dKfo5FFq8_0),.clk(gclk));
	jdff dff_A_euFG9zf55_0(.dout(w_dff_A_x39Ff9zt8_0),.din(w_dff_A_euFG9zf55_0),.clk(gclk));
	jdff dff_A_x39Ff9zt8_0(.dout(w_dff_A_meAbKCtT8_0),.din(w_dff_A_x39Ff9zt8_0),.clk(gclk));
	jdff dff_A_meAbKCtT8_0(.dout(w_dff_A_iZJ3QSDR9_0),.din(w_dff_A_meAbKCtT8_0),.clk(gclk));
	jdff dff_A_iZJ3QSDR9_0(.dout(w_dff_A_GYdczOMX1_0),.din(w_dff_A_iZJ3QSDR9_0),.clk(gclk));
	jdff dff_A_GYdczOMX1_0(.dout(w_dff_A_zaOeb0f63_0),.din(w_dff_A_GYdczOMX1_0),.clk(gclk));
	jdff dff_A_zaOeb0f63_0(.dout(w_dff_A_pwtacHqE4_0),.din(w_dff_A_zaOeb0f63_0),.clk(gclk));
	jdff dff_A_pwtacHqE4_0(.dout(w_dff_A_XuWS0maq8_0),.din(w_dff_A_pwtacHqE4_0),.clk(gclk));
	jdff dff_A_XuWS0maq8_0(.dout(w_dff_A_PYTOf91n7_0),.din(w_dff_A_XuWS0maq8_0),.clk(gclk));
	jdff dff_A_PYTOf91n7_0(.dout(w_dff_A_m7Rav7Rh8_0),.din(w_dff_A_PYTOf91n7_0),.clk(gclk));
	jdff dff_A_m7Rav7Rh8_0(.dout(w_dff_A_xyIOOBwo1_0),.din(w_dff_A_m7Rav7Rh8_0),.clk(gclk));
	jdff dff_A_xyIOOBwo1_0(.dout(sin11),.din(w_dff_A_xyIOOBwo1_0),.clk(gclk));
	jdff dff_A_5LHruE6g9_2(.dout(w_dff_A_XraBX9ax8_0),.din(w_dff_A_5LHruE6g9_2),.clk(gclk));
	jdff dff_A_XraBX9ax8_0(.dout(w_dff_A_36XP6H9o3_0),.din(w_dff_A_XraBX9ax8_0),.clk(gclk));
	jdff dff_A_36XP6H9o3_0(.dout(w_dff_A_oMdRGqlV4_0),.din(w_dff_A_36XP6H9o3_0),.clk(gclk));
	jdff dff_A_oMdRGqlV4_0(.dout(w_dff_A_jRegBd9L2_0),.din(w_dff_A_oMdRGqlV4_0),.clk(gclk));
	jdff dff_A_jRegBd9L2_0(.dout(w_dff_A_gQxxtX7L3_0),.din(w_dff_A_jRegBd9L2_0),.clk(gclk));
	jdff dff_A_gQxxtX7L3_0(.dout(w_dff_A_2G8L8kIx3_0),.din(w_dff_A_gQxxtX7L3_0),.clk(gclk));
	jdff dff_A_2G8L8kIx3_0(.dout(w_dff_A_0LDLR0aL2_0),.din(w_dff_A_2G8L8kIx3_0),.clk(gclk));
	jdff dff_A_0LDLR0aL2_0(.dout(w_dff_A_V8hz3nfq6_0),.din(w_dff_A_0LDLR0aL2_0),.clk(gclk));
	jdff dff_A_V8hz3nfq6_0(.dout(w_dff_A_KKZotsfK4_0),.din(w_dff_A_V8hz3nfq6_0),.clk(gclk));
	jdff dff_A_KKZotsfK4_0(.dout(w_dff_A_QETzy8Qf0_0),.din(w_dff_A_KKZotsfK4_0),.clk(gclk));
	jdff dff_A_QETzy8Qf0_0(.dout(w_dff_A_tC1zSLKx6_0),.din(w_dff_A_QETzy8Qf0_0),.clk(gclk));
	jdff dff_A_tC1zSLKx6_0(.dout(w_dff_A_kPOlxqHF4_0),.din(w_dff_A_tC1zSLKx6_0),.clk(gclk));
	jdff dff_A_kPOlxqHF4_0(.dout(w_dff_A_FiwSAyo31_0),.din(w_dff_A_kPOlxqHF4_0),.clk(gclk));
	jdff dff_A_FiwSAyo31_0(.dout(w_dff_A_eOmUKcvu1_0),.din(w_dff_A_FiwSAyo31_0),.clk(gclk));
	jdff dff_A_eOmUKcvu1_0(.dout(w_dff_A_FgYbu4IE2_0),.din(w_dff_A_eOmUKcvu1_0),.clk(gclk));
	jdff dff_A_FgYbu4IE2_0(.dout(w_dff_A_CX4aF0us2_0),.din(w_dff_A_FgYbu4IE2_0),.clk(gclk));
	jdff dff_A_CX4aF0us2_0(.dout(w_dff_A_Hfxu5oWq8_0),.din(w_dff_A_CX4aF0us2_0),.clk(gclk));
	jdff dff_A_Hfxu5oWq8_0(.dout(w_dff_A_btSXAvG23_0),.din(w_dff_A_Hfxu5oWq8_0),.clk(gclk));
	jdff dff_A_btSXAvG23_0(.dout(w_dff_A_QWZuBYSD7_0),.din(w_dff_A_btSXAvG23_0),.clk(gclk));
	jdff dff_A_QWZuBYSD7_0(.dout(sin12),.din(w_dff_A_QWZuBYSD7_0),.clk(gclk));
	jdff dff_A_oxEVAVgt4_2(.dout(w_dff_A_FPVKDFJ45_0),.din(w_dff_A_oxEVAVgt4_2),.clk(gclk));
	jdff dff_A_FPVKDFJ45_0(.dout(w_dff_A_ToSWAq2x5_0),.din(w_dff_A_FPVKDFJ45_0),.clk(gclk));
	jdff dff_A_ToSWAq2x5_0(.dout(w_dff_A_wM0OhjKk0_0),.din(w_dff_A_ToSWAq2x5_0),.clk(gclk));
	jdff dff_A_wM0OhjKk0_0(.dout(w_dff_A_V9Yf3nlK6_0),.din(w_dff_A_wM0OhjKk0_0),.clk(gclk));
	jdff dff_A_V9Yf3nlK6_0(.dout(w_dff_A_bHPpDfnj2_0),.din(w_dff_A_V9Yf3nlK6_0),.clk(gclk));
	jdff dff_A_bHPpDfnj2_0(.dout(w_dff_A_J67J2Nt24_0),.din(w_dff_A_bHPpDfnj2_0),.clk(gclk));
	jdff dff_A_J67J2Nt24_0(.dout(w_dff_A_Y5IUSRh22_0),.din(w_dff_A_J67J2Nt24_0),.clk(gclk));
	jdff dff_A_Y5IUSRh22_0(.dout(w_dff_A_WUHuYyqG9_0),.din(w_dff_A_Y5IUSRh22_0),.clk(gclk));
	jdff dff_A_WUHuYyqG9_0(.dout(w_dff_A_9w0Xae3d8_0),.din(w_dff_A_WUHuYyqG9_0),.clk(gclk));
	jdff dff_A_9w0Xae3d8_0(.dout(w_dff_A_PoAdZYf43_0),.din(w_dff_A_9w0Xae3d8_0),.clk(gclk));
	jdff dff_A_PoAdZYf43_0(.dout(w_dff_A_NfoXnuL88_0),.din(w_dff_A_PoAdZYf43_0),.clk(gclk));
	jdff dff_A_NfoXnuL88_0(.dout(w_dff_A_o6vZFeEC2_0),.din(w_dff_A_NfoXnuL88_0),.clk(gclk));
	jdff dff_A_o6vZFeEC2_0(.dout(w_dff_A_wAH8io2v1_0),.din(w_dff_A_o6vZFeEC2_0),.clk(gclk));
	jdff dff_A_wAH8io2v1_0(.dout(w_dff_A_ywLq8MK66_0),.din(w_dff_A_wAH8io2v1_0),.clk(gclk));
	jdff dff_A_ywLq8MK66_0(.dout(w_dff_A_u4gMFVF98_0),.din(w_dff_A_ywLq8MK66_0),.clk(gclk));
	jdff dff_A_u4gMFVF98_0(.dout(w_dff_A_Ge9anYdW7_0),.din(w_dff_A_u4gMFVF98_0),.clk(gclk));
	jdff dff_A_Ge9anYdW7_0(.dout(w_dff_A_OOy7QXUP8_0),.din(w_dff_A_Ge9anYdW7_0),.clk(gclk));
	jdff dff_A_OOy7QXUP8_0(.dout(sin13),.din(w_dff_A_OOy7QXUP8_0),.clk(gclk));
	jdff dff_A_CHdzBFmi0_2(.dout(w_dff_A_UnU6ipts8_0),.din(w_dff_A_CHdzBFmi0_2),.clk(gclk));
	jdff dff_A_UnU6ipts8_0(.dout(w_dff_A_URYwyff68_0),.din(w_dff_A_UnU6ipts8_0),.clk(gclk));
	jdff dff_A_URYwyff68_0(.dout(w_dff_A_DJO6BGWh1_0),.din(w_dff_A_URYwyff68_0),.clk(gclk));
	jdff dff_A_DJO6BGWh1_0(.dout(w_dff_A_XK0V8Yav0_0),.din(w_dff_A_DJO6BGWh1_0),.clk(gclk));
	jdff dff_A_XK0V8Yav0_0(.dout(w_dff_A_lrIuidol1_0),.din(w_dff_A_XK0V8Yav0_0),.clk(gclk));
	jdff dff_A_lrIuidol1_0(.dout(w_dff_A_8k3b3W493_0),.din(w_dff_A_lrIuidol1_0),.clk(gclk));
	jdff dff_A_8k3b3W493_0(.dout(w_dff_A_scJTSTg71_0),.din(w_dff_A_8k3b3W493_0),.clk(gclk));
	jdff dff_A_scJTSTg71_0(.dout(w_dff_A_X5d0iTYj7_0),.din(w_dff_A_scJTSTg71_0),.clk(gclk));
	jdff dff_A_X5d0iTYj7_0(.dout(w_dff_A_yaIwIwEV5_0),.din(w_dff_A_X5d0iTYj7_0),.clk(gclk));
	jdff dff_A_yaIwIwEV5_0(.dout(w_dff_A_mp6WrrJI0_0),.din(w_dff_A_yaIwIwEV5_0),.clk(gclk));
	jdff dff_A_mp6WrrJI0_0(.dout(w_dff_A_wFhcnsMx3_0),.din(w_dff_A_mp6WrrJI0_0),.clk(gclk));
	jdff dff_A_wFhcnsMx3_0(.dout(w_dff_A_xzfUSp979_0),.din(w_dff_A_wFhcnsMx3_0),.clk(gclk));
	jdff dff_A_xzfUSp979_0(.dout(w_dff_A_sdbpSfTh9_0),.din(w_dff_A_xzfUSp979_0),.clk(gclk));
	jdff dff_A_sdbpSfTh9_0(.dout(w_dff_A_8pzOy3UG5_0),.din(w_dff_A_sdbpSfTh9_0),.clk(gclk));
	jdff dff_A_8pzOy3UG5_0(.dout(w_dff_A_hEgTE9hf0_0),.din(w_dff_A_8pzOy3UG5_0),.clk(gclk));
	jdff dff_A_hEgTE9hf0_0(.dout(sin14),.din(w_dff_A_hEgTE9hf0_0),.clk(gclk));
	jdff dff_A_rLUmXsuL3_2(.dout(w_dff_A_otiGIucp1_0),.din(w_dff_A_rLUmXsuL3_2),.clk(gclk));
	jdff dff_A_otiGIucp1_0(.dout(w_dff_A_QCIAlclO5_0),.din(w_dff_A_otiGIucp1_0),.clk(gclk));
	jdff dff_A_QCIAlclO5_0(.dout(w_dff_A_PKNUWaTc8_0),.din(w_dff_A_QCIAlclO5_0),.clk(gclk));
	jdff dff_A_PKNUWaTc8_0(.dout(w_dff_A_tnvxfwEx6_0),.din(w_dff_A_PKNUWaTc8_0),.clk(gclk));
	jdff dff_A_tnvxfwEx6_0(.dout(w_dff_A_bI7eZstP8_0),.din(w_dff_A_tnvxfwEx6_0),.clk(gclk));
	jdff dff_A_bI7eZstP8_0(.dout(w_dff_A_LfD11Ul04_0),.din(w_dff_A_bI7eZstP8_0),.clk(gclk));
	jdff dff_A_LfD11Ul04_0(.dout(w_dff_A_uCEdhaHI9_0),.din(w_dff_A_LfD11Ul04_0),.clk(gclk));
	jdff dff_A_uCEdhaHI9_0(.dout(w_dff_A_VSNBlYSA8_0),.din(w_dff_A_uCEdhaHI9_0),.clk(gclk));
	jdff dff_A_VSNBlYSA8_0(.dout(w_dff_A_DunAigsW4_0),.din(w_dff_A_VSNBlYSA8_0),.clk(gclk));
	jdff dff_A_DunAigsW4_0(.dout(w_dff_A_ws1ZNx7D7_0),.din(w_dff_A_DunAigsW4_0),.clk(gclk));
	jdff dff_A_ws1ZNx7D7_0(.dout(w_dff_A_eQ2uXRjN7_0),.din(w_dff_A_ws1ZNx7D7_0),.clk(gclk));
	jdff dff_A_eQ2uXRjN7_0(.dout(w_dff_A_qkbQYpJS9_0),.din(w_dff_A_eQ2uXRjN7_0),.clk(gclk));
	jdff dff_A_qkbQYpJS9_0(.dout(w_dff_A_6w7bUJw38_0),.din(w_dff_A_qkbQYpJS9_0),.clk(gclk));
	jdff dff_A_6w7bUJw38_0(.dout(sin15),.din(w_dff_A_6w7bUJw38_0),.clk(gclk));
	jdff dff_A_J2WpamXl7_2(.dout(w_dff_A_SSc9x9V91_0),.din(w_dff_A_J2WpamXl7_2),.clk(gclk));
	jdff dff_A_SSc9x9V91_0(.dout(w_dff_A_RoJR0kUy8_0),.din(w_dff_A_SSc9x9V91_0),.clk(gclk));
	jdff dff_A_RoJR0kUy8_0(.dout(w_dff_A_VFhQUbqC4_0),.din(w_dff_A_RoJR0kUy8_0),.clk(gclk));
	jdff dff_A_VFhQUbqC4_0(.dout(w_dff_A_gKxJifTD3_0),.din(w_dff_A_VFhQUbqC4_0),.clk(gclk));
	jdff dff_A_gKxJifTD3_0(.dout(w_dff_A_zK6tjDpz5_0),.din(w_dff_A_gKxJifTD3_0),.clk(gclk));
	jdff dff_A_zK6tjDpz5_0(.dout(w_dff_A_2EczkCpu2_0),.din(w_dff_A_zK6tjDpz5_0),.clk(gclk));
	jdff dff_A_2EczkCpu2_0(.dout(w_dff_A_7dlymOGj7_0),.din(w_dff_A_2EczkCpu2_0),.clk(gclk));
	jdff dff_A_7dlymOGj7_0(.dout(w_dff_A_KcxQcDa58_0),.din(w_dff_A_7dlymOGj7_0),.clk(gclk));
	jdff dff_A_KcxQcDa58_0(.dout(w_dff_A_6qiLiz9K4_0),.din(w_dff_A_KcxQcDa58_0),.clk(gclk));
	jdff dff_A_6qiLiz9K4_0(.dout(w_dff_A_QV6JNCbe6_0),.din(w_dff_A_6qiLiz9K4_0),.clk(gclk));
	jdff dff_A_QV6JNCbe6_0(.dout(sin16),.din(w_dff_A_QV6JNCbe6_0),.clk(gclk));
	jdff dff_A_k0YYIuNo5_2(.dout(w_dff_A_7bgQ0bRC0_0),.din(w_dff_A_k0YYIuNo5_2),.clk(gclk));
	jdff dff_A_7bgQ0bRC0_0(.dout(w_dff_A_wxlMlu5M2_0),.din(w_dff_A_7bgQ0bRC0_0),.clk(gclk));
	jdff dff_A_wxlMlu5M2_0(.dout(w_dff_A_SCmN7kIq5_0),.din(w_dff_A_wxlMlu5M2_0),.clk(gclk));
	jdff dff_A_SCmN7kIq5_0(.dout(w_dff_A_GBCejgwR2_0),.din(w_dff_A_SCmN7kIq5_0),.clk(gclk));
	jdff dff_A_GBCejgwR2_0(.dout(w_dff_A_rLusq6RD4_0),.din(w_dff_A_GBCejgwR2_0),.clk(gclk));
	jdff dff_A_rLusq6RD4_0(.dout(w_dff_A_wOGxBmPA5_0),.din(w_dff_A_rLusq6RD4_0),.clk(gclk));
	jdff dff_A_wOGxBmPA5_0(.dout(w_dff_A_rqlcZPUQ3_0),.din(w_dff_A_wOGxBmPA5_0),.clk(gclk));
	jdff dff_A_rqlcZPUQ3_0(.dout(w_dff_A_wzXcXi204_0),.din(w_dff_A_rqlcZPUQ3_0),.clk(gclk));
	jdff dff_A_wzXcXi204_0(.dout(sin17),.din(w_dff_A_wzXcXi204_0),.clk(gclk));
	jdff dff_A_0nVz4h2P4_2(.dout(w_dff_A_7ztwvdHZ5_0),.din(w_dff_A_0nVz4h2P4_2),.clk(gclk));
	jdff dff_A_7ztwvdHZ5_0(.dout(w_dff_A_HxzPE9Ro9_0),.din(w_dff_A_7ztwvdHZ5_0),.clk(gclk));
	jdff dff_A_HxzPE9Ro9_0(.dout(w_dff_A_6itk3QDR1_0),.din(w_dff_A_HxzPE9Ro9_0),.clk(gclk));
	jdff dff_A_6itk3QDR1_0(.dout(w_dff_A_J1zHO9iV7_0),.din(w_dff_A_6itk3QDR1_0),.clk(gclk));
	jdff dff_A_J1zHO9iV7_0(.dout(w_dff_A_PHDW0HQK8_0),.din(w_dff_A_J1zHO9iV7_0),.clk(gclk));
	jdff dff_A_PHDW0HQK8_0(.dout(w_dff_A_cGXW2PwO3_0),.din(w_dff_A_PHDW0HQK8_0),.clk(gclk));
	jdff dff_A_cGXW2PwO3_0(.dout(sin18),.din(w_dff_A_cGXW2PwO3_0),.clk(gclk));
	jdff dff_A_Cw7elsfJ2_2(.dout(w_dff_A_SQqGAZ728_0),.din(w_dff_A_Cw7elsfJ2_2),.clk(gclk));
	jdff dff_A_SQqGAZ728_0(.dout(w_dff_A_ieToSDME3_0),.din(w_dff_A_SQqGAZ728_0),.clk(gclk));
	jdff dff_A_ieToSDME3_0(.dout(w_dff_A_r1o6n5ps1_0),.din(w_dff_A_ieToSDME3_0),.clk(gclk));
	jdff dff_A_r1o6n5ps1_0(.dout(w_dff_A_GC1Xlu628_0),.din(w_dff_A_r1o6n5ps1_0),.clk(gclk));
	jdff dff_A_GC1Xlu628_0(.dout(sin19),.din(w_dff_A_GC1Xlu628_0),.clk(gclk));
	jdff dff_A_gS2lI5Ue9_2(.dout(w_dff_A_G2ckHM4a8_0),.din(w_dff_A_gS2lI5Ue9_2),.clk(gclk));
	jdff dff_A_G2ckHM4a8_0(.dout(w_dff_A_xrK6u3Nq1_0),.din(w_dff_A_G2ckHM4a8_0),.clk(gclk));
	jdff dff_A_xrK6u3Nq1_0(.dout(w_dff_A_UG9OPTVc9_0),.din(w_dff_A_xrK6u3Nq1_0),.clk(gclk));
	jdff dff_A_UG9OPTVc9_0(.dout(sin20),.din(w_dff_A_UG9OPTVc9_0),.clk(gclk));
	jdff dff_A_TNSINLGv9_2(.dout(w_dff_A_mEOc6pxz8_0),.din(w_dff_A_TNSINLGv9_2),.clk(gclk));
	jdff dff_A_mEOc6pxz8_0(.dout(w_dff_A_S7Y49kXp0_0),.din(w_dff_A_mEOc6pxz8_0),.clk(gclk));
	jdff dff_A_S7Y49kXp0_0(.dout(sin21),.din(w_dff_A_S7Y49kXp0_0),.clk(gclk));
	jdff dff_A_HR8wY1806_2(.dout(w_dff_A_b1AKM4qo9_0),.din(w_dff_A_HR8wY1806_2),.clk(gclk));
	jdff dff_A_b1AKM4qo9_0(.dout(sin22),.din(w_dff_A_b1AKM4qo9_0),.clk(gclk));
endmodule

