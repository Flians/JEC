/*

c880:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jdff: 1147
	jand: 151
	jor: 122

Summary:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jdff: 1147
	jand: 151
	jor: 122

The maximum logic level gap of any gate:
	c880: 5
*/

module gf_c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n103;
	wire n104;
	wire n105;
	wire n107;
	wire n108;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n119;
	wire n120;
	wire n122;
	wire n123;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire[2:0] w_G1gat_0;
	wire[1:0] w_G1gat_1;
	wire[1:0] w_G8gat_0;
	wire[1:0] w_G13gat_0;
	wire[2:0] w_G17gat_0;
	wire[2:0] w_G17gat_1;
	wire[2:0] w_G17gat_2;
	wire[1:0] w_G26gat_0;
	wire[2:0] w_G29gat_0;
	wire[1:0] w_G36gat_0;
	wire[2:0] w_G42gat_0;
	wire[2:0] w_G42gat_1;
	wire[1:0] w_G42gat_2;
	wire[2:0] w_G51gat_0;
	wire[1:0] w_G51gat_1;
	wire[2:0] w_G55gat_0;
	wire[2:0] w_G59gat_0;
	wire[1:0] w_G59gat_1;
	wire[1:0] w_G68gat_0;
	wire[1:0] w_G75gat_0;
	wire[2:0] w_G80gat_0;
	wire[2:0] w_G91gat_0;
	wire[2:0] w_G96gat_0;
	wire[2:0] w_G101gat_0;
	wire[2:0] w_G106gat_0;
	wire[2:0] w_G111gat_0;
	wire[2:0] w_G116gat_0;
	wire[2:0] w_G121gat_0;
	wire[2:0] w_G126gat_0;
	wire[1:0] w_G130gat_0;
	wire[2:0] w_G138gat_0;
	wire[1:0] w_G138gat_1;
	wire[1:0] w_G143gat_0;
	wire[1:0] w_G146gat_0;
	wire[1:0] w_G149gat_0;
	wire[2:0] w_G153gat_0;
	wire[1:0] w_G156gat_0;
	wire[2:0] w_G159gat_0;
	wire[2:0] w_G159gat_1;
	wire[2:0] w_G165gat_0;
	wire[2:0] w_G165gat_1;
	wire[2:0] w_G171gat_0;
	wire[2:0] w_G171gat_1;
	wire[2:0] w_G177gat_0;
	wire[2:0] w_G177gat_1;
	wire[2:0] w_G183gat_0;
	wire[2:0] w_G183gat_1;
	wire[2:0] w_G189gat_0;
	wire[2:0] w_G189gat_1;
	wire[1:0] w_G189gat_2;
	wire[2:0] w_G195gat_0;
	wire[2:0] w_G195gat_1;
	wire[1:0] w_G195gat_2;
	wire[2:0] w_G201gat_0;
	wire[1:0] w_G201gat_1;
	wire[2:0] w_G210gat_0;
	wire[2:0] w_G210gat_1;
	wire[2:0] w_G210gat_2;
	wire[1:0] w_G210gat_3;
	wire[2:0] w_G219gat_0;
	wire[2:0] w_G219gat_1;
	wire[2:0] w_G219gat_2;
	wire[2:0] w_G219gat_3;
	wire[2:0] w_G228gat_0;
	wire[2:0] w_G228gat_1;
	wire[2:0] w_G228gat_2;
	wire[1:0] w_G228gat_3;
	wire[2:0] w_G237gat_0;
	wire[2:0] w_G237gat_1;
	wire[2:0] w_G237gat_2;
	wire[1:0] w_G237gat_3;
	wire[2:0] w_G246gat_0;
	wire[2:0] w_G246gat_1;
	wire[2:0] w_G246gat_2;
	wire[1:0] w_G246gat_3;
	wire[2:0] w_G255gat_0;
	wire[2:0] w_G261gat_0;
	wire[1:0] w_G268gat_0;
	wire[1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire[2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire[1:0] w_n86_0;
	wire[1:0] w_n88_0;
	wire[1:0] w_n92_0;
	wire[1:0] w_n93_0;
	wire[2:0] w_n95_0;
	wire[1:0] w_n97_0;
	wire[1:0] w_n99_0;
	wire[1:0] w_n101_0;
	wire[1:0] w_n103_0;
	wire[1:0] w_n104_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n109_0;
	wire[1:0] w_n111_0;
	wire[1:0] w_n113_0;
	wire[2:0] w_n119_0;
	wire[1:0] w_n122_0;
	wire[1:0] w_n144_0;
	wire[1:0] w_n146_0;
	wire[2:0] w_n148_0;
	wire[2:0] w_n148_1;
	wire[1:0] w_n149_0;
	wire[1:0] w_n151_0;
	wire[1:0] w_n152_0;
	wire[1:0] w_n162_0;
	wire[2:0] w_n164_0;
	wire[2:0] w_n164_1;
	wire[2:0] w_n164_2;
	wire[1:0] w_n164_3;
	wire[1:0] w_n167_0;
	wire[1:0] w_n168_0;
	wire[2:0] w_n170_0;
	wire[1:0] w_n170_1;
	wire[1:0] w_n173_0;
	wire[2:0] w_n178_0;
	wire[2:0] w_n178_1;
	wire[2:0] w_n178_2;
	wire[1:0] w_n178_3;
	wire[2:0] w_n181_0;
	wire[1:0] w_n185_0;
	wire[2:0] w_n197_0;
	wire[2:0] w_n198_0;
	wire[1:0] w_n200_0;
	wire[1:0] w_n209_0;
	wire[2:0] w_n218_0;
	wire[1:0] w_n218_1;
	wire[2:0] w_n219_0;
	wire[2:0] w_n222_0;
	wire[2:0] w_n233_0;
	wire[1:0] w_n233_1;
	wire[1:0] w_n234_0;
	wire[1:0] w_n235_0;
	wire[2:0] w_n239_0;
	wire[1:0] w_n239_1;
	wire[1:0] w_n240_0;
	wire[1:0] w_n241_0;
	wire[1:0] w_n242_0;
	wire[1:0] w_n245_0;
	wire[1:0] w_n247_0;
	wire[1:0] w_n249_0;
	wire[1:0] w_n258_0;
	wire[1:0] w_n260_0;
	wire[1:0] w_n262_0;
	wire[2:0] w_n267_0;
	wire[2:0] w_n285_0;
	wire[2:0] w_n303_0;
	wire[1:0] w_n303_1;
	wire[2:0] w_n306_0;
	wire[1:0] w_n306_1;
	wire[2:0] w_n311_0;
	wire[2:0] w_n311_1;
	wire[2:0] w_n319_0;
	wire[2:0] w_n319_1;
	wire[1:0] w_n320_0;
	wire[1:0] w_n321_0;
	wire[2:0] w_n327_0;
	wire[2:0] w_n327_1;
	wire[1:0] w_n328_0;
	wire[1:0] w_n329_0;
	wire[2:0] w_n335_0;
	wire[1:0] w_n335_1;
	wire[2:0] w_n336_0;
	wire[1:0] w_n339_0;
	wire[1:0] w_n343_0;
	wire[1:0] w_n346_0;
	wire[1:0] w_n348_0;
	wire[1:0] w_n350_0;
	wire[1:0] w_n352_0;
	wire[1:0] w_n355_0;
	wire[1:0] w_n361_0;
	wire[2:0] w_n377_0;
	wire[1:0] w_n391_0;
	wire[1:0] w_n393_0;
	wire[2:0] w_n404_0;
	wire[2:0] w_n420_0;
	wire w_dff_B_1CEGbPvb3_2;
	wire w_dff_B_31NqMquM7_1;
	wire w_dff_B_898klcWp2_1;
	wire w_dff_A_RoEms7Ki0_1;
	wire w_dff_A_93NRgkcP8_1;
	wire w_dff_B_ebNhaN5W2_1;
	wire w_dff_B_CPF8Woo24_1;
	wire w_dff_B_cLth2hkf3_1;
	wire w_dff_B_yptoowMS6_1;
	wire w_dff_B_LPpNpuYv6_1;
	wire w_dff_B_UEMNSjmT2_1;
	wire w_dff_B_whXXqEr29_1;
	wire w_dff_B_IW5aM6qg5_1;
	wire w_dff_B_fVDOO5gV5_0;
	wire w_dff_B_mmcesAxq8_0;
	wire w_dff_B_5hwMQP213_0;
	wire w_dff_B_GcyP0NqW6_0;
	wire w_dff_B_gEBb9dRg0_0;
	wire w_dff_B_i783zhWw9_0;
	wire w_dff_B_VhHJXHd58_0;
	wire w_dff_B_VwoFMJOR7_0;
	wire w_dff_B_YOAELoHn9_0;
	wire w_dff_B_Hs1qRRcX5_0;
	wire w_dff_B_OkIX0lT05_0;
	wire w_dff_B_L3FYPAHp2_0;
	wire w_dff_B_SjQqSxhC5_0;
	wire w_dff_B_U2Ez93Tr9_0;
	wire w_dff_B_DzqD2APM0_1;
	wire w_dff_B_ME7H3JVk1_1;
	wire w_dff_B_iNXNHolu3_1;
	wire w_dff_B_gAxZpEKN6_1;
	wire w_dff_B_xlWS6p896_1;
	wire w_dff_B_vCCuB4CT6_1;
	wire w_dff_B_QpUcM2BV6_1;
	wire w_dff_B_bKe4wP4T8_1;
	wire w_dff_B_UnLTmpaN7_1;
	wire w_dff_B_NI0cE1AZ1_1;
	wire w_dff_B_GnGBpPiK7_1;
	wire w_dff_B_8EEViAgp5_1;
	wire w_dff_B_ZBXRjinY4_1;
	wire w_dff_B_vpM9D0Nn1_1;
	wire w_dff_B_7gp16oMc7_1;
	wire w_dff_B_Rj3ZIoqq0_1;
	wire w_dff_B_CttyHu5X5_1;
	wire w_dff_B_eqnvoQfK6_1;
	wire w_dff_B_1zCmO3lA2_1;
	wire w_dff_B_mGP2rv5o3_1;
	wire w_dff_B_FL9O8gPR8_1;
	wire w_dff_B_df95UIfR2_0;
	wire w_dff_B_XuzvRLPn3_0;
	wire w_dff_B_stLYjEdZ3_0;
	wire w_dff_B_3zVDPLk09_0;
	wire w_dff_B_QzWvvx3q0_0;
	wire w_dff_B_4lmlfvqX7_0;
	wire w_dff_B_UUZuZzHr4_0;
	wire w_dff_B_cmR8wiw80_0;
	wire w_dff_A_11az7EPc0_1;
	wire w_dff_A_J0on60g63_1;
	wire w_dff_A_4XAIkLJo8_1;
	wire w_dff_A_xTzFV7qt0_1;
	wire w_dff_A_uGzJbVJk5_1;
	wire w_dff_A_rx4gjPAv9_1;
	wire w_dff_A_aAbtjdr84_1;
	wire w_dff_A_ttwvEnVp9_1;
	wire w_dff_A_WgetRk2g0_1;
	wire w_dff_A_y8Eld7Ju7_1;
	wire w_dff_B_XY0MeAbk0_1;
	wire w_dff_B_c9O0j8eg6_1;
	wire w_dff_B_NwbbVXk69_1;
	wire w_dff_B_H0Cw9gyn7_1;
	wire w_dff_B_wJjuf0yv8_1;
	wire w_dff_B_pzxGdjD11_1;
	wire w_dff_B_mOBbxzxg0_0;
	wire w_dff_B_05R5fqsH1_0;
	wire w_dff_B_1IxAMKWI8_0;
	wire w_dff_B_OdaqrOtz5_0;
	wire w_dff_A_RUXZGA5t8_0;
	wire w_dff_A_8ptVZXIC5_0;
	wire w_dff_A_gaBE8EBh3_0;
	wire w_dff_A_0EQwirwp1_1;
	wire w_dff_A_tfA2nGQm0_1;
	wire w_dff_A_2p3IiiEe1_1;
	wire w_dff_A_6phzMpUm2_1;
	wire w_dff_A_Vs6wtd3O9_1;
	wire w_dff_B_7Jcnxepb2_1;
	wire w_dff_B_wMUZqVJX6_0;
	wire w_dff_B_6yVM5fKy6_0;
	wire w_dff_B_IhgK8L7H9_0;
	wire w_dff_B_gyWb3mQN5_0;
	wire w_dff_B_qKue6jvL7_1;
	wire w_dff_B_JyDi3Oy99_1;
	wire w_dff_B_MpRywvLK8_1;
	wire w_dff_B_WsMdoAZy9_1;
	wire w_dff_B_RATKL9N39_1;
	wire w_dff_B_kw6UwvrJ0_1;
	wire w_dff_B_ETZZTpSk0_1;
	wire w_dff_B_ogepBvZs6_1;
	wire w_dff_B_HrlsXUcx3_0;
	wire w_dff_B_cuXdf9w35_0;
	wire w_dff_B_n54Jdcop5_0;
	wire w_dff_B_ykWxcPfT8_0;
	wire w_dff_B_0I3M9pmG9_0;
	wire w_dff_B_LiJqcHEa1_0;
	wire w_dff_A_m5dLRo3E2_1;
	wire w_dff_A_Z6oCp6y41_1;
	wire w_dff_A_22A5OXr00_1;
	wire w_dff_A_Rxc8T17A4_1;
	wire w_dff_A_5b2xuoH16_1;
	wire w_dff_B_uKBg6Jm14_1;
	wire w_dff_B_2C1W7kJe2_1;
	wire w_dff_B_uX9nyNKO7_1;
	wire w_dff_B_FAex2s4q4_1;
	wire w_dff_B_XxtknBJ05_0;
	wire w_dff_B_ENeW9ryo0_0;
	wire w_dff_B_kP6EvrmH0_1;
	wire w_dff_B_8LqnAwx22_0;
	wire w_dff_B_GA6yjg4Y7_0;
	wire w_dff_B_zNGHe30A7_0;
	wire w_dff_B_ebZatS749_0;
	wire w_dff_B_ol4EIhmR1_1;
	wire w_dff_B_9kS0Tl0Z8_1;
	wire w_dff_B_V2uSvaJJ9_1;
	wire w_dff_B_JNic7gWJ7_1;
	wire w_dff_B_unMdeZK19_1;
	wire w_dff_B_M3nn9zj39_1;
	wire w_dff_B_ZKiGkW802_1;
	wire w_dff_B_AjMpcyz35_1;
	wire w_dff_B_khiGMJkC6_0;
	wire w_dff_B_cTdvZy4r8_0;
	wire w_dff_B_WCKlEtiR0_0;
	wire w_dff_B_2a5z1Xjg8_0;
	wire w_dff_B_n8OiMxVB2_0;
	wire w_dff_B_mC5ZY7pu3_0;
	wire w_dff_A_EG9VRG8W6_1;
	wire w_dff_A_TDoDTVbA9_1;
	wire w_dff_A_pkqm1NpZ6_1;
	wire w_dff_B_fQmRPZON8_1;
	wire w_dff_B_T2BT045J4_1;
	wire w_dff_B_Vjnz68aJ2_1;
	wire w_dff_B_HHKzXRgK4_1;
	wire w_dff_B_PKTNXSdz9_1;
	wire w_dff_B_1fe2UGLo9_1;
	wire w_dff_B_uFzmVCRF6_1;
	wire w_dff_B_oqSPIjM86_1;
	wire w_dff_B_aGB5ctIR2_1;
	wire w_dff_B_zCKZstdA2_1;
	wire w_dff_B_EPFRqy7F8_1;
	wire w_dff_B_4i9kXI6q3_1;
	wire w_dff_B_SAkTrJKB8_1;
	wire w_dff_B_9yKBK2lv1_1;
	wire w_dff_B_jQQigADs9_1;
	wire w_dff_B_1ghF9F5c0_1;
	wire w_dff_B_fgtMIk5n0_1;
	wire w_dff_B_4xuD6Oz99_1;
	wire w_dff_B_Sl7Zzit09_1;
	wire w_dff_B_knfWUuIT3_1;
	wire w_dff_B_JYzYanh11_1;
	wire w_dff_B_jn2LKAOE3_1;
	wire w_dff_B_Il4C0t5C1_1;
	wire w_dff_B_6ZBnnazU6_1;
	wire w_dff_B_6zpwPUYv8_1;
	wire w_dff_B_0sXp9gMc4_1;
	wire w_dff_B_FAoYoW3d1_1;
	wire w_dff_B_b5qaLfel0_1;
	wire w_dff_B_uRMRSEKs8_1;
	wire w_dff_B_BqlEClB84_1;
	wire w_dff_B_1Tv7GAvm9_1;
	wire w_dff_B_ve0nPmlW8_0;
	wire w_dff_B_tgWSbjKB2_0;
	wire w_dff_B_Jq33RNee0_0;
	wire w_dff_B_uERczs310_0;
	wire w_dff_B_9mc8XRc13_0;
	wire w_dff_B_8VlGQYTN5_0;
	wire w_dff_B_1qVZahQd5_0;
	wire w_dff_B_cT7p5vUi3_0;
	wire w_dff_B_kLpPMk8B5_0;
	wire w_dff_B_AENKSLvw6_0;
	wire w_dff_B_9BGn4cHj0_0;
	wire w_dff_B_oN1vl44e4_0;
	wire w_dff_B_Bs7DS11W5_0;
	wire w_dff_A_Cu0EyjeM0_0;
	wire w_dff_A_BJqwCyrt5_0;
	wire w_dff_A_lfm1JmaT8_0;
	wire w_dff_A_k31Yre1t9_0;
	wire w_dff_A_EBaxjGJw3_0;
	wire w_dff_A_UFCUDzQm4_0;
	wire w_dff_A_fz5qyEiG5_0;
	wire w_dff_A_eG6iFr2p8_0;
	wire w_dff_A_cwaJ42z55_0;
	wire w_dff_A_qHxwdpt16_0;
	wire w_dff_B_zqoxhkzJ3_1;
	wire w_dff_B_yG6Jm40g3_1;
	wire w_dff_B_jJJgY1Qs3_1;
	wire w_dff_B_95RgYvRz4_1;
	wire w_dff_B_aHtzEbHB4_1;
	wire w_dff_B_PFNWSu7G1_1;
	wire w_dff_B_Yykectua0_1;
	wire w_dff_B_BLIkJKXs8_1;
	wire w_dff_A_UPjMzRRM7_0;
	wire w_dff_A_stdpmX2N9_0;
	wire w_dff_A_iPzLhe5Q3_0;
	wire w_dff_A_xM7THKaw2_0;
	wire w_dff_A_7eFcm9HF7_0;
	wire w_dff_A_of1xeFnv0_1;
	wire w_dff_A_2zxuqYs59_1;
	wire w_dff_A_ywjDpfpj5_1;
	wire w_dff_A_jnnl83Gv3_1;
	wire w_dff_A_YnXncBJ56_1;
	wire w_dff_A_2GrLUlwC4_0;
	wire w_dff_A_Fmz9ih9H1_0;
	wire w_dff_A_B01JyBuR4_0;
	wire w_dff_A_Yb8ZA5p08_0;
	wire w_dff_A_pxZ0xUpf1_0;
	wire w_dff_A_C7Mu9xf33_0;
	wire w_dff_A_OKZjSb8D3_0;
	wire w_dff_A_cbvdV27n2_0;
	wire w_dff_A_0Dvpp9520_0;
	wire w_dff_A_fs0rZYQO3_0;
	wire w_dff_B_BRCBa8Gm3_1;
	wire w_dff_B_dE3nxvlr2_1;
	wire w_dff_B_JhWLMC056_1;
	wire w_dff_B_JWUBqizD4_1;
	wire w_dff_B_hXbeFuTr8_1;
	wire w_dff_B_w0avvtP58_1;
	wire w_dff_B_lAvnDYCV9_1;
	wire w_dff_B_CCaDncC33_1;
	wire w_dff_B_nRcRGbWL5_1;
	wire w_dff_B_kSHNl5BN0_1;
	wire w_dff_B_udxFi3po4_1;
	wire w_dff_B_cgovtZgz8_1;
	wire w_dff_B_cwtaCgur6_1;
	wire w_dff_B_j1jZDTRW8_1;
	wire w_dff_B_tl4V774Y2_0;
	wire w_dff_B_9qAjwCpN3_0;
	wire w_dff_B_GgSowWm09_0;
	wire w_dff_B_u4XwBN3V3_0;
	wire w_dff_B_Qqh7uzFs6_0;
	wire w_dff_B_mbSjwtzG9_0;
	wire w_dff_B_Wei9aZmN0_0;
	wire w_dff_B_QgysHtIL2_0;
	wire w_dff_B_Zd8bgh8O6_0;
	wire w_dff_B_mHafxW2Q4_0;
	wire w_dff_B_CX3IjYz83_0;
	wire w_dff_B_iVt3tfbj1_0;
	wire w_dff_B_p8dNjgNM2_0;
	wire w_dff_B_DJB3hdRk1_1;
	wire w_dff_B_FJqerLoq1_1;
	wire w_dff_B_Wq865ogK6_1;
	wire w_dff_B_LewQBoAp5_1;
	wire w_dff_B_NeTiRv242_1;
	wire w_dff_B_spsy8lYm5_1;
	wire w_dff_B_pPASdmkn0_1;
	wire w_dff_B_Q5hMidMZ8_1;
	wire w_dff_B_6l3PGBbg8_1;
	wire w_dff_B_ntz2DTLr8_1;
	wire w_dff_B_gyQzON464_1;
	wire w_dff_B_uC21U4j09_1;
	wire w_dff_B_1zGjvSz99_1;
	wire w_dff_B_Odu7rsgL8_1;
	wire w_dff_B_CeDgb4uI5_1;
	wire w_dff_B_hLhf6NjV9_1;
	wire w_dff_B_0gP8RICC7_1;
	wire w_dff_B_CDBMehEJ7_1;
	wire w_dff_B_K4ubMvt41_1;
	wire w_dff_B_pVGD8yq74_1;
	wire w_dff_B_6mcDbINK2_1;
	wire w_dff_B_4BmzX0fv0_1;
	wire w_dff_B_kXtpPMaG3_1;
	wire w_dff_A_6XpegKSm4_1;
	wire w_dff_A_drOnVS6z3_1;
	wire w_dff_A_LrXIiMcv6_1;
	wire w_dff_A_yAmbt8ID9_1;
	wire w_dff_A_0jQ6sryO3_1;
	wire w_dff_A_o0i22IS56_1;
	wire w_dff_A_jv5mWzwL6_1;
	wire w_dff_A_ihPpej2Q0_1;
	wire w_dff_A_7JtItBnh3_1;
	wire w_dff_A_Zm3lozEW9_1;
	wire w_dff_A_3nGvN2zy2_1;
	wire w_dff_A_BdvaWRgm5_1;
	wire w_dff_A_drq8MwUV8_1;
	wire w_dff_A_oVQe4ZXh9_1;
	wire w_dff_A_zTsKiS1O7_1;
	wire w_dff_A_2m1P00Ww4_1;
	wire w_dff_A_nDwfb40U1_1;
	wire w_dff_A_bXrPZwFe6_1;
	wire w_dff_A_MgiaceAj4_1;
	wire w_dff_A_WYotL46y6_1;
	wire w_dff_A_d2Hob7nh7_1;
	wire w_dff_A_4ss6uSeZ6_1;
	wire w_dff_A_HHwTvurL0_1;
	wire w_dff_A_VinsUufh7_1;
	wire w_dff_A_QPcncT2h7_1;
	wire w_dff_B_9u6nPr194_1;
	wire w_dff_B_8D4hzEhG8_0;
	wire w_dff_B_rEqfqAFS6_0;
	wire w_dff_B_BPh8WUSn4_0;
	wire w_dff_B_H1YqvDCf7_0;
	wire w_dff_B_EUSsslwO7_0;
	wire w_dff_B_0Al4fIGv0_0;
	wire w_dff_B_aw9470NU3_0;
	wire w_dff_B_gZLslMqB6_0;
	wire w_dff_B_Jz4QAnE20_0;
	wire w_dff_B_CSH8IHe66_0;
	wire w_dff_B_IEinr5W55_0;
	wire w_dff_B_oBmZdDdv8_0;
	wire w_dff_A_VE65fi8p4_1;
	wire w_dff_A_8npv2VtM7_1;
	wire w_dff_A_NN5MZ7WJ6_1;
	wire w_dff_A_tVDnmAWv5_1;
	wire w_dff_A_I1W6iqkX5_1;
	wire w_dff_A_GXwDeevO2_1;
	wire w_dff_A_1kAzhMjp9_1;
	wire w_dff_A_hwuFFAAX3_1;
	wire w_dff_A_MOddnX0B8_1;
	wire w_dff_A_FfDxJoP55_1;
	wire w_dff_A_U6VAVltF6_1;
	wire w_dff_A_wKyYd6S56_1;
	wire w_dff_A_nZJIOFmZ7_1;
	wire w_dff_A_Wm4FoYEo2_1;
	wire w_dff_B_b71Job3Z5_1;
	wire w_dff_B_Sf1zdOW27_0;
	wire w_dff_B_LeYyGgHc9_0;
	wire w_dff_B_WWxggge34_0;
	wire w_dff_B_8nT4UyrV7_0;
	wire w_dff_B_eN03l9Bm9_0;
	wire w_dff_B_3ValmUWV0_0;
	wire w_dff_B_ZolByrk60_1;
	wire w_dff_B_wsv61f505_1;
	wire w_dff_B_J9Wx4gGl4_1;
	wire w_dff_B_G73jK7Yv0_1;
	wire w_dff_B_YZqZ1I5a4_1;
	wire w_dff_B_6zkGhcqR0_1;
	wire w_dff_B_iL7YsaSi3_1;
	wire w_dff_B_mmGwhevC0_1;
	wire w_dff_B_y9yv7Atf3_1;
	wire w_dff_B_otcIjMka3_1;
	wire w_dff_B_Y9GjR7lO0_1;
	wire w_dff_B_GbNwPoWg2_1;
	wire w_dff_B_kHNch1gY8_1;
	wire w_dff_B_RpbT6EdF9_0;
	wire w_dff_B_DX3c679I1_0;
	wire w_dff_B_MikbEnIR6_0;
	wire w_dff_B_WWSsA49G4_0;
	wire w_dff_B_MkiFlSdV1_0;
	wire w_dff_B_y4HYu6Jw1_0;
	wire w_dff_B_xlS5GCmq0_0;
	wire w_dff_B_J6Sg49TN7_0;
	wire w_dff_B_ckyUDNnz6_0;
	wire w_dff_B_aPkeSVf45_0;
	wire w_dff_B_U4V7GEKf5_0;
	wire w_dff_B_NiSVb9Os5_1;
	wire w_dff_B_V5DqC9ZO5_1;
	wire w_dff_B_NQHEajNl6_1;
	wire w_dff_B_fwR8nQXi6_1;
	wire w_dff_B_Z8eQGXLn4_1;
	wire w_dff_B_no5Sn7fN3_1;
	wire w_dff_B_zKyFHKTi2_1;
	wire w_dff_B_dt9sWZbE6_1;
	wire w_dff_B_Ma9DwKAm4_1;
	wire w_dff_B_FXd0XQD89_1;
	wire w_dff_B_c5FYvj8b9_1;
	wire w_dff_B_bPMLuo3p9_1;
	wire w_dff_B_el4TNwmN7_1;
	wire w_dff_B_ZGdEnHiH1_1;
	wire w_dff_B_bpbVVJxx7_1;
	wire w_dff_B_iQ7bSX4n0_1;
	wire w_dff_B_Qiyg8Xpl5_1;
	wire w_dff_B_V5OrcNKd5_1;
	wire w_dff_B_HjtU3Aed2_1;
	wire w_dff_A_nC3SVYna5_1;
	wire w_dff_A_2nvY5ech3_1;
	wire w_dff_A_vYh9QrKF0_1;
	wire w_dff_A_7EYB9jgz2_1;
	wire w_dff_A_rEl56Bl92_1;
	wire w_dff_A_F4wyE4ca0_1;
	wire w_dff_A_nDCqtvNd2_1;
	wire w_dff_A_0xAL95QH9_1;
	wire w_dff_A_XP5ba5uf3_1;
	wire w_dff_A_cY3IRWIR9_1;
	wire w_dff_A_byFM5CMs1_1;
	wire w_dff_A_lWkHPceK0_1;
	wire w_dff_A_uLw6UAGe3_1;
	wire w_dff_A_rJHttrSe5_1;
	wire w_dff_A_kPEQXXh86_1;
	wire w_dff_A_udFDzaU99_1;
	wire w_dff_A_ANfIQFMG9_1;
	wire w_dff_A_9mkipwhk5_1;
	wire w_dff_A_dqMb4v3t7_1;
	wire w_dff_A_YCTG0Q1d0_1;
	wire w_dff_A_C0tNwMXZ7_1;
	wire w_dff_B_KYrhI0hC1_1;
	wire w_dff_B_ACO85Wrf1_0;
	wire w_dff_B_k7CZ7hhD3_0;
	wire w_dff_B_qQoAygvn1_0;
	wire w_dff_B_yqPklDZu7_0;
	wire w_dff_B_f31QfJbB3_0;
	wire w_dff_B_w6CpIRLc4_0;
	wire w_dff_B_rV088fa16_0;
	wire w_dff_B_mwsxLrJF3_0;
	wire w_dff_B_cjMy5KA00_0;
	wire w_dff_B_cs5Ker5C6_0;
	wire w_dff_B_vuJxep6s2_0;
	wire w_dff_B_W5jbDRS45_0;
	wire w_dff_A_IwDjKkBE0_1;
	wire w_dff_A_3bZIFlVQ8_1;
	wire w_dff_A_FXkBUiM52_1;
	wire w_dff_A_F4txEN0w3_1;
	wire w_dff_A_dCTX42Ty0_1;
	wire w_dff_A_pg7rHJG33_1;
	wire w_dff_A_oL28DVCB8_1;
	wire w_dff_A_AfHaIRxi5_1;
	wire w_dff_A_flsEitT15_1;
	wire w_dff_A_LuxiEYsX8_1;
	wire w_dff_A_gX7i0XKC4_1;
	wire w_dff_A_xWZaWM6C1_1;
	wire w_dff_B_kmBlNeDa0_0;
	wire w_dff_B_bkn0FYDb9_0;
	wire w_dff_B_dJnYQKnp4_0;
	wire w_dff_B_lh2Yrq4M4_0;
	wire w_dff_B_Z9TYzfVw8_0;
	wire w_dff_A_3XFyiUAB4_0;
	wire w_dff_A_D50Szkfz6_0;
	wire w_dff_B_x2OqQQJj7_1;
	wire w_dff_B_xRtgmgyj1_1;
	wire w_dff_B_dcvMEqTw1_1;
	wire w_dff_B_HNAqs8C04_1;
	wire w_dff_B_s3mmBsKy9_1;
	wire w_dff_B_0SBp3vsu3_1;
	wire w_dff_B_vQPr47jz8_1;
	wire w_dff_B_18risy2H5_1;
	wire w_dff_B_kuM9YojE4_1;
	wire w_dff_B_mqO1nELF3_1;
	wire w_dff_B_4PayGcsh8_1;
	wire w_dff_B_MHy3BuVX4_1;
	wire w_dff_B_x5888I8n6_1;
	wire w_dff_B_Gbl7UWRP9_1;
	wire w_dff_B_74pt3QHk6_1;
	wire w_dff_B_tybF7BoW7_1;
	wire w_dff_B_J5ysfJUO0_1;
	wire w_dff_B_Fu1JlMXh1_1;
	wire w_dff_B_xWFVi4sX9_1;
	wire w_dff_B_fzwK6v1P7_1;
	wire w_dff_B_cvIQccYk8_1;
	wire w_dff_B_Ymb89kTl0_0;
	wire w_dff_A_6pwiBZiD1_1;
	wire w_dff_A_RWZmEWs59_1;
	wire w_dff_A_JONvI4Ah7_2;
	wire w_dff_A_GyAh0DSE4_2;
	wire w_dff_A_SI1dviB09_2;
	wire w_dff_A_IYzUJds28_2;
	wire w_dff_A_EMlu2N5b4_0;
	wire w_dff_A_Ti5cg5ph1_0;
	wire w_dff_A_PGDTSPWh0_0;
	wire w_dff_A_hdvXsXBp9_0;
	wire w_dff_A_MoIeqth39_0;
	wire w_dff_A_JtfTxExS7_0;
	wire w_dff_A_QzQoHkma3_0;
	wire w_dff_A_Ib2ld3B62_0;
	wire w_dff_A_k8q9eGSe7_0;
	wire w_dff_A_2HLhW8dn4_1;
	wire w_dff_B_nealyHUp2_3;
	wire w_dff_B_xtI4oHHV2_3;
	wire w_dff_B_bayc14bM7_3;
	wire w_dff_B_0i1sCJu34_3;
	wire w_dff_B_byz4GMMS8_3;
	wire w_dff_B_6th8OTEB6_3;
	wire w_dff_B_YsyELdkb6_3;
	wire w_dff_B_ADMuWfEC4_3;
	wire w_dff_B_CBt1BKL09_3;
	wire w_dff_B_ZbozWSWy9_3;
	wire w_dff_B_GMdIAMAk0_3;
	wire w_dff_B_HuHRgb4z3_3;
	wire w_dff_B_yd3rmF5e8_0;
	wire w_dff_B_tVoOs6xB3_0;
	wire w_dff_B_HnNJIOhJ6_0;
	wire w_dff_B_2B2v49to7_0;
	wire w_dff_B_rwgBmrGf7_0;
	wire w_dff_B_YwmusE7S0_0;
	wire w_dff_B_92mOriVu0_0;
	wire w_dff_B_cUIJ56Cx7_0;
	wire w_dff_B_eCn0yA8Z3_0;
	wire w_dff_B_sDhUd0Mh1_1;
	wire w_dff_B_hXqSAjS32_1;
	wire w_dff_B_PotbSWsY0_1;
	wire w_dff_B_lcAPsD593_1;
	wire w_dff_B_ffLRV7A62_1;
	wire w_dff_B_TsYMy0rj5_1;
	wire w_dff_B_7RhKTItA8_1;
	wire w_dff_B_BnHVhi8v1_1;
	wire w_dff_B_J3NRScyI2_1;
	wire w_dff_B_VDeR1XEv4_1;
	wire w_dff_B_VzH4R8Tb0_1;
	wire w_dff_B_HA636BSQ9_1;
	wire w_dff_B_oSafIrro8_1;
	wire w_dff_B_vIeKzdDZ5_1;
	wire w_dff_B_D2Y4UE0M3_1;
	wire w_dff_B_MMyIBFcg6_1;
	wire w_dff_B_fX5KxfZH6_1;
	wire w_dff_B_DPoa9dGu1_1;
	wire w_dff_B_oueMcbXP4_1;
	wire w_dff_B_iqUzzj4d5_1;
	wire w_dff_B_BWLpF0KT9_1;
	wire w_dff_B_dO6qtV3b4_1;
	wire w_dff_B_IEyFdywL9_1;
	wire w_dff_B_bjbKh9n43_1;
	wire w_dff_B_Y1UyWR7U8_1;
	wire w_dff_B_JwNGO53n3_1;
	wire w_dff_B_zVRLC9Ba5_1;
	wire w_dff_B_COuJfQxM1_1;
	wire w_dff_B_1yNXocHa2_1;
	wire w_dff_A_4cNoCPSg0_1;
	wire w_dff_B_uq5YB8iY8_2;
	wire w_dff_B_FB1pJWiG3_2;
	wire w_dff_B_zU9dKjYx9_2;
	wire w_dff_B_sqAbqZFa9_2;
	wire w_dff_B_aAin9rsL6_2;
	wire w_dff_B_U1QogUBc1_2;
	wire w_dff_B_J4gD7p7d8_2;
	wire w_dff_B_V3pVTEM05_2;
	wire w_dff_B_LL0ht2Ne4_2;
	wire w_dff_A_E5k1HrQO9_0;
	wire w_dff_B_VKIL1KgJ4_1;
	wire w_dff_B_uB5UaBTU2_3;
	wire w_dff_B_8JH9X9W86_3;
	wire w_dff_B_wCN4TqMH2_3;
	wire w_dff_B_9q4cAsx81_3;
	wire w_dff_B_mF65vmDV9_3;
	wire w_dff_B_V1UkLjfl8_3;
	wire w_dff_B_eKqibSVd7_3;
	wire w_dff_B_BEqYUOMv2_3;
	wire w_dff_A_CEQ0lxKp2_1;
	wire w_dff_A_qT6muqyn8_1;
	wire w_dff_A_ZuR8lNHC0_1;
	wire w_dff_A_C7z8XBoT4_1;
	wire w_dff_A_XJnaNOnP7_1;
	wire w_dff_A_w6ASu1417_1;
	wire w_dff_A_Zzzc8CrR8_1;
	wire w_dff_A_3nkQ5RB82_1;
	wire w_dff_A_dn19Lk7u3_1;
	wire w_dff_A_f8gnE0gU2_1;
	wire w_dff_A_JARPD4A55_1;
	wire w_dff_A_0VkJRlpF6_1;
	wire w_dff_A_XZk3ieHp2_1;
	wire w_dff_A_yN8XxgSW7_1;
	wire w_dff_A_i4ftW9cE8_1;
	wire w_dff_A_IrI6sxS90_1;
	wire w_dff_A_yanv0OM79_1;
	wire w_dff_A_npFGjXrQ4_1;
	wire w_dff_A_ktiDR8at9_1;
	wire w_dff_B_TpqTVJ4n0_2;
	wire w_dff_B_iJFi5h6D0_2;
	wire w_dff_B_vKcqEVzi0_2;
	wire w_dff_B_oEo3lIF12_2;
	wire w_dff_A_812H5gga4_0;
	wire w_dff_A_29hTzBdz1_0;
	wire w_dff_A_RHCq5V7U5_0;
	wire w_dff_A_GibsDc8A7_0;
	wire w_dff_A_THLsNrii0_0;
	wire w_dff_A_xLgms4vS7_0;
	wire w_dff_B_3De2OvN21_1;
	wire w_dff_B_9s0KUMA57_1;
	wire w_dff_B_5r88tqMS6_1;
	wire w_dff_B_pPLs2kKB7_1;
	wire w_dff_B_rEQ14hc79_1;
	wire w_dff_B_YPFORqkM5_1;
	wire w_dff_B_km6G1oom0_1;
	wire w_dff_B_jf0EZXZZ0_1;
	wire w_dff_A_qMP30cKL8_1;
	wire w_dff_A_ctMDOhS61_1;
	wire w_dff_A_KPw1I5xz5_1;
	wire w_dff_A_CjNlyoDA3_1;
	wire w_dff_A_OB9FY0mw8_1;
	wire w_dff_A_zCvbnzqH0_1;
	wire w_dff_A_ilpXpt4I6_1;
	wire w_dff_A_FEssNtyE2_1;
	wire w_dff_A_z7MgNYZq9_1;
	wire w_dff_B_RuFuQY6l2_2;
	wire w_dff_B_c9eL9yPE2_2;
	wire w_dff_B_9C246Ov72_2;
	wire w_dff_B_XhZnIYUG3_2;
	wire w_dff_A_4jVZ6Q4k0_2;
	wire w_dff_A_eyc1lp049_2;
	wire w_dff_A_vRECN8X80_0;
	wire w_dff_A_BXbPzA7g5_0;
	wire w_dff_A_mqntJa0Q9_0;
	wire w_dff_A_uAXpYeU64_0;
	wire w_dff_A_fHltFPqQ2_0;
	wire w_dff_A_A7xyoMr72_0;
	wire w_dff_A_k9lRbkI00_0;
	wire w_dff_B_lBgFsyx20_1;
	wire w_dff_B_UWSlXJpb0_1;
	wire w_dff_B_VMwBgffC5_1;
	wire w_dff_B_M1Co64tr0_1;
	wire w_dff_B_ARK7wgVa3_1;
	wire w_dff_B_B1TVZA8A8_1;
	wire w_dff_B_RLjpRnwm5_1;
	wire w_dff_B_packt20l1_1;
	wire w_dff_B_kH9XimPh4_1;
	wire w_dff_A_4KfbYxTX8_2;
	wire w_dff_A_a3hEkdSU9_2;
	wire w_dff_A_g8OKYjpm7_2;
	wire w_dff_A_dNObNzfW5_2;
	wire w_dff_A_C9AsslSj3_2;
	wire w_dff_A_TqEfXRn22_2;
	wire w_dff_A_pYcbskS19_2;
	wire w_dff_A_1VsQDjyT1_2;
	wire w_dff_A_I9q8PbWb9_2;
	wire w_dff_B_Adq0vX6W4_0;
	wire w_dff_B_njyr8vIk2_0;
	wire w_dff_B_Lpn9Z3KK6_0;
	wire w_dff_B_JG5eNFVF2_0;
	wire w_dff_B_3mYVtRII6_0;
	wire w_dff_B_2kQkNnHJ0_1;
	wire w_dff_B_phD424OH4_0;
	wire w_dff_B_DSR0Iwlk1_0;
	wire w_dff_B_vW0l3lgO9_0;
	wire w_dff_B_AVjAxP8g4_0;
	wire w_dff_B_O7Q7vZ1q1_0;
	wire w_dff_B_Hz9FnoPw5_0;
	wire w_dff_B_T7xEy7BW6_0;
	wire w_dff_B_WFxQdlRu6_0;
	wire w_dff_B_7YlY6QFn3_0;
	wire w_dff_B_nK1sqyT44_0;
	wire w_dff_B_oS9HL1Vp2_0;
	wire w_dff_B_fWNdO3uh7_0;
	wire w_dff_A_3vB0jX6m8_0;
	wire w_dff_A_ZkgXwSBz1_0;
	wire w_dff_A_PumeAMUn9_0;
	wire w_dff_A_AMi2o2DU1_0;
	wire w_dff_A_W951Bk605_0;
	wire w_dff_A_ROlnZwSd1_0;
	wire w_dff_A_ayTVddLw1_0;
	wire w_dff_A_26g6vfx57_0;
	wire w_dff_A_NULuFxEu5_0;
	wire w_dff_A_mAAVI44v4_0;
	wire w_dff_A_gDQHMYla4_0;
	wire w_dff_B_e8Cptkpo8_3;
	wire w_dff_B_Y6SQOTPq6_3;
	wire w_dff_B_mUnJNkGj4_3;
	wire w_dff_B_UmB4pous4_3;
	wire w_dff_B_fv5ELtF35_3;
	wire w_dff_B_fvAHvOyo3_3;
	wire w_dff_B_ysQSu4lh2_3;
	wire w_dff_B_bgjsFjNt8_3;
	wire w_dff_B_ZIZCD5EV5_3;
	wire w_dff_B_XMZ4bwEE7_0;
	wire w_dff_B_M9ufdmyz8_0;
	wire w_dff_B_b9KVB5Ps8_0;
	wire w_dff_B_Z2RNZhHl2_0;
	wire w_dff_B_D33PHtD84_0;
	wire w_dff_A_GMKVTrYB1_1;
	wire w_dff_B_eapsGmJZ7_2;
	wire w_dff_B_CRYdfOjP6_2;
	wire w_dff_B_mDG0AUJA2_2;
	wire w_dff_B_dNetj7Sz0_2;
	wire w_dff_B_X2HSRZXt6_1;
	wire w_dff_A_o84xzYsp9_1;
	wire w_dff_A_W9ACGTnI8_1;
	wire w_dff_A_GZc8ihL28_2;
	wire w_dff_A_2cGXA9CZ0_2;
	wire w_dff_A_ClR1RSNQ7_2;
	wire w_dff_A_tbx6V7qa2_0;
	wire w_dff_A_hCZC8D6S0_0;
	wire w_dff_B_AvgRFnk69_2;
	wire w_dff_B_cbwv2hc83_2;
	wire w_dff_B_XH2BfRRp4_2;
	wire w_dff_B_hBYn5AJP7_2;
	wire w_dff_A_c5h1KxxZ5_2;
	wire w_dff_A_0hz0x1rk4_0;
	wire w_dff_A_lzBRTOd43_0;
	wire w_dff_A_LuIFG4NY8_0;
	wire w_dff_A_OjtJI3LO3_0;
	wire w_dff_A_kNatINEV2_0;
	wire w_dff_A_ahb4I5EB5_0;
	wire w_dff_A_HKZnpPuc7_0;
	wire w_dff_A_gITBhv6J7_0;
	wire w_dff_A_squcgHag0_0;
	wire w_dff_A_Tfn9dkpY0_0;
	wire w_dff_A_hu1UzQuk0_0;
	wire w_dff_A_DDJjnWAb7_0;
	wire w_dff_A_wAENiHcK5_0;
	wire w_dff_A_BRk26rU56_0;
	wire w_dff_A_Kjt2lBi47_0;
	wire w_dff_A_I77dcwIH0_0;
	wire w_dff_A_lrcGNN8K0_0;
	wire w_dff_A_xqktSLiR8_0;
	wire w_dff_A_xyAdLGRP0_0;
	wire w_dff_A_mTfym79l9_0;
	wire w_dff_A_kKppd7Q86_0;
	wire w_dff_A_Coh57M5J7_0;
	wire w_dff_A_9kXdEFYu4_0;
	wire w_dff_A_ovCiETst6_0;
	wire w_dff_A_jlWpYqjF7_0;
	wire w_dff_A_YHZgzuPt7_2;
	wire w_dff_A_2pj7O4Oz1_0;
	wire w_dff_A_p5iXJXfI3_0;
	wire w_dff_A_kmHT3BLT7_0;
	wire w_dff_A_CBHOuStn6_0;
	wire w_dff_A_7jEBTaXk6_0;
	wire w_dff_A_fiGJKQ7K0_0;
	wire w_dff_A_t9yd53Aj8_0;
	wire w_dff_A_Z4cNUS6r7_0;
	wire w_dff_A_fJNDyBEI4_0;
	wire w_dff_A_jLWAwJhD5_0;
	wire w_dff_A_9GjkLUdN6_0;
	wire w_dff_A_RA0lXuQX4_0;
	wire w_dff_A_g9CnU2Mo3_0;
	wire w_dff_A_kTSVgl7x6_0;
	wire w_dff_A_aEuud5z42_0;
	wire w_dff_A_9wEAD8aZ8_0;
	wire w_dff_A_Kk07Xzig4_0;
	wire w_dff_A_j7h72xcg4_0;
	wire w_dff_A_s0ZNuBuv9_0;
	wire w_dff_A_8Ojp18G63_0;
	wire w_dff_A_VvWr8UZz5_0;
	wire w_dff_A_ycyIkFor0_0;
	wire w_dff_A_iPSVez904_0;
	wire w_dff_A_hjVCQoff5_0;
	wire w_dff_A_bXcbNNkp5_0;
	wire w_dff_A_7Fl3brhr8_2;
	wire w_dff_A_Vj7jclsq4_0;
	wire w_dff_A_PxxECmuW9_0;
	wire w_dff_A_QJMYOs5p5_0;
	wire w_dff_A_IFUgtrnu2_0;
	wire w_dff_A_NlNE6MGn6_0;
	wire w_dff_A_FRXKEXcd8_0;
	wire w_dff_A_H4UR5eXj1_0;
	wire w_dff_A_V18BWkYp0_0;
	wire w_dff_A_pln6gSJq9_0;
	wire w_dff_A_43AVfQz67_0;
	wire w_dff_A_h0mk5r0I2_0;
	wire w_dff_A_yylNi8HB5_0;
	wire w_dff_A_SMwMkbNL2_0;
	wire w_dff_A_5CimCWX73_0;
	wire w_dff_A_TVNGGGuQ7_0;
	wire w_dff_A_2YrnX8Nc4_0;
	wire w_dff_A_HSrhI1nk6_0;
	wire w_dff_A_yFiJAvbr8_0;
	wire w_dff_A_WzppOk8E1_0;
	wire w_dff_A_ZBK14rFI0_0;
	wire w_dff_A_T0ZiEYZJ3_0;
	wire w_dff_A_302dtReM9_0;
	wire w_dff_A_Zlz96OXR9_0;
	wire w_dff_A_6xOEEjyv3_0;
	wire w_dff_A_VsgpJBsG9_0;
	wire w_dff_A_5rAfykWU6_2;
	wire w_dff_A_CzzcoIrD4_0;
	wire w_dff_A_ex3mqZMD4_0;
	wire w_dff_A_NTp0Tono1_0;
	wire w_dff_A_hFM5zlto8_0;
	wire w_dff_A_onB6vq4B5_0;
	wire w_dff_A_p73G01dB3_0;
	wire w_dff_A_laiYJfCm3_0;
	wire w_dff_A_4uKSTSHW0_0;
	wire w_dff_A_CjUlM47D4_0;
	wire w_dff_A_oaxb6zZz4_0;
	wire w_dff_A_toC1T2xZ3_0;
	wire w_dff_A_vbgWhGs84_0;
	wire w_dff_A_FoUtZfni6_0;
	wire w_dff_A_2rpz6Gtd8_0;
	wire w_dff_A_ZLLxJkv58_0;
	wire w_dff_A_Yf09qgEI9_0;
	wire w_dff_A_LtbDNfuw2_0;
	wire w_dff_A_bPWhjKrN9_0;
	wire w_dff_A_UhhShjdn2_0;
	wire w_dff_A_YASDx3W27_0;
	wire w_dff_A_o26qZyEt8_0;
	wire w_dff_A_tPu3aBsV1_0;
	wire w_dff_A_njIE0DK75_0;
	wire w_dff_A_3H0m2vnj9_0;
	wire w_dff_A_EDknwrmB1_0;
	wire w_dff_A_U7VvD8Jc2_0;
	wire w_dff_A_9uEusv4s6_2;
	wire w_dff_A_TFLZaW9g7_0;
	wire w_dff_A_za17e4i92_0;
	wire w_dff_A_79NOVBLH2_0;
	wire w_dff_A_dnI1umAM1_0;
	wire w_dff_A_IWLYgiZ98_0;
	wire w_dff_A_CxcAPjgn3_0;
	wire w_dff_A_gSzj3tVD3_0;
	wire w_dff_A_mLO9Rlle0_0;
	wire w_dff_A_urBtdoC78_0;
	wire w_dff_A_oGNZ1BnE3_0;
	wire w_dff_A_BcXW1JCM7_0;
	wire w_dff_A_eyi3NToG8_0;
	wire w_dff_A_7y8vWWbu7_0;
	wire w_dff_A_DPDstFdz3_0;
	wire w_dff_A_kph5iynj7_0;
	wire w_dff_A_xHuqdW4u4_0;
	wire w_dff_A_l4n1jSio7_0;
	wire w_dff_A_9Z9W60q11_0;
	wire w_dff_A_OITfyRiK1_0;
	wire w_dff_A_mzda089A1_0;
	wire w_dff_A_WEcZ2iW12_0;
	wire w_dff_A_fWvJ53HN4_0;
	wire w_dff_A_HMXV228V9_0;
	wire w_dff_A_5GFHkcEq5_0;
	wire w_dff_A_Pjx5uvvz8_2;
	wire w_dff_A_kNXwVVQk5_0;
	wire w_dff_A_Hxt8a4OA8_0;
	wire w_dff_A_v6VoS3YZ6_0;
	wire w_dff_A_6jjTL19g2_0;
	wire w_dff_A_9NcwBcff5_0;
	wire w_dff_A_qXcqqucO9_0;
	wire w_dff_A_bfsNheRL0_0;
	wire w_dff_A_2TS8YV1G2_0;
	wire w_dff_A_P2jtaxxK0_0;
	wire w_dff_A_Opu76JVi5_0;
	wire w_dff_A_7kR1rqoC4_0;
	wire w_dff_A_xChkfXOo9_0;
	wire w_dff_A_CJ41juEX8_0;
	wire w_dff_A_gH9byscB2_0;
	wire w_dff_A_wcao1Hsz5_0;
	wire w_dff_A_rB6i93TA9_0;
	wire w_dff_A_CNjFLDeT7_0;
	wire w_dff_A_CZDy6jk95_0;
	wire w_dff_A_eU16c4oW0_0;
	wire w_dff_A_d03moyHC8_0;
	wire w_dff_A_jP557fHe5_0;
	wire w_dff_A_IfH9F0ig3_0;
	wire w_dff_A_tn1EyM9i3_2;
	wire w_dff_A_2jhrJeQb9_0;
	wire w_dff_A_hdL1ACui3_0;
	wire w_dff_A_7cAUZ44P4_0;
	wire w_dff_A_8u62kS8E6_0;
	wire w_dff_A_iOSMhwi01_0;
	wire w_dff_A_wOn50Mqd4_0;
	wire w_dff_A_RNp7315i2_0;
	wire w_dff_A_7P2Ns1h92_0;
	wire w_dff_A_yboWpnap3_0;
	wire w_dff_A_ok0x16gL1_0;
	wire w_dff_A_paKelJtN5_0;
	wire w_dff_A_4i6WhpPq2_0;
	wire w_dff_A_cJka9j9i7_0;
	wire w_dff_A_HiTtZQB10_0;
	wire w_dff_A_iCbNs5643_0;
	wire w_dff_A_YVZP8Hit7_0;
	wire w_dff_A_dnCHc4FG7_0;
	wire w_dff_A_X7ha8v5G5_0;
	wire w_dff_A_wLlaiJpM4_0;
	wire w_dff_A_v75tMy0o0_0;
	wire w_dff_A_3vbDz3c77_0;
	wire w_dff_A_twN5M79m5_0;
	wire w_dff_A_61AsB52f5_0;
	wire w_dff_A_tKl0CTRg3_0;
	wire w_dff_A_WVLP6Vxk8_2;
	wire w_dff_A_PWgPFtjU2_0;
	wire w_dff_A_uMzpYxq58_0;
	wire w_dff_A_3fyKWzI73_0;
	wire w_dff_A_AdPmfEQb9_0;
	wire w_dff_A_2wN7WGGz8_0;
	wire w_dff_A_zo38pquS9_0;
	wire w_dff_A_xaHe7qAy0_0;
	wire w_dff_A_seNgpSMG8_0;
	wire w_dff_A_DkpRyY655_0;
	wire w_dff_A_93sfPJ2V6_0;
	wire w_dff_A_rRBfyQMw1_0;
	wire w_dff_A_F0ncmQOy0_0;
	wire w_dff_A_p6Xv2Vj36_0;
	wire w_dff_A_roSWSQVY7_0;
	wire w_dff_A_3fhK9Hho3_0;
	wire w_dff_A_38EjjIEu3_0;
	wire w_dff_A_nDeH3VAR4_0;
	wire w_dff_A_OAwbyRkb3_0;
	wire w_dff_A_crCyPbkk3_0;
	wire w_dff_A_td5plFan6_0;
	wire w_dff_A_2mxWfBNh4_0;
	wire w_dff_A_lXlBCIey5_0;
	wire w_dff_A_Yj8tPGme5_0;
	wire w_dff_A_RghVUsn29_0;
	wire w_dff_A_f3B3tmMs4_2;
	wire w_dff_A_3vO6cYus4_0;
	wire w_dff_A_f4jjXWyO5_0;
	wire w_dff_A_zseyeVDx1_0;
	wire w_dff_A_rSMSIBmD0_0;
	wire w_dff_A_hYlZPvfI3_0;
	wire w_dff_A_3qK4F6kU9_0;
	wire w_dff_A_varSMzUI0_0;
	wire w_dff_A_lAkQP9w03_0;
	wire w_dff_A_nAITM0H65_0;
	wire w_dff_A_53GLPONo1_0;
	wire w_dff_A_OxOrGcbc3_0;
	wire w_dff_A_HFFcodYn2_0;
	wire w_dff_A_d3XfeB2A4_0;
	wire w_dff_A_WXqRxgAq9_0;
	wire w_dff_A_TAlcihmq7_0;
	wire w_dff_A_PDajkseE6_0;
	wire w_dff_A_xR2ntWuf3_0;
	wire w_dff_A_Ot6ZQt8L0_0;
	wire w_dff_A_cCjI2IwX6_0;
	wire w_dff_A_DlHsNY8J4_0;
	wire w_dff_A_kXFTkjuy4_0;
	wire w_dff_A_YNeUI7727_0;
	wire w_dff_A_M1qiqP2D8_0;
	wire w_dff_A_zpcNDc227_0;
	wire w_dff_A_zLSryDsq1_2;
	wire w_dff_A_X9BNpIy34_0;
	wire w_dff_A_ggggMBR32_0;
	wire w_dff_A_SAoG3qgB6_0;
	wire w_dff_A_1nbfXsTM0_0;
	wire w_dff_A_0XY46UUv1_0;
	wire w_dff_A_GphiGjuU7_0;
	wire w_dff_A_r6okzc7v7_0;
	wire w_dff_A_jMTnckTl7_0;
	wire w_dff_A_Yp44VbbJ0_0;
	wire w_dff_A_F3RrdjPz0_0;
	wire w_dff_A_Kk9XY2NS7_0;
	wire w_dff_A_dqJDGKUL5_0;
	wire w_dff_A_qvca6MJE9_0;
	wire w_dff_A_hFrwHAby2_0;
	wire w_dff_A_9ia8pK5b7_0;
	wire w_dff_A_f66Zlgwn4_0;
	wire w_dff_A_L8Iev85q9_0;
	wire w_dff_A_W9kaoHXd6_0;
	wire w_dff_A_e1IPzIUv1_0;
	wire w_dff_A_QvYRI3Qy8_0;
	wire w_dff_A_4TCN0c4I8_0;
	wire w_dff_A_p17Oa3ES5_0;
	wire w_dff_A_9OczA3Qo7_0;
	wire w_dff_A_MNV2tNp50_0;
	wire w_dff_A_ztAzJqOG4_0;
	wire w_dff_A_eJuXV8JT9_2;
	wire w_dff_A_NLYbL3sp8_0;
	wire w_dff_A_mecAV2dE2_0;
	wire w_dff_A_OspmI1xt8_0;
	wire w_dff_A_Kueb2dXJ4_0;
	wire w_dff_A_MMf1I3c55_0;
	wire w_dff_A_LoDKSHCH3_0;
	wire w_dff_A_9EmlGL5Z7_0;
	wire w_dff_A_xICStOLo1_0;
	wire w_dff_A_a4CYGuR08_0;
	wire w_dff_A_mBriqa6r7_0;
	wire w_dff_A_XSw3uw2i4_0;
	wire w_dff_A_25QxoFKl7_0;
	wire w_dff_A_Tcvo3xgU1_0;
	wire w_dff_A_ncoFE3At2_0;
	wire w_dff_A_LKN1qEfb6_0;
	wire w_dff_A_VvNGi9QZ6_0;
	wire w_dff_A_5905t9GQ3_0;
	wire w_dff_A_hgghZ0xo4_0;
	wire w_dff_A_JgolRGYL7_0;
	wire w_dff_A_Kg3BixOI0_0;
	wire w_dff_A_3LzS4Le53_0;
	wire w_dff_A_JNC0STpk8_0;
	wire w_dff_A_okknghdw6_1;
	wire w_dff_A_BbMXuhmh8_0;
	wire w_dff_A_PlmPaojf1_0;
	wire w_dff_A_xmbYEDkx2_0;
	wire w_dff_A_eOA6Pwj32_0;
	wire w_dff_A_glXFxzKQ9_0;
	wire w_dff_A_RZ6mZWeL9_0;
	wire w_dff_A_ZYHfgCxj7_0;
	wire w_dff_A_qS7pJICS4_0;
	wire w_dff_A_HEItSyrG1_0;
	wire w_dff_A_WSWvwix68_0;
	wire w_dff_A_TXcrylQe7_0;
	wire w_dff_A_zciIJX5T0_0;
	wire w_dff_A_eMkvwg2O6_0;
	wire w_dff_A_Tre5AUZR5_0;
	wire w_dff_A_2LlgYQZT8_0;
	wire w_dff_A_LK2iKSf28_0;
	wire w_dff_A_MJJPlJeh2_0;
	wire w_dff_A_VaY9n6zX4_0;
	wire w_dff_A_0wgGH0mP9_0;
	wire w_dff_A_heyu5tkl4_0;
	wire w_dff_A_DIc8uGqI6_0;
	wire w_dff_A_TJ3o8bmC6_0;
	wire w_dff_A_auIwklQa2_0;
	wire w_dff_A_MyMSigOS3_0;
	wire w_dff_A_JPpWur601_0;
	wire w_dff_A_SKkp85xP3_2;
	wire w_dff_A_cc31PMoT9_0;
	wire w_dff_A_9GZ1hK3I0_0;
	wire w_dff_A_4RkgZDEY2_0;
	wire w_dff_A_zDnCm8nu0_0;
	wire w_dff_A_ISbHSzu51_0;
	wire w_dff_A_zM8TL5qy7_0;
	wire w_dff_A_NbgrN2uM2_0;
	wire w_dff_A_oWrModiM8_0;
	wire w_dff_A_zj0JWWbJ9_0;
	wire w_dff_A_wpwEF8NO8_0;
	wire w_dff_A_Zgrdx8975_0;
	wire w_dff_A_uJSpuao87_0;
	wire w_dff_A_W6OqyxXw8_0;
	wire w_dff_A_oxz5g3aZ4_0;
	wire w_dff_A_sk6ExhNv7_0;
	wire w_dff_A_2hSo6UjF9_0;
	wire w_dff_A_gslfoMKd5_0;
	wire w_dff_A_YbN9g6Lz3_0;
	wire w_dff_A_lyd6BDC26_0;
	wire w_dff_A_Cy9RN5Ea9_0;
	wire w_dff_A_4acUKDlH8_0;
	wire w_dff_A_xPmhi39g0_0;
	wire w_dff_A_35oqKIZp5_2;
	wire w_dff_A_iaTm8Ie48_0;
	wire w_dff_A_BkKoa1Aj0_0;
	wire w_dff_A_ncJ6leYY4_0;
	wire w_dff_A_yRCu0ZN53_0;
	wire w_dff_A_86ZZKC897_0;
	wire w_dff_A_9yLVeOEW4_0;
	wire w_dff_A_NoBSmdu83_0;
	wire w_dff_A_EQv6kdJ69_0;
	wire w_dff_A_49GhB9GP3_0;
	wire w_dff_A_NejYa9Hm4_0;
	wire w_dff_A_mwi356Ei5_0;
	wire w_dff_A_4UK8dmLU4_0;
	wire w_dff_A_YjvQG4Vb9_0;
	wire w_dff_A_xMjtTQtq5_0;
	wire w_dff_A_xZBRDJea5_0;
	wire w_dff_A_8VmaL1QW4_0;
	wire w_dff_A_aLy163v86_0;
	wire w_dff_A_JLpcIygJ6_0;
	wire w_dff_A_JRNZfyNX8_0;
	wire w_dff_A_DUn2SYoX2_0;
	wire w_dff_A_SVIyMXnD0_0;
	wire w_dff_A_wMOjNUqD0_0;
	wire w_dff_A_XzrLJwvU7_2;
	wire w_dff_A_WGsUVzCW5_0;
	wire w_dff_A_f5vfj9Lo2_0;
	wire w_dff_A_GjJAyAxn3_0;
	wire w_dff_A_zf5aOjMK3_0;
	wire w_dff_A_fdnWkuQj8_0;
	wire w_dff_A_Vhcm3Vsi0_0;
	wire w_dff_A_xDrrMfif8_0;
	wire w_dff_A_n8DNWQXD0_0;
	wire w_dff_A_1PIGjyax6_0;
	wire w_dff_A_U4tjKopR2_0;
	wire w_dff_A_uPnkL4H75_0;
	wire w_dff_A_fRe3ziQ83_0;
	wire w_dff_A_nXQt28No0_0;
	wire w_dff_A_MR4rYd8Y2_0;
	wire w_dff_A_57kI9jKK2_0;
	wire w_dff_A_LJz7AEag5_0;
	wire w_dff_A_H1u2yFCu8_0;
	wire w_dff_A_hEiuQsy60_0;
	wire w_dff_A_Jp7BKBcE8_0;
	wire w_dff_A_JO5z6CfR0_0;
	wire w_dff_A_cjQoounO9_0;
	wire w_dff_A_nwMOwfqC9_0;
	wire w_dff_A_AVNYSklC9_0;
	wire w_dff_A_QCDFiWI29_0;
	wire w_dff_A_0PMn0hJB0_0;
	wire w_dff_A_GfrfYs7c3_2;
	wire w_dff_A_bOVUXuoD0_0;
	wire w_dff_A_Tt5IM3gC2_0;
	wire w_dff_A_vJllNvW37_0;
	wire w_dff_A_anvMCwWk5_0;
	wire w_dff_A_9ZpPBmDb3_0;
	wire w_dff_A_T13WJN8i9_0;
	wire w_dff_A_eB7DEgd49_0;
	wire w_dff_A_AS7pQGWR3_0;
	wire w_dff_A_LyhT3Z584_0;
	wire w_dff_A_6omjgayz8_0;
	wire w_dff_A_bwdaUsn80_0;
	wire w_dff_A_YdgMZpal5_0;
	wire w_dff_A_6I9W7B382_0;
	wire w_dff_A_lF7573D76_0;
	wire w_dff_A_HKn00WHx4_0;
	wire w_dff_A_Ki16IQvh5_0;
	wire w_dff_A_Os2j3Xf64_0;
	wire w_dff_A_kjS6n2Tj3_0;
	wire w_dff_A_OvIHAtGE4_0;
	wire w_dff_A_6DChSZZH1_0;
	wire w_dff_A_z77Qdrzb2_0;
	wire w_dff_A_tNGgaUHW5_0;
	wire w_dff_A_aqqygrba0_0;
	wire w_dff_A_V2xBhqVi9_2;
	wire w_dff_A_UhEno39s5_0;
	wire w_dff_A_H6ADwYna4_0;
	wire w_dff_A_UcMitI1C7_0;
	wire w_dff_A_aSVkd4Ff7_0;
	wire w_dff_A_1oP9gFMZ7_0;
	wire w_dff_A_OLmp3Pkl3_0;
	wire w_dff_A_cRGSIDc77_0;
	wire w_dff_A_k0rs1XpL1_0;
	wire w_dff_A_08Ksdl6U1_0;
	wire w_dff_A_5DBO5nBd9_0;
	wire w_dff_A_GnLSMS6k0_0;
	wire w_dff_A_YSOOJHDj7_0;
	wire w_dff_A_PqsA697P7_0;
	wire w_dff_A_u0ogulA74_0;
	wire w_dff_A_lJjyH7pR1_0;
	wire w_dff_A_GB8OJbKW5_0;
	wire w_dff_A_0VkPOqun0_0;
	wire w_dff_A_rTlckvfX8_0;
	wire w_dff_A_yJLFYMXo8_0;
	wire w_dff_A_W0LjnJ1Y3_0;
	wire w_dff_A_K9AScd5x5_0;
	wire w_dff_A_PdT8HLSw6_0;
	wire w_dff_A_rMOKO8Va0_0;
	wire w_dff_A_mActxA1q1_2;
	wire w_dff_A_mpNryBtD7_0;
	wire w_dff_A_lRTd2kHq2_0;
	wire w_dff_A_RO5XnqGe0_0;
	wire w_dff_A_ja5ECaDl7_0;
	wire w_dff_A_RujbHO2T6_0;
	wire w_dff_A_9MvXUAwN6_0;
	wire w_dff_A_ObNNLjWz3_0;
	wire w_dff_A_Q85dHfFR8_0;
	wire w_dff_A_CJ7l9IIl9_0;
	wire w_dff_A_vJ2mjGAW2_0;
	wire w_dff_A_EqBCNLti8_0;
	wire w_dff_A_3bWZAoto9_0;
	wire w_dff_A_60dQ0vME0_2;
	wire w_dff_A_FxINdpY90_0;
	wire w_dff_A_LAPyEJzi7_0;
	wire w_dff_A_cFpF1vaT8_0;
	wire w_dff_A_PigixGgt4_0;
	wire w_dff_A_3WOGSuKH6_0;
	wire w_dff_A_Tk06FzEK8_0;
	wire w_dff_A_mQZdZmLF8_0;
	wire w_dff_A_wy9iCPNA8_2;
	wire w_dff_A_CR6Atpxz3_0;
	wire w_dff_A_aiGWq3Ct5_0;
	wire w_dff_A_5AvoXO3C0_0;
	wire w_dff_A_Jekc0ell4_0;
	wire w_dff_A_EGaa7CQv5_0;
	wire w_dff_A_GkhGHBf64_0;
	wire w_dff_A_DtDmt0P51_0;
	wire w_dff_A_JMvGVQtW8_0;
	wire w_dff_A_F0uIHKDW3_0;
	wire w_dff_A_Sdrq4YvS9_2;
	wire w_dff_A_o1bfOnu03_0;
	wire w_dff_A_PwAQE4pJ6_0;
	wire w_dff_A_nNYK5rPu9_0;
	wire w_dff_A_b6zPkQoE0_0;
	wire w_dff_A_gyIhbuSH0_0;
	wire w_dff_A_sM8YiyDE4_0;
	wire w_dff_A_viukNfvi6_0;
	wire w_dff_A_N3sOEtk88_0;
	wire w_dff_A_k2mXTqrK8_0;
	wire w_dff_A_3DTwPGHW6_0;
	wire w_dff_A_mZEP9Xyo0_0;
	wire w_dff_A_qYIxtJuD1_2;
	wire w_dff_A_o4YoZEAw8_0;
	wire w_dff_A_gyc3Cwpg3_2;
	wire w_dff_A_ZsT733M38_0;
	wire w_dff_A_0IjuXLnU4_0;
	wire w_dff_A_02VidGkE4_0;
	wire w_dff_A_8ipjTEtQ4_0;
	wire w_dff_A_OP8VKc2T4_2;
	wire w_dff_A_ntucOagn6_0;
	wire w_dff_A_Ddccxeqd0_2;
	wire w_dff_A_FnkDKaHR4_0;
	wire w_dff_A_8gLXGBeE6_0;
	wire w_dff_A_rk1Nj5926_0;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(w_dff_A_c5h1KxxZ5_2),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(w_dff_A_YHZgzuPt7_2),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(w_dff_A_5rAfykWU6_2),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_n92_0[1]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_G17gat_2[2]),.dout(w_dff_A_9uEusv4s6_2),.clk(gclk));
	jnot g009(.din(w_G17gat_2[1]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G13gat_0[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G1gat_1[0]),.dout(n97),.clk(gclk));
	jnot g012(.din(w_G26gat_0[1]),.dout(n98),.clk(gclk));
	jor g013(.dina(n98),.dinb(w_n97_0[1]),.dout(n99),.clk(gclk));
	jor g014(.dina(w_n99_0[1]),.dinb(n96),.dout(n100),.clk(gclk));
	jor g015(.dina(n100),.dinb(w_n95_0[2]),.dout(n101),.clk(gclk));
	jor g016(.dina(w_n101_0[1]),.dinb(w_G390gat_0[1]),.dout(w_dff_A_Pjx5uvvz8_2),.clk(gclk));
	jnot g017(.din(w_G80gat_0[1]),.dout(n103),.clk(gclk));
	jand g018(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n104),.clk(gclk));
	jnot g019(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jor g020(.dina(n105),.dinb(w_n103_0[1]),.dout(w_dff_A_tn1EyM9i3_2),.clk(gclk));
	jnot g021(.din(w_G36gat_0[0]),.dout(n107),.clk(gclk));
	jnot g022(.din(w_G59gat_1[0]),.dout(n108),.clk(gclk));
	jor g023(.dina(w_n108_0[1]),.dinb(n107),.dout(n109),.clk(gclk));
	jor g024(.dina(w_n109_0[1]),.dinb(w_n103_0[0]),.dout(w_dff_A_WVLP6Vxk8_2),.clk(gclk));
	jnot g025(.din(w_G42gat_1[2]),.dout(n111),.clk(gclk));
	jor g026(.dina(w_n109_0[0]),.dinb(w_n111_0[1]),.dout(w_dff_A_f3B3tmMs4_2),.clk(gclk));
	jor g027(.dina(G88gat),.dinb(G87gat),.dout(n113),.clk(gclk));
	jand g028(.dina(w_n113_0[1]),.dinb(w_dff_B_31NqMquM7_1),.dout(w_dff_A_zLSryDsq1_2),.clk(gclk));
	jnot g029(.din(w_G390gat_0[0]),.dout(n115),.clk(gclk));
	jor g030(.dina(w_n101_0[0]),.dinb(w_dff_B_898klcWp2_1),.dout(w_dff_A_eJuXV8JT9_2),.clk(gclk));
	jand g031(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g033(.dina(w_n93_0[0]),.dinb(w_G55gat_0[2]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_n119_0[2]),.dinb(w_G29gat_0[0]),.dout(n120),.clk(gclk));
	jand g035(.dina(n120),.dinb(w_G68gat_0[1]),.dout(w_dff_A_SKkp85xP3_2),.clk(gclk));
	jand g036(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n122),.clk(gclk));
	jand g037(.dina(w_n119_0[1]),.dinb(G74gat),.dout(n123),.clk(gclk));
	jand g038(.dina(n123),.dinb(w_n122_0[1]),.dout(w_dff_A_35oqKIZp5_2),.clk(gclk));
	jand g039(.dina(w_n113_0[0]),.dinb(w_dff_B_ebNhaN5W2_1),.dout(w_dff_A_XzrLJwvU7_2),.clk(gclk));
	jxor g040(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n126),.clk(gclk));
	jxor g041(.dina(n126),.dinb(G135gat),.dout(n127),.clk(gclk));
	jxor g042(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n128),.clk(gclk));
	jxor g043(.dina(n128),.dinb(w_G130gat_0[1]),.dout(n129),.clk(gclk));
	jxor g044(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G126gat_0[2]),.dinb(w_G121gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(n131),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n129),.dout(n133),.clk(gclk));
	jxor g048(.dina(n133),.dinb(w_dff_B_CPF8Woo24_1),.dout(w_dff_A_GfrfYs7c3_2),.clk(gclk));
	jxor g049(.dina(w_G189gat_2[1]),.dinb(w_G183gat_1[2]),.dout(n135),.clk(gclk));
	jxor g050(.dina(n135),.dinb(G207gat),.dout(n136),.clk(gclk));
	jxor g051(.dina(w_G159gat_1[2]),.dinb(w_G130gat_0[0]),.dout(n137),.clk(gclk));
	jxor g052(.dina(n137),.dinb(w_G165gat_1[2]),.dout(n138),.clk(gclk));
	jxor g053(.dina(w_G177gat_1[2]),.dinb(w_G171gat_1[2]),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G201gat_1[1]),.dinb(w_G195gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n138),.dout(n142),.clk(gclk));
	jxor g057(.dina(n142),.dinb(w_dff_B_cLth2hkf3_1),.dout(w_dff_A_V2xBhqVi9_2),.clk(gclk));
	jnot g058(.din(w_G268gat_0[1]),.dout(n144),.clk(gclk));
	jand g059(.dina(w_G447gat_1),.dinb(w_G80gat_0[0]),.dout(n145),.clk(gclk));
	jand g060(.dina(n145),.dinb(w_n86_0[0]),.dout(n146),.clk(gclk));
	jand g061(.dina(w_n146_0[1]),.dinb(w_G55gat_0[1]),.dout(n147),.clk(gclk));
	jand g062(.dina(n147),.dinb(w_n144_0[1]),.dout(n148),.clk(gclk));
	jand g063(.dina(w_n111_0[0]),.dinb(w_n95_0[1]),.dout(n149),.clk(gclk));
	jnot g064(.din(w_n149_0[1]),.dout(n150),.clk(gclk));
	jand g065(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(w_G42gat_1[1]),.dinb(w_G17gat_2[0]),.dout(n152),.clk(gclk));
	jnot g067(.din(w_n152_0[1]),.dout(n153),.clk(gclk));
	jand g068(.dina(n153),.dinb(w_n151_0[1]),.dout(n154),.clk(gclk));
	jand g069(.dina(n154),.dinb(w_G447gat_0[2]),.dout(n155),.clk(gclk));
	jand g070(.dina(n155),.dinb(w_dff_B_X2HSRZXt6_1),.dout(n156),.clk(gclk));
	jnot g071(.din(w_n92_0[0]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n104_0[0]),.dinb(w_G42gat_1[0]),.dout(n158),.clk(gclk));
	jand g073(.dina(w_G51gat_1[0]),.dinb(w_G17gat_1[2]),.dout(n159),.clk(gclk));
	jnot g074(.din(n159),.dout(n160),.clk(gclk));
	jor g075(.dina(n160),.dinb(n158),.dout(n161),.clk(gclk));
	jor g076(.dina(n161),.dinb(n157),.dout(n162),.clk(gclk));
	jnot g077(.din(w_n162_0[1]),.dout(n163),.clk(gclk));
	jor g078(.dina(n163),.dinb(n156),.dout(n164),.clk(gclk));
	jand g079(.dina(w_n164_3[1]),.dinb(w_G126gat_0[1]),.dout(n165),.clk(gclk));
	jnot g080(.din(w_G156gat_0[0]),.dout(n166),.clk(gclk));
	jor g081(.dina(n166),.dinb(w_n108_0[0]),.dout(n167),.clk(gclk));
	jand g082(.dina(w_n167_0[1]),.dinb(w_G447gat_0[1]),.dout(n168),.clk(gclk));
	jand g083(.dina(w_n168_0[1]),.dinb(w_G17gat_1[1]),.dout(n169),.clk(gclk));
	jor g084(.dina(n169),.dinb(w_n97_0[0]),.dout(n170),.clk(gclk));
	jand g085(.dina(w_n170_1[1]),.dinb(w_G153gat_0[2]),.dout(n171),.clk(gclk));
	jor g086(.dina(w_dff_B_Ymb89kTl0_0),.dinb(n165),.dout(n172),.clk(gclk));
	jor g087(.dina(n172),.dinb(w_n148_1[2]),.dout(n173),.clk(gclk));
	jand g088(.dina(w_n173_0[1]),.dinb(w_G246gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_n122_0[0]),.dinb(w_G42gat_0[2]),.dout(n175),.clk(gclk));
	jand g090(.dina(G73gat),.dinb(G72gat),.dout(n176),.clk(gclk));
	jand g091(.dina(n176),.dinb(n175),.dout(n177),.clk(gclk));
	jand g092(.dina(n177),.dinb(w_n119_0[0]),.dout(n178),.clk(gclk));
	jand g093(.dina(w_n178_3[1]),.dinb(w_G201gat_1[0]),.dout(n179),.clk(gclk));
	jor g094(.dina(w_dff_B_U2Ez93Tr9_0),.dinb(n174),.dout(n180),.clk(gclk));
	jnot g095(.din(w_G201gat_0[2]),.dout(n181),.clk(gclk));
	jnot g096(.din(w_n148_1[1]),.dout(n182),.clk(gclk));
	jnot g097(.din(w_G126gat_0[0]),.dout(n183),.clk(gclk));
	jnot g098(.din(w_G51gat_0[2]),.dout(n184),.clk(gclk));
	jor g099(.dina(w_n99_0[0]),.dinb(n184),.dout(n185),.clk(gclk));
	jor g100(.dina(w_n152_0[0]),.dinb(w_n167_0[0]),.dout(n186),.clk(gclk));
	jor g101(.dina(n186),.dinb(w_n185_0[1]),.dout(n187),.clk(gclk));
	jor g102(.dina(n187),.dinb(w_n149_0[0]),.dout(n188),.clk(gclk));
	jand g103(.dina(w_n162_0[0]),.dinb(n188),.dout(n189),.clk(gclk));
	jor g104(.dina(n189),.dinb(n183),.dout(n190),.clk(gclk));
	jnot g105(.din(w_G153gat_0[1]),.dout(n191),.clk(gclk));
	jor g106(.dina(w_n151_0[0]),.dinb(w_n185_0[0]),.dout(n192),.clk(gclk));
	jor g107(.dina(n192),.dinb(w_n95_0[0]),.dout(n193),.clk(gclk));
	jand g108(.dina(n193),.dinb(w_G1gat_0[1]),.dout(n194),.clk(gclk));
	jor g109(.dina(n194),.dinb(n191),.dout(n195),.clk(gclk));
	jand g110(.dina(n195),.dinb(n190),.dout(n196),.clk(gclk));
	jand g111(.dina(n196),.dinb(w_dff_B_VKIL1KgJ4_1),.dout(n197),.clk(gclk));
	jxor g112(.dina(w_n197_0[2]),.dinb(w_n181_0[2]),.dout(n198),.clk(gclk));
	jand g113(.dina(w_n198_0[2]),.dinb(w_G228gat_3[1]),.dout(n199),.clk(gclk));
	jand g114(.dina(w_n173_0[0]),.dinb(w_G201gat_0[1]),.dout(n200),.clk(gclk));
	jand g115(.dina(w_n200_0[1]),.dinb(w_G237gat_3[1]),.dout(n201),.clk(gclk));
	jand g116(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n202),.clk(gclk));
	jand g117(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n203),.clk(gclk));
	jor g118(.dina(n203),.dinb(n202),.dout(n204),.clk(gclk));
	jor g119(.dina(w_dff_B_YOAELoHn9_0),.dinb(n201),.dout(n205),.clk(gclk));
	jor g120(.dina(n205),.dinb(w_dff_B_IW5aM6qg5_1),.dout(n206),.clk(gclk));
	jor g121(.dina(n206),.dinb(w_dff_B_whXXqEr29_1),.dout(n207),.clk(gclk));
	jor g122(.dina(w_n198_0[1]),.dinb(w_G261gat_0[2]),.dout(n208),.clk(gclk));
	jnot g123(.din(w_G261gat_0[1]),.dout(n209),.clk(gclk));
	jnot g124(.din(w_n198_0[0]),.dout(n210),.clk(gclk));
	jor g125(.dina(n210),.dinb(w_n209_0[1]),.dout(n211),.clk(gclk));
	jand g126(.dina(n211),.dinb(w_G219gat_3[2]),.dout(n212),.clk(gclk));
	jand g127(.dina(n212),.dinb(w_dff_B_LPpNpuYv6_1),.dout(n213),.clk(gclk));
	jor g128(.dina(n213),.dinb(n207),.dout(w_dff_A_mActxA1q1_2),.clk(gclk));
	jand g129(.dina(w_n164_3[0]),.dinb(w_G111gat_0[1]),.dout(n215),.clk(gclk));
	jand g130(.dina(w_n170_1[0]),.dinb(w_G143gat_0[1]),.dout(n216),.clk(gclk));
	jor g131(.dina(n216),.dinb(w_n148_1[0]),.dout(n217),.clk(gclk));
	jor g132(.dina(n217),.dinb(n215),.dout(n218),.clk(gclk));
	jxor g133(.dina(w_n218_1[1]),.dinb(w_G183gat_1[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n219_0[2]),.dinb(w_G228gat_3[0]),.dout(n220),.clk(gclk));
	jand g135(.dina(w_n178_3[0]),.dinb(w_G183gat_1[0]),.dout(n221),.clk(gclk));
	jand g136(.dina(w_n218_1[0]),.dinb(w_G183gat_0[2]),.dout(n222),.clk(gclk));
	jand g137(.dina(w_n222_0[2]),.dinb(w_G237gat_3[0]),.dout(n223),.clk(gclk));
	jand g138(.dina(w_n218_0[2]),.dinb(w_G246gat_3[0]),.dout(n224),.clk(gclk));
	jand g139(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n225),.clk(gclk));
	jor g140(.dina(w_dff_B_cmR8wiw80_0),.dinb(n224),.dout(n226),.clk(gclk));
	jor g141(.dina(n226),.dinb(n223),.dout(n227),.clk(gclk));
	jor g142(.dina(n227),.dinb(w_dff_B_FL9O8gPR8_1),.dout(n228),.clk(gclk));
	jor g143(.dina(n228),.dinb(w_dff_B_7gp16oMc7_1),.dout(n229),.clk(gclk));
	jand g144(.dina(w_n164_2[2]),.dinb(w_G116gat_0[1]),.dout(n230),.clk(gclk));
	jand g145(.dina(w_n170_0[2]),.dinb(w_G146gat_0[1]),.dout(n231),.clk(gclk));
	jor g146(.dina(n231),.dinb(w_n148_0[2]),.dout(n232),.clk(gclk));
	jor g147(.dina(n232),.dinb(n230),.dout(n233),.clk(gclk));
	jand g148(.dina(w_n233_1[1]),.dinb(w_G189gat_2[0]),.dout(n234),.clk(gclk));
	jor g149(.dina(w_n233_1[0]),.dinb(w_G189gat_1[2]),.dout(n235),.clk(gclk));
	jand g150(.dina(w_n164_2[1]),.dinb(w_G121gat_0[0]),.dout(n236),.clk(gclk));
	jand g151(.dina(w_n170_0[1]),.dinb(w_G149gat_0[1]),.dout(n237),.clk(gclk));
	jor g152(.dina(n237),.dinb(w_n148_0[1]),.dout(n238),.clk(gclk));
	jor g153(.dina(n238),.dinb(n236),.dout(n239),.clk(gclk));
	jand g154(.dina(w_n239_1[1]),.dinb(w_G195gat_2[0]),.dout(n240),.clk(gclk));
	jor g155(.dina(w_n239_1[0]),.dinb(w_G195gat_1[2]),.dout(n241),.clk(gclk));
	jand g156(.dina(w_n197_0[1]),.dinb(w_n181_0[1]),.dout(n242),.clk(gclk));
	jnot g157(.din(w_n242_0[1]),.dout(n243),.clk(gclk));
	jor g158(.dina(w_n200_0[0]),.dinb(w_G261gat_0[0]),.dout(n244),.clk(gclk));
	jand g159(.dina(n244),.dinb(n243),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n245_0[1]),.dinb(w_n241_0[1]),.dout(n246),.clk(gclk));
	jor g161(.dina(n246),.dinb(w_n240_0[1]),.dout(n247),.clk(gclk));
	jand g162(.dina(w_n247_0[1]),.dinb(w_n235_0[1]),.dout(n248),.clk(gclk));
	jor g163(.dina(n248),.dinb(w_n234_0[1]),.dout(n249),.clk(gclk));
	jor g164(.dina(w_n249_0[1]),.dinb(w_n219_0[1]),.dout(n250),.clk(gclk));
	jnot g165(.din(w_n219_0[0]),.dout(n251),.clk(gclk));
	jnot g166(.din(w_n234_0[0]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n235_0[0]),.dout(n253),.clk(gclk));
	jnot g168(.din(w_n240_0[0]),.dout(n254),.clk(gclk));
	jnot g169(.din(w_n241_0[0]),.dout(n255),.clk(gclk));
	jor g170(.dina(w_n197_0[0]),.dinb(w_n181_0[0]),.dout(n256),.clk(gclk));
	jand g171(.dina(n256),.dinb(w_n209_0[0]),.dout(n257),.clk(gclk));
	jor g172(.dina(n257),.dinb(w_n242_0[0]),.dout(n258),.clk(gclk));
	jor g173(.dina(w_n258_0[1]),.dinb(w_dff_B_1yNXocHa2_1),.dout(n259),.clk(gclk));
	jand g174(.dina(n259),.dinb(w_dff_B_zVRLC9Ba5_1),.dout(n260),.clk(gclk));
	jor g175(.dina(w_n260_0[1]),.dinb(w_dff_B_bjbKh9n43_1),.dout(n261),.clk(gclk));
	jand g176(.dina(n261),.dinb(w_dff_B_iqUzzj4d5_1),.dout(n262),.clk(gclk));
	jor g177(.dina(w_n262_0[1]),.dinb(w_dff_B_ZBXRjinY4_1),.dout(n263),.clk(gclk));
	jand g178(.dina(n263),.dinb(w_G219gat_3[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(n264),.dinb(w_dff_B_QpUcM2BV6_1),.dout(n265),.clk(gclk));
	jor g180(.dina(n265),.dinb(w_dff_B_vCCuB4CT6_1),.dout(w_dff_A_60dQ0vME0_2),.clk(gclk));
	jxor g181(.dina(w_n233_0[2]),.dinb(w_G189gat_1[1]),.dout(n267),.clk(gclk));
	jand g182(.dina(w_n267_0[2]),.dinb(w_G228gat_2[2]),.dout(n268),.clk(gclk));
	jand g183(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n269),.clk(gclk));
	jand g184(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n270),.clk(gclk));
	jor g185(.dina(n270),.dinb(w_G246gat_2[2]),.dout(n271),.clk(gclk));
	jand g186(.dina(w_dff_B_LiJqcHEa1_0),.dinb(w_n233_0[1]),.dout(n272),.clk(gclk));
	jor g187(.dina(n272),.dinb(w_dff_B_ogepBvZs6_1),.dout(n273),.clk(gclk));
	jand g188(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n274),.clk(gclk));
	jand g189(.dina(w_n178_2[2]),.dinb(w_G189gat_0[2]),.dout(n275),.clk(gclk));
	jor g190(.dina(n275),.dinb(n274),.dout(n276),.clk(gclk));
	jor g191(.dina(w_dff_B_gyWb3mQN5_0),.dinb(n273),.dout(n277),.clk(gclk));
	jor g192(.dina(n277),.dinb(w_dff_B_7Jcnxepb2_1),.dout(n278),.clk(gclk));
	jor g193(.dina(w_n267_0[1]),.dinb(w_n247_0[0]),.dout(n279),.clk(gclk));
	jnot g194(.din(w_n267_0[0]),.dout(n280),.clk(gclk));
	jor g195(.dina(w_dff_B_OdaqrOtz5_0),.dinb(w_n260_0[0]),.dout(n281),.clk(gclk));
	jand g196(.dina(n281),.dinb(w_G219gat_3[0]),.dout(n282),.clk(gclk));
	jand g197(.dina(n282),.dinb(w_dff_B_pzxGdjD11_1),.dout(n283),.clk(gclk));
	jor g198(.dina(n283),.dinb(w_dff_B_wJjuf0yv8_1),.dout(w_dff_A_wy9iCPNA8_2),.clk(gclk));
	jxor g199(.dina(w_n239_0[2]),.dinb(w_G195gat_1[1]),.dout(n285),.clk(gclk));
	jand g200(.dina(w_n285_0[2]),.dinb(w_G228gat_2[1]),.dout(n286),.clk(gclk));
	jand g201(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n287),.clk(gclk));
	jand g202(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n288),.clk(gclk));
	jor g203(.dina(n288),.dinb(w_G246gat_2[1]),.dout(n289),.clk(gclk));
	jand g204(.dina(w_dff_B_mC5ZY7pu3_0),.dinb(w_n239_0[1]),.dout(n290),.clk(gclk));
	jor g205(.dina(n290),.dinb(w_dff_B_AjMpcyz35_1),.dout(n291),.clk(gclk));
	jand g206(.dina(w_n178_2[1]),.dinb(w_G195gat_0[2]),.dout(n292),.clk(gclk));
	jand g207(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n293),.clk(gclk));
	jor g208(.dina(n293),.dinb(n292),.dout(n294),.clk(gclk));
	jor g209(.dina(w_dff_B_ebZatS749_0),.dinb(n291),.dout(n295),.clk(gclk));
	jor g210(.dina(n295),.dinb(w_dff_B_kP6EvrmH0_1),.dout(n296),.clk(gclk));
	jor g211(.dina(w_n285_0[1]),.dinb(w_n245_0[0]),.dout(n297),.clk(gclk));
	jnot g212(.din(w_n285_0[0]),.dout(n298),.clk(gclk));
	jor g213(.dina(w_dff_B_ENeW9ryo0_0),.dinb(w_n258_0[0]),.dout(n299),.clk(gclk));
	jand g214(.dina(n299),.dinb(w_G219gat_2[2]),.dout(n300),.clk(gclk));
	jand g215(.dina(n300),.dinb(w_dff_B_FAex2s4q4_1),.dout(n301),.clk(gclk));
	jor g216(.dina(n301),.dinb(w_dff_B_uX9nyNKO7_1),.dout(w_dff_A_Sdrq4YvS9_2),.clk(gclk));
	jand g217(.dina(w_n168_0[0]),.dinb(w_G55gat_0[0]),.dout(n303),.clk(gclk));
	jand g218(.dina(w_n303_1[1]),.dinb(w_G143gat_0[0]),.dout(n304),.clk(gclk));
	jand g219(.dina(w_n146_0[0]),.dinb(w_G17gat_1[0]),.dout(n305),.clk(gclk));
	jand g220(.dina(n305),.dinb(w_n144_0[0]),.dout(n306),.clk(gclk));
	jor g221(.dina(w_n306_1[1]),.dinb(w_dff_B_ZolByrk60_1),.dout(n307),.clk(gclk));
	jand g222(.dina(w_n164_2[0]),.dinb(w_G91gat_0[1]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n309),.clk(gclk));
	jor g224(.dina(w_dff_B_3ValmUWV0_0),.dinb(n308),.dout(n310),.clk(gclk));
	jor g225(.dina(n310),.dinb(w_dff_B_b71Job3Z5_1),.dout(n311),.clk(gclk));
	jand g226(.dina(w_n311_1[2]),.dinb(w_G159gat_1[1]),.dout(n312),.clk(gclk));
	jor g227(.dina(w_n311_1[1]),.dinb(w_G159gat_1[0]),.dout(n313),.clk(gclk));
	jand g228(.dina(w_n164_1[2]),.dinb(w_G96gat_0[1]),.dout(n314),.clk(gclk));
	jand g229(.dina(w_n303_1[0]),.dinb(w_G146gat_0[0]),.dout(n315),.clk(gclk));
	jand g230(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n316),.clk(gclk));
	jor g231(.dina(w_dff_B_Z9TYzfVw8_0),.dinb(n315),.dout(n317),.clk(gclk));
	jor g232(.dina(w_dff_B_kmBlNeDa0_0),.dinb(n314),.dout(n318),.clk(gclk));
	jor g233(.dina(n318),.dinb(w_n306_1[0]),.dout(n319),.clk(gclk));
	jand g234(.dina(w_n319_1[2]),.dinb(w_G165gat_1[1]),.dout(n320),.clk(gclk));
	jor g235(.dina(w_n319_1[1]),.dinb(w_G165gat_1[0]),.dout(n321),.clk(gclk));
	jand g236(.dina(w_n164_1[1]),.dinb(w_G101gat_0[1]),.dout(n322),.clk(gclk));
	jand g237(.dina(w_n303_0[2]),.dinb(w_G149gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n324),.clk(gclk));
	jor g239(.dina(w_dff_B_D33PHtD84_0),.dinb(n323),.dout(n325),.clk(gclk));
	jor g240(.dina(w_dff_B_XMZ4bwEE7_0),.dinb(n322),.dout(n326),.clk(gclk));
	jor g241(.dina(n326),.dinb(w_n306_0[2]),.dout(n327),.clk(gclk));
	jand g242(.dina(w_n327_1[2]),.dinb(w_G171gat_1[1]),.dout(n328),.clk(gclk));
	jor g243(.dina(w_n327_1[1]),.dinb(w_G171gat_1[0]),.dout(n329),.clk(gclk));
	jand g244(.dina(w_n164_1[0]),.dinb(w_G106gat_0[0]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n303_0[1]),.dinb(w_G153gat_0[0]),.dout(n331),.clk(gclk));
	jand g246(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n332),.clk(gclk));
	jor g247(.dina(w_dff_B_3mYVtRII6_0),.dinb(n331),.dout(n333),.clk(gclk));
	jor g248(.dina(w_dff_B_Adq0vX6W4_0),.dinb(n330),.dout(n334),.clk(gclk));
	jor g249(.dina(n334),.dinb(w_n306_0[1]),.dout(n335),.clk(gclk));
	jand g250(.dina(w_n335_1[1]),.dinb(w_G177gat_1[1]),.dout(n336),.clk(gclk));
	jnot g251(.din(w_G177gat_1[0]),.dout(n337),.clk(gclk));
	jnot g252(.din(w_n335_1[0]),.dout(n338),.clk(gclk));
	jand g253(.dina(n338),.dinb(w_dff_B_kH9XimPh4_1),.dout(n339),.clk(gclk));
	jnot g254(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jnot g255(.din(w_G183gat_0[1]),.dout(n341),.clk(gclk));
	jnot g256(.din(w_n218_0[1]),.dout(n342),.clk(gclk));
	jand g257(.dina(n342),.dinb(w_dff_B_jf0EZXZZ0_1),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n343_0[1]),.dout(n344),.clk(gclk));
	jand g259(.dina(w_n249_0[0]),.dinb(w_dff_B_cvIQccYk8_1),.dout(n345),.clk(gclk));
	jor g260(.dina(n345),.dinb(w_n222_0[1]),.dout(n346),.clk(gclk));
	jand g261(.dina(w_n346_0[1]),.dinb(w_dff_B_tybF7BoW7_1),.dout(n347),.clk(gclk));
	jor g262(.dina(n347),.dinb(w_n336_0[2]),.dout(n348),.clk(gclk));
	jand g263(.dina(w_n348_0[1]),.dinb(w_n329_0[1]),.dout(n349),.clk(gclk));
	jor g264(.dina(n349),.dinb(w_n328_0[1]),.dout(n350),.clk(gclk));
	jand g265(.dina(w_n350_0[1]),.dinb(w_n321_0[1]),.dout(n351),.clk(gclk));
	jor g266(.dina(n351),.dinb(w_n320_0[1]),.dout(n352),.clk(gclk));
	jand g267(.dina(w_n352_0[1]),.dinb(w_dff_B_uRMRSEKs8_1),.dout(n353),.clk(gclk));
	jor g268(.dina(n353),.dinb(w_dff_B_jQQigADs9_1),.dout(w_dff_A_qYIxtJuD1_2),.clk(gclk));
	jxor g269(.dina(w_n335_0[2]),.dinb(w_G177gat_0[2]),.dout(n355),.clk(gclk));
	jnot g270(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n346_0[0]),.dinb(w_G219gat_2[1]),.dout(n357),.clk(gclk));
	jand g272(.dina(n357),.dinb(w_dff_B_BLIkJKXs8_1),.dout(n358),.clk(gclk));
	jnot g273(.din(w_n222_0[0]),.dout(n359),.clk(gclk));
	jor g274(.dina(w_n262_0[0]),.dinb(w_n343_0[0]),.dout(n360),.clk(gclk));
	jand g275(.dina(n360),.dinb(w_dff_B_D2Y4UE0M3_1),.dout(n361),.clk(gclk));
	jand g276(.dina(w_n361_0[1]),.dinb(w_G219gat_2[0]),.dout(n362),.clk(gclk));
	jor g277(.dina(n362),.dinb(w_G228gat_2[0]),.dout(n363),.clk(gclk));
	jand g278(.dina(n363),.dinb(w_n355_0[0]),.dout(n364),.clk(gclk));
	jand g279(.dina(w_n336_0[1]),.dinb(w_G237gat_2[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_n335_0[1]),.dinb(w_G246gat_2[0]),.dout(n366),.clk(gclk));
	jand g281(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n367),.clk(gclk));
	jand g282(.dina(w_n178_2[0]),.dinb(w_G177gat_0[1]),.dout(n368),.clk(gclk));
	jor g283(.dina(n368),.dinb(n367),.dout(n369),.clk(gclk));
	jor g284(.dina(w_dff_B_Bs7DS11W5_0),.dinb(n366),.dout(n370),.clk(gclk));
	jor g285(.dina(n370),.dinb(n365),.dout(n371),.clk(gclk));
	jor g286(.dina(w_dff_B_kLpPMk8B5_0),.dinb(n364),.dout(n372),.clk(gclk));
	jor g287(.dina(n372),.dinb(w_dff_B_1Tv7GAvm9_1),.dout(w_dff_A_gyc3Cwpg3_2),.clk(gclk));
	jand g288(.dina(w_n311_1[0]),.dinb(w_G237gat_1[2]),.dout(n374),.clk(gclk));
	jor g289(.dina(n374),.dinb(w_n178_1[2]),.dout(n375),.clk(gclk));
	jand g290(.dina(n375),.dinb(w_G159gat_0[2]),.dout(n376),.clk(gclk));
	jxor g291(.dina(w_n311_0[2]),.dinb(w_G159gat_0[1]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_n377_0[2]),.dinb(w_G228gat_1[2]),.dout(n378),.clk(gclk));
	jand g293(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n379),.clk(gclk));
	jor g294(.dina(w_dff_B_oBmZdDdv8_0),.dinb(n378),.dout(n380),.clk(gclk));
	jand g295(.dina(w_n311_0[1]),.dinb(w_G246gat_1[2]),.dout(n381),.clk(gclk));
	jor g296(.dina(w_dff_B_rEqfqAFS6_0),.dinb(n380),.dout(n382),.clk(gclk));
	jor g297(.dina(n382),.dinb(w_dff_B_9u6nPr194_1),.dout(n383),.clk(gclk));
	jor g298(.dina(w_n377_0[1]),.dinb(w_n352_0[0]),.dout(n384),.clk(gclk));
	jnot g299(.din(w_n320_0[0]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n321_0[0]),.dout(n386),.clk(gclk));
	jnot g301(.din(w_n328_0[0]),.dout(n387),.clk(gclk));
	jnot g302(.din(w_n329_0[0]),.dout(n388),.clk(gclk));
	jnot g303(.din(w_n336_0[0]),.dout(n389),.clk(gclk));
	jor g304(.dina(w_n361_0[0]),.dinb(w_n339_0[0]),.dout(n390),.clk(gclk));
	jand g305(.dina(n390),.dinb(w_dff_B_BnHVhi8v1_1),.dout(n391),.clk(gclk));
	jor g306(.dina(w_n391_0[1]),.dinb(w_dff_B_HjtU3Aed2_1),.dout(n392),.clk(gclk));
	jand g307(.dina(n392),.dinb(w_dff_B_FXd0XQD89_1),.dout(n393),.clk(gclk));
	jor g308(.dina(w_n393_0[1]),.dinb(w_dff_B_kXtpPMaG3_1),.dout(n394),.clk(gclk));
	jand g309(.dina(n394),.dinb(w_dff_B_uC21U4j09_1),.dout(n395),.clk(gclk));
	jnot g310(.din(w_n377_0[0]),.dout(n396),.clk(gclk));
	jor g311(.dina(w_dff_B_p8dNjgNM2_0),.dinb(n395),.dout(n397),.clk(gclk));
	jand g312(.dina(n397),.dinb(w_G219gat_1[2]),.dout(n398),.clk(gclk));
	jand g313(.dina(n398),.dinb(w_dff_B_j1jZDTRW8_1),.dout(n399),.clk(gclk));
	jor g314(.dina(n399),.dinb(w_dff_B_cwtaCgur6_1),.dout(G878gat),.clk(gclk));
	jand g315(.dina(w_n319_1[0]),.dinb(w_G237gat_1[1]),.dout(n401),.clk(gclk));
	jor g316(.dina(n401),.dinb(w_n178_1[1]),.dout(n402),.clk(gclk));
	jand g317(.dina(n402),.dinb(w_G165gat_0[2]),.dout(n403),.clk(gclk));
	jxor g318(.dina(w_n319_0[2]),.dinb(w_G165gat_0[1]),.dout(n404),.clk(gclk));
	jand g319(.dina(w_n404_0[2]),.dinb(w_G228gat_1[1]),.dout(n405),.clk(gclk));
	jand g320(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n406),.clk(gclk));
	jor g321(.dina(w_dff_B_W5jbDRS45_0),.dinb(n405),.dout(n407),.clk(gclk));
	jand g322(.dina(w_n319_0[1]),.dinb(w_G246gat_1[1]),.dout(n408),.clk(gclk));
	jor g323(.dina(w_dff_B_k7CZ7hhD3_0),.dinb(n407),.dout(n409),.clk(gclk));
	jor g324(.dina(n409),.dinb(w_dff_B_KYrhI0hC1_1),.dout(n410),.clk(gclk));
	jor g325(.dina(w_n404_0[1]),.dinb(w_n350_0[0]),.dout(n411),.clk(gclk));
	jnot g326(.din(w_n404_0[0]),.dout(n412),.clk(gclk));
	jor g327(.dina(w_dff_B_U4V7GEKf5_0),.dinb(w_n393_0[0]),.dout(n413),.clk(gclk));
	jand g328(.dina(n413),.dinb(w_G219gat_1[1]),.dout(n414),.clk(gclk));
	jand g329(.dina(n414),.dinb(w_dff_B_kHNch1gY8_1),.dout(n415),.clk(gclk));
	jor g330(.dina(n415),.dinb(w_dff_B_GbNwPoWg2_1),.dout(w_dff_A_OP8VKc2T4_2),.clk(gclk));
	jand g331(.dina(w_n327_1[0]),.dinb(w_G237gat_1[0]),.dout(n417),.clk(gclk));
	jor g332(.dina(n417),.dinb(w_n178_1[0]),.dout(n418),.clk(gclk));
	jand g333(.dina(n418),.dinb(w_G171gat_0[2]),.dout(n419),.clk(gclk));
	jxor g334(.dina(w_n327_0[2]),.dinb(w_G171gat_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n420_0[2]),.dinb(w_G228gat_1[0]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jor g337(.dina(w_dff_B_fWNdO3uh7_0),.dinb(n421),.dout(n423),.clk(gclk));
	jand g338(.dina(w_n327_0[1]),.dinb(w_G246gat_1[0]),.dout(n424),.clk(gclk));
	jor g339(.dina(w_dff_B_DSR0Iwlk1_0),.dinb(n423),.dout(n425),.clk(gclk));
	jor g340(.dina(n425),.dinb(w_dff_B_2kQkNnHJ0_1),.dout(n426),.clk(gclk));
	jnot g341(.din(w_n420_0[1]),.dout(n427),.clk(gclk));
	jor g342(.dina(w_dff_B_eCn0yA8Z3_0),.dinb(w_n391_0[0]),.dout(n428),.clk(gclk));
	jor g343(.dina(w_n420_0[0]),.dinb(w_n348_0[0]),.dout(n429),.clk(gclk));
	jand g344(.dina(n429),.dinb(w_G219gat_1[0]),.dout(n430),.clk(gclk));
	jand g345(.dina(n430),.dinb(w_dff_B_mqO1nELF3_1),.dout(n431),.clk(gclk));
	jor g346(.dina(n431),.dinb(w_dff_B_kuM9YojE4_1),.dout(w_dff_A_Ddccxeqd0_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_G13gat_0[1]),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_G17gat_1[0]),.doutb(w_G17gat_1[1]),.doutc(w_G17gat_1[2]),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_G17gat_2[2]),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_G29gat_0[0]),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_G42gat_0[1]),.doutc(w_G42gat_0[2]),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_G42gat_1[0]),.doutb(w_G42gat_1[1]),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_G51gat_1[1]),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_G55gat_0[0]),.doutb(w_G55gat_0[1]),.doutc(w_G55gat_0[2]),.din(G55gat));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_G68gat_0[1]),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_G80gat_0[0]),.doutb(w_G80gat_0[1]),.doutc(w_G80gat_0[2]),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_G91gat_0[1]),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_G96gat_0[1]),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_G101gat_0[1]),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_G106gat_0[0]),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_G111gat_0[1]),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_G116gat_0[1]),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_G121gat_0[0]),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl3 jspl3_w_G126gat_0(.douta(w_G126gat_0[0]),.doutb(w_G126gat_0[1]),.doutc(w_G126gat_0[2]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_G130gat_0[1]),.din(G130gat));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_dff_A_z7MgNYZq9_1),.din(w_dff_B_XhZnIYUG3_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_dff_A_ktiDR8at9_1),.din(w_dff_B_oEo3lIF12_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_dff_A_GMKVTrYB1_1),.din(w_dff_B_dNetj7Sz0_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_G153gat_0[0]),.doutb(w_G153gat_0[1]),.doutc(w_G153gat_0[2]),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_G159gat_0[1]),.doutc(w_G159gat_0[2]),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_G159gat_1[0]),.doutb(w_G159gat_1[1]),.doutc(w_G159gat_1[2]),.din(w_G159gat_0[0]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_G165gat_0[1]),.doutc(w_G165gat_0[2]),.din(G165gat));
	jspl3 jspl3_w_G165gat_1(.douta(w_G165gat_1[0]),.doutb(w_G165gat_1[1]),.doutc(w_G165gat_1[2]),.din(w_G165gat_0[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_G177gat_0[1]),.doutc(w_G177gat_0[2]),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_G177gat_1[1]),.doutc(w_G177gat_1[2]),.din(w_G177gat_0[0]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_G183gat_0[2]),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_G183gat_1[0]),.doutb(w_G183gat_1[1]),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_G189gat_0[2]),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_G189gat_1[1]),.doutc(w_G189gat_1[2]),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_G189gat_2[0]),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_G195gat_0[2]),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_G195gat_1[1]),.doutc(w_G195gat_1[2]),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_G195gat_2[0]),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_G201gat_0[1]),.doutc(w_G201gat_0[2]),.din(G201gat));
	jspl jspl_w_G201gat_1(.douta(w_G201gat_1[0]),.doutb(w_G201gat_1[1]),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_k8q9eGSe7_0),.doutb(w_dff_A_2HLhW8dn4_1),.doutc(w_G219gat_0[2]),.din(w_dff_B_HuHRgb4z3_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_G219gat_1[0]),.doutb(w_dff_A_RWZmEWs59_1),.doutc(w_dff_A_IYzUJds28_2),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_7eFcm9HF7_0),.doutb(w_dff_A_YnXncBJ56_1),.doutc(w_G219gat_2[2]),.din(w_G219gat_0[1]));
	jspl3 jspl3_w_G219gat_3(.douta(w_dff_A_gaBE8EBh3_0),.doutb(w_dff_A_Vs6wtd3O9_1),.doutc(w_G219gat_3[2]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_dff_A_gDQHMYla4_0),.doutb(w_G228gat_0[1]),.doutc(w_G228gat_0[2]),.din(w_dff_B_ZIZCD5EV5_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_dff_A_qHxwdpt16_0),.doutb(w_G228gat_2[1]),.doutc(w_G228gat_2[2]),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_dff_A_y8Eld7Ju7_1),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_G237gat_0[0]),.doutb(w_G237gat_0[1]),.doutc(w_G237gat_0[2]),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_G237gat_2[0]),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_dff_A_J0on60g63_1),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_G246gat_0[0]),.doutb(w_G246gat_0[1]),.doutc(w_G246gat_0[2]),.din(G246gat));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_G246gat_2[0]),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_dff_A_11az7EPc0_1),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_G261gat_0[0]),.doutb(w_G261gat_0[1]),.doutc(w_G261gat_0[2]),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_dff_A_93NRgkcP8_1),.doutc(w_dff_A_7Fl3brhr8_2),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_dff_A_ClR1RSNQ7_2),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(w_dff_A_okknghdw6_1),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_dff_A_hCZC8D6S0_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n95_0(.douta(w_n95_0[0]),.doutb(w_n95_0[1]),.doutc(w_n95_0[2]),.din(n95));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.din(w_dff_B_1CEGbPvb3_2));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.din(n113));
	jspl3 jspl3_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.doutc(w_n119_0[2]),.din(n119));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.din(n122));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(w_dff_B_hBYn5AJP7_2));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_n148_1[0]),.doutb(w_n148_1[1]),.doutc(w_dff_A_eyc1lp049_2),.din(w_n148_0[0]));
	jspl jspl_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.din(n149));
	jspl jspl_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_n164_0[2]),.din(n164));
	jspl3 jspl3_w_n164_1(.douta(w_n164_1[0]),.doutb(w_n164_1[1]),.doutc(w_n164_1[2]),.din(w_n164_0[0]));
	jspl3 jspl3_w_n164_2(.douta(w_n164_2[0]),.doutb(w_n164_2[1]),.doutc(w_n164_2[2]),.din(w_n164_0[1]));
	jspl jspl_w_n164_3(.douta(w_n164_3[0]),.doutb(w_n164_3[1]),.din(w_n164_0[2]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n170_1(.douta(w_n170_1[0]),.doutb(w_n170_1[1]),.din(w_n170_0[0]));
	jspl jspl_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.din(n173));
	jspl3 jspl3_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.doutc(w_n178_0[2]),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_n178_1[1]),.doutc(w_n178_1[2]),.din(w_n178_0[0]));
	jspl3 jspl3_w_n178_2(.douta(w_n178_2[0]),.doutb(w_n178_2[1]),.doutc(w_n178_2[2]),.din(w_n178_0[1]));
	jspl jspl_w_n178_3(.douta(w_n178_3[0]),.doutb(w_n178_3[1]),.din(w_n178_0[2]));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(w_dff_B_BEqYUOMv2_3));
	jspl jspl_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.din(n185));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_n198_0[2]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_dff_A_4cNoCPSg0_1),.din(w_dff_B_LL0ht2Ne4_2));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_n218_0[2]),.din(n218));
	jspl jspl_w_n218_1(.douta(w_n218_1[0]),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl3 jspl3_w_n219_0(.douta(w_n219_0[0]),.doutb(w_dff_A_WgetRk2g0_1),.doutc(w_n219_0[2]),.din(n219));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_dff_A_FEssNtyE2_1),.doutc(w_n222_0[2]),.din(n222));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl jspl_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.din(w_n233_0[0]));
	jspl jspl_w_n234_0(.douta(w_n234_0[0]),.doutb(w_dff_A_npFGjXrQ4_1),.din(n234));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_dff_A_0VkJRlpF6_1),.din(n235));
	jspl3 jspl3_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.doutc(w_n239_0[2]),.din(n239));
	jspl jspl_w_n239_1(.douta(w_n239_1[0]),.doutb(w_n239_1[1]),.din(w_n239_0[0]));
	jspl jspl_w_n240_0(.douta(w_n240_0[0]),.doutb(w_dff_A_Zzzc8CrR8_1),.din(n240));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_dff_A_ZuR8lNHC0_1),.din(n241));
	jspl jspl_w_n242_0(.douta(w_dff_A_E5k1HrQO9_0),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.din(n258));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl jspl_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_dff_A_5b2xuoH16_1),.doutc(w_n267_0[2]),.din(n267));
	jspl3 jspl3_w_n285_0(.douta(w_n285_0[0]),.doutb(w_dff_A_pkqm1NpZ6_1),.doutc(w_n285_0[2]),.din(n285));
	jspl3 jspl3_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.doutc(w_n303_0[2]),.din(n303));
	jspl jspl_w_n303_1(.douta(w_n303_1[0]),.doutb(w_n303_1[1]),.din(w_n303_0[0]));
	jspl3 jspl3_w_n306_0(.douta(w_n306_0[0]),.doutb(w_dff_A_W9ACGTnI8_1),.doutc(w_dff_A_2cGXA9CZ0_2),.din(n306));
	jspl jspl_w_n306_1(.douta(w_dff_A_D50Szkfz6_0),.doutb(w_n306_1[1]),.din(w_n306_0[0]));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.doutc(w_n311_0[2]),.din(n311));
	jspl3 jspl3_w_n311_1(.douta(w_n311_1[0]),.doutb(w_n311_1[1]),.doutc(w_n311_1[2]),.din(w_n311_0[0]));
	jspl3 jspl3_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.doutc(w_n319_0[2]),.din(n319));
	jspl3 jspl3_w_n319_1(.douta(w_n319_1[0]),.doutb(w_n319_1[1]),.doutc(w_n319_1[2]),.din(w_n319_0[0]));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_dff_A_QPcncT2h7_1),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_dff_A_BdvaWRgm5_1),.din(n321));
	jspl3 jspl3_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.doutc(w_n327_0[2]),.din(n327));
	jspl3 jspl3_w_n327_1(.douta(w_n327_1[0]),.doutb(w_n327_1[1]),.doutc(w_n327_1[2]),.din(w_n327_0[0]));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_dff_A_C0tNwMXZ7_1),.din(n328));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_dff_A_cY3IRWIR9_1),.din(n329));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl jspl_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.din(w_n335_0[0]));
	jspl3 jspl3_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.doutc(w_dff_A_I9q8PbWb9_2),.din(n336));
	jspl jspl_w_n339_0(.douta(w_dff_A_k9lRbkI00_0),.doutb(w_n339_0[1]),.din(n339));
	jspl jspl_w_n343_0(.douta(w_dff_A_xLgms4vS7_0),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n352_0(.douta(w_n352_0[0]),.doutb(w_n352_0[1]),.din(n352));
	jspl jspl_w_n355_0(.douta(w_dff_A_fs0rZYQO3_0),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_dff_A_Wm4FoYEo2_1),.doutc(w_n377_0[2]),.din(n377));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(n391));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_dff_A_xWZaWM6C1_1),.doutc(w_n404_0[2]),.din(n404));
	jspl3 jspl3_w_n420_0(.douta(w_dff_A_mAAVI44v4_0),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jdff dff_B_1CEGbPvb3_2(.din(n103),.dout(w_dff_B_1CEGbPvb3_2),.clk(gclk));
	jdff dff_B_31NqMquM7_1(.din(G90gat),.dout(w_dff_B_31NqMquM7_1),.clk(gclk));
	jdff dff_B_898klcWp2_1(.din(n115),.dout(w_dff_B_898klcWp2_1),.clk(gclk));
	jdff dff_A_RoEms7Ki0_1(.dout(w_G390gat_0[1]),.din(w_dff_A_RoEms7Ki0_1),.clk(gclk));
	jdff dff_A_93NRgkcP8_1(.dout(w_dff_A_RoEms7Ki0_1),.din(w_dff_A_93NRgkcP8_1),.clk(gclk));
	jdff dff_B_ebNhaN5W2_1(.din(G89gat),.dout(w_dff_B_ebNhaN5W2_1),.clk(gclk));
	jdff dff_B_CPF8Woo24_1(.din(n127),.dout(w_dff_B_CPF8Woo24_1),.clk(gclk));
	jdff dff_B_cLth2hkf3_1(.din(n136),.dout(w_dff_B_cLth2hkf3_1),.clk(gclk));
	jdff dff_B_yptoowMS6_1(.din(n208),.dout(w_dff_B_yptoowMS6_1),.clk(gclk));
	jdff dff_B_LPpNpuYv6_1(.din(w_dff_B_yptoowMS6_1),.dout(w_dff_B_LPpNpuYv6_1),.clk(gclk));
	jdff dff_B_UEMNSjmT2_1(.din(n180),.dout(w_dff_B_UEMNSjmT2_1),.clk(gclk));
	jdff dff_B_whXXqEr29_1(.din(w_dff_B_UEMNSjmT2_1),.dout(w_dff_B_whXXqEr29_1),.clk(gclk));
	jdff dff_B_IW5aM6qg5_1(.din(n199),.dout(w_dff_B_IW5aM6qg5_1),.clk(gclk));
	jdff dff_B_fVDOO5gV5_0(.din(n204),.dout(w_dff_B_fVDOO5gV5_0),.clk(gclk));
	jdff dff_B_mmcesAxq8_0(.din(w_dff_B_fVDOO5gV5_0),.dout(w_dff_B_mmcesAxq8_0),.clk(gclk));
	jdff dff_B_5hwMQP213_0(.din(w_dff_B_mmcesAxq8_0),.dout(w_dff_B_5hwMQP213_0),.clk(gclk));
	jdff dff_B_GcyP0NqW6_0(.din(w_dff_B_5hwMQP213_0),.dout(w_dff_B_GcyP0NqW6_0),.clk(gclk));
	jdff dff_B_gEBb9dRg0_0(.din(w_dff_B_GcyP0NqW6_0),.dout(w_dff_B_gEBb9dRg0_0),.clk(gclk));
	jdff dff_B_i783zhWw9_0(.din(w_dff_B_gEBb9dRg0_0),.dout(w_dff_B_i783zhWw9_0),.clk(gclk));
	jdff dff_B_VhHJXHd58_0(.din(w_dff_B_i783zhWw9_0),.dout(w_dff_B_VhHJXHd58_0),.clk(gclk));
	jdff dff_B_VwoFMJOR7_0(.din(w_dff_B_VhHJXHd58_0),.dout(w_dff_B_VwoFMJOR7_0),.clk(gclk));
	jdff dff_B_YOAELoHn9_0(.din(w_dff_B_VwoFMJOR7_0),.dout(w_dff_B_YOAELoHn9_0),.clk(gclk));
	jdff dff_B_Hs1qRRcX5_0(.din(n179),.dout(w_dff_B_Hs1qRRcX5_0),.clk(gclk));
	jdff dff_B_OkIX0lT05_0(.din(w_dff_B_Hs1qRRcX5_0),.dout(w_dff_B_OkIX0lT05_0),.clk(gclk));
	jdff dff_B_L3FYPAHp2_0(.din(w_dff_B_OkIX0lT05_0),.dout(w_dff_B_L3FYPAHp2_0),.clk(gclk));
	jdff dff_B_SjQqSxhC5_0(.din(w_dff_B_L3FYPAHp2_0),.dout(w_dff_B_SjQqSxhC5_0),.clk(gclk));
	jdff dff_B_U2Ez93Tr9_0(.din(w_dff_B_SjQqSxhC5_0),.dout(w_dff_B_U2Ez93Tr9_0),.clk(gclk));
	jdff dff_B_DzqD2APM0_1(.din(n229),.dout(w_dff_B_DzqD2APM0_1),.clk(gclk));
	jdff dff_B_ME7H3JVk1_1(.din(w_dff_B_DzqD2APM0_1),.dout(w_dff_B_ME7H3JVk1_1),.clk(gclk));
	jdff dff_B_iNXNHolu3_1(.din(w_dff_B_ME7H3JVk1_1),.dout(w_dff_B_iNXNHolu3_1),.clk(gclk));
	jdff dff_B_gAxZpEKN6_1(.din(w_dff_B_iNXNHolu3_1),.dout(w_dff_B_gAxZpEKN6_1),.clk(gclk));
	jdff dff_B_xlWS6p896_1(.din(w_dff_B_gAxZpEKN6_1),.dout(w_dff_B_xlWS6p896_1),.clk(gclk));
	jdff dff_B_vCCuB4CT6_1(.din(w_dff_B_xlWS6p896_1),.dout(w_dff_B_vCCuB4CT6_1),.clk(gclk));
	jdff dff_B_QpUcM2BV6_1(.din(n250),.dout(w_dff_B_QpUcM2BV6_1),.clk(gclk));
	jdff dff_B_bKe4wP4T8_1(.din(n251),.dout(w_dff_B_bKe4wP4T8_1),.clk(gclk));
	jdff dff_B_UnLTmpaN7_1(.din(w_dff_B_bKe4wP4T8_1),.dout(w_dff_B_UnLTmpaN7_1),.clk(gclk));
	jdff dff_B_NI0cE1AZ1_1(.din(w_dff_B_UnLTmpaN7_1),.dout(w_dff_B_NI0cE1AZ1_1),.clk(gclk));
	jdff dff_B_GnGBpPiK7_1(.din(w_dff_B_NI0cE1AZ1_1),.dout(w_dff_B_GnGBpPiK7_1),.clk(gclk));
	jdff dff_B_8EEViAgp5_1(.din(w_dff_B_GnGBpPiK7_1),.dout(w_dff_B_8EEViAgp5_1),.clk(gclk));
	jdff dff_B_ZBXRjinY4_1(.din(w_dff_B_8EEViAgp5_1),.dout(w_dff_B_ZBXRjinY4_1),.clk(gclk));
	jdff dff_B_vpM9D0Nn1_1(.din(n220),.dout(w_dff_B_vpM9D0Nn1_1),.clk(gclk));
	jdff dff_B_7gp16oMc7_1(.din(w_dff_B_vpM9D0Nn1_1),.dout(w_dff_B_7gp16oMc7_1),.clk(gclk));
	jdff dff_B_Rj3ZIoqq0_1(.din(n221),.dout(w_dff_B_Rj3ZIoqq0_1),.clk(gclk));
	jdff dff_B_CttyHu5X5_1(.din(w_dff_B_Rj3ZIoqq0_1),.dout(w_dff_B_CttyHu5X5_1),.clk(gclk));
	jdff dff_B_eqnvoQfK6_1(.din(w_dff_B_CttyHu5X5_1),.dout(w_dff_B_eqnvoQfK6_1),.clk(gclk));
	jdff dff_B_1zCmO3lA2_1(.din(w_dff_B_eqnvoQfK6_1),.dout(w_dff_B_1zCmO3lA2_1),.clk(gclk));
	jdff dff_B_mGP2rv5o3_1(.din(w_dff_B_1zCmO3lA2_1),.dout(w_dff_B_mGP2rv5o3_1),.clk(gclk));
	jdff dff_B_FL9O8gPR8_1(.din(w_dff_B_mGP2rv5o3_1),.dout(w_dff_B_FL9O8gPR8_1),.clk(gclk));
	jdff dff_B_df95UIfR2_0(.din(n225),.dout(w_dff_B_df95UIfR2_0),.clk(gclk));
	jdff dff_B_XuzvRLPn3_0(.din(w_dff_B_df95UIfR2_0),.dout(w_dff_B_XuzvRLPn3_0),.clk(gclk));
	jdff dff_B_stLYjEdZ3_0(.din(w_dff_B_XuzvRLPn3_0),.dout(w_dff_B_stLYjEdZ3_0),.clk(gclk));
	jdff dff_B_3zVDPLk09_0(.din(w_dff_B_stLYjEdZ3_0),.dout(w_dff_B_3zVDPLk09_0),.clk(gclk));
	jdff dff_B_QzWvvx3q0_0(.din(w_dff_B_3zVDPLk09_0),.dout(w_dff_B_QzWvvx3q0_0),.clk(gclk));
	jdff dff_B_4lmlfvqX7_0(.din(w_dff_B_QzWvvx3q0_0),.dout(w_dff_B_4lmlfvqX7_0),.clk(gclk));
	jdff dff_B_UUZuZzHr4_0(.din(w_dff_B_4lmlfvqX7_0),.dout(w_dff_B_UUZuZzHr4_0),.clk(gclk));
	jdff dff_B_cmR8wiw80_0(.din(w_dff_B_UUZuZzHr4_0),.dout(w_dff_B_cmR8wiw80_0),.clk(gclk));
	jdff dff_A_11az7EPc0_1(.dout(w_G246gat_3[1]),.din(w_dff_A_11az7EPc0_1),.clk(gclk));
	jdff dff_A_J0on60g63_1(.dout(w_G237gat_3[1]),.din(w_dff_A_J0on60g63_1),.clk(gclk));
	jdff dff_A_4XAIkLJo8_1(.dout(w_n219_0[1]),.din(w_dff_A_4XAIkLJo8_1),.clk(gclk));
	jdff dff_A_xTzFV7qt0_1(.dout(w_dff_A_4XAIkLJo8_1),.din(w_dff_A_xTzFV7qt0_1),.clk(gclk));
	jdff dff_A_uGzJbVJk5_1(.dout(w_dff_A_xTzFV7qt0_1),.din(w_dff_A_uGzJbVJk5_1),.clk(gclk));
	jdff dff_A_rx4gjPAv9_1(.dout(w_dff_A_uGzJbVJk5_1),.din(w_dff_A_rx4gjPAv9_1),.clk(gclk));
	jdff dff_A_aAbtjdr84_1(.dout(w_dff_A_rx4gjPAv9_1),.din(w_dff_A_aAbtjdr84_1),.clk(gclk));
	jdff dff_A_ttwvEnVp9_1(.dout(w_dff_A_aAbtjdr84_1),.din(w_dff_A_ttwvEnVp9_1),.clk(gclk));
	jdff dff_A_WgetRk2g0_1(.dout(w_dff_A_ttwvEnVp9_1),.din(w_dff_A_WgetRk2g0_1),.clk(gclk));
	jdff dff_A_y8Eld7Ju7_1(.dout(w_G228gat_3[1]),.din(w_dff_A_y8Eld7Ju7_1),.clk(gclk));
	jdff dff_B_XY0MeAbk0_1(.din(n278),.dout(w_dff_B_XY0MeAbk0_1),.clk(gclk));
	jdff dff_B_c9O0j8eg6_1(.din(w_dff_B_XY0MeAbk0_1),.dout(w_dff_B_c9O0j8eg6_1),.clk(gclk));
	jdff dff_B_NwbbVXk69_1(.din(w_dff_B_c9O0j8eg6_1),.dout(w_dff_B_NwbbVXk69_1),.clk(gclk));
	jdff dff_B_H0Cw9gyn7_1(.din(w_dff_B_NwbbVXk69_1),.dout(w_dff_B_H0Cw9gyn7_1),.clk(gclk));
	jdff dff_B_wJjuf0yv8_1(.din(w_dff_B_H0Cw9gyn7_1),.dout(w_dff_B_wJjuf0yv8_1),.clk(gclk));
	jdff dff_B_pzxGdjD11_1(.din(n279),.dout(w_dff_B_pzxGdjD11_1),.clk(gclk));
	jdff dff_B_mOBbxzxg0_0(.din(n280),.dout(w_dff_B_mOBbxzxg0_0),.clk(gclk));
	jdff dff_B_05R5fqsH1_0(.din(w_dff_B_mOBbxzxg0_0),.dout(w_dff_B_05R5fqsH1_0),.clk(gclk));
	jdff dff_B_1IxAMKWI8_0(.din(w_dff_B_05R5fqsH1_0),.dout(w_dff_B_1IxAMKWI8_0),.clk(gclk));
	jdff dff_B_OdaqrOtz5_0(.din(w_dff_B_1IxAMKWI8_0),.dout(w_dff_B_OdaqrOtz5_0),.clk(gclk));
	jdff dff_A_RUXZGA5t8_0(.dout(w_G219gat_3[0]),.din(w_dff_A_RUXZGA5t8_0),.clk(gclk));
	jdff dff_A_8ptVZXIC5_0(.dout(w_dff_A_RUXZGA5t8_0),.din(w_dff_A_8ptVZXIC5_0),.clk(gclk));
	jdff dff_A_gaBE8EBh3_0(.dout(w_dff_A_8ptVZXIC5_0),.din(w_dff_A_gaBE8EBh3_0),.clk(gclk));
	jdff dff_A_0EQwirwp1_1(.dout(w_G219gat_3[1]),.din(w_dff_A_0EQwirwp1_1),.clk(gclk));
	jdff dff_A_tfA2nGQm0_1(.dout(w_dff_A_0EQwirwp1_1),.din(w_dff_A_tfA2nGQm0_1),.clk(gclk));
	jdff dff_A_2p3IiiEe1_1(.dout(w_dff_A_tfA2nGQm0_1),.din(w_dff_A_2p3IiiEe1_1),.clk(gclk));
	jdff dff_A_6phzMpUm2_1(.dout(w_dff_A_2p3IiiEe1_1),.din(w_dff_A_6phzMpUm2_1),.clk(gclk));
	jdff dff_A_Vs6wtd3O9_1(.dout(w_dff_A_6phzMpUm2_1),.din(w_dff_A_Vs6wtd3O9_1),.clk(gclk));
	jdff dff_B_7Jcnxepb2_1(.din(n268),.dout(w_dff_B_7Jcnxepb2_1),.clk(gclk));
	jdff dff_B_wMUZqVJX6_0(.din(n276),.dout(w_dff_B_wMUZqVJX6_0),.clk(gclk));
	jdff dff_B_6yVM5fKy6_0(.din(w_dff_B_wMUZqVJX6_0),.dout(w_dff_B_6yVM5fKy6_0),.clk(gclk));
	jdff dff_B_IhgK8L7H9_0(.din(w_dff_B_6yVM5fKy6_0),.dout(w_dff_B_IhgK8L7H9_0),.clk(gclk));
	jdff dff_B_gyWb3mQN5_0(.din(w_dff_B_IhgK8L7H9_0),.dout(w_dff_B_gyWb3mQN5_0),.clk(gclk));
	jdff dff_B_qKue6jvL7_1(.din(n269),.dout(w_dff_B_qKue6jvL7_1),.clk(gclk));
	jdff dff_B_JyDi3Oy99_1(.din(w_dff_B_qKue6jvL7_1),.dout(w_dff_B_JyDi3Oy99_1),.clk(gclk));
	jdff dff_B_MpRywvLK8_1(.din(w_dff_B_JyDi3Oy99_1),.dout(w_dff_B_MpRywvLK8_1),.clk(gclk));
	jdff dff_B_WsMdoAZy9_1(.din(w_dff_B_MpRywvLK8_1),.dout(w_dff_B_WsMdoAZy9_1),.clk(gclk));
	jdff dff_B_RATKL9N39_1(.din(w_dff_B_WsMdoAZy9_1),.dout(w_dff_B_RATKL9N39_1),.clk(gclk));
	jdff dff_B_kw6UwvrJ0_1(.din(w_dff_B_RATKL9N39_1),.dout(w_dff_B_kw6UwvrJ0_1),.clk(gclk));
	jdff dff_B_ETZZTpSk0_1(.din(w_dff_B_kw6UwvrJ0_1),.dout(w_dff_B_ETZZTpSk0_1),.clk(gclk));
	jdff dff_B_ogepBvZs6_1(.din(w_dff_B_ETZZTpSk0_1),.dout(w_dff_B_ogepBvZs6_1),.clk(gclk));
	jdff dff_B_HrlsXUcx3_0(.din(n271),.dout(w_dff_B_HrlsXUcx3_0),.clk(gclk));
	jdff dff_B_cuXdf9w35_0(.din(w_dff_B_HrlsXUcx3_0),.dout(w_dff_B_cuXdf9w35_0),.clk(gclk));
	jdff dff_B_n54Jdcop5_0(.din(w_dff_B_cuXdf9w35_0),.dout(w_dff_B_n54Jdcop5_0),.clk(gclk));
	jdff dff_B_ykWxcPfT8_0(.din(w_dff_B_n54Jdcop5_0),.dout(w_dff_B_ykWxcPfT8_0),.clk(gclk));
	jdff dff_B_0I3M9pmG9_0(.din(w_dff_B_ykWxcPfT8_0),.dout(w_dff_B_0I3M9pmG9_0),.clk(gclk));
	jdff dff_B_LiJqcHEa1_0(.din(w_dff_B_0I3M9pmG9_0),.dout(w_dff_B_LiJqcHEa1_0),.clk(gclk));
	jdff dff_A_m5dLRo3E2_1(.dout(w_n267_0[1]),.din(w_dff_A_m5dLRo3E2_1),.clk(gclk));
	jdff dff_A_Z6oCp6y41_1(.dout(w_dff_A_m5dLRo3E2_1),.din(w_dff_A_Z6oCp6y41_1),.clk(gclk));
	jdff dff_A_22A5OXr00_1(.dout(w_dff_A_Z6oCp6y41_1),.din(w_dff_A_22A5OXr00_1),.clk(gclk));
	jdff dff_A_Rxc8T17A4_1(.dout(w_dff_A_22A5OXr00_1),.din(w_dff_A_Rxc8T17A4_1),.clk(gclk));
	jdff dff_A_5b2xuoH16_1(.dout(w_dff_A_Rxc8T17A4_1),.din(w_dff_A_5b2xuoH16_1),.clk(gclk));
	jdff dff_B_uKBg6Jm14_1(.din(n296),.dout(w_dff_B_uKBg6Jm14_1),.clk(gclk));
	jdff dff_B_2C1W7kJe2_1(.din(w_dff_B_uKBg6Jm14_1),.dout(w_dff_B_2C1W7kJe2_1),.clk(gclk));
	jdff dff_B_uX9nyNKO7_1(.din(w_dff_B_2C1W7kJe2_1),.dout(w_dff_B_uX9nyNKO7_1),.clk(gclk));
	jdff dff_B_FAex2s4q4_1(.din(n297),.dout(w_dff_B_FAex2s4q4_1),.clk(gclk));
	jdff dff_B_XxtknBJ05_0(.din(n298),.dout(w_dff_B_XxtknBJ05_0),.clk(gclk));
	jdff dff_B_ENeW9ryo0_0(.din(w_dff_B_XxtknBJ05_0),.dout(w_dff_B_ENeW9ryo0_0),.clk(gclk));
	jdff dff_B_kP6EvrmH0_1(.din(n286),.dout(w_dff_B_kP6EvrmH0_1),.clk(gclk));
	jdff dff_B_8LqnAwx22_0(.din(n294),.dout(w_dff_B_8LqnAwx22_0),.clk(gclk));
	jdff dff_B_GA6yjg4Y7_0(.din(w_dff_B_8LqnAwx22_0),.dout(w_dff_B_GA6yjg4Y7_0),.clk(gclk));
	jdff dff_B_zNGHe30A7_0(.din(w_dff_B_GA6yjg4Y7_0),.dout(w_dff_B_zNGHe30A7_0),.clk(gclk));
	jdff dff_B_ebZatS749_0(.din(w_dff_B_zNGHe30A7_0),.dout(w_dff_B_ebZatS749_0),.clk(gclk));
	jdff dff_B_ol4EIhmR1_1(.din(n287),.dout(w_dff_B_ol4EIhmR1_1),.clk(gclk));
	jdff dff_B_9kS0Tl0Z8_1(.din(w_dff_B_ol4EIhmR1_1),.dout(w_dff_B_9kS0Tl0Z8_1),.clk(gclk));
	jdff dff_B_V2uSvaJJ9_1(.din(w_dff_B_9kS0Tl0Z8_1),.dout(w_dff_B_V2uSvaJJ9_1),.clk(gclk));
	jdff dff_B_JNic7gWJ7_1(.din(w_dff_B_V2uSvaJJ9_1),.dout(w_dff_B_JNic7gWJ7_1),.clk(gclk));
	jdff dff_B_unMdeZK19_1(.din(w_dff_B_JNic7gWJ7_1),.dout(w_dff_B_unMdeZK19_1),.clk(gclk));
	jdff dff_B_M3nn9zj39_1(.din(w_dff_B_unMdeZK19_1),.dout(w_dff_B_M3nn9zj39_1),.clk(gclk));
	jdff dff_B_ZKiGkW802_1(.din(w_dff_B_M3nn9zj39_1),.dout(w_dff_B_ZKiGkW802_1),.clk(gclk));
	jdff dff_B_AjMpcyz35_1(.din(w_dff_B_ZKiGkW802_1),.dout(w_dff_B_AjMpcyz35_1),.clk(gclk));
	jdff dff_B_khiGMJkC6_0(.din(n289),.dout(w_dff_B_khiGMJkC6_0),.clk(gclk));
	jdff dff_B_cTdvZy4r8_0(.din(w_dff_B_khiGMJkC6_0),.dout(w_dff_B_cTdvZy4r8_0),.clk(gclk));
	jdff dff_B_WCKlEtiR0_0(.din(w_dff_B_cTdvZy4r8_0),.dout(w_dff_B_WCKlEtiR0_0),.clk(gclk));
	jdff dff_B_2a5z1Xjg8_0(.din(w_dff_B_WCKlEtiR0_0),.dout(w_dff_B_2a5z1Xjg8_0),.clk(gclk));
	jdff dff_B_n8OiMxVB2_0(.din(w_dff_B_2a5z1Xjg8_0),.dout(w_dff_B_n8OiMxVB2_0),.clk(gclk));
	jdff dff_B_mC5ZY7pu3_0(.din(w_dff_B_n8OiMxVB2_0),.dout(w_dff_B_mC5ZY7pu3_0),.clk(gclk));
	jdff dff_A_EG9VRG8W6_1(.dout(w_n285_0[1]),.din(w_dff_A_EG9VRG8W6_1),.clk(gclk));
	jdff dff_A_TDoDTVbA9_1(.dout(w_dff_A_EG9VRG8W6_1),.din(w_dff_A_TDoDTVbA9_1),.clk(gclk));
	jdff dff_A_pkqm1NpZ6_1(.dout(w_dff_A_TDoDTVbA9_1),.din(w_dff_A_pkqm1NpZ6_1),.clk(gclk));
	jdff dff_B_fQmRPZON8_1(.din(n312),.dout(w_dff_B_fQmRPZON8_1),.clk(gclk));
	jdff dff_B_T2BT045J4_1(.din(w_dff_B_fQmRPZON8_1),.dout(w_dff_B_T2BT045J4_1),.clk(gclk));
	jdff dff_B_Vjnz68aJ2_1(.din(w_dff_B_T2BT045J4_1),.dout(w_dff_B_Vjnz68aJ2_1),.clk(gclk));
	jdff dff_B_HHKzXRgK4_1(.din(w_dff_B_Vjnz68aJ2_1),.dout(w_dff_B_HHKzXRgK4_1),.clk(gclk));
	jdff dff_B_PKTNXSdz9_1(.din(w_dff_B_HHKzXRgK4_1),.dout(w_dff_B_PKTNXSdz9_1),.clk(gclk));
	jdff dff_B_1fe2UGLo9_1(.din(w_dff_B_PKTNXSdz9_1),.dout(w_dff_B_1fe2UGLo9_1),.clk(gclk));
	jdff dff_B_uFzmVCRF6_1(.din(w_dff_B_1fe2UGLo9_1),.dout(w_dff_B_uFzmVCRF6_1),.clk(gclk));
	jdff dff_B_oqSPIjM86_1(.din(w_dff_B_uFzmVCRF6_1),.dout(w_dff_B_oqSPIjM86_1),.clk(gclk));
	jdff dff_B_aGB5ctIR2_1(.din(w_dff_B_oqSPIjM86_1),.dout(w_dff_B_aGB5ctIR2_1),.clk(gclk));
	jdff dff_B_zCKZstdA2_1(.din(w_dff_B_aGB5ctIR2_1),.dout(w_dff_B_zCKZstdA2_1),.clk(gclk));
	jdff dff_B_EPFRqy7F8_1(.din(w_dff_B_zCKZstdA2_1),.dout(w_dff_B_EPFRqy7F8_1),.clk(gclk));
	jdff dff_B_4i9kXI6q3_1(.din(w_dff_B_EPFRqy7F8_1),.dout(w_dff_B_4i9kXI6q3_1),.clk(gclk));
	jdff dff_B_SAkTrJKB8_1(.din(w_dff_B_4i9kXI6q3_1),.dout(w_dff_B_SAkTrJKB8_1),.clk(gclk));
	jdff dff_B_9yKBK2lv1_1(.din(w_dff_B_SAkTrJKB8_1),.dout(w_dff_B_9yKBK2lv1_1),.clk(gclk));
	jdff dff_B_jQQigADs9_1(.din(w_dff_B_9yKBK2lv1_1),.dout(w_dff_B_jQQigADs9_1),.clk(gclk));
	jdff dff_B_1ghF9F5c0_1(.din(n313),.dout(w_dff_B_1ghF9F5c0_1),.clk(gclk));
	jdff dff_B_fgtMIk5n0_1(.din(w_dff_B_1ghF9F5c0_1),.dout(w_dff_B_fgtMIk5n0_1),.clk(gclk));
	jdff dff_B_4xuD6Oz99_1(.din(w_dff_B_fgtMIk5n0_1),.dout(w_dff_B_4xuD6Oz99_1),.clk(gclk));
	jdff dff_B_Sl7Zzit09_1(.din(w_dff_B_4xuD6Oz99_1),.dout(w_dff_B_Sl7Zzit09_1),.clk(gclk));
	jdff dff_B_knfWUuIT3_1(.din(w_dff_B_Sl7Zzit09_1),.dout(w_dff_B_knfWUuIT3_1),.clk(gclk));
	jdff dff_B_JYzYanh11_1(.din(w_dff_B_knfWUuIT3_1),.dout(w_dff_B_JYzYanh11_1),.clk(gclk));
	jdff dff_B_jn2LKAOE3_1(.din(w_dff_B_JYzYanh11_1),.dout(w_dff_B_jn2LKAOE3_1),.clk(gclk));
	jdff dff_B_Il4C0t5C1_1(.din(w_dff_B_jn2LKAOE3_1),.dout(w_dff_B_Il4C0t5C1_1),.clk(gclk));
	jdff dff_B_6ZBnnazU6_1(.din(w_dff_B_Il4C0t5C1_1),.dout(w_dff_B_6ZBnnazU6_1),.clk(gclk));
	jdff dff_B_6zpwPUYv8_1(.din(w_dff_B_6ZBnnazU6_1),.dout(w_dff_B_6zpwPUYv8_1),.clk(gclk));
	jdff dff_B_0sXp9gMc4_1(.din(w_dff_B_6zpwPUYv8_1),.dout(w_dff_B_0sXp9gMc4_1),.clk(gclk));
	jdff dff_B_FAoYoW3d1_1(.din(w_dff_B_0sXp9gMc4_1),.dout(w_dff_B_FAoYoW3d1_1),.clk(gclk));
	jdff dff_B_b5qaLfel0_1(.din(w_dff_B_FAoYoW3d1_1),.dout(w_dff_B_b5qaLfel0_1),.clk(gclk));
	jdff dff_B_uRMRSEKs8_1(.din(w_dff_B_b5qaLfel0_1),.dout(w_dff_B_uRMRSEKs8_1),.clk(gclk));
	jdff dff_B_BqlEClB84_1(.din(n358),.dout(w_dff_B_BqlEClB84_1),.clk(gclk));
	jdff dff_B_1Tv7GAvm9_1(.din(w_dff_B_BqlEClB84_1),.dout(w_dff_B_1Tv7GAvm9_1),.clk(gclk));
	jdff dff_B_ve0nPmlW8_0(.din(n371),.dout(w_dff_B_ve0nPmlW8_0),.clk(gclk));
	jdff dff_B_tgWSbjKB2_0(.din(w_dff_B_ve0nPmlW8_0),.dout(w_dff_B_tgWSbjKB2_0),.clk(gclk));
	jdff dff_B_Jq33RNee0_0(.din(w_dff_B_tgWSbjKB2_0),.dout(w_dff_B_Jq33RNee0_0),.clk(gclk));
	jdff dff_B_uERczs310_0(.din(w_dff_B_Jq33RNee0_0),.dout(w_dff_B_uERczs310_0),.clk(gclk));
	jdff dff_B_9mc8XRc13_0(.din(w_dff_B_uERczs310_0),.dout(w_dff_B_9mc8XRc13_0),.clk(gclk));
	jdff dff_B_8VlGQYTN5_0(.din(w_dff_B_9mc8XRc13_0),.dout(w_dff_B_8VlGQYTN5_0),.clk(gclk));
	jdff dff_B_1qVZahQd5_0(.din(w_dff_B_8VlGQYTN5_0),.dout(w_dff_B_1qVZahQd5_0),.clk(gclk));
	jdff dff_B_cT7p5vUi3_0(.din(w_dff_B_1qVZahQd5_0),.dout(w_dff_B_cT7p5vUi3_0),.clk(gclk));
	jdff dff_B_kLpPMk8B5_0(.din(w_dff_B_cT7p5vUi3_0),.dout(w_dff_B_kLpPMk8B5_0),.clk(gclk));
	jdff dff_B_AENKSLvw6_0(.din(n369),.dout(w_dff_B_AENKSLvw6_0),.clk(gclk));
	jdff dff_B_9BGn4cHj0_0(.din(w_dff_B_AENKSLvw6_0),.dout(w_dff_B_9BGn4cHj0_0),.clk(gclk));
	jdff dff_B_oN1vl44e4_0(.din(w_dff_B_9BGn4cHj0_0),.dout(w_dff_B_oN1vl44e4_0),.clk(gclk));
	jdff dff_B_Bs7DS11W5_0(.din(w_dff_B_oN1vl44e4_0),.dout(w_dff_B_Bs7DS11W5_0),.clk(gclk));
	jdff dff_A_Cu0EyjeM0_0(.dout(w_G228gat_2[0]),.din(w_dff_A_Cu0EyjeM0_0),.clk(gclk));
	jdff dff_A_BJqwCyrt5_0(.dout(w_dff_A_Cu0EyjeM0_0),.din(w_dff_A_BJqwCyrt5_0),.clk(gclk));
	jdff dff_A_lfm1JmaT8_0(.dout(w_dff_A_BJqwCyrt5_0),.din(w_dff_A_lfm1JmaT8_0),.clk(gclk));
	jdff dff_A_k31Yre1t9_0(.dout(w_dff_A_lfm1JmaT8_0),.din(w_dff_A_k31Yre1t9_0),.clk(gclk));
	jdff dff_A_EBaxjGJw3_0(.dout(w_dff_A_k31Yre1t9_0),.din(w_dff_A_EBaxjGJw3_0),.clk(gclk));
	jdff dff_A_UFCUDzQm4_0(.dout(w_dff_A_EBaxjGJw3_0),.din(w_dff_A_UFCUDzQm4_0),.clk(gclk));
	jdff dff_A_fz5qyEiG5_0(.dout(w_dff_A_UFCUDzQm4_0),.din(w_dff_A_fz5qyEiG5_0),.clk(gclk));
	jdff dff_A_eG6iFr2p8_0(.dout(w_dff_A_fz5qyEiG5_0),.din(w_dff_A_eG6iFr2p8_0),.clk(gclk));
	jdff dff_A_cwaJ42z55_0(.dout(w_dff_A_eG6iFr2p8_0),.din(w_dff_A_cwaJ42z55_0),.clk(gclk));
	jdff dff_A_qHxwdpt16_0(.dout(w_dff_A_cwaJ42z55_0),.din(w_dff_A_qHxwdpt16_0),.clk(gclk));
	jdff dff_B_zqoxhkzJ3_1(.din(n356),.dout(w_dff_B_zqoxhkzJ3_1),.clk(gclk));
	jdff dff_B_yG6Jm40g3_1(.din(w_dff_B_zqoxhkzJ3_1),.dout(w_dff_B_yG6Jm40g3_1),.clk(gclk));
	jdff dff_B_jJJgY1Qs3_1(.din(w_dff_B_yG6Jm40g3_1),.dout(w_dff_B_jJJgY1Qs3_1),.clk(gclk));
	jdff dff_B_95RgYvRz4_1(.din(w_dff_B_jJJgY1Qs3_1),.dout(w_dff_B_95RgYvRz4_1),.clk(gclk));
	jdff dff_B_aHtzEbHB4_1(.din(w_dff_B_95RgYvRz4_1),.dout(w_dff_B_aHtzEbHB4_1),.clk(gclk));
	jdff dff_B_PFNWSu7G1_1(.din(w_dff_B_aHtzEbHB4_1),.dout(w_dff_B_PFNWSu7G1_1),.clk(gclk));
	jdff dff_B_Yykectua0_1(.din(w_dff_B_PFNWSu7G1_1),.dout(w_dff_B_Yykectua0_1),.clk(gclk));
	jdff dff_B_BLIkJKXs8_1(.din(w_dff_B_Yykectua0_1),.dout(w_dff_B_BLIkJKXs8_1),.clk(gclk));
	jdff dff_A_UPjMzRRM7_0(.dout(w_G219gat_2[0]),.din(w_dff_A_UPjMzRRM7_0),.clk(gclk));
	jdff dff_A_stdpmX2N9_0(.dout(w_dff_A_UPjMzRRM7_0),.din(w_dff_A_stdpmX2N9_0),.clk(gclk));
	jdff dff_A_iPzLhe5Q3_0(.dout(w_dff_A_stdpmX2N9_0),.din(w_dff_A_iPzLhe5Q3_0),.clk(gclk));
	jdff dff_A_xM7THKaw2_0(.dout(w_dff_A_iPzLhe5Q3_0),.din(w_dff_A_xM7THKaw2_0),.clk(gclk));
	jdff dff_A_7eFcm9HF7_0(.dout(w_dff_A_xM7THKaw2_0),.din(w_dff_A_7eFcm9HF7_0),.clk(gclk));
	jdff dff_A_of1xeFnv0_1(.dout(w_G219gat_2[1]),.din(w_dff_A_of1xeFnv0_1),.clk(gclk));
	jdff dff_A_2zxuqYs59_1(.dout(w_dff_A_of1xeFnv0_1),.din(w_dff_A_2zxuqYs59_1),.clk(gclk));
	jdff dff_A_ywjDpfpj5_1(.dout(w_dff_A_2zxuqYs59_1),.din(w_dff_A_ywjDpfpj5_1),.clk(gclk));
	jdff dff_A_jnnl83Gv3_1(.dout(w_dff_A_ywjDpfpj5_1),.din(w_dff_A_jnnl83Gv3_1),.clk(gclk));
	jdff dff_A_YnXncBJ56_1(.dout(w_dff_A_jnnl83Gv3_1),.din(w_dff_A_YnXncBJ56_1),.clk(gclk));
	jdff dff_A_2GrLUlwC4_0(.dout(w_n355_0[0]),.din(w_dff_A_2GrLUlwC4_0),.clk(gclk));
	jdff dff_A_Fmz9ih9H1_0(.dout(w_dff_A_2GrLUlwC4_0),.din(w_dff_A_Fmz9ih9H1_0),.clk(gclk));
	jdff dff_A_B01JyBuR4_0(.dout(w_dff_A_Fmz9ih9H1_0),.din(w_dff_A_B01JyBuR4_0),.clk(gclk));
	jdff dff_A_Yb8ZA5p08_0(.dout(w_dff_A_B01JyBuR4_0),.din(w_dff_A_Yb8ZA5p08_0),.clk(gclk));
	jdff dff_A_pxZ0xUpf1_0(.dout(w_dff_A_Yb8ZA5p08_0),.din(w_dff_A_pxZ0xUpf1_0),.clk(gclk));
	jdff dff_A_C7Mu9xf33_0(.dout(w_dff_A_pxZ0xUpf1_0),.din(w_dff_A_C7Mu9xf33_0),.clk(gclk));
	jdff dff_A_OKZjSb8D3_0(.dout(w_dff_A_C7Mu9xf33_0),.din(w_dff_A_OKZjSb8D3_0),.clk(gclk));
	jdff dff_A_cbvdV27n2_0(.dout(w_dff_A_OKZjSb8D3_0),.din(w_dff_A_cbvdV27n2_0),.clk(gclk));
	jdff dff_A_0Dvpp9520_0(.dout(w_dff_A_cbvdV27n2_0),.din(w_dff_A_0Dvpp9520_0),.clk(gclk));
	jdff dff_A_fs0rZYQO3_0(.dout(w_dff_A_0Dvpp9520_0),.din(w_dff_A_fs0rZYQO3_0),.clk(gclk));
	jdff dff_B_BRCBa8Gm3_1(.din(n383),.dout(w_dff_B_BRCBa8Gm3_1),.clk(gclk));
	jdff dff_B_dE3nxvlr2_1(.din(w_dff_B_BRCBa8Gm3_1),.dout(w_dff_B_dE3nxvlr2_1),.clk(gclk));
	jdff dff_B_JhWLMC056_1(.din(w_dff_B_dE3nxvlr2_1),.dout(w_dff_B_JhWLMC056_1),.clk(gclk));
	jdff dff_B_JWUBqizD4_1(.din(w_dff_B_JhWLMC056_1),.dout(w_dff_B_JWUBqizD4_1),.clk(gclk));
	jdff dff_B_hXbeFuTr8_1(.din(w_dff_B_JWUBqizD4_1),.dout(w_dff_B_hXbeFuTr8_1),.clk(gclk));
	jdff dff_B_w0avvtP58_1(.din(w_dff_B_hXbeFuTr8_1),.dout(w_dff_B_w0avvtP58_1),.clk(gclk));
	jdff dff_B_lAvnDYCV9_1(.din(w_dff_B_w0avvtP58_1),.dout(w_dff_B_lAvnDYCV9_1),.clk(gclk));
	jdff dff_B_CCaDncC33_1(.din(w_dff_B_lAvnDYCV9_1),.dout(w_dff_B_CCaDncC33_1),.clk(gclk));
	jdff dff_B_nRcRGbWL5_1(.din(w_dff_B_CCaDncC33_1),.dout(w_dff_B_nRcRGbWL5_1),.clk(gclk));
	jdff dff_B_kSHNl5BN0_1(.din(w_dff_B_nRcRGbWL5_1),.dout(w_dff_B_kSHNl5BN0_1),.clk(gclk));
	jdff dff_B_udxFi3po4_1(.din(w_dff_B_kSHNl5BN0_1),.dout(w_dff_B_udxFi3po4_1),.clk(gclk));
	jdff dff_B_cgovtZgz8_1(.din(w_dff_B_udxFi3po4_1),.dout(w_dff_B_cgovtZgz8_1),.clk(gclk));
	jdff dff_B_cwtaCgur6_1(.din(w_dff_B_cgovtZgz8_1),.dout(w_dff_B_cwtaCgur6_1),.clk(gclk));
	jdff dff_B_j1jZDTRW8_1(.din(n384),.dout(w_dff_B_j1jZDTRW8_1),.clk(gclk));
	jdff dff_B_tl4V774Y2_0(.din(n396),.dout(w_dff_B_tl4V774Y2_0),.clk(gclk));
	jdff dff_B_9qAjwCpN3_0(.din(w_dff_B_tl4V774Y2_0),.dout(w_dff_B_9qAjwCpN3_0),.clk(gclk));
	jdff dff_B_GgSowWm09_0(.din(w_dff_B_9qAjwCpN3_0),.dout(w_dff_B_GgSowWm09_0),.clk(gclk));
	jdff dff_B_u4XwBN3V3_0(.din(w_dff_B_GgSowWm09_0),.dout(w_dff_B_u4XwBN3V3_0),.clk(gclk));
	jdff dff_B_Qqh7uzFs6_0(.din(w_dff_B_u4XwBN3V3_0),.dout(w_dff_B_Qqh7uzFs6_0),.clk(gclk));
	jdff dff_B_mbSjwtzG9_0(.din(w_dff_B_Qqh7uzFs6_0),.dout(w_dff_B_mbSjwtzG9_0),.clk(gclk));
	jdff dff_B_Wei9aZmN0_0(.din(w_dff_B_mbSjwtzG9_0),.dout(w_dff_B_Wei9aZmN0_0),.clk(gclk));
	jdff dff_B_QgysHtIL2_0(.din(w_dff_B_Wei9aZmN0_0),.dout(w_dff_B_QgysHtIL2_0),.clk(gclk));
	jdff dff_B_Zd8bgh8O6_0(.din(w_dff_B_QgysHtIL2_0),.dout(w_dff_B_Zd8bgh8O6_0),.clk(gclk));
	jdff dff_B_mHafxW2Q4_0(.din(w_dff_B_Zd8bgh8O6_0),.dout(w_dff_B_mHafxW2Q4_0),.clk(gclk));
	jdff dff_B_CX3IjYz83_0(.din(w_dff_B_mHafxW2Q4_0),.dout(w_dff_B_CX3IjYz83_0),.clk(gclk));
	jdff dff_B_iVt3tfbj1_0(.din(w_dff_B_CX3IjYz83_0),.dout(w_dff_B_iVt3tfbj1_0),.clk(gclk));
	jdff dff_B_p8dNjgNM2_0(.din(w_dff_B_iVt3tfbj1_0),.dout(w_dff_B_p8dNjgNM2_0),.clk(gclk));
	jdff dff_B_DJB3hdRk1_1(.din(n385),.dout(w_dff_B_DJB3hdRk1_1),.clk(gclk));
	jdff dff_B_FJqerLoq1_1(.din(w_dff_B_DJB3hdRk1_1),.dout(w_dff_B_FJqerLoq1_1),.clk(gclk));
	jdff dff_B_Wq865ogK6_1(.din(w_dff_B_FJqerLoq1_1),.dout(w_dff_B_Wq865ogK6_1),.clk(gclk));
	jdff dff_B_LewQBoAp5_1(.din(w_dff_B_Wq865ogK6_1),.dout(w_dff_B_LewQBoAp5_1),.clk(gclk));
	jdff dff_B_NeTiRv242_1(.din(w_dff_B_LewQBoAp5_1),.dout(w_dff_B_NeTiRv242_1),.clk(gclk));
	jdff dff_B_spsy8lYm5_1(.din(w_dff_B_NeTiRv242_1),.dout(w_dff_B_spsy8lYm5_1),.clk(gclk));
	jdff dff_B_pPASdmkn0_1(.din(w_dff_B_spsy8lYm5_1),.dout(w_dff_B_pPASdmkn0_1),.clk(gclk));
	jdff dff_B_Q5hMidMZ8_1(.din(w_dff_B_pPASdmkn0_1),.dout(w_dff_B_Q5hMidMZ8_1),.clk(gclk));
	jdff dff_B_6l3PGBbg8_1(.din(w_dff_B_Q5hMidMZ8_1),.dout(w_dff_B_6l3PGBbg8_1),.clk(gclk));
	jdff dff_B_ntz2DTLr8_1(.din(w_dff_B_6l3PGBbg8_1),.dout(w_dff_B_ntz2DTLr8_1),.clk(gclk));
	jdff dff_B_gyQzON464_1(.din(w_dff_B_ntz2DTLr8_1),.dout(w_dff_B_gyQzON464_1),.clk(gclk));
	jdff dff_B_uC21U4j09_1(.din(w_dff_B_gyQzON464_1),.dout(w_dff_B_uC21U4j09_1),.clk(gclk));
	jdff dff_B_1zGjvSz99_1(.din(n386),.dout(w_dff_B_1zGjvSz99_1),.clk(gclk));
	jdff dff_B_Odu7rsgL8_1(.din(w_dff_B_1zGjvSz99_1),.dout(w_dff_B_Odu7rsgL8_1),.clk(gclk));
	jdff dff_B_CeDgb4uI5_1(.din(w_dff_B_Odu7rsgL8_1),.dout(w_dff_B_CeDgb4uI5_1),.clk(gclk));
	jdff dff_B_hLhf6NjV9_1(.din(w_dff_B_CeDgb4uI5_1),.dout(w_dff_B_hLhf6NjV9_1),.clk(gclk));
	jdff dff_B_0gP8RICC7_1(.din(w_dff_B_hLhf6NjV9_1),.dout(w_dff_B_0gP8RICC7_1),.clk(gclk));
	jdff dff_B_CDBMehEJ7_1(.din(w_dff_B_0gP8RICC7_1),.dout(w_dff_B_CDBMehEJ7_1),.clk(gclk));
	jdff dff_B_K4ubMvt41_1(.din(w_dff_B_CDBMehEJ7_1),.dout(w_dff_B_K4ubMvt41_1),.clk(gclk));
	jdff dff_B_pVGD8yq74_1(.din(w_dff_B_K4ubMvt41_1),.dout(w_dff_B_pVGD8yq74_1),.clk(gclk));
	jdff dff_B_6mcDbINK2_1(.din(w_dff_B_pVGD8yq74_1),.dout(w_dff_B_6mcDbINK2_1),.clk(gclk));
	jdff dff_B_4BmzX0fv0_1(.din(w_dff_B_6mcDbINK2_1),.dout(w_dff_B_4BmzX0fv0_1),.clk(gclk));
	jdff dff_B_kXtpPMaG3_1(.din(w_dff_B_4BmzX0fv0_1),.dout(w_dff_B_kXtpPMaG3_1),.clk(gclk));
	jdff dff_A_6XpegKSm4_1(.dout(w_n321_0[1]),.din(w_dff_A_6XpegKSm4_1),.clk(gclk));
	jdff dff_A_drOnVS6z3_1(.dout(w_dff_A_6XpegKSm4_1),.din(w_dff_A_drOnVS6z3_1),.clk(gclk));
	jdff dff_A_LrXIiMcv6_1(.dout(w_dff_A_drOnVS6z3_1),.din(w_dff_A_LrXIiMcv6_1),.clk(gclk));
	jdff dff_A_yAmbt8ID9_1(.dout(w_dff_A_LrXIiMcv6_1),.din(w_dff_A_yAmbt8ID9_1),.clk(gclk));
	jdff dff_A_0jQ6sryO3_1(.dout(w_dff_A_yAmbt8ID9_1),.din(w_dff_A_0jQ6sryO3_1),.clk(gclk));
	jdff dff_A_o0i22IS56_1(.dout(w_dff_A_0jQ6sryO3_1),.din(w_dff_A_o0i22IS56_1),.clk(gclk));
	jdff dff_A_jv5mWzwL6_1(.dout(w_dff_A_o0i22IS56_1),.din(w_dff_A_jv5mWzwL6_1),.clk(gclk));
	jdff dff_A_ihPpej2Q0_1(.dout(w_dff_A_jv5mWzwL6_1),.din(w_dff_A_ihPpej2Q0_1),.clk(gclk));
	jdff dff_A_7JtItBnh3_1(.dout(w_dff_A_ihPpej2Q0_1),.din(w_dff_A_7JtItBnh3_1),.clk(gclk));
	jdff dff_A_Zm3lozEW9_1(.dout(w_dff_A_7JtItBnh3_1),.din(w_dff_A_Zm3lozEW9_1),.clk(gclk));
	jdff dff_A_3nGvN2zy2_1(.dout(w_dff_A_Zm3lozEW9_1),.din(w_dff_A_3nGvN2zy2_1),.clk(gclk));
	jdff dff_A_BdvaWRgm5_1(.dout(w_dff_A_3nGvN2zy2_1),.din(w_dff_A_BdvaWRgm5_1),.clk(gclk));
	jdff dff_A_drq8MwUV8_1(.dout(w_n320_0[1]),.din(w_dff_A_drq8MwUV8_1),.clk(gclk));
	jdff dff_A_oVQe4ZXh9_1(.dout(w_dff_A_drq8MwUV8_1),.din(w_dff_A_oVQe4ZXh9_1),.clk(gclk));
	jdff dff_A_zTsKiS1O7_1(.dout(w_dff_A_oVQe4ZXh9_1),.din(w_dff_A_zTsKiS1O7_1),.clk(gclk));
	jdff dff_A_2m1P00Ww4_1(.dout(w_dff_A_zTsKiS1O7_1),.din(w_dff_A_2m1P00Ww4_1),.clk(gclk));
	jdff dff_A_nDwfb40U1_1(.dout(w_dff_A_2m1P00Ww4_1),.din(w_dff_A_nDwfb40U1_1),.clk(gclk));
	jdff dff_A_bXrPZwFe6_1(.dout(w_dff_A_nDwfb40U1_1),.din(w_dff_A_bXrPZwFe6_1),.clk(gclk));
	jdff dff_A_MgiaceAj4_1(.dout(w_dff_A_bXrPZwFe6_1),.din(w_dff_A_MgiaceAj4_1),.clk(gclk));
	jdff dff_A_WYotL46y6_1(.dout(w_dff_A_MgiaceAj4_1),.din(w_dff_A_WYotL46y6_1),.clk(gclk));
	jdff dff_A_d2Hob7nh7_1(.dout(w_dff_A_WYotL46y6_1),.din(w_dff_A_d2Hob7nh7_1),.clk(gclk));
	jdff dff_A_4ss6uSeZ6_1(.dout(w_dff_A_d2Hob7nh7_1),.din(w_dff_A_4ss6uSeZ6_1),.clk(gclk));
	jdff dff_A_HHwTvurL0_1(.dout(w_dff_A_4ss6uSeZ6_1),.din(w_dff_A_HHwTvurL0_1),.clk(gclk));
	jdff dff_A_VinsUufh7_1(.dout(w_dff_A_HHwTvurL0_1),.din(w_dff_A_VinsUufh7_1),.clk(gclk));
	jdff dff_A_QPcncT2h7_1(.dout(w_dff_A_VinsUufh7_1),.din(w_dff_A_QPcncT2h7_1),.clk(gclk));
	jdff dff_B_9u6nPr194_1(.din(n376),.dout(w_dff_B_9u6nPr194_1),.clk(gclk));
	jdff dff_B_8D4hzEhG8_0(.din(n381),.dout(w_dff_B_8D4hzEhG8_0),.clk(gclk));
	jdff dff_B_rEqfqAFS6_0(.din(w_dff_B_8D4hzEhG8_0),.dout(w_dff_B_rEqfqAFS6_0),.clk(gclk));
	jdff dff_B_BPh8WUSn4_0(.din(n379),.dout(w_dff_B_BPh8WUSn4_0),.clk(gclk));
	jdff dff_B_H1YqvDCf7_0(.din(w_dff_B_BPh8WUSn4_0),.dout(w_dff_B_H1YqvDCf7_0),.clk(gclk));
	jdff dff_B_EUSsslwO7_0(.din(w_dff_B_H1YqvDCf7_0),.dout(w_dff_B_EUSsslwO7_0),.clk(gclk));
	jdff dff_B_0Al4fIGv0_0(.din(w_dff_B_EUSsslwO7_0),.dout(w_dff_B_0Al4fIGv0_0),.clk(gclk));
	jdff dff_B_aw9470NU3_0(.din(w_dff_B_0Al4fIGv0_0),.dout(w_dff_B_aw9470NU3_0),.clk(gclk));
	jdff dff_B_gZLslMqB6_0(.din(w_dff_B_aw9470NU3_0),.dout(w_dff_B_gZLslMqB6_0),.clk(gclk));
	jdff dff_B_Jz4QAnE20_0(.din(w_dff_B_gZLslMqB6_0),.dout(w_dff_B_Jz4QAnE20_0),.clk(gclk));
	jdff dff_B_CSH8IHe66_0(.din(w_dff_B_Jz4QAnE20_0),.dout(w_dff_B_CSH8IHe66_0),.clk(gclk));
	jdff dff_B_IEinr5W55_0(.din(w_dff_B_CSH8IHe66_0),.dout(w_dff_B_IEinr5W55_0),.clk(gclk));
	jdff dff_B_oBmZdDdv8_0(.din(w_dff_B_IEinr5W55_0),.dout(w_dff_B_oBmZdDdv8_0),.clk(gclk));
	jdff dff_A_VE65fi8p4_1(.dout(w_n377_0[1]),.din(w_dff_A_VE65fi8p4_1),.clk(gclk));
	jdff dff_A_8npv2VtM7_1(.dout(w_dff_A_VE65fi8p4_1),.din(w_dff_A_8npv2VtM7_1),.clk(gclk));
	jdff dff_A_NN5MZ7WJ6_1(.dout(w_dff_A_8npv2VtM7_1),.din(w_dff_A_NN5MZ7WJ6_1),.clk(gclk));
	jdff dff_A_tVDnmAWv5_1(.dout(w_dff_A_NN5MZ7WJ6_1),.din(w_dff_A_tVDnmAWv5_1),.clk(gclk));
	jdff dff_A_I1W6iqkX5_1(.dout(w_dff_A_tVDnmAWv5_1),.din(w_dff_A_I1W6iqkX5_1),.clk(gclk));
	jdff dff_A_GXwDeevO2_1(.dout(w_dff_A_I1W6iqkX5_1),.din(w_dff_A_GXwDeevO2_1),.clk(gclk));
	jdff dff_A_1kAzhMjp9_1(.dout(w_dff_A_GXwDeevO2_1),.din(w_dff_A_1kAzhMjp9_1),.clk(gclk));
	jdff dff_A_hwuFFAAX3_1(.dout(w_dff_A_1kAzhMjp9_1),.din(w_dff_A_hwuFFAAX3_1),.clk(gclk));
	jdff dff_A_MOddnX0B8_1(.dout(w_dff_A_hwuFFAAX3_1),.din(w_dff_A_MOddnX0B8_1),.clk(gclk));
	jdff dff_A_FfDxJoP55_1(.dout(w_dff_A_MOddnX0B8_1),.din(w_dff_A_FfDxJoP55_1),.clk(gclk));
	jdff dff_A_U6VAVltF6_1(.dout(w_dff_A_FfDxJoP55_1),.din(w_dff_A_U6VAVltF6_1),.clk(gclk));
	jdff dff_A_wKyYd6S56_1(.dout(w_dff_A_U6VAVltF6_1),.din(w_dff_A_wKyYd6S56_1),.clk(gclk));
	jdff dff_A_nZJIOFmZ7_1(.dout(w_dff_A_wKyYd6S56_1),.din(w_dff_A_nZJIOFmZ7_1),.clk(gclk));
	jdff dff_A_Wm4FoYEo2_1(.dout(w_dff_A_nZJIOFmZ7_1),.din(w_dff_A_Wm4FoYEo2_1),.clk(gclk));
	jdff dff_B_b71Job3Z5_1(.din(n307),.dout(w_dff_B_b71Job3Z5_1),.clk(gclk));
	jdff dff_B_Sf1zdOW27_0(.din(n309),.dout(w_dff_B_Sf1zdOW27_0),.clk(gclk));
	jdff dff_B_LeYyGgHc9_0(.din(w_dff_B_Sf1zdOW27_0),.dout(w_dff_B_LeYyGgHc9_0),.clk(gclk));
	jdff dff_B_WWxggge34_0(.din(w_dff_B_LeYyGgHc9_0),.dout(w_dff_B_WWxggge34_0),.clk(gclk));
	jdff dff_B_8nT4UyrV7_0(.din(w_dff_B_WWxggge34_0),.dout(w_dff_B_8nT4UyrV7_0),.clk(gclk));
	jdff dff_B_eN03l9Bm9_0(.din(w_dff_B_8nT4UyrV7_0),.dout(w_dff_B_eN03l9Bm9_0),.clk(gclk));
	jdff dff_B_3ValmUWV0_0(.din(w_dff_B_eN03l9Bm9_0),.dout(w_dff_B_3ValmUWV0_0),.clk(gclk));
	jdff dff_B_ZolByrk60_1(.din(n304),.dout(w_dff_B_ZolByrk60_1),.clk(gclk));
	jdff dff_B_wsv61f505_1(.din(n410),.dout(w_dff_B_wsv61f505_1),.clk(gclk));
	jdff dff_B_J9Wx4gGl4_1(.din(w_dff_B_wsv61f505_1),.dout(w_dff_B_J9Wx4gGl4_1),.clk(gclk));
	jdff dff_B_G73jK7Yv0_1(.din(w_dff_B_J9Wx4gGl4_1),.dout(w_dff_B_G73jK7Yv0_1),.clk(gclk));
	jdff dff_B_YZqZ1I5a4_1(.din(w_dff_B_G73jK7Yv0_1),.dout(w_dff_B_YZqZ1I5a4_1),.clk(gclk));
	jdff dff_B_6zkGhcqR0_1(.din(w_dff_B_YZqZ1I5a4_1),.dout(w_dff_B_6zkGhcqR0_1),.clk(gclk));
	jdff dff_B_iL7YsaSi3_1(.din(w_dff_B_6zkGhcqR0_1),.dout(w_dff_B_iL7YsaSi3_1),.clk(gclk));
	jdff dff_B_mmGwhevC0_1(.din(w_dff_B_iL7YsaSi3_1),.dout(w_dff_B_mmGwhevC0_1),.clk(gclk));
	jdff dff_B_y9yv7Atf3_1(.din(w_dff_B_mmGwhevC0_1),.dout(w_dff_B_y9yv7Atf3_1),.clk(gclk));
	jdff dff_B_otcIjMka3_1(.din(w_dff_B_y9yv7Atf3_1),.dout(w_dff_B_otcIjMka3_1),.clk(gclk));
	jdff dff_B_Y9GjR7lO0_1(.din(w_dff_B_otcIjMka3_1),.dout(w_dff_B_Y9GjR7lO0_1),.clk(gclk));
	jdff dff_B_GbNwPoWg2_1(.din(w_dff_B_Y9GjR7lO0_1),.dout(w_dff_B_GbNwPoWg2_1),.clk(gclk));
	jdff dff_B_kHNch1gY8_1(.din(n411),.dout(w_dff_B_kHNch1gY8_1),.clk(gclk));
	jdff dff_B_RpbT6EdF9_0(.din(n412),.dout(w_dff_B_RpbT6EdF9_0),.clk(gclk));
	jdff dff_B_DX3c679I1_0(.din(w_dff_B_RpbT6EdF9_0),.dout(w_dff_B_DX3c679I1_0),.clk(gclk));
	jdff dff_B_MikbEnIR6_0(.din(w_dff_B_DX3c679I1_0),.dout(w_dff_B_MikbEnIR6_0),.clk(gclk));
	jdff dff_B_WWSsA49G4_0(.din(w_dff_B_MikbEnIR6_0),.dout(w_dff_B_WWSsA49G4_0),.clk(gclk));
	jdff dff_B_MkiFlSdV1_0(.din(w_dff_B_WWSsA49G4_0),.dout(w_dff_B_MkiFlSdV1_0),.clk(gclk));
	jdff dff_B_y4HYu6Jw1_0(.din(w_dff_B_MkiFlSdV1_0),.dout(w_dff_B_y4HYu6Jw1_0),.clk(gclk));
	jdff dff_B_xlS5GCmq0_0(.din(w_dff_B_y4HYu6Jw1_0),.dout(w_dff_B_xlS5GCmq0_0),.clk(gclk));
	jdff dff_B_J6Sg49TN7_0(.din(w_dff_B_xlS5GCmq0_0),.dout(w_dff_B_J6Sg49TN7_0),.clk(gclk));
	jdff dff_B_ckyUDNnz6_0(.din(w_dff_B_J6Sg49TN7_0),.dout(w_dff_B_ckyUDNnz6_0),.clk(gclk));
	jdff dff_B_aPkeSVf45_0(.din(w_dff_B_ckyUDNnz6_0),.dout(w_dff_B_aPkeSVf45_0),.clk(gclk));
	jdff dff_B_U4V7GEKf5_0(.din(w_dff_B_aPkeSVf45_0),.dout(w_dff_B_U4V7GEKf5_0),.clk(gclk));
	jdff dff_B_NiSVb9Os5_1(.din(n387),.dout(w_dff_B_NiSVb9Os5_1),.clk(gclk));
	jdff dff_B_V5DqC9ZO5_1(.din(w_dff_B_NiSVb9Os5_1),.dout(w_dff_B_V5DqC9ZO5_1),.clk(gclk));
	jdff dff_B_NQHEajNl6_1(.din(w_dff_B_V5DqC9ZO5_1),.dout(w_dff_B_NQHEajNl6_1),.clk(gclk));
	jdff dff_B_fwR8nQXi6_1(.din(w_dff_B_NQHEajNl6_1),.dout(w_dff_B_fwR8nQXi6_1),.clk(gclk));
	jdff dff_B_Z8eQGXLn4_1(.din(w_dff_B_fwR8nQXi6_1),.dout(w_dff_B_Z8eQGXLn4_1),.clk(gclk));
	jdff dff_B_no5Sn7fN3_1(.din(w_dff_B_Z8eQGXLn4_1),.dout(w_dff_B_no5Sn7fN3_1),.clk(gclk));
	jdff dff_B_zKyFHKTi2_1(.din(w_dff_B_no5Sn7fN3_1),.dout(w_dff_B_zKyFHKTi2_1),.clk(gclk));
	jdff dff_B_dt9sWZbE6_1(.din(w_dff_B_zKyFHKTi2_1),.dout(w_dff_B_dt9sWZbE6_1),.clk(gclk));
	jdff dff_B_Ma9DwKAm4_1(.din(w_dff_B_dt9sWZbE6_1),.dout(w_dff_B_Ma9DwKAm4_1),.clk(gclk));
	jdff dff_B_FXd0XQD89_1(.din(w_dff_B_Ma9DwKAm4_1),.dout(w_dff_B_FXd0XQD89_1),.clk(gclk));
	jdff dff_B_c5FYvj8b9_1(.din(n388),.dout(w_dff_B_c5FYvj8b9_1),.clk(gclk));
	jdff dff_B_bPMLuo3p9_1(.din(w_dff_B_c5FYvj8b9_1),.dout(w_dff_B_bPMLuo3p9_1),.clk(gclk));
	jdff dff_B_el4TNwmN7_1(.din(w_dff_B_bPMLuo3p9_1),.dout(w_dff_B_el4TNwmN7_1),.clk(gclk));
	jdff dff_B_ZGdEnHiH1_1(.din(w_dff_B_el4TNwmN7_1),.dout(w_dff_B_ZGdEnHiH1_1),.clk(gclk));
	jdff dff_B_bpbVVJxx7_1(.din(w_dff_B_ZGdEnHiH1_1),.dout(w_dff_B_bpbVVJxx7_1),.clk(gclk));
	jdff dff_B_iQ7bSX4n0_1(.din(w_dff_B_bpbVVJxx7_1),.dout(w_dff_B_iQ7bSX4n0_1),.clk(gclk));
	jdff dff_B_Qiyg8Xpl5_1(.din(w_dff_B_iQ7bSX4n0_1),.dout(w_dff_B_Qiyg8Xpl5_1),.clk(gclk));
	jdff dff_B_V5OrcNKd5_1(.din(w_dff_B_Qiyg8Xpl5_1),.dout(w_dff_B_V5OrcNKd5_1),.clk(gclk));
	jdff dff_B_HjtU3Aed2_1(.din(w_dff_B_V5OrcNKd5_1),.dout(w_dff_B_HjtU3Aed2_1),.clk(gclk));
	jdff dff_A_nC3SVYna5_1(.dout(w_n329_0[1]),.din(w_dff_A_nC3SVYna5_1),.clk(gclk));
	jdff dff_A_2nvY5ech3_1(.dout(w_dff_A_nC3SVYna5_1),.din(w_dff_A_2nvY5ech3_1),.clk(gclk));
	jdff dff_A_vYh9QrKF0_1(.dout(w_dff_A_2nvY5ech3_1),.din(w_dff_A_vYh9QrKF0_1),.clk(gclk));
	jdff dff_A_7EYB9jgz2_1(.dout(w_dff_A_vYh9QrKF0_1),.din(w_dff_A_7EYB9jgz2_1),.clk(gclk));
	jdff dff_A_rEl56Bl92_1(.dout(w_dff_A_7EYB9jgz2_1),.din(w_dff_A_rEl56Bl92_1),.clk(gclk));
	jdff dff_A_F4wyE4ca0_1(.dout(w_dff_A_rEl56Bl92_1),.din(w_dff_A_F4wyE4ca0_1),.clk(gclk));
	jdff dff_A_nDCqtvNd2_1(.dout(w_dff_A_F4wyE4ca0_1),.din(w_dff_A_nDCqtvNd2_1),.clk(gclk));
	jdff dff_A_0xAL95QH9_1(.dout(w_dff_A_nDCqtvNd2_1),.din(w_dff_A_0xAL95QH9_1),.clk(gclk));
	jdff dff_A_XP5ba5uf3_1(.dout(w_dff_A_0xAL95QH9_1),.din(w_dff_A_XP5ba5uf3_1),.clk(gclk));
	jdff dff_A_cY3IRWIR9_1(.dout(w_dff_A_XP5ba5uf3_1),.din(w_dff_A_cY3IRWIR9_1),.clk(gclk));
	jdff dff_A_byFM5CMs1_1(.dout(w_n328_0[1]),.din(w_dff_A_byFM5CMs1_1),.clk(gclk));
	jdff dff_A_lWkHPceK0_1(.dout(w_dff_A_byFM5CMs1_1),.din(w_dff_A_lWkHPceK0_1),.clk(gclk));
	jdff dff_A_uLw6UAGe3_1(.dout(w_dff_A_lWkHPceK0_1),.din(w_dff_A_uLw6UAGe3_1),.clk(gclk));
	jdff dff_A_rJHttrSe5_1(.dout(w_dff_A_uLw6UAGe3_1),.din(w_dff_A_rJHttrSe5_1),.clk(gclk));
	jdff dff_A_kPEQXXh86_1(.dout(w_dff_A_rJHttrSe5_1),.din(w_dff_A_kPEQXXh86_1),.clk(gclk));
	jdff dff_A_udFDzaU99_1(.dout(w_dff_A_kPEQXXh86_1),.din(w_dff_A_udFDzaU99_1),.clk(gclk));
	jdff dff_A_ANfIQFMG9_1(.dout(w_dff_A_udFDzaU99_1),.din(w_dff_A_ANfIQFMG9_1),.clk(gclk));
	jdff dff_A_9mkipwhk5_1(.dout(w_dff_A_ANfIQFMG9_1),.din(w_dff_A_9mkipwhk5_1),.clk(gclk));
	jdff dff_A_dqMb4v3t7_1(.dout(w_dff_A_9mkipwhk5_1),.din(w_dff_A_dqMb4v3t7_1),.clk(gclk));
	jdff dff_A_YCTG0Q1d0_1(.dout(w_dff_A_dqMb4v3t7_1),.din(w_dff_A_YCTG0Q1d0_1),.clk(gclk));
	jdff dff_A_C0tNwMXZ7_1(.dout(w_dff_A_YCTG0Q1d0_1),.din(w_dff_A_C0tNwMXZ7_1),.clk(gclk));
	jdff dff_B_KYrhI0hC1_1(.din(n403),.dout(w_dff_B_KYrhI0hC1_1),.clk(gclk));
	jdff dff_B_ACO85Wrf1_0(.din(n408),.dout(w_dff_B_ACO85Wrf1_0),.clk(gclk));
	jdff dff_B_k7CZ7hhD3_0(.din(w_dff_B_ACO85Wrf1_0),.dout(w_dff_B_k7CZ7hhD3_0),.clk(gclk));
	jdff dff_B_qQoAygvn1_0(.din(n406),.dout(w_dff_B_qQoAygvn1_0),.clk(gclk));
	jdff dff_B_yqPklDZu7_0(.din(w_dff_B_qQoAygvn1_0),.dout(w_dff_B_yqPklDZu7_0),.clk(gclk));
	jdff dff_B_f31QfJbB3_0(.din(w_dff_B_yqPklDZu7_0),.dout(w_dff_B_f31QfJbB3_0),.clk(gclk));
	jdff dff_B_w6CpIRLc4_0(.din(w_dff_B_f31QfJbB3_0),.dout(w_dff_B_w6CpIRLc4_0),.clk(gclk));
	jdff dff_B_rV088fa16_0(.din(w_dff_B_w6CpIRLc4_0),.dout(w_dff_B_rV088fa16_0),.clk(gclk));
	jdff dff_B_mwsxLrJF3_0(.din(w_dff_B_rV088fa16_0),.dout(w_dff_B_mwsxLrJF3_0),.clk(gclk));
	jdff dff_B_cjMy5KA00_0(.din(w_dff_B_mwsxLrJF3_0),.dout(w_dff_B_cjMy5KA00_0),.clk(gclk));
	jdff dff_B_cs5Ker5C6_0(.din(w_dff_B_cjMy5KA00_0),.dout(w_dff_B_cs5Ker5C6_0),.clk(gclk));
	jdff dff_B_vuJxep6s2_0(.din(w_dff_B_cs5Ker5C6_0),.dout(w_dff_B_vuJxep6s2_0),.clk(gclk));
	jdff dff_B_W5jbDRS45_0(.din(w_dff_B_vuJxep6s2_0),.dout(w_dff_B_W5jbDRS45_0),.clk(gclk));
	jdff dff_A_IwDjKkBE0_1(.dout(w_n404_0[1]),.din(w_dff_A_IwDjKkBE0_1),.clk(gclk));
	jdff dff_A_3bZIFlVQ8_1(.dout(w_dff_A_IwDjKkBE0_1),.din(w_dff_A_3bZIFlVQ8_1),.clk(gclk));
	jdff dff_A_FXkBUiM52_1(.dout(w_dff_A_3bZIFlVQ8_1),.din(w_dff_A_FXkBUiM52_1),.clk(gclk));
	jdff dff_A_F4txEN0w3_1(.dout(w_dff_A_FXkBUiM52_1),.din(w_dff_A_F4txEN0w3_1),.clk(gclk));
	jdff dff_A_dCTX42Ty0_1(.dout(w_dff_A_F4txEN0w3_1),.din(w_dff_A_dCTX42Ty0_1),.clk(gclk));
	jdff dff_A_pg7rHJG33_1(.dout(w_dff_A_dCTX42Ty0_1),.din(w_dff_A_pg7rHJG33_1),.clk(gclk));
	jdff dff_A_oL28DVCB8_1(.dout(w_dff_A_pg7rHJG33_1),.din(w_dff_A_oL28DVCB8_1),.clk(gclk));
	jdff dff_A_AfHaIRxi5_1(.dout(w_dff_A_oL28DVCB8_1),.din(w_dff_A_AfHaIRxi5_1),.clk(gclk));
	jdff dff_A_flsEitT15_1(.dout(w_dff_A_AfHaIRxi5_1),.din(w_dff_A_flsEitT15_1),.clk(gclk));
	jdff dff_A_LuxiEYsX8_1(.dout(w_dff_A_flsEitT15_1),.din(w_dff_A_LuxiEYsX8_1),.clk(gclk));
	jdff dff_A_gX7i0XKC4_1(.dout(w_dff_A_LuxiEYsX8_1),.din(w_dff_A_gX7i0XKC4_1),.clk(gclk));
	jdff dff_A_xWZaWM6C1_1(.dout(w_dff_A_gX7i0XKC4_1),.din(w_dff_A_xWZaWM6C1_1),.clk(gclk));
	jdff dff_B_kmBlNeDa0_0(.din(n317),.dout(w_dff_B_kmBlNeDa0_0),.clk(gclk));
	jdff dff_B_bkn0FYDb9_0(.din(n316),.dout(w_dff_B_bkn0FYDb9_0),.clk(gclk));
	jdff dff_B_dJnYQKnp4_0(.din(w_dff_B_bkn0FYDb9_0),.dout(w_dff_B_dJnYQKnp4_0),.clk(gclk));
	jdff dff_B_lh2Yrq4M4_0(.din(w_dff_B_dJnYQKnp4_0),.dout(w_dff_B_lh2Yrq4M4_0),.clk(gclk));
	jdff dff_B_Z9TYzfVw8_0(.din(w_dff_B_lh2Yrq4M4_0),.dout(w_dff_B_Z9TYzfVw8_0),.clk(gclk));
	jdff dff_A_3XFyiUAB4_0(.dout(w_n306_1[0]),.din(w_dff_A_3XFyiUAB4_0),.clk(gclk));
	jdff dff_A_D50Szkfz6_0(.dout(w_dff_A_3XFyiUAB4_0),.din(w_dff_A_D50Szkfz6_0),.clk(gclk));
	jdff dff_B_x2OqQQJj7_1(.din(n426),.dout(w_dff_B_x2OqQQJj7_1),.clk(gclk));
	jdff dff_B_xRtgmgyj1_1(.din(w_dff_B_x2OqQQJj7_1),.dout(w_dff_B_xRtgmgyj1_1),.clk(gclk));
	jdff dff_B_dcvMEqTw1_1(.din(w_dff_B_xRtgmgyj1_1),.dout(w_dff_B_dcvMEqTw1_1),.clk(gclk));
	jdff dff_B_HNAqs8C04_1(.din(w_dff_B_dcvMEqTw1_1),.dout(w_dff_B_HNAqs8C04_1),.clk(gclk));
	jdff dff_B_s3mmBsKy9_1(.din(w_dff_B_HNAqs8C04_1),.dout(w_dff_B_s3mmBsKy9_1),.clk(gclk));
	jdff dff_B_0SBp3vsu3_1(.din(w_dff_B_s3mmBsKy9_1),.dout(w_dff_B_0SBp3vsu3_1),.clk(gclk));
	jdff dff_B_vQPr47jz8_1(.din(w_dff_B_0SBp3vsu3_1),.dout(w_dff_B_vQPr47jz8_1),.clk(gclk));
	jdff dff_B_18risy2H5_1(.din(w_dff_B_vQPr47jz8_1),.dout(w_dff_B_18risy2H5_1),.clk(gclk));
	jdff dff_B_kuM9YojE4_1(.din(w_dff_B_18risy2H5_1),.dout(w_dff_B_kuM9YojE4_1),.clk(gclk));
	jdff dff_B_mqO1nELF3_1(.din(n428),.dout(w_dff_B_mqO1nELF3_1),.clk(gclk));
	jdff dff_B_4PayGcsh8_1(.din(n340),.dout(w_dff_B_4PayGcsh8_1),.clk(gclk));
	jdff dff_B_MHy3BuVX4_1(.din(w_dff_B_4PayGcsh8_1),.dout(w_dff_B_MHy3BuVX4_1),.clk(gclk));
	jdff dff_B_x5888I8n6_1(.din(w_dff_B_MHy3BuVX4_1),.dout(w_dff_B_x5888I8n6_1),.clk(gclk));
	jdff dff_B_Gbl7UWRP9_1(.din(w_dff_B_x5888I8n6_1),.dout(w_dff_B_Gbl7UWRP9_1),.clk(gclk));
	jdff dff_B_74pt3QHk6_1(.din(w_dff_B_Gbl7UWRP9_1),.dout(w_dff_B_74pt3QHk6_1),.clk(gclk));
	jdff dff_B_tybF7BoW7_1(.din(w_dff_B_74pt3QHk6_1),.dout(w_dff_B_tybF7BoW7_1),.clk(gclk));
	jdff dff_B_J5ysfJUO0_1(.din(n344),.dout(w_dff_B_J5ysfJUO0_1),.clk(gclk));
	jdff dff_B_Fu1JlMXh1_1(.din(w_dff_B_J5ysfJUO0_1),.dout(w_dff_B_Fu1JlMXh1_1),.clk(gclk));
	jdff dff_B_xWFVi4sX9_1(.din(w_dff_B_Fu1JlMXh1_1),.dout(w_dff_B_xWFVi4sX9_1),.clk(gclk));
	jdff dff_B_fzwK6v1P7_1(.din(w_dff_B_xWFVi4sX9_1),.dout(w_dff_B_fzwK6v1P7_1),.clk(gclk));
	jdff dff_B_cvIQccYk8_1(.din(w_dff_B_fzwK6v1P7_1),.dout(w_dff_B_cvIQccYk8_1),.clk(gclk));
	jdff dff_B_Ymb89kTl0_0(.din(n171),.dout(w_dff_B_Ymb89kTl0_0),.clk(gclk));
	jdff dff_A_6pwiBZiD1_1(.dout(w_G219gat_1[1]),.din(w_dff_A_6pwiBZiD1_1),.clk(gclk));
	jdff dff_A_RWZmEWs59_1(.dout(w_dff_A_6pwiBZiD1_1),.din(w_dff_A_RWZmEWs59_1),.clk(gclk));
	jdff dff_A_JONvI4Ah7_2(.dout(w_G219gat_1[2]),.din(w_dff_A_JONvI4Ah7_2),.clk(gclk));
	jdff dff_A_GyAh0DSE4_2(.dout(w_dff_A_JONvI4Ah7_2),.din(w_dff_A_GyAh0DSE4_2),.clk(gclk));
	jdff dff_A_SI1dviB09_2(.dout(w_dff_A_GyAh0DSE4_2),.din(w_dff_A_SI1dviB09_2),.clk(gclk));
	jdff dff_A_IYzUJds28_2(.dout(w_dff_A_SI1dviB09_2),.din(w_dff_A_IYzUJds28_2),.clk(gclk));
	jdff dff_A_EMlu2N5b4_0(.dout(w_G219gat_0[0]),.din(w_dff_A_EMlu2N5b4_0),.clk(gclk));
	jdff dff_A_Ti5cg5ph1_0(.dout(w_dff_A_EMlu2N5b4_0),.din(w_dff_A_Ti5cg5ph1_0),.clk(gclk));
	jdff dff_A_PGDTSPWh0_0(.dout(w_dff_A_Ti5cg5ph1_0),.din(w_dff_A_PGDTSPWh0_0),.clk(gclk));
	jdff dff_A_hdvXsXBp9_0(.dout(w_dff_A_PGDTSPWh0_0),.din(w_dff_A_hdvXsXBp9_0),.clk(gclk));
	jdff dff_A_MoIeqth39_0(.dout(w_dff_A_hdvXsXBp9_0),.din(w_dff_A_MoIeqth39_0),.clk(gclk));
	jdff dff_A_JtfTxExS7_0(.dout(w_dff_A_MoIeqth39_0),.din(w_dff_A_JtfTxExS7_0),.clk(gclk));
	jdff dff_A_QzQoHkma3_0(.dout(w_dff_A_JtfTxExS7_0),.din(w_dff_A_QzQoHkma3_0),.clk(gclk));
	jdff dff_A_Ib2ld3B62_0(.dout(w_dff_A_QzQoHkma3_0),.din(w_dff_A_Ib2ld3B62_0),.clk(gclk));
	jdff dff_A_k8q9eGSe7_0(.dout(w_dff_A_Ib2ld3B62_0),.din(w_dff_A_k8q9eGSe7_0),.clk(gclk));
	jdff dff_A_2HLhW8dn4_1(.dout(w_G219gat_0[1]),.din(w_dff_A_2HLhW8dn4_1),.clk(gclk));
	jdff dff_B_nealyHUp2_3(.din(G219gat),.dout(w_dff_B_nealyHUp2_3),.clk(gclk));
	jdff dff_B_xtI4oHHV2_3(.din(w_dff_B_nealyHUp2_3),.dout(w_dff_B_xtI4oHHV2_3),.clk(gclk));
	jdff dff_B_bayc14bM7_3(.din(w_dff_B_xtI4oHHV2_3),.dout(w_dff_B_bayc14bM7_3),.clk(gclk));
	jdff dff_B_0i1sCJu34_3(.din(w_dff_B_bayc14bM7_3),.dout(w_dff_B_0i1sCJu34_3),.clk(gclk));
	jdff dff_B_byz4GMMS8_3(.din(w_dff_B_0i1sCJu34_3),.dout(w_dff_B_byz4GMMS8_3),.clk(gclk));
	jdff dff_B_6th8OTEB6_3(.din(w_dff_B_byz4GMMS8_3),.dout(w_dff_B_6th8OTEB6_3),.clk(gclk));
	jdff dff_B_YsyELdkb6_3(.din(w_dff_B_6th8OTEB6_3),.dout(w_dff_B_YsyELdkb6_3),.clk(gclk));
	jdff dff_B_ADMuWfEC4_3(.din(w_dff_B_YsyELdkb6_3),.dout(w_dff_B_ADMuWfEC4_3),.clk(gclk));
	jdff dff_B_CBt1BKL09_3(.din(w_dff_B_ADMuWfEC4_3),.dout(w_dff_B_CBt1BKL09_3),.clk(gclk));
	jdff dff_B_ZbozWSWy9_3(.din(w_dff_B_CBt1BKL09_3),.dout(w_dff_B_ZbozWSWy9_3),.clk(gclk));
	jdff dff_B_GMdIAMAk0_3(.din(w_dff_B_ZbozWSWy9_3),.dout(w_dff_B_GMdIAMAk0_3),.clk(gclk));
	jdff dff_B_HuHRgb4z3_3(.din(w_dff_B_GMdIAMAk0_3),.dout(w_dff_B_HuHRgb4z3_3),.clk(gclk));
	jdff dff_B_yd3rmF5e8_0(.din(n427),.dout(w_dff_B_yd3rmF5e8_0),.clk(gclk));
	jdff dff_B_tVoOs6xB3_0(.din(w_dff_B_yd3rmF5e8_0),.dout(w_dff_B_tVoOs6xB3_0),.clk(gclk));
	jdff dff_B_HnNJIOhJ6_0(.din(w_dff_B_tVoOs6xB3_0),.dout(w_dff_B_HnNJIOhJ6_0),.clk(gclk));
	jdff dff_B_2B2v49to7_0(.din(w_dff_B_HnNJIOhJ6_0),.dout(w_dff_B_2B2v49to7_0),.clk(gclk));
	jdff dff_B_rwgBmrGf7_0(.din(w_dff_B_2B2v49to7_0),.dout(w_dff_B_rwgBmrGf7_0),.clk(gclk));
	jdff dff_B_YwmusE7S0_0(.din(w_dff_B_rwgBmrGf7_0),.dout(w_dff_B_YwmusE7S0_0),.clk(gclk));
	jdff dff_B_92mOriVu0_0(.din(w_dff_B_YwmusE7S0_0),.dout(w_dff_B_92mOriVu0_0),.clk(gclk));
	jdff dff_B_cUIJ56Cx7_0(.din(w_dff_B_92mOriVu0_0),.dout(w_dff_B_cUIJ56Cx7_0),.clk(gclk));
	jdff dff_B_eCn0yA8Z3_0(.din(w_dff_B_cUIJ56Cx7_0),.dout(w_dff_B_eCn0yA8Z3_0),.clk(gclk));
	jdff dff_B_sDhUd0Mh1_1(.din(n389),.dout(w_dff_B_sDhUd0Mh1_1),.clk(gclk));
	jdff dff_B_hXqSAjS32_1(.din(w_dff_B_sDhUd0Mh1_1),.dout(w_dff_B_hXqSAjS32_1),.clk(gclk));
	jdff dff_B_PotbSWsY0_1(.din(w_dff_B_hXqSAjS32_1),.dout(w_dff_B_PotbSWsY0_1),.clk(gclk));
	jdff dff_B_lcAPsD593_1(.din(w_dff_B_PotbSWsY0_1),.dout(w_dff_B_lcAPsD593_1),.clk(gclk));
	jdff dff_B_ffLRV7A62_1(.din(w_dff_B_lcAPsD593_1),.dout(w_dff_B_ffLRV7A62_1),.clk(gclk));
	jdff dff_B_TsYMy0rj5_1(.din(w_dff_B_ffLRV7A62_1),.dout(w_dff_B_TsYMy0rj5_1),.clk(gclk));
	jdff dff_B_7RhKTItA8_1(.din(w_dff_B_TsYMy0rj5_1),.dout(w_dff_B_7RhKTItA8_1),.clk(gclk));
	jdff dff_B_BnHVhi8v1_1(.din(w_dff_B_7RhKTItA8_1),.dout(w_dff_B_BnHVhi8v1_1),.clk(gclk));
	jdff dff_B_J3NRScyI2_1(.din(n359),.dout(w_dff_B_J3NRScyI2_1),.clk(gclk));
	jdff dff_B_VDeR1XEv4_1(.din(w_dff_B_J3NRScyI2_1),.dout(w_dff_B_VDeR1XEv4_1),.clk(gclk));
	jdff dff_B_VzH4R8Tb0_1(.din(w_dff_B_VDeR1XEv4_1),.dout(w_dff_B_VzH4R8Tb0_1),.clk(gclk));
	jdff dff_B_HA636BSQ9_1(.din(w_dff_B_VzH4R8Tb0_1),.dout(w_dff_B_HA636BSQ9_1),.clk(gclk));
	jdff dff_B_oSafIrro8_1(.din(w_dff_B_HA636BSQ9_1),.dout(w_dff_B_oSafIrro8_1),.clk(gclk));
	jdff dff_B_vIeKzdDZ5_1(.din(w_dff_B_oSafIrro8_1),.dout(w_dff_B_vIeKzdDZ5_1),.clk(gclk));
	jdff dff_B_D2Y4UE0M3_1(.din(w_dff_B_vIeKzdDZ5_1),.dout(w_dff_B_D2Y4UE0M3_1),.clk(gclk));
	jdff dff_B_MMyIBFcg6_1(.din(n252),.dout(w_dff_B_MMyIBFcg6_1),.clk(gclk));
	jdff dff_B_fX5KxfZH6_1(.din(w_dff_B_MMyIBFcg6_1),.dout(w_dff_B_fX5KxfZH6_1),.clk(gclk));
	jdff dff_B_DPoa9dGu1_1(.din(w_dff_B_fX5KxfZH6_1),.dout(w_dff_B_DPoa9dGu1_1),.clk(gclk));
	jdff dff_B_oueMcbXP4_1(.din(w_dff_B_DPoa9dGu1_1),.dout(w_dff_B_oueMcbXP4_1),.clk(gclk));
	jdff dff_B_iqUzzj4d5_1(.din(w_dff_B_oueMcbXP4_1),.dout(w_dff_B_iqUzzj4d5_1),.clk(gclk));
	jdff dff_B_BWLpF0KT9_1(.din(n253),.dout(w_dff_B_BWLpF0KT9_1),.clk(gclk));
	jdff dff_B_dO6qtV3b4_1(.din(w_dff_B_BWLpF0KT9_1),.dout(w_dff_B_dO6qtV3b4_1),.clk(gclk));
	jdff dff_B_IEyFdywL9_1(.din(w_dff_B_dO6qtV3b4_1),.dout(w_dff_B_IEyFdywL9_1),.clk(gclk));
	jdff dff_B_bjbKh9n43_1(.din(w_dff_B_IEyFdywL9_1),.dout(w_dff_B_bjbKh9n43_1),.clk(gclk));
	jdff dff_B_Y1UyWR7U8_1(.din(n254),.dout(w_dff_B_Y1UyWR7U8_1),.clk(gclk));
	jdff dff_B_JwNGO53n3_1(.din(w_dff_B_Y1UyWR7U8_1),.dout(w_dff_B_JwNGO53n3_1),.clk(gclk));
	jdff dff_B_zVRLC9Ba5_1(.din(w_dff_B_JwNGO53n3_1),.dout(w_dff_B_zVRLC9Ba5_1),.clk(gclk));
	jdff dff_B_COuJfQxM1_1(.din(n255),.dout(w_dff_B_COuJfQxM1_1),.clk(gclk));
	jdff dff_B_1yNXocHa2_1(.din(w_dff_B_COuJfQxM1_1),.dout(w_dff_B_1yNXocHa2_1),.clk(gclk));
	jdff dff_A_4cNoCPSg0_1(.dout(w_n209_0[1]),.din(w_dff_A_4cNoCPSg0_1),.clk(gclk));
	jdff dff_B_uq5YB8iY8_2(.din(n209),.dout(w_dff_B_uq5YB8iY8_2),.clk(gclk));
	jdff dff_B_FB1pJWiG3_2(.din(w_dff_B_uq5YB8iY8_2),.dout(w_dff_B_FB1pJWiG3_2),.clk(gclk));
	jdff dff_B_zU9dKjYx9_2(.din(w_dff_B_FB1pJWiG3_2),.dout(w_dff_B_zU9dKjYx9_2),.clk(gclk));
	jdff dff_B_sqAbqZFa9_2(.din(w_dff_B_zU9dKjYx9_2),.dout(w_dff_B_sqAbqZFa9_2),.clk(gclk));
	jdff dff_B_aAin9rsL6_2(.din(w_dff_B_sqAbqZFa9_2),.dout(w_dff_B_aAin9rsL6_2),.clk(gclk));
	jdff dff_B_U1QogUBc1_2(.din(w_dff_B_aAin9rsL6_2),.dout(w_dff_B_U1QogUBc1_2),.clk(gclk));
	jdff dff_B_J4gD7p7d8_2(.din(w_dff_B_U1QogUBc1_2),.dout(w_dff_B_J4gD7p7d8_2),.clk(gclk));
	jdff dff_B_V3pVTEM05_2(.din(w_dff_B_J4gD7p7d8_2),.dout(w_dff_B_V3pVTEM05_2),.clk(gclk));
	jdff dff_B_LL0ht2Ne4_2(.din(w_dff_B_V3pVTEM05_2),.dout(w_dff_B_LL0ht2Ne4_2),.clk(gclk));
	jdff dff_A_E5k1HrQO9_0(.dout(w_n242_0[0]),.din(w_dff_A_E5k1HrQO9_0),.clk(gclk));
	jdff dff_B_VKIL1KgJ4_1(.din(n182),.dout(w_dff_B_VKIL1KgJ4_1),.clk(gclk));
	jdff dff_B_uB5UaBTU2_3(.din(n181),.dout(w_dff_B_uB5UaBTU2_3),.clk(gclk));
	jdff dff_B_8JH9X9W86_3(.din(w_dff_B_uB5UaBTU2_3),.dout(w_dff_B_8JH9X9W86_3),.clk(gclk));
	jdff dff_B_wCN4TqMH2_3(.din(w_dff_B_8JH9X9W86_3),.dout(w_dff_B_wCN4TqMH2_3),.clk(gclk));
	jdff dff_B_9q4cAsx81_3(.din(w_dff_B_wCN4TqMH2_3),.dout(w_dff_B_9q4cAsx81_3),.clk(gclk));
	jdff dff_B_mF65vmDV9_3(.din(w_dff_B_9q4cAsx81_3),.dout(w_dff_B_mF65vmDV9_3),.clk(gclk));
	jdff dff_B_V1UkLjfl8_3(.din(w_dff_B_mF65vmDV9_3),.dout(w_dff_B_V1UkLjfl8_3),.clk(gclk));
	jdff dff_B_eKqibSVd7_3(.din(w_dff_B_V1UkLjfl8_3),.dout(w_dff_B_eKqibSVd7_3),.clk(gclk));
	jdff dff_B_BEqYUOMv2_3(.din(w_dff_B_eKqibSVd7_3),.dout(w_dff_B_BEqYUOMv2_3),.clk(gclk));
	jdff dff_A_CEQ0lxKp2_1(.dout(w_n241_0[1]),.din(w_dff_A_CEQ0lxKp2_1),.clk(gclk));
	jdff dff_A_qT6muqyn8_1(.dout(w_dff_A_CEQ0lxKp2_1),.din(w_dff_A_qT6muqyn8_1),.clk(gclk));
	jdff dff_A_ZuR8lNHC0_1(.dout(w_dff_A_qT6muqyn8_1),.din(w_dff_A_ZuR8lNHC0_1),.clk(gclk));
	jdff dff_A_C7z8XBoT4_1(.dout(w_n240_0[1]),.din(w_dff_A_C7z8XBoT4_1),.clk(gclk));
	jdff dff_A_XJnaNOnP7_1(.dout(w_dff_A_C7z8XBoT4_1),.din(w_dff_A_XJnaNOnP7_1),.clk(gclk));
	jdff dff_A_w6ASu1417_1(.dout(w_dff_A_XJnaNOnP7_1),.din(w_dff_A_w6ASu1417_1),.clk(gclk));
	jdff dff_A_Zzzc8CrR8_1(.dout(w_dff_A_w6ASu1417_1),.din(w_dff_A_Zzzc8CrR8_1),.clk(gclk));
	jdff dff_A_3nkQ5RB82_1(.dout(w_n235_0[1]),.din(w_dff_A_3nkQ5RB82_1),.clk(gclk));
	jdff dff_A_dn19Lk7u3_1(.dout(w_dff_A_3nkQ5RB82_1),.din(w_dff_A_dn19Lk7u3_1),.clk(gclk));
	jdff dff_A_f8gnE0gU2_1(.dout(w_dff_A_dn19Lk7u3_1),.din(w_dff_A_f8gnE0gU2_1),.clk(gclk));
	jdff dff_A_JARPD4A55_1(.dout(w_dff_A_f8gnE0gU2_1),.din(w_dff_A_JARPD4A55_1),.clk(gclk));
	jdff dff_A_0VkJRlpF6_1(.dout(w_dff_A_JARPD4A55_1),.din(w_dff_A_0VkJRlpF6_1),.clk(gclk));
	jdff dff_A_XZk3ieHp2_1(.dout(w_n234_0[1]),.din(w_dff_A_XZk3ieHp2_1),.clk(gclk));
	jdff dff_A_yN8XxgSW7_1(.dout(w_dff_A_XZk3ieHp2_1),.din(w_dff_A_yN8XxgSW7_1),.clk(gclk));
	jdff dff_A_i4ftW9cE8_1(.dout(w_dff_A_yN8XxgSW7_1),.din(w_dff_A_i4ftW9cE8_1),.clk(gclk));
	jdff dff_A_IrI6sxS90_1(.dout(w_dff_A_i4ftW9cE8_1),.din(w_dff_A_IrI6sxS90_1),.clk(gclk));
	jdff dff_A_yanv0OM79_1(.dout(w_dff_A_IrI6sxS90_1),.din(w_dff_A_yanv0OM79_1),.clk(gclk));
	jdff dff_A_npFGjXrQ4_1(.dout(w_dff_A_yanv0OM79_1),.din(w_dff_A_npFGjXrQ4_1),.clk(gclk));
	jdff dff_A_ktiDR8at9_1(.dout(w_G146gat_0[1]),.din(w_dff_A_ktiDR8at9_1),.clk(gclk));
	jdff dff_B_TpqTVJ4n0_2(.din(G146gat),.dout(w_dff_B_TpqTVJ4n0_2),.clk(gclk));
	jdff dff_B_iJFi5h6D0_2(.din(w_dff_B_TpqTVJ4n0_2),.dout(w_dff_B_iJFi5h6D0_2),.clk(gclk));
	jdff dff_B_vKcqEVzi0_2(.din(w_dff_B_iJFi5h6D0_2),.dout(w_dff_B_vKcqEVzi0_2),.clk(gclk));
	jdff dff_B_oEo3lIF12_2(.din(w_dff_B_vKcqEVzi0_2),.dout(w_dff_B_oEo3lIF12_2),.clk(gclk));
	jdff dff_A_812H5gga4_0(.dout(w_n343_0[0]),.din(w_dff_A_812H5gga4_0),.clk(gclk));
	jdff dff_A_29hTzBdz1_0(.dout(w_dff_A_812H5gga4_0),.din(w_dff_A_29hTzBdz1_0),.clk(gclk));
	jdff dff_A_RHCq5V7U5_0(.dout(w_dff_A_29hTzBdz1_0),.din(w_dff_A_RHCq5V7U5_0),.clk(gclk));
	jdff dff_A_GibsDc8A7_0(.dout(w_dff_A_RHCq5V7U5_0),.din(w_dff_A_GibsDc8A7_0),.clk(gclk));
	jdff dff_A_THLsNrii0_0(.dout(w_dff_A_GibsDc8A7_0),.din(w_dff_A_THLsNrii0_0),.clk(gclk));
	jdff dff_A_xLgms4vS7_0(.dout(w_dff_A_THLsNrii0_0),.din(w_dff_A_xLgms4vS7_0),.clk(gclk));
	jdff dff_B_3De2OvN21_1(.din(n341),.dout(w_dff_B_3De2OvN21_1),.clk(gclk));
	jdff dff_B_9s0KUMA57_1(.din(w_dff_B_3De2OvN21_1),.dout(w_dff_B_9s0KUMA57_1),.clk(gclk));
	jdff dff_B_5r88tqMS6_1(.din(w_dff_B_9s0KUMA57_1),.dout(w_dff_B_5r88tqMS6_1),.clk(gclk));
	jdff dff_B_pPLs2kKB7_1(.din(w_dff_B_5r88tqMS6_1),.dout(w_dff_B_pPLs2kKB7_1),.clk(gclk));
	jdff dff_B_rEQ14hc79_1(.din(w_dff_B_pPLs2kKB7_1),.dout(w_dff_B_rEQ14hc79_1),.clk(gclk));
	jdff dff_B_YPFORqkM5_1(.din(w_dff_B_rEQ14hc79_1),.dout(w_dff_B_YPFORqkM5_1),.clk(gclk));
	jdff dff_B_km6G1oom0_1(.din(w_dff_B_YPFORqkM5_1),.dout(w_dff_B_km6G1oom0_1),.clk(gclk));
	jdff dff_B_jf0EZXZZ0_1(.din(w_dff_B_km6G1oom0_1),.dout(w_dff_B_jf0EZXZZ0_1),.clk(gclk));
	jdff dff_A_qMP30cKL8_1(.dout(w_n222_0[1]),.din(w_dff_A_qMP30cKL8_1),.clk(gclk));
	jdff dff_A_ctMDOhS61_1(.dout(w_dff_A_qMP30cKL8_1),.din(w_dff_A_ctMDOhS61_1),.clk(gclk));
	jdff dff_A_KPw1I5xz5_1(.dout(w_dff_A_ctMDOhS61_1),.din(w_dff_A_KPw1I5xz5_1),.clk(gclk));
	jdff dff_A_CjNlyoDA3_1(.dout(w_dff_A_KPw1I5xz5_1),.din(w_dff_A_CjNlyoDA3_1),.clk(gclk));
	jdff dff_A_OB9FY0mw8_1(.dout(w_dff_A_CjNlyoDA3_1),.din(w_dff_A_OB9FY0mw8_1),.clk(gclk));
	jdff dff_A_zCvbnzqH0_1(.dout(w_dff_A_OB9FY0mw8_1),.din(w_dff_A_zCvbnzqH0_1),.clk(gclk));
	jdff dff_A_ilpXpt4I6_1(.dout(w_dff_A_zCvbnzqH0_1),.din(w_dff_A_ilpXpt4I6_1),.clk(gclk));
	jdff dff_A_FEssNtyE2_1(.dout(w_dff_A_ilpXpt4I6_1),.din(w_dff_A_FEssNtyE2_1),.clk(gclk));
	jdff dff_A_z7MgNYZq9_1(.dout(w_G143gat_0[1]),.din(w_dff_A_z7MgNYZq9_1),.clk(gclk));
	jdff dff_B_RuFuQY6l2_2(.din(G143gat),.dout(w_dff_B_RuFuQY6l2_2),.clk(gclk));
	jdff dff_B_c9eL9yPE2_2(.din(w_dff_B_RuFuQY6l2_2),.dout(w_dff_B_c9eL9yPE2_2),.clk(gclk));
	jdff dff_B_9C246Ov72_2(.din(w_dff_B_c9eL9yPE2_2),.dout(w_dff_B_9C246Ov72_2),.clk(gclk));
	jdff dff_B_XhZnIYUG3_2(.din(w_dff_B_9C246Ov72_2),.dout(w_dff_B_XhZnIYUG3_2),.clk(gclk));
	jdff dff_A_4jVZ6Q4k0_2(.dout(w_n148_1[2]),.din(w_dff_A_4jVZ6Q4k0_2),.clk(gclk));
	jdff dff_A_eyc1lp049_2(.dout(w_dff_A_4jVZ6Q4k0_2),.din(w_dff_A_eyc1lp049_2),.clk(gclk));
	jdff dff_A_vRECN8X80_0(.dout(w_n339_0[0]),.din(w_dff_A_vRECN8X80_0),.clk(gclk));
	jdff dff_A_BXbPzA7g5_0(.dout(w_dff_A_vRECN8X80_0),.din(w_dff_A_BXbPzA7g5_0),.clk(gclk));
	jdff dff_A_mqntJa0Q9_0(.dout(w_dff_A_BXbPzA7g5_0),.din(w_dff_A_mqntJa0Q9_0),.clk(gclk));
	jdff dff_A_uAXpYeU64_0(.dout(w_dff_A_mqntJa0Q9_0),.din(w_dff_A_uAXpYeU64_0),.clk(gclk));
	jdff dff_A_fHltFPqQ2_0(.dout(w_dff_A_uAXpYeU64_0),.din(w_dff_A_fHltFPqQ2_0),.clk(gclk));
	jdff dff_A_A7xyoMr72_0(.dout(w_dff_A_fHltFPqQ2_0),.din(w_dff_A_A7xyoMr72_0),.clk(gclk));
	jdff dff_A_k9lRbkI00_0(.dout(w_dff_A_A7xyoMr72_0),.din(w_dff_A_k9lRbkI00_0),.clk(gclk));
	jdff dff_B_lBgFsyx20_1(.din(n337),.dout(w_dff_B_lBgFsyx20_1),.clk(gclk));
	jdff dff_B_UWSlXJpb0_1(.din(w_dff_B_lBgFsyx20_1),.dout(w_dff_B_UWSlXJpb0_1),.clk(gclk));
	jdff dff_B_VMwBgffC5_1(.din(w_dff_B_UWSlXJpb0_1),.dout(w_dff_B_VMwBgffC5_1),.clk(gclk));
	jdff dff_B_M1Co64tr0_1(.din(w_dff_B_VMwBgffC5_1),.dout(w_dff_B_M1Co64tr0_1),.clk(gclk));
	jdff dff_B_ARK7wgVa3_1(.din(w_dff_B_M1Co64tr0_1),.dout(w_dff_B_ARK7wgVa3_1),.clk(gclk));
	jdff dff_B_B1TVZA8A8_1(.din(w_dff_B_ARK7wgVa3_1),.dout(w_dff_B_B1TVZA8A8_1),.clk(gclk));
	jdff dff_B_RLjpRnwm5_1(.din(w_dff_B_B1TVZA8A8_1),.dout(w_dff_B_RLjpRnwm5_1),.clk(gclk));
	jdff dff_B_packt20l1_1(.din(w_dff_B_RLjpRnwm5_1),.dout(w_dff_B_packt20l1_1),.clk(gclk));
	jdff dff_B_kH9XimPh4_1(.din(w_dff_B_packt20l1_1),.dout(w_dff_B_kH9XimPh4_1),.clk(gclk));
	jdff dff_A_4KfbYxTX8_2(.dout(w_n336_0[2]),.din(w_dff_A_4KfbYxTX8_2),.clk(gclk));
	jdff dff_A_a3hEkdSU9_2(.dout(w_dff_A_4KfbYxTX8_2),.din(w_dff_A_a3hEkdSU9_2),.clk(gclk));
	jdff dff_A_g8OKYjpm7_2(.dout(w_dff_A_a3hEkdSU9_2),.din(w_dff_A_g8OKYjpm7_2),.clk(gclk));
	jdff dff_A_dNObNzfW5_2(.dout(w_dff_A_g8OKYjpm7_2),.din(w_dff_A_dNObNzfW5_2),.clk(gclk));
	jdff dff_A_C9AsslSj3_2(.dout(w_dff_A_dNObNzfW5_2),.din(w_dff_A_C9AsslSj3_2),.clk(gclk));
	jdff dff_A_TqEfXRn22_2(.dout(w_dff_A_C9AsslSj3_2),.din(w_dff_A_TqEfXRn22_2),.clk(gclk));
	jdff dff_A_pYcbskS19_2(.dout(w_dff_A_TqEfXRn22_2),.din(w_dff_A_pYcbskS19_2),.clk(gclk));
	jdff dff_A_1VsQDjyT1_2(.dout(w_dff_A_pYcbskS19_2),.din(w_dff_A_1VsQDjyT1_2),.clk(gclk));
	jdff dff_A_I9q8PbWb9_2(.dout(w_dff_A_1VsQDjyT1_2),.din(w_dff_A_I9q8PbWb9_2),.clk(gclk));
	jdff dff_B_Adq0vX6W4_0(.din(n333),.dout(w_dff_B_Adq0vX6W4_0),.clk(gclk));
	jdff dff_B_njyr8vIk2_0(.din(n332),.dout(w_dff_B_njyr8vIk2_0),.clk(gclk));
	jdff dff_B_Lpn9Z3KK6_0(.din(w_dff_B_njyr8vIk2_0),.dout(w_dff_B_Lpn9Z3KK6_0),.clk(gclk));
	jdff dff_B_JG5eNFVF2_0(.din(w_dff_B_Lpn9Z3KK6_0),.dout(w_dff_B_JG5eNFVF2_0),.clk(gclk));
	jdff dff_B_3mYVtRII6_0(.din(w_dff_B_JG5eNFVF2_0),.dout(w_dff_B_3mYVtRII6_0),.clk(gclk));
	jdff dff_B_2kQkNnHJ0_1(.din(n419),.dout(w_dff_B_2kQkNnHJ0_1),.clk(gclk));
	jdff dff_B_phD424OH4_0(.din(n424),.dout(w_dff_B_phD424OH4_0),.clk(gclk));
	jdff dff_B_DSR0Iwlk1_0(.din(w_dff_B_phD424OH4_0),.dout(w_dff_B_DSR0Iwlk1_0),.clk(gclk));
	jdff dff_B_vW0l3lgO9_0(.din(n422),.dout(w_dff_B_vW0l3lgO9_0),.clk(gclk));
	jdff dff_B_AVjAxP8g4_0(.din(w_dff_B_vW0l3lgO9_0),.dout(w_dff_B_AVjAxP8g4_0),.clk(gclk));
	jdff dff_B_O7Q7vZ1q1_0(.din(w_dff_B_AVjAxP8g4_0),.dout(w_dff_B_O7Q7vZ1q1_0),.clk(gclk));
	jdff dff_B_Hz9FnoPw5_0(.din(w_dff_B_O7Q7vZ1q1_0),.dout(w_dff_B_Hz9FnoPw5_0),.clk(gclk));
	jdff dff_B_T7xEy7BW6_0(.din(w_dff_B_Hz9FnoPw5_0),.dout(w_dff_B_T7xEy7BW6_0),.clk(gclk));
	jdff dff_B_WFxQdlRu6_0(.din(w_dff_B_T7xEy7BW6_0),.dout(w_dff_B_WFxQdlRu6_0),.clk(gclk));
	jdff dff_B_7YlY6QFn3_0(.din(w_dff_B_WFxQdlRu6_0),.dout(w_dff_B_7YlY6QFn3_0),.clk(gclk));
	jdff dff_B_nK1sqyT44_0(.din(w_dff_B_7YlY6QFn3_0),.dout(w_dff_B_nK1sqyT44_0),.clk(gclk));
	jdff dff_B_oS9HL1Vp2_0(.din(w_dff_B_nK1sqyT44_0),.dout(w_dff_B_oS9HL1Vp2_0),.clk(gclk));
	jdff dff_B_fWNdO3uh7_0(.din(w_dff_B_oS9HL1Vp2_0),.dout(w_dff_B_fWNdO3uh7_0),.clk(gclk));
	jdff dff_A_3vB0jX6m8_0(.dout(w_n420_0[0]),.din(w_dff_A_3vB0jX6m8_0),.clk(gclk));
	jdff dff_A_ZkgXwSBz1_0(.dout(w_dff_A_3vB0jX6m8_0),.din(w_dff_A_ZkgXwSBz1_0),.clk(gclk));
	jdff dff_A_PumeAMUn9_0(.dout(w_dff_A_ZkgXwSBz1_0),.din(w_dff_A_PumeAMUn9_0),.clk(gclk));
	jdff dff_A_AMi2o2DU1_0(.dout(w_dff_A_PumeAMUn9_0),.din(w_dff_A_AMi2o2DU1_0),.clk(gclk));
	jdff dff_A_W951Bk605_0(.dout(w_dff_A_AMi2o2DU1_0),.din(w_dff_A_W951Bk605_0),.clk(gclk));
	jdff dff_A_ROlnZwSd1_0(.dout(w_dff_A_W951Bk605_0),.din(w_dff_A_ROlnZwSd1_0),.clk(gclk));
	jdff dff_A_ayTVddLw1_0(.dout(w_dff_A_ROlnZwSd1_0),.din(w_dff_A_ayTVddLw1_0),.clk(gclk));
	jdff dff_A_26g6vfx57_0(.dout(w_dff_A_ayTVddLw1_0),.din(w_dff_A_26g6vfx57_0),.clk(gclk));
	jdff dff_A_NULuFxEu5_0(.dout(w_dff_A_26g6vfx57_0),.din(w_dff_A_NULuFxEu5_0),.clk(gclk));
	jdff dff_A_mAAVI44v4_0(.dout(w_dff_A_NULuFxEu5_0),.din(w_dff_A_mAAVI44v4_0),.clk(gclk));
	jdff dff_A_gDQHMYla4_0(.dout(w_G228gat_0[0]),.din(w_dff_A_gDQHMYla4_0),.clk(gclk));
	jdff dff_B_e8Cptkpo8_3(.din(G228gat),.dout(w_dff_B_e8Cptkpo8_3),.clk(gclk));
	jdff dff_B_Y6SQOTPq6_3(.din(w_dff_B_e8Cptkpo8_3),.dout(w_dff_B_Y6SQOTPq6_3),.clk(gclk));
	jdff dff_B_mUnJNkGj4_3(.din(w_dff_B_Y6SQOTPq6_3),.dout(w_dff_B_mUnJNkGj4_3),.clk(gclk));
	jdff dff_B_UmB4pous4_3(.din(w_dff_B_mUnJNkGj4_3),.dout(w_dff_B_UmB4pous4_3),.clk(gclk));
	jdff dff_B_fv5ELtF35_3(.din(w_dff_B_UmB4pous4_3),.dout(w_dff_B_fv5ELtF35_3),.clk(gclk));
	jdff dff_B_fvAHvOyo3_3(.din(w_dff_B_fv5ELtF35_3),.dout(w_dff_B_fvAHvOyo3_3),.clk(gclk));
	jdff dff_B_ysQSu4lh2_3(.din(w_dff_B_fvAHvOyo3_3),.dout(w_dff_B_ysQSu4lh2_3),.clk(gclk));
	jdff dff_B_bgjsFjNt8_3(.din(w_dff_B_ysQSu4lh2_3),.dout(w_dff_B_bgjsFjNt8_3),.clk(gclk));
	jdff dff_B_ZIZCD5EV5_3(.din(w_dff_B_bgjsFjNt8_3),.dout(w_dff_B_ZIZCD5EV5_3),.clk(gclk));
	jdff dff_B_XMZ4bwEE7_0(.din(n325),.dout(w_dff_B_XMZ4bwEE7_0),.clk(gclk));
	jdff dff_B_M9ufdmyz8_0(.din(n324),.dout(w_dff_B_M9ufdmyz8_0),.clk(gclk));
	jdff dff_B_b9KVB5Ps8_0(.din(w_dff_B_M9ufdmyz8_0),.dout(w_dff_B_b9KVB5Ps8_0),.clk(gclk));
	jdff dff_B_Z2RNZhHl2_0(.din(w_dff_B_b9KVB5Ps8_0),.dout(w_dff_B_Z2RNZhHl2_0),.clk(gclk));
	jdff dff_B_D33PHtD84_0(.din(w_dff_B_Z2RNZhHl2_0),.dout(w_dff_B_D33PHtD84_0),.clk(gclk));
	jdff dff_A_GMKVTrYB1_1(.dout(w_G149gat_0[1]),.din(w_dff_A_GMKVTrYB1_1),.clk(gclk));
	jdff dff_B_eapsGmJZ7_2(.din(G149gat),.dout(w_dff_B_eapsGmJZ7_2),.clk(gclk));
	jdff dff_B_CRYdfOjP6_2(.din(w_dff_B_eapsGmJZ7_2),.dout(w_dff_B_CRYdfOjP6_2),.clk(gclk));
	jdff dff_B_mDG0AUJA2_2(.din(w_dff_B_CRYdfOjP6_2),.dout(w_dff_B_mDG0AUJA2_2),.clk(gclk));
	jdff dff_B_dNetj7Sz0_2(.din(w_dff_B_mDG0AUJA2_2),.dout(w_dff_B_dNetj7Sz0_2),.clk(gclk));
	jdff dff_B_X2HSRZXt6_1(.din(n150),.dout(w_dff_B_X2HSRZXt6_1),.clk(gclk));
	jdff dff_A_o84xzYsp9_1(.dout(w_n306_0[1]),.din(w_dff_A_o84xzYsp9_1),.clk(gclk));
	jdff dff_A_W9ACGTnI8_1(.dout(w_dff_A_o84xzYsp9_1),.din(w_dff_A_W9ACGTnI8_1),.clk(gclk));
	jdff dff_A_GZc8ihL28_2(.dout(w_n306_0[2]),.din(w_dff_A_GZc8ihL28_2),.clk(gclk));
	jdff dff_A_2cGXA9CZ0_2(.dout(w_dff_A_GZc8ihL28_2),.din(w_dff_A_2cGXA9CZ0_2),.clk(gclk));
	jdff dff_A_ClR1RSNQ7_2(.dout(w_G447gat_0[2]),.din(w_dff_A_ClR1RSNQ7_2),.clk(gclk));
	jdff dff_A_tbx6V7qa2_0(.dout(w_n86_0[0]),.din(w_dff_A_tbx6V7qa2_0),.clk(gclk));
	jdff dff_A_hCZC8D6S0_0(.dout(w_dff_A_tbx6V7qa2_0),.din(w_dff_A_hCZC8D6S0_0),.clk(gclk));
	jdff dff_B_AvgRFnk69_2(.din(n144),.dout(w_dff_B_AvgRFnk69_2),.clk(gclk));
	jdff dff_B_cbwv2hc83_2(.din(w_dff_B_AvgRFnk69_2),.dout(w_dff_B_cbwv2hc83_2),.clk(gclk));
	jdff dff_B_XH2BfRRp4_2(.din(w_dff_B_cbwv2hc83_2),.dout(w_dff_B_XH2BfRRp4_2),.clk(gclk));
	jdff dff_B_hBYn5AJP7_2(.din(w_dff_B_XH2BfRRp4_2),.dout(w_dff_B_hBYn5AJP7_2),.clk(gclk));
	jdff dff_A_c5h1KxxZ5_2(.dout(w_dff_A_0hz0x1rk4_0),.din(w_dff_A_c5h1KxxZ5_2),.clk(gclk));
	jdff dff_A_0hz0x1rk4_0(.dout(w_dff_A_lzBRTOd43_0),.din(w_dff_A_0hz0x1rk4_0),.clk(gclk));
	jdff dff_A_lzBRTOd43_0(.dout(w_dff_A_LuIFG4NY8_0),.din(w_dff_A_lzBRTOd43_0),.clk(gclk));
	jdff dff_A_LuIFG4NY8_0(.dout(w_dff_A_OjtJI3LO3_0),.din(w_dff_A_LuIFG4NY8_0),.clk(gclk));
	jdff dff_A_OjtJI3LO3_0(.dout(w_dff_A_kNatINEV2_0),.din(w_dff_A_OjtJI3LO3_0),.clk(gclk));
	jdff dff_A_kNatINEV2_0(.dout(w_dff_A_ahb4I5EB5_0),.din(w_dff_A_kNatINEV2_0),.clk(gclk));
	jdff dff_A_ahb4I5EB5_0(.dout(w_dff_A_HKZnpPuc7_0),.din(w_dff_A_ahb4I5EB5_0),.clk(gclk));
	jdff dff_A_HKZnpPuc7_0(.dout(w_dff_A_gITBhv6J7_0),.din(w_dff_A_HKZnpPuc7_0),.clk(gclk));
	jdff dff_A_gITBhv6J7_0(.dout(w_dff_A_squcgHag0_0),.din(w_dff_A_gITBhv6J7_0),.clk(gclk));
	jdff dff_A_squcgHag0_0(.dout(w_dff_A_Tfn9dkpY0_0),.din(w_dff_A_squcgHag0_0),.clk(gclk));
	jdff dff_A_Tfn9dkpY0_0(.dout(w_dff_A_hu1UzQuk0_0),.din(w_dff_A_Tfn9dkpY0_0),.clk(gclk));
	jdff dff_A_hu1UzQuk0_0(.dout(w_dff_A_DDJjnWAb7_0),.din(w_dff_A_hu1UzQuk0_0),.clk(gclk));
	jdff dff_A_DDJjnWAb7_0(.dout(w_dff_A_wAENiHcK5_0),.din(w_dff_A_DDJjnWAb7_0),.clk(gclk));
	jdff dff_A_wAENiHcK5_0(.dout(w_dff_A_BRk26rU56_0),.din(w_dff_A_wAENiHcK5_0),.clk(gclk));
	jdff dff_A_BRk26rU56_0(.dout(w_dff_A_Kjt2lBi47_0),.din(w_dff_A_BRk26rU56_0),.clk(gclk));
	jdff dff_A_Kjt2lBi47_0(.dout(w_dff_A_I77dcwIH0_0),.din(w_dff_A_Kjt2lBi47_0),.clk(gclk));
	jdff dff_A_I77dcwIH0_0(.dout(w_dff_A_lrcGNN8K0_0),.din(w_dff_A_I77dcwIH0_0),.clk(gclk));
	jdff dff_A_lrcGNN8K0_0(.dout(w_dff_A_xqktSLiR8_0),.din(w_dff_A_lrcGNN8K0_0),.clk(gclk));
	jdff dff_A_xqktSLiR8_0(.dout(w_dff_A_xyAdLGRP0_0),.din(w_dff_A_xqktSLiR8_0),.clk(gclk));
	jdff dff_A_xyAdLGRP0_0(.dout(w_dff_A_mTfym79l9_0),.din(w_dff_A_xyAdLGRP0_0),.clk(gclk));
	jdff dff_A_mTfym79l9_0(.dout(w_dff_A_kKppd7Q86_0),.din(w_dff_A_mTfym79l9_0),.clk(gclk));
	jdff dff_A_kKppd7Q86_0(.dout(w_dff_A_Coh57M5J7_0),.din(w_dff_A_kKppd7Q86_0),.clk(gclk));
	jdff dff_A_Coh57M5J7_0(.dout(w_dff_A_9kXdEFYu4_0),.din(w_dff_A_Coh57M5J7_0),.clk(gclk));
	jdff dff_A_9kXdEFYu4_0(.dout(w_dff_A_ovCiETst6_0),.din(w_dff_A_9kXdEFYu4_0),.clk(gclk));
	jdff dff_A_ovCiETst6_0(.dout(w_dff_A_jlWpYqjF7_0),.din(w_dff_A_ovCiETst6_0),.clk(gclk));
	jdff dff_A_jlWpYqjF7_0(.dout(G388gat),.din(w_dff_A_jlWpYqjF7_0),.clk(gclk));
	jdff dff_A_YHZgzuPt7_2(.dout(w_dff_A_2pj7O4Oz1_0),.din(w_dff_A_YHZgzuPt7_2),.clk(gclk));
	jdff dff_A_2pj7O4Oz1_0(.dout(w_dff_A_p5iXJXfI3_0),.din(w_dff_A_2pj7O4Oz1_0),.clk(gclk));
	jdff dff_A_p5iXJXfI3_0(.dout(w_dff_A_kmHT3BLT7_0),.din(w_dff_A_p5iXJXfI3_0),.clk(gclk));
	jdff dff_A_kmHT3BLT7_0(.dout(w_dff_A_CBHOuStn6_0),.din(w_dff_A_kmHT3BLT7_0),.clk(gclk));
	jdff dff_A_CBHOuStn6_0(.dout(w_dff_A_7jEBTaXk6_0),.din(w_dff_A_CBHOuStn6_0),.clk(gclk));
	jdff dff_A_7jEBTaXk6_0(.dout(w_dff_A_fiGJKQ7K0_0),.din(w_dff_A_7jEBTaXk6_0),.clk(gclk));
	jdff dff_A_fiGJKQ7K0_0(.dout(w_dff_A_t9yd53Aj8_0),.din(w_dff_A_fiGJKQ7K0_0),.clk(gclk));
	jdff dff_A_t9yd53Aj8_0(.dout(w_dff_A_Z4cNUS6r7_0),.din(w_dff_A_t9yd53Aj8_0),.clk(gclk));
	jdff dff_A_Z4cNUS6r7_0(.dout(w_dff_A_fJNDyBEI4_0),.din(w_dff_A_Z4cNUS6r7_0),.clk(gclk));
	jdff dff_A_fJNDyBEI4_0(.dout(w_dff_A_jLWAwJhD5_0),.din(w_dff_A_fJNDyBEI4_0),.clk(gclk));
	jdff dff_A_jLWAwJhD5_0(.dout(w_dff_A_9GjkLUdN6_0),.din(w_dff_A_jLWAwJhD5_0),.clk(gclk));
	jdff dff_A_9GjkLUdN6_0(.dout(w_dff_A_RA0lXuQX4_0),.din(w_dff_A_9GjkLUdN6_0),.clk(gclk));
	jdff dff_A_RA0lXuQX4_0(.dout(w_dff_A_g9CnU2Mo3_0),.din(w_dff_A_RA0lXuQX4_0),.clk(gclk));
	jdff dff_A_g9CnU2Mo3_0(.dout(w_dff_A_kTSVgl7x6_0),.din(w_dff_A_g9CnU2Mo3_0),.clk(gclk));
	jdff dff_A_kTSVgl7x6_0(.dout(w_dff_A_aEuud5z42_0),.din(w_dff_A_kTSVgl7x6_0),.clk(gclk));
	jdff dff_A_aEuud5z42_0(.dout(w_dff_A_9wEAD8aZ8_0),.din(w_dff_A_aEuud5z42_0),.clk(gclk));
	jdff dff_A_9wEAD8aZ8_0(.dout(w_dff_A_Kk07Xzig4_0),.din(w_dff_A_9wEAD8aZ8_0),.clk(gclk));
	jdff dff_A_Kk07Xzig4_0(.dout(w_dff_A_j7h72xcg4_0),.din(w_dff_A_Kk07Xzig4_0),.clk(gclk));
	jdff dff_A_j7h72xcg4_0(.dout(w_dff_A_s0ZNuBuv9_0),.din(w_dff_A_j7h72xcg4_0),.clk(gclk));
	jdff dff_A_s0ZNuBuv9_0(.dout(w_dff_A_8Ojp18G63_0),.din(w_dff_A_s0ZNuBuv9_0),.clk(gclk));
	jdff dff_A_8Ojp18G63_0(.dout(w_dff_A_VvWr8UZz5_0),.din(w_dff_A_8Ojp18G63_0),.clk(gclk));
	jdff dff_A_VvWr8UZz5_0(.dout(w_dff_A_ycyIkFor0_0),.din(w_dff_A_VvWr8UZz5_0),.clk(gclk));
	jdff dff_A_ycyIkFor0_0(.dout(w_dff_A_iPSVez904_0),.din(w_dff_A_ycyIkFor0_0),.clk(gclk));
	jdff dff_A_iPSVez904_0(.dout(w_dff_A_hjVCQoff5_0),.din(w_dff_A_iPSVez904_0),.clk(gclk));
	jdff dff_A_hjVCQoff5_0(.dout(w_dff_A_bXcbNNkp5_0),.din(w_dff_A_hjVCQoff5_0),.clk(gclk));
	jdff dff_A_bXcbNNkp5_0(.dout(G389gat),.din(w_dff_A_bXcbNNkp5_0),.clk(gclk));
	jdff dff_A_7Fl3brhr8_2(.dout(w_dff_A_Vj7jclsq4_0),.din(w_dff_A_7Fl3brhr8_2),.clk(gclk));
	jdff dff_A_Vj7jclsq4_0(.dout(w_dff_A_PxxECmuW9_0),.din(w_dff_A_Vj7jclsq4_0),.clk(gclk));
	jdff dff_A_PxxECmuW9_0(.dout(w_dff_A_QJMYOs5p5_0),.din(w_dff_A_PxxECmuW9_0),.clk(gclk));
	jdff dff_A_QJMYOs5p5_0(.dout(w_dff_A_IFUgtrnu2_0),.din(w_dff_A_QJMYOs5p5_0),.clk(gclk));
	jdff dff_A_IFUgtrnu2_0(.dout(w_dff_A_NlNE6MGn6_0),.din(w_dff_A_IFUgtrnu2_0),.clk(gclk));
	jdff dff_A_NlNE6MGn6_0(.dout(w_dff_A_FRXKEXcd8_0),.din(w_dff_A_NlNE6MGn6_0),.clk(gclk));
	jdff dff_A_FRXKEXcd8_0(.dout(w_dff_A_H4UR5eXj1_0),.din(w_dff_A_FRXKEXcd8_0),.clk(gclk));
	jdff dff_A_H4UR5eXj1_0(.dout(w_dff_A_V18BWkYp0_0),.din(w_dff_A_H4UR5eXj1_0),.clk(gclk));
	jdff dff_A_V18BWkYp0_0(.dout(w_dff_A_pln6gSJq9_0),.din(w_dff_A_V18BWkYp0_0),.clk(gclk));
	jdff dff_A_pln6gSJq9_0(.dout(w_dff_A_43AVfQz67_0),.din(w_dff_A_pln6gSJq9_0),.clk(gclk));
	jdff dff_A_43AVfQz67_0(.dout(w_dff_A_h0mk5r0I2_0),.din(w_dff_A_43AVfQz67_0),.clk(gclk));
	jdff dff_A_h0mk5r0I2_0(.dout(w_dff_A_yylNi8HB5_0),.din(w_dff_A_h0mk5r0I2_0),.clk(gclk));
	jdff dff_A_yylNi8HB5_0(.dout(w_dff_A_SMwMkbNL2_0),.din(w_dff_A_yylNi8HB5_0),.clk(gclk));
	jdff dff_A_SMwMkbNL2_0(.dout(w_dff_A_5CimCWX73_0),.din(w_dff_A_SMwMkbNL2_0),.clk(gclk));
	jdff dff_A_5CimCWX73_0(.dout(w_dff_A_TVNGGGuQ7_0),.din(w_dff_A_5CimCWX73_0),.clk(gclk));
	jdff dff_A_TVNGGGuQ7_0(.dout(w_dff_A_2YrnX8Nc4_0),.din(w_dff_A_TVNGGGuQ7_0),.clk(gclk));
	jdff dff_A_2YrnX8Nc4_0(.dout(w_dff_A_HSrhI1nk6_0),.din(w_dff_A_2YrnX8Nc4_0),.clk(gclk));
	jdff dff_A_HSrhI1nk6_0(.dout(w_dff_A_yFiJAvbr8_0),.din(w_dff_A_HSrhI1nk6_0),.clk(gclk));
	jdff dff_A_yFiJAvbr8_0(.dout(w_dff_A_WzppOk8E1_0),.din(w_dff_A_yFiJAvbr8_0),.clk(gclk));
	jdff dff_A_WzppOk8E1_0(.dout(w_dff_A_ZBK14rFI0_0),.din(w_dff_A_WzppOk8E1_0),.clk(gclk));
	jdff dff_A_ZBK14rFI0_0(.dout(w_dff_A_T0ZiEYZJ3_0),.din(w_dff_A_ZBK14rFI0_0),.clk(gclk));
	jdff dff_A_T0ZiEYZJ3_0(.dout(w_dff_A_302dtReM9_0),.din(w_dff_A_T0ZiEYZJ3_0),.clk(gclk));
	jdff dff_A_302dtReM9_0(.dout(w_dff_A_Zlz96OXR9_0),.din(w_dff_A_302dtReM9_0),.clk(gclk));
	jdff dff_A_Zlz96OXR9_0(.dout(w_dff_A_6xOEEjyv3_0),.din(w_dff_A_Zlz96OXR9_0),.clk(gclk));
	jdff dff_A_6xOEEjyv3_0(.dout(w_dff_A_VsgpJBsG9_0),.din(w_dff_A_6xOEEjyv3_0),.clk(gclk));
	jdff dff_A_VsgpJBsG9_0(.dout(G390gat),.din(w_dff_A_VsgpJBsG9_0),.clk(gclk));
	jdff dff_A_5rAfykWU6_2(.dout(w_dff_A_CzzcoIrD4_0),.din(w_dff_A_5rAfykWU6_2),.clk(gclk));
	jdff dff_A_CzzcoIrD4_0(.dout(w_dff_A_ex3mqZMD4_0),.din(w_dff_A_CzzcoIrD4_0),.clk(gclk));
	jdff dff_A_ex3mqZMD4_0(.dout(w_dff_A_NTp0Tono1_0),.din(w_dff_A_ex3mqZMD4_0),.clk(gclk));
	jdff dff_A_NTp0Tono1_0(.dout(w_dff_A_hFM5zlto8_0),.din(w_dff_A_NTp0Tono1_0),.clk(gclk));
	jdff dff_A_hFM5zlto8_0(.dout(w_dff_A_onB6vq4B5_0),.din(w_dff_A_hFM5zlto8_0),.clk(gclk));
	jdff dff_A_onB6vq4B5_0(.dout(w_dff_A_p73G01dB3_0),.din(w_dff_A_onB6vq4B5_0),.clk(gclk));
	jdff dff_A_p73G01dB3_0(.dout(w_dff_A_laiYJfCm3_0),.din(w_dff_A_p73G01dB3_0),.clk(gclk));
	jdff dff_A_laiYJfCm3_0(.dout(w_dff_A_4uKSTSHW0_0),.din(w_dff_A_laiYJfCm3_0),.clk(gclk));
	jdff dff_A_4uKSTSHW0_0(.dout(w_dff_A_CjUlM47D4_0),.din(w_dff_A_4uKSTSHW0_0),.clk(gclk));
	jdff dff_A_CjUlM47D4_0(.dout(w_dff_A_oaxb6zZz4_0),.din(w_dff_A_CjUlM47D4_0),.clk(gclk));
	jdff dff_A_oaxb6zZz4_0(.dout(w_dff_A_toC1T2xZ3_0),.din(w_dff_A_oaxb6zZz4_0),.clk(gclk));
	jdff dff_A_toC1T2xZ3_0(.dout(w_dff_A_vbgWhGs84_0),.din(w_dff_A_toC1T2xZ3_0),.clk(gclk));
	jdff dff_A_vbgWhGs84_0(.dout(w_dff_A_FoUtZfni6_0),.din(w_dff_A_vbgWhGs84_0),.clk(gclk));
	jdff dff_A_FoUtZfni6_0(.dout(w_dff_A_2rpz6Gtd8_0),.din(w_dff_A_FoUtZfni6_0),.clk(gclk));
	jdff dff_A_2rpz6Gtd8_0(.dout(w_dff_A_ZLLxJkv58_0),.din(w_dff_A_2rpz6Gtd8_0),.clk(gclk));
	jdff dff_A_ZLLxJkv58_0(.dout(w_dff_A_Yf09qgEI9_0),.din(w_dff_A_ZLLxJkv58_0),.clk(gclk));
	jdff dff_A_Yf09qgEI9_0(.dout(w_dff_A_LtbDNfuw2_0),.din(w_dff_A_Yf09qgEI9_0),.clk(gclk));
	jdff dff_A_LtbDNfuw2_0(.dout(w_dff_A_bPWhjKrN9_0),.din(w_dff_A_LtbDNfuw2_0),.clk(gclk));
	jdff dff_A_bPWhjKrN9_0(.dout(w_dff_A_UhhShjdn2_0),.din(w_dff_A_bPWhjKrN9_0),.clk(gclk));
	jdff dff_A_UhhShjdn2_0(.dout(w_dff_A_YASDx3W27_0),.din(w_dff_A_UhhShjdn2_0),.clk(gclk));
	jdff dff_A_YASDx3W27_0(.dout(w_dff_A_o26qZyEt8_0),.din(w_dff_A_YASDx3W27_0),.clk(gclk));
	jdff dff_A_o26qZyEt8_0(.dout(w_dff_A_tPu3aBsV1_0),.din(w_dff_A_o26qZyEt8_0),.clk(gclk));
	jdff dff_A_tPu3aBsV1_0(.dout(w_dff_A_njIE0DK75_0),.din(w_dff_A_tPu3aBsV1_0),.clk(gclk));
	jdff dff_A_njIE0DK75_0(.dout(w_dff_A_3H0m2vnj9_0),.din(w_dff_A_njIE0DK75_0),.clk(gclk));
	jdff dff_A_3H0m2vnj9_0(.dout(w_dff_A_EDknwrmB1_0),.din(w_dff_A_3H0m2vnj9_0),.clk(gclk));
	jdff dff_A_EDknwrmB1_0(.dout(w_dff_A_U7VvD8Jc2_0),.din(w_dff_A_EDknwrmB1_0),.clk(gclk));
	jdff dff_A_U7VvD8Jc2_0(.dout(G391gat),.din(w_dff_A_U7VvD8Jc2_0),.clk(gclk));
	jdff dff_A_9uEusv4s6_2(.dout(w_dff_A_TFLZaW9g7_0),.din(w_dff_A_9uEusv4s6_2),.clk(gclk));
	jdff dff_A_TFLZaW9g7_0(.dout(w_dff_A_za17e4i92_0),.din(w_dff_A_TFLZaW9g7_0),.clk(gclk));
	jdff dff_A_za17e4i92_0(.dout(w_dff_A_79NOVBLH2_0),.din(w_dff_A_za17e4i92_0),.clk(gclk));
	jdff dff_A_79NOVBLH2_0(.dout(w_dff_A_dnI1umAM1_0),.din(w_dff_A_79NOVBLH2_0),.clk(gclk));
	jdff dff_A_dnI1umAM1_0(.dout(w_dff_A_IWLYgiZ98_0),.din(w_dff_A_dnI1umAM1_0),.clk(gclk));
	jdff dff_A_IWLYgiZ98_0(.dout(w_dff_A_CxcAPjgn3_0),.din(w_dff_A_IWLYgiZ98_0),.clk(gclk));
	jdff dff_A_CxcAPjgn3_0(.dout(w_dff_A_gSzj3tVD3_0),.din(w_dff_A_CxcAPjgn3_0),.clk(gclk));
	jdff dff_A_gSzj3tVD3_0(.dout(w_dff_A_mLO9Rlle0_0),.din(w_dff_A_gSzj3tVD3_0),.clk(gclk));
	jdff dff_A_mLO9Rlle0_0(.dout(w_dff_A_urBtdoC78_0),.din(w_dff_A_mLO9Rlle0_0),.clk(gclk));
	jdff dff_A_urBtdoC78_0(.dout(w_dff_A_oGNZ1BnE3_0),.din(w_dff_A_urBtdoC78_0),.clk(gclk));
	jdff dff_A_oGNZ1BnE3_0(.dout(w_dff_A_BcXW1JCM7_0),.din(w_dff_A_oGNZ1BnE3_0),.clk(gclk));
	jdff dff_A_BcXW1JCM7_0(.dout(w_dff_A_eyi3NToG8_0),.din(w_dff_A_BcXW1JCM7_0),.clk(gclk));
	jdff dff_A_eyi3NToG8_0(.dout(w_dff_A_7y8vWWbu7_0),.din(w_dff_A_eyi3NToG8_0),.clk(gclk));
	jdff dff_A_7y8vWWbu7_0(.dout(w_dff_A_DPDstFdz3_0),.din(w_dff_A_7y8vWWbu7_0),.clk(gclk));
	jdff dff_A_DPDstFdz3_0(.dout(w_dff_A_kph5iynj7_0),.din(w_dff_A_DPDstFdz3_0),.clk(gclk));
	jdff dff_A_kph5iynj7_0(.dout(w_dff_A_xHuqdW4u4_0),.din(w_dff_A_kph5iynj7_0),.clk(gclk));
	jdff dff_A_xHuqdW4u4_0(.dout(w_dff_A_l4n1jSio7_0),.din(w_dff_A_xHuqdW4u4_0),.clk(gclk));
	jdff dff_A_l4n1jSio7_0(.dout(w_dff_A_9Z9W60q11_0),.din(w_dff_A_l4n1jSio7_0),.clk(gclk));
	jdff dff_A_9Z9W60q11_0(.dout(w_dff_A_OITfyRiK1_0),.din(w_dff_A_9Z9W60q11_0),.clk(gclk));
	jdff dff_A_OITfyRiK1_0(.dout(w_dff_A_mzda089A1_0),.din(w_dff_A_OITfyRiK1_0),.clk(gclk));
	jdff dff_A_mzda089A1_0(.dout(w_dff_A_WEcZ2iW12_0),.din(w_dff_A_mzda089A1_0),.clk(gclk));
	jdff dff_A_WEcZ2iW12_0(.dout(w_dff_A_fWvJ53HN4_0),.din(w_dff_A_WEcZ2iW12_0),.clk(gclk));
	jdff dff_A_fWvJ53HN4_0(.dout(w_dff_A_HMXV228V9_0),.din(w_dff_A_fWvJ53HN4_0),.clk(gclk));
	jdff dff_A_HMXV228V9_0(.dout(w_dff_A_5GFHkcEq5_0),.din(w_dff_A_HMXV228V9_0),.clk(gclk));
	jdff dff_A_5GFHkcEq5_0(.dout(G418gat),.din(w_dff_A_5GFHkcEq5_0),.clk(gclk));
	jdff dff_A_Pjx5uvvz8_2(.dout(w_dff_A_kNXwVVQk5_0),.din(w_dff_A_Pjx5uvvz8_2),.clk(gclk));
	jdff dff_A_kNXwVVQk5_0(.dout(w_dff_A_Hxt8a4OA8_0),.din(w_dff_A_kNXwVVQk5_0),.clk(gclk));
	jdff dff_A_Hxt8a4OA8_0(.dout(w_dff_A_v6VoS3YZ6_0),.din(w_dff_A_Hxt8a4OA8_0),.clk(gclk));
	jdff dff_A_v6VoS3YZ6_0(.dout(w_dff_A_6jjTL19g2_0),.din(w_dff_A_v6VoS3YZ6_0),.clk(gclk));
	jdff dff_A_6jjTL19g2_0(.dout(w_dff_A_9NcwBcff5_0),.din(w_dff_A_6jjTL19g2_0),.clk(gclk));
	jdff dff_A_9NcwBcff5_0(.dout(w_dff_A_qXcqqucO9_0),.din(w_dff_A_9NcwBcff5_0),.clk(gclk));
	jdff dff_A_qXcqqucO9_0(.dout(w_dff_A_bfsNheRL0_0),.din(w_dff_A_qXcqqucO9_0),.clk(gclk));
	jdff dff_A_bfsNheRL0_0(.dout(w_dff_A_2TS8YV1G2_0),.din(w_dff_A_bfsNheRL0_0),.clk(gclk));
	jdff dff_A_2TS8YV1G2_0(.dout(w_dff_A_P2jtaxxK0_0),.din(w_dff_A_2TS8YV1G2_0),.clk(gclk));
	jdff dff_A_P2jtaxxK0_0(.dout(w_dff_A_Opu76JVi5_0),.din(w_dff_A_P2jtaxxK0_0),.clk(gclk));
	jdff dff_A_Opu76JVi5_0(.dout(w_dff_A_7kR1rqoC4_0),.din(w_dff_A_Opu76JVi5_0),.clk(gclk));
	jdff dff_A_7kR1rqoC4_0(.dout(w_dff_A_xChkfXOo9_0),.din(w_dff_A_7kR1rqoC4_0),.clk(gclk));
	jdff dff_A_xChkfXOo9_0(.dout(w_dff_A_CJ41juEX8_0),.din(w_dff_A_xChkfXOo9_0),.clk(gclk));
	jdff dff_A_CJ41juEX8_0(.dout(w_dff_A_gH9byscB2_0),.din(w_dff_A_CJ41juEX8_0),.clk(gclk));
	jdff dff_A_gH9byscB2_0(.dout(w_dff_A_wcao1Hsz5_0),.din(w_dff_A_gH9byscB2_0),.clk(gclk));
	jdff dff_A_wcao1Hsz5_0(.dout(w_dff_A_rB6i93TA9_0),.din(w_dff_A_wcao1Hsz5_0),.clk(gclk));
	jdff dff_A_rB6i93TA9_0(.dout(w_dff_A_CNjFLDeT7_0),.din(w_dff_A_rB6i93TA9_0),.clk(gclk));
	jdff dff_A_CNjFLDeT7_0(.dout(w_dff_A_CZDy6jk95_0),.din(w_dff_A_CNjFLDeT7_0),.clk(gclk));
	jdff dff_A_CZDy6jk95_0(.dout(w_dff_A_eU16c4oW0_0),.din(w_dff_A_CZDy6jk95_0),.clk(gclk));
	jdff dff_A_eU16c4oW0_0(.dout(w_dff_A_d03moyHC8_0),.din(w_dff_A_eU16c4oW0_0),.clk(gclk));
	jdff dff_A_d03moyHC8_0(.dout(w_dff_A_jP557fHe5_0),.din(w_dff_A_d03moyHC8_0),.clk(gclk));
	jdff dff_A_jP557fHe5_0(.dout(w_dff_A_IfH9F0ig3_0),.din(w_dff_A_jP557fHe5_0),.clk(gclk));
	jdff dff_A_IfH9F0ig3_0(.dout(G419gat),.din(w_dff_A_IfH9F0ig3_0),.clk(gclk));
	jdff dff_A_tn1EyM9i3_2(.dout(w_dff_A_2jhrJeQb9_0),.din(w_dff_A_tn1EyM9i3_2),.clk(gclk));
	jdff dff_A_2jhrJeQb9_0(.dout(w_dff_A_hdL1ACui3_0),.din(w_dff_A_2jhrJeQb9_0),.clk(gclk));
	jdff dff_A_hdL1ACui3_0(.dout(w_dff_A_7cAUZ44P4_0),.din(w_dff_A_hdL1ACui3_0),.clk(gclk));
	jdff dff_A_7cAUZ44P4_0(.dout(w_dff_A_8u62kS8E6_0),.din(w_dff_A_7cAUZ44P4_0),.clk(gclk));
	jdff dff_A_8u62kS8E6_0(.dout(w_dff_A_iOSMhwi01_0),.din(w_dff_A_8u62kS8E6_0),.clk(gclk));
	jdff dff_A_iOSMhwi01_0(.dout(w_dff_A_wOn50Mqd4_0),.din(w_dff_A_iOSMhwi01_0),.clk(gclk));
	jdff dff_A_wOn50Mqd4_0(.dout(w_dff_A_RNp7315i2_0),.din(w_dff_A_wOn50Mqd4_0),.clk(gclk));
	jdff dff_A_RNp7315i2_0(.dout(w_dff_A_7P2Ns1h92_0),.din(w_dff_A_RNp7315i2_0),.clk(gclk));
	jdff dff_A_7P2Ns1h92_0(.dout(w_dff_A_yboWpnap3_0),.din(w_dff_A_7P2Ns1h92_0),.clk(gclk));
	jdff dff_A_yboWpnap3_0(.dout(w_dff_A_ok0x16gL1_0),.din(w_dff_A_yboWpnap3_0),.clk(gclk));
	jdff dff_A_ok0x16gL1_0(.dout(w_dff_A_paKelJtN5_0),.din(w_dff_A_ok0x16gL1_0),.clk(gclk));
	jdff dff_A_paKelJtN5_0(.dout(w_dff_A_4i6WhpPq2_0),.din(w_dff_A_paKelJtN5_0),.clk(gclk));
	jdff dff_A_4i6WhpPq2_0(.dout(w_dff_A_cJka9j9i7_0),.din(w_dff_A_4i6WhpPq2_0),.clk(gclk));
	jdff dff_A_cJka9j9i7_0(.dout(w_dff_A_HiTtZQB10_0),.din(w_dff_A_cJka9j9i7_0),.clk(gclk));
	jdff dff_A_HiTtZQB10_0(.dout(w_dff_A_iCbNs5643_0),.din(w_dff_A_HiTtZQB10_0),.clk(gclk));
	jdff dff_A_iCbNs5643_0(.dout(w_dff_A_YVZP8Hit7_0),.din(w_dff_A_iCbNs5643_0),.clk(gclk));
	jdff dff_A_YVZP8Hit7_0(.dout(w_dff_A_dnCHc4FG7_0),.din(w_dff_A_YVZP8Hit7_0),.clk(gclk));
	jdff dff_A_dnCHc4FG7_0(.dout(w_dff_A_X7ha8v5G5_0),.din(w_dff_A_dnCHc4FG7_0),.clk(gclk));
	jdff dff_A_X7ha8v5G5_0(.dout(w_dff_A_wLlaiJpM4_0),.din(w_dff_A_X7ha8v5G5_0),.clk(gclk));
	jdff dff_A_wLlaiJpM4_0(.dout(w_dff_A_v75tMy0o0_0),.din(w_dff_A_wLlaiJpM4_0),.clk(gclk));
	jdff dff_A_v75tMy0o0_0(.dout(w_dff_A_3vbDz3c77_0),.din(w_dff_A_v75tMy0o0_0),.clk(gclk));
	jdff dff_A_3vbDz3c77_0(.dout(w_dff_A_twN5M79m5_0),.din(w_dff_A_3vbDz3c77_0),.clk(gclk));
	jdff dff_A_twN5M79m5_0(.dout(w_dff_A_61AsB52f5_0),.din(w_dff_A_twN5M79m5_0),.clk(gclk));
	jdff dff_A_61AsB52f5_0(.dout(w_dff_A_tKl0CTRg3_0),.din(w_dff_A_61AsB52f5_0),.clk(gclk));
	jdff dff_A_tKl0CTRg3_0(.dout(G420gat),.din(w_dff_A_tKl0CTRg3_0),.clk(gclk));
	jdff dff_A_WVLP6Vxk8_2(.dout(w_dff_A_PWgPFtjU2_0),.din(w_dff_A_WVLP6Vxk8_2),.clk(gclk));
	jdff dff_A_PWgPFtjU2_0(.dout(w_dff_A_uMzpYxq58_0),.din(w_dff_A_PWgPFtjU2_0),.clk(gclk));
	jdff dff_A_uMzpYxq58_0(.dout(w_dff_A_3fyKWzI73_0),.din(w_dff_A_uMzpYxq58_0),.clk(gclk));
	jdff dff_A_3fyKWzI73_0(.dout(w_dff_A_AdPmfEQb9_0),.din(w_dff_A_3fyKWzI73_0),.clk(gclk));
	jdff dff_A_AdPmfEQb9_0(.dout(w_dff_A_2wN7WGGz8_0),.din(w_dff_A_AdPmfEQb9_0),.clk(gclk));
	jdff dff_A_2wN7WGGz8_0(.dout(w_dff_A_zo38pquS9_0),.din(w_dff_A_2wN7WGGz8_0),.clk(gclk));
	jdff dff_A_zo38pquS9_0(.dout(w_dff_A_xaHe7qAy0_0),.din(w_dff_A_zo38pquS9_0),.clk(gclk));
	jdff dff_A_xaHe7qAy0_0(.dout(w_dff_A_seNgpSMG8_0),.din(w_dff_A_xaHe7qAy0_0),.clk(gclk));
	jdff dff_A_seNgpSMG8_0(.dout(w_dff_A_DkpRyY655_0),.din(w_dff_A_seNgpSMG8_0),.clk(gclk));
	jdff dff_A_DkpRyY655_0(.dout(w_dff_A_93sfPJ2V6_0),.din(w_dff_A_DkpRyY655_0),.clk(gclk));
	jdff dff_A_93sfPJ2V6_0(.dout(w_dff_A_rRBfyQMw1_0),.din(w_dff_A_93sfPJ2V6_0),.clk(gclk));
	jdff dff_A_rRBfyQMw1_0(.dout(w_dff_A_F0ncmQOy0_0),.din(w_dff_A_rRBfyQMw1_0),.clk(gclk));
	jdff dff_A_F0ncmQOy0_0(.dout(w_dff_A_p6Xv2Vj36_0),.din(w_dff_A_F0ncmQOy0_0),.clk(gclk));
	jdff dff_A_p6Xv2Vj36_0(.dout(w_dff_A_roSWSQVY7_0),.din(w_dff_A_p6Xv2Vj36_0),.clk(gclk));
	jdff dff_A_roSWSQVY7_0(.dout(w_dff_A_3fhK9Hho3_0),.din(w_dff_A_roSWSQVY7_0),.clk(gclk));
	jdff dff_A_3fhK9Hho3_0(.dout(w_dff_A_38EjjIEu3_0),.din(w_dff_A_3fhK9Hho3_0),.clk(gclk));
	jdff dff_A_38EjjIEu3_0(.dout(w_dff_A_nDeH3VAR4_0),.din(w_dff_A_38EjjIEu3_0),.clk(gclk));
	jdff dff_A_nDeH3VAR4_0(.dout(w_dff_A_OAwbyRkb3_0),.din(w_dff_A_nDeH3VAR4_0),.clk(gclk));
	jdff dff_A_OAwbyRkb3_0(.dout(w_dff_A_crCyPbkk3_0),.din(w_dff_A_OAwbyRkb3_0),.clk(gclk));
	jdff dff_A_crCyPbkk3_0(.dout(w_dff_A_td5plFan6_0),.din(w_dff_A_crCyPbkk3_0),.clk(gclk));
	jdff dff_A_td5plFan6_0(.dout(w_dff_A_2mxWfBNh4_0),.din(w_dff_A_td5plFan6_0),.clk(gclk));
	jdff dff_A_2mxWfBNh4_0(.dout(w_dff_A_lXlBCIey5_0),.din(w_dff_A_2mxWfBNh4_0),.clk(gclk));
	jdff dff_A_lXlBCIey5_0(.dout(w_dff_A_Yj8tPGme5_0),.din(w_dff_A_lXlBCIey5_0),.clk(gclk));
	jdff dff_A_Yj8tPGme5_0(.dout(w_dff_A_RghVUsn29_0),.din(w_dff_A_Yj8tPGme5_0),.clk(gclk));
	jdff dff_A_RghVUsn29_0(.dout(G421gat),.din(w_dff_A_RghVUsn29_0),.clk(gclk));
	jdff dff_A_f3B3tmMs4_2(.dout(w_dff_A_3vO6cYus4_0),.din(w_dff_A_f3B3tmMs4_2),.clk(gclk));
	jdff dff_A_3vO6cYus4_0(.dout(w_dff_A_f4jjXWyO5_0),.din(w_dff_A_3vO6cYus4_0),.clk(gclk));
	jdff dff_A_f4jjXWyO5_0(.dout(w_dff_A_zseyeVDx1_0),.din(w_dff_A_f4jjXWyO5_0),.clk(gclk));
	jdff dff_A_zseyeVDx1_0(.dout(w_dff_A_rSMSIBmD0_0),.din(w_dff_A_zseyeVDx1_0),.clk(gclk));
	jdff dff_A_rSMSIBmD0_0(.dout(w_dff_A_hYlZPvfI3_0),.din(w_dff_A_rSMSIBmD0_0),.clk(gclk));
	jdff dff_A_hYlZPvfI3_0(.dout(w_dff_A_3qK4F6kU9_0),.din(w_dff_A_hYlZPvfI3_0),.clk(gclk));
	jdff dff_A_3qK4F6kU9_0(.dout(w_dff_A_varSMzUI0_0),.din(w_dff_A_3qK4F6kU9_0),.clk(gclk));
	jdff dff_A_varSMzUI0_0(.dout(w_dff_A_lAkQP9w03_0),.din(w_dff_A_varSMzUI0_0),.clk(gclk));
	jdff dff_A_lAkQP9w03_0(.dout(w_dff_A_nAITM0H65_0),.din(w_dff_A_lAkQP9w03_0),.clk(gclk));
	jdff dff_A_nAITM0H65_0(.dout(w_dff_A_53GLPONo1_0),.din(w_dff_A_nAITM0H65_0),.clk(gclk));
	jdff dff_A_53GLPONo1_0(.dout(w_dff_A_OxOrGcbc3_0),.din(w_dff_A_53GLPONo1_0),.clk(gclk));
	jdff dff_A_OxOrGcbc3_0(.dout(w_dff_A_HFFcodYn2_0),.din(w_dff_A_OxOrGcbc3_0),.clk(gclk));
	jdff dff_A_HFFcodYn2_0(.dout(w_dff_A_d3XfeB2A4_0),.din(w_dff_A_HFFcodYn2_0),.clk(gclk));
	jdff dff_A_d3XfeB2A4_0(.dout(w_dff_A_WXqRxgAq9_0),.din(w_dff_A_d3XfeB2A4_0),.clk(gclk));
	jdff dff_A_WXqRxgAq9_0(.dout(w_dff_A_TAlcihmq7_0),.din(w_dff_A_WXqRxgAq9_0),.clk(gclk));
	jdff dff_A_TAlcihmq7_0(.dout(w_dff_A_PDajkseE6_0),.din(w_dff_A_TAlcihmq7_0),.clk(gclk));
	jdff dff_A_PDajkseE6_0(.dout(w_dff_A_xR2ntWuf3_0),.din(w_dff_A_PDajkseE6_0),.clk(gclk));
	jdff dff_A_xR2ntWuf3_0(.dout(w_dff_A_Ot6ZQt8L0_0),.din(w_dff_A_xR2ntWuf3_0),.clk(gclk));
	jdff dff_A_Ot6ZQt8L0_0(.dout(w_dff_A_cCjI2IwX6_0),.din(w_dff_A_Ot6ZQt8L0_0),.clk(gclk));
	jdff dff_A_cCjI2IwX6_0(.dout(w_dff_A_DlHsNY8J4_0),.din(w_dff_A_cCjI2IwX6_0),.clk(gclk));
	jdff dff_A_DlHsNY8J4_0(.dout(w_dff_A_kXFTkjuy4_0),.din(w_dff_A_DlHsNY8J4_0),.clk(gclk));
	jdff dff_A_kXFTkjuy4_0(.dout(w_dff_A_YNeUI7727_0),.din(w_dff_A_kXFTkjuy4_0),.clk(gclk));
	jdff dff_A_YNeUI7727_0(.dout(w_dff_A_M1qiqP2D8_0),.din(w_dff_A_YNeUI7727_0),.clk(gclk));
	jdff dff_A_M1qiqP2D8_0(.dout(w_dff_A_zpcNDc227_0),.din(w_dff_A_M1qiqP2D8_0),.clk(gclk));
	jdff dff_A_zpcNDc227_0(.dout(G422gat),.din(w_dff_A_zpcNDc227_0),.clk(gclk));
	jdff dff_A_zLSryDsq1_2(.dout(w_dff_A_X9BNpIy34_0),.din(w_dff_A_zLSryDsq1_2),.clk(gclk));
	jdff dff_A_X9BNpIy34_0(.dout(w_dff_A_ggggMBR32_0),.din(w_dff_A_X9BNpIy34_0),.clk(gclk));
	jdff dff_A_ggggMBR32_0(.dout(w_dff_A_SAoG3qgB6_0),.din(w_dff_A_ggggMBR32_0),.clk(gclk));
	jdff dff_A_SAoG3qgB6_0(.dout(w_dff_A_1nbfXsTM0_0),.din(w_dff_A_SAoG3qgB6_0),.clk(gclk));
	jdff dff_A_1nbfXsTM0_0(.dout(w_dff_A_0XY46UUv1_0),.din(w_dff_A_1nbfXsTM0_0),.clk(gclk));
	jdff dff_A_0XY46UUv1_0(.dout(w_dff_A_GphiGjuU7_0),.din(w_dff_A_0XY46UUv1_0),.clk(gclk));
	jdff dff_A_GphiGjuU7_0(.dout(w_dff_A_r6okzc7v7_0),.din(w_dff_A_GphiGjuU7_0),.clk(gclk));
	jdff dff_A_r6okzc7v7_0(.dout(w_dff_A_jMTnckTl7_0),.din(w_dff_A_r6okzc7v7_0),.clk(gclk));
	jdff dff_A_jMTnckTl7_0(.dout(w_dff_A_Yp44VbbJ0_0),.din(w_dff_A_jMTnckTl7_0),.clk(gclk));
	jdff dff_A_Yp44VbbJ0_0(.dout(w_dff_A_F3RrdjPz0_0),.din(w_dff_A_Yp44VbbJ0_0),.clk(gclk));
	jdff dff_A_F3RrdjPz0_0(.dout(w_dff_A_Kk9XY2NS7_0),.din(w_dff_A_F3RrdjPz0_0),.clk(gclk));
	jdff dff_A_Kk9XY2NS7_0(.dout(w_dff_A_dqJDGKUL5_0),.din(w_dff_A_Kk9XY2NS7_0),.clk(gclk));
	jdff dff_A_dqJDGKUL5_0(.dout(w_dff_A_qvca6MJE9_0),.din(w_dff_A_dqJDGKUL5_0),.clk(gclk));
	jdff dff_A_qvca6MJE9_0(.dout(w_dff_A_hFrwHAby2_0),.din(w_dff_A_qvca6MJE9_0),.clk(gclk));
	jdff dff_A_hFrwHAby2_0(.dout(w_dff_A_9ia8pK5b7_0),.din(w_dff_A_hFrwHAby2_0),.clk(gclk));
	jdff dff_A_9ia8pK5b7_0(.dout(w_dff_A_f66Zlgwn4_0),.din(w_dff_A_9ia8pK5b7_0),.clk(gclk));
	jdff dff_A_f66Zlgwn4_0(.dout(w_dff_A_L8Iev85q9_0),.din(w_dff_A_f66Zlgwn4_0),.clk(gclk));
	jdff dff_A_L8Iev85q9_0(.dout(w_dff_A_W9kaoHXd6_0),.din(w_dff_A_L8Iev85q9_0),.clk(gclk));
	jdff dff_A_W9kaoHXd6_0(.dout(w_dff_A_e1IPzIUv1_0),.din(w_dff_A_W9kaoHXd6_0),.clk(gclk));
	jdff dff_A_e1IPzIUv1_0(.dout(w_dff_A_QvYRI3Qy8_0),.din(w_dff_A_e1IPzIUv1_0),.clk(gclk));
	jdff dff_A_QvYRI3Qy8_0(.dout(w_dff_A_4TCN0c4I8_0),.din(w_dff_A_QvYRI3Qy8_0),.clk(gclk));
	jdff dff_A_4TCN0c4I8_0(.dout(w_dff_A_p17Oa3ES5_0),.din(w_dff_A_4TCN0c4I8_0),.clk(gclk));
	jdff dff_A_p17Oa3ES5_0(.dout(w_dff_A_9OczA3Qo7_0),.din(w_dff_A_p17Oa3ES5_0),.clk(gclk));
	jdff dff_A_9OczA3Qo7_0(.dout(w_dff_A_MNV2tNp50_0),.din(w_dff_A_9OczA3Qo7_0),.clk(gclk));
	jdff dff_A_MNV2tNp50_0(.dout(w_dff_A_ztAzJqOG4_0),.din(w_dff_A_MNV2tNp50_0),.clk(gclk));
	jdff dff_A_ztAzJqOG4_0(.dout(G423gat),.din(w_dff_A_ztAzJqOG4_0),.clk(gclk));
	jdff dff_A_eJuXV8JT9_2(.dout(w_dff_A_NLYbL3sp8_0),.din(w_dff_A_eJuXV8JT9_2),.clk(gclk));
	jdff dff_A_NLYbL3sp8_0(.dout(w_dff_A_mecAV2dE2_0),.din(w_dff_A_NLYbL3sp8_0),.clk(gclk));
	jdff dff_A_mecAV2dE2_0(.dout(w_dff_A_OspmI1xt8_0),.din(w_dff_A_mecAV2dE2_0),.clk(gclk));
	jdff dff_A_OspmI1xt8_0(.dout(w_dff_A_Kueb2dXJ4_0),.din(w_dff_A_OspmI1xt8_0),.clk(gclk));
	jdff dff_A_Kueb2dXJ4_0(.dout(w_dff_A_MMf1I3c55_0),.din(w_dff_A_Kueb2dXJ4_0),.clk(gclk));
	jdff dff_A_MMf1I3c55_0(.dout(w_dff_A_LoDKSHCH3_0),.din(w_dff_A_MMf1I3c55_0),.clk(gclk));
	jdff dff_A_LoDKSHCH3_0(.dout(w_dff_A_9EmlGL5Z7_0),.din(w_dff_A_LoDKSHCH3_0),.clk(gclk));
	jdff dff_A_9EmlGL5Z7_0(.dout(w_dff_A_xICStOLo1_0),.din(w_dff_A_9EmlGL5Z7_0),.clk(gclk));
	jdff dff_A_xICStOLo1_0(.dout(w_dff_A_a4CYGuR08_0),.din(w_dff_A_xICStOLo1_0),.clk(gclk));
	jdff dff_A_a4CYGuR08_0(.dout(w_dff_A_mBriqa6r7_0),.din(w_dff_A_a4CYGuR08_0),.clk(gclk));
	jdff dff_A_mBriqa6r7_0(.dout(w_dff_A_XSw3uw2i4_0),.din(w_dff_A_mBriqa6r7_0),.clk(gclk));
	jdff dff_A_XSw3uw2i4_0(.dout(w_dff_A_25QxoFKl7_0),.din(w_dff_A_XSw3uw2i4_0),.clk(gclk));
	jdff dff_A_25QxoFKl7_0(.dout(w_dff_A_Tcvo3xgU1_0),.din(w_dff_A_25QxoFKl7_0),.clk(gclk));
	jdff dff_A_Tcvo3xgU1_0(.dout(w_dff_A_ncoFE3At2_0),.din(w_dff_A_Tcvo3xgU1_0),.clk(gclk));
	jdff dff_A_ncoFE3At2_0(.dout(w_dff_A_LKN1qEfb6_0),.din(w_dff_A_ncoFE3At2_0),.clk(gclk));
	jdff dff_A_LKN1qEfb6_0(.dout(w_dff_A_VvNGi9QZ6_0),.din(w_dff_A_LKN1qEfb6_0),.clk(gclk));
	jdff dff_A_VvNGi9QZ6_0(.dout(w_dff_A_5905t9GQ3_0),.din(w_dff_A_VvNGi9QZ6_0),.clk(gclk));
	jdff dff_A_5905t9GQ3_0(.dout(w_dff_A_hgghZ0xo4_0),.din(w_dff_A_5905t9GQ3_0),.clk(gclk));
	jdff dff_A_hgghZ0xo4_0(.dout(w_dff_A_JgolRGYL7_0),.din(w_dff_A_hgghZ0xo4_0),.clk(gclk));
	jdff dff_A_JgolRGYL7_0(.dout(w_dff_A_Kg3BixOI0_0),.din(w_dff_A_JgolRGYL7_0),.clk(gclk));
	jdff dff_A_Kg3BixOI0_0(.dout(w_dff_A_3LzS4Le53_0),.din(w_dff_A_Kg3BixOI0_0),.clk(gclk));
	jdff dff_A_3LzS4Le53_0(.dout(w_dff_A_JNC0STpk8_0),.din(w_dff_A_3LzS4Le53_0),.clk(gclk));
	jdff dff_A_JNC0STpk8_0(.dout(G446gat),.din(w_dff_A_JNC0STpk8_0),.clk(gclk));
	jdff dff_A_okknghdw6_1(.dout(w_dff_A_BbMXuhmh8_0),.din(w_dff_A_okknghdw6_1),.clk(gclk));
	jdff dff_A_BbMXuhmh8_0(.dout(w_dff_A_PlmPaojf1_0),.din(w_dff_A_BbMXuhmh8_0),.clk(gclk));
	jdff dff_A_PlmPaojf1_0(.dout(w_dff_A_xmbYEDkx2_0),.din(w_dff_A_PlmPaojf1_0),.clk(gclk));
	jdff dff_A_xmbYEDkx2_0(.dout(w_dff_A_eOA6Pwj32_0),.din(w_dff_A_xmbYEDkx2_0),.clk(gclk));
	jdff dff_A_eOA6Pwj32_0(.dout(w_dff_A_glXFxzKQ9_0),.din(w_dff_A_eOA6Pwj32_0),.clk(gclk));
	jdff dff_A_glXFxzKQ9_0(.dout(w_dff_A_RZ6mZWeL9_0),.din(w_dff_A_glXFxzKQ9_0),.clk(gclk));
	jdff dff_A_RZ6mZWeL9_0(.dout(w_dff_A_ZYHfgCxj7_0),.din(w_dff_A_RZ6mZWeL9_0),.clk(gclk));
	jdff dff_A_ZYHfgCxj7_0(.dout(w_dff_A_qS7pJICS4_0),.din(w_dff_A_ZYHfgCxj7_0),.clk(gclk));
	jdff dff_A_qS7pJICS4_0(.dout(w_dff_A_HEItSyrG1_0),.din(w_dff_A_qS7pJICS4_0),.clk(gclk));
	jdff dff_A_HEItSyrG1_0(.dout(w_dff_A_WSWvwix68_0),.din(w_dff_A_HEItSyrG1_0),.clk(gclk));
	jdff dff_A_WSWvwix68_0(.dout(w_dff_A_TXcrylQe7_0),.din(w_dff_A_WSWvwix68_0),.clk(gclk));
	jdff dff_A_TXcrylQe7_0(.dout(w_dff_A_zciIJX5T0_0),.din(w_dff_A_TXcrylQe7_0),.clk(gclk));
	jdff dff_A_zciIJX5T0_0(.dout(w_dff_A_eMkvwg2O6_0),.din(w_dff_A_zciIJX5T0_0),.clk(gclk));
	jdff dff_A_eMkvwg2O6_0(.dout(w_dff_A_Tre5AUZR5_0),.din(w_dff_A_eMkvwg2O6_0),.clk(gclk));
	jdff dff_A_Tre5AUZR5_0(.dout(w_dff_A_2LlgYQZT8_0),.din(w_dff_A_Tre5AUZR5_0),.clk(gclk));
	jdff dff_A_2LlgYQZT8_0(.dout(w_dff_A_LK2iKSf28_0),.din(w_dff_A_2LlgYQZT8_0),.clk(gclk));
	jdff dff_A_LK2iKSf28_0(.dout(w_dff_A_MJJPlJeh2_0),.din(w_dff_A_LK2iKSf28_0),.clk(gclk));
	jdff dff_A_MJJPlJeh2_0(.dout(w_dff_A_VaY9n6zX4_0),.din(w_dff_A_MJJPlJeh2_0),.clk(gclk));
	jdff dff_A_VaY9n6zX4_0(.dout(w_dff_A_0wgGH0mP9_0),.din(w_dff_A_VaY9n6zX4_0),.clk(gclk));
	jdff dff_A_0wgGH0mP9_0(.dout(w_dff_A_heyu5tkl4_0),.din(w_dff_A_0wgGH0mP9_0),.clk(gclk));
	jdff dff_A_heyu5tkl4_0(.dout(w_dff_A_DIc8uGqI6_0),.din(w_dff_A_heyu5tkl4_0),.clk(gclk));
	jdff dff_A_DIc8uGqI6_0(.dout(w_dff_A_TJ3o8bmC6_0),.din(w_dff_A_DIc8uGqI6_0),.clk(gclk));
	jdff dff_A_TJ3o8bmC6_0(.dout(w_dff_A_auIwklQa2_0),.din(w_dff_A_TJ3o8bmC6_0),.clk(gclk));
	jdff dff_A_auIwklQa2_0(.dout(w_dff_A_MyMSigOS3_0),.din(w_dff_A_auIwklQa2_0),.clk(gclk));
	jdff dff_A_MyMSigOS3_0(.dout(w_dff_A_JPpWur601_0),.din(w_dff_A_MyMSigOS3_0),.clk(gclk));
	jdff dff_A_JPpWur601_0(.dout(G447gat),.din(w_dff_A_JPpWur601_0),.clk(gclk));
	jdff dff_A_SKkp85xP3_2(.dout(w_dff_A_cc31PMoT9_0),.din(w_dff_A_SKkp85xP3_2),.clk(gclk));
	jdff dff_A_cc31PMoT9_0(.dout(w_dff_A_9GZ1hK3I0_0),.din(w_dff_A_cc31PMoT9_0),.clk(gclk));
	jdff dff_A_9GZ1hK3I0_0(.dout(w_dff_A_4RkgZDEY2_0),.din(w_dff_A_9GZ1hK3I0_0),.clk(gclk));
	jdff dff_A_4RkgZDEY2_0(.dout(w_dff_A_zDnCm8nu0_0),.din(w_dff_A_4RkgZDEY2_0),.clk(gclk));
	jdff dff_A_zDnCm8nu0_0(.dout(w_dff_A_ISbHSzu51_0),.din(w_dff_A_zDnCm8nu0_0),.clk(gclk));
	jdff dff_A_ISbHSzu51_0(.dout(w_dff_A_zM8TL5qy7_0),.din(w_dff_A_ISbHSzu51_0),.clk(gclk));
	jdff dff_A_zM8TL5qy7_0(.dout(w_dff_A_NbgrN2uM2_0),.din(w_dff_A_zM8TL5qy7_0),.clk(gclk));
	jdff dff_A_NbgrN2uM2_0(.dout(w_dff_A_oWrModiM8_0),.din(w_dff_A_NbgrN2uM2_0),.clk(gclk));
	jdff dff_A_oWrModiM8_0(.dout(w_dff_A_zj0JWWbJ9_0),.din(w_dff_A_oWrModiM8_0),.clk(gclk));
	jdff dff_A_zj0JWWbJ9_0(.dout(w_dff_A_wpwEF8NO8_0),.din(w_dff_A_zj0JWWbJ9_0),.clk(gclk));
	jdff dff_A_wpwEF8NO8_0(.dout(w_dff_A_Zgrdx8975_0),.din(w_dff_A_wpwEF8NO8_0),.clk(gclk));
	jdff dff_A_Zgrdx8975_0(.dout(w_dff_A_uJSpuao87_0),.din(w_dff_A_Zgrdx8975_0),.clk(gclk));
	jdff dff_A_uJSpuao87_0(.dout(w_dff_A_W6OqyxXw8_0),.din(w_dff_A_uJSpuao87_0),.clk(gclk));
	jdff dff_A_W6OqyxXw8_0(.dout(w_dff_A_oxz5g3aZ4_0),.din(w_dff_A_W6OqyxXw8_0),.clk(gclk));
	jdff dff_A_oxz5g3aZ4_0(.dout(w_dff_A_sk6ExhNv7_0),.din(w_dff_A_oxz5g3aZ4_0),.clk(gclk));
	jdff dff_A_sk6ExhNv7_0(.dout(w_dff_A_2hSo6UjF9_0),.din(w_dff_A_sk6ExhNv7_0),.clk(gclk));
	jdff dff_A_2hSo6UjF9_0(.dout(w_dff_A_gslfoMKd5_0),.din(w_dff_A_2hSo6UjF9_0),.clk(gclk));
	jdff dff_A_gslfoMKd5_0(.dout(w_dff_A_YbN9g6Lz3_0),.din(w_dff_A_gslfoMKd5_0),.clk(gclk));
	jdff dff_A_YbN9g6Lz3_0(.dout(w_dff_A_lyd6BDC26_0),.din(w_dff_A_YbN9g6Lz3_0),.clk(gclk));
	jdff dff_A_lyd6BDC26_0(.dout(w_dff_A_Cy9RN5Ea9_0),.din(w_dff_A_lyd6BDC26_0),.clk(gclk));
	jdff dff_A_Cy9RN5Ea9_0(.dout(w_dff_A_4acUKDlH8_0),.din(w_dff_A_Cy9RN5Ea9_0),.clk(gclk));
	jdff dff_A_4acUKDlH8_0(.dout(w_dff_A_xPmhi39g0_0),.din(w_dff_A_4acUKDlH8_0),.clk(gclk));
	jdff dff_A_xPmhi39g0_0(.dout(G448gat),.din(w_dff_A_xPmhi39g0_0),.clk(gclk));
	jdff dff_A_35oqKIZp5_2(.dout(w_dff_A_iaTm8Ie48_0),.din(w_dff_A_35oqKIZp5_2),.clk(gclk));
	jdff dff_A_iaTm8Ie48_0(.dout(w_dff_A_BkKoa1Aj0_0),.din(w_dff_A_iaTm8Ie48_0),.clk(gclk));
	jdff dff_A_BkKoa1Aj0_0(.dout(w_dff_A_ncJ6leYY4_0),.din(w_dff_A_BkKoa1Aj0_0),.clk(gclk));
	jdff dff_A_ncJ6leYY4_0(.dout(w_dff_A_yRCu0ZN53_0),.din(w_dff_A_ncJ6leYY4_0),.clk(gclk));
	jdff dff_A_yRCu0ZN53_0(.dout(w_dff_A_86ZZKC897_0),.din(w_dff_A_yRCu0ZN53_0),.clk(gclk));
	jdff dff_A_86ZZKC897_0(.dout(w_dff_A_9yLVeOEW4_0),.din(w_dff_A_86ZZKC897_0),.clk(gclk));
	jdff dff_A_9yLVeOEW4_0(.dout(w_dff_A_NoBSmdu83_0),.din(w_dff_A_9yLVeOEW4_0),.clk(gclk));
	jdff dff_A_NoBSmdu83_0(.dout(w_dff_A_EQv6kdJ69_0),.din(w_dff_A_NoBSmdu83_0),.clk(gclk));
	jdff dff_A_EQv6kdJ69_0(.dout(w_dff_A_49GhB9GP3_0),.din(w_dff_A_EQv6kdJ69_0),.clk(gclk));
	jdff dff_A_49GhB9GP3_0(.dout(w_dff_A_NejYa9Hm4_0),.din(w_dff_A_49GhB9GP3_0),.clk(gclk));
	jdff dff_A_NejYa9Hm4_0(.dout(w_dff_A_mwi356Ei5_0),.din(w_dff_A_NejYa9Hm4_0),.clk(gclk));
	jdff dff_A_mwi356Ei5_0(.dout(w_dff_A_4UK8dmLU4_0),.din(w_dff_A_mwi356Ei5_0),.clk(gclk));
	jdff dff_A_4UK8dmLU4_0(.dout(w_dff_A_YjvQG4Vb9_0),.din(w_dff_A_4UK8dmLU4_0),.clk(gclk));
	jdff dff_A_YjvQG4Vb9_0(.dout(w_dff_A_xMjtTQtq5_0),.din(w_dff_A_YjvQG4Vb9_0),.clk(gclk));
	jdff dff_A_xMjtTQtq5_0(.dout(w_dff_A_xZBRDJea5_0),.din(w_dff_A_xMjtTQtq5_0),.clk(gclk));
	jdff dff_A_xZBRDJea5_0(.dout(w_dff_A_8VmaL1QW4_0),.din(w_dff_A_xZBRDJea5_0),.clk(gclk));
	jdff dff_A_8VmaL1QW4_0(.dout(w_dff_A_aLy163v86_0),.din(w_dff_A_8VmaL1QW4_0),.clk(gclk));
	jdff dff_A_aLy163v86_0(.dout(w_dff_A_JLpcIygJ6_0),.din(w_dff_A_aLy163v86_0),.clk(gclk));
	jdff dff_A_JLpcIygJ6_0(.dout(w_dff_A_JRNZfyNX8_0),.din(w_dff_A_JLpcIygJ6_0),.clk(gclk));
	jdff dff_A_JRNZfyNX8_0(.dout(w_dff_A_DUn2SYoX2_0),.din(w_dff_A_JRNZfyNX8_0),.clk(gclk));
	jdff dff_A_DUn2SYoX2_0(.dout(w_dff_A_SVIyMXnD0_0),.din(w_dff_A_DUn2SYoX2_0),.clk(gclk));
	jdff dff_A_SVIyMXnD0_0(.dout(w_dff_A_wMOjNUqD0_0),.din(w_dff_A_SVIyMXnD0_0),.clk(gclk));
	jdff dff_A_wMOjNUqD0_0(.dout(G449gat),.din(w_dff_A_wMOjNUqD0_0),.clk(gclk));
	jdff dff_A_XzrLJwvU7_2(.dout(w_dff_A_WGsUVzCW5_0),.din(w_dff_A_XzrLJwvU7_2),.clk(gclk));
	jdff dff_A_WGsUVzCW5_0(.dout(w_dff_A_f5vfj9Lo2_0),.din(w_dff_A_WGsUVzCW5_0),.clk(gclk));
	jdff dff_A_f5vfj9Lo2_0(.dout(w_dff_A_GjJAyAxn3_0),.din(w_dff_A_f5vfj9Lo2_0),.clk(gclk));
	jdff dff_A_GjJAyAxn3_0(.dout(w_dff_A_zf5aOjMK3_0),.din(w_dff_A_GjJAyAxn3_0),.clk(gclk));
	jdff dff_A_zf5aOjMK3_0(.dout(w_dff_A_fdnWkuQj8_0),.din(w_dff_A_zf5aOjMK3_0),.clk(gclk));
	jdff dff_A_fdnWkuQj8_0(.dout(w_dff_A_Vhcm3Vsi0_0),.din(w_dff_A_fdnWkuQj8_0),.clk(gclk));
	jdff dff_A_Vhcm3Vsi0_0(.dout(w_dff_A_xDrrMfif8_0),.din(w_dff_A_Vhcm3Vsi0_0),.clk(gclk));
	jdff dff_A_xDrrMfif8_0(.dout(w_dff_A_n8DNWQXD0_0),.din(w_dff_A_xDrrMfif8_0),.clk(gclk));
	jdff dff_A_n8DNWQXD0_0(.dout(w_dff_A_1PIGjyax6_0),.din(w_dff_A_n8DNWQXD0_0),.clk(gclk));
	jdff dff_A_1PIGjyax6_0(.dout(w_dff_A_U4tjKopR2_0),.din(w_dff_A_1PIGjyax6_0),.clk(gclk));
	jdff dff_A_U4tjKopR2_0(.dout(w_dff_A_uPnkL4H75_0),.din(w_dff_A_U4tjKopR2_0),.clk(gclk));
	jdff dff_A_uPnkL4H75_0(.dout(w_dff_A_fRe3ziQ83_0),.din(w_dff_A_uPnkL4H75_0),.clk(gclk));
	jdff dff_A_fRe3ziQ83_0(.dout(w_dff_A_nXQt28No0_0),.din(w_dff_A_fRe3ziQ83_0),.clk(gclk));
	jdff dff_A_nXQt28No0_0(.dout(w_dff_A_MR4rYd8Y2_0),.din(w_dff_A_nXQt28No0_0),.clk(gclk));
	jdff dff_A_MR4rYd8Y2_0(.dout(w_dff_A_57kI9jKK2_0),.din(w_dff_A_MR4rYd8Y2_0),.clk(gclk));
	jdff dff_A_57kI9jKK2_0(.dout(w_dff_A_LJz7AEag5_0),.din(w_dff_A_57kI9jKK2_0),.clk(gclk));
	jdff dff_A_LJz7AEag5_0(.dout(w_dff_A_H1u2yFCu8_0),.din(w_dff_A_LJz7AEag5_0),.clk(gclk));
	jdff dff_A_H1u2yFCu8_0(.dout(w_dff_A_hEiuQsy60_0),.din(w_dff_A_H1u2yFCu8_0),.clk(gclk));
	jdff dff_A_hEiuQsy60_0(.dout(w_dff_A_Jp7BKBcE8_0),.din(w_dff_A_hEiuQsy60_0),.clk(gclk));
	jdff dff_A_Jp7BKBcE8_0(.dout(w_dff_A_JO5z6CfR0_0),.din(w_dff_A_Jp7BKBcE8_0),.clk(gclk));
	jdff dff_A_JO5z6CfR0_0(.dout(w_dff_A_cjQoounO9_0),.din(w_dff_A_JO5z6CfR0_0),.clk(gclk));
	jdff dff_A_cjQoounO9_0(.dout(w_dff_A_nwMOwfqC9_0),.din(w_dff_A_cjQoounO9_0),.clk(gclk));
	jdff dff_A_nwMOwfqC9_0(.dout(w_dff_A_AVNYSklC9_0),.din(w_dff_A_nwMOwfqC9_0),.clk(gclk));
	jdff dff_A_AVNYSklC9_0(.dout(w_dff_A_QCDFiWI29_0),.din(w_dff_A_AVNYSklC9_0),.clk(gclk));
	jdff dff_A_QCDFiWI29_0(.dout(w_dff_A_0PMn0hJB0_0),.din(w_dff_A_QCDFiWI29_0),.clk(gclk));
	jdff dff_A_0PMn0hJB0_0(.dout(G450gat),.din(w_dff_A_0PMn0hJB0_0),.clk(gclk));
	jdff dff_A_GfrfYs7c3_2(.dout(w_dff_A_bOVUXuoD0_0),.din(w_dff_A_GfrfYs7c3_2),.clk(gclk));
	jdff dff_A_bOVUXuoD0_0(.dout(w_dff_A_Tt5IM3gC2_0),.din(w_dff_A_bOVUXuoD0_0),.clk(gclk));
	jdff dff_A_Tt5IM3gC2_0(.dout(w_dff_A_vJllNvW37_0),.din(w_dff_A_Tt5IM3gC2_0),.clk(gclk));
	jdff dff_A_vJllNvW37_0(.dout(w_dff_A_anvMCwWk5_0),.din(w_dff_A_vJllNvW37_0),.clk(gclk));
	jdff dff_A_anvMCwWk5_0(.dout(w_dff_A_9ZpPBmDb3_0),.din(w_dff_A_anvMCwWk5_0),.clk(gclk));
	jdff dff_A_9ZpPBmDb3_0(.dout(w_dff_A_T13WJN8i9_0),.din(w_dff_A_9ZpPBmDb3_0),.clk(gclk));
	jdff dff_A_T13WJN8i9_0(.dout(w_dff_A_eB7DEgd49_0),.din(w_dff_A_T13WJN8i9_0),.clk(gclk));
	jdff dff_A_eB7DEgd49_0(.dout(w_dff_A_AS7pQGWR3_0),.din(w_dff_A_eB7DEgd49_0),.clk(gclk));
	jdff dff_A_AS7pQGWR3_0(.dout(w_dff_A_LyhT3Z584_0),.din(w_dff_A_AS7pQGWR3_0),.clk(gclk));
	jdff dff_A_LyhT3Z584_0(.dout(w_dff_A_6omjgayz8_0),.din(w_dff_A_LyhT3Z584_0),.clk(gclk));
	jdff dff_A_6omjgayz8_0(.dout(w_dff_A_bwdaUsn80_0),.din(w_dff_A_6omjgayz8_0),.clk(gclk));
	jdff dff_A_bwdaUsn80_0(.dout(w_dff_A_YdgMZpal5_0),.din(w_dff_A_bwdaUsn80_0),.clk(gclk));
	jdff dff_A_YdgMZpal5_0(.dout(w_dff_A_6I9W7B382_0),.din(w_dff_A_YdgMZpal5_0),.clk(gclk));
	jdff dff_A_6I9W7B382_0(.dout(w_dff_A_lF7573D76_0),.din(w_dff_A_6I9W7B382_0),.clk(gclk));
	jdff dff_A_lF7573D76_0(.dout(w_dff_A_HKn00WHx4_0),.din(w_dff_A_lF7573D76_0),.clk(gclk));
	jdff dff_A_HKn00WHx4_0(.dout(w_dff_A_Ki16IQvh5_0),.din(w_dff_A_HKn00WHx4_0),.clk(gclk));
	jdff dff_A_Ki16IQvh5_0(.dout(w_dff_A_Os2j3Xf64_0),.din(w_dff_A_Ki16IQvh5_0),.clk(gclk));
	jdff dff_A_Os2j3Xf64_0(.dout(w_dff_A_kjS6n2Tj3_0),.din(w_dff_A_Os2j3Xf64_0),.clk(gclk));
	jdff dff_A_kjS6n2Tj3_0(.dout(w_dff_A_OvIHAtGE4_0),.din(w_dff_A_kjS6n2Tj3_0),.clk(gclk));
	jdff dff_A_OvIHAtGE4_0(.dout(w_dff_A_6DChSZZH1_0),.din(w_dff_A_OvIHAtGE4_0),.clk(gclk));
	jdff dff_A_6DChSZZH1_0(.dout(w_dff_A_z77Qdrzb2_0),.din(w_dff_A_6DChSZZH1_0),.clk(gclk));
	jdff dff_A_z77Qdrzb2_0(.dout(w_dff_A_tNGgaUHW5_0),.din(w_dff_A_z77Qdrzb2_0),.clk(gclk));
	jdff dff_A_tNGgaUHW5_0(.dout(w_dff_A_aqqygrba0_0),.din(w_dff_A_tNGgaUHW5_0),.clk(gclk));
	jdff dff_A_aqqygrba0_0(.dout(G767gat),.din(w_dff_A_aqqygrba0_0),.clk(gclk));
	jdff dff_A_V2xBhqVi9_2(.dout(w_dff_A_UhEno39s5_0),.din(w_dff_A_V2xBhqVi9_2),.clk(gclk));
	jdff dff_A_UhEno39s5_0(.dout(w_dff_A_H6ADwYna4_0),.din(w_dff_A_UhEno39s5_0),.clk(gclk));
	jdff dff_A_H6ADwYna4_0(.dout(w_dff_A_UcMitI1C7_0),.din(w_dff_A_H6ADwYna4_0),.clk(gclk));
	jdff dff_A_UcMitI1C7_0(.dout(w_dff_A_aSVkd4Ff7_0),.din(w_dff_A_UcMitI1C7_0),.clk(gclk));
	jdff dff_A_aSVkd4Ff7_0(.dout(w_dff_A_1oP9gFMZ7_0),.din(w_dff_A_aSVkd4Ff7_0),.clk(gclk));
	jdff dff_A_1oP9gFMZ7_0(.dout(w_dff_A_OLmp3Pkl3_0),.din(w_dff_A_1oP9gFMZ7_0),.clk(gclk));
	jdff dff_A_OLmp3Pkl3_0(.dout(w_dff_A_cRGSIDc77_0),.din(w_dff_A_OLmp3Pkl3_0),.clk(gclk));
	jdff dff_A_cRGSIDc77_0(.dout(w_dff_A_k0rs1XpL1_0),.din(w_dff_A_cRGSIDc77_0),.clk(gclk));
	jdff dff_A_k0rs1XpL1_0(.dout(w_dff_A_08Ksdl6U1_0),.din(w_dff_A_k0rs1XpL1_0),.clk(gclk));
	jdff dff_A_08Ksdl6U1_0(.dout(w_dff_A_5DBO5nBd9_0),.din(w_dff_A_08Ksdl6U1_0),.clk(gclk));
	jdff dff_A_5DBO5nBd9_0(.dout(w_dff_A_GnLSMS6k0_0),.din(w_dff_A_5DBO5nBd9_0),.clk(gclk));
	jdff dff_A_GnLSMS6k0_0(.dout(w_dff_A_YSOOJHDj7_0),.din(w_dff_A_GnLSMS6k0_0),.clk(gclk));
	jdff dff_A_YSOOJHDj7_0(.dout(w_dff_A_PqsA697P7_0),.din(w_dff_A_YSOOJHDj7_0),.clk(gclk));
	jdff dff_A_PqsA697P7_0(.dout(w_dff_A_u0ogulA74_0),.din(w_dff_A_PqsA697P7_0),.clk(gclk));
	jdff dff_A_u0ogulA74_0(.dout(w_dff_A_lJjyH7pR1_0),.din(w_dff_A_u0ogulA74_0),.clk(gclk));
	jdff dff_A_lJjyH7pR1_0(.dout(w_dff_A_GB8OJbKW5_0),.din(w_dff_A_lJjyH7pR1_0),.clk(gclk));
	jdff dff_A_GB8OJbKW5_0(.dout(w_dff_A_0VkPOqun0_0),.din(w_dff_A_GB8OJbKW5_0),.clk(gclk));
	jdff dff_A_0VkPOqun0_0(.dout(w_dff_A_rTlckvfX8_0),.din(w_dff_A_0VkPOqun0_0),.clk(gclk));
	jdff dff_A_rTlckvfX8_0(.dout(w_dff_A_yJLFYMXo8_0),.din(w_dff_A_rTlckvfX8_0),.clk(gclk));
	jdff dff_A_yJLFYMXo8_0(.dout(w_dff_A_W0LjnJ1Y3_0),.din(w_dff_A_yJLFYMXo8_0),.clk(gclk));
	jdff dff_A_W0LjnJ1Y3_0(.dout(w_dff_A_K9AScd5x5_0),.din(w_dff_A_W0LjnJ1Y3_0),.clk(gclk));
	jdff dff_A_K9AScd5x5_0(.dout(w_dff_A_PdT8HLSw6_0),.din(w_dff_A_K9AScd5x5_0),.clk(gclk));
	jdff dff_A_PdT8HLSw6_0(.dout(w_dff_A_rMOKO8Va0_0),.din(w_dff_A_PdT8HLSw6_0),.clk(gclk));
	jdff dff_A_rMOKO8Va0_0(.dout(G768gat),.din(w_dff_A_rMOKO8Va0_0),.clk(gclk));
	jdff dff_A_mActxA1q1_2(.dout(w_dff_A_mpNryBtD7_0),.din(w_dff_A_mActxA1q1_2),.clk(gclk));
	jdff dff_A_mpNryBtD7_0(.dout(w_dff_A_lRTd2kHq2_0),.din(w_dff_A_mpNryBtD7_0),.clk(gclk));
	jdff dff_A_lRTd2kHq2_0(.dout(w_dff_A_RO5XnqGe0_0),.din(w_dff_A_lRTd2kHq2_0),.clk(gclk));
	jdff dff_A_RO5XnqGe0_0(.dout(w_dff_A_ja5ECaDl7_0),.din(w_dff_A_RO5XnqGe0_0),.clk(gclk));
	jdff dff_A_ja5ECaDl7_0(.dout(w_dff_A_RujbHO2T6_0),.din(w_dff_A_ja5ECaDl7_0),.clk(gclk));
	jdff dff_A_RujbHO2T6_0(.dout(w_dff_A_9MvXUAwN6_0),.din(w_dff_A_RujbHO2T6_0),.clk(gclk));
	jdff dff_A_9MvXUAwN6_0(.dout(w_dff_A_ObNNLjWz3_0),.din(w_dff_A_9MvXUAwN6_0),.clk(gclk));
	jdff dff_A_ObNNLjWz3_0(.dout(w_dff_A_Q85dHfFR8_0),.din(w_dff_A_ObNNLjWz3_0),.clk(gclk));
	jdff dff_A_Q85dHfFR8_0(.dout(w_dff_A_CJ7l9IIl9_0),.din(w_dff_A_Q85dHfFR8_0),.clk(gclk));
	jdff dff_A_CJ7l9IIl9_0(.dout(w_dff_A_vJ2mjGAW2_0),.din(w_dff_A_CJ7l9IIl9_0),.clk(gclk));
	jdff dff_A_vJ2mjGAW2_0(.dout(w_dff_A_EqBCNLti8_0),.din(w_dff_A_vJ2mjGAW2_0),.clk(gclk));
	jdff dff_A_EqBCNLti8_0(.dout(w_dff_A_3bWZAoto9_0),.din(w_dff_A_EqBCNLti8_0),.clk(gclk));
	jdff dff_A_3bWZAoto9_0(.dout(G850gat),.din(w_dff_A_3bWZAoto9_0),.clk(gclk));
	jdff dff_A_60dQ0vME0_2(.dout(w_dff_A_FxINdpY90_0),.din(w_dff_A_60dQ0vME0_2),.clk(gclk));
	jdff dff_A_FxINdpY90_0(.dout(w_dff_A_LAPyEJzi7_0),.din(w_dff_A_FxINdpY90_0),.clk(gclk));
	jdff dff_A_LAPyEJzi7_0(.dout(w_dff_A_cFpF1vaT8_0),.din(w_dff_A_LAPyEJzi7_0),.clk(gclk));
	jdff dff_A_cFpF1vaT8_0(.dout(w_dff_A_PigixGgt4_0),.din(w_dff_A_cFpF1vaT8_0),.clk(gclk));
	jdff dff_A_PigixGgt4_0(.dout(w_dff_A_3WOGSuKH6_0),.din(w_dff_A_PigixGgt4_0),.clk(gclk));
	jdff dff_A_3WOGSuKH6_0(.dout(w_dff_A_Tk06FzEK8_0),.din(w_dff_A_3WOGSuKH6_0),.clk(gclk));
	jdff dff_A_Tk06FzEK8_0(.dout(w_dff_A_mQZdZmLF8_0),.din(w_dff_A_Tk06FzEK8_0),.clk(gclk));
	jdff dff_A_mQZdZmLF8_0(.dout(G863gat),.din(w_dff_A_mQZdZmLF8_0),.clk(gclk));
	jdff dff_A_wy9iCPNA8_2(.dout(w_dff_A_CR6Atpxz3_0),.din(w_dff_A_wy9iCPNA8_2),.clk(gclk));
	jdff dff_A_CR6Atpxz3_0(.dout(w_dff_A_aiGWq3Ct5_0),.din(w_dff_A_CR6Atpxz3_0),.clk(gclk));
	jdff dff_A_aiGWq3Ct5_0(.dout(w_dff_A_5AvoXO3C0_0),.din(w_dff_A_aiGWq3Ct5_0),.clk(gclk));
	jdff dff_A_5AvoXO3C0_0(.dout(w_dff_A_Jekc0ell4_0),.din(w_dff_A_5AvoXO3C0_0),.clk(gclk));
	jdff dff_A_Jekc0ell4_0(.dout(w_dff_A_EGaa7CQv5_0),.din(w_dff_A_Jekc0ell4_0),.clk(gclk));
	jdff dff_A_EGaa7CQv5_0(.dout(w_dff_A_GkhGHBf64_0),.din(w_dff_A_EGaa7CQv5_0),.clk(gclk));
	jdff dff_A_GkhGHBf64_0(.dout(w_dff_A_DtDmt0P51_0),.din(w_dff_A_GkhGHBf64_0),.clk(gclk));
	jdff dff_A_DtDmt0P51_0(.dout(w_dff_A_JMvGVQtW8_0),.din(w_dff_A_DtDmt0P51_0),.clk(gclk));
	jdff dff_A_JMvGVQtW8_0(.dout(w_dff_A_F0uIHKDW3_0),.din(w_dff_A_JMvGVQtW8_0),.clk(gclk));
	jdff dff_A_F0uIHKDW3_0(.dout(G864gat),.din(w_dff_A_F0uIHKDW3_0),.clk(gclk));
	jdff dff_A_Sdrq4YvS9_2(.dout(w_dff_A_o1bfOnu03_0),.din(w_dff_A_Sdrq4YvS9_2),.clk(gclk));
	jdff dff_A_o1bfOnu03_0(.dout(w_dff_A_PwAQE4pJ6_0),.din(w_dff_A_o1bfOnu03_0),.clk(gclk));
	jdff dff_A_PwAQE4pJ6_0(.dout(w_dff_A_nNYK5rPu9_0),.din(w_dff_A_PwAQE4pJ6_0),.clk(gclk));
	jdff dff_A_nNYK5rPu9_0(.dout(w_dff_A_b6zPkQoE0_0),.din(w_dff_A_nNYK5rPu9_0),.clk(gclk));
	jdff dff_A_b6zPkQoE0_0(.dout(w_dff_A_gyIhbuSH0_0),.din(w_dff_A_b6zPkQoE0_0),.clk(gclk));
	jdff dff_A_gyIhbuSH0_0(.dout(w_dff_A_sM8YiyDE4_0),.din(w_dff_A_gyIhbuSH0_0),.clk(gclk));
	jdff dff_A_sM8YiyDE4_0(.dout(w_dff_A_viukNfvi6_0),.din(w_dff_A_sM8YiyDE4_0),.clk(gclk));
	jdff dff_A_viukNfvi6_0(.dout(w_dff_A_N3sOEtk88_0),.din(w_dff_A_viukNfvi6_0),.clk(gclk));
	jdff dff_A_N3sOEtk88_0(.dout(w_dff_A_k2mXTqrK8_0),.din(w_dff_A_N3sOEtk88_0),.clk(gclk));
	jdff dff_A_k2mXTqrK8_0(.dout(w_dff_A_3DTwPGHW6_0),.din(w_dff_A_k2mXTqrK8_0),.clk(gclk));
	jdff dff_A_3DTwPGHW6_0(.dout(w_dff_A_mZEP9Xyo0_0),.din(w_dff_A_3DTwPGHW6_0),.clk(gclk));
	jdff dff_A_mZEP9Xyo0_0(.dout(G865gat),.din(w_dff_A_mZEP9Xyo0_0),.clk(gclk));
	jdff dff_A_qYIxtJuD1_2(.dout(w_dff_A_o4YoZEAw8_0),.din(w_dff_A_qYIxtJuD1_2),.clk(gclk));
	jdff dff_A_o4YoZEAw8_0(.dout(G866gat),.din(w_dff_A_o4YoZEAw8_0),.clk(gclk));
	jdff dff_A_gyc3Cwpg3_2(.dout(w_dff_A_ZsT733M38_0),.din(w_dff_A_gyc3Cwpg3_2),.clk(gclk));
	jdff dff_A_ZsT733M38_0(.dout(w_dff_A_0IjuXLnU4_0),.din(w_dff_A_ZsT733M38_0),.clk(gclk));
	jdff dff_A_0IjuXLnU4_0(.dout(w_dff_A_02VidGkE4_0),.din(w_dff_A_0IjuXLnU4_0),.clk(gclk));
	jdff dff_A_02VidGkE4_0(.dout(w_dff_A_8ipjTEtQ4_0),.din(w_dff_A_02VidGkE4_0),.clk(gclk));
	jdff dff_A_8ipjTEtQ4_0(.dout(G874gat),.din(w_dff_A_8ipjTEtQ4_0),.clk(gclk));
	jdff dff_A_OP8VKc2T4_2(.dout(w_dff_A_ntucOagn6_0),.din(w_dff_A_OP8VKc2T4_2),.clk(gclk));
	jdff dff_A_ntucOagn6_0(.dout(G879gat),.din(w_dff_A_ntucOagn6_0),.clk(gclk));
	jdff dff_A_Ddccxeqd0_2(.dout(w_dff_A_FnkDKaHR4_0),.din(w_dff_A_Ddccxeqd0_2),.clk(gclk));
	jdff dff_A_FnkDKaHR4_0(.dout(w_dff_A_8gLXGBeE6_0),.din(w_dff_A_FnkDKaHR4_0),.clk(gclk));
	jdff dff_A_8gLXGBeE6_0(.dout(w_dff_A_rk1Nj5926_0),.din(w_dff_A_8gLXGBeE6_0),.clk(gclk));
	jdff dff_A_rk1Nj5926_0(.dout(G880gat),.din(w_dff_A_rk1Nj5926_0),.clk(gclk));
endmodule

