/*

c3540:
	jxor: 52
	jspl: 225
	jspl3: 338
	jnot: 188
	jdff: 381
	jand: 525
	jor: 352

Summary:
	jxor: 52
	jspl: 225
	jspl3: 338
	jnot: 188
	jdff: 381
	jand: 525
	jor: 352

The maximum logic level gap of any gate:
	c3540: 26
*/

module gf_c3540(gclk, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402);
	input gclk;
	input G1;
	input G13;
	input G20;
	input G33;
	input G41;
	input G45;
	input G50;
	input G58;
	input G68;
	input G77;
	input G87;
	input G97;
	input G107;
	input G116;
	input G124;
	input G125;
	input G128;
	input G132;
	input G137;
	input G143;
	input G150;
	input G159;
	input G169;
	input G179;
	input G190;
	input G200;
	input G213;
	input G222;
	input G223;
	input G226;
	input G232;
	input G238;
	input G244;
	input G250;
	input G257;
	input G264;
	input G270;
	input G274;
	input G283;
	input G294;
	input G303;
	input G311;
	input G317;
	input G322;
	input G326;
	input G329;
	input G330;
	input G343;
	input G1698;
	input G2897;
	output G353;
	output G355;
	output G361;
	output G358;
	output G351;
	output G372;
	output G369;
	output G399;
	output G364;
	output G396;
	output G384;
	output G367;
	output G387;
	output G393;
	output G390;
	output G378;
	output G375;
	output G381;
	output G407;
	output G409;
	output G405;
	output G402;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[1:0] w_G1_2;
	wire[2:0] w_G13_0;
	wire[2:0] w_G13_1;
	wire[1:0] w_G13_2;
	wire[2:0] w_G20_0;
	wire[2:0] w_G20_1;
	wire[2:0] w_G20_2;
	wire[2:0] w_G20_3;
	wire[2:0] w_G20_4;
	wire[2:0] w_G20_5;
	wire[2:0] w_G20_6;
	wire[2:0] w_G33_0;
	wire[2:0] w_G33_1;
	wire[2:0] w_G33_2;
	wire[2:0] w_G33_3;
	wire[2:0] w_G33_4;
	wire[2:0] w_G33_5;
	wire[2:0] w_G33_6;
	wire[2:0] w_G33_7;
	wire[2:0] w_G33_8;
	wire[2:0] w_G33_9;
	wire[2:0] w_G33_10;
	wire[2:0] w_G33_11;
	wire[2:0] w_G33_12;
	wire[2:0] w_G41_0;
	wire[2:0] w_G45_0;
	wire[1:0] w_G45_1;
	wire[2:0] w_G50_0;
	wire[2:0] w_G50_1;
	wire[2:0] w_G50_2;
	wire[2:0] w_G50_3;
	wire[2:0] w_G50_4;
	wire[2:0] w_G50_5;
	wire[2:0] w_G58_0;
	wire[2:0] w_G58_1;
	wire[2:0] w_G58_2;
	wire[2:0] w_G58_3;
	wire[2:0] w_G58_4;
	wire[2:0] w_G58_5;
	wire[2:0] w_G68_0;
	wire[2:0] w_G68_1;
	wire[2:0] w_G68_2;
	wire[2:0] w_G68_3;
	wire[2:0] w_G68_4;
	wire[2:0] w_G68_5;
	wire[2:0] w_G77_0;
	wire[2:0] w_G77_1;
	wire[2:0] w_G77_2;
	wire[2:0] w_G77_3;
	wire[2:0] w_G77_4;
	wire[2:0] w_G87_0;
	wire[2:0] w_G87_1;
	wire[2:0] w_G87_2;
	wire[2:0] w_G87_3;
	wire[2:0] w_G97_0;
	wire[2:0] w_G97_1;
	wire[2:0] w_G97_2;
	wire[2:0] w_G97_3;
	wire[2:0] w_G97_4;
	wire[2:0] w_G107_0;
	wire[2:0] w_G107_1;
	wire[2:0] w_G107_2;
	wire[2:0] w_G107_3;
	wire[1:0] w_G107_4;
	wire[2:0] w_G116_0;
	wire[2:0] w_G116_1;
	wire[2:0] w_G116_2;
	wire[2:0] w_G116_3;
	wire[2:0] w_G116_4;
	wire[2:0] w_G116_5;
	wire[1:0] w_G125_0;
	wire[2:0] w_G128_0;
	wire[2:0] w_G132_0;
	wire[1:0] w_G132_1;
	wire[2:0] w_G137_0;
	wire[2:0] w_G137_1;
	wire[2:0] w_G143_0;
	wire[2:0] w_G143_1;
	wire[1:0] w_G143_2;
	wire[2:0] w_G150_0;
	wire[2:0] w_G150_1;
	wire[2:0] w_G150_2;
	wire[1:0] w_G150_3;
	wire[2:0] w_G159_0;
	wire[2:0] w_G159_1;
	wire[2:0] w_G159_2;
	wire[2:0] w_G159_3;
	wire[2:0] w_G169_0;
	wire[2:0] w_G169_1;
	wire[2:0] w_G169_2;
	wire[1:0] w_G169_3;
	wire[2:0] w_G179_0;
	wire[2:0] w_G179_1;
	wire[2:0] w_G179_2;
	wire[2:0] w_G190_0;
	wire[2:0] w_G190_1;
	wire[2:0] w_G190_2;
	wire[2:0] w_G190_3;
	wire[2:0] w_G190_4;
	wire[2:0] w_G200_0;
	wire[2:0] w_G200_1;
	wire[2:0] w_G200_2;
	wire[1:0] w_G200_3;
	wire[2:0] w_G213_0;
	wire[1:0] w_G223_0;
	wire[2:0] w_G226_0;
	wire[2:0] w_G226_1;
	wire[2:0] w_G232_0;
	wire[2:0] w_G232_1;
	wire[2:0] w_G238_0;
	wire[2:0] w_G244_0;
	wire[1:0] w_G244_1;
	wire[2:0] w_G250_0;
	wire[2:0] w_G257_0;
	wire[2:0] w_G257_1;
	wire[2:0] w_G264_0;
	wire[2:0] w_G270_0;
	wire[2:0] w_G274_0;
	wire[2:0] w_G283_0;
	wire[2:0] w_G283_1;
	wire[2:0] w_G283_2;
	wire[2:0] w_G283_3;
	wire[2:0] w_G294_0;
	wire[2:0] w_G294_1;
	wire[2:0] w_G294_2;
	wire[1:0] w_G294_3;
	wire[2:0] w_G303_0;
	wire[2:0] w_G303_1;
	wire[2:0] w_G303_2;
	wire[2:0] w_G311_0;
	wire[2:0] w_G311_1;
	wire[2:0] w_G317_0;
	wire[1:0] w_G317_1;
	wire[2:0] w_G322_0;
	wire[1:0] w_G326_0;
	wire[2:0] w_G330_0;
	wire[1:0] w_G343_0;
	wire[2:0] w_G1698_0;
	wire w_G355_0;
	wire G355_fa_;
	wire w_G396_0;
	wire G396_fa_;
	wire w_G384_0;
	wire G384_fa_;
	wire[2:0] w_n72_0;
	wire[2:0] w_n72_1;
	wire[2:0] w_n73_0;
	wire[2:0] w_n73_1;
	wire[2:0] w_n73_2;
	wire[2:0] w_n74_0;
	wire[2:0] w_n74_1;
	wire[1:0] w_n74_2;
	wire[2:0] w_n75_0;
	wire[2:0] w_n75_1;
	wire[1:0] w_n75_2;
	wire[1:0] w_n76_0;
	wire[1:0] w_n77_0;
	wire[2:0] w_n79_0;
	wire[2:0] w_n79_1;
	wire[2:0] w_n80_0;
	wire[2:0] w_n80_1;
	wire[2:0] w_n81_0;
	wire[2:0] w_n81_1;
	wire[1:0] w_n81_2;
	wire[2:0] w_n84_0;
	wire[2:0] w_n84_1;
	wire[1:0] w_n85_0;
	wire[2:0] w_n86_0;
	wire[1:0] w_n89_0;
	wire[2:0] w_n90_0;
	wire[2:0] w_n91_0;
	wire[2:0] w_n91_1;
	wire[2:0] w_n94_0;
	wire[2:0] w_n96_0;
	wire[2:0] w_n105_0;
	wire[1:0] w_n105_1;
	wire[2:0] w_n111_0;
	wire[1:0] w_n112_0;
	wire[2:0] w_n118_0;
	wire[1:0] w_n120_0;
	wire[1:0] w_n126_0;
	wire[1:0] w_n130_0;
	wire[1:0] w_n134_0;
	wire[1:0] w_n137_0;
	wire[2:0] w_n139_0;
	wire[2:0] w_n139_1;
	wire[1:0] w_n140_0;
	wire[2:0] w_n141_0;
	wire[2:0] w_n141_1;
	wire[2:0] w_n141_2;
	wire[1:0] w_n141_3;
	wire[2:0] w_n142_0;
	wire[2:0] w_n142_1;
	wire[1:0] w_n142_2;
	wire[1:0] w_n143_0;
	wire[2:0] w_n144_0;
	wire[2:0] w_n144_1;
	wire[1:0] w_n144_2;
	wire[2:0] w_n147_0;
	wire[1:0] w_n148_0;
	wire[2:0] w_n151_0;
	wire[2:0] w_n151_1;
	wire[2:0] w_n151_2;
	wire[2:0] w_n151_3;
	wire[2:0] w_n151_4;
	wire[2:0] w_n151_5;
	wire[1:0] w_n151_6;
	wire[2:0] w_n152_0;
	wire[2:0] w_n153_0;
	wire[2:0] w_n153_1;
	wire[2:0] w_n153_2;
	wire[2:0] w_n153_3;
	wire[2:0] w_n153_4;
	wire[2:0] w_n153_5;
	wire[2:0] w_n153_6;
	wire[2:0] w_n153_7;
	wire[1:0] w_n153_8;
	wire[2:0] w_n161_0;
	wire[2:0] w_n163_0;
	wire[1:0] w_n163_1;
	wire[2:0] w_n164_0;
	wire[1:0] w_n165_0;
	wire[1:0] w_n167_0;
	wire[2:0] w_n168_0;
	wire[2:0] w_n168_1;
	wire[2:0] w_n168_2;
	wire[2:0] w_n168_3;
	wire[2:0] w_n168_4;
	wire[1:0] w_n168_5;
	wire[1:0] w_n169_0;
	wire[2:0] w_n170_0;
	wire[2:0] w_n172_0;
	wire[2:0] w_n172_1;
	wire[2:0] w_n172_2;
	wire[2:0] w_n172_3;
	wire[2:0] w_n172_4;
	wire[2:0] w_n173_0;
	wire[2:0] w_n173_1;
	wire[2:0] w_n173_2;
	wire[1:0] w_n173_3;
	wire[1:0] w_n176_0;
	wire[2:0] w_n177_0;
	wire[2:0] w_n177_1;
	wire[2:0] w_n182_0;
	wire[1:0] w_n182_1;
	wire[2:0] w_n186_0;
	wire[2:0] w_n186_1;
	wire[2:0] w_n189_0;
	wire[2:0] w_n189_1;
	wire[2:0] w_n189_2;
	wire[1:0] w_n190_0;
	wire[2:0] w_n192_0;
	wire[2:0] w_n198_0;
	wire[2:0] w_n199_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n202_0;
	wire[2:0] w_n205_0;
	wire[1:0] w_n205_1;
	wire[1:0] w_n207_0;
	wire[2:0] w_n212_0;
	wire[1:0] w_n212_1;
	wire[1:0] w_n213_0;
	wire[1:0] w_n215_0;
	wire[1:0] w_n218_0;
	wire[2:0] w_n224_0;
	wire[1:0] w_n224_1;
	wire[1:0] w_n225_0;
	wire[1:0] w_n229_0;
	wire[2:0] w_n234_0;
	wire[1:0] w_n234_1;
	wire[2:0] w_n237_0;
	wire[1:0] w_n238_0;
	wire[2:0] w_n242_0;
	wire[1:0] w_n243_0;
	wire[1:0] w_n247_0;
	wire[1:0] w_n250_0;
	wire[1:0] w_n251_0;
	wire[2:0] w_n255_0;
	wire[1:0] w_n255_1;
	wire[1:0] w_n256_0;
	wire[1:0] w_n257_0;
	wire[1:0] w_n259_0;
	wire[1:0] w_n260_0;
	wire[2:0] w_n261_0;
	wire[2:0] w_n261_1;
	wire[2:0] w_n262_0;
	wire[1:0] w_n269_0;
	wire[1:0] w_n272_0;
	wire[2:0] w_n279_0;
	wire[1:0] w_n279_1;
	wire[1:0] w_n282_0;
	wire[1:0] w_n283_0;
	wire[2:0] w_n292_0;
	wire[1:0] w_n298_0;
	wire[2:0] w_n308_0;
	wire[2:0] w_n308_1;
	wire[1:0] w_n309_0;
	wire[1:0] w_n310_0;
	wire[1:0] w_n312_0;
	wire[1:0] w_n313_0;
	wire[2:0] w_n315_0;
	wire[1:0] w_n321_0;
	wire[2:0] w_n323_0;
	wire[2:0] w_n330_0;
	wire[1:0] w_n333_0;
	wire[1:0] w_n334_0;
	wire[1:0] w_n344_0;
	wire[1:0] w_n347_0;
	wire[1:0] w_n348_0;
	wire[1:0] w_n349_0;
	wire[1:0] w_n350_0;
	wire[1:0] w_n351_0;
	wire[2:0] w_n352_0;
	wire[1:0] w_n352_1;
	wire[2:0] w_n354_0;
	wire[1:0] w_n354_1;
	wire[1:0] w_n355_0;
	wire[2:0] w_n356_0;
	wire[1:0] w_n356_1;
	wire[1:0] w_n357_0;
	wire[2:0] w_n367_0;
	wire[1:0] w_n367_1;
	wire[1:0] w_n370_0;
	wire[1:0] w_n375_0;
	wire[1:0] w_n378_0;
	wire[2:0] w_n383_0;
	wire[2:0] w_n387_0;
	wire[2:0] w_n388_0;
	wire[2:0] w_n388_1;
	wire[1:0] w_n388_2;
	wire[1:0] w_n394_0;
	wire[1:0] w_n395_0;
	wire[2:0] w_n404_0;
	wire[1:0] w_n405_0;
	wire[1:0] w_n407_0;
	wire[2:0] w_n414_0;
	wire[2:0] w_n417_0;
	wire[1:0] w_n420_0;
	wire[1:0] w_n425_0;
	wire[1:0] w_n426_0;
	wire[1:0] w_n428_0;
	wire[1:0] w_n430_0;
	wire[1:0] w_n435_0;
	wire[2:0] w_n439_0;
	wire[1:0] w_n441_0;
	wire[1:0] w_n445_0;
	wire[1:0] w_n450_0;
	wire[1:0] w_n452_0;
	wire[1:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[1:0] w_n465_0;
	wire[1:0] w_n472_0;
	wire[1:0] w_n473_0;
	wire[2:0] w_n482_0;
	wire[1:0] w_n483_0;
	wire[1:0] w_n494_0;
	wire[1:0] w_n499_0;
	wire[1:0] w_n500_0;
	wire[2:0] w_n503_0;
	wire[2:0] w_n507_0;
	wire[2:0] w_n507_1;
	wire[1:0] w_n507_2;
	wire[1:0] w_n511_0;
	wire[1:0] w_n512_0;
	wire[2:0] w_n514_0;
	wire[1:0] w_n514_1;
	wire[1:0] w_n520_0;
	wire[1:0] w_n533_0;
	wire[1:0] w_n534_0;
	wire[1:0] w_n541_0;
	wire[1:0] w_n542_0;
	wire[1:0] w_n543_0;
	wire[1:0] w_n544_0;
	wire[1:0] w_n548_0;
	wire[1:0] w_n550_0;
	wire[1:0] w_n551_0;
	wire[1:0] w_n559_0;
	wire[1:0] w_n562_0;
	wire[2:0] w_n566_0;
	wire[1:0] w_n566_1;
	wire[2:0] w_n567_0;
	wire[2:0] w_n567_1;
	wire[2:0] w_n567_2;
	wire[2:0] w_n567_3;
	wire[2:0] w_n567_4;
	wire[1:0] w_n567_5;
	wire[1:0] w_n569_0;
	wire[1:0] w_n570_0;
	wire[2:0] w_n571_0;
	wire[2:0] w_n571_1;
	wire[1:0] w_n571_2;
	wire[2:0] w_n572_0;
	wire[1:0] w_n573_0;
	wire[1:0] w_n574_0;
	wire[2:0] w_n576_0;
	wire[1:0] w_n577_0;
	wire[2:0] w_n579_0;
	wire[1:0] w_n579_1;
	wire[2:0] w_n580_0;
	wire[1:0] w_n582_0;
	wire[1:0] w_n584_0;
	wire[1:0] w_n598_0;
	wire[2:0] w_n600_0;
	wire[2:0] w_n600_1;
	wire[2:0] w_n601_0;
	wire[1:0] w_n602_0;
	wire[2:0] w_n604_0;
	wire[2:0] w_n604_1;
	wire[2:0] w_n604_2;
	wire[2:0] w_n605_0;
	wire[2:0] w_n613_0;
	wire[2:0] w_n613_1;
	wire[2:0] w_n614_0;
	wire[2:0] w_n614_1;
	wire[2:0] w_n614_2;
	wire[2:0] w_n614_3;
	wire[2:0] w_n614_4;
	wire[1:0] w_n614_5;
	wire[2:0] w_n618_0;
	wire[2:0] w_n618_1;
	wire[1:0] w_n618_2;
	wire[2:0] w_n619_0;
	wire[2:0] w_n620_0;
	wire[1:0] w_n622_0;
	wire[1:0] w_n624_0;
	wire[2:0] w_n626_0;
	wire[1:0] w_n628_0;
	wire[2:0] w_n629_0;
	wire[2:0] w_n629_1;
	wire[2:0] w_n629_2;
	wire[2:0] w_n629_3;
	wire[2:0] w_n629_4;
	wire[1:0] w_n629_5;
	wire[1:0] w_n630_0;
	wire[1:0] w_n632_0;
	wire[2:0] w_n633_0;
	wire[2:0] w_n633_1;
	wire[2:0] w_n633_2;
	wire[2:0] w_n633_3;
	wire[2:0] w_n633_4;
	wire[2:0] w_n633_5;
	wire[1:0] w_n633_6;
	wire[1:0] w_n634_0;
	wire[1:0] w_n637_0;
	wire[2:0] w_n638_0;
	wire[2:0] w_n638_1;
	wire[2:0] w_n638_2;
	wire[2:0] w_n638_3;
	wire[2:0] w_n638_4;
	wire[2:0] w_n638_5;
	wire[2:0] w_n638_6;
	wire[1:0] w_n638_7;
	wire[2:0] w_n640_0;
	wire[2:0] w_n640_1;
	wire[2:0] w_n640_2;
	wire[2:0] w_n640_3;
	wire[2:0] w_n640_4;
	wire[2:0] w_n640_5;
	wire[2:0] w_n640_6;
	wire[1:0] w_n640_7;
	wire[2:0] w_n646_0;
	wire[2:0] w_n646_1;
	wire[2:0] w_n646_2;
	wire[2:0] w_n646_3;
	wire[2:0] w_n646_4;
	wire[2:0] w_n646_5;
	wire[2:0] w_n646_6;
	wire[1:0] w_n646_7;
	wire[2:0] w_n648_0;
	wire[2:0] w_n648_1;
	wire[2:0] w_n648_2;
	wire[2:0] w_n648_3;
	wire[1:0] w_n648_4;
	wire[1:0] w_n649_0;
	wire[1:0] w_n650_0;
	wire[2:0] w_n651_0;
	wire[2:0] w_n651_1;
	wire[2:0] w_n651_2;
	wire[2:0] w_n651_3;
	wire[2:0] w_n651_4;
	wire[2:0] w_n651_5;
	wire[2:0] w_n651_6;
	wire[1:0] w_n651_7;
	wire[2:0] w_n653_0;
	wire[2:0] w_n653_1;
	wire[2:0] w_n653_2;
	wire[2:0] w_n653_3;
	wire[2:0] w_n653_4;
	wire[2:0] w_n653_5;
	wire[2:0] w_n653_6;
	wire[1:0] w_n653_7;
	wire[2:0] w_n680_0;
	wire[2:0] w_n680_1;
	wire[2:0] w_n680_2;
	wire[2:0] w_n680_3;
	wire[1:0] w_n680_4;
	wire[1:0] w_n682_0;
	wire[2:0] w_n684_0;
	wire[1:0] w_n685_0;
	wire[2:0] w_n690_0;
	wire[1:0] w_n690_1;
	wire[1:0] w_n692_0;
	wire[2:0] w_n703_0;
	wire[1:0] w_n703_1;
	wire[1:0] w_n704_0;
	wire[1:0] w_n718_0;
	wire[1:0] w_n733_0;
	wire[2:0] w_n741_0;
	wire[1:0] w_n741_1;
	wire[1:0] w_n748_0;
	wire[1:0] w_n754_0;
	wire[1:0] w_n759_0;
	wire[1:0] w_n766_0;
	wire[2:0] w_n767_0;
	wire[1:0] w_n767_1;
	wire[2:0] w_n771_0;
	wire[1:0] w_n771_1;
	wire[1:0] w_n772_0;
	wire[1:0] w_n773_0;
	wire[1:0] w_n775_0;
	wire[1:0] w_n777_0;
	wire[1:0] w_n782_0;
	wire[1:0] w_n798_0;
	wire[2:0] w_n802_0;
	wire[1:0] w_n817_0;
	wire[1:0] w_n830_0;
	wire[1:0] w_n833_0;
	wire[2:0] w_n845_0;
	wire[1:0] w_n855_0;
	wire[1:0] w_n860_0;
	wire[1:0] w_n861_0;
	wire[2:0] w_n863_0;
	wire[2:0] w_n869_0;
	wire[1:0] w_n873_0;
	wire[1:0] w_n875_0;
	wire[1:0] w_n884_0;
	wire[1:0] w_n887_0;
	wire[2:0] w_n937_0;
	wire[1:0] w_n959_0;
	wire[2:0] w_n987_0;
	wire[2:0] w_n1029_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1036_0;
	wire[1:0] w_n1039_0;
	wire[1:0] w_n1040_0;
	wire[1:0] w_n1041_0;
	wire[1:0] w_n1043_0;
	wire[1:0] w_n1044_0;
	wire[1:0] w_n1045_0;
	wire[1:0] w_n1048_0;
	wire[2:0] w_n1053_0;
	wire[1:0] w_n1056_0;
	wire[1:0] w_n1062_0;
	wire[1:0] w_n1091_0;
	wire[2:0] w_n1114_0;
	wire[2:0] w_n1159_0;
	wire[1:0] w_n1161_0;
	wire[1:0] w_n1164_0;
	wire[1:0] w_n1168_0;
	wire[1:0] w_n1170_0;
	wire[1:0] w_n1177_0;
	wire[1:0] w_n1178_0;
	wire[1:0] w_n1179_0;
	wire[1:0] w_n1184_0;
	wire w_dff_B_xHjQUWcM6_1;
	wire w_dff_B_VjmlfsDy9_1;
	wire w_dff_B_Mt4cKI405_1;
	wire w_dff_B_HQ7X0MvH1_1;
	wire w_dff_B_22bVWtfL0_1;
	wire w_dff_B_2TT2DMn67_1;
	wire w_dff_B_QVk4dQrZ1_1;
	wire w_dff_B_oLBQvcT41_1;
	wire w_dff_B_kwkvJeIU9_1;
	wire w_dff_B_TGoVpYEx6_1;
	wire w_dff_B_Fk2wDTnf3_1;
	wire w_dff_B_5snqWQgf3_1;
	wire w_dff_B_634dszOY3_1;
	wire w_dff_B_6pWQF2Zt3_1;
	wire w_dff_B_A7SfOkGb4_1;
	wire w_dff_B_J0H42DkE9_1;
	wire w_dff_B_sccYniaQ7_1;
	wire w_dff_B_IexGRyFg3_1;
	wire w_dff_B_ueFBhWi45_1;
	wire w_dff_B_u0KPQAqv5_0;
	wire w_dff_B_2GVCeahx4_0;
	wire w_dff_B_WysWk24V4_0;
	wire w_dff_B_FOEMFtkR0_0;
	wire w_dff_B_BylPbcSb9_0;
	wire w_dff_B_SCuwsZ4y1_0;
	wire w_dff_B_UOhUKV8Q1_0;
	wire w_dff_B_urnAEHxh0_0;
	wire w_dff_B_1ST408VS9_0;
	wire w_dff_B_RDDKxhKt5_0;
	wire w_dff_B_DTkC4zXD7_0;
	wire w_dff_B_MnaE5uDC8_0;
	wire w_dff_B_VnxhVx6Z9_0;
	wire w_dff_B_Gcvpk43x2_0;
	wire w_dff_B_9oyPHs7g1_0;
	wire w_dff_B_OQBD1u0p4_0;
	wire w_dff_B_Q2OW7rOi7_0;
	wire w_dff_B_q6bNldw60_1;
	wire w_dff_B_l3lZnQLq9_1;
	wire w_dff_B_jnLKg6zc8_1;
	wire w_dff_B_YQWUqsGM8_1;
	wire w_dff_B_xqUFUO7K0_1;
	wire w_dff_B_QMLcvk0t1_1;
	wire w_dff_B_rfz4CH6Q5_1;
	wire w_dff_B_AWJ7WFQe3_1;
	wire w_dff_B_ta9doG5X1_1;
	wire w_dff_B_2aULs05t3_1;
	wire w_dff_B_1e8Tsy3Y7_1;
	wire w_dff_B_jriraDas1_1;
	wire w_dff_B_lzlWFihn9_1;
	wire w_dff_B_0solhEAT9_1;
	wire w_dff_B_JlIj0nb70_1;
	wire w_dff_B_9hCywfez2_1;
	wire w_dff_B_TpzJBJHo9_1;
	wire w_dff_B_03WS732s8_1;
	wire w_dff_B_X6R4aNGE6_1;
	wire w_dff_B_L8RNaC5U4_1;
	wire w_dff_B_81gzoYDd3_1;
	wire w_dff_B_8rdXXyPZ7_1;
	wire w_dff_B_QhvOIY9O8_1;
	wire w_dff_B_eGGmHCC48_1;
	wire w_dff_B_lXd2Awnt0_1;
	wire w_dff_B_bOsBCVpY4_1;
	wire w_dff_B_prp0mfij9_1;
	wire w_dff_B_j8FbVouI0_1;
	wire w_dff_B_mu9n9ilP0_1;
	wire w_dff_B_0ZaFb6Dc1_1;
	wire w_dff_B_c7VrnfJj6_0;
	wire w_dff_B_9zpnASnZ7_0;
	wire w_dff_B_muoYqJAP6_1;
	wire w_dff_B_zWiukuNG3_1;
	wire w_dff_B_WdUXIHfI8_1;
	wire w_dff_B_exGhWo893_1;
	wire w_dff_B_KuRzPd3r4_1;
	wire w_dff_B_jPnidbuk4_1;
	wire w_dff_B_WGNNI6Js1_1;
	wire w_dff_B_e9ZR4Lw22_1;
	wire w_dff_B_jZtfpIr95_1;
	wire w_dff_B_Ut40zb8L0_1;
	wire w_dff_B_Gedsz2kC2_1;
	wire w_dff_B_ACEyuKxm7_1;
	wire w_dff_B_6lU5nar68_1;
	wire w_dff_B_T2cfWnkw0_1;
	wire w_dff_B_IdKWaz1P7_1;
	wire w_dff_B_EtTGXOoa6_1;
	wire w_dff_B_Gb5dMDpc1_1;
	wire w_dff_B_DvcwlsgN3_1;
	wire w_dff_B_xHL8CGM99_1;
	wire w_dff_B_3uApdKyi9_1;
	wire w_dff_B_7ldL9vkR7_1;
	wire w_dff_B_yGM9w70N1_1;
	wire w_dff_B_vqt2ixL65_1;
	wire w_dff_B_SLNhhTuD3_1;
	wire w_dff_B_wCBFBJ289_1;
	wire w_dff_B_r16mdVyf5_1;
	wire w_dff_B_R0y0XQyz9_1;
	wire w_dff_B_mV3DpgdJ3_1;
	wire w_dff_B_71ZeuXyD3_1;
	wire w_dff_B_ieRAh7pn1_1;
	wire w_dff_B_jgDIuOm97_1;
	wire w_dff_B_0qLziPTL0_1;
	wire w_dff_B_KHiWN5fs7_1;
	wire w_dff_B_Kwx5Zzrv2_1;
	wire w_dff_B_BLn13hMk0_1;
	wire w_dff_B_cBrdFfoY9_1;
	wire w_dff_B_xpplfx8y9_1;
	wire w_dff_B_TpYVZ56u7_1;
	wire w_dff_B_Lk0aWGUz5_1;
	wire w_dff_B_vNB21VeQ7_1;
	wire w_dff_B_TueIlBv25_1;
	wire w_dff_B_ZHeLmu9d1_1;
	wire w_dff_B_wOe0PS6z4_1;
	wire w_dff_B_4oi2hvdW4_1;
	wire w_dff_B_DJfgBu7q6_1;
	wire w_dff_B_wJFwYcwK6_1;
	wire w_dff_B_zsuITUe04_1;
	wire w_dff_B_PgYY4vUx7_1;
	wire w_dff_B_tyELKyBq2_1;
	wire w_dff_B_ROu1pqix5_1;
	wire w_dff_B_PC9xXn8s6_1;
	wire w_dff_B_C4JZ1NsH6_1;
	wire w_dff_A_1cQEWpcD0_0;
	wire w_dff_A_nEeQ9yMU7_0;
	wire w_dff_A_BhJhL6gc7_0;
	wire w_dff_A_0bqHEcZ56_1;
	wire w_dff_A_5UrYmzix0_1;
	wire w_dff_B_lHnJ19Zu1_2;
	wire w_dff_B_HFykTtMo5_2;
	wire w_dff_B_nAxUj1iK8_1;
	wire w_dff_B_FAEdZJEp2_2;
	wire w_dff_B_tXLhldf20_2;
	wire w_dff_B_gUkXXbu39_2;
	wire w_dff_B_HpHtOqHA3_2;
	wire w_dff_B_DNikSduU6_1;
	wire w_dff_B_pETUV4B08_0;
	wire w_dff_B_CyQrIu989_0;
	wire w_dff_B_P6gvEx497_0;
	wire w_dff_B_BdB41wc63_0;
	wire w_dff_B_QI4QLR1u6_0;
	wire w_dff_A_z3QgeTlH5_0;
	wire w_dff_A_rykcEi9w2_2;
	wire w_dff_A_7tXAyvIc9_0;
	wire w_dff_A_sJ26Vx1O7_0;
	wire w_dff_A_J6sjkAqq8_0;
	wire w_dff_A_bvAV8NCD6_0;
	wire w_dff_A_78xeVvM67_0;
	wire w_dff_A_8ZrYs9dv9_0;
	wire w_dff_A_q9YlF5aK2_0;
	wire w_dff_A_aCiwPFen2_0;
	wire w_dff_A_BrII8quO0_0;
	wire w_dff_A_BNxYVpX82_0;
	wire w_dff_A_pLGlTChb9_0;
	wire w_dff_A_wlGAPGV14_0;
	wire w_dff_A_ACPekjjV3_0;
	wire w_dff_A_XW192r1e4_0;
	wire w_dff_A_Ov05VS1I6_0;
	wire w_dff_A_Ehf5bj7o1_0;
	wire w_dff_A_BCEjLeVG1_0;
	wire w_dff_A_Na8c8buW1_0;
	wire w_dff_A_9nOBslLD0_0;
	wire w_dff_A_TxiSdO7Q1_0;
	wire w_dff_A_0PKeuSai9_0;
	wire w_dff_A_vBFf419J5_0;
	wire w_dff_A_Bc4lmPKi8_0;
	wire w_dff_A_RDsEoRlQ8_0;
	wire w_dff_A_EQGyNptT1_0;
	wire w_dff_A_2ex2bB0s2_0;
	wire w_dff_A_iY0rTqRq8_1;
	wire w_dff_A_lYvf9yv19_0;
	wire w_dff_A_aAa5JjEc7_0;
	wire w_dff_A_Fhngsv7p4_0;
	wire w_dff_A_IiXeey773_0;
	wire w_dff_A_sbaw8oi15_0;
	wire w_dff_A_wCgExy7V3_0;
	wire w_dff_A_a7QWWlo49_0;
	wire w_dff_A_97MhZySN7_0;
	wire w_dff_A_fXNCu55L5_0;
	wire w_dff_A_noLTKY9K1_0;
	wire w_dff_A_s8ZpllIO5_0;
	wire w_dff_A_rRYQwDuV9_0;
	wire w_dff_A_wVhcwU9y1_0;
	wire w_dff_A_AA0t5bqS3_0;
	wire w_dff_A_x8DSkExS1_0;
	wire w_dff_A_2rCmqjTR3_0;
	wire w_dff_A_pzAxV5YN0_0;
	wire w_dff_A_1pWOxKmm2_0;
	wire w_dff_A_vXqGkER71_0;
	wire w_dff_A_74NmZsTt6_0;
	wire w_dff_A_NUL87zGZ7_0;
	wire w_dff_A_HwuPOGwD1_0;
	wire w_dff_A_VgBe6X6X6_0;
	wire w_dff_A_k0bEhgrd6_0;
	wire w_dff_A_87qaW5RV8_0;
	wire w_dff_A_oQ8HNp3w4_0;
	wire w_dff_A_n7f1N90w6_0;
	wire w_dff_A_tGv9QlUg2_2;
	wire w_dff_A_3x64q4q06_0;
	wire w_dff_A_8zTbKcVM5_0;
	wire w_dff_A_WcRpnLv47_0;
	wire w_dff_A_VWMlx0DM4_0;
	wire w_dff_A_SRswPu2g9_0;
	wire w_dff_A_dsW8gz3d1_0;
	wire w_dff_A_9nxvnyL83_0;
	wire w_dff_A_rjysqVXr3_0;
	wire w_dff_A_1MMwLd568_0;
	wire w_dff_A_mplGl4XJ4_0;
	wire w_dff_A_RBGPa3Sa1_0;
	wire w_dff_A_JJoZgGzJ0_0;
	wire w_dff_A_1ERsv94T0_0;
	wire w_dff_A_zuCevQOC5_0;
	wire w_dff_A_8uszQAbC5_0;
	wire w_dff_A_C8aYFkpA1_0;
	wire w_dff_A_nsIxJLQ78_0;
	wire w_dff_A_zXV78VOh4_0;
	wire w_dff_A_Zhpbic7e7_0;
	wire w_dff_A_WZikTYSU2_0;
	wire w_dff_A_UJ6dkv765_0;
	wire w_dff_A_iNnPeafG1_0;
	wire w_dff_A_FASwSrM37_2;
	wire w_dff_A_dces0ZHC1_0;
	wire w_dff_A_RT13c4cr8_0;
	wire w_dff_A_2TFo5LhC0_0;
	wire w_dff_A_o5jm3Mm81_0;
	wire w_dff_A_meQoZqRp6_0;
	wire w_dff_A_o0Dkscnh8_0;
	wire w_dff_A_FU0qnnH58_0;
	wire w_dff_A_YQCi2RKZ1_0;
	wire w_dff_A_1Lyz008O0_0;
	wire w_dff_A_dn3jklqc2_0;
	wire w_dff_A_IzrKkmJm6_0;
	wire w_dff_A_RgvbBbXO7_0;
	wire w_dff_A_d6UYDttH1_0;
	wire w_dff_A_q7kUgwte7_0;
	wire w_dff_A_78s6Bmiz5_0;
	wire w_dff_A_XSQYp8zp7_0;
	wire w_dff_A_XQDd9TfH3_0;
	wire w_dff_A_ORBJJzze9_0;
	wire w_dff_A_p0KFPyrp9_0;
	wire w_dff_A_2fEjbVbc3_0;
	wire w_dff_A_klDGG1qC4_0;
	wire w_dff_A_dbikGQN51_0;
	wire w_dff_A_4JGf5plu9_0;
	wire w_dff_A_mZS3SlCI8_0;
	wire w_dff_A_w2ewmxbD2_0;
	wire w_dff_A_aHt6RkCZ8_2;
	wire w_dff_A_9kbngka28_0;
	wire w_dff_A_IYTSwjoI4_0;
	wire w_dff_A_qqrfy9M99_0;
	wire w_dff_A_oaVQbbEI6_0;
	wire w_dff_A_kXgogSIG3_0;
	wire w_dff_A_WNT0POCn7_0;
	wire w_dff_A_nqoJYSNL1_0;
	wire w_dff_A_cYsBGSsA7_0;
	wire w_dff_A_B2x7IUKZ3_0;
	wire w_dff_A_8Y6CJ15X6_0;
	wire w_dff_A_dd4MIhLH5_0;
	wire w_dff_A_2mCLAEP53_0;
	wire w_dff_A_301Oya3x9_0;
	wire w_dff_A_l4Z1rTCC8_0;
	wire w_dff_A_0MT9M76Q4_0;
	wire w_dff_A_vzCd2yne5_0;
	wire w_dff_A_Md6n8JZm6_0;
	wire w_dff_A_Gzgq586f7_0;
	wire w_dff_A_TSk4U95C5_0;
	wire w_dff_A_78grfziF7_0;
	wire w_dff_A_8gwvzG3Y4_0;
	wire w_dff_A_gQ4ywcus0_0;
	wire w_dff_A_OWR7LLM93_0;
	wire w_dff_A_3yZSjYJI9_0;
	wire w_dff_A_Vf4sBJ6B5_0;
	wire w_dff_A_GiPrHPkG6_0;
	wire w_dff_A_iZwOYoxD1_2;
	wire w_dff_A_nxynkYd86_0;
	wire w_dff_A_1Yf1Nag91_0;
	wire w_dff_A_L48ZhFEL1_0;
	wire w_dff_A_V1RyywYX5_0;
	wire w_dff_A_mPPi4LPU7_0;
	wire w_dff_A_r0rYql7X9_0;
	wire w_dff_A_WbN5nSJi3_0;
	wire w_dff_A_AaYTQQIO4_0;
	wire w_dff_A_di5db3TJ7_0;
	wire w_dff_A_YExiTsD20_0;
	wire w_dff_A_GNI49PoX8_0;
	wire w_dff_A_PUvCBNmy8_0;
	wire w_dff_A_e0vPEeNW9_0;
	wire w_dff_A_UNMIhmVW3_2;
	wire w_dff_A_W573gzgN9_0;
	wire w_dff_A_NMw2Zrv26_0;
	wire w_dff_A_JjnjHTSU2_0;
	wire w_dff_A_Xxem4AfI3_0;
	wire w_dff_A_grmmOweH7_0;
	wire w_dff_A_ACA69HnV9_0;
	wire w_dff_A_wpYTuy680_0;
	wire w_dff_A_KuWfMyM55_0;
	wire w_dff_A_ivu8aHFk6_0;
	wire w_dff_A_hAuOoFWj5_0;
	wire w_dff_A_fr52rNKf2_0;
	wire w_dff_A_74kv90FR7_2;
	wire w_dff_A_cjS2pxn31_0;
	wire w_dff_A_WueOsCzZ7_0;
	wire w_dff_A_oGhCCwGG8_0;
	wire w_dff_A_OKllOvWW4_0;
	wire w_dff_A_QdQBOA8w3_0;
	wire w_dff_A_Slg7fNet9_0;
	wire w_dff_A_MqE4mDbP7_0;
	wire w_dff_A_kDZ2kY0h4_0;
	wire w_dff_A_puLJejtV0_0;
	wire w_dff_A_XdftFSS88_0;
	wire w_dff_A_pcZx37y88_0;
	wire w_dff_A_CwM31BKC3_0;
	wire w_dff_A_uNfvpnLU7_0;
	wire w_dff_A_oGQbtTGb6_2;
	wire w_dff_A_u4Y6Oiym5_0;
	wire w_dff_A_z1roqDWs3_0;
	wire w_dff_A_qTzjGlMH7_0;
	wire w_dff_A_NfmaXxh35_0;
	wire w_dff_A_TS3mP57A5_0;
	wire w_dff_A_Hn3wW3cl6_0;
	wire w_dff_A_vDJgBnJw7_0;
	wire w_dff_A_iBMZlcHm8_0;
	wire w_dff_A_OMDYSKow2_1;
	wire w_dff_A_CLoWoswO9_0;
	wire w_dff_A_1GY6J38V1_0;
	wire w_dff_A_UfW6VExg5_0;
	wire w_dff_A_ZSKi4e2b8_0;
	wire w_dff_A_3UYy6rT51_0;
	wire w_dff_A_qvaVkxqt4_0;
	wire w_dff_A_v1DjgLVT8_0;
	wire w_dff_A_x0Ej28Hs0_0;
	wire w_dff_A_CbRgsCRD0_0;
	wire w_dff_A_UjOfFQLK5_0;
	wire w_dff_A_IB1KoBEj5_0;
	wire w_dff_A_1fhjShhg7_0;
	wire w_dff_A_BIzCn8732_1;
	wire w_dff_A_NnaKXWZx5_0;
	wire w_dff_A_KyS9Hjs93_0;
	wire w_dff_A_0g3CbZTa8_0;
	wire w_dff_A_1M87rgWm2_0;
	wire w_dff_A_DErI4UT83_0;
	wire w_dff_A_VTfJQwGE2_0;
	wire w_dff_A_t0bPdXfN7_0;
	wire w_dff_A_a1Iu7cw04_2;
	wire w_dff_A_y1N5lnv53_0;
	wire w_dff_A_dVxtIZAd8_0;
	wire w_dff_A_g97xnSVg6_0;
	wire w_dff_A_C82QFasT6_0;
	wire w_dff_A_qyQ4axtJ9_0;
	wire w_dff_A_T6L90GSH9_0;
	wire w_dff_A_PSsr8Fhy0_1;
	wire w_dff_A_gudd3lGr8_0;
	wire w_dff_A_tdXo1ibK4_0;
	wire w_dff_A_wlwNzbXG0_0;
	wire w_dff_A_2O09XMK62_0;
	wire w_dff_A_Gw1BjGpo0_0;
	wire w_dff_A_6yoiM3mB4_1;
	wire w_dff_A_bHnA99PJ1_0;
	wire w_dff_A_YTjfZZFu2_0;
	wire w_dff_A_NVctI2WS2_0;
	wire w_dff_A_oDfHDQeK2_0;
	wire w_dff_A_46DSCL1y5_0;
	wire w_dff_A_jfdPnZ8C5_0;
	wire w_dff_A_6xuJbluM3_1;
	wire w_dff_A_DrYpNYYV3_0;
	wire w_dff_A_dmHlHfbC2_0;
	wire w_dff_A_ayDuw0Rr3_0;
	wire w_dff_A_dMyhEWA48_0;
	wire w_dff_A_XsSApLM01_0;
	wire w_dff_A_tByJlnk29_1;
	wire w_dff_A_5eXJgyL09_0;
	wire w_dff_A_1WDh2ufO5_0;
	wire w_dff_A_arVy5Q4o0_0;
	wire w_dff_A_F97UfJu59_1;
	wire w_dff_A_yAIUZYfb7_0;
	wire w_dff_A_bGBEGjHA2_0;
	wire w_dff_A_QYZeNjaj8_0;
	wire w_dff_A_07wqAPrM9_1;
	wire w_dff_A_2L7PwvHK6_0;
	wire w_dff_A_9uTwBV9l3_0;
	wire w_dff_A_BXTsnPBU4_0;
	wire w_dff_A_eICaxmaI2_1;
	wire w_dff_A_LcUuZJrn4_2;
	wire w_dff_A_OigxRcUw0_0;
	jnot g0000(.din(w_G77_4[2]),.dout(n72),.clk(gclk));
	jnot g0001(.din(w_G50_5[2]),.dout(n73),.clk(gclk));
	jnot g0002(.din(w_G58_5[2]),.dout(n74),.clk(gclk));
	jnot g0003(.din(w_G68_5[2]),.dout(n75),.clk(gclk));
	jand g0004(.dina(w_n75_2[1]),.dinb(w_n74_2[1]),.dout(n76),.clk(gclk));
	jand g0005(.dina(w_n76_0[1]),.dinb(w_n73_2[2]),.dout(n77),.clk(gclk));
	jand g0006(.dina(w_n77_0[1]),.dinb(w_n72_1[2]),.dout(w_dff_A_rykcEi9w2_2),.clk(gclk));
	jnot g0007(.din(w_G87_3[2]),.dout(n79),.clk(gclk));
	jnot g0008(.din(w_G97_4[2]),.dout(n80),.clk(gclk));
	jnot g0009(.din(w_G107_4[1]),.dout(n81),.clk(gclk));
	jand g0010(.dina(w_n81_2[1]),.dinb(w_n80_1[2]),.dout(n82),.clk(gclk));
	jor g0011(.dina(n82),.dinb(w_n79_1[2]),.dout(G355_fa_),.clk(gclk));
	jnot g0012(.din(w_G250_0[2]),.dout(n84),.clk(gclk));
	jnot g0013(.din(w_G257_1[2]),.dout(n85),.clk(gclk));
	jnot g0014(.din(w_G264_0[2]),.dout(n86),.clk(gclk));
	jand g0015(.dina(w_n86_0[2]),.dinb(w_n85_0[1]),.dout(n87),.clk(gclk));
	jor g0016(.dina(n87),.dinb(w_n84_1[2]),.dout(n88),.clk(gclk));
	jnot g0017(.din(w_G13_2[1]),.dout(n89),.clk(gclk));
	jand g0018(.dina(w_n89_0[1]),.dinb(w_G1_2[1]),.dout(n90),.clk(gclk));
	jand g0019(.dina(w_n90_0[2]),.dinb(w_G20_6[2]),.dout(n91),.clk(gclk));
	jand g0020(.dina(w_n91_1[2]),.dinb(n88),.dout(n92),.clk(gclk));
	jor g0021(.dina(w_n85_0[0]),.dinb(w_n80_1[1]),.dout(n93),.clk(gclk));
	jnot g0022(.din(w_G244_1[1]),.dout(n94),.clk(gclk));
	jor g0023(.dina(w_n94_0[2]),.dinb(w_n72_1[1]),.dout(n95),.clk(gclk));
	jnot g0024(.din(w_G238_0[2]),.dout(n96),.clk(gclk));
	jor g0025(.dina(w_n96_0[2]),.dinb(w_n75_2[0]),.dout(n97),.clk(gclk));
	jand g0026(.dina(n97),.dinb(n95),.dout(n98),.clk(gclk));
	jnot g0027(.din(w_G226_1[2]),.dout(n99),.clk(gclk));
	jor g0028(.dina(n99),.dinb(w_n73_2[1]),.dout(n100),.clk(gclk));
	jand g0029(.dina(n100),.dinb(n98),.dout(n101),.clk(gclk));
	jand g0030(.dina(n101),.dinb(n93),.dout(n102),.clk(gclk));
	jnot g0031(.din(w_G232_1[2]),.dout(n103),.clk(gclk));
	jor g0032(.dina(n103),.dinb(w_n74_2[0]),.dout(n104),.clk(gclk));
	jnot g0033(.din(w_G116_5[2]),.dout(n105),.clk(gclk));
	jnot g0034(.din(w_G270_0[2]),.dout(n106),.clk(gclk));
	jor g0035(.dina(n106),.dinb(w_n105_1[1]),.dout(n107),.clk(gclk));
	jand g0036(.dina(n107),.dinb(n104),.dout(n108),.clk(gclk));
	jor g0037(.dina(w_n86_0[1]),.dinb(w_n81_2[0]),.dout(n109),.clk(gclk));
	jand g0038(.dina(n109),.dinb(n108),.dout(n110),.clk(gclk));
	jand g0039(.dina(w_G20_6[1]),.dinb(w_G1_2[0]),.dout(n111),.clk(gclk));
	jnot g0040(.din(w_n111_0[2]),.dout(n112),.clk(gclk));
	jor g0041(.dina(w_n84_1[1]),.dinb(w_n79_1[1]),.dout(n113),.clk(gclk));
	jand g0042(.dina(n113),.dinb(w_n112_0[1]),.dout(n114),.clk(gclk));
	jand g0043(.dina(n114),.dinb(n110),.dout(n115),.clk(gclk));
	jand g0044(.dina(n115),.dinb(n102),.dout(n116),.clk(gclk));
	jnot g0045(.din(w_n76_0[0]),.dout(n117),.clk(gclk));
	jand g0046(.dina(n117),.dinb(w_G50_5[1]),.dout(n118),.clk(gclk));
	jnot g0047(.din(w_n118_0[2]),.dout(n119),.clk(gclk));
	jand g0048(.dina(w_n111_0[1]),.dinb(w_G13_2[0]),.dout(n120),.clk(gclk));
	jand g0049(.dina(w_n120_0[1]),.dinb(n119),.dout(n121),.clk(gclk));
	jor g0050(.dina(n121),.dinb(n116),.dout(n122),.clk(gclk));
	jor g0051(.dina(n122),.dinb(w_dff_B_Mt4cKI405_1),.dout(w_dff_A_tGv9QlUg2_2),.clk(gclk));
	jxor g0052(.dina(w_G270_0[1]),.dinb(w_n86_0[0]),.dout(n124),.clk(gclk));
	jxor g0053(.dina(w_G257_1[1]),.dinb(w_G250_0[1]),.dout(n125),.clk(gclk));
	jxor g0054(.dina(n125),.dinb(n124),.dout(n126),.clk(gclk));
	jnot g0055(.din(w_n126_0[1]),.dout(n127),.clk(gclk));
	jxor g0056(.dina(w_G244_1[0]),.dinb(w_n96_0[1]),.dout(n128),.clk(gclk));
	jxor g0057(.dina(w_G232_1[1]),.dinb(w_G226_1[1]),.dout(n129),.clk(gclk));
	jxor g0058(.dina(n129),.dinb(n128),.dout(n130),.clk(gclk));
	jxor g0059(.dina(w_n130_0[1]),.dinb(n127),.dout(w_dff_A_FASwSrM37_2),.clk(gclk));
	jxor g0060(.dina(w_G58_5[1]),.dinb(w_G50_5[0]),.dout(n132),.clk(gclk));
	jxor g0061(.dina(w_G77_4[1]),.dinb(w_G68_5[1]),.dout(n133),.clk(gclk));
	jxor g0062(.dina(n133),.dinb(n132),.dout(n134),.clk(gclk));
	jxor g0063(.dina(w_G116_5[1]),.dinb(w_n81_1[2]),.dout(n135),.clk(gclk));
	jxor g0064(.dina(w_G97_4[1]),.dinb(w_G87_3[1]),.dout(n136),.clk(gclk));
	jxor g0065(.dina(n136),.dinb(n135),.dout(n137),.clk(gclk));
	jxor g0066(.dina(w_n137_0[1]),.dinb(w_n134_0[1]),.dout(w_dff_A_aHt6RkCZ8_2),.clk(gclk));
	jand g0067(.dina(w_G13_1[2]),.dinb(w_G1_1[2]),.dout(n139),.clk(gclk));
	jand g0068(.dina(w_n111_0[0]),.dinb(w_G33_12[2]),.dout(n140),.clk(gclk));
	jor g0069(.dina(w_n140_0[1]),.dinb(w_n139_1[2]),.dout(n141),.clk(gclk));
	jnot g0070(.din(w_G1_1[1]),.dout(n142),.clk(gclk));
	jand g0071(.dina(w_G13_1[1]),.dinb(w_n142_2[1]),.dout(n143),.clk(gclk));
	jand g0072(.dina(w_n143_0[1]),.dinb(w_G20_6[0]),.dout(n144),.clk(gclk));
	jor g0073(.dina(w_n144_2[1]),.dinb(w_n141_3[1]),.dout(n145),.clk(gclk));
	jand g0074(.dina(w_G33_12[1]),.dinb(w_n142_2[0]),.dout(n146),.clk(gclk));
	jor g0075(.dina(n146),.dinb(n145),.dout(n147),.clk(gclk));
	jnot g0076(.din(w_n147_0[2]),.dout(n148),.clk(gclk));
	jand g0077(.dina(w_n148_0[1]),.dinb(w_G116_5[0]),.dout(n149),.clk(gclk));
	jand g0078(.dina(w_G116_4[2]),.dinb(w_G20_5[2]),.dout(n150),.clk(gclk));
	jnot g0079(.din(w_G20_5[1]),.dout(n151),.clk(gclk));
	jand g0080(.dina(w_G283_3[2]),.dinb(w_G33_12[0]),.dout(n152),.clk(gclk));
	jnot g0081(.din(w_G33_11[2]),.dout(n153),.clk(gclk));
	jand g0082(.dina(w_G97_4[0]),.dinb(w_n153_8[1]),.dout(n154),.clk(gclk));
	jor g0083(.dina(n154),.dinb(w_n152_0[2]),.dout(n155),.clk(gclk));
	jand g0084(.dina(n155),.dinb(w_n151_6[1]),.dout(n156),.clk(gclk));
	jor g0085(.dina(n156),.dinb(n150),.dout(n157),.clk(gclk));
	jand g0086(.dina(n157),.dinb(w_n141_3[0]),.dout(n158),.clk(gclk));
	jand g0087(.dina(w_n144_2[0]),.dinb(w_n105_1[0]),.dout(n159),.clk(gclk));
	jor g0088(.dina(n159),.dinb(n158),.dout(n160),.clk(gclk));
	jor g0089(.dina(n160),.dinb(n149),.dout(n161),.clk(gclk));
	jnot g0090(.din(w_n161_0[2]),.dout(n162),.clk(gclk));
	jnot g0091(.din(w_G41_0[2]),.dout(n163),.clk(gclk));
	jand g0092(.dina(w_G45_1[1]),.dinb(w_n142_1[2]),.dout(n164),.clk(gclk));
	jand g0093(.dina(w_n164_0[2]),.dinb(w_n163_1[1]),.dout(n165),.clk(gclk));
	jnot g0094(.din(w_n139_1[1]),.dout(n166),.clk(gclk));
	jand g0095(.dina(w_G41_0[1]),.dinb(w_G33_11[1]),.dout(n167),.clk(gclk));
	jor g0096(.dina(w_n167_0[1]),.dinb(n166),.dout(n168),.clk(gclk));
	jand g0097(.dina(w_n168_5[1]),.dinb(w_G274_0[2]),.dout(n169),.clk(gclk));
	jand g0098(.dina(w_n169_0[1]),.dinb(w_n165_0[1]),.dout(n170),.clk(gclk));
	jnot g0099(.din(w_n167_0[0]),.dout(n171),.clk(gclk));
	jand g0100(.dina(n171),.dinb(w_n139_1[0]),.dout(n172),.clk(gclk));
	jand g0101(.dina(w_G1698_0[2]),.dinb(w_n153_8[0]),.dout(n173),.clk(gclk));
	jand g0102(.dina(w_n173_3[1]),.dinb(w_G264_0[1]),.dout(n174),.clk(gclk));
	jand g0103(.dina(w_G303_2[2]),.dinb(w_G33_11[0]),.dout(n175),.clk(gclk));
	jnot g0104(.din(w_G1698_0[1]),.dout(n176),.clk(gclk));
	jand g0105(.dina(w_n176_0[1]),.dinb(w_n153_7[2]),.dout(n177),.clk(gclk));
	jand g0106(.dina(w_n177_1[2]),.dinb(w_G257_1[0]),.dout(n178),.clk(gclk));
	jor g0107(.dina(n178),.dinb(n175),.dout(n179),.clk(gclk));
	jor g0108(.dina(n179),.dinb(n174),.dout(n180),.clk(gclk));
	jand g0109(.dina(n180),.dinb(w_n172_4[2]),.dout(n181),.clk(gclk));
	jnot g0110(.din(w_n165_0[0]),.dout(n182),.clk(gclk));
	jand g0111(.dina(w_n168_5[0]),.dinb(w_G270_0[0]),.dout(n183),.clk(gclk));
	jand g0112(.dina(n183),.dinb(w_n182_1[1]),.dout(n184),.clk(gclk));
	jor g0113(.dina(n184),.dinb(n181),.dout(n185),.clk(gclk));
	jor g0114(.dina(n185),.dinb(w_n170_0[2]),.dout(n186),.clk(gclk));
	jand g0115(.dina(w_n186_1[2]),.dinb(w_G169_3[1]),.dout(n187),.clk(gclk));
	jnot g0116(.din(n187),.dout(n188),.clk(gclk));
	jnot g0117(.din(w_G179_2[2]),.dout(n189),.clk(gclk));
	jor g0118(.dina(w_n186_1[1]),.dinb(w_n189_2[2]),.dout(n190),.clk(gclk));
	jand g0119(.dina(w_n190_0[1]),.dinb(n188),.dout(n191),.clk(gclk));
	jor g0120(.dina(n191),.dinb(n162),.dout(n192),.clk(gclk));
	jand g0121(.dina(w_n186_1[0]),.dinb(w_G200_3[1]),.dout(n193),.clk(gclk));
	jnot g0122(.din(w_n186_0[2]),.dout(n194),.clk(gclk));
	jand g0123(.dina(n194),.dinb(w_G190_4[2]),.dout(n195),.clk(gclk));
	jor g0124(.dina(n195),.dinb(w_n161_0[1]),.dout(n196),.clk(gclk));
	jor g0125(.dina(n196),.dinb(n193),.dout(n197),.clk(gclk));
	jand g0126(.dina(n197),.dinb(w_n192_0[2]),.dout(n198),.clk(gclk));
	jnot g0127(.din(w_G169_3[0]),.dout(n199),.clk(gclk));
	jand g0128(.dina(w_n168_4[2]),.dinb(w_G264_0[0]),.dout(n200),.clk(gclk));
	jand g0129(.dina(n200),.dinb(w_n182_1[0]),.dout(n201),.clk(gclk));
	jand g0130(.dina(w_n173_3[0]),.dinb(w_G257_0[2]),.dout(n202),.clk(gclk));
	jand g0131(.dina(w_G294_3[1]),.dinb(w_G33_10[2]),.dout(n203),.clk(gclk));
	jnot g0132(.din(n203),.dout(n204),.clk(gclk));
	jor g0133(.dina(w_G1698_0[0]),.dinb(w_G33_10[1]),.dout(n205),.clk(gclk));
	jor g0134(.dina(w_n205_1[1]),.dinb(w_n84_1[0]),.dout(n206),.clk(gclk));
	jand g0135(.dina(n206),.dinb(n204),.dout(n207),.clk(gclk));
	jnot g0136(.din(w_n207_0[1]),.dout(n208),.clk(gclk));
	jor g0137(.dina(n208),.dinb(w_n202_0[1]),.dout(n209),.clk(gclk));
	jand g0138(.dina(n209),.dinb(w_n172_4[1]),.dout(n210),.clk(gclk));
	jor g0139(.dina(n210),.dinb(w_n170_0[1]),.dout(n211),.clk(gclk));
	jor g0140(.dina(n211),.dinb(w_n201_0[1]),.dout(n212),.clk(gclk));
	jand g0141(.dina(w_n212_1[1]),.dinb(w_n199_0[2]),.dout(n213),.clk(gclk));
	jand g0142(.dina(w_n148_0[0]),.dinb(w_G107_4[0]),.dout(n214),.clk(gclk));
	jor g0143(.dina(w_n140_0[0]),.dinb(w_G13_1[0]),.dout(n215),.clk(gclk));
	jand g0144(.dina(w_n81_1[1]),.dinb(w_G20_5[0]),.dout(n216),.clk(gclk));
	jand g0145(.dina(n216),.dinb(w_n215_0[1]),.dout(n217),.clk(gclk));
	jand g0146(.dina(w_G116_4[1]),.dinb(w_G33_10[0]),.dout(n218),.clk(gclk));
	jand g0147(.dina(w_G87_3[0]),.dinb(w_n153_7[1]),.dout(n219),.clk(gclk));
	jor g0148(.dina(n219),.dinb(w_n218_0[1]),.dout(n220),.clk(gclk));
	jand g0149(.dina(n220),.dinb(w_n141_2[2]),.dout(n221),.clk(gclk));
	jand g0150(.dina(n221),.dinb(w_n151_6[0]),.dout(n222),.clk(gclk));
	jor g0151(.dina(n222),.dinb(n217),.dout(n223),.clk(gclk));
	jor g0152(.dina(n223),.dinb(n214),.dout(n224),.clk(gclk));
	jnot g0153(.din(w_n224_1[1]),.dout(n225),.clk(gclk));
	jnot g0154(.din(w_n201_0[0]),.dout(n226),.clk(gclk));
	jnot g0155(.din(w_G274_0[1]),.dout(n227),.clk(gclk));
	jor g0156(.dina(w_n172_4[0]),.dinb(n227),.dout(n228),.clk(gclk));
	jor g0157(.dina(n228),.dinb(w_n182_0[2]),.dout(n229),.clk(gclk));
	jnot g0158(.din(w_n202_0[0]),.dout(n230),.clk(gclk));
	jand g0159(.dina(w_n207_0[0]),.dinb(n230),.dout(n231),.clk(gclk));
	jor g0160(.dina(n231),.dinb(w_n168_4[1]),.dout(n232),.clk(gclk));
	jand g0161(.dina(n232),.dinb(w_n229_0[1]),.dout(n233),.clk(gclk));
	jand g0162(.dina(n233),.dinb(n226),.dout(n234),.clk(gclk));
	jand g0163(.dina(w_n234_1[1]),.dinb(w_n189_2[1]),.dout(n235),.clk(gclk));
	jor g0164(.dina(n235),.dinb(w_n225_0[1]),.dout(n236),.clk(gclk));
	jor g0165(.dina(n236),.dinb(w_n213_0[1]),.dout(n237),.clk(gclk));
	jand g0166(.dina(w_n234_1[0]),.dinb(w_G190_4[1]),.dout(n238),.clk(gclk));
	jand g0167(.dina(w_n212_1[0]),.dinb(w_G200_3[0]),.dout(n239),.clk(gclk));
	jor g0168(.dina(n239),.dinb(w_n224_1[0]),.dout(n240),.clk(gclk));
	jor g0169(.dina(n240),.dinb(w_n238_0[1]),.dout(n241),.clk(gclk));
	jand g0170(.dina(n241),.dinb(w_n237_0[2]),.dout(n242),.clk(gclk));
	jand g0171(.dina(w_n173_2[2]),.dinb(w_G244_0[2]),.dout(n243),.clk(gclk));
	jnot g0172(.din(w_n243_0[1]),.dout(n244),.clk(gclk));
	jnot g0173(.din(w_n218_0[0]),.dout(n245),.clk(gclk));
	jor g0174(.dina(w_n205_1[0]),.dinb(w_n96_0[0]),.dout(n246),.clk(gclk));
	jand g0175(.dina(n246),.dinb(n245),.dout(n247),.clk(gclk));
	jand g0176(.dina(w_n247_0[1]),.dinb(n244),.dout(n248),.clk(gclk));
	jand g0177(.dina(n248),.dinb(w_n172_3[2]),.dout(n249),.clk(gclk));
	jor g0178(.dina(w_n164_0[1]),.dinb(w_n84_0[2]),.dout(n250),.clk(gclk));
	jand g0179(.dina(w_n164_0[0]),.dinb(w_G274_0[0]),.dout(n251),.clk(gclk));
	jnot g0180(.din(w_n251_0[1]),.dout(n252),.clk(gclk));
	jand g0181(.dina(n252),.dinb(w_n250_0[1]),.dout(n253),.clk(gclk));
	jand g0182(.dina(n253),.dinb(w_n168_4[0]),.dout(n254),.clk(gclk));
	jor g0183(.dina(n254),.dinb(n249),.dout(n255),.clk(gclk));
	jand g0184(.dina(w_n255_1[1]),.dinb(w_n189_2[0]),.dout(n256),.clk(gclk));
	jor g0185(.dina(w_n147_0[1]),.dinb(w_n79_1[0]),.dout(n257),.clk(gclk));
	jand g0186(.dina(w_n80_1[0]),.dinb(w_n79_0[2]),.dout(n258),.clk(gclk));
	jand g0187(.dina(n258),.dinb(w_n81_1[0]),.dout(n259),.clk(gclk));
	jand g0188(.dina(w_n259_0[1]),.dinb(w_G20_4[2]),.dout(n260),.clk(gclk));
	jnot g0189(.din(w_n141_2[1]),.dout(n261),.clk(gclk));
	jand g0190(.dina(w_G97_3[2]),.dinb(w_G33_9[2]),.dout(n262),.clk(gclk));
	jnot g0191(.din(w_n262_0[2]),.dout(n263),.clk(gclk));
	jor g0192(.dina(w_n75_1[2]),.dinb(w_G33_9[1]),.dout(n264),.clk(gclk));
	jand g0193(.dina(n264),.dinb(w_n151_5[2]),.dout(n265),.clk(gclk));
	jand g0194(.dina(n265),.dinb(n263),.dout(n266),.clk(gclk));
	jor g0195(.dina(n266),.dinb(w_n261_1[2]),.dout(n267),.clk(gclk));
	jor g0196(.dina(n267),.dinb(w_n260_0[1]),.dout(n268),.clk(gclk));
	jand g0197(.dina(w_n144_1[2]),.dinb(w_n79_0[1]),.dout(n269),.clk(gclk));
	jnot g0198(.din(w_n269_0[1]),.dout(n270),.clk(gclk));
	jand g0199(.dina(n270),.dinb(n268),.dout(n271),.clk(gclk));
	jand g0200(.dina(n271),.dinb(w_n257_0[1]),.dout(n272),.clk(gclk));
	jnot g0201(.din(w_n247_0[0]),.dout(n273),.clk(gclk));
	jor g0202(.dina(n273),.dinb(w_n243_0[0]),.dout(n274),.clk(gclk));
	jor g0203(.dina(n274),.dinb(w_n168_3[2]),.dout(n275),.clk(gclk));
	jnot g0204(.din(w_n250_0[0]),.dout(n276),.clk(gclk));
	jor g0205(.dina(w_n251_0[0]),.dinb(n276),.dout(n277),.clk(gclk));
	jor g0206(.dina(n277),.dinb(w_n172_3[1]),.dout(n278),.clk(gclk));
	jand g0207(.dina(n278),.dinb(n275),.dout(n279),.clk(gclk));
	jand g0208(.dina(w_n279_1[1]),.dinb(w_n199_0[1]),.dout(n280),.clk(gclk));
	jor g0209(.dina(n280),.dinb(w_n272_0[1]),.dout(n281),.clk(gclk));
	jor g0210(.dina(n281),.dinb(w_n256_0[1]),.dout(n282),.clk(gclk));
	jand g0211(.dina(w_n279_1[0]),.dinb(w_G200_2[2]),.dout(n283),.clk(gclk));
	jnot g0212(.din(w_n257_0[0]),.dout(n284),.clk(gclk));
	jnot g0213(.din(w_n260_0[0]),.dout(n285),.clk(gclk));
	jand g0214(.dina(w_G68_5[0]),.dinb(w_n153_7[0]),.dout(n286),.clk(gclk));
	jor g0215(.dina(n286),.dinb(w_G20_4[1]),.dout(n287),.clk(gclk));
	jor g0216(.dina(n287),.dinb(w_n262_0[1]),.dout(n288),.clk(gclk));
	jand g0217(.dina(n288),.dinb(w_n141_2[0]),.dout(n289),.clk(gclk));
	jand g0218(.dina(n289),.dinb(n285),.dout(n290),.clk(gclk));
	jor g0219(.dina(w_n269_0[0]),.dinb(n290),.dout(n291),.clk(gclk));
	jor g0220(.dina(n291),.dinb(n284),.dout(n292),.clk(gclk));
	jand g0221(.dina(w_n255_1[0]),.dinb(w_G190_4[0]),.dout(n293),.clk(gclk));
	jor g0222(.dina(n293),.dinb(w_n292_0[2]),.dout(n294),.clk(gclk));
	jor g0223(.dina(n294),.dinb(w_n283_0[1]),.dout(n295),.clk(gclk));
	jand g0224(.dina(n295),.dinb(w_n282_0[1]),.dout(n296),.clk(gclk));
	jand g0225(.dina(w_n168_3[1]),.dinb(w_G257_0[1]),.dout(n297),.clk(gclk));
	jand g0226(.dina(n297),.dinb(w_n182_0[1]),.dout(n298),.clk(gclk));
	jnot g0227(.din(w_n298_0[1]),.dout(n299),.clk(gclk));
	jor g0228(.dina(w_n176_0[0]),.dinb(w_G33_9[0]),.dout(n300),.clk(gclk));
	jor g0229(.dina(n300),.dinb(w_n84_0[1]),.dout(n301),.clk(gclk));
	jnot g0230(.din(w_n152_0[1]),.dout(n302),.clk(gclk));
	jor g0231(.dina(w_n205_0[2]),.dinb(w_n94_0[1]),.dout(n303),.clk(gclk));
	jand g0232(.dina(n303),.dinb(n302),.dout(n304),.clk(gclk));
	jand g0233(.dina(n304),.dinb(n301),.dout(n305),.clk(gclk));
	jor g0234(.dina(n305),.dinb(w_n168_3[0]),.dout(n306),.clk(gclk));
	jand g0235(.dina(n306),.dinb(w_n229_0[0]),.dout(n307),.clk(gclk));
	jand g0236(.dina(n307),.dinb(n299),.dout(n308),.clk(gclk));
	jand g0237(.dina(w_n308_1[2]),.dinb(w_G190_3[2]),.dout(n309),.clk(gclk));
	jor g0238(.dina(w_n147_0[0]),.dinb(w_n80_0[2]),.dout(n310),.clk(gclk));
	jnot g0239(.din(w_n310_0[1]),.dout(n311),.clk(gclk));
	jxor g0240(.dina(w_G107_3[2]),.dinb(w_G97_3[1]),.dout(n312),.clk(gclk));
	jand g0241(.dina(w_n312_0[1]),.dinb(w_G20_4[0]),.dout(n313),.clk(gclk));
	jnot g0242(.din(w_n313_0[1]),.dout(n314),.clk(gclk));
	jand g0243(.dina(w_G107_3[1]),.dinb(w_G33_8[2]),.dout(n315),.clk(gclk));
	jand g0244(.dina(w_G77_4[0]),.dinb(w_n153_6[2]),.dout(n316),.clk(gclk));
	jor g0245(.dina(n316),.dinb(w_G20_3[2]),.dout(n317),.clk(gclk));
	jor g0246(.dina(n317),.dinb(w_n315_0[2]),.dout(n318),.clk(gclk));
	jand g0247(.dina(n318),.dinb(w_n141_1[2]),.dout(n319),.clk(gclk));
	jand g0248(.dina(n319),.dinb(n314),.dout(n320),.clk(gclk));
	jand g0249(.dina(w_n144_1[1]),.dinb(w_n80_0[1]),.dout(n321),.clk(gclk));
	jor g0250(.dina(w_n321_0[1]),.dinb(n320),.dout(n322),.clk(gclk));
	jor g0251(.dina(n322),.dinb(n311),.dout(n323),.clk(gclk));
	jand g0252(.dina(w_n173_2[1]),.dinb(w_G250_0[0]),.dout(n324),.clk(gclk));
	jand g0253(.dina(w_n177_1[1]),.dinb(w_G244_0[1]),.dout(n325),.clk(gclk));
	jor g0254(.dina(n325),.dinb(w_n152_0[0]),.dout(n326),.clk(gclk));
	jor g0255(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jand g0256(.dina(n327),.dinb(w_n172_3[0]),.dout(n328),.clk(gclk));
	jor g0257(.dina(n328),.dinb(w_n170_0[0]),.dout(n329),.clk(gclk));
	jor g0258(.dina(n329),.dinb(w_n298_0[0]),.dout(n330),.clk(gclk));
	jand g0259(.dina(w_n330_0[2]),.dinb(w_G200_2[1]),.dout(n331),.clk(gclk));
	jor g0260(.dina(n331),.dinb(w_n323_0[2]),.dout(n332),.clk(gclk));
	jor g0261(.dina(n332),.dinb(w_n309_0[1]),.dout(n333),.clk(gclk));
	jor g0262(.dina(w_n308_1[1]),.dinb(w_G169_2[2]),.dout(n334),.clk(gclk));
	jnot g0263(.din(w_n334_0[1]),.dout(n335),.clk(gclk));
	jnot g0264(.din(w_n315_0[1]),.dout(n336),.clk(gclk));
	jor g0265(.dina(w_n72_1[0]),.dinb(w_G33_8[1]),.dout(n337),.clk(gclk));
	jand g0266(.dina(n337),.dinb(w_n151_5[1]),.dout(n338),.clk(gclk));
	jand g0267(.dina(n338),.dinb(n336),.dout(n339),.clk(gclk));
	jor g0268(.dina(n339),.dinb(w_n261_1[1]),.dout(n340),.clk(gclk));
	jor g0269(.dina(n340),.dinb(w_n313_0[0]),.dout(n341),.clk(gclk));
	jnot g0270(.din(w_n321_0[0]),.dout(n342),.clk(gclk));
	jand g0271(.dina(n342),.dinb(n341),.dout(n343),.clk(gclk));
	jand g0272(.dina(n343),.dinb(w_n310_0[0]),.dout(n344),.clk(gclk));
	jand g0273(.dina(w_n308_1[0]),.dinb(w_n189_1[2]),.dout(n345),.clk(gclk));
	jor g0274(.dina(n345),.dinb(w_n344_0[1]),.dout(n346),.clk(gclk));
	jor g0275(.dina(n346),.dinb(n335),.dout(n347),.clk(gclk));
	jand g0276(.dina(w_n347_0[1]),.dinb(w_n333_0[1]),.dout(n348),.clk(gclk));
	jand g0277(.dina(w_n348_0[1]),.dinb(n296),.dout(n349),.clk(gclk));
	jand g0278(.dina(w_n349_0[1]),.dinb(w_n242_0[2]),.dout(n350),.clk(gclk));
	jand g0279(.dina(w_n350_0[1]),.dinb(w_n198_0[2]),.dout(n351),.clk(gclk));
	jnot g0280(.din(w_G45_1[0]),.dout(n352),.clk(gclk));
	jand g0281(.dina(w_n352_1[1]),.dinb(w_n163_1[0]),.dout(n353),.clk(gclk));
	jor g0282(.dina(n353),.dinb(w_G1_1[0]),.dout(n354),.clk(gclk));
	jnot g0283(.din(w_n354_1[1]),.dout(n355),.clk(gclk));
	jand g0284(.dina(w_n355_0[1]),.dinb(w_n169_0[0]),.dout(n356),.clk(gclk));
	jnot g0285(.din(w_n356_1[1]),.dout(n357),.clk(gclk));
	jand g0286(.dina(w_n173_2[0]),.dinb(w_G238_0[1]),.dout(n358),.clk(gclk));
	jand g0287(.dina(w_n177_1[0]),.dinb(w_G232_1[0]),.dout(n359),.clk(gclk));
	jor g0288(.dina(n359),.dinb(w_n315_0[0]),.dout(n360),.clk(gclk));
	jor g0289(.dina(n360),.dinb(n358),.dout(n361),.clk(gclk));
	jand g0290(.dina(n361),.dinb(w_n172_2[2]),.dout(n362),.clk(gclk));
	jnot g0291(.din(n362),.dout(n363),.clk(gclk));
	jor g0292(.dina(w_n355_0[0]),.dinb(w_n94_0[0]),.dout(n364),.clk(gclk));
	jor g0293(.dina(n364),.dinb(w_n172_2[1]),.dout(n365),.clk(gclk));
	jand g0294(.dina(n365),.dinb(n363),.dout(n366),.clk(gclk));
	jand g0295(.dina(n366),.dinb(w_n357_0[1]),.dout(n367),.clk(gclk));
	jnot g0296(.din(w_n367_1[1]),.dout(n368),.clk(gclk));
	jand g0297(.dina(n368),.dinb(w_n199_0[0]),.dout(n369),.clk(gclk));
	jand g0298(.dina(w_G87_2[2]),.dinb(w_G33_8[0]),.dout(n370),.clk(gclk));
	jand g0299(.dina(w_G58_5[0]),.dinb(w_n153_6[1]),.dout(n371),.clk(gclk));
	jor g0300(.dina(n371),.dinb(w_n370_0[1]),.dout(n372),.clk(gclk));
	jand g0301(.dina(n372),.dinb(w_n151_5[0]),.dout(n373),.clk(gclk));
	jand g0302(.dina(n373),.dinb(w_n141_1[1]),.dout(n374),.clk(gclk));
	jand g0303(.dina(w_n139_0[2]),.dinb(w_n151_4[2]),.dout(n375),.clk(gclk));
	jnot g0304(.din(w_n375_0[1]),.dout(n376),.clk(gclk));
	jand g0305(.dina(w_G20_3[1]),.dinb(w_n142_1[1]),.dout(n377),.clk(gclk));
	jnot g0306(.din(n377),.dout(n378),.clk(gclk));
	jand g0307(.dina(w_n378_0[1]),.dinb(w_G77_3[2]),.dout(n379),.clk(gclk));
	jand g0308(.dina(n379),.dinb(n376),.dout(n380),.clk(gclk));
	jand g0309(.dina(w_n144_1[0]),.dinb(w_n72_0[2]),.dout(n381),.clk(gclk));
	jor g0310(.dina(n381),.dinb(n380),.dout(n382),.clk(gclk));
	jor g0311(.dina(n382),.dinb(n374),.dout(n383),.clk(gclk));
	jnot g0312(.din(w_n383_0[2]),.dout(n384),.clk(gclk));
	jand g0313(.dina(w_n367_1[0]),.dinb(w_n189_1[1]),.dout(n385),.clk(gclk));
	jor g0314(.dina(n385),.dinb(n384),.dout(n386),.clk(gclk));
	jor g0315(.dina(n386),.dinb(n369),.dout(n387),.clk(gclk));
	jnot g0316(.din(w_G200_2[0]),.dout(n388),.clk(gclk));
	jor g0317(.dina(w_n367_0[2]),.dinb(w_n388_2[1]),.dout(n389),.clk(gclk));
	jnot g0318(.din(n389),.dout(n390),.clk(gclk));
	jand g0319(.dina(w_n367_0[1]),.dinb(w_G190_3[1]),.dout(n391),.clk(gclk));
	jor g0320(.dina(n391),.dinb(w_n383_0[1]),.dout(n392),.clk(gclk));
	jor g0321(.dina(n392),.dinb(n390),.dout(n393),.clk(gclk));
	jand g0322(.dina(n393),.dinb(w_n387_0[2]),.dout(n394),.clk(gclk));
	jnot g0323(.din(w_n394_0[1]),.dout(n395),.clk(gclk));
	jand g0324(.dina(w_n168_2[2]),.dinb(w_G238_0[0]),.dout(n396),.clk(gclk));
	jand g0325(.dina(n396),.dinb(w_n354_1[0]),.dout(n397),.clk(gclk));
	jand g0326(.dina(w_n173_1[2]),.dinb(w_G232_0[2]),.dout(n398),.clk(gclk));
	jand g0327(.dina(w_n177_0[2]),.dinb(w_G226_1[0]),.dout(n399),.clk(gclk));
	jor g0328(.dina(n399),.dinb(w_n262_0[0]),.dout(n400),.clk(gclk));
	jor g0329(.dina(n400),.dinb(n398),.dout(n401),.clk(gclk));
	jand g0330(.dina(n401),.dinb(w_n172_2[0]),.dout(n402),.clk(gclk));
	jor g0331(.dina(n402),.dinb(w_n356_1[0]),.dout(n403),.clk(gclk));
	jor g0332(.dina(n403),.dinb(n397),.dout(n404),.clk(gclk));
	jnot g0333(.din(w_n404_0[2]),.dout(n405),.clk(gclk));
	jor g0334(.dina(w_n405_0[1]),.dinb(w_G169_2[1]),.dout(n406),.clk(gclk));
	jand g0335(.dina(w_G77_3[1]),.dinb(w_G33_7[2]),.dout(n407),.clk(gclk));
	jand g0336(.dina(w_G50_4[2]),.dinb(w_n153_6[0]),.dout(n408),.clk(gclk));
	jor g0337(.dina(n408),.dinb(w_n407_0[1]),.dout(n409),.clk(gclk));
	jand g0338(.dina(n409),.dinb(w_n141_1[0]),.dout(n410),.clk(gclk));
	jand g0339(.dina(n410),.dinb(w_n151_4[1]),.dout(n411),.clk(gclk));
	jand g0340(.dina(w_n75_1[1]),.dinb(w_G20_3[0]),.dout(n412),.clk(gclk));
	jand g0341(.dina(n412),.dinb(w_n215_0[0]),.dout(n413),.clk(gclk));
	jand g0342(.dina(w_n378_0[0]),.dinb(w_n261_1[0]),.dout(n414),.clk(gclk));
	jand g0343(.dina(w_n414_0[2]),.dinb(w_G68_4[2]),.dout(n415),.clk(gclk));
	jor g0344(.dina(n415),.dinb(n413),.dout(n416),.clk(gclk));
	jor g0345(.dina(n416),.dinb(n411),.dout(n417),.clk(gclk));
	jor g0346(.dina(w_n404_0[1]),.dinb(w_G179_2[1]),.dout(n418),.clk(gclk));
	jand g0347(.dina(n418),.dinb(w_n417_0[2]),.dout(n419),.clk(gclk));
	jand g0348(.dina(n419),.dinb(n406),.dout(n420),.clk(gclk));
	jand g0349(.dina(w_n405_0[0]),.dinb(w_G190_3[0]),.dout(n421),.clk(gclk));
	jand g0350(.dina(w_n404_0[0]),.dinb(w_G200_1[2]),.dout(n422),.clk(gclk));
	jor g0351(.dina(n422),.dinb(w_n417_0[1]),.dout(n423),.clk(gclk));
	jor g0352(.dina(n423),.dinb(n421),.dout(n424),.clk(gclk));
	jnot g0353(.din(n424),.dout(n425),.clk(gclk));
	jor g0354(.dina(w_n425_0[1]),.dinb(w_n420_0[1]),.dout(n426),.clk(gclk));
	jand g0355(.dina(w_n168_2[1]),.dinb(w_G226_0[2]),.dout(n427),.clk(gclk));
	jand g0356(.dina(n427),.dinb(w_n354_0[2]),.dout(n428),.clk(gclk));
	jnot g0357(.din(w_n428_0[1]),.dout(n429),.clk(gclk));
	jand g0358(.dina(w_n173_1[1]),.dinb(w_G223_0[1]),.dout(n430),.clk(gclk));
	jnot g0359(.din(w_n430_0[1]),.dout(n431),.clk(gclk));
	jnot g0360(.din(w_n407_0[0]),.dout(n432),.clk(gclk));
	jnot g0361(.din(G222),.dout(n433),.clk(gclk));
	jor g0362(.dina(w_n205_0[1]),.dinb(n433),.dout(n434),.clk(gclk));
	jand g0363(.dina(n434),.dinb(n432),.dout(n435),.clk(gclk));
	jand g0364(.dina(w_n435_0[1]),.dinb(n431),.dout(n436),.clk(gclk));
	jor g0365(.dina(n436),.dinb(w_n168_2[0]),.dout(n437),.clk(gclk));
	jand g0366(.dina(n437),.dinb(w_n357_0[0]),.dout(n438),.clk(gclk));
	jand g0367(.dina(n438),.dinb(n429),.dout(n439),.clk(gclk));
	jor g0368(.dina(w_n439_0[2]),.dinb(w_G169_2[0]),.dout(n440),.clk(gclk));
	jand g0369(.dina(w_G33_7[1]),.dinb(w_n151_4[0]),.dout(n441),.clk(gclk));
	jand g0370(.dina(w_n441_0[1]),.dinb(w_G58_4[2]),.dout(n442),.clk(gclk));
	jnot g0371(.din(n442),.dout(n443),.clk(gclk));
	jor g0372(.dina(w_n77_0[0]),.dinb(w_n151_3[2]),.dout(n444),.clk(gclk));
	jand g0373(.dina(w_n153_5[2]),.dinb(w_n151_3[1]),.dout(n445),.clk(gclk));
	jand g0374(.dina(w_n445_0[1]),.dinb(w_G150_3[1]),.dout(n446),.clk(gclk));
	jnot g0375(.din(n446),.dout(n447),.clk(gclk));
	jand g0376(.dina(n447),.dinb(n444),.dout(n448),.clk(gclk));
	jand g0377(.dina(n448),.dinb(n443),.dout(n449),.clk(gclk));
	jor g0378(.dina(n449),.dinb(w_n261_0[2]),.dout(n450),.clk(gclk));
	jnot g0379(.din(w_n450_0[1]),.dout(n451),.clk(gclk));
	jnot g0380(.din(w_n144_0[2]),.dout(n452),.clk(gclk));
	jand g0381(.dina(w_n452_0[1]),.dinb(w_n73_2[0]),.dout(n453),.clk(gclk));
	jnot g0382(.din(n453),.dout(n454),.clk(gclk));
	jor g0383(.dina(w_n414_0[1]),.dinb(w_n73_1[2]),.dout(n455),.clk(gclk));
	jand g0384(.dina(n455),.dinb(n454),.dout(n456),.clk(gclk));
	jor g0385(.dina(w_n456_0[1]),.dinb(n451),.dout(n457),.clk(gclk));
	jnot g0386(.din(w_n435_0[0]),.dout(n458),.clk(gclk));
	jor g0387(.dina(n458),.dinb(w_n430_0[0]),.dout(n459),.clk(gclk));
	jand g0388(.dina(n459),.dinb(w_n172_1[2]),.dout(n460),.clk(gclk));
	jor g0389(.dina(n460),.dinb(w_n356_0[2]),.dout(n461),.clk(gclk));
	jor g0390(.dina(n461),.dinb(w_n428_0[0]),.dout(n462),.clk(gclk));
	jor g0391(.dina(n462),.dinb(w_G179_2[0]),.dout(n463),.clk(gclk));
	jand g0392(.dina(n463),.dinb(w_n457_0[1]),.dout(n464),.clk(gclk));
	jand g0393(.dina(n464),.dinb(n440),.dout(n465),.clk(gclk));
	jand g0394(.dina(w_n439_0[1]),.dinb(w_G190_2[2]),.dout(n466),.clk(gclk));
	jnot g0395(.din(n466),.dout(n467),.clk(gclk));
	jnot g0396(.din(w_n456_0[0]),.dout(n468),.clk(gclk));
	jand g0397(.dina(n468),.dinb(w_n450_0[0]),.dout(n469),.clk(gclk));
	jor g0398(.dina(w_n439_0[0]),.dinb(w_n388_2[0]),.dout(n470),.clk(gclk));
	jand g0399(.dina(n470),.dinb(n469),.dout(n471),.clk(gclk));
	jand g0400(.dina(n471),.dinb(n467),.dout(n472),.clk(gclk));
	jor g0401(.dina(w_n472_0[1]),.dinb(w_n465_0[1]),.dout(n473),.clk(gclk));
	jand g0402(.dina(w_n168_1[2]),.dinb(w_G232_0[1]),.dout(n474),.clk(gclk));
	jand g0403(.dina(n474),.dinb(w_n354_0[1]),.dout(n475),.clk(gclk));
	jand g0404(.dina(w_n173_1[0]),.dinb(w_G226_0[1]),.dout(n476),.clk(gclk));
	jand g0405(.dina(w_n177_0[1]),.dinb(w_G223_0[0]),.dout(n477),.clk(gclk));
	jor g0406(.dina(n477),.dinb(w_n370_0[0]),.dout(n478),.clk(gclk));
	jor g0407(.dina(n478),.dinb(n476),.dout(n479),.clk(gclk));
	jand g0408(.dina(n479),.dinb(w_n172_1[1]),.dout(n480),.clk(gclk));
	jor g0409(.dina(n480),.dinb(w_n356_0[1]),.dout(n481),.clk(gclk));
	jor g0410(.dina(n481),.dinb(n475),.dout(n482),.clk(gclk));
	jnot g0411(.din(w_n482_0[2]),.dout(n483),.clk(gclk));
	jor g0412(.dina(w_n483_0[1]),.dinb(w_G169_1[2]),.dout(n484),.clk(gclk));
	jnot g0413(.din(w_G159_3[2]),.dout(n485),.clk(gclk));
	jnot g0414(.din(w_n445_0[0]),.dout(n486),.clk(gclk));
	jor g0415(.dina(n486),.dinb(n485),.dout(n487),.clk(gclk));
	jxor g0416(.dina(w_G68_4[1]),.dinb(w_G58_4[1]),.dout(n488),.clk(gclk));
	jor g0417(.dina(n488),.dinb(w_n151_3[0]),.dout(n489),.clk(gclk));
	jand g0418(.dina(w_n441_0[0]),.dinb(w_G68_4[0]),.dout(n490),.clk(gclk));
	jnot g0419(.din(n490),.dout(n491),.clk(gclk));
	jand g0420(.dina(n491),.dinb(n489),.dout(n492),.clk(gclk));
	jand g0421(.dina(n492),.dinb(n487),.dout(n493),.clk(gclk));
	jor g0422(.dina(n493),.dinb(w_n261_0[1]),.dout(n494),.clk(gclk));
	jnot g0423(.din(w_n494_0[1]),.dout(n495),.clk(gclk));
	jand g0424(.dina(w_n452_0[0]),.dinb(w_n74_1[2]),.dout(n496),.clk(gclk));
	jnot g0425(.din(n496),.dout(n497),.clk(gclk));
	jor g0426(.dina(w_n414_0[0]),.dinb(w_n74_1[1]),.dout(n498),.clk(gclk));
	jand g0427(.dina(n498),.dinb(n497),.dout(n499),.clk(gclk));
	jor g0428(.dina(w_n499_0[1]),.dinb(n495),.dout(n500),.clk(gclk));
	jor g0429(.dina(w_n482_0[1]),.dinb(w_G179_1[2]),.dout(n501),.clk(gclk));
	jand g0430(.dina(n501),.dinb(w_n500_0[1]),.dout(n502),.clk(gclk));
	jand g0431(.dina(n502),.dinb(n484),.dout(n503),.clk(gclk));
	jor g0432(.dina(w_n483_0[0]),.dinb(w_n388_1[2]),.dout(n504),.clk(gclk));
	jnot g0433(.din(w_n499_0[0]),.dout(n505),.clk(gclk));
	jand g0434(.dina(n505),.dinb(w_n494_0[0]),.dout(n506),.clk(gclk));
	jnot g0435(.din(w_G190_2[1]),.dout(n507),.clk(gclk));
	jor g0436(.dina(w_n482_0[0]),.dinb(w_n507_2[1]),.dout(n508),.clk(gclk));
	jand g0437(.dina(n508),.dinb(n506),.dout(n509),.clk(gclk));
	jand g0438(.dina(n509),.dinb(n504),.dout(n510),.clk(gclk));
	jor g0439(.dina(n510),.dinb(w_n503_0[2]),.dout(n511),.clk(gclk));
	jor g0440(.dina(w_n511_0[1]),.dinb(w_n473_0[1]),.dout(n512),.clk(gclk));
	jor g0441(.dina(w_n512_0[1]),.dinb(w_n426_0[1]),.dout(n513),.clk(gclk));
	jor g0442(.dina(n513),.dinb(w_n395_0[1]),.dout(n514),.clk(gclk));
	jnot g0443(.din(w_n514_1[1]),.dout(n515),.clk(gclk));
	jand g0444(.dina(n515),.dinb(w_n351_0[1]),.dout(w_dff_A_iZwOYoxD1_2),.clk(gclk));
	jnot g0445(.din(w_n213_0[0]),.dout(n517),.clk(gclk));
	jor g0446(.dina(w_n212_0[2]),.dinb(w_G179_1[1]),.dout(n518),.clk(gclk));
	jand g0447(.dina(n518),.dinb(w_n224_0[2]),.dout(n519),.clk(gclk));
	jand g0448(.dina(n519),.dinb(n517),.dout(n520),.clk(gclk));
	jnot g0449(.din(w_n238_0[0]),.dout(n521),.clk(gclk));
	jor g0450(.dina(w_n234_0[2]),.dinb(w_n388_1[1]),.dout(n522),.clk(gclk));
	jand g0451(.dina(n522),.dinb(w_n225_0[0]),.dout(n523),.clk(gclk));
	jand g0452(.dina(n523),.dinb(n521),.dout(n524),.clk(gclk));
	jor g0453(.dina(n524),.dinb(w_n520_0[1]),.dout(n525),.clk(gclk));
	jnot g0454(.din(w_n256_0[0]),.dout(n526),.clk(gclk));
	jor g0455(.dina(w_n255_0[2]),.dinb(w_G169_1[1]),.dout(n527),.clk(gclk));
	jand g0456(.dina(n527),.dinb(w_n292_0[1]),.dout(n528),.clk(gclk));
	jand g0457(.dina(n528),.dinb(n526),.dout(n529),.clk(gclk));
	jnot g0458(.din(w_n283_0[0]),.dout(n530),.clk(gclk));
	jor g0459(.dina(w_n279_0[2]),.dinb(w_n507_2[0]),.dout(n531),.clk(gclk));
	jand g0460(.dina(n531),.dinb(w_n272_0[0]),.dout(n532),.clk(gclk));
	jand g0461(.dina(n532),.dinb(n530),.dout(n533),.clk(gclk));
	jor g0462(.dina(w_n533_0[1]),.dinb(n529),.dout(n534),.clk(gclk));
	jnot g0463(.din(w_n309_0[0]),.dout(n535),.clk(gclk));
	jor g0464(.dina(w_n308_0[2]),.dinb(w_n388_1[0]),.dout(n536),.clk(gclk));
	jand g0465(.dina(n536),.dinb(w_n344_0[0]),.dout(n537),.clk(gclk));
	jand g0466(.dina(n537),.dinb(n535),.dout(n538),.clk(gclk));
	jor g0467(.dina(w_n330_0[1]),.dinb(w_G179_1[0]),.dout(n539),.clk(gclk));
	jand g0468(.dina(n539),.dinb(w_n323_0[1]),.dout(n540),.clk(gclk));
	jand g0469(.dina(n540),.dinb(w_n334_0[0]),.dout(n541),.clk(gclk));
	jor g0470(.dina(w_n541_0[1]),.dinb(n538),.dout(n542),.clk(gclk));
	jor g0471(.dina(w_n542_0[1]),.dinb(w_n534_0[1]),.dout(n543),.clk(gclk));
	jor g0472(.dina(w_n543_0[1]),.dinb(n525),.dout(n544),.clk(gclk));
	jor g0473(.dina(w_n544_0[1]),.dinb(w_n192_0[1]),.dout(n545),.clk(gclk));
	jor g0474(.dina(w_n543_0[0]),.dinb(w_n237_0[1]),.dout(n546),.clk(gclk));
	jor g0475(.dina(w_n347_0[0]),.dinb(w_n533_0[0]),.dout(n547),.clk(gclk));
	jand g0476(.dina(n547),.dinb(w_n282_0[0]),.dout(n548),.clk(gclk));
	jand g0477(.dina(w_n548_0[1]),.dinb(n546),.dout(n549),.clk(gclk));
	jand g0478(.dina(n549),.dinb(n545),.dout(n550),.clk(gclk));
	jor g0479(.dina(w_n550_0[1]),.dinb(w_n514_1[0]),.dout(n551),.clk(gclk));
	jnot g0480(.din(w_n551_0[1]),.dout(n552),.clk(gclk));
	jnot g0481(.din(w_n472_0[0]),.dout(n553),.clk(gclk));
	jand g0482(.dina(w_n503_0[1]),.dinb(n553),.dout(n554),.clk(gclk));
	jnot g0483(.din(n554),.dout(n555),.clk(gclk));
	jnot g0484(.din(w_n465_0[0]),.dout(n556),.clk(gclk));
	jnot g0485(.din(w_n420_0[0]),.dout(n557),.clk(gclk));
	jor g0486(.dina(w_n425_0[0]),.dinb(w_n387_0[1]),.dout(n558),.clk(gclk));
	jand g0487(.dina(n558),.dinb(n557),.dout(n559),.clk(gclk));
	jor g0488(.dina(w_n559_0[1]),.dinb(w_n512_0[0]),.dout(n560),.clk(gclk));
	jand g0489(.dina(n560),.dinb(n556),.dout(n561),.clk(gclk));
	jand g0490(.dina(n561),.dinb(n555),.dout(n562),.clk(gclk));
	jnot g0491(.din(w_n562_0[1]),.dout(n563),.clk(gclk));
	jor g0492(.dina(n563),.dinb(n552),.dout(w_dff_A_UNMIhmVW3_2),.clk(gclk));
	jand g0493(.dina(w_n143_0[0]),.dinb(w_G213_0[2]),.dout(n565),.clk(gclk));
	jand g0494(.dina(n565),.dinb(w_n151_2[2]),.dout(n566),.clk(gclk));
	jand g0495(.dina(w_n566_1[1]),.dinb(w_G343_0[1]),.dout(n567),.clk(gclk));
	jor g0496(.dina(w_n567_5[1]),.dinb(w_n237_0[0]),.dout(n568),.clk(gclk));
	jnot g0497(.din(n568),.dout(n569),.clk(gclk));
	jnot g0498(.din(w_n192_0[0]),.dout(n570),.clk(gclk));
	jnot g0499(.din(w_n567_5[0]),.dout(n571),.clk(gclk));
	jand g0500(.dina(w_n571_2[1]),.dinb(w_n570_0[1]),.dout(n572),.clk(gclk));
	jand g0501(.dina(w_n572_0[2]),.dinb(w_n242_0[1]),.dout(n573),.clk(gclk));
	jor g0502(.dina(w_n573_0[1]),.dinb(w_n569_0[1]),.dout(n574),.clk(gclk));
	jand g0503(.dina(w_n567_4[2]),.dinb(w_n161_0[0]),.dout(n575),.clk(gclk));
	jxor g0504(.dina(n575),.dinb(w_n198_0[1]),.dout(n576),.clk(gclk));
	jand g0505(.dina(w_n576_0[2]),.dinb(w_G330_0[2]),.dout(n577),.clk(gclk));
	jand g0506(.dina(w_n567_4[1]),.dinb(w_n224_0[1]),.dout(n578),.clk(gclk));
	jxor g0507(.dina(n578),.dinb(w_n242_0[0]),.dout(n579),.clk(gclk));
	jand g0508(.dina(w_n579_1[1]),.dinb(w_n577_0[1]),.dout(n580),.clk(gclk));
	jor g0509(.dina(w_n580_0[2]),.dinb(w_n574_0[1]),.dout(w_dff_A_74kv90FR7_2),.clk(gclk));
	jand g0510(.dina(w_n91_1[1]),.dinb(w_n163_0[2]),.dout(n582),.clk(gclk));
	jand g0511(.dina(w_n582_0[1]),.dinb(w_n118_0[1]),.dout(n583),.clk(gclk));
	jor g0512(.dina(w_n567_4[0]),.dinb(w_n550_0[0]),.dout(n584),.clk(gclk));
	jnot g0513(.din(w_n198_0[0]),.dout(n585),.clk(gclk));
	jor g0514(.dina(w_n544_0[0]),.dinb(n585),.dout(n586),.clk(gclk));
	jand g0515(.dina(w_n571_2[0]),.dinb(n586),.dout(n587),.clk(gclk));
	jnot g0516(.din(w_n190_0[0]),.dout(n588),.clk(gclk));
	jand g0517(.dina(w_n308_0[1]),.dinb(w_n255_0[1]),.dout(n589),.clk(gclk));
	jand g0518(.dina(n589),.dinb(n588),.dout(n590),.clk(gclk));
	jand g0519(.dina(n590),.dinb(w_n234_0[1]),.dout(n591),.clk(gclk));
	jand g0520(.dina(w_n279_0[1]),.dinb(w_n189_1[0]),.dout(n592),.clk(gclk));
	jand g0521(.dina(n592),.dinb(w_n330_0[0]),.dout(n593),.clk(gclk));
	jand g0522(.dina(n593),.dinb(w_n186_0[1]),.dout(n594),.clk(gclk));
	jand g0523(.dina(n594),.dinb(w_n212_0[1]),.dout(n595),.clk(gclk));
	jor g0524(.dina(n595),.dinb(w_n571_1[2]),.dout(n596),.clk(gclk));
	jor g0525(.dina(n596),.dinb(n591),.dout(n597),.clk(gclk));
	jand g0526(.dina(n597),.dinb(w_G330_0[1]),.dout(n598),.clk(gclk));
	jnot g0527(.din(w_n598_0[1]),.dout(n599),.clk(gclk));
	jor g0528(.dina(n599),.dinb(n587),.dout(n600),.clk(gclk));
	jand g0529(.dina(w_n600_1[2]),.dinb(w_n584_0[1]),.dout(n601),.clk(gclk));
	jnot g0530(.din(w_n601_0[2]),.dout(n602),.clk(gclk));
	jand g0531(.dina(w_n602_0[1]),.dinb(w_n142_1[0]),.dout(n603),.clk(gclk));
	jnot g0532(.din(w_n582_0[0]),.dout(n604),.clk(gclk));
	jand g0533(.dina(w_n259_0[0]),.dinb(w_n105_0[2]),.dout(n605),.clk(gclk));
	jand g0534(.dina(w_n605_0[2]),.dinb(w_G1_0[2]),.dout(n606),.clk(gclk));
	jand g0535(.dina(n606),.dinb(w_n604_2[2]),.dout(n607),.clk(gclk));
	jor g0536(.dina(n607),.dinb(n603),.dout(n608),.clk(gclk));
	jor g0537(.dina(n608),.dinb(w_dff_B_ueFBhWi45_1),.dout(w_dff_A_oGQbtTGb6_2),.clk(gclk));
	jand g0538(.dina(w_G45_0[2]),.dinb(w_G13_0[2]),.dout(n610),.clk(gclk));
	jand g0539(.dina(n610),.dinb(w_n151_2[1]),.dout(n611),.clk(gclk));
	jor g0540(.dina(n611),.dinb(w_n142_0[2]),.dout(n612),.clk(gclk));
	jnot g0541(.din(n612),.dout(n613),.clk(gclk));
	jand g0542(.dina(w_n613_1[2]),.dinb(w_n604_2[1]),.dout(n614),.clk(gclk));
	jnot g0543(.din(w_n614_5[1]),.dout(n615),.clk(gclk));
	jxor g0544(.dina(w_n576_0[1]),.dinb(w_G330_0[0]),.dout(n616),.clk(gclk));
	jand g0545(.dina(n616),.dinb(n615),.dout(n617),.clk(gclk));
	jand g0546(.dina(w_n153_5[1]),.dinb(w_n89_0[0]),.dout(n618),.clk(gclk));
	jand g0547(.dina(w_n618_2[1]),.dinb(w_n151_2[0]),.dout(n619),.clk(gclk));
	jnot g0548(.din(w_n619_0[2]),.dout(n620),.clk(gclk));
	jor g0549(.dina(w_n620_0[2]),.dinb(w_n576_0[0]),.dout(n621),.clk(gclk));
	jand g0550(.dina(w_n507_1[2]),.dinb(w_G20_2[2]),.dout(n622),.clk(gclk));
	jnot g0551(.din(w_n622_0[1]),.dout(n623),.clk(gclk));
	jand g0552(.dina(w_G200_1[1]),.dinb(w_G20_2[1]),.dout(n624),.clk(gclk));
	jnot g0553(.din(w_n624_0[1]),.dout(n625),.clk(gclk));
	jand g0554(.dina(w_G179_0[2]),.dinb(w_G20_2[0]),.dout(n626),.clk(gclk));
	jnot g0555(.din(w_n626_0[2]),.dout(n627),.clk(gclk));
	jand g0556(.dina(n627),.dinb(n625),.dout(n628),.clk(gclk));
	jand g0557(.dina(w_n628_0[1]),.dinb(n623),.dout(n629),.clk(gclk));
	jand g0558(.dina(w_n629_5[1]),.dinb(w_G97_3[0]),.dout(n630),.clk(gclk));
	jnot g0559(.din(w_n630_0[1]),.dout(n631),.clk(gclk));
	jand g0560(.dina(w_n624_0[0]),.dinb(w_n189_0[2]),.dout(n632),.clk(gclk));
	jand g0561(.dina(w_n632_0[1]),.dinb(w_G190_2[0]),.dout(n633),.clk(gclk));
	jand g0562(.dina(w_n633_6[1]),.dinb(w_G87_2[1]),.dout(n634),.clk(gclk));
	jnot g0563(.din(w_n634_0[1]),.dout(n635),.clk(gclk));
	jand g0564(.dina(n635),.dinb(n631),.dout(n636),.clk(gclk));
	jand g0565(.dina(w_n626_0[1]),.dinb(w_n388_0[2]),.dout(n637),.clk(gclk));
	jand g0566(.dina(w_n637_0[1]),.dinb(w_n507_1[1]),.dout(n638),.clk(gclk));
	jand g0567(.dina(w_n638_7[1]),.dinb(w_G77_3[0]),.dout(n639),.clk(gclk));
	jand g0568(.dina(w_n628_0[0]),.dinb(w_n622_0[0]),.dout(n640),.clk(gclk));
	jand g0569(.dina(w_n640_7[1]),.dinb(w_G159_3[1]),.dout(n641),.clk(gclk));
	jor g0570(.dina(n641),.dinb(n639),.dout(n642),.clk(gclk));
	jor g0571(.dina(n642),.dinb(w_G33_7[0]),.dout(n643),.clk(gclk));
	jnot g0572(.din(n643),.dout(n644),.clk(gclk));
	jand g0573(.dina(n644),.dinb(n636),.dout(n645),.clk(gclk));
	jand g0574(.dina(w_n637_0[0]),.dinb(w_G190_1[2]),.dout(n646),.clk(gclk));
	jand g0575(.dina(w_n646_7[1]),.dinb(w_G58_4[0]),.dout(n647),.clk(gclk));
	jand g0576(.dina(w_n632_0[0]),.dinb(w_n507_1[0]),.dout(n648),.clk(gclk));
	jand g0577(.dina(w_n648_4[1]),.dinb(w_G107_3[0]),.dout(n649),.clk(gclk));
	jand g0578(.dina(w_n626_0[0]),.dinb(w_G200_1[0]),.dout(n650),.clk(gclk));
	jand g0579(.dina(w_n650_0[1]),.dinb(w_G190_1[1]),.dout(n651),.clk(gclk));
	jand g0580(.dina(w_n651_7[1]),.dinb(w_G50_4[1]),.dout(n652),.clk(gclk));
	jand g0581(.dina(w_n650_0[0]),.dinb(w_n507_0[2]),.dout(n653),.clk(gclk));
	jand g0582(.dina(w_n653_7[1]),.dinb(w_G68_3[2]),.dout(n654),.clk(gclk));
	jor g0583(.dina(n654),.dinb(n652),.dout(n655),.clk(gclk));
	jor g0584(.dina(n655),.dinb(w_n649_0[1]),.dout(n656),.clk(gclk));
	jor g0585(.dina(n656),.dinb(n647),.dout(n657),.clk(gclk));
	jnot g0586(.din(n657),.dout(n658),.clk(gclk));
	jand g0587(.dina(n658),.dinb(n645),.dout(n659),.clk(gclk));
	jnot g0588(.din(n659),.dout(n660),.clk(gclk));
	jand g0589(.dina(w_n646_7[0]),.dinb(w_G322_0[2]),.dout(n661),.clk(gclk));
	jand g0590(.dina(w_n633_6[0]),.dinb(w_G303_2[1]),.dout(n662),.clk(gclk));
	jand g0591(.dina(w_n629_5[0]),.dinb(w_G294_3[0]),.dout(n663),.clk(gclk));
	jor g0592(.dina(n663),.dinb(n662),.dout(n664),.clk(gclk));
	jand g0593(.dina(w_n651_7[0]),.dinb(w_G326_0[1]),.dout(n665),.clk(gclk));
	jor g0594(.dina(n665),.dinb(n664),.dout(n666),.clk(gclk));
	jand g0595(.dina(w_n640_7[0]),.dinb(G329),.dout(n667),.clk(gclk));
	jor g0596(.dina(n667),.dinb(w_n153_5[0]),.dout(n668),.clk(gclk));
	jand g0597(.dina(w_n638_7[0]),.dinb(w_G311_1[2]),.dout(n669),.clk(gclk));
	jand g0598(.dina(w_n653_7[0]),.dinb(w_G317_1[1]),.dout(n670),.clk(gclk));
	jor g0599(.dina(n670),.dinb(n669),.dout(n671),.clk(gclk));
	jand g0600(.dina(w_n648_4[0]),.dinb(w_G283_3[1]),.dout(n672),.clk(gclk));
	jor g0601(.dina(n672),.dinb(n671),.dout(n673),.clk(gclk));
	jor g0602(.dina(n673),.dinb(n668),.dout(n674),.clk(gclk));
	jor g0603(.dina(n674),.dinb(n666),.dout(n675),.clk(gclk));
	jor g0604(.dina(n675),.dinb(n661),.dout(n676),.clk(gclk));
	jand g0605(.dina(n676),.dinb(n660),.dout(n677),.clk(gclk));
	jand g0606(.dina(w_n139_0[1]),.dinb(w_G169_1[0]),.dout(n678),.clk(gclk));
	jor g0607(.dina(n678),.dinb(w_n375_0[0]),.dout(n679),.clk(gclk));
	jnot g0608(.din(n679),.dout(n680),.clk(gclk));
	jor g0609(.dina(w_n680_4[1]),.dinb(n677),.dout(n681),.clk(gclk));
	jand g0610(.dina(w_n680_4[0]),.dinb(w_n620_0[1]),.dout(n682),.clk(gclk));
	jor g0611(.dina(w_n134_0[0]),.dinb(w_n352_1[0]),.dout(n683),.clk(gclk));
	jand g0612(.dina(w_n91_1[0]),.dinb(w_G33_6[2]),.dout(n684),.clk(gclk));
	jnot g0613(.din(w_n684_0[2]),.dout(n685),.clk(gclk));
	jand g0614(.dina(w_n118_0[0]),.dinb(w_n352_0[2]),.dout(n686),.clk(gclk));
	jor g0615(.dina(n686),.dinb(w_n685_0[1]),.dout(n687),.clk(gclk));
	jnot g0616(.din(n687),.dout(n688),.clk(gclk));
	jand g0617(.dina(n688),.dinb(n683),.dout(n689),.clk(gclk));
	jnot g0618(.din(w_n91_0[2]),.dout(n690),.clk(gclk));
	jand g0619(.dina(w_n690_1[1]),.dinb(w_n105_0[1]),.dout(n691),.clk(gclk));
	jand g0620(.dina(w_n91_0[1]),.dinb(w_n153_4[2]),.dout(n692),.clk(gclk));
	jand g0621(.dina(w_n692_0[1]),.dinb(w_G355_0),.dout(n693),.clk(gclk));
	jor g0622(.dina(n693),.dinb(n691),.dout(n694),.clk(gclk));
	jor g0623(.dina(w_dff_B_QI4QLR1u6_0),.dinb(n689),.dout(n695),.clk(gclk));
	jand g0624(.dina(n695),.dinb(w_n682_0[1]),.dout(n696),.clk(gclk));
	jnot g0625(.din(n696),.dout(n697),.clk(gclk));
	jand g0626(.dina(w_dff_B_P6gvEx497_0),.dinb(n681),.dout(n698),.clk(gclk));
	jand g0627(.dina(w_dff_B_pETUV4B08_0),.dinb(n621),.dout(n699),.clk(gclk));
	jand g0628(.dina(n699),.dinb(w_n614_5[0]),.dout(n700),.clk(gclk));
	jor g0629(.dina(n700),.dinb(w_dff_B_DNikSduU6_1),.dout(G396_fa_),.clk(gclk));
	jand g0630(.dina(w_n567_3[2]),.dinb(w_n383_0[0]),.dout(n702),.clk(gclk));
	jxor g0631(.dina(n702),.dinb(w_n394_0[0]),.dout(n703),.clk(gclk));
	jnot g0632(.din(w_n703_1[1]),.dout(n704),.clk(gclk));
	jand g0633(.dina(w_n704_0[1]),.dinb(w_n618_2[0]),.dout(n705),.clk(gclk));
	jnot g0634(.din(n705),.dout(n706),.clk(gclk));
	jand g0635(.dina(w_n653_6[2]),.dinb(w_G150_3[0]),.dout(n707),.clk(gclk));
	jand g0636(.dina(w_n651_6[2]),.dinb(w_G137_1[2]),.dout(n708),.clk(gclk));
	jand g0637(.dina(w_n633_5[2]),.dinb(w_G50_4[0]),.dout(n709),.clk(gclk));
	jor g0638(.dina(n709),.dinb(n708),.dout(n710),.clk(gclk));
	jand g0639(.dina(w_n646_6[2]),.dinb(w_G143_2[1]),.dout(n711),.clk(gclk));
	jor g0640(.dina(n711),.dinb(n710),.dout(n712),.clk(gclk));
	jor g0641(.dina(n712),.dinb(n707),.dout(n713),.clk(gclk));
	jand g0642(.dina(w_n638_6[2]),.dinb(w_G159_3[0]),.dout(n714),.clk(gclk));
	jand g0643(.dina(w_n640_6[2]),.dinb(w_G132_1[1]),.dout(n715),.clk(gclk));
	jor g0644(.dina(n715),.dinb(n714),.dout(n716),.clk(gclk));
	jand g0645(.dina(w_n629_4[2]),.dinb(w_G58_3[2]),.dout(n717),.clk(gclk));
	jand g0646(.dina(w_n648_3[2]),.dinb(w_G68_3[1]),.dout(n718),.clk(gclk));
	jor g0647(.dina(w_n718_0[1]),.dinb(n717),.dout(n719),.clk(gclk));
	jor g0648(.dina(n719),.dinb(w_G33_6[1]),.dout(n720),.clk(gclk));
	jor g0649(.dina(n720),.dinb(n716),.dout(n721),.clk(gclk));
	jor g0650(.dina(n721),.dinb(n713),.dout(n722),.clk(gclk));
	jand g0651(.dina(w_n653_6[1]),.dinb(w_G283_3[0]),.dout(n723),.clk(gclk));
	jand g0652(.dina(w_n640_6[1]),.dinb(w_G311_1[1]),.dout(n724),.clk(gclk));
	jor g0653(.dina(n724),.dinb(n723),.dout(n725),.clk(gclk));
	jand g0654(.dina(w_n633_5[1]),.dinb(w_G107_2[2]),.dout(n726),.clk(gclk));
	jor g0655(.dina(n726),.dinb(w_n630_0[0]),.dout(n727),.clk(gclk));
	jor g0656(.dina(n727),.dinb(n725),.dout(n728),.clk(gclk));
	jand g0657(.dina(w_n646_6[1]),.dinb(w_G294_2[2]),.dout(n729),.clk(gclk));
	jand g0658(.dina(w_n638_6[1]),.dinb(w_G116_4[0]),.dout(n730),.clk(gclk));
	jor g0659(.dina(n730),.dinb(n729),.dout(n731),.clk(gclk));
	jand g0660(.dina(w_n651_6[1]),.dinb(w_G303_2[0]),.dout(n732),.clk(gclk));
	jand g0661(.dina(w_n648_3[1]),.dinb(w_G87_2[0]),.dout(n733),.clk(gclk));
	jor g0662(.dina(w_n733_0[1]),.dinb(n732),.dout(n734),.clk(gclk));
	jor g0663(.dina(n734),.dinb(n731),.dout(n735),.clk(gclk));
	jor g0664(.dina(n735),.dinb(n728),.dout(n736),.clk(gclk));
	jor g0665(.dina(n736),.dinb(w_n153_4[1]),.dout(n737),.clk(gclk));
	jand g0666(.dina(n737),.dinb(n722),.dout(n738),.clk(gclk));
	jor g0667(.dina(n738),.dinb(w_n680_3[2]),.dout(n739),.clk(gclk));
	jnot g0668(.din(w_n618_1[2]),.dout(n740),.clk(gclk));
	jand g0669(.dina(w_n680_3[1]),.dinb(n740),.dout(n741),.clk(gclk));
	jand g0670(.dina(w_n741_1[1]),.dinb(w_n72_0[1]),.dout(n742),.clk(gclk));
	jnot g0671(.din(n742),.dout(n743),.clk(gclk));
	jand g0672(.dina(n743),.dinb(n739),.dout(n744),.clk(gclk));
	jand g0673(.dina(n744),.dinb(w_n614_4[2]),.dout(n745),.clk(gclk));
	jand g0674(.dina(n745),.dinb(n706),.dout(n746),.clk(gclk));
	jnot g0675(.din(n746),.dout(n747),.clk(gclk));
	jor g0676(.dina(w_n584_0[0]),.dinb(w_n395_0[0]),.dout(n748),.clk(gclk));
	jand g0677(.dina(w_n350_0[0]),.dinb(w_n570_0[0]),.dout(n749),.clk(gclk));
	jand g0678(.dina(w_n349_0[0]),.dinb(w_n520_0[0]),.dout(n750),.clk(gclk));
	jnot g0679(.din(w_n548_0[0]),.dout(n751),.clk(gclk));
	jor g0680(.dina(n751),.dinb(n750),.dout(n752),.clk(gclk));
	jor g0681(.dina(n752),.dinb(n749),.dout(n753),.clk(gclk));
	jand g0682(.dina(w_n571_1[1]),.dinb(n753),.dout(n754),.clk(gclk));
	jor g0683(.dina(w_n703_1[0]),.dinb(w_n754_0[1]),.dout(n755),.clk(gclk));
	jand g0684(.dina(n755),.dinb(w_n748_0[1]),.dout(n756),.clk(gclk));
	jxor g0685(.dina(n756),.dinb(w_n600_1[1]),.dout(n757),.clk(gclk));
	jor g0686(.dina(n757),.dinb(w_n614_4[1]),.dout(n758),.clk(gclk));
	jand g0687(.dina(n758),.dinb(n747),.dout(n759),.clk(gclk));
	jnot g0688(.din(w_n759_0[1]),.dout(G384_fa_),.clk(gclk));
	jnot g0689(.din(w_n90_0[1]),.dout(n761),.clk(gclk));
	jand g0690(.dina(w_n112_0[0]),.dinb(n761),.dout(n762),.clk(gclk));
	jnot g0691(.din(w_n566_1[0]),.dout(n763),.clk(gclk));
	jand g0692(.dina(n763),.dinb(w_n503_0[0]),.dout(n764),.clk(gclk));
	jand g0693(.dina(w_n566_0[2]),.dinb(w_n500_0[0]),.dout(n765),.clk(gclk));
	jxor g0694(.dina(n765),.dinb(w_n511_0[0]),.dout(n766),.clk(gclk));
	jnot g0695(.din(w_n766_0[1]),.dout(n767),.clk(gclk));
	jor g0696(.dina(w_n567_3[1]),.dinb(w_n559_0[0]),.dout(n768),.clk(gclk));
	jnot g0697(.din(n768),.dout(n769),.clk(gclk));
	jand g0698(.dina(w_n567_3[0]),.dinb(w_n417_0[0]),.dout(n770),.clk(gclk));
	jxor g0699(.dina(n770),.dinb(w_n426_0[0]),.dout(n771),.clk(gclk));
	jnot g0700(.din(w_n771_1[1]),.dout(n772),.clk(gclk));
	jand g0701(.dina(w_n772_0[1]),.dinb(w_n703_0[2]),.dout(n773),.clk(gclk));
	jand g0702(.dina(w_n773_0[1]),.dinb(w_n754_0[0]),.dout(n774),.clk(gclk));
	jor g0703(.dina(n774),.dinb(n769),.dout(n775),.clk(gclk));
	jand g0704(.dina(w_n775_0[1]),.dinb(w_n767_1[1]),.dout(n776),.clk(gclk));
	jor g0705(.dina(n776),.dinb(n764),.dout(n777),.clk(gclk));
	jand g0706(.dina(w_n773_0[0]),.dinb(w_n767_1[0]),.dout(n778),.clk(gclk));
	jxor g0707(.dina(n778),.dinb(w_n514_0[2]),.dout(n779),.clk(gclk));
	jor g0708(.dina(n779),.dinb(w_n600_1[0]),.dout(n780),.clk(gclk));
	jor g0709(.dina(w_n567_2[2]),.dinb(w_n551_0[0]),.dout(n781),.clk(gclk));
	jand g0710(.dina(n781),.dinb(w_n562_0[0]),.dout(n782),.clk(gclk));
	jxor g0711(.dina(w_n782_0[1]),.dinb(n780),.dout(n783),.clk(gclk));
	jxor g0712(.dina(n783),.dinb(w_n777_0[1]),.dout(n784),.clk(gclk));
	jand g0713(.dina(n784),.dinb(n762),.dout(n785),.clk(gclk));
	jor g0714(.dina(w_n75_1[0]),.dinb(w_n74_1[0]),.dout(n786),.clk(gclk));
	jand g0715(.dina(n786),.dinb(w_G77_2[2]),.dout(n787),.clk(gclk));
	jor g0716(.dina(n787),.dinb(w_n73_1[1]),.dout(n788),.clk(gclk));
	jand g0717(.dina(w_G58_3[1]),.dinb(w_G50_3[2]),.dout(n789),.clk(gclk));
	jor g0718(.dina(n789),.dinb(w_G68_3[0]),.dout(n790),.clk(gclk));
	jand g0719(.dina(n790),.dinb(w_n90_0[0]),.dout(n791),.clk(gclk));
	jand g0720(.dina(n791),.dinb(n788),.dout(n792),.clk(gclk));
	jand g0721(.dina(w_n312_0[0]),.dinb(w_n120_0[0]),.dout(n793),.clk(gclk));
	jand g0722(.dina(n793),.dinb(w_G116_3[2]),.dout(n794),.clk(gclk));
	jor g0723(.dina(n794),.dinb(n792),.dout(n795),.clk(gclk));
	jor g0724(.dina(w_dff_B_Q2OW7rOi7_0),.dinb(n785),.dout(w_dff_A_a1Iu7cw04_2),.clk(gclk));
	jand g0725(.dina(w_n567_2[1]),.dinb(w_n292_0[0]),.dout(n797),.clk(gclk));
	jxor g0726(.dina(n797),.dinb(w_n534_0[0]),.dout(n798),.clk(gclk));
	jand g0727(.dina(w_n798_0[1]),.dinb(w_n619_0[1]),.dout(n799),.clk(gclk));
	jnot g0728(.din(n799),.dout(n800),.clk(gclk));
	jand g0729(.dina(w_n684_0[1]),.dinb(w_n126_0[0]),.dout(n801),.clk(gclk));
	jnot g0730(.din(w_n682_0[0]),.dout(n802),.clk(gclk));
	jand g0731(.dina(w_n690_1[0]),.dinb(w_G87_1[2]),.dout(n803),.clk(gclk));
	jor g0732(.dina(n803),.dinb(w_n802_0[2]),.dout(n804),.clk(gclk));
	jor g0733(.dina(n804),.dinb(n801),.dout(n805),.clk(gclk));
	jand g0734(.dina(n805),.dinb(w_n614_4[0]),.dout(n806),.clk(gclk));
	jand g0735(.dina(w_n646_6[0]),.dinb(w_G303_1[2]),.dout(n807),.clk(gclk));
	jand g0736(.dina(w_n638_6[0]),.dinb(w_G283_2[2]),.dout(n808),.clk(gclk));
	jor g0737(.dina(n808),.dinb(n807),.dout(n809),.clk(gclk));
	jand g0738(.dina(w_n651_6[0]),.dinb(w_G311_1[0]),.dout(n810),.clk(gclk));
	jand g0739(.dina(w_n633_5[0]),.dinb(w_G116_3[1]),.dout(n811),.clk(gclk));
	jor g0740(.dina(n811),.dinb(n810),.dout(n812),.clk(gclk));
	jand g0741(.dina(w_n653_6[0]),.dinb(w_G294_2[1]),.dout(n813),.clk(gclk));
	jand g0742(.dina(w_n640_6[0]),.dinb(w_G317_1[0]),.dout(n814),.clk(gclk));
	jor g0743(.dina(n814),.dinb(n813),.dout(n815),.clk(gclk));
	jand g0744(.dina(w_n629_4[1]),.dinb(w_G107_2[1]),.dout(n816),.clk(gclk));
	jand g0745(.dina(w_n648_3[0]),.dinb(w_G97_2[2]),.dout(n817),.clk(gclk));
	jor g0746(.dina(w_n817_0[1]),.dinb(n816),.dout(n818),.clk(gclk));
	jor g0747(.dina(n818),.dinb(n815),.dout(n819),.clk(gclk));
	jor g0748(.dina(n819),.dinb(n812),.dout(n820),.clk(gclk));
	jor g0749(.dina(n820),.dinb(n809),.dout(n821),.clk(gclk));
	jand g0750(.dina(n821),.dinb(w_G33_6[0]),.dout(n822),.clk(gclk));
	jand g0751(.dina(w_n638_5[2]),.dinb(w_G50_3[1]),.dout(n823),.clk(gclk));
	jand g0752(.dina(w_n640_5[2]),.dinb(w_G137_1[1]),.dout(n824),.clk(gclk));
	jor g0753(.dina(n824),.dinb(n823),.dout(n825),.clk(gclk));
	jand g0754(.dina(w_n651_5[2]),.dinb(w_G143_2[0]),.dout(n826),.clk(gclk));
	jand g0755(.dina(w_n653_5[2]),.dinb(w_G159_2[2]),.dout(n827),.clk(gclk));
	jor g0756(.dina(n827),.dinb(n826),.dout(n828),.clk(gclk));
	jand g0757(.dina(w_n633_4[2]),.dinb(w_G58_3[0]),.dout(n829),.clk(gclk));
	jand g0758(.dina(w_n629_4[0]),.dinb(w_G68_2[2]),.dout(n830),.clk(gclk));
	jor g0759(.dina(w_n830_0[1]),.dinb(n829),.dout(n831),.clk(gclk));
	jand g0760(.dina(w_n646_5[2]),.dinb(w_G150_2[2]),.dout(n832),.clk(gclk));
	jand g0761(.dina(w_n648_2[2]),.dinb(w_G77_2[1]),.dout(n833),.clk(gclk));
	jor g0762(.dina(w_n833_0[1]),.dinb(n832),.dout(n834),.clk(gclk));
	jor g0763(.dina(n834),.dinb(n831),.dout(n835),.clk(gclk));
	jor g0764(.dina(n835),.dinb(n828),.dout(n836),.clk(gclk));
	jor g0765(.dina(n836),.dinb(n825),.dout(n837),.clk(gclk));
	jand g0766(.dina(n837),.dinb(w_n153_4[0]),.dout(n838),.clk(gclk));
	jor g0767(.dina(n838),.dinb(n822),.dout(n839),.clk(gclk));
	jor g0768(.dina(n839),.dinb(w_n680_3[0]),.dout(n840),.clk(gclk));
	jand g0769(.dina(n840),.dinb(n806),.dout(n841),.clk(gclk));
	jand g0770(.dina(n841),.dinb(n800),.dout(n842),.clk(gclk));
	jnot g0771(.din(n842),.dout(n843),.clk(gclk));
	jand g0772(.dina(w_n567_2[0]),.dinb(w_n323_0[0]),.dout(n844),.clk(gclk));
	jxor g0773(.dina(n844),.dinb(w_n542_0[0]),.dout(n845),.clk(gclk));
	jnot g0774(.din(w_n845_0[2]),.dout(n846),.clk(gclk));
	jand g0775(.dina(n846),.dinb(w_n580_0[1]),.dout(n847),.clk(gclk));
	jand g0776(.dina(w_n571_1[0]),.dinb(w_n541_0[0]),.dout(n848),.clk(gclk));
	jand g0777(.dina(w_n579_1[0]),.dinb(w_n348_0[0]),.dout(n849),.clk(gclk));
	jand g0778(.dina(n849),.dinb(w_n572_0[1]),.dout(n850),.clk(gclk));
	jand g0779(.dina(w_n569_0[0]),.dinb(w_n333_0[0]),.dout(n851),.clk(gclk));
	jor g0780(.dina(n851),.dinb(n850),.dout(n852),.clk(gclk));
	jor g0781(.dina(n852),.dinb(n848),.dout(n853),.clk(gclk));
	jxor g0782(.dina(n853),.dinb(w_n798_0[0]),.dout(n854),.clk(gclk));
	jxor g0783(.dina(n854),.dinb(n847),.dout(n855),.clk(gclk));
	jor g0784(.dina(w_n855_0[1]),.dinb(w_n613_1[1]),.dout(n856),.clk(gclk));
	jnot g0785(.din(w_n573_0[0]),.dout(n857),.clk(gclk));
	jor g0786(.dina(w_n579_0[2]),.dinb(w_n572_0[0]),.dout(n858),.clk(gclk));
	jand g0787(.dina(n858),.dinb(n857),.dout(n859),.clk(gclk));
	jxor g0788(.dina(n859),.dinb(w_n577_0[0]),.dout(n860),.clk(gclk));
	jnot g0789(.din(w_n860_0[1]),.dout(n861),.clk(gclk));
	jxor g0790(.dina(w_n580_0[0]),.dinb(w_n574_0[0]),.dout(n862),.clk(gclk));
	jxor g0791(.dina(n862),.dinb(w_n845_0[1]),.dout(n863),.clk(gclk));
	jor g0792(.dina(w_n863_0[2]),.dinb(w_n861_0[1]),.dout(n864),.clk(gclk));
	jand g0793(.dina(n864),.dinb(w_n601_0[1]),.dout(n865),.clk(gclk));
	jor g0794(.dina(w_n855_0[0]),.dinb(w_n604_2[0]),.dout(n866),.clk(gclk));
	jor g0795(.dina(n866),.dinb(n865),.dout(n867),.clk(gclk));
	jand g0796(.dina(n867),.dinb(n856),.dout(n868),.clk(gclk));
	jand g0797(.dina(n868),.dinb(n843),.dout(n869),.clk(gclk));
	jnot g0798(.din(w_n869_0[2]),.dout(w_dff_A_PSsr8Fhy0_1),.clk(gclk));
	jor g0799(.dina(w_n602_0[0]),.dinb(w_n604_1[2]),.dout(n871),.clk(gclk));
	jand g0800(.dina(n871),.dinb(w_n861_0[0]),.dout(n872),.clk(gclk));
	jand g0801(.dina(w_n860_0[0]),.dinb(w_n601_0[0]),.dout(n873),.clk(gclk));
	jand g0802(.dina(w_n873_0[1]),.dinb(w_n613_1[0]),.dout(n874),.clk(gclk));
	jor g0803(.dina(n874),.dinb(w_n614_3[2]),.dout(n875),.clk(gclk));
	jor g0804(.dina(w_n875_0[1]),.dinb(n872),.dout(n876),.clk(gclk));
	jor g0805(.dina(w_n620_0[0]),.dinb(w_n579_0[1]),.dout(n877),.clk(gclk));
	jand g0806(.dina(w_n653_5[1]),.dinb(w_G58_2[2]),.dout(n878),.clk(gclk));
	jand g0807(.dina(w_n638_5[1]),.dinb(w_G68_2[1]),.dout(n879),.clk(gclk));
	jor g0808(.dina(n879),.dinb(w_n817_0[0]),.dout(n880),.clk(gclk));
	jor g0809(.dina(n880),.dinb(w_G33_5[2]),.dout(n881),.clk(gclk));
	jor g0810(.dina(n881),.dinb(n878),.dout(n882),.clk(gclk));
	jnot g0811(.din(n882),.dout(n883),.clk(gclk));
	jand g0812(.dina(w_n629_3[2]),.dinb(w_G87_1[1]),.dout(n884),.clk(gclk));
	jnot g0813(.din(w_n884_0[1]),.dout(n885),.clk(gclk));
	jand g0814(.dina(w_n633_4[1]),.dinb(w_G77_2[0]),.dout(n886),.clk(gclk));
	jnot g0815(.din(n886),.dout(n887),.clk(gclk));
	jand g0816(.dina(w_n887_0[1]),.dinb(n885),.dout(n888),.clk(gclk));
	jand g0817(.dina(w_n646_5[1]),.dinb(w_G50_3[0]),.dout(n889),.clk(gclk));
	jand g0818(.dina(w_n640_5[1]),.dinb(w_G150_2[1]),.dout(n890),.clk(gclk));
	jor g0819(.dina(n890),.dinb(n889),.dout(n891),.clk(gclk));
	jand g0820(.dina(w_n651_5[1]),.dinb(w_G159_2[1]),.dout(n892),.clk(gclk));
	jor g0821(.dina(n892),.dinb(n891),.dout(n893),.clk(gclk));
	jnot g0822(.din(n893),.dout(n894),.clk(gclk));
	jand g0823(.dina(n894),.dinb(n888),.dout(n895),.clk(gclk));
	jand g0824(.dina(n895),.dinb(n883),.dout(n896),.clk(gclk));
	jnot g0825(.din(n896),.dout(n897),.clk(gclk));
	jand g0826(.dina(w_n653_5[0]),.dinb(w_G311_0[2]),.dout(n898),.clk(gclk));
	jand g0827(.dina(w_n633_4[0]),.dinb(w_G294_2[0]),.dout(n899),.clk(gclk));
	jand g0828(.dina(w_n629_3[1]),.dinb(w_G283_2[1]),.dout(n900),.clk(gclk));
	jor g0829(.dina(n900),.dinb(n899),.dout(n901),.clk(gclk));
	jand g0830(.dina(w_n651_5[0]),.dinb(w_G322_0[1]),.dout(n902),.clk(gclk));
	jand g0831(.dina(w_n640_5[0]),.dinb(w_G326_0[0]),.dout(n903),.clk(gclk));
	jor g0832(.dina(n903),.dinb(n902),.dout(n904),.clk(gclk));
	jor g0833(.dina(n904),.dinb(n901),.dout(n905),.clk(gclk));
	jand g0834(.dina(w_n638_5[0]),.dinb(w_G303_1[1]),.dout(n906),.clk(gclk));
	jand g0835(.dina(w_n648_2[1]),.dinb(w_G116_3[0]),.dout(n907),.clk(gclk));
	jor g0836(.dina(n907),.dinb(n906),.dout(n908),.clk(gclk));
	jand g0837(.dina(w_n646_5[0]),.dinb(w_G317_0[2]),.dout(n909),.clk(gclk));
	jor g0838(.dina(n909),.dinb(n908),.dout(n910),.clk(gclk));
	jor g0839(.dina(n910),.dinb(w_n153_3[2]),.dout(n911),.clk(gclk));
	jor g0840(.dina(n911),.dinb(n905),.dout(n912),.clk(gclk));
	jor g0841(.dina(n912),.dinb(n898),.dout(n913),.clk(gclk));
	jand g0842(.dina(n913),.dinb(n897),.dout(n914),.clk(gclk));
	jor g0843(.dina(n914),.dinb(w_n680_2[2]),.dout(n915),.clk(gclk));
	jand g0844(.dina(w_n690_0[2]),.dinb(w_n81_0[2]),.dout(n916),.clk(gclk));
	jnot g0845(.din(n916),.dout(n917),.clk(gclk));
	jnot g0846(.din(w_n605_0[1]),.dout(n918),.clk(gclk));
	jand g0847(.dina(w_n692_0[0]),.dinb(n918),.dout(n919),.clk(gclk));
	jnot g0848(.din(n919),.dout(n920),.clk(gclk));
	jand g0849(.dina(w_n130_0[0]),.dinb(w_G45_0[1]),.dout(n921),.clk(gclk));
	jor g0850(.dina(n921),.dinb(w_n685_0[0]),.dout(n922),.clk(gclk));
	jand g0851(.dina(n922),.dinb(n920),.dout(n923),.clk(gclk));
	jand g0852(.dina(w_G77_1[2]),.dinb(w_G68_2[0]),.dout(n924),.clk(gclk));
	jnot g0853(.din(n924),.dout(n925),.clk(gclk));
	jand g0854(.dina(w_G58_2[1]),.dinb(w_n73_1[0]),.dout(n926),.clk(gclk));
	jand g0855(.dina(n926),.dinb(n925),.dout(n927),.clk(gclk));
	jand g0856(.dina(n927),.dinb(w_n605_0[0]),.dout(n928),.clk(gclk));
	jand g0857(.dina(n928),.dinb(w_n352_0[1]),.dout(n929),.clk(gclk));
	jor g0858(.dina(n929),.dinb(n923),.dout(n930),.clk(gclk));
	jand g0859(.dina(n930),.dinb(n917),.dout(n931),.clk(gclk));
	jor g0860(.dina(n931),.dinb(w_n802_0[1]),.dout(n932),.clk(gclk));
	jand g0861(.dina(n932),.dinb(n915),.dout(n933),.clk(gclk));
	jand g0862(.dina(n933),.dinb(n877),.dout(n934),.clk(gclk));
	jand g0863(.dina(n934),.dinb(w_n614_3[1]),.dout(n935),.clk(gclk));
	jnot g0864(.din(n935),.dout(n936),.clk(gclk));
	jand g0865(.dina(n936),.dinb(n876),.dout(n937),.clk(gclk));
	jnot g0866(.din(w_n937_0[2]),.dout(w_dff_A_6yoiM3mB4_1),.clk(gclk));
	jnot g0867(.din(w_n863_0[1]),.dout(n939),.clk(gclk));
	jnot g0868(.din(w_n873_0[0]),.dout(n940),.clk(gclk));
	jor g0869(.dina(n940),.dinb(n939),.dout(n941),.clk(gclk));
	jor g0870(.dina(n941),.dinb(w_n604_1[1]),.dout(n942),.clk(gclk));
	jor g0871(.dina(w_n875_0[0]),.dinb(w_n863_0[0]),.dout(n943),.clk(gclk));
	jand g0872(.dina(w_n845_0[0]),.dinb(w_n619_0[0]),.dout(n944),.clk(gclk));
	jnot g0873(.din(n944),.dout(n945),.clk(gclk));
	jand g0874(.dina(w_n690_0[1]),.dinb(w_G97_2[1]),.dout(n946),.clk(gclk));
	jand g0875(.dina(w_n684_0[0]),.dinb(w_n137_0[0]),.dout(n947),.clk(gclk));
	jor g0876(.dina(n947),.dinb(w_n802_0[0]),.dout(n948),.clk(gclk));
	jor g0877(.dina(n948),.dinb(n946),.dout(n949),.clk(gclk));
	jand g0878(.dina(w_n653_4[2]),.dinb(w_G50_2[2]),.dout(n950),.clk(gclk));
	jand g0879(.dina(w_n638_4[2]),.dinb(w_G58_2[0]),.dout(n951),.clk(gclk));
	jor g0880(.dina(n951),.dinb(n950),.dout(n952),.clk(gclk));
	jand g0881(.dina(w_n646_4[2]),.dinb(w_G159_2[0]),.dout(n953),.clk(gclk));
	jand g0882(.dina(w_n633_3[2]),.dinb(w_G68_1[2]),.dout(n954),.clk(gclk));
	jor g0883(.dina(n954),.dinb(n953),.dout(n955),.clk(gclk));
	jand g0884(.dina(w_n651_4[2]),.dinb(w_G150_2[0]),.dout(n956),.clk(gclk));
	jor g0885(.dina(n956),.dinb(w_n733_0[0]),.dout(n957),.clk(gclk));
	jand g0886(.dina(w_n640_4[2]),.dinb(w_G143_1[2]),.dout(n958),.clk(gclk));
	jand g0887(.dina(w_n629_3[0]),.dinb(w_G77_1[1]),.dout(n959),.clk(gclk));
	jor g0888(.dina(w_n959_0[1]),.dinb(n958),.dout(n960),.clk(gclk));
	jor g0889(.dina(n960),.dinb(n957),.dout(n961),.clk(gclk));
	jor g0890(.dina(n961),.dinb(n955),.dout(n962),.clk(gclk));
	jor g0891(.dina(n962),.dinb(n952),.dout(n963),.clk(gclk));
	jand g0892(.dina(n963),.dinb(w_n153_3[1]),.dout(n964),.clk(gclk));
	jand g0893(.dina(w_n638_4[1]),.dinb(w_G294_1[2]),.dout(n965),.clk(gclk));
	jand g0894(.dina(w_n640_4[1]),.dinb(w_G322_0[0]),.dout(n966),.clk(gclk));
	jor g0895(.dina(n966),.dinb(n965),.dout(n967),.clk(gclk));
	jand g0896(.dina(w_n646_4[1]),.dinb(w_G311_0[1]),.dout(n968),.clk(gclk));
	jand g0897(.dina(w_n651_4[1]),.dinb(w_G317_0[1]),.dout(n969),.clk(gclk));
	jor g0898(.dina(n969),.dinb(n968),.dout(n970),.clk(gclk));
	jand g0899(.dina(w_n653_4[1]),.dinb(w_G303_1[0]),.dout(n971),.clk(gclk));
	jor g0900(.dina(n971),.dinb(w_n649_0[0]),.dout(n972),.clk(gclk));
	jor g0901(.dina(n972),.dinb(n970),.dout(n973),.clk(gclk));
	jand g0902(.dina(w_n633_3[1]),.dinb(w_G283_2[0]),.dout(n974),.clk(gclk));
	jand g0903(.dina(w_n629_2[2]),.dinb(w_G116_2[2]),.dout(n975),.clk(gclk));
	jor g0904(.dina(n975),.dinb(n974),.dout(n976),.clk(gclk));
	jor g0905(.dina(n976),.dinb(n973),.dout(n977),.clk(gclk));
	jor g0906(.dina(n977),.dinb(n967),.dout(n978),.clk(gclk));
	jand g0907(.dina(n978),.dinb(w_G33_5[1]),.dout(n979),.clk(gclk));
	jor g0908(.dina(n979),.dinb(w_n680_2[1]),.dout(n980),.clk(gclk));
	jor g0909(.dina(n980),.dinb(n964),.dout(n981),.clk(gclk));
	jand g0910(.dina(n981),.dinb(w_n614_3[0]),.dout(n982),.clk(gclk));
	jand g0911(.dina(n982),.dinb(n949),.dout(n983),.clk(gclk));
	jand g0912(.dina(n983),.dinb(n945),.dout(n984),.clk(gclk));
	jnot g0913(.din(n984),.dout(n985),.clk(gclk));
	jand g0914(.dina(n985),.dinb(n943),.dout(n986),.clk(gclk));
	jand g0915(.dina(n986),.dinb(n942),.dout(n987),.clk(gclk));
	jnot g0916(.din(w_n987_0[2]),.dout(w_dff_A_6xuJbluM3_1),.clk(gclk));
	jand g0917(.dina(w_n766_0[0]),.dinb(w_n618_1[1]),.dout(n989),.clk(gclk));
	jnot g0918(.din(n989),.dout(n990),.clk(gclk));
	jand g0919(.dina(w_n651_4[0]),.dinb(w_G128_0[2]),.dout(n991),.clk(gclk));
	jand g0920(.dina(w_n640_4[0]),.dinb(w_G125_0[1]),.dout(n992),.clk(gclk));
	jor g0921(.dina(n992),.dinb(n991),.dout(n993),.clk(gclk));
	jand g0922(.dina(w_n648_2[0]),.dinb(w_G50_2[1]),.dout(n994),.clk(gclk));
	jand g0923(.dina(w_n653_4[0]),.dinb(w_G137_1[0]),.dout(n995),.clk(gclk));
	jor g0924(.dina(n995),.dinb(n994),.dout(n996),.clk(gclk));
	jor g0925(.dina(n996),.dinb(w_G33_5[0]),.dout(n997),.clk(gclk));
	jor g0926(.dina(n997),.dinb(n993),.dout(n998),.clk(gclk));
	jand g0927(.dina(w_n638_4[0]),.dinb(w_G143_1[1]),.dout(n999),.clk(gclk));
	jand g0928(.dina(w_n633_3[0]),.dinb(w_G150_1[2]),.dout(n1000),.clk(gclk));
	jand g0929(.dina(w_n629_2[1]),.dinb(w_G159_1[2]),.dout(n1001),.clk(gclk));
	jand g0930(.dina(w_n646_4[0]),.dinb(w_G132_1[0]),.dout(n1002),.clk(gclk));
	jor g0931(.dina(n1002),.dinb(n1001),.dout(n1003),.clk(gclk));
	jor g0932(.dina(n1003),.dinb(n1000),.dout(n1004),.clk(gclk));
	jor g0933(.dina(n1004),.dinb(n999),.dout(n1005),.clk(gclk));
	jor g0934(.dina(n1005),.dinb(n998),.dout(n1006),.clk(gclk));
	jand g0935(.dina(w_n651_3[2]),.dinb(w_G283_1[2]),.dout(n1007),.clk(gclk));
	jand g0936(.dina(w_n638_3[2]),.dinb(w_G97_2[0]),.dout(n1008),.clk(gclk));
	jor g0937(.dina(n1008),.dinb(w_n153_3[0]),.dout(n1009),.clk(gclk));
	jor g0938(.dina(n1009),.dinb(n1007),.dout(n1010),.clk(gclk));
	jand g0939(.dina(w_n646_3[2]),.dinb(w_G116_2[1]),.dout(n1011),.clk(gclk));
	jand g0940(.dina(w_n640_3[2]),.dinb(w_G294_1[1]),.dout(n1012),.clk(gclk));
	jor g0941(.dina(n1012),.dinb(n1011),.dout(n1013),.clk(gclk));
	jand g0942(.dina(w_n653_3[2]),.dinb(w_G107_2[0]),.dout(n1014),.clk(gclk));
	jor g0943(.dina(n1014),.dinb(w_n634_0[0]),.dout(n1015),.clk(gclk));
	jor g0944(.dina(n1015),.dinb(n1013),.dout(n1016),.clk(gclk));
	jor g0945(.dina(n1016),.dinb(n1010),.dout(n1017),.clk(gclk));
	jor g0946(.dina(n1017),.dinb(w_n959_0[0]),.dout(n1018),.clk(gclk));
	jor g0947(.dina(n1018),.dinb(w_n718_0[0]),.dout(n1019),.clk(gclk));
	jand g0948(.dina(n1019),.dinb(n1006),.dout(n1020),.clk(gclk));
	jor g0949(.dina(n1020),.dinb(w_n680_2[0]),.dout(n1021),.clk(gclk));
	jand g0950(.dina(w_n741_1[0]),.dinb(w_n74_0[2]),.dout(n1022),.clk(gclk));
	jnot g0951(.din(n1022),.dout(n1023),.clk(gclk));
	jand g0952(.dina(n1023),.dinb(n1021),.dout(n1024),.clk(gclk));
	jand g0953(.dina(n1024),.dinb(w_n614_2[2]),.dout(n1025),.clk(gclk));
	jand g0954(.dina(n1025),.dinb(n990),.dout(n1026),.clk(gclk));
	jnot g0955(.din(n1026),.dout(n1027),.clk(gclk));
	jor g0956(.dina(w_n600_0[2]),.dinb(w_n514_0[1]),.dout(n1028),.clk(gclk));
	jand g0957(.dina(n1028),.dinb(w_n782_0[0]),.dout(n1029),.clk(gclk));
	jnot g0958(.din(w_n387_0[0]),.dout(n1030),.clk(gclk));
	jand g0959(.dina(w_n571_0[2]),.dinb(n1030),.dout(n1031),.clk(gclk));
	jnot g0960(.din(n1031),.dout(n1032),.clk(gclk));
	jand g0961(.dina(n1032),.dinb(w_n748_0[0]),.dout(n1033),.clk(gclk));
	jor g0962(.dina(w_n567_1[2]),.dinb(w_n351_0[0]),.dout(n1034),.clk(gclk));
	jand g0963(.dina(w_n598_0[0]),.dinb(n1034),.dout(n1035),.clk(gclk));
	jand g0964(.dina(w_n703_0[1]),.dinb(n1035),.dout(n1036),.clk(gclk));
	jxor g0965(.dina(w_n1036_0[1]),.dinb(w_n771_1[0]),.dout(n1037),.clk(gclk));
	jxor g0966(.dina(n1037),.dinb(w_n1033_0[1]),.dout(n1038),.clk(gclk));
	jand g0967(.dina(n1038),.dinb(w_n1029_0[2]),.dout(n1039),.clk(gclk));
	jor g0968(.dina(w_n1039_0[1]),.dinb(w_n604_1[0]),.dout(n1040),.clk(gclk));
	jand g0969(.dina(w_n1040_0[1]),.dinb(w_n613_0[2]),.dout(n1041),.clk(gclk));
	jor g0970(.dina(w_n704_0[0]),.dinb(w_n600_0[1]),.dout(n1042),.clk(gclk));
	jor g0971(.dina(n1042),.dinb(w_n771_0[2]),.dout(n1043),.clk(gclk));
	jxor g0972(.dina(w_n775_0[0]),.dinb(w_n767_0[2]),.dout(n1044),.clk(gclk));
	jxor g0973(.dina(w_n1044_0[1]),.dinb(w_n1043_0[1]),.dout(n1045),.clk(gclk));
	jor g0974(.dina(w_n1045_0[1]),.dinb(w_n1041_0[1]),.dout(n1046),.clk(gclk));
	jnot g0975(.din(w_n1039_0[0]),.dout(n1047),.clk(gclk));
	jnot g0976(.din(w_n1043_0[0]),.dout(n1048),.clk(gclk));
	jxor g0977(.dina(w_n1044_0[0]),.dinb(w_n1048_0[1]),.dout(n1049),.clk(gclk));
	jor g0978(.dina(n1049),.dinb(w_n604_0[2]),.dout(n1050),.clk(gclk));
	jor g0979(.dina(n1050),.dinb(n1047),.dout(n1051),.clk(gclk));
	jand g0980(.dina(n1051),.dinb(n1046),.dout(n1052),.clk(gclk));
	jand g0981(.dina(n1052),.dinb(n1027),.dout(n1053),.clk(gclk));
	jnot g0982(.din(w_n1053_0[2]),.dout(w_dff_A_tByJlnk29_1),.clk(gclk));
	jxor g0983(.dina(w_n1036_0[0]),.dinb(w_n772_0[0]),.dout(n1055),.clk(gclk));
	jxor g0984(.dina(n1055),.dinb(w_n1033_0[0]),.dout(n1056),.clk(gclk));
	jor g0985(.dina(w_n1045_0[0]),.dinb(w_n1056_0[1]),.dout(n1057),.clk(gclk));
	jand g0986(.dina(w_n1029_0[1]),.dinb(w_n613_0[1]),.dout(n1058),.clk(gclk));
	jand g0987(.dina(n1058),.dinb(n1057),.dout(n1059),.clk(gclk));
	jand g0988(.dina(w_n1048_0[0]),.dinb(w_n767_0[1]),.dout(n1060),.clk(gclk));
	jand g0989(.dina(w_n566_0[1]),.dinb(w_n457_0[0]),.dout(n1061),.clk(gclk));
	jxor g0990(.dina(n1061),.dinb(w_n473_0[0]),.dout(n1062),.clk(gclk));
	jxor g0991(.dina(w_n1062_0[1]),.dinb(w_n777_0[0]),.dout(n1063),.clk(gclk));
	jxor g0992(.dina(n1063),.dinb(n1060),.dout(n1064),.clk(gclk));
	jor g0993(.dina(n1064),.dinb(n1059),.dout(n1065),.clk(gclk));
	jor g0994(.dina(n1065),.dinb(w_n614_2[1]),.dout(n1066),.clk(gclk));
	jand g0995(.dina(w_n1062_0[0]),.dinb(w_n618_1[0]),.dout(n1067),.clk(gclk));
	jnot g0996(.din(n1067),.dout(n1068),.clk(gclk));
	jand g0997(.dina(w_G50_2[0]),.dinb(w_G41_0[0]),.dout(n1069),.clk(gclk));
	jor g0998(.dina(n1069),.dinb(w_n680_1[2]),.dout(n1070),.clk(gclk));
	jand g0999(.dina(w_n638_3[1]),.dinb(w_G137_0[2]),.dout(n1071),.clk(gclk));
	jand g1000(.dina(w_n633_2[2]),.dinb(w_G143_1[0]),.dout(n1072),.clk(gclk));
	jand g1001(.dina(w_n651_3[1]),.dinb(w_G125_0[0]),.dout(n1073),.clk(gclk));
	jor g1002(.dina(n1073),.dinb(n1072),.dout(n1074),.clk(gclk));
	jor g1003(.dina(n1074),.dinb(n1071),.dout(n1075),.clk(gclk));
	jand g1004(.dina(w_n640_3[1]),.dinb(G124),.dout(n1076),.clk(gclk));
	jand g1005(.dina(w_n629_2[0]),.dinb(w_G150_1[1]),.dout(n1077),.clk(gclk));
	jand g1006(.dina(w_n646_3[1]),.dinb(w_G128_0[1]),.dout(n1078),.clk(gclk));
	jor g1007(.dina(n1078),.dinb(n1077),.dout(n1079),.clk(gclk));
	jor g1008(.dina(n1079),.dinb(n1076),.dout(n1080),.clk(gclk));
	jand g1009(.dina(w_n648_1[2]),.dinb(w_G159_1[1]),.dout(n1081),.clk(gclk));
	jand g1010(.dina(w_n653_3[1]),.dinb(w_G132_0[2]),.dout(n1082),.clk(gclk));
	jor g1011(.dina(n1082),.dinb(n1081),.dout(n1083),.clk(gclk));
	jor g1012(.dina(n1083),.dinb(w_G33_4[2]),.dout(n1084),.clk(gclk));
	jor g1013(.dina(n1084),.dinb(n1080),.dout(n1085),.clk(gclk));
	jor g1014(.dina(n1085),.dinb(n1075),.dout(n1086),.clk(gclk));
	jand g1015(.dina(w_n653_3[0]),.dinb(w_G97_1[2]),.dout(n1087),.clk(gclk));
	jand g1016(.dina(w_n646_3[0]),.dinb(w_G107_1[2]),.dout(n1088),.clk(gclk));
	jor g1017(.dina(n1088),.dinb(n1087),.dout(n1089),.clk(gclk));
	jnot g1018(.din(n1089),.dout(n1090),.clk(gclk));
	jand g1019(.dina(w_n648_1[1]),.dinb(w_G58_1[2]),.dout(n1091),.clk(gclk));
	jnot g1020(.din(w_n1091_0[1]),.dout(n1092),.clk(gclk));
	jand g1021(.dina(n1092),.dinb(w_n887_0[0]),.dout(n1093),.clk(gclk));
	jand g1022(.dina(n1093),.dinb(n1090),.dout(n1094),.clk(gclk));
	jand g1023(.dina(w_n640_3[0]),.dinb(w_G283_1[1]),.dout(n1095),.clk(gclk));
	jor g1024(.dina(n1095),.dinb(w_n830_0[0]),.dout(n1096),.clk(gclk));
	jand g1025(.dina(w_n651_3[0]),.dinb(w_G116_2[0]),.dout(n1097),.clk(gclk));
	jand g1026(.dina(w_n638_3[0]),.dinb(w_G87_1[0]),.dout(n1098),.clk(gclk));
	jor g1027(.dina(n1098),.dinb(n1097),.dout(n1099),.clk(gclk));
	jor g1028(.dina(n1099),.dinb(n1096),.dout(n1100),.clk(gclk));
	jnot g1029(.din(n1100),.dout(n1101),.clk(gclk));
	jand g1030(.dina(n1101),.dinb(n1094),.dout(n1102),.clk(gclk));
	jand g1031(.dina(n1102),.dinb(w_G33_4[1]),.dout(n1103),.clk(gclk));
	jnot g1032(.din(n1103),.dout(n1104),.clk(gclk));
	jand g1033(.dina(n1104),.dinb(n1086),.dout(n1105),.clk(gclk));
	jand g1034(.dina(n1105),.dinb(w_n163_0[1]),.dout(n1106),.clk(gclk));
	jor g1035(.dina(n1106),.dinb(n1070),.dout(n1107),.clk(gclk));
	jand g1036(.dina(w_n741_0[2]),.dinb(w_n73_0[2]),.dout(n1108),.clk(gclk));
	jnot g1037(.din(n1108),.dout(n1109),.clk(gclk));
	jand g1038(.dina(n1109),.dinb(n1107),.dout(n1110),.clk(gclk));
	jand g1039(.dina(n1110),.dinb(n1068),.dout(n1111),.clk(gclk));
	jand g1040(.dina(n1111),.dinb(w_n614_2[0]),.dout(n1112),.clk(gclk));
	jnot g1041(.din(n1112),.dout(n1113),.clk(gclk));
	jand g1042(.dina(n1113),.dinb(n1066),.dout(n1114),.clk(gclk));
	jnot g1043(.din(w_n1114_0[2]),.dout(w_dff_A_F97UfJu59_1),.clk(gclk));
	jand g1044(.dina(w_n771_0[1]),.dinb(w_n618_0[2]),.dout(n1116),.clk(gclk));
	jnot g1045(.din(n1116),.dout(n1117),.clk(gclk));
	jand g1046(.dina(w_n646_2[2]),.dinb(w_G283_1[0]),.dout(n1118),.clk(gclk));
	jand g1047(.dina(w_n633_2[1]),.dinb(w_G97_1[1]),.dout(n1119),.clk(gclk));
	jand g1048(.dina(w_n653_2[2]),.dinb(w_G116_1[2]),.dout(n1120),.clk(gclk));
	jor g1049(.dina(n1120),.dinb(n1119),.dout(n1121),.clk(gclk));
	jand g1050(.dina(w_n640_2[2]),.dinb(w_G303_0[2]),.dout(n1122),.clk(gclk));
	jor g1051(.dina(n1122),.dinb(n1121),.dout(n1123),.clk(gclk));
	jor g1052(.dina(n1123),.dinb(n1118),.dout(n1124),.clk(gclk));
	jor g1053(.dina(w_n884_0[0]),.dinb(w_n833_0[0]),.dout(n1125),.clk(gclk));
	jand g1054(.dina(w_n651_2[2]),.dinb(w_G294_1[0]),.dout(n1126),.clk(gclk));
	jand g1055(.dina(w_n638_2[2]),.dinb(w_G107_1[1]),.dout(n1127),.clk(gclk));
	jor g1056(.dina(n1127),.dinb(n1126),.dout(n1128),.clk(gclk));
	jor g1057(.dina(n1128),.dinb(w_n153_2[2]),.dout(n1129),.clk(gclk));
	jor g1058(.dina(n1129),.dinb(n1125),.dout(n1130),.clk(gclk));
	jor g1059(.dina(n1130),.dinb(n1124),.dout(n1131),.clk(gclk));
	jand g1060(.dina(w_n646_2[1]),.dinb(w_G137_0[1]),.dout(n1132),.clk(gclk));
	jand g1061(.dina(w_n633_2[0]),.dinb(w_G159_1[0]),.dout(n1133),.clk(gclk));
	jand g1062(.dina(w_n638_2[1]),.dinb(w_G150_1[0]),.dout(n1134),.clk(gclk));
	jor g1063(.dina(n1134),.dinb(n1133),.dout(n1135),.clk(gclk));
	jand g1064(.dina(w_n651_2[1]),.dinb(w_G132_0[1]),.dout(n1136),.clk(gclk));
	jand g1065(.dina(w_n629_1[2]),.dinb(w_G50_1[2]),.dout(n1137),.clk(gclk));
	jor g1066(.dina(n1137),.dinb(w_n1091_0[0]),.dout(n1138),.clk(gclk));
	jor g1067(.dina(n1138),.dinb(n1136),.dout(n1139),.clk(gclk));
	jand g1068(.dina(w_n653_2[1]),.dinb(w_G143_0[2]),.dout(n1140),.clk(gclk));
	jand g1069(.dina(w_n640_2[1]),.dinb(w_G128_0[0]),.dout(n1141),.clk(gclk));
	jor g1070(.dina(n1141),.dinb(n1140),.dout(n1142),.clk(gclk));
	jor g1071(.dina(n1142),.dinb(w_G33_4[0]),.dout(n1143),.clk(gclk));
	jor g1072(.dina(n1143),.dinb(n1139),.dout(n1144),.clk(gclk));
	jor g1073(.dina(n1144),.dinb(n1135),.dout(n1145),.clk(gclk));
	jor g1074(.dina(n1145),.dinb(n1132),.dout(n1146),.clk(gclk));
	jand g1075(.dina(n1146),.dinb(n1131),.dout(n1147),.clk(gclk));
	jor g1076(.dina(n1147),.dinb(w_n680_1[1]),.dout(n1148),.clk(gclk));
	jand g1077(.dina(w_n741_0[1]),.dinb(w_n75_0[2]),.dout(n1149),.clk(gclk));
	jnot g1078(.din(n1149),.dout(n1150),.clk(gclk));
	jand g1079(.dina(n1150),.dinb(n1148),.dout(n1151),.clk(gclk));
	jand g1080(.dina(n1151),.dinb(n1117),.dout(n1152),.clk(gclk));
	jand g1081(.dina(n1152),.dinb(w_n614_1[2]),.dout(n1153),.clk(gclk));
	jnot g1082(.din(n1153),.dout(n1154),.clk(gclk));
	jor g1083(.dina(w_n1041_0[0]),.dinb(w_n1056_0[0]),.dout(n1155),.clk(gclk));
	jnot g1084(.din(w_n1029_0[0]),.dout(n1156),.clk(gclk));
	jor g1085(.dina(w_n1040_0[0]),.dinb(n1156),.dout(n1157),.clk(gclk));
	jand g1086(.dina(n1157),.dinb(n1155),.dout(n1158),.clk(gclk));
	jand g1087(.dina(n1158),.dinb(n1154),.dout(n1159),.clk(gclk));
	jnot g1088(.din(w_n1159_0[2]),.dout(w_dff_A_07wqAPrM9_1),.clk(gclk));
	jand g1089(.dina(w_n1114_0[1]),.dinb(w_n1053_0[1]),.dout(n1161),.clk(gclk));
	jand g1090(.dina(w_n1159_0[1]),.dinb(w_n759_0[0]),.dout(n1162),.clk(gclk));
	jand g1091(.dina(w_n987_0[1]),.dinb(w_n869_0[1]),.dout(n1163),.clk(gclk));
	jnot g1092(.din(w_G396_0),.dout(n1164),.clk(gclk));
	jand g1093(.dina(w_n937_0[1]),.dinb(w_n1164_0[1]),.dout(n1165),.clk(gclk));
	jand g1094(.dina(w_dff_B_9zpnASnZ7_0),.dinb(n1163),.dout(n1166),.clk(gclk));
	jand g1095(.dina(w_dff_B_c7VrnfJj6_0),.dinb(n1162),.dout(n1167),.clk(gclk));
	jand g1096(.dina(n1167),.dinb(w_n1161_0[1]),.dout(n1168),.clk(gclk));
	jnot g1097(.din(w_n1168_0[1]),.dout(w_dff_A_eICaxmaI2_1),.clk(gclk));
	jnot g1098(.din(w_G343_0[0]),.dout(n1170),.clk(gclk));
	jand g1099(.dina(w_n1161_0[0]),.dinb(w_n1170_0[1]),.dout(n1171),.clk(gclk));
	jnot g1100(.din(w_G213_0[1]),.dout(n1172),.clk(gclk));
	jor g1101(.dina(w_n1168_0[0]),.dinb(w_dff_B_0ZaFb6Dc1_1),.dout(n1173),.clk(gclk));
	jor g1102(.dina(n1173),.dinb(w_dff_B_l3lZnQLq9_1),.dout(G409),.clk(gclk));
	jxor g1103(.dina(w_n937_0[0]),.dinb(w_n1164_0[0]),.dout(n1175),.clk(gclk));
	jxor g1104(.dina(w_n987_0[0]),.dinb(w_n869_0[0]),.dout(n1176),.clk(gclk));
	jxor g1105(.dina(n1176),.dinb(w_dff_B_nAxUj1iK8_1),.dout(n1177),.clk(gclk));
	jand g1106(.dina(w_n1170_0[0]),.dinb(w_G213_0[0]),.dout(n1178),.clk(gclk));
	jxor g1107(.dina(w_n1159_0[0]),.dinb(w_G384_0),.dout(n1179),.clk(gclk));
	jxor g1108(.dina(w_n1179_0[1]),.dinb(w_dff_B_C4JZ1NsH6_1),.dout(n1180),.clk(gclk));
	jand g1109(.dina(n1180),.dinb(w_n1178_0[1]),.dout(n1181),.clk(gclk));
	jnot g1110(.din(w_n1178_0[0]),.dout(n1182),.clk(gclk));
	jxor g1111(.dina(w_n1114_0[0]),.dinb(w_n1053_0[0]),.dout(n1183),.clk(gclk));
	jxor g1112(.dina(n1183),.dinb(w_n1179_0[0]),.dout(n1184),.clk(gclk));
	jand g1113(.dina(w_n1184_0[1]),.dinb(w_dff_B_wCBFBJ289_1),.dout(n1185),.clk(gclk));
	jor g1114(.dina(n1185),.dinb(n1181),.dout(n1186),.clk(gclk));
	jxor g1115(.dina(n1186),.dinb(w_n1177_0[1]),.dout(G405),.clk(gclk));
	jxor g1116(.dina(w_n1184_0[0]),.dinb(w_n1177_0[0]),.dout(w_dff_A_LcUuZJrn4_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G13_0(.douta(w_G13_0[0]),.doutb(w_G13_0[1]),.doutc(w_G13_0[2]),.din(G13));
	jspl3 jspl3_w_G13_1(.douta(w_G13_1[0]),.doutb(w_G13_1[1]),.doutc(w_G13_1[2]),.din(w_G13_0[0]));
	jspl jspl_w_G13_2(.douta(w_G13_2[0]),.doutb(w_G13_2[1]),.din(w_G13_0[1]));
	jspl3 jspl3_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.doutc(w_G20_0[2]),.din(G20));
	jspl3 jspl3_w_G20_1(.douta(w_G20_1[0]),.doutb(w_G20_1[1]),.doutc(w_G20_1[2]),.din(w_G20_0[0]));
	jspl3 jspl3_w_G20_2(.douta(w_G20_2[0]),.doutb(w_G20_2[1]),.doutc(w_G20_2[2]),.din(w_G20_0[1]));
	jspl3 jspl3_w_G20_3(.douta(w_G20_3[0]),.doutb(w_G20_3[1]),.doutc(w_G20_3[2]),.din(w_G20_0[2]));
	jspl3 jspl3_w_G20_4(.douta(w_G20_4[0]),.doutb(w_G20_4[1]),.doutc(w_G20_4[2]),.din(w_G20_1[0]));
	jspl3 jspl3_w_G20_5(.douta(w_G20_5[0]),.doutb(w_G20_5[1]),.doutc(w_G20_5[2]),.din(w_G20_1[1]));
	jspl3 jspl3_w_G20_6(.douta(w_G20_6[0]),.doutb(w_G20_6[1]),.doutc(w_G20_6[2]),.din(w_G20_1[2]));
	jspl3 jspl3_w_G33_0(.douta(w_G33_0[0]),.doutb(w_G33_0[1]),.doutc(w_G33_0[2]),.din(G33));
	jspl3 jspl3_w_G33_1(.douta(w_G33_1[0]),.doutb(w_G33_1[1]),.doutc(w_G33_1[2]),.din(w_G33_0[0]));
	jspl3 jspl3_w_G33_2(.douta(w_G33_2[0]),.doutb(w_G33_2[1]),.doutc(w_G33_2[2]),.din(w_G33_0[1]));
	jspl3 jspl3_w_G33_3(.douta(w_G33_3[0]),.doutb(w_G33_3[1]),.doutc(w_G33_3[2]),.din(w_G33_0[2]));
	jspl3 jspl3_w_G33_4(.douta(w_G33_4[0]),.doutb(w_G33_4[1]),.doutc(w_G33_4[2]),.din(w_G33_1[0]));
	jspl3 jspl3_w_G33_5(.douta(w_G33_5[0]),.doutb(w_G33_5[1]),.doutc(w_G33_5[2]),.din(w_G33_1[1]));
	jspl3 jspl3_w_G33_6(.douta(w_G33_6[0]),.doutb(w_G33_6[1]),.doutc(w_G33_6[2]),.din(w_G33_1[2]));
	jspl3 jspl3_w_G33_7(.douta(w_G33_7[0]),.doutb(w_G33_7[1]),.doutc(w_G33_7[2]),.din(w_G33_2[0]));
	jspl3 jspl3_w_G33_8(.douta(w_G33_8[0]),.doutb(w_G33_8[1]),.doutc(w_G33_8[2]),.din(w_G33_2[1]));
	jspl3 jspl3_w_G33_9(.douta(w_G33_9[0]),.doutb(w_G33_9[1]),.doutc(w_G33_9[2]),.din(w_G33_2[2]));
	jspl3 jspl3_w_G33_10(.douta(w_G33_10[0]),.doutb(w_G33_10[1]),.doutc(w_G33_10[2]),.din(w_G33_3[0]));
	jspl3 jspl3_w_G33_11(.douta(w_G33_11[0]),.doutb(w_G33_11[1]),.doutc(w_G33_11[2]),.din(w_G33_3[1]));
	jspl3 jspl3_w_G33_12(.douta(w_G33_12[0]),.doutb(w_G33_12[1]),.doutc(w_G33_12[2]),.din(w_G33_3[2]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_G41_0[1]),.doutc(w_G41_0[2]),.din(G41));
	jspl3 jspl3_w_G45_0(.douta(w_G45_0[0]),.doutb(w_G45_0[1]),.doutc(w_G45_0[2]),.din(G45));
	jspl jspl_w_G45_1(.douta(w_G45_1[0]),.doutb(w_G45_1[1]),.din(w_G45_0[0]));
	jspl3 jspl3_w_G50_0(.douta(w_G50_0[0]),.doutb(w_G50_0[1]),.doutc(w_G50_0[2]),.din(G50));
	jspl3 jspl3_w_G50_1(.douta(w_G50_1[0]),.doutb(w_G50_1[1]),.doutc(w_G50_1[2]),.din(w_G50_0[0]));
	jspl3 jspl3_w_G50_2(.douta(w_G50_2[0]),.doutb(w_G50_2[1]),.doutc(w_G50_2[2]),.din(w_G50_0[1]));
	jspl3 jspl3_w_G50_3(.douta(w_G50_3[0]),.doutb(w_G50_3[1]),.doutc(w_G50_3[2]),.din(w_G50_0[2]));
	jspl3 jspl3_w_G50_4(.douta(w_G50_4[0]),.doutb(w_G50_4[1]),.doutc(w_G50_4[2]),.din(w_G50_1[0]));
	jspl3 jspl3_w_G50_5(.douta(w_G50_5[0]),.doutb(w_G50_5[1]),.doutc(w_G50_5[2]),.din(w_G50_1[1]));
	jspl3 jspl3_w_G58_0(.douta(w_G58_0[0]),.doutb(w_G58_0[1]),.doutc(w_G58_0[2]),.din(G58));
	jspl3 jspl3_w_G58_1(.douta(w_G58_1[0]),.doutb(w_G58_1[1]),.doutc(w_G58_1[2]),.din(w_G58_0[0]));
	jspl3 jspl3_w_G58_2(.douta(w_G58_2[0]),.doutb(w_G58_2[1]),.doutc(w_G58_2[2]),.din(w_G58_0[1]));
	jspl3 jspl3_w_G58_3(.douta(w_G58_3[0]),.doutb(w_G58_3[1]),.doutc(w_G58_3[2]),.din(w_G58_0[2]));
	jspl3 jspl3_w_G58_4(.douta(w_G58_4[0]),.doutb(w_G58_4[1]),.doutc(w_G58_4[2]),.din(w_G58_1[0]));
	jspl3 jspl3_w_G58_5(.douta(w_G58_5[0]),.doutb(w_G58_5[1]),.doutc(w_G58_5[2]),.din(w_G58_1[1]));
	jspl3 jspl3_w_G68_0(.douta(w_G68_0[0]),.doutb(w_G68_0[1]),.doutc(w_G68_0[2]),.din(G68));
	jspl3 jspl3_w_G68_1(.douta(w_G68_1[0]),.doutb(w_G68_1[1]),.doutc(w_G68_1[2]),.din(w_G68_0[0]));
	jspl3 jspl3_w_G68_2(.douta(w_G68_2[0]),.doutb(w_G68_2[1]),.doutc(w_G68_2[2]),.din(w_G68_0[1]));
	jspl3 jspl3_w_G68_3(.douta(w_G68_3[0]),.doutb(w_G68_3[1]),.doutc(w_G68_3[2]),.din(w_G68_0[2]));
	jspl3 jspl3_w_G68_4(.douta(w_G68_4[0]),.doutb(w_G68_4[1]),.doutc(w_G68_4[2]),.din(w_G68_1[0]));
	jspl3 jspl3_w_G68_5(.douta(w_G68_5[0]),.doutb(w_G68_5[1]),.doutc(w_G68_5[2]),.din(w_G68_1[1]));
	jspl3 jspl3_w_G77_0(.douta(w_G77_0[0]),.doutb(w_G77_0[1]),.doutc(w_G77_0[2]),.din(G77));
	jspl3 jspl3_w_G77_1(.douta(w_G77_1[0]),.doutb(w_G77_1[1]),.doutc(w_G77_1[2]),.din(w_G77_0[0]));
	jspl3 jspl3_w_G77_2(.douta(w_G77_2[0]),.doutb(w_G77_2[1]),.doutc(w_G77_2[2]),.din(w_G77_0[1]));
	jspl3 jspl3_w_G77_3(.douta(w_G77_3[0]),.doutb(w_G77_3[1]),.doutc(w_G77_3[2]),.din(w_G77_0[2]));
	jspl3 jspl3_w_G77_4(.douta(w_G77_4[0]),.doutb(w_G77_4[1]),.doutc(w_G77_4[2]),.din(w_G77_1[0]));
	jspl3 jspl3_w_G87_0(.douta(w_G87_0[0]),.doutb(w_G87_0[1]),.doutc(w_G87_0[2]),.din(G87));
	jspl3 jspl3_w_G87_1(.douta(w_G87_1[0]),.doutb(w_G87_1[1]),.doutc(w_G87_1[2]),.din(w_G87_0[0]));
	jspl3 jspl3_w_G87_2(.douta(w_G87_2[0]),.doutb(w_G87_2[1]),.doutc(w_G87_2[2]),.din(w_G87_0[1]));
	jspl3 jspl3_w_G87_3(.douta(w_G87_3[0]),.doutb(w_G87_3[1]),.doutc(w_G87_3[2]),.din(w_G87_0[2]));
	jspl3 jspl3_w_G97_0(.douta(w_G97_0[0]),.doutb(w_G97_0[1]),.doutc(w_G97_0[2]),.din(G97));
	jspl3 jspl3_w_G97_1(.douta(w_G97_1[0]),.doutb(w_G97_1[1]),.doutc(w_G97_1[2]),.din(w_G97_0[0]));
	jspl3 jspl3_w_G97_2(.douta(w_G97_2[0]),.doutb(w_G97_2[1]),.doutc(w_G97_2[2]),.din(w_G97_0[1]));
	jspl3 jspl3_w_G97_3(.douta(w_G97_3[0]),.doutb(w_G97_3[1]),.doutc(w_G97_3[2]),.din(w_G97_0[2]));
	jspl3 jspl3_w_G97_4(.douta(w_G97_4[0]),.doutb(w_G97_4[1]),.doutc(w_G97_4[2]),.din(w_G97_1[0]));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_G107_0[1]),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G107_1(.douta(w_G107_1[0]),.doutb(w_G107_1[1]),.doutc(w_G107_1[2]),.din(w_G107_0[0]));
	jspl3 jspl3_w_G107_2(.douta(w_G107_2[0]),.doutb(w_G107_2[1]),.doutc(w_G107_2[2]),.din(w_G107_0[1]));
	jspl3 jspl3_w_G107_3(.douta(w_G107_3[0]),.doutb(w_G107_3[1]),.doutc(w_G107_3[2]),.din(w_G107_0[2]));
	jspl jspl_w_G107_4(.douta(w_G107_4[0]),.doutb(w_G107_4[1]),.din(w_G107_1[0]));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G116_1(.douta(w_G116_1[0]),.doutb(w_G116_1[1]),.doutc(w_G116_1[2]),.din(w_G116_0[0]));
	jspl3 jspl3_w_G116_2(.douta(w_G116_2[0]),.doutb(w_G116_2[1]),.doutc(w_G116_2[2]),.din(w_G116_0[1]));
	jspl3 jspl3_w_G116_3(.douta(w_G116_3[0]),.doutb(w_G116_3[1]),.doutc(w_G116_3[2]),.din(w_G116_0[2]));
	jspl3 jspl3_w_G116_4(.douta(w_G116_4[0]),.doutb(w_G116_4[1]),.doutc(w_G116_4[2]),.din(w_G116_1[0]));
	jspl3 jspl3_w_G116_5(.douta(w_G116_5[0]),.doutb(w_G116_5[1]),.doutc(w_G116_5[2]),.din(w_G116_1[1]));
	jspl jspl_w_G125_0(.douta(w_G125_0[0]),.doutb(w_G125_0[1]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(G128));
	jspl3 jspl3_w_G132_0(.douta(w_G132_0[0]),.doutb(w_G132_0[1]),.doutc(w_G132_0[2]),.din(G132));
	jspl jspl_w_G132_1(.douta(w_G132_1[0]),.doutb(w_G132_1[1]),.din(w_G132_0[0]));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_G137_1[0]),.doutb(w_G137_1[1]),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(G143));
	jspl3 jspl3_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.doutc(w_G143_1[2]),.din(w_G143_0[0]));
	jspl jspl_w_G143_2(.douta(w_G143_2[0]),.doutb(w_G143_2[1]),.din(w_G143_0[1]));
	jspl3 jspl3_w_G150_0(.douta(w_G150_0[0]),.doutb(w_G150_0[1]),.doutc(w_G150_0[2]),.din(G150));
	jspl3 jspl3_w_G150_1(.douta(w_G150_1[0]),.doutb(w_G150_1[1]),.doutc(w_G150_1[2]),.din(w_G150_0[0]));
	jspl3 jspl3_w_G150_2(.douta(w_G150_2[0]),.doutb(w_G150_2[1]),.doutc(w_G150_2[2]),.din(w_G150_0[1]));
	jspl jspl_w_G150_3(.douta(w_G150_3[0]),.doutb(w_G150_3[1]),.din(w_G150_0[2]));
	jspl3 jspl3_w_G159_0(.douta(w_G159_0[0]),.doutb(w_G159_0[1]),.doutc(w_G159_0[2]),.din(G159));
	jspl3 jspl3_w_G159_1(.douta(w_G159_1[0]),.doutb(w_G159_1[1]),.doutc(w_G159_1[2]),.din(w_G159_0[0]));
	jspl3 jspl3_w_G159_2(.douta(w_G159_2[0]),.doutb(w_G159_2[1]),.doutc(w_G159_2[2]),.din(w_G159_0[1]));
	jspl3 jspl3_w_G159_3(.douta(w_G159_3[0]),.doutb(w_G159_3[1]),.doutc(w_G159_3[2]),.din(w_G159_0[2]));
	jspl3 jspl3_w_G169_0(.douta(w_G169_0[0]),.doutb(w_G169_0[1]),.doutc(w_G169_0[2]),.din(G169));
	jspl3 jspl3_w_G169_1(.douta(w_G169_1[0]),.doutb(w_G169_1[1]),.doutc(w_G169_1[2]),.din(w_G169_0[0]));
	jspl3 jspl3_w_G169_2(.douta(w_G169_2[0]),.doutb(w_G169_2[1]),.doutc(w_G169_2[2]),.din(w_G169_0[1]));
	jspl jspl_w_G169_3(.douta(w_G169_3[0]),.doutb(w_G169_3[1]),.din(w_G169_0[2]));
	jspl3 jspl3_w_G179_0(.douta(w_G179_0[0]),.doutb(w_G179_0[1]),.doutc(w_G179_0[2]),.din(G179));
	jspl3 jspl3_w_G179_1(.douta(w_G179_1[0]),.doutb(w_G179_1[1]),.doutc(w_G179_1[2]),.din(w_G179_0[0]));
	jspl3 jspl3_w_G179_2(.douta(w_G179_2[0]),.doutb(w_G179_2[1]),.doutc(w_G179_2[2]),.din(w_G179_0[1]));
	jspl3 jspl3_w_G190_0(.douta(w_G190_0[0]),.doutb(w_G190_0[1]),.doutc(w_G190_0[2]),.din(G190));
	jspl3 jspl3_w_G190_1(.douta(w_G190_1[0]),.doutb(w_G190_1[1]),.doutc(w_G190_1[2]),.din(w_G190_0[0]));
	jspl3 jspl3_w_G190_2(.douta(w_G190_2[0]),.doutb(w_G190_2[1]),.doutc(w_G190_2[2]),.din(w_G190_0[1]));
	jspl3 jspl3_w_G190_3(.douta(w_G190_3[0]),.doutb(w_G190_3[1]),.doutc(w_G190_3[2]),.din(w_G190_0[2]));
	jspl3 jspl3_w_G190_4(.douta(w_G190_4[0]),.doutb(w_G190_4[1]),.doutc(w_G190_4[2]),.din(w_G190_1[0]));
	jspl3 jspl3_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.doutc(w_G200_0[2]),.din(G200));
	jspl3 jspl3_w_G200_1(.douta(w_G200_1[0]),.doutb(w_G200_1[1]),.doutc(w_G200_1[2]),.din(w_G200_0[0]));
	jspl3 jspl3_w_G200_2(.douta(w_G200_2[0]),.doutb(w_G200_2[1]),.doutc(w_G200_2[2]),.din(w_G200_0[1]));
	jspl jspl_w_G200_3(.douta(w_G200_3[0]),.doutb(w_G200_3[1]),.din(w_G200_0[2]));
	jspl3 jspl3_w_G213_0(.douta(w_G213_0[0]),.doutb(w_G213_0[1]),.doutc(w_G213_0[2]),.din(G213));
	jspl jspl_w_G223_0(.douta(w_G223_0[0]),.doutb(w_G223_0[1]),.din(G223));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_G226_0[2]),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_G226_1[0]),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G232_0(.douta(w_G232_0[0]),.doutb(w_G232_0[1]),.doutc(w_G232_0[2]),.din(G232));
	jspl3 jspl3_w_G232_1(.douta(w_G232_1[0]),.doutb(w_G232_1[1]),.doutc(w_G232_1[2]),.din(w_G232_0[0]));
	jspl3 jspl3_w_G238_0(.douta(w_G238_0[0]),.doutb(w_G238_0[1]),.doutc(w_G238_0[2]),.din(G238));
	jspl3 jspl3_w_G244_0(.douta(w_G244_0[0]),.doutb(w_G244_0[1]),.doutc(w_G244_0[2]),.din(G244));
	jspl jspl_w_G244_1(.douta(w_G244_1[0]),.doutb(w_G244_1[1]),.din(w_G244_0[0]));
	jspl3 jspl3_w_G250_0(.douta(w_G250_0[0]),.doutb(w_G250_0[1]),.doutc(w_G250_0[2]),.din(G250));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_G257_0[2]),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_G257_1[0]),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G264_0(.douta(w_G264_0[0]),.doutb(w_G264_0[1]),.doutc(w_G264_0[2]),.din(G264));
	jspl3 jspl3_w_G270_0(.douta(w_G270_0[0]),.doutb(w_G270_0[1]),.doutc(w_G270_0[2]),.din(G270));
	jspl3 jspl3_w_G274_0(.douta(w_G274_0[0]),.doutb(w_G274_0[1]),.doutc(w_G274_0[2]),.din(G274));
	jspl3 jspl3_w_G283_0(.douta(w_G283_0[0]),.doutb(w_G283_0[1]),.doutc(w_G283_0[2]),.din(G283));
	jspl3 jspl3_w_G283_1(.douta(w_G283_1[0]),.doutb(w_G283_1[1]),.doutc(w_G283_1[2]),.din(w_G283_0[0]));
	jspl3 jspl3_w_G283_2(.douta(w_G283_2[0]),.doutb(w_G283_2[1]),.doutc(w_G283_2[2]),.din(w_G283_0[1]));
	jspl3 jspl3_w_G283_3(.douta(w_G283_3[0]),.doutb(w_G283_3[1]),.doutc(w_G283_3[2]),.din(w_G283_0[2]));
	jspl3 jspl3_w_G294_0(.douta(w_G294_0[0]),.doutb(w_G294_0[1]),.doutc(w_G294_0[2]),.din(G294));
	jspl3 jspl3_w_G294_1(.douta(w_G294_1[0]),.doutb(w_G294_1[1]),.doutc(w_G294_1[2]),.din(w_G294_0[0]));
	jspl3 jspl3_w_G294_2(.douta(w_G294_2[0]),.doutb(w_G294_2[1]),.doutc(w_G294_2[2]),.din(w_G294_0[1]));
	jspl jspl_w_G294_3(.douta(w_G294_3[0]),.doutb(w_G294_3[1]),.din(w_G294_0[2]));
	jspl3 jspl3_w_G303_0(.douta(w_G303_0[0]),.doutb(w_G303_0[1]),.doutc(w_G303_0[2]),.din(G303));
	jspl3 jspl3_w_G303_1(.douta(w_G303_1[0]),.doutb(w_G303_1[1]),.doutc(w_G303_1[2]),.din(w_G303_0[0]));
	jspl3 jspl3_w_G303_2(.douta(w_G303_2[0]),.doutb(w_G303_2[1]),.doutc(w_G303_2[2]),.din(w_G303_0[1]));
	jspl3 jspl3_w_G311_0(.douta(w_G311_0[0]),.doutb(w_G311_0[1]),.doutc(w_G311_0[2]),.din(G311));
	jspl3 jspl3_w_G311_1(.douta(w_G311_1[0]),.doutb(w_G311_1[1]),.doutc(w_G311_1[2]),.din(w_G311_0[0]));
	jspl3 jspl3_w_G317_0(.douta(w_G317_0[0]),.doutb(w_G317_0[1]),.doutc(w_G317_0[2]),.din(G317));
	jspl jspl_w_G317_1(.douta(w_G317_1[0]),.doutb(w_G317_1[1]),.din(w_G317_0[0]));
	jspl3 jspl3_w_G322_0(.douta(w_G322_0[0]),.doutb(w_G322_0[1]),.doutc(w_G322_0[2]),.din(G322));
	jspl jspl_w_G326_0(.douta(w_G326_0[0]),.doutb(w_G326_0[1]),.din(G326));
	jspl3 jspl3_w_G330_0(.douta(w_G330_0[0]),.doutb(w_G330_0[1]),.doutc(w_G330_0[2]),.din(G330));
	jspl jspl_w_G343_0(.douta(w_G343_0[0]),.doutb(w_G343_0[1]),.din(G343));
	jspl3 jspl3_w_G1698_0(.douta(w_G1698_0[0]),.doutb(w_G1698_0[1]),.doutc(w_G1698_0[2]),.din(G1698));
	jspl jspl_w_G355_0(.douta(w_dff_A_z3QgeTlH5_0),.doutb(w_dff_A_iY0rTqRq8_1),.din(G355_fa_));
	jspl jspl_w_G396_0(.douta(w_G396_0),.doutb(w_dff_A_OMDYSKow2_1),.din(G396_fa_));
	jspl jspl_w_G384_0(.douta(w_dff_A_BhJhL6gc7_0),.doutb(w_dff_A_BIzCn8732_1),.din(G384_fa_));
	jspl3 jspl3_w_n72_0(.douta(w_n72_0[0]),.doutb(w_n72_0[1]),.doutc(w_n72_0[2]),.din(n72));
	jspl3 jspl3_w_n72_1(.douta(w_n72_1[0]),.doutb(w_n72_1[1]),.doutc(w_n72_1[2]),.din(w_n72_0[0]));
	jspl3 jspl3_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.doutc(w_n73_0[2]),.din(n73));
	jspl3 jspl3_w_n73_1(.douta(w_n73_1[0]),.doutb(w_n73_1[1]),.doutc(w_n73_1[2]),.din(w_n73_0[0]));
	jspl3 jspl3_w_n73_2(.douta(w_n73_2[0]),.doutb(w_n73_2[1]),.doutc(w_n73_2[2]),.din(w_n73_0[1]));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl3 jspl3_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.doutc(w_n74_1[2]),.din(w_n74_0[0]));
	jspl jspl_w_n74_2(.douta(w_n74_2[0]),.doutb(w_n74_2[1]),.din(w_n74_0[1]));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.doutc(w_n75_0[2]),.din(n75));
	jspl3 jspl3_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.doutc(w_n75_1[2]),.din(w_n75_0[0]));
	jspl jspl_w_n75_2(.douta(w_n75_2[0]),.doutb(w_n75_2[1]),.din(w_n75_0[1]));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.din(n76));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl3 jspl3_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.doutc(w_n79_0[2]),.din(n79));
	jspl3 jspl3_w_n79_1(.douta(w_n79_1[0]),.doutb(w_n79_1[1]),.doutc(w_n79_1[2]),.din(w_n79_0[0]));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.doutc(w_n80_0[2]),.din(n80));
	jspl3 jspl3_w_n80_1(.douta(w_n80_1[0]),.doutb(w_n80_1[1]),.doutc(w_n80_1[2]),.din(w_n80_0[0]));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl3 jspl3_w_n81_1(.douta(w_n81_1[0]),.doutb(w_n81_1[1]),.doutc(w_n81_1[2]),.din(w_n81_0[0]));
	jspl jspl_w_n81_2(.douta(w_n81_2[0]),.doutb(w_n81_2[1]),.din(w_n81_0[1]));
	jspl3 jspl3_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.doutc(w_n84_0[2]),.din(n84));
	jspl3 jspl3_w_n84_1(.douta(w_n84_1[0]),.doutb(w_n84_1[1]),.doutc(w_n84_1[2]),.din(w_n84_0[0]));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl3 jspl3_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.doutc(w_n86_0[2]),.din(n86));
	jspl jspl_w_n89_0(.douta(w_n89_0[0]),.doutb(w_n89_0[1]),.din(n89));
	jspl3 jspl3_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.doutc(w_n91_0[2]),.din(n91));
	jspl3 jspl3_w_n91_1(.douta(w_n91_1[0]),.doutb(w_n91_1[1]),.doutc(w_n91_1[2]),.din(w_n91_0[0]));
	jspl3 jspl3_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.doutc(w_n96_0[2]),.din(n96));
	jspl3 jspl3_w_n105_0(.douta(w_n105_0[0]),.doutb(w_n105_0[1]),.doutc(w_n105_0[2]),.din(n105));
	jspl jspl_w_n105_1(.douta(w_n105_1[0]),.doutb(w_n105_1[1]),.din(w_n105_0[0]));
	jspl3 jspl3_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.doutc(w_n111_0[2]),.din(n111));
	jspl jspl_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.din(n126));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.din(n130));
	jspl jspl_w_n134_0(.douta(w_n134_0[0]),.doutb(w_n134_0[1]),.din(n134));
	jspl jspl_w_n137_0(.douta(w_n137_0[0]),.doutb(w_n137_0[1]),.din(n137));
	jspl3 jspl3_w_n139_0(.douta(w_n139_0[0]),.doutb(w_n139_0[1]),.doutc(w_n139_0[2]),.din(n139));
	jspl3 jspl3_w_n139_1(.douta(w_n139_1[0]),.doutb(w_n139_1[1]),.doutc(w_n139_1[2]),.din(w_n139_0[0]));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl3 jspl3_w_n141_1(.douta(w_n141_1[0]),.doutb(w_n141_1[1]),.doutc(w_n141_1[2]),.din(w_n141_0[0]));
	jspl3 jspl3_w_n141_2(.douta(w_n141_2[0]),.doutb(w_n141_2[1]),.doutc(w_n141_2[2]),.din(w_n141_0[1]));
	jspl jspl_w_n141_3(.douta(w_n141_3[0]),.doutb(w_n141_3[1]),.din(w_n141_0[2]));
	jspl3 jspl3_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.doutc(w_n142_0[2]),.din(n142));
	jspl3 jspl3_w_n142_1(.douta(w_n142_1[0]),.doutb(w_n142_1[1]),.doutc(w_n142_1[2]),.din(w_n142_0[0]));
	jspl jspl_w_n142_2(.douta(w_n142_2[0]),.doutb(w_n142_2[1]),.din(w_n142_0[1]));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n144_1(.douta(w_n144_1[0]),.doutb(w_n144_1[1]),.doutc(w_n144_1[2]),.din(w_n144_0[0]));
	jspl jspl_w_n144_2(.douta(w_n144_2[0]),.doutb(w_n144_2[1]),.din(w_n144_0[1]));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl jspl_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.din(n148));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_n151_1[1]),.doutc(w_n151_1[2]),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_n151_2[0]),.doutb(w_n151_2[1]),.doutc(w_n151_2[2]),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_n151_3[0]),.doutb(w_n151_3[1]),.doutc(w_n151_3[2]),.din(w_n151_0[2]));
	jspl3 jspl3_w_n151_4(.douta(w_n151_4[0]),.doutb(w_n151_4[1]),.doutc(w_n151_4[2]),.din(w_n151_1[0]));
	jspl3 jspl3_w_n151_5(.douta(w_n151_5[0]),.doutb(w_n151_5[1]),.doutc(w_n151_5[2]),.din(w_n151_1[1]));
	jspl jspl_w_n151_6(.douta(w_n151_6[0]),.doutb(w_n151_6[1]),.din(w_n151_1[2]));
	jspl3 jspl3_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.doutc(w_n152_0[2]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.doutc(w_n153_1[2]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n153_2(.douta(w_n153_2[0]),.doutb(w_n153_2[1]),.doutc(w_n153_2[2]),.din(w_n153_0[1]));
	jspl3 jspl3_w_n153_3(.douta(w_n153_3[0]),.doutb(w_n153_3[1]),.doutc(w_n153_3[2]),.din(w_n153_0[2]));
	jspl3 jspl3_w_n153_4(.douta(w_n153_4[0]),.doutb(w_n153_4[1]),.doutc(w_n153_4[2]),.din(w_n153_1[0]));
	jspl3 jspl3_w_n153_5(.douta(w_n153_5[0]),.doutb(w_n153_5[1]),.doutc(w_n153_5[2]),.din(w_n153_1[1]));
	jspl3 jspl3_w_n153_6(.douta(w_n153_6[0]),.doutb(w_n153_6[1]),.doutc(w_n153_6[2]),.din(w_n153_1[2]));
	jspl3 jspl3_w_n153_7(.douta(w_n153_7[0]),.doutb(w_n153_7[1]),.doutc(w_n153_7[2]),.din(w_n153_2[0]));
	jspl jspl_w_n153_8(.douta(w_n153_8[0]),.doutb(w_n153_8[1]),.din(w_n153_2[1]));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_n163_0[2]),.din(n163));
	jspl jspl_w_n163_1(.douta(w_n163_1[0]),.doutb(w_n163_1[1]),.din(w_n163_0[0]));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_n164_0[2]),.din(n164));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(n165));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl3 jspl3_w_n168_1(.douta(w_n168_1[0]),.doutb(w_n168_1[1]),.doutc(w_n168_1[2]),.din(w_n168_0[0]));
	jspl3 jspl3_w_n168_2(.douta(w_n168_2[0]),.doutb(w_n168_2[1]),.doutc(w_n168_2[2]),.din(w_n168_0[1]));
	jspl3 jspl3_w_n168_3(.douta(w_n168_3[0]),.doutb(w_n168_3[1]),.doutc(w_n168_3[2]),.din(w_n168_0[2]));
	jspl3 jspl3_w_n168_4(.douta(w_n168_4[0]),.doutb(w_n168_4[1]),.doutc(w_n168_4[2]),.din(w_n168_1[0]));
	jspl jspl_w_n168_5(.douta(w_n168_5[0]),.doutb(w_n168_5[1]),.din(w_n168_1[1]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl3 jspl3_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.doutc(w_n172_0[2]),.din(n172));
	jspl3 jspl3_w_n172_1(.douta(w_n172_1[0]),.doutb(w_n172_1[1]),.doutc(w_n172_1[2]),.din(w_n172_0[0]));
	jspl3 jspl3_w_n172_2(.douta(w_n172_2[0]),.doutb(w_n172_2[1]),.doutc(w_n172_2[2]),.din(w_n172_0[1]));
	jspl3 jspl3_w_n172_3(.douta(w_n172_3[0]),.doutb(w_n172_3[1]),.doutc(w_n172_3[2]),.din(w_n172_0[2]));
	jspl3 jspl3_w_n172_4(.douta(w_n172_4[0]),.doutb(w_n172_4[1]),.doutc(w_n172_4[2]),.din(w_n172_1[0]));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl3 jspl3_w_n173_1(.douta(w_n173_1[0]),.doutb(w_n173_1[1]),.doutc(w_n173_1[2]),.din(w_n173_0[0]));
	jspl3 jspl3_w_n173_2(.douta(w_n173_2[0]),.doutb(w_n173_2[1]),.doutc(w_n173_2[2]),.din(w_n173_0[1]));
	jspl jspl_w_n173_3(.douta(w_n173_3[0]),.doutb(w_n173_3[1]),.din(w_n173_0[2]));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.doutc(w_n177_0[2]),.din(n177));
	jspl3 jspl3_w_n177_1(.douta(w_n177_1[0]),.doutb(w_n177_1[1]),.doutc(w_n177_1[2]),.din(w_n177_0[0]));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl jspl_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.doutc(w_n186_0[2]),.din(n186));
	jspl3 jspl3_w_n186_1(.douta(w_n186_1[0]),.doutb(w_n186_1[1]),.doutc(w_n186_1[2]),.din(w_n186_0[0]));
	jspl3 jspl3_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.doutc(w_n189_0[2]),.din(n189));
	jspl3 jspl3_w_n189_1(.douta(w_n189_1[0]),.doutb(w_n189_1[1]),.doutc(w_n189_1[2]),.din(w_n189_0[0]));
	jspl3 jspl3_w_n189_2(.douta(w_n189_2[0]),.doutb(w_n189_2[1]),.doutc(w_n189_2[2]),.din(w_n189_0[1]));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.doutc(w_n192_0[2]),.din(n192));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_n198_0[2]),.din(n198));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.doutc(w_n199_0[2]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(n202));
	jspl3 jspl3_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.doutc(w_n205_0[2]),.din(n205));
	jspl jspl_w_n205_1(.douta(w_n205_1[0]),.doutb(w_n205_1[1]),.din(w_n205_0[0]));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl3 jspl3_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.doutc(w_n212_0[2]),.din(n212));
	jspl jspl_w_n212_1(.douta(w_n212_1[0]),.doutb(w_n212_1[1]),.din(w_n212_0[0]));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl jspl_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.din(n215));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.doutc(w_n224_0[2]),.din(n224));
	jspl jspl_w_n224_1(.douta(w_n224_1[0]),.doutb(w_n224_1[1]),.din(w_n224_0[0]));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(n225));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.din(n229));
	jspl3 jspl3_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.doutc(w_n234_0[2]),.din(n234));
	jspl jspl_w_n234_1(.douta(w_n234_1[0]),.doutb(w_n234_1[1]),.din(w_n234_0[0]));
	jspl3 jspl3_w_n237_0(.douta(w_n237_0[0]),.doutb(w_n237_0[1]),.doutc(w_n237_0[2]),.din(n237));
	jspl jspl_w_n238_0(.douta(w_n238_0[0]),.doutb(w_n238_0[1]),.din(n238));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl jspl_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.din(n243));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.din(n251));
	jspl3 jspl3_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.doutc(w_n255_0[2]),.din(n255));
	jspl jspl_w_n255_1(.douta(w_n255_1[0]),.doutb(w_n255_1[1]),.din(w_n255_0[0]));
	jspl jspl_w_n256_0(.douta(w_n256_0[0]),.doutb(w_n256_0[1]),.din(n256));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl3 jspl3_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.doutc(w_n261_0[2]),.din(n261));
	jspl3 jspl3_w_n261_1(.douta(w_n261_1[0]),.doutb(w_n261_1[1]),.doutc(w_n261_1[2]),.din(w_n261_0[0]));
	jspl3 jspl3_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.doutc(w_n262_0[2]),.din(n262));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.din(n269));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl3 jspl3_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.doutc(w_n279_0[2]),.din(n279));
	jspl jspl_w_n279_1(.douta(w_n279_1[0]),.doutb(w_n279_1[1]),.din(w_n279_0[0]));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.din(n283));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.din(n298));
	jspl3 jspl3_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.doutc(w_n308_0[2]),.din(n308));
	jspl3 jspl3_w_n308_1(.douta(w_n308_1[0]),.doutb(w_n308_1[1]),.doutc(w_n308_1[2]),.din(w_n308_0[0]));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(n309));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(n310));
	jspl jspl_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.din(n312));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.doutc(w_n315_0[2]),.din(n315));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.din(n321));
	jspl3 jspl3_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.doutc(w_n323_0[2]),.din(n323));
	jspl3 jspl3_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.doutc(w_n330_0[2]),.din(n330));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl jspl_w_n344_0(.douta(w_n344_0[0]),.doutb(w_n344_0[1]),.din(n344));
	jspl jspl_w_n347_0(.douta(w_n347_0[0]),.doutb(w_n347_0[1]),.din(n347));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n351_0(.douta(w_n351_0[0]),.doutb(w_n351_0[1]),.din(n351));
	jspl3 jspl3_w_n352_0(.douta(w_n352_0[0]),.doutb(w_n352_0[1]),.doutc(w_n352_0[2]),.din(n352));
	jspl jspl_w_n352_1(.douta(w_n352_1[0]),.doutb(w_n352_1[1]),.din(w_n352_0[0]));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_n354_0[2]),.din(n354));
	jspl jspl_w_n354_1(.douta(w_n354_1[0]),.doutb(w_n354_1[1]),.din(w_n354_0[0]));
	jspl jspl_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.din(n355));
	jspl3 jspl3_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.doutc(w_n356_0[2]),.din(n356));
	jspl jspl_w_n356_1(.douta(w_n356_1[0]),.doutb(w_n356_1[1]),.din(w_n356_0[0]));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl jspl_w_n367_1(.douta(w_n367_1[0]),.doutb(w_n367_1[1]),.din(w_n367_0[0]));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(n370));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl jspl_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.din(n378));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_n388_0[2]),.din(n388));
	jspl3 jspl3_w_n388_1(.douta(w_n388_1[0]),.doutb(w_n388_1[1]),.doutc(w_n388_1[2]),.din(w_n388_0[0]));
	jspl jspl_w_n388_2(.douta(w_n388_2[0]),.doutb(w_n388_2[1]),.din(w_n388_0[1]));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n395_0(.douta(w_n395_0[0]),.doutb(w_n395_0[1]),.din(n395));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl3 jspl3_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.doutc(w_n414_0[2]),.din(n414));
	jspl3 jspl3_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.doutc(w_n417_0[2]),.din(n417));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.din(n420));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl jspl_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.din(n428));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.doutc(w_n439_0[2]),.din(n439));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n450_0(.douta(w_n450_0[0]),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl jspl_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.din(n473));
	jspl3 jspl3_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.doutc(w_n482_0[2]),.din(n482));
	jspl jspl_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(n499));
	jspl jspl_w_n500_0(.douta(w_n500_0[0]),.doutb(w_n500_0[1]),.din(n500));
	jspl3 jspl3_w_n503_0(.douta(w_n503_0[0]),.doutb(w_n503_0[1]),.doutc(w_n503_0[2]),.din(n503));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl jspl_w_n507_2(.douta(w_n507_2[0]),.doutb(w_n507_2[1]),.din(w_n507_0[1]));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl3 jspl3_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.doutc(w_n514_0[2]),.din(n514));
	jspl jspl_w_n514_1(.douta(w_n514_1[0]),.doutb(w_n514_1[1]),.din(w_n514_0[0]));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_n559_0[1]),.din(n559));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl jspl_w_n566_1(.douta(w_n566_1[0]),.doutb(w_n566_1[1]),.din(w_n566_0[0]));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl3 jspl3_w_n567_1(.douta(w_n567_1[0]),.doutb(w_n567_1[1]),.doutc(w_n567_1[2]),.din(w_n567_0[0]));
	jspl3 jspl3_w_n567_2(.douta(w_n567_2[0]),.doutb(w_n567_2[1]),.doutc(w_n567_2[2]),.din(w_n567_0[1]));
	jspl3 jspl3_w_n567_3(.douta(w_n567_3[0]),.doutb(w_n567_3[1]),.doutc(w_n567_3[2]),.din(w_n567_0[2]));
	jspl3 jspl3_w_n567_4(.douta(w_n567_4[0]),.doutb(w_n567_4[1]),.doutc(w_n567_4[2]),.din(w_n567_1[0]));
	jspl jspl_w_n567_5(.douta(w_n567_5[0]),.doutb(w_n567_5[1]),.din(w_n567_1[1]));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.din(n569));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_n571_0[2]),.din(n571));
	jspl3 jspl3_w_n571_1(.douta(w_n571_1[0]),.doutb(w_n571_1[1]),.doutc(w_n571_1[2]),.din(w_n571_0[0]));
	jspl jspl_w_n571_2(.douta(w_n571_2[0]),.doutb(w_n571_2[1]),.din(w_n571_0[1]));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl jspl_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.din(n573));
	jspl jspl_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.din(n574));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(n577));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.doutc(w_n579_0[2]),.din(n579));
	jspl jspl_w_n579_1(.douta(w_n579_1[0]),.doutb(w_n579_1[1]),.din(w_n579_0[0]));
	jspl3 jspl3_w_n580_0(.douta(w_n580_0[0]),.doutb(w_n580_0[1]),.doutc(w_n580_0[2]),.din(n580));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl3 jspl3_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.doutc(w_n600_0[2]),.din(n600));
	jspl3 jspl3_w_n600_1(.douta(w_n600_1[0]),.doutb(w_n600_1[1]),.doutc(w_n600_1[2]),.din(w_n600_0[0]));
	jspl3 jspl3_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.doutc(w_n601_0[2]),.din(n601));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.doutc(w_n604_0[2]),.din(n604));
	jspl3 jspl3_w_n604_1(.douta(w_n604_1[0]),.doutb(w_n604_1[1]),.doutc(w_n604_1[2]),.din(w_n604_0[0]));
	jspl3 jspl3_w_n604_2(.douta(w_n604_2[0]),.doutb(w_n604_2[1]),.doutc(w_n604_2[2]),.din(w_n604_0[1]));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.doutc(w_n613_1[2]),.din(w_n613_0[0]));
	jspl3 jspl3_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.doutc(w_n614_0[2]),.din(n614));
	jspl3 jspl3_w_n614_1(.douta(w_n614_1[0]),.doutb(w_n614_1[1]),.doutc(w_n614_1[2]),.din(w_n614_0[0]));
	jspl3 jspl3_w_n614_2(.douta(w_n614_2[0]),.doutb(w_n614_2[1]),.doutc(w_n614_2[2]),.din(w_n614_0[1]));
	jspl3 jspl3_w_n614_3(.douta(w_n614_3[0]),.doutb(w_n614_3[1]),.doutc(w_n614_3[2]),.din(w_n614_0[2]));
	jspl3 jspl3_w_n614_4(.douta(w_n614_4[0]),.doutb(w_n614_4[1]),.doutc(w_n614_4[2]),.din(w_n614_1[0]));
	jspl jspl_w_n614_5(.douta(w_n614_5[0]),.doutb(w_n614_5[1]),.din(w_n614_1[1]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl3 jspl3_w_n618_1(.douta(w_n618_1[0]),.doutb(w_n618_1[1]),.doutc(w_n618_1[2]),.din(w_n618_0[0]));
	jspl jspl_w_n618_2(.douta(w_n618_2[0]),.doutb(w_n618_2[1]),.din(w_n618_0[1]));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.doutc(w_n620_0[2]),.din(n620));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl3 jspl3_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.doutc(w_n626_0[2]),.din(n626));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(n628));
	jspl3 jspl3_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.doutc(w_n629_0[2]),.din(n629));
	jspl3 jspl3_w_n629_1(.douta(w_n629_1[0]),.doutb(w_n629_1[1]),.doutc(w_n629_1[2]),.din(w_n629_0[0]));
	jspl3 jspl3_w_n629_2(.douta(w_n629_2[0]),.doutb(w_n629_2[1]),.doutc(w_n629_2[2]),.din(w_n629_0[1]));
	jspl3 jspl3_w_n629_3(.douta(w_n629_3[0]),.doutb(w_n629_3[1]),.doutc(w_n629_3[2]),.din(w_n629_0[2]));
	jspl3 jspl3_w_n629_4(.douta(w_n629_4[0]),.doutb(w_n629_4[1]),.doutc(w_n629_4[2]),.din(w_n629_1[0]));
	jspl jspl_w_n629_5(.douta(w_n629_5[0]),.doutb(w_n629_5[1]),.din(w_n629_1[1]));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl3 jspl3_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.doutc(w_n633_0[2]),.din(n633));
	jspl3 jspl3_w_n633_1(.douta(w_n633_1[0]),.doutb(w_n633_1[1]),.doutc(w_n633_1[2]),.din(w_n633_0[0]));
	jspl3 jspl3_w_n633_2(.douta(w_n633_2[0]),.doutb(w_n633_2[1]),.doutc(w_n633_2[2]),.din(w_n633_0[1]));
	jspl3 jspl3_w_n633_3(.douta(w_n633_3[0]),.doutb(w_n633_3[1]),.doutc(w_n633_3[2]),.din(w_n633_0[2]));
	jspl3 jspl3_w_n633_4(.douta(w_n633_4[0]),.doutb(w_n633_4[1]),.doutc(w_n633_4[2]),.din(w_n633_1[0]));
	jspl3 jspl3_w_n633_5(.douta(w_n633_5[0]),.doutb(w_n633_5[1]),.doutc(w_n633_5[2]),.din(w_n633_1[1]));
	jspl jspl_w_n633_6(.douta(w_n633_6[0]),.doutb(w_n633_6[1]),.din(w_n633_1[2]));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(n637));
	jspl3 jspl3_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.doutc(w_n638_0[2]),.din(n638));
	jspl3 jspl3_w_n638_1(.douta(w_n638_1[0]),.doutb(w_n638_1[1]),.doutc(w_n638_1[2]),.din(w_n638_0[0]));
	jspl3 jspl3_w_n638_2(.douta(w_n638_2[0]),.doutb(w_n638_2[1]),.doutc(w_n638_2[2]),.din(w_n638_0[1]));
	jspl3 jspl3_w_n638_3(.douta(w_n638_3[0]),.doutb(w_n638_3[1]),.doutc(w_n638_3[2]),.din(w_n638_0[2]));
	jspl3 jspl3_w_n638_4(.douta(w_n638_4[0]),.doutb(w_n638_4[1]),.doutc(w_n638_4[2]),.din(w_n638_1[0]));
	jspl3 jspl3_w_n638_5(.douta(w_n638_5[0]),.doutb(w_n638_5[1]),.doutc(w_n638_5[2]),.din(w_n638_1[1]));
	jspl3 jspl3_w_n638_6(.douta(w_n638_6[0]),.doutb(w_n638_6[1]),.doutc(w_n638_6[2]),.din(w_n638_1[2]));
	jspl jspl_w_n638_7(.douta(w_n638_7[0]),.doutb(w_n638_7[1]),.din(w_n638_2[0]));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl3 jspl3_w_n640_2(.douta(w_n640_2[0]),.doutb(w_n640_2[1]),.doutc(w_n640_2[2]),.din(w_n640_0[1]));
	jspl3 jspl3_w_n640_3(.douta(w_n640_3[0]),.doutb(w_n640_3[1]),.doutc(w_n640_3[2]),.din(w_n640_0[2]));
	jspl3 jspl3_w_n640_4(.douta(w_n640_4[0]),.doutb(w_n640_4[1]),.doutc(w_n640_4[2]),.din(w_n640_1[0]));
	jspl3 jspl3_w_n640_5(.douta(w_n640_5[0]),.doutb(w_n640_5[1]),.doutc(w_n640_5[2]),.din(w_n640_1[1]));
	jspl3 jspl3_w_n640_6(.douta(w_n640_6[0]),.doutb(w_n640_6[1]),.doutc(w_n640_6[2]),.din(w_n640_1[2]));
	jspl jspl_w_n640_7(.douta(w_n640_7[0]),.doutb(w_n640_7[1]),.din(w_n640_2[0]));
	jspl3 jspl3_w_n646_0(.douta(w_n646_0[0]),.doutb(w_n646_0[1]),.doutc(w_n646_0[2]),.din(n646));
	jspl3 jspl3_w_n646_1(.douta(w_n646_1[0]),.doutb(w_n646_1[1]),.doutc(w_n646_1[2]),.din(w_n646_0[0]));
	jspl3 jspl3_w_n646_2(.douta(w_n646_2[0]),.doutb(w_n646_2[1]),.doutc(w_n646_2[2]),.din(w_n646_0[1]));
	jspl3 jspl3_w_n646_3(.douta(w_n646_3[0]),.doutb(w_n646_3[1]),.doutc(w_n646_3[2]),.din(w_n646_0[2]));
	jspl3 jspl3_w_n646_4(.douta(w_n646_4[0]),.doutb(w_n646_4[1]),.doutc(w_n646_4[2]),.din(w_n646_1[0]));
	jspl3 jspl3_w_n646_5(.douta(w_n646_5[0]),.doutb(w_n646_5[1]),.doutc(w_n646_5[2]),.din(w_n646_1[1]));
	jspl3 jspl3_w_n646_6(.douta(w_n646_6[0]),.doutb(w_n646_6[1]),.doutc(w_n646_6[2]),.din(w_n646_1[2]));
	jspl jspl_w_n646_7(.douta(w_n646_7[0]),.doutb(w_n646_7[1]),.din(w_n646_2[0]));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.doutc(w_n648_0[2]),.din(n648));
	jspl3 jspl3_w_n648_1(.douta(w_n648_1[0]),.doutb(w_n648_1[1]),.doutc(w_n648_1[2]),.din(w_n648_0[0]));
	jspl3 jspl3_w_n648_2(.douta(w_n648_2[0]),.doutb(w_n648_2[1]),.doutc(w_n648_2[2]),.din(w_n648_0[1]));
	jspl3 jspl3_w_n648_3(.douta(w_n648_3[0]),.doutb(w_n648_3[1]),.doutc(w_n648_3[2]),.din(w_n648_0[2]));
	jspl jspl_w_n648_4(.douta(w_n648_4[0]),.doutb(w_n648_4[1]),.din(w_n648_1[0]));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.doutc(w_n651_0[2]),.din(n651));
	jspl3 jspl3_w_n651_1(.douta(w_n651_1[0]),.doutb(w_n651_1[1]),.doutc(w_n651_1[2]),.din(w_n651_0[0]));
	jspl3 jspl3_w_n651_2(.douta(w_n651_2[0]),.doutb(w_n651_2[1]),.doutc(w_n651_2[2]),.din(w_n651_0[1]));
	jspl3 jspl3_w_n651_3(.douta(w_n651_3[0]),.doutb(w_n651_3[1]),.doutc(w_n651_3[2]),.din(w_n651_0[2]));
	jspl3 jspl3_w_n651_4(.douta(w_n651_4[0]),.doutb(w_n651_4[1]),.doutc(w_n651_4[2]),.din(w_n651_1[0]));
	jspl3 jspl3_w_n651_5(.douta(w_n651_5[0]),.doutb(w_n651_5[1]),.doutc(w_n651_5[2]),.din(w_n651_1[1]));
	jspl3 jspl3_w_n651_6(.douta(w_n651_6[0]),.doutb(w_n651_6[1]),.doutc(w_n651_6[2]),.din(w_n651_1[2]));
	jspl jspl_w_n651_7(.douta(w_n651_7[0]),.doutb(w_n651_7[1]),.din(w_n651_2[0]));
	jspl3 jspl3_w_n653_0(.douta(w_n653_0[0]),.doutb(w_n653_0[1]),.doutc(w_n653_0[2]),.din(n653));
	jspl3 jspl3_w_n653_1(.douta(w_n653_1[0]),.doutb(w_n653_1[1]),.doutc(w_n653_1[2]),.din(w_n653_0[0]));
	jspl3 jspl3_w_n653_2(.douta(w_n653_2[0]),.doutb(w_n653_2[1]),.doutc(w_n653_2[2]),.din(w_n653_0[1]));
	jspl3 jspl3_w_n653_3(.douta(w_n653_3[0]),.doutb(w_n653_3[1]),.doutc(w_n653_3[2]),.din(w_n653_0[2]));
	jspl3 jspl3_w_n653_4(.douta(w_n653_4[0]),.doutb(w_n653_4[1]),.doutc(w_n653_4[2]),.din(w_n653_1[0]));
	jspl3 jspl3_w_n653_5(.douta(w_n653_5[0]),.doutb(w_n653_5[1]),.doutc(w_n653_5[2]),.din(w_n653_1[1]));
	jspl3 jspl3_w_n653_6(.douta(w_n653_6[0]),.doutb(w_n653_6[1]),.doutc(w_n653_6[2]),.din(w_n653_1[2]));
	jspl jspl_w_n653_7(.douta(w_n653_7[0]),.doutb(w_n653_7[1]),.din(w_n653_2[0]));
	jspl3 jspl3_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.doutc(w_n680_0[2]),.din(n680));
	jspl3 jspl3_w_n680_1(.douta(w_n680_1[0]),.doutb(w_n680_1[1]),.doutc(w_n680_1[2]),.din(w_n680_0[0]));
	jspl3 jspl3_w_n680_2(.douta(w_n680_2[0]),.doutb(w_n680_2[1]),.doutc(w_n680_2[2]),.din(w_n680_0[1]));
	jspl3 jspl3_w_n680_3(.douta(w_n680_3[0]),.doutb(w_n680_3[1]),.doutc(w_n680_3[2]),.din(w_n680_0[2]));
	jspl jspl_w_n680_4(.douta(w_n680_4[0]),.doutb(w_n680_4[1]),.din(w_n680_1[0]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl3 jspl3_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.doutc(w_n684_0[2]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl3 jspl3_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.doutc(w_n690_0[2]),.din(n690));
	jspl jspl_w_n690_1(.douta(w_n690_1[0]),.doutb(w_n690_1[1]),.din(w_n690_0[0]));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.din(n692));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n703_1(.douta(w_n703_1[0]),.doutb(w_n703_1[1]),.din(w_n703_0[0]));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.din(n718));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n741_1(.douta(w_n741_1[0]),.doutb(w_n741_1[1]),.din(w_n741_0[0]));
	jspl jspl_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.din(n748));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n766_0(.douta(w_n766_0[0]),.doutb(w_n766_0[1]),.din(n766));
	jspl3 jspl3_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.doutc(w_n767_0[2]),.din(n767));
	jspl jspl_w_n767_1(.douta(w_n767_1[0]),.doutb(w_n767_1[1]),.din(w_n767_0[0]));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_n771_0[2]),.din(n771));
	jspl jspl_w_n771_1(.douta(w_n771_1[0]),.doutb(w_n771_1[1]),.din(w_n771_0[0]));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.din(n798));
	jspl3 jspl3_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.doutc(w_n802_0[2]),.din(n802));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(n817));
	jspl jspl_w_n830_0(.douta(w_n830_0[0]),.doutb(w_n830_0[1]),.din(n830));
	jspl jspl_w_n833_0(.douta(w_n833_0[0]),.doutb(w_n833_0[1]),.din(n833));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.doutc(w_n845_0[2]),.din(n845));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(n861));
	jspl3 jspl3_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.doutc(w_n863_0[2]),.din(n863));
	jspl3 jspl3_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.doutc(w_n869_0[2]),.din(n869));
	jspl jspl_w_n873_0(.douta(w_n873_0[0]),.doutb(w_n873_0[1]),.din(n873));
	jspl jspl_w_n875_0(.douta(w_n875_0[0]),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.din(n887));
	jspl3 jspl3_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.doutc(w_n937_0[2]),.din(n937));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(n959));
	jspl3 jspl3_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.doutc(w_n987_0[2]),.din(n987));
	jspl3 jspl3_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.doutc(w_n1029_0[2]),.din(n1029));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1036_0(.douta(w_n1036_0[0]),.doutb(w_n1036_0[1]),.din(n1036));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.din(n1039));
	jspl jspl_w_n1040_0(.douta(w_n1040_0[0]),.doutb(w_n1040_0[1]),.din(n1040));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(n1043));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(n1044));
	jspl jspl_w_n1045_0(.douta(w_n1045_0[0]),.doutb(w_n1045_0[1]),.din(n1045));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(n1048));
	jspl3 jspl3_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.doutc(w_n1053_0[2]),.din(n1053));
	jspl jspl_w_n1056_0(.douta(w_n1056_0[0]),.doutb(w_n1056_0[1]),.din(n1056));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.din(n1062));
	jspl jspl_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.din(n1091));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl3 jspl3_w_n1159_0(.douta(w_n1159_0[0]),.doutb(w_n1159_0[1]),.doutc(w_n1159_0[2]),.din(n1159));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(n1161));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(w_dff_B_HpHtOqHA3_2));
	jspl jspl_w_n1168_0(.douta(w_n1168_0[0]),.doutb(w_n1168_0[1]),.din(n1168));
	jspl jspl_w_n1170_0(.douta(w_n1170_0[0]),.doutb(w_n1170_0[1]),.din(n1170));
	jspl jspl_w_n1177_0(.douta(w_n1177_0[0]),.doutb(w_dff_A_5UrYmzix0_1),.din(w_dff_B_HFykTtMo5_2));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.din(n1178));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.din(n1184));
	jdff dff_B_xHjQUWcM6_1(.din(n92),.dout(w_dff_B_xHjQUWcM6_1),.clk(gclk));
	jdff dff_B_VjmlfsDy9_1(.din(w_dff_B_xHjQUWcM6_1),.dout(w_dff_B_VjmlfsDy9_1),.clk(gclk));
	jdff dff_B_Mt4cKI405_1(.din(w_dff_B_VjmlfsDy9_1),.dout(w_dff_B_Mt4cKI405_1),.clk(gclk));
	jdff dff_B_HQ7X0MvH1_1(.din(n583),.dout(w_dff_B_HQ7X0MvH1_1),.clk(gclk));
	jdff dff_B_22bVWtfL0_1(.din(w_dff_B_HQ7X0MvH1_1),.dout(w_dff_B_22bVWtfL0_1),.clk(gclk));
	jdff dff_B_2TT2DMn67_1(.din(w_dff_B_22bVWtfL0_1),.dout(w_dff_B_2TT2DMn67_1),.clk(gclk));
	jdff dff_B_QVk4dQrZ1_1(.din(w_dff_B_2TT2DMn67_1),.dout(w_dff_B_QVk4dQrZ1_1),.clk(gclk));
	jdff dff_B_oLBQvcT41_1(.din(w_dff_B_QVk4dQrZ1_1),.dout(w_dff_B_oLBQvcT41_1),.clk(gclk));
	jdff dff_B_kwkvJeIU9_1(.din(w_dff_B_oLBQvcT41_1),.dout(w_dff_B_kwkvJeIU9_1),.clk(gclk));
	jdff dff_B_TGoVpYEx6_1(.din(w_dff_B_kwkvJeIU9_1),.dout(w_dff_B_TGoVpYEx6_1),.clk(gclk));
	jdff dff_B_Fk2wDTnf3_1(.din(w_dff_B_TGoVpYEx6_1),.dout(w_dff_B_Fk2wDTnf3_1),.clk(gclk));
	jdff dff_B_5snqWQgf3_1(.din(w_dff_B_Fk2wDTnf3_1),.dout(w_dff_B_5snqWQgf3_1),.clk(gclk));
	jdff dff_B_634dszOY3_1(.din(w_dff_B_5snqWQgf3_1),.dout(w_dff_B_634dszOY3_1),.clk(gclk));
	jdff dff_B_6pWQF2Zt3_1(.din(w_dff_B_634dszOY3_1),.dout(w_dff_B_6pWQF2Zt3_1),.clk(gclk));
	jdff dff_B_A7SfOkGb4_1(.din(w_dff_B_6pWQF2Zt3_1),.dout(w_dff_B_A7SfOkGb4_1),.clk(gclk));
	jdff dff_B_J0H42DkE9_1(.din(w_dff_B_A7SfOkGb4_1),.dout(w_dff_B_J0H42DkE9_1),.clk(gclk));
	jdff dff_B_sccYniaQ7_1(.din(w_dff_B_J0H42DkE9_1),.dout(w_dff_B_sccYniaQ7_1),.clk(gclk));
	jdff dff_B_IexGRyFg3_1(.din(w_dff_B_sccYniaQ7_1),.dout(w_dff_B_IexGRyFg3_1),.clk(gclk));
	jdff dff_B_ueFBhWi45_1(.din(w_dff_B_IexGRyFg3_1),.dout(w_dff_B_ueFBhWi45_1),.clk(gclk));
	jdff dff_B_u0KPQAqv5_0(.din(n795),.dout(w_dff_B_u0KPQAqv5_0),.clk(gclk));
	jdff dff_B_2GVCeahx4_0(.din(w_dff_B_u0KPQAqv5_0),.dout(w_dff_B_2GVCeahx4_0),.clk(gclk));
	jdff dff_B_WysWk24V4_0(.din(w_dff_B_2GVCeahx4_0),.dout(w_dff_B_WysWk24V4_0),.clk(gclk));
	jdff dff_B_FOEMFtkR0_0(.din(w_dff_B_WysWk24V4_0),.dout(w_dff_B_FOEMFtkR0_0),.clk(gclk));
	jdff dff_B_BylPbcSb9_0(.din(w_dff_B_FOEMFtkR0_0),.dout(w_dff_B_BylPbcSb9_0),.clk(gclk));
	jdff dff_B_SCuwsZ4y1_0(.din(w_dff_B_BylPbcSb9_0),.dout(w_dff_B_SCuwsZ4y1_0),.clk(gclk));
	jdff dff_B_UOhUKV8Q1_0(.din(w_dff_B_SCuwsZ4y1_0),.dout(w_dff_B_UOhUKV8Q1_0),.clk(gclk));
	jdff dff_B_urnAEHxh0_0(.din(w_dff_B_UOhUKV8Q1_0),.dout(w_dff_B_urnAEHxh0_0),.clk(gclk));
	jdff dff_B_1ST408VS9_0(.din(w_dff_B_urnAEHxh0_0),.dout(w_dff_B_1ST408VS9_0),.clk(gclk));
	jdff dff_B_RDDKxhKt5_0(.din(w_dff_B_1ST408VS9_0),.dout(w_dff_B_RDDKxhKt5_0),.clk(gclk));
	jdff dff_B_DTkC4zXD7_0(.din(w_dff_B_RDDKxhKt5_0),.dout(w_dff_B_DTkC4zXD7_0),.clk(gclk));
	jdff dff_B_MnaE5uDC8_0(.din(w_dff_B_DTkC4zXD7_0),.dout(w_dff_B_MnaE5uDC8_0),.clk(gclk));
	jdff dff_B_VnxhVx6Z9_0(.din(w_dff_B_MnaE5uDC8_0),.dout(w_dff_B_VnxhVx6Z9_0),.clk(gclk));
	jdff dff_B_Gcvpk43x2_0(.din(w_dff_B_VnxhVx6Z9_0),.dout(w_dff_B_Gcvpk43x2_0),.clk(gclk));
	jdff dff_B_9oyPHs7g1_0(.din(w_dff_B_Gcvpk43x2_0),.dout(w_dff_B_9oyPHs7g1_0),.clk(gclk));
	jdff dff_B_OQBD1u0p4_0(.din(w_dff_B_9oyPHs7g1_0),.dout(w_dff_B_OQBD1u0p4_0),.clk(gclk));
	jdff dff_B_Q2OW7rOi7_0(.din(w_dff_B_OQBD1u0p4_0),.dout(w_dff_B_Q2OW7rOi7_0),.clk(gclk));
	jdff dff_B_q6bNldw60_1(.din(n1171),.dout(w_dff_B_q6bNldw60_1),.clk(gclk));
	jdff dff_B_l3lZnQLq9_1(.din(w_dff_B_q6bNldw60_1),.dout(w_dff_B_l3lZnQLq9_1),.clk(gclk));
	jdff dff_B_jnLKg6zc8_1(.din(n1172),.dout(w_dff_B_jnLKg6zc8_1),.clk(gclk));
	jdff dff_B_YQWUqsGM8_1(.din(w_dff_B_jnLKg6zc8_1),.dout(w_dff_B_YQWUqsGM8_1),.clk(gclk));
	jdff dff_B_xqUFUO7K0_1(.din(w_dff_B_YQWUqsGM8_1),.dout(w_dff_B_xqUFUO7K0_1),.clk(gclk));
	jdff dff_B_QMLcvk0t1_1(.din(w_dff_B_xqUFUO7K0_1),.dout(w_dff_B_QMLcvk0t1_1),.clk(gclk));
	jdff dff_B_rfz4CH6Q5_1(.din(w_dff_B_QMLcvk0t1_1),.dout(w_dff_B_rfz4CH6Q5_1),.clk(gclk));
	jdff dff_B_AWJ7WFQe3_1(.din(w_dff_B_rfz4CH6Q5_1),.dout(w_dff_B_AWJ7WFQe3_1),.clk(gclk));
	jdff dff_B_ta9doG5X1_1(.din(w_dff_B_AWJ7WFQe3_1),.dout(w_dff_B_ta9doG5X1_1),.clk(gclk));
	jdff dff_B_2aULs05t3_1(.din(w_dff_B_ta9doG5X1_1),.dout(w_dff_B_2aULs05t3_1),.clk(gclk));
	jdff dff_B_1e8Tsy3Y7_1(.din(w_dff_B_2aULs05t3_1),.dout(w_dff_B_1e8Tsy3Y7_1),.clk(gclk));
	jdff dff_B_jriraDas1_1(.din(w_dff_B_1e8Tsy3Y7_1),.dout(w_dff_B_jriraDas1_1),.clk(gclk));
	jdff dff_B_lzlWFihn9_1(.din(w_dff_B_jriraDas1_1),.dout(w_dff_B_lzlWFihn9_1),.clk(gclk));
	jdff dff_B_0solhEAT9_1(.din(w_dff_B_lzlWFihn9_1),.dout(w_dff_B_0solhEAT9_1),.clk(gclk));
	jdff dff_B_JlIj0nb70_1(.din(w_dff_B_0solhEAT9_1),.dout(w_dff_B_JlIj0nb70_1),.clk(gclk));
	jdff dff_B_9hCywfez2_1(.din(w_dff_B_JlIj0nb70_1),.dout(w_dff_B_9hCywfez2_1),.clk(gclk));
	jdff dff_B_TpzJBJHo9_1(.din(w_dff_B_9hCywfez2_1),.dout(w_dff_B_TpzJBJHo9_1),.clk(gclk));
	jdff dff_B_03WS732s8_1(.din(w_dff_B_TpzJBJHo9_1),.dout(w_dff_B_03WS732s8_1),.clk(gclk));
	jdff dff_B_X6R4aNGE6_1(.din(w_dff_B_03WS732s8_1),.dout(w_dff_B_X6R4aNGE6_1),.clk(gclk));
	jdff dff_B_L8RNaC5U4_1(.din(w_dff_B_X6R4aNGE6_1),.dout(w_dff_B_L8RNaC5U4_1),.clk(gclk));
	jdff dff_B_81gzoYDd3_1(.din(w_dff_B_L8RNaC5U4_1),.dout(w_dff_B_81gzoYDd3_1),.clk(gclk));
	jdff dff_B_8rdXXyPZ7_1(.din(w_dff_B_81gzoYDd3_1),.dout(w_dff_B_8rdXXyPZ7_1),.clk(gclk));
	jdff dff_B_QhvOIY9O8_1(.din(w_dff_B_8rdXXyPZ7_1),.dout(w_dff_B_QhvOIY9O8_1),.clk(gclk));
	jdff dff_B_eGGmHCC48_1(.din(w_dff_B_QhvOIY9O8_1),.dout(w_dff_B_eGGmHCC48_1),.clk(gclk));
	jdff dff_B_lXd2Awnt0_1(.din(w_dff_B_eGGmHCC48_1),.dout(w_dff_B_lXd2Awnt0_1),.clk(gclk));
	jdff dff_B_bOsBCVpY4_1(.din(w_dff_B_lXd2Awnt0_1),.dout(w_dff_B_bOsBCVpY4_1),.clk(gclk));
	jdff dff_B_prp0mfij9_1(.din(w_dff_B_bOsBCVpY4_1),.dout(w_dff_B_prp0mfij9_1),.clk(gclk));
	jdff dff_B_j8FbVouI0_1(.din(w_dff_B_prp0mfij9_1),.dout(w_dff_B_j8FbVouI0_1),.clk(gclk));
	jdff dff_B_mu9n9ilP0_1(.din(w_dff_B_j8FbVouI0_1),.dout(w_dff_B_mu9n9ilP0_1),.clk(gclk));
	jdff dff_B_0ZaFb6Dc1_1(.din(w_dff_B_mu9n9ilP0_1),.dout(w_dff_B_0ZaFb6Dc1_1),.clk(gclk));
	jdff dff_B_c7VrnfJj6_0(.din(n1166),.dout(w_dff_B_c7VrnfJj6_0),.clk(gclk));
	jdff dff_B_9zpnASnZ7_0(.din(n1165),.dout(w_dff_B_9zpnASnZ7_0),.clk(gclk));
	jdff dff_B_muoYqJAP6_1(.din(n1182),.dout(w_dff_B_muoYqJAP6_1),.clk(gclk));
	jdff dff_B_zWiukuNG3_1(.din(w_dff_B_muoYqJAP6_1),.dout(w_dff_B_zWiukuNG3_1),.clk(gclk));
	jdff dff_B_WdUXIHfI8_1(.din(w_dff_B_zWiukuNG3_1),.dout(w_dff_B_WdUXIHfI8_1),.clk(gclk));
	jdff dff_B_exGhWo893_1(.din(w_dff_B_WdUXIHfI8_1),.dout(w_dff_B_exGhWo893_1),.clk(gclk));
	jdff dff_B_KuRzPd3r4_1(.din(w_dff_B_exGhWo893_1),.dout(w_dff_B_KuRzPd3r4_1),.clk(gclk));
	jdff dff_B_jPnidbuk4_1(.din(w_dff_B_KuRzPd3r4_1),.dout(w_dff_B_jPnidbuk4_1),.clk(gclk));
	jdff dff_B_WGNNI6Js1_1(.din(w_dff_B_jPnidbuk4_1),.dout(w_dff_B_WGNNI6Js1_1),.clk(gclk));
	jdff dff_B_e9ZR4Lw22_1(.din(w_dff_B_WGNNI6Js1_1),.dout(w_dff_B_e9ZR4Lw22_1),.clk(gclk));
	jdff dff_B_jZtfpIr95_1(.din(w_dff_B_e9ZR4Lw22_1),.dout(w_dff_B_jZtfpIr95_1),.clk(gclk));
	jdff dff_B_Ut40zb8L0_1(.din(w_dff_B_jZtfpIr95_1),.dout(w_dff_B_Ut40zb8L0_1),.clk(gclk));
	jdff dff_B_Gedsz2kC2_1(.din(w_dff_B_Ut40zb8L0_1),.dout(w_dff_B_Gedsz2kC2_1),.clk(gclk));
	jdff dff_B_ACEyuKxm7_1(.din(w_dff_B_Gedsz2kC2_1),.dout(w_dff_B_ACEyuKxm7_1),.clk(gclk));
	jdff dff_B_6lU5nar68_1(.din(w_dff_B_ACEyuKxm7_1),.dout(w_dff_B_6lU5nar68_1),.clk(gclk));
	jdff dff_B_T2cfWnkw0_1(.din(w_dff_B_6lU5nar68_1),.dout(w_dff_B_T2cfWnkw0_1),.clk(gclk));
	jdff dff_B_IdKWaz1P7_1(.din(w_dff_B_T2cfWnkw0_1),.dout(w_dff_B_IdKWaz1P7_1),.clk(gclk));
	jdff dff_B_EtTGXOoa6_1(.din(w_dff_B_IdKWaz1P7_1),.dout(w_dff_B_EtTGXOoa6_1),.clk(gclk));
	jdff dff_B_Gb5dMDpc1_1(.din(w_dff_B_EtTGXOoa6_1),.dout(w_dff_B_Gb5dMDpc1_1),.clk(gclk));
	jdff dff_B_DvcwlsgN3_1(.din(w_dff_B_Gb5dMDpc1_1),.dout(w_dff_B_DvcwlsgN3_1),.clk(gclk));
	jdff dff_B_xHL8CGM99_1(.din(w_dff_B_DvcwlsgN3_1),.dout(w_dff_B_xHL8CGM99_1),.clk(gclk));
	jdff dff_B_3uApdKyi9_1(.din(w_dff_B_xHL8CGM99_1),.dout(w_dff_B_3uApdKyi9_1),.clk(gclk));
	jdff dff_B_7ldL9vkR7_1(.din(w_dff_B_3uApdKyi9_1),.dout(w_dff_B_7ldL9vkR7_1),.clk(gclk));
	jdff dff_B_yGM9w70N1_1(.din(w_dff_B_7ldL9vkR7_1),.dout(w_dff_B_yGM9w70N1_1),.clk(gclk));
	jdff dff_B_vqt2ixL65_1(.din(w_dff_B_yGM9w70N1_1),.dout(w_dff_B_vqt2ixL65_1),.clk(gclk));
	jdff dff_B_SLNhhTuD3_1(.din(w_dff_B_vqt2ixL65_1),.dout(w_dff_B_SLNhhTuD3_1),.clk(gclk));
	jdff dff_B_wCBFBJ289_1(.din(w_dff_B_SLNhhTuD3_1),.dout(w_dff_B_wCBFBJ289_1),.clk(gclk));
	jdff dff_B_r16mdVyf5_1(.din(G2897),.dout(w_dff_B_r16mdVyf5_1),.clk(gclk));
	jdff dff_B_R0y0XQyz9_1(.din(w_dff_B_r16mdVyf5_1),.dout(w_dff_B_R0y0XQyz9_1),.clk(gclk));
	jdff dff_B_mV3DpgdJ3_1(.din(w_dff_B_R0y0XQyz9_1),.dout(w_dff_B_mV3DpgdJ3_1),.clk(gclk));
	jdff dff_B_71ZeuXyD3_1(.din(w_dff_B_mV3DpgdJ3_1),.dout(w_dff_B_71ZeuXyD3_1),.clk(gclk));
	jdff dff_B_ieRAh7pn1_1(.din(w_dff_B_71ZeuXyD3_1),.dout(w_dff_B_ieRAh7pn1_1),.clk(gclk));
	jdff dff_B_jgDIuOm97_1(.din(w_dff_B_ieRAh7pn1_1),.dout(w_dff_B_jgDIuOm97_1),.clk(gclk));
	jdff dff_B_0qLziPTL0_1(.din(w_dff_B_jgDIuOm97_1),.dout(w_dff_B_0qLziPTL0_1),.clk(gclk));
	jdff dff_B_KHiWN5fs7_1(.din(w_dff_B_0qLziPTL0_1),.dout(w_dff_B_KHiWN5fs7_1),.clk(gclk));
	jdff dff_B_Kwx5Zzrv2_1(.din(w_dff_B_KHiWN5fs7_1),.dout(w_dff_B_Kwx5Zzrv2_1),.clk(gclk));
	jdff dff_B_BLn13hMk0_1(.din(w_dff_B_Kwx5Zzrv2_1),.dout(w_dff_B_BLn13hMk0_1),.clk(gclk));
	jdff dff_B_cBrdFfoY9_1(.din(w_dff_B_BLn13hMk0_1),.dout(w_dff_B_cBrdFfoY9_1),.clk(gclk));
	jdff dff_B_xpplfx8y9_1(.din(w_dff_B_cBrdFfoY9_1),.dout(w_dff_B_xpplfx8y9_1),.clk(gclk));
	jdff dff_B_TpYVZ56u7_1(.din(w_dff_B_xpplfx8y9_1),.dout(w_dff_B_TpYVZ56u7_1),.clk(gclk));
	jdff dff_B_Lk0aWGUz5_1(.din(w_dff_B_TpYVZ56u7_1),.dout(w_dff_B_Lk0aWGUz5_1),.clk(gclk));
	jdff dff_B_vNB21VeQ7_1(.din(w_dff_B_Lk0aWGUz5_1),.dout(w_dff_B_vNB21VeQ7_1),.clk(gclk));
	jdff dff_B_TueIlBv25_1(.din(w_dff_B_vNB21VeQ7_1),.dout(w_dff_B_TueIlBv25_1),.clk(gclk));
	jdff dff_B_ZHeLmu9d1_1(.din(w_dff_B_TueIlBv25_1),.dout(w_dff_B_ZHeLmu9d1_1),.clk(gclk));
	jdff dff_B_wOe0PS6z4_1(.din(w_dff_B_ZHeLmu9d1_1),.dout(w_dff_B_wOe0PS6z4_1),.clk(gclk));
	jdff dff_B_4oi2hvdW4_1(.din(w_dff_B_wOe0PS6z4_1),.dout(w_dff_B_4oi2hvdW4_1),.clk(gclk));
	jdff dff_B_DJfgBu7q6_1(.din(w_dff_B_4oi2hvdW4_1),.dout(w_dff_B_DJfgBu7q6_1),.clk(gclk));
	jdff dff_B_wJFwYcwK6_1(.din(w_dff_B_DJfgBu7q6_1),.dout(w_dff_B_wJFwYcwK6_1),.clk(gclk));
	jdff dff_B_zsuITUe04_1(.din(w_dff_B_wJFwYcwK6_1),.dout(w_dff_B_zsuITUe04_1),.clk(gclk));
	jdff dff_B_PgYY4vUx7_1(.din(w_dff_B_zsuITUe04_1),.dout(w_dff_B_PgYY4vUx7_1),.clk(gclk));
	jdff dff_B_tyELKyBq2_1(.din(w_dff_B_PgYY4vUx7_1),.dout(w_dff_B_tyELKyBq2_1),.clk(gclk));
	jdff dff_B_ROu1pqix5_1(.din(w_dff_B_tyELKyBq2_1),.dout(w_dff_B_ROu1pqix5_1),.clk(gclk));
	jdff dff_B_PC9xXn8s6_1(.din(w_dff_B_ROu1pqix5_1),.dout(w_dff_B_PC9xXn8s6_1),.clk(gclk));
	jdff dff_B_C4JZ1NsH6_1(.din(w_dff_B_PC9xXn8s6_1),.dout(w_dff_B_C4JZ1NsH6_1),.clk(gclk));
	jdff dff_A_1cQEWpcD0_0(.dout(w_G384_0),.din(w_dff_A_1cQEWpcD0_0),.clk(gclk));
	jdff dff_A_nEeQ9yMU7_0(.dout(w_dff_A_1cQEWpcD0_0),.din(w_dff_A_nEeQ9yMU7_0),.clk(gclk));
	jdff dff_A_BhJhL6gc7_0(.dout(w_dff_A_nEeQ9yMU7_0),.din(w_dff_A_BhJhL6gc7_0),.clk(gclk));
	jdff dff_A_0bqHEcZ56_1(.dout(w_n1177_0[1]),.din(w_dff_A_0bqHEcZ56_1),.clk(gclk));
	jdff dff_A_5UrYmzix0_1(.dout(w_dff_A_0bqHEcZ56_1),.din(w_dff_A_5UrYmzix0_1),.clk(gclk));
	jdff dff_B_lHnJ19Zu1_2(.din(n1177),.dout(w_dff_B_lHnJ19Zu1_2),.clk(gclk));
	jdff dff_B_HFykTtMo5_2(.din(w_dff_B_lHnJ19Zu1_2),.dout(w_dff_B_HFykTtMo5_2),.clk(gclk));
	jdff dff_B_nAxUj1iK8_1(.din(n1175),.dout(w_dff_B_nAxUj1iK8_1),.clk(gclk));
	jdff dff_B_FAEdZJEp2_2(.din(n1164),.dout(w_dff_B_FAEdZJEp2_2),.clk(gclk));
	jdff dff_B_tXLhldf20_2(.din(w_dff_B_FAEdZJEp2_2),.dout(w_dff_B_tXLhldf20_2),.clk(gclk));
	jdff dff_B_gUkXXbu39_2(.din(w_dff_B_tXLhldf20_2),.dout(w_dff_B_gUkXXbu39_2),.clk(gclk));
	jdff dff_B_HpHtOqHA3_2(.din(w_dff_B_gUkXXbu39_2),.dout(w_dff_B_HpHtOqHA3_2),.clk(gclk));
	jdff dff_B_DNikSduU6_1(.din(n617),.dout(w_dff_B_DNikSduU6_1),.clk(gclk));
	jdff dff_B_pETUV4B08_0(.din(n698),.dout(w_dff_B_pETUV4B08_0),.clk(gclk));
	jdff dff_B_CyQrIu989_0(.din(n697),.dout(w_dff_B_CyQrIu989_0),.clk(gclk));
	jdff dff_B_P6gvEx497_0(.din(w_dff_B_CyQrIu989_0),.dout(w_dff_B_P6gvEx497_0),.clk(gclk));
	jdff dff_B_BdB41wc63_0(.din(n694),.dout(w_dff_B_BdB41wc63_0),.clk(gclk));
	jdff dff_B_QI4QLR1u6_0(.din(w_dff_B_BdB41wc63_0),.dout(w_dff_B_QI4QLR1u6_0),.clk(gclk));
	jdff dff_A_z3QgeTlH5_0(.dout(w_G355_0),.din(w_dff_A_z3QgeTlH5_0),.clk(gclk));
	jdff dff_A_rykcEi9w2_2(.dout(w_dff_A_7tXAyvIc9_0),.din(w_dff_A_rykcEi9w2_2),.clk(gclk));
	jdff dff_A_7tXAyvIc9_0(.dout(w_dff_A_sJ26Vx1O7_0),.din(w_dff_A_7tXAyvIc9_0),.clk(gclk));
	jdff dff_A_sJ26Vx1O7_0(.dout(w_dff_A_J6sjkAqq8_0),.din(w_dff_A_sJ26Vx1O7_0),.clk(gclk));
	jdff dff_A_J6sjkAqq8_0(.dout(w_dff_A_bvAV8NCD6_0),.din(w_dff_A_J6sjkAqq8_0),.clk(gclk));
	jdff dff_A_bvAV8NCD6_0(.dout(w_dff_A_78xeVvM67_0),.din(w_dff_A_bvAV8NCD6_0),.clk(gclk));
	jdff dff_A_78xeVvM67_0(.dout(w_dff_A_8ZrYs9dv9_0),.din(w_dff_A_78xeVvM67_0),.clk(gclk));
	jdff dff_A_8ZrYs9dv9_0(.dout(w_dff_A_q9YlF5aK2_0),.din(w_dff_A_8ZrYs9dv9_0),.clk(gclk));
	jdff dff_A_q9YlF5aK2_0(.dout(w_dff_A_aCiwPFen2_0),.din(w_dff_A_q9YlF5aK2_0),.clk(gclk));
	jdff dff_A_aCiwPFen2_0(.dout(w_dff_A_BrII8quO0_0),.din(w_dff_A_aCiwPFen2_0),.clk(gclk));
	jdff dff_A_BrII8quO0_0(.dout(w_dff_A_BNxYVpX82_0),.din(w_dff_A_BrII8quO0_0),.clk(gclk));
	jdff dff_A_BNxYVpX82_0(.dout(w_dff_A_pLGlTChb9_0),.din(w_dff_A_BNxYVpX82_0),.clk(gclk));
	jdff dff_A_pLGlTChb9_0(.dout(w_dff_A_wlGAPGV14_0),.din(w_dff_A_pLGlTChb9_0),.clk(gclk));
	jdff dff_A_wlGAPGV14_0(.dout(w_dff_A_ACPekjjV3_0),.din(w_dff_A_wlGAPGV14_0),.clk(gclk));
	jdff dff_A_ACPekjjV3_0(.dout(w_dff_A_XW192r1e4_0),.din(w_dff_A_ACPekjjV3_0),.clk(gclk));
	jdff dff_A_XW192r1e4_0(.dout(w_dff_A_Ov05VS1I6_0),.din(w_dff_A_XW192r1e4_0),.clk(gclk));
	jdff dff_A_Ov05VS1I6_0(.dout(w_dff_A_Ehf5bj7o1_0),.din(w_dff_A_Ov05VS1I6_0),.clk(gclk));
	jdff dff_A_Ehf5bj7o1_0(.dout(w_dff_A_BCEjLeVG1_0),.din(w_dff_A_Ehf5bj7o1_0),.clk(gclk));
	jdff dff_A_BCEjLeVG1_0(.dout(w_dff_A_Na8c8buW1_0),.din(w_dff_A_BCEjLeVG1_0),.clk(gclk));
	jdff dff_A_Na8c8buW1_0(.dout(w_dff_A_9nOBslLD0_0),.din(w_dff_A_Na8c8buW1_0),.clk(gclk));
	jdff dff_A_9nOBslLD0_0(.dout(w_dff_A_TxiSdO7Q1_0),.din(w_dff_A_9nOBslLD0_0),.clk(gclk));
	jdff dff_A_TxiSdO7Q1_0(.dout(w_dff_A_0PKeuSai9_0),.din(w_dff_A_TxiSdO7Q1_0),.clk(gclk));
	jdff dff_A_0PKeuSai9_0(.dout(w_dff_A_vBFf419J5_0),.din(w_dff_A_0PKeuSai9_0),.clk(gclk));
	jdff dff_A_vBFf419J5_0(.dout(w_dff_A_Bc4lmPKi8_0),.din(w_dff_A_vBFf419J5_0),.clk(gclk));
	jdff dff_A_Bc4lmPKi8_0(.dout(w_dff_A_RDsEoRlQ8_0),.din(w_dff_A_Bc4lmPKi8_0),.clk(gclk));
	jdff dff_A_RDsEoRlQ8_0(.dout(w_dff_A_EQGyNptT1_0),.din(w_dff_A_RDsEoRlQ8_0),.clk(gclk));
	jdff dff_A_EQGyNptT1_0(.dout(w_dff_A_2ex2bB0s2_0),.din(w_dff_A_EQGyNptT1_0),.clk(gclk));
	jdff dff_A_2ex2bB0s2_0(.dout(G353),.din(w_dff_A_2ex2bB0s2_0),.clk(gclk));
	jdff dff_A_iY0rTqRq8_1(.dout(w_dff_A_lYvf9yv19_0),.din(w_dff_A_iY0rTqRq8_1),.clk(gclk));
	jdff dff_A_lYvf9yv19_0(.dout(w_dff_A_aAa5JjEc7_0),.din(w_dff_A_lYvf9yv19_0),.clk(gclk));
	jdff dff_A_aAa5JjEc7_0(.dout(w_dff_A_Fhngsv7p4_0),.din(w_dff_A_aAa5JjEc7_0),.clk(gclk));
	jdff dff_A_Fhngsv7p4_0(.dout(w_dff_A_IiXeey773_0),.din(w_dff_A_Fhngsv7p4_0),.clk(gclk));
	jdff dff_A_IiXeey773_0(.dout(w_dff_A_sbaw8oi15_0),.din(w_dff_A_IiXeey773_0),.clk(gclk));
	jdff dff_A_sbaw8oi15_0(.dout(w_dff_A_wCgExy7V3_0),.din(w_dff_A_sbaw8oi15_0),.clk(gclk));
	jdff dff_A_wCgExy7V3_0(.dout(w_dff_A_a7QWWlo49_0),.din(w_dff_A_wCgExy7V3_0),.clk(gclk));
	jdff dff_A_a7QWWlo49_0(.dout(w_dff_A_97MhZySN7_0),.din(w_dff_A_a7QWWlo49_0),.clk(gclk));
	jdff dff_A_97MhZySN7_0(.dout(w_dff_A_fXNCu55L5_0),.din(w_dff_A_97MhZySN7_0),.clk(gclk));
	jdff dff_A_fXNCu55L5_0(.dout(w_dff_A_noLTKY9K1_0),.din(w_dff_A_fXNCu55L5_0),.clk(gclk));
	jdff dff_A_noLTKY9K1_0(.dout(w_dff_A_s8ZpllIO5_0),.din(w_dff_A_noLTKY9K1_0),.clk(gclk));
	jdff dff_A_s8ZpllIO5_0(.dout(w_dff_A_rRYQwDuV9_0),.din(w_dff_A_s8ZpllIO5_0),.clk(gclk));
	jdff dff_A_rRYQwDuV9_0(.dout(w_dff_A_wVhcwU9y1_0),.din(w_dff_A_rRYQwDuV9_0),.clk(gclk));
	jdff dff_A_wVhcwU9y1_0(.dout(w_dff_A_AA0t5bqS3_0),.din(w_dff_A_wVhcwU9y1_0),.clk(gclk));
	jdff dff_A_AA0t5bqS3_0(.dout(w_dff_A_x8DSkExS1_0),.din(w_dff_A_AA0t5bqS3_0),.clk(gclk));
	jdff dff_A_x8DSkExS1_0(.dout(w_dff_A_2rCmqjTR3_0),.din(w_dff_A_x8DSkExS1_0),.clk(gclk));
	jdff dff_A_2rCmqjTR3_0(.dout(w_dff_A_pzAxV5YN0_0),.din(w_dff_A_2rCmqjTR3_0),.clk(gclk));
	jdff dff_A_pzAxV5YN0_0(.dout(w_dff_A_1pWOxKmm2_0),.din(w_dff_A_pzAxV5YN0_0),.clk(gclk));
	jdff dff_A_1pWOxKmm2_0(.dout(w_dff_A_vXqGkER71_0),.din(w_dff_A_1pWOxKmm2_0),.clk(gclk));
	jdff dff_A_vXqGkER71_0(.dout(w_dff_A_74NmZsTt6_0),.din(w_dff_A_vXqGkER71_0),.clk(gclk));
	jdff dff_A_74NmZsTt6_0(.dout(w_dff_A_NUL87zGZ7_0),.din(w_dff_A_74NmZsTt6_0),.clk(gclk));
	jdff dff_A_NUL87zGZ7_0(.dout(w_dff_A_HwuPOGwD1_0),.din(w_dff_A_NUL87zGZ7_0),.clk(gclk));
	jdff dff_A_HwuPOGwD1_0(.dout(w_dff_A_VgBe6X6X6_0),.din(w_dff_A_HwuPOGwD1_0),.clk(gclk));
	jdff dff_A_VgBe6X6X6_0(.dout(w_dff_A_k0bEhgrd6_0),.din(w_dff_A_VgBe6X6X6_0),.clk(gclk));
	jdff dff_A_k0bEhgrd6_0(.dout(w_dff_A_87qaW5RV8_0),.din(w_dff_A_k0bEhgrd6_0),.clk(gclk));
	jdff dff_A_87qaW5RV8_0(.dout(w_dff_A_oQ8HNp3w4_0),.din(w_dff_A_87qaW5RV8_0),.clk(gclk));
	jdff dff_A_oQ8HNp3w4_0(.dout(w_dff_A_n7f1N90w6_0),.din(w_dff_A_oQ8HNp3w4_0),.clk(gclk));
	jdff dff_A_n7f1N90w6_0(.dout(G355),.din(w_dff_A_n7f1N90w6_0),.clk(gclk));
	jdff dff_A_tGv9QlUg2_2(.dout(w_dff_A_3x64q4q06_0),.din(w_dff_A_tGv9QlUg2_2),.clk(gclk));
	jdff dff_A_3x64q4q06_0(.dout(w_dff_A_8zTbKcVM5_0),.din(w_dff_A_3x64q4q06_0),.clk(gclk));
	jdff dff_A_8zTbKcVM5_0(.dout(w_dff_A_WcRpnLv47_0),.din(w_dff_A_8zTbKcVM5_0),.clk(gclk));
	jdff dff_A_WcRpnLv47_0(.dout(w_dff_A_VWMlx0DM4_0),.din(w_dff_A_WcRpnLv47_0),.clk(gclk));
	jdff dff_A_VWMlx0DM4_0(.dout(w_dff_A_SRswPu2g9_0),.din(w_dff_A_VWMlx0DM4_0),.clk(gclk));
	jdff dff_A_SRswPu2g9_0(.dout(w_dff_A_dsW8gz3d1_0),.din(w_dff_A_SRswPu2g9_0),.clk(gclk));
	jdff dff_A_dsW8gz3d1_0(.dout(w_dff_A_9nxvnyL83_0),.din(w_dff_A_dsW8gz3d1_0),.clk(gclk));
	jdff dff_A_9nxvnyL83_0(.dout(w_dff_A_rjysqVXr3_0),.din(w_dff_A_9nxvnyL83_0),.clk(gclk));
	jdff dff_A_rjysqVXr3_0(.dout(w_dff_A_1MMwLd568_0),.din(w_dff_A_rjysqVXr3_0),.clk(gclk));
	jdff dff_A_1MMwLd568_0(.dout(w_dff_A_mplGl4XJ4_0),.din(w_dff_A_1MMwLd568_0),.clk(gclk));
	jdff dff_A_mplGl4XJ4_0(.dout(w_dff_A_RBGPa3Sa1_0),.din(w_dff_A_mplGl4XJ4_0),.clk(gclk));
	jdff dff_A_RBGPa3Sa1_0(.dout(w_dff_A_JJoZgGzJ0_0),.din(w_dff_A_RBGPa3Sa1_0),.clk(gclk));
	jdff dff_A_JJoZgGzJ0_0(.dout(w_dff_A_1ERsv94T0_0),.din(w_dff_A_JJoZgGzJ0_0),.clk(gclk));
	jdff dff_A_1ERsv94T0_0(.dout(w_dff_A_zuCevQOC5_0),.din(w_dff_A_1ERsv94T0_0),.clk(gclk));
	jdff dff_A_zuCevQOC5_0(.dout(w_dff_A_8uszQAbC5_0),.din(w_dff_A_zuCevQOC5_0),.clk(gclk));
	jdff dff_A_8uszQAbC5_0(.dout(w_dff_A_C8aYFkpA1_0),.din(w_dff_A_8uszQAbC5_0),.clk(gclk));
	jdff dff_A_C8aYFkpA1_0(.dout(w_dff_A_nsIxJLQ78_0),.din(w_dff_A_C8aYFkpA1_0),.clk(gclk));
	jdff dff_A_nsIxJLQ78_0(.dout(w_dff_A_zXV78VOh4_0),.din(w_dff_A_nsIxJLQ78_0),.clk(gclk));
	jdff dff_A_zXV78VOh4_0(.dout(w_dff_A_Zhpbic7e7_0),.din(w_dff_A_zXV78VOh4_0),.clk(gclk));
	jdff dff_A_Zhpbic7e7_0(.dout(w_dff_A_WZikTYSU2_0),.din(w_dff_A_Zhpbic7e7_0),.clk(gclk));
	jdff dff_A_WZikTYSU2_0(.dout(w_dff_A_UJ6dkv765_0),.din(w_dff_A_WZikTYSU2_0),.clk(gclk));
	jdff dff_A_UJ6dkv765_0(.dout(w_dff_A_iNnPeafG1_0),.din(w_dff_A_UJ6dkv765_0),.clk(gclk));
	jdff dff_A_iNnPeafG1_0(.dout(G361),.din(w_dff_A_iNnPeafG1_0),.clk(gclk));
	jdff dff_A_FASwSrM37_2(.dout(w_dff_A_dces0ZHC1_0),.din(w_dff_A_FASwSrM37_2),.clk(gclk));
	jdff dff_A_dces0ZHC1_0(.dout(w_dff_A_RT13c4cr8_0),.din(w_dff_A_dces0ZHC1_0),.clk(gclk));
	jdff dff_A_RT13c4cr8_0(.dout(w_dff_A_2TFo5LhC0_0),.din(w_dff_A_RT13c4cr8_0),.clk(gclk));
	jdff dff_A_2TFo5LhC0_0(.dout(w_dff_A_o5jm3Mm81_0),.din(w_dff_A_2TFo5LhC0_0),.clk(gclk));
	jdff dff_A_o5jm3Mm81_0(.dout(w_dff_A_meQoZqRp6_0),.din(w_dff_A_o5jm3Mm81_0),.clk(gclk));
	jdff dff_A_meQoZqRp6_0(.dout(w_dff_A_o0Dkscnh8_0),.din(w_dff_A_meQoZqRp6_0),.clk(gclk));
	jdff dff_A_o0Dkscnh8_0(.dout(w_dff_A_FU0qnnH58_0),.din(w_dff_A_o0Dkscnh8_0),.clk(gclk));
	jdff dff_A_FU0qnnH58_0(.dout(w_dff_A_YQCi2RKZ1_0),.din(w_dff_A_FU0qnnH58_0),.clk(gclk));
	jdff dff_A_YQCi2RKZ1_0(.dout(w_dff_A_1Lyz008O0_0),.din(w_dff_A_YQCi2RKZ1_0),.clk(gclk));
	jdff dff_A_1Lyz008O0_0(.dout(w_dff_A_dn3jklqc2_0),.din(w_dff_A_1Lyz008O0_0),.clk(gclk));
	jdff dff_A_dn3jklqc2_0(.dout(w_dff_A_IzrKkmJm6_0),.din(w_dff_A_dn3jklqc2_0),.clk(gclk));
	jdff dff_A_IzrKkmJm6_0(.dout(w_dff_A_RgvbBbXO7_0),.din(w_dff_A_IzrKkmJm6_0),.clk(gclk));
	jdff dff_A_RgvbBbXO7_0(.dout(w_dff_A_d6UYDttH1_0),.din(w_dff_A_RgvbBbXO7_0),.clk(gclk));
	jdff dff_A_d6UYDttH1_0(.dout(w_dff_A_q7kUgwte7_0),.din(w_dff_A_d6UYDttH1_0),.clk(gclk));
	jdff dff_A_q7kUgwte7_0(.dout(w_dff_A_78s6Bmiz5_0),.din(w_dff_A_q7kUgwte7_0),.clk(gclk));
	jdff dff_A_78s6Bmiz5_0(.dout(w_dff_A_XSQYp8zp7_0),.din(w_dff_A_78s6Bmiz5_0),.clk(gclk));
	jdff dff_A_XSQYp8zp7_0(.dout(w_dff_A_XQDd9TfH3_0),.din(w_dff_A_XSQYp8zp7_0),.clk(gclk));
	jdff dff_A_XQDd9TfH3_0(.dout(w_dff_A_ORBJJzze9_0),.din(w_dff_A_XQDd9TfH3_0),.clk(gclk));
	jdff dff_A_ORBJJzze9_0(.dout(w_dff_A_p0KFPyrp9_0),.din(w_dff_A_ORBJJzze9_0),.clk(gclk));
	jdff dff_A_p0KFPyrp9_0(.dout(w_dff_A_2fEjbVbc3_0),.din(w_dff_A_p0KFPyrp9_0),.clk(gclk));
	jdff dff_A_2fEjbVbc3_0(.dout(w_dff_A_klDGG1qC4_0),.din(w_dff_A_2fEjbVbc3_0),.clk(gclk));
	jdff dff_A_klDGG1qC4_0(.dout(w_dff_A_dbikGQN51_0),.din(w_dff_A_klDGG1qC4_0),.clk(gclk));
	jdff dff_A_dbikGQN51_0(.dout(w_dff_A_4JGf5plu9_0),.din(w_dff_A_dbikGQN51_0),.clk(gclk));
	jdff dff_A_4JGf5plu9_0(.dout(w_dff_A_mZS3SlCI8_0),.din(w_dff_A_4JGf5plu9_0),.clk(gclk));
	jdff dff_A_mZS3SlCI8_0(.dout(w_dff_A_w2ewmxbD2_0),.din(w_dff_A_mZS3SlCI8_0),.clk(gclk));
	jdff dff_A_w2ewmxbD2_0(.dout(G358),.din(w_dff_A_w2ewmxbD2_0),.clk(gclk));
	jdff dff_A_aHt6RkCZ8_2(.dout(w_dff_A_9kbngka28_0),.din(w_dff_A_aHt6RkCZ8_2),.clk(gclk));
	jdff dff_A_9kbngka28_0(.dout(w_dff_A_IYTSwjoI4_0),.din(w_dff_A_9kbngka28_0),.clk(gclk));
	jdff dff_A_IYTSwjoI4_0(.dout(w_dff_A_qqrfy9M99_0),.din(w_dff_A_IYTSwjoI4_0),.clk(gclk));
	jdff dff_A_qqrfy9M99_0(.dout(w_dff_A_oaVQbbEI6_0),.din(w_dff_A_qqrfy9M99_0),.clk(gclk));
	jdff dff_A_oaVQbbEI6_0(.dout(w_dff_A_kXgogSIG3_0),.din(w_dff_A_oaVQbbEI6_0),.clk(gclk));
	jdff dff_A_kXgogSIG3_0(.dout(w_dff_A_WNT0POCn7_0),.din(w_dff_A_kXgogSIG3_0),.clk(gclk));
	jdff dff_A_WNT0POCn7_0(.dout(w_dff_A_nqoJYSNL1_0),.din(w_dff_A_WNT0POCn7_0),.clk(gclk));
	jdff dff_A_nqoJYSNL1_0(.dout(w_dff_A_cYsBGSsA7_0),.din(w_dff_A_nqoJYSNL1_0),.clk(gclk));
	jdff dff_A_cYsBGSsA7_0(.dout(w_dff_A_B2x7IUKZ3_0),.din(w_dff_A_cYsBGSsA7_0),.clk(gclk));
	jdff dff_A_B2x7IUKZ3_0(.dout(w_dff_A_8Y6CJ15X6_0),.din(w_dff_A_B2x7IUKZ3_0),.clk(gclk));
	jdff dff_A_8Y6CJ15X6_0(.dout(w_dff_A_dd4MIhLH5_0),.din(w_dff_A_8Y6CJ15X6_0),.clk(gclk));
	jdff dff_A_dd4MIhLH5_0(.dout(w_dff_A_2mCLAEP53_0),.din(w_dff_A_dd4MIhLH5_0),.clk(gclk));
	jdff dff_A_2mCLAEP53_0(.dout(w_dff_A_301Oya3x9_0),.din(w_dff_A_2mCLAEP53_0),.clk(gclk));
	jdff dff_A_301Oya3x9_0(.dout(w_dff_A_l4Z1rTCC8_0),.din(w_dff_A_301Oya3x9_0),.clk(gclk));
	jdff dff_A_l4Z1rTCC8_0(.dout(w_dff_A_0MT9M76Q4_0),.din(w_dff_A_l4Z1rTCC8_0),.clk(gclk));
	jdff dff_A_0MT9M76Q4_0(.dout(w_dff_A_vzCd2yne5_0),.din(w_dff_A_0MT9M76Q4_0),.clk(gclk));
	jdff dff_A_vzCd2yne5_0(.dout(w_dff_A_Md6n8JZm6_0),.din(w_dff_A_vzCd2yne5_0),.clk(gclk));
	jdff dff_A_Md6n8JZm6_0(.dout(w_dff_A_Gzgq586f7_0),.din(w_dff_A_Md6n8JZm6_0),.clk(gclk));
	jdff dff_A_Gzgq586f7_0(.dout(w_dff_A_TSk4U95C5_0),.din(w_dff_A_Gzgq586f7_0),.clk(gclk));
	jdff dff_A_TSk4U95C5_0(.dout(w_dff_A_78grfziF7_0),.din(w_dff_A_TSk4U95C5_0),.clk(gclk));
	jdff dff_A_78grfziF7_0(.dout(w_dff_A_8gwvzG3Y4_0),.din(w_dff_A_78grfziF7_0),.clk(gclk));
	jdff dff_A_8gwvzG3Y4_0(.dout(w_dff_A_gQ4ywcus0_0),.din(w_dff_A_8gwvzG3Y4_0),.clk(gclk));
	jdff dff_A_gQ4ywcus0_0(.dout(w_dff_A_OWR7LLM93_0),.din(w_dff_A_gQ4ywcus0_0),.clk(gclk));
	jdff dff_A_OWR7LLM93_0(.dout(w_dff_A_3yZSjYJI9_0),.din(w_dff_A_OWR7LLM93_0),.clk(gclk));
	jdff dff_A_3yZSjYJI9_0(.dout(w_dff_A_Vf4sBJ6B5_0),.din(w_dff_A_3yZSjYJI9_0),.clk(gclk));
	jdff dff_A_Vf4sBJ6B5_0(.dout(w_dff_A_GiPrHPkG6_0),.din(w_dff_A_Vf4sBJ6B5_0),.clk(gclk));
	jdff dff_A_GiPrHPkG6_0(.dout(G351),.din(w_dff_A_GiPrHPkG6_0),.clk(gclk));
	jdff dff_A_iZwOYoxD1_2(.dout(w_dff_A_nxynkYd86_0),.din(w_dff_A_iZwOYoxD1_2),.clk(gclk));
	jdff dff_A_nxynkYd86_0(.dout(w_dff_A_1Yf1Nag91_0),.din(w_dff_A_nxynkYd86_0),.clk(gclk));
	jdff dff_A_1Yf1Nag91_0(.dout(w_dff_A_L48ZhFEL1_0),.din(w_dff_A_1Yf1Nag91_0),.clk(gclk));
	jdff dff_A_L48ZhFEL1_0(.dout(w_dff_A_V1RyywYX5_0),.din(w_dff_A_L48ZhFEL1_0),.clk(gclk));
	jdff dff_A_V1RyywYX5_0(.dout(w_dff_A_mPPi4LPU7_0),.din(w_dff_A_V1RyywYX5_0),.clk(gclk));
	jdff dff_A_mPPi4LPU7_0(.dout(w_dff_A_r0rYql7X9_0),.din(w_dff_A_mPPi4LPU7_0),.clk(gclk));
	jdff dff_A_r0rYql7X9_0(.dout(w_dff_A_WbN5nSJi3_0),.din(w_dff_A_r0rYql7X9_0),.clk(gclk));
	jdff dff_A_WbN5nSJi3_0(.dout(w_dff_A_AaYTQQIO4_0),.din(w_dff_A_WbN5nSJi3_0),.clk(gclk));
	jdff dff_A_AaYTQQIO4_0(.dout(w_dff_A_di5db3TJ7_0),.din(w_dff_A_AaYTQQIO4_0),.clk(gclk));
	jdff dff_A_di5db3TJ7_0(.dout(w_dff_A_YExiTsD20_0),.din(w_dff_A_di5db3TJ7_0),.clk(gclk));
	jdff dff_A_YExiTsD20_0(.dout(w_dff_A_GNI49PoX8_0),.din(w_dff_A_YExiTsD20_0),.clk(gclk));
	jdff dff_A_GNI49PoX8_0(.dout(w_dff_A_PUvCBNmy8_0),.din(w_dff_A_GNI49PoX8_0),.clk(gclk));
	jdff dff_A_PUvCBNmy8_0(.dout(w_dff_A_e0vPEeNW9_0),.din(w_dff_A_PUvCBNmy8_0),.clk(gclk));
	jdff dff_A_e0vPEeNW9_0(.dout(G372),.din(w_dff_A_e0vPEeNW9_0),.clk(gclk));
	jdff dff_A_UNMIhmVW3_2(.dout(w_dff_A_W573gzgN9_0),.din(w_dff_A_UNMIhmVW3_2),.clk(gclk));
	jdff dff_A_W573gzgN9_0(.dout(w_dff_A_NMw2Zrv26_0),.din(w_dff_A_W573gzgN9_0),.clk(gclk));
	jdff dff_A_NMw2Zrv26_0(.dout(w_dff_A_JjnjHTSU2_0),.din(w_dff_A_NMw2Zrv26_0),.clk(gclk));
	jdff dff_A_JjnjHTSU2_0(.dout(w_dff_A_Xxem4AfI3_0),.din(w_dff_A_JjnjHTSU2_0),.clk(gclk));
	jdff dff_A_Xxem4AfI3_0(.dout(w_dff_A_grmmOweH7_0),.din(w_dff_A_Xxem4AfI3_0),.clk(gclk));
	jdff dff_A_grmmOweH7_0(.dout(w_dff_A_ACA69HnV9_0),.din(w_dff_A_grmmOweH7_0),.clk(gclk));
	jdff dff_A_ACA69HnV9_0(.dout(w_dff_A_wpYTuy680_0),.din(w_dff_A_ACA69HnV9_0),.clk(gclk));
	jdff dff_A_wpYTuy680_0(.dout(w_dff_A_KuWfMyM55_0),.din(w_dff_A_wpYTuy680_0),.clk(gclk));
	jdff dff_A_KuWfMyM55_0(.dout(w_dff_A_ivu8aHFk6_0),.din(w_dff_A_KuWfMyM55_0),.clk(gclk));
	jdff dff_A_ivu8aHFk6_0(.dout(w_dff_A_hAuOoFWj5_0),.din(w_dff_A_ivu8aHFk6_0),.clk(gclk));
	jdff dff_A_hAuOoFWj5_0(.dout(w_dff_A_fr52rNKf2_0),.din(w_dff_A_hAuOoFWj5_0),.clk(gclk));
	jdff dff_A_fr52rNKf2_0(.dout(G369),.din(w_dff_A_fr52rNKf2_0),.clk(gclk));
	jdff dff_A_74kv90FR7_2(.dout(w_dff_A_cjS2pxn31_0),.din(w_dff_A_74kv90FR7_2),.clk(gclk));
	jdff dff_A_cjS2pxn31_0(.dout(w_dff_A_WueOsCzZ7_0),.din(w_dff_A_cjS2pxn31_0),.clk(gclk));
	jdff dff_A_WueOsCzZ7_0(.dout(w_dff_A_oGhCCwGG8_0),.din(w_dff_A_WueOsCzZ7_0),.clk(gclk));
	jdff dff_A_oGhCCwGG8_0(.dout(w_dff_A_OKllOvWW4_0),.din(w_dff_A_oGhCCwGG8_0),.clk(gclk));
	jdff dff_A_OKllOvWW4_0(.dout(w_dff_A_QdQBOA8w3_0),.din(w_dff_A_OKllOvWW4_0),.clk(gclk));
	jdff dff_A_QdQBOA8w3_0(.dout(w_dff_A_Slg7fNet9_0),.din(w_dff_A_QdQBOA8w3_0),.clk(gclk));
	jdff dff_A_Slg7fNet9_0(.dout(w_dff_A_MqE4mDbP7_0),.din(w_dff_A_Slg7fNet9_0),.clk(gclk));
	jdff dff_A_MqE4mDbP7_0(.dout(w_dff_A_kDZ2kY0h4_0),.din(w_dff_A_MqE4mDbP7_0),.clk(gclk));
	jdff dff_A_kDZ2kY0h4_0(.dout(w_dff_A_puLJejtV0_0),.din(w_dff_A_kDZ2kY0h4_0),.clk(gclk));
	jdff dff_A_puLJejtV0_0(.dout(w_dff_A_XdftFSS88_0),.din(w_dff_A_puLJejtV0_0),.clk(gclk));
	jdff dff_A_XdftFSS88_0(.dout(w_dff_A_pcZx37y88_0),.din(w_dff_A_XdftFSS88_0),.clk(gclk));
	jdff dff_A_pcZx37y88_0(.dout(w_dff_A_CwM31BKC3_0),.din(w_dff_A_pcZx37y88_0),.clk(gclk));
	jdff dff_A_CwM31BKC3_0(.dout(w_dff_A_uNfvpnLU7_0),.din(w_dff_A_CwM31BKC3_0),.clk(gclk));
	jdff dff_A_uNfvpnLU7_0(.dout(G399),.din(w_dff_A_uNfvpnLU7_0),.clk(gclk));
	jdff dff_A_oGQbtTGb6_2(.dout(w_dff_A_u4Y6Oiym5_0),.din(w_dff_A_oGQbtTGb6_2),.clk(gclk));
	jdff dff_A_u4Y6Oiym5_0(.dout(w_dff_A_z1roqDWs3_0),.din(w_dff_A_u4Y6Oiym5_0),.clk(gclk));
	jdff dff_A_z1roqDWs3_0(.dout(w_dff_A_qTzjGlMH7_0),.din(w_dff_A_z1roqDWs3_0),.clk(gclk));
	jdff dff_A_qTzjGlMH7_0(.dout(w_dff_A_NfmaXxh35_0),.din(w_dff_A_qTzjGlMH7_0),.clk(gclk));
	jdff dff_A_NfmaXxh35_0(.dout(w_dff_A_TS3mP57A5_0),.din(w_dff_A_NfmaXxh35_0),.clk(gclk));
	jdff dff_A_TS3mP57A5_0(.dout(w_dff_A_Hn3wW3cl6_0),.din(w_dff_A_TS3mP57A5_0),.clk(gclk));
	jdff dff_A_Hn3wW3cl6_0(.dout(w_dff_A_vDJgBnJw7_0),.din(w_dff_A_Hn3wW3cl6_0),.clk(gclk));
	jdff dff_A_vDJgBnJw7_0(.dout(w_dff_A_iBMZlcHm8_0),.din(w_dff_A_vDJgBnJw7_0),.clk(gclk));
	jdff dff_A_iBMZlcHm8_0(.dout(G364),.din(w_dff_A_iBMZlcHm8_0),.clk(gclk));
	jdff dff_A_OMDYSKow2_1(.dout(w_dff_A_CLoWoswO9_0),.din(w_dff_A_OMDYSKow2_1),.clk(gclk));
	jdff dff_A_CLoWoswO9_0(.dout(w_dff_A_1GY6J38V1_0),.din(w_dff_A_CLoWoswO9_0),.clk(gclk));
	jdff dff_A_1GY6J38V1_0(.dout(w_dff_A_UfW6VExg5_0),.din(w_dff_A_1GY6J38V1_0),.clk(gclk));
	jdff dff_A_UfW6VExg5_0(.dout(w_dff_A_ZSKi4e2b8_0),.din(w_dff_A_UfW6VExg5_0),.clk(gclk));
	jdff dff_A_ZSKi4e2b8_0(.dout(w_dff_A_3UYy6rT51_0),.din(w_dff_A_ZSKi4e2b8_0),.clk(gclk));
	jdff dff_A_3UYy6rT51_0(.dout(w_dff_A_qvaVkxqt4_0),.din(w_dff_A_3UYy6rT51_0),.clk(gclk));
	jdff dff_A_qvaVkxqt4_0(.dout(w_dff_A_v1DjgLVT8_0),.din(w_dff_A_qvaVkxqt4_0),.clk(gclk));
	jdff dff_A_v1DjgLVT8_0(.dout(w_dff_A_x0Ej28Hs0_0),.din(w_dff_A_v1DjgLVT8_0),.clk(gclk));
	jdff dff_A_x0Ej28Hs0_0(.dout(w_dff_A_CbRgsCRD0_0),.din(w_dff_A_x0Ej28Hs0_0),.clk(gclk));
	jdff dff_A_CbRgsCRD0_0(.dout(w_dff_A_UjOfFQLK5_0),.din(w_dff_A_CbRgsCRD0_0),.clk(gclk));
	jdff dff_A_UjOfFQLK5_0(.dout(w_dff_A_IB1KoBEj5_0),.din(w_dff_A_UjOfFQLK5_0),.clk(gclk));
	jdff dff_A_IB1KoBEj5_0(.dout(w_dff_A_1fhjShhg7_0),.din(w_dff_A_IB1KoBEj5_0),.clk(gclk));
	jdff dff_A_1fhjShhg7_0(.dout(G396),.din(w_dff_A_1fhjShhg7_0),.clk(gclk));
	jdff dff_A_BIzCn8732_1(.dout(w_dff_A_NnaKXWZx5_0),.din(w_dff_A_BIzCn8732_1),.clk(gclk));
	jdff dff_A_NnaKXWZx5_0(.dout(w_dff_A_KyS9Hjs93_0),.din(w_dff_A_NnaKXWZx5_0),.clk(gclk));
	jdff dff_A_KyS9Hjs93_0(.dout(w_dff_A_0g3CbZTa8_0),.din(w_dff_A_KyS9Hjs93_0),.clk(gclk));
	jdff dff_A_0g3CbZTa8_0(.dout(w_dff_A_1M87rgWm2_0),.din(w_dff_A_0g3CbZTa8_0),.clk(gclk));
	jdff dff_A_1M87rgWm2_0(.dout(w_dff_A_DErI4UT83_0),.din(w_dff_A_1M87rgWm2_0),.clk(gclk));
	jdff dff_A_DErI4UT83_0(.dout(w_dff_A_VTfJQwGE2_0),.din(w_dff_A_DErI4UT83_0),.clk(gclk));
	jdff dff_A_VTfJQwGE2_0(.dout(w_dff_A_t0bPdXfN7_0),.din(w_dff_A_VTfJQwGE2_0),.clk(gclk));
	jdff dff_A_t0bPdXfN7_0(.dout(G384),.din(w_dff_A_t0bPdXfN7_0),.clk(gclk));
	jdff dff_A_a1Iu7cw04_2(.dout(w_dff_A_y1N5lnv53_0),.din(w_dff_A_a1Iu7cw04_2),.clk(gclk));
	jdff dff_A_y1N5lnv53_0(.dout(w_dff_A_dVxtIZAd8_0),.din(w_dff_A_y1N5lnv53_0),.clk(gclk));
	jdff dff_A_dVxtIZAd8_0(.dout(w_dff_A_g97xnSVg6_0),.din(w_dff_A_dVxtIZAd8_0),.clk(gclk));
	jdff dff_A_g97xnSVg6_0(.dout(w_dff_A_C82QFasT6_0),.din(w_dff_A_g97xnSVg6_0),.clk(gclk));
	jdff dff_A_C82QFasT6_0(.dout(w_dff_A_qyQ4axtJ9_0),.din(w_dff_A_C82QFasT6_0),.clk(gclk));
	jdff dff_A_qyQ4axtJ9_0(.dout(w_dff_A_T6L90GSH9_0),.din(w_dff_A_qyQ4axtJ9_0),.clk(gclk));
	jdff dff_A_T6L90GSH9_0(.dout(G367),.din(w_dff_A_T6L90GSH9_0),.clk(gclk));
	jdff dff_A_PSsr8Fhy0_1(.dout(w_dff_A_gudd3lGr8_0),.din(w_dff_A_PSsr8Fhy0_1),.clk(gclk));
	jdff dff_A_gudd3lGr8_0(.dout(w_dff_A_tdXo1ibK4_0),.din(w_dff_A_gudd3lGr8_0),.clk(gclk));
	jdff dff_A_tdXo1ibK4_0(.dout(w_dff_A_wlwNzbXG0_0),.din(w_dff_A_tdXo1ibK4_0),.clk(gclk));
	jdff dff_A_wlwNzbXG0_0(.dout(w_dff_A_2O09XMK62_0),.din(w_dff_A_wlwNzbXG0_0),.clk(gclk));
	jdff dff_A_2O09XMK62_0(.dout(w_dff_A_Gw1BjGpo0_0),.din(w_dff_A_2O09XMK62_0),.clk(gclk));
	jdff dff_A_Gw1BjGpo0_0(.dout(G387),.din(w_dff_A_Gw1BjGpo0_0),.clk(gclk));
	jdff dff_A_6yoiM3mB4_1(.dout(w_dff_A_bHnA99PJ1_0),.din(w_dff_A_6yoiM3mB4_1),.clk(gclk));
	jdff dff_A_bHnA99PJ1_0(.dout(w_dff_A_YTjfZZFu2_0),.din(w_dff_A_bHnA99PJ1_0),.clk(gclk));
	jdff dff_A_YTjfZZFu2_0(.dout(w_dff_A_NVctI2WS2_0),.din(w_dff_A_YTjfZZFu2_0),.clk(gclk));
	jdff dff_A_NVctI2WS2_0(.dout(w_dff_A_oDfHDQeK2_0),.din(w_dff_A_NVctI2WS2_0),.clk(gclk));
	jdff dff_A_oDfHDQeK2_0(.dout(w_dff_A_46DSCL1y5_0),.din(w_dff_A_oDfHDQeK2_0),.clk(gclk));
	jdff dff_A_46DSCL1y5_0(.dout(w_dff_A_jfdPnZ8C5_0),.din(w_dff_A_46DSCL1y5_0),.clk(gclk));
	jdff dff_A_jfdPnZ8C5_0(.dout(G393),.din(w_dff_A_jfdPnZ8C5_0),.clk(gclk));
	jdff dff_A_6xuJbluM3_1(.dout(w_dff_A_DrYpNYYV3_0),.din(w_dff_A_6xuJbluM3_1),.clk(gclk));
	jdff dff_A_DrYpNYYV3_0(.dout(w_dff_A_dmHlHfbC2_0),.din(w_dff_A_DrYpNYYV3_0),.clk(gclk));
	jdff dff_A_dmHlHfbC2_0(.dout(w_dff_A_ayDuw0Rr3_0),.din(w_dff_A_dmHlHfbC2_0),.clk(gclk));
	jdff dff_A_ayDuw0Rr3_0(.dout(w_dff_A_dMyhEWA48_0),.din(w_dff_A_ayDuw0Rr3_0),.clk(gclk));
	jdff dff_A_dMyhEWA48_0(.dout(w_dff_A_XsSApLM01_0),.din(w_dff_A_dMyhEWA48_0),.clk(gclk));
	jdff dff_A_XsSApLM01_0(.dout(G390),.din(w_dff_A_XsSApLM01_0),.clk(gclk));
	jdff dff_A_tByJlnk29_1(.dout(w_dff_A_5eXJgyL09_0),.din(w_dff_A_tByJlnk29_1),.clk(gclk));
	jdff dff_A_5eXJgyL09_0(.dout(w_dff_A_1WDh2ufO5_0),.din(w_dff_A_5eXJgyL09_0),.clk(gclk));
	jdff dff_A_1WDh2ufO5_0(.dout(w_dff_A_arVy5Q4o0_0),.din(w_dff_A_1WDh2ufO5_0),.clk(gclk));
	jdff dff_A_arVy5Q4o0_0(.dout(G378),.din(w_dff_A_arVy5Q4o0_0),.clk(gclk));
	jdff dff_A_F97UfJu59_1(.dout(w_dff_A_yAIUZYfb7_0),.din(w_dff_A_F97UfJu59_1),.clk(gclk));
	jdff dff_A_yAIUZYfb7_0(.dout(w_dff_A_bGBEGjHA2_0),.din(w_dff_A_yAIUZYfb7_0),.clk(gclk));
	jdff dff_A_bGBEGjHA2_0(.dout(w_dff_A_QYZeNjaj8_0),.din(w_dff_A_bGBEGjHA2_0),.clk(gclk));
	jdff dff_A_QYZeNjaj8_0(.dout(G375),.din(w_dff_A_QYZeNjaj8_0),.clk(gclk));
	jdff dff_A_07wqAPrM9_1(.dout(w_dff_A_2L7PwvHK6_0),.din(w_dff_A_07wqAPrM9_1),.clk(gclk));
	jdff dff_A_2L7PwvHK6_0(.dout(w_dff_A_9uTwBV9l3_0),.din(w_dff_A_2L7PwvHK6_0),.clk(gclk));
	jdff dff_A_9uTwBV9l3_0(.dout(w_dff_A_BXTsnPBU4_0),.din(w_dff_A_9uTwBV9l3_0),.clk(gclk));
	jdff dff_A_BXTsnPBU4_0(.dout(G381),.din(w_dff_A_BXTsnPBU4_0),.clk(gclk));
	jdff dff_A_eICaxmaI2_1(.dout(G407),.din(w_dff_A_eICaxmaI2_1),.clk(gclk));
	jdff dff_A_LcUuZJrn4_2(.dout(w_dff_A_OigxRcUw0_0),.din(w_dff_A_LcUuZJrn4_2),.clk(gclk));
	jdff dff_A_OigxRcUw0_0(.dout(G402),.din(w_dff_A_OigxRcUw0_0),.clk(gclk));
endmodule

