/*

c1908:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jcb: 102
	jdff: 813
	jand: 128

Summary:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jcb: 102
	jdff: 813
	jand: 128
*/

module c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n188;
	wire n189;
	wire n190;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n202;
	wire n204;
	wire n205;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n222;
	wire n224;
	wire n225;
	wire n226;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire [2:0] w_G101_0;
	wire [2:0] w_G104_0;
	wire [2:0] w_G107_0;
	wire [2:0] w_G110_0;
	wire [1:0] w_G110_1;
	wire [1:0] w_G113_0;
	wire [2:0] w_G116_0;
	wire [2:0] w_G119_0;
	wire [2:0] w_G122_0;
	wire [1:0] w_G122_1;
	wire [2:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [1:0] w_G128_1;
	wire [1:0] w_G131_0;
	wire [2:0] w_G134_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G140_0;
	wire [2:0] w_G143_0;
	wire [1:0] w_G143_1;
	wire [2:0] w_G146_0;
	wire [2:0] w_G210_0;
	wire [1:0] w_G214_0;
	wire [2:0] w_G217_0;
	wire [1:0] w_G221_0;
	wire [1:0] w_G224_0;
	wire [1:0] w_G227_0;
	wire [2:0] w_G234_0;
	wire [2:0] w_G237_0;
	wire [2:0] w_G469_0;
	wire [1:0] w_G472_0;
	wire [2:0] w_G475_0;
	wire [2:0] w_G478_0;
	wire [2:0] w_G902_0;
	wire [2:0] w_G902_1;
	wire [2:0] w_G902_2;
	wire [2:0] w_G902_3;
	wire [2:0] w_G952_0;
	wire [2:0] w_G953_0;
	wire [2:0] w_G953_1;
	wire [1:0] w_n59_0;
	wire [2:0] w_n60_0;
	wire [2:0] w_n61_0;
	wire [2:0] w_n61_1;
	wire [2:0] w_n61_2;
	wire [2:0] w_n61_3;
	wire [1:0] w_n62_0;
	wire [1:0] w_n67_0;
	wire [1:0] w_n68_0;
	wire [2:0] w_n70_0;
	wire [2:0] w_n70_1;
	wire [2:0] w_n70_2;
	wire [1:0] w_n70_3;
	wire [1:0] w_n71_0;
	wire [1:0] w_n73_0;
	wire [2:0] w_n74_0;
	wire [1:0] w_n74_1;
	wire [1:0] w_n77_0;
	wire [1:0] w_n79_0;
	wire [2:0] w_n81_0;
	wire [1:0] w_n82_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n86_0;
	wire [2:0] w_n90_0;
	wire [2:0] w_n92_0;
	wire [2:0] w_n92_1;
	wire [2:0] w_n93_0;
	wire [1:0] w_n94_0;
	wire [2:0] w_n95_0;
	wire [2:0] w_n96_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [2:0] w_n107_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n109_0;
	wire [2:0] w_n110_0;
	wire [2:0] w_n112_0;
	wire [1:0] w_n112_1;
	wire [2:0] w_n117_0;
	wire [1:0] w_n118_0;
	wire [1:0] w_n119_0;
	wire [1:0] w_n120_0;
	wire [2:0] w_n121_0;
	wire [1:0] w_n121_1;
	wire [1:0] w_n122_0;
	wire [2:0] w_n130_0;
	wire [1:0] w_n131_0;
	wire [2:0] w_n132_0;
	wire [2:0] w_n141_0;
	wire [1:0] w_n142_0;
	wire [2:0] w_n143_0;
	wire [1:0] w_n143_1;
	wire [2:0] w_n144_0;
	wire [2:0] w_n144_1;
	wire [1:0] w_n145_0;
	wire [1:0] w_n146_0;
	wire [1:0] w_n147_0;
	wire [2:0] w_n151_0;
	wire [1:0] w_n152_0;
	wire [2:0] w_n153_0;
	wire [2:0] w_n154_0;
	wire [1:0] w_n154_1;
	wire [2:0] w_n155_0;
	wire [1:0] w_n156_0;
	wire [2:0] w_n158_0;
	wire [1:0] w_n158_1;
	wire [2:0] w_n159_0;
	wire [1:0] w_n159_1;
	wire [1:0] w_n160_0;
	wire [2:0] w_n161_0;
	wire [1:0] w_n162_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n164_0;
	wire [2:0] w_n166_0;
	wire [1:0] w_n166_1;
	wire [1:0] w_n167_0;
	wire [2:0] w_n168_0;
	wire [1:0] w_n169_0;
	wire [1:0] w_n172_0;
	wire [2:0] w_n174_0;
	wire [1:0] w_n174_1;
	wire [1:0] w_n175_0;
	wire [1:0] w_n177_0;
	wire [2:0] w_n179_0;
	wire [1:0] w_n180_0;
	wire [2:0] w_n181_0;
	wire [2:0] w_n183_0;
	wire [2:0] w_n184_0;
	wire [1:0] w_n184_1;
	wire [2:0] w_n185_0;
	wire [1:0] w_n186_0;
	wire [2:0] w_n188_0;
	wire [1:0] w_n189_0;
	wire [1:0] w_n190_0;
	wire [2:0] w_n192_0;
	wire [1:0] w_n193_0;
	wire [2:0] w_n196_0;
	wire [2:0] w_n197_0;
	wire [1:0] w_n197_1;
	wire [2:0] w_n198_0;
	wire [1:0] w_n198_1;
	wire [1:0] w_n199_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n202_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n210_0;
	wire [1:0] w_n212_0;
	wire [1:0] w_n213_0;
	wire [2:0] w_n216_0;
	wire [2:0] w_n217_0;
	wire [2:0] w_n218_0;
	wire [1:0] w_n218_1;
	wire [1:0] w_n219_0;
	wire [1:0] w_n220_0;
	wire [1:0] w_n222_0;
	wire [1:0] w_n226_0;
	wire [1:0] w_n228_0;
	wire [2:0] w_n244_0;
	wire [2:0] w_n244_1;
	wire [2:0] w_n244_2;
	wire [1:0] w_n252_0;
	wire [2:0] w_n253_0;
	wire [2:0] w_n254_0;
	wire [1:0] w_n254_1;
	wire [2:0] w_n273_0;
	wire [1:0] w_n274_0;
	wire [1:0] w_n275_0;
	wire [2:0] w_n276_0;
	wire [1:0] w_n276_1;
	wire [1:0] w_n277_0;
	wire [1:0] w_n278_0;
	wire [1:0] w_n280_0;
	wire [2:0] w_n281_0;
	wire [1:0] w_n282_0;
	wire [1:0] w_n286_0;
	wire [2:0] w_n288_0;
	wire [1:0] w_n289_0;
	wire [2:0] w_n290_0;
	wire [1:0] w_n291_0;
	wire [1:0] w_n295_0;
	wire [1:0] w_n308_0;
	wire [1:0] w_n309_0;
	wire [2:0] w_n311_0;
	wire [2:0] w_n314_0;
	wire [1:0] w_n315_0;
	wire [1:0] w_n318_0;
	wire [1:0] w_n325_0;
	wire [1:0] w_n334_0;
	wire [2:0] w_n335_0;
	wire [2:0] w_n335_1;
	wire [1:0] w_n335_2;
	wire [1:0] w_n336_0;
	wire [2:0] w_n340_0;
	wire [2:0] w_n340_1;
	wire [1:0] w_n340_2;
	wire [1:0] w_n346_0;
	wire [1:0] w_n355_0;
	wire [1:0] w_n364_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n395_0;
	wire w_dff_B_qIklqYuI8_0;
	wire w_dff_B_aMa4dRVW8_0;
	wire w_dff_B_KZlQMPHE0_0;
	wire w_dff_B_UUkHKZoh3_1;
	wire w_dff_B_Ko9Q0Ouk9_0;
	wire w_dff_B_qLE4qJCR1_0;
	wire w_dff_B_DTiGo68Z0_0;
	wire w_dff_B_x3X379eF2_2;
	wire w_dff_B_Leox0wox6_0;
	wire w_dff_B_X5b1YLFJ7_1;
	wire w_dff_B_PbRkO0Ib6_1;
	wire w_dff_B_tZb0ThWF1_1;
	wire w_dff_B_p3Y1KmNo3_1;
	wire w_dff_B_0kPGg72q9_1;
	wire w_dff_B_AIw4y7yr9_1;
	wire w_dff_B_wKrwOjjf4_1;
	wire w_dff_B_4JD1duB90_1;
	wire w_dff_B_XpMiKSVd3_0;
	wire w_dff_B_nPgonPMr5_0;
	wire w_dff_B_8MNJWJOr5_0;
	wire w_dff_B_S46GJT483_0;
	wire w_dff_B_eOBnwvJ22_0;
	wire w_dff_B_L8DhmnAe5_0;
	wire w_dff_B_rVCYKYF15_0;
	wire w_dff_B_P2noYk0w1_0;
	wire w_dff_B_KHL9ZZiS4_0;
	wire w_dff_B_vX93nVos8_0;
	wire w_dff_B_IWsozdop8_0;
	wire w_dff_B_qvJFveWg6_0;
	wire w_dff_A_XiONjEUM2_0;
	wire w_dff_A_YqtWxJyX4_0;
	wire w_dff_A_aTaWS9d60_0;
	wire w_dff_A_mfUZGYf69_0;
	wire w_dff_A_xl8xkgtH0_0;
	wire w_dff_A_fIajYCHH2_0;
	wire w_dff_A_xQK1tryG4_0;
	wire w_dff_A_MMdwnign8_0;
	wire w_dff_A_AvyULZ1F5_0;
	wire w_dff_A_q6qdmp4l7_0;
	wire w_dff_A_4KWj67gY2_0;
	wire w_dff_B_4gSGPn0c7_1;
	wire w_dff_B_PftEIhlQ2_1;
	wire w_dff_B_4cv6HsYs4_1;
	wire w_dff_B_HhksMVJk3_1;
	wire w_dff_B_8HdxeRHo2_1;
	wire w_dff_B_tcwanO0x6_1;
	wire w_dff_B_z6Nu5UI97_1;
	wire w_dff_B_TsqBpAWs7_1;
	wire w_dff_B_h6Hshl8r8_0;
	wire w_dff_B_lnTU46Ef4_0;
	wire w_dff_B_tCzDTeqT0_0;
	wire w_dff_B_YUMKxQk66_0;
	wire w_dff_B_6aPnnOYi4_0;
	wire w_dff_B_iYRoJbsl9_0;
	wire w_dff_B_SOQaeGBi5_0;
	wire w_dff_B_BpIB3ZO56_0;
	wire w_dff_B_QebjCnVd4_0;
	wire w_dff_B_LVGe939C6_0;
	wire w_dff_B_TQD91yn85_0;
	wire w_dff_B_G06qirAy6_0;
	wire w_dff_A_eMp0VwuS4_0;
	wire w_dff_A_geepDOnh4_0;
	wire w_dff_A_B9UNNt9x7_0;
	wire w_dff_A_snupMABS2_0;
	wire w_dff_A_9D0fOy2s0_0;
	wire w_dff_A_m8HZVMo33_0;
	wire w_dff_A_6Y4fJwgq7_0;
	wire w_dff_A_F3YcPR6V1_0;
	wire w_dff_A_VmV5FVrD4_0;
	wire w_dff_A_JUVxXoti1_0;
	wire w_dff_A_PhNOj6iL2_0;
	wire w_dff_B_gzcYmuB61_1;
	wire w_dff_B_395PlfaZ4_1;
	wire w_dff_B_F8Bk1z935_1;
	wire w_dff_B_RR7Uxxnl8_1;
	wire w_dff_B_ZeVdFJOw8_1;
	wire w_dff_B_VX07fHe10_1;
	wire w_dff_B_GfWWVd2B8_1;
	wire w_dff_B_0cRPFybT1_1;
	wire w_dff_B_DTXxkQbj7_0;
	wire w_dff_B_1McTIwJt3_0;
	wire w_dff_B_Jw0Z8M1B9_0;
	wire w_dff_B_Vz6Vlum58_0;
	wire w_dff_B_dINI8ZUP3_0;
	wire w_dff_B_Qivm8uCV2_0;
	wire w_dff_B_eF2q1hLQ7_0;
	wire w_dff_B_TY6vQDrg4_0;
	wire w_dff_B_PhZkkJJa1_0;
	wire w_dff_B_NzZ5V3kN8_0;
	wire w_dff_B_Wjf4zQ7n9_0;
	wire w_dff_B_s2kl1zm84_0;
	wire w_dff_A_bzQR8LFP0_0;
	wire w_dff_A_gc8R2JtK2_0;
	wire w_dff_A_d7zF79lz3_0;
	wire w_dff_A_nQ6aHKOg1_0;
	wire w_dff_A_dm8tWFpL6_0;
	wire w_dff_A_umN1t3SI3_0;
	wire w_dff_A_6Wfwcwbb4_0;
	wire w_dff_A_fxG2Bkiq3_0;
	wire w_dff_A_22BpD5M60_0;
	wire w_dff_A_imeOIfBC3_0;
	wire w_dff_A_Wi2sX6WX9_0;
	wire w_dff_B_0A5AnHRJ6_1;
	wire w_dff_B_IWOnRHmV8_1;
	wire w_dff_B_vd7RZRZQ4_1;
	wire w_dff_B_1teWePyF9_1;
	wire w_dff_B_si90QFER0_1;
	wire w_dff_B_icu8dmV40_1;
	wire w_dff_B_Q4gWqjTo5_1;
	wire w_dff_B_GUcOIG9m7_1;
	wire w_dff_B_evOaY06v4_0;
	wire w_dff_B_KlX3RWNc3_0;
	wire w_dff_B_cW3URVOS0_0;
	wire w_dff_B_tbqvdAG68_0;
	wire w_dff_B_r836DeSm9_0;
	wire w_dff_B_YnFkwijJ8_0;
	wire w_dff_B_23WNmQWq8_0;
	wire w_dff_B_kZOWN7u47_0;
	wire w_dff_B_S7jUhja64_0;
	wire w_dff_B_bubJ0FPE4_0;
	wire w_dff_B_jC8nVPTV4_0;
	wire w_dff_B_iVxIWCT72_0;
	wire w_dff_A_7tlowIyn2_0;
	wire w_dff_A_zHbC0nEr4_0;
	wire w_dff_A_3E0vZNI53_0;
	wire w_dff_A_NkVginFn0_0;
	wire w_dff_A_xkvxwhXk6_0;
	wire w_dff_A_RmdZkWv63_0;
	wire w_dff_A_hooEpd6B0_0;
	wire w_dff_A_VATPqFss2_0;
	wire w_dff_A_CdbqV4wH7_0;
	wire w_dff_A_oB3bxZdb5_0;
	wire w_dff_A_I6BHAfxa8_0;
	wire w_dff_B_zKKZ3OEc9_1;
	wire w_dff_B_MgoIaZ0d6_1;
	wire w_dff_B_rQ3APO7a0_0;
	wire w_dff_B_2Vc9FAdH3_0;
	wire w_dff_B_dIHTQlUc5_0;
	wire w_dff_B_pMAnzE9l5_0;
	wire w_dff_B_ZNW43P2h7_0;
	wire w_dff_B_8dkfrdX51_0;
	wire w_dff_B_wSvcQ8VG9_0;
	wire w_dff_B_n5BItyIC8_0;
	wire w_dff_B_knUKdgrF7_0;
	wire w_dff_B_jTCA9YDL5_0;
	wire w_dff_B_NcuqmW5k8_0;
	wire w_dff_B_2KeNDtYV1_0;
	wire w_dff_A_rHrGhwGm6_0;
	wire w_dff_A_VtiVWISb2_1;
	wire w_dff_A_SjSFDZ172_1;
	wire w_dff_A_HnDKh3SD2_1;
	wire w_dff_A_LVohhpl28_1;
	wire w_dff_A_jotmuWdv7_1;
	wire w_dff_A_NwbRj9zl4_1;
	wire w_dff_A_RkMChSBt7_1;
	wire w_dff_A_aTKAHHWz1_1;
	wire w_dff_A_UxttpmSE7_1;
	wire w_dff_A_b4AgwyJ03_1;
	wire w_dff_A_TL2yhSof4_1;
	wire w_dff_B_X55qSwQ59_1;
	wire w_dff_B_6i9ei40a9_1;
	wire w_dff_B_BE0wj4rv4_1;
	wire w_dff_B_UnDnEvbz5_1;
	wire w_dff_B_65ZOrPmx6_1;
	wire w_dff_B_FQDpFeNo3_1;
	wire w_dff_B_nA4SKkqB7_1;
	wire w_dff_B_DIgbkSqt5_1;
	wire w_dff_B_yLSdhCZv3_1;
	wire w_dff_B_h1QunbAe8_1;
	wire w_dff_B_EtETzIiC2_1;
	wire w_dff_B_3U02k0zt1_1;
	wire w_dff_B_FpHpHvB37_1;
	wire w_dff_B_29L0AqtW3_0;
	wire w_dff_B_f1rGZROM0_0;
	wire w_dff_B_CXPGAOjp9_0;
	wire w_dff_B_x6buodD33_0;
	wire w_dff_B_m7Ig0zAD1_0;
	wire w_dff_B_lOepdcUX9_0;
	wire w_dff_B_czWIJref1_0;
	wire w_dff_B_gcUtwAsh1_0;
	wire w_dff_B_mbzieB0G6_0;
	wire w_dff_B_QZkuKSeL6_0;
	wire w_dff_B_4UcDNbX05_0;
	wire w_dff_B_h3nV6xkx4_0;
	wire w_dff_B_kxufNpK89_0;
	wire w_dff_B_BcqZbD243_0;
	wire w_dff_B_HE0CuCCN0_0;
	wire w_dff_B_gssPliqy2_0;
	wire w_dff_B_J7xJxTDd6_0;
	wire w_dff_B_vzeYRoUh1_0;
	wire w_dff_B_Crwz3Alx7_0;
	wire w_dff_B_WVAZna0S0_0;
	wire w_dff_B_61pLk6yF7_0;
	wire w_dff_B_PdPedVg21_1;
	wire w_dff_B_suVRAECO2_1;
	wire w_dff_B_022ZCcFP7_1;
	wire w_dff_B_dBRpNvDI0_0;
	wire w_dff_B_VVOSGF3B5_0;
	wire w_dff_B_VFhQmT8V3_0;
	wire w_dff_B_Gn09emKO0_0;
	wire w_dff_B_ImpSVUN95_0;
	wire w_dff_B_v0Qnln3h1_0;
	wire w_dff_B_8vxcRGM88_0;
	wire w_dff_B_vSf3deVJ8_0;
	wire w_dff_B_ox8kK8oC3_0;
	wire w_dff_B_OCWgBTbT0_0;
	wire w_dff_B_QcpHiPlY3_0;
	wire w_dff_B_y5Ms6zHM2_0;
	wire w_dff_A_TTLwkGB22_0;
	wire w_dff_A_kenMqaJC9_0;
	wire w_dff_A_o6iHd4wS5_0;
	wire w_dff_A_GfqyIOPq1_0;
	wire w_dff_A_PGts8FVS1_0;
	wire w_dff_A_1wJHQT8i1_2;
	wire w_dff_A_LcBlZ9aX5_2;
	wire w_dff_A_Fa2UMt9f5_2;
	wire w_dff_B_axGrS3Iv1_3;
	wire w_dff_B_nI5fi7wz8_0;
	wire w_dff_A_8rWjRxp07_0;
	wire w_dff_B_dSziAO2Z1_0;
	wire w_dff_A_BNL5dXN84_0;
	wire w_dff_A_prYlLrbr6_2;
	wire w_dff_A_2B8NSCZf5_2;
	wire w_dff_A_Vd29EL2O1_0;
	wire w_dff_A_dA8Bc4bg1_0;
	wire w_dff_B_7SPTAqeQ4_3;
	wire w_dff_A_7t150ZsV1_0;
	wire w_dff_A_1wrvM3uX4_1;
	wire w_dff_A_YONZmBkR0_0;
	wire w_dff_A_zs3zT8BU7_2;
	wire w_dff_A_8YxqbqHk9_0;
	wire w_dff_A_3qPQklFW8_1;
	wire w_dff_A_3cSJ8hMY5_2;
	wire w_dff_A_pod2XMWh3_2;
	wire w_dff_A_STNXeMv85_1;
	wire w_dff_A_QYAUMjpJ2_1;
	wire w_dff_A_G1aJbt6l0_1;
	wire w_dff_A_WtZesN640_1;
	wire w_dff_A_e2uwbNNi9_1;
	wire w_dff_A_3PBly9OT4_2;
	wire w_dff_A_SKE5l9Sv3_2;
	wire w_dff_A_P22dRqlb4_2;
	wire w_dff_A_5Xc59Xal7_2;
	wire w_dff_A_HQSc0RKe9_2;
	wire w_dff_B_o5OKE4Qy5_3;
	wire w_dff_B_cNBx2DoW7_3;
	wire w_dff_B_YudUmxXw9_3;
	wire w_dff_B_Fb0mb4rz9_3;
	wire w_dff_B_IQIZtJwg9_3;
	wire w_dff_B_cT0aTmBS3_3;
	wire w_dff_B_H5glYabS3_3;
	wire w_dff_B_gIQ4yZ628_3;
	wire w_dff_B_ijbgwGBd3_3;
	wire w_dff_B_hmP7Xgvq0_3;
	wire w_dff_B_SAdMQ8W21_3;
	wire w_dff_B_mOt15Rct5_3;
	wire w_dff_B_yh0Ff1q94_1;
	wire w_dff_B_tEU1EZhI4_1;
	wire w_dff_B_uQkA5nfM7_1;
	wire w_dff_B_TsgPsMYj5_1;
	wire w_dff_B_msmgJLvC1_1;
	wire w_dff_B_c6CCa8PK5_1;
	wire w_dff_B_dqsrEPo56_1;
	wire w_dff_B_Czv2JzUB9_1;
	wire w_dff_B_sqnk2SLN1_0;
	wire w_dff_B_Rzr8Ywb19_0;
	wire w_dff_B_DxmhlZKD5_0;
	wire w_dff_B_ODSuntNp6_0;
	wire w_dff_B_SBkrtyXU0_0;
	wire w_dff_B_onb1ImyF2_0;
	wire w_dff_B_a6crvk4w2_0;
	wire w_dff_B_pNSd7VtP8_0;
	wire w_dff_B_kR6XVgw99_0;
	wire w_dff_B_k8RBcNYk9_0;
	wire w_dff_B_fA13W3LH0_0;
	wire w_dff_B_AjK9z4Zd6_0;
	wire w_dff_A_QW8XngQV8_0;
	wire w_dff_A_lMNyvMra4_0;
	wire w_dff_A_z1un55ZR9_0;
	wire w_dff_A_ENPr6b0i8_0;
	wire w_dff_A_o4kweXGV0_0;
	wire w_dff_A_5pDU0vH70_0;
	wire w_dff_A_3bvbr5rV8_0;
	wire w_dff_A_gGaJ42v52_0;
	wire w_dff_A_y7tY9tcx0_0;
	wire w_dff_A_s8mRo0vA3_0;
	wire w_dff_A_CTbbxFKx9_0;
	wire w_dff_B_4Ceh4tJ99_0;
	wire w_dff_B_UCJLGiV16_0;
	wire w_dff_B_SoUsOi0K6_0;
	wire w_dff_B_dRAP4BFq1_0;
	wire w_dff_B_u1v0oDzC5_0;
	wire w_dff_A_Co56wZdW7_1;
	wire w_dff_B_syV6dGNo7_1;
	wire w_dff_A_1OKfejET8_1;
	wire w_dff_A_KJgL8d3N4_2;
	wire w_dff_A_0Epgjh5R4_2;
	wire w_dff_B_9C0m26qy5_3;
	wire w_dff_B_01Sj3U7Z8_3;
	wire w_dff_B_KxqXcm3f6_1;
	wire w_dff_A_ytS0m6ve3_0;
	wire w_dff_A_1QG9NFcn5_2;
	wire w_dff_B_YxBQv0KS6_3;
	wire w_dff_A_WliHaTzo1_1;
	wire w_dff_B_Hc8yxGjE5_3;
	wire w_dff_A_AYIUsmw50_0;
	wire w_dff_A_3t72QqKb7_0;
	wire w_dff_A_inl9Q56b6_1;
	wire w_dff_A_vPrrgWUx2_1;
	wire w_dff_B_xaq43RIw5_0;
	wire w_dff_B_acby1dGc9_0;
	wire w_dff_B_jMQCyKhi9_0;
	wire w_dff_B_vdJpMGfu1_1;
	wire w_dff_A_fQQWn7ir4_0;
	wire w_dff_A_GFsw4uTu9_0;
	wire w_dff_B_IzJsr9a93_1;
	wire w_dff_B_Jkj5CeEG9_0;
	wire w_dff_B_AypWXcsc5_0;
	wire w_dff_B_nlL1oXQa2_0;
	wire w_dff_A_wPCGl1qU9_1;
	wire w_dff_B_xmAMFAiU6_0;
	wire w_dff_A_0TVHd13F1_0;
	wire w_dff_B_ElRGm0qY9_2;
	wire w_dff_A_FApMqmB96_2;
	wire w_dff_B_HhfOLex49_3;
	wire w_dff_A_F5N597V85_0;
	wire w_dff_A_oIpNTQ8z8_0;
	wire w_dff_A_KQ9LXcof3_1;
	wire w_dff_A_BbZgDHH93_0;
	wire w_dff_A_S0id8zff3_0;
	wire w_dff_A_c9ksjVia9_2;
	wire w_dff_A_psk5xJCz6_1;
	wire w_dff_A_JH53DPRX5_2;
	wire w_dff_B_9jxaQbhS9_1;
	wire w_dff_B_qhZi3BqZ7_1;
	wire w_dff_B_2nYgILi63_1;
	wire w_dff_B_WPWpcJ4S9_1;
	wire w_dff_B_N9MFRpiV9_1;
	wire w_dff_B_opegiqZu4_0;
	wire w_dff_B_ESBooY621_0;
	wire w_dff_A_E9HyUkut8_0;
	wire w_dff_A_EnfNjDbK7_0;
	wire w_dff_A_lqMR1kOK2_0;
	wire w_dff_A_yLpA6jkf7_0;
	wire w_dff_A_xqBNKJBb9_0;
	wire w_dff_A_EkgqexoQ7_0;
	wire w_dff_A_Fc7Heav51_0;
	wire w_dff_A_clZThNqh3_1;
	wire w_dff_B_U6R6kNON7_3;
	wire w_dff_A_xLqE1JzG5_1;
	wire w_dff_A_9ptEOAnV7_2;
	wire w_dff_B_dEIbBMUA1_1;
	wire w_dff_B_wGZVrejg7_1;
	wire w_dff_B_DSYPtOPP9_1;
	wire w_dff_B_oRFGlCql2_1;
	wire w_dff_B_rSVmiRJ22_1;
	wire w_dff_A_ihBmT6X81_0;
	wire w_dff_A_6RqHY63b9_0;
	wire w_dff_A_3caWganY0_0;
	wire w_dff_A_GEDPlgqP4_0;
	wire w_dff_A_TZAWdQve4_0;
	wire w_dff_A_U9qEaIsr8_0;
	wire w_dff_A_qQswp3Rc4_0;
	wire w_dff_A_1WZ6LAoB7_0;
	wire w_dff_B_qSEcbz4e4_1;
	wire w_dff_B_NZNl7SDx2_1;
	wire w_dff_B_2iYyE76X8_0;
	wire w_dff_A_YtbwLOvK1_1;
	wire w_dff_A_fqFOCZqU4_1;
	wire w_dff_A_iSz2xtx77_1;
	wire w_dff_A_9cDS0aSX6_1;
	wire w_dff_A_dFfHpZLB9_1;
	wire w_dff_A_a4VxBFAt6_1;
	wire w_dff_A_eHwbqypz2_0;
	wire w_dff_A_lbJ74lRp3_0;
	wire w_dff_A_xy84moId2_0;
	wire w_dff_A_c4AWVLou1_0;
	wire w_dff_A_ZMRlQDSQ9_0;
	wire w_dff_A_7x47ZWu61_0;
	wire w_dff_A_Ub33pQGe3_0;
	wire w_dff_A_YhyKNndE6_0;
	wire w_dff_B_hOZClFAs5_1;
	wire w_dff_B_SM4MwVuM7_1;
	wire w_dff_B_m6YuB7hj4_1;
	wire w_dff_B_I98vDFqU9_0;
	wire w_dff_A_2n2Yxywx8_1;
	wire w_dff_A_y8KKYUSx4_1;
	wire w_dff_A_R6Id4wSI8_1;
	wire w_dff_A_X96W8BW71_1;
	wire w_dff_A_mqmHQGXz3_1;
	wire w_dff_A_3qplDVlv4_1;
	wire w_dff_B_MrzhAbhq1_3;
	wire w_dff_B_fNgSMBRA9_3;
	wire w_dff_A_9QmyvYKP1_0;
	wire w_dff_A_S4xbV8Hs5_0;
	wire w_dff_A_okHa4Bzi7_1;
	wire w_dff_A_Ro2hpgkn1_1;
	wire w_dff_B_4mOGeCqi9_1;
	wire w_dff_B_qE8bWmkO5_1;
	wire w_dff_B_YR1gWoKv7_1;
	wire w_dff_A_iIfVa4Dt5_1;
	wire w_dff_A_0XuJysZd7_1;
	wire w_dff_A_Dylii5uV1_1;
	wire w_dff_A_dJZKeeg89_1;
	wire w_dff_A_jkYG3eLP8_1;
	wire w_dff_A_Sgcd4f6U3_1;
	wire w_dff_A_n5qQQkyW4_1;
	wire w_dff_A_D7oeaaDe2_1;
	wire w_dff_A_cgWO6s0e3_1;
	wire w_dff_A_TqnVoeS69_1;
	wire w_dff_A_wcUY13iH0_1;
	wire w_dff_A_kSzVm8uM8_1;
	wire w_dff_A_ukeACLI76_1;
	wire w_dff_A_yB2Frsr14_1;
	wire w_dff_A_I0rpjgeH9_1;
	wire w_dff_A_Pigc28xR3_1;
	wire w_dff_A_7kAo5nXh7_1;
	wire w_dff_A_dg4Yy4wf7_1;
	wire w_dff_A_sfXzP4f65_1;
	wire w_dff_B_fdscj1JI9_3;
	wire w_dff_B_JPJZpma22_1;
	wire w_dff_B_CwepJYR72_2;
	wire w_dff_A_vYcfVLIy1_1;
	wire w_dff_A_zqYekie86_2;
	wire w_dff_A_gjC2y7aA7_2;
	wire w_dff_A_CqgGQlX77_1;
	wire w_dff_A_4PhKBgEt9_1;
	wire w_dff_A_XoSdplwf8_1;
	wire w_dff_A_vQqJWAqS3_1;
	wire w_dff_A_jSMj55om2_1;
	wire w_dff_A_PiOiHVkx0_1;
	wire w_dff_A_zI8VUVET9_0;
	wire w_dff_B_qg1uBTWy8_2;
	wire w_dff_B_RgNxSbqc4_2;
	wire w_dff_B_OPpNW5H85_2;
	wire w_dff_A_kaVXNc8z2_1;
	wire w_dff_A_VehClCCv1_1;
	wire w_dff_A_pMkwi8aY5_2;
	wire w_dff_A_lvYd21NF1_2;
	wire w_dff_A_MOEusTo60_2;
	wire w_dff_A_Imz1djx30_0;
	wire w_dff_A_sOHgbdgu6_0;
	wire w_dff_A_nPdhDemH2_0;
	wire w_dff_A_FeuGXCMF4_0;
	wire w_dff_A_wiDoK8v92_0;
	wire w_dff_A_FnkGLtEb5_0;
	wire w_dff_B_HLA88eNZ3_1;
	wire w_dff_B_1y5pYWzk4_1;
	wire w_dff_B_WHlG6HFB2_1;
	wire w_dff_B_VVnMqQBO2_0;
	wire w_dff_B_qzwN81lV1_0;
	wire w_dff_B_iJOcSZc75_0;
	wire w_dff_A_X1VyPlIh4_2;
	wire w_dff_A_Q0YPYRrC2_2;
	wire w_dff_A_ImAltbNP0_2;
	wire w_dff_A_9Q4mYpeZ7_2;
	wire w_dff_A_WAdGVKVL0_0;
	wire w_dff_A_kwNRHKi92_0;
	wire w_dff_A_oD3XMy220_0;
	wire w_dff_A_DsDVFYKP5_0;
	wire w_dff_A_IacUM4se0_0;
	wire w_dff_A_Q0UtPfUY9_0;
	wire w_dff_A_WTPZk5ac1_0;
	wire w_dff_A_G9Z0dt8A8_0;
	wire w_dff_A_4Pgu4pSc6_0;
	wire w_dff_A_dj1IMBKV3_2;
	wire w_dff_A_cWvGkUWR9_2;
	wire w_dff_A_001YZGUH6_2;
	wire w_dff_A_1Clx8xz59_2;
	wire w_dff_A_CN1DHKJk6_1;
	wire w_dff_A_uMjKPJT36_2;
	wire w_dff_B_bhRoY6r93_3;
	wire w_dff_B_wPr0VNwI5_1;
	wire w_dff_B_E6QzsEVb9_1;
	wire w_dff_B_gK1ELPSS8_1;
	wire w_dff_B_z2HNY8DT5_1;
	wire w_dff_B_b35UPb6X8_1;
	wire w_dff_A_SAYqYeAA6_0;
	wire w_dff_A_PSWQlojB4_0;
	wire w_dff_A_HW16vTXj7_0;
	wire w_dff_A_I7WEYVly6_0;
	wire w_dff_A_9B813XqM8_0;
	wire w_dff_A_B3Rzr5Ie7_0;
	wire w_dff_A_6dDmuJIW0_0;
	wire w_dff_A_PHCmtKUe5_0;
	wire w_dff_B_occ79nkz0_1;
	wire w_dff_B_XF7aPHFI7_1;
	wire w_dff_B_XwWUbyaA9_2;
	wire w_dff_A_2Pwe5xD42_0;
	wire w_dff_A_ob64nq451_0;
	wire w_dff_A_dIDDNrYK9_0;
	wire w_dff_A_G7RP05tB1_0;
	wire w_dff_A_s7KsCvYc6_0;
	wire w_dff_A_Pm5qag2M2_0;
	wire w_dff_A_D9thSa8h3_0;
	wire w_dff_A_c0MtNqIm1_0;
	wire w_dff_A_vIZevEEt4_0;
	wire w_dff_A_wig9lR7E1_0;
	wire w_dff_A_NaXfPu0L9_0;
	wire w_dff_A_1T56NcLb3_0;
	wire w_dff_A_CmI19uGM8_2;
	wire w_dff_A_UKa6iSEb7_2;
	wire w_dff_A_GL32B1qB5_2;
	wire w_dff_A_V9o54ueu7_2;
	wire w_dff_A_hABQ7jQC6_2;
	wire w_dff_A_wRghbfZ99_2;
	wire w_dff_B_R5NvZTUM2_2;
	wire w_dff_B_ZtOJtenl6_2;
	wire w_dff_B_mjWg5OmM2_2;
	wire w_dff_B_iXVu6Lhd7_2;
	wire w_dff_A_kLuhzMdc3_0;
	wire w_dff_A_gnm3weAu1_0;
	wire w_dff_A_hR1qtTLz2_0;
	wire w_dff_A_YXptWKBs5_0;
	wire w_dff_A_vi6JzD1y3_0;
	wire w_dff_B_nwK763Rc6_1;
	wire w_dff_A_fW8uNh8t5_0;
	wire w_dff_A_ulwh2wrP4_0;
	wire w_dff_A_e1f2Foyk0_0;
	wire w_dff_A_4wBYh1qH1_0;
	wire w_dff_A_gsFWYLBg9_1;
	wire w_dff_A_El32Yq4F9_2;
	wire w_dff_A_BVXrdtrh1_1;
	wire w_dff_A_epkGa6cy4_1;
	wire w_dff_A_71NluWUL3_1;
	wire w_dff_B_5iqB7ot68_1;
	wire w_dff_B_HwDtq9ba8_1;
	wire w_dff_B_jNMOTHPc9_1;
	wire w_dff_B_PFrBXyXU6_1;
	wire w_dff_A_YzWqgtEM3_0;
	wire w_dff_A_OmQqO8tT0_0;
	wire w_dff_A_AjiuBpna8_0;
	wire w_dff_A_Nid2gwQV2_0;
	wire w_dff_A_WBaCJjy50_0;
	wire w_dff_A_TMVH4ehc8_0;
	wire w_dff_A_J7D7C9zu3_0;
	wire w_dff_A_A4XgrKl65_0;
	wire w_dff_B_SLrfBU200_1;
	wire w_dff_A_kOlMzfbA4_0;
	wire w_dff_A_VqhBz2OE9_0;
	wire w_dff_A_bDnFGNFv6_0;
	wire w_dff_A_ztGTFqxF8_0;
	wire w_dff_A_rwGRa3Gc2_0;
	wire w_dff_A_4yRaVz2j3_0;
	wire w_dff_A_Ofm4sO5M1_0;
	wire w_dff_A_ZCPcl85m3_0;
	wire w_dff_A_VNRUGPVX2_0;
	wire w_dff_A_EmibUZNn8_0;
	wire w_dff_A_ZN1uhVPD6_0;
	wire w_dff_A_TZgUmoyB5_0;
	wire w_dff_A_oqaEsJhU9_1;
	wire w_dff_A_7RDDJqxm0_1;
	wire w_dff_B_j8NchfuQ0_2;
	wire w_dff_A_acQ6BEHC1_0;
	wire w_dff_A_B4KoY9132_0;
	wire w_dff_A_7GwyrfkY4_0;
	wire w_dff_A_U9yKmZmb1_0;
	wire w_dff_A_xzGsgmxU6_0;
	wire w_dff_A_YDczaK3y5_0;
	wire w_dff_A_BrdlmCpc2_0;
	wire w_dff_A_ALXZVDQY9_0;
	wire w_dff_A_KazlaGO74_0;
	wire w_dff_A_8dtt8jhM9_0;
	wire w_dff_B_xd96ETnW8_1;
	wire w_dff_A_JlWKuqRR8_0;
	wire w_dff_A_eHbWDQ225_0;
	wire w_dff_A_derTroX22_0;
	wire w_dff_A_EWZZk98l8_0;
	wire w_dff_A_XxAhpcdm3_0;
	wire w_dff_A_BgBLwZxo2_0;
	wire w_dff_A_dLiz0d3b6_0;
	wire w_dff_A_3En41kxw5_0;
	wire w_dff_A_4O1YrcTA3_0;
	wire w_dff_A_gHPRsLIL2_0;
	wire w_dff_A_XFy2QIpz0_0;
	wire w_dff_A_GJISJ8Pl9_0;
	wire w_dff_A_GC5GjNp01_0;
	wire w_dff_A_P1HxWyZA5_0;
	wire w_dff_A_qVYgheDy9_0;
	wire w_dff_A_5TNbuzRu1_0;
	wire w_dff_A_3FDNVewa7_0;
	wire w_dff_A_6kPDtOT71_0;
	wire w_dff_A_yjAX5vwI9_0;
	wire w_dff_A_W6H8pUiF4_0;
	wire w_dff_A_yHUWdIBR4_0;
	wire w_dff_A_3LXgP0c93_0;
	wire w_dff_A_jwEtlGrS2_1;
	wire w_dff_A_zNv4tfBu4_1;
	wire w_dff_A_9DdSNxao3_1;
	wire w_dff_A_2GK19s0i0_1;
	wire w_dff_A_z650O9AP3_1;
	wire w_dff_A_UIemolCt2_1;
	wire w_dff_A_F7YPdviM6_1;
	wire w_dff_A_iIVvANJ47_1;
	wire w_dff_A_K4wuwk3z8_1;
	wire w_dff_A_EzXFpg7j1_1;
	wire w_dff_A_GSjoSRex1_1;
	wire w_dff_A_BTA3jP3j7_1;
	wire w_dff_A_9hMkmGVH8_1;
	wire w_dff_A_XdZ53zG34_1;
	wire w_dff_A_ny2tcttW0_2;
	wire w_dff_A_ABcTzrzq6_1;
	wire w_dff_A_WVPUjYEs2_1;
	wire w_dff_A_yy4fQQUe6_1;
	wire w_dff_A_J15qkT5W3_1;
	wire w_dff_A_4oX8d2lL8_1;
	wire w_dff_A_zcGxgUb23_1;
	wire w_dff_A_vtlyfzYp8_1;
	wire w_dff_A_75rzG71e3_1;
	wire w_dff_A_IwoBo1on5_1;
	wire w_dff_A_iFccukDN9_1;
	wire w_dff_A_EGB9BWmx9_1;
	wire w_dff_A_dRvqBBIl1_1;
	wire w_dff_A_XBzWfh0L6_1;
	wire w_dff_A_rrns76VM5_1;
	wire w_dff_A_EpIsYTrm1_1;
	wire w_dff_A_MZFvmqbH6_1;
	wire w_dff_A_6Y0SRe8A8_1;
	wire w_dff_A_TYclLP6L4_1;
	wire w_dff_A_QMLcamct7_1;
	wire w_dff_A_cRoJLPQA3_1;
	wire w_dff_A_JXaWVVBu4_1;
	wire w_dff_A_XNAk2NZk7_1;
	wire w_dff_A_3kGUtjRt9_1;
	wire w_dff_A_rV874PmD9_1;
	wire w_dff_A_xZ7tDhxY8_1;
	wire w_dff_A_VN6hA1Nm1_1;
	wire w_dff_A_8wjsgzGh7_0;
	wire w_dff_A_lcM2ykDn8_0;
	wire w_dff_A_8166cvVF4_0;
	wire w_dff_A_PvPANHgX4_0;
	wire w_dff_A_vvtOcw8v3_0;
	wire w_dff_A_4sr6rX5J6_0;
	wire w_dff_A_6kKjIGKo4_1;
	wire w_dff_A_dpZiBVzy7_1;
	wire w_dff_A_DQ7uY5mP0_1;
	wire w_dff_A_wjDOrDyr6_1;
	wire w_dff_A_sFH2u8nm8_1;
	wire w_dff_A_yUMrUTrr4_1;
	wire w_dff_A_HhxTUasi1_2;
	wire w_dff_A_ZD40DTeX6_2;
	wire w_dff_A_xkE8FqOR1_2;
	wire w_dff_A_xFZzRMFV9_2;
	wire w_dff_A_XV0vLJNQ4_2;
	wire w_dff_A_9cQh8x9l0_2;
	wire w_dff_A_oa6Wi5jE0_2;
	wire w_dff_A_Xr5gq0lD3_0;
	wire w_dff_A_H0g2eFmb7_0;
	wire w_dff_A_jc4OPAdb0_0;
	wire w_dff_A_op7mq9RO8_0;
	wire w_dff_A_drDN8AOp0_0;
	wire w_dff_A_mtDt0H3R5_0;
	wire w_dff_A_SAgvGc9c8_0;
	wire w_dff_A_xEf78y8R0_0;
	wire w_dff_B_pbx0NWAq9_0;
	wire w_dff_B_2dX0KMoU9_2;
	wire w_dff_A_rN4PWyHm5_0;
	wire w_dff_A_eZ42Bc6Y4_0;
	wire w_dff_A_S1QrIG7Q1_0;
	wire w_dff_A_NLhFgFi00_0;
	wire w_dff_A_YvTB9ISE9_0;
	wire w_dff_A_YJnwZ44V1_0;
	wire w_dff_A_FwqwMjRY3_0;
	wire w_dff_A_OjNuXhHU0_0;
	wire w_dff_A_NQ4qOvEp7_0;
	wire w_dff_A_EHVgwXFq4_0;
	wire w_dff_A_jKJOKbtK3_0;
	wire w_dff_A_IGaND4c64_1;
	wire w_dff_A_714Enl0P3_1;
	wire w_dff_A_wNfGWoYm2_1;
	wire w_dff_A_iVbfdqdV1_1;
	wire w_dff_A_aInKHHQv8_1;
	wire w_dff_A_eVyqfnfQ6_1;
	wire w_dff_A_P4RmtLTS0_1;
	wire w_dff_A_zAQi7Tox5_1;
	wire w_dff_A_1N14BGgV1_1;
	wire w_dff_A_ZwgU9lFw0_1;
	wire w_dff_A_WfePsrL82_1;
	wire w_dff_A_fHj8Qlmy9_1;
	wire w_dff_A_O2HRP7rs9_1;
	wire w_dff_A_Gm5PiSKX9_2;
	wire w_dff_A_mn6ZkUyT0_2;
	wire w_dff_A_tbhiNONq6_2;
	wire w_dff_A_B3td6LzI6_2;
	wire w_dff_A_tLjjikdm6_2;
	wire w_dff_A_V3aEJJsO6_2;
	wire w_dff_A_toKElB6Y4_2;
	wire w_dff_A_RPDo84dn2_2;
	wire w_dff_A_4yWKP1v25_2;
	wire w_dff_A_EMIIOYeM7_2;
	wire w_dff_A_BJKAFMm76_2;
	wire w_dff_A_gX385W5s1_2;
	wire w_dff_A_ddUKeo2G2_2;
	wire w_dff_A_ylYDucCB8_0;
	wire w_dff_A_EKld3pcg0_0;
	wire w_dff_A_q0nHAXmV4_0;
	wire w_dff_A_AmEHrhQV6_0;
	wire w_dff_A_VqRIrjjA9_0;
	wire w_dff_A_GwJqMgDY6_0;
	wire w_dff_A_EMfXk32e9_0;
	wire w_dff_A_tumOYY1B4_0;
	wire w_dff_A_F4JAuFmx3_0;
	wire w_dff_A_SPqektBu0_0;
	wire w_dff_B_IWk5oVRb7_3;
	wire w_dff_A_qveKPsB94_0;
	wire w_dff_A_vL4OBC3h5_0;
	wire w_dff_A_Y3muUcoT4_0;
	wire w_dff_A_x2Bd3gdv0_0;
	wire w_dff_A_AgN90Q0G7_0;
	wire w_dff_A_LMaFAXdJ1_0;
	wire w_dff_A_0QVct4Pr0_0;
	wire w_dff_A_nWq8BmDO8_0;
	wire w_dff_A_rBOdxVvI0_0;
	wire w_dff_A_QRMLf8KU3_0;
	wire w_dff_A_lrpOe7On2_0;
	wire w_dff_A_wOPgZHQT5_0;
	wire w_dff_A_pGIcC5Nb1_0;
	wire w_dff_A_9Dj2fXD11_0;
	wire w_dff_A_MWREZoIe4_0;
	wire w_dff_A_xhKX1fZa1_0;
	wire w_dff_A_5ZpvOOzI4_0;
	wire w_dff_A_0F0hN5Xy2_0;
	wire w_dff_A_Nck09PbR6_0;
	wire w_dff_A_Q0GO04VI3_0;
	wire w_dff_A_XfJSyxlP7_0;
	wire w_dff_A_Xx0hi9WI9_0;
	wire w_dff_A_tyrBzHzI7_0;
	wire w_dff_A_LJf4yOhf3_0;
	wire w_dff_A_CSNq7BSX8_0;
	wire w_dff_A_QsWjfle73_0;
	wire w_dff_A_7JFzegV06_0;
	wire w_dff_A_EisgLbwD9_0;
	wire w_dff_A_dkxi518c3_0;
	wire w_dff_A_AmCo4Aej2_0;
	wire w_dff_A_W1qqONbB1_0;
	wire w_dff_A_q1A0qZEl3_0;
	wire w_dff_A_OutWcRG95_0;
	wire w_dff_A_Vz1GAtqw7_0;
	wire w_dff_B_5VKQOKOj0_1;
	wire w_dff_A_tla3SoKu1_0;
	wire w_dff_A_wKtR7sIw7_0;
	wire w_dff_A_PQ10YjKH9_0;
	wire w_dff_A_lGmpFOEn6_0;
	wire w_dff_A_xEvKF5tx7_0;
	wire w_dff_A_ocggoty87_0;
	wire w_dff_A_uAEfHOzT4_0;
	wire w_dff_A_gS0TxkNc8_0;
	wire w_dff_A_rtLv1IwE6_0;
	wire w_dff_A_U7aYvUsJ2_0;
	wire w_dff_A_y2O5yMa80_0;
	wire w_dff_A_IqzNrTTb5_0;
	wire w_dff_A_uNgtkKv92_1;
	wire w_dff_A_WZhKdfIf8_1;
	wire w_dff_A_FG0UcSXU9_1;
	wire w_dff_A_hGLNjpR19_1;
	wire w_dff_A_LeXS26RJ4_1;
	wire w_dff_A_HDM9xbZg1_1;
	wire w_dff_A_ThyI4IAu2_1;
	wire w_dff_A_leaLF7tD6_1;
	wire w_dff_A_Ung9iAtf2_1;
	wire w_dff_A_bE9whqp88_1;
	wire w_dff_A_McHXRgtX7_1;
	wire w_dff_A_P79p6jqT7_2;
	wire w_dff_A_JRAGx0Nq6_0;
	wire w_dff_A_ff2iXvSU5_1;
	wire w_dff_A_XazWRSaf1_1;
	wire w_dff_A_DzTql2697_1;
	wire w_dff_A_mFRkDpYh1_1;
	wire w_dff_A_5JyVBdS30_1;
	wire w_dff_A_FgbG6MNU9_1;
	wire w_dff_A_abkQUR1R5_1;
	wire w_dff_A_zbqQPR770_1;
	wire w_dff_A_PrTlXV8E9_1;
	wire w_dff_A_xYyJJ0060_1;
	wire w_dff_A_MwfhDWU89_1;
	wire w_dff_A_Ieji7Bl78_1;
	wire w_dff_A_B1IMyYbE1_1;
	wire w_dff_A_VGCYIe8S6_0;
	wire w_dff_A_ZvLVeX474_0;
	wire w_dff_A_s0APKqXo3_0;
	wire w_dff_A_3GO2tmR13_0;
	wire w_dff_A_imf2LaAW7_0;
	wire w_dff_A_hdFgw2bm0_0;
	wire w_dff_A_wiZeESvy6_0;
	wire w_dff_A_LStv0DhR0_0;
	wire w_dff_A_LL4W1OTT3_0;
	wire w_dff_A_uCchKFyL9_0;
	wire w_dff_A_NvTiZtab6_0;
	wire w_dff_A_3hDjbJ9a1_0;
	wire w_dff_A_zgTcLVob3_0;
	wire w_dff_A_RS764XpV0_0;
	wire w_dff_A_s1PP3tVz0_0;
	wire w_dff_A_h1DWEH6k2_0;
	wire w_dff_A_xyaU7Rad7_0;
	wire w_dff_A_k3ndl7Y64_0;
	wire w_dff_A_tb5KwVXj3_0;
	wire w_dff_A_XvgoQNPf8_0;
	wire w_dff_A_5iRqOBHK5_0;
	wire w_dff_A_VfRoeoli6_0;
	wire w_dff_A_FNCOujbh5_2;
	wire w_dff_A_seMvB0Zz0_2;
	wire w_dff_B_Yb2Y004C3_3;
	wire w_dff_A_WPSsL5Ei1_0;
	wire w_dff_A_5OzUNPNt7_0;
	wire w_dff_A_q6HbcHHl6_0;
	wire w_dff_A_xKJatb3f9_0;
	wire w_dff_A_OFPz05A60_0;
	wire w_dff_A_60LGZOKg3_0;
	wire w_dff_A_Y07P36u01_0;
	wire w_dff_A_CWvdlzJN9_0;
	wire w_dff_A_bnBL7SIz9_0;
	wire w_dff_A_ZwmTRFwx9_0;
	wire w_dff_A_LdSlPXbY0_0;
	jnot g000(.din(w_G146_0[2]),.dout(n58),.clk(gclk));
	jxor g001(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n59),.clk(gclk));
	jxor g002(.dina(w_n59_0[1]),.dinb(n58),.dout(n60),.clk(gclk));
	jnot g003(.din(w_G953_1[2]),.dout(n61),.clk(gclk));
	jand g004(.dina(w_n61_3[2]),.dinb(w_G234_0[2]),.dout(n62),.clk(gclk));
	jand g005(.dina(w_n62_0[1]),.dinb(w_G221_0[1]),.dout(n63),.clk(gclk));
	jxor g006(.dina(n63),.dinb(w_G137_0[2]),.dout(n64),.clk(gclk));
	jxor g007(.dina(w_G128_1[1]),.dinb(w_G119_0[2]),.dout(n65),.clk(gclk));
	jxor g008(.dina(w_dff_B_iJOcSZc75_0),.dinb(n64),.dout(n66),.clk(gclk));
	jxor g009(.dina(n66),.dinb(w_G110_1[1]),.dout(n67),.clk(gclk));
	jxor g010(.dina(w_n67_0[1]),.dinb(w_n60_0[2]),.dout(n68),.clk(gclk));
	jcb g011(.dina(w_n68_0[1]),.dinb(w_G902_3[2]),.dout(n69));
	jnot g012(.din(w_G902_3[1]),.dout(n70),.clk(gclk));
	jand g013(.dina(w_n70_3[1]),.dinb(w_G234_0[1]),.dout(n71),.clk(gclk));
	jnot g014(.din(w_n71_0[1]),.dout(n72),.clk(gclk));
	jand g015(.dina(n72),.dinb(w_G217_0[2]),.dout(n73),.clk(gclk));
	jxor g016(.dina(w_n73_0[1]),.dinb(n69),.dout(n74),.clk(gclk));
	jnot g017(.din(w_G134_0[2]),.dout(n75),.clk(gclk));
	jxor g018(.dina(w_G137_0[1]),.dinb(n75),.dout(n76),.clk(gclk));
	jnot g019(.din(w_G131_0[1]),.dout(n77),.clk(gclk));
	jxor g020(.dina(w_G146_0[1]),.dinb(w_G143_1[1]),.dout(n78),.clk(gclk));
	jxor g021(.dina(n78),.dinb(w_G128_1[0]),.dout(n79),.clk(gclk));
	jxor g022(.dina(w_n79_0[1]),.dinb(w_n77_0[1]),.dout(n80),.clk(gclk));
	jxor g023(.dina(n80),.dinb(w_dff_B_5VKQOKOj0_1),.dout(n81),.clk(gclk));
	jnot g024(.din(w_G113_0[1]),.dout(n82),.clk(gclk));
	jxor g025(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g026(.dina(n83),.dinb(w_n82_0[1]),.dout(n84),.clk(gclk));
	jnot g027(.din(w_G210_0[2]),.dout(n85),.clk(gclk));
	jcb g028(.dina(w_G953_1[1]),.dinb(w_G237_0[2]),.dout(n86));
	jcb g029(.dina(w_n86_0[1]),.dinb(n85),.dout(n87));
	jxor g030(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g031(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g032(.dina(w_dff_B_pbx0NWAq9_0),.dinb(w_n81_0[2]),.dout(n90),.clk(gclk));
	jand g033(.dina(w_n90_0[2]),.dinb(w_n70_3[0]),.dout(n91),.clk(gclk));
	jxor g034(.dina(n91),.dinb(w_G472_0[1]),.dout(n92),.clk(gclk));
	jand g035(.dina(w_n92_1[2]),.dinb(w_n74_1[1]),.dout(n93),.clk(gclk));
	jcb g036(.dina(w_G902_3[0]),.dinb(w_G237_0[1]),.dout(n94));
	jand g037(.dina(w_n94_0[1]),.dinb(w_G214_0[1]),.dout(n95),.clk(gclk));
	jnot g038(.din(w_n95_0[2]),.dout(n96),.clk(gclk));
	jand g039(.dina(w_n94_0[0]),.dinb(w_G210_0[1]),.dout(n97),.clk(gclk));
	jnot g040(.din(w_G110_1[0]),.dout(n98),.clk(gclk));
	jxor g041(.dina(w_G122_1[1]),.dinb(n98),.dout(n99),.clk(gclk));
	jxor g042(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n100),.clk(gclk));
	jxor g043(.dina(n100),.dinb(w_G101_0[1]),.dout(n101),.clk(gclk));
	jxor g044(.dina(w_n101_0[1]),.dinb(w_n84_0[0]),.dout(n102),.clk(gclk));
	jxor g045(.dina(n102),.dinb(w_dff_B_xd96ETnW8_1),.dout(n103),.clk(gclk));
	jand g046(.dina(w_n61_3[1]),.dinb(w_G224_0[1]),.dout(n104),.clk(gclk));
	jxor g047(.dina(w_n79_0[0]),.dinb(w_G125_0[1]),.dout(n105),.clk(gclk));
	jxor g048(.dina(n105),.dinb(w_dff_B_SLrfBU200_1),.dout(n106),.clk(gclk));
	jxor g049(.dina(n106),.dinb(w_n103_0[1]),.dout(n107),.clk(gclk));
	jand g050(.dina(w_n107_0[2]),.dinb(w_n70_2[2]),.dout(n108),.clk(gclk));
	jxor g051(.dina(w_n108_0[1]),.dinb(w_n97_0[1]),.dout(n109),.clk(gclk));
	jand g052(.dina(w_n109_0[1]),.dinb(w_n96_0[2]),.dout(n110),.clk(gclk));
	jnot g053(.din(w_G221_0[0]),.dout(n111),.clk(gclk));
	jcb g054(.dina(w_n71_0[0]),.dinb(w_dff_B_nwK763Rc6_1),.dout(n112));
	jxor g055(.dina(w_G140_0[1]),.dinb(w_G110_0[2]),.dout(n113),.clk(gclk));
	jand g056(.dina(w_n61_3[0]),.dinb(w_G227_0[1]),.dout(n114),.clk(gclk));
	jxor g057(.dina(n114),.dinb(w_n101_0[0]),.dout(n115),.clk(gclk));
	jxor g058(.dina(n115),.dinb(w_dff_B_XF7aPHFI7_1),.dout(n116),.clk(gclk));
	jxor g059(.dina(n116),.dinb(w_n81_0[1]),.dout(n117),.clk(gclk));
	jand g060(.dina(w_n117_0[2]),.dinb(w_n70_2[1]),.dout(n118),.clk(gclk));
	jxor g061(.dina(w_n118_0[1]),.dinb(w_G469_0[2]),.dout(n119),.clk(gclk));
	jand g062(.dina(w_n119_0[1]),.dinb(w_n112_1[1]),.dout(n120),.clk(gclk));
	jand g063(.dina(w_n120_0[1]),.dinb(w_n110_0[2]),.dout(n121),.clk(gclk));
	jand g064(.dina(w_n121_1[1]),.dinb(w_n93_0[2]),.dout(n122),.clk(gclk));
	jnot g065(.din(w_G478_0[2]),.dout(n123),.clk(gclk));
	jxor g066(.dina(w_G143_1[0]),.dinb(w_G128_0[2]),.dout(n124),.clk(gclk));
	jand g067(.dina(w_n62_0[0]),.dinb(w_G217_0[1]),.dout(n125),.clk(gclk));
	jxor g068(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n126),.clk(gclk));
	jxor g069(.dina(w_G134_0[1]),.dinb(w_G107_0[1]),.dout(n127),.clk(gclk));
	jxor g070(.dina(n127),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g071(.dina(w_dff_B_I98vDFqU9_0),.dinb(n125),.dout(n129),.clk(gclk));
	jxor g072(.dina(n129),.dinb(w_dff_B_m6YuB7hj4_1),.dout(n130),.clk(gclk));
	jand g073(.dina(w_n130_0[2]),.dinb(w_n70_2[0]),.dout(n131),.clk(gclk));
	jxor g074(.dina(w_n131_0[1]),.dinb(w_dff_B_N9MFRpiV9_1),.dout(n132),.clk(gclk));
	jnot g075(.din(w_G475_0[2]),.dout(n133),.clk(gclk));
	jxor g076(.dina(w_G143_0[2]),.dinb(w_n77_0[0]),.dout(n134),.clk(gclk));
	jxor g077(.dina(w_G122_0[2]),.dinb(w_n82_0[0]),.dout(n135),.clk(gclk));
	jxor g078(.dina(n135),.dinb(w_G104_0[1]),.dout(n136),.clk(gclk));
	jnot g079(.din(w_G214_0[0]),.dout(n137),.clk(gclk));
	jcb g080(.dina(w_n86_0[0]),.dinb(n137),.dout(n138));
	jxor g081(.dina(w_dff_B_2iYyE76X8_0),.dinb(w_n60_0[1]),.dout(n139),.clk(gclk));
	jxor g082(.dina(n139),.dinb(n136),.dout(n140),.clk(gclk));
	jxor g083(.dina(n140),.dinb(w_dff_B_NZNl7SDx2_1),.dout(n141),.clk(gclk));
	jand g084(.dina(w_n141_0[2]),.dinb(w_n70_1[2]),.dout(n142),.clk(gclk));
	jxor g085(.dina(w_n142_0[1]),.dinb(w_dff_B_rSVmiRJ22_1),.dout(n143),.clk(gclk));
	jand g086(.dina(w_n143_1[1]),.dinb(w_n132_0[2]),.dout(n144),.clk(gclk));
	jcb g087(.dina(w_n61_2[2]),.dinb(w_dff_B_JPJZpma22_1),.dout(n145));
	jand g088(.dina(w_G237_0[0]),.dinb(w_G234_0[0]),.dout(n146),.clk(gclk));
	jcb g089(.dina(w_n146_0[1]),.dinb(w_n70_1[1]),.dout(n147));
	jcb g090(.dina(w_n147_0[1]),.dinb(w_n145_0[1]),.dout(n148));
	jnot g091(.din(w_n146_0[0]),.dout(n149),.clk(gclk));
	jand g092(.dina(w_n61_2[1]),.dinb(w_G952_0[2]),.dout(n150),.clk(gclk));
	jand g093(.dina(n150),.dinb(n149),.dout(n151),.clk(gclk));
	jnot g094(.din(w_n151_0[2]),.dout(n152),.clk(gclk));
	jand g095(.dina(w_n152_0[1]),.dinb(w_dff_B_YR1gWoKv7_1),.dout(n153),.clk(gclk));
	jnot g096(.din(w_n153_0[2]),.dout(n154),.clk(gclk));
	jand g097(.dina(w_n154_1[1]),.dinb(w_n144_1[2]),.dout(n155),.clk(gclk));
	jand g098(.dina(w_n155_0[2]),.dinb(w_n122_0[1]),.dout(n156),.clk(gclk));
	jxor g099(.dina(w_n156_0[1]),.dinb(w_G101_0[0]),.dout(G3),.clk(gclk));
	jnot g100(.din(w_n92_1[1]),.dout(n158),.clk(gclk));
	jand g101(.dina(w_n158_1[1]),.dinb(w_n74_1[0]),.dout(n159),.clk(gclk));
	jand g102(.dina(w_n159_1[1]),.dinb(w_n121_1[0]),.dout(n160),.clk(gclk));
	jxor g103(.dina(w_n142_0[0]),.dinb(w_G475_0[1]),.dout(n161),.clk(gclk));
	jand g104(.dina(w_n161_0[2]),.dinb(w_n132_0[1]),.dout(n162),.clk(gclk));
	jand g105(.dina(w_n162_0[1]),.dinb(w_n154_1[0]),.dout(n163),.clk(gclk));
	jand g106(.dina(w_n163_0[2]),.dinb(w_n160_0[1]),.dout(n164),.clk(gclk));
	jxor g107(.dina(w_n164_0[1]),.dinb(w_G104_0[0]),.dout(G6),.clk(gclk));
	jxor g108(.dina(w_n131_0[0]),.dinb(w_G478_0[1]),.dout(n166),.clk(gclk));
	jand g109(.dina(w_n143_1[0]),.dinb(w_n166_1[1]),.dout(n167),.clk(gclk));
	jand g110(.dina(w_n167_0[1]),.dinb(w_n154_0[2]),.dout(n168),.clk(gclk));
	jand g111(.dina(w_n168_0[2]),.dinb(w_n160_0[0]),.dout(n169),.clk(gclk));
	jxor g112(.dina(w_n169_0[1]),.dinb(w_G107_0[0]),.dout(G9),.clk(gclk));
	jnot g113(.din(w_n60_0[0]),.dout(n171),.clk(gclk));
	jxor g114(.dina(w_n67_0[0]),.dinb(w_dff_B_WHlG6HFB2_1),.dout(n172),.clk(gclk));
	jand g115(.dina(w_n172_0[1]),.dinb(w_n70_1[0]),.dout(n173),.clk(gclk));
	jxor g116(.dina(w_n73_0[0]),.dinb(n173),.dout(n174),.clk(gclk));
	jand g117(.dina(w_n158_1[0]),.dinb(w_n174_1[1]),.dout(n175),.clk(gclk));
	jand g118(.dina(w_n175_0[1]),.dinb(w_n155_0[1]),.dout(n176),.clk(gclk));
	jand g119(.dina(n176),.dinb(w_n121_0[2]),.dout(n177),.clk(gclk));
	jxor g120(.dina(w_n177_0[1]),.dinb(w_G110_0[1]),.dout(G12),.clk(gclk));
	jand g121(.dina(w_n92_1[0]),.dinb(w_n174_1[0]),.dout(n179),.clk(gclk));
	jand g122(.dina(w_n179_0[2]),.dinb(w_n121_0[1]),.dout(n180),.clk(gclk));
	jcb g123(.dina(w_n61_2[0]),.dinb(w_dff_B_vdJpMGfu1_1),.dout(n181));
	jcb g124(.dina(w_n181_0[2]),.dinb(w_n147_0[0]),.dout(n182));
	jand g125(.dina(w_dff_B_jMQCyKhi9_0),.dinb(w_n152_0[0]),.dout(n183),.clk(gclk));
	jnot g126(.din(w_n183_0[2]),.dout(n184),.clk(gclk));
	jand g127(.dina(w_n184_1[1]),.dinb(w_n167_0[0]),.dout(n185),.clk(gclk));
	jand g128(.dina(w_n185_0[2]),.dinb(w_n180_0[1]),.dout(n186),.clk(gclk));
	jxor g129(.dina(w_n186_0[1]),.dinb(w_G128_0[1]),.dout(G30),.clk(gclk));
	jand g130(.dina(w_n161_0[1]),.dinb(w_n166_1[0]),.dout(n188),.clk(gclk));
	jand g131(.dina(w_n188_0[2]),.dinb(w_n184_1[0]),.dout(n189),.clk(gclk));
	jand g132(.dina(w_n189_0[1]),.dinb(w_n122_0[0]),.dout(n190),.clk(gclk));
	jxor g133(.dina(w_n190_0[1]),.dinb(w_G143_0[1]),.dout(G45),.clk(gclk));
	jand g134(.dina(w_n184_0[2]),.dinb(w_n162_0[0]),.dout(n192),.clk(gclk));
	jand g135(.dina(w_n192_0[2]),.dinb(w_n180_0[0]),.dout(n193),.clk(gclk));
	jxor g136(.dina(w_n193_0[1]),.dinb(w_G146_0[0]),.dout(G48),.clk(gclk));
	jnot g137(.din(w_G469_0[1]),.dout(n195),.clk(gclk));
	jxor g138(.dina(w_n118_0[0]),.dinb(w_dff_B_b35UPb6X8_1),.dout(n196),.clk(gclk));
	jand g139(.dina(w_n196_0[2]),.dinb(w_n112_1[0]),.dout(n197),.clk(gclk));
	jand g140(.dina(w_n197_1[1]),.dinb(w_n110_0[1]),.dout(n198),.clk(gclk));
	jand g141(.dina(w_n198_1[1]),.dinb(w_n93_0[1]),.dout(n199),.clk(gclk));
	jand g142(.dina(w_n199_0[1]),.dinb(w_n163_0[1]),.dout(n200),.clk(gclk));
	jxor g143(.dina(w_n200_0[1]),.dinb(w_G113_0[0]),.dout(G15),.clk(gclk));
	jand g144(.dina(w_n199_0[0]),.dinb(w_n168_0[1]),.dout(n202),.clk(gclk));
	jxor g145(.dina(w_n202_0[1]),.dinb(w_G116_0[0]),.dout(G18),.clk(gclk));
	jand g146(.dina(w_n198_1[0]),.dinb(w_n179_0[1]),.dout(n204),.clk(gclk));
	jand g147(.dina(n204),.dinb(w_n155_0[0]),.dout(n205),.clk(gclk));
	jxor g148(.dina(w_n205_0[1]),.dinb(w_G119_0[0]),.dout(G21),.clk(gclk));
	jand g149(.dina(w_n197_1[0]),.dinb(w_n159_1[0]),.dout(n207),.clk(gclk));
	jand g150(.dina(w_n154_0[1]),.dinb(w_n110_0[0]),.dout(n208),.clk(gclk));
	jand g151(.dina(n208),.dinb(w_n188_0[1]),.dout(n209),.clk(gclk));
	jand g152(.dina(n209),.dinb(w_n207_0[1]),.dout(n210),.clk(gclk));
	jxor g153(.dina(w_n210_0[1]),.dinb(w_G122_0[1]),.dout(G24),.clk(gclk));
	jand g154(.dina(w_n192_0[1]),.dinb(w_n175_0[0]),.dout(n212),.clk(gclk));
	jand g155(.dina(w_n212_0[1]),.dinb(w_n198_0[2]),.dout(n213),.clk(gclk));
	jxor g156(.dina(w_n213_0[1]),.dinb(w_G125_0[0]),.dout(G27),.clk(gclk));
	jnot g157(.din(w_n97_0[0]),.dout(n215),.clk(gclk));
	jxor g158(.dina(w_n108_0[0]),.dinb(w_dff_B_PFrBXyXU6_1),.dout(n216),.clk(gclk));
	jand g159(.dina(w_n216_0[2]),.dinb(w_n96_0[1]),.dout(n217),.clk(gclk));
	jand g160(.dina(w_n217_0[2]),.dinb(w_n120_0[0]),.dout(n218),.clk(gclk));
	jand g161(.dina(w_n218_1[1]),.dinb(w_n93_0[0]),.dout(n219),.clk(gclk));
	jand g162(.dina(w_n219_0[1]),.dinb(w_n192_0[0]),.dout(n220),.clk(gclk));
	jxor g163(.dina(w_n220_0[1]),.dinb(w_G131_0[0]),.dout(G33),.clk(gclk));
	jand g164(.dina(w_n219_0[0]),.dinb(w_n185_0[1]),.dout(n222),.clk(gclk));
	jxor g165(.dina(w_n222_0[1]),.dinb(w_G134_0[0]),.dout(G36),.clk(gclk));
	jand g166(.dina(w_n184_0[1]),.dinb(w_n144_1[1]),.dout(n224),.clk(gclk));
	jand g167(.dina(w_dff_B_y5Ms6zHM2_0),.dinb(w_n179_0[0]),.dout(n225),.clk(gclk));
	jand g168(.dina(n225),.dinb(w_n218_1[0]),.dout(n226),.clk(gclk));
	jxor g169(.dina(w_n226_0[1]),.dinb(w_G137_0[0]),.dout(G39),.clk(gclk));
	jand g170(.dina(w_n218_0[2]),.dinb(w_n212_0[0]),.dout(n228),.clk(gclk));
	jxor g171(.dina(w_n228_0[1]),.dinb(w_G140_0[0]),.dout(G42),.clk(gclk));
	jcb g172(.dina(w_n177_0[0]),.dinb(w_n169_0[0]),.dout(n230));
	jcb g173(.dina(w_n202_0[0]),.dinb(w_n164_0[0]),.dout(n231));
	jcb g174(.dina(w_dff_B_dSziAO2Z1_0),.dinb(n230),.dout(n232));
	jcb g175(.dina(w_n205_0[0]),.dinb(w_n156_0[0]),.dout(n233));
	jcb g176(.dina(w_n210_0[0]),.dinb(w_n200_0[0]),.dout(n234));
	jcb g177(.dina(w_dff_B_nI5fi7wz8_0),.dinb(n233),.dout(n235));
	jcb g178(.dina(n235),.dinb(n232),.dout(n236));
	jcb g179(.dina(w_n220_0[0]),.dinb(w_n193_0[0]),.dout(n237));
	jcb g180(.dina(w_n222_0[0]),.dinb(w_n186_0[0]),.dout(n238));
	jcb g181(.dina(n238),.dinb(n237),.dout(n239));
	jcb g182(.dina(w_n228_0[0]),.dinb(w_n190_0[0]),.dout(n240));
	jcb g183(.dina(w_n226_0[0]),.dinb(w_n213_0[0]),.dout(n241));
	jcb g184(.dina(n241),.dinb(n240),.dout(n242));
	jcb g185(.dina(n242),.dinb(n239),.dout(n243));
	jcb g186(.dina(n243),.dinb(n236),.dout(n244));
	jcb g187(.dina(w_n218_0[1]),.dinb(w_n198_0[1]),.dout(n245));
	jand g188(.dina(n245),.dinb(w_n144_1[0]),.dout(n246),.clk(gclk));
	jand g189(.dina(w_n217_0[1]),.dinb(w_n197_0[2]),.dout(n247),.clk(gclk));
	jxor g190(.dina(w_n143_0[2]),.dinb(w_n132_0[0]),.dout(n248),.clk(gclk));
	jand g191(.dina(w_dff_B_Leox0wox6_0),.dinb(n247),.dout(n249),.clk(gclk));
	jcb g192(.dina(n249),.dinb(n246),.dout(n250));
	jand g193(.dina(n250),.dinb(w_n159_0[2]),.dout(n251),.clk(gclk));
	jand g194(.dina(w_n217_0[0]),.dinb(w_n144_0[2]),.dout(n252),.clk(gclk));
	jcb g195(.dina(w_n92_0[2]),.dinb(w_n174_0[2]),.dout(n253));
	jcb g196(.dina(w_n158_0[2]),.dinb(w_n74_0[2]),.dout(n254));
	jand g197(.dina(w_n197_0[1]),.dinb(w_n254_1[1]),.dout(n255),.clk(gclk));
	jand g198(.dina(n255),.dinb(w_n253_0[2]),.dout(n256),.clk(gclk));
	jand g199(.dina(n256),.dinb(w_n252_0[1]),.dout(n257),.clk(gclk));
	jcb g200(.dina(n257),.dinb(n251),.dout(n258));
	jand g201(.dina(n258),.dinb(w_n151_0[1]),.dout(n259),.clk(gclk));
	jxor g202(.dina(w_n112_0[2]),.dinb(w_n96_0[0]),.dout(n260),.clk(gclk));
	jand g203(.dina(n260),.dinb(w_n151_0[0]),.dout(n261),.clk(gclk));
	jand g204(.dina(w_dff_B_DTiGo68Z0_0),.dinb(w_n196_0[1]),.dout(n262),.clk(gclk));
	jand g205(.dina(n262),.dinb(w_n216_0[1]),.dout(n263),.clk(gclk));
	jand g206(.dina(w_n159_0[1]),.dinb(w_n144_0[1]),.dout(n264),.clk(gclk));
	jand g207(.dina(n264),.dinb(w_dff_B_UUkHKZoh3_1),.dout(n265),.clk(gclk));
	jcb g208(.dina(w_dff_B_KZlQMPHE0_0),.dinb(n259),.dout(n266));
	jcb g209(.dina(n266),.dinb(w_n244_2[2]),.dout(n267));
	jand g210(.dina(n267),.dinb(w_G952_0[1]),.dout(n268),.clk(gclk));
	jand g211(.dina(w_n252_0[0]),.dinb(w_n207_0[0]),.dout(n269),.clk(gclk));
	jcb g212(.dina(n269),.dinb(w_G953_1[0]),.dout(n270));
	jcb g213(.dina(w_dff_B_aMa4dRVW8_0),.dinb(n268),.dout(G75));
	jnot g214(.din(w_n107_0[1]),.dout(n272),.clk(gclk));
	jcb g215(.dina(w_n216_0[0]),.dinb(w_n95_0[1]),.dout(n273));
	jnot g216(.din(w_n112_0[1]),.dout(n274),.clk(gclk));
	jcb g217(.dina(w_n196_0[0]),.dinb(w_n274_0[1]),.dout(n275));
	jcb g218(.dina(w_n275_0[1]),.dinb(w_n273_0[2]),.dout(n276));
	jcb g219(.dina(w_n253_0[1]),.dinb(w_n276_1[1]),.dout(n277));
	jnot g220(.din(w_n168_0[0]),.dout(n278),.clk(gclk));
	jcb g221(.dina(w_n278_0[1]),.dinb(w_n277_0[1]),.dout(n279));
	jcb g222(.dina(w_n161_0[0]),.dinb(w_n166_0[2]),.dout(n280));
	jcb g223(.dina(w_n153_0[1]),.dinb(w_n280_0[1]),.dout(n281));
	jcb g224(.dina(w_n92_0[1]),.dinb(w_n74_0[1]),.dout(n282));
	jcb g225(.dina(w_n282_0[1]),.dinb(w_n281_0[2]),.dout(n283));
	jcb g226(.dina(n283),.dinb(w_n276_1[0]),.dout(n284));
	jand g227(.dina(w_dff_B_ESBooY621_0),.dinb(n279),.dout(n285),.clk(gclk));
	jnot g228(.din(w_n163_0[0]),.dout(n286),.clk(gclk));
	jcb g229(.dina(w_n286_0[1]),.dinb(w_n277_0[0]),.dout(n287));
	jcb g230(.dina(w_n158_0[1]),.dinb(w_n174_0[1]),.dout(n288));
	jcb g231(.dina(w_n119_0[0]),.dinb(w_n274_0[0]),.dout(n289));
	jcb g232(.dina(w_n289_0[1]),.dinb(w_n273_0[1]),.dout(n290));
	jcb g233(.dina(w_n290_0[2]),.dinb(w_n288_0[2]),.dout(n291));
	jcb g234(.dina(w_n291_0[1]),.dinb(w_n278_0[0]),.dout(n292));
	jand g235(.dina(n292),.dinb(n287),.dout(n293),.clk(gclk));
	jand g236(.dina(n293),.dinb(n285),.dout(n294),.clk(gclk));
	jcb g237(.dina(w_n276_0[2]),.dinb(w_n288_0[1]),.dout(n295));
	jcb g238(.dina(w_n281_0[1]),.dinb(w_n295_0[1]),.dout(n296));
	jcb g239(.dina(w_n290_0[1]),.dinb(w_n254_1[0]),.dout(n297));
	jcb g240(.dina(n297),.dinb(w_n281_0[0]),.dout(n298));
	jand g241(.dina(w_dff_B_xmAMFAiU6_0),.dinb(n296),.dout(n299),.clk(gclk));
	jcb g242(.dina(w_n291_0[0]),.dinb(w_n286_0[0]),.dout(n300));
	jcb g243(.dina(w_n289_0[0]),.dinb(w_n253_0[0]),.dout(n301));
	jnot g244(.din(w_n188_0[0]),.dout(n302),.clk(gclk));
	jcb g245(.dina(w_n153_0[0]),.dinb(w_n273_0[0]),.dout(n303));
	jcb g246(.dina(w_dff_B_nlL1oXQa2_0),.dinb(n302),.dout(n304));
	jcb g247(.dina(n304),.dinb(n301),.dout(n305));
	jand g248(.dina(w_dff_B_Jkj5CeEG9_0),.dinb(n300),.dout(n306),.clk(gclk));
	jand g249(.dina(n306),.dinb(w_dff_B_IzJsr9a93_1),.dout(n307),.clk(gclk));
	jand g250(.dina(n307),.dinb(n294),.dout(n308),.clk(gclk));
	jcb g251(.dina(w_n254_0[2]),.dinb(w_n276_0[1]),.dout(n309));
	jcb g252(.dina(w_n143_0[1]),.dinb(w_n166_0[1]),.dout(n310));
	jcb g253(.dina(w_n183_0[1]),.dinb(n310),.dout(n311));
	jcb g254(.dina(w_n311_0[2]),.dinb(w_n309_0[1]),.dout(n312));
	jcb g255(.dina(w_n109_0[0]),.dinb(w_n95_0[0]),.dout(n313));
	jcb g256(.dina(n313),.dinb(w_n275_0[0]),.dout(n314));
	jcb g257(.dina(w_n314_0[2]),.dinb(w_n288_0[0]),.dout(n315));
	jcb g258(.dina(w_n315_0[1]),.dinb(w_n311_0[1]),.dout(n316));
	jand g259(.dina(n316),.dinb(w_dff_B_KxqXcm3f6_1),.dout(n317),.clk(gclk));
	jnot g260(.din(w_n185_0[0]),.dout(n318),.clk(gclk));
	jcb g261(.dina(w_n318_0[1]),.dinb(w_n309_0[0]),.dout(n319));
	jcb g262(.dina(w_n315_0[0]),.dinb(w_n318_0[0]),.dout(n320));
	jand g263(.dina(n320),.dinb(n319),.dout(n321),.clk(gclk));
	jand g264(.dina(n321),.dinb(w_dff_B_syV6dGNo7_1),.dout(n322),.clk(gclk));
	jnot g265(.din(w_n189_0[0]),.dout(n323),.clk(gclk));
	jcb g266(.dina(n323),.dinb(w_n295_0[0]),.dout(n324));
	jcb g267(.dina(w_n311_0[0]),.dinb(w_n282_0[0]),.dout(n325));
	jcb g268(.dina(w_n314_0[1]),.dinb(w_n325_0[1]),.dout(n326));
	jand g269(.dina(w_dff_B_u1v0oDzC5_0),.dinb(n324),.dout(n327),.clk(gclk));
	jcb g270(.dina(w_n325_0[0]),.dinb(w_n290_0[0]),.dout(n328));
	jcb g271(.dina(w_n183_0[0]),.dinb(w_n280_0[0]),.dout(n329));
	jcb g272(.dina(w_dff_B_SoUsOi0K6_0),.dinb(w_n254_0[1]),.dout(n330));
	jcb g273(.dina(n330),.dinb(w_n314_0[0]),.dout(n331));
	jand g274(.dina(n331),.dinb(n328),.dout(n332),.clk(gclk));
	jand g275(.dina(w_dff_B_UCJLGiV16_0),.dinb(n327),.dout(n333),.clk(gclk));
	jand g276(.dina(n333),.dinb(n322),.dout(n334),.clk(gclk));
	jand g277(.dina(w_n334_0[1]),.dinb(w_n308_0[1]),.dout(n335),.clk(gclk));
	jand g278(.dina(w_G902_2[2]),.dinb(w_G210_0[0]),.dout(n336),.clk(gclk));
	jnot g279(.din(w_n336_0[1]),.dout(n337),.clk(gclk));
	jcb g280(.dina(w_dff_B_qvJFveWg6_0),.dinb(w_n335_2[1]),.dout(n338));
	jcb g281(.dina(n338),.dinb(w_dff_B_4JD1duB90_1),.dout(n339));
	jcb g282(.dina(w_n61_1[2]),.dinb(w_G952_0[0]),.dout(n340));
	jand g283(.dina(w_n336_0[0]),.dinb(w_n244_2[1]),.dout(n341),.clk(gclk));
	jcb g284(.dina(n341),.dinb(w_n107_0[0]),.dout(n342));
	jand g285(.dina(n342),.dinb(w_n340_2[1]),.dout(n343),.clk(gclk));
	jand g286(.dina(n343),.dinb(n339),.dout(G51),.clk(gclk));
	jnot g287(.din(w_n117_0[1]),.dout(n345),.clk(gclk));
	jand g288(.dina(w_G902_2[1]),.dinb(w_G469_0[0]),.dout(n346),.clk(gclk));
	jnot g289(.din(w_n346_0[1]),.dout(n347),.clk(gclk));
	jcb g290(.dina(w_dff_B_G06qirAy6_0),.dinb(w_n335_2[0]),.dout(n348));
	jcb g291(.dina(n348),.dinb(w_dff_B_TsqBpAWs7_1),.dout(n349));
	jand g292(.dina(w_n346_0[0]),.dinb(w_n244_2[0]),.dout(n350),.clk(gclk));
	jcb g293(.dina(n350),.dinb(w_n117_0[0]),.dout(n351));
	jand g294(.dina(n351),.dinb(w_n340_2[0]),.dout(n352),.clk(gclk));
	jand g295(.dina(n352),.dinb(n349),.dout(G54),.clk(gclk));
	jnot g296(.din(w_n141_0[1]),.dout(n354),.clk(gclk));
	jand g297(.dina(w_G902_2[0]),.dinb(w_G475_0[0]),.dout(n355),.clk(gclk));
	jnot g298(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jcb g299(.dina(w_dff_B_s2kl1zm84_0),.dinb(w_n335_1[2]),.dout(n357));
	jcb g300(.dina(n357),.dinb(w_dff_B_0cRPFybT1_1),.dout(n358));
	jand g301(.dina(w_n355_0[0]),.dinb(w_n244_1[2]),.dout(n359),.clk(gclk));
	jcb g302(.dina(n359),.dinb(w_n141_0[0]),.dout(n360));
	jand g303(.dina(n360),.dinb(w_n340_1[2]),.dout(n361),.clk(gclk));
	jand g304(.dina(n361),.dinb(n358),.dout(G60),.clk(gclk));
	jnot g305(.din(w_n130_0[1]),.dout(n363),.clk(gclk));
	jand g306(.dina(w_G902_1[2]),.dinb(w_G478_0[0]),.dout(n364),.clk(gclk));
	jnot g307(.din(w_n364_0[1]),.dout(n365),.clk(gclk));
	jcb g308(.dina(w_dff_B_iVxIWCT72_0),.dinb(w_n335_1[1]),.dout(n366));
	jcb g309(.dina(n366),.dinb(w_dff_B_GUcOIG9m7_1),.dout(n367));
	jand g310(.dina(w_n364_0[0]),.dinb(w_n244_1[1]),.dout(n368),.clk(gclk));
	jcb g311(.dina(n368),.dinb(w_n130_0[0]),.dout(n369));
	jand g312(.dina(n369),.dinb(w_n340_1[1]),.dout(n370),.clk(gclk));
	jand g313(.dina(n370),.dinb(n367),.dout(G63),.clk(gclk));
	jand g314(.dina(w_G902_1[1]),.dinb(w_G217_0[0]),.dout(n372),.clk(gclk));
	jand g315(.dina(w_n372_0[1]),.dinb(w_n244_1[0]),.dout(n373),.clk(gclk));
	jcb g316(.dina(n373),.dinb(w_n172_0[0]),.dout(n374));
	jnot g317(.din(w_n372_0[0]),.dout(n375),.clk(gclk));
	jcb g318(.dina(w_dff_B_2KeNDtYV1_0),.dinb(w_n335_1[0]),.dout(n376));
	jcb g319(.dina(n376),.dinb(w_n68_0[0]),.dout(n377));
	jand g320(.dina(n377),.dinb(w_n340_1[0]),.dout(n378),.clk(gclk));
	jand g321(.dina(n378),.dinb(w_dff_B_MgoIaZ0d6_1),.dout(G66),.clk(gclk));
	jnot g322(.din(w_n145_0[0]),.dout(n380),.clk(gclk));
	jcb g323(.dina(w_n308_0[0]),.dinb(w_G953_0[2]),.dout(n381));
	jcb g324(.dina(w_n61_1[1]),.dinb(w_G224_0[0]),.dout(n382));
	jand g325(.dina(w_dff_B_h3nV6xkx4_0),.dinb(n381),.dout(n383),.clk(gclk));
	jxor g326(.dina(n383),.dinb(w_n103_0[0]),.dout(n384),.clk(gclk));
	jcb g327(.dina(n384),.dinb(w_dff_B_FpHpHvB37_1),.dout(G69));
	jcb g328(.dina(w_n334_0[0]),.dinb(w_G953_0[1]),.dout(n386));
	jcb g329(.dina(w_n61_1[0]),.dinb(w_G227_0[0]),.dout(n387));
	jand g330(.dina(n387),.dinb(w_n181_0[1]),.dout(n388),.clk(gclk));
	jand g331(.dina(w_dff_B_QcpHiPlY3_0),.dinb(n386),.dout(n389),.clk(gclk));
	jnot g332(.din(w_n181_0[0]),.dout(n390),.clk(gclk));
	jxor g333(.dina(w_n81_0[0]),.dinb(w_n59_0[0]),.dout(n391),.clk(gclk));
	jcb g334(.dina(n391),.dinb(w_dff_B_022ZCcFP7_1),.dout(n392));
	jxor g335(.dina(w_dff_B_61pLk6yF7_0),.dinb(n389),.dout(G72),.clk(gclk));
	jnot g336(.din(w_n90_0[1]),.dout(n394),.clk(gclk));
	jand g337(.dina(w_G902_1[0]),.dinb(w_G472_0[0]),.dout(n395),.clk(gclk));
	jnot g338(.din(w_n395_0[1]),.dout(n396),.clk(gclk));
	jcb g339(.dina(w_dff_B_AjK9z4Zd6_0),.dinb(w_n335_0[2]),.dout(n397));
	jcb g340(.dina(n397),.dinb(w_dff_B_Czv2JzUB9_1),.dout(n398));
	jand g341(.dina(w_n395_0[0]),.dinb(w_n244_0[2]),.dout(n399),.clk(gclk));
	jcb g342(.dina(n399),.dinb(w_n90_0[0]),.dout(n400));
	jand g343(.dina(n400),.dinb(w_n340_0[2]),.dout(n401),.clk(gclk));
	jand g344(.dina(n401),.dinb(n398),.dout(G57),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_dff_A_SPqektBu0_0),.doutb(w_G101_0[1]),.doutc(w_G101_0[2]),.din(w_dff_B_IWk5oVRb7_3));
	jspl3 jspl3_w_G104_0(.douta(w_dff_A_3LXgP0c93_0),.doutb(w_dff_A_zNv4tfBu4_1),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_dff_A_XFy2QIpz0_0),.doutb(w_G107_0[1]),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_G110_0[0]),.doutb(w_dff_A_6Y0SRe8A8_1),.doutc(w_G110_0[2]),.din(G110));
	jspl jspl_w_G110_1(.douta(w_G110_1[0]),.doutb(w_dff_A_4oX8d2lL8_1),.din(w_G110_0[0]));
	jspl jspl_w_G113_0(.douta(w_dff_A_Vz1GAtqw7_0),.doutb(w_G113_0[1]),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_dff_A_tyrBzHzI7_0),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_dff_A_wOPgZHQT5_0),.doutb(w_G119_0[1]),.doutc(w_G119_0[2]),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_dff_A_XdZ53zG34_1),.doutc(w_dff_A_ny2tcttW0_2),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_dff_A_9DdSNxao3_1),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_dff_A_TZgUmoyB5_0),.doutb(w_dff_A_7RDDJqxm0_1),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_dff_A_Ieji7Bl78_1),.doutc(w_G128_0[2]),.din(G128));
	jspl jspl_w_G128_1(.douta(w_dff_A_JRAGx0Nq6_0),.doutb(w_G128_1[1]),.din(w_G128_0[0]));
	jspl jspl_w_G131_0(.douta(w_dff_A_NvTiZtab6_0),.doutb(w_G131_0[1]),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_dff_A_LdSlPXbY0_0),.doutb(w_G134_0[1]),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_VfRoeoli6_0),.doutb(w_G137_0[1]),.doutc(w_dff_A_seMvB0Zz0_2),.din(w_dff_B_Yb2Y004C3_3));
	jspl3 jspl3_w_G140_0(.douta(w_dff_A_1T56NcLb3_0),.doutb(w_G140_0[1]),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_dff_A_McHXRgtX7_1),.doutc(w_dff_A_P79p6jqT7_2),.din(G143));
	jspl jspl_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.din(w_G143_0[0]));
	jspl3 jspl3_w_G146_0(.douta(w_dff_A_IqzNrTTb5_0),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(G146));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_G210_0[2]),.din(G210));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_G214_0[1]),.din(G214));
	jspl3 jspl3_w_G217_0(.douta(w_G217_0[0]),.doutb(w_dff_A_VehClCCv1_1),.doutc(w_dff_A_MOEusTo60_2),.din(G217));
	jspl jspl_w_G221_0(.douta(w_G221_0[0]),.doutb(w_dff_A_epkGa6cy4_1),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_G224_0[1]),.din(w_dff_B_j8NchfuQ0_2));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_G227_0[1]),.din(w_dff_B_XwWUbyaA9_2));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_dff_A_gsFWYLBg9_1),.doutc(w_dff_A_El32Yq4F9_2),.din(G234));
	jspl3 jspl3_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.doutc(w_G237_0[2]),.din(G237));
	jspl3 jspl3_w_G469_0(.douta(w_G469_0[0]),.doutb(w_G469_0[1]),.doutc(w_dff_A_wRghbfZ99_2),.din(G469));
	jspl jspl_w_G472_0(.douta(w_G472_0[0]),.doutb(w_dff_A_PiOiHVkx0_1),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_dff_A_a4VxBFAt6_1),.doutc(w_G475_0[2]),.din(G475));
	jspl3 jspl3_w_G478_0(.douta(w_G478_0[0]),.doutb(w_dff_A_3qplDVlv4_1),.doutc(w_G478_0[2]),.din(G478));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_G902_0[2]),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_G902_1[1]),.doutc(w_G902_1[2]),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_G902_2[1]),.doutc(w_G902_2[2]),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_G902_3[0]),.doutb(w_G902_3[1]),.doutc(w_dff_A_oa6Wi5jE0_2),.din(w_G902_0[2]));
	jspl3 jspl3_w_G952_0(.douta(w_G952_0[0]),.doutb(w_dff_A_sfXzP4f65_1),.doutc(w_G952_0[2]),.din(w_dff_B_fdscj1JI9_3));
	jspl3 jspl3_w_G953_0(.douta(w_G953_0[0]),.doutb(w_dff_A_O2HRP7rs9_1),.doutc(w_dff_A_ddUKeo2G2_2),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_dff_A_jKJOKbtK3_0),.doutb(w_G953_1[1]),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl jspl_w_n59_0(.douta(w_dff_A_oD3XMy220_0),.doutb(w_n59_0[1]),.din(n59));
	jspl3 jspl3_w_n60_0(.douta(w_n60_0[0]),.doutb(w_n60_0[1]),.doutc(w_dff_A_9Q4mYpeZ7_2),.din(n60));
	jspl3 jspl3_w_n61_0(.douta(w_n61_0[0]),.doutb(w_n61_0[1]),.doutc(w_n61_0[2]),.din(n61));
	jspl3 jspl3_w_n61_1(.douta(w_n61_1[0]),.doutb(w_n61_1[1]),.doutc(w_n61_1[2]),.din(w_n61_0[0]));
	jspl3 jspl3_w_n61_2(.douta(w_n61_2[0]),.doutb(w_n61_2[1]),.doutc(w_n61_2[2]),.din(w_n61_0[1]));
	jspl3 jspl3_w_n61_3(.douta(w_n61_3[0]),.doutb(w_n61_3[1]),.doutc(w_n61_3[2]),.din(w_n61_0[2]));
	jspl jspl_w_n62_0(.douta(w_n62_0[0]),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n68_0(.douta(w_dff_A_Fc7Heav51_0),.doutb(w_n68_0[1]),.din(n68));
	jspl3 jspl3_w_n70_0(.douta(w_n70_0[0]),.doutb(w_dff_A_JXaWVVBu4_1),.doutc(w_n70_0[2]),.din(n70));
	jspl3 jspl3_w_n70_1(.douta(w_dff_A_4Pgu4pSc6_0),.doutb(w_n70_1[1]),.doutc(w_dff_A_1Clx8xz59_2),.din(w_n70_0[0]));
	jspl3 jspl3_w_n70_2(.douta(w_n70_2[0]),.doutb(w_n70_2[1]),.doutc(w_n70_2[2]),.din(w_n70_0[1]));
	jspl jspl_w_n70_3(.douta(w_dff_A_4wBYh1qH1_0),.doutb(w_n70_3[1]),.din(w_n70_0[2]));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n73_0(.douta(w_dff_A_zI8VUVET9_0),.doutb(w_n73_0[1]),.din(w_dff_B_OPpNW5H85_2));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_dff_A_B1IMyYbE1_1),.din(n77));
	jspl jspl_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.din(n79));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl jspl_w_n82_0(.douta(w_n82_0[0]),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(w_dff_B_2dX0KMoU9_2));
	jspl3 jspl3_w_n90_0(.douta(w_dff_A_xEf78y8R0_0),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_dff_A_vYcfVLIy1_1),.doutc(w_dff_A_gjC2y7aA7_2),.din(n92));
	jspl3 jspl3_w_n92_1(.douta(w_dff_A_S0id8zff3_0),.doutb(w_n92_1[1]),.doutc(w_dff_A_c9ksjVia9_2),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n95_0(.douta(w_dff_A_4sr6rX5J6_0),.doutb(w_dff_A_yUMrUTrr4_1),.doutc(w_n95_0[2]),.din(n95));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_dff_A_e2uwbNNi9_1),.doutc(w_dff_A_HQSc0RKe9_2),.din(n96));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_dff_A_VN6hA1Nm1_1),.din(n97));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_dff_A_8dtt8jhM9_0),.doutb(w_n103_0[1]),.din(n103));
	jspl3 jspl3_w_n107_0(.douta(w_dff_A_A4XgrKl65_0),.doutb(w_n107_0[1]),.doutc(w_n107_0[2]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.doutc(w_n110_0[2]),.din(n110));
	jspl3 jspl3_w_n112_0(.douta(w_dff_A_vi6JzD1y3_0),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl jspl_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_dff_A_PHCmtKUe5_0),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_dff_A_3qPQklFW8_1),.doutc(w_dff_A_pod2XMWh3_2),.din(n121));
	jspl jspl_w_n121_1(.douta(w_n121_1[0]),.doutb(w_n121_1[1]),.din(w_n121_0[0]));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.din(n122));
	jspl3 jspl3_w_n130_0(.douta(w_dff_A_YhyKNndE6_0),.doutb(w_n130_0[1]),.doutc(w_n130_0[2]),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n141_0(.douta(w_dff_A_1WZ6LAoB7_0),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl3 jspl3_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.doutc(w_n143_0[2]),.din(n143));
	jspl jspl_w_n143_1(.douta(w_n143_1[0]),.doutb(w_n143_1[1]),.din(w_n143_0[0]));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_dff_A_1wrvM3uX4_1),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n144_1(.douta(w_dff_A_7t150ZsV1_0),.doutb(w_n144_1[1]),.doutc(w_n144_1[2]),.din(w_n144_0[0]));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_D7oeaaDe2_1),.doutc(w_n151_0[2]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_dff_A_S4xbV8Hs5_0),.doutb(w_dff_A_Ro2hpgkn1_1),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_n154_0[2]),.din(w_dff_B_fNgSMBRA9_3));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl3 jspl3_w_n155_0(.douta(w_dff_A_dA8Bc4bg1_0),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(w_dff_B_7SPTAqeQ4_3));
	jspl jspl_w_n156_0(.douta(w_dff_A_8rWjRxp07_0),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n158_0(.douta(w_n158_0[0]),.doutb(w_dff_A_KQ9LXcof3_1),.doutc(w_n158_0[2]),.din(n158));
	jspl jspl_w_n158_1(.douta(w_dff_A_8YxqbqHk9_0),.doutb(w_n158_1[1]),.din(w_n158_0[0]));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_dff_A_zs3zT8BU7_2),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_dff_A_psk5xJCz6_1),.doutc(w_dff_A_JH53DPRX5_2),.din(n163));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl jspl_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.din(w_n166_0[0]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_dff_A_xLqE1JzG5_1),.doutc(w_dff_A_9ptEOAnV7_2),.din(n168));
	jspl jspl_w_n169_0(.douta(w_dff_A_YONZmBkR0_0),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n172_0(.douta(w_dff_A_FnkGLtEb5_0),.doutb(w_n172_0[1]),.din(n172));
	jspl3 jspl3_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.doutc(w_n174_0[2]),.din(n174));
	jspl jspl_w_n174_1(.douta(w_n174_1[0]),.doutb(w_n174_1[1]),.din(w_n174_0[0]));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_n179_0[1]),.doutc(w_n179_0[2]),.din(n179));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n183_0(.douta(w_dff_A_3t72QqKb7_0),.doutb(w_dff_A_vPrrgWUx2_1),.doutc(w_n183_0[2]),.din(n183));
	jspl3 jspl3_w_n184_0(.douta(w_n184_0[0]),.doutb(w_n184_0[1]),.doutc(w_n184_0[2]),.din(w_dff_B_01Sj3U7Z8_3));
	jspl jspl_w_n184_1(.douta(w_n184_1[0]),.doutb(w_n184_1[1]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_dff_A_1OKfejET8_1),.doutc(w_dff_A_0Epgjh5R4_2),.din(n185));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl3 jspl3_w_n188_0(.douta(w_n188_0[0]),.doutb(w_dff_A_wPCGl1qU9_1),.doutc(w_n188_0[2]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_dff_A_Co56wZdW7_1),.din(n189));
	jspl jspl_w_n190_0(.douta(w_dff_A_TTLwkGB22_0),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.doutc(w_dff_A_Fa2UMt9f5_2),.din(w_dff_B_axGrS3Iv1_3));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.din(n193));
	jspl3 jspl3_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.doutc(w_n196_0[2]),.din(n196));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_dff_A_Vd29EL2O1_0),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_dff_A_2B8NSCZf5_2),.din(n198));
	jspl jspl_w_n198_1(.douta(w_dff_A_BNL5dXN84_0),.doutb(w_n198_1[1]),.din(w_n198_0[0]));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_dff_A_71NluWUL3_1),.doutc(w_n216_0[2]),.din(n216));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_dff_A_LcBlZ9aX5_2),.din(n218));
	jspl jspl_w_n218_1(.douta(w_dff_A_PGts8FVS1_0),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_dff_A_o6iHd4wS5_0),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n222_0(.douta(w_dff_A_kenMqaJC9_0),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl3 jspl3_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.doutc(w_n244_0[2]),.din(n244));
	jspl3 jspl3_w_n244_1(.douta(w_n244_1[0]),.doutb(w_n244_1[1]),.doutc(w_n244_1[2]),.din(w_n244_0[0]));
	jspl3 jspl3_w_n244_2(.douta(w_n244_2[0]),.doutb(w_n244_2[1]),.doutc(w_n244_2[2]),.din(w_n244_0[1]));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(w_dff_B_x3X379eF2_2));
	jspl3 jspl3_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.doutc(w_n253_0[2]),.din(n253));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl jspl_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.doutc(w_n273_0[2]),.din(n273));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(w_dff_B_iXVu6Lhd7_2));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl3 jspl3_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.doutc(w_dff_A_uMjKPJT36_2),.din(w_dff_B_bhRoY6r93_3));
	jspl jspl_w_n276_1(.douta(w_n276_1[0]),.doutb(w_dff_A_CN1DHKJk6_1),.din(w_n276_0[0]));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(w_dff_B_CwepJYR72_2));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(n278));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n281_0(.douta(w_n281_0[0]),.doutb(w_dff_A_clZThNqh3_1),.doutc(w_n281_0[2]),.din(w_dff_B_U6R6kNON7_3));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(n286));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n289_0(.douta(w_dff_A_oIpNTQ8z8_0),.doutb(w_n289_0[1]),.din(n289));
	jspl3 jspl3_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.doutc(w_dff_A_FApMqmB96_2),.din(w_dff_B_HhfOLex49_3));
	jspl jspl_w_n291_0(.douta(w_n291_0[0]),.doutb(w_n291_0[1]),.din(w_dff_B_ElRGm0qY9_2));
	jspl jspl_w_n295_0(.douta(w_dff_A_0TVHd13F1_0),.doutb(w_n295_0[1]),.din(n295));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_dff_A_GFsw4uTu9_0),.doutb(w_n309_0[1]),.din(n309));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_dff_A_WliHaTzo1_1),.doutc(w_n311_0[2]),.din(w_dff_B_Hc8yxGjE5_3));
	jspl3 jspl3_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.doutc(w_dff_A_1QG9NFcn5_2),.din(w_dff_B_YxBQv0KS6_3));
	jspl jspl_w_n315_0(.douta(w_dff_A_ytS0m6ve3_0),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.doutc(w_n335_1[2]),.din(w_n335_0[0]));
	jspl jspl_w_n335_2(.douta(w_n335_2[0]),.doutb(w_n335_2[1]),.din(w_n335_0[1]));
	jspl jspl_w_n336_0(.douta(w_dff_A_4KWj67gY2_0),.doutb(w_n336_0[1]),.din(n336));
	jspl3 jspl3_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.doutc(w_n340_0[2]),.din(w_dff_B_mOt15Rct5_3));
	jspl3 jspl3_w_n340_1(.douta(w_dff_A_rHrGhwGm6_0),.doutb(w_n340_1[1]),.doutc(w_n340_1[2]),.din(w_n340_0[0]));
	jspl jspl_w_n340_2(.douta(w_n340_2[0]),.doutb(w_n340_2[1]),.din(w_n340_0[1]));
	jspl jspl_w_n346_0(.douta(w_dff_A_PhNOj6iL2_0),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n355_0(.douta(w_dff_A_Wi2sX6WX9_0),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n364_0(.douta(w_dff_A_I6BHAfxa8_0),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_TL2yhSof4_1),.din(n372));
	jspl jspl_w_n395_0(.douta(w_dff_A_CTbbxFKx9_0),.doutb(w_n395_0[1]),.din(n395));
	jdff dff_B_qIklqYuI8_0(.din(n270),.dout(w_dff_B_qIklqYuI8_0),.clk(gclk));
	jdff dff_B_aMa4dRVW8_0(.din(w_dff_B_qIklqYuI8_0),.dout(w_dff_B_aMa4dRVW8_0),.clk(gclk));
	jdff dff_B_KZlQMPHE0_0(.din(n265),.dout(w_dff_B_KZlQMPHE0_0),.clk(gclk));
	jdff dff_B_UUkHKZoh3_1(.din(n263),.dout(w_dff_B_UUkHKZoh3_1),.clk(gclk));
	jdff dff_B_Ko9Q0Ouk9_0(.din(n261),.dout(w_dff_B_Ko9Q0Ouk9_0),.clk(gclk));
	jdff dff_B_qLE4qJCR1_0(.din(w_dff_B_Ko9Q0Ouk9_0),.dout(w_dff_B_qLE4qJCR1_0),.clk(gclk));
	jdff dff_B_DTiGo68Z0_0(.din(w_dff_B_qLE4qJCR1_0),.dout(w_dff_B_DTiGo68Z0_0),.clk(gclk));
	jdff dff_B_x3X379eF2_2(.din(n252),.dout(w_dff_B_x3X379eF2_2),.clk(gclk));
	jdff dff_B_Leox0wox6_0(.din(n248),.dout(w_dff_B_Leox0wox6_0),.clk(gclk));
	jdff dff_B_X5b1YLFJ7_1(.din(n272),.dout(w_dff_B_X5b1YLFJ7_1),.clk(gclk));
	jdff dff_B_PbRkO0Ib6_1(.din(w_dff_B_X5b1YLFJ7_1),.dout(w_dff_B_PbRkO0Ib6_1),.clk(gclk));
	jdff dff_B_tZb0ThWF1_1(.din(w_dff_B_PbRkO0Ib6_1),.dout(w_dff_B_tZb0ThWF1_1),.clk(gclk));
	jdff dff_B_p3Y1KmNo3_1(.din(w_dff_B_tZb0ThWF1_1),.dout(w_dff_B_p3Y1KmNo3_1),.clk(gclk));
	jdff dff_B_0kPGg72q9_1(.din(w_dff_B_p3Y1KmNo3_1),.dout(w_dff_B_0kPGg72q9_1),.clk(gclk));
	jdff dff_B_AIw4y7yr9_1(.din(w_dff_B_0kPGg72q9_1),.dout(w_dff_B_AIw4y7yr9_1),.clk(gclk));
	jdff dff_B_wKrwOjjf4_1(.din(w_dff_B_AIw4y7yr9_1),.dout(w_dff_B_wKrwOjjf4_1),.clk(gclk));
	jdff dff_B_4JD1duB90_1(.din(w_dff_B_wKrwOjjf4_1),.dout(w_dff_B_4JD1duB90_1),.clk(gclk));
	jdff dff_B_XpMiKSVd3_0(.din(n337),.dout(w_dff_B_XpMiKSVd3_0),.clk(gclk));
	jdff dff_B_nPgonPMr5_0(.din(w_dff_B_XpMiKSVd3_0),.dout(w_dff_B_nPgonPMr5_0),.clk(gclk));
	jdff dff_B_8MNJWJOr5_0(.din(w_dff_B_nPgonPMr5_0),.dout(w_dff_B_8MNJWJOr5_0),.clk(gclk));
	jdff dff_B_S46GJT483_0(.din(w_dff_B_8MNJWJOr5_0),.dout(w_dff_B_S46GJT483_0),.clk(gclk));
	jdff dff_B_eOBnwvJ22_0(.din(w_dff_B_S46GJT483_0),.dout(w_dff_B_eOBnwvJ22_0),.clk(gclk));
	jdff dff_B_L8DhmnAe5_0(.din(w_dff_B_eOBnwvJ22_0),.dout(w_dff_B_L8DhmnAe5_0),.clk(gclk));
	jdff dff_B_rVCYKYF15_0(.din(w_dff_B_L8DhmnAe5_0),.dout(w_dff_B_rVCYKYF15_0),.clk(gclk));
	jdff dff_B_P2noYk0w1_0(.din(w_dff_B_rVCYKYF15_0),.dout(w_dff_B_P2noYk0w1_0),.clk(gclk));
	jdff dff_B_KHL9ZZiS4_0(.din(w_dff_B_P2noYk0w1_0),.dout(w_dff_B_KHL9ZZiS4_0),.clk(gclk));
	jdff dff_B_vX93nVos8_0(.din(w_dff_B_KHL9ZZiS4_0),.dout(w_dff_B_vX93nVos8_0),.clk(gclk));
	jdff dff_B_IWsozdop8_0(.din(w_dff_B_vX93nVos8_0),.dout(w_dff_B_IWsozdop8_0),.clk(gclk));
	jdff dff_B_qvJFveWg6_0(.din(w_dff_B_IWsozdop8_0),.dout(w_dff_B_qvJFveWg6_0),.clk(gclk));
	jdff dff_A_XiONjEUM2_0(.dout(w_n336_0[0]),.din(w_dff_A_XiONjEUM2_0),.clk(gclk));
	jdff dff_A_YqtWxJyX4_0(.dout(w_dff_A_XiONjEUM2_0),.din(w_dff_A_YqtWxJyX4_0),.clk(gclk));
	jdff dff_A_aTaWS9d60_0(.dout(w_dff_A_YqtWxJyX4_0),.din(w_dff_A_aTaWS9d60_0),.clk(gclk));
	jdff dff_A_mfUZGYf69_0(.dout(w_dff_A_aTaWS9d60_0),.din(w_dff_A_mfUZGYf69_0),.clk(gclk));
	jdff dff_A_xl8xkgtH0_0(.dout(w_dff_A_mfUZGYf69_0),.din(w_dff_A_xl8xkgtH0_0),.clk(gclk));
	jdff dff_A_fIajYCHH2_0(.dout(w_dff_A_xl8xkgtH0_0),.din(w_dff_A_fIajYCHH2_0),.clk(gclk));
	jdff dff_A_xQK1tryG4_0(.dout(w_dff_A_fIajYCHH2_0),.din(w_dff_A_xQK1tryG4_0),.clk(gclk));
	jdff dff_A_MMdwnign8_0(.dout(w_dff_A_xQK1tryG4_0),.din(w_dff_A_MMdwnign8_0),.clk(gclk));
	jdff dff_A_AvyULZ1F5_0(.dout(w_dff_A_MMdwnign8_0),.din(w_dff_A_AvyULZ1F5_0),.clk(gclk));
	jdff dff_A_q6qdmp4l7_0(.dout(w_dff_A_AvyULZ1F5_0),.din(w_dff_A_q6qdmp4l7_0),.clk(gclk));
	jdff dff_A_4KWj67gY2_0(.dout(w_dff_A_q6qdmp4l7_0),.din(w_dff_A_4KWj67gY2_0),.clk(gclk));
	jdff dff_B_4gSGPn0c7_1(.din(n345),.dout(w_dff_B_4gSGPn0c7_1),.clk(gclk));
	jdff dff_B_PftEIhlQ2_1(.din(w_dff_B_4gSGPn0c7_1),.dout(w_dff_B_PftEIhlQ2_1),.clk(gclk));
	jdff dff_B_4cv6HsYs4_1(.din(w_dff_B_PftEIhlQ2_1),.dout(w_dff_B_4cv6HsYs4_1),.clk(gclk));
	jdff dff_B_HhksMVJk3_1(.din(w_dff_B_4cv6HsYs4_1),.dout(w_dff_B_HhksMVJk3_1),.clk(gclk));
	jdff dff_B_8HdxeRHo2_1(.din(w_dff_B_HhksMVJk3_1),.dout(w_dff_B_8HdxeRHo2_1),.clk(gclk));
	jdff dff_B_tcwanO0x6_1(.din(w_dff_B_8HdxeRHo2_1),.dout(w_dff_B_tcwanO0x6_1),.clk(gclk));
	jdff dff_B_z6Nu5UI97_1(.din(w_dff_B_tcwanO0x6_1),.dout(w_dff_B_z6Nu5UI97_1),.clk(gclk));
	jdff dff_B_TsqBpAWs7_1(.din(w_dff_B_z6Nu5UI97_1),.dout(w_dff_B_TsqBpAWs7_1),.clk(gclk));
	jdff dff_B_h6Hshl8r8_0(.din(n347),.dout(w_dff_B_h6Hshl8r8_0),.clk(gclk));
	jdff dff_B_lnTU46Ef4_0(.din(w_dff_B_h6Hshl8r8_0),.dout(w_dff_B_lnTU46Ef4_0),.clk(gclk));
	jdff dff_B_tCzDTeqT0_0(.din(w_dff_B_lnTU46Ef4_0),.dout(w_dff_B_tCzDTeqT0_0),.clk(gclk));
	jdff dff_B_YUMKxQk66_0(.din(w_dff_B_tCzDTeqT0_0),.dout(w_dff_B_YUMKxQk66_0),.clk(gclk));
	jdff dff_B_6aPnnOYi4_0(.din(w_dff_B_YUMKxQk66_0),.dout(w_dff_B_6aPnnOYi4_0),.clk(gclk));
	jdff dff_B_iYRoJbsl9_0(.din(w_dff_B_6aPnnOYi4_0),.dout(w_dff_B_iYRoJbsl9_0),.clk(gclk));
	jdff dff_B_SOQaeGBi5_0(.din(w_dff_B_iYRoJbsl9_0),.dout(w_dff_B_SOQaeGBi5_0),.clk(gclk));
	jdff dff_B_BpIB3ZO56_0(.din(w_dff_B_SOQaeGBi5_0),.dout(w_dff_B_BpIB3ZO56_0),.clk(gclk));
	jdff dff_B_QebjCnVd4_0(.din(w_dff_B_BpIB3ZO56_0),.dout(w_dff_B_QebjCnVd4_0),.clk(gclk));
	jdff dff_B_LVGe939C6_0(.din(w_dff_B_QebjCnVd4_0),.dout(w_dff_B_LVGe939C6_0),.clk(gclk));
	jdff dff_B_TQD91yn85_0(.din(w_dff_B_LVGe939C6_0),.dout(w_dff_B_TQD91yn85_0),.clk(gclk));
	jdff dff_B_G06qirAy6_0(.din(w_dff_B_TQD91yn85_0),.dout(w_dff_B_G06qirAy6_0),.clk(gclk));
	jdff dff_A_eMp0VwuS4_0(.dout(w_n346_0[0]),.din(w_dff_A_eMp0VwuS4_0),.clk(gclk));
	jdff dff_A_geepDOnh4_0(.dout(w_dff_A_eMp0VwuS4_0),.din(w_dff_A_geepDOnh4_0),.clk(gclk));
	jdff dff_A_B9UNNt9x7_0(.dout(w_dff_A_geepDOnh4_0),.din(w_dff_A_B9UNNt9x7_0),.clk(gclk));
	jdff dff_A_snupMABS2_0(.dout(w_dff_A_B9UNNt9x7_0),.din(w_dff_A_snupMABS2_0),.clk(gclk));
	jdff dff_A_9D0fOy2s0_0(.dout(w_dff_A_snupMABS2_0),.din(w_dff_A_9D0fOy2s0_0),.clk(gclk));
	jdff dff_A_m8HZVMo33_0(.dout(w_dff_A_9D0fOy2s0_0),.din(w_dff_A_m8HZVMo33_0),.clk(gclk));
	jdff dff_A_6Y4fJwgq7_0(.dout(w_dff_A_m8HZVMo33_0),.din(w_dff_A_6Y4fJwgq7_0),.clk(gclk));
	jdff dff_A_F3YcPR6V1_0(.dout(w_dff_A_6Y4fJwgq7_0),.din(w_dff_A_F3YcPR6V1_0),.clk(gclk));
	jdff dff_A_VmV5FVrD4_0(.dout(w_dff_A_F3YcPR6V1_0),.din(w_dff_A_VmV5FVrD4_0),.clk(gclk));
	jdff dff_A_JUVxXoti1_0(.dout(w_dff_A_VmV5FVrD4_0),.din(w_dff_A_JUVxXoti1_0),.clk(gclk));
	jdff dff_A_PhNOj6iL2_0(.dout(w_dff_A_JUVxXoti1_0),.din(w_dff_A_PhNOj6iL2_0),.clk(gclk));
	jdff dff_B_gzcYmuB61_1(.din(n354),.dout(w_dff_B_gzcYmuB61_1),.clk(gclk));
	jdff dff_B_395PlfaZ4_1(.din(w_dff_B_gzcYmuB61_1),.dout(w_dff_B_395PlfaZ4_1),.clk(gclk));
	jdff dff_B_F8Bk1z935_1(.din(w_dff_B_395PlfaZ4_1),.dout(w_dff_B_F8Bk1z935_1),.clk(gclk));
	jdff dff_B_RR7Uxxnl8_1(.din(w_dff_B_F8Bk1z935_1),.dout(w_dff_B_RR7Uxxnl8_1),.clk(gclk));
	jdff dff_B_ZeVdFJOw8_1(.din(w_dff_B_RR7Uxxnl8_1),.dout(w_dff_B_ZeVdFJOw8_1),.clk(gclk));
	jdff dff_B_VX07fHe10_1(.din(w_dff_B_ZeVdFJOw8_1),.dout(w_dff_B_VX07fHe10_1),.clk(gclk));
	jdff dff_B_GfWWVd2B8_1(.din(w_dff_B_VX07fHe10_1),.dout(w_dff_B_GfWWVd2B8_1),.clk(gclk));
	jdff dff_B_0cRPFybT1_1(.din(w_dff_B_GfWWVd2B8_1),.dout(w_dff_B_0cRPFybT1_1),.clk(gclk));
	jdff dff_B_DTXxkQbj7_0(.din(n356),.dout(w_dff_B_DTXxkQbj7_0),.clk(gclk));
	jdff dff_B_1McTIwJt3_0(.din(w_dff_B_DTXxkQbj7_0),.dout(w_dff_B_1McTIwJt3_0),.clk(gclk));
	jdff dff_B_Jw0Z8M1B9_0(.din(w_dff_B_1McTIwJt3_0),.dout(w_dff_B_Jw0Z8M1B9_0),.clk(gclk));
	jdff dff_B_Vz6Vlum58_0(.din(w_dff_B_Jw0Z8M1B9_0),.dout(w_dff_B_Vz6Vlum58_0),.clk(gclk));
	jdff dff_B_dINI8ZUP3_0(.din(w_dff_B_Vz6Vlum58_0),.dout(w_dff_B_dINI8ZUP3_0),.clk(gclk));
	jdff dff_B_Qivm8uCV2_0(.din(w_dff_B_dINI8ZUP3_0),.dout(w_dff_B_Qivm8uCV2_0),.clk(gclk));
	jdff dff_B_eF2q1hLQ7_0(.din(w_dff_B_Qivm8uCV2_0),.dout(w_dff_B_eF2q1hLQ7_0),.clk(gclk));
	jdff dff_B_TY6vQDrg4_0(.din(w_dff_B_eF2q1hLQ7_0),.dout(w_dff_B_TY6vQDrg4_0),.clk(gclk));
	jdff dff_B_PhZkkJJa1_0(.din(w_dff_B_TY6vQDrg4_0),.dout(w_dff_B_PhZkkJJa1_0),.clk(gclk));
	jdff dff_B_NzZ5V3kN8_0(.din(w_dff_B_PhZkkJJa1_0),.dout(w_dff_B_NzZ5V3kN8_0),.clk(gclk));
	jdff dff_B_Wjf4zQ7n9_0(.din(w_dff_B_NzZ5V3kN8_0),.dout(w_dff_B_Wjf4zQ7n9_0),.clk(gclk));
	jdff dff_B_s2kl1zm84_0(.din(w_dff_B_Wjf4zQ7n9_0),.dout(w_dff_B_s2kl1zm84_0),.clk(gclk));
	jdff dff_A_bzQR8LFP0_0(.dout(w_n355_0[0]),.din(w_dff_A_bzQR8LFP0_0),.clk(gclk));
	jdff dff_A_gc8R2JtK2_0(.dout(w_dff_A_bzQR8LFP0_0),.din(w_dff_A_gc8R2JtK2_0),.clk(gclk));
	jdff dff_A_d7zF79lz3_0(.dout(w_dff_A_gc8R2JtK2_0),.din(w_dff_A_d7zF79lz3_0),.clk(gclk));
	jdff dff_A_nQ6aHKOg1_0(.dout(w_dff_A_d7zF79lz3_0),.din(w_dff_A_nQ6aHKOg1_0),.clk(gclk));
	jdff dff_A_dm8tWFpL6_0(.dout(w_dff_A_nQ6aHKOg1_0),.din(w_dff_A_dm8tWFpL6_0),.clk(gclk));
	jdff dff_A_umN1t3SI3_0(.dout(w_dff_A_dm8tWFpL6_0),.din(w_dff_A_umN1t3SI3_0),.clk(gclk));
	jdff dff_A_6Wfwcwbb4_0(.dout(w_dff_A_umN1t3SI3_0),.din(w_dff_A_6Wfwcwbb4_0),.clk(gclk));
	jdff dff_A_fxG2Bkiq3_0(.dout(w_dff_A_6Wfwcwbb4_0),.din(w_dff_A_fxG2Bkiq3_0),.clk(gclk));
	jdff dff_A_22BpD5M60_0(.dout(w_dff_A_fxG2Bkiq3_0),.din(w_dff_A_22BpD5M60_0),.clk(gclk));
	jdff dff_A_imeOIfBC3_0(.dout(w_dff_A_22BpD5M60_0),.din(w_dff_A_imeOIfBC3_0),.clk(gclk));
	jdff dff_A_Wi2sX6WX9_0(.dout(w_dff_A_imeOIfBC3_0),.din(w_dff_A_Wi2sX6WX9_0),.clk(gclk));
	jdff dff_B_0A5AnHRJ6_1(.din(n363),.dout(w_dff_B_0A5AnHRJ6_1),.clk(gclk));
	jdff dff_B_IWOnRHmV8_1(.din(w_dff_B_0A5AnHRJ6_1),.dout(w_dff_B_IWOnRHmV8_1),.clk(gclk));
	jdff dff_B_vd7RZRZQ4_1(.din(w_dff_B_IWOnRHmV8_1),.dout(w_dff_B_vd7RZRZQ4_1),.clk(gclk));
	jdff dff_B_1teWePyF9_1(.din(w_dff_B_vd7RZRZQ4_1),.dout(w_dff_B_1teWePyF9_1),.clk(gclk));
	jdff dff_B_si90QFER0_1(.din(w_dff_B_1teWePyF9_1),.dout(w_dff_B_si90QFER0_1),.clk(gclk));
	jdff dff_B_icu8dmV40_1(.din(w_dff_B_si90QFER0_1),.dout(w_dff_B_icu8dmV40_1),.clk(gclk));
	jdff dff_B_Q4gWqjTo5_1(.din(w_dff_B_icu8dmV40_1),.dout(w_dff_B_Q4gWqjTo5_1),.clk(gclk));
	jdff dff_B_GUcOIG9m7_1(.din(w_dff_B_Q4gWqjTo5_1),.dout(w_dff_B_GUcOIG9m7_1),.clk(gclk));
	jdff dff_B_evOaY06v4_0(.din(n365),.dout(w_dff_B_evOaY06v4_0),.clk(gclk));
	jdff dff_B_KlX3RWNc3_0(.din(w_dff_B_evOaY06v4_0),.dout(w_dff_B_KlX3RWNc3_0),.clk(gclk));
	jdff dff_B_cW3URVOS0_0(.din(w_dff_B_KlX3RWNc3_0),.dout(w_dff_B_cW3URVOS0_0),.clk(gclk));
	jdff dff_B_tbqvdAG68_0(.din(w_dff_B_cW3URVOS0_0),.dout(w_dff_B_tbqvdAG68_0),.clk(gclk));
	jdff dff_B_r836DeSm9_0(.din(w_dff_B_tbqvdAG68_0),.dout(w_dff_B_r836DeSm9_0),.clk(gclk));
	jdff dff_B_YnFkwijJ8_0(.din(w_dff_B_r836DeSm9_0),.dout(w_dff_B_YnFkwijJ8_0),.clk(gclk));
	jdff dff_B_23WNmQWq8_0(.din(w_dff_B_YnFkwijJ8_0),.dout(w_dff_B_23WNmQWq8_0),.clk(gclk));
	jdff dff_B_kZOWN7u47_0(.din(w_dff_B_23WNmQWq8_0),.dout(w_dff_B_kZOWN7u47_0),.clk(gclk));
	jdff dff_B_S7jUhja64_0(.din(w_dff_B_kZOWN7u47_0),.dout(w_dff_B_S7jUhja64_0),.clk(gclk));
	jdff dff_B_bubJ0FPE4_0(.din(w_dff_B_S7jUhja64_0),.dout(w_dff_B_bubJ0FPE4_0),.clk(gclk));
	jdff dff_B_jC8nVPTV4_0(.din(w_dff_B_bubJ0FPE4_0),.dout(w_dff_B_jC8nVPTV4_0),.clk(gclk));
	jdff dff_B_iVxIWCT72_0(.din(w_dff_B_jC8nVPTV4_0),.dout(w_dff_B_iVxIWCT72_0),.clk(gclk));
	jdff dff_A_7tlowIyn2_0(.dout(w_n364_0[0]),.din(w_dff_A_7tlowIyn2_0),.clk(gclk));
	jdff dff_A_zHbC0nEr4_0(.dout(w_dff_A_7tlowIyn2_0),.din(w_dff_A_zHbC0nEr4_0),.clk(gclk));
	jdff dff_A_3E0vZNI53_0(.dout(w_dff_A_zHbC0nEr4_0),.din(w_dff_A_3E0vZNI53_0),.clk(gclk));
	jdff dff_A_NkVginFn0_0(.dout(w_dff_A_3E0vZNI53_0),.din(w_dff_A_NkVginFn0_0),.clk(gclk));
	jdff dff_A_xkvxwhXk6_0(.dout(w_dff_A_NkVginFn0_0),.din(w_dff_A_xkvxwhXk6_0),.clk(gclk));
	jdff dff_A_RmdZkWv63_0(.dout(w_dff_A_xkvxwhXk6_0),.din(w_dff_A_RmdZkWv63_0),.clk(gclk));
	jdff dff_A_hooEpd6B0_0(.dout(w_dff_A_RmdZkWv63_0),.din(w_dff_A_hooEpd6B0_0),.clk(gclk));
	jdff dff_A_VATPqFss2_0(.dout(w_dff_A_hooEpd6B0_0),.din(w_dff_A_VATPqFss2_0),.clk(gclk));
	jdff dff_A_CdbqV4wH7_0(.dout(w_dff_A_VATPqFss2_0),.din(w_dff_A_CdbqV4wH7_0),.clk(gclk));
	jdff dff_A_oB3bxZdb5_0(.dout(w_dff_A_CdbqV4wH7_0),.din(w_dff_A_oB3bxZdb5_0),.clk(gclk));
	jdff dff_A_I6BHAfxa8_0(.dout(w_dff_A_oB3bxZdb5_0),.din(w_dff_A_I6BHAfxa8_0),.clk(gclk));
	jdff dff_B_zKKZ3OEc9_1(.din(n374),.dout(w_dff_B_zKKZ3OEc9_1),.clk(gclk));
	jdff dff_B_MgoIaZ0d6_1(.din(w_dff_B_zKKZ3OEc9_1),.dout(w_dff_B_MgoIaZ0d6_1),.clk(gclk));
	jdff dff_B_rQ3APO7a0_0(.din(n375),.dout(w_dff_B_rQ3APO7a0_0),.clk(gclk));
	jdff dff_B_2Vc9FAdH3_0(.din(w_dff_B_rQ3APO7a0_0),.dout(w_dff_B_2Vc9FAdH3_0),.clk(gclk));
	jdff dff_B_dIHTQlUc5_0(.din(w_dff_B_2Vc9FAdH3_0),.dout(w_dff_B_dIHTQlUc5_0),.clk(gclk));
	jdff dff_B_pMAnzE9l5_0(.din(w_dff_B_dIHTQlUc5_0),.dout(w_dff_B_pMAnzE9l5_0),.clk(gclk));
	jdff dff_B_ZNW43P2h7_0(.din(w_dff_B_pMAnzE9l5_0),.dout(w_dff_B_ZNW43P2h7_0),.clk(gclk));
	jdff dff_B_8dkfrdX51_0(.din(w_dff_B_ZNW43P2h7_0),.dout(w_dff_B_8dkfrdX51_0),.clk(gclk));
	jdff dff_B_wSvcQ8VG9_0(.din(w_dff_B_8dkfrdX51_0),.dout(w_dff_B_wSvcQ8VG9_0),.clk(gclk));
	jdff dff_B_n5BItyIC8_0(.din(w_dff_B_wSvcQ8VG9_0),.dout(w_dff_B_n5BItyIC8_0),.clk(gclk));
	jdff dff_B_knUKdgrF7_0(.din(w_dff_B_n5BItyIC8_0),.dout(w_dff_B_knUKdgrF7_0),.clk(gclk));
	jdff dff_B_jTCA9YDL5_0(.din(w_dff_B_knUKdgrF7_0),.dout(w_dff_B_jTCA9YDL5_0),.clk(gclk));
	jdff dff_B_NcuqmW5k8_0(.din(w_dff_B_jTCA9YDL5_0),.dout(w_dff_B_NcuqmW5k8_0),.clk(gclk));
	jdff dff_B_2KeNDtYV1_0(.din(w_dff_B_NcuqmW5k8_0),.dout(w_dff_B_2KeNDtYV1_0),.clk(gclk));
	jdff dff_A_rHrGhwGm6_0(.dout(w_n340_1[0]),.din(w_dff_A_rHrGhwGm6_0),.clk(gclk));
	jdff dff_A_VtiVWISb2_1(.dout(w_n372_0[1]),.din(w_dff_A_VtiVWISb2_1),.clk(gclk));
	jdff dff_A_SjSFDZ172_1(.dout(w_dff_A_VtiVWISb2_1),.din(w_dff_A_SjSFDZ172_1),.clk(gclk));
	jdff dff_A_HnDKh3SD2_1(.dout(w_dff_A_SjSFDZ172_1),.din(w_dff_A_HnDKh3SD2_1),.clk(gclk));
	jdff dff_A_LVohhpl28_1(.dout(w_dff_A_HnDKh3SD2_1),.din(w_dff_A_LVohhpl28_1),.clk(gclk));
	jdff dff_A_jotmuWdv7_1(.dout(w_dff_A_LVohhpl28_1),.din(w_dff_A_jotmuWdv7_1),.clk(gclk));
	jdff dff_A_NwbRj9zl4_1(.dout(w_dff_A_jotmuWdv7_1),.din(w_dff_A_NwbRj9zl4_1),.clk(gclk));
	jdff dff_A_RkMChSBt7_1(.dout(w_dff_A_NwbRj9zl4_1),.din(w_dff_A_RkMChSBt7_1),.clk(gclk));
	jdff dff_A_aTKAHHWz1_1(.dout(w_dff_A_RkMChSBt7_1),.din(w_dff_A_aTKAHHWz1_1),.clk(gclk));
	jdff dff_A_UxttpmSE7_1(.dout(w_dff_A_aTKAHHWz1_1),.din(w_dff_A_UxttpmSE7_1),.clk(gclk));
	jdff dff_A_b4AgwyJ03_1(.dout(w_dff_A_UxttpmSE7_1),.din(w_dff_A_b4AgwyJ03_1),.clk(gclk));
	jdff dff_A_TL2yhSof4_1(.dout(w_dff_A_b4AgwyJ03_1),.din(w_dff_A_TL2yhSof4_1),.clk(gclk));
	jdff dff_B_X55qSwQ59_1(.din(n380),.dout(w_dff_B_X55qSwQ59_1),.clk(gclk));
	jdff dff_B_6i9ei40a9_1(.din(w_dff_B_X55qSwQ59_1),.dout(w_dff_B_6i9ei40a9_1),.clk(gclk));
	jdff dff_B_BE0wj4rv4_1(.din(w_dff_B_6i9ei40a9_1),.dout(w_dff_B_BE0wj4rv4_1),.clk(gclk));
	jdff dff_B_UnDnEvbz5_1(.din(w_dff_B_BE0wj4rv4_1),.dout(w_dff_B_UnDnEvbz5_1),.clk(gclk));
	jdff dff_B_65ZOrPmx6_1(.din(w_dff_B_UnDnEvbz5_1),.dout(w_dff_B_65ZOrPmx6_1),.clk(gclk));
	jdff dff_B_FQDpFeNo3_1(.din(w_dff_B_65ZOrPmx6_1),.dout(w_dff_B_FQDpFeNo3_1),.clk(gclk));
	jdff dff_B_nA4SKkqB7_1(.din(w_dff_B_FQDpFeNo3_1),.dout(w_dff_B_nA4SKkqB7_1),.clk(gclk));
	jdff dff_B_DIgbkSqt5_1(.din(w_dff_B_nA4SKkqB7_1),.dout(w_dff_B_DIgbkSqt5_1),.clk(gclk));
	jdff dff_B_yLSdhCZv3_1(.din(w_dff_B_DIgbkSqt5_1),.dout(w_dff_B_yLSdhCZv3_1),.clk(gclk));
	jdff dff_B_h1QunbAe8_1(.din(w_dff_B_yLSdhCZv3_1),.dout(w_dff_B_h1QunbAe8_1),.clk(gclk));
	jdff dff_B_EtETzIiC2_1(.din(w_dff_B_h1QunbAe8_1),.dout(w_dff_B_EtETzIiC2_1),.clk(gclk));
	jdff dff_B_3U02k0zt1_1(.din(w_dff_B_EtETzIiC2_1),.dout(w_dff_B_3U02k0zt1_1),.clk(gclk));
	jdff dff_B_FpHpHvB37_1(.din(w_dff_B_3U02k0zt1_1),.dout(w_dff_B_FpHpHvB37_1),.clk(gclk));
	jdff dff_B_29L0AqtW3_0(.din(n382),.dout(w_dff_B_29L0AqtW3_0),.clk(gclk));
	jdff dff_B_f1rGZROM0_0(.din(w_dff_B_29L0AqtW3_0),.dout(w_dff_B_f1rGZROM0_0),.clk(gclk));
	jdff dff_B_CXPGAOjp9_0(.din(w_dff_B_f1rGZROM0_0),.dout(w_dff_B_CXPGAOjp9_0),.clk(gclk));
	jdff dff_B_x6buodD33_0(.din(w_dff_B_CXPGAOjp9_0),.dout(w_dff_B_x6buodD33_0),.clk(gclk));
	jdff dff_B_m7Ig0zAD1_0(.din(w_dff_B_x6buodD33_0),.dout(w_dff_B_m7Ig0zAD1_0),.clk(gclk));
	jdff dff_B_lOepdcUX9_0(.din(w_dff_B_m7Ig0zAD1_0),.dout(w_dff_B_lOepdcUX9_0),.clk(gclk));
	jdff dff_B_czWIJref1_0(.din(w_dff_B_lOepdcUX9_0),.dout(w_dff_B_czWIJref1_0),.clk(gclk));
	jdff dff_B_gcUtwAsh1_0(.din(w_dff_B_czWIJref1_0),.dout(w_dff_B_gcUtwAsh1_0),.clk(gclk));
	jdff dff_B_mbzieB0G6_0(.din(w_dff_B_gcUtwAsh1_0),.dout(w_dff_B_mbzieB0G6_0),.clk(gclk));
	jdff dff_B_QZkuKSeL6_0(.din(w_dff_B_mbzieB0G6_0),.dout(w_dff_B_QZkuKSeL6_0),.clk(gclk));
	jdff dff_B_4UcDNbX05_0(.din(w_dff_B_QZkuKSeL6_0),.dout(w_dff_B_4UcDNbX05_0),.clk(gclk));
	jdff dff_B_h3nV6xkx4_0(.din(w_dff_B_4UcDNbX05_0),.dout(w_dff_B_h3nV6xkx4_0),.clk(gclk));
	jdff dff_B_kxufNpK89_0(.din(n392),.dout(w_dff_B_kxufNpK89_0),.clk(gclk));
	jdff dff_B_BcqZbD243_0(.din(w_dff_B_kxufNpK89_0),.dout(w_dff_B_BcqZbD243_0),.clk(gclk));
	jdff dff_B_HE0CuCCN0_0(.din(w_dff_B_BcqZbD243_0),.dout(w_dff_B_HE0CuCCN0_0),.clk(gclk));
	jdff dff_B_gssPliqy2_0(.din(w_dff_B_HE0CuCCN0_0),.dout(w_dff_B_gssPliqy2_0),.clk(gclk));
	jdff dff_B_J7xJxTDd6_0(.din(w_dff_B_gssPliqy2_0),.dout(w_dff_B_J7xJxTDd6_0),.clk(gclk));
	jdff dff_B_vzeYRoUh1_0(.din(w_dff_B_J7xJxTDd6_0),.dout(w_dff_B_vzeYRoUh1_0),.clk(gclk));
	jdff dff_B_Crwz3Alx7_0(.din(w_dff_B_vzeYRoUh1_0),.dout(w_dff_B_Crwz3Alx7_0),.clk(gclk));
	jdff dff_B_WVAZna0S0_0(.din(w_dff_B_Crwz3Alx7_0),.dout(w_dff_B_WVAZna0S0_0),.clk(gclk));
	jdff dff_B_61pLk6yF7_0(.din(w_dff_B_WVAZna0S0_0),.dout(w_dff_B_61pLk6yF7_0),.clk(gclk));
	jdff dff_B_PdPedVg21_1(.din(n390),.dout(w_dff_B_PdPedVg21_1),.clk(gclk));
	jdff dff_B_suVRAECO2_1(.din(w_dff_B_PdPedVg21_1),.dout(w_dff_B_suVRAECO2_1),.clk(gclk));
	jdff dff_B_022ZCcFP7_1(.din(w_dff_B_suVRAECO2_1),.dout(w_dff_B_022ZCcFP7_1),.clk(gclk));
	jdff dff_B_dBRpNvDI0_0(.din(n388),.dout(w_dff_B_dBRpNvDI0_0),.clk(gclk));
	jdff dff_B_VVOSGF3B5_0(.din(w_dff_B_dBRpNvDI0_0),.dout(w_dff_B_VVOSGF3B5_0),.clk(gclk));
	jdff dff_B_VFhQmT8V3_0(.din(w_dff_B_VVOSGF3B5_0),.dout(w_dff_B_VFhQmT8V3_0),.clk(gclk));
	jdff dff_B_Gn09emKO0_0(.din(w_dff_B_VFhQmT8V3_0),.dout(w_dff_B_Gn09emKO0_0),.clk(gclk));
	jdff dff_B_ImpSVUN95_0(.din(w_dff_B_Gn09emKO0_0),.dout(w_dff_B_ImpSVUN95_0),.clk(gclk));
	jdff dff_B_v0Qnln3h1_0(.din(w_dff_B_ImpSVUN95_0),.dout(w_dff_B_v0Qnln3h1_0),.clk(gclk));
	jdff dff_B_8vxcRGM88_0(.din(w_dff_B_v0Qnln3h1_0),.dout(w_dff_B_8vxcRGM88_0),.clk(gclk));
	jdff dff_B_vSf3deVJ8_0(.din(w_dff_B_8vxcRGM88_0),.dout(w_dff_B_vSf3deVJ8_0),.clk(gclk));
	jdff dff_B_ox8kK8oC3_0(.din(w_dff_B_vSf3deVJ8_0),.dout(w_dff_B_ox8kK8oC3_0),.clk(gclk));
	jdff dff_B_OCWgBTbT0_0(.din(w_dff_B_ox8kK8oC3_0),.dout(w_dff_B_OCWgBTbT0_0),.clk(gclk));
	jdff dff_B_QcpHiPlY3_0(.din(w_dff_B_OCWgBTbT0_0),.dout(w_dff_B_QcpHiPlY3_0),.clk(gclk));
	jdff dff_B_y5Ms6zHM2_0(.din(n224),.dout(w_dff_B_y5Ms6zHM2_0),.clk(gclk));
	jdff dff_A_TTLwkGB22_0(.dout(w_n190_0[0]),.din(w_dff_A_TTLwkGB22_0),.clk(gclk));
	jdff dff_A_kenMqaJC9_0(.dout(w_n222_0[0]),.din(w_dff_A_kenMqaJC9_0),.clk(gclk));
	jdff dff_A_o6iHd4wS5_0(.dout(w_n220_0[0]),.din(w_dff_A_o6iHd4wS5_0),.clk(gclk));
	jdff dff_A_GfqyIOPq1_0(.dout(w_n218_1[0]),.din(w_dff_A_GfqyIOPq1_0),.clk(gclk));
	jdff dff_A_PGts8FVS1_0(.dout(w_dff_A_GfqyIOPq1_0),.din(w_dff_A_PGts8FVS1_0),.clk(gclk));
	jdff dff_A_1wJHQT8i1_2(.dout(w_n218_0[2]),.din(w_dff_A_1wJHQT8i1_2),.clk(gclk));
	jdff dff_A_LcBlZ9aX5_2(.dout(w_dff_A_1wJHQT8i1_2),.din(w_dff_A_LcBlZ9aX5_2),.clk(gclk));
	jdff dff_A_Fa2UMt9f5_2(.dout(w_n192_0[2]),.din(w_dff_A_Fa2UMt9f5_2),.clk(gclk));
	jdff dff_B_axGrS3Iv1_3(.din(n192),.dout(w_dff_B_axGrS3Iv1_3),.clk(gclk));
	jdff dff_B_nI5fi7wz8_0(.din(n234),.dout(w_dff_B_nI5fi7wz8_0),.clk(gclk));
	jdff dff_A_8rWjRxp07_0(.dout(w_n156_0[0]),.din(w_dff_A_8rWjRxp07_0),.clk(gclk));
	jdff dff_B_dSziAO2Z1_0(.din(n231),.dout(w_dff_B_dSziAO2Z1_0),.clk(gclk));
	jdff dff_A_BNL5dXN84_0(.dout(w_n198_1[0]),.din(w_dff_A_BNL5dXN84_0),.clk(gclk));
	jdff dff_A_prYlLrbr6_2(.dout(w_n198_0[2]),.din(w_dff_A_prYlLrbr6_2),.clk(gclk));
	jdff dff_A_2B8NSCZf5_2(.dout(w_dff_A_prYlLrbr6_2),.din(w_dff_A_2B8NSCZf5_2),.clk(gclk));
	jdff dff_A_Vd29EL2O1_0(.dout(w_n197_1[0]),.din(w_dff_A_Vd29EL2O1_0),.clk(gclk));
	jdff dff_A_dA8Bc4bg1_0(.dout(w_n155_0[0]),.din(w_dff_A_dA8Bc4bg1_0),.clk(gclk));
	jdff dff_B_7SPTAqeQ4_3(.din(n155),.dout(w_dff_B_7SPTAqeQ4_3),.clk(gclk));
	jdff dff_A_7t150ZsV1_0(.dout(w_n144_1[0]),.din(w_dff_A_7t150ZsV1_0),.clk(gclk));
	jdff dff_A_1wrvM3uX4_1(.dout(w_n144_0[1]),.din(w_dff_A_1wrvM3uX4_1),.clk(gclk));
	jdff dff_A_YONZmBkR0_0(.dout(w_n169_0[0]),.din(w_dff_A_YONZmBkR0_0),.clk(gclk));
	jdff dff_A_zs3zT8BU7_2(.dout(w_n159_0[2]),.din(w_dff_A_zs3zT8BU7_2),.clk(gclk));
	jdff dff_A_8YxqbqHk9_0(.dout(w_n158_1[0]),.din(w_dff_A_8YxqbqHk9_0),.clk(gclk));
	jdff dff_A_3qPQklFW8_1(.dout(w_n121_0[1]),.din(w_dff_A_3qPQklFW8_1),.clk(gclk));
	jdff dff_A_3cSJ8hMY5_2(.dout(w_n121_0[2]),.din(w_dff_A_3cSJ8hMY5_2),.clk(gclk));
	jdff dff_A_pod2XMWh3_2(.dout(w_dff_A_3cSJ8hMY5_2),.din(w_dff_A_pod2XMWh3_2),.clk(gclk));
	jdff dff_A_STNXeMv85_1(.dout(w_n96_0[1]),.din(w_dff_A_STNXeMv85_1),.clk(gclk));
	jdff dff_A_QYAUMjpJ2_1(.dout(w_dff_A_STNXeMv85_1),.din(w_dff_A_QYAUMjpJ2_1),.clk(gclk));
	jdff dff_A_G1aJbt6l0_1(.dout(w_dff_A_QYAUMjpJ2_1),.din(w_dff_A_G1aJbt6l0_1),.clk(gclk));
	jdff dff_A_WtZesN640_1(.dout(w_dff_A_G1aJbt6l0_1),.din(w_dff_A_WtZesN640_1),.clk(gclk));
	jdff dff_A_e2uwbNNi9_1(.dout(w_dff_A_WtZesN640_1),.din(w_dff_A_e2uwbNNi9_1),.clk(gclk));
	jdff dff_A_3PBly9OT4_2(.dout(w_n96_0[2]),.din(w_dff_A_3PBly9OT4_2),.clk(gclk));
	jdff dff_A_SKE5l9Sv3_2(.dout(w_dff_A_3PBly9OT4_2),.din(w_dff_A_SKE5l9Sv3_2),.clk(gclk));
	jdff dff_A_P22dRqlb4_2(.dout(w_dff_A_SKE5l9Sv3_2),.din(w_dff_A_P22dRqlb4_2),.clk(gclk));
	jdff dff_A_5Xc59Xal7_2(.dout(w_dff_A_P22dRqlb4_2),.din(w_dff_A_5Xc59Xal7_2),.clk(gclk));
	jdff dff_A_HQSc0RKe9_2(.dout(w_dff_A_5Xc59Xal7_2),.din(w_dff_A_HQSc0RKe9_2),.clk(gclk));
	jdff dff_B_o5OKE4Qy5_3(.din(n340),.dout(w_dff_B_o5OKE4Qy5_3),.clk(gclk));
	jdff dff_B_cNBx2DoW7_3(.din(w_dff_B_o5OKE4Qy5_3),.dout(w_dff_B_cNBx2DoW7_3),.clk(gclk));
	jdff dff_B_YudUmxXw9_3(.din(w_dff_B_cNBx2DoW7_3),.dout(w_dff_B_YudUmxXw9_3),.clk(gclk));
	jdff dff_B_Fb0mb4rz9_3(.din(w_dff_B_YudUmxXw9_3),.dout(w_dff_B_Fb0mb4rz9_3),.clk(gclk));
	jdff dff_B_IQIZtJwg9_3(.din(w_dff_B_Fb0mb4rz9_3),.dout(w_dff_B_IQIZtJwg9_3),.clk(gclk));
	jdff dff_B_cT0aTmBS3_3(.din(w_dff_B_IQIZtJwg9_3),.dout(w_dff_B_cT0aTmBS3_3),.clk(gclk));
	jdff dff_B_H5glYabS3_3(.din(w_dff_B_cT0aTmBS3_3),.dout(w_dff_B_H5glYabS3_3),.clk(gclk));
	jdff dff_B_gIQ4yZ628_3(.din(w_dff_B_H5glYabS3_3),.dout(w_dff_B_gIQ4yZ628_3),.clk(gclk));
	jdff dff_B_ijbgwGBd3_3(.din(w_dff_B_gIQ4yZ628_3),.dout(w_dff_B_ijbgwGBd3_3),.clk(gclk));
	jdff dff_B_hmP7Xgvq0_3(.din(w_dff_B_ijbgwGBd3_3),.dout(w_dff_B_hmP7Xgvq0_3),.clk(gclk));
	jdff dff_B_SAdMQ8W21_3(.din(w_dff_B_hmP7Xgvq0_3),.dout(w_dff_B_SAdMQ8W21_3),.clk(gclk));
	jdff dff_B_mOt15Rct5_3(.din(w_dff_B_SAdMQ8W21_3),.dout(w_dff_B_mOt15Rct5_3),.clk(gclk));
	jdff dff_B_yh0Ff1q94_1(.din(n394),.dout(w_dff_B_yh0Ff1q94_1),.clk(gclk));
	jdff dff_B_tEU1EZhI4_1(.din(w_dff_B_yh0Ff1q94_1),.dout(w_dff_B_tEU1EZhI4_1),.clk(gclk));
	jdff dff_B_uQkA5nfM7_1(.din(w_dff_B_tEU1EZhI4_1),.dout(w_dff_B_uQkA5nfM7_1),.clk(gclk));
	jdff dff_B_TsgPsMYj5_1(.din(w_dff_B_uQkA5nfM7_1),.dout(w_dff_B_TsgPsMYj5_1),.clk(gclk));
	jdff dff_B_msmgJLvC1_1(.din(w_dff_B_TsgPsMYj5_1),.dout(w_dff_B_msmgJLvC1_1),.clk(gclk));
	jdff dff_B_c6CCa8PK5_1(.din(w_dff_B_msmgJLvC1_1),.dout(w_dff_B_c6CCa8PK5_1),.clk(gclk));
	jdff dff_B_dqsrEPo56_1(.din(w_dff_B_c6CCa8PK5_1),.dout(w_dff_B_dqsrEPo56_1),.clk(gclk));
	jdff dff_B_Czv2JzUB9_1(.din(w_dff_B_dqsrEPo56_1),.dout(w_dff_B_Czv2JzUB9_1),.clk(gclk));
	jdff dff_B_sqnk2SLN1_0(.din(n396),.dout(w_dff_B_sqnk2SLN1_0),.clk(gclk));
	jdff dff_B_Rzr8Ywb19_0(.din(w_dff_B_sqnk2SLN1_0),.dout(w_dff_B_Rzr8Ywb19_0),.clk(gclk));
	jdff dff_B_DxmhlZKD5_0(.din(w_dff_B_Rzr8Ywb19_0),.dout(w_dff_B_DxmhlZKD5_0),.clk(gclk));
	jdff dff_B_ODSuntNp6_0(.din(w_dff_B_DxmhlZKD5_0),.dout(w_dff_B_ODSuntNp6_0),.clk(gclk));
	jdff dff_B_SBkrtyXU0_0(.din(w_dff_B_ODSuntNp6_0),.dout(w_dff_B_SBkrtyXU0_0),.clk(gclk));
	jdff dff_B_onb1ImyF2_0(.din(w_dff_B_SBkrtyXU0_0),.dout(w_dff_B_onb1ImyF2_0),.clk(gclk));
	jdff dff_B_a6crvk4w2_0(.din(w_dff_B_onb1ImyF2_0),.dout(w_dff_B_a6crvk4w2_0),.clk(gclk));
	jdff dff_B_pNSd7VtP8_0(.din(w_dff_B_a6crvk4w2_0),.dout(w_dff_B_pNSd7VtP8_0),.clk(gclk));
	jdff dff_B_kR6XVgw99_0(.din(w_dff_B_pNSd7VtP8_0),.dout(w_dff_B_kR6XVgw99_0),.clk(gclk));
	jdff dff_B_k8RBcNYk9_0(.din(w_dff_B_kR6XVgw99_0),.dout(w_dff_B_k8RBcNYk9_0),.clk(gclk));
	jdff dff_B_fA13W3LH0_0(.din(w_dff_B_k8RBcNYk9_0),.dout(w_dff_B_fA13W3LH0_0),.clk(gclk));
	jdff dff_B_AjK9z4Zd6_0(.din(w_dff_B_fA13W3LH0_0),.dout(w_dff_B_AjK9z4Zd6_0),.clk(gclk));
	jdff dff_A_QW8XngQV8_0(.dout(w_n395_0[0]),.din(w_dff_A_QW8XngQV8_0),.clk(gclk));
	jdff dff_A_lMNyvMra4_0(.dout(w_dff_A_QW8XngQV8_0),.din(w_dff_A_lMNyvMra4_0),.clk(gclk));
	jdff dff_A_z1un55ZR9_0(.dout(w_dff_A_lMNyvMra4_0),.din(w_dff_A_z1un55ZR9_0),.clk(gclk));
	jdff dff_A_ENPr6b0i8_0(.dout(w_dff_A_z1un55ZR9_0),.din(w_dff_A_ENPr6b0i8_0),.clk(gclk));
	jdff dff_A_o4kweXGV0_0(.dout(w_dff_A_ENPr6b0i8_0),.din(w_dff_A_o4kweXGV0_0),.clk(gclk));
	jdff dff_A_5pDU0vH70_0(.dout(w_dff_A_o4kweXGV0_0),.din(w_dff_A_5pDU0vH70_0),.clk(gclk));
	jdff dff_A_3bvbr5rV8_0(.dout(w_dff_A_5pDU0vH70_0),.din(w_dff_A_3bvbr5rV8_0),.clk(gclk));
	jdff dff_A_gGaJ42v52_0(.dout(w_dff_A_3bvbr5rV8_0),.din(w_dff_A_gGaJ42v52_0),.clk(gclk));
	jdff dff_A_y7tY9tcx0_0(.dout(w_dff_A_gGaJ42v52_0),.din(w_dff_A_y7tY9tcx0_0),.clk(gclk));
	jdff dff_A_s8mRo0vA3_0(.dout(w_dff_A_y7tY9tcx0_0),.din(w_dff_A_s8mRo0vA3_0),.clk(gclk));
	jdff dff_A_CTbbxFKx9_0(.dout(w_dff_A_s8mRo0vA3_0),.din(w_dff_A_CTbbxFKx9_0),.clk(gclk));
	jdff dff_B_4Ceh4tJ99_0(.din(n332),.dout(w_dff_B_4Ceh4tJ99_0),.clk(gclk));
	jdff dff_B_UCJLGiV16_0(.din(w_dff_B_4Ceh4tJ99_0),.dout(w_dff_B_UCJLGiV16_0),.clk(gclk));
	jdff dff_B_SoUsOi0K6_0(.din(n329),.dout(w_dff_B_SoUsOi0K6_0),.clk(gclk));
	jdff dff_B_dRAP4BFq1_0(.din(n326),.dout(w_dff_B_dRAP4BFq1_0),.clk(gclk));
	jdff dff_B_u1v0oDzC5_0(.din(w_dff_B_dRAP4BFq1_0),.dout(w_dff_B_u1v0oDzC5_0),.clk(gclk));
	jdff dff_A_Co56wZdW7_1(.dout(w_n189_0[1]),.din(w_dff_A_Co56wZdW7_1),.clk(gclk));
	jdff dff_B_syV6dGNo7_1(.din(n317),.dout(w_dff_B_syV6dGNo7_1),.clk(gclk));
	jdff dff_A_1OKfejET8_1(.dout(w_n185_0[1]),.din(w_dff_A_1OKfejET8_1),.clk(gclk));
	jdff dff_A_KJgL8d3N4_2(.dout(w_n185_0[2]),.din(w_dff_A_KJgL8d3N4_2),.clk(gclk));
	jdff dff_A_0Epgjh5R4_2(.dout(w_dff_A_KJgL8d3N4_2),.din(w_dff_A_0Epgjh5R4_2),.clk(gclk));
	jdff dff_B_9C0m26qy5_3(.din(n184),.dout(w_dff_B_9C0m26qy5_3),.clk(gclk));
	jdff dff_B_01Sj3U7Z8_3(.din(w_dff_B_9C0m26qy5_3),.dout(w_dff_B_01Sj3U7Z8_3),.clk(gclk));
	jdff dff_B_KxqXcm3f6_1(.din(n312),.dout(w_dff_B_KxqXcm3f6_1),.clk(gclk));
	jdff dff_A_ytS0m6ve3_0(.dout(w_n315_0[0]),.din(w_dff_A_ytS0m6ve3_0),.clk(gclk));
	jdff dff_A_1QG9NFcn5_2(.dout(w_n314_0[2]),.din(w_dff_A_1QG9NFcn5_2),.clk(gclk));
	jdff dff_B_YxBQv0KS6_3(.din(n314),.dout(w_dff_B_YxBQv0KS6_3),.clk(gclk));
	jdff dff_A_WliHaTzo1_1(.dout(w_n311_0[1]),.din(w_dff_A_WliHaTzo1_1),.clk(gclk));
	jdff dff_B_Hc8yxGjE5_3(.din(n311),.dout(w_dff_B_Hc8yxGjE5_3),.clk(gclk));
	jdff dff_A_AYIUsmw50_0(.dout(w_n183_0[0]),.din(w_dff_A_AYIUsmw50_0),.clk(gclk));
	jdff dff_A_3t72QqKb7_0(.dout(w_dff_A_AYIUsmw50_0),.din(w_dff_A_3t72QqKb7_0),.clk(gclk));
	jdff dff_A_inl9Q56b6_1(.dout(w_n183_0[1]),.din(w_dff_A_inl9Q56b6_1),.clk(gclk));
	jdff dff_A_vPrrgWUx2_1(.dout(w_dff_A_inl9Q56b6_1),.din(w_dff_A_vPrrgWUx2_1),.clk(gclk));
	jdff dff_B_xaq43RIw5_0(.din(n182),.dout(w_dff_B_xaq43RIw5_0),.clk(gclk));
	jdff dff_B_acby1dGc9_0(.din(w_dff_B_xaq43RIw5_0),.dout(w_dff_B_acby1dGc9_0),.clk(gclk));
	jdff dff_B_jMQCyKhi9_0(.din(w_dff_B_acby1dGc9_0),.dout(w_dff_B_jMQCyKhi9_0),.clk(gclk));
	jdff dff_B_vdJpMGfu1_1(.din(G900),.dout(w_dff_B_vdJpMGfu1_1),.clk(gclk));
	jdff dff_A_fQQWn7ir4_0(.dout(w_n309_0[0]),.din(w_dff_A_fQQWn7ir4_0),.clk(gclk));
	jdff dff_A_GFsw4uTu9_0(.dout(w_dff_A_fQQWn7ir4_0),.din(w_dff_A_GFsw4uTu9_0),.clk(gclk));
	jdff dff_B_IzJsr9a93_1(.din(n299),.dout(w_dff_B_IzJsr9a93_1),.clk(gclk));
	jdff dff_B_Jkj5CeEG9_0(.din(n305),.dout(w_dff_B_Jkj5CeEG9_0),.clk(gclk));
	jdff dff_B_AypWXcsc5_0(.din(n303),.dout(w_dff_B_AypWXcsc5_0),.clk(gclk));
	jdff dff_B_nlL1oXQa2_0(.din(w_dff_B_AypWXcsc5_0),.dout(w_dff_B_nlL1oXQa2_0),.clk(gclk));
	jdff dff_A_wPCGl1qU9_1(.dout(w_n188_0[1]),.din(w_dff_A_wPCGl1qU9_1),.clk(gclk));
	jdff dff_B_xmAMFAiU6_0(.din(n298),.dout(w_dff_B_xmAMFAiU6_0),.clk(gclk));
	jdff dff_A_0TVHd13F1_0(.dout(w_n295_0[0]),.din(w_dff_A_0TVHd13F1_0),.clk(gclk));
	jdff dff_B_ElRGm0qY9_2(.din(n291),.dout(w_dff_B_ElRGm0qY9_2),.clk(gclk));
	jdff dff_A_FApMqmB96_2(.dout(w_n290_0[2]),.din(w_dff_A_FApMqmB96_2),.clk(gclk));
	jdff dff_B_HhfOLex49_3(.din(n290),.dout(w_dff_B_HhfOLex49_3),.clk(gclk));
	jdff dff_A_F5N597V85_0(.dout(w_n289_0[0]),.din(w_dff_A_F5N597V85_0),.clk(gclk));
	jdff dff_A_oIpNTQ8z8_0(.dout(w_dff_A_F5N597V85_0),.din(w_dff_A_oIpNTQ8z8_0),.clk(gclk));
	jdff dff_A_KQ9LXcof3_1(.dout(w_n158_0[1]),.din(w_dff_A_KQ9LXcof3_1),.clk(gclk));
	jdff dff_A_BbZgDHH93_0(.dout(w_n92_1[0]),.din(w_dff_A_BbZgDHH93_0),.clk(gclk));
	jdff dff_A_S0id8zff3_0(.dout(w_dff_A_BbZgDHH93_0),.din(w_dff_A_S0id8zff3_0),.clk(gclk));
	jdff dff_A_c9ksjVia9_2(.dout(w_n92_1[2]),.din(w_dff_A_c9ksjVia9_2),.clk(gclk));
	jdff dff_A_psk5xJCz6_1(.dout(w_n163_0[1]),.din(w_dff_A_psk5xJCz6_1),.clk(gclk));
	jdff dff_A_JH53DPRX5_2(.dout(w_n163_0[2]),.din(w_dff_A_JH53DPRX5_2),.clk(gclk));
	jdff dff_B_9jxaQbhS9_1(.din(n123),.dout(w_dff_B_9jxaQbhS9_1),.clk(gclk));
	jdff dff_B_qhZi3BqZ7_1(.din(w_dff_B_9jxaQbhS9_1),.dout(w_dff_B_qhZi3BqZ7_1),.clk(gclk));
	jdff dff_B_2nYgILi63_1(.din(w_dff_B_qhZi3BqZ7_1),.dout(w_dff_B_2nYgILi63_1),.clk(gclk));
	jdff dff_B_WPWpcJ4S9_1(.din(w_dff_B_2nYgILi63_1),.dout(w_dff_B_WPWpcJ4S9_1),.clk(gclk));
	jdff dff_B_N9MFRpiV9_1(.din(w_dff_B_WPWpcJ4S9_1),.dout(w_dff_B_N9MFRpiV9_1),.clk(gclk));
	jdff dff_B_opegiqZu4_0(.din(n284),.dout(w_dff_B_opegiqZu4_0),.clk(gclk));
	jdff dff_B_ESBooY621_0(.din(w_dff_B_opegiqZu4_0),.dout(w_dff_B_ESBooY621_0),.clk(gclk));
	jdff dff_A_E9HyUkut8_0(.dout(w_n68_0[0]),.din(w_dff_A_E9HyUkut8_0),.clk(gclk));
	jdff dff_A_EnfNjDbK7_0(.dout(w_dff_A_E9HyUkut8_0),.din(w_dff_A_EnfNjDbK7_0),.clk(gclk));
	jdff dff_A_lqMR1kOK2_0(.dout(w_dff_A_EnfNjDbK7_0),.din(w_dff_A_lqMR1kOK2_0),.clk(gclk));
	jdff dff_A_yLpA6jkf7_0(.dout(w_dff_A_lqMR1kOK2_0),.din(w_dff_A_yLpA6jkf7_0),.clk(gclk));
	jdff dff_A_xqBNKJBb9_0(.dout(w_dff_A_yLpA6jkf7_0),.din(w_dff_A_xqBNKJBb9_0),.clk(gclk));
	jdff dff_A_EkgqexoQ7_0(.dout(w_dff_A_xqBNKJBb9_0),.din(w_dff_A_EkgqexoQ7_0),.clk(gclk));
	jdff dff_A_Fc7Heav51_0(.dout(w_dff_A_EkgqexoQ7_0),.din(w_dff_A_Fc7Heav51_0),.clk(gclk));
	jdff dff_A_clZThNqh3_1(.dout(w_n281_0[1]),.din(w_dff_A_clZThNqh3_1),.clk(gclk));
	jdff dff_B_U6R6kNON7_3(.din(n281),.dout(w_dff_B_U6R6kNON7_3),.clk(gclk));
	jdff dff_A_xLqE1JzG5_1(.dout(w_n168_0[1]),.din(w_dff_A_xLqE1JzG5_1),.clk(gclk));
	jdff dff_A_9ptEOAnV7_2(.dout(w_n168_0[2]),.din(w_dff_A_9ptEOAnV7_2),.clk(gclk));
	jdff dff_B_dEIbBMUA1_1(.din(n133),.dout(w_dff_B_dEIbBMUA1_1),.clk(gclk));
	jdff dff_B_wGZVrejg7_1(.din(w_dff_B_dEIbBMUA1_1),.dout(w_dff_B_wGZVrejg7_1),.clk(gclk));
	jdff dff_B_DSYPtOPP9_1(.din(w_dff_B_wGZVrejg7_1),.dout(w_dff_B_DSYPtOPP9_1),.clk(gclk));
	jdff dff_B_oRFGlCql2_1(.din(w_dff_B_DSYPtOPP9_1),.dout(w_dff_B_oRFGlCql2_1),.clk(gclk));
	jdff dff_B_rSVmiRJ22_1(.din(w_dff_B_oRFGlCql2_1),.dout(w_dff_B_rSVmiRJ22_1),.clk(gclk));
	jdff dff_A_ihBmT6X81_0(.dout(w_n141_0[0]),.din(w_dff_A_ihBmT6X81_0),.clk(gclk));
	jdff dff_A_6RqHY63b9_0(.dout(w_dff_A_ihBmT6X81_0),.din(w_dff_A_6RqHY63b9_0),.clk(gclk));
	jdff dff_A_3caWganY0_0(.dout(w_dff_A_6RqHY63b9_0),.din(w_dff_A_3caWganY0_0),.clk(gclk));
	jdff dff_A_GEDPlgqP4_0(.dout(w_dff_A_3caWganY0_0),.din(w_dff_A_GEDPlgqP4_0),.clk(gclk));
	jdff dff_A_TZAWdQve4_0(.dout(w_dff_A_GEDPlgqP4_0),.din(w_dff_A_TZAWdQve4_0),.clk(gclk));
	jdff dff_A_U9qEaIsr8_0(.dout(w_dff_A_TZAWdQve4_0),.din(w_dff_A_U9qEaIsr8_0),.clk(gclk));
	jdff dff_A_qQswp3Rc4_0(.dout(w_dff_A_U9qEaIsr8_0),.din(w_dff_A_qQswp3Rc4_0),.clk(gclk));
	jdff dff_A_1WZ6LAoB7_0(.dout(w_dff_A_qQswp3Rc4_0),.din(w_dff_A_1WZ6LAoB7_0),.clk(gclk));
	jdff dff_B_qSEcbz4e4_1(.din(n134),.dout(w_dff_B_qSEcbz4e4_1),.clk(gclk));
	jdff dff_B_NZNl7SDx2_1(.din(w_dff_B_qSEcbz4e4_1),.dout(w_dff_B_NZNl7SDx2_1),.clk(gclk));
	jdff dff_B_2iYyE76X8_0(.din(n138),.dout(w_dff_B_2iYyE76X8_0),.clk(gclk));
	jdff dff_A_YtbwLOvK1_1(.dout(w_G475_0[1]),.din(w_dff_A_YtbwLOvK1_1),.clk(gclk));
	jdff dff_A_fqFOCZqU4_1(.dout(w_dff_A_YtbwLOvK1_1),.din(w_dff_A_fqFOCZqU4_1),.clk(gclk));
	jdff dff_A_iSz2xtx77_1(.dout(w_dff_A_fqFOCZqU4_1),.din(w_dff_A_iSz2xtx77_1),.clk(gclk));
	jdff dff_A_9cDS0aSX6_1(.dout(w_dff_A_iSz2xtx77_1),.din(w_dff_A_9cDS0aSX6_1),.clk(gclk));
	jdff dff_A_dFfHpZLB9_1(.dout(w_dff_A_9cDS0aSX6_1),.din(w_dff_A_dFfHpZLB9_1),.clk(gclk));
	jdff dff_A_a4VxBFAt6_1(.dout(w_dff_A_dFfHpZLB9_1),.din(w_dff_A_a4VxBFAt6_1),.clk(gclk));
	jdff dff_A_eHwbqypz2_0(.dout(w_n130_0[0]),.din(w_dff_A_eHwbqypz2_0),.clk(gclk));
	jdff dff_A_lbJ74lRp3_0(.dout(w_dff_A_eHwbqypz2_0),.din(w_dff_A_lbJ74lRp3_0),.clk(gclk));
	jdff dff_A_xy84moId2_0(.dout(w_dff_A_lbJ74lRp3_0),.din(w_dff_A_xy84moId2_0),.clk(gclk));
	jdff dff_A_c4AWVLou1_0(.dout(w_dff_A_xy84moId2_0),.din(w_dff_A_c4AWVLou1_0),.clk(gclk));
	jdff dff_A_ZMRlQDSQ9_0(.dout(w_dff_A_c4AWVLou1_0),.din(w_dff_A_ZMRlQDSQ9_0),.clk(gclk));
	jdff dff_A_7x47ZWu61_0(.dout(w_dff_A_ZMRlQDSQ9_0),.din(w_dff_A_7x47ZWu61_0),.clk(gclk));
	jdff dff_A_Ub33pQGe3_0(.dout(w_dff_A_7x47ZWu61_0),.din(w_dff_A_Ub33pQGe3_0),.clk(gclk));
	jdff dff_A_YhyKNndE6_0(.dout(w_dff_A_Ub33pQGe3_0),.din(w_dff_A_YhyKNndE6_0),.clk(gclk));
	jdff dff_B_hOZClFAs5_1(.din(n124),.dout(w_dff_B_hOZClFAs5_1),.clk(gclk));
	jdff dff_B_SM4MwVuM7_1(.din(w_dff_B_hOZClFAs5_1),.dout(w_dff_B_SM4MwVuM7_1),.clk(gclk));
	jdff dff_B_m6YuB7hj4_1(.din(w_dff_B_SM4MwVuM7_1),.dout(w_dff_B_m6YuB7hj4_1),.clk(gclk));
	jdff dff_B_I98vDFqU9_0(.din(n128),.dout(w_dff_B_I98vDFqU9_0),.clk(gclk));
	jdff dff_A_2n2Yxywx8_1(.dout(w_G478_0[1]),.din(w_dff_A_2n2Yxywx8_1),.clk(gclk));
	jdff dff_A_y8KKYUSx4_1(.dout(w_dff_A_2n2Yxywx8_1),.din(w_dff_A_y8KKYUSx4_1),.clk(gclk));
	jdff dff_A_R6Id4wSI8_1(.dout(w_dff_A_y8KKYUSx4_1),.din(w_dff_A_R6Id4wSI8_1),.clk(gclk));
	jdff dff_A_X96W8BW71_1(.dout(w_dff_A_R6Id4wSI8_1),.din(w_dff_A_X96W8BW71_1),.clk(gclk));
	jdff dff_A_mqmHQGXz3_1(.dout(w_dff_A_X96W8BW71_1),.din(w_dff_A_mqmHQGXz3_1),.clk(gclk));
	jdff dff_A_3qplDVlv4_1(.dout(w_dff_A_mqmHQGXz3_1),.din(w_dff_A_3qplDVlv4_1),.clk(gclk));
	jdff dff_B_MrzhAbhq1_3(.din(n154),.dout(w_dff_B_MrzhAbhq1_3),.clk(gclk));
	jdff dff_B_fNgSMBRA9_3(.din(w_dff_B_MrzhAbhq1_3),.dout(w_dff_B_fNgSMBRA9_3),.clk(gclk));
	jdff dff_A_9QmyvYKP1_0(.dout(w_n153_0[0]),.din(w_dff_A_9QmyvYKP1_0),.clk(gclk));
	jdff dff_A_S4xbV8Hs5_0(.dout(w_dff_A_9QmyvYKP1_0),.din(w_dff_A_S4xbV8Hs5_0),.clk(gclk));
	jdff dff_A_okHa4Bzi7_1(.dout(w_n153_0[1]),.din(w_dff_A_okHa4Bzi7_1),.clk(gclk));
	jdff dff_A_Ro2hpgkn1_1(.dout(w_dff_A_okHa4Bzi7_1),.din(w_dff_A_Ro2hpgkn1_1),.clk(gclk));
	jdff dff_B_4mOGeCqi9_1(.din(n148),.dout(w_dff_B_4mOGeCqi9_1),.clk(gclk));
	jdff dff_B_qE8bWmkO5_1(.din(w_dff_B_4mOGeCqi9_1),.dout(w_dff_B_qE8bWmkO5_1),.clk(gclk));
	jdff dff_B_YR1gWoKv7_1(.din(w_dff_B_qE8bWmkO5_1),.dout(w_dff_B_YR1gWoKv7_1),.clk(gclk));
	jdff dff_A_iIfVa4Dt5_1(.dout(w_n151_0[1]),.din(w_dff_A_iIfVa4Dt5_1),.clk(gclk));
	jdff dff_A_0XuJysZd7_1(.dout(w_dff_A_iIfVa4Dt5_1),.din(w_dff_A_0XuJysZd7_1),.clk(gclk));
	jdff dff_A_Dylii5uV1_1(.dout(w_dff_A_0XuJysZd7_1),.din(w_dff_A_Dylii5uV1_1),.clk(gclk));
	jdff dff_A_dJZKeeg89_1(.dout(w_dff_A_Dylii5uV1_1),.din(w_dff_A_dJZKeeg89_1),.clk(gclk));
	jdff dff_A_jkYG3eLP8_1(.dout(w_dff_A_dJZKeeg89_1),.din(w_dff_A_jkYG3eLP8_1),.clk(gclk));
	jdff dff_A_Sgcd4f6U3_1(.dout(w_dff_A_jkYG3eLP8_1),.din(w_dff_A_Sgcd4f6U3_1),.clk(gclk));
	jdff dff_A_n5qQQkyW4_1(.dout(w_dff_A_Sgcd4f6U3_1),.din(w_dff_A_n5qQQkyW4_1),.clk(gclk));
	jdff dff_A_D7oeaaDe2_1(.dout(w_dff_A_n5qQQkyW4_1),.din(w_dff_A_D7oeaaDe2_1),.clk(gclk));
	jdff dff_A_cgWO6s0e3_1(.dout(w_G952_0[1]),.din(w_dff_A_cgWO6s0e3_1),.clk(gclk));
	jdff dff_A_TqnVoeS69_1(.dout(w_dff_A_cgWO6s0e3_1),.din(w_dff_A_TqnVoeS69_1),.clk(gclk));
	jdff dff_A_wcUY13iH0_1(.dout(w_dff_A_TqnVoeS69_1),.din(w_dff_A_wcUY13iH0_1),.clk(gclk));
	jdff dff_A_kSzVm8uM8_1(.dout(w_dff_A_wcUY13iH0_1),.din(w_dff_A_kSzVm8uM8_1),.clk(gclk));
	jdff dff_A_ukeACLI76_1(.dout(w_dff_A_kSzVm8uM8_1),.din(w_dff_A_ukeACLI76_1),.clk(gclk));
	jdff dff_A_yB2Frsr14_1(.dout(w_dff_A_ukeACLI76_1),.din(w_dff_A_yB2Frsr14_1),.clk(gclk));
	jdff dff_A_I0rpjgeH9_1(.dout(w_dff_A_yB2Frsr14_1),.din(w_dff_A_I0rpjgeH9_1),.clk(gclk));
	jdff dff_A_Pigc28xR3_1(.dout(w_dff_A_I0rpjgeH9_1),.din(w_dff_A_Pigc28xR3_1),.clk(gclk));
	jdff dff_A_7kAo5nXh7_1(.dout(w_dff_A_Pigc28xR3_1),.din(w_dff_A_7kAo5nXh7_1),.clk(gclk));
	jdff dff_A_dg4Yy4wf7_1(.dout(w_dff_A_7kAo5nXh7_1),.din(w_dff_A_dg4Yy4wf7_1),.clk(gclk));
	jdff dff_A_sfXzP4f65_1(.dout(w_dff_A_dg4Yy4wf7_1),.din(w_dff_A_sfXzP4f65_1),.clk(gclk));
	jdff dff_B_fdscj1JI9_3(.din(G952),.dout(w_dff_B_fdscj1JI9_3),.clk(gclk));
	jdff dff_B_JPJZpma22_1(.din(G898),.dout(w_dff_B_JPJZpma22_1),.clk(gclk));
	jdff dff_B_CwepJYR72_2(.din(n277),.dout(w_dff_B_CwepJYR72_2),.clk(gclk));
	jdff dff_A_vYcfVLIy1_1(.dout(w_n92_0[1]),.din(w_dff_A_vYcfVLIy1_1),.clk(gclk));
	jdff dff_A_zqYekie86_2(.dout(w_n92_0[2]),.din(w_dff_A_zqYekie86_2),.clk(gclk));
	jdff dff_A_gjC2y7aA7_2(.dout(w_dff_A_zqYekie86_2),.din(w_dff_A_gjC2y7aA7_2),.clk(gclk));
	jdff dff_A_CqgGQlX77_1(.dout(w_G472_0[1]),.din(w_dff_A_CqgGQlX77_1),.clk(gclk));
	jdff dff_A_4PhKBgEt9_1(.dout(w_dff_A_CqgGQlX77_1),.din(w_dff_A_4PhKBgEt9_1),.clk(gclk));
	jdff dff_A_XoSdplwf8_1(.dout(w_dff_A_4PhKBgEt9_1),.din(w_dff_A_XoSdplwf8_1),.clk(gclk));
	jdff dff_A_vQqJWAqS3_1(.dout(w_dff_A_XoSdplwf8_1),.din(w_dff_A_vQqJWAqS3_1),.clk(gclk));
	jdff dff_A_jSMj55om2_1(.dout(w_dff_A_vQqJWAqS3_1),.din(w_dff_A_jSMj55om2_1),.clk(gclk));
	jdff dff_A_PiOiHVkx0_1(.dout(w_dff_A_jSMj55om2_1),.din(w_dff_A_PiOiHVkx0_1),.clk(gclk));
	jdff dff_A_zI8VUVET9_0(.dout(w_n73_0[0]),.din(w_dff_A_zI8VUVET9_0),.clk(gclk));
	jdff dff_B_qg1uBTWy8_2(.din(n73),.dout(w_dff_B_qg1uBTWy8_2),.clk(gclk));
	jdff dff_B_RgNxSbqc4_2(.din(w_dff_B_qg1uBTWy8_2),.dout(w_dff_B_RgNxSbqc4_2),.clk(gclk));
	jdff dff_B_OPpNW5H85_2(.din(w_dff_B_RgNxSbqc4_2),.dout(w_dff_B_OPpNW5H85_2),.clk(gclk));
	jdff dff_A_kaVXNc8z2_1(.dout(w_G217_0[1]),.din(w_dff_A_kaVXNc8z2_1),.clk(gclk));
	jdff dff_A_VehClCCv1_1(.dout(w_dff_A_kaVXNc8z2_1),.din(w_dff_A_VehClCCv1_1),.clk(gclk));
	jdff dff_A_pMkwi8aY5_2(.dout(w_G217_0[2]),.din(w_dff_A_pMkwi8aY5_2),.clk(gclk));
	jdff dff_A_lvYd21NF1_2(.dout(w_dff_A_pMkwi8aY5_2),.din(w_dff_A_lvYd21NF1_2),.clk(gclk));
	jdff dff_A_MOEusTo60_2(.dout(w_dff_A_lvYd21NF1_2),.din(w_dff_A_MOEusTo60_2),.clk(gclk));
	jdff dff_A_Imz1djx30_0(.dout(w_n172_0[0]),.din(w_dff_A_Imz1djx30_0),.clk(gclk));
	jdff dff_A_sOHgbdgu6_0(.dout(w_dff_A_Imz1djx30_0),.din(w_dff_A_sOHgbdgu6_0),.clk(gclk));
	jdff dff_A_nPdhDemH2_0(.dout(w_dff_A_sOHgbdgu6_0),.din(w_dff_A_nPdhDemH2_0),.clk(gclk));
	jdff dff_A_FeuGXCMF4_0(.dout(w_dff_A_nPdhDemH2_0),.din(w_dff_A_FeuGXCMF4_0),.clk(gclk));
	jdff dff_A_wiDoK8v92_0(.dout(w_dff_A_FeuGXCMF4_0),.din(w_dff_A_wiDoK8v92_0),.clk(gclk));
	jdff dff_A_FnkGLtEb5_0(.dout(w_dff_A_wiDoK8v92_0),.din(w_dff_A_FnkGLtEb5_0),.clk(gclk));
	jdff dff_B_HLA88eNZ3_1(.din(n171),.dout(w_dff_B_HLA88eNZ3_1),.clk(gclk));
	jdff dff_B_1y5pYWzk4_1(.din(w_dff_B_HLA88eNZ3_1),.dout(w_dff_B_1y5pYWzk4_1),.clk(gclk));
	jdff dff_B_WHlG6HFB2_1(.din(w_dff_B_1y5pYWzk4_1),.dout(w_dff_B_WHlG6HFB2_1),.clk(gclk));
	jdff dff_B_VVnMqQBO2_0(.din(n65),.dout(w_dff_B_VVnMqQBO2_0),.clk(gclk));
	jdff dff_B_qzwN81lV1_0(.din(w_dff_B_VVnMqQBO2_0),.dout(w_dff_B_qzwN81lV1_0),.clk(gclk));
	jdff dff_B_iJOcSZc75_0(.din(w_dff_B_qzwN81lV1_0),.dout(w_dff_B_iJOcSZc75_0),.clk(gclk));
	jdff dff_A_X1VyPlIh4_2(.dout(w_n60_0[2]),.din(w_dff_A_X1VyPlIh4_2),.clk(gclk));
	jdff dff_A_Q0YPYRrC2_2(.dout(w_dff_A_X1VyPlIh4_2),.din(w_dff_A_Q0YPYRrC2_2),.clk(gclk));
	jdff dff_A_ImAltbNP0_2(.dout(w_dff_A_Q0YPYRrC2_2),.din(w_dff_A_ImAltbNP0_2),.clk(gclk));
	jdff dff_A_9Q4mYpeZ7_2(.dout(w_dff_A_ImAltbNP0_2),.din(w_dff_A_9Q4mYpeZ7_2),.clk(gclk));
	jdff dff_A_WAdGVKVL0_0(.dout(w_n59_0[0]),.din(w_dff_A_WAdGVKVL0_0),.clk(gclk));
	jdff dff_A_kwNRHKi92_0(.dout(w_dff_A_WAdGVKVL0_0),.din(w_dff_A_kwNRHKi92_0),.clk(gclk));
	jdff dff_A_oD3XMy220_0(.dout(w_dff_A_kwNRHKi92_0),.din(w_dff_A_oD3XMy220_0),.clk(gclk));
	jdff dff_A_DsDVFYKP5_0(.dout(w_n70_1[0]),.din(w_dff_A_DsDVFYKP5_0),.clk(gclk));
	jdff dff_A_IacUM4se0_0(.dout(w_dff_A_DsDVFYKP5_0),.din(w_dff_A_IacUM4se0_0),.clk(gclk));
	jdff dff_A_Q0UtPfUY9_0(.dout(w_dff_A_IacUM4se0_0),.din(w_dff_A_Q0UtPfUY9_0),.clk(gclk));
	jdff dff_A_WTPZk5ac1_0(.dout(w_dff_A_Q0UtPfUY9_0),.din(w_dff_A_WTPZk5ac1_0),.clk(gclk));
	jdff dff_A_G9Z0dt8A8_0(.dout(w_dff_A_WTPZk5ac1_0),.din(w_dff_A_G9Z0dt8A8_0),.clk(gclk));
	jdff dff_A_4Pgu4pSc6_0(.dout(w_dff_A_G9Z0dt8A8_0),.din(w_dff_A_4Pgu4pSc6_0),.clk(gclk));
	jdff dff_A_dj1IMBKV3_2(.dout(w_n70_1[2]),.din(w_dff_A_dj1IMBKV3_2),.clk(gclk));
	jdff dff_A_cWvGkUWR9_2(.dout(w_dff_A_dj1IMBKV3_2),.din(w_dff_A_cWvGkUWR9_2),.clk(gclk));
	jdff dff_A_001YZGUH6_2(.dout(w_dff_A_cWvGkUWR9_2),.din(w_dff_A_001YZGUH6_2),.clk(gclk));
	jdff dff_A_1Clx8xz59_2(.dout(w_dff_A_001YZGUH6_2),.din(w_dff_A_1Clx8xz59_2),.clk(gclk));
	jdff dff_A_CN1DHKJk6_1(.dout(w_n276_1[1]),.din(w_dff_A_CN1DHKJk6_1),.clk(gclk));
	jdff dff_A_uMjKPJT36_2(.dout(w_n276_0[2]),.din(w_dff_A_uMjKPJT36_2),.clk(gclk));
	jdff dff_B_bhRoY6r93_3(.din(n276),.dout(w_dff_B_bhRoY6r93_3),.clk(gclk));
	jdff dff_B_wPr0VNwI5_1(.din(n195),.dout(w_dff_B_wPr0VNwI5_1),.clk(gclk));
	jdff dff_B_E6QzsEVb9_1(.din(w_dff_B_wPr0VNwI5_1),.dout(w_dff_B_E6QzsEVb9_1),.clk(gclk));
	jdff dff_B_gK1ELPSS8_1(.din(w_dff_B_E6QzsEVb9_1),.dout(w_dff_B_gK1ELPSS8_1),.clk(gclk));
	jdff dff_B_z2HNY8DT5_1(.din(w_dff_B_gK1ELPSS8_1),.dout(w_dff_B_z2HNY8DT5_1),.clk(gclk));
	jdff dff_B_b35UPb6X8_1(.din(w_dff_B_z2HNY8DT5_1),.dout(w_dff_B_b35UPb6X8_1),.clk(gclk));
	jdff dff_A_SAYqYeAA6_0(.dout(w_n117_0[0]),.din(w_dff_A_SAYqYeAA6_0),.clk(gclk));
	jdff dff_A_PSWQlojB4_0(.dout(w_dff_A_SAYqYeAA6_0),.din(w_dff_A_PSWQlojB4_0),.clk(gclk));
	jdff dff_A_HW16vTXj7_0(.dout(w_dff_A_PSWQlojB4_0),.din(w_dff_A_HW16vTXj7_0),.clk(gclk));
	jdff dff_A_I7WEYVly6_0(.dout(w_dff_A_HW16vTXj7_0),.din(w_dff_A_I7WEYVly6_0),.clk(gclk));
	jdff dff_A_9B813XqM8_0(.dout(w_dff_A_I7WEYVly6_0),.din(w_dff_A_9B813XqM8_0),.clk(gclk));
	jdff dff_A_B3Rzr5Ie7_0(.dout(w_dff_A_9B813XqM8_0),.din(w_dff_A_B3Rzr5Ie7_0),.clk(gclk));
	jdff dff_A_6dDmuJIW0_0(.dout(w_dff_A_B3Rzr5Ie7_0),.din(w_dff_A_6dDmuJIW0_0),.clk(gclk));
	jdff dff_A_PHCmtKUe5_0(.dout(w_dff_A_6dDmuJIW0_0),.din(w_dff_A_PHCmtKUe5_0),.clk(gclk));
	jdff dff_B_occ79nkz0_1(.din(n113),.dout(w_dff_B_occ79nkz0_1),.clk(gclk));
	jdff dff_B_XF7aPHFI7_1(.din(w_dff_B_occ79nkz0_1),.dout(w_dff_B_XF7aPHFI7_1),.clk(gclk));
	jdff dff_B_XwWUbyaA9_2(.din(G227),.dout(w_dff_B_XwWUbyaA9_2),.clk(gclk));
	jdff dff_A_2Pwe5xD42_0(.dout(w_G140_0[0]),.din(w_dff_A_2Pwe5xD42_0),.clk(gclk));
	jdff dff_A_ob64nq451_0(.dout(w_dff_A_2Pwe5xD42_0),.din(w_dff_A_ob64nq451_0),.clk(gclk));
	jdff dff_A_dIDDNrYK9_0(.dout(w_dff_A_ob64nq451_0),.din(w_dff_A_dIDDNrYK9_0),.clk(gclk));
	jdff dff_A_G7RP05tB1_0(.dout(w_dff_A_dIDDNrYK9_0),.din(w_dff_A_G7RP05tB1_0),.clk(gclk));
	jdff dff_A_s7KsCvYc6_0(.dout(w_dff_A_G7RP05tB1_0),.din(w_dff_A_s7KsCvYc6_0),.clk(gclk));
	jdff dff_A_Pm5qag2M2_0(.dout(w_dff_A_s7KsCvYc6_0),.din(w_dff_A_Pm5qag2M2_0),.clk(gclk));
	jdff dff_A_D9thSa8h3_0(.dout(w_dff_A_Pm5qag2M2_0),.din(w_dff_A_D9thSa8h3_0),.clk(gclk));
	jdff dff_A_c0MtNqIm1_0(.dout(w_dff_A_D9thSa8h3_0),.din(w_dff_A_c0MtNqIm1_0),.clk(gclk));
	jdff dff_A_vIZevEEt4_0(.dout(w_dff_A_c0MtNqIm1_0),.din(w_dff_A_vIZevEEt4_0),.clk(gclk));
	jdff dff_A_wig9lR7E1_0(.dout(w_dff_A_vIZevEEt4_0),.din(w_dff_A_wig9lR7E1_0),.clk(gclk));
	jdff dff_A_NaXfPu0L9_0(.dout(w_dff_A_wig9lR7E1_0),.din(w_dff_A_NaXfPu0L9_0),.clk(gclk));
	jdff dff_A_1T56NcLb3_0(.dout(w_dff_A_NaXfPu0L9_0),.din(w_dff_A_1T56NcLb3_0),.clk(gclk));
	jdff dff_A_CmI19uGM8_2(.dout(w_G469_0[2]),.din(w_dff_A_CmI19uGM8_2),.clk(gclk));
	jdff dff_A_UKa6iSEb7_2(.dout(w_dff_A_CmI19uGM8_2),.din(w_dff_A_UKa6iSEb7_2),.clk(gclk));
	jdff dff_A_GL32B1qB5_2(.dout(w_dff_A_UKa6iSEb7_2),.din(w_dff_A_GL32B1qB5_2),.clk(gclk));
	jdff dff_A_V9o54ueu7_2(.dout(w_dff_A_GL32B1qB5_2),.din(w_dff_A_V9o54ueu7_2),.clk(gclk));
	jdff dff_A_hABQ7jQC6_2(.dout(w_dff_A_V9o54ueu7_2),.din(w_dff_A_hABQ7jQC6_2),.clk(gclk));
	jdff dff_A_wRghbfZ99_2(.dout(w_dff_A_hABQ7jQC6_2),.din(w_dff_A_wRghbfZ99_2),.clk(gclk));
	jdff dff_B_R5NvZTUM2_2(.din(n274),.dout(w_dff_B_R5NvZTUM2_2),.clk(gclk));
	jdff dff_B_ZtOJtenl6_2(.din(w_dff_B_R5NvZTUM2_2),.dout(w_dff_B_ZtOJtenl6_2),.clk(gclk));
	jdff dff_B_mjWg5OmM2_2(.din(w_dff_B_ZtOJtenl6_2),.dout(w_dff_B_mjWg5OmM2_2),.clk(gclk));
	jdff dff_B_iXVu6Lhd7_2(.din(w_dff_B_mjWg5OmM2_2),.dout(w_dff_B_iXVu6Lhd7_2),.clk(gclk));
	jdff dff_A_kLuhzMdc3_0(.dout(w_n112_0[0]),.din(w_dff_A_kLuhzMdc3_0),.clk(gclk));
	jdff dff_A_gnm3weAu1_0(.dout(w_dff_A_kLuhzMdc3_0),.din(w_dff_A_gnm3weAu1_0),.clk(gclk));
	jdff dff_A_hR1qtTLz2_0(.dout(w_dff_A_gnm3weAu1_0),.din(w_dff_A_hR1qtTLz2_0),.clk(gclk));
	jdff dff_A_YXptWKBs5_0(.dout(w_dff_A_hR1qtTLz2_0),.din(w_dff_A_YXptWKBs5_0),.clk(gclk));
	jdff dff_A_vi6JzD1y3_0(.dout(w_dff_A_YXptWKBs5_0),.din(w_dff_A_vi6JzD1y3_0),.clk(gclk));
	jdff dff_B_nwK763Rc6_1(.din(n111),.dout(w_dff_B_nwK763Rc6_1),.clk(gclk));
	jdff dff_A_fW8uNh8t5_0(.dout(w_n70_3[0]),.din(w_dff_A_fW8uNh8t5_0),.clk(gclk));
	jdff dff_A_ulwh2wrP4_0(.dout(w_dff_A_fW8uNh8t5_0),.din(w_dff_A_ulwh2wrP4_0),.clk(gclk));
	jdff dff_A_e1f2Foyk0_0(.dout(w_dff_A_ulwh2wrP4_0),.din(w_dff_A_e1f2Foyk0_0),.clk(gclk));
	jdff dff_A_4wBYh1qH1_0(.dout(w_dff_A_e1f2Foyk0_0),.din(w_dff_A_4wBYh1qH1_0),.clk(gclk));
	jdff dff_A_gsFWYLBg9_1(.dout(w_G234_0[1]),.din(w_dff_A_gsFWYLBg9_1),.clk(gclk));
	jdff dff_A_El32Yq4F9_2(.dout(w_G234_0[2]),.din(w_dff_A_El32Yq4F9_2),.clk(gclk));
	jdff dff_A_BVXrdtrh1_1(.dout(w_G221_0[1]),.din(w_dff_A_BVXrdtrh1_1),.clk(gclk));
	jdff dff_A_epkGa6cy4_1(.dout(w_dff_A_BVXrdtrh1_1),.din(w_dff_A_epkGa6cy4_1),.clk(gclk));
	jdff dff_A_71NluWUL3_1(.dout(w_n216_0[1]),.din(w_dff_A_71NluWUL3_1),.clk(gclk));
	jdff dff_B_5iqB7ot68_1(.din(n215),.dout(w_dff_B_5iqB7ot68_1),.clk(gclk));
	jdff dff_B_HwDtq9ba8_1(.din(w_dff_B_5iqB7ot68_1),.dout(w_dff_B_HwDtq9ba8_1),.clk(gclk));
	jdff dff_B_jNMOTHPc9_1(.din(w_dff_B_HwDtq9ba8_1),.dout(w_dff_B_jNMOTHPc9_1),.clk(gclk));
	jdff dff_B_PFrBXyXU6_1(.din(w_dff_B_jNMOTHPc9_1),.dout(w_dff_B_PFrBXyXU6_1),.clk(gclk));
	jdff dff_A_YzWqgtEM3_0(.dout(w_n107_0[0]),.din(w_dff_A_YzWqgtEM3_0),.clk(gclk));
	jdff dff_A_OmQqO8tT0_0(.dout(w_dff_A_YzWqgtEM3_0),.din(w_dff_A_OmQqO8tT0_0),.clk(gclk));
	jdff dff_A_AjiuBpna8_0(.dout(w_dff_A_OmQqO8tT0_0),.din(w_dff_A_AjiuBpna8_0),.clk(gclk));
	jdff dff_A_Nid2gwQV2_0(.dout(w_dff_A_AjiuBpna8_0),.din(w_dff_A_Nid2gwQV2_0),.clk(gclk));
	jdff dff_A_WBaCJjy50_0(.dout(w_dff_A_Nid2gwQV2_0),.din(w_dff_A_WBaCJjy50_0),.clk(gclk));
	jdff dff_A_TMVH4ehc8_0(.dout(w_dff_A_WBaCJjy50_0),.din(w_dff_A_TMVH4ehc8_0),.clk(gclk));
	jdff dff_A_J7D7C9zu3_0(.dout(w_dff_A_TMVH4ehc8_0),.din(w_dff_A_J7D7C9zu3_0),.clk(gclk));
	jdff dff_A_A4XgrKl65_0(.dout(w_dff_A_J7D7C9zu3_0),.din(w_dff_A_A4XgrKl65_0),.clk(gclk));
	jdff dff_B_SLrfBU200_1(.din(n104),.dout(w_dff_B_SLrfBU200_1),.clk(gclk));
	jdff dff_A_kOlMzfbA4_0(.dout(w_G125_0[0]),.din(w_dff_A_kOlMzfbA4_0),.clk(gclk));
	jdff dff_A_VqhBz2OE9_0(.dout(w_dff_A_kOlMzfbA4_0),.din(w_dff_A_VqhBz2OE9_0),.clk(gclk));
	jdff dff_A_bDnFGNFv6_0(.dout(w_dff_A_VqhBz2OE9_0),.din(w_dff_A_bDnFGNFv6_0),.clk(gclk));
	jdff dff_A_ztGTFqxF8_0(.dout(w_dff_A_bDnFGNFv6_0),.din(w_dff_A_ztGTFqxF8_0),.clk(gclk));
	jdff dff_A_rwGRa3Gc2_0(.dout(w_dff_A_ztGTFqxF8_0),.din(w_dff_A_rwGRa3Gc2_0),.clk(gclk));
	jdff dff_A_4yRaVz2j3_0(.dout(w_dff_A_rwGRa3Gc2_0),.din(w_dff_A_4yRaVz2j3_0),.clk(gclk));
	jdff dff_A_Ofm4sO5M1_0(.dout(w_dff_A_4yRaVz2j3_0),.din(w_dff_A_Ofm4sO5M1_0),.clk(gclk));
	jdff dff_A_ZCPcl85m3_0(.dout(w_dff_A_Ofm4sO5M1_0),.din(w_dff_A_ZCPcl85m3_0),.clk(gclk));
	jdff dff_A_VNRUGPVX2_0(.dout(w_dff_A_ZCPcl85m3_0),.din(w_dff_A_VNRUGPVX2_0),.clk(gclk));
	jdff dff_A_EmibUZNn8_0(.dout(w_dff_A_VNRUGPVX2_0),.din(w_dff_A_EmibUZNn8_0),.clk(gclk));
	jdff dff_A_ZN1uhVPD6_0(.dout(w_dff_A_EmibUZNn8_0),.din(w_dff_A_ZN1uhVPD6_0),.clk(gclk));
	jdff dff_A_TZgUmoyB5_0(.dout(w_dff_A_ZN1uhVPD6_0),.din(w_dff_A_TZgUmoyB5_0),.clk(gclk));
	jdff dff_A_oqaEsJhU9_1(.dout(w_G125_0[1]),.din(w_dff_A_oqaEsJhU9_1),.clk(gclk));
	jdff dff_A_7RDDJqxm0_1(.dout(w_dff_A_oqaEsJhU9_1),.din(w_dff_A_7RDDJqxm0_1),.clk(gclk));
	jdff dff_B_j8NchfuQ0_2(.din(G224),.dout(w_dff_B_j8NchfuQ0_2),.clk(gclk));
	jdff dff_A_acQ6BEHC1_0(.dout(w_n103_0[0]),.din(w_dff_A_acQ6BEHC1_0),.clk(gclk));
	jdff dff_A_B4KoY9132_0(.dout(w_dff_A_acQ6BEHC1_0),.din(w_dff_A_B4KoY9132_0),.clk(gclk));
	jdff dff_A_7GwyrfkY4_0(.dout(w_dff_A_B4KoY9132_0),.din(w_dff_A_7GwyrfkY4_0),.clk(gclk));
	jdff dff_A_U9yKmZmb1_0(.dout(w_dff_A_7GwyrfkY4_0),.din(w_dff_A_U9yKmZmb1_0),.clk(gclk));
	jdff dff_A_xzGsgmxU6_0(.dout(w_dff_A_U9yKmZmb1_0),.din(w_dff_A_xzGsgmxU6_0),.clk(gclk));
	jdff dff_A_YDczaK3y5_0(.dout(w_dff_A_xzGsgmxU6_0),.din(w_dff_A_YDczaK3y5_0),.clk(gclk));
	jdff dff_A_BrdlmCpc2_0(.dout(w_dff_A_YDczaK3y5_0),.din(w_dff_A_BrdlmCpc2_0),.clk(gclk));
	jdff dff_A_ALXZVDQY9_0(.dout(w_dff_A_BrdlmCpc2_0),.din(w_dff_A_ALXZVDQY9_0),.clk(gclk));
	jdff dff_A_KazlaGO74_0(.dout(w_dff_A_ALXZVDQY9_0),.din(w_dff_A_KazlaGO74_0),.clk(gclk));
	jdff dff_A_8dtt8jhM9_0(.dout(w_dff_A_KazlaGO74_0),.din(w_dff_A_8dtt8jhM9_0),.clk(gclk));
	jdff dff_B_xd96ETnW8_1(.din(n99),.dout(w_dff_B_xd96ETnW8_1),.clk(gclk));
	jdff dff_A_JlWKuqRR8_0(.dout(w_G107_0[0]),.din(w_dff_A_JlWKuqRR8_0),.clk(gclk));
	jdff dff_A_eHbWDQ225_0(.dout(w_dff_A_JlWKuqRR8_0),.din(w_dff_A_eHbWDQ225_0),.clk(gclk));
	jdff dff_A_derTroX22_0(.dout(w_dff_A_eHbWDQ225_0),.din(w_dff_A_derTroX22_0),.clk(gclk));
	jdff dff_A_EWZZk98l8_0(.dout(w_dff_A_derTroX22_0),.din(w_dff_A_EWZZk98l8_0),.clk(gclk));
	jdff dff_A_XxAhpcdm3_0(.dout(w_dff_A_EWZZk98l8_0),.din(w_dff_A_XxAhpcdm3_0),.clk(gclk));
	jdff dff_A_BgBLwZxo2_0(.dout(w_dff_A_XxAhpcdm3_0),.din(w_dff_A_BgBLwZxo2_0),.clk(gclk));
	jdff dff_A_dLiz0d3b6_0(.dout(w_dff_A_BgBLwZxo2_0),.din(w_dff_A_dLiz0d3b6_0),.clk(gclk));
	jdff dff_A_3En41kxw5_0(.dout(w_dff_A_dLiz0d3b6_0),.din(w_dff_A_3En41kxw5_0),.clk(gclk));
	jdff dff_A_4O1YrcTA3_0(.dout(w_dff_A_3En41kxw5_0),.din(w_dff_A_4O1YrcTA3_0),.clk(gclk));
	jdff dff_A_gHPRsLIL2_0(.dout(w_dff_A_4O1YrcTA3_0),.din(w_dff_A_gHPRsLIL2_0),.clk(gclk));
	jdff dff_A_XFy2QIpz0_0(.dout(w_dff_A_gHPRsLIL2_0),.din(w_dff_A_XFy2QIpz0_0),.clk(gclk));
	jdff dff_A_GJISJ8Pl9_0(.dout(w_G104_0[0]),.din(w_dff_A_GJISJ8Pl9_0),.clk(gclk));
	jdff dff_A_GC5GjNp01_0(.dout(w_dff_A_GJISJ8Pl9_0),.din(w_dff_A_GC5GjNp01_0),.clk(gclk));
	jdff dff_A_P1HxWyZA5_0(.dout(w_dff_A_GC5GjNp01_0),.din(w_dff_A_P1HxWyZA5_0),.clk(gclk));
	jdff dff_A_qVYgheDy9_0(.dout(w_dff_A_P1HxWyZA5_0),.din(w_dff_A_qVYgheDy9_0),.clk(gclk));
	jdff dff_A_5TNbuzRu1_0(.dout(w_dff_A_qVYgheDy9_0),.din(w_dff_A_5TNbuzRu1_0),.clk(gclk));
	jdff dff_A_3FDNVewa7_0(.dout(w_dff_A_5TNbuzRu1_0),.din(w_dff_A_3FDNVewa7_0),.clk(gclk));
	jdff dff_A_6kPDtOT71_0(.dout(w_dff_A_3FDNVewa7_0),.din(w_dff_A_6kPDtOT71_0),.clk(gclk));
	jdff dff_A_yjAX5vwI9_0(.dout(w_dff_A_6kPDtOT71_0),.din(w_dff_A_yjAX5vwI9_0),.clk(gclk));
	jdff dff_A_W6H8pUiF4_0(.dout(w_dff_A_yjAX5vwI9_0),.din(w_dff_A_W6H8pUiF4_0),.clk(gclk));
	jdff dff_A_yHUWdIBR4_0(.dout(w_dff_A_W6H8pUiF4_0),.din(w_dff_A_yHUWdIBR4_0),.clk(gclk));
	jdff dff_A_3LXgP0c93_0(.dout(w_dff_A_yHUWdIBR4_0),.din(w_dff_A_3LXgP0c93_0),.clk(gclk));
	jdff dff_A_jwEtlGrS2_1(.dout(w_G104_0[1]),.din(w_dff_A_jwEtlGrS2_1),.clk(gclk));
	jdff dff_A_zNv4tfBu4_1(.dout(w_dff_A_jwEtlGrS2_1),.din(w_dff_A_zNv4tfBu4_1),.clk(gclk));
	jdff dff_A_9DdSNxao3_1(.dout(w_G122_1[1]),.din(w_dff_A_9DdSNxao3_1),.clk(gclk));
	jdff dff_A_2GK19s0i0_1(.dout(w_G122_0[1]),.din(w_dff_A_2GK19s0i0_1),.clk(gclk));
	jdff dff_A_z650O9AP3_1(.dout(w_dff_A_2GK19s0i0_1),.din(w_dff_A_z650O9AP3_1),.clk(gclk));
	jdff dff_A_UIemolCt2_1(.dout(w_dff_A_z650O9AP3_1),.din(w_dff_A_UIemolCt2_1),.clk(gclk));
	jdff dff_A_F7YPdviM6_1(.dout(w_dff_A_UIemolCt2_1),.din(w_dff_A_F7YPdviM6_1),.clk(gclk));
	jdff dff_A_iIVvANJ47_1(.dout(w_dff_A_F7YPdviM6_1),.din(w_dff_A_iIVvANJ47_1),.clk(gclk));
	jdff dff_A_K4wuwk3z8_1(.dout(w_dff_A_iIVvANJ47_1),.din(w_dff_A_K4wuwk3z8_1),.clk(gclk));
	jdff dff_A_EzXFpg7j1_1(.dout(w_dff_A_K4wuwk3z8_1),.din(w_dff_A_EzXFpg7j1_1),.clk(gclk));
	jdff dff_A_GSjoSRex1_1(.dout(w_dff_A_EzXFpg7j1_1),.din(w_dff_A_GSjoSRex1_1),.clk(gclk));
	jdff dff_A_BTA3jP3j7_1(.dout(w_dff_A_GSjoSRex1_1),.din(w_dff_A_BTA3jP3j7_1),.clk(gclk));
	jdff dff_A_9hMkmGVH8_1(.dout(w_dff_A_BTA3jP3j7_1),.din(w_dff_A_9hMkmGVH8_1),.clk(gclk));
	jdff dff_A_XdZ53zG34_1(.dout(w_dff_A_9hMkmGVH8_1),.din(w_dff_A_XdZ53zG34_1),.clk(gclk));
	jdff dff_A_ny2tcttW0_2(.dout(w_G122_0[2]),.din(w_dff_A_ny2tcttW0_2),.clk(gclk));
	jdff dff_A_ABcTzrzq6_1(.dout(w_G110_1[1]),.din(w_dff_A_ABcTzrzq6_1),.clk(gclk));
	jdff dff_A_WVPUjYEs2_1(.dout(w_dff_A_ABcTzrzq6_1),.din(w_dff_A_WVPUjYEs2_1),.clk(gclk));
	jdff dff_A_yy4fQQUe6_1(.dout(w_dff_A_WVPUjYEs2_1),.din(w_dff_A_yy4fQQUe6_1),.clk(gclk));
	jdff dff_A_J15qkT5W3_1(.dout(w_dff_A_yy4fQQUe6_1),.din(w_dff_A_J15qkT5W3_1),.clk(gclk));
	jdff dff_A_4oX8d2lL8_1(.dout(w_dff_A_J15qkT5W3_1),.din(w_dff_A_4oX8d2lL8_1),.clk(gclk));
	jdff dff_A_zcGxgUb23_1(.dout(w_G110_0[1]),.din(w_dff_A_zcGxgUb23_1),.clk(gclk));
	jdff dff_A_vtlyfzYp8_1(.dout(w_dff_A_zcGxgUb23_1),.din(w_dff_A_vtlyfzYp8_1),.clk(gclk));
	jdff dff_A_75rzG71e3_1(.dout(w_dff_A_vtlyfzYp8_1),.din(w_dff_A_75rzG71e3_1),.clk(gclk));
	jdff dff_A_IwoBo1on5_1(.dout(w_dff_A_75rzG71e3_1),.din(w_dff_A_IwoBo1on5_1),.clk(gclk));
	jdff dff_A_iFccukDN9_1(.dout(w_dff_A_IwoBo1on5_1),.din(w_dff_A_iFccukDN9_1),.clk(gclk));
	jdff dff_A_EGB9BWmx9_1(.dout(w_dff_A_iFccukDN9_1),.din(w_dff_A_EGB9BWmx9_1),.clk(gclk));
	jdff dff_A_dRvqBBIl1_1(.dout(w_dff_A_EGB9BWmx9_1),.din(w_dff_A_dRvqBBIl1_1),.clk(gclk));
	jdff dff_A_XBzWfh0L6_1(.dout(w_dff_A_dRvqBBIl1_1),.din(w_dff_A_XBzWfh0L6_1),.clk(gclk));
	jdff dff_A_rrns76VM5_1(.dout(w_dff_A_XBzWfh0L6_1),.din(w_dff_A_rrns76VM5_1),.clk(gclk));
	jdff dff_A_EpIsYTrm1_1(.dout(w_dff_A_rrns76VM5_1),.din(w_dff_A_EpIsYTrm1_1),.clk(gclk));
	jdff dff_A_MZFvmqbH6_1(.dout(w_dff_A_EpIsYTrm1_1),.din(w_dff_A_MZFvmqbH6_1),.clk(gclk));
	jdff dff_A_6Y0SRe8A8_1(.dout(w_dff_A_MZFvmqbH6_1),.din(w_dff_A_6Y0SRe8A8_1),.clk(gclk));
	jdff dff_A_TYclLP6L4_1(.dout(w_n70_0[1]),.din(w_dff_A_TYclLP6L4_1),.clk(gclk));
	jdff dff_A_QMLcamct7_1(.dout(w_dff_A_TYclLP6L4_1),.din(w_dff_A_QMLcamct7_1),.clk(gclk));
	jdff dff_A_cRoJLPQA3_1(.dout(w_dff_A_QMLcamct7_1),.din(w_dff_A_cRoJLPQA3_1),.clk(gclk));
	jdff dff_A_JXaWVVBu4_1(.dout(w_dff_A_cRoJLPQA3_1),.din(w_dff_A_JXaWVVBu4_1),.clk(gclk));
	jdff dff_A_XNAk2NZk7_1(.dout(w_n97_0[1]),.din(w_dff_A_XNAk2NZk7_1),.clk(gclk));
	jdff dff_A_3kGUtjRt9_1(.dout(w_dff_A_XNAk2NZk7_1),.din(w_dff_A_3kGUtjRt9_1),.clk(gclk));
	jdff dff_A_rV874PmD9_1(.dout(w_dff_A_3kGUtjRt9_1),.din(w_dff_A_rV874PmD9_1),.clk(gclk));
	jdff dff_A_xZ7tDhxY8_1(.dout(w_dff_A_rV874PmD9_1),.din(w_dff_A_xZ7tDhxY8_1),.clk(gclk));
	jdff dff_A_VN6hA1Nm1_1(.dout(w_dff_A_xZ7tDhxY8_1),.din(w_dff_A_VN6hA1Nm1_1),.clk(gclk));
	jdff dff_A_8wjsgzGh7_0(.dout(w_n95_0[0]),.din(w_dff_A_8wjsgzGh7_0),.clk(gclk));
	jdff dff_A_lcM2ykDn8_0(.dout(w_dff_A_8wjsgzGh7_0),.din(w_dff_A_lcM2ykDn8_0),.clk(gclk));
	jdff dff_A_8166cvVF4_0(.dout(w_dff_A_lcM2ykDn8_0),.din(w_dff_A_8166cvVF4_0),.clk(gclk));
	jdff dff_A_PvPANHgX4_0(.dout(w_dff_A_8166cvVF4_0),.din(w_dff_A_PvPANHgX4_0),.clk(gclk));
	jdff dff_A_vvtOcw8v3_0(.dout(w_dff_A_PvPANHgX4_0),.din(w_dff_A_vvtOcw8v3_0),.clk(gclk));
	jdff dff_A_4sr6rX5J6_0(.dout(w_dff_A_vvtOcw8v3_0),.din(w_dff_A_4sr6rX5J6_0),.clk(gclk));
	jdff dff_A_6kKjIGKo4_1(.dout(w_n95_0[1]),.din(w_dff_A_6kKjIGKo4_1),.clk(gclk));
	jdff dff_A_dpZiBVzy7_1(.dout(w_dff_A_6kKjIGKo4_1),.din(w_dff_A_dpZiBVzy7_1),.clk(gclk));
	jdff dff_A_DQ7uY5mP0_1(.dout(w_dff_A_dpZiBVzy7_1),.din(w_dff_A_DQ7uY5mP0_1),.clk(gclk));
	jdff dff_A_wjDOrDyr6_1(.dout(w_dff_A_DQ7uY5mP0_1),.din(w_dff_A_wjDOrDyr6_1),.clk(gclk));
	jdff dff_A_sFH2u8nm8_1(.dout(w_dff_A_wjDOrDyr6_1),.din(w_dff_A_sFH2u8nm8_1),.clk(gclk));
	jdff dff_A_yUMrUTrr4_1(.dout(w_dff_A_sFH2u8nm8_1),.din(w_dff_A_yUMrUTrr4_1),.clk(gclk));
	jdff dff_A_HhxTUasi1_2(.dout(w_G902_3[2]),.din(w_dff_A_HhxTUasi1_2),.clk(gclk));
	jdff dff_A_ZD40DTeX6_2(.dout(w_dff_A_HhxTUasi1_2),.din(w_dff_A_ZD40DTeX6_2),.clk(gclk));
	jdff dff_A_xkE8FqOR1_2(.dout(w_dff_A_ZD40DTeX6_2),.din(w_dff_A_xkE8FqOR1_2),.clk(gclk));
	jdff dff_A_xFZzRMFV9_2(.dout(w_dff_A_xkE8FqOR1_2),.din(w_dff_A_xFZzRMFV9_2),.clk(gclk));
	jdff dff_A_XV0vLJNQ4_2(.dout(w_dff_A_xFZzRMFV9_2),.din(w_dff_A_XV0vLJNQ4_2),.clk(gclk));
	jdff dff_A_9cQh8x9l0_2(.dout(w_dff_A_XV0vLJNQ4_2),.din(w_dff_A_9cQh8x9l0_2),.clk(gclk));
	jdff dff_A_oa6Wi5jE0_2(.dout(w_dff_A_9cQh8x9l0_2),.din(w_dff_A_oa6Wi5jE0_2),.clk(gclk));
	jdff dff_A_Xr5gq0lD3_0(.dout(w_n90_0[0]),.din(w_dff_A_Xr5gq0lD3_0),.clk(gclk));
	jdff dff_A_H0g2eFmb7_0(.dout(w_dff_A_Xr5gq0lD3_0),.din(w_dff_A_H0g2eFmb7_0),.clk(gclk));
	jdff dff_A_jc4OPAdb0_0(.dout(w_dff_A_H0g2eFmb7_0),.din(w_dff_A_jc4OPAdb0_0),.clk(gclk));
	jdff dff_A_op7mq9RO8_0(.dout(w_dff_A_jc4OPAdb0_0),.din(w_dff_A_op7mq9RO8_0),.clk(gclk));
	jdff dff_A_drDN8AOp0_0(.dout(w_dff_A_op7mq9RO8_0),.din(w_dff_A_drDN8AOp0_0),.clk(gclk));
	jdff dff_A_mtDt0H3R5_0(.dout(w_dff_A_drDN8AOp0_0),.din(w_dff_A_mtDt0H3R5_0),.clk(gclk));
	jdff dff_A_SAgvGc9c8_0(.dout(w_dff_A_mtDt0H3R5_0),.din(w_dff_A_SAgvGc9c8_0),.clk(gclk));
	jdff dff_A_xEf78y8R0_0(.dout(w_dff_A_SAgvGc9c8_0),.din(w_dff_A_xEf78y8R0_0),.clk(gclk));
	jdff dff_B_pbx0NWAq9_0(.din(n89),.dout(w_dff_B_pbx0NWAq9_0),.clk(gclk));
	jdff dff_B_2dX0KMoU9_2(.din(n86),.dout(w_dff_B_2dX0KMoU9_2),.clk(gclk));
	jdff dff_A_rN4PWyHm5_0(.dout(w_G953_1[0]),.din(w_dff_A_rN4PWyHm5_0),.clk(gclk));
	jdff dff_A_eZ42Bc6Y4_0(.dout(w_dff_A_rN4PWyHm5_0),.din(w_dff_A_eZ42Bc6Y4_0),.clk(gclk));
	jdff dff_A_S1QrIG7Q1_0(.dout(w_dff_A_eZ42Bc6Y4_0),.din(w_dff_A_S1QrIG7Q1_0),.clk(gclk));
	jdff dff_A_NLhFgFi00_0(.dout(w_dff_A_S1QrIG7Q1_0),.din(w_dff_A_NLhFgFi00_0),.clk(gclk));
	jdff dff_A_YvTB9ISE9_0(.dout(w_dff_A_NLhFgFi00_0),.din(w_dff_A_YvTB9ISE9_0),.clk(gclk));
	jdff dff_A_YJnwZ44V1_0(.dout(w_dff_A_YvTB9ISE9_0),.din(w_dff_A_YJnwZ44V1_0),.clk(gclk));
	jdff dff_A_FwqwMjRY3_0(.dout(w_dff_A_YJnwZ44V1_0),.din(w_dff_A_FwqwMjRY3_0),.clk(gclk));
	jdff dff_A_OjNuXhHU0_0(.dout(w_dff_A_FwqwMjRY3_0),.din(w_dff_A_OjNuXhHU0_0),.clk(gclk));
	jdff dff_A_NQ4qOvEp7_0(.dout(w_dff_A_OjNuXhHU0_0),.din(w_dff_A_NQ4qOvEp7_0),.clk(gclk));
	jdff dff_A_EHVgwXFq4_0(.dout(w_dff_A_NQ4qOvEp7_0),.din(w_dff_A_EHVgwXFq4_0),.clk(gclk));
	jdff dff_A_jKJOKbtK3_0(.dout(w_dff_A_EHVgwXFq4_0),.din(w_dff_A_jKJOKbtK3_0),.clk(gclk));
	jdff dff_A_IGaND4c64_1(.dout(w_G953_0[1]),.din(w_dff_A_IGaND4c64_1),.clk(gclk));
	jdff dff_A_714Enl0P3_1(.dout(w_dff_A_IGaND4c64_1),.din(w_dff_A_714Enl0P3_1),.clk(gclk));
	jdff dff_A_wNfGWoYm2_1(.dout(w_dff_A_714Enl0P3_1),.din(w_dff_A_wNfGWoYm2_1),.clk(gclk));
	jdff dff_A_iVbfdqdV1_1(.dout(w_dff_A_wNfGWoYm2_1),.din(w_dff_A_iVbfdqdV1_1),.clk(gclk));
	jdff dff_A_aInKHHQv8_1(.dout(w_dff_A_iVbfdqdV1_1),.din(w_dff_A_aInKHHQv8_1),.clk(gclk));
	jdff dff_A_eVyqfnfQ6_1(.dout(w_dff_A_aInKHHQv8_1),.din(w_dff_A_eVyqfnfQ6_1),.clk(gclk));
	jdff dff_A_P4RmtLTS0_1(.dout(w_dff_A_eVyqfnfQ6_1),.din(w_dff_A_P4RmtLTS0_1),.clk(gclk));
	jdff dff_A_zAQi7Tox5_1(.dout(w_dff_A_P4RmtLTS0_1),.din(w_dff_A_zAQi7Tox5_1),.clk(gclk));
	jdff dff_A_1N14BGgV1_1(.dout(w_dff_A_zAQi7Tox5_1),.din(w_dff_A_1N14BGgV1_1),.clk(gclk));
	jdff dff_A_ZwgU9lFw0_1(.dout(w_dff_A_1N14BGgV1_1),.din(w_dff_A_ZwgU9lFw0_1),.clk(gclk));
	jdff dff_A_WfePsrL82_1(.dout(w_dff_A_ZwgU9lFw0_1),.din(w_dff_A_WfePsrL82_1),.clk(gclk));
	jdff dff_A_fHj8Qlmy9_1(.dout(w_dff_A_WfePsrL82_1),.din(w_dff_A_fHj8Qlmy9_1),.clk(gclk));
	jdff dff_A_O2HRP7rs9_1(.dout(w_dff_A_fHj8Qlmy9_1),.din(w_dff_A_O2HRP7rs9_1),.clk(gclk));
	jdff dff_A_Gm5PiSKX9_2(.dout(w_G953_0[2]),.din(w_dff_A_Gm5PiSKX9_2),.clk(gclk));
	jdff dff_A_mn6ZkUyT0_2(.dout(w_dff_A_Gm5PiSKX9_2),.din(w_dff_A_mn6ZkUyT0_2),.clk(gclk));
	jdff dff_A_tbhiNONq6_2(.dout(w_dff_A_mn6ZkUyT0_2),.din(w_dff_A_tbhiNONq6_2),.clk(gclk));
	jdff dff_A_B3td6LzI6_2(.dout(w_dff_A_tbhiNONq6_2),.din(w_dff_A_B3td6LzI6_2),.clk(gclk));
	jdff dff_A_tLjjikdm6_2(.dout(w_dff_A_B3td6LzI6_2),.din(w_dff_A_tLjjikdm6_2),.clk(gclk));
	jdff dff_A_V3aEJJsO6_2(.dout(w_dff_A_tLjjikdm6_2),.din(w_dff_A_V3aEJJsO6_2),.clk(gclk));
	jdff dff_A_toKElB6Y4_2(.dout(w_dff_A_V3aEJJsO6_2),.din(w_dff_A_toKElB6Y4_2),.clk(gclk));
	jdff dff_A_RPDo84dn2_2(.dout(w_dff_A_toKElB6Y4_2),.din(w_dff_A_RPDo84dn2_2),.clk(gclk));
	jdff dff_A_4yWKP1v25_2(.dout(w_dff_A_RPDo84dn2_2),.din(w_dff_A_4yWKP1v25_2),.clk(gclk));
	jdff dff_A_EMIIOYeM7_2(.dout(w_dff_A_4yWKP1v25_2),.din(w_dff_A_EMIIOYeM7_2),.clk(gclk));
	jdff dff_A_BJKAFMm76_2(.dout(w_dff_A_EMIIOYeM7_2),.din(w_dff_A_BJKAFMm76_2),.clk(gclk));
	jdff dff_A_gX385W5s1_2(.dout(w_dff_A_BJKAFMm76_2),.din(w_dff_A_gX385W5s1_2),.clk(gclk));
	jdff dff_A_ddUKeo2G2_2(.dout(w_dff_A_gX385W5s1_2),.din(w_dff_A_ddUKeo2G2_2),.clk(gclk));
	jdff dff_A_ylYDucCB8_0(.dout(w_G101_0[0]),.din(w_dff_A_ylYDucCB8_0),.clk(gclk));
	jdff dff_A_EKld3pcg0_0(.dout(w_dff_A_ylYDucCB8_0),.din(w_dff_A_EKld3pcg0_0),.clk(gclk));
	jdff dff_A_q0nHAXmV4_0(.dout(w_dff_A_EKld3pcg0_0),.din(w_dff_A_q0nHAXmV4_0),.clk(gclk));
	jdff dff_A_AmEHrhQV6_0(.dout(w_dff_A_q0nHAXmV4_0),.din(w_dff_A_AmEHrhQV6_0),.clk(gclk));
	jdff dff_A_VqRIrjjA9_0(.dout(w_dff_A_AmEHrhQV6_0),.din(w_dff_A_VqRIrjjA9_0),.clk(gclk));
	jdff dff_A_GwJqMgDY6_0(.dout(w_dff_A_VqRIrjjA9_0),.din(w_dff_A_GwJqMgDY6_0),.clk(gclk));
	jdff dff_A_EMfXk32e9_0(.dout(w_dff_A_GwJqMgDY6_0),.din(w_dff_A_EMfXk32e9_0),.clk(gclk));
	jdff dff_A_tumOYY1B4_0(.dout(w_dff_A_EMfXk32e9_0),.din(w_dff_A_tumOYY1B4_0),.clk(gclk));
	jdff dff_A_F4JAuFmx3_0(.dout(w_dff_A_tumOYY1B4_0),.din(w_dff_A_F4JAuFmx3_0),.clk(gclk));
	jdff dff_A_SPqektBu0_0(.dout(w_dff_A_F4JAuFmx3_0),.din(w_dff_A_SPqektBu0_0),.clk(gclk));
	jdff dff_B_IWk5oVRb7_3(.din(G101),.dout(w_dff_B_IWk5oVRb7_3),.clk(gclk));
	jdff dff_A_qveKPsB94_0(.dout(w_G119_0[0]),.din(w_dff_A_qveKPsB94_0),.clk(gclk));
	jdff dff_A_vL4OBC3h5_0(.dout(w_dff_A_qveKPsB94_0),.din(w_dff_A_vL4OBC3h5_0),.clk(gclk));
	jdff dff_A_Y3muUcoT4_0(.dout(w_dff_A_vL4OBC3h5_0),.din(w_dff_A_Y3muUcoT4_0),.clk(gclk));
	jdff dff_A_x2Bd3gdv0_0(.dout(w_dff_A_Y3muUcoT4_0),.din(w_dff_A_x2Bd3gdv0_0),.clk(gclk));
	jdff dff_A_AgN90Q0G7_0(.dout(w_dff_A_x2Bd3gdv0_0),.din(w_dff_A_AgN90Q0G7_0),.clk(gclk));
	jdff dff_A_LMaFAXdJ1_0(.dout(w_dff_A_AgN90Q0G7_0),.din(w_dff_A_LMaFAXdJ1_0),.clk(gclk));
	jdff dff_A_0QVct4Pr0_0(.dout(w_dff_A_LMaFAXdJ1_0),.din(w_dff_A_0QVct4Pr0_0),.clk(gclk));
	jdff dff_A_nWq8BmDO8_0(.dout(w_dff_A_0QVct4Pr0_0),.din(w_dff_A_nWq8BmDO8_0),.clk(gclk));
	jdff dff_A_rBOdxVvI0_0(.dout(w_dff_A_nWq8BmDO8_0),.din(w_dff_A_rBOdxVvI0_0),.clk(gclk));
	jdff dff_A_QRMLf8KU3_0(.dout(w_dff_A_rBOdxVvI0_0),.din(w_dff_A_QRMLf8KU3_0),.clk(gclk));
	jdff dff_A_lrpOe7On2_0(.dout(w_dff_A_QRMLf8KU3_0),.din(w_dff_A_lrpOe7On2_0),.clk(gclk));
	jdff dff_A_wOPgZHQT5_0(.dout(w_dff_A_lrpOe7On2_0),.din(w_dff_A_wOPgZHQT5_0),.clk(gclk));
	jdff dff_A_pGIcC5Nb1_0(.dout(w_G116_0[0]),.din(w_dff_A_pGIcC5Nb1_0),.clk(gclk));
	jdff dff_A_9Dj2fXD11_0(.dout(w_dff_A_pGIcC5Nb1_0),.din(w_dff_A_9Dj2fXD11_0),.clk(gclk));
	jdff dff_A_MWREZoIe4_0(.dout(w_dff_A_9Dj2fXD11_0),.din(w_dff_A_MWREZoIe4_0),.clk(gclk));
	jdff dff_A_xhKX1fZa1_0(.dout(w_dff_A_MWREZoIe4_0),.din(w_dff_A_xhKX1fZa1_0),.clk(gclk));
	jdff dff_A_5ZpvOOzI4_0(.dout(w_dff_A_xhKX1fZa1_0),.din(w_dff_A_5ZpvOOzI4_0),.clk(gclk));
	jdff dff_A_0F0hN5Xy2_0(.dout(w_dff_A_5ZpvOOzI4_0),.din(w_dff_A_0F0hN5Xy2_0),.clk(gclk));
	jdff dff_A_Nck09PbR6_0(.dout(w_dff_A_0F0hN5Xy2_0),.din(w_dff_A_Nck09PbR6_0),.clk(gclk));
	jdff dff_A_Q0GO04VI3_0(.dout(w_dff_A_Nck09PbR6_0),.din(w_dff_A_Q0GO04VI3_0),.clk(gclk));
	jdff dff_A_XfJSyxlP7_0(.dout(w_dff_A_Q0GO04VI3_0),.din(w_dff_A_XfJSyxlP7_0),.clk(gclk));
	jdff dff_A_Xx0hi9WI9_0(.dout(w_dff_A_XfJSyxlP7_0),.din(w_dff_A_Xx0hi9WI9_0),.clk(gclk));
	jdff dff_A_tyrBzHzI7_0(.dout(w_dff_A_Xx0hi9WI9_0),.din(w_dff_A_tyrBzHzI7_0),.clk(gclk));
	jdff dff_A_LJf4yOhf3_0(.dout(w_G113_0[0]),.din(w_dff_A_LJf4yOhf3_0),.clk(gclk));
	jdff dff_A_CSNq7BSX8_0(.dout(w_dff_A_LJf4yOhf3_0),.din(w_dff_A_CSNq7BSX8_0),.clk(gclk));
	jdff dff_A_QsWjfle73_0(.dout(w_dff_A_CSNq7BSX8_0),.din(w_dff_A_QsWjfle73_0),.clk(gclk));
	jdff dff_A_7JFzegV06_0(.dout(w_dff_A_QsWjfle73_0),.din(w_dff_A_7JFzegV06_0),.clk(gclk));
	jdff dff_A_EisgLbwD9_0(.dout(w_dff_A_7JFzegV06_0),.din(w_dff_A_EisgLbwD9_0),.clk(gclk));
	jdff dff_A_dkxi518c3_0(.dout(w_dff_A_EisgLbwD9_0),.din(w_dff_A_dkxi518c3_0),.clk(gclk));
	jdff dff_A_AmCo4Aej2_0(.dout(w_dff_A_dkxi518c3_0),.din(w_dff_A_AmCo4Aej2_0),.clk(gclk));
	jdff dff_A_W1qqONbB1_0(.dout(w_dff_A_AmCo4Aej2_0),.din(w_dff_A_W1qqONbB1_0),.clk(gclk));
	jdff dff_A_q1A0qZEl3_0(.dout(w_dff_A_W1qqONbB1_0),.din(w_dff_A_q1A0qZEl3_0),.clk(gclk));
	jdff dff_A_OutWcRG95_0(.dout(w_dff_A_q1A0qZEl3_0),.din(w_dff_A_OutWcRG95_0),.clk(gclk));
	jdff dff_A_Vz1GAtqw7_0(.dout(w_dff_A_OutWcRG95_0),.din(w_dff_A_Vz1GAtqw7_0),.clk(gclk));
	jdff dff_B_5VKQOKOj0_1(.din(n76),.dout(w_dff_B_5VKQOKOj0_1),.clk(gclk));
	jdff dff_A_tla3SoKu1_0(.dout(w_G146_0[0]),.din(w_dff_A_tla3SoKu1_0),.clk(gclk));
	jdff dff_A_wKtR7sIw7_0(.dout(w_dff_A_tla3SoKu1_0),.din(w_dff_A_wKtR7sIw7_0),.clk(gclk));
	jdff dff_A_PQ10YjKH9_0(.dout(w_dff_A_wKtR7sIw7_0),.din(w_dff_A_PQ10YjKH9_0),.clk(gclk));
	jdff dff_A_lGmpFOEn6_0(.dout(w_dff_A_PQ10YjKH9_0),.din(w_dff_A_lGmpFOEn6_0),.clk(gclk));
	jdff dff_A_xEvKF5tx7_0(.dout(w_dff_A_lGmpFOEn6_0),.din(w_dff_A_xEvKF5tx7_0),.clk(gclk));
	jdff dff_A_ocggoty87_0(.dout(w_dff_A_xEvKF5tx7_0),.din(w_dff_A_ocggoty87_0),.clk(gclk));
	jdff dff_A_uAEfHOzT4_0(.dout(w_dff_A_ocggoty87_0),.din(w_dff_A_uAEfHOzT4_0),.clk(gclk));
	jdff dff_A_gS0TxkNc8_0(.dout(w_dff_A_uAEfHOzT4_0),.din(w_dff_A_gS0TxkNc8_0),.clk(gclk));
	jdff dff_A_rtLv1IwE6_0(.dout(w_dff_A_gS0TxkNc8_0),.din(w_dff_A_rtLv1IwE6_0),.clk(gclk));
	jdff dff_A_U7aYvUsJ2_0(.dout(w_dff_A_rtLv1IwE6_0),.din(w_dff_A_U7aYvUsJ2_0),.clk(gclk));
	jdff dff_A_y2O5yMa80_0(.dout(w_dff_A_U7aYvUsJ2_0),.din(w_dff_A_y2O5yMa80_0),.clk(gclk));
	jdff dff_A_IqzNrTTb5_0(.dout(w_dff_A_y2O5yMa80_0),.din(w_dff_A_IqzNrTTb5_0),.clk(gclk));
	jdff dff_A_uNgtkKv92_1(.dout(w_G143_0[1]),.din(w_dff_A_uNgtkKv92_1),.clk(gclk));
	jdff dff_A_WZhKdfIf8_1(.dout(w_dff_A_uNgtkKv92_1),.din(w_dff_A_WZhKdfIf8_1),.clk(gclk));
	jdff dff_A_FG0UcSXU9_1(.dout(w_dff_A_WZhKdfIf8_1),.din(w_dff_A_FG0UcSXU9_1),.clk(gclk));
	jdff dff_A_hGLNjpR19_1(.dout(w_dff_A_FG0UcSXU9_1),.din(w_dff_A_hGLNjpR19_1),.clk(gclk));
	jdff dff_A_LeXS26RJ4_1(.dout(w_dff_A_hGLNjpR19_1),.din(w_dff_A_LeXS26RJ4_1),.clk(gclk));
	jdff dff_A_HDM9xbZg1_1(.dout(w_dff_A_LeXS26RJ4_1),.din(w_dff_A_HDM9xbZg1_1),.clk(gclk));
	jdff dff_A_ThyI4IAu2_1(.dout(w_dff_A_HDM9xbZg1_1),.din(w_dff_A_ThyI4IAu2_1),.clk(gclk));
	jdff dff_A_leaLF7tD6_1(.dout(w_dff_A_ThyI4IAu2_1),.din(w_dff_A_leaLF7tD6_1),.clk(gclk));
	jdff dff_A_Ung9iAtf2_1(.dout(w_dff_A_leaLF7tD6_1),.din(w_dff_A_Ung9iAtf2_1),.clk(gclk));
	jdff dff_A_bE9whqp88_1(.dout(w_dff_A_Ung9iAtf2_1),.din(w_dff_A_bE9whqp88_1),.clk(gclk));
	jdff dff_A_McHXRgtX7_1(.dout(w_dff_A_bE9whqp88_1),.din(w_dff_A_McHXRgtX7_1),.clk(gclk));
	jdff dff_A_P79p6jqT7_2(.dout(w_G143_0[2]),.din(w_dff_A_P79p6jqT7_2),.clk(gclk));
	jdff dff_A_JRAGx0Nq6_0(.dout(w_G128_1[0]),.din(w_dff_A_JRAGx0Nq6_0),.clk(gclk));
	jdff dff_A_ff2iXvSU5_1(.dout(w_G128_0[1]),.din(w_dff_A_ff2iXvSU5_1),.clk(gclk));
	jdff dff_A_XazWRSaf1_1(.dout(w_dff_A_ff2iXvSU5_1),.din(w_dff_A_XazWRSaf1_1),.clk(gclk));
	jdff dff_A_DzTql2697_1(.dout(w_dff_A_XazWRSaf1_1),.din(w_dff_A_DzTql2697_1),.clk(gclk));
	jdff dff_A_mFRkDpYh1_1(.dout(w_dff_A_DzTql2697_1),.din(w_dff_A_mFRkDpYh1_1),.clk(gclk));
	jdff dff_A_5JyVBdS30_1(.dout(w_dff_A_mFRkDpYh1_1),.din(w_dff_A_5JyVBdS30_1),.clk(gclk));
	jdff dff_A_FgbG6MNU9_1(.dout(w_dff_A_5JyVBdS30_1),.din(w_dff_A_FgbG6MNU9_1),.clk(gclk));
	jdff dff_A_abkQUR1R5_1(.dout(w_dff_A_FgbG6MNU9_1),.din(w_dff_A_abkQUR1R5_1),.clk(gclk));
	jdff dff_A_zbqQPR770_1(.dout(w_dff_A_abkQUR1R5_1),.din(w_dff_A_zbqQPR770_1),.clk(gclk));
	jdff dff_A_PrTlXV8E9_1(.dout(w_dff_A_zbqQPR770_1),.din(w_dff_A_PrTlXV8E9_1),.clk(gclk));
	jdff dff_A_xYyJJ0060_1(.dout(w_dff_A_PrTlXV8E9_1),.din(w_dff_A_xYyJJ0060_1),.clk(gclk));
	jdff dff_A_MwfhDWU89_1(.dout(w_dff_A_xYyJJ0060_1),.din(w_dff_A_MwfhDWU89_1),.clk(gclk));
	jdff dff_A_Ieji7Bl78_1(.dout(w_dff_A_MwfhDWU89_1),.din(w_dff_A_Ieji7Bl78_1),.clk(gclk));
	jdff dff_A_B1IMyYbE1_1(.dout(w_n77_0[1]),.din(w_dff_A_B1IMyYbE1_1),.clk(gclk));
	jdff dff_A_VGCYIe8S6_0(.dout(w_G131_0[0]),.din(w_dff_A_VGCYIe8S6_0),.clk(gclk));
	jdff dff_A_ZvLVeX474_0(.dout(w_dff_A_VGCYIe8S6_0),.din(w_dff_A_ZvLVeX474_0),.clk(gclk));
	jdff dff_A_s0APKqXo3_0(.dout(w_dff_A_ZvLVeX474_0),.din(w_dff_A_s0APKqXo3_0),.clk(gclk));
	jdff dff_A_3GO2tmR13_0(.dout(w_dff_A_s0APKqXo3_0),.din(w_dff_A_3GO2tmR13_0),.clk(gclk));
	jdff dff_A_imf2LaAW7_0(.dout(w_dff_A_3GO2tmR13_0),.din(w_dff_A_imf2LaAW7_0),.clk(gclk));
	jdff dff_A_hdFgw2bm0_0(.dout(w_dff_A_imf2LaAW7_0),.din(w_dff_A_hdFgw2bm0_0),.clk(gclk));
	jdff dff_A_wiZeESvy6_0(.dout(w_dff_A_hdFgw2bm0_0),.din(w_dff_A_wiZeESvy6_0),.clk(gclk));
	jdff dff_A_LStv0DhR0_0(.dout(w_dff_A_wiZeESvy6_0),.din(w_dff_A_LStv0DhR0_0),.clk(gclk));
	jdff dff_A_LL4W1OTT3_0(.dout(w_dff_A_LStv0DhR0_0),.din(w_dff_A_LL4W1OTT3_0),.clk(gclk));
	jdff dff_A_uCchKFyL9_0(.dout(w_dff_A_LL4W1OTT3_0),.din(w_dff_A_uCchKFyL9_0),.clk(gclk));
	jdff dff_A_NvTiZtab6_0(.dout(w_dff_A_uCchKFyL9_0),.din(w_dff_A_NvTiZtab6_0),.clk(gclk));
	jdff dff_A_3hDjbJ9a1_0(.dout(w_G137_0[0]),.din(w_dff_A_3hDjbJ9a1_0),.clk(gclk));
	jdff dff_A_zgTcLVob3_0(.dout(w_dff_A_3hDjbJ9a1_0),.din(w_dff_A_zgTcLVob3_0),.clk(gclk));
	jdff dff_A_RS764XpV0_0(.dout(w_dff_A_zgTcLVob3_0),.din(w_dff_A_RS764XpV0_0),.clk(gclk));
	jdff dff_A_s1PP3tVz0_0(.dout(w_dff_A_RS764XpV0_0),.din(w_dff_A_s1PP3tVz0_0),.clk(gclk));
	jdff dff_A_h1DWEH6k2_0(.dout(w_dff_A_s1PP3tVz0_0),.din(w_dff_A_h1DWEH6k2_0),.clk(gclk));
	jdff dff_A_xyaU7Rad7_0(.dout(w_dff_A_h1DWEH6k2_0),.din(w_dff_A_xyaU7Rad7_0),.clk(gclk));
	jdff dff_A_k3ndl7Y64_0(.dout(w_dff_A_xyaU7Rad7_0),.din(w_dff_A_k3ndl7Y64_0),.clk(gclk));
	jdff dff_A_tb5KwVXj3_0(.dout(w_dff_A_k3ndl7Y64_0),.din(w_dff_A_tb5KwVXj3_0),.clk(gclk));
	jdff dff_A_XvgoQNPf8_0(.dout(w_dff_A_tb5KwVXj3_0),.din(w_dff_A_XvgoQNPf8_0),.clk(gclk));
	jdff dff_A_5iRqOBHK5_0(.dout(w_dff_A_XvgoQNPf8_0),.din(w_dff_A_5iRqOBHK5_0),.clk(gclk));
	jdff dff_A_VfRoeoli6_0(.dout(w_dff_A_5iRqOBHK5_0),.din(w_dff_A_VfRoeoli6_0),.clk(gclk));
	jdff dff_A_FNCOujbh5_2(.dout(w_G137_0[2]),.din(w_dff_A_FNCOujbh5_2),.clk(gclk));
	jdff dff_A_seMvB0Zz0_2(.dout(w_dff_A_FNCOujbh5_2),.din(w_dff_A_seMvB0Zz0_2),.clk(gclk));
	jdff dff_B_Yb2Y004C3_3(.din(G137),.dout(w_dff_B_Yb2Y004C3_3),.clk(gclk));
	jdff dff_A_WPSsL5Ei1_0(.dout(w_G134_0[0]),.din(w_dff_A_WPSsL5Ei1_0),.clk(gclk));
	jdff dff_A_5OzUNPNt7_0(.dout(w_dff_A_WPSsL5Ei1_0),.din(w_dff_A_5OzUNPNt7_0),.clk(gclk));
	jdff dff_A_q6HbcHHl6_0(.dout(w_dff_A_5OzUNPNt7_0),.din(w_dff_A_q6HbcHHl6_0),.clk(gclk));
	jdff dff_A_xKJatb3f9_0(.dout(w_dff_A_q6HbcHHl6_0),.din(w_dff_A_xKJatb3f9_0),.clk(gclk));
	jdff dff_A_OFPz05A60_0(.dout(w_dff_A_xKJatb3f9_0),.din(w_dff_A_OFPz05A60_0),.clk(gclk));
	jdff dff_A_60LGZOKg3_0(.dout(w_dff_A_OFPz05A60_0),.din(w_dff_A_60LGZOKg3_0),.clk(gclk));
	jdff dff_A_Y07P36u01_0(.dout(w_dff_A_60LGZOKg3_0),.din(w_dff_A_Y07P36u01_0),.clk(gclk));
	jdff dff_A_CWvdlzJN9_0(.dout(w_dff_A_Y07P36u01_0),.din(w_dff_A_CWvdlzJN9_0),.clk(gclk));
	jdff dff_A_bnBL7SIz9_0(.dout(w_dff_A_CWvdlzJN9_0),.din(w_dff_A_bnBL7SIz9_0),.clk(gclk));
	jdff dff_A_ZwmTRFwx9_0(.dout(w_dff_A_bnBL7SIz9_0),.din(w_dff_A_ZwmTRFwx9_0),.clk(gclk));
	jdff dff_A_LdSlPXbY0_0(.dout(w_dff_A_ZwmTRFwx9_0),.din(w_dff_A_LdSlPXbY0_0),.clk(gclk));
endmodule

