// Benchmark "top" written by ABC on Wed May 27 23:34:26 2020

module top ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , a16 ,
    a17 , a18 , a19 , a20 , a21 , a22 , a23 , a24 ,
    a25 , a26 , a27 , a28 , a29 , a30 , a31 , a32 ,
    a33 , a34 , a35 , a36 , a37 , a38 , a39 , a40 ,
    a41 , a42 , a43 , a44 , a45 , a46 , a47 , a48 ,
    a49 , a50 , a51 , a52 , a53 , a54 , a55 , a56 ,
    a57 , a58 , a59 , a60 , a61 , a62 , a63 , a64 ,
    a65 , a66 , a67 , a68 , a69 , a70 , a71 , a72 ,
    a73 , a74 , a75 , a76 , a77 , a78 , a79 , a80 ,
    a81 , a82 , a83 , a84 , a85 , a86 , a87 , a88 ,
    a89 , a90 , a91 , a92 , a93 , a94 , a95 , a96 ,
    a97 , a98 , a99 , a100 , a101 , a102 , a103 ,
    a104 , a105 , a106 , a107 , a108 , a109 , a110 ,
    a111 , a112 , a113 , a114 , a115 , a116 , a117 ,
    a118 , a119 , a120 , a121 , a122 , a123 , a124 ,
    a125 , a126 , a127 , shift0 , shift1 , shift2 ,
    shift3 , shift4 , shift5 , shift6 ,
    result0 , result1 , result2 , result3 , result4 ,
    result5 , result6 , result7 , result8 , result9 ,
    result10 , result11 , result12 , result13 , result14 ,
    result15 , result16 , result17 , result18 , result19 ,
    result20 , result21 , result22 , result23 , result24 ,
    result25 , result26 , result27 , result28 , result29 ,
    result30 , result31 , result32 , result33 , result34 ,
    result35 , result36 , result37 , result38 , result39 ,
    result40 , result41 , result42 , result43 , result44 ,
    result45 , result46 , result47 , result48 , result49 ,
    result50 , result51 , result52 , result53 , result54 ,
    result55 , result56 , result57 , result58 , result59 ,
    result60 , result61 , result62 , result63 , result64 ,
    result65 , result66 , result67 , result68 , result69 ,
    result70 , result71 , result72 , result73 , result74 ,
    result75 , result76 , result77 , result78 , result79 ,
    result80 , result81 , result82 , result83 , result84 ,
    result85 , result86 , result87 , result88 , result89 ,
    result90 , result91 , result92 , result93 , result94 ,
    result95 , result96 , result97 , result98 , result99 ,
    result100 , result101 , result102 , result103 ,
    result104 , result105 , result106 , result107 ,
    result108 , result109 , result110 , result111 ,
    result112 , result113 , result114 , result115 ,
    result116 , result117 , result118 , result119 ,
    result120 , result121 , result122 , result123 ,
    result124 , result125 , result126 , result127   );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    a16 , a17 , a18 , a19 , a20 , a21 , a22 , a23 ,
    a24 , a25 , a26 , a27 , a28 , a29 , a30 , a31 ,
    a32 , a33 , a34 , a35 , a36 , a37 , a38 , a39 ,
    a40 , a41 , a42 , a43 , a44 , a45 , a46 , a47 ,
    a48 , a49 , a50 , a51 , a52 , a53 , a54 , a55 ,
    a56 , a57 , a58 , a59 , a60 , a61 , a62 , a63 ,
    a64 , a65 , a66 , a67 , a68 , a69 , a70 , a71 ,
    a72 , a73 , a74 , a75 , a76 , a77 , a78 , a79 ,
    a80 , a81 , a82 , a83 , a84 , a85 , a86 , a87 ,
    a88 , a89 , a90 , a91 , a92 , a93 , a94 , a95 ,
    a96 , a97 , a98 , a99 , a100 , a101 , a102 ,
    a103 , a104 , a105 , a106 , a107 , a108 , a109 ,
    a110 , a111 , a112 , a113 , a114 , a115 , a116 ,
    a117 , a118 , a119 , a120 , a121 , a122 , a123 ,
    a124 , a125 , a126 , a127 , shift0 , shift1 ,
    shift2 , shift3 , shift4 , shift5 , shift6 ;
  output result0 , result1 , result2 , result3 , result4 ,
    result5 , result6 , result7 , result8 , result9 ,
    result10 , result11 , result12 , result13 , result14 ,
    result15 , result16 , result17 , result18 , result19 ,
    result20 , result21 , result22 , result23 , result24 ,
    result25 , result26 , result27 , result28 , result29 ,
    result30 , result31 , result32 , result33 , result34 ,
    result35 , result36 , result37 , result38 , result39 ,
    result40 , result41 , result42 , result43 , result44 ,
    result45 , result46 , result47 , result48 , result49 ,
    result50 , result51 , result52 , result53 , result54 ,
    result55 , result56 , result57 , result58 , result59 ,
    result60 , result61 , result62 , result63 , result64 ,
    result65 , result66 , result67 , result68 , result69 ,
    result70 , result71 , result72 , result73 , result74 ,
    result75 , result76 , result77 , result78 , result79 ,
    result80 , result81 , result82 , result83 , result84 ,
    result85 , result86 , result87 , result88 , result89 ,
    result90 , result91 , result92 , result93 , result94 ,
    result95 , result96 , result97 , result98 , result99 ,
    result100 , result101 , result102 , result103 ,
    result104 , result105 , result106 , result107 ,
    result108 , result109 , result110 , result111 ,
    result112 , result113 , result114 , result115 ,
    result116 , result117 , result118 , result119 ,
    result120 , result121 , result122 , result123 ,
    result124 , result125 , result126 , result127 ;
  wire n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
    n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
    n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
    n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
    n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
    n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
    n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
    n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
    n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
    n2339, n2340, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
    n2442, n2443, n2444, n2445, n2446, n2447, n2449, n2450, n2451, n2452,
    n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2823, n2824,
    n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
    n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
    n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3095, n3096, n3097, n3098, n3099, n3100,
    n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
    n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
    n3143, n3144, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
    n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3231, n3232, n3234, n3235, n3237, n3238, n3240, n3241,
    n3243, n3244, n3246, n3247, n3249, n3250, n3252, n3253, n3255, n3256,
    n3258, n3259, n3261, n3262, n3264, n3265, n3267, n3268, n3270, n3271,
    n3273, n3274, n3276, n3277, n3279, n3280, n3282, n3283, n3285, n3286,
    n3288, n3289, n3291, n3292, n3294, n3295, n3297, n3298, n3300, n3301,
    n3303, n3304, n3306, n3307, n3309, n3310, n3312, n3313, n3315, n3316,
    n3318, n3319, n3321, n3322, n3324, n3325, n3327, n3328, n3330, n3331,
    n3333, n3334, n3336, n3337, n3339, n3340, n3342, n3343, n3345, n3346,
    n3348, n3349, n3351, n3352, n3354, n3355, n3357, n3358, n3360, n3361,
    n3363, n3364, n3366, n3367, n3369, n3370, n3372, n3373, n3375, n3376,
    n3378, n3379, n3381, n3382, n3384, n3385, n3387, n3388, n3390, n3391,
    n3393, n3394, n3396, n3397, n3399, n3400, n3402, n3403, n3405, n3406,
    n3408, n3409, n3411, n3412, n3414, n3415, n3417, n3418, n3420, n3421;
  jnot g0000(.din(shift6 ), .dout(n263));
  jnot g0001(.din(shift2 ), .dout(n264));
  jnot g0002(.din(shift3 ), .dout(n265));
  jand g0003(.dina(n265), .dinb(n264), .dout(n266));
  jand g0004(.dina(shift0 ), .dinb(a79 ), .dout(n267));
  jor  g0005(.dina(n267), .dinb(shift1 ), .dout(n268));
  jnot g0006(.din(shift1 ), .dout(n269));
  jnot g0007(.din(shift0 ), .dout(n270));
  jand g0008(.dina(n270), .dinb(a78 ), .dout(n271));
  jor  g0009(.dina(n271), .dinb(n269), .dout(n272));
  jand g0010(.dina(n272), .dinb(n268), .dout(n273));
  jand g0011(.dina(shift0 ), .dinb(a77 ), .dout(n274));
  jand g0012(.dina(n274), .dinb(shift1 ), .dout(n275));
  jand g0013(.dina(n270), .dinb(a80 ), .dout(n276));
  jand g0014(.dina(n276), .dinb(n269), .dout(n277));
  jor  g0015(.dina(n277), .dinb(n275), .dout(n278));
  jor  g0016(.dina(n278), .dinb(n273), .dout(n279));
  jand g0017(.dina(n279), .dinb(n266), .dout(n280));
  jand g0018(.dina(shift3 ), .dinb(n264), .dout(n281));
  jand g0019(.dina(shift0 ), .dinb(a71 ), .dout(n282));
  jor  g0020(.dina(n282), .dinb(shift1 ), .dout(n283));
  jand g0021(.dina(n270), .dinb(a70 ), .dout(n284));
  jor  g0022(.dina(n284), .dinb(n269), .dout(n285));
  jand g0023(.dina(n285), .dinb(n283), .dout(n286));
  jand g0024(.dina(shift0 ), .dinb(a69 ), .dout(n287));
  jand g0025(.dina(n287), .dinb(shift1 ), .dout(n288));
  jand g0026(.dina(n270), .dinb(a72 ), .dout(n289));
  jand g0027(.dina(n289), .dinb(n269), .dout(n290));
  jor  g0028(.dina(n290), .dinb(n288), .dout(n291));
  jor  g0029(.dina(n291), .dinb(n286), .dout(n292));
  jand g0030(.dina(n292), .dinb(n281), .dout(n293));
  jor  g0031(.dina(n293), .dinb(n280), .dout(n294));
  jand g0032(.dina(n265), .dinb(shift2 ), .dout(n295));
  jand g0033(.dina(shift0 ), .dinb(a75 ), .dout(n296));
  jor  g0034(.dina(n296), .dinb(shift1 ), .dout(n297));
  jand g0035(.dina(n270), .dinb(a74 ), .dout(n298));
  jor  g0036(.dina(n298), .dinb(n269), .dout(n299));
  jand g0037(.dina(n299), .dinb(n297), .dout(n300));
  jand g0038(.dina(shift0 ), .dinb(a73 ), .dout(n301));
  jand g0039(.dina(n301), .dinb(shift1 ), .dout(n302));
  jand g0040(.dina(n270), .dinb(a76 ), .dout(n303));
  jand g0041(.dina(n303), .dinb(n269), .dout(n304));
  jor  g0042(.dina(n304), .dinb(n302), .dout(n305));
  jor  g0043(.dina(n305), .dinb(n300), .dout(n306));
  jand g0044(.dina(n306), .dinb(n295), .dout(n307));
  jand g0045(.dina(shift3 ), .dinb(shift2 ), .dout(n308));
  jand g0046(.dina(shift0 ), .dinb(a67 ), .dout(n309));
  jor  g0047(.dina(n309), .dinb(shift1 ), .dout(n310));
  jand g0048(.dina(n270), .dinb(a66 ), .dout(n311));
  jor  g0049(.dina(n311), .dinb(n269), .dout(n312));
  jand g0050(.dina(n312), .dinb(n310), .dout(n313));
  jand g0051(.dina(shift0 ), .dinb(a65 ), .dout(n314));
  jand g0052(.dina(n314), .dinb(shift1 ), .dout(n315));
  jand g0053(.dina(n270), .dinb(a68 ), .dout(n316));
  jand g0054(.dina(n316), .dinb(n269), .dout(n317));
  jor  g0055(.dina(n317), .dinb(n315), .dout(n318));
  jor  g0056(.dina(n318), .dinb(n313), .dout(n319));
  jand g0057(.dina(n319), .dinb(n308), .dout(n320));
  jor  g0058(.dina(n320), .dinb(n307), .dout(n321));
  jor  g0059(.dina(n321), .dinb(n294), .dout(n322));
  jand g0060(.dina(shift5 ), .dinb(shift4 ), .dout(n323));
  jand g0061(.dina(n323), .dinb(n322), .dout(n324));
  jand g0062(.dina(shift0 ), .dinb(a111 ), .dout(n325));
  jor  g0063(.dina(n325), .dinb(shift1 ), .dout(n326));
  jand g0064(.dina(n270), .dinb(a110 ), .dout(n327));
  jor  g0065(.dina(n327), .dinb(n269), .dout(n328));
  jand g0066(.dina(n328), .dinb(n326), .dout(n329));
  jand g0067(.dina(shift0 ), .dinb(a109 ), .dout(n330));
  jand g0068(.dina(n330), .dinb(shift1 ), .dout(n331));
  jand g0069(.dina(n270), .dinb(a112 ), .dout(n332));
  jand g0070(.dina(n332), .dinb(n269), .dout(n333));
  jor  g0071(.dina(n333), .dinb(n331), .dout(n334));
  jor  g0072(.dina(n334), .dinb(n329), .dout(n335));
  jand g0073(.dina(n335), .dinb(n266), .dout(n336));
  jand g0074(.dina(shift0 ), .dinb(a103 ), .dout(n337));
  jor  g0075(.dina(n337), .dinb(shift1 ), .dout(n338));
  jand g0076(.dina(n270), .dinb(a102 ), .dout(n339));
  jor  g0077(.dina(n339), .dinb(n269), .dout(n340));
  jand g0078(.dina(n340), .dinb(n338), .dout(n341));
  jand g0079(.dina(shift0 ), .dinb(a101 ), .dout(n342));
  jand g0080(.dina(n342), .dinb(shift1 ), .dout(n343));
  jand g0081(.dina(n270), .dinb(a104 ), .dout(n344));
  jand g0082(.dina(n344), .dinb(n269), .dout(n345));
  jor  g0083(.dina(n345), .dinb(n343), .dout(n346));
  jor  g0084(.dina(n346), .dinb(n341), .dout(n347));
  jand g0085(.dina(n347), .dinb(n281), .dout(n348));
  jor  g0086(.dina(n348), .dinb(n336), .dout(n349));
  jand g0087(.dina(shift0 ), .dinb(a107 ), .dout(n350));
  jor  g0088(.dina(n350), .dinb(shift1 ), .dout(n351));
  jand g0089(.dina(n270), .dinb(a106 ), .dout(n352));
  jor  g0090(.dina(n352), .dinb(n269), .dout(n353));
  jand g0091(.dina(n353), .dinb(n351), .dout(n354));
  jand g0092(.dina(shift0 ), .dinb(a105 ), .dout(n355));
  jand g0093(.dina(n355), .dinb(shift1 ), .dout(n356));
  jand g0094(.dina(n270), .dinb(a108 ), .dout(n357));
  jand g0095(.dina(n357), .dinb(n269), .dout(n358));
  jor  g0096(.dina(n358), .dinb(n356), .dout(n359));
  jor  g0097(.dina(n359), .dinb(n354), .dout(n360));
  jand g0098(.dina(n360), .dinb(n295), .dout(n361));
  jand g0099(.dina(shift0 ), .dinb(a99 ), .dout(n362));
  jor  g0100(.dina(n362), .dinb(shift1 ), .dout(n363));
  jand g0101(.dina(n270), .dinb(a98 ), .dout(n364));
  jor  g0102(.dina(n364), .dinb(n269), .dout(n365));
  jand g0103(.dina(n365), .dinb(n363), .dout(n366));
  jand g0104(.dina(shift0 ), .dinb(a97 ), .dout(n367));
  jand g0105(.dina(n367), .dinb(shift1 ), .dout(n368));
  jand g0106(.dina(n270), .dinb(a100 ), .dout(n369));
  jand g0107(.dina(n369), .dinb(n269), .dout(n370));
  jor  g0108(.dina(n370), .dinb(n368), .dout(n371));
  jor  g0109(.dina(n371), .dinb(n366), .dout(n372));
  jand g0110(.dina(n372), .dinb(n308), .dout(n373));
  jor  g0111(.dina(n373), .dinb(n361), .dout(n374));
  jor  g0112(.dina(n374), .dinb(n349), .dout(n375));
  jnot g0113(.din(shift5 ), .dout(n376));
  jand g0114(.dina(n376), .dinb(shift4 ), .dout(n377));
  jand g0115(.dina(n377), .dinb(n375), .dout(n378));
  jor  g0116(.dina(n378), .dinb(n324), .dout(n379));
  jand g0117(.dina(shift0 ), .dinb(a95 ), .dout(n380));
  jor  g0118(.dina(n380), .dinb(shift1 ), .dout(n381));
  jand g0119(.dina(n270), .dinb(a94 ), .dout(n382));
  jor  g0120(.dina(n382), .dinb(n269), .dout(n383));
  jand g0121(.dina(n383), .dinb(n381), .dout(n384));
  jand g0122(.dina(shift0 ), .dinb(a93 ), .dout(n385));
  jand g0123(.dina(n385), .dinb(shift1 ), .dout(n386));
  jand g0124(.dina(n270), .dinb(a96 ), .dout(n387));
  jand g0125(.dina(n387), .dinb(n269), .dout(n388));
  jor  g0126(.dina(n388), .dinb(n386), .dout(n389));
  jor  g0127(.dina(n389), .dinb(n384), .dout(n390));
  jand g0128(.dina(n390), .dinb(n266), .dout(n391));
  jand g0129(.dina(shift0 ), .dinb(a87 ), .dout(n392));
  jor  g0130(.dina(n392), .dinb(shift1 ), .dout(n393));
  jand g0131(.dina(n270), .dinb(a86 ), .dout(n394));
  jor  g0132(.dina(n394), .dinb(n269), .dout(n395));
  jand g0133(.dina(n395), .dinb(n393), .dout(n396));
  jand g0134(.dina(shift0 ), .dinb(a85 ), .dout(n397));
  jand g0135(.dina(n397), .dinb(shift1 ), .dout(n398));
  jand g0136(.dina(n270), .dinb(a88 ), .dout(n399));
  jand g0137(.dina(n399), .dinb(n269), .dout(n400));
  jor  g0138(.dina(n400), .dinb(n398), .dout(n401));
  jor  g0139(.dina(n401), .dinb(n396), .dout(n402));
  jand g0140(.dina(n402), .dinb(n281), .dout(n403));
  jor  g0141(.dina(n403), .dinb(n391), .dout(n404));
  jand g0142(.dina(shift0 ), .dinb(a91 ), .dout(n405));
  jor  g0143(.dina(n405), .dinb(shift1 ), .dout(n406));
  jand g0144(.dina(n270), .dinb(a90 ), .dout(n407));
  jor  g0145(.dina(n407), .dinb(n269), .dout(n408));
  jand g0146(.dina(n408), .dinb(n406), .dout(n409));
  jand g0147(.dina(shift0 ), .dinb(a89 ), .dout(n410));
  jand g0148(.dina(n410), .dinb(shift1 ), .dout(n411));
  jand g0149(.dina(n270), .dinb(a92 ), .dout(n412));
  jand g0150(.dina(n412), .dinb(n269), .dout(n413));
  jor  g0151(.dina(n413), .dinb(n411), .dout(n414));
  jor  g0152(.dina(n414), .dinb(n409), .dout(n415));
  jand g0153(.dina(n415), .dinb(n295), .dout(n416));
  jand g0154(.dina(shift0 ), .dinb(a83 ), .dout(n417));
  jor  g0155(.dina(n417), .dinb(shift1 ), .dout(n418));
  jand g0156(.dina(n270), .dinb(a82 ), .dout(n419));
  jor  g0157(.dina(n419), .dinb(n269), .dout(n420));
  jand g0158(.dina(n420), .dinb(n418), .dout(n421));
  jand g0159(.dina(shift0 ), .dinb(a81 ), .dout(n422));
  jand g0160(.dina(n422), .dinb(shift1 ), .dout(n423));
  jand g0161(.dina(n270), .dinb(a84 ), .dout(n424));
  jand g0162(.dina(n424), .dinb(n269), .dout(n425));
  jor  g0163(.dina(n425), .dinb(n423), .dout(n426));
  jor  g0164(.dina(n426), .dinb(n421), .dout(n427));
  jand g0165(.dina(n427), .dinb(n308), .dout(n428));
  jor  g0166(.dina(n428), .dinb(n416), .dout(n429));
  jor  g0167(.dina(n429), .dinb(n404), .dout(n430));
  jnot g0168(.din(shift4 ), .dout(n431));
  jand g0169(.dina(shift5 ), .dinb(n431), .dout(n432));
  jand g0170(.dina(n432), .dinb(n430), .dout(n433));
  jand g0171(.dina(shift0 ), .dinb(a127 ), .dout(n434));
  jor  g0172(.dina(n434), .dinb(shift1 ), .dout(n435));
  jand g0173(.dina(n270), .dinb(a126 ), .dout(n436));
  jor  g0174(.dina(n436), .dinb(n269), .dout(n437));
  jand g0175(.dina(n437), .dinb(n435), .dout(n438));
  jand g0176(.dina(shift0 ), .dinb(a125 ), .dout(n439));
  jand g0177(.dina(n439), .dinb(shift1 ), .dout(n440));
  jand g0178(.dina(n270), .dinb(a0 ), .dout(n441));
  jand g0179(.dina(n441), .dinb(n269), .dout(n442));
  jor  g0180(.dina(n442), .dinb(n440), .dout(n443));
  jor  g0181(.dina(n443), .dinb(n438), .dout(n444));
  jand g0182(.dina(n444), .dinb(n266), .dout(n445));
  jand g0183(.dina(shift0 ), .dinb(a119 ), .dout(n446));
  jor  g0184(.dina(n446), .dinb(shift1 ), .dout(n447));
  jand g0185(.dina(n270), .dinb(a118 ), .dout(n448));
  jor  g0186(.dina(n448), .dinb(n269), .dout(n449));
  jand g0187(.dina(n449), .dinb(n447), .dout(n450));
  jand g0188(.dina(shift0 ), .dinb(a117 ), .dout(n451));
  jand g0189(.dina(n451), .dinb(shift1 ), .dout(n452));
  jand g0190(.dina(n270), .dinb(a120 ), .dout(n453));
  jand g0191(.dina(n453), .dinb(n269), .dout(n454));
  jor  g0192(.dina(n454), .dinb(n452), .dout(n455));
  jor  g0193(.dina(n455), .dinb(n450), .dout(n456));
  jand g0194(.dina(n456), .dinb(n281), .dout(n457));
  jor  g0195(.dina(n457), .dinb(n445), .dout(n458));
  jand g0196(.dina(shift0 ), .dinb(a123 ), .dout(n459));
  jor  g0197(.dina(n459), .dinb(shift1 ), .dout(n460));
  jand g0198(.dina(n270), .dinb(a122 ), .dout(n461));
  jor  g0199(.dina(n461), .dinb(n269), .dout(n462));
  jand g0200(.dina(n462), .dinb(n460), .dout(n463));
  jand g0201(.dina(shift0 ), .dinb(a121 ), .dout(n464));
  jand g0202(.dina(n464), .dinb(shift1 ), .dout(n465));
  jand g0203(.dina(n270), .dinb(a124 ), .dout(n466));
  jand g0204(.dina(n466), .dinb(n269), .dout(n467));
  jor  g0205(.dina(n467), .dinb(n465), .dout(n468));
  jor  g0206(.dina(n468), .dinb(n463), .dout(n469));
  jand g0207(.dina(n469), .dinb(n295), .dout(n470));
  jand g0208(.dina(shift0 ), .dinb(a115 ), .dout(n471));
  jor  g0209(.dina(n471), .dinb(shift1 ), .dout(n472));
  jand g0210(.dina(n270), .dinb(a114 ), .dout(n473));
  jor  g0211(.dina(n473), .dinb(n269), .dout(n474));
  jand g0212(.dina(n474), .dinb(n472), .dout(n475));
  jand g0213(.dina(shift0 ), .dinb(a113 ), .dout(n476));
  jand g0214(.dina(n476), .dinb(shift1 ), .dout(n477));
  jand g0215(.dina(n270), .dinb(a116 ), .dout(n478));
  jand g0216(.dina(n478), .dinb(n269), .dout(n479));
  jor  g0217(.dina(n479), .dinb(n477), .dout(n480));
  jor  g0218(.dina(n480), .dinb(n475), .dout(n481));
  jand g0219(.dina(n481), .dinb(n308), .dout(n482));
  jor  g0220(.dina(n482), .dinb(n470), .dout(n483));
  jor  g0221(.dina(n483), .dinb(n458), .dout(n484));
  jand g0222(.dina(n376), .dinb(n431), .dout(n485));
  jand g0223(.dina(n485), .dinb(n484), .dout(n486));
  jor  g0224(.dina(n486), .dinb(n433), .dout(n487));
  jor  g0225(.dina(n487), .dinb(n379), .dout(n488));
  jand g0226(.dina(n488), .dinb(n263), .dout(n489));
  jand g0227(.dina(shift0 ), .dinb(a15 ), .dout(n490));
  jor  g0228(.dina(n490), .dinb(shift1 ), .dout(n491));
  jand g0229(.dina(n270), .dinb(a14 ), .dout(n492));
  jor  g0230(.dina(n492), .dinb(n269), .dout(n493));
  jand g0231(.dina(n493), .dinb(n491), .dout(n494));
  jand g0232(.dina(shift0 ), .dinb(a13 ), .dout(n495));
  jand g0233(.dina(n495), .dinb(shift1 ), .dout(n496));
  jand g0234(.dina(n270), .dinb(a16 ), .dout(n497));
  jand g0235(.dina(n497), .dinb(n269), .dout(n498));
  jor  g0236(.dina(n498), .dinb(n496), .dout(n499));
  jor  g0237(.dina(n499), .dinb(n494), .dout(n500));
  jand g0238(.dina(n500), .dinb(n266), .dout(n501));
  jand g0239(.dina(shift0 ), .dinb(a7 ), .dout(n502));
  jor  g0240(.dina(n502), .dinb(shift1 ), .dout(n503));
  jand g0241(.dina(n270), .dinb(a6 ), .dout(n504));
  jor  g0242(.dina(n504), .dinb(n269), .dout(n505));
  jand g0243(.dina(n505), .dinb(n503), .dout(n506));
  jand g0244(.dina(shift0 ), .dinb(a5 ), .dout(n507));
  jand g0245(.dina(n507), .dinb(shift1 ), .dout(n508));
  jand g0246(.dina(n270), .dinb(a8 ), .dout(n509));
  jand g0247(.dina(n509), .dinb(n269), .dout(n510));
  jor  g0248(.dina(n510), .dinb(n508), .dout(n511));
  jor  g0249(.dina(n511), .dinb(n506), .dout(n512));
  jand g0250(.dina(n512), .dinb(n281), .dout(n513));
  jor  g0251(.dina(n513), .dinb(n501), .dout(n514));
  jand g0252(.dina(shift0 ), .dinb(a11 ), .dout(n515));
  jor  g0253(.dina(n515), .dinb(shift1 ), .dout(n516));
  jand g0254(.dina(n270), .dinb(a10 ), .dout(n517));
  jor  g0255(.dina(n517), .dinb(n269), .dout(n518));
  jand g0256(.dina(n518), .dinb(n516), .dout(n519));
  jand g0257(.dina(shift0 ), .dinb(a9 ), .dout(n520));
  jand g0258(.dina(n520), .dinb(shift1 ), .dout(n521));
  jand g0259(.dina(n270), .dinb(a12 ), .dout(n522));
  jand g0260(.dina(n522), .dinb(n269), .dout(n523));
  jor  g0261(.dina(n523), .dinb(n521), .dout(n524));
  jor  g0262(.dina(n524), .dinb(n519), .dout(n525));
  jand g0263(.dina(n525), .dinb(n295), .dout(n526));
  jand g0264(.dina(shift0 ), .dinb(a3 ), .dout(n527));
  jor  g0265(.dina(n527), .dinb(shift1 ), .dout(n528));
  jand g0266(.dina(n270), .dinb(a2 ), .dout(n529));
  jor  g0267(.dina(n529), .dinb(n269), .dout(n530));
  jand g0268(.dina(n530), .dinb(n528), .dout(n531));
  jand g0269(.dina(shift0 ), .dinb(a1 ), .dout(n532));
  jand g0270(.dina(n532), .dinb(shift1 ), .dout(n533));
  jand g0271(.dina(n270), .dinb(a4 ), .dout(n534));
  jand g0272(.dina(n534), .dinb(n269), .dout(n535));
  jor  g0273(.dina(n535), .dinb(n533), .dout(n536));
  jor  g0274(.dina(n536), .dinb(n531), .dout(n537));
  jand g0275(.dina(n537), .dinb(n308), .dout(n538));
  jor  g0276(.dina(n538), .dinb(n526), .dout(n539));
  jor  g0277(.dina(n539), .dinb(n514), .dout(n540));
  jand g0278(.dina(n540), .dinb(n323), .dout(n541));
  jand g0279(.dina(shift0 ), .dinb(a47 ), .dout(n542));
  jor  g0280(.dina(n542), .dinb(shift1 ), .dout(n543));
  jand g0281(.dina(n270), .dinb(a46 ), .dout(n544));
  jor  g0282(.dina(n544), .dinb(n269), .dout(n545));
  jand g0283(.dina(n545), .dinb(n543), .dout(n546));
  jand g0284(.dina(shift0 ), .dinb(a45 ), .dout(n547));
  jand g0285(.dina(n547), .dinb(shift1 ), .dout(n548));
  jand g0286(.dina(n270), .dinb(a48 ), .dout(n549));
  jand g0287(.dina(n549), .dinb(n269), .dout(n550));
  jor  g0288(.dina(n550), .dinb(n548), .dout(n551));
  jor  g0289(.dina(n551), .dinb(n546), .dout(n552));
  jand g0290(.dina(n552), .dinb(n266), .dout(n553));
  jand g0291(.dina(n270), .dinb(a40 ), .dout(n554));
  jand g0292(.dina(shift0 ), .dinb(a39 ), .dout(n555));
  jor  g0293(.dina(n555), .dinb(n554), .dout(n556));
  jand g0294(.dina(n556), .dinb(n269), .dout(n557));
  jand g0295(.dina(n270), .dinb(a38 ), .dout(n558));
  jand g0296(.dina(shift0 ), .dinb(a37 ), .dout(n559));
  jor  g0297(.dina(n559), .dinb(n558), .dout(n560));
  jand g0298(.dina(n560), .dinb(shift1 ), .dout(n561));
  jor  g0299(.dina(n561), .dinb(n557), .dout(n562));
  jand g0300(.dina(n562), .dinb(n281), .dout(n563));
  jor  g0301(.dina(n563), .dinb(n553), .dout(n564));
  jand g0302(.dina(shift0 ), .dinb(a43 ), .dout(n565));
  jor  g0303(.dina(n565), .dinb(shift1 ), .dout(n566));
  jand g0304(.dina(n270), .dinb(a42 ), .dout(n567));
  jor  g0305(.dina(n567), .dinb(n269), .dout(n568));
  jand g0306(.dina(n568), .dinb(n566), .dout(n569));
  jand g0307(.dina(shift0 ), .dinb(a41 ), .dout(n570));
  jand g0308(.dina(n570), .dinb(shift1 ), .dout(n571));
  jand g0309(.dina(n270), .dinb(a44 ), .dout(n572));
  jand g0310(.dina(n572), .dinb(n269), .dout(n573));
  jor  g0311(.dina(n573), .dinb(n571), .dout(n574));
  jor  g0312(.dina(n574), .dinb(n569), .dout(n575));
  jand g0313(.dina(n575), .dinb(n295), .dout(n576));
  jand g0314(.dina(shift0 ), .dinb(a35 ), .dout(n577));
  jor  g0315(.dina(n577), .dinb(shift1 ), .dout(n578));
  jand g0316(.dina(n270), .dinb(a34 ), .dout(n579));
  jor  g0317(.dina(n579), .dinb(n269), .dout(n580));
  jand g0318(.dina(n580), .dinb(n578), .dout(n581));
  jand g0319(.dina(shift0 ), .dinb(a33 ), .dout(n582));
  jand g0320(.dina(n582), .dinb(shift1 ), .dout(n583));
  jand g0321(.dina(n270), .dinb(a36 ), .dout(n584));
  jand g0322(.dina(n584), .dinb(n269), .dout(n585));
  jor  g0323(.dina(n585), .dinb(n583), .dout(n586));
  jor  g0324(.dina(n586), .dinb(n581), .dout(n587));
  jand g0325(.dina(n587), .dinb(n308), .dout(n588));
  jor  g0326(.dina(n588), .dinb(n576), .dout(n589));
  jor  g0327(.dina(n589), .dinb(n564), .dout(n590));
  jand g0328(.dina(n590), .dinb(n377), .dout(n591));
  jor  g0329(.dina(n591), .dinb(n541), .dout(n592));
  jand g0330(.dina(shift0 ), .dinb(a31 ), .dout(n593));
  jor  g0331(.dina(n593), .dinb(shift1 ), .dout(n594));
  jand g0332(.dina(n270), .dinb(a30 ), .dout(n595));
  jor  g0333(.dina(n595), .dinb(n269), .dout(n596));
  jand g0334(.dina(n596), .dinb(n594), .dout(n597));
  jand g0335(.dina(shift0 ), .dinb(a29 ), .dout(n598));
  jand g0336(.dina(n598), .dinb(shift1 ), .dout(n599));
  jand g0337(.dina(n270), .dinb(a32 ), .dout(n600));
  jand g0338(.dina(n600), .dinb(n269), .dout(n601));
  jor  g0339(.dina(n601), .dinb(n599), .dout(n602));
  jor  g0340(.dina(n602), .dinb(n597), .dout(n603));
  jand g0341(.dina(n603), .dinb(n266), .dout(n604));
  jand g0342(.dina(shift0 ), .dinb(a23 ), .dout(n605));
  jor  g0343(.dina(n605), .dinb(shift1 ), .dout(n606));
  jand g0344(.dina(n270), .dinb(a22 ), .dout(n607));
  jor  g0345(.dina(n607), .dinb(n269), .dout(n608));
  jand g0346(.dina(n608), .dinb(n606), .dout(n609));
  jand g0347(.dina(shift0 ), .dinb(a21 ), .dout(n610));
  jand g0348(.dina(n610), .dinb(shift1 ), .dout(n611));
  jand g0349(.dina(n270), .dinb(a24 ), .dout(n612));
  jand g0350(.dina(n612), .dinb(n269), .dout(n613));
  jor  g0351(.dina(n613), .dinb(n611), .dout(n614));
  jor  g0352(.dina(n614), .dinb(n609), .dout(n615));
  jand g0353(.dina(n615), .dinb(n281), .dout(n616));
  jor  g0354(.dina(n616), .dinb(n604), .dout(n617));
  jand g0355(.dina(shift0 ), .dinb(a27 ), .dout(n618));
  jor  g0356(.dina(n618), .dinb(shift1 ), .dout(n619));
  jand g0357(.dina(n270), .dinb(a26 ), .dout(n620));
  jor  g0358(.dina(n620), .dinb(n269), .dout(n621));
  jand g0359(.dina(n621), .dinb(n619), .dout(n622));
  jand g0360(.dina(shift0 ), .dinb(a25 ), .dout(n623));
  jand g0361(.dina(n623), .dinb(shift1 ), .dout(n624));
  jand g0362(.dina(n270), .dinb(a28 ), .dout(n625));
  jand g0363(.dina(n625), .dinb(n269), .dout(n626));
  jor  g0364(.dina(n626), .dinb(n624), .dout(n627));
  jor  g0365(.dina(n627), .dinb(n622), .dout(n628));
  jand g0366(.dina(n628), .dinb(n295), .dout(n629));
  jand g0367(.dina(shift0 ), .dinb(a19 ), .dout(n630));
  jor  g0368(.dina(n630), .dinb(shift1 ), .dout(n631));
  jand g0369(.dina(n270), .dinb(a18 ), .dout(n632));
  jor  g0370(.dina(n632), .dinb(n269), .dout(n633));
  jand g0371(.dina(n633), .dinb(n631), .dout(n634));
  jand g0372(.dina(shift0 ), .dinb(a17 ), .dout(n635));
  jand g0373(.dina(n635), .dinb(shift1 ), .dout(n636));
  jand g0374(.dina(n270), .dinb(a20 ), .dout(n637));
  jand g0375(.dina(n637), .dinb(n269), .dout(n638));
  jor  g0376(.dina(n638), .dinb(n636), .dout(n639));
  jor  g0377(.dina(n639), .dinb(n634), .dout(n640));
  jand g0378(.dina(n640), .dinb(n308), .dout(n641));
  jor  g0379(.dina(n641), .dinb(n629), .dout(n642));
  jor  g0380(.dina(n642), .dinb(n617), .dout(n643));
  jand g0381(.dina(n643), .dinb(n432), .dout(n644));
  jand g0382(.dina(shift0 ), .dinb(a63 ), .dout(n645));
  jor  g0383(.dina(n645), .dinb(shift1 ), .dout(n646));
  jand g0384(.dina(n270), .dinb(a62 ), .dout(n647));
  jor  g0385(.dina(n647), .dinb(n269), .dout(n648));
  jand g0386(.dina(n648), .dinb(n646), .dout(n649));
  jand g0387(.dina(shift0 ), .dinb(a61 ), .dout(n650));
  jand g0388(.dina(n650), .dinb(shift1 ), .dout(n651));
  jand g0389(.dina(n270), .dinb(a64 ), .dout(n652));
  jand g0390(.dina(n652), .dinb(n269), .dout(n653));
  jor  g0391(.dina(n653), .dinb(n651), .dout(n654));
  jor  g0392(.dina(n654), .dinb(n649), .dout(n655));
  jand g0393(.dina(n655), .dinb(n266), .dout(n656));
  jand g0394(.dina(shift0 ), .dinb(a55 ), .dout(n657));
  jor  g0395(.dina(n657), .dinb(shift1 ), .dout(n658));
  jand g0396(.dina(n270), .dinb(a54 ), .dout(n659));
  jor  g0397(.dina(n659), .dinb(n269), .dout(n660));
  jand g0398(.dina(n660), .dinb(n658), .dout(n661));
  jand g0399(.dina(shift0 ), .dinb(a53 ), .dout(n662));
  jand g0400(.dina(n662), .dinb(shift1 ), .dout(n663));
  jand g0401(.dina(n270), .dinb(a56 ), .dout(n664));
  jand g0402(.dina(n664), .dinb(n269), .dout(n665));
  jor  g0403(.dina(n665), .dinb(n663), .dout(n666));
  jor  g0404(.dina(n666), .dinb(n661), .dout(n667));
  jand g0405(.dina(n667), .dinb(n281), .dout(n668));
  jor  g0406(.dina(n668), .dinb(n656), .dout(n669));
  jand g0407(.dina(shift0 ), .dinb(a59 ), .dout(n670));
  jor  g0408(.dina(n670), .dinb(shift1 ), .dout(n671));
  jand g0409(.dina(n270), .dinb(a58 ), .dout(n672));
  jor  g0410(.dina(n672), .dinb(n269), .dout(n673));
  jand g0411(.dina(n673), .dinb(n671), .dout(n674));
  jand g0412(.dina(shift0 ), .dinb(a57 ), .dout(n675));
  jand g0413(.dina(n675), .dinb(shift1 ), .dout(n676));
  jand g0414(.dina(n270), .dinb(a60 ), .dout(n677));
  jand g0415(.dina(n677), .dinb(n269), .dout(n678));
  jor  g0416(.dina(n678), .dinb(n676), .dout(n679));
  jor  g0417(.dina(n679), .dinb(n674), .dout(n680));
  jand g0418(.dina(n680), .dinb(n295), .dout(n681));
  jand g0419(.dina(shift0 ), .dinb(a51 ), .dout(n682));
  jor  g0420(.dina(n682), .dinb(shift1 ), .dout(n683));
  jand g0421(.dina(n270), .dinb(a50 ), .dout(n684));
  jor  g0422(.dina(n684), .dinb(n269), .dout(n685));
  jand g0423(.dina(n685), .dinb(n683), .dout(n686));
  jand g0424(.dina(shift0 ), .dinb(a49 ), .dout(n687));
  jand g0425(.dina(n687), .dinb(shift1 ), .dout(n688));
  jand g0426(.dina(n270), .dinb(a52 ), .dout(n689));
  jand g0427(.dina(n689), .dinb(n269), .dout(n690));
  jor  g0428(.dina(n690), .dinb(n688), .dout(n691));
  jor  g0429(.dina(n691), .dinb(n686), .dout(n692));
  jand g0430(.dina(n692), .dinb(n308), .dout(n693));
  jor  g0431(.dina(n693), .dinb(n681), .dout(n694));
  jor  g0432(.dina(n694), .dinb(n669), .dout(n695));
  jand g0433(.dina(n695), .dinb(n485), .dout(n696));
  jor  g0434(.dina(n696), .dinb(n644), .dout(n697));
  jor  g0435(.dina(n697), .dinb(n592), .dout(n698));
  jand g0436(.dina(n698), .dinb(shift6 ), .dout(n699));
  jor  g0437(.dina(n699), .dinb(n489), .dout(result0 ));
  jor  g0438(.dina(n270), .dinb(a78 ), .dout(n701));
  jor  g0439(.dina(shift0 ), .dinb(a79 ), .dout(n702));
  jand g0440(.dina(n702), .dinb(n701), .dout(n703));
  jor  g0441(.dina(n703), .dinb(n269), .dout(n704));
  jor  g0442(.dina(n270), .dinb(a80 ), .dout(n705));
  jor  g0443(.dina(shift0 ), .dinb(a81 ), .dout(n706));
  jand g0444(.dina(n706), .dinb(n705), .dout(n707));
  jor  g0445(.dina(n707), .dinb(shift1 ), .dout(n708));
  jand g0446(.dina(n708), .dinb(n704), .dout(n709));
  jand g0447(.dina(n709), .dinb(n266), .dout(n710));
  jor  g0448(.dina(n270), .dinb(a70 ), .dout(n711));
  jor  g0449(.dina(shift0 ), .dinb(a71 ), .dout(n712));
  jand g0450(.dina(n712), .dinb(n711), .dout(n713));
  jor  g0451(.dina(n713), .dinb(n269), .dout(n714));
  jor  g0452(.dina(n270), .dinb(a72 ), .dout(n715));
  jor  g0453(.dina(shift0 ), .dinb(a73 ), .dout(n716));
  jand g0454(.dina(n716), .dinb(n715), .dout(n717));
  jor  g0455(.dina(n717), .dinb(shift1 ), .dout(n718));
  jand g0456(.dina(n718), .dinb(n714), .dout(n719));
  jand g0457(.dina(n719), .dinb(n281), .dout(n720));
  jor  g0458(.dina(n720), .dinb(n710), .dout(n721));
  jor  g0459(.dina(n270), .dinb(a74 ), .dout(n722));
  jor  g0460(.dina(shift0 ), .dinb(a75 ), .dout(n723));
  jand g0461(.dina(n723), .dinb(n722), .dout(n724));
  jor  g0462(.dina(n724), .dinb(n269), .dout(n725));
  jor  g0463(.dina(n270), .dinb(a76 ), .dout(n726));
  jor  g0464(.dina(shift0 ), .dinb(a77 ), .dout(n727));
  jand g0465(.dina(n727), .dinb(n726), .dout(n728));
  jor  g0466(.dina(n728), .dinb(shift1 ), .dout(n729));
  jand g0467(.dina(n729), .dinb(n725), .dout(n730));
  jand g0468(.dina(n730), .dinb(n295), .dout(n731));
  jor  g0469(.dina(n270), .dinb(a66 ), .dout(n732));
  jor  g0470(.dina(shift0 ), .dinb(a67 ), .dout(n733));
  jand g0471(.dina(n733), .dinb(n732), .dout(n734));
  jor  g0472(.dina(n734), .dinb(n269), .dout(n735));
  jor  g0473(.dina(n270), .dinb(a68 ), .dout(n736));
  jor  g0474(.dina(shift0 ), .dinb(a69 ), .dout(n737));
  jand g0475(.dina(n737), .dinb(n736), .dout(n738));
  jor  g0476(.dina(n738), .dinb(shift1 ), .dout(n739));
  jand g0477(.dina(n739), .dinb(n735), .dout(n740));
  jand g0478(.dina(n740), .dinb(n308), .dout(n741));
  jor  g0479(.dina(n741), .dinb(n731), .dout(n742));
  jor  g0480(.dina(n742), .dinb(n721), .dout(n743));
  jand g0481(.dina(n743), .dinb(n323), .dout(n744));
  jor  g0482(.dina(n270), .dinb(a110 ), .dout(n745));
  jor  g0483(.dina(shift0 ), .dinb(a111 ), .dout(n746));
  jand g0484(.dina(n746), .dinb(n745), .dout(n747));
  jor  g0485(.dina(n747), .dinb(n269), .dout(n748));
  jor  g0486(.dina(n270), .dinb(a112 ), .dout(n749));
  jor  g0487(.dina(shift0 ), .dinb(a113 ), .dout(n750));
  jand g0488(.dina(n750), .dinb(n749), .dout(n751));
  jor  g0489(.dina(n751), .dinb(shift1 ), .dout(n752));
  jand g0490(.dina(n752), .dinb(n748), .dout(n753));
  jand g0491(.dina(n753), .dinb(n266), .dout(n754));
  jor  g0492(.dina(n270), .dinb(a102 ), .dout(n755));
  jor  g0493(.dina(shift0 ), .dinb(a103 ), .dout(n756));
  jand g0494(.dina(n756), .dinb(n755), .dout(n757));
  jor  g0495(.dina(n757), .dinb(n269), .dout(n758));
  jor  g0496(.dina(n270), .dinb(a104 ), .dout(n759));
  jor  g0497(.dina(shift0 ), .dinb(a105 ), .dout(n760));
  jand g0498(.dina(n760), .dinb(n759), .dout(n761));
  jor  g0499(.dina(n761), .dinb(shift1 ), .dout(n762));
  jand g0500(.dina(n762), .dinb(n758), .dout(n763));
  jand g0501(.dina(n763), .dinb(n281), .dout(n764));
  jor  g0502(.dina(n764), .dinb(n754), .dout(n765));
  jor  g0503(.dina(n270), .dinb(a106 ), .dout(n766));
  jor  g0504(.dina(shift0 ), .dinb(a107 ), .dout(n767));
  jand g0505(.dina(n767), .dinb(n766), .dout(n768));
  jor  g0506(.dina(n768), .dinb(n269), .dout(n769));
  jor  g0507(.dina(n270), .dinb(a108 ), .dout(n770));
  jor  g0508(.dina(shift0 ), .dinb(a109 ), .dout(n771));
  jand g0509(.dina(n771), .dinb(n770), .dout(n772));
  jor  g0510(.dina(n772), .dinb(shift1 ), .dout(n773));
  jand g0511(.dina(n773), .dinb(n769), .dout(n774));
  jand g0512(.dina(n774), .dinb(n295), .dout(n775));
  jor  g0513(.dina(n270), .dinb(a98 ), .dout(n776));
  jor  g0514(.dina(shift0 ), .dinb(a99 ), .dout(n777));
  jand g0515(.dina(n777), .dinb(n776), .dout(n778));
  jor  g0516(.dina(n778), .dinb(n269), .dout(n779));
  jor  g0517(.dina(n270), .dinb(a100 ), .dout(n780));
  jor  g0518(.dina(shift0 ), .dinb(a101 ), .dout(n781));
  jand g0519(.dina(n781), .dinb(n780), .dout(n782));
  jor  g0520(.dina(n782), .dinb(shift1 ), .dout(n783));
  jand g0521(.dina(n783), .dinb(n779), .dout(n784));
  jand g0522(.dina(n784), .dinb(n308), .dout(n785));
  jor  g0523(.dina(n785), .dinb(n775), .dout(n786));
  jor  g0524(.dina(n786), .dinb(n765), .dout(n787));
  jand g0525(.dina(n787), .dinb(n377), .dout(n788));
  jor  g0526(.dina(n788), .dinb(n744), .dout(n789));
  jor  g0527(.dina(n270), .dinb(a94 ), .dout(n790));
  jor  g0528(.dina(shift0 ), .dinb(a95 ), .dout(n791));
  jand g0529(.dina(n791), .dinb(n790), .dout(n792));
  jor  g0530(.dina(n792), .dinb(n269), .dout(n793));
  jor  g0531(.dina(n270), .dinb(a96 ), .dout(n794));
  jor  g0532(.dina(shift0 ), .dinb(a97 ), .dout(n795));
  jand g0533(.dina(n795), .dinb(n794), .dout(n796));
  jor  g0534(.dina(n796), .dinb(shift1 ), .dout(n797));
  jand g0535(.dina(n797), .dinb(n793), .dout(n798));
  jand g0536(.dina(n798), .dinb(n266), .dout(n799));
  jor  g0537(.dina(n270), .dinb(a86 ), .dout(n800));
  jor  g0538(.dina(shift0 ), .dinb(a87 ), .dout(n801));
  jand g0539(.dina(n801), .dinb(n800), .dout(n802));
  jor  g0540(.dina(n802), .dinb(n269), .dout(n803));
  jor  g0541(.dina(n270), .dinb(a88 ), .dout(n804));
  jor  g0542(.dina(shift0 ), .dinb(a89 ), .dout(n805));
  jand g0543(.dina(n805), .dinb(n804), .dout(n806));
  jor  g0544(.dina(n806), .dinb(shift1 ), .dout(n807));
  jand g0545(.dina(n807), .dinb(n803), .dout(n808));
  jand g0546(.dina(n808), .dinb(n281), .dout(n809));
  jor  g0547(.dina(n809), .dinb(n799), .dout(n810));
  jor  g0548(.dina(n270), .dinb(a90 ), .dout(n811));
  jor  g0549(.dina(shift0 ), .dinb(a91 ), .dout(n812));
  jand g0550(.dina(n812), .dinb(n811), .dout(n813));
  jor  g0551(.dina(n813), .dinb(n269), .dout(n814));
  jor  g0552(.dina(n270), .dinb(a92 ), .dout(n815));
  jor  g0553(.dina(shift0 ), .dinb(a93 ), .dout(n816));
  jand g0554(.dina(n816), .dinb(n815), .dout(n817));
  jor  g0555(.dina(n817), .dinb(shift1 ), .dout(n818));
  jand g0556(.dina(n818), .dinb(n814), .dout(n819));
  jand g0557(.dina(n819), .dinb(n295), .dout(n820));
  jor  g0558(.dina(n270), .dinb(a82 ), .dout(n821));
  jor  g0559(.dina(shift0 ), .dinb(a83 ), .dout(n822));
  jand g0560(.dina(n822), .dinb(n821), .dout(n823));
  jor  g0561(.dina(n823), .dinb(n269), .dout(n824));
  jor  g0562(.dina(n270), .dinb(a84 ), .dout(n825));
  jor  g0563(.dina(shift0 ), .dinb(a85 ), .dout(n826));
  jand g0564(.dina(n826), .dinb(n825), .dout(n827));
  jor  g0565(.dina(n827), .dinb(shift1 ), .dout(n828));
  jand g0566(.dina(n828), .dinb(n824), .dout(n829));
  jand g0567(.dina(n829), .dinb(n308), .dout(n830));
  jor  g0568(.dina(n830), .dinb(n820), .dout(n831));
  jor  g0569(.dina(n831), .dinb(n810), .dout(n832));
  jand g0570(.dina(n832), .dinb(n432), .dout(n833));
  jor  g0571(.dina(n270), .dinb(a126 ), .dout(n834));
  jor  g0572(.dina(shift0 ), .dinb(a127 ), .dout(n835));
  jand g0573(.dina(n835), .dinb(n834), .dout(n836));
  jor  g0574(.dina(n836), .dinb(n269), .dout(n837));
  jor  g0575(.dina(n270), .dinb(a0 ), .dout(n838));
  jor  g0576(.dina(shift0 ), .dinb(a1 ), .dout(n839));
  jand g0577(.dina(n839), .dinb(n838), .dout(n840));
  jor  g0578(.dina(n840), .dinb(shift1 ), .dout(n841));
  jand g0579(.dina(n841), .dinb(n837), .dout(n842));
  jand g0580(.dina(n842), .dinb(n266), .dout(n843));
  jor  g0581(.dina(n270), .dinb(a118 ), .dout(n844));
  jor  g0582(.dina(shift0 ), .dinb(a119 ), .dout(n845));
  jand g0583(.dina(n845), .dinb(n844), .dout(n846));
  jor  g0584(.dina(n846), .dinb(n269), .dout(n847));
  jor  g0585(.dina(n270), .dinb(a120 ), .dout(n848));
  jor  g0586(.dina(shift0 ), .dinb(a121 ), .dout(n849));
  jand g0587(.dina(n849), .dinb(n848), .dout(n850));
  jor  g0588(.dina(n850), .dinb(shift1 ), .dout(n851));
  jand g0589(.dina(n851), .dinb(n847), .dout(n852));
  jand g0590(.dina(n852), .dinb(n281), .dout(n853));
  jor  g0591(.dina(n853), .dinb(n843), .dout(n854));
  jor  g0592(.dina(n270), .dinb(a122 ), .dout(n855));
  jor  g0593(.dina(shift0 ), .dinb(a123 ), .dout(n856));
  jand g0594(.dina(n856), .dinb(n855), .dout(n857));
  jor  g0595(.dina(n857), .dinb(n269), .dout(n858));
  jor  g0596(.dina(n270), .dinb(a124 ), .dout(n859));
  jor  g0597(.dina(shift0 ), .dinb(a125 ), .dout(n860));
  jand g0598(.dina(n860), .dinb(n859), .dout(n861));
  jor  g0599(.dina(n861), .dinb(shift1 ), .dout(n862));
  jand g0600(.dina(n862), .dinb(n858), .dout(n863));
  jand g0601(.dina(n863), .dinb(n295), .dout(n864));
  jor  g0602(.dina(n270), .dinb(a114 ), .dout(n865));
  jor  g0603(.dina(shift0 ), .dinb(a115 ), .dout(n866));
  jand g0604(.dina(n866), .dinb(n865), .dout(n867));
  jor  g0605(.dina(n867), .dinb(n269), .dout(n868));
  jor  g0606(.dina(n270), .dinb(a116 ), .dout(n869));
  jor  g0607(.dina(shift0 ), .dinb(a117 ), .dout(n870));
  jand g0608(.dina(n870), .dinb(n869), .dout(n871));
  jor  g0609(.dina(n871), .dinb(shift1 ), .dout(n872));
  jand g0610(.dina(n872), .dinb(n868), .dout(n873));
  jand g0611(.dina(n873), .dinb(n308), .dout(n874));
  jor  g0612(.dina(n874), .dinb(n864), .dout(n875));
  jor  g0613(.dina(n875), .dinb(n854), .dout(n876));
  jand g0614(.dina(n876), .dinb(n485), .dout(n877));
  jor  g0615(.dina(n877), .dinb(n833), .dout(n878));
  jor  g0616(.dina(n878), .dinb(n789), .dout(n879));
  jand g0617(.dina(n879), .dinb(n263), .dout(n880));
  jor  g0618(.dina(n270), .dinb(a62 ), .dout(n881));
  jor  g0619(.dina(shift0 ), .dinb(a63 ), .dout(n882));
  jand g0620(.dina(n882), .dinb(n881), .dout(n883));
  jor  g0621(.dina(n883), .dinb(n269), .dout(n884));
  jor  g0622(.dina(n270), .dinb(a64 ), .dout(n885));
  jor  g0623(.dina(shift0 ), .dinb(a65 ), .dout(n886));
  jand g0624(.dina(n886), .dinb(n885), .dout(n887));
  jor  g0625(.dina(n887), .dinb(shift1 ), .dout(n888));
  jand g0626(.dina(n888), .dinb(n884), .dout(n889));
  jand g0627(.dina(n889), .dinb(n266), .dout(n890));
  jor  g0628(.dina(n270), .dinb(a54 ), .dout(n891));
  jor  g0629(.dina(shift0 ), .dinb(a55 ), .dout(n892));
  jand g0630(.dina(n892), .dinb(n891), .dout(n893));
  jor  g0631(.dina(n893), .dinb(n269), .dout(n894));
  jor  g0632(.dina(n270), .dinb(a56 ), .dout(n895));
  jor  g0633(.dina(shift0 ), .dinb(a57 ), .dout(n896));
  jand g0634(.dina(n896), .dinb(n895), .dout(n897));
  jor  g0635(.dina(n897), .dinb(shift1 ), .dout(n898));
  jand g0636(.dina(n898), .dinb(n894), .dout(n899));
  jand g0637(.dina(n899), .dinb(n281), .dout(n900));
  jor  g0638(.dina(n900), .dinb(n890), .dout(n901));
  jor  g0639(.dina(n270), .dinb(a58 ), .dout(n902));
  jor  g0640(.dina(shift0 ), .dinb(a59 ), .dout(n903));
  jand g0641(.dina(n903), .dinb(n902), .dout(n904));
  jor  g0642(.dina(n904), .dinb(n269), .dout(n905));
  jor  g0643(.dina(n270), .dinb(a60 ), .dout(n906));
  jor  g0644(.dina(shift0 ), .dinb(a61 ), .dout(n907));
  jand g0645(.dina(n907), .dinb(n906), .dout(n908));
  jor  g0646(.dina(n908), .dinb(shift1 ), .dout(n909));
  jand g0647(.dina(n909), .dinb(n905), .dout(n910));
  jand g0648(.dina(n910), .dinb(n295), .dout(n911));
  jor  g0649(.dina(n270), .dinb(a50 ), .dout(n912));
  jor  g0650(.dina(shift0 ), .dinb(a51 ), .dout(n913));
  jand g0651(.dina(n913), .dinb(n912), .dout(n914));
  jor  g0652(.dina(n914), .dinb(n269), .dout(n915));
  jor  g0653(.dina(n270), .dinb(a52 ), .dout(n916));
  jor  g0654(.dina(shift0 ), .dinb(a53 ), .dout(n917));
  jand g0655(.dina(n917), .dinb(n916), .dout(n918));
  jor  g0656(.dina(n918), .dinb(shift1 ), .dout(n919));
  jand g0657(.dina(n919), .dinb(n915), .dout(n920));
  jand g0658(.dina(n920), .dinb(n308), .dout(n921));
  jor  g0659(.dina(n921), .dinb(n911), .dout(n922));
  jor  g0660(.dina(n922), .dinb(n901), .dout(n923));
  jand g0661(.dina(n923), .dinb(n485), .dout(n924));
  jor  g0662(.dina(n270), .dinb(a30 ), .dout(n925));
  jor  g0663(.dina(shift0 ), .dinb(a31 ), .dout(n926));
  jand g0664(.dina(n926), .dinb(n925), .dout(n927));
  jor  g0665(.dina(n927), .dinb(n269), .dout(n928));
  jor  g0666(.dina(n270), .dinb(a32 ), .dout(n929));
  jor  g0667(.dina(shift0 ), .dinb(a33 ), .dout(n930));
  jand g0668(.dina(n930), .dinb(n929), .dout(n931));
  jor  g0669(.dina(n931), .dinb(shift1 ), .dout(n932));
  jand g0670(.dina(n932), .dinb(n928), .dout(n933));
  jand g0671(.dina(n933), .dinb(n266), .dout(n934));
  jor  g0672(.dina(n270), .dinb(a22 ), .dout(n935));
  jor  g0673(.dina(shift0 ), .dinb(a23 ), .dout(n936));
  jand g0674(.dina(n936), .dinb(n935), .dout(n937));
  jor  g0675(.dina(n937), .dinb(n269), .dout(n938));
  jor  g0676(.dina(n270), .dinb(a24 ), .dout(n939));
  jor  g0677(.dina(shift0 ), .dinb(a25 ), .dout(n940));
  jand g0678(.dina(n940), .dinb(n939), .dout(n941));
  jor  g0679(.dina(n941), .dinb(shift1 ), .dout(n942));
  jand g0680(.dina(n942), .dinb(n938), .dout(n943));
  jand g0681(.dina(n943), .dinb(n281), .dout(n944));
  jor  g0682(.dina(n944), .dinb(n934), .dout(n945));
  jor  g0683(.dina(n270), .dinb(a26 ), .dout(n946));
  jor  g0684(.dina(shift0 ), .dinb(a27 ), .dout(n947));
  jand g0685(.dina(n947), .dinb(n946), .dout(n948));
  jor  g0686(.dina(n948), .dinb(n269), .dout(n949));
  jor  g0687(.dina(n270), .dinb(a28 ), .dout(n950));
  jor  g0688(.dina(shift0 ), .dinb(a29 ), .dout(n951));
  jand g0689(.dina(n951), .dinb(n950), .dout(n952));
  jor  g0690(.dina(n952), .dinb(shift1 ), .dout(n953));
  jand g0691(.dina(n953), .dinb(n949), .dout(n954));
  jand g0692(.dina(n954), .dinb(n295), .dout(n955));
  jor  g0693(.dina(n270), .dinb(a18 ), .dout(n956));
  jor  g0694(.dina(shift0 ), .dinb(a19 ), .dout(n957));
  jand g0695(.dina(n957), .dinb(n956), .dout(n958));
  jor  g0696(.dina(n958), .dinb(n269), .dout(n959));
  jor  g0697(.dina(n270), .dinb(a20 ), .dout(n960));
  jor  g0698(.dina(shift0 ), .dinb(a21 ), .dout(n961));
  jand g0699(.dina(n961), .dinb(n960), .dout(n962));
  jor  g0700(.dina(n962), .dinb(shift1 ), .dout(n963));
  jand g0701(.dina(n963), .dinb(n959), .dout(n964));
  jand g0702(.dina(n964), .dinb(n308), .dout(n965));
  jor  g0703(.dina(n965), .dinb(n955), .dout(n966));
  jor  g0704(.dina(n966), .dinb(n945), .dout(n967));
  jand g0705(.dina(n967), .dinb(n432), .dout(n968));
  jor  g0706(.dina(n968), .dinb(n924), .dout(n969));
  jor  g0707(.dina(n270), .dinb(a14 ), .dout(n970));
  jor  g0708(.dina(shift0 ), .dinb(a15 ), .dout(n971));
  jand g0709(.dina(n971), .dinb(n970), .dout(n972));
  jor  g0710(.dina(n972), .dinb(n269), .dout(n973));
  jor  g0711(.dina(n270), .dinb(a16 ), .dout(n974));
  jor  g0712(.dina(shift0 ), .dinb(a17 ), .dout(n975));
  jand g0713(.dina(n975), .dinb(n974), .dout(n976));
  jor  g0714(.dina(n976), .dinb(shift1 ), .dout(n977));
  jand g0715(.dina(n977), .dinb(n973), .dout(n978));
  jand g0716(.dina(n978), .dinb(n266), .dout(n979));
  jor  g0717(.dina(n270), .dinb(a6 ), .dout(n980));
  jor  g0718(.dina(shift0 ), .dinb(a7 ), .dout(n981));
  jand g0719(.dina(n981), .dinb(n980), .dout(n982));
  jor  g0720(.dina(n982), .dinb(n269), .dout(n983));
  jor  g0721(.dina(n270), .dinb(a8 ), .dout(n984));
  jor  g0722(.dina(shift0 ), .dinb(a9 ), .dout(n985));
  jand g0723(.dina(n985), .dinb(n984), .dout(n986));
  jor  g0724(.dina(n986), .dinb(shift1 ), .dout(n987));
  jand g0725(.dina(n987), .dinb(n983), .dout(n988));
  jand g0726(.dina(n988), .dinb(n281), .dout(n989));
  jor  g0727(.dina(n989), .dinb(n979), .dout(n990));
  jor  g0728(.dina(n270), .dinb(a10 ), .dout(n991));
  jor  g0729(.dina(shift0 ), .dinb(a11 ), .dout(n992));
  jand g0730(.dina(n992), .dinb(n991), .dout(n993));
  jor  g0731(.dina(n993), .dinb(n269), .dout(n994));
  jor  g0732(.dina(n270), .dinb(a12 ), .dout(n995));
  jor  g0733(.dina(shift0 ), .dinb(a13 ), .dout(n996));
  jand g0734(.dina(n996), .dinb(n995), .dout(n997));
  jor  g0735(.dina(n997), .dinb(shift1 ), .dout(n998));
  jand g0736(.dina(n998), .dinb(n994), .dout(n999));
  jand g0737(.dina(n999), .dinb(n295), .dout(n1000));
  jor  g0738(.dina(n270), .dinb(a2 ), .dout(n1001));
  jor  g0739(.dina(shift0 ), .dinb(a3 ), .dout(n1002));
  jand g0740(.dina(n1002), .dinb(n1001), .dout(n1003));
  jor  g0741(.dina(n1003), .dinb(n269), .dout(n1004));
  jor  g0742(.dina(n270), .dinb(a4 ), .dout(n1005));
  jor  g0743(.dina(shift0 ), .dinb(a5 ), .dout(n1006));
  jand g0744(.dina(n1006), .dinb(n1005), .dout(n1007));
  jor  g0745(.dina(n1007), .dinb(shift1 ), .dout(n1008));
  jand g0746(.dina(n1008), .dinb(n1004), .dout(n1009));
  jand g0747(.dina(n1009), .dinb(n308), .dout(n1010));
  jor  g0748(.dina(n1010), .dinb(n1000), .dout(n1011));
  jor  g0749(.dina(n1011), .dinb(n990), .dout(n1012));
  jand g0750(.dina(n1012), .dinb(n323), .dout(n1013));
  jor  g0751(.dina(n270), .dinb(a48 ), .dout(n1014));
  jor  g0752(.dina(shift0 ), .dinb(a49 ), .dout(n1015));
  jand g0753(.dina(n1015), .dinb(n1014), .dout(n1016));
  jand g0754(.dina(n1016), .dinb(n269), .dout(n1017));
  jand g0755(.dina(n270), .dinb(a47 ), .dout(n1018));
  jand g0756(.dina(shift0 ), .dinb(a46 ), .dout(n1019));
  jor  g0757(.dina(n1019), .dinb(n1018), .dout(n1020));
  jand g0758(.dina(n1020), .dinb(shift1 ), .dout(n1021));
  jor  g0759(.dina(n1021), .dinb(n1017), .dout(n1022));
  jand g0760(.dina(n1022), .dinb(n266), .dout(n1023));
  jand g0761(.dina(n270), .dinb(a39 ), .dout(n1024));
  jor  g0762(.dina(n1024), .dinb(n269), .dout(n1025));
  jand g0763(.dina(n270), .dinb(a41 ), .dout(n1026));
  jor  g0764(.dina(n1026), .dinb(shift1 ), .dout(n1027));
  jand g0765(.dina(n1027), .dinb(n1025), .dout(n1028));
  jand g0766(.dina(shift0 ), .dinb(a38 ), .dout(n1029));
  jand g0767(.dina(n1029), .dinb(shift1 ), .dout(n1030));
  jand g0768(.dina(shift0 ), .dinb(a40 ), .dout(n1031));
  jand g0769(.dina(n1031), .dinb(n269), .dout(n1032));
  jor  g0770(.dina(n1032), .dinb(n1030), .dout(n1033));
  jor  g0771(.dina(n1033), .dinb(n1028), .dout(n1034));
  jand g0772(.dina(n1034), .dinb(n281), .dout(n1035));
  jor  g0773(.dina(n1035), .dinb(n1023), .dout(n1036));
  jand g0774(.dina(shift0 ), .dinb(a44 ), .dout(n1037));
  jor  g0775(.dina(n1037), .dinb(shift1 ), .dout(n1038));
  jand g0776(.dina(n270), .dinb(a43 ), .dout(n1039));
  jor  g0777(.dina(n1039), .dinb(n269), .dout(n1040));
  jand g0778(.dina(n1040), .dinb(n1038), .dout(n1041));
  jand g0779(.dina(shift0 ), .dinb(a42 ), .dout(n1042));
  jand g0780(.dina(n1042), .dinb(shift1 ), .dout(n1043));
  jand g0781(.dina(n270), .dinb(a45 ), .dout(n1044));
  jand g0782(.dina(n1044), .dinb(n269), .dout(n1045));
  jor  g0783(.dina(n1045), .dinb(n1043), .dout(n1046));
  jor  g0784(.dina(n1046), .dinb(n1041), .dout(n1047));
  jand g0785(.dina(n1047), .dinb(n295), .dout(n1048));
  jor  g0786(.dina(n270), .dinb(a34 ), .dout(n1049));
  jor  g0787(.dina(shift0 ), .dinb(a35 ), .dout(n1050));
  jand g0788(.dina(n1050), .dinb(n1049), .dout(n1051));
  jor  g0789(.dina(n1051), .dinb(n269), .dout(n1052));
  jor  g0790(.dina(n270), .dinb(a36 ), .dout(n1053));
  jor  g0791(.dina(shift0 ), .dinb(a37 ), .dout(n1054));
  jand g0792(.dina(n1054), .dinb(n1053), .dout(n1055));
  jor  g0793(.dina(n1055), .dinb(shift1 ), .dout(n1056));
  jand g0794(.dina(n1056), .dinb(n1052), .dout(n1057));
  jand g0795(.dina(n1057), .dinb(n308), .dout(n1058));
  jor  g0796(.dina(n1058), .dinb(n1048), .dout(n1059));
  jor  g0797(.dina(n1059), .dinb(n1036), .dout(n1060));
  jand g0798(.dina(n1060), .dinb(n377), .dout(n1061));
  jor  g0799(.dina(n1061), .dinb(n1013), .dout(n1062));
  jor  g0800(.dina(n1062), .dinb(n969), .dout(n1063));
  jand g0801(.dina(n1063), .dinb(shift6 ), .dout(n1064));
  jor  g0802(.dina(n1064), .dinb(n880), .dout(result1 ));
  jor  g0803(.dina(n419), .dinb(shift1 ), .dout(n1066));
  jor  g0804(.dina(n267), .dinb(n269), .dout(n1067));
  jand g0805(.dina(n1067), .dinb(n1066), .dout(n1068));
  jand g0806(.dina(n276), .dinb(shift1 ), .dout(n1069));
  jand g0807(.dina(n422), .dinb(n269), .dout(n1070));
  jor  g0808(.dina(n1070), .dinb(n1069), .dout(n1071));
  jor  g0809(.dina(n1071), .dinb(n1068), .dout(n1072));
  jand g0810(.dina(n1072), .dinb(n266), .dout(n1073));
  jor  g0811(.dina(n298), .dinb(shift1 ), .dout(n1074));
  jor  g0812(.dina(n282), .dinb(n269), .dout(n1075));
  jand g0813(.dina(n1075), .dinb(n1074), .dout(n1076));
  jand g0814(.dina(n289), .dinb(shift1 ), .dout(n1077));
  jand g0815(.dina(n301), .dinb(n269), .dout(n1078));
  jor  g0816(.dina(n1078), .dinb(n1077), .dout(n1079));
  jor  g0817(.dina(n1079), .dinb(n1076), .dout(n1080));
  jand g0818(.dina(n1080), .dinb(n281), .dout(n1081));
  jor  g0819(.dina(n1081), .dinb(n1073), .dout(n1082));
  jor  g0820(.dina(n271), .dinb(shift1 ), .dout(n1083));
  jor  g0821(.dina(n296), .dinb(n269), .dout(n1084));
  jand g0822(.dina(n1084), .dinb(n1083), .dout(n1085));
  jand g0823(.dina(n303), .dinb(shift1 ), .dout(n1086));
  jand g0824(.dina(n274), .dinb(n269), .dout(n1087));
  jor  g0825(.dina(n1087), .dinb(n1086), .dout(n1088));
  jor  g0826(.dina(n1088), .dinb(n1085), .dout(n1089));
  jand g0827(.dina(n1089), .dinb(n295), .dout(n1090));
  jor  g0828(.dina(n284), .dinb(shift1 ), .dout(n1091));
  jor  g0829(.dina(n309), .dinb(n269), .dout(n1092));
  jand g0830(.dina(n1092), .dinb(n1091), .dout(n1093));
  jand g0831(.dina(n316), .dinb(shift1 ), .dout(n1094));
  jand g0832(.dina(n287), .dinb(n269), .dout(n1095));
  jor  g0833(.dina(n1095), .dinb(n1094), .dout(n1096));
  jor  g0834(.dina(n1096), .dinb(n1093), .dout(n1097));
  jand g0835(.dina(n1097), .dinb(n308), .dout(n1098));
  jor  g0836(.dina(n1098), .dinb(n1090), .dout(n1099));
  jor  g0837(.dina(n1099), .dinb(n1082), .dout(n1100));
  jand g0838(.dina(n1100), .dinb(n323), .dout(n1101));
  jor  g0839(.dina(n473), .dinb(shift1 ), .dout(n1102));
  jor  g0840(.dina(n325), .dinb(n269), .dout(n1103));
  jand g0841(.dina(n1103), .dinb(n1102), .dout(n1104));
  jand g0842(.dina(n332), .dinb(shift1 ), .dout(n1105));
  jand g0843(.dina(n476), .dinb(n269), .dout(n1106));
  jor  g0844(.dina(n1106), .dinb(n1105), .dout(n1107));
  jor  g0845(.dina(n1107), .dinb(n1104), .dout(n1108));
  jand g0846(.dina(n1108), .dinb(n266), .dout(n1109));
  jor  g0847(.dina(n352), .dinb(shift1 ), .dout(n1110));
  jor  g0848(.dina(n337), .dinb(n269), .dout(n1111));
  jand g0849(.dina(n1111), .dinb(n1110), .dout(n1112));
  jand g0850(.dina(n344), .dinb(shift1 ), .dout(n1113));
  jand g0851(.dina(n355), .dinb(n269), .dout(n1114));
  jor  g0852(.dina(n1114), .dinb(n1113), .dout(n1115));
  jor  g0853(.dina(n1115), .dinb(n1112), .dout(n1116));
  jand g0854(.dina(n1116), .dinb(n281), .dout(n1117));
  jor  g0855(.dina(n1117), .dinb(n1109), .dout(n1118));
  jor  g0856(.dina(n327), .dinb(shift1 ), .dout(n1119));
  jor  g0857(.dina(n350), .dinb(n269), .dout(n1120));
  jand g0858(.dina(n1120), .dinb(n1119), .dout(n1121));
  jand g0859(.dina(n357), .dinb(shift1 ), .dout(n1122));
  jand g0860(.dina(n330), .dinb(n269), .dout(n1123));
  jor  g0861(.dina(n1123), .dinb(n1122), .dout(n1124));
  jor  g0862(.dina(n1124), .dinb(n1121), .dout(n1125));
  jand g0863(.dina(n1125), .dinb(n295), .dout(n1126));
  jor  g0864(.dina(n339), .dinb(shift1 ), .dout(n1127));
  jor  g0865(.dina(n362), .dinb(n269), .dout(n1128));
  jand g0866(.dina(n1128), .dinb(n1127), .dout(n1129));
  jand g0867(.dina(n369), .dinb(shift1 ), .dout(n1130));
  jand g0868(.dina(n342), .dinb(n269), .dout(n1131));
  jor  g0869(.dina(n1131), .dinb(n1130), .dout(n1132));
  jor  g0870(.dina(n1132), .dinb(n1129), .dout(n1133));
  jand g0871(.dina(n1133), .dinb(n308), .dout(n1134));
  jor  g0872(.dina(n1134), .dinb(n1126), .dout(n1135));
  jor  g0873(.dina(n1135), .dinb(n1118), .dout(n1136));
  jand g0874(.dina(n1136), .dinb(n377), .dout(n1137));
  jor  g0875(.dina(n1137), .dinb(n1101), .dout(n1138));
  jor  g0876(.dina(n364), .dinb(shift1 ), .dout(n1139));
  jor  g0877(.dina(n380), .dinb(n269), .dout(n1140));
  jand g0878(.dina(n1140), .dinb(n1139), .dout(n1141));
  jand g0879(.dina(n387), .dinb(shift1 ), .dout(n1142));
  jand g0880(.dina(n367), .dinb(n269), .dout(n1143));
  jor  g0881(.dina(n1143), .dinb(n1142), .dout(n1144));
  jor  g0882(.dina(n1144), .dinb(n1141), .dout(n1145));
  jand g0883(.dina(n1145), .dinb(n266), .dout(n1146));
  jor  g0884(.dina(n407), .dinb(shift1 ), .dout(n1147));
  jor  g0885(.dina(n392), .dinb(n269), .dout(n1148));
  jand g0886(.dina(n1148), .dinb(n1147), .dout(n1149));
  jand g0887(.dina(n399), .dinb(shift1 ), .dout(n1150));
  jand g0888(.dina(n410), .dinb(n269), .dout(n1151));
  jor  g0889(.dina(n1151), .dinb(n1150), .dout(n1152));
  jor  g0890(.dina(n1152), .dinb(n1149), .dout(n1153));
  jand g0891(.dina(n1153), .dinb(n281), .dout(n1154));
  jor  g0892(.dina(n1154), .dinb(n1146), .dout(n1155));
  jor  g0893(.dina(n382), .dinb(shift1 ), .dout(n1156));
  jor  g0894(.dina(n405), .dinb(n269), .dout(n1157));
  jand g0895(.dina(n1157), .dinb(n1156), .dout(n1158));
  jand g0896(.dina(n412), .dinb(shift1 ), .dout(n1159));
  jand g0897(.dina(n385), .dinb(n269), .dout(n1160));
  jor  g0898(.dina(n1160), .dinb(n1159), .dout(n1161));
  jor  g0899(.dina(n1161), .dinb(n1158), .dout(n1162));
  jand g0900(.dina(n1162), .dinb(n295), .dout(n1163));
  jor  g0901(.dina(n394), .dinb(shift1 ), .dout(n1164));
  jor  g0902(.dina(n417), .dinb(n269), .dout(n1165));
  jand g0903(.dina(n1165), .dinb(n1164), .dout(n1166));
  jand g0904(.dina(n424), .dinb(shift1 ), .dout(n1167));
  jand g0905(.dina(n397), .dinb(n269), .dout(n1168));
  jor  g0906(.dina(n1168), .dinb(n1167), .dout(n1169));
  jor  g0907(.dina(n1169), .dinb(n1166), .dout(n1170));
  jand g0908(.dina(n1170), .dinb(n308), .dout(n1171));
  jor  g0909(.dina(n1171), .dinb(n1163), .dout(n1172));
  jor  g0910(.dina(n1172), .dinb(n1155), .dout(n1173));
  jand g0911(.dina(n1173), .dinb(n432), .dout(n1174));
  jor  g0912(.dina(n529), .dinb(shift1 ), .dout(n1175));
  jor  g0913(.dina(n434), .dinb(n269), .dout(n1176));
  jand g0914(.dina(n1176), .dinb(n1175), .dout(n1177));
  jand g0915(.dina(n441), .dinb(shift1 ), .dout(n1178));
  jand g0916(.dina(n532), .dinb(n269), .dout(n1179));
  jor  g0917(.dina(n1179), .dinb(n1178), .dout(n1180));
  jor  g0918(.dina(n1180), .dinb(n1177), .dout(n1181));
  jand g0919(.dina(n1181), .dinb(n266), .dout(n1182));
  jor  g0920(.dina(n461), .dinb(shift1 ), .dout(n1183));
  jor  g0921(.dina(n446), .dinb(n269), .dout(n1184));
  jand g0922(.dina(n1184), .dinb(n1183), .dout(n1185));
  jand g0923(.dina(n453), .dinb(shift1 ), .dout(n1186));
  jand g0924(.dina(n464), .dinb(n269), .dout(n1187));
  jor  g0925(.dina(n1187), .dinb(n1186), .dout(n1188));
  jor  g0926(.dina(n1188), .dinb(n1185), .dout(n1189));
  jand g0927(.dina(n1189), .dinb(n281), .dout(n1190));
  jor  g0928(.dina(n1190), .dinb(n1182), .dout(n1191));
  jor  g0929(.dina(n436), .dinb(shift1 ), .dout(n1192));
  jor  g0930(.dina(n459), .dinb(n269), .dout(n1193));
  jand g0931(.dina(n1193), .dinb(n1192), .dout(n1194));
  jand g0932(.dina(n466), .dinb(shift1 ), .dout(n1195));
  jand g0933(.dina(n439), .dinb(n269), .dout(n1196));
  jor  g0934(.dina(n1196), .dinb(n1195), .dout(n1197));
  jor  g0935(.dina(n1197), .dinb(n1194), .dout(n1198));
  jand g0936(.dina(n1198), .dinb(n295), .dout(n1199));
  jor  g0937(.dina(n448), .dinb(shift1 ), .dout(n1200));
  jor  g0938(.dina(n471), .dinb(n269), .dout(n1201));
  jand g0939(.dina(n1201), .dinb(n1200), .dout(n1202));
  jand g0940(.dina(n478), .dinb(shift1 ), .dout(n1203));
  jand g0941(.dina(n451), .dinb(n269), .dout(n1204));
  jor  g0942(.dina(n1204), .dinb(n1203), .dout(n1205));
  jor  g0943(.dina(n1205), .dinb(n1202), .dout(n1206));
  jand g0944(.dina(n1206), .dinb(n308), .dout(n1207));
  jor  g0945(.dina(n1207), .dinb(n1199), .dout(n1208));
  jor  g0946(.dina(n1208), .dinb(n1191), .dout(n1209));
  jand g0947(.dina(n1209), .dinb(n485), .dout(n1210));
  jor  g0948(.dina(n1210), .dinb(n1174), .dout(n1211));
  jor  g0949(.dina(n1211), .dinb(n1138), .dout(n1212));
  jand g0950(.dina(n1212), .dinb(n263), .dout(n1213));
  jor  g0951(.dina(n311), .dinb(shift1 ), .dout(n1214));
  jor  g0952(.dina(n645), .dinb(n269), .dout(n1215));
  jand g0953(.dina(n1215), .dinb(n1214), .dout(n1216));
  jand g0954(.dina(n652), .dinb(shift1 ), .dout(n1217));
  jand g0955(.dina(n314), .dinb(n269), .dout(n1218));
  jor  g0956(.dina(n1218), .dinb(n1217), .dout(n1219));
  jor  g0957(.dina(n1219), .dinb(n1216), .dout(n1220));
  jand g0958(.dina(n1220), .dinb(n266), .dout(n1221));
  jor  g0959(.dina(n672), .dinb(shift1 ), .dout(n1222));
  jor  g0960(.dina(n657), .dinb(n269), .dout(n1223));
  jand g0961(.dina(n1223), .dinb(n1222), .dout(n1224));
  jand g0962(.dina(n664), .dinb(shift1 ), .dout(n1225));
  jand g0963(.dina(n675), .dinb(n269), .dout(n1226));
  jor  g0964(.dina(n1226), .dinb(n1225), .dout(n1227));
  jor  g0965(.dina(n1227), .dinb(n1224), .dout(n1228));
  jand g0966(.dina(n1228), .dinb(n281), .dout(n1229));
  jor  g0967(.dina(n1229), .dinb(n1221), .dout(n1230));
  jor  g0968(.dina(n647), .dinb(shift1 ), .dout(n1231));
  jor  g0969(.dina(n670), .dinb(n269), .dout(n1232));
  jand g0970(.dina(n1232), .dinb(n1231), .dout(n1233));
  jand g0971(.dina(n677), .dinb(shift1 ), .dout(n1234));
  jand g0972(.dina(n650), .dinb(n269), .dout(n1235));
  jor  g0973(.dina(n1235), .dinb(n1234), .dout(n1236));
  jor  g0974(.dina(n1236), .dinb(n1233), .dout(n1237));
  jand g0975(.dina(n1237), .dinb(n295), .dout(n1238));
  jor  g0976(.dina(n659), .dinb(shift1 ), .dout(n1239));
  jor  g0977(.dina(n682), .dinb(n269), .dout(n1240));
  jand g0978(.dina(n1240), .dinb(n1239), .dout(n1241));
  jand g0979(.dina(n689), .dinb(shift1 ), .dout(n1242));
  jand g0980(.dina(n662), .dinb(n269), .dout(n1243));
  jor  g0981(.dina(n1243), .dinb(n1242), .dout(n1244));
  jor  g0982(.dina(n1244), .dinb(n1241), .dout(n1245));
  jand g0983(.dina(n1245), .dinb(n308), .dout(n1246));
  jor  g0984(.dina(n1246), .dinb(n1238), .dout(n1247));
  jor  g0985(.dina(n1247), .dinb(n1230), .dout(n1248));
  jand g0986(.dina(n1248), .dinb(n485), .dout(n1249));
  jor  g0987(.dina(n579), .dinb(shift1 ), .dout(n1250));
  jor  g0988(.dina(n593), .dinb(n269), .dout(n1251));
  jand g0989(.dina(n1251), .dinb(n1250), .dout(n1252));
  jand g0990(.dina(n600), .dinb(shift1 ), .dout(n1253));
  jand g0991(.dina(n582), .dinb(n269), .dout(n1254));
  jor  g0992(.dina(n1254), .dinb(n1253), .dout(n1255));
  jor  g0993(.dina(n1255), .dinb(n1252), .dout(n1256));
  jand g0994(.dina(n1256), .dinb(n266), .dout(n1257));
  jor  g0995(.dina(n620), .dinb(shift1 ), .dout(n1258));
  jor  g0996(.dina(n605), .dinb(n269), .dout(n1259));
  jand g0997(.dina(n1259), .dinb(n1258), .dout(n1260));
  jand g0998(.dina(n612), .dinb(shift1 ), .dout(n1261));
  jand g0999(.dina(n623), .dinb(n269), .dout(n1262));
  jor  g1000(.dina(n1262), .dinb(n1261), .dout(n1263));
  jor  g1001(.dina(n1263), .dinb(n1260), .dout(n1264));
  jand g1002(.dina(n1264), .dinb(n281), .dout(n1265));
  jor  g1003(.dina(n1265), .dinb(n1257), .dout(n1266));
  jor  g1004(.dina(n595), .dinb(shift1 ), .dout(n1267));
  jor  g1005(.dina(n618), .dinb(n269), .dout(n1268));
  jand g1006(.dina(n1268), .dinb(n1267), .dout(n1269));
  jand g1007(.dina(n625), .dinb(shift1 ), .dout(n1270));
  jand g1008(.dina(n598), .dinb(n269), .dout(n1271));
  jor  g1009(.dina(n1271), .dinb(n1270), .dout(n1272));
  jor  g1010(.dina(n1272), .dinb(n1269), .dout(n1273));
  jand g1011(.dina(n1273), .dinb(n295), .dout(n1274));
  jor  g1012(.dina(n607), .dinb(shift1 ), .dout(n1275));
  jor  g1013(.dina(n630), .dinb(n269), .dout(n1276));
  jand g1014(.dina(n1276), .dinb(n1275), .dout(n1277));
  jand g1015(.dina(n637), .dinb(shift1 ), .dout(n1278));
  jand g1016(.dina(n610), .dinb(n269), .dout(n1279));
  jor  g1017(.dina(n1279), .dinb(n1278), .dout(n1280));
  jor  g1018(.dina(n1280), .dinb(n1277), .dout(n1281));
  jand g1019(.dina(n1281), .dinb(n308), .dout(n1282));
  jor  g1020(.dina(n1282), .dinb(n1274), .dout(n1283));
  jor  g1021(.dina(n1283), .dinb(n1266), .dout(n1284));
  jand g1022(.dina(n1284), .dinb(n432), .dout(n1285));
  jor  g1023(.dina(n1285), .dinb(n1249), .dout(n1286));
  jor  g1024(.dina(n632), .dinb(shift1 ), .dout(n1287));
  jor  g1025(.dina(n490), .dinb(n269), .dout(n1288));
  jand g1026(.dina(n1288), .dinb(n1287), .dout(n1289));
  jand g1027(.dina(n497), .dinb(shift1 ), .dout(n1290));
  jand g1028(.dina(n635), .dinb(n269), .dout(n1291));
  jor  g1029(.dina(n1291), .dinb(n1290), .dout(n1292));
  jor  g1030(.dina(n1292), .dinb(n1289), .dout(n1293));
  jand g1031(.dina(n1293), .dinb(n266), .dout(n1294));
  jor  g1032(.dina(n517), .dinb(shift1 ), .dout(n1295));
  jor  g1033(.dina(n502), .dinb(n269), .dout(n1296));
  jand g1034(.dina(n1296), .dinb(n1295), .dout(n1297));
  jand g1035(.dina(n509), .dinb(shift1 ), .dout(n1298));
  jand g1036(.dina(n520), .dinb(n269), .dout(n1299));
  jor  g1037(.dina(n1299), .dinb(n1298), .dout(n1300));
  jor  g1038(.dina(n1300), .dinb(n1297), .dout(n1301));
  jand g1039(.dina(n1301), .dinb(n281), .dout(n1302));
  jor  g1040(.dina(n1302), .dinb(n1294), .dout(n1303));
  jor  g1041(.dina(n492), .dinb(shift1 ), .dout(n1304));
  jor  g1042(.dina(n515), .dinb(n269), .dout(n1305));
  jand g1043(.dina(n1305), .dinb(n1304), .dout(n1306));
  jand g1044(.dina(n522), .dinb(shift1 ), .dout(n1307));
  jand g1045(.dina(n495), .dinb(n269), .dout(n1308));
  jor  g1046(.dina(n1308), .dinb(n1307), .dout(n1309));
  jor  g1047(.dina(n1309), .dinb(n1306), .dout(n1310));
  jand g1048(.dina(n1310), .dinb(n295), .dout(n1311));
  jor  g1049(.dina(n504), .dinb(shift1 ), .dout(n1312));
  jor  g1050(.dina(n527), .dinb(n269), .dout(n1313));
  jand g1051(.dina(n1313), .dinb(n1312), .dout(n1314));
  jand g1052(.dina(n534), .dinb(shift1 ), .dout(n1315));
  jand g1053(.dina(n507), .dinb(n269), .dout(n1316));
  jor  g1054(.dina(n1316), .dinb(n1315), .dout(n1317));
  jor  g1055(.dina(n1317), .dinb(n1314), .dout(n1318));
  jand g1056(.dina(n1318), .dinb(n308), .dout(n1319));
  jor  g1057(.dina(n1319), .dinb(n1311), .dout(n1320));
  jor  g1058(.dina(n1320), .dinb(n1303), .dout(n1321));
  jand g1059(.dina(n1321), .dinb(n323), .dout(n1322));
  jor  g1060(.dina(n684), .dinb(shift1 ), .dout(n1323));
  jor  g1061(.dina(n542), .dinb(n269), .dout(n1324));
  jand g1062(.dina(n1324), .dinb(n1323), .dout(n1325));
  jand g1063(.dina(n549), .dinb(shift1 ), .dout(n1326));
  jand g1064(.dina(n687), .dinb(n269), .dout(n1327));
  jor  g1065(.dina(n1327), .dinb(n1326), .dout(n1328));
  jor  g1066(.dina(n1328), .dinb(n1325), .dout(n1329));
  jand g1067(.dina(n1329), .dinb(n266), .dout(n1330));
  jor  g1068(.dina(n555), .dinb(n269), .dout(n1331));
  jor  g1069(.dina(n570), .dinb(shift1 ), .dout(n1332));
  jand g1070(.dina(n1332), .dinb(n1331), .dout(n1333));
  jand g1071(.dina(n554), .dinb(shift1 ), .dout(n1334));
  jand g1072(.dina(n567), .dinb(n269), .dout(n1335));
  jor  g1073(.dina(n1335), .dinb(n1334), .dout(n1336));
  jor  g1074(.dina(n1336), .dinb(n1333), .dout(n1337));
  jand g1075(.dina(n1337), .dinb(n281), .dout(n1338));
  jor  g1076(.dina(n1338), .dinb(n1330), .dout(n1339));
  jor  g1077(.dina(n547), .dinb(shift1 ), .dout(n1340));
  jor  g1078(.dina(n572), .dinb(n269), .dout(n1341));
  jand g1079(.dina(n1341), .dinb(n1340), .dout(n1342));
  jand g1080(.dina(n565), .dinb(shift1 ), .dout(n1343));
  jand g1081(.dina(n544), .dinb(n269), .dout(n1344));
  jor  g1082(.dina(n1344), .dinb(n1343), .dout(n1345));
  jor  g1083(.dina(n1345), .dinb(n1342), .dout(n1346));
  jand g1084(.dina(n1346), .dinb(n295), .dout(n1347));
  jor  g1085(.dina(n558), .dinb(shift1 ), .dout(n1348));
  jor  g1086(.dina(n577), .dinb(n269), .dout(n1349));
  jand g1087(.dina(n1349), .dinb(n1348), .dout(n1350));
  jand g1088(.dina(n584), .dinb(shift1 ), .dout(n1351));
  jand g1089(.dina(n559), .dinb(n269), .dout(n1352));
  jor  g1090(.dina(n1352), .dinb(n1351), .dout(n1353));
  jor  g1091(.dina(n1353), .dinb(n1350), .dout(n1354));
  jand g1092(.dina(n1354), .dinb(n308), .dout(n1355));
  jor  g1093(.dina(n1355), .dinb(n1347), .dout(n1356));
  jor  g1094(.dina(n1356), .dinb(n1339), .dout(n1357));
  jand g1095(.dina(n1357), .dinb(n377), .dout(n1358));
  jor  g1096(.dina(n1358), .dinb(n1322), .dout(n1359));
  jor  g1097(.dina(n1359), .dinb(n1286), .dout(n1360));
  jand g1098(.dina(n1360), .dinb(shift6 ), .dout(n1361));
  jor  g1099(.dina(n1361), .dinb(n1213), .dout(result2 ));
  jor  g1100(.dina(n751), .dinb(n269), .dout(n1363));
  jor  g1101(.dina(n867), .dinb(shift1 ), .dout(n1364));
  jand g1102(.dina(n1364), .dinb(n1363), .dout(n1365));
  jand g1103(.dina(n1365), .dinb(n266), .dout(n1366));
  jor  g1104(.dina(n761), .dinb(n269), .dout(n1367));
  jor  g1105(.dina(n768), .dinb(shift1 ), .dout(n1368));
  jand g1106(.dina(n1368), .dinb(n1367), .dout(n1369));
  jand g1107(.dina(n1369), .dinb(n281), .dout(n1370));
  jor  g1108(.dina(n1370), .dinb(n1366), .dout(n1371));
  jor  g1109(.dina(n772), .dinb(n269), .dout(n1372));
  jor  g1110(.dina(n747), .dinb(shift1 ), .dout(n1373));
  jand g1111(.dina(n1373), .dinb(n1372), .dout(n1374));
  jand g1112(.dina(n1374), .dinb(n295), .dout(n1375));
  jor  g1113(.dina(n782), .dinb(n269), .dout(n1376));
  jor  g1114(.dina(n757), .dinb(shift1 ), .dout(n1377));
  jand g1115(.dina(n1377), .dinb(n1376), .dout(n1378));
  jand g1116(.dina(n1378), .dinb(n308), .dout(n1379));
  jor  g1117(.dina(n1379), .dinb(n1375), .dout(n1380));
  jor  g1118(.dina(n1380), .dinb(n1371), .dout(n1381));
  jand g1119(.dina(n1381), .dinb(n377), .dout(n1382));
  jor  g1120(.dina(n707), .dinb(n269), .dout(n1383));
  jor  g1121(.dina(n823), .dinb(shift1 ), .dout(n1384));
  jand g1122(.dina(n1384), .dinb(n1383), .dout(n1385));
  jand g1123(.dina(n1385), .dinb(n266), .dout(n1386));
  jor  g1124(.dina(n717), .dinb(n269), .dout(n1387));
  jor  g1125(.dina(n724), .dinb(shift1 ), .dout(n1388));
  jand g1126(.dina(n1388), .dinb(n1387), .dout(n1389));
  jand g1127(.dina(n1389), .dinb(n281), .dout(n1390));
  jor  g1128(.dina(n1390), .dinb(n1386), .dout(n1391));
  jor  g1129(.dina(n728), .dinb(n269), .dout(n1392));
  jor  g1130(.dina(n703), .dinb(shift1 ), .dout(n1393));
  jand g1131(.dina(n1393), .dinb(n1392), .dout(n1394));
  jand g1132(.dina(n1394), .dinb(n295), .dout(n1395));
  jor  g1133(.dina(n738), .dinb(n269), .dout(n1396));
  jor  g1134(.dina(n713), .dinb(shift1 ), .dout(n1397));
  jand g1135(.dina(n1397), .dinb(n1396), .dout(n1398));
  jand g1136(.dina(n1398), .dinb(n308), .dout(n1399));
  jor  g1137(.dina(n1399), .dinb(n1395), .dout(n1400));
  jor  g1138(.dina(n1400), .dinb(n1391), .dout(n1401));
  jand g1139(.dina(n1401), .dinb(n323), .dout(n1402));
  jor  g1140(.dina(n1402), .dinb(n1382), .dout(n1403));
  jor  g1141(.dina(n796), .dinb(n269), .dout(n1404));
  jor  g1142(.dina(n778), .dinb(shift1 ), .dout(n1405));
  jand g1143(.dina(n1405), .dinb(n1404), .dout(n1406));
  jand g1144(.dina(n1406), .dinb(n266), .dout(n1407));
  jor  g1145(.dina(n806), .dinb(n269), .dout(n1408));
  jor  g1146(.dina(n813), .dinb(shift1 ), .dout(n1409));
  jand g1147(.dina(n1409), .dinb(n1408), .dout(n1410));
  jand g1148(.dina(n1410), .dinb(n281), .dout(n1411));
  jor  g1149(.dina(n1411), .dinb(n1407), .dout(n1412));
  jor  g1150(.dina(n817), .dinb(n269), .dout(n1413));
  jor  g1151(.dina(n792), .dinb(shift1 ), .dout(n1414));
  jand g1152(.dina(n1414), .dinb(n1413), .dout(n1415));
  jand g1153(.dina(n1415), .dinb(n295), .dout(n1416));
  jor  g1154(.dina(n827), .dinb(n269), .dout(n1417));
  jor  g1155(.dina(n802), .dinb(shift1 ), .dout(n1418));
  jand g1156(.dina(n1418), .dinb(n1417), .dout(n1419));
  jand g1157(.dina(n1419), .dinb(n308), .dout(n1420));
  jor  g1158(.dina(n1420), .dinb(n1416), .dout(n1421));
  jor  g1159(.dina(n1421), .dinb(n1412), .dout(n1422));
  jand g1160(.dina(n1422), .dinb(n432), .dout(n1423));
  jor  g1161(.dina(n840), .dinb(n269), .dout(n1424));
  jor  g1162(.dina(n1003), .dinb(shift1 ), .dout(n1425));
  jand g1163(.dina(n1425), .dinb(n1424), .dout(n1426));
  jand g1164(.dina(n1426), .dinb(n266), .dout(n1427));
  jor  g1165(.dina(n850), .dinb(n269), .dout(n1428));
  jor  g1166(.dina(n857), .dinb(shift1 ), .dout(n1429));
  jand g1167(.dina(n1429), .dinb(n1428), .dout(n1430));
  jand g1168(.dina(n1430), .dinb(n281), .dout(n1431));
  jor  g1169(.dina(n1431), .dinb(n1427), .dout(n1432));
  jor  g1170(.dina(n861), .dinb(n269), .dout(n1433));
  jor  g1171(.dina(n836), .dinb(shift1 ), .dout(n1434));
  jand g1172(.dina(n1434), .dinb(n1433), .dout(n1435));
  jand g1173(.dina(n1435), .dinb(n295), .dout(n1436));
  jor  g1174(.dina(n871), .dinb(n269), .dout(n1437));
  jor  g1175(.dina(n846), .dinb(shift1 ), .dout(n1438));
  jand g1176(.dina(n1438), .dinb(n1437), .dout(n1439));
  jand g1177(.dina(n1439), .dinb(n308), .dout(n1440));
  jor  g1178(.dina(n1440), .dinb(n1436), .dout(n1441));
  jor  g1179(.dina(n1441), .dinb(n1432), .dout(n1442));
  jand g1180(.dina(n1442), .dinb(n485), .dout(n1443));
  jor  g1181(.dina(n1443), .dinb(n1423), .dout(n1444));
  jor  g1182(.dina(n1444), .dinb(n1403), .dout(n1445));
  jand g1183(.dina(n1445), .dinb(n263), .dout(n1446));
  jor  g1184(.dina(n887), .dinb(n269), .dout(n1447));
  jor  g1185(.dina(n734), .dinb(shift1 ), .dout(n1448));
  jand g1186(.dina(n1448), .dinb(n1447), .dout(n1449));
  jand g1187(.dina(n1449), .dinb(n266), .dout(n1450));
  jor  g1188(.dina(n897), .dinb(n269), .dout(n1451));
  jor  g1189(.dina(n904), .dinb(shift1 ), .dout(n1452));
  jand g1190(.dina(n1452), .dinb(n1451), .dout(n1453));
  jand g1191(.dina(n1453), .dinb(n281), .dout(n1454));
  jor  g1192(.dina(n1454), .dinb(n1450), .dout(n1455));
  jor  g1193(.dina(n908), .dinb(n269), .dout(n1456));
  jor  g1194(.dina(n883), .dinb(shift1 ), .dout(n1457));
  jand g1195(.dina(n1457), .dinb(n1456), .dout(n1458));
  jand g1196(.dina(n1458), .dinb(n295), .dout(n1459));
  jor  g1197(.dina(n918), .dinb(n269), .dout(n1460));
  jor  g1198(.dina(n893), .dinb(shift1 ), .dout(n1461));
  jand g1199(.dina(n1461), .dinb(n1460), .dout(n1462));
  jand g1200(.dina(n1462), .dinb(n308), .dout(n1463));
  jor  g1201(.dina(n1463), .dinb(n1459), .dout(n1464));
  jor  g1202(.dina(n1464), .dinb(n1455), .dout(n1465));
  jand g1203(.dina(n1465), .dinb(n485), .dout(n1466));
  jor  g1204(.dina(n931), .dinb(n269), .dout(n1467));
  jor  g1205(.dina(n1051), .dinb(shift1 ), .dout(n1468));
  jand g1206(.dina(n1468), .dinb(n1467), .dout(n1469));
  jand g1207(.dina(n1469), .dinb(n266), .dout(n1470));
  jor  g1208(.dina(n941), .dinb(n269), .dout(n1471));
  jor  g1209(.dina(n948), .dinb(shift1 ), .dout(n1472));
  jand g1210(.dina(n1472), .dinb(n1471), .dout(n1473));
  jand g1211(.dina(n1473), .dinb(n281), .dout(n1474));
  jor  g1212(.dina(n1474), .dinb(n1470), .dout(n1475));
  jor  g1213(.dina(n952), .dinb(n269), .dout(n1476));
  jor  g1214(.dina(n927), .dinb(shift1 ), .dout(n1477));
  jand g1215(.dina(n1477), .dinb(n1476), .dout(n1478));
  jand g1216(.dina(n1478), .dinb(n295), .dout(n1479));
  jor  g1217(.dina(n962), .dinb(n269), .dout(n1480));
  jor  g1218(.dina(n937), .dinb(shift1 ), .dout(n1481));
  jand g1219(.dina(n1481), .dinb(n1480), .dout(n1482));
  jand g1220(.dina(n1482), .dinb(n308), .dout(n1483));
  jor  g1221(.dina(n1483), .dinb(n1479), .dout(n1484));
  jor  g1222(.dina(n1484), .dinb(n1475), .dout(n1485));
  jand g1223(.dina(n1485), .dinb(n432), .dout(n1486));
  jor  g1224(.dina(n1486), .dinb(n1466), .dout(n1487));
  jor  g1225(.dina(n1016), .dinb(n269), .dout(n1488));
  jor  g1226(.dina(n914), .dinb(shift1 ), .dout(n1489));
  jand g1227(.dina(n1489), .dinb(n1488), .dout(n1490));
  jand g1228(.dina(n1490), .dinb(n266), .dout(n1491));
  jor  g1229(.dina(n1031), .dinb(n1026), .dout(n1492));
  jand g1230(.dina(n1492), .dinb(shift1 ), .dout(n1493));
  jor  g1231(.dina(n1042), .dinb(n1039), .dout(n1494));
  jand g1232(.dina(n1494), .dinb(n269), .dout(n1495));
  jor  g1233(.dina(n1495), .dinb(n1493), .dout(n1496));
  jand g1234(.dina(n1496), .dinb(n281), .dout(n1497));
  jor  g1235(.dina(n1497), .dinb(n1491), .dout(n1498));
  jor  g1236(.dina(n1019), .dinb(shift1 ), .dout(n1499));
  jor  g1237(.dina(n1044), .dinb(n269), .dout(n1500));
  jand g1238(.dina(n1500), .dinb(n1499), .dout(n1501));
  jand g1239(.dina(n1037), .dinb(shift1 ), .dout(n1502));
  jand g1240(.dina(n1018), .dinb(n269), .dout(n1503));
  jor  g1241(.dina(n1503), .dinb(n1502), .dout(n1504));
  jor  g1242(.dina(n1504), .dinb(n1501), .dout(n1505));
  jand g1243(.dina(n1505), .dinb(n295), .dout(n1506));
  jand g1244(.dina(n1055), .dinb(shift1 ), .dout(n1507));
  jor  g1245(.dina(n1029), .dinb(n1024), .dout(n1508));
  jand g1246(.dina(n1508), .dinb(n269), .dout(n1509));
  jor  g1247(.dina(n1509), .dinb(n1507), .dout(n1510));
  jand g1248(.dina(n1510), .dinb(n308), .dout(n1511));
  jor  g1249(.dina(n1511), .dinb(n1506), .dout(n1512));
  jor  g1250(.dina(n1512), .dinb(n1498), .dout(n1513));
  jand g1251(.dina(n1513), .dinb(n377), .dout(n1514));
  jor  g1252(.dina(n976), .dinb(n269), .dout(n1515));
  jor  g1253(.dina(n958), .dinb(shift1 ), .dout(n1516));
  jand g1254(.dina(n1516), .dinb(n1515), .dout(n1517));
  jand g1255(.dina(n1517), .dinb(n266), .dout(n1518));
  jor  g1256(.dina(n986), .dinb(n269), .dout(n1519));
  jor  g1257(.dina(n993), .dinb(shift1 ), .dout(n1520));
  jand g1258(.dina(n1520), .dinb(n1519), .dout(n1521));
  jand g1259(.dina(n1521), .dinb(n281), .dout(n1522));
  jor  g1260(.dina(n1522), .dinb(n1518), .dout(n1523));
  jor  g1261(.dina(n997), .dinb(n269), .dout(n1524));
  jor  g1262(.dina(n972), .dinb(shift1 ), .dout(n1525));
  jand g1263(.dina(n1525), .dinb(n1524), .dout(n1526));
  jand g1264(.dina(n1526), .dinb(n295), .dout(n1527));
  jor  g1265(.dina(n1007), .dinb(n269), .dout(n1528));
  jor  g1266(.dina(n982), .dinb(shift1 ), .dout(n1529));
  jand g1267(.dina(n1529), .dinb(n1528), .dout(n1530));
  jand g1268(.dina(n1530), .dinb(n308), .dout(n1531));
  jor  g1269(.dina(n1531), .dinb(n1527), .dout(n1532));
  jor  g1270(.dina(n1532), .dinb(n1523), .dout(n1533));
  jand g1271(.dina(n1533), .dinb(n323), .dout(n1534));
  jor  g1272(.dina(n1534), .dinb(n1514), .dout(n1535));
  jor  g1273(.dina(n1535), .dinb(n1487), .dout(n1536));
  jand g1274(.dina(n1536), .dinb(shift6 ), .dout(n1537));
  jor  g1275(.dina(n1537), .dinb(n1446), .dout(result3 ));
  jand g1276(.dina(n427), .dinb(n266), .dout(n1539));
  jand g1277(.dina(n306), .dinb(n281), .dout(n1540));
  jor  g1278(.dina(n1540), .dinb(n1539), .dout(n1541));
  jand g1279(.dina(n295), .dinb(n279), .dout(n1542));
  jand g1280(.dina(n308), .dinb(n292), .dout(n1543));
  jor  g1281(.dina(n1543), .dinb(n1542), .dout(n1544));
  jor  g1282(.dina(n1544), .dinb(n1541), .dout(n1545));
  jand g1283(.dina(n1545), .dinb(n323), .dout(n1546));
  jand g1284(.dina(n481), .dinb(n266), .dout(n1547));
  jand g1285(.dina(n360), .dinb(n281), .dout(n1548));
  jor  g1286(.dina(n1548), .dinb(n1547), .dout(n1549));
  jand g1287(.dina(n335), .dinb(n295), .dout(n1550));
  jand g1288(.dina(n347), .dinb(n308), .dout(n1551));
  jor  g1289(.dina(n1551), .dinb(n1550), .dout(n1552));
  jor  g1290(.dina(n1552), .dinb(n1549), .dout(n1553));
  jand g1291(.dina(n1553), .dinb(n377), .dout(n1554));
  jor  g1292(.dina(n1554), .dinb(n1546), .dout(n1555));
  jand g1293(.dina(n372), .dinb(n266), .dout(n1556));
  jand g1294(.dina(n415), .dinb(n281), .dout(n1557));
  jor  g1295(.dina(n1557), .dinb(n1556), .dout(n1558));
  jand g1296(.dina(n390), .dinb(n295), .dout(n1559));
  jand g1297(.dina(n402), .dinb(n308), .dout(n1560));
  jor  g1298(.dina(n1560), .dinb(n1559), .dout(n1561));
  jor  g1299(.dina(n1561), .dinb(n1558), .dout(n1562));
  jand g1300(.dina(n1562), .dinb(n432), .dout(n1563));
  jand g1301(.dina(n537), .dinb(n266), .dout(n1564));
  jand g1302(.dina(n469), .dinb(n281), .dout(n1565));
  jor  g1303(.dina(n1565), .dinb(n1564), .dout(n1566));
  jand g1304(.dina(n444), .dinb(n295), .dout(n1567));
  jand g1305(.dina(n456), .dinb(n308), .dout(n1568));
  jor  g1306(.dina(n1568), .dinb(n1567), .dout(n1569));
  jor  g1307(.dina(n1569), .dinb(n1566), .dout(n1570));
  jand g1308(.dina(n1570), .dinb(n485), .dout(n1571));
  jor  g1309(.dina(n1571), .dinb(n1563), .dout(n1572));
  jor  g1310(.dina(n1572), .dinb(n1555), .dout(n1573));
  jand g1311(.dina(n1573), .dinb(n263), .dout(n1574));
  jand g1312(.dina(n692), .dinb(n266), .dout(n1575));
  jand g1313(.dina(n575), .dinb(n281), .dout(n1576));
  jor  g1314(.dina(n1576), .dinb(n1575), .dout(n1577));
  jand g1315(.dina(n552), .dinb(n295), .dout(n1578));
  jand g1316(.dina(n562), .dinb(n308), .dout(n1579));
  jor  g1317(.dina(n1579), .dinb(n1578), .dout(n1580));
  jor  g1318(.dina(n1580), .dinb(n1577), .dout(n1581));
  jand g1319(.dina(n1581), .dinb(n377), .dout(n1582));
  jand g1320(.dina(n640), .dinb(n266), .dout(n1583));
  jand g1321(.dina(n525), .dinb(n281), .dout(n1584));
  jor  g1322(.dina(n1584), .dinb(n1583), .dout(n1585));
  jand g1323(.dina(n500), .dinb(n295), .dout(n1586));
  jand g1324(.dina(n512), .dinb(n308), .dout(n1587));
  jor  g1325(.dina(n1587), .dinb(n1586), .dout(n1588));
  jor  g1326(.dina(n1588), .dinb(n1585), .dout(n1589));
  jand g1327(.dina(n1589), .dinb(n323), .dout(n1590));
  jor  g1328(.dina(n1590), .dinb(n1582), .dout(n1591));
  jand g1329(.dina(n319), .dinb(n266), .dout(n1592));
  jand g1330(.dina(n680), .dinb(n281), .dout(n1593));
  jor  g1331(.dina(n1593), .dinb(n1592), .dout(n1594));
  jand g1332(.dina(n655), .dinb(n295), .dout(n1595));
  jand g1333(.dina(n667), .dinb(n308), .dout(n1596));
  jor  g1334(.dina(n1596), .dinb(n1595), .dout(n1597));
  jor  g1335(.dina(n1597), .dinb(n1594), .dout(n1598));
  jand g1336(.dina(n1598), .dinb(n485), .dout(n1599));
  jand g1337(.dina(n587), .dinb(n266), .dout(n1600));
  jand g1338(.dina(n628), .dinb(n281), .dout(n1601));
  jor  g1339(.dina(n1601), .dinb(n1600), .dout(n1602));
  jand g1340(.dina(n603), .dinb(n295), .dout(n1603));
  jand g1341(.dina(n615), .dinb(n308), .dout(n1604));
  jor  g1342(.dina(n1604), .dinb(n1603), .dout(n1605));
  jor  g1343(.dina(n1605), .dinb(n1602), .dout(n1606));
  jand g1344(.dina(n1606), .dinb(n432), .dout(n1607));
  jor  g1345(.dina(n1607), .dinb(n1599), .dout(n1608));
  jor  g1346(.dina(n1608), .dinb(n1591), .dout(n1609));
  jand g1347(.dina(n1609), .dinb(shift6 ), .dout(n1610));
  jor  g1348(.dina(n1610), .dinb(n1574), .dout(result4 ));
  jand g1349(.dina(n829), .dinb(n266), .dout(n1612));
  jand g1350(.dina(n730), .dinb(n281), .dout(n1613));
  jor  g1351(.dina(n1613), .dinb(n1612), .dout(n1614));
  jand g1352(.dina(n709), .dinb(n295), .dout(n1615));
  jand g1353(.dina(n719), .dinb(n308), .dout(n1616));
  jor  g1354(.dina(n1616), .dinb(n1615), .dout(n1617));
  jor  g1355(.dina(n1617), .dinb(n1614), .dout(n1618));
  jand g1356(.dina(n1618), .dinb(n323), .dout(n1619));
  jand g1357(.dina(n873), .dinb(n266), .dout(n1620));
  jand g1358(.dina(n774), .dinb(n281), .dout(n1621));
  jor  g1359(.dina(n1621), .dinb(n1620), .dout(n1622));
  jand g1360(.dina(n753), .dinb(n295), .dout(n1623));
  jand g1361(.dina(n763), .dinb(n308), .dout(n1624));
  jor  g1362(.dina(n1624), .dinb(n1623), .dout(n1625));
  jor  g1363(.dina(n1625), .dinb(n1622), .dout(n1626));
  jand g1364(.dina(n1626), .dinb(n377), .dout(n1627));
  jor  g1365(.dina(n1627), .dinb(n1619), .dout(n1628));
  jand g1366(.dina(n784), .dinb(n266), .dout(n1629));
  jand g1367(.dina(n819), .dinb(n281), .dout(n1630));
  jor  g1368(.dina(n1630), .dinb(n1629), .dout(n1631));
  jand g1369(.dina(n798), .dinb(n295), .dout(n1632));
  jand g1370(.dina(n808), .dinb(n308), .dout(n1633));
  jor  g1371(.dina(n1633), .dinb(n1632), .dout(n1634));
  jor  g1372(.dina(n1634), .dinb(n1631), .dout(n1635));
  jand g1373(.dina(n1635), .dinb(n432), .dout(n1636));
  jand g1374(.dina(n1009), .dinb(n266), .dout(n1637));
  jand g1375(.dina(n863), .dinb(n281), .dout(n1638));
  jor  g1376(.dina(n1638), .dinb(n1637), .dout(n1639));
  jand g1377(.dina(n842), .dinb(n295), .dout(n1640));
  jand g1378(.dina(n852), .dinb(n308), .dout(n1641));
  jor  g1379(.dina(n1641), .dinb(n1640), .dout(n1642));
  jor  g1380(.dina(n1642), .dinb(n1639), .dout(n1643));
  jand g1381(.dina(n1643), .dinb(n485), .dout(n1644));
  jor  g1382(.dina(n1644), .dinb(n1636), .dout(n1645));
  jor  g1383(.dina(n1645), .dinb(n1628), .dout(n1646));
  jand g1384(.dina(n1646), .dinb(n263), .dout(n1647));
  jand g1385(.dina(n920), .dinb(n266), .dout(n1648));
  jand g1386(.dina(n1047), .dinb(n281), .dout(n1649));
  jor  g1387(.dina(n1649), .dinb(n1648), .dout(n1650));
  jand g1388(.dina(n1022), .dinb(n295), .dout(n1651));
  jand g1389(.dina(n1034), .dinb(n308), .dout(n1652));
  jor  g1390(.dina(n1652), .dinb(n1651), .dout(n1653));
  jor  g1391(.dina(n1653), .dinb(n1650), .dout(n1654));
  jand g1392(.dina(n1654), .dinb(n377), .dout(n1655));
  jand g1393(.dina(n964), .dinb(n266), .dout(n1656));
  jand g1394(.dina(n999), .dinb(n281), .dout(n1657));
  jor  g1395(.dina(n1657), .dinb(n1656), .dout(n1658));
  jand g1396(.dina(n978), .dinb(n295), .dout(n1659));
  jand g1397(.dina(n988), .dinb(n308), .dout(n1660));
  jor  g1398(.dina(n1660), .dinb(n1659), .dout(n1661));
  jor  g1399(.dina(n1661), .dinb(n1658), .dout(n1662));
  jand g1400(.dina(n1662), .dinb(n323), .dout(n1663));
  jor  g1401(.dina(n1663), .dinb(n1655), .dout(n1664));
  jand g1402(.dina(n740), .dinb(n266), .dout(n1665));
  jand g1403(.dina(n910), .dinb(n281), .dout(n1666));
  jor  g1404(.dina(n1666), .dinb(n1665), .dout(n1667));
  jand g1405(.dina(n889), .dinb(n295), .dout(n1668));
  jand g1406(.dina(n899), .dinb(n308), .dout(n1669));
  jor  g1407(.dina(n1669), .dinb(n1668), .dout(n1670));
  jor  g1408(.dina(n1670), .dinb(n1667), .dout(n1671));
  jand g1409(.dina(n1671), .dinb(n485), .dout(n1672));
  jand g1410(.dina(n1057), .dinb(n266), .dout(n1673));
  jand g1411(.dina(n954), .dinb(n281), .dout(n1674));
  jor  g1412(.dina(n1674), .dinb(n1673), .dout(n1675));
  jand g1413(.dina(n933), .dinb(n295), .dout(n1676));
  jand g1414(.dina(n943), .dinb(n308), .dout(n1677));
  jor  g1415(.dina(n1677), .dinb(n1676), .dout(n1678));
  jor  g1416(.dina(n1678), .dinb(n1675), .dout(n1679));
  jand g1417(.dina(n1679), .dinb(n432), .dout(n1680));
  jor  g1418(.dina(n1680), .dinb(n1672), .dout(n1681));
  jor  g1419(.dina(n1681), .dinb(n1664), .dout(n1682));
  jand g1420(.dina(n1682), .dinb(shift6 ), .dout(n1683));
  jor  g1421(.dina(n1683), .dinb(n1647), .dout(result5 ));
  jand g1422(.dina(n1170), .dinb(n266), .dout(n1685));
  jand g1423(.dina(n1089), .dinb(n281), .dout(n1686));
  jor  g1424(.dina(n1686), .dinb(n1685), .dout(n1687));
  jand g1425(.dina(n1072), .dinb(n295), .dout(n1688));
  jand g1426(.dina(n1080), .dinb(n308), .dout(n1689));
  jor  g1427(.dina(n1689), .dinb(n1688), .dout(n1690));
  jor  g1428(.dina(n1690), .dinb(n1687), .dout(n1691));
  jand g1429(.dina(n1691), .dinb(n323), .dout(n1692));
  jand g1430(.dina(n1206), .dinb(n266), .dout(n1693));
  jand g1431(.dina(n1125), .dinb(n281), .dout(n1694));
  jor  g1432(.dina(n1694), .dinb(n1693), .dout(n1695));
  jand g1433(.dina(n1108), .dinb(n295), .dout(n1696));
  jand g1434(.dina(n1116), .dinb(n308), .dout(n1697));
  jor  g1435(.dina(n1697), .dinb(n1696), .dout(n1698));
  jor  g1436(.dina(n1698), .dinb(n1695), .dout(n1699));
  jand g1437(.dina(n1699), .dinb(n377), .dout(n1700));
  jor  g1438(.dina(n1700), .dinb(n1692), .dout(n1701));
  jand g1439(.dina(n1133), .dinb(n266), .dout(n1702));
  jand g1440(.dina(n1162), .dinb(n281), .dout(n1703));
  jor  g1441(.dina(n1703), .dinb(n1702), .dout(n1704));
  jand g1442(.dina(n1145), .dinb(n295), .dout(n1705));
  jand g1443(.dina(n1153), .dinb(n308), .dout(n1706));
  jor  g1444(.dina(n1706), .dinb(n1705), .dout(n1707));
  jor  g1445(.dina(n1707), .dinb(n1704), .dout(n1708));
  jand g1446(.dina(n1708), .dinb(n432), .dout(n1709));
  jand g1447(.dina(n1318), .dinb(n266), .dout(n1710));
  jand g1448(.dina(n1198), .dinb(n281), .dout(n1711));
  jor  g1449(.dina(n1711), .dinb(n1710), .dout(n1712));
  jand g1450(.dina(n1181), .dinb(n295), .dout(n1713));
  jand g1451(.dina(n1189), .dinb(n308), .dout(n1714));
  jor  g1452(.dina(n1714), .dinb(n1713), .dout(n1715));
  jor  g1453(.dina(n1715), .dinb(n1712), .dout(n1716));
  jand g1454(.dina(n1716), .dinb(n485), .dout(n1717));
  jor  g1455(.dina(n1717), .dinb(n1709), .dout(n1718));
  jor  g1456(.dina(n1718), .dinb(n1701), .dout(n1719));
  jand g1457(.dina(n1719), .dinb(n263), .dout(n1720));
  jand g1458(.dina(n1245), .dinb(n266), .dout(n1721));
  jand g1459(.dina(n1346), .dinb(n281), .dout(n1722));
  jor  g1460(.dina(n1722), .dinb(n1721), .dout(n1723));
  jand g1461(.dina(n1329), .dinb(n295), .dout(n1724));
  jand g1462(.dina(n1337), .dinb(n308), .dout(n1725));
  jor  g1463(.dina(n1725), .dinb(n1724), .dout(n1726));
  jor  g1464(.dina(n1726), .dinb(n1723), .dout(n1727));
  jand g1465(.dina(n1727), .dinb(n377), .dout(n1728));
  jand g1466(.dina(n1281), .dinb(n266), .dout(n1729));
  jand g1467(.dina(n1310), .dinb(n281), .dout(n1730));
  jor  g1468(.dina(n1730), .dinb(n1729), .dout(n1731));
  jand g1469(.dina(n1293), .dinb(n295), .dout(n1732));
  jand g1470(.dina(n1301), .dinb(n308), .dout(n1733));
  jor  g1471(.dina(n1733), .dinb(n1732), .dout(n1734));
  jor  g1472(.dina(n1734), .dinb(n1731), .dout(n1735));
  jand g1473(.dina(n1735), .dinb(n323), .dout(n1736));
  jor  g1474(.dina(n1736), .dinb(n1728), .dout(n1737));
  jand g1475(.dina(n1097), .dinb(n266), .dout(n1738));
  jand g1476(.dina(n1237), .dinb(n281), .dout(n1739));
  jor  g1477(.dina(n1739), .dinb(n1738), .dout(n1740));
  jand g1478(.dina(n1220), .dinb(n295), .dout(n1741));
  jand g1479(.dina(n1228), .dinb(n308), .dout(n1742));
  jor  g1480(.dina(n1742), .dinb(n1741), .dout(n1743));
  jor  g1481(.dina(n1743), .dinb(n1740), .dout(n1744));
  jand g1482(.dina(n1744), .dinb(n485), .dout(n1745));
  jand g1483(.dina(n1354), .dinb(n266), .dout(n1746));
  jand g1484(.dina(n1273), .dinb(n281), .dout(n1747));
  jor  g1485(.dina(n1747), .dinb(n1746), .dout(n1748));
  jand g1486(.dina(n1256), .dinb(n295), .dout(n1749));
  jand g1487(.dina(n1264), .dinb(n308), .dout(n1750));
  jor  g1488(.dina(n1750), .dinb(n1749), .dout(n1751));
  jor  g1489(.dina(n1751), .dinb(n1748), .dout(n1752));
  jand g1490(.dina(n1752), .dinb(n432), .dout(n1753));
  jor  g1491(.dina(n1753), .dinb(n1745), .dout(n1754));
  jor  g1492(.dina(n1754), .dinb(n1737), .dout(n1755));
  jand g1493(.dina(n1755), .dinb(shift6 ), .dout(n1756));
  jor  g1494(.dina(n1756), .dinb(n1720), .dout(result6 ));
  jand g1495(.dina(n1419), .dinb(n266), .dout(n1758));
  jand g1496(.dina(n1394), .dinb(n281), .dout(n1759));
  jor  g1497(.dina(n1759), .dinb(n1758), .dout(n1760));
  jand g1498(.dina(n1385), .dinb(n295), .dout(n1761));
  jand g1499(.dina(n1389), .dinb(n308), .dout(n1762));
  jor  g1500(.dina(n1762), .dinb(n1761), .dout(n1763));
  jor  g1501(.dina(n1763), .dinb(n1760), .dout(n1764));
  jand g1502(.dina(n1764), .dinb(n323), .dout(n1765));
  jand g1503(.dina(n1439), .dinb(n266), .dout(n1766));
  jand g1504(.dina(n1374), .dinb(n281), .dout(n1767));
  jor  g1505(.dina(n1767), .dinb(n1766), .dout(n1768));
  jand g1506(.dina(n1365), .dinb(n295), .dout(n1769));
  jand g1507(.dina(n1369), .dinb(n308), .dout(n1770));
  jor  g1508(.dina(n1770), .dinb(n1769), .dout(n1771));
  jor  g1509(.dina(n1771), .dinb(n1768), .dout(n1772));
  jand g1510(.dina(n1772), .dinb(n377), .dout(n1773));
  jor  g1511(.dina(n1773), .dinb(n1765), .dout(n1774));
  jand g1512(.dina(n1378), .dinb(n266), .dout(n1775));
  jand g1513(.dina(n1415), .dinb(n281), .dout(n1776));
  jor  g1514(.dina(n1776), .dinb(n1775), .dout(n1777));
  jand g1515(.dina(n1406), .dinb(n295), .dout(n1778));
  jand g1516(.dina(n1410), .dinb(n308), .dout(n1779));
  jor  g1517(.dina(n1779), .dinb(n1778), .dout(n1780));
  jor  g1518(.dina(n1780), .dinb(n1777), .dout(n1781));
  jand g1519(.dina(n1781), .dinb(n432), .dout(n1782));
  jand g1520(.dina(n1530), .dinb(n266), .dout(n1783));
  jand g1521(.dina(n1435), .dinb(n281), .dout(n1784));
  jor  g1522(.dina(n1784), .dinb(n1783), .dout(n1785));
  jand g1523(.dina(n1426), .dinb(n295), .dout(n1786));
  jand g1524(.dina(n1430), .dinb(n308), .dout(n1787));
  jor  g1525(.dina(n1787), .dinb(n1786), .dout(n1788));
  jor  g1526(.dina(n1788), .dinb(n1785), .dout(n1789));
  jand g1527(.dina(n1789), .dinb(n485), .dout(n1790));
  jor  g1528(.dina(n1790), .dinb(n1782), .dout(n1791));
  jor  g1529(.dina(n1791), .dinb(n1774), .dout(n1792));
  jand g1530(.dina(n1792), .dinb(n263), .dout(n1793));
  jand g1531(.dina(n1490), .dinb(n295), .dout(n1794));
  jand g1532(.dina(n1462), .dinb(n266), .dout(n1795));
  jor  g1533(.dina(n1795), .dinb(n1794), .dout(n1796));
  jand g1534(.dina(n1505), .dinb(n281), .dout(n1797));
  jand g1535(.dina(n1496), .dinb(n308), .dout(n1798));
  jor  g1536(.dina(n1798), .dinb(n1797), .dout(n1799));
  jor  g1537(.dina(n1799), .dinb(n1796), .dout(n1800));
  jand g1538(.dina(n1800), .dinb(n377), .dout(n1801));
  jand g1539(.dina(n1482), .dinb(n266), .dout(n1802));
  jand g1540(.dina(n1526), .dinb(n281), .dout(n1803));
  jor  g1541(.dina(n1803), .dinb(n1802), .dout(n1804));
  jand g1542(.dina(n1517), .dinb(n295), .dout(n1805));
  jand g1543(.dina(n1521), .dinb(n308), .dout(n1806));
  jor  g1544(.dina(n1806), .dinb(n1805), .dout(n1807));
  jor  g1545(.dina(n1807), .dinb(n1804), .dout(n1808));
  jand g1546(.dina(n1808), .dinb(n323), .dout(n1809));
  jor  g1547(.dina(n1809), .dinb(n1801), .dout(n1810));
  jand g1548(.dina(n1398), .dinb(n266), .dout(n1811));
  jand g1549(.dina(n1458), .dinb(n281), .dout(n1812));
  jor  g1550(.dina(n1812), .dinb(n1811), .dout(n1813));
  jand g1551(.dina(n1449), .dinb(n295), .dout(n1814));
  jand g1552(.dina(n1453), .dinb(n308), .dout(n1815));
  jor  g1553(.dina(n1815), .dinb(n1814), .dout(n1816));
  jor  g1554(.dina(n1816), .dinb(n1813), .dout(n1817));
  jand g1555(.dina(n1817), .dinb(n485), .dout(n1818));
  jand g1556(.dina(n1510), .dinb(n266), .dout(n1819));
  jand g1557(.dina(n1478), .dinb(n281), .dout(n1820));
  jor  g1558(.dina(n1820), .dinb(n1819), .dout(n1821));
  jand g1559(.dina(n1469), .dinb(n295), .dout(n1822));
  jand g1560(.dina(n1473), .dinb(n308), .dout(n1823));
  jor  g1561(.dina(n1823), .dinb(n1822), .dout(n1824));
  jor  g1562(.dina(n1824), .dinb(n1821), .dout(n1825));
  jand g1563(.dina(n1825), .dinb(n432), .dout(n1826));
  jor  g1564(.dina(n1826), .dinb(n1818), .dout(n1827));
  jor  g1565(.dina(n1827), .dinb(n1810), .dout(n1828));
  jand g1566(.dina(n1828), .dinb(shift6 ), .dout(n1829));
  jor  g1567(.dina(n1829), .dinb(n1793), .dout(result7 ));
  jand g1568(.dina(n402), .dinb(n266), .dout(n1831));
  jand g1569(.dina(n281), .dinb(n279), .dout(n1832));
  jor  g1570(.dina(n1832), .dinb(n1831), .dout(n1833));
  jand g1571(.dina(n427), .dinb(n295), .dout(n1834));
  jand g1572(.dina(n308), .dinb(n306), .dout(n1835));
  jor  g1573(.dina(n1835), .dinb(n1834), .dout(n1836));
  jor  g1574(.dina(n1836), .dinb(n1833), .dout(n1837));
  jand g1575(.dina(n1837), .dinb(n323), .dout(n1838));
  jand g1576(.dina(n456), .dinb(n266), .dout(n1839));
  jand g1577(.dina(n335), .dinb(n281), .dout(n1840));
  jor  g1578(.dina(n1840), .dinb(n1839), .dout(n1841));
  jand g1579(.dina(n481), .dinb(n295), .dout(n1842));
  jand g1580(.dina(n360), .dinb(n308), .dout(n1843));
  jor  g1581(.dina(n1843), .dinb(n1842), .dout(n1844));
  jor  g1582(.dina(n1844), .dinb(n1841), .dout(n1845));
  jand g1583(.dina(n1845), .dinb(n377), .dout(n1846));
  jor  g1584(.dina(n1846), .dinb(n1838), .dout(n1847));
  jand g1585(.dina(n347), .dinb(n266), .dout(n1848));
  jand g1586(.dina(n390), .dinb(n281), .dout(n1849));
  jor  g1587(.dina(n1849), .dinb(n1848), .dout(n1850));
  jand g1588(.dina(n372), .dinb(n295), .dout(n1851));
  jand g1589(.dina(n415), .dinb(n308), .dout(n1852));
  jor  g1590(.dina(n1852), .dinb(n1851), .dout(n1853));
  jor  g1591(.dina(n1853), .dinb(n1850), .dout(n1854));
  jand g1592(.dina(n1854), .dinb(n432), .dout(n1855));
  jand g1593(.dina(n512), .dinb(n266), .dout(n1856));
  jand g1594(.dina(n444), .dinb(n281), .dout(n1857));
  jor  g1595(.dina(n1857), .dinb(n1856), .dout(n1858));
  jand g1596(.dina(n537), .dinb(n295), .dout(n1859));
  jand g1597(.dina(n469), .dinb(n308), .dout(n1860));
  jor  g1598(.dina(n1860), .dinb(n1859), .dout(n1861));
  jor  g1599(.dina(n1861), .dinb(n1858), .dout(n1862));
  jand g1600(.dina(n1862), .dinb(n485), .dout(n1863));
  jor  g1601(.dina(n1863), .dinb(n1855), .dout(n1864));
  jor  g1602(.dina(n1864), .dinb(n1847), .dout(n1865));
  jand g1603(.dina(n1865), .dinb(n263), .dout(n1866));
  jand g1604(.dina(n667), .dinb(n266), .dout(n1867));
  jand g1605(.dina(n552), .dinb(n281), .dout(n1868));
  jor  g1606(.dina(n1868), .dinb(n1867), .dout(n1869));
  jand g1607(.dina(n692), .dinb(n295), .dout(n1870));
  jand g1608(.dina(n575), .dinb(n308), .dout(n1871));
  jor  g1609(.dina(n1871), .dinb(n1870), .dout(n1872));
  jor  g1610(.dina(n1872), .dinb(n1869), .dout(n1873));
  jand g1611(.dina(n1873), .dinb(n377), .dout(n1874));
  jand g1612(.dina(n615), .dinb(n266), .dout(n1875));
  jand g1613(.dina(n500), .dinb(n281), .dout(n1876));
  jor  g1614(.dina(n1876), .dinb(n1875), .dout(n1877));
  jand g1615(.dina(n640), .dinb(n295), .dout(n1878));
  jand g1616(.dina(n525), .dinb(n308), .dout(n1879));
  jor  g1617(.dina(n1879), .dinb(n1878), .dout(n1880));
  jor  g1618(.dina(n1880), .dinb(n1877), .dout(n1881));
  jand g1619(.dina(n1881), .dinb(n323), .dout(n1882));
  jor  g1620(.dina(n1882), .dinb(n1874), .dout(n1883));
  jand g1621(.dina(n292), .dinb(n266), .dout(n1884));
  jand g1622(.dina(n655), .dinb(n281), .dout(n1885));
  jor  g1623(.dina(n1885), .dinb(n1884), .dout(n1886));
  jand g1624(.dina(n319), .dinb(n295), .dout(n1887));
  jand g1625(.dina(n680), .dinb(n308), .dout(n1888));
  jor  g1626(.dina(n1888), .dinb(n1887), .dout(n1889));
  jor  g1627(.dina(n1889), .dinb(n1886), .dout(n1890));
  jand g1628(.dina(n1890), .dinb(n485), .dout(n1891));
  jand g1629(.dina(n562), .dinb(n266), .dout(n1892));
  jand g1630(.dina(n603), .dinb(n281), .dout(n1893));
  jor  g1631(.dina(n1893), .dinb(n1892), .dout(n1894));
  jand g1632(.dina(n587), .dinb(n295), .dout(n1895));
  jand g1633(.dina(n628), .dinb(n308), .dout(n1896));
  jor  g1634(.dina(n1896), .dinb(n1895), .dout(n1897));
  jor  g1635(.dina(n1897), .dinb(n1894), .dout(n1898));
  jand g1636(.dina(n1898), .dinb(n432), .dout(n1899));
  jor  g1637(.dina(n1899), .dinb(n1891), .dout(n1900));
  jor  g1638(.dina(n1900), .dinb(n1883), .dout(n1901));
  jand g1639(.dina(n1901), .dinb(shift6 ), .dout(n1902));
  jor  g1640(.dina(n1902), .dinb(n1866), .dout(result8 ));
  jand g1641(.dina(n808), .dinb(n266), .dout(n1904));
  jand g1642(.dina(n709), .dinb(n281), .dout(n1905));
  jor  g1643(.dina(n1905), .dinb(n1904), .dout(n1906));
  jand g1644(.dina(n829), .dinb(n295), .dout(n1907));
  jand g1645(.dina(n730), .dinb(n308), .dout(n1908));
  jor  g1646(.dina(n1908), .dinb(n1907), .dout(n1909));
  jor  g1647(.dina(n1909), .dinb(n1906), .dout(n1910));
  jand g1648(.dina(n1910), .dinb(n323), .dout(n1911));
  jand g1649(.dina(n852), .dinb(n266), .dout(n1912));
  jand g1650(.dina(n753), .dinb(n281), .dout(n1913));
  jor  g1651(.dina(n1913), .dinb(n1912), .dout(n1914));
  jand g1652(.dina(n873), .dinb(n295), .dout(n1915));
  jand g1653(.dina(n774), .dinb(n308), .dout(n1916));
  jor  g1654(.dina(n1916), .dinb(n1915), .dout(n1917));
  jor  g1655(.dina(n1917), .dinb(n1914), .dout(n1918));
  jand g1656(.dina(n1918), .dinb(n377), .dout(n1919));
  jor  g1657(.dina(n1919), .dinb(n1911), .dout(n1920));
  jand g1658(.dina(n763), .dinb(n266), .dout(n1921));
  jand g1659(.dina(n798), .dinb(n281), .dout(n1922));
  jor  g1660(.dina(n1922), .dinb(n1921), .dout(n1923));
  jand g1661(.dina(n784), .dinb(n295), .dout(n1924));
  jand g1662(.dina(n819), .dinb(n308), .dout(n1925));
  jor  g1663(.dina(n1925), .dinb(n1924), .dout(n1926));
  jor  g1664(.dina(n1926), .dinb(n1923), .dout(n1927));
  jand g1665(.dina(n1927), .dinb(n432), .dout(n1928));
  jand g1666(.dina(n988), .dinb(n266), .dout(n1929));
  jand g1667(.dina(n842), .dinb(n281), .dout(n1930));
  jor  g1668(.dina(n1930), .dinb(n1929), .dout(n1931));
  jand g1669(.dina(n1009), .dinb(n295), .dout(n1932));
  jand g1670(.dina(n863), .dinb(n308), .dout(n1933));
  jor  g1671(.dina(n1933), .dinb(n1932), .dout(n1934));
  jor  g1672(.dina(n1934), .dinb(n1931), .dout(n1935));
  jand g1673(.dina(n1935), .dinb(n485), .dout(n1936));
  jor  g1674(.dina(n1936), .dinb(n1928), .dout(n1937));
  jor  g1675(.dina(n1937), .dinb(n1920), .dout(n1938));
  jand g1676(.dina(n1938), .dinb(n263), .dout(n1939));
  jand g1677(.dina(n899), .dinb(n266), .dout(n1940));
  jand g1678(.dina(n1022), .dinb(n281), .dout(n1941));
  jor  g1679(.dina(n1941), .dinb(n1940), .dout(n1942));
  jand g1680(.dina(n920), .dinb(n295), .dout(n1943));
  jand g1681(.dina(n1047), .dinb(n308), .dout(n1944));
  jor  g1682(.dina(n1944), .dinb(n1943), .dout(n1945));
  jor  g1683(.dina(n1945), .dinb(n1942), .dout(n1946));
  jand g1684(.dina(n1946), .dinb(n377), .dout(n1947));
  jand g1685(.dina(n943), .dinb(n266), .dout(n1948));
  jand g1686(.dina(n978), .dinb(n281), .dout(n1949));
  jor  g1687(.dina(n1949), .dinb(n1948), .dout(n1950));
  jand g1688(.dina(n964), .dinb(n295), .dout(n1951));
  jand g1689(.dina(n999), .dinb(n308), .dout(n1952));
  jor  g1690(.dina(n1952), .dinb(n1951), .dout(n1953));
  jor  g1691(.dina(n1953), .dinb(n1950), .dout(n1954));
  jand g1692(.dina(n1954), .dinb(n323), .dout(n1955));
  jor  g1693(.dina(n1955), .dinb(n1947), .dout(n1956));
  jand g1694(.dina(n719), .dinb(n266), .dout(n1957));
  jand g1695(.dina(n889), .dinb(n281), .dout(n1958));
  jor  g1696(.dina(n1958), .dinb(n1957), .dout(n1959));
  jand g1697(.dina(n740), .dinb(n295), .dout(n1960));
  jand g1698(.dina(n910), .dinb(n308), .dout(n1961));
  jor  g1699(.dina(n1961), .dinb(n1960), .dout(n1962));
  jor  g1700(.dina(n1962), .dinb(n1959), .dout(n1963));
  jand g1701(.dina(n1963), .dinb(n485), .dout(n1964));
  jand g1702(.dina(n1034), .dinb(n266), .dout(n1965));
  jand g1703(.dina(n933), .dinb(n281), .dout(n1966));
  jor  g1704(.dina(n1966), .dinb(n1965), .dout(n1967));
  jand g1705(.dina(n1057), .dinb(n295), .dout(n1968));
  jand g1706(.dina(n954), .dinb(n308), .dout(n1969));
  jor  g1707(.dina(n1969), .dinb(n1968), .dout(n1970));
  jor  g1708(.dina(n1970), .dinb(n1967), .dout(n1971));
  jand g1709(.dina(n1971), .dinb(n432), .dout(n1972));
  jor  g1710(.dina(n1972), .dinb(n1964), .dout(n1973));
  jor  g1711(.dina(n1973), .dinb(n1956), .dout(n1974));
  jand g1712(.dina(n1974), .dinb(shift6 ), .dout(n1975));
  jor  g1713(.dina(n1975), .dinb(n1939), .dout(result9 ));
  jand g1714(.dina(n1153), .dinb(n266), .dout(n1977));
  jand g1715(.dina(n1072), .dinb(n281), .dout(n1978));
  jor  g1716(.dina(n1978), .dinb(n1977), .dout(n1979));
  jand g1717(.dina(n1170), .dinb(n295), .dout(n1980));
  jand g1718(.dina(n1089), .dinb(n308), .dout(n1981));
  jor  g1719(.dina(n1981), .dinb(n1980), .dout(n1982));
  jor  g1720(.dina(n1982), .dinb(n1979), .dout(n1983));
  jand g1721(.dina(n1983), .dinb(n323), .dout(n1984));
  jand g1722(.dina(n1189), .dinb(n266), .dout(n1985));
  jand g1723(.dina(n1108), .dinb(n281), .dout(n1986));
  jor  g1724(.dina(n1986), .dinb(n1985), .dout(n1987));
  jand g1725(.dina(n1206), .dinb(n295), .dout(n1988));
  jand g1726(.dina(n1125), .dinb(n308), .dout(n1989));
  jor  g1727(.dina(n1989), .dinb(n1988), .dout(n1990));
  jor  g1728(.dina(n1990), .dinb(n1987), .dout(n1991));
  jand g1729(.dina(n1991), .dinb(n377), .dout(n1992));
  jor  g1730(.dina(n1992), .dinb(n1984), .dout(n1993));
  jand g1731(.dina(n1116), .dinb(n266), .dout(n1994));
  jand g1732(.dina(n1145), .dinb(n281), .dout(n1995));
  jor  g1733(.dina(n1995), .dinb(n1994), .dout(n1996));
  jand g1734(.dina(n1133), .dinb(n295), .dout(n1997));
  jand g1735(.dina(n1162), .dinb(n308), .dout(n1998));
  jor  g1736(.dina(n1998), .dinb(n1997), .dout(n1999));
  jor  g1737(.dina(n1999), .dinb(n1996), .dout(n2000));
  jand g1738(.dina(n2000), .dinb(n432), .dout(n2001));
  jand g1739(.dina(n1301), .dinb(n266), .dout(n2002));
  jand g1740(.dina(n1181), .dinb(n281), .dout(n2003));
  jor  g1741(.dina(n2003), .dinb(n2002), .dout(n2004));
  jand g1742(.dina(n1318), .dinb(n295), .dout(n2005));
  jand g1743(.dina(n1198), .dinb(n308), .dout(n2006));
  jor  g1744(.dina(n2006), .dinb(n2005), .dout(n2007));
  jor  g1745(.dina(n2007), .dinb(n2004), .dout(n2008));
  jand g1746(.dina(n2008), .dinb(n485), .dout(n2009));
  jor  g1747(.dina(n2009), .dinb(n2001), .dout(n2010));
  jor  g1748(.dina(n2010), .dinb(n1993), .dout(n2011));
  jand g1749(.dina(n2011), .dinb(n263), .dout(n2012));
  jand g1750(.dina(n1228), .dinb(n266), .dout(n2013));
  jand g1751(.dina(n1329), .dinb(n281), .dout(n2014));
  jor  g1752(.dina(n2014), .dinb(n2013), .dout(n2015));
  jand g1753(.dina(n1245), .dinb(n295), .dout(n2016));
  jand g1754(.dina(n1346), .dinb(n308), .dout(n2017));
  jor  g1755(.dina(n2017), .dinb(n2016), .dout(n2018));
  jor  g1756(.dina(n2018), .dinb(n2015), .dout(n2019));
  jand g1757(.dina(n2019), .dinb(n377), .dout(n2020));
  jand g1758(.dina(n1264), .dinb(n266), .dout(n2021));
  jand g1759(.dina(n1293), .dinb(n281), .dout(n2022));
  jor  g1760(.dina(n2022), .dinb(n2021), .dout(n2023));
  jand g1761(.dina(n1281), .dinb(n295), .dout(n2024));
  jand g1762(.dina(n1310), .dinb(n308), .dout(n2025));
  jor  g1763(.dina(n2025), .dinb(n2024), .dout(n2026));
  jor  g1764(.dina(n2026), .dinb(n2023), .dout(n2027));
  jand g1765(.dina(n2027), .dinb(n323), .dout(n2028));
  jor  g1766(.dina(n2028), .dinb(n2020), .dout(n2029));
  jand g1767(.dina(n1080), .dinb(n266), .dout(n2030));
  jand g1768(.dina(n1220), .dinb(n281), .dout(n2031));
  jor  g1769(.dina(n2031), .dinb(n2030), .dout(n2032));
  jand g1770(.dina(n1097), .dinb(n295), .dout(n2033));
  jand g1771(.dina(n1237), .dinb(n308), .dout(n2034));
  jor  g1772(.dina(n2034), .dinb(n2033), .dout(n2035));
  jor  g1773(.dina(n2035), .dinb(n2032), .dout(n2036));
  jand g1774(.dina(n2036), .dinb(n485), .dout(n2037));
  jand g1775(.dina(n1337), .dinb(n266), .dout(n2038));
  jand g1776(.dina(n1256), .dinb(n281), .dout(n2039));
  jor  g1777(.dina(n2039), .dinb(n2038), .dout(n2040));
  jand g1778(.dina(n1354), .dinb(n295), .dout(n2041));
  jand g1779(.dina(n1273), .dinb(n308), .dout(n2042));
  jor  g1780(.dina(n2042), .dinb(n2041), .dout(n2043));
  jor  g1781(.dina(n2043), .dinb(n2040), .dout(n2044));
  jand g1782(.dina(n2044), .dinb(n432), .dout(n2045));
  jor  g1783(.dina(n2045), .dinb(n2037), .dout(n2046));
  jor  g1784(.dina(n2046), .dinb(n2029), .dout(n2047));
  jand g1785(.dina(n2047), .dinb(shift6 ), .dout(n2048));
  jor  g1786(.dina(n2048), .dinb(n2012), .dout(result10 ));
  jand g1787(.dina(n1410), .dinb(n266), .dout(n2050));
  jand g1788(.dina(n1385), .dinb(n281), .dout(n2051));
  jor  g1789(.dina(n2051), .dinb(n2050), .dout(n2052));
  jand g1790(.dina(n1419), .dinb(n295), .dout(n2053));
  jand g1791(.dina(n1394), .dinb(n308), .dout(n2054));
  jor  g1792(.dina(n2054), .dinb(n2053), .dout(n2055));
  jor  g1793(.dina(n2055), .dinb(n2052), .dout(n2056));
  jand g1794(.dina(n2056), .dinb(n323), .dout(n2057));
  jand g1795(.dina(n1430), .dinb(n266), .dout(n2058));
  jand g1796(.dina(n1365), .dinb(n281), .dout(n2059));
  jor  g1797(.dina(n2059), .dinb(n2058), .dout(n2060));
  jand g1798(.dina(n1439), .dinb(n295), .dout(n2061));
  jand g1799(.dina(n1374), .dinb(n308), .dout(n2062));
  jor  g1800(.dina(n2062), .dinb(n2061), .dout(n2063));
  jor  g1801(.dina(n2063), .dinb(n2060), .dout(n2064));
  jand g1802(.dina(n2064), .dinb(n377), .dout(n2065));
  jor  g1803(.dina(n2065), .dinb(n2057), .dout(n2066));
  jand g1804(.dina(n1369), .dinb(n266), .dout(n2067));
  jand g1805(.dina(n1406), .dinb(n281), .dout(n2068));
  jor  g1806(.dina(n2068), .dinb(n2067), .dout(n2069));
  jand g1807(.dina(n1378), .dinb(n295), .dout(n2070));
  jand g1808(.dina(n1415), .dinb(n308), .dout(n2071));
  jor  g1809(.dina(n2071), .dinb(n2070), .dout(n2072));
  jor  g1810(.dina(n2072), .dinb(n2069), .dout(n2073));
  jand g1811(.dina(n2073), .dinb(n432), .dout(n2074));
  jand g1812(.dina(n1521), .dinb(n266), .dout(n2075));
  jand g1813(.dina(n1426), .dinb(n281), .dout(n2076));
  jor  g1814(.dina(n2076), .dinb(n2075), .dout(n2077));
  jand g1815(.dina(n1530), .dinb(n295), .dout(n2078));
  jand g1816(.dina(n1435), .dinb(n308), .dout(n2079));
  jor  g1817(.dina(n2079), .dinb(n2078), .dout(n2080));
  jor  g1818(.dina(n2080), .dinb(n2077), .dout(n2081));
  jand g1819(.dina(n2081), .dinb(n485), .dout(n2082));
  jor  g1820(.dina(n2082), .dinb(n2074), .dout(n2083));
  jor  g1821(.dina(n2083), .dinb(n2066), .dout(n2084));
  jand g1822(.dina(n2084), .dinb(n263), .dout(n2085));
  jand g1823(.dina(n1453), .dinb(n266), .dout(n2086));
  jand g1824(.dina(n1462), .dinb(n295), .dout(n2087));
  jor  g1825(.dina(n2087), .dinb(n2086), .dout(n2088));
  jand g1826(.dina(n1490), .dinb(n281), .dout(n2089));
  jand g1827(.dina(n1505), .dinb(n308), .dout(n2090));
  jor  g1828(.dina(n2090), .dinb(n2089), .dout(n2091));
  jor  g1829(.dina(n2091), .dinb(n2088), .dout(n2092));
  jand g1830(.dina(n2092), .dinb(n377), .dout(n2093));
  jand g1831(.dina(n1473), .dinb(n266), .dout(n2094));
  jand g1832(.dina(n1517), .dinb(n281), .dout(n2095));
  jor  g1833(.dina(n2095), .dinb(n2094), .dout(n2096));
  jand g1834(.dina(n1482), .dinb(n295), .dout(n2097));
  jand g1835(.dina(n1526), .dinb(n308), .dout(n2098));
  jor  g1836(.dina(n2098), .dinb(n2097), .dout(n2099));
  jor  g1837(.dina(n2099), .dinb(n2096), .dout(n2100));
  jand g1838(.dina(n2100), .dinb(n323), .dout(n2101));
  jor  g1839(.dina(n2101), .dinb(n2093), .dout(n2102));
  jand g1840(.dina(n1389), .dinb(n266), .dout(n2103));
  jand g1841(.dina(n1449), .dinb(n281), .dout(n2104));
  jor  g1842(.dina(n2104), .dinb(n2103), .dout(n2105));
  jand g1843(.dina(n1398), .dinb(n295), .dout(n2106));
  jand g1844(.dina(n1458), .dinb(n308), .dout(n2107));
  jor  g1845(.dina(n2107), .dinb(n2106), .dout(n2108));
  jor  g1846(.dina(n2108), .dinb(n2105), .dout(n2109));
  jand g1847(.dina(n2109), .dinb(n485), .dout(n2110));
  jand g1848(.dina(n1496), .dinb(n266), .dout(n2111));
  jand g1849(.dina(n1469), .dinb(n281), .dout(n2112));
  jor  g1850(.dina(n2112), .dinb(n2111), .dout(n2113));
  jand g1851(.dina(n1510), .dinb(n295), .dout(n2114));
  jand g1852(.dina(n1478), .dinb(n308), .dout(n2115));
  jor  g1853(.dina(n2115), .dinb(n2114), .dout(n2116));
  jor  g1854(.dina(n2116), .dinb(n2113), .dout(n2117));
  jand g1855(.dina(n2117), .dinb(n432), .dout(n2118));
  jor  g1856(.dina(n2118), .dinb(n2110), .dout(n2119));
  jor  g1857(.dina(n2119), .dinb(n2102), .dout(n2120));
  jand g1858(.dina(n2120), .dinb(shift6 ), .dout(n2121));
  jor  g1859(.dina(n2121), .dinb(n2085), .dout(result11 ));
  jand g1860(.dina(n415), .dinb(n266), .dout(n2123));
  jand g1861(.dina(n427), .dinb(n281), .dout(n2124));
  jor  g1862(.dina(n2124), .dinb(n2123), .dout(n2125));
  jand g1863(.dina(n402), .dinb(n295), .dout(n2126));
  jand g1864(.dina(n308), .dinb(n279), .dout(n2127));
  jor  g1865(.dina(n2127), .dinb(n2126), .dout(n2128));
  jor  g1866(.dina(n2128), .dinb(n2125), .dout(n2129));
  jand g1867(.dina(n2129), .dinb(n323), .dout(n2130));
  jand g1868(.dina(n469), .dinb(n266), .dout(n2131));
  jand g1869(.dina(n481), .dinb(n281), .dout(n2132));
  jor  g1870(.dina(n2132), .dinb(n2131), .dout(n2133));
  jand g1871(.dina(n456), .dinb(n295), .dout(n2134));
  jand g1872(.dina(n335), .dinb(n308), .dout(n2135));
  jor  g1873(.dina(n2135), .dinb(n2134), .dout(n2136));
  jor  g1874(.dina(n2136), .dinb(n2133), .dout(n2137));
  jand g1875(.dina(n2137), .dinb(n377), .dout(n2138));
  jor  g1876(.dina(n2138), .dinb(n2130), .dout(n2139));
  jand g1877(.dina(n360), .dinb(n266), .dout(n2140));
  jand g1878(.dina(n372), .dinb(n281), .dout(n2141));
  jor  g1879(.dina(n2141), .dinb(n2140), .dout(n2142));
  jand g1880(.dina(n347), .dinb(n295), .dout(n2143));
  jand g1881(.dina(n390), .dinb(n308), .dout(n2144));
  jor  g1882(.dina(n2144), .dinb(n2143), .dout(n2145));
  jor  g1883(.dina(n2145), .dinb(n2142), .dout(n2146));
  jand g1884(.dina(n2146), .dinb(n432), .dout(n2147));
  jand g1885(.dina(n525), .dinb(n266), .dout(n2148));
  jand g1886(.dina(n537), .dinb(n281), .dout(n2149));
  jor  g1887(.dina(n2149), .dinb(n2148), .dout(n2150));
  jand g1888(.dina(n512), .dinb(n295), .dout(n2151));
  jand g1889(.dina(n444), .dinb(n308), .dout(n2152));
  jor  g1890(.dina(n2152), .dinb(n2151), .dout(n2153));
  jor  g1891(.dina(n2153), .dinb(n2150), .dout(n2154));
  jand g1892(.dina(n2154), .dinb(n485), .dout(n2155));
  jor  g1893(.dina(n2155), .dinb(n2147), .dout(n2156));
  jor  g1894(.dina(n2156), .dinb(n2139), .dout(n2157));
  jand g1895(.dina(n2157), .dinb(n263), .dout(n2158));
  jand g1896(.dina(n680), .dinb(n266), .dout(n2159));
  jand g1897(.dina(n692), .dinb(n281), .dout(n2160));
  jor  g1898(.dina(n2160), .dinb(n2159), .dout(n2161));
  jand g1899(.dina(n667), .dinb(n295), .dout(n2162));
  jand g1900(.dina(n552), .dinb(n308), .dout(n2163));
  jor  g1901(.dina(n2163), .dinb(n2162), .dout(n2164));
  jor  g1902(.dina(n2164), .dinb(n2161), .dout(n2165));
  jand g1903(.dina(n2165), .dinb(n377), .dout(n2166));
  jand g1904(.dina(n628), .dinb(n266), .dout(n2167));
  jand g1905(.dina(n640), .dinb(n281), .dout(n2168));
  jor  g1906(.dina(n2168), .dinb(n2167), .dout(n2169));
  jand g1907(.dina(n615), .dinb(n295), .dout(n2170));
  jand g1908(.dina(n500), .dinb(n308), .dout(n2171));
  jor  g1909(.dina(n2171), .dinb(n2170), .dout(n2172));
  jor  g1910(.dina(n2172), .dinb(n2169), .dout(n2173));
  jand g1911(.dina(n2173), .dinb(n323), .dout(n2174));
  jor  g1912(.dina(n2174), .dinb(n2166), .dout(n2175));
  jand g1913(.dina(n306), .dinb(n266), .dout(n2176));
  jand g1914(.dina(n319), .dinb(n281), .dout(n2177));
  jor  g1915(.dina(n2177), .dinb(n2176), .dout(n2178));
  jand g1916(.dina(n295), .dinb(n292), .dout(n2179));
  jand g1917(.dina(n655), .dinb(n308), .dout(n2180));
  jor  g1918(.dina(n2180), .dinb(n2179), .dout(n2181));
  jor  g1919(.dina(n2181), .dinb(n2178), .dout(n2182));
  jand g1920(.dina(n2182), .dinb(n485), .dout(n2183));
  jand g1921(.dina(n575), .dinb(n266), .dout(n2184));
  jand g1922(.dina(n587), .dinb(n281), .dout(n2185));
  jor  g1923(.dina(n2185), .dinb(n2184), .dout(n2186));
  jand g1924(.dina(n562), .dinb(n295), .dout(n2187));
  jand g1925(.dina(n603), .dinb(n308), .dout(n2188));
  jor  g1926(.dina(n2188), .dinb(n2187), .dout(n2189));
  jor  g1927(.dina(n2189), .dinb(n2186), .dout(n2190));
  jand g1928(.dina(n2190), .dinb(n432), .dout(n2191));
  jor  g1929(.dina(n2191), .dinb(n2183), .dout(n2192));
  jor  g1930(.dina(n2192), .dinb(n2175), .dout(n2193));
  jand g1931(.dina(n2193), .dinb(shift6 ), .dout(n2194));
  jor  g1932(.dina(n2194), .dinb(n2158), .dout(result12 ));
  jand g1933(.dina(n819), .dinb(n266), .dout(n2196));
  jand g1934(.dina(n829), .dinb(n281), .dout(n2197));
  jor  g1935(.dina(n2197), .dinb(n2196), .dout(n2198));
  jand g1936(.dina(n808), .dinb(n295), .dout(n2199));
  jand g1937(.dina(n709), .dinb(n308), .dout(n2200));
  jor  g1938(.dina(n2200), .dinb(n2199), .dout(n2201));
  jor  g1939(.dina(n2201), .dinb(n2198), .dout(n2202));
  jand g1940(.dina(n2202), .dinb(n323), .dout(n2203));
  jand g1941(.dina(n863), .dinb(n266), .dout(n2204));
  jand g1942(.dina(n873), .dinb(n281), .dout(n2205));
  jor  g1943(.dina(n2205), .dinb(n2204), .dout(n2206));
  jand g1944(.dina(n852), .dinb(n295), .dout(n2207));
  jand g1945(.dina(n753), .dinb(n308), .dout(n2208));
  jor  g1946(.dina(n2208), .dinb(n2207), .dout(n2209));
  jor  g1947(.dina(n2209), .dinb(n2206), .dout(n2210));
  jand g1948(.dina(n2210), .dinb(n377), .dout(n2211));
  jor  g1949(.dina(n2211), .dinb(n2203), .dout(n2212));
  jand g1950(.dina(n774), .dinb(n266), .dout(n2213));
  jand g1951(.dina(n784), .dinb(n281), .dout(n2214));
  jor  g1952(.dina(n2214), .dinb(n2213), .dout(n2215));
  jand g1953(.dina(n763), .dinb(n295), .dout(n2216));
  jand g1954(.dina(n798), .dinb(n308), .dout(n2217));
  jor  g1955(.dina(n2217), .dinb(n2216), .dout(n2218));
  jor  g1956(.dina(n2218), .dinb(n2215), .dout(n2219));
  jand g1957(.dina(n2219), .dinb(n432), .dout(n2220));
  jand g1958(.dina(n999), .dinb(n266), .dout(n2221));
  jand g1959(.dina(n1009), .dinb(n281), .dout(n2222));
  jor  g1960(.dina(n2222), .dinb(n2221), .dout(n2223));
  jand g1961(.dina(n988), .dinb(n295), .dout(n2224));
  jand g1962(.dina(n842), .dinb(n308), .dout(n2225));
  jor  g1963(.dina(n2225), .dinb(n2224), .dout(n2226));
  jor  g1964(.dina(n2226), .dinb(n2223), .dout(n2227));
  jand g1965(.dina(n2227), .dinb(n485), .dout(n2228));
  jor  g1966(.dina(n2228), .dinb(n2220), .dout(n2229));
  jor  g1967(.dina(n2229), .dinb(n2212), .dout(n2230));
  jand g1968(.dina(n2230), .dinb(n263), .dout(n2231));
  jand g1969(.dina(n910), .dinb(n266), .dout(n2232));
  jand g1970(.dina(n920), .dinb(n281), .dout(n2233));
  jor  g1971(.dina(n2233), .dinb(n2232), .dout(n2234));
  jand g1972(.dina(n899), .dinb(n295), .dout(n2235));
  jand g1973(.dina(n1022), .dinb(n308), .dout(n2236));
  jor  g1974(.dina(n2236), .dinb(n2235), .dout(n2237));
  jor  g1975(.dina(n2237), .dinb(n2234), .dout(n2238));
  jand g1976(.dina(n2238), .dinb(n377), .dout(n2239));
  jand g1977(.dina(n954), .dinb(n266), .dout(n2240));
  jand g1978(.dina(n964), .dinb(n281), .dout(n2241));
  jor  g1979(.dina(n2241), .dinb(n2240), .dout(n2242));
  jand g1980(.dina(n943), .dinb(n295), .dout(n2243));
  jand g1981(.dina(n978), .dinb(n308), .dout(n2244));
  jor  g1982(.dina(n2244), .dinb(n2243), .dout(n2245));
  jor  g1983(.dina(n2245), .dinb(n2242), .dout(n2246));
  jand g1984(.dina(n2246), .dinb(n323), .dout(n2247));
  jor  g1985(.dina(n2247), .dinb(n2239), .dout(n2248));
  jand g1986(.dina(n730), .dinb(n266), .dout(n2249));
  jand g1987(.dina(n740), .dinb(n281), .dout(n2250));
  jor  g1988(.dina(n2250), .dinb(n2249), .dout(n2251));
  jand g1989(.dina(n719), .dinb(n295), .dout(n2252));
  jand g1990(.dina(n889), .dinb(n308), .dout(n2253));
  jor  g1991(.dina(n2253), .dinb(n2252), .dout(n2254));
  jor  g1992(.dina(n2254), .dinb(n2251), .dout(n2255));
  jand g1993(.dina(n2255), .dinb(n485), .dout(n2256));
  jand g1994(.dina(n1047), .dinb(n266), .dout(n2257));
  jand g1995(.dina(n1057), .dinb(n281), .dout(n2258));
  jor  g1996(.dina(n2258), .dinb(n2257), .dout(n2259));
  jand g1997(.dina(n1034), .dinb(n295), .dout(n2260));
  jand g1998(.dina(n933), .dinb(n308), .dout(n2261));
  jor  g1999(.dina(n2261), .dinb(n2260), .dout(n2262));
  jor  g2000(.dina(n2262), .dinb(n2259), .dout(n2263));
  jand g2001(.dina(n2263), .dinb(n432), .dout(n2264));
  jor  g2002(.dina(n2264), .dinb(n2256), .dout(n2265));
  jor  g2003(.dina(n2265), .dinb(n2248), .dout(n2266));
  jand g2004(.dina(n2266), .dinb(shift6 ), .dout(n2267));
  jor  g2005(.dina(n2267), .dinb(n2231), .dout(result13 ));
  jand g2006(.dina(n1162), .dinb(n266), .dout(n2269));
  jand g2007(.dina(n1170), .dinb(n281), .dout(n2270));
  jor  g2008(.dina(n2270), .dinb(n2269), .dout(n2271));
  jand g2009(.dina(n1153), .dinb(n295), .dout(n2272));
  jand g2010(.dina(n1072), .dinb(n308), .dout(n2273));
  jor  g2011(.dina(n2273), .dinb(n2272), .dout(n2274));
  jor  g2012(.dina(n2274), .dinb(n2271), .dout(n2275));
  jand g2013(.dina(n2275), .dinb(n323), .dout(n2276));
  jand g2014(.dina(n1198), .dinb(n266), .dout(n2277));
  jand g2015(.dina(n1206), .dinb(n281), .dout(n2278));
  jor  g2016(.dina(n2278), .dinb(n2277), .dout(n2279));
  jand g2017(.dina(n1189), .dinb(n295), .dout(n2280));
  jand g2018(.dina(n1108), .dinb(n308), .dout(n2281));
  jor  g2019(.dina(n2281), .dinb(n2280), .dout(n2282));
  jor  g2020(.dina(n2282), .dinb(n2279), .dout(n2283));
  jand g2021(.dina(n2283), .dinb(n377), .dout(n2284));
  jor  g2022(.dina(n2284), .dinb(n2276), .dout(n2285));
  jand g2023(.dina(n1125), .dinb(n266), .dout(n2286));
  jand g2024(.dina(n1133), .dinb(n281), .dout(n2287));
  jor  g2025(.dina(n2287), .dinb(n2286), .dout(n2288));
  jand g2026(.dina(n1116), .dinb(n295), .dout(n2289));
  jand g2027(.dina(n1145), .dinb(n308), .dout(n2290));
  jor  g2028(.dina(n2290), .dinb(n2289), .dout(n2291));
  jor  g2029(.dina(n2291), .dinb(n2288), .dout(n2292));
  jand g2030(.dina(n2292), .dinb(n432), .dout(n2293));
  jand g2031(.dina(n1310), .dinb(n266), .dout(n2294));
  jand g2032(.dina(n1318), .dinb(n281), .dout(n2295));
  jor  g2033(.dina(n2295), .dinb(n2294), .dout(n2296));
  jand g2034(.dina(n1301), .dinb(n295), .dout(n2297));
  jand g2035(.dina(n1181), .dinb(n308), .dout(n2298));
  jor  g2036(.dina(n2298), .dinb(n2297), .dout(n2299));
  jor  g2037(.dina(n2299), .dinb(n2296), .dout(n2300));
  jand g2038(.dina(n2300), .dinb(n485), .dout(n2301));
  jor  g2039(.dina(n2301), .dinb(n2293), .dout(n2302));
  jor  g2040(.dina(n2302), .dinb(n2285), .dout(n2303));
  jand g2041(.dina(n2303), .dinb(n263), .dout(n2304));
  jand g2042(.dina(n1237), .dinb(n266), .dout(n2305));
  jand g2043(.dina(n1245), .dinb(n281), .dout(n2306));
  jor  g2044(.dina(n2306), .dinb(n2305), .dout(n2307));
  jand g2045(.dina(n1228), .dinb(n295), .dout(n2308));
  jand g2046(.dina(n1329), .dinb(n308), .dout(n2309));
  jor  g2047(.dina(n2309), .dinb(n2308), .dout(n2310));
  jor  g2048(.dina(n2310), .dinb(n2307), .dout(n2311));
  jand g2049(.dina(n2311), .dinb(n377), .dout(n2312));
  jand g2050(.dina(n1273), .dinb(n266), .dout(n2313));
  jand g2051(.dina(n1281), .dinb(n281), .dout(n2314));
  jor  g2052(.dina(n2314), .dinb(n2313), .dout(n2315));
  jand g2053(.dina(n1264), .dinb(n295), .dout(n2316));
  jand g2054(.dina(n1293), .dinb(n308), .dout(n2317));
  jor  g2055(.dina(n2317), .dinb(n2316), .dout(n2318));
  jor  g2056(.dina(n2318), .dinb(n2315), .dout(n2319));
  jand g2057(.dina(n2319), .dinb(n323), .dout(n2320));
  jor  g2058(.dina(n2320), .dinb(n2312), .dout(n2321));
  jand g2059(.dina(n1089), .dinb(n266), .dout(n2322));
  jand g2060(.dina(n1097), .dinb(n281), .dout(n2323));
  jor  g2061(.dina(n2323), .dinb(n2322), .dout(n2324));
  jand g2062(.dina(n1080), .dinb(n295), .dout(n2325));
  jand g2063(.dina(n1220), .dinb(n308), .dout(n2326));
  jor  g2064(.dina(n2326), .dinb(n2325), .dout(n2327));
  jor  g2065(.dina(n2327), .dinb(n2324), .dout(n2328));
  jand g2066(.dina(n2328), .dinb(n485), .dout(n2329));
  jand g2067(.dina(n1346), .dinb(n266), .dout(n2330));
  jand g2068(.dina(n1354), .dinb(n281), .dout(n2331));
  jor  g2069(.dina(n2331), .dinb(n2330), .dout(n2332));
  jand g2070(.dina(n1337), .dinb(n295), .dout(n2333));
  jand g2071(.dina(n1256), .dinb(n308), .dout(n2334));
  jor  g2072(.dina(n2334), .dinb(n2333), .dout(n2335));
  jor  g2073(.dina(n2335), .dinb(n2332), .dout(n2336));
  jand g2074(.dina(n2336), .dinb(n432), .dout(n2337));
  jor  g2075(.dina(n2337), .dinb(n2329), .dout(n2338));
  jor  g2076(.dina(n2338), .dinb(n2321), .dout(n2339));
  jand g2077(.dina(n2339), .dinb(shift6 ), .dout(n2340));
  jor  g2078(.dina(n2340), .dinb(n2304), .dout(result14 ));
  jand g2079(.dina(n1415), .dinb(n266), .dout(n2342));
  jand g2080(.dina(n1419), .dinb(n281), .dout(n2343));
  jor  g2081(.dina(n2343), .dinb(n2342), .dout(n2344));
  jand g2082(.dina(n1410), .dinb(n295), .dout(n2345));
  jand g2083(.dina(n1385), .dinb(n308), .dout(n2346));
  jor  g2084(.dina(n2346), .dinb(n2345), .dout(n2347));
  jor  g2085(.dina(n2347), .dinb(n2344), .dout(n2348));
  jand g2086(.dina(n2348), .dinb(n323), .dout(n2349));
  jand g2087(.dina(n1435), .dinb(n266), .dout(n2350));
  jand g2088(.dina(n1439), .dinb(n281), .dout(n2351));
  jor  g2089(.dina(n2351), .dinb(n2350), .dout(n2352));
  jand g2090(.dina(n1430), .dinb(n295), .dout(n2353));
  jand g2091(.dina(n1365), .dinb(n308), .dout(n2354));
  jor  g2092(.dina(n2354), .dinb(n2353), .dout(n2355));
  jor  g2093(.dina(n2355), .dinb(n2352), .dout(n2356));
  jand g2094(.dina(n2356), .dinb(n377), .dout(n2357));
  jor  g2095(.dina(n2357), .dinb(n2349), .dout(n2358));
  jand g2096(.dina(n1374), .dinb(n266), .dout(n2359));
  jand g2097(.dina(n1378), .dinb(n281), .dout(n2360));
  jor  g2098(.dina(n2360), .dinb(n2359), .dout(n2361));
  jand g2099(.dina(n1369), .dinb(n295), .dout(n2362));
  jand g2100(.dina(n1406), .dinb(n308), .dout(n2363));
  jor  g2101(.dina(n2363), .dinb(n2362), .dout(n2364));
  jor  g2102(.dina(n2364), .dinb(n2361), .dout(n2365));
  jand g2103(.dina(n2365), .dinb(n432), .dout(n2366));
  jand g2104(.dina(n1526), .dinb(n266), .dout(n2367));
  jand g2105(.dina(n1530), .dinb(n281), .dout(n2368));
  jor  g2106(.dina(n2368), .dinb(n2367), .dout(n2369));
  jand g2107(.dina(n1521), .dinb(n295), .dout(n2370));
  jand g2108(.dina(n1426), .dinb(n308), .dout(n2371));
  jor  g2109(.dina(n2371), .dinb(n2370), .dout(n2372));
  jor  g2110(.dina(n2372), .dinb(n2369), .dout(n2373));
  jand g2111(.dina(n2373), .dinb(n485), .dout(n2374));
  jor  g2112(.dina(n2374), .dinb(n2366), .dout(n2375));
  jor  g2113(.dina(n2375), .dinb(n2358), .dout(n2376));
  jand g2114(.dina(n2376), .dinb(n263), .dout(n2377));
  jand g2115(.dina(n1458), .dinb(n266), .dout(n2378));
  jand g2116(.dina(n1462), .dinb(n281), .dout(n2379));
  jor  g2117(.dina(n2379), .dinb(n2378), .dout(n2380));
  jand g2118(.dina(n1453), .dinb(n295), .dout(n2381));
  jand g2119(.dina(n1490), .dinb(n308), .dout(n2382));
  jor  g2120(.dina(n2382), .dinb(n2381), .dout(n2383));
  jor  g2121(.dina(n2383), .dinb(n2380), .dout(n2384));
  jand g2122(.dina(n2384), .dinb(n377), .dout(n2385));
  jand g2123(.dina(n1478), .dinb(n266), .dout(n2386));
  jand g2124(.dina(n1482), .dinb(n281), .dout(n2387));
  jor  g2125(.dina(n2387), .dinb(n2386), .dout(n2388));
  jand g2126(.dina(n1473), .dinb(n295), .dout(n2389));
  jand g2127(.dina(n1517), .dinb(n308), .dout(n2390));
  jor  g2128(.dina(n2390), .dinb(n2389), .dout(n2391));
  jor  g2129(.dina(n2391), .dinb(n2388), .dout(n2392));
  jand g2130(.dina(n2392), .dinb(n323), .dout(n2393));
  jor  g2131(.dina(n2393), .dinb(n2385), .dout(n2394));
  jand g2132(.dina(n1394), .dinb(n266), .dout(n2395));
  jand g2133(.dina(n1398), .dinb(n281), .dout(n2396));
  jor  g2134(.dina(n2396), .dinb(n2395), .dout(n2397));
  jand g2135(.dina(n1389), .dinb(n295), .dout(n2398));
  jand g2136(.dina(n1449), .dinb(n308), .dout(n2399));
  jor  g2137(.dina(n2399), .dinb(n2398), .dout(n2400));
  jor  g2138(.dina(n2400), .dinb(n2397), .dout(n2401));
  jand g2139(.dina(n2401), .dinb(n485), .dout(n2402));
  jand g2140(.dina(n1505), .dinb(n266), .dout(n2403));
  jand g2141(.dina(n1510), .dinb(n281), .dout(n2404));
  jor  g2142(.dina(n2404), .dinb(n2403), .dout(n2405));
  jand g2143(.dina(n1496), .dinb(n295), .dout(n2406));
  jand g2144(.dina(n1469), .dinb(n308), .dout(n2407));
  jor  g2145(.dina(n2407), .dinb(n2406), .dout(n2408));
  jor  g2146(.dina(n2408), .dinb(n2405), .dout(n2409));
  jand g2147(.dina(n2409), .dinb(n432), .dout(n2410));
  jor  g2148(.dina(n2410), .dinb(n2402), .dout(n2411));
  jor  g2149(.dina(n2411), .dinb(n2394), .dout(n2412));
  jand g2150(.dina(n2412), .dinb(shift6 ), .dout(n2413));
  jor  g2151(.dina(n2413), .dinb(n2377), .dout(result15 ));
  jand g2152(.dina(n430), .dinb(n323), .dout(n2415));
  jand g2153(.dina(n484), .dinb(n377), .dout(n2416));
  jor  g2154(.dina(n2416), .dinb(n2415), .dout(n2417));
  jand g2155(.dina(n432), .dinb(n375), .dout(n2418));
  jand g2156(.dina(n540), .dinb(n485), .dout(n2419));
  jor  g2157(.dina(n2419), .dinb(n2418), .dout(n2420));
  jor  g2158(.dina(n2420), .dinb(n2417), .dout(n2421));
  jand g2159(.dina(n2421), .dinb(n263), .dout(n2422));
  jand g2160(.dina(n485), .dinb(n322), .dout(n2423));
  jand g2161(.dina(n590), .dinb(n432), .dout(n2424));
  jor  g2162(.dina(n2424), .dinb(n2423), .dout(n2425));
  jand g2163(.dina(n643), .dinb(n323), .dout(n2426));
  jand g2164(.dina(n695), .dinb(n377), .dout(n2427));
  jor  g2165(.dina(n2427), .dinb(n2426), .dout(n2428));
  jor  g2166(.dina(n2428), .dinb(n2425), .dout(n2429));
  jand g2167(.dina(n2429), .dinb(shift6 ), .dout(n2430));
  jor  g2168(.dina(n2430), .dinb(n2422), .dout(result16 ));
  jand g2169(.dina(n832), .dinb(n323), .dout(n2432));
  jand g2170(.dina(n876), .dinb(n377), .dout(n2433));
  jor  g2171(.dina(n2433), .dinb(n2432), .dout(n2434));
  jand g2172(.dina(n787), .dinb(n432), .dout(n2435));
  jand g2173(.dina(n1012), .dinb(n485), .dout(n2436));
  jor  g2174(.dina(n2436), .dinb(n2435), .dout(n2437));
  jor  g2175(.dina(n2437), .dinb(n2434), .dout(n2438));
  jand g2176(.dina(n2438), .dinb(n263), .dout(n2439));
  jand g2177(.dina(n923), .dinb(n377), .dout(n2440));
  jand g2178(.dina(n967), .dinb(n323), .dout(n2441));
  jor  g2179(.dina(n2441), .dinb(n2440), .dout(n2442));
  jand g2180(.dina(n743), .dinb(n485), .dout(n2443));
  jand g2181(.dina(n1060), .dinb(n432), .dout(n2444));
  jor  g2182(.dina(n2444), .dinb(n2443), .dout(n2445));
  jor  g2183(.dina(n2445), .dinb(n2442), .dout(n2446));
  jand g2184(.dina(n2446), .dinb(shift6 ), .dout(n2447));
  jor  g2185(.dina(n2447), .dinb(n2439), .dout(result17 ));
  jand g2186(.dina(n1173), .dinb(n323), .dout(n2449));
  jand g2187(.dina(n1209), .dinb(n377), .dout(n2450));
  jor  g2188(.dina(n2450), .dinb(n2449), .dout(n2451));
  jand g2189(.dina(n1136), .dinb(n432), .dout(n2452));
  jand g2190(.dina(n1321), .dinb(n485), .dout(n2453));
  jor  g2191(.dina(n2453), .dinb(n2452), .dout(n2454));
  jor  g2192(.dina(n2454), .dinb(n2451), .dout(n2455));
  jand g2193(.dina(n2455), .dinb(n263), .dout(n2456));
  jand g2194(.dina(n1248), .dinb(n377), .dout(n2457));
  jand g2195(.dina(n1284), .dinb(n323), .dout(n2458));
  jor  g2196(.dina(n2458), .dinb(n2457), .dout(n2459));
  jand g2197(.dina(n1100), .dinb(n485), .dout(n2460));
  jand g2198(.dina(n1357), .dinb(n432), .dout(n2461));
  jor  g2199(.dina(n2461), .dinb(n2460), .dout(n2462));
  jor  g2200(.dina(n2462), .dinb(n2459), .dout(n2463));
  jand g2201(.dina(n2463), .dinb(shift6 ), .dout(n2464));
  jor  g2202(.dina(n2464), .dinb(n2456), .dout(result18 ));
  jand g2203(.dina(n1381), .dinb(n432), .dout(n2466));
  jand g2204(.dina(n1533), .dinb(n485), .dout(n2467));
  jor  g2205(.dina(n2467), .dinb(n2466), .dout(n2468));
  jand g2206(.dina(n1422), .dinb(n323), .dout(n2469));
  jand g2207(.dina(n1442), .dinb(n377), .dout(n2470));
  jor  g2208(.dina(n2470), .dinb(n2469), .dout(n2471));
  jor  g2209(.dina(n2471), .dinb(n2468), .dout(n2472));
  jand g2210(.dina(n2472), .dinb(n263), .dout(n2473));
  jand g2211(.dina(n1465), .dinb(n377), .dout(n2474));
  jand g2212(.dina(n1513), .dinb(n432), .dout(n2475));
  jor  g2213(.dina(n2475), .dinb(n2474), .dout(n2476));
  jand g2214(.dina(n1401), .dinb(n485), .dout(n2477));
  jand g2215(.dina(n1485), .dinb(n323), .dout(n2478));
  jor  g2216(.dina(n2478), .dinb(n2477), .dout(n2479));
  jor  g2217(.dina(n2479), .dinb(n2476), .dout(n2480));
  jand g2218(.dina(n2480), .dinb(shift6 ), .dout(n2481));
  jor  g2219(.dina(n2481), .dinb(n2473), .dout(result19 ));
  jand g2220(.dina(n1562), .dinb(n323), .dout(n2483));
  jand g2221(.dina(n1570), .dinb(n377), .dout(n2484));
  jor  g2222(.dina(n2484), .dinb(n2483), .dout(n2485));
  jand g2223(.dina(n1553), .dinb(n432), .dout(n2486));
  jand g2224(.dina(n1589), .dinb(n485), .dout(n2487));
  jor  g2225(.dina(n2487), .dinb(n2486), .dout(n2488));
  jor  g2226(.dina(n2488), .dinb(n2485), .dout(n2489));
  jand g2227(.dina(n2489), .dinb(n263), .dout(n2490));
  jand g2228(.dina(n1545), .dinb(n485), .dout(n2491));
  jand g2229(.dina(n1598), .dinb(n377), .dout(n2492));
  jor  g2230(.dina(n2492), .dinb(n2491), .dout(n2493));
  jand g2231(.dina(n1581), .dinb(n432), .dout(n2494));
  jand g2232(.dina(n1606), .dinb(n323), .dout(n2495));
  jor  g2233(.dina(n2495), .dinb(n2494), .dout(n2496));
  jor  g2234(.dina(n2496), .dinb(n2493), .dout(n2497));
  jand g2235(.dina(n2497), .dinb(shift6 ), .dout(n2498));
  jor  g2236(.dina(n2498), .dinb(n2490), .dout(result20 ));
  jand g2237(.dina(n1635), .dinb(n323), .dout(n2500));
  jand g2238(.dina(n1643), .dinb(n377), .dout(n2501));
  jor  g2239(.dina(n2501), .dinb(n2500), .dout(n2502));
  jand g2240(.dina(n1626), .dinb(n432), .dout(n2503));
  jand g2241(.dina(n1662), .dinb(n485), .dout(n2504));
  jor  g2242(.dina(n2504), .dinb(n2503), .dout(n2505));
  jor  g2243(.dina(n2505), .dinb(n2502), .dout(n2506));
  jand g2244(.dina(n2506), .dinb(n263), .dout(n2507));
  jand g2245(.dina(n1618), .dinb(n485), .dout(n2508));
  jand g2246(.dina(n1671), .dinb(n377), .dout(n2509));
  jor  g2247(.dina(n2509), .dinb(n2508), .dout(n2510));
  jand g2248(.dina(n1654), .dinb(n432), .dout(n2511));
  jand g2249(.dina(n1679), .dinb(n323), .dout(n2512));
  jor  g2250(.dina(n2512), .dinb(n2511), .dout(n2513));
  jor  g2251(.dina(n2513), .dinb(n2510), .dout(n2514));
  jand g2252(.dina(n2514), .dinb(shift6 ), .dout(n2515));
  jor  g2253(.dina(n2515), .dinb(n2507), .dout(result21 ));
  jand g2254(.dina(n1708), .dinb(n323), .dout(n2517));
  jand g2255(.dina(n1716), .dinb(n377), .dout(n2518));
  jor  g2256(.dina(n2518), .dinb(n2517), .dout(n2519));
  jand g2257(.dina(n1699), .dinb(n432), .dout(n2520));
  jand g2258(.dina(n1735), .dinb(n485), .dout(n2521));
  jor  g2259(.dina(n2521), .dinb(n2520), .dout(n2522));
  jor  g2260(.dina(n2522), .dinb(n2519), .dout(n2523));
  jand g2261(.dina(n2523), .dinb(n263), .dout(n2524));
  jand g2262(.dina(n1691), .dinb(n485), .dout(n2525));
  jand g2263(.dina(n1744), .dinb(n377), .dout(n2526));
  jor  g2264(.dina(n2526), .dinb(n2525), .dout(n2527));
  jand g2265(.dina(n1727), .dinb(n432), .dout(n2528));
  jand g2266(.dina(n1752), .dinb(n323), .dout(n2529));
  jor  g2267(.dina(n2529), .dinb(n2528), .dout(n2530));
  jor  g2268(.dina(n2530), .dinb(n2527), .dout(n2531));
  jand g2269(.dina(n2531), .dinb(shift6 ), .dout(n2532));
  jor  g2270(.dina(n2532), .dinb(n2524), .dout(result22 ));
  jand g2271(.dina(n1781), .dinb(n323), .dout(n2534));
  jand g2272(.dina(n1772), .dinb(n432), .dout(n2535));
  jor  g2273(.dina(n2535), .dinb(n2534), .dout(n2536));
  jand g2274(.dina(n1808), .dinb(n485), .dout(n2537));
  jand g2275(.dina(n1789), .dinb(n377), .dout(n2538));
  jor  g2276(.dina(n2538), .dinb(n2537), .dout(n2539));
  jor  g2277(.dina(n2539), .dinb(n2536), .dout(n2540));
  jand g2278(.dina(n2540), .dinb(n263), .dout(n2541));
  jand g2279(.dina(n1800), .dinb(n432), .dout(n2542));
  jand g2280(.dina(n1764), .dinb(n485), .dout(n2543));
  jor  g2281(.dina(n2543), .dinb(n2542), .dout(n2544));
  jand g2282(.dina(n1817), .dinb(n377), .dout(n2545));
  jand g2283(.dina(n1825), .dinb(n323), .dout(n2546));
  jor  g2284(.dina(n2546), .dinb(n2545), .dout(n2547));
  jor  g2285(.dina(n2547), .dinb(n2544), .dout(n2548));
  jand g2286(.dina(n2548), .dinb(shift6 ), .dout(n2549));
  jor  g2287(.dina(n2549), .dinb(n2541), .dout(result23 ));
  jand g2288(.dina(n1854), .dinb(n323), .dout(n2551));
  jand g2289(.dina(n1845), .dinb(n432), .dout(n2552));
  jor  g2290(.dina(n2552), .dinb(n2551), .dout(n2553));
  jand g2291(.dina(n1881), .dinb(n485), .dout(n2554));
  jand g2292(.dina(n1862), .dinb(n377), .dout(n2555));
  jor  g2293(.dina(n2555), .dinb(n2554), .dout(n2556));
  jor  g2294(.dina(n2556), .dinb(n2553), .dout(n2557));
  jand g2295(.dina(n2557), .dinb(n263), .dout(n2558));
  jand g2296(.dina(n1873), .dinb(n432), .dout(n2559));
  jand g2297(.dina(n1837), .dinb(n485), .dout(n2560));
  jor  g2298(.dina(n2560), .dinb(n2559), .dout(n2561));
  jand g2299(.dina(n1890), .dinb(n377), .dout(n2562));
  jand g2300(.dina(n1898), .dinb(n323), .dout(n2563));
  jor  g2301(.dina(n2563), .dinb(n2562), .dout(n2564));
  jor  g2302(.dina(n2564), .dinb(n2561), .dout(n2565));
  jand g2303(.dina(n2565), .dinb(shift6 ), .dout(n2566));
  jor  g2304(.dina(n2566), .dinb(n2558), .dout(result24 ));
  jand g2305(.dina(n1927), .dinb(n323), .dout(n2568));
  jand g2306(.dina(n1918), .dinb(n432), .dout(n2569));
  jor  g2307(.dina(n2569), .dinb(n2568), .dout(n2570));
  jand g2308(.dina(n1954), .dinb(n485), .dout(n2571));
  jand g2309(.dina(n1935), .dinb(n377), .dout(n2572));
  jor  g2310(.dina(n2572), .dinb(n2571), .dout(n2573));
  jor  g2311(.dina(n2573), .dinb(n2570), .dout(n2574));
  jand g2312(.dina(n2574), .dinb(n263), .dout(n2575));
  jand g2313(.dina(n1946), .dinb(n432), .dout(n2576));
  jand g2314(.dina(n1910), .dinb(n485), .dout(n2577));
  jor  g2315(.dina(n2577), .dinb(n2576), .dout(n2578));
  jand g2316(.dina(n1963), .dinb(n377), .dout(n2579));
  jand g2317(.dina(n1971), .dinb(n323), .dout(n2580));
  jor  g2318(.dina(n2580), .dinb(n2579), .dout(n2581));
  jor  g2319(.dina(n2581), .dinb(n2578), .dout(n2582));
  jand g2320(.dina(n2582), .dinb(shift6 ), .dout(n2583));
  jor  g2321(.dina(n2583), .dinb(n2575), .dout(result25 ));
  jand g2322(.dina(n2000), .dinb(n323), .dout(n2585));
  jand g2323(.dina(n2008), .dinb(n377), .dout(n2586));
  jor  g2324(.dina(n2586), .dinb(n2585), .dout(n2587));
  jand g2325(.dina(n1991), .dinb(n432), .dout(n2588));
  jand g2326(.dina(n2027), .dinb(n485), .dout(n2589));
  jor  g2327(.dina(n2589), .dinb(n2588), .dout(n2590));
  jor  g2328(.dina(n2590), .dinb(n2587), .dout(n2591));
  jand g2329(.dina(n2591), .dinb(n263), .dout(n2592));
  jand g2330(.dina(n2019), .dinb(n432), .dout(n2593));
  jand g2331(.dina(n1983), .dinb(n485), .dout(n2594));
  jor  g2332(.dina(n2594), .dinb(n2593), .dout(n2595));
  jand g2333(.dina(n2036), .dinb(n377), .dout(n2596));
  jand g2334(.dina(n2044), .dinb(n323), .dout(n2597));
  jor  g2335(.dina(n2597), .dinb(n2596), .dout(n2598));
  jor  g2336(.dina(n2598), .dinb(n2595), .dout(n2599));
  jand g2337(.dina(n2599), .dinb(shift6 ), .dout(n2600));
  jor  g2338(.dina(n2600), .dinb(n2592), .dout(result26 ));
  jand g2339(.dina(n2073), .dinb(n323), .dout(n2602));
  jand g2340(.dina(n2081), .dinb(n377), .dout(n2603));
  jor  g2341(.dina(n2603), .dinb(n2602), .dout(n2604));
  jand g2342(.dina(n2064), .dinb(n432), .dout(n2605));
  jand g2343(.dina(n2100), .dinb(n485), .dout(n2606));
  jor  g2344(.dina(n2606), .dinb(n2605), .dout(n2607));
  jor  g2345(.dina(n2607), .dinb(n2604), .dout(n2608));
  jand g2346(.dina(n2608), .dinb(n263), .dout(n2609));
  jand g2347(.dina(n2092), .dinb(n432), .dout(n2610));
  jand g2348(.dina(n2056), .dinb(n485), .dout(n2611));
  jor  g2349(.dina(n2611), .dinb(n2610), .dout(n2612));
  jand g2350(.dina(n2109), .dinb(n377), .dout(n2613));
  jand g2351(.dina(n2117), .dinb(n323), .dout(n2614));
  jor  g2352(.dina(n2614), .dinb(n2613), .dout(n2615));
  jor  g2353(.dina(n2615), .dinb(n2612), .dout(n2616));
  jand g2354(.dina(n2616), .dinb(shift6 ), .dout(n2617));
  jor  g2355(.dina(n2617), .dinb(n2609), .dout(result27 ));
  jand g2356(.dina(n2146), .dinb(n323), .dout(n2619));
  jand g2357(.dina(n2154), .dinb(n377), .dout(n2620));
  jor  g2358(.dina(n2620), .dinb(n2619), .dout(n2621));
  jand g2359(.dina(n2137), .dinb(n432), .dout(n2622));
  jand g2360(.dina(n2173), .dinb(n485), .dout(n2623));
  jor  g2361(.dina(n2623), .dinb(n2622), .dout(n2624));
  jor  g2362(.dina(n2624), .dinb(n2621), .dout(n2625));
  jand g2363(.dina(n2625), .dinb(n263), .dout(n2626));
  jand g2364(.dina(n2165), .dinb(n432), .dout(n2627));
  jand g2365(.dina(n2129), .dinb(n485), .dout(n2628));
  jor  g2366(.dina(n2628), .dinb(n2627), .dout(n2629));
  jand g2367(.dina(n2182), .dinb(n377), .dout(n2630));
  jand g2368(.dina(n2190), .dinb(n323), .dout(n2631));
  jor  g2369(.dina(n2631), .dinb(n2630), .dout(n2632));
  jor  g2370(.dina(n2632), .dinb(n2629), .dout(n2633));
  jand g2371(.dina(n2633), .dinb(shift6 ), .dout(n2634));
  jor  g2372(.dina(n2634), .dinb(n2626), .dout(result28 ));
  jand g2373(.dina(n2219), .dinb(n323), .dout(n2636));
  jand g2374(.dina(n2227), .dinb(n377), .dout(n2637));
  jor  g2375(.dina(n2637), .dinb(n2636), .dout(n2638));
  jand g2376(.dina(n2210), .dinb(n432), .dout(n2639));
  jand g2377(.dina(n2246), .dinb(n485), .dout(n2640));
  jor  g2378(.dina(n2640), .dinb(n2639), .dout(n2641));
  jor  g2379(.dina(n2641), .dinb(n2638), .dout(n2642));
  jand g2380(.dina(n2642), .dinb(n263), .dout(n2643));
  jand g2381(.dina(n2238), .dinb(n432), .dout(n2644));
  jand g2382(.dina(n2202), .dinb(n485), .dout(n2645));
  jor  g2383(.dina(n2645), .dinb(n2644), .dout(n2646));
  jand g2384(.dina(n2255), .dinb(n377), .dout(n2647));
  jand g2385(.dina(n2263), .dinb(n323), .dout(n2648));
  jor  g2386(.dina(n2648), .dinb(n2647), .dout(n2649));
  jor  g2387(.dina(n2649), .dinb(n2646), .dout(n2650));
  jand g2388(.dina(n2650), .dinb(shift6 ), .dout(n2651));
  jor  g2389(.dina(n2651), .dinb(n2643), .dout(result29 ));
  jand g2390(.dina(n2292), .dinb(n323), .dout(n2653));
  jand g2391(.dina(n2300), .dinb(n377), .dout(n2654));
  jor  g2392(.dina(n2654), .dinb(n2653), .dout(n2655));
  jand g2393(.dina(n2283), .dinb(n432), .dout(n2656));
  jand g2394(.dina(n2319), .dinb(n485), .dout(n2657));
  jor  g2395(.dina(n2657), .dinb(n2656), .dout(n2658));
  jor  g2396(.dina(n2658), .dinb(n2655), .dout(n2659));
  jand g2397(.dina(n2659), .dinb(n263), .dout(n2660));
  jand g2398(.dina(n2311), .dinb(n432), .dout(n2661));
  jand g2399(.dina(n2275), .dinb(n485), .dout(n2662));
  jor  g2400(.dina(n2662), .dinb(n2661), .dout(n2663));
  jand g2401(.dina(n2328), .dinb(n377), .dout(n2664));
  jand g2402(.dina(n2336), .dinb(n323), .dout(n2665));
  jor  g2403(.dina(n2665), .dinb(n2664), .dout(n2666));
  jor  g2404(.dina(n2666), .dinb(n2663), .dout(n2667));
  jand g2405(.dina(n2667), .dinb(shift6 ), .dout(n2668));
  jor  g2406(.dina(n2668), .dinb(n2660), .dout(result30 ));
  jand g2407(.dina(n2365), .dinb(n323), .dout(n2670));
  jand g2408(.dina(n2373), .dinb(n377), .dout(n2671));
  jor  g2409(.dina(n2671), .dinb(n2670), .dout(n2672));
  jand g2410(.dina(n2356), .dinb(n432), .dout(n2673));
  jand g2411(.dina(n2392), .dinb(n485), .dout(n2674));
  jor  g2412(.dina(n2674), .dinb(n2673), .dout(n2675));
  jor  g2413(.dina(n2675), .dinb(n2672), .dout(n2676));
  jand g2414(.dina(n2676), .dinb(n263), .dout(n2677));
  jand g2415(.dina(n2384), .dinb(n432), .dout(n2678));
  jand g2416(.dina(n2348), .dinb(n485), .dout(n2679));
  jor  g2417(.dina(n2679), .dinb(n2678), .dout(n2680));
  jand g2418(.dina(n2401), .dinb(n377), .dout(n2681));
  jand g2419(.dina(n2409), .dinb(n323), .dout(n2682));
  jor  g2420(.dina(n2682), .dinb(n2681), .dout(n2683));
  jor  g2421(.dina(n2683), .dinb(n2680), .dout(n2684));
  jand g2422(.dina(n2684), .dinb(shift6 ), .dout(n2685));
  jor  g2423(.dina(n2685), .dinb(n2677), .dout(result31 ));
  jand g2424(.dina(n375), .dinb(n323), .dout(n2687));
  jand g2425(.dina(n540), .dinb(n377), .dout(n2688));
  jor  g2426(.dina(n2688), .dinb(n2687), .dout(n2689));
  jand g2427(.dina(n484), .dinb(n432), .dout(n2690));
  jand g2428(.dina(n643), .dinb(n485), .dout(n2691));
  jor  g2429(.dina(n2691), .dinb(n2690), .dout(n2692));
  jor  g2430(.dina(n2692), .dinb(n2689), .dout(n2693));
  jand g2431(.dina(n2693), .dinb(n263), .dout(n2694));
  jand g2432(.dina(n377), .dinb(n322), .dout(n2695));
  jand g2433(.dina(n590), .dinb(n323), .dout(n2696));
  jor  g2434(.dina(n2696), .dinb(n2695), .dout(n2697));
  jand g2435(.dina(n485), .dinb(n430), .dout(n2698));
  jand g2436(.dina(n695), .dinb(n432), .dout(n2699));
  jor  g2437(.dina(n2699), .dinb(n2698), .dout(n2700));
  jor  g2438(.dina(n2700), .dinb(n2697), .dout(n2701));
  jand g2439(.dina(n2701), .dinb(shift6 ), .dout(n2702));
  jor  g2440(.dina(n2702), .dinb(n2694), .dout(result32 ));
  jand g2441(.dina(n787), .dinb(n323), .dout(n2704));
  jand g2442(.dina(n1012), .dinb(n377), .dout(n2705));
  jor  g2443(.dina(n2705), .dinb(n2704), .dout(n2706));
  jand g2444(.dina(n876), .dinb(n432), .dout(n2707));
  jand g2445(.dina(n967), .dinb(n485), .dout(n2708));
  jor  g2446(.dina(n2708), .dinb(n2707), .dout(n2709));
  jor  g2447(.dina(n2709), .dinb(n2706), .dout(n2710));
  jand g2448(.dina(n2710), .dinb(n263), .dout(n2711));
  jand g2449(.dina(n923), .dinb(n432), .dout(n2712));
  jand g2450(.dina(n832), .dinb(n485), .dout(n2713));
  jor  g2451(.dina(n2713), .dinb(n2712), .dout(n2714));
  jand g2452(.dina(n743), .dinb(n377), .dout(n2715));
  jand g2453(.dina(n1060), .dinb(n323), .dout(n2716));
  jor  g2454(.dina(n2716), .dinb(n2715), .dout(n2717));
  jor  g2455(.dina(n2717), .dinb(n2714), .dout(n2718));
  jand g2456(.dina(n2718), .dinb(shift6 ), .dout(n2719));
  jor  g2457(.dina(n2719), .dinb(n2711), .dout(result33 ));
  jand g2458(.dina(n1136), .dinb(n323), .dout(n2721));
  jand g2459(.dina(n1321), .dinb(n377), .dout(n2722));
  jor  g2460(.dina(n2722), .dinb(n2721), .dout(n2723));
  jand g2461(.dina(n1209), .dinb(n432), .dout(n2724));
  jand g2462(.dina(n1284), .dinb(n485), .dout(n2725));
  jor  g2463(.dina(n2725), .dinb(n2724), .dout(n2726));
  jor  g2464(.dina(n2726), .dinb(n2723), .dout(n2727));
  jand g2465(.dina(n2727), .dinb(n263), .dout(n2728));
  jand g2466(.dina(n1248), .dinb(n432), .dout(n2729));
  jand g2467(.dina(n1173), .dinb(n485), .dout(n2730));
  jor  g2468(.dina(n2730), .dinb(n2729), .dout(n2731));
  jand g2469(.dina(n1100), .dinb(n377), .dout(n2732));
  jand g2470(.dina(n1357), .dinb(n323), .dout(n2733));
  jor  g2471(.dina(n2733), .dinb(n2732), .dout(n2734));
  jor  g2472(.dina(n2734), .dinb(n2731), .dout(n2735));
  jand g2473(.dina(n2735), .dinb(shift6 ), .dout(n2736));
  jor  g2474(.dina(n2736), .dinb(n2728), .dout(result34 ));
  jand g2475(.dina(n1381), .dinb(n323), .dout(n2738));
  jand g2476(.dina(n1533), .dinb(n377), .dout(n2739));
  jor  g2477(.dina(n2739), .dinb(n2738), .dout(n2740));
  jand g2478(.dina(n1485), .dinb(n485), .dout(n2741));
  jand g2479(.dina(n1442), .dinb(n432), .dout(n2742));
  jor  g2480(.dina(n2742), .dinb(n2741), .dout(n2743));
  jor  g2481(.dina(n2743), .dinb(n2740), .dout(n2744));
  jand g2482(.dina(n2744), .dinb(n263), .dout(n2745));
  jand g2483(.dina(n1465), .dinb(n432), .dout(n2746));
  jand g2484(.dina(n1401), .dinb(n377), .dout(n2747));
  jor  g2485(.dina(n2747), .dinb(n2746), .dout(n2748));
  jand g2486(.dina(n1422), .dinb(n485), .dout(n2749));
  jand g2487(.dina(n1513), .dinb(n323), .dout(n2750));
  jor  g2488(.dina(n2750), .dinb(n2749), .dout(n2751));
  jor  g2489(.dina(n2751), .dinb(n2748), .dout(n2752));
  jand g2490(.dina(n2752), .dinb(shift6 ), .dout(n2753));
  jor  g2491(.dina(n2753), .dinb(n2745), .dout(result35 ));
  jand g2492(.dina(n1553), .dinb(n323), .dout(n2755));
  jand g2493(.dina(n1589), .dinb(n377), .dout(n2756));
  jor  g2494(.dina(n2756), .dinb(n2755), .dout(n2757));
  jand g2495(.dina(n1570), .dinb(n432), .dout(n2758));
  jand g2496(.dina(n1606), .dinb(n485), .dout(n2759));
  jor  g2497(.dina(n2759), .dinb(n2758), .dout(n2760));
  jor  g2498(.dina(n2760), .dinb(n2757), .dout(n2761));
  jand g2499(.dina(n2761), .dinb(n263), .dout(n2762));
  jand g2500(.dina(n1545), .dinb(n377), .dout(n2763));
  jand g2501(.dina(n1581), .dinb(n323), .dout(n2764));
  jor  g2502(.dina(n2764), .dinb(n2763), .dout(n2765));
  jand g2503(.dina(n1562), .dinb(n485), .dout(n2766));
  jand g2504(.dina(n1598), .dinb(n432), .dout(n2767));
  jor  g2505(.dina(n2767), .dinb(n2766), .dout(n2768));
  jor  g2506(.dina(n2768), .dinb(n2765), .dout(n2769));
  jand g2507(.dina(n2769), .dinb(shift6 ), .dout(n2770));
  jor  g2508(.dina(n2770), .dinb(n2762), .dout(result36 ));
  jand g2509(.dina(n1626), .dinb(n323), .dout(n2772));
  jand g2510(.dina(n1662), .dinb(n377), .dout(n2773));
  jor  g2511(.dina(n2773), .dinb(n2772), .dout(n2774));
  jand g2512(.dina(n1643), .dinb(n432), .dout(n2775));
  jand g2513(.dina(n1679), .dinb(n485), .dout(n2776));
  jor  g2514(.dina(n2776), .dinb(n2775), .dout(n2777));
  jor  g2515(.dina(n2777), .dinb(n2774), .dout(n2778));
  jand g2516(.dina(n2778), .dinb(n263), .dout(n2779));
  jand g2517(.dina(n1618), .dinb(n377), .dout(n2780));
  jand g2518(.dina(n1654), .dinb(n323), .dout(n2781));
  jor  g2519(.dina(n2781), .dinb(n2780), .dout(n2782));
  jand g2520(.dina(n1635), .dinb(n485), .dout(n2783));
  jand g2521(.dina(n1671), .dinb(n432), .dout(n2784));
  jor  g2522(.dina(n2784), .dinb(n2783), .dout(n2785));
  jor  g2523(.dina(n2785), .dinb(n2782), .dout(n2786));
  jand g2524(.dina(n2786), .dinb(shift6 ), .dout(n2787));
  jor  g2525(.dina(n2787), .dinb(n2779), .dout(result37 ));
  jand g2526(.dina(n1699), .dinb(n323), .dout(n2789));
  jand g2527(.dina(n1735), .dinb(n377), .dout(n2790));
  jor  g2528(.dina(n2790), .dinb(n2789), .dout(n2791));
  jand g2529(.dina(n1716), .dinb(n432), .dout(n2792));
  jand g2530(.dina(n1752), .dinb(n485), .dout(n2793));
  jor  g2531(.dina(n2793), .dinb(n2792), .dout(n2794));
  jor  g2532(.dina(n2794), .dinb(n2791), .dout(n2795));
  jand g2533(.dina(n2795), .dinb(n263), .dout(n2796));
  jand g2534(.dina(n1691), .dinb(n377), .dout(n2797));
  jand g2535(.dina(n1727), .dinb(n323), .dout(n2798));
  jor  g2536(.dina(n2798), .dinb(n2797), .dout(n2799));
  jand g2537(.dina(n1708), .dinb(n485), .dout(n2800));
  jand g2538(.dina(n1744), .dinb(n432), .dout(n2801));
  jor  g2539(.dina(n2801), .dinb(n2800), .dout(n2802));
  jor  g2540(.dina(n2802), .dinb(n2799), .dout(n2803));
  jand g2541(.dina(n2803), .dinb(shift6 ), .dout(n2804));
  jor  g2542(.dina(n2804), .dinb(n2796), .dout(result38 ));
  jand g2543(.dina(n1808), .dinb(n377), .dout(n2806));
  jand g2544(.dina(n1772), .dinb(n323), .dout(n2807));
  jor  g2545(.dina(n2807), .dinb(n2806), .dout(n2808));
  jand g2546(.dina(n1825), .dinb(n485), .dout(n2809));
  jand g2547(.dina(n1789), .dinb(n432), .dout(n2810));
  jor  g2548(.dina(n2810), .dinb(n2809), .dout(n2811));
  jor  g2549(.dina(n2811), .dinb(n2808), .dout(n2812));
  jand g2550(.dina(n2812), .dinb(n263), .dout(n2813));
  jand g2551(.dina(n1800), .dinb(n323), .dout(n2814));
  jand g2552(.dina(n1764), .dinb(n377), .dout(n2815));
  jor  g2553(.dina(n2815), .dinb(n2814), .dout(n2816));
  jand g2554(.dina(n1817), .dinb(n432), .dout(n2817));
  jand g2555(.dina(n1781), .dinb(n485), .dout(n2818));
  jor  g2556(.dina(n2818), .dinb(n2817), .dout(n2819));
  jor  g2557(.dina(n2819), .dinb(n2816), .dout(n2820));
  jand g2558(.dina(n2820), .dinb(shift6 ), .dout(n2821));
  jor  g2559(.dina(n2821), .dinb(n2813), .dout(result39 ));
  jand g2560(.dina(n1881), .dinb(n377), .dout(n2823));
  jand g2561(.dina(n1845), .dinb(n323), .dout(n2824));
  jor  g2562(.dina(n2824), .dinb(n2823), .dout(n2825));
  jand g2563(.dina(n1898), .dinb(n485), .dout(n2826));
  jand g2564(.dina(n1862), .dinb(n432), .dout(n2827));
  jor  g2565(.dina(n2827), .dinb(n2826), .dout(n2828));
  jor  g2566(.dina(n2828), .dinb(n2825), .dout(n2829));
  jand g2567(.dina(n2829), .dinb(n263), .dout(n2830));
  jand g2568(.dina(n1873), .dinb(n323), .dout(n2831));
  jand g2569(.dina(n1837), .dinb(n377), .dout(n2832));
  jor  g2570(.dina(n2832), .dinb(n2831), .dout(n2833));
  jand g2571(.dina(n1890), .dinb(n432), .dout(n2834));
  jand g2572(.dina(n1854), .dinb(n485), .dout(n2835));
  jor  g2573(.dina(n2835), .dinb(n2834), .dout(n2836));
  jor  g2574(.dina(n2836), .dinb(n2833), .dout(n2837));
  jand g2575(.dina(n2837), .dinb(shift6 ), .dout(n2838));
  jor  g2576(.dina(n2838), .dinb(n2830), .dout(result40 ));
  jand g2577(.dina(n1954), .dinb(n377), .dout(n2840));
  jand g2578(.dina(n1918), .dinb(n323), .dout(n2841));
  jor  g2579(.dina(n2841), .dinb(n2840), .dout(n2842));
  jand g2580(.dina(n1971), .dinb(n485), .dout(n2843));
  jand g2581(.dina(n1935), .dinb(n432), .dout(n2844));
  jor  g2582(.dina(n2844), .dinb(n2843), .dout(n2845));
  jor  g2583(.dina(n2845), .dinb(n2842), .dout(n2846));
  jand g2584(.dina(n2846), .dinb(n263), .dout(n2847));
  jand g2585(.dina(n1946), .dinb(n323), .dout(n2848));
  jand g2586(.dina(n1910), .dinb(n377), .dout(n2849));
  jor  g2587(.dina(n2849), .dinb(n2848), .dout(n2850));
  jand g2588(.dina(n1963), .dinb(n432), .dout(n2851));
  jand g2589(.dina(n1927), .dinb(n485), .dout(n2852));
  jor  g2590(.dina(n2852), .dinb(n2851), .dout(n2853));
  jor  g2591(.dina(n2853), .dinb(n2850), .dout(n2854));
  jand g2592(.dina(n2854), .dinb(shift6 ), .dout(n2855));
  jor  g2593(.dina(n2855), .dinb(n2847), .dout(result41 ));
  jand g2594(.dina(n1991), .dinb(n323), .dout(n2857));
  jand g2595(.dina(n2027), .dinb(n377), .dout(n2858));
  jor  g2596(.dina(n2858), .dinb(n2857), .dout(n2859));
  jand g2597(.dina(n2008), .dinb(n432), .dout(n2860));
  jand g2598(.dina(n2044), .dinb(n485), .dout(n2861));
  jor  g2599(.dina(n2861), .dinb(n2860), .dout(n2862));
  jor  g2600(.dina(n2862), .dinb(n2859), .dout(n2863));
  jand g2601(.dina(n2863), .dinb(n263), .dout(n2864));
  jand g2602(.dina(n2019), .dinb(n323), .dout(n2865));
  jand g2603(.dina(n1983), .dinb(n377), .dout(n2866));
  jor  g2604(.dina(n2866), .dinb(n2865), .dout(n2867));
  jand g2605(.dina(n2036), .dinb(n432), .dout(n2868));
  jand g2606(.dina(n2000), .dinb(n485), .dout(n2869));
  jor  g2607(.dina(n2869), .dinb(n2868), .dout(n2870));
  jor  g2608(.dina(n2870), .dinb(n2867), .dout(n2871));
  jand g2609(.dina(n2871), .dinb(shift6 ), .dout(n2872));
  jor  g2610(.dina(n2872), .dinb(n2864), .dout(result42 ));
  jand g2611(.dina(n2064), .dinb(n323), .dout(n2874));
  jand g2612(.dina(n2100), .dinb(n377), .dout(n2875));
  jor  g2613(.dina(n2875), .dinb(n2874), .dout(n2876));
  jand g2614(.dina(n2081), .dinb(n432), .dout(n2877));
  jand g2615(.dina(n2117), .dinb(n485), .dout(n2878));
  jor  g2616(.dina(n2878), .dinb(n2877), .dout(n2879));
  jor  g2617(.dina(n2879), .dinb(n2876), .dout(n2880));
  jand g2618(.dina(n2880), .dinb(n263), .dout(n2881));
  jand g2619(.dina(n2092), .dinb(n323), .dout(n2882));
  jand g2620(.dina(n2056), .dinb(n377), .dout(n2883));
  jor  g2621(.dina(n2883), .dinb(n2882), .dout(n2884));
  jand g2622(.dina(n2109), .dinb(n432), .dout(n2885));
  jand g2623(.dina(n2073), .dinb(n485), .dout(n2886));
  jor  g2624(.dina(n2886), .dinb(n2885), .dout(n2887));
  jor  g2625(.dina(n2887), .dinb(n2884), .dout(n2888));
  jand g2626(.dina(n2888), .dinb(shift6 ), .dout(n2889));
  jor  g2627(.dina(n2889), .dinb(n2881), .dout(result43 ));
  jand g2628(.dina(n2137), .dinb(n323), .dout(n2891));
  jand g2629(.dina(n2173), .dinb(n377), .dout(n2892));
  jor  g2630(.dina(n2892), .dinb(n2891), .dout(n2893));
  jand g2631(.dina(n2154), .dinb(n432), .dout(n2894));
  jand g2632(.dina(n2190), .dinb(n485), .dout(n2895));
  jor  g2633(.dina(n2895), .dinb(n2894), .dout(n2896));
  jor  g2634(.dina(n2896), .dinb(n2893), .dout(n2897));
  jand g2635(.dina(n2897), .dinb(n263), .dout(n2898));
  jand g2636(.dina(n2165), .dinb(n323), .dout(n2899));
  jand g2637(.dina(n2129), .dinb(n377), .dout(n2900));
  jor  g2638(.dina(n2900), .dinb(n2899), .dout(n2901));
  jand g2639(.dina(n2182), .dinb(n432), .dout(n2902));
  jand g2640(.dina(n2146), .dinb(n485), .dout(n2903));
  jor  g2641(.dina(n2903), .dinb(n2902), .dout(n2904));
  jor  g2642(.dina(n2904), .dinb(n2901), .dout(n2905));
  jand g2643(.dina(n2905), .dinb(shift6 ), .dout(n2906));
  jor  g2644(.dina(n2906), .dinb(n2898), .dout(result44 ));
  jand g2645(.dina(n2210), .dinb(n323), .dout(n2908));
  jand g2646(.dina(n2246), .dinb(n377), .dout(n2909));
  jor  g2647(.dina(n2909), .dinb(n2908), .dout(n2910));
  jand g2648(.dina(n2227), .dinb(n432), .dout(n2911));
  jand g2649(.dina(n2263), .dinb(n485), .dout(n2912));
  jor  g2650(.dina(n2912), .dinb(n2911), .dout(n2913));
  jor  g2651(.dina(n2913), .dinb(n2910), .dout(n2914));
  jand g2652(.dina(n2914), .dinb(n263), .dout(n2915));
  jand g2653(.dina(n2238), .dinb(n323), .dout(n2916));
  jand g2654(.dina(n2202), .dinb(n377), .dout(n2917));
  jor  g2655(.dina(n2917), .dinb(n2916), .dout(n2918));
  jand g2656(.dina(n2255), .dinb(n432), .dout(n2919));
  jand g2657(.dina(n2219), .dinb(n485), .dout(n2920));
  jor  g2658(.dina(n2920), .dinb(n2919), .dout(n2921));
  jor  g2659(.dina(n2921), .dinb(n2918), .dout(n2922));
  jand g2660(.dina(n2922), .dinb(shift6 ), .dout(n2923));
  jor  g2661(.dina(n2923), .dinb(n2915), .dout(result45 ));
  jand g2662(.dina(n2283), .dinb(n323), .dout(n2925));
  jand g2663(.dina(n2319), .dinb(n377), .dout(n2926));
  jor  g2664(.dina(n2926), .dinb(n2925), .dout(n2927));
  jand g2665(.dina(n2300), .dinb(n432), .dout(n2928));
  jand g2666(.dina(n2336), .dinb(n485), .dout(n2929));
  jor  g2667(.dina(n2929), .dinb(n2928), .dout(n2930));
  jor  g2668(.dina(n2930), .dinb(n2927), .dout(n2931));
  jand g2669(.dina(n2931), .dinb(n263), .dout(n2932));
  jand g2670(.dina(n2311), .dinb(n323), .dout(n2933));
  jand g2671(.dina(n2275), .dinb(n377), .dout(n2934));
  jor  g2672(.dina(n2934), .dinb(n2933), .dout(n2935));
  jand g2673(.dina(n2328), .dinb(n432), .dout(n2936));
  jand g2674(.dina(n2292), .dinb(n485), .dout(n2937));
  jor  g2675(.dina(n2937), .dinb(n2936), .dout(n2938));
  jor  g2676(.dina(n2938), .dinb(n2935), .dout(n2939));
  jand g2677(.dina(n2939), .dinb(shift6 ), .dout(n2940));
  jor  g2678(.dina(n2940), .dinb(n2932), .dout(result46 ));
  jand g2679(.dina(n2356), .dinb(n323), .dout(n2942));
  jand g2680(.dina(n2392), .dinb(n377), .dout(n2943));
  jor  g2681(.dina(n2943), .dinb(n2942), .dout(n2944));
  jand g2682(.dina(n2373), .dinb(n432), .dout(n2945));
  jand g2683(.dina(n2409), .dinb(n485), .dout(n2946));
  jor  g2684(.dina(n2946), .dinb(n2945), .dout(n2947));
  jor  g2685(.dina(n2947), .dinb(n2944), .dout(n2948));
  jand g2686(.dina(n2948), .dinb(n263), .dout(n2949));
  jand g2687(.dina(n2384), .dinb(n323), .dout(n2950));
  jand g2688(.dina(n2348), .dinb(n377), .dout(n2951));
  jor  g2689(.dina(n2951), .dinb(n2950), .dout(n2952));
  jand g2690(.dina(n2401), .dinb(n432), .dout(n2953));
  jand g2691(.dina(n2365), .dinb(n485), .dout(n2954));
  jor  g2692(.dina(n2954), .dinb(n2953), .dout(n2955));
  jor  g2693(.dina(n2955), .dinb(n2952), .dout(n2956));
  jand g2694(.dina(n2956), .dinb(shift6 ), .dout(n2957));
  jor  g2695(.dina(n2957), .dinb(n2949), .dout(result47 ));
  jand g2696(.dina(n484), .dinb(n323), .dout(n2959));
  jand g2697(.dina(n643), .dinb(n377), .dout(n2960));
  jor  g2698(.dina(n2960), .dinb(n2959), .dout(n2961));
  jand g2699(.dina(n540), .dinb(n432), .dout(n2962));
  jand g2700(.dina(n590), .dinb(n485), .dout(n2963));
  jor  g2701(.dina(n2963), .dinb(n2962), .dout(n2964));
  jor  g2702(.dina(n2964), .dinb(n2961), .dout(n2965));
  jand g2703(.dina(n2965), .dinb(n263), .dout(n2966));
  jand g2704(.dina(n432), .dinb(n322), .dout(n2967));
  jand g2705(.dina(n485), .dinb(n375), .dout(n2968));
  jor  g2706(.dina(n2968), .dinb(n2967), .dout(n2969));
  jand g2707(.dina(n430), .dinb(n377), .dout(n2970));
  jand g2708(.dina(n695), .dinb(n323), .dout(n2971));
  jor  g2709(.dina(n2971), .dinb(n2970), .dout(n2972));
  jor  g2710(.dina(n2972), .dinb(n2969), .dout(n2973));
  jand g2711(.dina(n2973), .dinb(shift6 ), .dout(n2974));
  jor  g2712(.dina(n2974), .dinb(n2966), .dout(result48 ));
  jand g2713(.dina(n876), .dinb(n323), .dout(n2976));
  jand g2714(.dina(n967), .dinb(n377), .dout(n2977));
  jor  g2715(.dina(n2977), .dinb(n2976), .dout(n2978));
  jand g2716(.dina(n1012), .dinb(n432), .dout(n2979));
  jand g2717(.dina(n1060), .dinb(n485), .dout(n2980));
  jor  g2718(.dina(n2980), .dinb(n2979), .dout(n2981));
  jor  g2719(.dina(n2981), .dinb(n2978), .dout(n2982));
  jand g2720(.dina(n2982), .dinb(n263), .dout(n2983));
  jand g2721(.dina(n923), .dinb(n323), .dout(n2984));
  jand g2722(.dina(n832), .dinb(n377), .dout(n2985));
  jor  g2723(.dina(n2985), .dinb(n2984), .dout(n2986));
  jand g2724(.dina(n743), .dinb(n432), .dout(n2987));
  jand g2725(.dina(n787), .dinb(n485), .dout(n2988));
  jor  g2726(.dina(n2988), .dinb(n2987), .dout(n2989));
  jor  g2727(.dina(n2989), .dinb(n2986), .dout(n2990));
  jand g2728(.dina(n2990), .dinb(shift6 ), .dout(n2991));
  jor  g2729(.dina(n2991), .dinb(n2983), .dout(result49 ));
  jand g2730(.dina(n1209), .dinb(n323), .dout(n2993));
  jand g2731(.dina(n1284), .dinb(n377), .dout(n2994));
  jor  g2732(.dina(n2994), .dinb(n2993), .dout(n2995));
  jand g2733(.dina(n1321), .dinb(n432), .dout(n2996));
  jand g2734(.dina(n1357), .dinb(n485), .dout(n2997));
  jor  g2735(.dina(n2997), .dinb(n2996), .dout(n2998));
  jor  g2736(.dina(n2998), .dinb(n2995), .dout(n2999));
  jand g2737(.dina(n2999), .dinb(n263), .dout(n3000));
  jand g2738(.dina(n1248), .dinb(n323), .dout(n3001));
  jand g2739(.dina(n1173), .dinb(n377), .dout(n3002));
  jor  g2740(.dina(n3002), .dinb(n3001), .dout(n3003));
  jand g2741(.dina(n1100), .dinb(n432), .dout(n3004));
  jand g2742(.dina(n1136), .dinb(n485), .dout(n3005));
  jor  g2743(.dina(n3005), .dinb(n3004), .dout(n3006));
  jor  g2744(.dina(n3006), .dinb(n3003), .dout(n3007));
  jand g2745(.dina(n3007), .dinb(shift6 ), .dout(n3008));
  jor  g2746(.dina(n3008), .dinb(n3000), .dout(result50 ));
  jand g2747(.dina(n1513), .dinb(n485), .dout(n3010));
  jand g2748(.dina(n1533), .dinb(n432), .dout(n3011));
  jor  g2749(.dina(n3011), .dinb(n3010), .dout(n3012));
  jand g2750(.dina(n1485), .dinb(n377), .dout(n3013));
  jand g2751(.dina(n1442), .dinb(n323), .dout(n3014));
  jor  g2752(.dina(n3014), .dinb(n3013), .dout(n3015));
  jor  g2753(.dina(n3015), .dinb(n3012), .dout(n3016));
  jand g2754(.dina(n3016), .dinb(n263), .dout(n3017));
  jand g2755(.dina(n1465), .dinb(n323), .dout(n3018));
  jand g2756(.dina(n1422), .dinb(n377), .dout(n3019));
  jor  g2757(.dina(n3019), .dinb(n3018), .dout(n3020));
  jand g2758(.dina(n1381), .dinb(n485), .dout(n3021));
  jand g2759(.dina(n1401), .dinb(n432), .dout(n3022));
  jor  g2760(.dina(n3022), .dinb(n3021), .dout(n3023));
  jor  g2761(.dina(n3023), .dinb(n3020), .dout(n3024));
  jand g2762(.dina(n3024), .dinb(shift6 ), .dout(n3025));
  jor  g2763(.dina(n3025), .dinb(n3017), .dout(result51 ));
  jand g2764(.dina(n1581), .dinb(n485), .dout(n3027));
  jand g2765(.dina(n1589), .dinb(n432), .dout(n3028));
  jor  g2766(.dina(n3028), .dinb(n3027), .dout(n3029));
  jand g2767(.dina(n1570), .dinb(n323), .dout(n3030));
  jand g2768(.dina(n1606), .dinb(n377), .dout(n3031));
  jor  g2769(.dina(n3031), .dinb(n3030), .dout(n3032));
  jor  g2770(.dina(n3032), .dinb(n3029), .dout(n3033));
  jand g2771(.dina(n3033), .dinb(n263), .dout(n3034));
  jand g2772(.dina(n1545), .dinb(n432), .dout(n3035));
  jand g2773(.dina(n1598), .dinb(n323), .dout(n3036));
  jor  g2774(.dina(n3036), .dinb(n3035), .dout(n3037));
  jand g2775(.dina(n1562), .dinb(n377), .dout(n3038));
  jand g2776(.dina(n1553), .dinb(n485), .dout(n3039));
  jor  g2777(.dina(n3039), .dinb(n3038), .dout(n3040));
  jor  g2778(.dina(n3040), .dinb(n3037), .dout(n3041));
  jand g2779(.dina(n3041), .dinb(shift6 ), .dout(n3042));
  jor  g2780(.dina(n3042), .dinb(n3034), .dout(result52 ));
  jand g2781(.dina(n1654), .dinb(n485), .dout(n3044));
  jand g2782(.dina(n1662), .dinb(n432), .dout(n3045));
  jor  g2783(.dina(n3045), .dinb(n3044), .dout(n3046));
  jand g2784(.dina(n1643), .dinb(n323), .dout(n3047));
  jand g2785(.dina(n1679), .dinb(n377), .dout(n3048));
  jor  g2786(.dina(n3048), .dinb(n3047), .dout(n3049));
  jor  g2787(.dina(n3049), .dinb(n3046), .dout(n3050));
  jand g2788(.dina(n3050), .dinb(n263), .dout(n3051));
  jand g2789(.dina(n1618), .dinb(n432), .dout(n3052));
  jand g2790(.dina(n1671), .dinb(n323), .dout(n3053));
  jor  g2791(.dina(n3053), .dinb(n3052), .dout(n3054));
  jand g2792(.dina(n1635), .dinb(n377), .dout(n3055));
  jand g2793(.dina(n1626), .dinb(n485), .dout(n3056));
  jor  g2794(.dina(n3056), .dinb(n3055), .dout(n3057));
  jor  g2795(.dina(n3057), .dinb(n3054), .dout(n3058));
  jand g2796(.dina(n3058), .dinb(shift6 ), .dout(n3059));
  jor  g2797(.dina(n3059), .dinb(n3051), .dout(result53 ));
  jand g2798(.dina(n1727), .dinb(n485), .dout(n3061));
  jand g2799(.dina(n1735), .dinb(n432), .dout(n3062));
  jor  g2800(.dina(n3062), .dinb(n3061), .dout(n3063));
  jand g2801(.dina(n1716), .dinb(n323), .dout(n3064));
  jand g2802(.dina(n1752), .dinb(n377), .dout(n3065));
  jor  g2803(.dina(n3065), .dinb(n3064), .dout(n3066));
  jor  g2804(.dina(n3066), .dinb(n3063), .dout(n3067));
  jand g2805(.dina(n3067), .dinb(n263), .dout(n3068));
  jand g2806(.dina(n1691), .dinb(n432), .dout(n3069));
  jand g2807(.dina(n1744), .dinb(n323), .dout(n3070));
  jor  g2808(.dina(n3070), .dinb(n3069), .dout(n3071));
  jand g2809(.dina(n1708), .dinb(n377), .dout(n3072));
  jand g2810(.dina(n1699), .dinb(n485), .dout(n3073));
  jor  g2811(.dina(n3073), .dinb(n3072), .dout(n3074));
  jor  g2812(.dina(n3074), .dinb(n3071), .dout(n3075));
  jand g2813(.dina(n3075), .dinb(shift6 ), .dout(n3076));
  jor  g2814(.dina(n3076), .dinb(n3068), .dout(result54 ));
  jand g2815(.dina(n1800), .dinb(n485), .dout(n3078));
  jand g2816(.dina(n1825), .dinb(n377), .dout(n3079));
  jor  g2817(.dina(n3079), .dinb(n3078), .dout(n3080));
  jand g2818(.dina(n1808), .dinb(n432), .dout(n3081));
  jand g2819(.dina(n1789), .dinb(n323), .dout(n3082));
  jor  g2820(.dina(n3082), .dinb(n3081), .dout(n3083));
  jor  g2821(.dina(n3083), .dinb(n3080), .dout(n3084));
  jand g2822(.dina(n3084), .dinb(n263), .dout(n3085));
  jand g2823(.dina(n1817), .dinb(n323), .dout(n3086));
  jand g2824(.dina(n1781), .dinb(n377), .dout(n3087));
  jor  g2825(.dina(n3087), .dinb(n3086), .dout(n3088));
  jand g2826(.dina(n1764), .dinb(n432), .dout(n3089));
  jand g2827(.dina(n1772), .dinb(n485), .dout(n3090));
  jor  g2828(.dina(n3090), .dinb(n3089), .dout(n3091));
  jor  g2829(.dina(n3091), .dinb(n3088), .dout(n3092));
  jand g2830(.dina(n3092), .dinb(shift6 ), .dout(n3093));
  jor  g2831(.dina(n3093), .dinb(n3085), .dout(result55 ));
  jand g2832(.dina(n1873), .dinb(n485), .dout(n3095));
  jand g2833(.dina(n1898), .dinb(n377), .dout(n3096));
  jor  g2834(.dina(n3096), .dinb(n3095), .dout(n3097));
  jand g2835(.dina(n1881), .dinb(n432), .dout(n3098));
  jand g2836(.dina(n1862), .dinb(n323), .dout(n3099));
  jor  g2837(.dina(n3099), .dinb(n3098), .dout(n3100));
  jor  g2838(.dina(n3100), .dinb(n3097), .dout(n3101));
  jand g2839(.dina(n3101), .dinb(n263), .dout(n3102));
  jand g2840(.dina(n1890), .dinb(n323), .dout(n3103));
  jand g2841(.dina(n1854), .dinb(n377), .dout(n3104));
  jor  g2842(.dina(n3104), .dinb(n3103), .dout(n3105));
  jand g2843(.dina(n1837), .dinb(n432), .dout(n3106));
  jand g2844(.dina(n1845), .dinb(n485), .dout(n3107));
  jor  g2845(.dina(n3107), .dinb(n3106), .dout(n3108));
  jor  g2846(.dina(n3108), .dinb(n3105), .dout(n3109));
  jand g2847(.dina(n3109), .dinb(shift6 ), .dout(n3110));
  jor  g2848(.dina(n3110), .dinb(n3102), .dout(result56 ));
  jand g2849(.dina(n1946), .dinb(n485), .dout(n3112));
  jand g2850(.dina(n1971), .dinb(n377), .dout(n3113));
  jor  g2851(.dina(n3113), .dinb(n3112), .dout(n3114));
  jand g2852(.dina(n1954), .dinb(n432), .dout(n3115));
  jand g2853(.dina(n1935), .dinb(n323), .dout(n3116));
  jor  g2854(.dina(n3116), .dinb(n3115), .dout(n3117));
  jor  g2855(.dina(n3117), .dinb(n3114), .dout(n3118));
  jand g2856(.dina(n3118), .dinb(n263), .dout(n3119));
  jand g2857(.dina(n1963), .dinb(n323), .dout(n3120));
  jand g2858(.dina(n1927), .dinb(n377), .dout(n3121));
  jor  g2859(.dina(n3121), .dinb(n3120), .dout(n3122));
  jand g2860(.dina(n1910), .dinb(n432), .dout(n3123));
  jand g2861(.dina(n1918), .dinb(n485), .dout(n3124));
  jor  g2862(.dina(n3124), .dinb(n3123), .dout(n3125));
  jor  g2863(.dina(n3125), .dinb(n3122), .dout(n3126));
  jand g2864(.dina(n3126), .dinb(shift6 ), .dout(n3127));
  jor  g2865(.dina(n3127), .dinb(n3119), .dout(result57 ));
  jand g2866(.dina(n2019), .dinb(n485), .dout(n3129));
  jand g2867(.dina(n2027), .dinb(n432), .dout(n3130));
  jor  g2868(.dina(n3130), .dinb(n3129), .dout(n3131));
  jand g2869(.dina(n2008), .dinb(n323), .dout(n3132));
  jand g2870(.dina(n2044), .dinb(n377), .dout(n3133));
  jor  g2871(.dina(n3133), .dinb(n3132), .dout(n3134));
  jor  g2872(.dina(n3134), .dinb(n3131), .dout(n3135));
  jand g2873(.dina(n3135), .dinb(n263), .dout(n3136));
  jand g2874(.dina(n2036), .dinb(n323), .dout(n3137));
  jand g2875(.dina(n2000), .dinb(n377), .dout(n3138));
  jor  g2876(.dina(n3138), .dinb(n3137), .dout(n3139));
  jand g2877(.dina(n1983), .dinb(n432), .dout(n3140));
  jand g2878(.dina(n1991), .dinb(n485), .dout(n3141));
  jor  g2879(.dina(n3141), .dinb(n3140), .dout(n3142));
  jor  g2880(.dina(n3142), .dinb(n3139), .dout(n3143));
  jand g2881(.dina(n3143), .dinb(shift6 ), .dout(n3144));
  jor  g2882(.dina(n3144), .dinb(n3136), .dout(result58 ));
  jand g2883(.dina(n2092), .dinb(n485), .dout(n3146));
  jand g2884(.dina(n2100), .dinb(n432), .dout(n3147));
  jor  g2885(.dina(n3147), .dinb(n3146), .dout(n3148));
  jand g2886(.dina(n2081), .dinb(n323), .dout(n3149));
  jand g2887(.dina(n2117), .dinb(n377), .dout(n3150));
  jor  g2888(.dina(n3150), .dinb(n3149), .dout(n3151));
  jor  g2889(.dina(n3151), .dinb(n3148), .dout(n3152));
  jand g2890(.dina(n3152), .dinb(n263), .dout(n3153));
  jand g2891(.dina(n2109), .dinb(n323), .dout(n3154));
  jand g2892(.dina(n2073), .dinb(n377), .dout(n3155));
  jor  g2893(.dina(n3155), .dinb(n3154), .dout(n3156));
  jand g2894(.dina(n2056), .dinb(n432), .dout(n3157));
  jand g2895(.dina(n2064), .dinb(n485), .dout(n3158));
  jor  g2896(.dina(n3158), .dinb(n3157), .dout(n3159));
  jor  g2897(.dina(n3159), .dinb(n3156), .dout(n3160));
  jand g2898(.dina(n3160), .dinb(shift6 ), .dout(n3161));
  jor  g2899(.dina(n3161), .dinb(n3153), .dout(result59 ));
  jand g2900(.dina(n2165), .dinb(n485), .dout(n3163));
  jand g2901(.dina(n2173), .dinb(n432), .dout(n3164));
  jor  g2902(.dina(n3164), .dinb(n3163), .dout(n3165));
  jand g2903(.dina(n2154), .dinb(n323), .dout(n3166));
  jand g2904(.dina(n2190), .dinb(n377), .dout(n3167));
  jor  g2905(.dina(n3167), .dinb(n3166), .dout(n3168));
  jor  g2906(.dina(n3168), .dinb(n3165), .dout(n3169));
  jand g2907(.dina(n3169), .dinb(n263), .dout(n3170));
  jand g2908(.dina(n2182), .dinb(n323), .dout(n3171));
  jand g2909(.dina(n2146), .dinb(n377), .dout(n3172));
  jor  g2910(.dina(n3172), .dinb(n3171), .dout(n3173));
  jand g2911(.dina(n2129), .dinb(n432), .dout(n3174));
  jand g2912(.dina(n2137), .dinb(n485), .dout(n3175));
  jor  g2913(.dina(n3175), .dinb(n3174), .dout(n3176));
  jor  g2914(.dina(n3176), .dinb(n3173), .dout(n3177));
  jand g2915(.dina(n3177), .dinb(shift6 ), .dout(n3178));
  jor  g2916(.dina(n3178), .dinb(n3170), .dout(result60 ));
  jand g2917(.dina(n2238), .dinb(n485), .dout(n3180));
  jand g2918(.dina(n2246), .dinb(n432), .dout(n3181));
  jor  g2919(.dina(n3181), .dinb(n3180), .dout(n3182));
  jand g2920(.dina(n2227), .dinb(n323), .dout(n3183));
  jand g2921(.dina(n2263), .dinb(n377), .dout(n3184));
  jor  g2922(.dina(n3184), .dinb(n3183), .dout(n3185));
  jor  g2923(.dina(n3185), .dinb(n3182), .dout(n3186));
  jand g2924(.dina(n3186), .dinb(n263), .dout(n3187));
  jand g2925(.dina(n2255), .dinb(n323), .dout(n3188));
  jand g2926(.dina(n2219), .dinb(n377), .dout(n3189));
  jor  g2927(.dina(n3189), .dinb(n3188), .dout(n3190));
  jand g2928(.dina(n2202), .dinb(n432), .dout(n3191));
  jand g2929(.dina(n2210), .dinb(n485), .dout(n3192));
  jor  g2930(.dina(n3192), .dinb(n3191), .dout(n3193));
  jor  g2931(.dina(n3193), .dinb(n3190), .dout(n3194));
  jand g2932(.dina(n3194), .dinb(shift6 ), .dout(n3195));
  jor  g2933(.dina(n3195), .dinb(n3187), .dout(result61 ));
  jand g2934(.dina(n2311), .dinb(n485), .dout(n3197));
  jand g2935(.dina(n2319), .dinb(n432), .dout(n3198));
  jor  g2936(.dina(n3198), .dinb(n3197), .dout(n3199));
  jand g2937(.dina(n2300), .dinb(n323), .dout(n3200));
  jand g2938(.dina(n2336), .dinb(n377), .dout(n3201));
  jor  g2939(.dina(n3201), .dinb(n3200), .dout(n3202));
  jor  g2940(.dina(n3202), .dinb(n3199), .dout(n3203));
  jand g2941(.dina(n3203), .dinb(n263), .dout(n3204));
  jand g2942(.dina(n2328), .dinb(n323), .dout(n3205));
  jand g2943(.dina(n2292), .dinb(n377), .dout(n3206));
  jor  g2944(.dina(n3206), .dinb(n3205), .dout(n3207));
  jand g2945(.dina(n2275), .dinb(n432), .dout(n3208));
  jand g2946(.dina(n2283), .dinb(n485), .dout(n3209));
  jor  g2947(.dina(n3209), .dinb(n3208), .dout(n3210));
  jor  g2948(.dina(n3210), .dinb(n3207), .dout(n3211));
  jand g2949(.dina(n3211), .dinb(shift6 ), .dout(n3212));
  jor  g2950(.dina(n3212), .dinb(n3204), .dout(result62 ));
  jand g2951(.dina(n2384), .dinb(n485), .dout(n3214));
  jand g2952(.dina(n2392), .dinb(n432), .dout(n3215));
  jor  g2953(.dina(n3215), .dinb(n3214), .dout(n3216));
  jand g2954(.dina(n2373), .dinb(n323), .dout(n3217));
  jand g2955(.dina(n2409), .dinb(n377), .dout(n3218));
  jor  g2956(.dina(n3218), .dinb(n3217), .dout(n3219));
  jor  g2957(.dina(n3219), .dinb(n3216), .dout(n3220));
  jand g2958(.dina(n3220), .dinb(n263), .dout(n3221));
  jand g2959(.dina(n2401), .dinb(n323), .dout(n3222));
  jand g2960(.dina(n2365), .dinb(n377), .dout(n3223));
  jor  g2961(.dina(n3223), .dinb(n3222), .dout(n3224));
  jand g2962(.dina(n2348), .dinb(n432), .dout(n3225));
  jand g2963(.dina(n2356), .dinb(n485), .dout(n3226));
  jor  g2964(.dina(n3226), .dinb(n3225), .dout(n3227));
  jor  g2965(.dina(n3227), .dinb(n3224), .dout(n3228));
  jand g2966(.dina(n3228), .dinb(shift6 ), .dout(n3229));
  jor  g2967(.dina(n3229), .dinb(n3221), .dout(result63 ));
  jand g2968(.dina(n698), .dinb(n263), .dout(n3231));
  jand g2969(.dina(n488), .dinb(shift6 ), .dout(n3232));
  jor  g2970(.dina(n3232), .dinb(n3231), .dout(result64 ));
  jand g2971(.dina(n1063), .dinb(n263), .dout(n3234));
  jand g2972(.dina(n879), .dinb(shift6 ), .dout(n3235));
  jor  g2973(.dina(n3235), .dinb(n3234), .dout(result65 ));
  jand g2974(.dina(n1360), .dinb(n263), .dout(n3237));
  jand g2975(.dina(n1212), .dinb(shift6 ), .dout(n3238));
  jor  g2976(.dina(n3238), .dinb(n3237), .dout(result66 ));
  jand g2977(.dina(n1536), .dinb(n263), .dout(n3240));
  jand g2978(.dina(n1445), .dinb(shift6 ), .dout(n3241));
  jor  g2979(.dina(n3241), .dinb(n3240), .dout(result67 ));
  jand g2980(.dina(n1609), .dinb(n263), .dout(n3243));
  jand g2981(.dina(n1573), .dinb(shift6 ), .dout(n3244));
  jor  g2982(.dina(n3244), .dinb(n3243), .dout(result68 ));
  jand g2983(.dina(n1682), .dinb(n263), .dout(n3246));
  jand g2984(.dina(n1646), .dinb(shift6 ), .dout(n3247));
  jor  g2985(.dina(n3247), .dinb(n3246), .dout(result69 ));
  jand g2986(.dina(n1755), .dinb(n263), .dout(n3249));
  jand g2987(.dina(n1719), .dinb(shift6 ), .dout(n3250));
  jor  g2988(.dina(n3250), .dinb(n3249), .dout(result70 ));
  jand g2989(.dina(n1828), .dinb(n263), .dout(n3252));
  jand g2990(.dina(n1792), .dinb(shift6 ), .dout(n3253));
  jor  g2991(.dina(n3253), .dinb(n3252), .dout(result71 ));
  jand g2992(.dina(n1901), .dinb(n263), .dout(n3255));
  jand g2993(.dina(n1865), .dinb(shift6 ), .dout(n3256));
  jor  g2994(.dina(n3256), .dinb(n3255), .dout(result72 ));
  jand g2995(.dina(n1974), .dinb(n263), .dout(n3258));
  jand g2996(.dina(n1938), .dinb(shift6 ), .dout(n3259));
  jor  g2997(.dina(n3259), .dinb(n3258), .dout(result73 ));
  jand g2998(.dina(n2047), .dinb(n263), .dout(n3261));
  jand g2999(.dina(n2011), .dinb(shift6 ), .dout(n3262));
  jor  g3000(.dina(n3262), .dinb(n3261), .dout(result74 ));
  jand g3001(.dina(n2120), .dinb(n263), .dout(n3264));
  jand g3002(.dina(n2084), .dinb(shift6 ), .dout(n3265));
  jor  g3003(.dina(n3265), .dinb(n3264), .dout(result75 ));
  jand g3004(.dina(n2193), .dinb(n263), .dout(n3267));
  jand g3005(.dina(n2157), .dinb(shift6 ), .dout(n3268));
  jor  g3006(.dina(n3268), .dinb(n3267), .dout(result76 ));
  jand g3007(.dina(n2266), .dinb(n263), .dout(n3270));
  jand g3008(.dina(n2230), .dinb(shift6 ), .dout(n3271));
  jor  g3009(.dina(n3271), .dinb(n3270), .dout(result77 ));
  jand g3010(.dina(n2339), .dinb(n263), .dout(n3273));
  jand g3011(.dina(n2303), .dinb(shift6 ), .dout(n3274));
  jor  g3012(.dina(n3274), .dinb(n3273), .dout(result78 ));
  jand g3013(.dina(n2412), .dinb(n263), .dout(n3276));
  jand g3014(.dina(n2376), .dinb(shift6 ), .dout(n3277));
  jor  g3015(.dina(n3277), .dinb(n3276), .dout(result79 ));
  jand g3016(.dina(n2429), .dinb(n263), .dout(n3279));
  jand g3017(.dina(n2421), .dinb(shift6 ), .dout(n3280));
  jor  g3018(.dina(n3280), .dinb(n3279), .dout(result80 ));
  jand g3019(.dina(n2446), .dinb(n263), .dout(n3282));
  jand g3020(.dina(n2438), .dinb(shift6 ), .dout(n3283));
  jor  g3021(.dina(n3283), .dinb(n3282), .dout(result81 ));
  jand g3022(.dina(n2463), .dinb(n263), .dout(n3285));
  jand g3023(.dina(n2455), .dinb(shift6 ), .dout(n3286));
  jor  g3024(.dina(n3286), .dinb(n3285), .dout(result82 ));
  jand g3025(.dina(n2480), .dinb(n263), .dout(n3288));
  jand g3026(.dina(n2472), .dinb(shift6 ), .dout(n3289));
  jor  g3027(.dina(n3289), .dinb(n3288), .dout(result83 ));
  jand g3028(.dina(n2497), .dinb(n263), .dout(n3291));
  jand g3029(.dina(n2489), .dinb(shift6 ), .dout(n3292));
  jor  g3030(.dina(n3292), .dinb(n3291), .dout(result84 ));
  jand g3031(.dina(n2514), .dinb(n263), .dout(n3294));
  jand g3032(.dina(n2506), .dinb(shift6 ), .dout(n3295));
  jor  g3033(.dina(n3295), .dinb(n3294), .dout(result85 ));
  jand g3034(.dina(n2531), .dinb(n263), .dout(n3297));
  jand g3035(.dina(n2523), .dinb(shift6 ), .dout(n3298));
  jor  g3036(.dina(n3298), .dinb(n3297), .dout(result86 ));
  jand g3037(.dina(n2548), .dinb(n263), .dout(n3300));
  jand g3038(.dina(n2540), .dinb(shift6 ), .dout(n3301));
  jor  g3039(.dina(n3301), .dinb(n3300), .dout(result87 ));
  jand g3040(.dina(n2565), .dinb(n263), .dout(n3303));
  jand g3041(.dina(n2557), .dinb(shift6 ), .dout(n3304));
  jor  g3042(.dina(n3304), .dinb(n3303), .dout(result88 ));
  jand g3043(.dina(n2582), .dinb(n263), .dout(n3306));
  jand g3044(.dina(n2574), .dinb(shift6 ), .dout(n3307));
  jor  g3045(.dina(n3307), .dinb(n3306), .dout(result89 ));
  jand g3046(.dina(n2599), .dinb(n263), .dout(n3309));
  jand g3047(.dina(n2591), .dinb(shift6 ), .dout(n3310));
  jor  g3048(.dina(n3310), .dinb(n3309), .dout(result90 ));
  jand g3049(.dina(n2616), .dinb(n263), .dout(n3312));
  jand g3050(.dina(n2608), .dinb(shift6 ), .dout(n3313));
  jor  g3051(.dina(n3313), .dinb(n3312), .dout(result91 ));
  jand g3052(.dina(n2633), .dinb(n263), .dout(n3315));
  jand g3053(.dina(n2625), .dinb(shift6 ), .dout(n3316));
  jor  g3054(.dina(n3316), .dinb(n3315), .dout(result92 ));
  jand g3055(.dina(n2650), .dinb(n263), .dout(n3318));
  jand g3056(.dina(n2642), .dinb(shift6 ), .dout(n3319));
  jor  g3057(.dina(n3319), .dinb(n3318), .dout(result93 ));
  jand g3058(.dina(n2667), .dinb(n263), .dout(n3321));
  jand g3059(.dina(n2659), .dinb(shift6 ), .dout(n3322));
  jor  g3060(.dina(n3322), .dinb(n3321), .dout(result94 ));
  jand g3061(.dina(n2684), .dinb(n263), .dout(n3324));
  jand g3062(.dina(n2676), .dinb(shift6 ), .dout(n3325));
  jor  g3063(.dina(n3325), .dinb(n3324), .dout(result95 ));
  jand g3064(.dina(n2701), .dinb(n263), .dout(n3327));
  jand g3065(.dina(n2693), .dinb(shift6 ), .dout(n3328));
  jor  g3066(.dina(n3328), .dinb(n3327), .dout(result96 ));
  jand g3067(.dina(n2718), .dinb(n263), .dout(n3330));
  jand g3068(.dina(n2710), .dinb(shift6 ), .dout(n3331));
  jor  g3069(.dina(n3331), .dinb(n3330), .dout(result97 ));
  jand g3070(.dina(n2735), .dinb(n263), .dout(n3333));
  jand g3071(.dina(n2727), .dinb(shift6 ), .dout(n3334));
  jor  g3072(.dina(n3334), .dinb(n3333), .dout(result98 ));
  jand g3073(.dina(n2752), .dinb(n263), .dout(n3336));
  jand g3074(.dina(n2744), .dinb(shift6 ), .dout(n3337));
  jor  g3075(.dina(n3337), .dinb(n3336), .dout(result99 ));
  jand g3076(.dina(n2769), .dinb(n263), .dout(n3339));
  jand g3077(.dina(n2761), .dinb(shift6 ), .dout(n3340));
  jor  g3078(.dina(n3340), .dinb(n3339), .dout(result100 ));
  jand g3079(.dina(n2786), .dinb(n263), .dout(n3342));
  jand g3080(.dina(n2778), .dinb(shift6 ), .dout(n3343));
  jor  g3081(.dina(n3343), .dinb(n3342), .dout(result101 ));
  jand g3082(.dina(n2803), .dinb(n263), .dout(n3345));
  jand g3083(.dina(n2795), .dinb(shift6 ), .dout(n3346));
  jor  g3084(.dina(n3346), .dinb(n3345), .dout(result102 ));
  jand g3085(.dina(n2820), .dinb(n263), .dout(n3348));
  jand g3086(.dina(n2812), .dinb(shift6 ), .dout(n3349));
  jor  g3087(.dina(n3349), .dinb(n3348), .dout(result103 ));
  jand g3088(.dina(n2837), .dinb(n263), .dout(n3351));
  jand g3089(.dina(n2829), .dinb(shift6 ), .dout(n3352));
  jor  g3090(.dina(n3352), .dinb(n3351), .dout(result104 ));
  jand g3091(.dina(n2854), .dinb(n263), .dout(n3354));
  jand g3092(.dina(n2846), .dinb(shift6 ), .dout(n3355));
  jor  g3093(.dina(n3355), .dinb(n3354), .dout(result105 ));
  jand g3094(.dina(n2871), .dinb(n263), .dout(n3357));
  jand g3095(.dina(n2863), .dinb(shift6 ), .dout(n3358));
  jor  g3096(.dina(n3358), .dinb(n3357), .dout(result106 ));
  jand g3097(.dina(n2888), .dinb(n263), .dout(n3360));
  jand g3098(.dina(n2880), .dinb(shift6 ), .dout(n3361));
  jor  g3099(.dina(n3361), .dinb(n3360), .dout(result107 ));
  jand g3100(.dina(n2905), .dinb(n263), .dout(n3363));
  jand g3101(.dina(n2897), .dinb(shift6 ), .dout(n3364));
  jor  g3102(.dina(n3364), .dinb(n3363), .dout(result108 ));
  jand g3103(.dina(n2922), .dinb(n263), .dout(n3366));
  jand g3104(.dina(n2914), .dinb(shift6 ), .dout(n3367));
  jor  g3105(.dina(n3367), .dinb(n3366), .dout(result109 ));
  jand g3106(.dina(n2939), .dinb(n263), .dout(n3369));
  jand g3107(.dina(n2931), .dinb(shift6 ), .dout(n3370));
  jor  g3108(.dina(n3370), .dinb(n3369), .dout(result110 ));
  jand g3109(.dina(n2956), .dinb(n263), .dout(n3372));
  jand g3110(.dina(n2948), .dinb(shift6 ), .dout(n3373));
  jor  g3111(.dina(n3373), .dinb(n3372), .dout(result111 ));
  jand g3112(.dina(n2973), .dinb(n263), .dout(n3375));
  jand g3113(.dina(n2965), .dinb(shift6 ), .dout(n3376));
  jor  g3114(.dina(n3376), .dinb(n3375), .dout(result112 ));
  jand g3115(.dina(n2990), .dinb(n263), .dout(n3378));
  jand g3116(.dina(n2982), .dinb(shift6 ), .dout(n3379));
  jor  g3117(.dina(n3379), .dinb(n3378), .dout(result113 ));
  jand g3118(.dina(n3007), .dinb(n263), .dout(n3381));
  jand g3119(.dina(n2999), .dinb(shift6 ), .dout(n3382));
  jor  g3120(.dina(n3382), .dinb(n3381), .dout(result114 ));
  jand g3121(.dina(n3024), .dinb(n263), .dout(n3384));
  jand g3122(.dina(n3016), .dinb(shift6 ), .dout(n3385));
  jor  g3123(.dina(n3385), .dinb(n3384), .dout(result115 ));
  jand g3124(.dina(n3041), .dinb(n263), .dout(n3387));
  jand g3125(.dina(n3033), .dinb(shift6 ), .dout(n3388));
  jor  g3126(.dina(n3388), .dinb(n3387), .dout(result116 ));
  jand g3127(.dina(n3058), .dinb(n263), .dout(n3390));
  jand g3128(.dina(n3050), .dinb(shift6 ), .dout(n3391));
  jor  g3129(.dina(n3391), .dinb(n3390), .dout(result117 ));
  jand g3130(.dina(n3075), .dinb(n263), .dout(n3393));
  jand g3131(.dina(n3067), .dinb(shift6 ), .dout(n3394));
  jor  g3132(.dina(n3394), .dinb(n3393), .dout(result118 ));
  jand g3133(.dina(n3092), .dinb(n263), .dout(n3396));
  jand g3134(.dina(n3084), .dinb(shift6 ), .dout(n3397));
  jor  g3135(.dina(n3397), .dinb(n3396), .dout(result119 ));
  jand g3136(.dina(n3109), .dinb(n263), .dout(n3399));
  jand g3137(.dina(n3101), .dinb(shift6 ), .dout(n3400));
  jor  g3138(.dina(n3400), .dinb(n3399), .dout(result120 ));
  jand g3139(.dina(n3126), .dinb(n263), .dout(n3402));
  jand g3140(.dina(n3118), .dinb(shift6 ), .dout(n3403));
  jor  g3141(.dina(n3403), .dinb(n3402), .dout(result121 ));
  jand g3142(.dina(n3143), .dinb(n263), .dout(n3405));
  jand g3143(.dina(n3135), .dinb(shift6 ), .dout(n3406));
  jor  g3144(.dina(n3406), .dinb(n3405), .dout(result122 ));
  jand g3145(.dina(n3160), .dinb(n263), .dout(n3408));
  jand g3146(.dina(n3152), .dinb(shift6 ), .dout(n3409));
  jor  g3147(.dina(n3409), .dinb(n3408), .dout(result123 ));
  jand g3148(.dina(n3177), .dinb(n263), .dout(n3411));
  jand g3149(.dina(n3169), .dinb(shift6 ), .dout(n3412));
  jor  g3150(.dina(n3412), .dinb(n3411), .dout(result124 ));
  jand g3151(.dina(n3194), .dinb(n263), .dout(n3414));
  jand g3152(.dina(n3186), .dinb(shift6 ), .dout(n3415));
  jor  g3153(.dina(n3415), .dinb(n3414), .dout(result125 ));
  jand g3154(.dina(n3211), .dinb(n263), .dout(n3417));
  jand g3155(.dina(n3203), .dinb(shift6 ), .dout(n3418));
  jor  g3156(.dina(n3418), .dinb(n3417), .dout(result126 ));
  jand g3157(.dina(n3228), .dinb(n263), .dout(n3420));
  jand g3158(.dina(n3220), .dinb(shift6 ), .dout(n3421));
  jor  g3159(.dina(n3421), .dinb(n3420), .dout(result127 ));
endmodule


