/*
gf_c7552:
	jxor: 242
	jspl: 295
	jspl3: 359
	jnot: 215
	jdff: 6368
	jor: 391
	jand: 479

Summary:
	jxor: 242
	jspl: 295
	jspl3: 359
	jnot: 215
	jdff: 6368
	jor: 391
	jand: 479

The maximum logic level gap of any gate:
	gf_c7552: 35
*/

module gf_c7552(gclk, G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526, G4528, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399);
	input gclk;
	input G1;
	input G5;
	input G9;
	input G12;
	input G15;
	input G18;
	input G23;
	input G26;
	input G29;
	input G32;
	input G35;
	input G38;
	input G41;
	input G44;
	input G47;
	input G50;
	input G53;
	input G54;
	input G55;
	input G56;
	input G57;
	input G58;
	input G59;
	input G60;
	input G61;
	input G62;
	input G63;
	input G64;
	input G65;
	input G66;
	input G69;
	input G70;
	input G73;
	input G74;
	input G75;
	input G76;
	input G77;
	input G78;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G84;
	input G85;
	input G86;
	input G87;
	input G88;
	input G89;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G110;
	input G111;
	input G112;
	input G113;
	input G114;
	input G115;
	input G118;
	input G121;
	input G124;
	input G127;
	input G130;
	input G133;
	input G134;
	input G135;
	input G138;
	input G141;
	input G144;
	input G147;
	input G150;
	input G151;
	input G152;
	input G153;
	input G154;
	input G155;
	input G156;
	input G157;
	input G158;
	input G159;
	input G160;
	input G161;
	input G162;
	input G163;
	input G164;
	input G165;
	input G166;
	input G167;
	input G168;
	input G169;
	input G170;
	input G171;
	input G172;
	input G173;
	input G174;
	input G175;
	input G176;
	input G177;
	input G178;
	input G179;
	input G180;
	input G181;
	input G182;
	input G183;
	input G184;
	input G185;
	input G186;
	input G187;
	input G188;
	input G189;
	input G190;
	input G191;
	input G192;
	input G193;
	input G194;
	input G195;
	input G196;
	input G197;
	input G198;
	input G199;
	input G200;
	input G201;
	input G202;
	input G203;
	input G204;
	input G205;
	input G206;
	input G207;
	input G208;
	input G209;
	input G210;
	input G211;
	input G212;
	input G213;
	input G214;
	input G215;
	input G216;
	input G217;
	input G218;
	input G219;
	input G220;
	input G221;
	input G222;
	input G223;
	input G224;
	input G225;
	input G226;
	input G227;
	input G228;
	input G229;
	input G230;
	input G231;
	input G232;
	input G233;
	input G234;
	input G235;
	input G236;
	input G237;
	input G238;
	input G239;
	input G240;
	input G339;
	input G1197;
	input G1455;
	input G1459;
	input G1462;
	input G1469;
	input G1480;
	input G1486;
	input G1492;
	input G1496;
	input G2204;
	input G2208;
	input G2211;
	input G2218;
	input G2224;
	input G2230;
	input G2236;
	input G2239;
	input G2247;
	input G2253;
	input G2256;
	input G3698;
	input G3701;
	input G3705;
	input G3711;
	input G3717;
	input G3723;
	input G3729;
	input G3737;
	input G3743;
	input G3749;
	input G4393;
	input G4394;
	input G4400;
	input G4405;
	input G4410;
	input G4415;
	input G4420;
	input G4427;
	input G4432;
	input G4437;
	input G4526;
	input G4528;
	output G2;
	output G3;
	output G450;
	output G448;
	output G444;
	output G442;
	output G440;
	output G438;
	output G496;
	output G494;
	output G492;
	output G490;
	output G488;
	output G486;
	output G484;
	output G482;
	output G480;
	output G560;
	output G542;
	output G558;
	output G556;
	output G554;
	output G552;
	output G550;
	output G548;
	output G546;
	output G544;
	output G540;
	output G538;
	output G536;
	output G534;
	output G532;
	output G530;
	output G528;
	output G526;
	output G524;
	output G279;
	output G436;
	output G478;
	output G522;
	output G402;
	output G404;
	output G406;
	output G408;
	output G410;
	output G432;
	output G446;
	output G284;
	output G286;
	output G289;
	output G292;
	output G341;
	output G281;
	output G453;
	output G278;
	output G373;
	output G246;
	output G258;
	output G264;
	output G270;
	output G388;
	output G391;
	output G394;
	output G397;
	output G376;
	output G379;
	output G382;
	output G385;
	output G412;
	output G414;
	output G416;
	output G249;
	output G295;
	output G324;
	output G252;
	output G276;
	output G310;
	output G313;
	output G316;
	output G319;
	output G327;
	output G330;
	output G333;
	output G336;
	output G418;
	output G273;
	output G298;
	output G301;
	output G304;
	output G307;
	output G344;
	output G422;
	output G469;
	output G419;
	output G471;
	output G359;
	output G362;
	output G365;
	output G368;
	output G347;
	output G350;
	output G353;
	output G356;
	output G321;
	output G338;
	output G370;
	output G399;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n347;
	wire n348;
	wire n349;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1082;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1102;
	wire n1103;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1356;
	wire n1357;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1384;
	wire n1385;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1399;
	wire n1400;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1413;
	wire n1414;
	wire n1416;
	wire n1417;
	wire n1419;
	wire n1421;
	wire n1423;
	wire n1424;
	wire n1426;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [2:0] w_G5_0;
	wire [1:0] w_G5_1;
	wire [2:0] w_G15_0;
	wire [2:0] w_G18_0;
	wire [2:0] w_G18_1;
	wire [2:0] w_G18_2;
	wire [2:0] w_G18_3;
	wire [2:0] w_G18_4;
	wire [2:0] w_G18_5;
	wire [2:0] w_G18_6;
	wire [2:0] w_G18_7;
	wire [2:0] w_G18_8;
	wire [2:0] w_G18_9;
	wire [2:0] w_G18_10;
	wire [2:0] w_G18_11;
	wire [2:0] w_G18_12;
	wire [2:0] w_G18_13;
	wire [2:0] w_G18_14;
	wire [2:0] w_G18_15;
	wire [2:0] w_G18_16;
	wire [2:0] w_G18_17;
	wire [2:0] w_G18_18;
	wire [2:0] w_G18_19;
	wire [2:0] w_G18_20;
	wire [2:0] w_G18_21;
	wire [2:0] w_G18_22;
	wire [2:0] w_G18_23;
	wire [2:0] w_G18_24;
	wire [2:0] w_G18_25;
	wire [2:0] w_G18_26;
	wire [2:0] w_G18_27;
	wire [2:0] w_G18_28;
	wire [2:0] w_G18_29;
	wire [2:0] w_G18_30;
	wire [2:0] w_G18_31;
	wire [2:0] w_G18_32;
	wire [2:0] w_G18_33;
	wire [2:0] w_G18_34;
	wire [2:0] w_G18_35;
	wire [2:0] w_G18_36;
	wire [2:0] w_G18_37;
	wire [2:0] w_G18_38;
	wire [2:0] w_G18_39;
	wire [2:0] w_G18_40;
	wire [2:0] w_G18_41;
	wire [2:0] w_G18_42;
	wire [2:0] w_G18_43;
	wire [2:0] w_G18_44;
	wire [2:0] w_G18_45;
	wire [2:0] w_G18_46;
	wire [2:0] w_G18_47;
	wire [2:0] w_G18_48;
	wire [2:0] w_G18_49;
	wire [1:0] w_G29_0;
	wire [2:0] w_G38_0;
	wire [2:0] w_G38_1;
	wire [2:0] w_G38_2;
	wire [1:0] w_G41_0;
	wire [1:0] w_G70_0;
	wire [1:0] w_G89_0;
	wire [2:0] w_G106_0;
	wire [1:0] w_G106_1;
	wire [1:0] w_G209_0;
	wire [1:0] w_G238_0;
	wire [2:0] w_G1455_0;
	wire [1:0] w_G1459_0;
	wire [1:0] w_G1462_0;
	wire [1:0] w_G1469_0;
	wire [2:0] w_G1480_0;
	wire [1:0] w_G1486_0;
	wire [2:0] w_G1492_0;
	wire [1:0] w_G1492_1;
	wire [2:0] w_G1496_0;
	wire [1:0] w_G1496_1;
	wire [2:0] w_G2204_0;
	wire [1:0] w_G2208_0;
	wire [2:0] w_G2211_0;
	wire [2:0] w_G2218_0;
	wire [2:0] w_G2224_0;
	wire [1:0] w_G2224_1;
	wire [2:0] w_G2230_0;
	wire [2:0] w_G2236_0;
	wire [2:0] w_G2239_0;
	wire [1:0] w_G2239_1;
	wire [2:0] w_G2247_0;
	wire [2:0] w_G2253_0;
	wire [1:0] w_G2256_0;
	wire [1:0] w_G3698_0;
	wire [2:0] w_G3701_0;
	wire [1:0] w_G3701_1;
	wire [2:0] w_G3705_0;
	wire [2:0] w_G3705_1;
	wire [1:0] w_G3711_0;
	wire [2:0] w_G3717_0;
	wire [2:0] w_G3723_0;
	wire [2:0] w_G3729_0;
	wire [1:0] w_G3729_1;
	wire [2:0] w_G3737_0;
	wire [2:0] w_G3743_0;
	wire [2:0] w_G3749_0;
	wire [1:0] w_G4393_0;
	wire [2:0] w_G4394_0;
	wire [1:0] w_G4394_1;
	wire [2:0] w_G4400_0;
	wire [1:0] w_G4400_1;
	wire [2:0] w_G4405_0;
	wire [1:0] w_G4405_1;
	wire [2:0] w_G4410_0;
	wire [2:0] w_G4415_0;
	wire [1:0] w_G4415_1;
	wire [2:0] w_G4420_0;
	wire [1:0] w_G4420_1;
	wire [2:0] w_G4427_0;
	wire [2:0] w_G4432_0;
	wire [2:0] w_G4437_0;
	wire [2:0] w_G4526_0;
	wire [2:0] w_G4526_1;
	wire [2:0] w_G4526_2;
	wire [2:0] w_G4528_0;
	wire w_G404_0;
	wire G404_fa_;
	wire w_G406_0;
	wire G406_fa_;
	wire w_G408_0;
	wire G408_fa_;
	wire w_G410_0;
	wire G410_fa_;
	wire w_G412_0;
	wire G412_fa_;
	wire w_G414_0;
	wire G414_fa_;
	wire w_G416_0;
	wire G416_fa_;
	wire w_G252_0;
	wire G252_fa_;
	wire [1:0] w_n345_0;
	wire [1:0] w_n347_0;
	wire [1:0] w_n349_0;
	wire [1:0] w_n353_0;
	wire [2:0] w_n354_0;
	wire [2:0] w_n355_0;
	wire [2:0] w_n355_1;
	wire [2:0] w_n355_2;
	wire [2:0] w_n355_3;
	wire [2:0] w_n355_4;
	wire [2:0] w_n355_5;
	wire [2:0] w_n355_6;
	wire [2:0] w_n355_7;
	wire [2:0] w_n355_8;
	wire [2:0] w_n355_9;
	wire [2:0] w_n355_10;
	wire [2:0] w_n355_11;
	wire [2:0] w_n355_12;
	wire [2:0] w_n355_13;
	wire [2:0] w_n355_14;
	wire [2:0] w_n355_15;
	wire [2:0] w_n355_16;
	wire [2:0] w_n355_17;
	wire [2:0] w_n355_18;
	wire [2:0] w_n355_19;
	wire [2:0] w_n355_20;
	wire [2:0] w_n355_21;
	wire [2:0] w_n355_22;
	wire [2:0] w_n355_23;
	wire [2:0] w_n355_24;
	wire [2:0] w_n355_25;
	wire [2:0] w_n355_26;
	wire [2:0] w_n355_27;
	wire [2:0] w_n355_28;
	wire [2:0] w_n355_29;
	wire [2:0] w_n355_30;
	wire [2:0] w_n355_31;
	wire [2:0] w_n355_32;
	wire [2:0] w_n355_33;
	wire [2:0] w_n355_34;
	wire [2:0] w_n355_35;
	wire [1:0] w_n357_0;
	wire [1:0] w_n358_0;
	wire [2:0] w_n359_0;
	wire [1:0] w_n359_1;
	wire [2:0] w_n361_0;
	wire [2:0] w_n362_0;
	wire [2:0] w_n363_0;
	wire [2:0] w_n364_0;
	wire [2:0] w_n366_0;
	wire [1:0] w_n367_0;
	wire [1:0] w_n368_0;
	wire [1:0] w_n369_0;
	wire [2:0] w_n370_0;
	wire [2:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [2:0] w_n373_0;
	wire [2:0] w_n373_1;
	wire [2:0] w_n373_2;
	wire [2:0] w_n373_3;
	wire [2:0] w_n373_4;
	wire [2:0] w_n373_5;
	wire [2:0] w_n373_6;
	wire [2:0] w_n373_7;
	wire [2:0] w_n373_8;
	wire [2:0] w_n373_9;
	wire [1:0] w_n374_0;
	wire [2:0] w_n375_0;
	wire [2:0] w_n377_0;
	wire [2:0] w_n377_1;
	wire [1:0] w_n378_0;
	wire [2:0] w_n379_0;
	wire [1:0] w_n380_0;
	wire [2:0] w_n383_0;
	wire [1:0] w_n385_0;
	wire [1:0] w_n386_0;
	wire [2:0] w_n387_0;
	wire [1:0] w_n387_1;
	wire [2:0] w_n388_0;
	wire [2:0] w_n388_1;
	wire [2:0] w_n389_0;
	wire [1:0] w_n389_1;
	wire [2:0] w_n391_0;
	wire [2:0] w_n392_0;
	wire [2:0] w_n393_0;
	wire [1:0] w_n393_1;
	wire [1:0] w_n394_0;
	wire [2:0] w_n395_0;
	wire [1:0] w_n395_1;
	wire [2:0] w_n396_0;
	wire [2:0] w_n396_1;
	wire [1:0] w_n397_0;
	wire [2:0] w_n405_0;
	wire [1:0] w_n407_0;
	wire [2:0] w_n409_0;
	wire [1:0] w_n409_1;
	wire [2:0] w_n411_0;
	wire [1:0] w_n411_1;
	wire [2:0] w_n413_0;
	wire [1:0] w_n413_1;
	wire [2:0] w_n414_0;
	wire [1:0] w_n414_1;
	wire [1:0] w_n415_0;
	wire [2:0] w_n416_0;
	wire [1:0] w_n418_0;
	wire [1:0] w_n419_0;
	wire [1:0] w_n420_0;
	wire [2:0] w_n421_0;
	wire [1:0] w_n422_0;
	wire [2:0] w_n423_0;
	wire [1:0] w_n424_0;
	wire [2:0] w_n425_0;
	wire [1:0] w_n425_1;
	wire [2:0] w_n426_0;
	wire [1:0] w_n427_0;
	wire [2:0] w_n428_0;
	wire [2:0] w_n429_0;
	wire [1:0] w_n430_0;
	wire [1:0] w_n431_0;
	wire [2:0] w_n432_0;
	wire [2:0] w_n433_0;
	wire [2:0] w_n433_1;
	wire [1:0] w_n434_0;
	wire [1:0] w_n435_0;
	wire [2:0] w_n436_0;
	wire [2:0] w_n437_0;
	wire [1:0] w_n438_0;
	wire [1:0] w_n440_0;
	wire [2:0] w_n444_0;
	wire [2:0] w_n445_0;
	wire [2:0] w_n447_0;
	wire [2:0] w_n449_0;
	wire [1:0] w_n449_1;
	wire [2:0] w_n450_0;
	wire [2:0] w_n451_0;
	wire [2:0] w_n453_0;
	wire [1:0] w_n453_1;
	wire [2:0] w_n456_0;
	wire [1:0] w_n457_0;
	wire [2:0] w_n459_0;
	wire [2:0] w_n460_0;
	wire [2:0] w_n460_1;
	wire [2:0] w_n462_0;
	wire [2:0] w_n463_0;
	wire [1:0] w_n463_1;
	wire [2:0] w_n464_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n466_0;
	wire [1:0] w_n467_0;
	wire [2:0] w_n469_0;
	wire [1:0] w_n469_1;
	wire [2:0] w_n470_0;
	wire [2:0] w_n471_0;
	wire [1:0] w_n472_0;
	wire [2:0] w_n474_0;
	wire [2:0] w_n475_0;
	wire [2:0] w_n476_0;
	wire [1:0] w_n477_0;
	wire [2:0] w_n479_0;
	wire [1:0] w_n479_1;
	wire [2:0] w_n480_0;
	wire [1:0] w_n480_1;
	wire [1:0] w_n481_0;
	wire [1:0] w_n485_0;
	wire [1:0] w_n486_0;
	wire [2:0] w_n487_0;
	wire [2:0] w_n489_0;
	wire [2:0] w_n491_0;
	wire [1:0] w_n491_1;
	wire [2:0] w_n495_0;
	wire [1:0] w_n495_1;
	wire [2:0] w_n496_0;
	wire [2:0] w_n497_0;
	wire [1:0] w_n497_1;
	wire [1:0] w_n499_0;
	wire [1:0] w_n500_0;
	wire [2:0] w_n501_0;
	wire [1:0] w_n503_0;
	wire [2:0] w_n504_0;
	wire [1:0] w_n504_1;
	wire [1:0] w_n505_0;
	wire [1:0] w_n507_0;
	wire [2:0] w_n509_0;
	wire [1:0] w_n511_0;
	wire [2:0] w_n512_0;
	wire [2:0] w_n513_0;
	wire [1:0] w_n513_1;
	wire [1:0] w_n514_0;
	wire [1:0] w_n516_0;
	wire [2:0] w_n517_0;
	wire [1:0] w_n517_1;
	wire [2:0] w_n518_0;
	wire [2:0] w_n518_1;
	wire [1:0] w_n520_0;
	wire [1:0] w_n522_0;
	wire [2:0] w_n523_0;
	wire [2:0] w_n524_0;
	wire [2:0] w_n524_1;
	wire [2:0] w_n526_0;
	wire [1:0] w_n528_0;
	wire [1:0] w_n530_0;
	wire [2:0] w_n531_0;
	wire [1:0] w_n531_1;
	wire [2:0] w_n536_0;
	wire [1:0] w_n538_0;
	wire [2:0] w_n539_0;
	wire [1:0] w_n539_1;
	wire [1:0] w_n544_0;
	wire [1:0] w_n546_0;
	wire [2:0] w_n547_0;
	wire [1:0] w_n547_1;
	wire [1:0] w_n548_0;
	wire [1:0] w_n550_0;
	wire [1:0] w_n552_0;
	wire [1:0] w_n554_0;
	wire [2:0] w_n555_0;
	wire [1:0] w_n555_1;
	wire [2:0] w_n556_0;
	wire [1:0] w_n558_0;
	wire [1:0] w_n560_0;
	wire [1:0] w_n562_0;
	wire [2:0] w_n563_0;
	wire [1:0] w_n563_1;
	wire [2:0] w_n564_0;
	wire [1:0] w_n565_0;
	wire [2:0] w_n566_0;
	wire [2:0] w_n568_0;
	wire [2:0] w_n570_0;
	wire [2:0] w_n570_1;
	wire [2:0] w_n572_0;
	wire [1:0] w_n572_1;
	wire [2:0] w_n573_0;
	wire [1:0] w_n573_1;
	wire [2:0] w_n574_0;
	wire [2:0] w_n575_0;
	wire [1:0] w_n575_1;
	wire [2:0] w_n576_0;
	wire [1:0] w_n577_0;
	wire [2:0] w_n578_0;
	wire [2:0] w_n580_0;
	wire [2:0] w_n581_0;
	wire [2:0] w_n582_0;
	wire [1:0] w_n584_0;
	wire [2:0] w_n585_0;
	wire [1:0] w_n585_1;
	wire [2:0] w_n586_0;
	wire [1:0] w_n588_0;
	wire [2:0] w_n590_0;
	wire [1:0] w_n592_0;
	wire [2:0] w_n593_0;
	wire [1:0] w_n593_1;
	wire [2:0] w_n594_0;
	wire [2:0] w_n595_0;
	wire [1:0] w_n597_0;
	wire [2:0] w_n598_0;
	wire [1:0] w_n598_1;
	wire [2:0] w_n599_0;
	wire [1:0] w_n600_0;
	wire [1:0] w_n602_0;
	wire [2:0] w_n603_0;
	wire [1:0] w_n603_1;
	wire [1:0] w_n604_0;
	wire [2:0] w_n605_0;
	wire [1:0] w_n609_0;
	wire [1:0] w_n610_0;
	wire [1:0] w_n612_0;
	wire [2:0] w_n613_0;
	wire [2:0] w_n615_0;
	wire [1:0] w_n616_0;
	wire [2:0] w_n618_0;
	wire [2:0] w_n619_0;
	wire [2:0] w_n622_0;
	wire [1:0] w_n624_0;
	wire [2:0] w_n625_0;
	wire [1:0] w_n625_1;
	wire [2:0] w_n626_0;
	wire [1:0] w_n626_1;
	wire [2:0] w_n627_0;
	wire [1:0] w_n629_0;
	wire [2:0] w_n630_0;
	wire [2:0] w_n631_0;
	wire [2:0] w_n632_0;
	wire [1:0] w_n632_1;
	wire [1:0] w_n634_0;
	wire [2:0] w_n635_0;
	wire [1:0] w_n635_1;
	wire [2:0] w_n636_0;
	wire [2:0] w_n641_0;
	wire [2:0] w_n642_0;
	wire [1:0] w_n644_0;
	wire [1:0] w_n645_0;
	wire [1:0] w_n646_0;
	wire [1:0] w_n647_0;
	wire [1:0] w_n649_0;
	wire [1:0] w_n651_0;
	wire [1:0] w_n652_0;
	wire [1:0] w_n653_0;
	wire [2:0] w_n654_0;
	wire [1:0] w_n655_0;
	wire [1:0] w_n656_0;
	wire [2:0] w_n657_0;
	wire [1:0] w_n659_0;
	wire [2:0] w_n660_0;
	wire [2:0] w_n661_0;
	wire [1:0] w_n662_0;
	wire [2:0] w_n663_0;
	wire [1:0] w_n663_1;
	wire [1:0] w_n664_0;
	wire [1:0] w_n666_0;
	wire [1:0] w_n669_0;
	wire [1:0] w_n671_0;
	wire [2:0] w_n673_0;
	wire [1:0] w_n674_0;
	wire [2:0] w_n676_0;
	wire [1:0] w_n678_0;
	wire [2:0] w_n680_0;
	wire [2:0] w_n680_1;
	wire [2:0] w_n680_2;
	wire [1:0] w_n682_0;
	wire [1:0] w_n683_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n689_0;
	wire [1:0] w_n690_0;
	wire [1:0] w_n693_0;
	wire [1:0] w_n694_0;
	wire [1:0] w_n695_0;
	wire [1:0] w_n696_0;
	wire [1:0] w_n698_0;
	wire [2:0] w_n700_0;
	wire [1:0] w_n700_1;
	wire [2:0] w_n703_0;
	wire [2:0] w_n703_1;
	wire [1:0] w_n705_0;
	wire [2:0] w_n707_0;
	wire [2:0] w_n707_1;
	wire [2:0] w_n709_0;
	wire [1:0] w_n709_1;
	wire [2:0] w_n711_0;
	wire [1:0] w_n711_1;
	wire [2:0] w_n712_0;
	wire [1:0] w_n713_0;
	wire [2:0] w_n715_0;
	wire [1:0] w_n715_1;
	wire [2:0] w_n718_0;
	wire [1:0] w_n719_0;
	wire [2:0] w_n720_0;
	wire [2:0] w_n723_0;
	wire [1:0] w_n724_0;
	wire [1:0] w_n725_0;
	wire [2:0] w_n726_0;
	wire [1:0] w_n726_1;
	wire [2:0] w_n729_0;
	wire [1:0] w_n729_1;
	wire [2:0] w_n734_0;
	wire [1:0] w_n736_0;
	wire [2:0] w_n737_0;
	wire [1:0] w_n737_1;
	wire [2:0] w_n741_0;
	wire [1:0] w_n741_1;
	wire [1:0] w_n743_0;
	wire [2:0] w_n744_0;
	wire [2:0] w_n747_0;
	wire [1:0] w_n749_0;
	wire [1:0] w_n754_0;
	wire [2:0] w_n755_0;
	wire [1:0] w_n755_1;
	wire [2:0] w_n758_0;
	wire [1:0] w_n758_1;
	wire [1:0] w_n760_0;
	wire [2:0] w_n761_0;
	wire [2:0] w_n764_0;
	wire [1:0] w_n766_0;
	wire [1:0] w_n767_0;
	wire [2:0] w_n768_0;
	wire [2:0] w_n772_0;
	wire [1:0] w_n773_0;
	wire [1:0] w_n774_0;
	wire [1:0] w_n775_0;
	wire [2:0] w_n776_0;
	wire [2:0] w_n780_0;
	wire [1:0] w_n781_0;
	wire [2:0] w_n796_0;
	wire [1:0] w_n796_1;
	wire [2:0] w_n800_0;
	wire [1:0] w_n800_1;
	wire [2:0] w_n803_0;
	wire [2:0] w_n806_0;
	wire [1:0] w_n808_0;
	wire [2:0] w_n810_0;
	wire [1:0] w_n810_1;
	wire [2:0] w_n814_0;
	wire [1:0] w_n814_1;
	wire [2:0] w_n817_0;
	wire [2:0] w_n820_0;
	wire [1:0] w_n822_0;
	wire [2:0] w_n824_0;
	wire [2:0] w_n827_0;
	wire [2:0] w_n845_0;
	wire [1:0] w_n845_1;
	wire [2:0] w_n848_0;
	wire [1:0] w_n848_1;
	wire [2:0] w_n851_0;
	wire [2:0] w_n854_0;
	wire [1:0] w_n856_0;
	wire [2:0] w_n858_0;
	wire [2:0] w_n862_0;
	wire [1:0] w_n863_0;
	wire [1:0] w_n864_0;
	wire [2:0] w_n866_0;
	wire [2:0] w_n870_0;
	wire [1:0] w_n871_0;
	wire [2:0] w_n885_0;
	wire [2:0] w_n888_0;
	wire [2:0] w_n891_0;
	wire [2:0] w_n894_0;
	wire [1:0] w_n895_0;
	wire [2:0] w_n900_0;
	wire [2:0] w_n903_0;
	wire [1:0] w_n905_0;
	wire [2:0] w_n916_0;
	wire [2:0] w_n919_0;
	wire [2:0] w_n926_0;
	wire [2:0] w_n930_0;
	wire [2:0] w_n935_0;
	wire [2:0] w_n938_0;
	wire [2:0] w_n944_0;
	wire [2:0] w_n947_0;
	wire [2:0] w_n950_0;
	wire [1:0] w_n950_1;
	wire [2:0] w_n953_0;
	wire [1:0] w_n953_1;
	wire [2:0] w_n966_0;
	wire [2:0] w_n970_0;
	wire [2:0] w_n973_0;
	wire [1:0] w_n973_1;
	wire [2:0] w_n977_0;
	wire [1:0] w_n977_1;
	wire [2:0] w_n980_0;
	wire [2:0] w_n983_0;
	wire [1:0] w_n985_0;
	wire [2:0] w_n987_0;
	wire [2:0] w_n991_0;
	wire [1:0] w_n992_0;
	wire [2:0] w_n995_0;
	wire [2:0] w_n999_0;
	wire [1:0] w_n1000_0;
	wire [1:0] w_n1003_0;
	wire [1:0] w_n1007_0;
	wire [1:0] w_n1008_0;
	wire [1:0] w_n1042_0;
	wire [2:0] w_n1059_0;
	wire [2:0] w_n1067_0;
	wire [2:0] w_n1069_0;
	wire [1:0] w_n1070_0;
	wire [1:0] w_n1073_0;
	wire [1:0] w_n1078_0;
	wire [2:0] w_n1084_0;
	wire [1:0] w_n1086_0;
	wire [1:0] w_n1090_0;
	wire [2:0] w_n1092_0;
	wire [2:0] w_n1094_0;
	wire [1:0] w_n1096_0;
	wire [1:0] w_n1099_0;
	wire [1:0] w_n1105_0;
	wire [1:0] w_n1106_0;
	wire [1:0] w_n1108_0;
	wire [1:0] w_n1113_0;
	wire [1:0] w_n1118_0;
	wire [1:0] w_n1127_0;
	wire [1:0] w_n1137_0;
	wire [1:0] w_n1150_0;
	wire [1:0] w_n1172_0;
	wire [1:0] w_n1307_0;
	wire [1:0] w_n1308_0;
	wire [1:0] w_n1309_0;
	wire [1:0] w_n1310_0;
	wire [2:0] w_n1312_0;
	wire [1:0] w_n1312_1;
	wire [1:0] w_n1316_0;
	wire [1:0] w_n1317_0;
	wire [2:0] w_n1321_0;
	wire [1:0] w_n1321_1;
	wire [1:0] w_n1323_0;
	wire [1:0] w_n1333_0;
	wire [2:0] w_n1337_0;
	wire [1:0] w_n1337_1;
	wire [2:0] w_n1340_0;
	wire [1:0] w_n1343_0;
	wire [1:0] w_n1344_0;
	wire [1:0] w_n1359_0;
	wire [1:0] w_n1364_0;
	wire [1:0] w_n1369_0;
	wire [1:0] w_n1370_0;
	wire [1:0] w_n1372_0;
	wire [1:0] w_n1387_0;
	wire [1:0] w_n1388_0;
	wire [1:0] w_n1396_0;
	wire [1:0] w_n1402_0;
	wire [1:0] w_n1408_0;
	wire [1:0] w_n1419_0;
	wire [1:0] w_n1426_0;
	wire [1:0] w_n1431_0;
	wire [1:0] w_n1433_0;
	wire [1:0] w_n1440_0;
	wire [2:0] w_n1452_0;
	wire [1:0] w_n1458_0;
	wire [1:0] w_n1486_0;
	wire [1:0] w_n1492_0;
	wire [1:0] w_n1506_0;
	wire [1:0] w_n1511_0;
	wire [1:0] w_n1518_0;
	wire [1:0] w_n1529_0;
	wire [1:0] w_n1531_0;
	wire [1:0] w_n1534_0;
	wire [1:0] w_n1536_0;
	wire [1:0] w_n1543_0;
	wire [1:0] w_n1554_0;
	wire [2:0] w_n1562_0;
	wire [1:0] w_n1587_0;
	wire [1:0] w_n1597_0;
	wire [1:0] w_n1605_0;
	wire [1:0] w_n1607_0;
	wire [1:0] w_n1610_0;
	wire [1:0] w_n1620_0;
	wire [1:0] w_n1624_0;
	wire w_dff_A_n9g5SFgC7_0;
	wire w_dff_A_7au7tv7s7_1;
	wire w_dff_A_QQzWuTYo3_2;
	wire w_dff_B_eVb1uE7h3_2;
	wire w_dff_B_QW2NFVLj0_0;
	wire w_dff_B_iv2qALu13_1;
	wire w_dff_B_JL3Uxk8f4_1;
	wire w_dff_B_nVkUxcQh2_1;
	wire w_dff_B_dZFVaLSq9_1;
	wire w_dff_B_bxUYwUlW2_1;
	wire w_dff_B_rFvENq0u8_1;
	wire w_dff_B_hlzU7xKp9_1;
	wire w_dff_B_crLpbJdd3_1;
	wire w_dff_B_7ugGyDHY8_1;
	wire w_dff_B_aM0y4fTl0_1;
	wire w_dff_B_oKopyVDu0_1;
	wire w_dff_B_VzZUjfJJ3_1;
	wire w_dff_B_LysNLlf65_1;
	wire w_dff_B_ZSK9EZ2f6_1;
	wire w_dff_B_w359KRXJ1_1;
	wire w_dff_B_QDqV3Viq0_1;
	wire w_dff_B_izIiGylm2_1;
	wire w_dff_B_BQCItuAB9_1;
	wire w_dff_B_8HFHMBLa2_0;
	wire w_dff_B_Fh2BoDEf2_0;
	wire w_dff_B_LVM4weCC0_0;
	wire w_dff_B_gW8CMy1h9_0;
	wire w_dff_B_cxf56XXI2_0;
	wire w_dff_B_EALYBs6j4_0;
	wire w_dff_B_RfPtmtFx6_0;
	wire w_dff_B_HNUnMUZf5_0;
	wire w_dff_B_3yh1LDUD9_0;
	wire w_dff_B_rPsERgDg4_0;
	wire w_dff_B_6aWEYUU27_0;
	wire w_dff_B_2gyqvWcx3_0;
	wire w_dff_B_OJFaf4C45_0;
	wire w_dff_B_agc9kbSX2_0;
	wire w_dff_B_QhklNHYJ1_0;
	wire w_dff_B_4OlEFcVr6_0;
	wire w_dff_B_UWyCibH59_1;
	wire w_dff_B_8JBo7MtE0_1;
	wire w_dff_B_2JDqAnWF6_1;
	wire w_dff_B_PNmrDce39_1;
	wire w_dff_B_aLZtl6TB0_1;
	wire w_dff_B_PVYmZCkK3_1;
	wire w_dff_B_rhWpG1sa2_1;
	wire w_dff_B_LOovrd8T7_1;
	wire w_dff_B_gMtGkkf78_1;
	wire w_dff_B_Xgr1Rhsw9_0;
	wire w_dff_B_QB02PcLq1_0;
	wire w_dff_B_oatz0fpB2_0;
	wire w_dff_B_XQf3rFE19_0;
	wire w_dff_B_vxvH3OFK4_0;
	wire w_dff_B_GrPooNUC1_0;
	wire w_dff_B_OfgiU85C0_0;
	wire w_dff_B_qPumAjg09_0;
	wire w_dff_B_V0LyciSs5_0;
	wire w_dff_B_Ka3Cw3Gj3_0;
	wire w_dff_B_BJYVUQtv6_0;
	wire w_dff_B_GSjd4Lz08_0;
	wire w_dff_B_OQGKkDLd6_0;
	wire w_dff_B_uRaaM5jN4_0;
	wire w_dff_B_Q0RK8VJb7_0;
	wire w_dff_B_RtWilZ243_0;
	wire w_dff_B_g3X5V15h0_0;
	wire w_dff_B_nKOYJWaS6_1;
	wire w_dff_B_akVBs4rW7_1;
	wire w_dff_A_etnL63KJ2_0;
	wire w_dff_B_2PwnoF0C9_1;
	wire w_dff_B_BGoAAQot9_1;
	wire w_dff_B_mjwidCI77_1;
	wire w_dff_B_V9nMdID11_1;
	wire w_dff_B_tYdbC80R0_1;
	wire w_dff_B_TH4u9rLa8_1;
	wire w_dff_B_lAxSjQ1s9_1;
	wire w_dff_B_5FUHYWFc4_1;
	wire w_dff_B_En9U1VzK2_1;
	wire w_dff_B_N2JrJOuG9_1;
	wire w_dff_B_BlWityMK6_1;
	wire w_dff_B_jwk2BptA6_1;
	wire w_dff_B_zPqGfzw23_1;
	wire w_dff_B_RbCkI6so9_1;
	wire w_dff_B_q2ed6MJC2_1;
	wire w_dff_B_3dj0ESMk7_1;
	wire w_dff_B_Ly1Pwmrj8_1;
	wire w_dff_B_b8V7jSAR0_1;
	wire w_dff_B_ISYftX5M2_1;
	wire w_dff_B_OJlOckdU6_1;
	wire w_dff_B_3UocEI9x1_1;
	wire w_dff_B_Zltogmk66_1;
	wire w_dff_B_aGNbQitz5_1;
	wire w_dff_B_tGTEbQFu9_1;
	wire w_dff_B_t4PbNbjN9_1;
	wire w_dff_B_k4zYkSZL1_1;
	wire w_dff_B_pQAnTvFN7_1;
	wire w_dff_B_o6SHvsb31_1;
	wire w_dff_B_17DmmvCM8_1;
	wire w_dff_B_gbMbJoQG1_1;
	wire w_dff_B_CFcAvKLj6_0;
	wire w_dff_B_rQbrq56t8_0;
	wire w_dff_B_HmzUSUyA1_0;
	wire w_dff_B_QXc6b5cQ2_0;
	wire w_dff_B_X0FCGtHk4_0;
	wire w_dff_B_PRKVWczS3_0;
	wire w_dff_B_FDHQqxPH7_0;
	wire w_dff_B_CdpEen625_0;
	wire w_dff_B_h5sEIVQ94_0;
	wire w_dff_B_hIYWDFIz8_0;
	wire w_dff_B_JQlIRtgm7_0;
	wire w_dff_B_dHo87xgk2_0;
	wire w_dff_B_1QSc33RG0_0;
	wire w_dff_B_DWOeTdVH9_0;
	wire w_dff_B_A988JWCx6_0;
	wire w_dff_B_Wrw5Hqd19_0;
	wire w_dff_B_udaqWIxX2_1;
	wire w_dff_B_UtZYf41y7_1;
	wire w_dff_B_SnWwyTbr1_1;
	wire w_dff_B_DeBSnkJO1_1;
	wire w_dff_B_Ibq7IEn14_1;
	wire w_dff_B_V5letM908_1;
	wire w_dff_B_xZ4Xqwaj8_1;
	wire w_dff_B_DR71AT8P1_1;
	wire w_dff_B_1HW4sbfE6_1;
	wire w_dff_B_hqillBlo1_1;
	wire w_dff_B_jilyhg740_1;
	wire w_dff_B_kU0byQFR8_1;
	wire w_dff_B_Sx1uNu5a3_1;
	wire w_dff_B_dZGAQpab0_1;
	wire w_dff_B_xLdrZaIi8_1;
	wire w_dff_B_JqCmj6pN7_1;
	wire w_dff_B_4Wuzp8db7_1;
	wire w_dff_B_wZtY4F0h6_1;
	wire w_dff_B_LWD6H3D95_1;
	wire w_dff_B_FyyDFzm21_1;
	wire w_dff_B_hSbRrYUw8_1;
	wire w_dff_B_UAu2N2p05_1;
	wire w_dff_B_hDBXXTch2_1;
	wire w_dff_B_6ZZMi8gg9_1;
	wire w_dff_B_bp3JTHAO6_0;
	wire w_dff_B_VOa6mjkz4_0;
	wire w_dff_B_obl5F4as6_0;
	wire w_dff_B_gcpaaMQq6_0;
	wire w_dff_B_C5z9MrMH0_0;
	wire w_dff_B_F25zxsnW1_0;
	wire w_dff_B_xfLNtrgX0_0;
	wire w_dff_B_hNdKFqWY8_0;
	wire w_dff_B_w78BfbYk0_0;
	wire w_dff_B_IN28J2OI0_0;
	wire w_dff_B_g0IXKYU45_0;
	wire w_dff_B_4iCGeQns8_0;
	wire w_dff_B_Cz8YghvD9_0;
	wire w_dff_B_cuMzDEww9_0;
	wire w_dff_B_1fYsCXVZ7_0;
	wire w_dff_B_RuudyVQP2_0;
	wire w_dff_B_ZkmYrJx73_1;
	wire w_dff_B_fNbtVY718_1;
	wire w_dff_B_PkOzYPwq0_0;
	wire w_dff_A_ZGaBYqMV5_1;
	wire w_dff_A_K0UyC9ij2_1;
	wire w_dff_B_7UnKPXbe2_0;
	wire w_dff_B_AysCa2sL2_1;
	wire w_dff_A_hL4QtHdo2_1;
	wire w_dff_B_9uMlF7Ay0_2;
	wire w_dff_B_tsEoyIJd7_1;
	wire w_dff_B_dobygOqp2_1;
	wire w_dff_B_TSRR2EAS2_1;
	wire w_dff_B_br1cFjSc2_1;
	wire w_dff_B_m7N8lvTH8_1;
	wire w_dff_B_XLCg4Vxz6_1;
	wire w_dff_A_Jl51lhWb4_1;
	wire w_dff_A_YFJq84cV2_1;
	wire w_dff_A_UCuGhZcJ5_1;
	wire w_dff_A_lttAXzVh7_1;
	wire w_dff_B_wyZkRwqg1_3;
	wire w_dff_B_WFFcg9b19_3;
	wire w_dff_B_GjJNepL59_3;
	wire w_dff_B_3Y7CzIhi9_3;
	wire w_dff_B_5FjumPSY2_3;
	wire w_dff_B_lnJSQtNq1_3;
	wire w_dff_B_VYBVRL0s7_3;
	wire w_dff_B_cshPhwWY7_3;
	wire w_dff_B_fAR5PAi63_3;
	wire w_dff_B_Tstrbp4H5_3;
	wire w_dff_B_gwZrCtHh3_3;
	wire w_dff_B_ecySOCm87_3;
	wire w_dff_B_rYNRIiR07_3;
	wire w_dff_B_KfHtvRn50_3;
	wire w_dff_B_AnFO0cLV7_3;
	wire w_dff_B_qLiOIZ6E7_3;
	wire w_dff_B_36q99d5L1_3;
	wire w_dff_B_jN5ZtIgq2_3;
	wire w_dff_B_Z4txTq0q7_3;
	wire w_dff_B_CNLUHhKi7_3;
	wire w_dff_B_iTjKjlLP6_3;
	wire w_dff_B_NWmhIE741_3;
	wire w_dff_B_moekdsPF3_3;
	wire w_dff_B_47SaYpgW2_3;
	wire w_dff_B_Xp7qq0Vb4_0;
	wire w_dff_B_XwvYcmZv1_1;
	wire w_dff_B_1KBvtN5y0_1;
	wire w_dff_B_Z1MCnMhS5_1;
	wire w_dff_B_8p0wyfGX5_1;
	wire w_dff_B_BTItQeXr3_1;
	wire w_dff_B_GcJ6Qs3N9_1;
	wire w_dff_B_F2Ipz71k2_1;
	wire w_dff_B_Dnilearv7_1;
	wire w_dff_B_GanduZdd6_1;
	wire w_dff_B_OL0A4bTl4_1;
	wire w_dff_B_vEEIB46e3_1;
	wire w_dff_B_lxQHE9iJ3_1;
	wire w_dff_B_YGEwG3Zv8_1;
	wire w_dff_B_oZNzsOXp5_1;
	wire w_dff_B_PzZ9sjmD6_1;
	wire w_dff_B_jDmQfozV5_1;
	wire w_dff_B_OQxyPvgY5_1;
	wire w_dff_B_HZJ6luck2_1;
	wire w_dff_B_iu6b9rUm6_1;
	wire w_dff_B_kEcfKRZY5_1;
	wire w_dff_B_nnbLFFhQ7_1;
	wire w_dff_B_ypHWpTQ32_1;
	wire w_dff_B_LxQ2xTZx8_1;
	wire w_dff_B_6sAumDgf3_1;
	wire w_dff_B_kfwgKews0_1;
	wire w_dff_B_7Dn82H1x6_1;
	wire w_dff_B_jStP1M7t8_1;
	wire w_dff_B_tOhu7D1u7_1;
	wire w_dff_B_Mag9w8OI4_1;
	wire w_dff_B_ZdJKHoFX8_1;
	wire w_dff_B_lx5nZqAc0_1;
	wire w_dff_B_Oo0QY9Ih6_1;
	wire w_dff_B_QJBBCxc72_1;
	wire w_dff_B_ttWn3OQ39_1;
	wire w_dff_B_7TZ60Xwn9_1;
	wire w_dff_B_ZgiK9XAF4_1;
	wire w_dff_B_Plyq66uC2_1;
	wire w_dff_B_uNYCFD427_1;
	wire w_dff_B_P2UJUTcZ8_1;
	wire w_dff_B_YTkSdiyG8_1;
	wire w_dff_B_hoqQbiCM6_1;
	wire w_dff_B_8Nz34Ps88_0;
	wire w_dff_B_RF3upjcN2_0;
	wire w_dff_B_JB2wzUzL0_0;
	wire w_dff_B_sQ5WW1bI7_0;
	wire w_dff_B_Cwm1zvf69_0;
	wire w_dff_B_kKSLLmd88_0;
	wire w_dff_B_lh8VyK5u1_0;
	wire w_dff_B_B2omcMka9_0;
	wire w_dff_B_23Ep1ycX0_0;
	wire w_dff_B_otYfyN7k6_0;
	wire w_dff_B_mFzj0fnV1_0;
	wire w_dff_B_JQsr2JeB4_0;
	wire w_dff_B_QNMsegxi0_1;
	wire w_dff_B_PNhe6DRF0_1;
	wire w_dff_B_AwPlcsak5_1;
	wire w_dff_B_jorYkMEJ4_1;
	wire w_dff_B_Hhr9qj9p0_0;
	wire w_dff_B_fKc0yDPw9_0;
	wire w_dff_B_bLFA0pqD5_1;
	wire w_dff_B_vETxS4Ly4_0;
	wire w_dff_B_1vllwRkt2_0;
	wire w_dff_B_4bXAa7Qs8_0;
	wire w_dff_B_Z2MGMkkr8_1;
	wire w_dff_B_e3nt4qMF6_1;
	wire w_dff_B_34isNXdR2_1;
	wire w_dff_B_3JTNGUfp6_1;
	wire w_dff_B_iSDLFJwX9_1;
	wire w_dff_B_ge5PWEz40_0;
	wire w_dff_B_ZDcraaM70_0;
	wire w_dff_B_HgrYxgY77_0;
	wire w_dff_A_wbodIdqm6_0;
	wire w_dff_A_EAfLFRDE2_0;
	wire w_dff_A_ZZF8lVze4_0;
	wire w_dff_A_A4sJ5E0u2_0;
	wire w_dff_B_Ah2aUiDQ3_1;
	wire w_dff_A_ezWMIB7q9_0;
	wire w_dff_A_N3BsIWX12_1;
	wire w_dff_A_RhqxIhuS9_1;
	wire w_dff_B_83cBPOSs0_2;
	wire w_dff_B_sdDMOuXZ9_0;
	wire w_dff_B_LEgRd1n37_0;
	wire w_dff_B_P0OTCDOI4_0;
	wire w_dff_B_zkNYjj430_0;
	wire w_dff_B_tnYWgAfx1_0;
	wire w_dff_B_uZ9L45DT7_0;
	wire w_dff_B_orv1wjnb3_1;
	wire w_dff_B_CNN3Tmiw0_0;
	wire w_dff_B_4kWLMhoZ9_0;
	wire w_dff_B_xFBDYDCS7_0;
	wire w_dff_B_JdUiZGCi0_0;
	wire w_dff_B_3bJApQEN4_0;
	wire w_dff_B_estVN0us2_0;
	wire w_dff_B_NehKFbxp0_0;
	wire w_dff_B_9iZzCCub3_0;
	wire w_dff_B_CidzbUxa3_0;
	wire w_dff_B_MapM6INs9_0;
	wire w_dff_B_BppfZCnu1_0;
	wire w_dff_B_Nz54HwJD5_0;
	wire w_dff_B_ID7XDYqu7_0;
	wire w_dff_B_DwOjqOiE3_0;
	wire w_dff_B_k180PTCX8_0;
	wire w_dff_B_gxkXCOrE5_0;
	wire w_dff_B_zxf4LBxI1_0;
	wire w_dff_B_nggOTCOy9_0;
	wire w_dff_B_bo2wYj5S3_1;
	wire w_dff_B_q6EnlDxl3_1;
	wire w_dff_B_ZauRDTiH8_1;
	wire w_dff_B_wRFYCBmU5_0;
	wire w_dff_B_1SRk8rnZ7_0;
	wire w_dff_B_RnXkE3it4_0;
	wire w_dff_B_BNFVeHPN2_0;
	wire w_dff_A_ZZDYvtpd2_0;
	wire w_dff_A_fwEvooYQ0_0;
	wire w_dff_B_xCGAEQP75_0;
	wire w_dff_B_R2ssDfRx2_1;
	wire w_dff_A_Ig6Jd2UU0_1;
	wire w_dff_A_RuXzwzZo6_1;
	wire w_dff_B_s5Hp0cC17_1;
	wire w_dff_B_y6tAviAl7_1;
	wire w_dff_B_eQadKVK99_1;
	wire w_dff_B_QOmj15Uf4_1;
	wire w_dff_B_c06RZygx3_1;
	wire w_dff_B_sjOvuJzq8_1;
	wire w_dff_B_OaYYyJIi8_1;
	wire w_dff_B_YYagu3qC3_1;
	wire w_dff_B_PNEekTyH5_1;
	wire w_dff_B_fUtICkG03_1;
	wire w_dff_B_NQhm448A5_1;
	wire w_dff_B_26CUA39Z9_1;
	wire w_dff_B_tnretszl7_1;
	wire w_dff_B_YnwHMZT42_1;
	wire w_dff_B_sfp0FJc35_1;
	wire w_dff_B_j8VXcBKN6_1;
	wire w_dff_B_b2IvIusC6_1;
	wire w_dff_B_PAWkJtJY9_1;
	wire w_dff_B_v8NiatIJ7_1;
	wire w_dff_B_j67HeSxg9_1;
	wire w_dff_B_rk62XQu75_1;
	wire w_dff_B_Yyae2c6K8_1;
	wire w_dff_B_PzBMoEd49_1;
	wire w_dff_B_IPsu51sy8_1;
	wire w_dff_B_YCx18kfC2_1;
	wire w_dff_B_EBsTKoK00_1;
	wire w_dff_B_Biz1UDPJ3_1;
	wire w_dff_B_5rz7YNcP1_1;
	wire w_dff_B_veDgjCRN8_1;
	wire w_dff_B_LlzMOLUu9_1;
	wire w_dff_B_jKGlioYE1_1;
	wire w_dff_B_r3vDdZ8X0_1;
	wire w_dff_B_3AZH8EsJ1_1;
	wire w_dff_B_TIhj8ilP0_1;
	wire w_dff_B_zAuZVIdH9_1;
	wire w_dff_B_mHSbwIWC5_1;
	wire w_dff_B_r0Yh98b39_1;
	wire w_dff_B_lEZTA7sg4_1;
	wire w_dff_B_Ib8tCxxr1_1;
	wire w_dff_B_YW26d8oN5_1;
	wire w_dff_B_gtvralSJ4_1;
	wire w_dff_B_50cW6R5h5_1;
	wire w_dff_B_9vv4BaAl1_1;
	wire w_dff_B_lT7YcpLB1_1;
	wire w_dff_B_RDORgMqD4_1;
	wire w_dff_B_ALJ4lXBz2_1;
	wire w_dff_B_LX7CG5Qt4_1;
	wire w_dff_B_LZwkqAo59_1;
	wire w_dff_B_1DLfnPfQ1_1;
	wire w_dff_B_EcLzNYaP2_1;
	wire w_dff_B_5DVjiJ859_1;
	wire w_dff_B_97LKRyJs4_1;
	wire w_dff_B_hy9CQt7z0_1;
	wire w_dff_B_JDntq90E5_1;
	wire w_dff_B_Vk81izGt4_1;
	wire w_dff_B_ahLpG0yz2_2;
	wire w_dff_B_A8Ubha8d9_2;
	wire w_dff_B_Pfp9khLw3_2;
	wire w_dff_B_JRXQ9fNn1_2;
	wire w_dff_B_IIjiu3Bv2_2;
	wire w_dff_B_oLXc25eD2_2;
	wire w_dff_B_HiNlUkE01_2;
	wire w_dff_B_wsUnivT46_2;
	wire w_dff_B_fsDYXqJj3_2;
	wire w_dff_B_cLBQPQYd8_2;
	wire w_dff_B_6NYEkpyw4_2;
	wire w_dff_B_Xzmf6IqD8_2;
	wire w_dff_B_YNLKOk187_2;
	wire w_dff_B_eQvRwRHh1_2;
	wire w_dff_B_LlkwaQ854_2;
	wire w_dff_B_ofEo3QIb5_2;
	wire w_dff_B_sOpolSFo4_2;
	wire w_dff_B_sqbqov2b6_2;
	wire w_dff_B_zQFllWNM0_2;
	wire w_dff_B_cRySGfZj1_2;
	wire w_dff_B_x3F9zCXM5_2;
	wire w_dff_B_Iwz6rXXn2_2;
	wire w_dff_B_2wAmErmz5_2;
	wire w_dff_B_nPlACwd95_2;
	wire w_dff_B_FfWgKOYy4_2;
	wire w_dff_B_1ul6ytrd7_2;
	wire w_dff_B_C7pro73t8_2;
	wire w_dff_B_xetpYuPs7_2;
	wire w_dff_B_eapPgTTJ3_2;
	wire w_dff_B_Nsi5X4a68_2;
	wire w_dff_B_Bh2we42W7_2;
	wire w_dff_B_ZQeZ26oA8_2;
	wire w_dff_B_XFy51k1n4_2;
	wire w_dff_B_0Ktn2SDL8_2;
	wire w_dff_B_V0recqrJ1_2;
	wire w_dff_B_3cYDWd4q5_2;
	wire w_dff_B_cCwouaHD3_2;
	wire w_dff_B_zOLsnwPo4_2;
	wire w_dff_B_TW8d3bdG2_2;
	wire w_dff_B_ZAW1SaQB6_2;
	wire w_dff_B_XL2DLYm64_2;
	wire w_dff_B_vOkVqBPd0_2;
	wire w_dff_B_N2PZ3a1Q0_2;
	wire w_dff_B_SH94kbda1_2;
	wire w_dff_B_4a0rIBNL6_2;
	wire w_dff_B_Gor3mNL25_2;
	wire w_dff_B_7vaA25NE1_2;
	wire w_dff_B_0YPyJ8Uc4_2;
	wire w_dff_B_aXUwLWky9_2;
	wire w_dff_B_2eIhZ2w12_2;
	wire w_dff_B_C4w7ZstR7_2;
	wire w_dff_B_JjtbViYg2_2;
	wire w_dff_B_vGWTtvqL1_2;
	wire w_dff_B_7ZadreeO3_2;
	wire w_dff_B_agoTf6pK2_2;
	wire w_dff_B_lCJ7p6YX6_2;
	wire w_dff_B_rqPDnjiC8_2;
	wire w_dff_B_vuxAlKJW3_2;
	wire w_dff_B_gm6zH1U62_2;
	wire w_dff_B_rYSpOFRW4_2;
	wire w_dff_B_nnIPsxnx3_1;
	wire w_dff_B_oJ3uk5Yu9_1;
	wire w_dff_B_5GBMW2tW7_1;
	wire w_dff_B_SQrA1Ldx3_1;
	wire w_dff_B_QfoNWJZa1_1;
	wire w_dff_B_jZ1VNd3j9_1;
	wire w_dff_B_zbpEuFZc3_1;
	wire w_dff_B_6neiXGcZ2_1;
	wire w_dff_B_WsznJuhN4_1;
	wire w_dff_B_D3ju29x52_1;
	wire w_dff_B_NRiDnaVs1_0;
	wire w_dff_B_xYAtRbtz9_0;
	wire w_dff_B_0P283q1G0_0;
	wire w_dff_B_DwLSuusb8_0;
	wire w_dff_B_e5eFDp330_0;
	wire w_dff_B_qNU6KT989_0;
	wire w_dff_B_hU40mBNJ5_0;
	wire w_dff_B_rfMi1FXX7_0;
	wire w_dff_B_nYIWO4Zh3_0;
	wire w_dff_B_qZ37TkEr6_0;
	wire w_dff_B_iO12gpId8_1;
	wire w_dff_B_hETOkRjX2_0;
	wire w_dff_B_7CjXRu199_1;
	wire w_dff_B_MEpDpiEk0_1;
	wire w_dff_B_jhQ9ZwHH8_1;
	wire w_dff_B_r4wVXBmI4_1;
	wire w_dff_B_ElLWtjbo3_1;
	wire w_dff_B_yxh4zwZu0_0;
	wire w_dff_B_DruvH7gb4_0;
	wire w_dff_B_VqDCOUdL7_0;
	wire w_dff_B_T8lypvRC0_0;
	wire w_dff_B_L7MDHylB8_1;
	wire w_dff_B_gX7dCrmQ4_0;
	wire w_dff_B_8KC414ka4_1;
	wire w_dff_B_oSRhgFo17_1;
	wire w_dff_B_cxn5ESvY5_1;
	wire w_dff_B_31ztlG9W9_1;
	wire w_dff_B_LCvwGGe99_0;
	wire w_dff_B_jXbhs1Ts2_0;
	wire w_dff_B_gg1Pz5RC7_0;
	wire w_dff_B_dxTagTcf8_0;
	wire w_dff_B_8NSQiVkX4_1;
	wire w_dff_B_pwJz712V9_1;
	wire w_dff_B_9OoVwt040_0;
	wire w_dff_B_78xqVym44_0;
	wire w_dff_B_VCPo7aj54_0;
	wire w_dff_B_HI17SWLs1_0;
	wire w_dff_B_xlnYYd9P9_0;
	wire w_dff_B_rilexsIN7_0;
	wire w_dff_B_ACptuE0V4_0;
	wire w_dff_B_lVJBxmwj6_0;
	wire w_dff_B_8afCptDr6_0;
	wire w_dff_B_neYfZjv58_0;
	wire w_dff_A_dvAMxUoN8_0;
	wire w_dff_B_XobirX4R6_0;
	wire w_dff_B_bqA7wn954_1;
	wire w_dff_B_wiIQHOaU6_1;
	wire w_dff_B_bWgIHx2K6_1;
	wire w_dff_B_yr36TW4i6_1;
	wire w_dff_B_9B07w0IG3_1;
	wire w_dff_A_kPtUaf2H8_0;
	wire w_dff_A_PpFG70SJ1_0;
	wire w_dff_B_X6BYXpZV8_0;
	wire w_dff_A_kCiJr1094_0;
	wire w_dff_A_2hx7wOQO9_0;
	wire w_dff_B_LdDA1UfB9_0;
	wire w_dff_B_q4LyJ9mr1_0;
	wire w_dff_A_8Cb6vKBt0_2;
	wire w_dff_B_IC7aNWb99_0;
	wire w_dff_B_4OUwLuKY1_1;
	wire w_dff_B_9v9MOOrH2_1;
	wire w_dff_B_mVGGaIz23_0;
	wire w_dff_A_9BgNPRCU5_1;
	wire w_dff_B_mTocefGd9_0;
	wire w_dff_B_lnZwKp530_0;
	wire w_dff_B_CwWHlkEl2_0;
	wire w_dff_B_fT6cpS2r5_0;
	wire w_dff_B_NfZNRfxe8_0;
	wire w_dff_B_fFR3xlQT2_0;
	wire w_dff_B_XXe0m7kV4_0;
	wire w_dff_B_cQLPEVoP8_0;
	wire w_dff_B_dnkm3fBP6_0;
	wire w_dff_B_fV89OfNc8_0;
	wire w_dff_B_g6xz6nVJ6_0;
	wire w_dff_B_bxk0bZM88_0;
	wire w_dff_B_MxQHdMvy2_0;
	wire w_dff_B_ZKWIEJTp2_0;
	wire w_dff_B_9SokRwpu0_0;
	wire w_dff_B_9bgLBXQJ9_0;
	wire w_dff_B_Jrk5eOK59_0;
	wire w_dff_B_1rrGnPMp2_0;
	wire w_dff_B_5YrEWmCa8_0;
	wire w_dff_B_4nTjbmam1_0;
	wire w_dff_B_tC5oChiN6_0;
	wire w_dff_B_q9i22s8O9_0;
	wire w_dff_A_ZFgUO11s5_0;
	wire w_dff_B_4s9IArk87_0;
	wire w_dff_A_ERBY7ag16_0;
	wire w_dff_B_gRr2QMWX6_1;
	wire w_dff_B_Y00uvtA76_1;
	wire w_dff_B_VaOgOo7R7_0;
	wire w_dff_B_FIx2mURg1_0;
	wire w_dff_B_U8wghQvY4_0;
	wire w_dff_B_KVIsyAul7_0;
	wire w_dff_B_oVCXBg7B5_0;
	wire w_dff_B_PknzMfj32_0;
	wire w_dff_B_suekqKZF4_0;
	wire w_dff_A_Cid0r0AO1_0;
	wire w_dff_A_RIAEFIVh8_2;
	wire w_dff_A_1ikDeAhx6_2;
	wire w_dff_B_UT7DX8AU3_1;
	wire w_dff_B_mmKU2qf88_1;
	wire w_dff_B_hIfhACI74_0;
	wire w_dff_A_HQPL7rNf1_0;
	wire w_dff_B_lmDZK8E89_0;
	wire w_dff_B_VAnidCBK9_1;
	wire w_dff_A_t7Tf8XrA0_1;
	wire w_dff_B_8rIQAGib9_0;
	wire w_dff_B_UQfx4r7m6_0;
	wire w_dff_B_l3G4sekk1_0;
	wire w_dff_B_i1Wnk4No1_0;
	wire w_dff_B_sQF7XcW14_0;
	wire w_dff_B_VMN7qhTg7_0;
	wire w_dff_B_bTJoSfQD1_0;
	wire w_dff_B_LWRHO66N8_1;
	wire w_dff_A_6HllCUn99_0;
	wire w_dff_B_DjGqyaxc6_0;
	wire w_dff_B_GVGkWjOU8_0;
	wire w_dff_A_rNjZUdEz4_0;
	wire w_dff_B_erXJUqiE4_0;
	wire w_dff_B_jCyB9P0P2_0;
	wire w_dff_B_LTj0zE0V5_0;
	wire w_dff_B_6S7kVID85_0;
	wire w_dff_B_bEl0xenY5_0;
	wire w_dff_B_K8YkDxMJ7_0;
	wire w_dff_B_kX1qkxWd0_0;
	wire w_dff_B_ZDQVdoiT8_0;
	wire w_dff_B_6S4NPvSl2_0;
	wire w_dff_B_hZpeGKhD7_0;
	wire w_dff_B_LlYTllIS2_0;
	wire w_dff_B_aJMHWVVK0_0;
	wire w_dff_B_IHKWq1ZS2_0;
	wire w_dff_B_Q1fKgDge9_0;
	wire w_dff_B_eweljXyV3_0;
	wire w_dff_B_motdm5k38_0;
	wire w_dff_B_NXZo4Vpb7_0;
	wire w_dff_A_RwjGpHMx3_0;
	wire w_dff_B_MevoUuZj5_0;
	wire w_dff_B_rZiy9hkI1_0;
	wire w_dff_B_7harNJMF0_3;
	wire w_dff_B_8OB2MLuA2_3;
	wire w_dff_B_YnPVhjWc0_3;
	wire w_dff_B_eu4nILTo8_3;
	wire w_dff_B_Vk2AVHSq9_3;
	wire w_dff_B_LJJj8OGw5_3;
	wire w_dff_B_HIa3BgOe6_3;
	wire w_dff_B_JgJYS9W98_3;
	wire w_dff_B_ESPycNKz5_3;
	wire w_dff_B_yWHsUTY29_3;
	wire w_dff_B_0gzNXEkO3_3;
	wire w_dff_B_VvcJRpKe3_3;
	wire w_dff_B_Pf0PwEVi3_3;
	wire w_dff_B_WPCQJIqE3_3;
	wire w_dff_B_58YVGJTN1_3;
	wire w_dff_B_MdRPCVhl7_3;
	wire w_dff_B_Oew8zBW70_3;
	wire w_dff_B_w0Mvhv1d9_3;
	wire w_dff_B_c8js4H3A1_3;
	wire w_dff_B_MBpvApYr2_3;
	wire w_dff_B_6rziHhf50_3;
	wire w_dff_B_YeNXfyw63_3;
	wire w_dff_B_yOSJnDMg0_3;
	wire w_dff_B_U4aXV4h35_3;
	wire w_dff_B_qEa75UDU2_3;
	wire w_dff_B_GVWJ8yq63_3;
	wire w_dff_B_zSMpWHB00_3;
	wire w_dff_B_v4tQL05P7_3;
	wire w_dff_B_Jl9eAITO4_3;
	wire w_dff_B_E0sjvPnC4_3;
	wire w_dff_B_jz4mq0wf2_3;
	wire w_dff_B_htuktq9e4_3;
	wire w_dff_B_cHzQtCIR4_3;
	wire w_dff_B_jHOlOr462_3;
	wire w_dff_B_ZQL03hyj8_0;
	wire w_dff_B_twlXeJ7q4_1;
	wire w_dff_B_XtVTCOOT6_1;
	wire w_dff_B_0ajKQru93_1;
	wire w_dff_B_mObBsoMl9_1;
	wire w_dff_B_5NRuV43X0_1;
	wire w_dff_B_T6QZYIjE6_1;
	wire w_dff_B_z2e1mNPa3_1;
	wire w_dff_B_JDGzKElI0_1;
	wire w_dff_B_jZweMMIS4_1;
	wire w_dff_B_rmHqHeNi5_1;
	wire w_dff_B_tkqYSXQp0_1;
	wire w_dff_B_JyJLMoj38_1;
	wire w_dff_B_NOccPzQb0_1;
	wire w_dff_B_h6faLEoc9_1;
	wire w_dff_B_DpojqN0o5_1;
	wire w_dff_B_PERSpz908_1;
	wire w_dff_B_Lpz9wFYH3_1;
	wire w_dff_B_iBF0zSIX9_1;
	wire w_dff_B_yEufKW7X7_1;
	wire w_dff_B_fq0e9X9X7_1;
	wire w_dff_B_FJr2wMqf2_1;
	wire w_dff_B_03xCJqGp8_1;
	wire w_dff_B_sVVjQfj48_1;
	wire w_dff_B_BKunGsue7_1;
	wire w_dff_B_8R73yoEh1_1;
	wire w_dff_B_qjyl5HXG2_1;
	wire w_dff_B_7EXr7k8h9_1;
	wire w_dff_B_0IJlOyoJ7_1;
	wire w_dff_B_sUkka6jM2_1;
	wire w_dff_B_RSrplJz97_1;
	wire w_dff_B_q3iB6P8T0_1;
	wire w_dff_B_gBVPGCjC2_1;
	wire w_dff_B_PO5zx7vC7_1;
	wire w_dff_B_5a4TbPj14_1;
	wire w_dff_A_HBTyAc6I7_0;
	wire w_dff_A_eMHmEffM2_0;
	wire w_dff_A_5RNSaOsB4_0;
	wire w_dff_A_7QrLGILF0_0;
	wire w_dff_A_UqDAvpNu7_0;
	wire w_dff_A_08piZveL4_0;
	wire w_dff_A_GLjZCPGx4_0;
	wire w_dff_A_dGsttuS78_0;
	wire w_dff_A_R3LwgNdi5_0;
	wire w_dff_A_z2ZIgc8r4_0;
	wire w_dff_A_DYkcfs9h4_0;
	wire w_dff_A_9ULzOk1L2_0;
	wire w_dff_A_a9dCG73h6_0;
	wire w_dff_A_V3cVFiR18_0;
	wire w_dff_A_xwI6hixk2_0;
	wire w_dff_A_83rLeqmB9_0;
	wire w_dff_A_XXUM6CNb9_0;
	wire w_dff_A_5zaQv1Fu1_0;
	wire w_dff_A_migGWQ6K0_0;
	wire w_dff_A_lbXWVGxB4_0;
	wire w_dff_A_uo4fPLGn1_0;
	wire w_dff_A_9v7X2MgY2_0;
	wire w_dff_A_zh8uifpR5_0;
	wire w_dff_A_XDFsk4m49_0;
	wire w_dff_A_t8tGgAvN9_0;
	wire w_dff_A_IvULAnd04_0;
	wire w_dff_A_5inUDP0s4_0;
	wire w_dff_A_lDbIQf1M1_0;
	wire w_dff_A_TLi6Ey8p3_0;
	wire w_dff_A_C4WFfANq9_0;
	wire w_dff_A_UID0nzDd2_0;
	wire w_dff_A_brOidayp1_0;
	wire w_dff_A_1NxDNOAD3_0;
	wire w_dff_A_wVLQgSOY1_0;
	wire w_dff_A_ihZcVA6G5_1;
	wire w_dff_A_BHKCSiIk4_0;
	wire w_dff_A_2FSUKeD00_0;
	wire w_dff_A_cEOHc9J08_1;
	wire w_dff_A_ehSBP0Yb4_1;
	wire w_dff_B_q0LQ1LIh0_3;
	wire w_dff_B_E7JCIvke2_3;
	wire w_dff_B_wMLwoEFJ5_3;
	wire w_dff_B_FFS9hwVn0_3;
	wire w_dff_B_Gj4y2JOc4_3;
	wire w_dff_B_6PjPud009_3;
	wire w_dff_B_0Zy8qH1L9_3;
	wire w_dff_B_mHJbPJ679_3;
	wire w_dff_B_tBka5SwJ4_3;
	wire w_dff_B_DdEpOIuM5_3;
	wire w_dff_B_RerjznoS2_3;
	wire w_dff_B_6iBaV3qT7_3;
	wire w_dff_B_y2IhB3Wx2_3;
	wire w_dff_B_JFyCRsdG0_3;
	wire w_dff_B_KuS2jGWu0_3;
	wire w_dff_B_xuvGn3c46_3;
	wire w_dff_B_pc5SgHtI1_3;
	wire w_dff_B_xUOIYxBN4_3;
	wire w_dff_B_DVHmYXEY2_3;
	wire w_dff_B_vEQQW6vH5_3;
	wire w_dff_B_0TcigI3U1_3;
	wire w_dff_B_AlUWaXrM6_3;
	wire w_dff_B_UJ55DKDV2_3;
	wire w_dff_B_adZOlTAc3_3;
	wire w_dff_B_ZtTqyoaC8_3;
	wire w_dff_B_IIYzzFNh4_3;
	wire w_dff_B_XKCGeKdu6_3;
	wire w_dff_B_xIIADPOF8_3;
	wire w_dff_B_pKKk1fqI5_3;
	wire w_dff_B_3UxzEWLV4_3;
	wire w_dff_B_otunNgPD3_3;
	wire w_dff_B_nxbVmBxn9_3;
	wire w_dff_B_gPMZX7B71_1;
	wire w_dff_A_DpxLS1m19_2;
	wire w_dff_B_Uq11c23E3_3;
	wire w_dff_B_QhcL4qzt4_3;
	wire w_dff_B_1mfOWhPf0_3;
	wire w_dff_B_Rosh9z2W5_3;
	wire w_dff_B_LvtAVJsN0_3;
	wire w_dff_B_3RjnZiL48_3;
	wire w_dff_B_rPE1qjcr5_3;
	wire w_dff_B_a8fbWRL04_3;
	wire w_dff_B_epQU5li38_3;
	wire w_dff_B_FeAzPCQL2_3;
	wire w_dff_B_ZLhaZyTj5_3;
	wire w_dff_B_UOMizGQl3_3;
	wire w_dff_B_Zf7VFlvj9_3;
	wire w_dff_B_PlUhUOXm0_3;
	wire w_dff_B_7fTbE3Qs0_3;
	wire w_dff_B_140LrTg14_3;
	wire w_dff_B_meu9KNNh7_3;
	wire w_dff_B_MlF8rQDI4_3;
	wire w_dff_B_p1VP9w0V4_3;
	wire w_dff_B_laQWJH2k2_3;
	wire w_dff_B_nh8BRbDh6_3;
	wire w_dff_B_VLp3duVg2_3;
	wire w_dff_B_jIgyEFNl8_3;
	wire w_dff_B_LO4dsblm8_3;
	wire w_dff_B_ofiOtxJx9_3;
	wire w_dff_B_12GJp60D6_3;
	wire w_dff_B_tCs5qjH55_3;
	wire w_dff_B_FlfoBxZO6_3;
	wire w_dff_B_et4NPvVk8_3;
	wire w_dff_B_85JHcCmn5_3;
	wire w_dff_B_8iLpfF7G6_3;
	wire w_dff_B_93hIVo6c5_3;
	wire w_dff_B_GwLzA4Vi2_3;
	wire w_dff_B_ICQHecuV9_3;
	wire w_dff_B_wWZk4Lds0_1;
	wire w_dff_B_wJv8Z09L0_1;
	wire w_dff_B_KGtdqV2A3_1;
	wire w_dff_B_5tREL57K7_1;
	wire w_dff_B_RF5t2aVj9_1;
	wire w_dff_B_WcJaMcar2_1;
	wire w_dff_B_LQia12gc9_1;
	wire w_dff_B_feOQWGXI5_0;
	wire w_dff_B_9nxREcP01_0;
	wire w_dff_B_GBOVEWZc9_0;
	wire w_dff_B_yZhpUOE74_0;
	wire w_dff_B_q5H8wVDo8_0;
	wire w_dff_B_4SapPi330_0;
	wire w_dff_B_qSPEZmw36_0;
	wire w_dff_B_PKJyVjaC7_0;
	wire w_dff_B_1pLUySZd3_0;
	wire w_dff_B_qZd0qqtg9_0;
	wire w_dff_B_zb3Fl8IE9_0;
	wire w_dff_B_nBniW0zQ0_0;
	wire w_dff_B_oQY7Vf4N0_0;
	wire w_dff_B_hvJq30dk8_0;
	wire w_dff_B_NDmSaG2h9_0;
	wire w_dff_B_9Ijh9dG00_0;
	wire w_dff_B_TK2VkFiS0_0;
	wire w_dff_B_12HAZl668_0;
	wire w_dff_B_oSPfDfeT1_0;
	wire w_dff_B_3A12Cw1k7_0;
	wire w_dff_B_1NZYUUDW3_0;
	wire w_dff_B_DxnJ7JMd7_0;
	wire w_dff_B_ruU84gPK4_0;
	wire w_dff_B_D5dEVWu88_0;
	wire w_dff_B_8vozDF7V2_0;
	wire w_dff_B_5qcoIMpU2_0;
	wire w_dff_B_Ca4LTnJZ4_0;
	wire w_dff_B_gIhRgRjM1_0;
	wire w_dff_B_Zt8ILZVx8_0;
	wire w_dff_B_gUUhPHdx0_0;
	wire w_dff_B_mhhPRSfj5_0;
	wire w_dff_B_x2Z9RvSJ7_0;
	wire w_dff_B_ElOjTrJk8_0;
	wire w_dff_B_6a3XpskK7_0;
	wire w_dff_B_bLwZTJWi7_0;
	wire w_dff_B_OUDgAJoO4_0;
	wire w_dff_B_rwukpntz1_0;
	wire w_dff_B_9FbwB4DN9_0;
	wire w_dff_B_4EJ33MHl7_0;
	wire w_dff_B_reTKQ3Mt8_0;
	wire w_dff_B_GQZn4cF11_0;
	wire w_dff_B_AXN5zYGA4_0;
	wire w_dff_B_2738FR838_0;
	wire w_dff_B_mQA7HCfO5_0;
	wire w_dff_B_8fkx1HXv7_0;
	wire w_dff_B_HGeN4flO9_0;
	wire w_dff_B_u2t1JI6M1_0;
	wire w_dff_B_Jbq6DmhX3_0;
	wire w_dff_B_rqNvkiyT5_0;
	wire w_dff_B_80hPncZ95_0;
	wire w_dff_B_S7F6LStF1_0;
	wire w_dff_B_BRMmmpfL0_0;
	wire w_dff_B_nRPVgKWW5_0;
	wire w_dff_B_8kAVW8gB0_0;
	wire w_dff_B_GmWRTMoa6_0;
	wire w_dff_B_d4kiu3Y44_0;
	wire w_dff_B_GfyjoT731_0;
	wire w_dff_B_hephm8TV5_0;
	wire w_dff_B_mxWw4cXU4_0;
	wire w_dff_B_JFGY0C2l5_0;
	wire w_dff_B_ACIfsFgv6_0;
	wire w_dff_B_oAbW667H2_0;
	wire w_dff_B_Rsfrln7j2_0;
	wire w_dff_B_8IkfZdUQ2_0;
	wire w_dff_B_jZ7TKH3V2_0;
	wire w_dff_B_ICu2GORB2_0;
	wire w_dff_B_dNevHoGM4_0;
	wire w_dff_B_W25aDOCw2_0;
	wire w_dff_B_uJpGYrPR3_0;
	wire w_dff_B_7mnuJ1KH0_0;
	wire w_dff_B_s4mshVr45_0;
	wire w_dff_B_INOpmN2v9_0;
	wire w_dff_B_PL1JEJ9U9_1;
	wire w_dff_B_1FyWNS501_0;
	wire w_dff_B_NozrAiAC0_0;
	wire w_dff_B_b9b3rXR82_0;
	wire w_dff_B_KYND4Y7A2_0;
	wire w_dff_B_ew9BjGEv2_1;
	wire w_dff_B_8MmWqEbC1_1;
	wire w_dff_B_yv0IKcgm6_0;
	wire w_dff_B_N2OCdIRW9_0;
	wire w_dff_B_xpKKAL3M3_0;
	wire w_dff_B_lc2rTYBf5_0;
	wire w_dff_A_719EER1D0_0;
	wire w_dff_A_OjBgAxHs3_0;
	wire w_dff_A_W0PFkf9e6_0;
	wire w_dff_A_TtsvZyKe2_0;
	wire w_dff_A_gbJB54ha2_2;
	wire w_dff_A_PzrwB98c9_2;
	wire w_dff_A_7oZDXmlx4_2;
	wire w_dff_A_krkk7XAh3_1;
	wire w_dff_A_aBj6fkYF0_2;
	wire w_dff_A_2zKwrxka1_2;
	wire w_dff_A_HUrhjDSj0_2;
	wire w_dff_A_beI3AcAP1_2;
	wire w_dff_A_QhrjhUhk6_2;
	wire w_dff_A_5r8eP85j4_2;
	wire w_dff_A_WEP0MKFF0_2;
	wire w_dff_A_YrUKhixG1_2;
	wire w_dff_A_eIOkxsDs3_2;
	wire w_dff_A_q5O3GhCj0_2;
	wire w_dff_A_LsF4A0HY3_2;
	wire w_dff_A_jtg43NQK5_2;
	wire w_dff_A_7yNIHFGd2_2;
	wire w_dff_A_QcorbPoi1_2;
	wire w_dff_A_ePWatc187_2;
	wire w_dff_A_XQE8hrzm9_2;
	wire w_dff_A_gUPboYWa9_2;
	wire w_dff_A_t7SZ7ibq3_2;
	wire w_dff_A_i00KGOL32_2;
	wire w_dff_A_HvtO3RM12_2;
	wire w_dff_A_jJI5G6gM5_2;
	wire w_dff_B_VayDGo799_3;
	wire w_dff_B_rDo5NBVx2_3;
	wire w_dff_B_tof5vAxJ8_3;
	wire w_dff_B_ijaMgSks0_0;
	wire w_dff_B_3rEMfBpF3_0;
	wire w_dff_B_hK5XbLPc3_0;
	wire w_dff_B_bzBj97qH0_0;
	wire w_dff_B_GAaUEI6x9_0;
	wire w_dff_B_Mv1xrPiQ3_0;
	wire w_dff_B_r8l9RA577_0;
	wire w_dff_B_ChH0EEBX8_0;
	wire w_dff_B_BSKntXx67_0;
	wire w_dff_B_77aDa9LM9_0;
	wire w_dff_B_UtGWPSW14_0;
	wire w_dff_B_B4SL31yq2_0;
	wire w_dff_B_zfRgEin34_0;
	wire w_dff_B_86m7VksF8_0;
	wire w_dff_B_5avHTFlS5_0;
	wire w_dff_B_UAJSjZ4p4_0;
	wire w_dff_B_xP21tEYM0_0;
	wire w_dff_B_fYPvapMd8_0;
	wire w_dff_B_NGsbwMpe2_0;
	wire w_dff_B_4HAgZNzg2_1;
	wire w_dff_B_nuGxlRcY6_0;
	wire w_dff_B_V51AO53A2_0;
	wire w_dff_B_pUYv3kJb8_0;
	wire w_dff_B_8p8f9pN02_0;
	wire w_dff_B_eDA1cr683_0;
	wire w_dff_B_2NVuRVOw5_0;
	wire w_dff_B_Hr4UWyl12_0;
	wire w_dff_B_CXgMz9647_0;
	wire w_dff_B_OERe5ODg6_0;
	wire w_dff_B_ImMSh5TZ2_0;
	wire w_dff_B_QaXdQIWl1_0;
	wire w_dff_B_1YZVfkZN3_0;
	wire w_dff_B_6rUDTuxD3_0;
	wire w_dff_B_6lcabkyl5_0;
	wire w_dff_B_YhVmrNL97_0;
	wire w_dff_B_mSlToNXx6_0;
	wire w_dff_B_MefwuRR94_0;
	wire w_dff_B_3xR3Qjsu8_0;
	wire w_dff_B_wgTQbKLv9_0;
	wire w_dff_B_MG03m1yT9_0;
	wire w_dff_B_hYjjC3xx1_0;
	wire w_dff_B_kGTsVbyO2_0;
	wire w_dff_B_bZewYbaQ4_0;
	wire w_dff_B_Jyi5VW8h0_1;
	wire w_dff_A_ND9Xw4v67_1;
	wire w_dff_A_x46G1Kg41_1;
	wire w_dff_A_mBJj3KzO0_1;
	wire w_dff_A_YbNCaeJ37_1;
	wire w_dff_A_oTD6dlzB2_1;
	wire w_dff_A_OgqFqi3b7_1;
	wire w_dff_A_Ou7NyWKl8_1;
	wire w_dff_A_Y6s8OPQO9_1;
	wire w_dff_A_2VYW4K1v6_1;
	wire w_dff_A_7fH6kUON8_1;
	wire w_dff_A_cevX7o0u9_1;
	wire w_dff_A_b4P4GOG36_1;
	wire w_dff_A_tEyVDrMj6_1;
	wire w_dff_A_zVfKWdjQ9_1;
	wire w_dff_A_CAAk2uRn9_1;
	wire w_dff_A_PIqAJi5a8_1;
	wire w_dff_A_3NmO94mg2_1;
	wire w_dff_A_3IP9oUZD1_1;
	wire w_dff_A_qc6uFhI29_1;
	wire w_dff_A_fQOs5RJI0_1;
	wire w_dff_A_cHkkuZrw5_1;
	wire w_dff_A_yBrlKAMT0_1;
	wire w_dff_A_L37J9nCp5_1;
	wire w_dff_A_Xlj8jfvv7_1;
	wire w_dff_A_LPFnN2Nq5_1;
	wire w_dff_A_UTUX7qT57_0;
	wire w_dff_A_aqmJyNgr3_0;
	wire w_dff_B_M4BynVLC9_2;
	wire w_dff_B_cUsg1qKh9_2;
	wire w_dff_B_0E7z0d090_2;
	wire w_dff_B_34c1KuyF5_2;
	wire w_dff_B_7Lz0IC683_0;
	wire w_dff_B_Tq42sKlL7_0;
	wire w_dff_B_QJJewbSj4_0;
	wire w_dff_B_1AgZ3Bjn8_0;
	wire w_dff_B_whGa9iPH5_0;
	wire w_dff_B_1AnSKQfI2_0;
	wire w_dff_B_REgLsSAk6_0;
	wire w_dff_B_yoFNMVqF6_0;
	wire w_dff_B_LO8MsGPn6_0;
	wire w_dff_B_MPZomksl0_0;
	wire w_dff_B_qPloL37m9_0;
	wire w_dff_B_EQRiOYtZ7_0;
	wire w_dff_B_5qvJ2mKi1_0;
	wire w_dff_B_VEzlivPG9_0;
	wire w_dff_B_luoQV8yu9_0;
	wire w_dff_B_l96kWJPL1_0;
	wire w_dff_B_lT3Pp4zg7_0;
	wire w_dff_B_JykNhceB1_0;
	wire w_dff_B_JwRnG0pd9_0;
	wire w_dff_A_8AxGSzgb4_1;
	wire w_dff_A_GAnxm2I85_1;
	wire w_dff_A_t9iASt3X5_1;
	wire w_dff_A_zV6UWLfI6_1;
	wire w_dff_A_7y77P9SC0_1;
	wire w_dff_A_2RVeAT833_1;
	wire w_dff_A_e9Go8sPr9_1;
	wire w_dff_A_HxTrJinE0_1;
	wire w_dff_A_nYkfMcrM3_1;
	wire w_dff_A_hbPUZvC87_1;
	wire w_dff_A_OZqdLF5D0_1;
	wire w_dff_A_dEH2fRdO4_1;
	wire w_dff_A_aspEWJ8J4_1;
	wire w_dff_A_UPBiKVTm1_1;
	wire w_dff_A_mxFMN0K67_1;
	wire w_dff_A_r997vqh18_1;
	wire w_dff_A_en48fLNx7_1;
	wire w_dff_A_eIgdf5oS8_1;
	wire w_dff_A_b6NpkqnL3_1;
	wire w_dff_A_l9fYWk477_1;
	wire w_dff_A_keEUnYQ00_1;
	wire w_dff_A_M7KmyMdH9_0;
	wire w_dff_A_tpY9nJRG5_0;
	wire w_dff_A_FNA0fCSX4_0;
	wire w_dff_A_cnEMWUXq2_0;
	wire w_dff_A_JkaivZjF0_0;
	wire w_dff_A_OEgsPleW8_0;
	wire w_dff_A_l1KiWBJ80_0;
	wire w_dff_A_7L673EWa7_0;
	wire w_dff_A_QgYzijuN2_0;
	wire w_dff_A_Edtt8bzm2_0;
	wire w_dff_A_bcSouc1D2_0;
	wire w_dff_A_36YJjSOi8_0;
	wire w_dff_A_cC7PaEWc9_0;
	wire w_dff_A_CaRJ8C2P2_0;
	wire w_dff_A_AR8wxLEs0_0;
	wire w_dff_A_Uv5lnRWA8_0;
	wire w_dff_A_iMxzCyTs2_0;
	wire w_dff_A_xpiY8Ufd5_0;
	wire w_dff_A_liH9GRf56_0;
	wire w_dff_A_9gO6g7tX7_0;
	wire w_dff_A_msS3zn0b7_0;
	wire w_dff_B_OnYKiijy7_1;
	wire w_dff_B_BwhpK7Re8_1;
	wire w_dff_B_u7raKxTd3_1;
	wire w_dff_B_p95jurqh9_1;
	wire w_dff_B_rIxcZSoR5_1;
	wire w_dff_B_i4G7rVJD8_1;
	wire w_dff_B_28qkGFQB2_1;
	wire w_dff_A_UHdhm1WF6_1;
	wire w_dff_A_ThXDYTK74_1;
	wire w_dff_A_wahFABi94_1;
	wire w_dff_A_qhGdko7W8_1;
	wire w_dff_A_oh1B2yho0_1;
	wire w_dff_A_StSoeVLD8_1;
	wire w_dff_B_oiF3CoFo6_0;
	wire w_dff_B_K5OSU1ID5_0;
	wire w_dff_B_uYuGoqJ38_0;
	wire w_dff_B_5A1JMwbV0_0;
	wire w_dff_B_Bib73DXc3_0;
	wire w_dff_B_gxFZF1cC6_0;
	wire w_dff_B_T1a1nCr90_0;
	wire w_dff_B_cmmUvgXQ2_0;
	wire w_dff_B_VcA1N3op7_0;
	wire w_dff_B_DpD6zRwG4_0;
	wire w_dff_B_9EtzbZrf0_0;
	wire w_dff_B_shyeRnQy5_0;
	wire w_dff_B_SzAEIMD45_0;
	wire w_dff_B_Dkxpceow1_0;
	wire w_dff_B_ir71D0UF7_0;
	wire w_dff_B_6iJ4ZQlC5_0;
	wire w_dff_B_R6auYvqy2_0;
	wire w_dff_B_Nrh579qe2_0;
	wire w_dff_B_iVnIzRsb0_1;
	wire w_dff_B_rUCszkdl1_0;
	wire w_dff_B_IKQhlY9y6_0;
	wire w_dff_B_RGnY6viN6_0;
	wire w_dff_B_sJYrScQ83_0;
	wire w_dff_B_YpX15TpO5_0;
	wire w_dff_B_1MTnPnjM5_0;
	wire w_dff_B_9wr4v2i46_0;
	wire w_dff_B_7M0PEGo79_0;
	wire w_dff_B_myCTkUXi8_0;
	wire w_dff_A_QNIvOtTH5_2;
	wire w_dff_A_4pDBzIkj8_0;
	wire w_dff_A_AoXjLKEa2_0;
	wire w_dff_A_0RqgLhFE7_0;
	wire w_dff_A_AV8fO8in9_1;
	wire w_dff_A_GEC2RqG04_0;
	wire w_dff_B_k6xiZitH3_2;
	wire w_dff_B_h91Oegy59_2;
	wire w_dff_B_ceZN13d44_2;
	wire w_dff_B_gItFd5wj3_2;
	wire w_dff_B_UaCCBgEI4_2;
	wire w_dff_B_6cX0yVnW7_2;
	wire w_dff_B_yeZl5t8Z9_2;
	wire w_dff_B_n59tdYKQ9_2;
	wire w_dff_B_GB5UhtBF0_1;
	wire w_dff_A_JsrNYtsM8_0;
	wire w_dff_A_XrVfKjOm6_0;
	wire w_dff_A_HXEhRKtJ6_2;
	wire w_dff_A_TygEWVQm6_2;
	wire w_dff_A_om8WZW3x7_2;
	wire w_dff_A_jj8FWGRv1_0;
	wire w_dff_A_5EyIJLb49_2;
	wire w_dff_A_z84Sivjb7_2;
	wire w_dff_A_0Ti9dv7b3_2;
	wire w_dff_A_FQOPaHzv0_0;
	wire w_dff_A_sWXvFQX26_2;
	wire w_dff_B_kXl7AKD53_1;
	wire w_dff_B_gXPd4Jwn9_1;
	wire w_dff_B_skhcZKns8_1;
	wire w_dff_B_3MxGaw4F7_1;
	wire w_dff_B_1leuiOL64_1;
	wire w_dff_B_6za001C86_1;
	wire w_dff_B_1VpL3ITN8_1;
	wire w_dff_B_GP6CBlmT3_1;
	wire w_dff_A_2scM1JL69_0;
	wire w_dff_A_HT7AMlND8_0;
	wire w_dff_A_3ny3aAEH1_0;
	wire w_dff_A_Wp3jAbI40_0;
	wire w_dff_A_5spAxOzI6_0;
	wire w_dff_A_19uBMY4k7_0;
	wire w_dff_A_7ylir7V19_0;
	wire w_dff_A_clLEDIGw9_0;
	wire w_dff_A_ePeB584u3_0;
	wire w_dff_A_CT1Zwr7E6_0;
	wire w_dff_A_NA3emlrz5_0;
	wire w_dff_A_1tUvtlUT3_0;
	wire w_dff_A_7EcG6Nh41_0;
	wire w_dff_A_4n9Cq2BZ1_0;
	wire w_dff_A_xbcpzsOe3_0;
	wire w_dff_A_pWnRGosz6_0;
	wire w_dff_A_Nfs8BZD57_0;
	wire w_dff_A_fVC9dVDB5_0;
	wire w_dff_A_9jIclCX84_0;
	wire w_dff_A_G9eBYFVB8_0;
	wire w_dff_A_73VINfOf7_0;
	wire w_dff_A_q4Rcgtd79_0;
	wire w_dff_A_VuJDRYHz4_0;
	wire w_dff_A_PFxXQQEF3_0;
	wire w_dff_A_biG1YBpe4_0;
	wire w_dff_A_UOo25iMB9_0;
	wire w_dff_A_2DWOwWGn1_0;
	wire w_dff_A_otJcy7zp3_0;
	wire w_dff_A_P3Kbsd9q8_0;
	wire w_dff_A_9QatQ9tk9_0;
	wire w_dff_A_SiChp53D2_2;
	wire w_dff_A_OpQKdVDa4_2;
	wire w_dff_A_CsClAuT21_2;
	wire w_dff_A_iNggLAeh1_2;
	wire w_dff_A_khjwgLvX2_2;
	wire w_dff_B_4URZCTKT2_1;
	wire w_dff_B_IIRAvDTi4_1;
	wire w_dff_B_H9669h9Z1_1;
	wire w_dff_B_XCrdcWAr7_1;
	wire w_dff_B_MScwB68L7_1;
	wire w_dff_B_n5I8J8zb3_1;
	wire w_dff_B_VecfdJva2_1;
	wire w_dff_B_lmdSCRQa8_1;
	wire w_dff_B_dQLeCAFX5_1;
	wire w_dff_B_52g9Ls848_1;
	wire w_dff_B_NATieFFa3_1;
	wire w_dff_B_2ZjSOoZk1_1;
	wire w_dff_B_K565x8eR5_1;
	wire w_dff_B_jJYMotSy6_1;
	wire w_dff_B_DPT6iVDN3_1;
	wire w_dff_B_2Rq562tP6_1;
	wire w_dff_B_v5OaJ4Ow5_1;
	wire w_dff_B_1eXPyZuP0_1;
	wire w_dff_B_2yN8lW562_1;
	wire w_dff_B_4bfEc6Q59_1;
	wire w_dff_B_iKOJSfaE1_1;
	wire w_dff_B_OBsVua4Z4_1;
	wire w_dff_B_dUJDzBcM6_1;
	wire w_dff_B_YoHRC7kQ1_1;
	wire w_dff_B_KUJFyn363_1;
	wire w_dff_B_a0A0R9iS4_1;
	wire w_dff_B_iBqu3Y7d7_1;
	wire w_dff_B_57n7TXKg3_1;
	wire w_dff_B_EzkNbk9Z3_1;
	wire w_dff_B_YaANBgLp9_1;
	wire w_dff_B_QwCIe8H74_1;
	wire w_dff_B_zAPGi7sQ9_0;
	wire w_dff_B_kpcEDEf08_0;
	wire w_dff_B_cxTFnbYF4_0;
	wire w_dff_B_uPPHhfSG4_0;
	wire w_dff_B_XK8ll53l8_0;
	wire w_dff_B_azRK4Jwg0_0;
	wire w_dff_B_QVinhlI20_0;
	wire w_dff_B_rawBPdkp5_0;
	wire w_dff_B_fexPNuMS8_0;
	wire w_dff_B_MaMLRemh2_0;
	wire w_dff_B_A901igYJ6_0;
	wire w_dff_B_dxs6qdP81_0;
	wire w_dff_B_LVMcigG42_0;
	wire w_dff_B_EOpICpsq9_0;
	wire w_dff_B_sA3whaAc2_0;
	wire w_dff_B_gvLAsJf49_0;
	wire w_dff_B_vfS4H3GJ8_0;
	wire w_dff_B_IU8FPb0D3_0;
	wire w_dff_B_3IfdK66J1_0;
	wire w_dff_B_AHUCtzZZ4_0;
	wire w_dff_B_VG3jWbMU3_1;
	wire w_dff_B_Wz9LiyGS3_1;
	wire w_dff_B_xStXXyDX5_0;
	wire w_dff_B_8C6OP5B58_0;
	wire w_dff_B_EkJW2d739_0;
	wire w_dff_B_GfHZKRgn0_0;
	wire w_dff_B_7TJ07BqD6_0;
	wire w_dff_A_FGO3VwDe7_1;
	wire w_dff_A_4GxBDFuK5_1;
	wire w_dff_A_9Dandry36_1;
	wire w_dff_A_WsZgq4ld1_1;
	wire w_dff_A_62agWQZ76_1;
	wire w_dff_A_AquFdCbi3_1;
	wire w_dff_A_FE4fiykW8_1;
	wire w_dff_A_pOPNpuih6_1;
	wire w_dff_A_A4OjkDoC9_1;
	wire w_dff_A_96IQSY3P0_1;
	wire w_dff_A_rcEpXCLT9_1;
	wire w_dff_A_FueC69Vb4_1;
	wire w_dff_A_VZSUXcJR1_1;
	wire w_dff_A_XdQMZGYT8_1;
	wire w_dff_A_KKXS9DGc4_1;
	wire w_dff_A_iEOT29u52_1;
	wire w_dff_A_xhJreGxM4_1;
	wire w_dff_A_5rZqYOZF2_1;
	wire w_dff_A_JMGaejtI5_1;
	wire w_dff_A_6kHtavVd7_1;
	wire w_dff_A_BtTuPcIS1_1;
	wire w_dff_A_VTtE4p5y2_1;
	wire w_dff_A_aMUHQ7Iu9_1;
	wire w_dff_A_G14UZ7Ts8_1;
	wire w_dff_A_xuCJl1nq8_1;
	wire w_dff_B_6dr2HROu8_0;
	wire w_dff_B_CJN2F4J86_0;
	wire w_dff_B_6Xm9GNkp1_0;
	wire w_dff_B_jvy3VoAt6_1;
	wire w_dff_B_iTP5sQCM5_1;
	wire w_dff_B_SFXMS2uJ4_1;
	wire w_dff_B_qVejruuc3_1;
	wire w_dff_B_zpFoqYh97_1;
	wire w_dff_A_qQNwmH5o6_1;
	wire w_dff_A_nVFKisTE2_1;
	wire w_dff_A_ktLMMZcL7_1;
	wire w_dff_A_SLotKsRL8_1;
	wire w_dff_A_EzpjlKyO6_1;
	wire w_dff_A_HfGWA7UL9_1;
	wire w_dff_A_hKV06LHL6_1;
	wire w_dff_A_7nE0DL139_1;
	wire w_dff_A_YmS8dCMC5_1;
	wire w_dff_A_UbIBYy1D3_1;
	wire w_dff_A_k0dx8DWQ3_1;
	wire w_dff_A_0m2DTqYc6_1;
	wire w_dff_A_TCvrdDZE9_1;
	wire w_dff_A_7Ayixigf7_1;
	wire w_dff_A_Iq0hghM34_1;
	wire w_dff_A_nYKAr1b15_1;
	wire w_dff_A_ARd6ITmS7_1;
	wire w_dff_A_GXlCHxSq3_1;
	wire w_dff_A_1i44VYq57_1;
	wire w_dff_A_xdS4xNOl2_1;
	wire w_dff_A_6GealkN51_1;
	wire w_dff_A_OQiWABd12_1;
	wire w_dff_B_H8oXmmA94_2;
	wire w_dff_A_nfikk4AQ6_0;
	wire w_dff_A_lkcE2c0P4_0;
	wire w_dff_A_qxMPcfHI4_0;
	wire w_dff_A_h4etcT9V1_0;
	wire w_dff_A_iWAGMO7h6_0;
	wire w_dff_B_bFGdTcFl7_1;
	wire w_dff_B_uktRUa4U6_1;
	wire w_dff_B_yPB3bYIt8_1;
	wire w_dff_B_SnoR0ISc2_1;
	wire w_dff_B_a6kOW1KS8_1;
	wire w_dff_B_mZtiIKQf2_1;
	wire w_dff_B_pZ9D4wAW0_1;
	wire w_dff_B_GclWk9i40_1;
	wire w_dff_B_NEiHFAHC2_1;
	wire w_dff_B_aR29EeWm8_1;
	wire w_dff_B_URtq9owT4_1;
	wire w_dff_B_4g3291wX8_1;
	wire w_dff_B_X2fhvDj11_1;
	wire w_dff_B_JJ2mHynC8_1;
	wire w_dff_B_gUZoFocb4_1;
	wire w_dff_B_GFxji9EJ8_1;
	wire w_dff_B_HE4ZSF592_1;
	wire w_dff_B_48tK7MUN0_1;
	wire w_dff_B_Su3kwOrT5_1;
	wire w_dff_B_DkS7F9ki1_1;
	wire w_dff_B_OiLJXAWd0_1;
	wire w_dff_B_jet4qFZK3_1;
	wire w_dff_B_0LPA7P8j1_1;
	wire w_dff_B_lInV46iW7_1;
	wire w_dff_B_8xwmUzaQ2_1;
	wire w_dff_B_sn5wKndL8_1;
	wire w_dff_B_k4OnJtg44_1;
	wire w_dff_B_zmbOQOvP3_1;
	wire w_dff_B_U3fnmt7e9_1;
	wire w_dff_B_PXcm5kGH7_1;
	wire w_dff_B_Du06je7b1_1;
	wire w_dff_B_4e5OsMwi1_1;
	wire w_dff_B_Nt7kok2D2_1;
	wire w_dff_B_LHcp6NtL3_1;
	wire w_dff_B_s0BKhxcC7_1;
	wire w_dff_B_uXUOpUnp0_1;
	wire w_dff_B_IuDRgzOw6_1;
	wire w_dff_B_iX6HCfrX8_1;
	wire w_dff_B_TkAQmy2F6_1;
	wire w_dff_B_HZP9cHmN3_1;
	wire w_dff_B_SErHn3Co3_1;
	wire w_dff_B_a5KWdw619_1;
	wire w_dff_B_6nfR4x0N9_1;
	wire w_dff_B_oqP1e4z64_1;
	wire w_dff_B_HrBH1RxL0_1;
	wire w_dff_B_yxSWqYma7_1;
	wire w_dff_B_o8Emg5SK9_1;
	wire w_dff_B_Rktz6AM47_1;
	wire w_dff_B_0QIdrxkI4_1;
	wire w_dff_B_Cf7HDrTi8_1;
	wire w_dff_B_ZsIJhXav8_1;
	wire w_dff_B_MpGPcPli1_1;
	wire w_dff_B_QxqAoEww1_1;
	wire w_dff_B_usKxzaUL4_1;
	wire w_dff_B_vp9A2Y2X7_1;
	wire w_dff_B_cESwo7Oj0_1;
	wire w_dff_B_R69Topu95_1;
	wire w_dff_B_67skyuQZ3_1;
	wire w_dff_B_AxBhauOz4_1;
	wire w_dff_B_KEgrpVWj1_1;
	wire w_dff_B_8zSm99nB1_1;
	wire w_dff_B_gPFETUWy8_1;
	wire w_dff_B_BQXFmObV5_1;
	wire w_dff_B_pKtYLJ7Z5_1;
	wire w_dff_B_wV0BdER56_1;
	wire w_dff_B_JPv22FWC9_1;
	wire w_dff_B_XnJiykrU9_1;
	wire w_dff_B_FL6Sb9Lk6_1;
	wire w_dff_B_T0wtvQYU4_1;
	wire w_dff_B_cCF5SyOg4_1;
	wire w_dff_B_KX9axuSC7_1;
	wire w_dff_B_NOkpmACW8_1;
	wire w_dff_B_Jb6RIUga0_1;
	wire w_dff_B_vdkrFCYN1_1;
	wire w_dff_B_ZsqlCYh01_1;
	wire w_dff_B_rnCe3Ork8_1;
	wire w_dff_B_k128GXOQ4_1;
	wire w_dff_B_8v1f5lu64_1;
	wire w_dff_B_qDMTBvTM4_1;
	wire w_dff_B_RpTJ8ne29_1;
	wire w_dff_B_AshLw6qE3_1;
	wire w_dff_B_Tc9xDrxg9_1;
	wire w_dff_B_5mxyAtXC7_1;
	wire w_dff_B_nrRkeC0n1_1;
	wire w_dff_B_sJ1BlAHw3_1;
	wire w_dff_B_NgtP7nAb7_1;
	wire w_dff_B_rae1xR3N7_1;
	wire w_dff_B_IK8yuc0C4_1;
	wire w_dff_B_3kuzFPr53_1;
	wire w_dff_B_CyWgGN208_1;
	wire w_dff_B_NNvIj3sz2_1;
	wire w_dff_B_qnAH5L7I0_1;
	wire w_dff_B_RgWgAMLJ0_1;
	wire w_dff_B_Jrt6afgO4_1;
	wire w_dff_B_4gExAVhN2_1;
	wire w_dff_B_lwVZCQWe7_1;
	wire w_dff_B_nd1RsLIr9_1;
	wire w_dff_B_HCXKnUV56_1;
	wire w_dff_B_44gYAvYT5_1;
	wire w_dff_B_ODsjwKZU9_1;
	wire w_dff_B_ohRFURxK8_1;
	wire w_dff_B_hw8qqWUl6_1;
	wire w_dff_B_ZFrDDfpJ6_1;
	wire w_dff_B_D5IQZtkR1_1;
	wire w_dff_B_UPCU2CmB6_1;
	wire w_dff_B_u6yzwprT5_1;
	wire w_dff_B_BonRRWPv8_1;
	wire w_dff_B_77XlgZEc1_1;
	wire w_dff_B_Akr6oeE66_1;
	wire w_dff_B_D03abrMJ9_1;
	wire w_dff_B_8lvX44m70_1;
	wire w_dff_B_MQlJAE9M7_1;
	wire w_dff_B_NAgtVxZD0_1;
	wire w_dff_B_Y5YldpcH8_1;
	wire w_dff_B_DP4CX1mM1_1;
	wire w_dff_B_5tklbAaM3_1;
	wire w_dff_B_Byl5Z62t8_1;
	wire w_dff_B_ytgcOuN60_1;
	wire w_dff_B_0kADtmeq4_1;
	wire w_dff_B_u6FH1tbz5_1;
	wire w_dff_B_jW935lNA8_1;
	wire w_dff_B_rLGvwbtD6_1;
	wire w_dff_B_nlH3rkY76_1;
	wire w_dff_B_i7s5kYnd1_1;
	wire w_dff_B_wYoPpZ6N7_1;
	wire w_dff_B_YTdOoUHr3_1;
	wire w_dff_B_e52IBdTD4_1;
	wire w_dff_B_j0QpTQHF5_1;
	wire w_dff_B_TOdfTB2l7_1;
	wire w_dff_B_rHabs0Ds3_1;
	wire w_dff_B_xlnIwjUB5_1;
	wire w_dff_B_epeUJmat6_1;
	wire w_dff_B_3bOwUSDR6_1;
	wire w_dff_B_7oCASZGe3_1;
	wire w_dff_B_4VyW49zX9_1;
	wire w_dff_B_pk97WiTA1_1;
	wire w_dff_B_xZKYKqV27_1;
	wire w_dff_B_Mz1q1YI47_1;
	wire w_dff_B_o1XJSCTh3_1;
	wire w_dff_B_IGC0S6jD6_1;
	wire w_dff_B_aTPdqReg6_1;
	wire w_dff_B_vxIYgitq5_1;
	wire w_dff_B_ZXtwGK773_1;
	wire w_dff_B_2iFnCUuU8_1;
	wire w_dff_B_RsyCdviq3_1;
	wire w_dff_B_nfriTmIm4_1;
	wire w_dff_B_oO0jZObY5_1;
	wire w_dff_B_BrvrR8gC2_1;
	wire w_dff_B_LJxHPsYZ4_1;
	wire w_dff_B_luDCltd93_1;
	wire w_dff_B_jDfHQxtX6_1;
	wire w_dff_B_padfVtME6_1;
	wire w_dff_B_YNsgfuEa4_1;
	wire w_dff_B_ySbCi0UA4_1;
	wire w_dff_B_sT2LG1VA4_1;
	wire w_dff_B_VkuhmvWQ4_1;
	wire w_dff_B_weELPwBH8_1;
	wire w_dff_B_MoK8K3V77_1;
	wire w_dff_B_aFiCM8Xa7_1;
	wire w_dff_B_RmXhfKrA5_1;
	wire w_dff_B_A9342yTM3_1;
	wire w_dff_B_DuUQPFvb7_1;
	wire w_dff_B_uo74DPz82_1;
	wire w_dff_B_PncgLYtv6_1;
	wire w_dff_B_1oMPnq7s8_1;
	wire w_dff_B_Y4voQsKt4_1;
	wire w_dff_B_6ZOy3w3J2_1;
	wire w_dff_B_OcKKJx5L0_1;
	wire w_dff_B_MLZPxglE7_1;
	wire w_dff_B_1H8NVeIm3_1;
	wire w_dff_B_ikio3lpP7_1;
	wire w_dff_A_IuxooMrp3_0;
	wire w_dff_B_g5yGYdSh2_2;
	wire w_dff_B_roBgkliS7_2;
	wire w_dff_B_5yXtPHCI4_2;
	wire w_dff_B_czORjX8i6_2;
	wire w_dff_B_vkNiYCuI6_2;
	wire w_dff_B_AamhJqBS7_2;
	wire w_dff_B_omN9lnRC1_2;
	wire w_dff_B_BvWSSrzu4_2;
	wire w_dff_B_V4gj3nKw4_2;
	wire w_dff_B_SMP7N7Ck0_2;
	wire w_dff_B_Up4m6slZ1_2;
	wire w_dff_B_UrTGNWhK7_2;
	wire w_dff_B_mBdl030i6_2;
	wire w_dff_B_8pQKnd758_2;
	wire w_dff_B_6ObSEDAw4_2;
	wire w_dff_B_KGY4CxUr5_2;
	wire w_dff_B_qXfQcp5F7_2;
	wire w_dff_B_Y5woxDGt8_2;
	wire w_dff_B_AGhvN9KA2_0;
	wire w_dff_B_0gJncxEk9_0;
	wire w_dff_B_AdBgfhpW3_0;
	wire w_dff_B_0TCVwuZs8_0;
	wire w_dff_B_rfKLOvf55_0;
	wire w_dff_B_05v4G4EF4_0;
	wire w_dff_B_FOqQI0gV0_0;
	wire w_dff_B_8ImvVHjO3_0;
	wire w_dff_B_X2YReIlf9_0;
	wire w_dff_B_LZXWKBZ50_0;
	wire w_dff_B_9xnFQAWl5_0;
	wire w_dff_B_98YENKx82_0;
	wire w_dff_B_E4vM521R1_0;
	wire w_dff_B_L07YgFGf5_0;
	wire w_dff_B_svOPQ0IX8_0;
	wire w_dff_B_XoqK1Qrf7_0;
	wire w_dff_B_mNVELAZ65_0;
	wire w_dff_B_wNjScP6a2_0;
	wire w_dff_B_F1pYMPkp7_0;
	wire w_dff_B_f6SH1Swa5_0;
	wire w_dff_B_QktJqICt2_0;
	wire w_dff_B_sF6oPbsM6_0;
	wire w_dff_B_5kIPSHbN4_0;
	wire w_dff_B_4T9BR8210_0;
	wire w_dff_B_Kzz4PDiU8_0;
	wire w_dff_B_nODN7bvz1_0;
	wire w_dff_A_gwZYhnKO5_1;
	wire w_dff_A_RvPdg9DA4_1;
	wire w_dff_A_r5vwT7TT8_1;
	wire w_dff_A_0EY8Gc0Y3_1;
	wire w_dff_A_L9KEOYBB9_1;
	wire w_dff_A_m5ViydYv5_1;
	wire w_dff_A_yoPZSWl13_1;
	wire w_dff_A_qWKx2dOq8_1;
	wire w_dff_B_eFgGSVwm2_1;
	wire w_dff_B_0FngQeLD3_1;
	wire w_dff_A_eZXnlpvS8_1;
	wire w_dff_A_6h3bIYF37_1;
	wire w_dff_A_7VYmYoYr9_1;
	wire w_dff_A_2poalKMA2_1;
	wire w_dff_A_KIx2VHi19_1;
	wire w_dff_A_5cO6ktaw9_1;
	wire w_dff_A_JejYPRDo3_1;
	wire w_dff_A_wCJ2uaZ43_1;
	wire w_dff_A_6xxYKv2a0_1;
	wire w_dff_A_tylyX5up8_1;
	wire w_dff_A_EZadv2aC4_1;
	wire w_dff_A_K311HNM89_1;
	wire w_dff_A_3pwP2hv86_1;
	wire w_dff_A_4NJksY3z7_1;
	wire w_dff_A_1Mj12XJM8_1;
	wire w_dff_A_fEZDBPaJ9_1;
	wire w_dff_A_9ZwlWKzu7_1;
	wire w_dff_A_BZTD7tpw2_1;
	wire w_dff_A_qjjDobR02_1;
	wire w_dff_A_OjhF358c0_1;
	wire w_dff_A_Tz7kdlG23_1;
	wire w_dff_A_9McRTXCu6_1;
	wire w_dff_A_XBoqCcEx7_1;
	wire w_dff_A_fdzOriLl1_1;
	wire w_dff_A_vYHgwxc30_1;
	wire w_dff_A_PZw6Hh9P7_1;
	wire w_dff_A_jarPTf8q0_1;
	wire w_dff_A_Mo5ZWezW7_1;
	wire w_dff_B_AnofVKPO2_2;
	wire w_dff_B_lJ5QNjnV4_2;
	wire w_dff_A_g92e85O21_2;
	wire w_dff_A_aglXCVb96_2;
	wire w_dff_A_YWRAjuvE8_2;
	wire w_dff_A_i34odZJ98_2;
	wire w_dff_A_3uf1oS8C3_2;
	wire w_dff_A_fYTI9cJ48_2;
	wire w_dff_A_AevRGeN78_2;
	wire w_dff_A_3J8NWZDi6_2;
	wire w_dff_A_TnqrOvdt0_2;
	wire w_dff_A_51aRyeB72_2;
	wire w_dff_A_woUc07xg0_2;
	wire w_dff_A_IjzyheDb7_2;
	wire w_dff_A_CxhTikps9_2;
	wire w_dff_A_MQNbCX390_2;
	wire w_dff_A_UE8spiDH8_2;
	wire w_dff_A_qrthNcPY3_2;
	wire w_dff_A_nXS0nba76_2;
	wire w_dff_A_W52wLRxE4_2;
	wire w_dff_A_jRNRbCtR5_2;
	wire w_dff_A_v90dEzJ47_2;
	wire w_dff_A_DvqT2GfO2_2;
	wire w_dff_A_gAZ44v0g8_2;
	wire w_dff_A_C5SgrmPL0_2;
	wire w_dff_B_Xzk5kxbQ0_1;
	wire w_dff_B_EDueLPXN5_1;
	wire w_dff_B_pYGNNO9i9_1;
	wire w_dff_B_9j5IoNto8_1;
	wire w_dff_B_RWZ0nrv75_1;
	wire w_dff_B_erbnnowH2_1;
	wire w_dff_B_R04qSkmn0_1;
	wire w_dff_B_ZQDWXIqq6_1;
	wire w_dff_B_Cw6wK2kq0_1;
	wire w_dff_A_BrJEZedj3_2;
	wire w_dff_A_HHPEyq3M9_2;
	wire w_dff_A_CJL8xyZz6_2;
	wire w_dff_A_dVODatoS0_2;
	wire w_dff_A_oU1ZM55K8_2;
	wire w_dff_A_sGjIIncj7_2;
	wire w_dff_A_6llkRCZ02_2;
	wire w_dff_A_SIOtIOml7_2;
	wire w_dff_A_glWGlEd73_2;
	wire w_dff_A_Cgz9fZJ48_2;
	wire w_dff_A_OILiBMmN9_2;
	wire w_dff_A_XSWRAldS2_2;
	wire w_dff_A_9HBIlFH77_2;
	wire w_dff_A_skJRAPsS0_2;
	wire w_dff_A_SPi4HDhp5_2;
	wire w_dff_A_LoqPWNol5_2;
	wire w_dff_A_UUzoMG4o9_2;
	wire w_dff_A_lhgEor1P6_2;
	wire w_dff_A_zMNFwiqL0_2;
	wire w_dff_A_jYck3y3b9_2;
	wire w_dff_A_2NPYQQ0K2_2;
	wire w_dff_A_BzExDJok8_2;
	wire w_dff_A_lXNnTDcK2_2;
	wire w_dff_A_r0jkB8Pt3_2;
	wire w_dff_A_Amuwpa848_2;
	wire w_dff_B_ip9tF0zH7_1;
	wire w_dff_A_0KsNRUZ00_0;
	wire w_dff_A_Vzst1tsa8_1;
	wire w_dff_A_HW0CNNaM1_1;
	wire w_dff_A_LiijGa0q0_1;
	wire w_dff_A_Rk8SrjUc5_1;
	wire w_dff_A_DSp4yWnr1_1;
	wire w_dff_A_LmdZapYT8_1;
	wire w_dff_A_Q4snMDE10_1;
	wire w_dff_A_nczq2ASh7_1;
	wire w_dff_A_rqdMaNH98_1;
	wire w_dff_A_K1SvHrs10_1;
	wire w_dff_A_Z4gY4QN91_1;
	wire w_dff_A_v3e3znSJ6_1;
	wire w_dff_A_986pFOJR1_1;
	wire w_dff_A_5DzojULb4_1;
	wire w_dff_A_Wrp4ADXB5_1;
	wire w_dff_A_EKEE6Tlo2_1;
	wire w_dff_A_b7NjEgFW8_1;
	wire w_dff_A_A9wfmooN6_1;
	wire w_dff_A_mTKAX2b75_1;
	wire w_dff_A_Z0DGIgll9_1;
	wire w_dff_A_Xxub7PmQ3_1;
	wire w_dff_A_Pq2XUUwU2_1;
	wire w_dff_A_jcUCBrq45_1;
	wire w_dff_A_dkolpX118_1;
	wire w_dff_A_njsPvHKF3_1;
	wire w_dff_A_hbAV5I5r2_1;
	wire w_dff_A_RhSNtQ7o7_1;
	wire w_dff_A_vHpQMJM47_1;
	wire w_dff_A_Apmk8SeQ1_1;
	wire w_dff_A_BhdubKHE1_1;
	wire w_dff_A_5xjHTlCY6_1;
	wire w_dff_A_nsaHze9V0_1;
	wire w_dff_B_bZf3Y5AV4_0;
	wire w_dff_A_rOTyxRsQ1_0;
	wire w_dff_A_BBzGkKiJ5_0;
	wire w_dff_A_ueWiOO963_1;
	wire w_dff_A_oj1IjktD9_1;
	wire w_dff_A_MChL85tW9_0;
	wire w_dff_A_XMXSjf4L9_0;
	wire w_dff_A_UyLnJLpV5_0;
	wire w_dff_A_XvxZdTNf7_0;
	wire w_dff_A_wx8BE9BM7_0;
	wire w_dff_B_SYp4AUKk5_2;
	wire w_dff_A_5XFw2BK36_0;
	wire w_dff_A_qqy3ED7z2_0;
	wire w_dff_A_GpfuqmSP6_1;
	wire w_dff_A_JXnlarNW9_1;
	wire w_dff_A_j3rjMdM79_0;
	wire w_dff_A_SRJSWJeu4_2;
	wire w_dff_A_vKP5qq0L8_0;
	wire w_dff_A_t6sCCjTH2_0;
	wire w_dff_A_p5p2AGaa0_2;
	wire w_dff_A_zbGCICaN3_2;
	wire w_dff_A_eO1qbKxK0_2;
	wire w_dff_A_bSvOCi7B0_2;
	wire w_dff_A_TP1DRJpF5_2;
	wire w_dff_A_zxZQCvQJ6_2;
	wire w_dff_A_idthlT9g4_2;
	wire w_dff_A_kjpjMtHF4_0;
	wire w_dff_A_tkqNoS2v5_0;
	wire w_dff_B_a909KlhV4_0;
	wire w_dff_A_X1TuwsZf3_1;
	wire w_dff_A_nuxPCBOz4_1;
	wire w_dff_A_FM3mH6a44_2;
	wire w_dff_A_fWSAdVKo6_2;
	wire w_dff_B_dxI4Drpe8_1;
	wire w_dff_B_pmThCi3D0_1;
	wire w_dff_B_iAKDS9Hl0_1;
	wire w_dff_B_fLkGQpSK7_1;
	wire w_dff_B_ouyj905a4_1;
	wire w_dff_B_wsYh0W1j6_1;
	wire w_dff_B_s7kfYvyR7_1;
	wire w_dff_B_djipIL9X3_1;
	wire w_dff_B_HaqvBl8E4_1;
	wire w_dff_B_3wgKmfbH2_1;
	wire w_dff_B_g1HA1iMZ8_1;
	wire w_dff_B_hV6BjzUi4_1;
	wire w_dff_B_gLD3NANP0_1;
	wire w_dff_B_6uYLmdzp6_1;
	wire w_dff_B_1XOwPlP90_1;
	wire w_dff_B_jhN7ONri7_1;
	wire w_dff_B_jQqlgt9b9_1;
	wire w_dff_B_eOrW3sMd4_1;
	wire w_dff_B_ivJcWUpd4_1;
	wire w_dff_B_A9ljM3pL5_0;
	wire w_dff_B_vWTXuyzV1_0;
	wire w_dff_B_gFmnUpz72_0;
	wire w_dff_B_5hs3d9dS8_0;
	wire w_dff_B_glKRk3gR5_0;
	wire w_dff_B_9rtOB0Lq3_0;
	wire w_dff_B_3yjIZrto9_0;
	wire w_dff_B_O2veVFGl5_0;
	wire w_dff_B_7TVa7QrY6_0;
	wire w_dff_B_sagEw58q7_0;
	wire w_dff_B_c6HAdUaN2_0;
	wire w_dff_B_lAEfoLb51_0;
	wire w_dff_B_n6A6nBpW3_0;
	wire w_dff_B_pce0MwIA2_0;
	wire w_dff_A_I7xDzB0S6_0;
	wire w_dff_A_cNv0txgm3_0;
	wire w_dff_A_aoVUsHNH4_0;
	wire w_dff_A_uMMjXF7A7_0;
	wire w_dff_A_jRglSfii3_0;
	wire w_dff_A_5hsSyzRu8_0;
	wire w_dff_A_aXu3DKeP5_0;
	wire w_dff_A_nmfzxFhA3_0;
	wire w_dff_A_USPKJ8132_0;
	wire w_dff_A_X2pZoTDj5_0;
	wire w_dff_A_f4xdTZ1k0_0;
	wire w_dff_A_Rszs5hxt9_0;
	wire w_dff_A_0C7stwN52_0;
	wire w_dff_A_JicpSNRF3_0;
	wire w_dff_A_b1VtYyyq2_0;
	wire w_dff_B_4l6EjjZ92_1;
	wire w_dff_B_4mONRwjK5_1;
	wire w_dff_B_2OvdcqoQ8_1;
	wire w_dff_B_tWHvgilG5_1;
	wire w_dff_B_j3c8LBmL0_1;
	wire w_dff_B_NRkqAHc08_1;
	wire w_dff_B_UU5OWMm29_1;
	wire w_dff_B_FF9BiwNp5_1;
	wire w_dff_B_ydLvFe607_1;
	wire w_dff_B_OaK0ATQs6_1;
	wire w_dff_B_BkLkavyk7_1;
	wire w_dff_B_xt3rlacS3_1;
	wire w_dff_B_Nb90LzJ29_1;
	wire w_dff_B_xEI4AJRJ0_1;
	wire w_dff_B_BuNIFx2m3_1;
	wire w_dff_B_uwJGeuQo2_1;
	wire w_dff_B_fLrw1hNJ4_1;
	wire w_dff_B_KpiQnyyo5_1;
	wire w_dff_B_4YOywbhc6_1;
	wire w_dff_B_pE2wBYNa4_1;
	wire w_dff_B_ZCvoo7Hx9_1;
	wire w_dff_B_pW0r1VbN2_1;
	wire w_dff_B_ZnnPsRxJ0_1;
	wire w_dff_B_MQNi7O0W7_1;
	wire w_dff_B_aoeJBiiz8_1;
	wire w_dff_B_P0hiPupE3_1;
	wire w_dff_B_HR0JZQQm7_1;
	wire w_dff_B_BPWMRp4e6_1;
	wire w_dff_B_hD6mkblq0_1;
	wire w_dff_B_bOk8bYvH9_1;
	wire w_dff_B_sBFOXOMN7_1;
	wire w_dff_B_vvQeQ9IZ6_1;
	wire w_dff_B_KrkYt20q1_1;
	wire w_dff_B_qToOmZvf7_1;
	wire w_dff_A_4AY1VK1h7_1;
	wire w_dff_A_OiCKnY8w5_1;
	wire w_dff_A_e0Ejqhux7_1;
	wire w_dff_A_5h6Q7F6G2_1;
	wire w_dff_A_kBBqhWdO2_1;
	wire w_dff_A_A1dL6dWk5_1;
	wire w_dff_A_n0BAAhXE8_1;
	wire w_dff_A_8vjMpDMc9_1;
	wire w_dff_A_F3FI9HFu1_1;
	wire w_dff_A_bUTvmJwf9_1;
	wire w_dff_A_W6Q6hwAB4_1;
	wire w_dff_A_CcYGYwLY7_1;
	wire w_dff_A_UGw49bNO0_1;
	wire w_dff_A_elMZDeJw5_1;
	wire w_dff_A_IATSXNEX0_1;
	wire w_dff_A_7TcVFsax4_1;
	wire w_dff_A_YY9Wa9DR3_1;
	wire w_dff_A_wAQ3i3Jc9_1;
	wire w_dff_A_6rMMNjas3_1;
	wire w_dff_A_mysvAp8W3_0;
	wire w_dff_A_W2jLkjl70_0;
	wire w_dff_A_wBl7ND0M6_0;
	wire w_dff_A_1kHYwltR7_0;
	wire w_dff_A_wVENETGK6_0;
	wire w_dff_A_9T32hcbM6_0;
	wire w_dff_A_cIucq7oY5_0;
	wire w_dff_A_DIfLTP544_0;
	wire w_dff_A_FEqIZsnq9_0;
	wire w_dff_A_EurOJcZ53_0;
	wire w_dff_A_8oSIy0W82_0;
	wire w_dff_A_4nbLLgR66_0;
	wire w_dff_A_N0awK1a70_0;
	wire w_dff_A_hY21ZafV7_0;
	wire w_dff_A_4jEY70Uv7_0;
	wire w_dff_A_hVdWN37r8_0;
	wire w_dff_A_bZG6rCt02_0;
	wire w_dff_A_j8Yyd3C18_0;
	wire w_dff_A_TytrfGEn0_0;
	wire w_dff_A_nQGtR75U2_0;
	wire w_dff_A_wXmX0e7m5_1;
	wire w_dff_A_dhNvzuby7_1;
	wire w_dff_A_DJqP3u7M2_1;
	wire w_dff_A_7Fqir6Uc3_1;
	wire w_dff_A_lRaNFEFP2_1;
	wire w_dff_A_4lf6tUkl5_1;
	wire w_dff_A_xVpNistd5_1;
	wire w_dff_A_4Q0HkovC8_1;
	wire w_dff_A_05cVpLKY5_1;
	wire w_dff_A_I3EHgkKR5_1;
	wire w_dff_A_TDuqIGv35_1;
	wire w_dff_A_H5Du67Uf9_1;
	wire w_dff_A_4FXWiXsM1_1;
	wire w_dff_A_DavtVEpX0_1;
	wire w_dff_A_Cfo0Ft2p4_1;
	wire w_dff_A_92OGamdW0_1;
	wire w_dff_A_lUlKWWju8_1;
	wire w_dff_A_IsUwWonB5_1;
	wire w_dff_A_ZAjNNJfD7_1;
	wire w_dff_A_1VSTvnbX6_1;
	wire w_dff_A_gHh1LAwz8_1;
	wire w_dff_A_RxW72wH48_1;
	wire w_dff_A_pV3i2Oqw1_1;
	wire w_dff_A_rZ0hgTC95_1;
	wire w_dff_A_hQTC4fE15_1;
	wire w_dff_A_mslwNtHw0_1;
	wire w_dff_A_ijRyzMBZ9_1;
	wire w_dff_A_wlVkLV6h4_1;
	wire w_dff_A_yWUIeNXJ3_1;
	wire w_dff_A_pQb2xkDp4_1;
	wire w_dff_A_8yZtTeNR1_1;
	wire w_dff_A_HSRsi5bl1_1;
	wire w_dff_A_cFUZ2Tor7_1;
	wire w_dff_A_3YjeGyEk6_1;
	wire w_dff_A_kodrTzqj5_1;
	wire w_dff_A_lMCx3fHi1_1;
	wire w_dff_A_ySDlUllu3_1;
	wire w_dff_A_fNRZdPWU1_1;
	wire w_dff_A_wmgdaXR69_1;
	wire w_dff_A_AJ2RaLHq2_1;
	wire w_dff_A_ZHrf0Wum6_1;
	wire w_dff_A_tIa5nNvV2_1;
	wire w_dff_A_g1XOuA2k6_1;
	wire w_dff_A_5RRLB7Y64_1;
	wire w_dff_A_CpQPaSC28_1;
	wire w_dff_A_BTgskNrm5_1;
	wire w_dff_A_4IMIwSgI0_1;
	wire w_dff_A_8XtrJMHW8_1;
	wire w_dff_A_FXU8MAlH3_1;
	wire w_dff_A_pfxgqJCX4_1;
	wire w_dff_A_nNkPY3zj6_1;
	wire w_dff_A_2CeUZ8G02_1;
	wire w_dff_A_mRi2UOy46_1;
	wire w_dff_A_bxcvZCMb8_1;
	wire w_dff_A_ELfkE1sR4_1;
	wire w_dff_A_SzNhROO54_1;
	wire w_dff_A_YKcXgaSB9_1;
	wire w_dff_A_2h3sDGq20_0;
	wire w_dff_A_xQp4L2oT1_0;
	wire w_dff_A_lP7LBitw2_0;
	wire w_dff_A_NeiOiegw4_0;
	wire w_dff_A_YCAS7qFR3_0;
	wire w_dff_A_aVVmcqqy9_0;
	wire w_dff_A_xqJnR9AY2_0;
	wire w_dff_A_5pBWwoNE3_0;
	wire w_dff_A_3Y0zYfS50_0;
	wire w_dff_A_QA8uoGzG6_0;
	wire w_dff_A_Ei0Pduxf5_0;
	wire w_dff_A_AzQzgRyV6_0;
	wire w_dff_A_tVVeXCWX9_0;
	wire w_dff_A_M04ERNrn8_0;
	wire w_dff_A_DURmX0lG4_0;
	wire w_dff_A_HshRxNag0_0;
	wire w_dff_A_qnv7e2B19_0;
	wire w_dff_A_M68AdHPb8_0;
	wire w_dff_A_IHcVICTS5_0;
	wire w_dff_B_tus5eRkm1_1;
	wire w_dff_B_eAXF9DqD6_1;
	wire w_dff_B_gyQ2zbRa9_1;
	wire w_dff_A_tuc5fw9a7_0;
	wire w_dff_A_IS805HAQ7_0;
	wire w_dff_A_UFxIPcbP1_0;
	wire w_dff_A_yetBByJb6_0;
	wire w_dff_A_ZQPQV9Ht5_0;
	wire w_dff_A_fDVTvTrs4_0;
	wire w_dff_A_LR0mbwcR8_0;
	wire w_dff_A_WnKG3TWf8_0;
	wire w_dff_A_x4xG804r2_0;
	wire w_dff_A_rXbJPyvP6_0;
	wire w_dff_A_YUovUFfc3_0;
	wire w_dff_A_oDpyawyB1_0;
	wire w_dff_A_J66xRmJJ2_0;
	wire w_dff_A_bvfMJeKd6_0;
	wire w_dff_A_qbs6oP5o0_0;
	wire w_dff_A_mMtwPRWV7_0;
	wire w_dff_A_9hRxczGh1_0;
	wire w_dff_A_2OlbOgEd7_0;
	wire w_dff_A_U03xe2o77_0;
	wire w_dff_B_Yv1yDio26_1;
	wire w_dff_B_GMRm2J0a2_1;
	wire w_dff_A_DgLoT3Cl6_0;
	wire w_dff_A_EeUnnpzw5_0;
	wire w_dff_A_heQPLmxD8_0;
	wire w_dff_A_HhlvpK5i5_2;
	wire w_dff_A_8J2edwd05_2;
	wire w_dff_A_wEhkXbVQ8_1;
	wire w_dff_A_hoEmSdRR5_1;
	wire w_dff_A_Yqac6JF91_1;
	wire w_dff_A_cQq5FWtM1_1;
	wire w_dff_A_kkyJwqUr4_1;
	wire w_dff_A_MVluvxhh8_1;
	wire w_dff_A_JqRgh5A39_1;
	wire w_dff_A_XAPlT4QL3_1;
	wire w_dff_A_uH5x4HXz4_1;
	wire w_dff_A_JDkxCPk02_1;
	wire w_dff_A_EU9PD6dJ6_1;
	wire w_dff_A_nlTJAkyk4_1;
	wire w_dff_A_ihrt3K1E9_1;
	wire w_dff_A_Xijo1cgG4_1;
	wire w_dff_A_dkJWDnAp9_1;
	wire w_dff_A_28sMcNK85_1;
	wire w_dff_A_OMaqpi0d6_1;
	wire w_dff_A_j1cVR0RX7_1;
	wire w_dff_A_ks5Qe54q5_1;
	wire w_dff_A_4dWtdapo3_1;
	wire w_dff_A_zpqqx4lL9_1;
	wire w_dff_A_xLymxBEh4_1;
	wire w_dff_A_FquwOoCd0_1;
	wire w_dff_A_JIc1SOCK2_1;
	wire w_dff_A_GqDk9loR0_0;
	wire w_dff_A_4Le9nGDZ9_0;
	wire w_dff_A_OS89iIST8_0;
	wire w_dff_A_MBUxQrmc6_0;
	wire w_dff_A_oFywIdMs1_0;
	wire w_dff_A_GRSvb2ma3_0;
	wire w_dff_A_VLOtDGPW1_0;
	wire w_dff_A_5ucflLL96_0;
	wire w_dff_A_zZEu0zwH3_0;
	wire w_dff_A_s0PqEE7h4_0;
	wire w_dff_A_bsGkyXTe7_0;
	wire w_dff_A_3b34rWmF2_0;
	wire w_dff_A_zJq1VtZc4_0;
	wire w_dff_A_66Rg3Y1y9_0;
	wire w_dff_A_ScUGOy2X8_0;
	wire w_dff_A_dKUNbawA1_0;
	wire w_dff_A_a5IIealN0_0;
	wire w_dff_A_uNdcLaJw2_0;
	wire w_dff_A_Nm6jfFKM7_0;
	wire w_dff_A_ONH35l2Y7_0;
	wire w_dff_A_99OCfEXo9_0;
	wire w_dff_A_NTePZsvj2_0;
	wire w_dff_A_7x6e1Cwz1_2;
	wire w_dff_A_h0mCwTHF4_2;
	wire w_dff_A_a2L6b9wV5_2;
	wire w_dff_A_RIidhpSp9_2;
	wire w_dff_A_FUPkHfDt6_2;
	wire w_dff_A_Z8wG2pGa3_2;
	wire w_dff_A_3nBVnkpo2_2;
	wire w_dff_A_y1aQQWlZ6_2;
	wire w_dff_A_1vWIW1Rv9_2;
	wire w_dff_A_UpnmtUR61_2;
	wire w_dff_A_99gaBX5H7_2;
	wire w_dff_A_SJJq44Bw8_2;
	wire w_dff_A_uc3cELp54_2;
	wire w_dff_A_s8lCTllk8_2;
	wire w_dff_A_17Tjddwp7_2;
	wire w_dff_A_tNy0GlAU6_2;
	wire w_dff_A_zr4HOGbH2_2;
	wire w_dff_A_zVRQU6PJ5_2;
	wire w_dff_A_t0EtXzjT4_2;
	wire w_dff_A_dymjYP6Y2_2;
	wire w_dff_A_E2nBjFEw2_2;
	wire w_dff_A_SKdSkvRK0_2;
	wire w_dff_A_oyn8YtEy2_2;
	wire w_dff_B_tvoDF4FO0_0;
	wire w_dff_B_0RG5tioS2_0;
	wire w_dff_A_tpcB4Xpz7_1;
	wire w_dff_A_kyLWR7fF2_1;
	wire w_dff_A_WCVFLqku1_2;
	wire w_dff_A_O9ZEuD0F3_2;
	wire w_dff_A_cxp9Ss3B8_1;
	wire w_dff_A_M4kje5Xf9_1;
	wire w_dff_A_6v2Rtka73_1;
	wire w_dff_A_SR3YcPDr8_1;
	wire w_dff_A_PFQbUgFH1_1;
	wire w_dff_A_Th03vIP36_1;
	wire w_dff_A_ZKmtSBG20_1;
	wire w_dff_A_RkLwn8DP2_1;
	wire w_dff_A_TTpxHY2E4_1;
	wire w_dff_A_C2fZkQEP0_1;
	wire w_dff_A_0xmRz43N0_1;
	wire w_dff_A_2RU396mk8_1;
	wire w_dff_A_jNqaqBZC6_1;
	wire w_dff_A_jJlfJYnV6_1;
	wire w_dff_A_jN5FDuS95_1;
	wire w_dff_A_nyXxN85x1_1;
	wire w_dff_A_EZt5qb8B7_1;
	wire w_dff_A_7X9AVkNe8_1;
	wire w_dff_A_iQ8Yl5Ej1_1;
	wire w_dff_A_ROcfoLcr4_1;
	wire w_dff_A_vSmminsJ0_1;
	wire w_dff_A_NUDMmJ1L5_1;
	wire w_dff_A_a5HHw5Zd5_1;
	wire w_dff_A_o38x5oMh6_1;
	wire w_dff_A_VmET2hKb8_1;
	wire w_dff_A_YNAHWE8k5_1;
	wire w_dff_A_y5Wqknl02_1;
	wire w_dff_A_UgbKSko40_1;
	wire w_dff_A_mti1uzGy6_1;
	wire w_dff_B_MQuA8mp51_0;
	wire w_dff_B_i95EsnAB8_0;
	wire w_dff_A_J2I59kpR2_1;
	wire w_dff_A_KfIMhN2W7_1;
	wire w_dff_A_ZJQ3nsOw6_2;
	wire w_dff_A_vtutKMai1_2;
	wire w_dff_A_sRfhcl926_1;
	wire w_dff_A_ihW1BRz73_1;
	wire w_dff_A_XHsNrMzL4_1;
	wire w_dff_A_MCNX1YCM4_1;
	wire w_dff_A_K2FeAn602_1;
	wire w_dff_A_lkVNIif41_1;
	wire w_dff_A_5OAbYRuu6_1;
	wire w_dff_A_m59Tvl0e4_1;
	wire w_dff_A_3B1BqbPB2_1;
	wire w_dff_A_KcalhAAw7_1;
	wire w_dff_A_126Nwlt32_1;
	wire w_dff_A_8gbLF7Hy3_1;
	wire w_dff_A_8R3nUI8J7_1;
	wire w_dff_A_XbsvL4823_1;
	wire w_dff_A_9xyuKzU62_1;
	wire w_dff_A_sqdGKtFa8_1;
	wire w_dff_A_1KBnA3xU1_1;
	wire w_dff_A_JrGpFuJX4_1;
	wire w_dff_A_vkXhnAcW9_1;
	wire w_dff_A_oxU45Yxl4_1;
	wire w_dff_A_XhlpIIz80_1;
	wire w_dff_A_EKDNYNzA3_1;
	wire w_dff_A_S6jx6gYA3_1;
	wire w_dff_A_Z31eQSZF6_1;
	wire w_dff_A_DZZnkvIi2_1;
	wire w_dff_A_9cFfsQxC2_1;
	wire w_dff_A_qogrGZcT3_1;
	wire w_dff_A_O3raPL9z5_1;
	wire w_dff_A_5A8AnfSW3_1;
	wire w_dff_A_PvTO2xKm6_2;
	wire w_dff_A_u8HoK95L0_1;
	wire w_dff_B_s4eA4dZI1_0;
	wire w_dff_B_FXRdcySs7_0;
	wire w_dff_B_1p7mmdux0_2;
	wire w_dff_B_JpelzHeC9_2;
	wire w_dff_A_M8I6GfXi6_0;
	wire w_dff_A_NQpzEZHc9_0;
	wire w_dff_A_ihlNcuCP0_0;
	wire w_dff_A_hBAC02z23_0;
	wire w_dff_A_cjpTw9ug5_1;
	wire w_dff_B_VNDBVOTU3_2;
	wire w_dff_B_RtRPpRmP0_2;
	wire w_dff_B_VqLeReC87_2;
	wire w_dff_B_La6GKKE27_2;
	wire w_dff_A_HnBWU2jf4_1;
	wire w_dff_A_1Vt5rRGr6_1;
	wire w_dff_A_Dgt347V98_1;
	wire w_dff_A_aLjvMWy45_1;
	wire w_dff_A_nwifDyRU6_1;
	wire w_dff_A_M8CUetKr4_1;
	wire w_dff_A_UffxN78d5_1;
	wire w_dff_A_p7TklzM11_1;
	wire w_dff_A_lu1XPUva1_1;
	wire w_dff_A_xUke9Sjr9_1;
	wire w_dff_A_N7g21i1s1_1;
	wire w_dff_A_ZS28p3fN6_1;
	wire w_dff_A_76zefZ4f4_1;
	wire w_dff_A_hVXxn5s43_1;
	wire w_dff_A_vvj5LD029_1;
	wire w_dff_A_FR1jVPtN9_1;
	wire w_dff_A_6A0JHep92_1;
	wire w_dff_A_0VlJsJY14_1;
	wire w_dff_A_IBc3Xsp34_1;
	wire w_dff_A_VlQXuF739_1;
	wire w_dff_A_zq2jNuoz6_1;
	wire w_dff_A_BWZ39dDq9_1;
	wire w_dff_A_xPtfVNsz4_1;
	wire w_dff_A_Bu5drJXT4_1;
	wire w_dff_A_z48JbY1H5_1;
	wire w_dff_A_4UQNzWyN7_1;
	wire w_dff_A_TYg8Tdpr4_0;
	wire w_dff_A_jMkhOUGu5_0;
	wire w_dff_A_9ygve7a99_0;
	wire w_dff_A_bDWqOgy68_0;
	wire w_dff_A_4wlQ1R3V9_0;
	wire w_dff_A_h1X0O4xv7_0;
	wire w_dff_A_3zzVk0uX3_0;
	wire w_dff_A_RI2R0slG6_0;
	wire w_dff_A_aZaxS6Bx2_0;
	wire w_dff_A_H1S0Lj2M4_0;
	wire w_dff_A_GRgmCoC55_0;
	wire w_dff_A_qQkC2sPC0_0;
	wire w_dff_A_hEXqIV035_0;
	wire w_dff_A_CAsVwaVG4_0;
	wire w_dff_A_ntPRJ1Yt2_0;
	wire w_dff_A_UfHD95A03_0;
	wire w_dff_A_xwjjFYpY0_0;
	wire w_dff_A_HY38IcR00_0;
	wire w_dff_A_lgy4JPt34_0;
	wire w_dff_A_vL5RymjX7_0;
	wire w_dff_A_dhVN3lCB6_0;
	wire w_dff_A_prACCyXJ7_0;
	wire w_dff_A_rz6XL2OO5_0;
	wire w_dff_A_u4ZDMtqK4_0;
	wire w_dff_A_28w2Jigz5_0;
	wire w_dff_A_cP91ZrdY0_0;
	wire w_dff_A_ADIvEDMc5_0;
	wire w_dff_A_NO57E4si4_0;
	wire w_dff_A_31WWWRHU3_1;
	wire w_dff_A_1aLQFsMz9_1;
	wire w_dff_A_QVBtoqvc1_1;
	wire w_dff_A_xC4ZM0WA6_2;
	wire w_dff_A_QF1WnZsW7_2;
	wire w_dff_A_Dujt7ChK9_2;
	wire w_dff_A_iJUqX09N6_2;
	wire w_dff_A_g2m1xBFl8_1;
	wire w_dff_A_B0oME9l07_1;
	wire w_dff_A_9jqs9Xlx5_1;
	wire w_dff_A_uaDqfkQw2_1;
	wire w_dff_A_IvlrDlFz0_1;
	wire w_dff_A_vWMoivkc3_1;
	wire w_dff_A_OU0AZkxh6_1;
	wire w_dff_A_hOFzT9tM4_1;
	wire w_dff_A_kXitvI2w6_1;
	wire w_dff_A_kEHsHiiy8_1;
	wire w_dff_A_igPE98EO4_1;
	wire w_dff_A_MdzvNzrV6_1;
	wire w_dff_A_FhSiNrK38_1;
	wire w_dff_A_aH8OxooQ2_1;
	wire w_dff_A_Qu7i0AOX5_1;
	wire w_dff_A_KUTh1DLr8_1;
	wire w_dff_A_Ua2Ycfdy6_1;
	wire w_dff_A_gHT68AVI8_1;
	wire w_dff_A_qNbB8PSW1_1;
	wire w_dff_A_pmqbbcJL1_1;
	wire w_dff_A_X9cBIOx54_1;
	wire w_dff_A_5Z81xz2U1_2;
	wire w_dff_A_LnyJASmM1_2;
	wire w_dff_A_j0ldxZUh0_2;
	wire w_dff_A_HIduge0I7_2;
	wire w_dff_A_l6iDbYvx2_2;
	wire w_dff_B_ROfqi5sd5_1;
	wire w_dff_A_r9uNt09E4_0;
	wire w_dff_A_rkdl9ovW0_0;
	wire w_dff_A_RK9WZi2Q1_0;
	wire w_dff_A_43ymp5HH0_0;
	wire w_dff_A_PlUjBCk18_0;
	wire w_dff_A_nalhsrNs8_0;
	wire w_dff_A_gTodIcZt1_0;
	wire w_dff_A_0c4x3L2H1_0;
	wire w_dff_A_8Wunz3Gz6_0;
	wire w_dff_A_F96IB2Yj5_0;
	wire w_dff_A_cVlb8Lai2_0;
	wire w_dff_A_q4kPMBVf3_0;
	wire w_dff_A_7ecolecs9_0;
	wire w_dff_A_dLJrDbS01_0;
	wire w_dff_A_YNLs3Fpt1_0;
	wire w_dff_A_nWYj38gu5_0;
	wire w_dff_A_fjHQlS0k7_0;
	wire w_dff_A_FmFN1t1E6_0;
	wire w_dff_A_07zxERxa6_0;
	wire w_dff_A_hE3TMeAi0_0;
	wire w_dff_A_vf7Phuzu2_0;
	wire w_dff_A_1k4KbDb68_0;
	wire w_dff_A_wAN75iSl7_0;
	wire w_dff_A_YRBUIWw11_0;
	wire w_dff_A_9lgaDUz22_0;
	wire w_dff_A_HkY0Ozwo5_0;
	wire w_dff_A_pC9SxTcg1_0;
	wire w_dff_A_wPtHeeCc1_0;
	wire w_dff_A_3ZpI47qr9_1;
	wire w_dff_A_bFQNGcgB9_1;
	wire w_dff_A_MZshv5gh3_1;
	wire w_dff_A_TwH1swP31_1;
	wire w_dff_A_8HORNGw25_1;
	wire w_dff_A_xFMB9gpv5_1;
	wire w_dff_A_5NdSYsBJ7_1;
	wire w_dff_A_vcR82Vn03_1;
	wire w_dff_A_reVZ7qnZ6_1;
	wire w_dff_A_DrHrwRI04_1;
	wire w_dff_A_tbLMEGHm9_1;
	wire w_dff_A_0u21JPMa1_1;
	wire w_dff_A_9W78x3VH4_1;
	wire w_dff_A_oHtssPdj0_1;
	wire w_dff_A_C2oswGKJ7_1;
	wire w_dff_A_ez8dfd7Z7_1;
	wire w_dff_A_V8dlpBUk4_1;
	wire w_dff_A_y6e35GZE3_1;
	wire w_dff_A_YErLJ0Y63_1;
	wire w_dff_A_JWPlhfRX4_1;
	wire w_dff_A_oghk7Wwo4_1;
	wire w_dff_A_ZE5QrrRW7_1;
	wire w_dff_A_jiaZanyy9_1;
	wire w_dff_A_qTxX4T0S2_1;
	wire w_dff_A_Ni3xbxCS0_1;
	wire w_dff_A_D5Uy5jKu4_1;
	wire w_dff_A_6Hqpq9og1_1;
	wire w_dff_A_hi7zk1CR7_1;
	wire w_dff_A_LF35YLmI6_1;
	wire w_dff_A_zcRclED08_1;
	wire w_dff_A_fJ6Z2Fym0_1;
	wire w_dff_A_H6YW1Fir0_1;
	wire w_dff_A_ELfZLHUX2_1;
	wire w_dff_A_tbc2fNk24_2;
	wire w_dff_A_ZO8xir4g0_2;
	wire w_dff_A_llcSN2BG4_2;
	wire w_dff_A_pUa3w54x3_2;
	wire w_dff_A_g3dRlHVv4_2;
	wire w_dff_A_4iMejImJ9_2;
	wire w_dff_A_9WxyhcV15_2;
	wire w_dff_B_4ktNGoya8_0;
	wire w_dff_B_W1sljb7y0_0;
	wire w_dff_A_K55uznzv1_1;
	wire w_dff_A_JnxynNQZ7_1;
	wire w_dff_A_iSt3pmoL4_2;
	wire w_dff_A_fzA0RuAB8_2;
	wire w_dff_A_62mwjYD83_1;
	wire w_dff_A_KHSdDUvG7_1;
	wire w_dff_A_WpstJHKE4_1;
	wire w_dff_A_cqRjat6f7_1;
	wire w_dff_A_tqesnuAW6_1;
	wire w_dff_B_1NhAGwVz7_0;
	wire w_dff_B_K5txonfB4_3;
	wire w_dff_B_ZTy8EqPV4_3;
	wire w_dff_A_MbeNTaRo8_2;
	wire w_dff_A_VqFYbCB53_2;
	wire w_dff_A_tg13M2sT7_2;
	wire w_dff_A_6XrtcXTY6_2;
	wire w_dff_A_jPNMqTsu8_2;
	wire w_dff_A_iMez3pks7_2;
	wire w_dff_A_ZwyOmiDg8_2;
	wire w_dff_A_1pWxHSlY1_2;
	wire w_dff_A_JDyQ9ai18_2;
	wire w_dff_A_iR6B7duH2_2;
	wire w_dff_A_OaDpa0iQ4_2;
	wire w_dff_A_dyS1aMqS3_2;
	wire w_dff_A_6pCGcHdt6_2;
	wire w_dff_A_yYbDhjX34_2;
	wire w_dff_A_hQ8yQrNP2_2;
	wire w_dff_A_41mxgmIB7_2;
	wire w_dff_A_pYHGwCkf2_2;
	wire w_dff_A_2D8usgXT5_2;
	wire w_dff_A_hYOCOZMz8_2;
	wire w_dff_A_FQOKUYsv5_2;
	wire w_dff_A_BfJp3bsu6_2;
	wire w_dff_A_yOGMEFVi3_2;
	wire w_dff_B_bEDm3zYn1_1;
	wire w_dff_B_BiI0ZTCU1_1;
	wire w_dff_A_wjKWvZBb3_0;
	wire w_dff_A_dJgKxRIC5_0;
	wire w_dff_A_1ZBRyKC30_0;
	wire w_dff_A_cVv02Nlj1_0;
	wire w_dff_A_rRkeo3GP2_0;
	wire w_dff_A_bldm7o9G6_0;
	wire w_dff_A_sBerXbpX6_0;
	wire w_dff_A_kEVfi8W48_0;
	wire w_dff_A_itbCi6411_0;
	wire w_dff_A_ePQy4ze88_0;
	wire w_dff_A_gpQCK13v9_0;
	wire w_dff_A_VgxrRdz78_0;
	wire w_dff_A_2ObhRrl09_0;
	wire w_dff_A_2D63Mkir0_0;
	wire w_dff_A_ssscaKOB5_0;
	wire w_dff_A_YYVbMTHo0_0;
	wire w_dff_A_YoUP7csR4_0;
	wire w_dff_A_RHxQU68j4_0;
	wire w_dff_A_Ol441Uz21_0;
	wire w_dff_A_bxayRSXS9_0;
	wire w_dff_A_KChkSnBZ2_0;
	wire w_dff_A_YDSTlRFl9_0;
	wire w_dff_B_pVUVu6oE9_1;
	wire w_dff_B_VEsaFXyh2_1;
	wire w_dff_B_2P3d0CEE3_1;
	wire w_dff_A_Yx4risHu8_1;
	wire w_dff_A_LPyXdJn96_1;
	wire w_dff_A_YRV2LOo14_1;
	wire w_dff_A_jPrX1cbm8_1;
	wire w_dff_A_BQ09mqDV6_1;
	wire w_dff_A_hnGbZB4c2_1;
	wire w_dff_A_LoWAeYgW8_1;
	wire w_dff_A_aga1Qr7U6_1;
	wire w_dff_A_E6b3rdbL2_1;
	wire w_dff_A_H2JKbEBc0_1;
	wire w_dff_A_tHGxxEfW7_1;
	wire w_dff_A_SV50TXc59_1;
	wire w_dff_A_ZCa0qgEb5_1;
	wire w_dff_A_seWYdYZu5_1;
	wire w_dff_A_esdau1Ez5_1;
	wire w_dff_A_88KGpDJV7_1;
	wire w_dff_A_sKYU1zDx5_1;
	wire w_dff_A_o83YnuwY8_1;
	wire w_dff_A_Tp2bWoNb3_1;
	wire w_dff_A_hXMuAwq23_1;
	wire w_dff_A_aNHrWs2m3_1;
	wire w_dff_A_DCRuM31d7_1;
	wire w_dff_A_cYntFtSi4_1;
	wire w_dff_A_kiwYSKer5_1;
	wire w_dff_A_DBXmQNFG7_1;
	wire w_dff_A_7PWrwykw5_1;
	wire w_dff_A_tVTt4gd04_1;
	wire w_dff_A_gLGe0Teh8_1;
	wire w_dff_A_9zluSdTd1_1;
	wire w_dff_A_tlvcJgdQ4_1;
	wire w_dff_A_SJerHwCp5_1;
	wire w_dff_A_O0RnGL9Z6_1;
	wire w_dff_A_8c5mLC0Q5_1;
	wire w_dff_A_iUP3jbLH0_1;
	wire w_dff_A_iLH3P6Ny7_1;
	wire w_dff_A_iraFo22z3_1;
	wire w_dff_A_BIz3xtaL1_1;
	wire w_dff_A_9wo9M0UM2_1;
	wire w_dff_A_ZlWK9vG67_1;
	wire w_dff_A_mrAwvEfd2_1;
	wire w_dff_A_RW5hLxVc4_1;
	wire w_dff_A_5WviFnyq4_1;
	wire w_dff_A_Pmjqmfgp6_1;
	wire w_dff_A_cW8swT584_1;
	wire w_dff_A_yiEcr5Fi0_1;
	wire w_dff_A_7fMavj4h1_1;
	wire w_dff_A_kMawKvbe0_1;
	wire w_dff_A_Wj9KDVlV5_1;
	wire w_dff_A_GxaZnX183_1;
	wire w_dff_A_Wdxvnsr97_1;
	wire w_dff_A_nRvZGQid1_1;
	wire w_dff_A_vlI9QMAP8_1;
	wire w_dff_A_mfUBjL8h2_1;
	wire w_dff_A_jGvha8wF0_2;
	wire w_dff_A_kggdpM1j0_0;
	wire w_dff_A_0oJUP1386_0;
	wire w_dff_A_k5pLKUhv3_0;
	wire w_dff_A_mJqz6rnL6_0;
	wire w_dff_A_PDW4LpkL6_0;
	wire w_dff_A_OmW5Xfae5_0;
	wire w_dff_A_EA2hOLsY0_0;
	wire w_dff_A_WbU7slYa3_0;
	wire w_dff_A_d7qouoRC9_0;
	wire w_dff_A_1P1smI3R2_0;
	wire w_dff_A_Fg6V4p2y1_0;
	wire w_dff_A_ydOLMp6N6_0;
	wire w_dff_A_EmUjLuic3_0;
	wire w_dff_A_LUvcrnHy4_0;
	wire w_dff_A_QTbTcMfe2_0;
	wire w_dff_A_xjM7abYy4_0;
	wire w_dff_A_g46lyfAZ5_0;
	wire w_dff_A_AiEyQROX8_0;
	wire w_dff_A_XEDLWGuX6_0;
	wire w_dff_A_S0iiNFFp4_0;
	wire w_dff_A_sXogL2F34_0;
	wire w_dff_A_Hf4XiKpk9_0;
	wire w_dff_A_gl02tlid9_0;
	wire w_dff_A_2G7fOMRi7_0;
	wire w_dff_A_b9i0mVPX4_0;
	wire w_dff_A_387xNCBw7_1;
	wire w_dff_A_mTJizaas6_1;
	wire w_dff_A_eBFFZHSR0_1;
	wire w_dff_A_m7l1VNKy0_1;
	wire w_dff_A_lbqrYRH56_1;
	wire w_dff_A_2RPepJyl2_1;
	wire w_dff_A_vsDihIaw3_1;
	wire w_dff_A_HR0oxJQG8_1;
	wire w_dff_A_euFO73gY0_1;
	wire w_dff_A_y5wHyyBy4_1;
	wire w_dff_A_bTwg9hed6_1;
	wire w_dff_A_PUmlXlX87_1;
	wire w_dff_A_Tmg5YTKb6_1;
	wire w_dff_A_z8vE3lil5_1;
	wire w_dff_A_Uu017SPj2_1;
	wire w_dff_A_SMs7wOsT4_1;
	wire w_dff_A_ozyoaQiE6_1;
	wire w_dff_A_ItrCI28u1_1;
	wire w_dff_A_LY8xMpdE4_1;
	wire w_dff_A_w6LFbHZM6_1;
	wire w_dff_A_ydoMcFHd3_1;
	wire w_dff_A_zMW1l7rV8_1;
	wire w_dff_A_pWMSAPij5_1;
	wire w_dff_A_ERRnKHiM3_1;
	wire w_dff_A_GVpSceM11_1;
	wire w_dff_A_R1lrvgxA0_1;
	wire w_dff_A_ixPLp55g3_0;
	wire w_dff_A_Dxy3LhG70_0;
	wire w_dff_B_wEA3Mhyp8_0;
	wire w_dff_B_q2wugx5I4_2;
	wire w_dff_B_59IVopTg7_2;
	wire w_dff_A_3wBuw7q61_2;
	wire w_dff_A_nKOwR62T0_2;
	wire w_dff_A_AUMhxIV25_2;
	wire w_dff_A_LcmCCn9p0_2;
	wire w_dff_A_pAmu6KRT6_0;
	wire w_dff_A_BdNNkt7t5_0;
	wire w_dff_A_GVtHqrqw2_0;
	wire w_dff_A_zema3Pci6_0;
	wire w_dff_A_pbkPyzqZ3_0;
	wire w_dff_A_1snCvRQM9_0;
	wire w_dff_A_fvnDjC625_0;
	wire w_dff_A_u8A8dzar6_0;
	wire w_dff_A_xPZ30kMI6_0;
	wire w_dff_A_igY3nnvL2_0;
	wire w_dff_A_F5ZTxqAJ1_0;
	wire w_dff_A_MTgprWJy7_0;
	wire w_dff_A_G0bKuq5s8_0;
	wire w_dff_A_RYW8Liwf4_0;
	wire w_dff_A_NOoDreEn2_0;
	wire w_dff_A_jnJX9vzc5_0;
	wire w_dff_A_sH9JF1vV8_0;
	wire w_dff_A_NrXAo8iN2_0;
	wire w_dff_A_KCGuJm2B2_0;
	wire w_dff_A_kfLL1v7W8_0;
	wire w_dff_A_GgfWM8fP3_0;
	wire w_dff_A_Qqjm0Ki83_0;
	wire w_dff_A_2aihjCnZ1_0;
	wire w_dff_A_elxtFNZ21_0;
	wire w_dff_A_c7ZQRUbS3_0;
	wire w_dff_A_Ar18Dr8B6_0;
	wire w_dff_A_cd83q31D9_0;
	wire w_dff_A_OuOmfGs39_0;
	wire w_dff_A_UYjlfQK17_2;
	wire w_dff_A_YLcjpomc1_2;
	wire w_dff_A_yvXqhH371_2;
	wire w_dff_A_ky3EWdLW5_2;
	wire w_dff_A_9FBXsJ5D7_0;
	wire w_dff_A_rZYiXbkz5_0;
	wire w_dff_B_F1xHy1Kr0_0;
	wire w_dff_B_aLOuqT6y1_2;
	wire w_dff_B_qfxNow3q4_2;
	wire w_dff_A_09Rzbv0n9_1;
	wire w_dff_A_zEQnSkvr7_1;
	wire w_dff_A_xGnoXxZc2_1;
	wire w_dff_A_sg9lbXIo8_1;
	wire w_dff_A_H6LTrRNq3_1;
	wire w_dff_A_suG4h3MQ2_1;
	wire w_dff_A_XwqpMb7r3_1;
	wire w_dff_A_gr4pZuZk5_1;
	wire w_dff_A_Zezn3gTG3_1;
	wire w_dff_A_79D3nSYZ5_1;
	wire w_dff_A_0m4mJ7o25_1;
	wire w_dff_A_RMSrkFxh6_1;
	wire w_dff_A_CmqjsdPN6_1;
	wire w_dff_A_fll1kGTT8_1;
	wire w_dff_A_4E0of3rE9_1;
	wire w_dff_A_moFGrM1t2_1;
	wire w_dff_A_Mjxs4LXI1_1;
	wire w_dff_A_36A6DOYl2_1;
	wire w_dff_A_zF5Nd7pD3_1;
	wire w_dff_A_RwvSeBfy3_1;
	wire w_dff_A_5gnAqyom9_1;
	wire w_dff_A_DhltJnR27_1;
	wire w_dff_A_cPYjnrig9_1;
	wire w_dff_A_hrEXM8FB1_1;
	wire w_dff_A_xddUA2Jw4_1;
	wire w_dff_A_cXhmlniw5_1;
	wire w_dff_A_1Ymh6j8A3_1;
	wire w_dff_A_YUTW2DAO3_1;
	wire w_dff_A_9gVNd9nX7_2;
	wire w_dff_A_4arLlfmD9_0;
	wire w_dff_A_Etqypq3F7_0;
	wire w_dff_B_8UG59Vca7_0;
	wire w_dff_A_QX1Bx6I01_1;
	wire w_dff_A_Ggj1yM443_1;
	wire w_dff_A_HTMGDVHZ1_2;
	wire w_dff_A_K5ZBCKeC9_2;
	wire w_dff_A_DY0byoKN3_1;
	wire w_dff_A_poaqWqFO4_1;
	wire w_dff_A_otUmM6eA6_1;
	wire w_dff_A_Pn0AJcb18_1;
	wire w_dff_A_baD3Q3CB8_1;
	wire w_dff_A_1R9bhMXu3_1;
	wire w_dff_A_wWKFtqNt8_1;
	wire w_dff_A_71pj1lpB6_1;
	wire w_dff_A_ryRSPHHA3_1;
	wire w_dff_A_KavIGZoi1_1;
	wire w_dff_A_OjjPaYin5_1;
	wire w_dff_A_49iVaXPm4_1;
	wire w_dff_A_uL3r89oo2_1;
	wire w_dff_A_K5wvCeqg4_1;
	wire w_dff_A_8GZUAg3f1_1;
	wire w_dff_A_y6Lu6vUt2_1;
	wire w_dff_A_yWVwfS0b3_1;
	wire w_dff_A_uSkAOhDH6_1;
	wire w_dff_A_yh9jPnZQ7_1;
	wire w_dff_A_CAjnkr406_1;
	wire w_dff_A_bZpG9w7x0_1;
	wire w_dff_A_3nTGLdvQ8_1;
	wire w_dff_A_Tqr5ye7V0_1;
	wire w_dff_A_MrxSu1Kd1_1;
	wire w_dff_A_z8TgFc517_1;
	wire w_dff_A_iYFIVBXd1_1;
	wire w_dff_A_CKmlYBeT8_1;
	wire w_dff_A_Lq8qeYY98_1;
	wire w_dff_A_AY0Ygbpn0_1;
	wire w_dff_A_tR2DfjdY3_1;
	wire w_dff_A_udk0DvfK8_1;
	wire w_dff_A_fHouZqGt3_1;
	wire w_dff_A_C5gFqW8C7_2;
	wire w_dff_A_AzhajSGA9_2;
	wire w_dff_A_anWRxKrp5_2;
	wire w_dff_A_CEBS9loZ4_2;
	wire w_dff_A_zWpz9K373_2;
	wire w_dff_A_tS34ImiE8_2;
	wire w_dff_A_i9BEr20I3_2;
	wire w_dff_A_6BNDKbQJ5_2;
	wire w_dff_A_wHvaS5eP5_2;
	wire w_dff_A_2UJBnGw15_2;
	wire w_dff_A_YHYPlSnV9_2;
	wire w_dff_A_NmpRpQDc7_2;
	wire w_dff_A_IIb8Gdv16_2;
	wire w_dff_A_QwKkJGS42_2;
	wire w_dff_A_FpE1NfNw5_2;
	wire w_dff_A_ZAXYdkzJ8_2;
	wire w_dff_A_b3I5VCR79_2;
	wire w_dff_A_M8tnH8qC1_2;
	wire w_dff_A_TzFzFNrV6_2;
	wire w_dff_A_xkqkMJMN6_2;
	wire w_dff_A_jvauE3K24_2;
	wire w_dff_A_QQKBQqh65_2;
	wire w_dff_A_tUUVP2Vy9_2;
	wire w_dff_A_BHs6HxvU7_2;
	wire w_dff_A_VmcHDvd72_2;
	wire w_dff_A_U6iUWgwA8_2;
	wire w_dff_A_FNcJlQLL3_2;
	wire w_dff_A_wqPvJ2r96_2;
	wire w_dff_A_JPCot2ZB7_1;
	wire w_dff_A_L7qavIXQ2_1;
	wire w_dff_A_AbUAfjVv8_1;
	wire w_dff_A_0vjlAh087_1;
	wire w_dff_A_rbzNotZQ9_1;
	wire w_dff_A_LIx7qTrD6_1;
	wire w_dff_A_TH2h2Jyo1_1;
	wire w_dff_A_63KIUd6P4_1;
	wire w_dff_A_LytSijHB7_1;
	wire w_dff_A_T6Pw4CQE5_1;
	wire w_dff_A_FecUEcXq0_1;
	wire w_dff_A_jfqI3rik3_1;
	wire w_dff_A_2VydCtZr7_1;
	wire w_dff_A_RwDE5Bnv0_1;
	wire w_dff_A_3wkFOEgy6_1;
	wire w_dff_A_r1jNPOol5_1;
	wire w_dff_A_qv6uDbQW6_1;
	wire w_dff_A_IxbBvkpg9_1;
	wire w_dff_A_nM5uXi1V4_1;
	wire w_dff_A_xs1WsFzi4_1;
	wire w_dff_A_h2OQWkcC5_1;
	wire w_dff_A_ZW4vS40h0_1;
	wire w_dff_A_BrYgqhBT2_1;
	wire w_dff_A_WVcPQJbm0_1;
	wire w_dff_A_lFLkfp0b5_1;
	wire w_dff_A_y8sCxpDE5_1;
	wire w_dff_A_vKkxQUhC6_1;
	wire w_dff_A_mXJSl3Zk9_1;
	wire w_dff_A_6GHje0Ez4_1;
	wire w_dff_A_HvRZD6YI7_0;
	wire w_dff_A_3oLcbMUW2_0;
	wire w_dff_B_KrwkUrhI8_0;
	wire w_dff_A_GKk1bp1A7_1;
	wire w_dff_A_J5y6YU0r4_1;
	wire w_dff_A_dIpyqVQs2_2;
	wire w_dff_A_fzPZDmtX3_2;
	wire w_dff_A_bUrptudo5_1;
	wire w_dff_A_aAH0WpaF9_1;
	wire w_dff_A_lNPuLJKy0_1;
	wire w_dff_A_8RIx3fbU2_1;
	wire w_dff_A_40hxMOXx5_1;
	wire w_dff_A_Tfq0k3aS0_1;
	wire w_dff_A_rLdU8sJG5_1;
	wire w_dff_A_GsibDraX6_1;
	wire w_dff_A_QlKpmL7l1_1;
	wire w_dff_A_idxDFid54_1;
	wire w_dff_A_pFynIBHc3_1;
	wire w_dff_A_KylSvzqG0_1;
	wire w_dff_A_JRn941Bw9_1;
	wire w_dff_A_hnYhUgvT6_1;
	wire w_dff_A_bKtJ0jLs3_1;
	wire w_dff_A_Lf6bnXpT7_1;
	wire w_dff_A_EsfkNbea7_1;
	wire w_dff_A_eRFKiswX8_1;
	wire w_dff_A_sHTJBg2x2_1;
	wire w_dff_A_zBdsHkwr0_1;
	wire w_dff_A_24gcnJs55_1;
	wire w_dff_A_2yoa0Xmg3_1;
	wire w_dff_A_I5NxoADI0_1;
	wire w_dff_A_dWsgIMZl3_1;
	wire w_dff_A_W9XIvgWl1_1;
	wire w_dff_A_5avsFQRR6_1;
	wire w_dff_A_huoydXMQ2_1;
	wire w_dff_A_hYt7MMz02_1;
	wire w_dff_A_NlVCp1mj4_1;
	wire w_dff_A_O4cQ5JZr6_1;
	wire w_dff_A_SKbTFCZj2_1;
	wire w_dff_A_1zVdYsML7_1;
	wire w_dff_A_rGde2L1r5_0;
	wire w_dff_A_zj7Wtcb85_0;
	wire w_dff_B_vxvT3Qbl3_0;
	wire w_dff_A_ZmpSsmGr0_1;
	wire w_dff_A_DY0VH9bL9_1;
	wire w_dff_A_w1WJmkCq5_2;
	wire w_dff_A_4u7xADtA8_2;
	wire w_dff_A_ob5eTzHp9_2;
	wire w_dff_A_3RoiRSzn7_2;
	wire w_dff_A_1guXg5S94_2;
	wire w_dff_A_lACnqkSy8_2;
	wire w_dff_B_ZagUfvbl0_0;
	wire w_dff_B_wPxDIRJ71_2;
	wire w_dff_B_8TkpM3NK2_2;
	wire w_dff_A_hV1GeVxG4_0;
	wire w_dff_A_B1dGCImi7_0;
	wire w_dff_A_jwPzA63V8_0;
	wire w_dff_A_Ooh0LBXd5_0;
	wire w_dff_B_03bsOFBl3_1;
	wire w_dff_B_65zW7JSU8_1;
	wire w_dff_B_dDmxprc12_1;
	wire w_dff_B_3SWdjrQz8_1;
	wire w_dff_B_lEXq7Dmk5_1;
	wire w_dff_B_q2YQNKPl0_1;
	wire w_dff_B_84g7pzSx1_1;
	wire w_dff_B_UsAZKtNS6_1;
	wire w_dff_B_7H7EWBKK6_1;
	wire w_dff_B_C6KzTMwc7_1;
	wire w_dff_B_r0ROCC9s4_1;
	wire w_dff_B_IjIqbyHH4_1;
	wire w_dff_B_flmF78nX9_1;
	wire w_dff_B_aofrh8mi9_1;
	wire w_dff_B_c6sAlVSH7_1;
	wire w_dff_B_sqaBfIcu0_0;
	wire w_dff_B_Ao6mYGi31_0;
	wire w_dff_B_UuW7iBjA1_0;
	wire w_dff_B_zXwjkqDF0_0;
	wire w_dff_B_WYToY6Qz7_0;
	wire w_dff_B_iiTVZbst1_0;
	wire w_dff_B_dWg3EtNZ9_0;
	wire w_dff_B_2ddakiyz8_0;
	wire w_dff_B_23s7cY9T8_0;
	wire w_dff_B_v0dM5hOn8_0;
	wire w_dff_B_qgka1V8r4_0;
	wire w_dff_B_cVuH9BZP5_1;
	wire w_dff_B_USdYKckw6_1;
	wire w_dff_B_uWWG181A2_0;
	wire w_dff_B_rnq9dnf40_0;
	wire w_dff_B_aqxciPkK8_0;
	wire w_dff_B_zcygb30n6_0;
	wire w_dff_B_jjk4JYtM5_0;
	wire w_dff_B_mORKMFCh6_0;
	wire w_dff_B_zwd4YUXK8_0;
	wire w_dff_A_PAVCvIjB5_0;
	wire w_dff_A_OgBIZFUB7_0;
	wire w_dff_A_mN0ce6hD7_0;
	wire w_dff_A_jWx3Jy360_0;
	wire w_dff_A_sNwyBztz9_0;
	wire w_dff_A_mwdLIJc12_0;
	wire w_dff_A_uzD2hOmg0_0;
	wire w_dff_A_CNVqdke96_1;
	wire w_dff_A_XjAjlG513_1;
	wire w_dff_A_whqrPRhn5_1;
	wire w_dff_A_hZU2Twyh5_1;
	wire w_dff_A_4UNpTZPn2_1;
	wire w_dff_A_bqsqtYaC7_1;
	wire w_dff_A_BGKrLFec7_1;
	wire w_dff_B_uLmvtIRD8_0;
	wire w_dff_B_Rvwz1Ntt5_0;
	wire w_dff_B_I4GYQyWz0_0;
	wire w_dff_B_FFuF2WM68_0;
	wire w_dff_A_eZkA2yIW6_1;
	wire w_dff_A_IjDgqFsP6_1;
	wire w_dff_A_05DUFI563_1;
	wire w_dff_A_WPxaR21L2_1;
	wire w_dff_A_K8H2s6xj3_1;
	wire w_dff_A_MWmQHqrw8_1;
	wire w_dff_A_H227V6P77_1;
	wire w_dff_B_qwYIpRNY4_1;
	wire w_dff_B_oUKrvhW93_1;
	wire w_dff_B_yJorNVda5_1;
	wire w_dff_B_mp19wXpG4_1;
	wire w_dff_B_j7ri32Ll5_1;
	wire w_dff_B_rqgIY5ES8_1;
	wire w_dff_B_EKprS7Q16_0;
	wire w_dff_B_bGDSMlsM5_0;
	wire w_dff_B_CnVb1Lwf1_0;
	wire w_dff_A_TabvV23X2_1;
	wire w_dff_A_vswOw34m7_1;
	wire w_dff_A_M1TycP0p7_1;
	wire w_dff_A_dfIKLkOG9_1;
	wire w_dff_A_DdevqCW49_1;
	wire w_dff_A_MLEKQuC59_1;
	wire w_dff_A_ngUTuCte4_1;
	wire w_dff_A_x3DqQd8p4_1;
	wire w_dff_A_Sg5V6eJQ8_1;
	wire w_dff_A_o9f56Jhc7_1;
	wire w_dff_A_39Do16BY4_1;
	wire w_dff_A_ahBHxoSc6_1;
	wire w_dff_A_n6i6XZTi2_1;
	wire w_dff_A_oWXDgH8R3_1;
	wire w_dff_A_07VbPBFq4_1;
	wire w_dff_B_1eGYARXL9_0;
	wire w_dff_B_JC4Q6jwA2_0;
	wire w_dff_B_wwtBx1AL7_1;
	wire w_dff_B_Zd7shYUE7_1;
	wire w_dff_B_4RDfK5419_1;
	wire w_dff_B_cpxQha6Z2_1;
	wire w_dff_B_kyDp6uk88_1;
	wire w_dff_B_oJVVuy8x8_1;
	wire w_dff_B_SEwrgOtF6_1;
	wire w_dff_B_NudPdGMP0_1;
	wire w_dff_B_tVNopkYn6_1;
	wire w_dff_B_eDtWO0qj3_1;
	wire w_dff_B_hMF0gLGw1_1;
	wire w_dff_B_R7AEYJd50_1;
	wire w_dff_B_eZ81QOBf4_0;
	wire w_dff_A_3BncMQJW6_1;
	wire w_dff_B_4FNzd9Pc5_2;
	wire w_dff_B_24mtxUlb8_2;
	wire w_dff_B_kBZpwD7o1_0;
	wire w_dff_B_hm3K74fN6_0;
	wire w_dff_B_XEqBx23A8_0;
	wire w_dff_B_4xMheUue8_0;
	wire w_dff_B_FkQP94Gv6_0;
	wire w_dff_B_CO0nfNWu6_1;
	wire w_dff_B_QDA88Cd25_1;
	wire w_dff_B_EU2ykJhL3_1;
	wire w_dff_A_h2VvtMUM2_0;
	wire w_dff_A_WMngvtCD5_0;
	wire w_dff_A_mRLmi6Zn1_0;
	wire w_dff_A_W85UgazU7_0;
	wire w_dff_A_9CJyk6me6_1;
	wire w_dff_A_JfAr3Uyd2_1;
	wire w_dff_A_aTcH09wp5_1;
	wire w_dff_A_pHS2QGSq2_1;
	wire w_dff_A_ipZqOBiQ8_1;
	wire w_dff_A_oTx87bls5_1;
	wire w_dff_A_iqqYYH0K0_1;
	wire w_dff_A_vygkvrDe7_1;
	wire w_dff_A_bRsDcaSe0_1;
	wire w_dff_A_TF5cqGEb7_1;
	wire w_dff_A_8IWkgJBx5_1;
	wire w_dff_A_LoRLtfpl3_1;
	wire w_dff_A_UEjyKK6E7_1;
	wire w_dff_A_TR24fotw6_1;
	wire w_dff_A_tVeRf5z89_1;
	wire w_dff_A_mdctKRx36_1;
	wire w_dff_B_uMxn8nPI8_0;
	wire w_dff_B_0VGiGqZB7_0;
	wire w_dff_B_M3G9IcnN5_0;
	wire w_dff_B_mrMzToCv7_0;
	wire w_dff_B_bLVqyfKW6_0;
	wire w_dff_B_d6WT5pj18_0;
	wire w_dff_B_qoeLEU5k2_0;
	wire w_dff_A_qdiTRg3f2_1;
	wire w_dff_A_PVUmlWos8_1;
	wire w_dff_A_reUXqUeJ4_1;
	wire w_dff_A_5EqcL14M4_1;
	wire w_dff_A_HQovdrkH7_1;
	wire w_dff_A_5tmnPJWJ9_1;
	wire w_dff_A_cZzw0s9p4_1;
	wire w_dff_A_VqPGuDRg5_1;
	wire w_dff_A_mnaXM1OV5_1;
	wire w_dff_A_XV4JvTtJ0_1;
	wire w_dff_A_WknRXqOa9_1;
	wire w_dff_A_X0XqqPhE6_1;
	wire w_dff_A_EdZdUDdb8_1;
	wire w_dff_A_NXxsCLP79_1;
	wire w_dff_A_Clg8QBrH5_1;
	wire w_dff_A_JRCBIb8S9_1;
	wire w_dff_A_ML0wQCZb4_1;
	wire w_dff_A_9g0Gj25A9_1;
	wire w_dff_A_WmUiygcc7_1;
	wire w_dff_A_NRvr2xNV3_1;
	wire w_dff_B_XkcTUA521_2;
	wire w_dff_A_FmgsxsHO6_2;
	wire w_dff_B_Wb2jObOc6_1;
	wire w_dff_B_K91H5ioU1_0;
	wire w_dff_A_pdW84Udt4_0;
	wire w_dff_A_KG5akhGz9_0;
	wire w_dff_A_CtKtQLz32_2;
	wire w_dff_A_qIxN32vE1_2;
	wire w_dff_A_9VwgKFyQ5_1;
	wire w_dff_A_Rph632JF4_1;
	wire w_dff_A_ruSKVlVn2_1;
	wire w_dff_A_bdb0wrOh4_1;
	wire w_dff_A_cUYEEm9U4_1;
	wire w_dff_A_Y9db0dxp5_1;
	wire w_dff_A_cAcLb03K7_1;
	wire w_dff_A_VKnKUEpK1_1;
	wire w_dff_A_MH9i3ecq1_1;
	wire w_dff_A_CFcnAxKv8_1;
	wire w_dff_A_3dSPtnlF5_1;
	wire w_dff_A_PlV3Rsls8_1;
	wire w_dff_A_rWD19SEB3_1;
	wire w_dff_A_0q8P4K7e5_1;
	wire w_dff_A_jlJRbxIg0_1;
	wire w_dff_A_VPXYOjKq6_1;
	wire w_dff_A_sLEVuBb67_1;
	wire w_dff_A_PzXjsi4a4_1;
	wire w_dff_A_KfWFhUva8_1;
	wire w_dff_A_sEhCQmEg5_1;
	wire w_dff_A_gcnzPzKn1_0;
	wire w_dff_A_gxjgvuVr0_1;
	wire w_dff_A_P1G8j8sL8_1;
	wire w_dff_A_OmPDAgAM1_1;
	wire w_dff_A_woM42a805_1;
	wire w_dff_A_Mz2LidRZ3_1;
	wire w_dff_A_QtMsrQbs7_1;
	wire w_dff_A_qGmwrrV43_1;
	wire w_dff_A_u2yqOSGB8_1;
	wire w_dff_A_FuSfG6mH8_1;
	wire w_dff_A_uEB1B4xG0_1;
	wire w_dff_A_qi908Ma83_1;
	wire w_dff_A_A9YZY4lC3_1;
	wire w_dff_A_vKpHolfe5_1;
	wire w_dff_A_ilokYAdb2_1;
	wire w_dff_A_xxYf9NAS1_1;
	wire w_dff_B_X5UPQFDB0_0;
	wire w_dff_A_NbdGURKy2_0;
	wire w_dff_A_Sv7nSz9l8_0;
	wire w_dff_A_FFXW9yYQ2_0;
	wire w_dff_A_tFkBshhu5_0;
	wire w_dff_A_SPOO0Qee5_0;
	wire w_dff_A_dLaasbX10_0;
	wire w_dff_A_ACfXfwOd5_0;
	wire w_dff_A_OKGU5iSW0_0;
	wire w_dff_A_HWnCfUvs6_0;
	wire w_dff_A_qa8Kysc94_0;
	wire w_dff_A_WSlPrr977_0;
	wire w_dff_A_AMiEeM2x1_0;
	wire w_dff_A_4KU2qdNu9_0;
	wire w_dff_A_cP1V2UuK0_0;
	wire w_dff_A_EgStRu3Z1_0;
	wire w_dff_A_fZaJ32m37_0;
	wire w_dff_A_DoHWcUNe7_0;
	wire w_dff_A_RF0FdYnX6_0;
	wire w_dff_B_0gubTSiJ7_1;
	wire w_dff_A_X3wpJNbL7_2;
	wire w_dff_A_xa0iUHlC0_2;
	wire w_dff_A_F4pBuDFz7_2;
	wire w_dff_A_3WTyAe7S4_2;
	wire w_dff_A_6C1fHsB43_2;
	wire w_dff_A_ndzhgdq44_2;
	wire w_dff_A_8oZU5jxL3_2;
	wire w_dff_A_YXHTOKGL7_2;
	wire w_dff_A_nxsvG44V5_2;
	wire w_dff_A_GkxlOikL3_2;
	wire w_dff_A_RiUiXrFZ1_2;
	wire w_dff_A_n5DF96ap2_2;
	wire w_dff_A_egbsKCSp0_2;
	wire w_dff_A_bGYEB6pl8_2;
	wire w_dff_A_0Z6mcsHj6_2;
	wire w_dff_A_tnuH08Or1_2;
	wire w_dff_A_rPeFpmjZ9_2;
	wire w_dff_A_WpnNlCOD7_0;
	wire w_dff_A_lIoSxRE81_0;
	wire w_dff_A_V1kp8t771_0;
	wire w_dff_A_7QRC78JY0_0;
	wire w_dff_A_Lw0NA0X93_0;
	wire w_dff_A_UZoUoleR8_0;
	wire w_dff_A_E761DXP95_0;
	wire w_dff_A_QaSYnA678_0;
	wire w_dff_A_eUgnv7qh7_0;
	wire w_dff_A_m9MJl1UE7_0;
	wire w_dff_A_5U7xi0fk0_0;
	wire w_dff_A_PzPvBfxc1_0;
	wire w_dff_A_VU7ydF1Q8_0;
	wire w_dff_A_eUTDHlIA4_0;
	wire w_dff_A_txV26H1W3_0;
	wire w_dff_A_zSSjrwjo9_0;
	wire w_dff_A_6BYmRLtj1_0;
	wire w_dff_A_lCny2K5N7_0;
	wire w_dff_B_1BBgLLMX6_1;
	wire w_dff_B_ZDKRkgen7_0;
	wire w_dff_B_DR692JWO3_2;
	wire w_dff_B_o50higMX4_2;
	wire w_dff_A_GhDTW6uW7_0;
	wire w_dff_A_yfxtB0Mj6_0;
	wire w_dff_A_5gr2MZxc3_0;
	wire w_dff_A_QOT75w8e3_0;
	wire w_dff_B_hfhO92eX9_1;
	wire w_dff_B_Tf4sktAQ5_0;
	wire w_dff_B_RoOexd8W5_2;
	wire w_dff_B_s3BtrIMB0_2;
	wire w_dff_A_9ccwibTO2_1;
	wire w_dff_B_xsOrJPyQ6_2;
	wire w_dff_A_OJnxlWYq1_2;
	wire w_dff_A_qSmO3sxM0_2;
	wire w_dff_A_9LQtxqQs0_2;
	wire w_dff_A_cyokqCZy9_2;
	wire w_dff_A_VgXoLfYa4_2;
	wire w_dff_B_S7QK8PnQ1_1;
	wire w_dff_B_GlAauAlX5_0;
	wire w_dff_A_4t9OGUoO9_1;
	wire w_dff_A_ze2TbJmO2_1;
	wire w_dff_A_McacbpMI7_2;
	wire w_dff_A_DSMLlou83_2;
	wire w_dff_A_lhwAhZoi6_1;
	wire w_dff_A_QUdhUQBY9_1;
	wire w_dff_A_AzityleY0_1;
	wire w_dff_A_ttAswpf56_1;
	wire w_dff_A_TLQRb0oS4_1;
	wire w_dff_A_fojp8nj44_1;
	wire w_dff_A_TiY8jbIF4_1;
	wire w_dff_A_Uy6kw2GG4_1;
	wire w_dff_A_QAA4dzyl1_1;
	wire w_dff_A_icwwhiNp2_1;
	wire w_dff_A_BzJeaHSw9_1;
	wire w_dff_A_O2xbLzO42_1;
	wire w_dff_A_qmdxOz5k3_1;
	wire w_dff_B_a6OhZh6Y1_1;
	wire w_dff_B_f82gaWqz6_1;
	wire w_dff_B_tH0iE8Zk9_1;
	wire w_dff_B_1xEumEkB4_1;
	wire w_dff_B_qjwCuMP90_1;
	wire w_dff_B_0H8kGMJe9_1;
	wire w_dff_B_0osHwrEi3_1;
	wire w_dff_B_zL3CkYRw0_1;
	wire w_dff_B_w5dep8MM1_1;
	wire w_dff_B_14DQgkg33_1;
	wire w_dff_B_iS5JGtt31_1;
	wire w_dff_B_1LTYs2VH4_1;
	wire w_dff_B_CXbr2tSP6_1;
	wire w_dff_B_6gyHgv593_1;
	wire w_dff_B_o9pz9yqM5_1;
	wire w_dff_A_7qvt01Gw7_1;
	wire w_dff_A_EeAwhK9t6_1;
	wire w_dff_A_jVlUQMio7_1;
	wire w_dff_A_HybwZxUB0_1;
	wire w_dff_A_45QPxJd27_1;
	wire w_dff_A_9zizjlgD3_1;
	wire w_dff_A_a2DMK6Mh4_1;
	wire w_dff_B_yiMi5WIJ2_1;
	wire w_dff_B_RPzbXaBE0_1;
	wire w_dff_B_oicmsVBS8_1;
	wire w_dff_B_EEYomzKA0_1;
	wire w_dff_B_Z9Yjz69g1_1;
	wire w_dff_B_nPL5O5D18_1;
	wire w_dff_B_aKKKoBAO2_1;
	wire w_dff_B_Me8b3bQA0_1;
	wire w_dff_B_zoefxJOB6_1;
	wire w_dff_B_oRD1y27v5_1;
	wire w_dff_B_Hit352gK4_1;
	wire w_dff_B_LBb1e79w3_1;
	wire w_dff_B_Md0cH27z3_1;
	wire w_dff_A_j7Vpwvjf1_0;
	wire w_dff_A_nMqu4bjN2_0;
	wire w_dff_A_cU02PYpS4_0;
	wire w_dff_A_RgqDsN3a3_0;
	wire w_dff_A_6Lo7wcKL3_0;
	wire w_dff_A_2ImJFL3k4_0;
	wire w_dff_A_BrNc2Zwt0_0;
	wire w_dff_A_ZB5F9ZHS6_0;
	wire w_dff_A_wY4cOqzB6_0;
	wire w_dff_A_ujQXfP9L6_0;
	wire w_dff_A_TRgHmW7P3_0;
	wire w_dff_A_h6jXJq6t3_1;
	wire w_dff_A_MhbFbLx72_1;
	wire w_dff_A_KdPodqNV8_1;
	wire w_dff_A_a4AEExw83_1;
	wire w_dff_A_fuN38Th80_1;
	wire w_dff_A_XYunfvvK4_1;
	wire w_dff_A_CIq3GO9s4_1;
	wire w_dff_A_4NkmOesI3_1;
	wire w_dff_A_gxjmdQNJ1_1;
	wire w_dff_A_BfOUIvdr8_1;
	wire w_dff_A_nbD5zfLn8_1;
	wire w_dff_A_Nx1p4Kpj3_1;
	wire w_dff_A_DfWVp4ef4_1;
	wire w_dff_A_MGkzqXCE2_1;
	wire w_dff_A_hFM6fXmV7_1;
	wire w_dff_A_kkEaQzo72_2;
	wire w_dff_A_md8RtMPF9_2;
	wire w_dff_A_9H7CSzP19_0;
	wire w_dff_A_oQuHNRS80_1;
	wire w_dff_A_R95kl5eb2_2;
	wire w_dff_A_gKKIKIjz5_2;
	wire w_dff_A_dGv0HnBV7_2;
	wire w_dff_A_xtbKG4df1_0;
	wire w_dff_A_itcAS2LG7_0;
	wire w_dff_A_VWIuIhjw6_0;
	wire w_dff_A_u9hrOZe56_0;
	wire w_dff_A_HAQrLaVw1_0;
	wire w_dff_A_E4QIsxER2_1;
	wire w_dff_A_QisLD6h50_1;
	wire w_dff_A_GngKVSlr5_1;
	wire w_dff_A_yLqtJmZL3_1;
	wire w_dff_A_3WoZ6Qs11_1;
	wire w_dff_A_aMyWZKbS1_1;
	wire w_dff_A_oKs18H4K4_1;
	wire w_dff_B_iS4GFBys8_2;
	wire w_dff_B_OC3cbWcf6_2;
	wire w_dff_B_hsmlqB6f6_2;
	wire w_dff_B_7CLyjbwD3_2;
	wire w_dff_B_6GTJuSD64_2;
	wire w_dff_B_qZe0Y4ZI8_2;
	wire w_dff_B_yU4cyUmK7_2;
	wire w_dff_B_jm3SBMPv0_2;
	wire w_dff_A_V9Yu8TzO9_0;
	wire w_dff_A_QQEgXUCX7_0;
	wire w_dff_A_Ydu3eo0F2_0;
	wire w_dff_A_nVS25w047_0;
	wire w_dff_A_XWCBOf1L4_0;
	wire w_dff_A_13P1wu2X7_0;
	wire w_dff_A_ljIFcQ6O6_0;
	wire w_dff_A_fcEi5dX74_2;
	wire w_dff_A_pFRmMylo5_2;
	wire w_dff_A_Y0RvLGZH2_2;
	wire w_dff_A_addw5Elf2_2;
	wire w_dff_A_aOM5wPos3_2;
	wire w_dff_A_a0xwW19R2_2;
	wire w_dff_A_m7BPBVeD9_2;
	wire w_dff_A_pglbKG1h6_2;
	wire w_dff_A_PQfki17f3_2;
	wire w_dff_A_BbqT1xbR5_2;
	wire w_dff_A_2EevMicO9_2;
	wire w_dff_A_j45oVpwh7_0;
	wire w_dff_A_jiux9eNi8_0;
	wire w_dff_A_bplawuSj0_0;
	wire w_dff_A_y4JmTDcA8_0;
	wire w_dff_A_WfVSZ6Rn1_0;
	wire w_dff_A_amHkDlX56_0;
	wire w_dff_A_IYP4Qtpr2_0;
	wire w_dff_A_f47I2eI74_1;
	wire w_dff_A_9iXGh8Hf9_1;
	wire w_dff_A_rXPU0POp2_1;
	wire w_dff_A_YSOuSMyB4_1;
	wire w_dff_A_HwNhSJvh4_1;
	wire w_dff_A_eYogqwxd6_1;
	wire w_dff_A_VANahx7h4_1;
	wire w_dff_A_q7M6kJU42_1;
	wire w_dff_A_q4eSgDJJ1_1;
	wire w_dff_A_vULS35Ya7_1;
	wire w_dff_A_vjUkS9AR4_1;
	wire w_dff_A_nSimRdzg0_1;
	wire w_dff_A_m1xlhcAx1_0;
	wire w_dff_A_eWSBL3Rl6_1;
	wire w_dff_A_tDpN4mup8_1;
	wire w_dff_A_IvD4zRpv4_1;
	wire w_dff_A_STxpAMYJ6_1;
	wire w_dff_A_Zz1qrTBt0_1;
	wire w_dff_A_UPRVCcTd1_1;
	wire w_dff_A_GWv2Ifkk4_1;
	wire w_dff_A_3n4UuHX64_1;
	wire w_dff_A_eXxIkS7S1_1;
	wire w_dff_A_rVEXEA3D4_1;
	wire w_dff_A_f10blSsZ4_1;
	wire w_dff_A_mqsdTUsB8_1;
	wire w_dff_A_yJoL8IxM9_1;
	wire w_dff_A_pnN4e0tt2_1;
	wire w_dff_A_icuiq9cj9_1;
	wire w_dff_A_Jy21ZVUD4_1;
	wire w_dff_B_lncsuzpc2_1;
	wire w_dff_B_NdacBAVQ8_0;
	wire w_dff_B_MCOGhzGZ9_2;
	wire w_dff_B_JLLYtHSi6_2;
	wire w_dff_A_jsUAqiQy4_0;
	wire w_dff_A_Nwk7wgF06_0;
	wire w_dff_A_5POAQ0Lp3_0;
	wire w_dff_A_KsBxcwTl2_0;
	wire w_dff_B_eBTD6XLU8_1;
	wire w_dff_B_VTqLAKE61_0;
	wire w_dff_A_fD6XjZkR4_1;
	wire w_dff_A_hOgeOUPF7_1;
	wire w_dff_A_wLnxcjBH0_2;
	wire w_dff_A_iC5C8OjB4_2;
	wire w_dff_A_DeYJNhYT6_1;
	wire w_dff_A_YXAAON592_1;
	wire w_dff_A_yT4V3izG7_1;
	wire w_dff_A_RQNKq2ED1_1;
	wire w_dff_A_H1TkR1ev1_0;
	wire w_dff_A_w25X416A8_0;
	wire w_dff_A_lUCU7CAt0_0;
	wire w_dff_A_VOURb8ns2_0;
	wire w_dff_A_Q1cYFrFu1_0;
	wire w_dff_A_xwFz6suw3_0;
	wire w_dff_A_e9mg32bY4_0;
	wire w_dff_A_kGhswp7n5_0;
	wire w_dff_A_XH39Dzng4_0;
	wire w_dff_A_UhNbnvkD5_0;
	wire w_dff_A_F7SLceJQ5_0;
	wire w_dff_A_fviSfmSJ5_0;
	wire w_dff_A_LqCO2wEt1_0;
	wire w_dff_A_L8Jt8ksO4_0;
	wire w_dff_A_4y45Qwkg8_0;
	wire w_dff_A_yAcqsvcv1_0;
	wire w_dff_A_hnsfD6Wa9_0;
	wire w_dff_A_Ec1vrAUN4_0;
	wire w_dff_A_Q4gWlfxQ5_0;
	wire w_dff_A_tc4wjIme4_0;
	wire w_dff_A_WKkDVb398_0;
	wire w_dff_A_zWBuL2iM5_0;
	wire w_dff_A_7nbNurT41_0;
	wire w_dff_A_1UPCQan38_0;
	wire w_dff_A_Db3vSDXQ2_0;
	wire w_dff_A_fgRorDQ94_0;
	wire w_dff_A_834GmKxn6_0;
	wire w_dff_A_mr411PyE1_2;
	wire w_dff_A_diwNUycN8_2;
	wire w_dff_A_z8Of0bIP4_2;
	wire w_dff_A_cL81nsjY6_2;
	wire w_dff_A_i3EjHGms9_2;
	wire w_dff_A_65K3OV268_2;
	wire w_dff_A_eq2zt1Y13_2;
	wire w_dff_A_OtOJedEa0_2;
	wire w_dff_A_TBsNULbG4_2;
	wire w_dff_A_7AA5fqZw8_2;
	wire w_dff_A_AzHJQS0M2_2;
	wire w_dff_A_eg8aB7iI1_2;
	wire w_dff_A_rGfyodch6_2;
	wire w_dff_A_vgM6wKl89_2;
	wire w_dff_B_zfeiiKV59_1;
	wire w_dff_B_B9vMYkRe1_0;
	wire w_dff_B_qmQ8RXc35_2;
	wire w_dff_B_mbNgPm2M9_2;
	wire w_dff_A_fBS8ixlD8_2;
	wire w_dff_A_UaorlTs97_2;
	wire w_dff_A_WWwU03BM3_2;
	wire w_dff_A_E5eUml0l6_2;
	wire w_dff_A_YjrnoYQ10_1;
	wire w_dff_A_6V5Tyu9B5_1;
	wire w_dff_A_IrR3M08e7_1;
	wire w_dff_A_CjzTuaok6_1;
	wire w_dff_A_Ai8doFeD4_1;
	wire w_dff_A_B4W2SeIN8_1;
	wire w_dff_A_h7He2goE9_1;
	wire w_dff_A_C3wFZKjy1_1;
	wire w_dff_A_aoA6KkSh8_1;
	wire w_dff_A_lwRixicT2_1;
	wire w_dff_A_JcXsaGgX0_1;
	wire w_dff_A_kkzKgLQU8_1;
	wire w_dff_A_ytGAotxk2_1;
	wire w_dff_A_UbRdQzBQ3_1;
	wire w_dff_A_FI0vtvFW6_1;
	wire w_dff_A_XafuP8tA7_1;
	wire w_dff_B_Ay4BhMt72_1;
	wire w_dff_B_d32fgfP58_0;
	wire w_dff_B_XMHt8AVL9_2;
	wire w_dff_B_o3YYZP3c6_2;
	wire w_dff_A_psUMw5Bv8_0;
	wire w_dff_A_ew2MzLwk9_0;
	wire w_dff_A_8ek1yGCB3_0;
	wire w_dff_A_pTOs2fBc6_0;
	wire w_dff_A_6MdOfsxL0_0;
	wire w_dff_A_AIIYD2so7_0;
	wire w_dff_A_REoYckIc9_0;
	wire w_dff_A_KUOvir0x7_0;
	wire w_dff_A_d40E8XcC7_0;
	wire w_dff_A_ynijqlNQ3_0;
	wire w_dff_A_Kpdj06vu8_0;
	wire w_dff_A_7xQjhrrT7_0;
	wire w_dff_A_INjiewfE2_0;
	wire w_dff_A_ejd5kZHd0_0;
	wire w_dff_A_6p5yPW499_0;
	wire w_dff_A_4AXJbFjP3_0;
	wire w_dff_A_gvkPwK1R6_0;
	wire w_dff_A_hguD7QRp5_0;
	wire w_dff_A_tYjulFFW0_1;
	wire w_dff_A_txsL6BBs8_1;
	wire w_dff_A_zkIvd3R72_1;
	wire w_dff_A_iDFAnv7Y7_2;
	wire w_dff_A_Pvhb6ZV98_2;
	wire w_dff_B_S8Z1ZWjF1_3;
	wire w_dff_B_w0b9mGea6_3;
	wire w_dff_B_hpaCQnrD8_1;
	wire w_dff_B_zO4tm7vU4_0;
	wire w_dff_B_TXLOIQC71_2;
	wire w_dff_B_6kXN9UvO1_2;
	wire w_dff_A_a3ffRSgg9_0;
	wire w_dff_A_nM7jgZub7_0;
	wire w_dff_A_I120n9PQ1_0;
	wire w_dff_A_9AKXfkfi4_0;
	wire w_dff_B_aV689boM3_1;
	wire w_dff_B_EMrRo1jj1_1;
	wire w_dff_B_LFNDJRb97_1;
	wire w_dff_B_PaXEQWEA3_1;
	wire w_dff_B_yKZFxwnm6_1;
	wire w_dff_B_8AhLXQQP6_1;
	wire w_dff_B_MdLgWlRM9_1;
	wire w_dff_B_xiawR7N49_1;
	wire w_dff_B_T6NLPMsr0_1;
	wire w_dff_B_VXnoGf3b7_1;
	wire w_dff_B_XvmBW3hC8_1;
	wire w_dff_B_skb62kuA6_1;
	wire w_dff_B_P7LsQFV40_1;
	wire w_dff_B_DN46X9li4_1;
	wire w_dff_B_W5HpanmD0_1;
	wire w_dff_B_FNWAFQOO8_1;
	wire w_dff_B_xZN7lzeh2_1;
	wire w_dff_B_arJKPxfw8_1;
	wire w_dff_A_2ydoM0Lz3_0;
	wire w_dff_A_0Q5F53ju8_0;
	wire w_dff_A_eGfvfQ5k5_0;
	wire w_dff_A_sYy0gg4E5_1;
	wire w_dff_A_HTS5qAX63_1;
	wire w_dff_A_rWmUNWKg4_1;
	wire w_dff_A_1qpZwEpq4_1;
	wire w_dff_A_fj54Z1BF9_1;
	wire w_dff_A_HL8nOjL58_1;
	wire w_dff_A_dzxADrtF4_1;
	wire w_dff_A_U4zVM82Y9_0;
	wire w_dff_A_n9LvWGKt4_0;
	wire w_dff_A_M2ofONVP6_0;
	wire w_dff_A_p6MopZZu3_0;
	wire w_dff_A_ahdM1dSZ2_0;
	wire w_dff_A_Z2ePpNmk0_0;
	wire w_dff_A_TutWKrlk6_0;
	wire w_dff_A_npGINIGV7_0;
	wire w_dff_A_iIlM0pb63_0;
	wire w_dff_A_SApXtcds4_0;
	wire w_dff_A_I8ZCmTMw6_0;
	wire w_dff_A_zL1CMt5T3_1;
	wire w_dff_A_zdNmMN4z5_1;
	wire w_dff_A_Kutyw1wQ0_1;
	wire w_dff_A_cVl90BdP7_1;
	wire w_dff_A_tWk0h5Mk6_1;
	wire w_dff_A_ONqJEs5t9_1;
	wire w_dff_A_2RymdssX3_1;
	wire w_dff_A_gnpfGqTm5_1;
	wire w_dff_A_JJmyLzV54_1;
	wire w_dff_A_7g1m9XmN6_1;
	wire w_dff_A_MTC5u9nW3_1;
	wire w_dff_A_Kvr04JiN4_1;
	wire w_dff_A_UOjkKZjf8_1;
	wire w_dff_A_vf1lO32r1_2;
	wire w_dff_A_I6NJZyvv3_2;
	wire w_dff_A_tpefdaWu0_2;
	wire w_dff_A_xg2SzjY73_2;
	wire w_dff_A_HtcKTuk79_2;
	wire w_dff_A_z767cB1A0_2;
	wire w_dff_A_LwSPtd0c8_2;
	wire w_dff_A_68v2XJIJ9_2;
	wire w_dff_A_uNmMGJuS4_2;
	wire w_dff_A_Sm5KmY0V8_2;
	wire w_dff_A_zAvLW0qS0_2;
	wire w_dff_A_3mdVLWpU8_2;
	wire w_dff_A_Jif3DlyP9_2;
	wire w_dff_B_sazdHijE6_0;
	wire w_dff_B_SrJEm8ST2_0;
	wire w_dff_B_Q71OLlIm8_0;
	wire w_dff_B_yLAvauhF0_0;
	wire w_dff_B_roJCGVcF8_0;
	wire w_dff_B_8LVKQobM8_0;
	wire w_dff_B_bzKPX9cf4_0;
	wire w_dff_B_d1aAI8ly4_0;
	wire w_dff_B_Az2yaSxJ4_0;
	wire w_dff_B_ozeg8SWK8_0;
	wire w_dff_B_dE3sVdpW8_0;
	wire w_dff_B_N05BqhbP3_1;
	wire w_dff_B_NIqczoov3_1;
	wire w_dff_B_qI4S16l17_1;
	wire w_dff_A_3xDhesA69_0;
	wire w_dff_A_o1ibeUd56_0;
	wire w_dff_B_pLSfkFdq2_0;
	wire w_dff_B_r2mzG9rG0_0;
	wire w_dff_B_6dtNDip40_1;
	wire w_dff_B_9hQjcZU16_1;
	wire w_dff_B_pGs50NTd7_1;
	wire w_dff_B_9fCmHICZ8_0;
	wire w_dff_B_2NxGL0PU0_0;
	wire w_dff_B_oOQZMAY02_0;
	wire w_dff_B_uBDpo2xi1_0;
	wire w_dff_B_fEle8DqW2_0;
	wire w_dff_A_T9LZAj526_0;
	wire w_dff_A_OtQD0IBF3_0;
	wire w_dff_A_6NPsbDMG0_0;
	wire w_dff_B_5Ifwxcif7_0;
	wire w_dff_A_UWlumCSz6_0;
	wire w_dff_A_r61HzQDy6_0;
	wire w_dff_A_tf5p52Ec4_0;
	wire w_dff_A_dPrAgsv13_0;
	wire w_dff_A_dOaRQNjy6_0;
	wire w_dff_B_NWmQF8Ab9_0;
	wire w_dff_B_YtMXNCep7_1;
	wire w_dff_A_cU7m0Lw71_1;
	wire w_dff_B_w8rOjI4n1_2;
	wire w_dff_B_3XopZPmy5_0;
	wire w_dff_B_vR2uCBVR6_0;
	wire w_dff_B_3KXtXQqc2_0;
	wire w_dff_B_ZmV7R1xK6_0;
	wire w_dff_B_0XqqsElB1_0;
	wire w_dff_A_LuCcrrTp7_1;
	wire w_dff_A_YmjYPiIJ5_1;
	wire w_dff_A_4RzCVLNv9_1;
	wire w_dff_A_RvvrxBSi0_1;
	wire w_dff_A_C86U8i2H1_1;
	wire w_dff_A_b9c2Mbgn9_1;
	wire w_dff_A_r3qnJ5C00_1;
	wire w_dff_A_QtZCvjht7_1;
	wire w_dff_A_BZUMQKgO2_1;
	wire w_dff_A_Da3PXiuw3_1;
	wire w_dff_A_GpkEY0jh0_1;
	wire w_dff_A_J8hwEzkF8_1;
	wire w_dff_A_xIQ7gbAj8_1;
	wire w_dff_A_HG3c8mgp8_1;
	wire w_dff_A_9j1YVS9y4_1;
	wire w_dff_B_9MsAzG8q7_1;
	wire w_dff_B_Q8FR69JP3_1;
	wire w_dff_A_SXs6JVZ94_0;
	wire w_dff_A_Av51p9Z88_0;
	wire w_dff_A_3GBMsHpT0_0;
	wire w_dff_A_h8BPYLPv4_0;
	wire w_dff_A_4HO5pGpq3_0;
	wire w_dff_B_R97nAaRo7_1;
	wire w_dff_B_1aY1013Z9_1;
	wire w_dff_A_Rq9lncRI9_0;
	wire w_dff_A_tPE7GcZP7_0;
	wire w_dff_A_2CcqA3Wp5_1;
	wire w_dff_A_A4Tkes5G2_1;
	wire w_dff_A_5mzia1uA7_1;
	wire w_dff_A_TNobmL449_1;
	wire w_dff_A_AZoqO2o88_1;
	wire w_dff_A_tYXA1acM7_1;
	wire w_dff_A_794GiRhN5_1;
	wire w_dff_A_gnJKtLYn9_1;
	wire w_dff_A_0KXMix2R7_1;
	wire w_dff_A_a6MHcINx3_0;
	wire w_dff_A_P0ECXsiM0_0;
	wire w_dff_A_K58WcmBV6_0;
	wire w_dff_A_f7lECtP44_0;
	wire w_dff_A_9nNDEB4q5_0;
	wire w_dff_A_tvzVDIrl0_0;
	wire w_dff_A_4odcy0QT3_0;
	wire w_dff_A_emGEHPlv5_0;
	wire w_dff_A_FLmQyZFF2_0;
	wire w_dff_A_eybIkGQx0_0;
	wire w_dff_A_dDpbM4O12_1;
	wire w_dff_A_L6t83EmZ4_1;
	wire w_dff_A_fzUHu6em2_1;
	wire w_dff_A_6BKBDSwR7_1;
	wire w_dff_A_S8jMWJYh0_1;
	wire w_dff_A_baKVXvgD7_1;
	wire w_dff_A_LVitKlWq9_1;
	wire w_dff_A_HZOXCUEY6_1;
	wire w_dff_A_wlaO9dSU5_1;
	wire w_dff_A_bykxBIGm9_1;
	wire w_dff_A_7SqSx9tl8_1;
	wire w_dff_A_kmmA1FoC8_1;
	wire w_dff_A_R7HIKgfX4_2;
	wire w_dff_B_vH4nvQFC5_1;
	wire w_dff_B_AjURoX3e3_1;
	wire w_dff_B_H3ACOtNF0_1;
	wire w_dff_B_KOksx7kp3_1;
	wire w_dff_A_Bwoqm0jQ7_0;
	wire w_dff_A_9oJWk3Pj8_0;
	wire w_dff_A_nBMtiG5B5_0;
	wire w_dff_B_eLWVEYyq7_2;
	wire w_dff_A_UqyDJu4D5_1;
	wire w_dff_A_Icd7JuWI5_1;
	wire w_dff_A_RwBj1TKk8_1;
	wire w_dff_A_kXj7iwpq7_1;
	wire w_dff_A_yUGoHWWg2_2;
	wire w_dff_B_pTaV3zpz2_1;
	wire w_dff_A_kF5LMZdN8_1;
	wire w_dff_A_A1OPI00p8_1;
	wire w_dff_A_v4wmxwJL6_2;
	wire w_dff_A_2GrllwjR3_2;
	wire w_dff_A_PZOFBsFT3_0;
	wire w_dff_A_kjJgJEyu9_0;
	wire w_dff_A_UjSvI0Ny8_0;
	wire w_dff_B_5lt25F7C8_2;
	wire w_dff_B_uoIN38tW4_2;
	wire w_dff_B_aEhxahxj8_2;
	wire w_dff_A_Rkv4QTmw4_0;
	wire w_dff_A_dEMNL1jD3_1;
	wire w_dff_A_dlGEQ5aM2_1;
	wire w_dff_B_uHsnKISb7_3;
	wire w_dff_B_HCaRfry94_3;
	wire w_dff_B_CHuIJ1FZ5_3;
	wire w_dff_B_YKTqkjlu3_3;
	wire w_dff_B_GBC6tgsS0_3;
	wire w_dff_B_fNNYFwtv6_3;
	wire w_dff_B_vRBwmbzP8_3;
	wire w_dff_B_Zzbkcf9B6_3;
	wire w_dff_B_jM3c1MzT9_3;
	wire w_dff_B_EsOLP7h00_3;
	wire w_dff_B_18wAMXjE5_3;
	wire w_dff_A_ZB8TSSX78_0;
	wire w_dff_A_e4bLKr3j3_0;
	wire w_dff_A_C5lxxWGP2_0;
	wire w_dff_A_SFO0hwky9_0;
	wire w_dff_A_NT4AtEq80_0;
	wire w_dff_A_fQAJd3EL8_0;
	wire w_dff_A_5yjwNBpz2_0;
	wire w_dff_A_SelS453N1_0;
	wire w_dff_A_qrO3UpGs9_0;
	wire w_dff_A_p2bKUdqv7_0;
	wire w_dff_A_WH1e1dBZ8_0;
	wire w_dff_A_4Iu5KSXc9_0;
	wire w_dff_A_rkpjtdP25_0;
	wire w_dff_A_WgW83LfH5_0;
	wire w_dff_A_XxhC2lv49_2;
	wire w_dff_A_KjHWuwaD6_2;
	wire w_dff_A_wROp01Cy2_2;
	wire w_dff_A_N2XdCU0N8_2;
	wire w_dff_A_vIdPQ6qN6_2;
	wire w_dff_A_kaQKAcE87_1;
	wire w_dff_A_pQu3n5bo0_1;
	wire w_dff_A_rof2vaeC3_1;
	wire w_dff_A_KzlUK4uX4_1;
	wire w_dff_A_AAVX09nF5_1;
	wire w_dff_A_WFnPfGsW1_2;
	wire w_dff_A_9fMpdCo01_2;
	wire w_dff_A_xeuuFKas7_2;
	wire w_dff_A_n39KGL7a6_2;
	wire w_dff_A_1wZzwL965_2;
	wire w_dff_A_GbpiApuL1_2;
	wire w_dff_A_iubDQSNR7_2;
	wire w_dff_A_zIkDMXcZ8_2;
	wire w_dff_A_8se1Bysi3_2;
	wire w_dff_A_dKJHBT0a7_2;
	wire w_dff_A_5gsDfRXy5_2;
	wire w_dff_A_CThn5KxT9_2;
	wire w_dff_A_M4E1PaT90_2;
	wire w_dff_B_B17T1vBb1_0;
	wire w_dff_B_ivaSIiH18_0;
	wire w_dff_B_x4WMh0ub5_1;
	wire w_dff_B_mGxIXwGq5_1;
	wire w_dff_B_JV2A6PtL3_0;
	wire w_dff_A_aUsyYBN80_0;
	wire w_dff_A_iag1hkad3_0;
	wire w_dff_A_8w9F53vG1_1;
	wire w_dff_A_9ZEcId8N2_1;
	wire w_dff_A_pQHBUbia0_2;
	wire w_dff_A_agWuWEKK0_2;
	wire w_dff_A_xCO3wEwh1_1;
	wire w_dff_A_X7auKSNU3_1;
	wire w_dff_A_LkTghKlY6_1;
	wire w_dff_A_VZOYcmTX5_1;
	wire w_dff_A_TrvEIaVe4_1;
	wire w_dff_A_nwt7supn4_1;
	wire w_dff_A_QRLz4kkM9_1;
	wire w_dff_A_ge2KhoMZ4_1;
	wire w_dff_A_6QjljWL94_1;
	wire w_dff_B_bDqZolpk9_2;
	wire w_dff_B_BXVAVGHI5_2;
	wire w_dff_A_NJ16sLVB1_1;
	wire w_dff_A_PWYghY9h1_1;
	wire w_dff_B_XqLl8wJC5_2;
	wire w_dff_B_tJHYdyLG7_2;
	wire w_dff_B_0Y1cWcdy6_1;
	wire w_dff_B_Vz2Xni5H6_0;
	wire w_dff_A_C4MMxLEe2_1;
	wire w_dff_A_pDhCs61i9_1;
	wire w_dff_A_1GwjxuQt0_1;
	wire w_dff_A_ggo8CN6V0_1;
	wire w_dff_A_689w9I3n8_1;
	wire w_dff_A_K5ZrTf5f6_2;
	wire w_dff_A_Hn9NuiWs7_2;
	wire w_dff_A_oezZcvdH4_2;
	wire w_dff_A_rewglPAF1_2;
	wire w_dff_A_kvJ3T86d4_2;
	wire w_dff_A_fJWjDWHI5_2;
	wire w_dff_A_QGWFhGrH0_2;
	wire w_dff_A_kWpWYWT03_2;
	wire w_dff_A_fO1wqDCy3_2;
	wire w_dff_A_rXWtukPu0_2;
	wire w_dff_A_WRFvq4cH9_2;
	wire w_dff_A_zIaVZtZh8_2;
	wire w_dff_B_izFmWNtm7_1;
	wire w_dff_B_pbQHyWMd6_0;
	wire w_dff_A_10QKI3Aw8_0;
	wire w_dff_A_bSEYi0OK8_0;
	wire w_dff_A_zKkWUVVK3_2;
	wire w_dff_A_ouNZOQcj1_2;
	wire w_dff_A_WlxqNpyP9_1;
	wire w_dff_A_JwtNIGmY0_1;
	wire w_dff_A_ysaxURk58_1;
	wire w_dff_A_zBnmxytd5_1;
	wire w_dff_A_pDtEMtL68_1;
	wire w_dff_A_O7Jo6SXl6_1;
	wire w_dff_A_3wySArqs6_1;
	wire w_dff_A_NYHHFhxm7_1;
	wire w_dff_A_KayMGbHT1_1;
	wire w_dff_A_lLFT9WMi5_1;
	wire w_dff_A_wKof2ftZ0_1;
	wire w_dff_A_Zpy5zA207_1;
	wire w_dff_A_ym1Eibhz7_1;
	wire w_dff_B_lULSSn2v6_1;
	wire w_dff_B_0p2ojq8i8_0;
	wire w_dff_A_SsXq4vV18_2;
	wire w_dff_A_fzEbCmmv1_2;
	wire w_dff_A_Myy3nlgI8_2;
	wire w_dff_A_Uq2Gp1T96_2;
	wire w_dff_A_IcAFC0mS5_1;
	wire w_dff_A_EZ39tuNI9_1;
	wire w_dff_A_OCosiyvZ4_1;
	wire w_dff_A_BUTLgfjH3_1;
	wire w_dff_A_AP5bIcxU3_1;
	wire w_dff_A_FtDVlJMR1_1;
	wire w_dff_A_CqddQdSg5_1;
	wire w_dff_A_JN1pSXGJ2_1;
	wire w_dff_A_kCk5ZQvw1_1;
	wire w_dff_A_eNTiblVA7_1;
	wire w_dff_B_dqPP4jvQ7_2;
	wire w_dff_B_XueDhB7k7_1;
	wire w_dff_B_XAFmI2px1_0;
	wire w_dff_A_G4DRRie31_1;
	wire w_dff_A_hKABPv192_1;
	wire w_dff_A_SqMPRcZC1_2;
	wire w_dff_A_OtRZhWkL0_2;
	wire w_dff_A_BuLXbkO42_1;
	wire w_dff_A_7NPCYtjt2_1;
	wire w_dff_A_cHu6eCAS9_1;
	wire w_dff_A_wq8328gB9_1;
	wire w_dff_B_LtWNy6fy1_1;
	wire w_dff_B_rO78xemd1_1;
	wire w_dff_B_QrSECUrD8_1;
	wire w_dff_B_t2W9AHbf2_1;
	wire w_dff_B_xEOXWKi15_1;
	wire w_dff_B_bqNfjuoh2_1;
	wire w_dff_B_iuGSE1wl9_1;
	wire w_dff_B_bxk3BgJ65_1;
	wire w_dff_B_45VyFlQB5_1;
	wire w_dff_B_ZdHS22Za8_1;
	wire w_dff_B_Tjb98FfF9_1;
	wire w_dff_B_8t3jpyCn9_1;
	wire w_dff_B_q4V9eCAW1_1;
	wire w_dff_A_cysCXh4O1_1;
	wire w_dff_A_bU3HxgH34_1;
	wire w_dff_A_FTVzuvmY1_1;
	wire w_dff_A_Ynu68b1n4_1;
	wire w_dff_A_PDijplF23_1;
	wire w_dff_A_OGbbccXe7_1;
	wire w_dff_A_FuBjQKpz4_1;
	wire w_dff_A_reYAtjlZ6_1;
	wire w_dff_A_6P3ypGPy3_1;
	wire w_dff_A_NUufaEzV0_1;
	wire w_dff_A_2vpKgsog9_1;
	wire w_dff_A_ce8Cg8FA8_1;
	wire w_dff_A_qPcqFAnM7_2;
	wire w_dff_A_b96WBDRe8_2;
	wire w_dff_A_JmNaSGB24_2;
	wire w_dff_A_zA6O4Agt9_2;
	wire w_dff_A_XI4CKZxJ1_0;
	wire w_dff_A_kG63O8gK8_0;
	wire w_dff_A_hkHSszR17_0;
	wire w_dff_A_nJFI4ewU7_0;
	wire w_dff_A_tgb0i89Y2_0;
	wire w_dff_A_0e2A0Xbb2_0;
	wire w_dff_A_vjFv8mU73_0;
	wire w_dff_A_wcqp9dnb6_0;
	wire w_dff_A_9aQUFTwP0_0;
	wire w_dff_A_9fFv3bbF7_1;
	wire w_dff_A_ryOVwv122_1;
	wire w_dff_A_uuO3hIu62_1;
	wire w_dff_A_lAilQdBT7_1;
	wire w_dff_A_igMw3oUG4_1;
	wire w_dff_A_LWSNA2DT0_1;
	wire w_dff_A_wGTAaL9u6_1;
	wire w_dff_A_5np9xzlW8_0;
	wire w_dff_B_ddE4oc3f2_2;
	wire w_dff_B_IrzrFxNw3_2;
	wire w_dff_A_I66KZtkK6_1;
	wire w_dff_A_vpPwzcMV9_1;
	wire w_dff_A_Xub83BwO5_1;
	wire w_dff_A_Q4gslOok1_1;
	wire w_dff_A_VjQZaMGs4_1;
	wire w_dff_B_NUMZYu669_3;
	wire w_dff_A_tj16hwk92_0;
	wire w_dff_A_3SL7naHL2_0;
	wire w_dff_A_L4pp5dTu2_0;
	wire w_dff_A_4z0juuWj9_0;
	wire w_dff_A_eorgmWoP0_2;
	wire w_dff_A_EIYJuf6S6_2;
	wire w_dff_A_YPFFoyh43_2;
	wire w_dff_A_V0MKqD0R2_2;
	wire w_dff_A_zSq0MprW8_2;
	wire w_dff_A_w8ug4njh8_2;
	wire w_dff_A_8QWeCkZB8_0;
	wire w_dff_A_qoaZTQKb9_0;
	wire w_dff_A_8u8zz0hI7_0;
	wire w_dff_B_bRLAOsI35_3;
	wire w_dff_A_ox4zSsWX7_0;
	wire w_dff_A_8S7dEa0i4_1;
	wire w_dff_A_Pqsjnv4v5_0;
	wire w_dff_A_xcezbmkX0_1;
	wire w_dff_A_ueHqDwNa9_1;
	wire w_dff_A_J7rztvn01_1;
	wire w_dff_A_gg61SxAS4_1;
	wire w_dff_A_ZKNFV40b0_2;
	wire w_dff_A_fEUrzPyw6_2;
	wire w_dff_B_C6xg2Z3Z4_1;
	wire w_dff_B_imc1wVcA6_0;
	wire w_dff_A_h8yjWpDz5_1;
	wire w_dff_A_xz0LDdqJ7_0;
	wire w_dff_A_oKX0JHAy5_0;
	wire w_dff_A_CKSZqIIO0_2;
	wire w_dff_A_nAx8PBdD7_2;
	wire w_dff_A_EtjwFWbC2_1;
	wire w_dff_A_xJI09LtI7_1;
	wire w_dff_A_DkSJbuj46_1;
	wire w_dff_A_J8W2vvAm2_1;
	wire w_dff_A_9Y44Fhkp4_1;
	wire w_dff_A_EXP6f9nN5_1;
	wire w_dff_A_tikeZxdx1_1;
	wire w_dff_A_WtEFTgVK8_2;
	wire w_dff_A_6fV3kaxC7_2;
	wire w_dff_A_FSv2gqVb9_2;
	wire w_dff_B_eSI8rUsk5_1;
	wire w_dff_B_qWV7iYu50_0;
	wire w_dff_A_9I9RuQo60_1;
	wire w_dff_A_imEWMNjW5_1;
	wire w_dff_A_lZJY7RlZ8_2;
	wire w_dff_A_woTKomL55_2;
	wire w_dff_A_1G0kWD285_1;
	wire w_dff_A_hyOa1aWo8_1;
	wire w_dff_A_PNL2GcxS9_1;
	wire w_dff_A_x0EMkzxd8_1;
	wire w_dff_A_jObMJrur8_0;
	wire w_dff_A_mKzlczDt4_0;
	wire w_dff_A_KtpsS1Dp0_0;
	wire w_dff_A_KEHmf4lu0_0;
	wire w_dff_A_Gs5W5Cso5_0;
	wire w_dff_A_ZBMCsjP81_0;
	wire w_dff_A_DhWvulUT0_0;
	wire w_dff_A_iimobAsk6_0;
	wire w_dff_A_3kVY6l0E9_0;
	wire w_dff_A_XNShdIJK8_1;
	wire w_dff_A_haP4sgFU1_1;
	wire w_dff_A_Qcljl5nJ4_1;
	wire w_dff_A_wND6vBd05_1;
	wire w_dff_B_A084MN4E7_1;
	wire w_dff_B_uNyvENmp2_0;
	wire w_dff_A_sd1wNqVa8_2;
	wire w_dff_A_QttmMOPF5_1;
	wire w_dff_A_Ovq9bdPh2_1;
	wire w_dff_A_zoLh1nev8_2;
	wire w_dff_A_erNsfYQU8_2;
	wire w_dff_A_nAynoQZb3_1;
	wire w_dff_A_8rwikamZ4_1;
	wire w_dff_A_OQjVDZsr1_1;
	wire w_dff_A_RgggCuSl6_1;
	wire w_dff_A_StDwqhMe5_1;
	wire w_dff_A_SeHU1hgo8_0;
	wire w_dff_A_T3vqXCwM2_0;
	wire w_dff_A_KoxgZOEF1_0;
	wire w_dff_A_bWecyCwf2_0;
	wire w_dff_A_AzJeX3xC8_0;
	wire w_dff_A_sL5HqlXH6_0;
	wire w_dff_A_jEGO6G9f3_0;
	wire w_dff_A_ol50RqS85_0;
	wire w_dff_A_V7E4IWB67_0;
	wire w_dff_A_WAdk7IEB6_0;
	wire w_dff_A_VOrFJZH17_0;
	wire w_dff_A_2mO9BGRa1_0;
	wire w_dff_A_7MkaPO6t1_0;
	wire w_dff_A_yGAzjzMr3_0;
	wire w_dff_A_QldLZweh7_0;
	wire w_dff_A_LRwXOCGr6_0;
	wire w_dff_A_cUxzD6Z81_0;
	wire w_dff_A_w1EMWtID4_0;
	wire w_dff_A_ICd6E9qD0_0;
	wire w_dff_A_Iewlz38u3_0;
	wire w_dff_A_UpIfp7D50_0;
	wire w_dff_A_TTQnkFMr2_0;
	wire w_dff_A_u2fcHUyK2_0;
	wire w_dff_A_KLwZPYX23_0;
	wire w_dff_A_YP5NO6vp6_0;
	wire w_dff_A_gV3La4kk8_0;
	wire w_dff_A_eB55MZVj0_0;
	wire w_dff_A_hKEjw8si9_0;
	wire w_dff_A_TGt4jsAn4_0;
	wire w_dff_A_fe7BH65t8_0;
	wire w_dff_A_NxO8nnaY3_0;
	wire w_dff_A_zwJRnC6v8_0;
	wire w_dff_A_5W9wWePd1_0;
	wire w_dff_A_WjqOJxsZ7_0;
	wire w_dff_A_7qk2mgLd2_0;
	wire w_dff_A_KhKWKH7s8_0;
	wire w_dff_A_3r7eKSVv3_0;
	wire w_dff_A_lnaQpt5X0_1;
	wire w_dff_A_akETpjd88_0;
	wire w_dff_A_BRWlUsTg0_0;
	wire w_dff_A_jbhnCSo23_0;
	wire w_dff_A_CvAgXfbh8_0;
	wire w_dff_A_JOO9heH96_0;
	wire w_dff_A_cb9wsTnb1_0;
	wire w_dff_A_H4a7cb6z9_0;
	wire w_dff_A_0h2NUQrw5_0;
	wire w_dff_A_Er9z4s6r0_0;
	wire w_dff_A_nuuhhDUB4_0;
	wire w_dff_A_Y0tSrl9Y2_0;
	wire w_dff_A_c3mtIW6s2_0;
	wire w_dff_A_ZAyTBcY43_0;
	wire w_dff_A_Jb4htPzv0_0;
	wire w_dff_A_Kno6wHgd8_0;
	wire w_dff_A_asZ4ybZH5_0;
	wire w_dff_A_JcMTuyK20_0;
	wire w_dff_A_E9klAfIO8_0;
	wire w_dff_A_aFhFIG2k8_0;
	wire w_dff_A_pC5ZSHLp6_0;
	wire w_dff_A_dcZZo00o8_0;
	wire w_dff_A_57l2aB2k0_0;
	wire w_dff_A_cZa7Y2LU5_0;
	wire w_dff_A_VtBhzFD22_0;
	wire w_dff_A_ZEnx1QJh6_0;
	wire w_dff_A_4lPC5YK68_0;
	wire w_dff_A_vR5xfdH05_0;
	wire w_dff_A_5pce0cdr3_0;
	wire w_dff_A_ULxU10nX0_0;
	wire w_dff_A_vRm0XJat8_0;
	wire w_dff_A_NoNuQYZl5_0;
	wire w_dff_A_kqJI1BYN8_0;
	wire w_dff_A_33yiYwlA9_0;
	wire w_dff_A_FetlggL45_0;
	wire w_dff_A_qErBFBCE0_0;
	wire w_dff_A_h2R4569f1_0;
	wire w_dff_A_Ka7CPswc2_0;
	wire w_dff_A_nByzfYml7_1;
	wire w_dff_A_J2dNTYMk9_0;
	wire w_dff_A_JlQzPGxX6_0;
	wire w_dff_A_hNT8dqZ58_0;
	wire w_dff_A_RilbSa9c8_0;
	wire w_dff_A_92Y45FwU6_0;
	wire w_dff_A_r1OWdJB38_0;
	wire w_dff_A_d3Oa4mE99_0;
	wire w_dff_A_m8qSEMKx5_0;
	wire w_dff_A_Kol595Eo5_0;
	wire w_dff_A_JTDHGrp79_0;
	wire w_dff_A_uwkSKMaW8_0;
	wire w_dff_A_vfBdUksM7_0;
	wire w_dff_A_02ugSumQ8_0;
	wire w_dff_A_7VOvqwFU2_0;
	wire w_dff_A_ZBMacSA12_0;
	wire w_dff_A_MugumP369_0;
	wire w_dff_A_1giOurUF3_0;
	wire w_dff_A_cor92Twd7_0;
	wire w_dff_A_3AHtEvjq0_0;
	wire w_dff_A_oDe15tqa7_0;
	wire w_dff_A_LzM80Iw81_0;
	wire w_dff_A_O3R5Eqsw7_0;
	wire w_dff_A_ax8DhLVl6_0;
	wire w_dff_A_XmvNloMl0_0;
	wire w_dff_A_v7bhiMPO1_0;
	wire w_dff_A_b14A3KCN9_0;
	wire w_dff_A_A8Uh0u299_0;
	wire w_dff_A_3vw78fWU2_0;
	wire w_dff_A_IVFV1qeD7_0;
	wire w_dff_A_cDn6Vza06_0;
	wire w_dff_A_U3Ur1uFB9_0;
	wire w_dff_A_gjmkPsRA6_0;
	wire w_dff_A_bm8orVMl7_0;
	wire w_dff_A_eTtD0IZL0_0;
	wire w_dff_A_v33XOql27_0;
	wire w_dff_A_mSnL3nEr0_0;
	wire w_dff_A_PC9rFL5d2_0;
	wire w_dff_A_X1gH7vPc7_1;
	wire w_dff_A_ydkh7xRL8_0;
	wire w_dff_A_FCvaEbTU9_0;
	wire w_dff_A_yJcuvwvd0_0;
	wire w_dff_A_CLlJzujA7_0;
	wire w_dff_A_25TzLaDL2_0;
	wire w_dff_A_GCGFgT1b1_0;
	wire w_dff_A_svYKQF5g5_0;
	wire w_dff_A_7bwT5q4B2_0;
	wire w_dff_A_cfzUSbMH7_0;
	wire w_dff_A_zverzQER2_0;
	wire w_dff_A_0N9Zz3165_0;
	wire w_dff_A_q3lNx0fH3_0;
	wire w_dff_A_S9xkrVUq0_0;
	wire w_dff_A_KzOr32x21_0;
	wire w_dff_A_cbP674Kv9_0;
	wire w_dff_A_atdhSgYQ0_0;
	wire w_dff_A_XEooD6Y84_0;
	wire w_dff_A_PMEDLE3F2_0;
	wire w_dff_A_unq1obuO9_0;
	wire w_dff_A_9pChAC9s5_0;
	wire w_dff_A_OxLpBcm77_0;
	wire w_dff_A_DNwDOW2w1_0;
	wire w_dff_A_MmIfOmpd2_0;
	wire w_dff_A_UhhXUQQY4_0;
	wire w_dff_A_xN8E6Ghb2_0;
	wire w_dff_A_PXYf0dZq4_0;
	wire w_dff_A_hfN5wi7i8_0;
	wire w_dff_A_oPajINVY9_0;
	wire w_dff_A_pnYtcv6T3_0;
	wire w_dff_A_YkqGDftS9_0;
	wire w_dff_A_RtToPjVr3_0;
	wire w_dff_A_ilREnJUH4_0;
	wire w_dff_A_FeK7bATw0_0;
	wire w_dff_A_lKYIe5Vw6_0;
	wire w_dff_A_wWOuanCo7_0;
	wire w_dff_A_E4l51J4X3_0;
	wire w_dff_A_f9ECAxSt3_0;
	wire w_dff_A_uLsdXGj77_1;
	wire w_dff_A_NX1FLLKx8_0;
	wire w_dff_A_i1fIY9VA9_0;
	wire w_dff_A_vinnMVKQ3_0;
	wire w_dff_A_Z6MLrGcd7_0;
	wire w_dff_A_8HtCx68v9_0;
	wire w_dff_A_gZq3zVus4_0;
	wire w_dff_A_l7tOmevN2_0;
	wire w_dff_A_OgqSDkSL2_0;
	wire w_dff_A_lPJuA1QS4_0;
	wire w_dff_A_nn0FKwip9_0;
	wire w_dff_A_NsBrquGu9_0;
	wire w_dff_A_CSnJrBrw5_0;
	wire w_dff_A_gP7CTIag1_0;
	wire w_dff_A_L5iHt3dr8_0;
	wire w_dff_A_K6JvbFWp4_0;
	wire w_dff_A_9fcGjbCy8_0;
	wire w_dff_A_wS6cb22j4_0;
	wire w_dff_A_GX3cdPUI3_0;
	wire w_dff_A_Lkvpz61y5_0;
	wire w_dff_A_GQehuQGn9_0;
	wire w_dff_A_BMg5TUVv2_0;
	wire w_dff_A_wZ2f8pTL6_0;
	wire w_dff_A_83ZOiplb4_0;
	wire w_dff_A_cE5GgqAB8_0;
	wire w_dff_A_GgNHQkRp9_0;
	wire w_dff_A_vIWR0YOL4_0;
	wire w_dff_A_w0W6kF634_0;
	wire w_dff_A_8os3EzAM6_0;
	wire w_dff_A_7nuPcMTJ8_0;
	wire w_dff_A_fXIeBo3c7_0;
	wire w_dff_A_DTuzhzlB3_0;
	wire w_dff_A_vbAbtqJV7_0;
	wire w_dff_A_FDpsTSAO0_0;
	wire w_dff_A_3PMa9iHI6_0;
	wire w_dff_A_cPOODtLB6_0;
	wire w_dff_A_cH04DPs96_0;
	wire w_dff_A_ybJM6jXC5_0;
	wire w_dff_A_2l1hqVy46_1;
	wire w_dff_A_9d3UVCu13_0;
	wire w_dff_A_KGfjFnLn0_0;
	wire w_dff_A_Z6Fss6RC9_0;
	wire w_dff_A_tf6WkaWM4_0;
	wire w_dff_A_Jau20yRE0_0;
	wire w_dff_A_H4CrkWjr8_0;
	wire w_dff_A_qMt4R6XX4_0;
	wire w_dff_A_tRWnFen94_0;
	wire w_dff_A_pPyLbdqA5_0;
	wire w_dff_A_aFPXLgXY1_0;
	wire w_dff_A_8MX3tftK2_0;
	wire w_dff_A_mSxr0lMG2_0;
	wire w_dff_A_CAYi5kPi8_0;
	wire w_dff_A_tk7VeiD46_0;
	wire w_dff_A_2YjvvqZ29_0;
	wire w_dff_A_oYZRwpwO7_0;
	wire w_dff_A_dic5qb4a4_0;
	wire w_dff_A_OmWpxsGv9_0;
	wire w_dff_A_bZp5g0I93_0;
	wire w_dff_A_kinliT5j2_0;
	wire w_dff_A_5Hc9Ldb98_0;
	wire w_dff_A_Dwc2Xno58_0;
	wire w_dff_A_rmc3rdFx6_0;
	wire w_dff_A_3HQ4aECa5_0;
	wire w_dff_A_6L5t83EB3_0;
	wire w_dff_A_jNTqtUKP1_0;
	wire w_dff_A_e5cC8NpR5_0;
	wire w_dff_A_vFOy2fyY4_0;
	wire w_dff_A_8EL24QTX0_0;
	wire w_dff_A_nqbQipO56_0;
	wire w_dff_A_5cxFsShh1_0;
	wire w_dff_A_nowipb605_0;
	wire w_dff_A_SHE8aMfO7_0;
	wire w_dff_A_5wO5d7hK3_0;
	wire w_dff_A_dfNJmO6F8_0;
	wire w_dff_A_q2Ks7Jvr8_0;
	wire w_dff_A_2rX7MfhW7_0;
	wire w_dff_A_HiWLfWKP7_1;
	wire w_dff_A_0UCvrhVi4_0;
	wire w_dff_A_n8cv8puG5_0;
	wire w_dff_A_RYvqZK1l1_0;
	wire w_dff_A_ENzhW5jK9_0;
	wire w_dff_A_dVMDnWrn3_0;
	wire w_dff_A_8e1c2y0W5_0;
	wire w_dff_A_xRJmrmeE0_0;
	wire w_dff_A_ATMFP5mw9_0;
	wire w_dff_A_fNIQnVzC4_0;
	wire w_dff_A_C12bCA4o3_0;
	wire w_dff_A_8ZbMhV4i6_0;
	wire w_dff_A_y9pz8Om91_0;
	wire w_dff_A_9NF812NG2_0;
	wire w_dff_A_iqBQPIcQ3_0;
	wire w_dff_A_RCkWIBlx8_0;
	wire w_dff_A_bY3ubHh02_0;
	wire w_dff_A_QfxCFLnc7_0;
	wire w_dff_A_xfmKH9L01_0;
	wire w_dff_A_KpNIUVEs0_0;
	wire w_dff_A_MIrF1B9i2_0;
	wire w_dff_A_HzGvQglx0_0;
	wire w_dff_A_4twZSC3O2_0;
	wire w_dff_A_kSagvAEW3_0;
	wire w_dff_A_IolfRFdE2_0;
	wire w_dff_A_GriAU1Pt1_0;
	wire w_dff_A_667x8J2q8_0;
	wire w_dff_A_vLmPdVaY4_0;
	wire w_dff_A_9cXdnejb2_0;
	wire w_dff_A_c9vUUgNJ6_0;
	wire w_dff_A_dSk0q1FY6_0;
	wire w_dff_A_p8LBrKaF4_0;
	wire w_dff_A_LmEwFyAl4_0;
	wire w_dff_A_ipSodC7T5_0;
	wire w_dff_A_frVC1RHd9_0;
	wire w_dff_A_9SQwtwIr4_0;
	wire w_dff_A_pYiQIiIQ6_0;
	wire w_dff_A_S2TA1OUr4_0;
	wire w_dff_A_kvGxlUzO4_1;
	wire w_dff_A_HQiO5ttM3_0;
	wire w_dff_A_wDMwpEe39_0;
	wire w_dff_A_D25LVPdq9_0;
	wire w_dff_A_LdqQ8GS96_0;
	wire w_dff_A_g5SNYsFV2_0;
	wire w_dff_A_7VIbVF2i0_0;
	wire w_dff_A_u5gsozjE8_0;
	wire w_dff_A_bYkPkdv60_0;
	wire w_dff_A_h6GV5PaT1_0;
	wire w_dff_A_5GOGn6aE4_0;
	wire w_dff_A_4RwAOoPy3_0;
	wire w_dff_A_PO8kIc2X7_0;
	wire w_dff_A_G0oO1yNn5_0;
	wire w_dff_A_wcG2Op2J1_0;
	wire w_dff_A_GH70SxUr8_0;
	wire w_dff_A_CcWFvBEL0_0;
	wire w_dff_A_sf5jpRQu8_0;
	wire w_dff_A_0WgsX7tT0_0;
	wire w_dff_A_nnPg39Tz2_0;
	wire w_dff_A_SHnaC6LD5_0;
	wire w_dff_A_WaTtFhQm2_0;
	wire w_dff_A_hD38IotZ8_0;
	wire w_dff_A_rGzf70ts7_0;
	wire w_dff_A_xRDBuaYF9_0;
	wire w_dff_A_xcQvfbi58_0;
	wire w_dff_A_SQGo8CdU4_0;
	wire w_dff_A_LWbBRtU55_0;
	wire w_dff_A_SvM85YHX4_0;
	wire w_dff_A_c7snQ1q51_0;
	wire w_dff_A_14omzql55_0;
	wire w_dff_A_uIKWQI7U1_0;
	wire w_dff_A_GTQTm0DE4_0;
	wire w_dff_A_wYryfeQU2_0;
	wire w_dff_A_R2ME4zqR4_0;
	wire w_dff_A_V5LgGH9N4_0;
	wire w_dff_A_wCgTN6nU2_0;
	wire w_dff_A_pp9IsZJP3_0;
	wire w_dff_A_fKxVyEvG8_1;
	wire w_dff_A_F92hdeRJ0_0;
	wire w_dff_A_lh4qTxSA6_0;
	wire w_dff_A_Lj4aZEHl3_0;
	wire w_dff_A_Ch9i7imW9_0;
	wire w_dff_A_kCkxOE5N3_0;
	wire w_dff_A_dnWzRb6X7_0;
	wire w_dff_A_2SrkhawT5_0;
	wire w_dff_A_J4ggTXvG5_0;
	wire w_dff_A_laU8SMs35_0;
	wire w_dff_A_z1f7J1W22_0;
	wire w_dff_A_FsoH9K6T3_0;
	wire w_dff_A_IoUyw4J14_0;
	wire w_dff_A_QURQmPgQ3_0;
	wire w_dff_A_aLGroFPl3_0;
	wire w_dff_A_LfcpGE3l3_0;
	wire w_dff_A_EqJmcoBQ9_0;
	wire w_dff_A_LUMKoF214_0;
	wire w_dff_A_3yUQLkN69_0;
	wire w_dff_A_bqDVKuKK3_0;
	wire w_dff_A_SAUFHYGW9_0;
	wire w_dff_A_TAfyRZJC0_0;
	wire w_dff_A_LBPJll499_0;
	wire w_dff_A_c2nudf8R7_0;
	wire w_dff_A_KcmDLKqn1_0;
	wire w_dff_A_s16URw4I2_0;
	wire w_dff_A_5JPYUQsM5_0;
	wire w_dff_A_Idu8qWNB6_0;
	wire w_dff_A_1WWExI6x8_0;
	wire w_dff_A_0mnoZRSQ5_0;
	wire w_dff_A_CF2GSWek0_0;
	wire w_dff_A_VQpVfuAR4_0;
	wire w_dff_A_e170Ure11_0;
	wire w_dff_A_3VILppcH7_0;
	wire w_dff_A_l4NAm9en6_0;
	wire w_dff_A_fDmTOJTi1_0;
	wire w_dff_A_hph6m4e00_0;
	wire w_dff_A_PSZgYxFA9_0;
	wire w_dff_A_AcwEvtBl8_1;
	wire w_dff_A_6OWjTLXC6_0;
	wire w_dff_A_rpdzzsy26_0;
	wire w_dff_A_RRnxiAJm6_0;
	wire w_dff_A_Prlg8BjP1_0;
	wire w_dff_A_3bCnMy7x4_0;
	wire w_dff_A_LGjH8Pn65_0;
	wire w_dff_A_VYde3mL26_0;
	wire w_dff_A_aBaFFw074_0;
	wire w_dff_A_YqWJ6E5b9_0;
	wire w_dff_A_ZRs2QVpA7_0;
	wire w_dff_A_9oebRl9I6_0;
	wire w_dff_A_hpjYXzxN6_0;
	wire w_dff_A_OBgwRlmI9_0;
	wire w_dff_A_EnWHsSSQ6_0;
	wire w_dff_A_ZqKAs4xj1_0;
	wire w_dff_A_mcCDbzoh3_0;
	wire w_dff_A_4APlkpIW4_0;
	wire w_dff_A_yGrE6SZE2_0;
	wire w_dff_A_ch7R156V2_0;
	wire w_dff_A_bbSEe4Wi5_0;
	wire w_dff_A_ebmEU7UJ1_0;
	wire w_dff_A_ww67YbTu2_0;
	wire w_dff_A_HNskSIVu3_0;
	wire w_dff_A_VKUvB8OA4_0;
	wire w_dff_A_XE5PC3Zx2_0;
	wire w_dff_A_iRRtSOHo3_0;
	wire w_dff_A_UhSxZrF77_0;
	wire w_dff_A_kTeJyuOT2_0;
	wire w_dff_A_vWv3fmiR5_0;
	wire w_dff_A_w1lbupO53_0;
	wire w_dff_A_nBVCXKhB1_0;
	wire w_dff_A_QbV8s2JN4_0;
	wire w_dff_A_0d02QCDj3_0;
	wire w_dff_A_Cy6LBfrM8_0;
	wire w_dff_A_K8hUt43B8_0;
	wire w_dff_A_JecLXnvU4_0;
	wire w_dff_A_NGD2okon1_0;
	wire w_dff_A_z4lHrBEn5_1;
	wire w_dff_A_wMXkQfNZ7_0;
	wire w_dff_A_PIHhjbMF1_0;
	wire w_dff_A_7XwEtK6h9_0;
	wire w_dff_A_VeQmwW8d0_0;
	wire w_dff_A_1IcuaTuF8_0;
	wire w_dff_A_Q0bxyaBG9_0;
	wire w_dff_A_AC23EK8I0_0;
	wire w_dff_A_1YFYwp1q0_0;
	wire w_dff_A_0uSb1EZf5_0;
	wire w_dff_A_fba7M4lh6_0;
	wire w_dff_A_1V4bVSun7_0;
	wire w_dff_A_GWUFa7EB2_0;
	wire w_dff_A_ydN3znsn0_0;
	wire w_dff_A_Wwalok0z5_0;
	wire w_dff_A_hVfJakKe3_0;
	wire w_dff_A_c6vz4bpA5_0;
	wire w_dff_A_eAhWjZ4y4_0;
	wire w_dff_A_5QBs58y93_0;
	wire w_dff_A_QME7xHGK3_0;
	wire w_dff_A_KUCDi4qU8_0;
	wire w_dff_A_bKhBPAJF1_0;
	wire w_dff_A_M1Vyk1d97_0;
	wire w_dff_A_n9aHY8JG4_0;
	wire w_dff_A_jnuSaW5o8_0;
	wire w_dff_A_WUqwmtjw0_0;
	wire w_dff_A_KQt9Ye494_0;
	wire w_dff_A_mNYPkUIT3_0;
	wire w_dff_A_WPAyqyhM6_0;
	wire w_dff_A_sDJbfh4v8_0;
	wire w_dff_A_eF4yq6ZG2_0;
	wire w_dff_A_rRUU0rwy4_0;
	wire w_dff_A_SRz56pQD2_0;
	wire w_dff_A_U23LyN9s0_0;
	wire w_dff_A_houm0qa04_0;
	wire w_dff_A_EWxXOe9A8_0;
	wire w_dff_A_RA96IEze4_0;
	wire w_dff_A_8oeq2vBk5_0;
	wire w_dff_A_36IIFIIA7_1;
	wire w_dff_A_FkmA8tq38_0;
	wire w_dff_A_9aGlH3DO0_0;
	wire w_dff_A_lMSm5W6U6_0;
	wire w_dff_A_prz6a1sx7_0;
	wire w_dff_A_3cQzEwjl6_0;
	wire w_dff_A_A3wrVfxj6_0;
	wire w_dff_A_ngJ6Fizn9_0;
	wire w_dff_A_ePkytt8P6_0;
	wire w_dff_A_nKeN6kf55_0;
	wire w_dff_A_ukFQpkC67_0;
	wire w_dff_A_9wB1IUS94_0;
	wire w_dff_A_0sQPsP7I3_0;
	wire w_dff_A_IYpIvJiJ2_0;
	wire w_dff_A_OvqoPMTn3_0;
	wire w_dff_A_9QwibUCc8_0;
	wire w_dff_A_R1ICejDp3_0;
	wire w_dff_A_oN2D5d8m5_0;
	wire w_dff_A_YuYOUTou0_0;
	wire w_dff_A_U6BGYJb88_0;
	wire w_dff_A_47TVOq246_0;
	wire w_dff_A_PbVCMIuH5_0;
	wire w_dff_A_ufFMvqlb0_0;
	wire w_dff_A_1M54oIVD0_0;
	wire w_dff_A_BrK1dTY31_0;
	wire w_dff_A_YaIfHXcC6_0;
	wire w_dff_A_gcwgr0Rl8_0;
	wire w_dff_A_ybpOetFU3_0;
	wire w_dff_A_6hEOK7Eq8_0;
	wire w_dff_A_4Yhz2anG0_0;
	wire w_dff_A_zRVHWq2I9_0;
	wire w_dff_A_32HSNbuY5_0;
	wire w_dff_A_xA2Dcb131_0;
	wire w_dff_A_cd7WkMJc1_0;
	wire w_dff_A_P6yfV3Ci3_0;
	wire w_dff_A_DKS9rln26_0;
	wire w_dff_A_gKtsmjWV7_0;
	wire w_dff_A_Kcmhynvt0_0;
	wire w_dff_A_DXzas7OV3_1;
	wire w_dff_A_DitevIQt4_0;
	wire w_dff_A_gXqQdEKN7_0;
	wire w_dff_A_cqb7lCs85_0;
	wire w_dff_A_KZ6waLow6_0;
	wire w_dff_A_KeltLhp16_0;
	wire w_dff_A_Wt7Ebn225_0;
	wire w_dff_A_mlvYLxPi1_0;
	wire w_dff_A_M0xobwCI7_0;
	wire w_dff_A_D25uNUG66_0;
	wire w_dff_A_Cn9l1ycb3_0;
	wire w_dff_A_nYnI3YW30_0;
	wire w_dff_A_XlR2KVD69_0;
	wire w_dff_A_lFNeG9137_0;
	wire w_dff_A_7s3CsHRd6_0;
	wire w_dff_A_szt6NtZ92_0;
	wire w_dff_A_AQOP14g49_0;
	wire w_dff_A_aC1yb7r84_0;
	wire w_dff_A_0AJZRDpq0_0;
	wire w_dff_A_IOWH5kqj7_0;
	wire w_dff_A_CuRnAuZp7_0;
	wire w_dff_A_O6yepDJU3_0;
	wire w_dff_A_lkxaeDzS6_0;
	wire w_dff_A_oPkwPXyi7_0;
	wire w_dff_A_M3HGtLT02_0;
	wire w_dff_A_F3Ojr0sb4_0;
	wire w_dff_A_7Xl7WXQP8_0;
	wire w_dff_A_KsFnX82u9_0;
	wire w_dff_A_5KInHmCx2_0;
	wire w_dff_A_MSMhMbcC5_0;
	wire w_dff_A_lEu24tQd8_0;
	wire w_dff_A_6FfYaLH39_0;
	wire w_dff_A_NT84FmHo9_0;
	wire w_dff_A_2fnemDXS9_0;
	wire w_dff_A_hADZS1ol7_0;
	wire w_dff_A_HFGnETG61_0;
	wire w_dff_A_J3VE4y9D9_0;
	wire w_dff_A_oSWjikhs8_0;
	wire w_dff_A_8wLrcBEf7_1;
	wire w_dff_A_MBtpf6nG4_0;
	wire w_dff_A_zTds5Dbw1_0;
	wire w_dff_A_dLAi06If4_0;
	wire w_dff_A_i9I3egDZ9_0;
	wire w_dff_A_5gnGIPUa4_0;
	wire w_dff_A_7Nvh6Vgj4_0;
	wire w_dff_A_erCiyXWt7_0;
	wire w_dff_A_TYHneHoA3_0;
	wire w_dff_A_FWqguuIS8_0;
	wire w_dff_A_Kz9cUupp4_0;
	wire w_dff_A_LhcF0VFA1_0;
	wire w_dff_A_TWLJK79o0_0;
	wire w_dff_A_AhAOzCav7_0;
	wire w_dff_A_pJDYz61E3_0;
	wire w_dff_A_MgswgbaL1_0;
	wire w_dff_A_mBbmJr9x4_0;
	wire w_dff_A_mwi9elKe0_0;
	wire w_dff_A_8h8XM6yw7_0;
	wire w_dff_A_0Fb1Z5739_0;
	wire w_dff_A_QdUUU36t8_0;
	wire w_dff_A_UZ1PALCw1_0;
	wire w_dff_A_K0ll3kxt0_0;
	wire w_dff_A_tdS0yNrO9_0;
	wire w_dff_A_fUBM5kay7_0;
	wire w_dff_A_1LCeM0fm7_0;
	wire w_dff_A_a6FGzUCU1_0;
	wire w_dff_A_cDyH5COV3_0;
	wire w_dff_A_anFDywGS0_0;
	wire w_dff_A_PqpMyNmQ3_0;
	wire w_dff_A_NJDgWsIe4_0;
	wire w_dff_A_A4NiK8Pt5_0;
	wire w_dff_A_JZ2xUKIN3_0;
	wire w_dff_A_wjYWRq041_0;
	wire w_dff_A_RCutgdgV5_0;
	wire w_dff_A_RuGhyXir1_0;
	wire w_dff_A_MySFxhTV8_0;
	wire w_dff_A_es4GlcNn2_0;
	wire w_dff_A_0XQfGMjy7_1;
	wire w_dff_A_GmWmMbMS4_0;
	wire w_dff_A_xfon8w0f5_0;
	wire w_dff_A_dpXPvg7D6_0;
	wire w_dff_A_CVj0Pjvs7_0;
	wire w_dff_A_qAfRDUAY1_0;
	wire w_dff_A_QfNvzWUm6_0;
	wire w_dff_A_eNVXP6yO2_0;
	wire w_dff_A_OLvJPhHz4_0;
	wire w_dff_A_hcvwTh5I5_0;
	wire w_dff_A_bCeKO90o8_0;
	wire w_dff_A_s8ITB5Uc1_0;
	wire w_dff_A_RjgeXgxr9_0;
	wire w_dff_A_u3rMyb6D9_0;
	wire w_dff_A_Tn0hMPUG9_0;
	wire w_dff_A_SWymwAb43_0;
	wire w_dff_A_bzW8e2QY6_0;
	wire w_dff_A_siXEcYW97_0;
	wire w_dff_A_Ecx6SjWU4_0;
	wire w_dff_A_VwCWuPYR3_0;
	wire w_dff_A_eZclCqGA6_0;
	wire w_dff_A_jL2jo5bH9_0;
	wire w_dff_A_AOQ49JsI8_0;
	wire w_dff_A_iZMLTyxH9_0;
	wire w_dff_A_oKnyiuwN2_0;
	wire w_dff_A_9fE7aXkZ7_0;
	wire w_dff_A_H9OV5D8P3_0;
	wire w_dff_A_tS1YKY697_0;
	wire w_dff_A_CDkfbcBc1_0;
	wire w_dff_A_b8Mrjkzo9_0;
	wire w_dff_A_efP6I1qo1_0;
	wire w_dff_A_Ty0eUYJ12_0;
	wire w_dff_A_xDMHUktA4_0;
	wire w_dff_A_mDxoQrm45_0;
	wire w_dff_A_uCFJA9Sx9_0;
	wire w_dff_A_xQXYupyA1_0;
	wire w_dff_A_vNexCwex3_0;
	wire w_dff_A_gZjphLfx4_0;
	wire w_dff_A_azIhLlon4_1;
	wire w_dff_A_aX7lGb0V6_0;
	wire w_dff_A_BVr18Mkg6_0;
	wire w_dff_A_7IjS7lU89_0;
	wire w_dff_A_f0wHBvQ86_0;
	wire w_dff_A_5gzUUM279_0;
	wire w_dff_A_nTOv59km5_0;
	wire w_dff_A_O0HAABJw1_0;
	wire w_dff_A_aOl1XXUs2_0;
	wire w_dff_A_fhLYO8NA7_0;
	wire w_dff_A_xaMWc1gD3_0;
	wire w_dff_A_SyVGQfqx2_0;
	wire w_dff_A_19Y0Xrxv7_0;
	wire w_dff_A_QXfnmOgn3_0;
	wire w_dff_A_MDxKriLN4_0;
	wire w_dff_A_KwSkPwEL1_0;
	wire w_dff_A_fGAuh8jG0_0;
	wire w_dff_A_Vl3eqJhC7_0;
	wire w_dff_A_9JF6gBlC6_0;
	wire w_dff_A_3wCsGf8m6_0;
	wire w_dff_A_E5FGXIej3_0;
	wire w_dff_A_vuSVhI3f8_0;
	wire w_dff_A_sgL9W5m90_0;
	wire w_dff_A_lgmrrzQR3_0;
	wire w_dff_A_jvqZIyvX9_0;
	wire w_dff_A_92QMTkZo8_0;
	wire w_dff_A_DhptXEy64_0;
	wire w_dff_A_kbsjlWvv7_0;
	wire w_dff_A_xMmYfnOj8_0;
	wire w_dff_A_GRJr3iAi0_0;
	wire w_dff_A_ZWEhvrVo6_0;
	wire w_dff_A_UP7ljwom8_0;
	wire w_dff_A_uvrF2HIT8_0;
	wire w_dff_A_lWV9yiZL0_0;
	wire w_dff_A_I2oZQKlL1_0;
	wire w_dff_A_Z2UxhWsj7_0;
	wire w_dff_A_IjTnKPUP4_0;
	wire w_dff_A_0bdAFRdb1_0;
	wire w_dff_A_OfRm1bFs5_1;
	wire w_dff_A_6KmIy3PK6_0;
	wire w_dff_A_aYfHaKv06_0;
	wire w_dff_A_ZejgaIp97_0;
	wire w_dff_A_yzGc5Yw31_0;
	wire w_dff_A_xqMcAvkU1_0;
	wire w_dff_A_R59MYq8p2_0;
	wire w_dff_A_tiPOHG574_0;
	wire w_dff_A_zkTwiCE67_0;
	wire w_dff_A_2Z5sOrnG3_0;
	wire w_dff_A_0g1jZ2Ei2_0;
	wire w_dff_A_sxPu2aiE8_0;
	wire w_dff_A_qXHISY2e5_0;
	wire w_dff_A_5V6AmOpN0_0;
	wire w_dff_A_IeZXgIph9_0;
	wire w_dff_A_6HeGVw1M1_0;
	wire w_dff_A_bxVfAVKx8_0;
	wire w_dff_A_UF25iH2F4_0;
	wire w_dff_A_7lydPKM67_0;
	wire w_dff_A_12i31rrE7_0;
	wire w_dff_A_aZccxvds0_0;
	wire w_dff_A_Jg6GTRmk2_0;
	wire w_dff_A_uO8ThcsR6_0;
	wire w_dff_A_ryiJoZyX0_0;
	wire w_dff_A_x43oecP31_0;
	wire w_dff_A_LcnKBECF8_0;
	wire w_dff_A_askDIDOz1_0;
	wire w_dff_A_yp5eiI6D2_0;
	wire w_dff_A_0pgN7H7a9_0;
	wire w_dff_A_J0Cl8Llt1_0;
	wire w_dff_A_MsnsuOBh0_0;
	wire w_dff_A_JlaKHGbb1_0;
	wire w_dff_A_7H0JS3R56_0;
	wire w_dff_A_S70F4loh0_0;
	wire w_dff_A_L0KI4wXP4_0;
	wire w_dff_A_NrQNIThS3_0;
	wire w_dff_A_B7IuYAhl5_0;
	wire w_dff_A_M8AkHDF90_0;
	wire w_dff_A_4CAs5RJf1_1;
	wire w_dff_A_QMx2GvSa2_0;
	wire w_dff_A_pSrOzuj04_0;
	wire w_dff_A_w6mjS1H76_0;
	wire w_dff_A_KIIoL9qz8_0;
	wire w_dff_A_geGPXntj4_0;
	wire w_dff_A_8ZxDRM5e6_0;
	wire w_dff_A_Jn6DX5Do3_0;
	wire w_dff_A_Q8F5g7S29_0;
	wire w_dff_A_UxBbbfbk4_0;
	wire w_dff_A_AjFpM39c8_0;
	wire w_dff_A_1m3PDwZa2_0;
	wire w_dff_A_vmH4HACf8_0;
	wire w_dff_A_xwXVKDmV3_0;
	wire w_dff_A_eAEiSS7W8_0;
	wire w_dff_A_YO3aOyis2_0;
	wire w_dff_A_8tlymgnb3_0;
	wire w_dff_A_kZWwcbLK3_0;
	wire w_dff_A_QN2zhAZ00_0;
	wire w_dff_A_Iw8tVeJe3_0;
	wire w_dff_A_A3NyS7Sa5_0;
	wire w_dff_A_4b5jcwNx0_0;
	wire w_dff_A_sch38MpP0_0;
	wire w_dff_A_oTwkmGe08_0;
	wire w_dff_A_zgtpWmSx4_0;
	wire w_dff_A_4x3UBLSF8_0;
	wire w_dff_A_yxhFuPQj5_0;
	wire w_dff_A_OLMT80EA4_0;
	wire w_dff_A_8owFwn9k2_0;
	wire w_dff_A_XP7bJKId0_0;
	wire w_dff_A_5aZy4HNv7_0;
	wire w_dff_A_s5UK2fwQ1_0;
	wire w_dff_A_dIiYmdtN4_0;
	wire w_dff_A_OZgHfJat0_0;
	wire w_dff_A_4XJbp7bv6_0;
	wire w_dff_A_gPxA2HPg8_0;
	wire w_dff_A_pGa0lBVM3_0;
	wire w_dff_A_L3bN9oRH5_0;
	wire w_dff_A_C0h2PJSo2_1;
	wire w_dff_A_3ZlSs3ql0_0;
	wire w_dff_A_u4y4jl7v3_0;
	wire w_dff_A_s6AQ10ey3_0;
	wire w_dff_A_nxrKI0JN5_0;
	wire w_dff_A_4ln3jjCC8_0;
	wire w_dff_A_5Yh2akrM3_0;
	wire w_dff_A_yFRi18p44_0;
	wire w_dff_A_oYyNcA7M6_0;
	wire w_dff_A_oNu8gdjv7_0;
	wire w_dff_A_RTGOMqj45_0;
	wire w_dff_A_9SOpOpus0_0;
	wire w_dff_A_ABGEGEJA6_0;
	wire w_dff_A_SIe8LqtX6_0;
	wire w_dff_A_iVpJPaOb8_0;
	wire w_dff_A_6BmYJTgU8_0;
	wire w_dff_A_GrpZCmGt9_0;
	wire w_dff_A_Ij9f2J918_0;
	wire w_dff_A_RLU4wszg0_0;
	wire w_dff_A_LgTtKnGd6_0;
	wire w_dff_A_6anem5Lo0_0;
	wire w_dff_A_we5WbZM39_0;
	wire w_dff_A_2CQsupRd5_0;
	wire w_dff_A_ps2xr9Xj4_0;
	wire w_dff_A_O9lqSmp91_0;
	wire w_dff_A_WVvNACZO4_0;
	wire w_dff_A_Vk368qoA7_0;
	wire w_dff_A_7zsfv1wu5_0;
	wire w_dff_A_bLGWfnQL5_0;
	wire w_dff_A_dAcC6USf3_0;
	wire w_dff_A_JIUqB4bi5_0;
	wire w_dff_A_vEfoIVrU5_0;
	wire w_dff_A_4ED88eQB2_0;
	wire w_dff_A_fptj2er38_0;
	wire w_dff_A_hPEzMaVO1_0;
	wire w_dff_A_TttMYAGY1_0;
	wire w_dff_A_0ZNHaH8t7_0;
	wire w_dff_A_1kvOQdXn9_0;
	wire w_dff_A_pxhHMs847_1;
	wire w_dff_A_VsW5jftS6_0;
	wire w_dff_A_JgySY6F13_0;
	wire w_dff_A_9sVR3Bsm9_0;
	wire w_dff_A_4IHpVARz4_0;
	wire w_dff_A_jeD6TjU52_0;
	wire w_dff_A_udeU1dBJ2_0;
	wire w_dff_A_WadM1TZy1_0;
	wire w_dff_A_iG0Oa1QY8_0;
	wire w_dff_A_yqICLXAO0_0;
	wire w_dff_A_XR9DT6Ab2_0;
	wire w_dff_A_W7zwRZey1_0;
	wire w_dff_A_5CeLt9wu6_0;
	wire w_dff_A_zCdns82z9_0;
	wire w_dff_A_o19kE1385_0;
	wire w_dff_A_CRP9tPGI1_0;
	wire w_dff_A_BYt7de0p9_0;
	wire w_dff_A_uR1WvLjb3_0;
	wire w_dff_A_3dSBGSdb4_0;
	wire w_dff_A_PYstLBrc4_0;
	wire w_dff_A_qS2eEVGC4_0;
	wire w_dff_A_rO4RnK5C1_0;
	wire w_dff_A_iTjdMU746_0;
	wire w_dff_A_iBVr8gmg1_0;
	wire w_dff_A_TNdRy4995_0;
	wire w_dff_A_bdntXmWL8_0;
	wire w_dff_A_C6YvucMg7_0;
	wire w_dff_A_5jVqDDGp3_0;
	wire w_dff_A_Ofw10gvI4_0;
	wire w_dff_A_lYmDq50Z4_0;
	wire w_dff_A_hsfvckSQ1_0;
	wire w_dff_A_LBYiaKUj8_0;
	wire w_dff_A_ecvZcZ1M3_0;
	wire w_dff_A_cK3SquUy9_0;
	wire w_dff_A_AO3odD4Z5_0;
	wire w_dff_A_pDZLOiEj7_0;
	wire w_dff_A_GjZBSWIH4_0;
	wire w_dff_A_Im9h7vRQ0_0;
	wire w_dff_A_PaiAskYr6_1;
	wire w_dff_A_PEa039RS9_0;
	wire w_dff_A_HjVD2Ytw1_0;
	wire w_dff_A_yT9STdds6_0;
	wire w_dff_A_RFgEf2nd3_0;
	wire w_dff_A_NzQEx5ya8_0;
	wire w_dff_A_kikej6Xq9_0;
	wire w_dff_A_h2d6Zx2W3_0;
	wire w_dff_A_LCDAcrbe1_0;
	wire w_dff_A_fMLPRsZ55_0;
	wire w_dff_A_7aDMI00h7_0;
	wire w_dff_A_SFh5HPZa5_0;
	wire w_dff_A_Mm7RvVhS7_0;
	wire w_dff_A_Jpov4B8I8_0;
	wire w_dff_A_cjL4xQIG5_0;
	wire w_dff_A_PSSwYHHx5_0;
	wire w_dff_A_2oZDLeZX0_0;
	wire w_dff_A_4KsZuqwr2_0;
	wire w_dff_A_iwURB6rR4_0;
	wire w_dff_A_h5hsiT301_0;
	wire w_dff_A_EAP9Fzxq8_0;
	wire w_dff_A_MTzjLy4Z3_0;
	wire w_dff_A_QyV2OEZm1_0;
	wire w_dff_A_LzccGiWz1_0;
	wire w_dff_A_4z79Vr0M3_0;
	wire w_dff_A_Mq503fkA3_0;
	wire w_dff_A_jZeqrxm32_0;
	wire w_dff_A_czPnHY5l5_0;
	wire w_dff_A_6O0aTqTv1_0;
	wire w_dff_A_pjbuSGrh8_0;
	wire w_dff_A_hCIu31mj5_0;
	wire w_dff_A_L8q86LG33_0;
	wire w_dff_A_lBlhLQ2q3_0;
	wire w_dff_A_7udL8dx51_0;
	wire w_dff_A_UKvZ8OJJ2_0;
	wire w_dff_A_XrhJPh4c1_0;
	wire w_dff_A_SPebHgFh5_0;
	wire w_dff_A_FWlxy7J35_0;
	wire w_dff_A_Nu4uyITW4_1;
	wire w_dff_A_KYGZMWuo6_0;
	wire w_dff_A_V4M1shWF4_0;
	wire w_dff_A_mYA8b5aI6_0;
	wire w_dff_A_rOxpbbnc1_0;
	wire w_dff_A_uIPU12619_0;
	wire w_dff_A_4uOo96oq0_0;
	wire w_dff_A_oUpgZ5rd5_0;
	wire w_dff_A_yN3MoL568_0;
	wire w_dff_A_Szwxe2ap6_0;
	wire w_dff_A_pMU5co2v7_0;
	wire w_dff_A_XbsXp4Hc6_0;
	wire w_dff_A_6zhj1UlZ9_0;
	wire w_dff_A_PYzorhCM0_0;
	wire w_dff_A_IpYh18977_0;
	wire w_dff_A_WJTv4oxh6_0;
	wire w_dff_A_7zD783ES2_0;
	wire w_dff_A_THVfvlSd4_0;
	wire w_dff_A_8k2dkvxx0_0;
	wire w_dff_A_pVcpbkyG8_0;
	wire w_dff_A_jcA1LeCl9_0;
	wire w_dff_A_ER5x3I9I6_0;
	wire w_dff_A_cDRioxeM9_0;
	wire w_dff_A_ABZ6XXaD7_0;
	wire w_dff_A_gZZUu6lb2_0;
	wire w_dff_A_sLQNeUj59_0;
	wire w_dff_A_ceg1PngX7_0;
	wire w_dff_A_w16ZXeoN1_0;
	wire w_dff_A_oagw8f2y1_0;
	wire w_dff_A_CqzgH1EY3_0;
	wire w_dff_A_wrhauYB39_0;
	wire w_dff_A_tQKxpYIC2_0;
	wire w_dff_A_RzdnuyV65_0;
	wire w_dff_A_aH1I6zrz7_0;
	wire w_dff_A_TRsc783g3_0;
	wire w_dff_A_im4eF1Z26_0;
	wire w_dff_A_jd4bV5Tj0_0;
	wire w_dff_A_JKCsMSY77_0;
	wire w_dff_A_Ol3YBVCw1_1;
	wire w_dff_A_3xSYrUPJ1_0;
	wire w_dff_A_SUusDXpc7_0;
	wire w_dff_A_UOfqOoHs5_0;
	wire w_dff_A_qsE9DeKb3_0;
	wire w_dff_A_HuUsKLXL9_0;
	wire w_dff_A_g31GadDR8_0;
	wire w_dff_A_FdiocZBN3_0;
	wire w_dff_A_FMYTCX8M9_0;
	wire w_dff_A_nF5Gf2cQ6_0;
	wire w_dff_A_55I86xLm8_0;
	wire w_dff_A_mACA9E8N1_0;
	wire w_dff_A_V49O5pIP8_0;
	wire w_dff_A_9SMjUDta9_0;
	wire w_dff_A_a9xdFmh85_0;
	wire w_dff_A_9lYXErQp7_0;
	wire w_dff_A_C5MZFXZ75_0;
	wire w_dff_A_bpCqdoll5_0;
	wire w_dff_A_L4yJ4DLO0_0;
	wire w_dff_A_QPFjJrQi9_0;
	wire w_dff_A_fEJvXimn8_0;
	wire w_dff_A_5IUykv0K0_0;
	wire w_dff_A_VsHqff184_0;
	wire w_dff_A_0UGzpnuI2_0;
	wire w_dff_A_zjP89fBS5_0;
	wire w_dff_A_6QF1TzX20_0;
	wire w_dff_A_jZB9fzoP3_0;
	wire w_dff_A_57zNAon70_0;
	wire w_dff_A_bwdy6hBL9_0;
	wire w_dff_A_MAliRglB3_0;
	wire w_dff_A_qiO91mHu9_0;
	wire w_dff_A_GFjYQP9P8_0;
	wire w_dff_A_8oHigkgq9_0;
	wire w_dff_A_B7zQoqDe2_0;
	wire w_dff_A_wk72eYIK2_0;
	wire w_dff_A_C0aK5UtC3_0;
	wire w_dff_A_3Ntfvrp73_0;
	wire w_dff_A_9BShlmBg5_0;
	wire w_dff_A_vskJrkeb7_1;
	wire w_dff_A_UXRGTtyt8_0;
	wire w_dff_A_IkSHepBD2_0;
	wire w_dff_A_zFEDy7cc2_0;
	wire w_dff_A_rA0VUDm33_0;
	wire w_dff_A_xiplURXD8_0;
	wire w_dff_A_8mkM6KpS5_0;
	wire w_dff_A_PR9l0QZ11_0;
	wire w_dff_A_SEXLDF4N1_0;
	wire w_dff_A_KBiiob3w8_0;
	wire w_dff_A_9WPEtNDk8_0;
	wire w_dff_A_KJ3QnQ0p9_0;
	wire w_dff_A_lktW1RCq9_0;
	wire w_dff_A_vqgQ8fcO2_0;
	wire w_dff_A_3gaC2I0l1_0;
	wire w_dff_A_u4c3Jyrf9_0;
	wire w_dff_A_e5XpNalE0_0;
	wire w_dff_A_haPEPRUE0_0;
	wire w_dff_A_5836id9O3_0;
	wire w_dff_A_DiVwlFmt9_0;
	wire w_dff_A_vTIAIXSj4_0;
	wire w_dff_A_VPgE7vpf6_0;
	wire w_dff_A_AXCSkW7H8_0;
	wire w_dff_A_GQlxiqb36_0;
	wire w_dff_A_fvYAw2d11_0;
	wire w_dff_A_fzBALfbb9_0;
	wire w_dff_A_z5Ba6lRk8_0;
	wire w_dff_A_RwwqTgD14_0;
	wire w_dff_A_JSUOVrrD5_0;
	wire w_dff_A_P6epez6C6_0;
	wire w_dff_A_wp7nBcW56_0;
	wire w_dff_A_wKKZ6bcq6_0;
	wire w_dff_A_orWLLVAh9_0;
	wire w_dff_A_oPsjac513_0;
	wire w_dff_A_onglniyU2_0;
	wire w_dff_A_eZ0JpgUC2_0;
	wire w_dff_A_ZIEpFpLb1_0;
	wire w_dff_A_JpkdzXt20_0;
	wire w_dff_A_RaK8syet9_1;
	wire w_dff_A_Pb0FOVEH6_0;
	wire w_dff_A_cNh3RjrQ9_0;
	wire w_dff_A_ubaG4VGD3_0;
	wire w_dff_A_L3uNG30D4_0;
	wire w_dff_A_IBFinrlo6_0;
	wire w_dff_A_CXm6vD924_0;
	wire w_dff_A_Ko6wFLrb9_0;
	wire w_dff_A_O95VmH619_0;
	wire w_dff_A_FuicjDch4_0;
	wire w_dff_A_9zh2Pvub1_0;
	wire w_dff_A_5B7ZAKeH5_0;
	wire w_dff_A_kyiH4Rgi2_0;
	wire w_dff_A_R6e2XuF09_0;
	wire w_dff_A_BaCSXDmo4_0;
	wire w_dff_A_xk4RxYvX4_0;
	wire w_dff_A_LcaHG0SP1_0;
	wire w_dff_A_E7OIItkO5_0;
	wire w_dff_A_TMCGoWJI1_0;
	wire w_dff_A_cRBGF4Ah5_0;
	wire w_dff_A_wAmiWsAq9_0;
	wire w_dff_A_OPHZwJFJ1_0;
	wire w_dff_A_2HsX3HrD8_0;
	wire w_dff_A_y8o5wT4a7_0;
	wire w_dff_A_ocYDhLiT6_0;
	wire w_dff_A_qdlBs3d92_0;
	wire w_dff_A_egPTUtCl0_0;
	wire w_dff_A_2qERvLwG6_0;
	wire w_dff_A_Rfq5qPW86_0;
	wire w_dff_A_PbSay1IH1_0;
	wire w_dff_A_YJjrWvDO5_0;
	wire w_dff_A_ICQVzuXr5_0;
	wire w_dff_A_PjGBXlrt5_0;
	wire w_dff_A_KEQio50c4_0;
	wire w_dff_A_cw6n8IGT6_0;
	wire w_dff_A_SOWjsBFD4_0;
	wire w_dff_A_e5wWdgSw4_0;
	wire w_dff_A_kzLLaeop0_0;
	wire w_dff_A_rcmF46MD0_1;
	wire w_dff_A_TIKAjhuU9_0;
	wire w_dff_A_ZRN1dQRs5_0;
	wire w_dff_A_myDFnknc2_0;
	wire w_dff_A_Pr60PBI84_0;
	wire w_dff_A_v9xMhqA74_0;
	wire w_dff_A_sTaudX3u8_0;
	wire w_dff_A_WkRKEYxj7_0;
	wire w_dff_A_8p3Y9tIm7_0;
	wire w_dff_A_63qalUZc9_0;
	wire w_dff_A_Y0gpKUP46_0;
	wire w_dff_A_Nl6H9Dbz0_0;
	wire w_dff_A_VBNYUmul2_0;
	wire w_dff_A_OZfGCYwu9_0;
	wire w_dff_A_cJtEl5kD8_0;
	wire w_dff_A_iEHPrY3h4_0;
	wire w_dff_A_hmaNOJpJ2_0;
	wire w_dff_A_UPoEbzff2_0;
	wire w_dff_A_JGzFKfVt4_0;
	wire w_dff_A_RAiL0qDq9_0;
	wire w_dff_A_xq0VoqIJ2_0;
	wire w_dff_A_OyMd5xR60_0;
	wire w_dff_A_JmEGPCpi9_0;
	wire w_dff_A_gJSuG6s35_0;
	wire w_dff_A_ARddEvWE7_0;
	wire w_dff_A_DbDzDBwI0_0;
	wire w_dff_A_Lupy8mqA7_0;
	wire w_dff_A_0VTU5TVu6_0;
	wire w_dff_A_SDITtrK46_0;
	wire w_dff_A_FVF7AGru3_0;
	wire w_dff_A_ICynjAzX7_0;
	wire w_dff_A_66klPyMA8_0;
	wire w_dff_A_V3PxxPoI9_0;
	wire w_dff_A_1cnWBF4V9_0;
	wire w_dff_A_ycaRZFlL9_0;
	wire w_dff_A_pbDOYEnG0_0;
	wire w_dff_A_bX0Ptm3l1_0;
	wire w_dff_A_ObZeEgSA1_0;
	wire w_dff_A_dxxPtiY89_1;
	wire w_dff_A_G97i5TXp7_0;
	wire w_dff_A_VHRF8OEO2_0;
	wire w_dff_A_I3eEu5BT4_0;
	wire w_dff_A_0ANP60F64_0;
	wire w_dff_A_PmBYg4Oq2_0;
	wire w_dff_A_XfqgMaMf9_0;
	wire w_dff_A_QdgbZmrm1_0;
	wire w_dff_A_b1Dk2QaW7_0;
	wire w_dff_A_yuhXJrgn8_0;
	wire w_dff_A_wxgERnc01_0;
	wire w_dff_A_T692Kb5M9_0;
	wire w_dff_A_E21QNLKS4_0;
	wire w_dff_A_W4iO5Nsn4_0;
	wire w_dff_A_eGycNfi15_0;
	wire w_dff_A_nW0dzScY3_0;
	wire w_dff_A_Outscrxx1_0;
	wire w_dff_A_VMIh675L0_0;
	wire w_dff_A_ORckzife0_0;
	wire w_dff_A_uxMBtKj98_0;
	wire w_dff_A_EvTsR43w5_0;
	wire w_dff_A_POHudtj46_0;
	wire w_dff_A_Cn5eg88Q0_0;
	wire w_dff_A_kCv8v0yV1_0;
	wire w_dff_A_BkYbtoU89_0;
	wire w_dff_A_2s01hytV1_0;
	wire w_dff_A_x0MQOnZ92_0;
	wire w_dff_A_YFmCDhea8_0;
	wire w_dff_A_JE7Bxocw3_0;
	wire w_dff_A_MSq3OtVs5_0;
	wire w_dff_A_LVicT9iL1_0;
	wire w_dff_A_yykhCNPr0_0;
	wire w_dff_A_kbhJRXdQ6_0;
	wire w_dff_A_2tqiUYdu1_0;
	wire w_dff_A_DKAYhMC89_0;
	wire w_dff_A_bjHWOuXD7_0;
	wire w_dff_A_RDsF7P6a8_0;
	wire w_dff_A_QYJkjfVl0_0;
	wire w_dff_A_k9lEreo95_1;
	wire w_dff_A_0nwAKcp88_0;
	wire w_dff_A_jGNhNoDc3_0;
	wire w_dff_A_ejCxPrz08_0;
	wire w_dff_A_w4MTPZZ84_0;
	wire w_dff_A_Sgf2csNq0_0;
	wire w_dff_A_8cjCODhm6_0;
	wire w_dff_A_DreVlXB93_0;
	wire w_dff_A_QvaNNxVW7_0;
	wire w_dff_A_Eae8EmhX1_0;
	wire w_dff_A_KDUKBNT96_0;
	wire w_dff_A_CJS2jRgH4_0;
	wire w_dff_A_0pg6gr2N2_0;
	wire w_dff_A_rUgAKxQk2_0;
	wire w_dff_A_F62ckR6d5_0;
	wire w_dff_A_hqze5srK4_0;
	wire w_dff_A_DYinpXFB0_0;
	wire w_dff_A_USTYARax8_0;
	wire w_dff_A_weaCHrdm0_0;
	wire w_dff_A_lIvf3hr91_0;
	wire w_dff_A_uy2MvhMz9_0;
	wire w_dff_A_4Non3de70_0;
	wire w_dff_A_MPeLjYBn4_0;
	wire w_dff_A_VpYkl1ja7_0;
	wire w_dff_A_uRS1m2v22_0;
	wire w_dff_A_dcCxrZNW1_0;
	wire w_dff_A_Zx2B5KrL4_0;
	wire w_dff_A_qJJSCMbZ0_0;
	wire w_dff_A_XFyMPW0X9_0;
	wire w_dff_A_B7epnpWG3_0;
	wire w_dff_A_JUZHmBjy2_0;
	wire w_dff_A_VXZs3TAF0_0;
	wire w_dff_A_MAqTSXBt9_0;
	wire w_dff_A_QOjK9iD20_0;
	wire w_dff_A_U2EDWbT94_0;
	wire w_dff_A_KkTw2BSX2_0;
	wire w_dff_A_CP1kEolh0_0;
	wire w_dff_A_19ElGh7A7_0;
	wire w_dff_A_OvoAegEm6_1;
	wire w_dff_A_ydkyoe2X6_0;
	wire w_dff_A_wh0eUoIo5_0;
	wire w_dff_A_7d98hpyX4_0;
	wire w_dff_A_rgZN6Zkb7_0;
	wire w_dff_A_xVug889p9_0;
	wire w_dff_A_ZZBzL6wA1_0;
	wire w_dff_A_GpDI3p6U6_0;
	wire w_dff_A_aVuUX56V4_0;
	wire w_dff_A_qwj7MtCH2_0;
	wire w_dff_A_X6n74ntP7_0;
	wire w_dff_A_M2xpWZOp0_0;
	wire w_dff_A_KrfvbOPY0_0;
	wire w_dff_A_mZ4nhya30_0;
	wire w_dff_A_KhIoE2iT8_0;
	wire w_dff_A_Ujr24iPF8_0;
	wire w_dff_A_B8fAShn17_0;
	wire w_dff_A_Ih6dd4rl0_0;
	wire w_dff_A_raRKZkES9_0;
	wire w_dff_A_yIUv6Glp2_0;
	wire w_dff_A_NWV0efjI5_0;
	wire w_dff_A_5vsPEcrY6_0;
	wire w_dff_A_yuhaGSUP4_0;
	wire w_dff_A_WbIpVahl1_0;
	wire w_dff_A_5nQjm3KJ8_0;
	wire w_dff_A_mbRarS1g5_0;
	wire w_dff_A_N5QgfnDu5_0;
	wire w_dff_A_Pb2yFNHE9_0;
	wire w_dff_A_Czc2e6Vp5_0;
	wire w_dff_A_hKmT7x8c4_0;
	wire w_dff_A_DDidJ2n95_0;
	wire w_dff_A_I59aTpTO1_0;
	wire w_dff_A_18OEmnbb0_0;
	wire w_dff_A_L3RXcbDh0_0;
	wire w_dff_A_4I5IVXMF3_0;
	wire w_dff_A_EWOwMrOK0_0;
	wire w_dff_A_0VpkrRIy8_0;
	wire w_dff_A_y10T6j0N4_0;
	wire w_dff_A_tWFx69fK7_1;
	wire w_dff_A_rBXTNuUt5_0;
	wire w_dff_A_o1iutIEO7_0;
	wire w_dff_A_gOWLBNeg9_0;
	wire w_dff_A_UGtPa2xC2_0;
	wire w_dff_A_nNwuuTzu5_0;
	wire w_dff_A_cqqhmPMK6_0;
	wire w_dff_A_ikMW08vh6_0;
	wire w_dff_A_RU6Ktixm8_0;
	wire w_dff_A_RlfKC6hj9_0;
	wire w_dff_A_fNk6dXlS5_0;
	wire w_dff_A_EYhkACvk6_0;
	wire w_dff_A_KdJX0QZ25_0;
	wire w_dff_A_TV58zjAa9_0;
	wire w_dff_A_zBTMu70L5_0;
	wire w_dff_A_EsETY64J9_0;
	wire w_dff_A_xvGjPyfh0_0;
	wire w_dff_A_65jCh6314_0;
	wire w_dff_A_yY971RDm1_0;
	wire w_dff_A_wcM56EJB3_0;
	wire w_dff_A_tFAjRxPB6_0;
	wire w_dff_A_QHXXRhc95_0;
	wire w_dff_A_FzEdkxbu0_0;
	wire w_dff_A_dmwX4KAX6_0;
	wire w_dff_A_LZUxxINK8_0;
	wire w_dff_A_XqCnE4RS6_0;
	wire w_dff_A_234JKLKH4_0;
	wire w_dff_A_g1iWwlxg0_0;
	wire w_dff_A_OyIrr8827_0;
	wire w_dff_A_6vm2bBBs2_0;
	wire w_dff_A_W5AHB6tU7_0;
	wire w_dff_A_dQ0E8VZA2_0;
	wire w_dff_A_OTO4CLrO6_0;
	wire w_dff_A_hBNXpWWr1_0;
	wire w_dff_A_k2jTy2Qw9_0;
	wire w_dff_A_JtbBrwXu8_0;
	wire w_dff_A_PxN5ufQQ4_0;
	wire w_dff_A_IRFD80KQ9_0;
	wire w_dff_A_WpSOD8rp3_1;
	wire w_dff_A_CdT4sQSo2_0;
	wire w_dff_A_HMHE3DiA7_0;
	wire w_dff_A_x67nYRTP7_0;
	wire w_dff_A_mcfY7cTk4_0;
	wire w_dff_A_fSiYOQJI0_0;
	wire w_dff_A_38EpSSyU5_0;
	wire w_dff_A_g6CO0Dzi9_0;
	wire w_dff_A_00OqCLVW3_0;
	wire w_dff_A_TsAWrXEj4_0;
	wire w_dff_A_IlTOizfN3_0;
	wire w_dff_A_RISActYd1_0;
	wire w_dff_A_H5j4OuP52_0;
	wire w_dff_A_adGiQ2RC5_0;
	wire w_dff_A_FiyPuiCJ2_0;
	wire w_dff_A_XFCBeme97_0;
	wire w_dff_A_CkcwRHEs5_0;
	wire w_dff_A_Tv2cXZev3_0;
	wire w_dff_A_J507qUcA2_0;
	wire w_dff_A_MEHbksYP3_0;
	wire w_dff_A_GjJV2pwR2_0;
	wire w_dff_A_a93uWquw8_0;
	wire w_dff_A_eYCmwouk4_0;
	wire w_dff_A_AFiznRLh2_0;
	wire w_dff_A_h5VXymDw1_0;
	wire w_dff_A_TZ63m7H05_0;
	wire w_dff_A_hrfWgdWW8_0;
	wire w_dff_A_UgHRdBhH4_0;
	wire w_dff_A_B6M3UwiU8_0;
	wire w_dff_A_FR305U978_0;
	wire w_dff_A_GWB1OvPB0_0;
	wire w_dff_A_1KLeYKf19_0;
	wire w_dff_A_pA7G6NbE5_0;
	wire w_dff_A_FOwIA3GO4_0;
	wire w_dff_A_3Lcnqqwp8_0;
	wire w_dff_A_qi1yUlle9_0;
	wire w_dff_A_g93qrmQt4_0;
	wire w_dff_A_lMOuGJNH0_0;
	wire w_dff_A_0Bt12MFX2_1;
	wire w_dff_A_rz54Zfzl8_0;
	wire w_dff_A_QOlJGFcz9_0;
	wire w_dff_A_mMDuSWno3_0;
	wire w_dff_A_HKdk1ZV48_0;
	wire w_dff_A_u2bfEMbj0_0;
	wire w_dff_A_wn1z2M069_0;
	wire w_dff_A_BQyIudlE2_0;
	wire w_dff_A_UuF8KJMG0_0;
	wire w_dff_A_vrQXckRA3_0;
	wire w_dff_A_htRr66EF8_0;
	wire w_dff_A_tPtjB26c0_0;
	wire w_dff_A_A0nrnv027_0;
	wire w_dff_A_cBlnpneQ5_0;
	wire w_dff_A_sGINlGaG2_0;
	wire w_dff_A_9ejt6TRu9_0;
	wire w_dff_A_FTc2yuNf2_0;
	wire w_dff_A_Qo0qyAeu0_0;
	wire w_dff_A_GYg1aoAD3_0;
	wire w_dff_A_oUYbyAmX5_0;
	wire w_dff_A_v2oLe0R57_0;
	wire w_dff_A_wfmD05pD2_0;
	wire w_dff_A_Q70oevZG8_0;
	wire w_dff_A_j9sDj5rm9_0;
	wire w_dff_A_W7AnjYws3_0;
	wire w_dff_A_Y0mNZce09_0;
	wire w_dff_A_hQAGEpKD2_0;
	wire w_dff_A_vQBBfBVH8_0;
	wire w_dff_A_LpnxXwLD7_0;
	wire w_dff_A_MWFhbBBb3_0;
	wire w_dff_A_Ns6dSFxd8_0;
	wire w_dff_A_A3DMHh212_0;
	wire w_dff_A_Gorq8wbJ5_0;
	wire w_dff_A_WotqE8j32_0;
	wire w_dff_A_wD6MLlh62_0;
	wire w_dff_A_IHPxW33Q6_0;
	wire w_dff_A_thYjKvrw5_0;
	wire w_dff_A_SfYhXbFh8_0;
	wire w_dff_A_Btoykzj63_1;
	wire w_dff_A_DBPTFWA46_0;
	wire w_dff_A_1iZsiXTt0_0;
	wire w_dff_A_10uOhHhX1_0;
	wire w_dff_A_BKq4JrHR1_0;
	wire w_dff_A_Ptj17vIZ4_0;
	wire w_dff_A_7lme9fO97_0;
	wire w_dff_A_6QkS7RX48_0;
	wire w_dff_A_GO9a7j7J8_0;
	wire w_dff_A_93u88cEs6_0;
	wire w_dff_A_05SoZ6GH4_0;
	wire w_dff_A_MS2eqpsR2_0;
	wire w_dff_A_PXDy0tFB9_0;
	wire w_dff_A_GvDIfDeg8_0;
	wire w_dff_A_BvgvXHtP6_0;
	wire w_dff_A_tDA1uXjO3_0;
	wire w_dff_A_uJD1uhaZ6_0;
	wire w_dff_A_l6BGa1Kh6_0;
	wire w_dff_A_1h69Ug5y4_0;
	wire w_dff_A_lGcKFsVI7_0;
	wire w_dff_A_gP1jGYPA2_0;
	wire w_dff_A_9pX1HmKe5_0;
	wire w_dff_A_OgPKySg30_0;
	wire w_dff_A_WW5Y83WK3_0;
	wire w_dff_A_fb7eTxiX1_0;
	wire w_dff_A_tuH7XCB63_0;
	wire w_dff_A_eJFWAKch7_0;
	wire w_dff_A_2cYrZ14W2_0;
	wire w_dff_A_Gzc1oqwx2_0;
	wire w_dff_A_sJdCtwPd5_0;
	wire w_dff_A_UkTyILvP7_0;
	wire w_dff_A_1WsKbfvO8_0;
	wire w_dff_A_cSIiDGfg7_0;
	wire w_dff_A_uTekU42l4_0;
	wire w_dff_A_lxZTtf413_0;
	wire w_dff_A_86D7dpH85_0;
	wire w_dff_A_phxFdKTc5_0;
	wire w_dff_A_wiS1sg8g9_0;
	wire w_dff_A_Mp0c0e9T0_1;
	wire w_dff_A_QAN1kA3n9_0;
	wire w_dff_A_ZLWJaSWH5_0;
	wire w_dff_A_9iINOz5i0_0;
	wire w_dff_A_UHSRuxXA0_0;
	wire w_dff_A_bobjiQpk6_0;
	wire w_dff_A_06zGBEtv9_0;
	wire w_dff_A_zawuMBcn0_0;
	wire w_dff_A_LHrGMtDa1_0;
	wire w_dff_A_YmhHv6QF0_0;
	wire w_dff_A_vZ6Yf7Ir1_0;
	wire w_dff_A_UW4jf6w40_0;
	wire w_dff_A_1vubCZQV2_0;
	wire w_dff_A_jrvG67F59_0;
	wire w_dff_A_gK1eM2kv2_0;
	wire w_dff_A_IIAWXZjE5_0;
	wire w_dff_A_Cwa9wFxL1_0;
	wire w_dff_A_nA96BF973_0;
	wire w_dff_A_V3UQUgxY9_0;
	wire w_dff_A_E4GdjO9Q8_0;
	wire w_dff_A_tAHhD5eq9_0;
	wire w_dff_A_bHB88nvE1_0;
	wire w_dff_A_9XwpDm3b1_0;
	wire w_dff_A_kCFIHhXa8_0;
	wire w_dff_A_tOIP03Re8_0;
	wire w_dff_A_dyv9nxPW5_0;
	wire w_dff_A_xKrQk2kV3_0;
	wire w_dff_A_aa9KrGIT1_0;
	wire w_dff_A_kbFOTB0W7_0;
	wire w_dff_A_69HdGNk67_0;
	wire w_dff_A_1YYDhmyB3_0;
	wire w_dff_A_lOghKWBG3_0;
	wire w_dff_A_CcIk14aE8_0;
	wire w_dff_A_qh42paZS2_0;
	wire w_dff_A_9kBu6i9W7_0;
	wire w_dff_A_RkerbP610_0;
	wire w_dff_A_Pzq9DuDH9_0;
	wire w_dff_A_qWJuqif76_0;
	wire w_dff_A_ReeCzHam0_1;
	wire w_dff_A_VAtd6ojO6_0;
	wire w_dff_A_fgLIz7579_0;
	wire w_dff_A_e6psGgm19_0;
	wire w_dff_A_HU1Er5R40_0;
	wire w_dff_A_p0ejQOe19_0;
	wire w_dff_A_OakH9ahz8_0;
	wire w_dff_A_namE0PEt9_0;
	wire w_dff_A_bKBHiHXY7_0;
	wire w_dff_A_5JS1xSX60_0;
	wire w_dff_A_BdGG74w49_0;
	wire w_dff_A_LxevbDgk3_0;
	wire w_dff_A_dyX5QeVm6_0;
	wire w_dff_A_7wrVGsvS6_0;
	wire w_dff_A_mdvTV2M94_0;
	wire w_dff_A_ZOXB797B5_0;
	wire w_dff_A_XqDhwwTU2_0;
	wire w_dff_A_FN2meJcS4_0;
	wire w_dff_A_UWDI1rcn2_0;
	wire w_dff_A_nQ5FjT9j2_0;
	wire w_dff_A_VMdq6R6P3_0;
	wire w_dff_A_UcPK5xLx8_0;
	wire w_dff_A_VaMgQ7rf1_0;
	wire w_dff_A_3KRlIzmx2_0;
	wire w_dff_A_1iZOStDw8_0;
	wire w_dff_A_WlBN6Pna2_0;
	wire w_dff_A_wYWfktBK4_0;
	wire w_dff_A_c278mtd82_0;
	wire w_dff_A_6Kt4kC7J3_0;
	wire w_dff_A_JxCayiBq8_0;
	wire w_dff_A_2EzZnyBp1_0;
	wire w_dff_A_tJsHhYII5_0;
	wire w_dff_A_BDPAqsf18_0;
	wire w_dff_A_LDtMW9hx8_0;
	wire w_dff_A_9K7Cq7G98_0;
	wire w_dff_A_vSWIXsnq3_0;
	wire w_dff_A_JsxhfXln5_0;
	wire w_dff_A_R8bl4UCH7_0;
	wire w_dff_A_wNDkqV9X6_1;
	wire w_dff_A_r0WQzJi04_0;
	wire w_dff_A_L7TZ5b2t1_0;
	wire w_dff_A_S8GueEaO6_0;
	wire w_dff_A_d2iAScxU8_0;
	wire w_dff_A_PeyvzLzQ4_0;
	wire w_dff_A_ajzfxveW1_0;
	wire w_dff_A_Iy9YAmz36_0;
	wire w_dff_A_W35tNQns1_0;
	wire w_dff_A_lWT33Ufv7_0;
	wire w_dff_A_ScI156pN7_0;
	wire w_dff_A_FAqIWjmC6_0;
	wire w_dff_A_fyOoPG2X5_0;
	wire w_dff_A_3OgmrwKD1_0;
	wire w_dff_A_Fs0ju9HF8_0;
	wire w_dff_A_uCWLPIYQ2_0;
	wire w_dff_A_LW9T8MCW7_0;
	wire w_dff_A_IYKKslCv1_0;
	wire w_dff_A_4nNAy4ns5_0;
	wire w_dff_A_oCRZZGWp7_0;
	wire w_dff_A_XsdgfgUC7_0;
	wire w_dff_A_xABX73f49_0;
	wire w_dff_A_zyGl4EHl4_0;
	wire w_dff_A_e3Ydfltt6_0;
	wire w_dff_A_Y83BffQe9_0;
	wire w_dff_A_sKtdNFkT7_0;
	wire w_dff_A_tJtXXvJM5_0;
	wire w_dff_A_stbY7ACb3_0;
	wire w_dff_A_mHiYY7PV6_0;
	wire w_dff_A_pxrAQ3mi1_0;
	wire w_dff_A_vDJsEelS6_0;
	wire w_dff_A_nMMYk4NR7_0;
	wire w_dff_A_f6L6XOUy6_0;
	wire w_dff_A_7l4D5zCO0_0;
	wire w_dff_A_TooqVmUK2_0;
	wire w_dff_A_fTxHXQjX8_0;
	wire w_dff_A_HTCSvGZZ3_0;
	wire w_dff_A_4hC2oC508_0;
	wire w_dff_A_TnC3fYtR3_1;
	wire w_dff_A_OusjvvD54_0;
	wire w_dff_A_X91AlhYc5_0;
	wire w_dff_A_MyYDfWOG7_0;
	wire w_dff_A_Ugd1jy1D7_0;
	wire w_dff_A_DkDYaxly0_0;
	wire w_dff_A_CUQTXiKE8_0;
	wire w_dff_A_7NUqq3zw5_0;
	wire w_dff_A_vLtl5ggm3_0;
	wire w_dff_A_njdB9fOO3_0;
	wire w_dff_A_fCkscxnd0_0;
	wire w_dff_A_IqkPXJAb0_0;
	wire w_dff_A_er7grrb98_0;
	wire w_dff_A_OKNEDAyD6_0;
	wire w_dff_A_aaO32Qjc1_0;
	wire w_dff_A_j6ckGRFj5_0;
	wire w_dff_A_j9CNGlJS8_0;
	wire w_dff_A_qJBXjZCB1_0;
	wire w_dff_A_K2dViIzc0_0;
	wire w_dff_A_RxcO7qo52_0;
	wire w_dff_A_RUL3SLqx6_0;
	wire w_dff_A_DlqLsbAj3_0;
	wire w_dff_A_VAF0i8ZA2_0;
	wire w_dff_A_aWDQUBIU0_0;
	wire w_dff_A_ojutfHwt4_0;
	wire w_dff_A_mPYCv19x1_0;
	wire w_dff_A_8hb3iYw81_0;
	wire w_dff_A_3zIjocPC5_0;
	wire w_dff_A_PypNKC9r3_0;
	wire w_dff_A_xW0JxjF53_0;
	wire w_dff_A_4VMtYlsa4_0;
	wire w_dff_A_ivYYIrsJ4_0;
	wire w_dff_A_ftxL8Nqp4_0;
	wire w_dff_A_q3D0uZNR4_0;
	wire w_dff_A_wB1HIsRx4_0;
	wire w_dff_A_TqJ2Mjfy5_0;
	wire w_dff_A_Uj2ECwpB9_0;
	wire w_dff_A_Xetz9aSM4_0;
	wire w_dff_A_3rxkWg5S9_1;
	wire w_dff_A_LE2rjmPW1_0;
	wire w_dff_A_QytUHVI58_0;
	wire w_dff_A_KorsMJiw9_0;
	wire w_dff_A_pgbKMHN99_0;
	wire w_dff_A_BXE8Vq7z6_0;
	wire w_dff_A_04mTBibP3_0;
	wire w_dff_A_KaB9jzjV7_0;
	wire w_dff_A_9pC5nFss3_0;
	wire w_dff_A_CwEBZBp51_0;
	wire w_dff_A_l9Vh7Do05_0;
	wire w_dff_A_vOvfAFlI4_0;
	wire w_dff_A_YIdbzm4r7_0;
	wire w_dff_A_mZUaz71h5_0;
	wire w_dff_A_HPPW8HyZ8_0;
	wire w_dff_A_wR0eZlHq0_0;
	wire w_dff_A_rimFFKaY6_0;
	wire w_dff_A_RkKW1rvY3_0;
	wire w_dff_A_QhWst42O8_0;
	wire w_dff_A_PKO1MUXk5_0;
	wire w_dff_A_OwNzPaYB5_0;
	wire w_dff_A_7UITA4t27_0;
	wire w_dff_A_CXJqxKHW3_0;
	wire w_dff_A_I73LU5FT4_0;
	wire w_dff_A_4ltZu5ML1_0;
	wire w_dff_A_9Tkyn4VC7_0;
	wire w_dff_A_Lg4ALZlf9_0;
	wire w_dff_A_hKpMjOIw7_0;
	wire w_dff_A_nLo2os3J5_0;
	wire w_dff_A_KA2T3DwW2_0;
	wire w_dff_A_f4BbQmFp5_0;
	wire w_dff_A_K06CakgD0_0;
	wire w_dff_A_eKKYvRWU5_0;
	wire w_dff_A_YHgJ9OAa6_0;
	wire w_dff_A_qtR2F5Pr4_0;
	wire w_dff_A_zKxJyPZ97_0;
	wire w_dff_A_xK5nuJMO5_0;
	wire w_dff_A_NIFIvBQ92_0;
	wire w_dff_A_VGhsnYzH9_1;
	wire w_dff_A_k0kxFyxg5_0;
	wire w_dff_A_0Kub6lVs4_0;
	wire w_dff_A_vpkqxgEZ9_0;
	wire w_dff_A_3D01UMmf6_0;
	wire w_dff_A_EHtETE1Z0_0;
	wire w_dff_A_Pv3fbyyt1_0;
	wire w_dff_A_4E9fniZY7_0;
	wire w_dff_A_MYc4JEl05_0;
	wire w_dff_A_oe8rHOUi9_0;
	wire w_dff_A_OWaAt6vZ5_0;
	wire w_dff_A_jkL1XRRL0_0;
	wire w_dff_A_pOnNXAhg8_0;
	wire w_dff_A_MNOt3Rpk5_0;
	wire w_dff_A_8bnmCgFn2_0;
	wire w_dff_A_GFqcIxkx0_0;
	wire w_dff_A_hK3okQKZ0_0;
	wire w_dff_A_6zYNJLny9_0;
	wire w_dff_A_MEoDZomE2_0;
	wire w_dff_A_JnNj51JT8_0;
	wire w_dff_A_JprOozQS7_0;
	wire w_dff_A_Ip0iVPii6_0;
	wire w_dff_A_R0sbkSL78_0;
	wire w_dff_A_tllcEnYY0_0;
	wire w_dff_A_0tEM0fhe1_0;
	wire w_dff_A_SMqhLXjc6_0;
	wire w_dff_A_qgBiWEHo1_0;
	wire w_dff_A_Fp9Uf06n7_0;
	wire w_dff_A_nSo6I93q6_0;
	wire w_dff_A_acXF0J0C6_0;
	wire w_dff_A_VCkrEa8s3_0;
	wire w_dff_A_dJHNVGkm4_0;
	wire w_dff_A_cgUuihUD0_0;
	wire w_dff_A_ntG72hgR0_0;
	wire w_dff_A_uYXQn4582_0;
	wire w_dff_A_28I0bMga3_0;
	wire w_dff_A_FIyxzINt4_0;
	wire w_dff_A_dMSxsxpb2_0;
	wire w_dff_A_JFXSKKkp5_1;
	wire w_dff_A_KmRG8YSZ8_0;
	wire w_dff_A_Hmd9HzlN3_0;
	wire w_dff_A_cjGxqako2_0;
	wire w_dff_A_tyW7NXjR8_0;
	wire w_dff_A_aWyQiUHD4_0;
	wire w_dff_A_CBYYRz818_0;
	wire w_dff_A_Rf3WrN775_0;
	wire w_dff_A_tgxb4eBv7_0;
	wire w_dff_A_astaUZVK0_0;
	wire w_dff_A_EbzHxp4j0_0;
	wire w_dff_A_TbGuQqq25_0;
	wire w_dff_A_dns6CZ698_0;
	wire w_dff_A_5nmK8d0p2_0;
	wire w_dff_A_OQJ8q4XR8_0;
	wire w_dff_A_AWSAZYem2_0;
	wire w_dff_A_k3YahAFL4_0;
	wire w_dff_A_56F7Au5a4_0;
	wire w_dff_A_zlQKHLze9_0;
	wire w_dff_A_kxFPVAmC5_0;
	wire w_dff_A_cUiNiaLE9_0;
	wire w_dff_A_LqlnNlhh8_0;
	wire w_dff_A_EoJ7s8AD2_0;
	wire w_dff_A_XVGMf8mF1_0;
	wire w_dff_A_xhiXXSCI6_0;
	wire w_dff_A_RsnUzjIM7_0;
	wire w_dff_A_nubtNemo2_0;
	wire w_dff_A_nEZtyRX62_0;
	wire w_dff_A_ME7rmiYF4_0;
	wire w_dff_A_Z058oID48_0;
	wire w_dff_A_wOc3JKWb7_0;
	wire w_dff_A_oIxqCI0V0_0;
	wire w_dff_A_i0LZDUdt2_0;
	wire w_dff_A_WHKvjddF5_0;
	wire w_dff_A_m07byV5r5_0;
	wire w_dff_A_0Lf6114F7_0;
	wire w_dff_A_MEU3uGmb7_0;
	wire w_dff_A_Vj3nW6U86_0;
	wire w_dff_A_158BVJfx5_2;
	wire w_dff_A_CLL2gg4d5_0;
	wire w_dff_A_9oE5xXgH8_0;
	wire w_dff_A_5Dm0OX310_0;
	wire w_dff_A_xacIzu1s5_0;
	wire w_dff_A_pemjsvk11_0;
	wire w_dff_A_VZZHPRUb7_0;
	wire w_dff_A_CFT6vBDo3_0;
	wire w_dff_A_b8zK4la92_0;
	wire w_dff_A_3Xb9YTFB0_0;
	wire w_dff_A_3sKgfhgL1_0;
	wire w_dff_A_miJLNjiY1_0;
	wire w_dff_A_Ih7lLUxj2_0;
	wire w_dff_A_wZ1HvS8d8_0;
	wire w_dff_A_8D0Z7R2P1_0;
	wire w_dff_A_ku5aXqcm2_0;
	wire w_dff_A_j4LrhcMD0_0;
	wire w_dff_A_RCMzzZ511_0;
	wire w_dff_A_ZmeHSxo71_0;
	wire w_dff_A_MNGIbMlA0_0;
	wire w_dff_A_EySmUv1b4_0;
	wire w_dff_A_fkQkFkf26_0;
	wire w_dff_A_QC3yvEuU0_0;
	wire w_dff_A_mOYl6UFY1_0;
	wire w_dff_A_nh36QvYs6_0;
	wire w_dff_A_etqlJ6TU7_0;
	wire w_dff_A_NjIgqH7Q1_0;
	wire w_dff_A_TGmHPZnS2_0;
	wire w_dff_A_EEN8P03i3_0;
	wire w_dff_A_rl3A3UPi4_0;
	wire w_dff_A_bYRWAxlR4_0;
	wire w_dff_A_o4VX0bgv8_0;
	wire w_dff_A_iRGSMRKl2_0;
	wire w_dff_A_Md8CSjuT2_0;
	wire w_dff_A_sYVzjdXt8_0;
	wire w_dff_A_J7k3LctK6_0;
	wire w_dff_A_FVVC0TFo0_0;
	wire w_dff_A_kWgYBNDK3_0;
	wire w_dff_A_GynMmCSi4_1;
	wire w_dff_A_vj1i6Q4W4_0;
	wire w_dff_A_9iyTVvLU4_0;
	wire w_dff_A_BIS7cSYb4_0;
	wire w_dff_A_DSrrF1LD0_0;
	wire w_dff_A_VIcrETCE7_0;
	wire w_dff_A_ZWUV3q6f1_0;
	wire w_dff_A_TJ3rlJPR7_0;
	wire w_dff_A_88fEcWo73_0;
	wire w_dff_A_e4qr6Kim1_0;
	wire w_dff_A_DIRzeKGR5_0;
	wire w_dff_A_qqwVFXsz4_0;
	wire w_dff_A_xqHEpXaw2_0;
	wire w_dff_A_WY0X2efS1_0;
	wire w_dff_A_hJ3ZGWct2_0;
	wire w_dff_A_nawroWYY6_0;
	wire w_dff_A_aTs9Zv9f3_0;
	wire w_dff_A_q8GdOi1s4_0;
	wire w_dff_A_VvfLsch44_0;
	wire w_dff_A_XimVxw858_0;
	wire w_dff_A_667T2w5h1_0;
	wire w_dff_A_HR4KjMBJ0_0;
	wire w_dff_A_0RwHo2li2_0;
	wire w_dff_A_JcJogVNy6_0;
	wire w_dff_A_YAUbcyV69_0;
	wire w_dff_A_Gs4iSEBu7_0;
	wire w_dff_A_Pkj2Y5nd5_0;
	wire w_dff_A_WFMLinim1_0;
	wire w_dff_A_RcIwekHA4_0;
	wire w_dff_A_0xaU0Cuh0_0;
	wire w_dff_A_HTAEPPW28_0;
	wire w_dff_A_Rdlf2Vif7_0;
	wire w_dff_A_PXw3ExlL2_0;
	wire w_dff_A_aCpWcBb56_0;
	wire w_dff_A_CpcPe3Hn7_0;
	wire w_dff_A_ao8jql5i9_0;
	wire w_dff_A_QtSapZun2_1;
	wire w_dff_A_Ni8tMVZk0_0;
	wire w_dff_A_Yr13wJqq8_0;
	wire w_dff_A_5HzB6MDS0_0;
	wire w_dff_A_Mmh4FKkW1_0;
	wire w_dff_A_NUUm0Deu7_0;
	wire w_dff_A_Eg47cOYr6_0;
	wire w_dff_A_DHI7KS9M8_0;
	wire w_dff_A_vF4yevS25_0;
	wire w_dff_A_a2Re9Td98_0;
	wire w_dff_A_rtUhi4762_0;
	wire w_dff_A_9rU4JBHW4_0;
	wire w_dff_A_EbPVg9GJ5_0;
	wire w_dff_A_tXaxjFRS5_0;
	wire w_dff_A_1etpoojM9_0;
	wire w_dff_A_ffGf5HGF1_0;
	wire w_dff_A_mdA6x57w6_0;
	wire w_dff_A_pM1xlMzH9_0;
	wire w_dff_A_BQVMZrRw0_0;
	wire w_dff_A_qB8ix4dM5_0;
	wire w_dff_A_UckGQ84b8_0;
	wire w_dff_A_3DyiCViY7_0;
	wire w_dff_A_lI64x69H9_0;
	wire w_dff_A_xABE00sC0_0;
	wire w_dff_A_9ifPF6r31_0;
	wire w_dff_A_aUxtXqlF6_0;
	wire w_dff_A_rsRX30xy1_0;
	wire w_dff_A_FHMB4Ax24_0;
	wire w_dff_A_4XAdbL8E9_0;
	wire w_dff_A_61Kaltr52_0;
	wire w_dff_A_xLSKHv535_0;
	wire w_dff_A_QUvfsMu10_0;
	wire w_dff_A_k9lcU8oD2_0;
	wire w_dff_A_SeTd8ZPF5_0;
	wire w_dff_A_G0pdch835_0;
	wire w_dff_A_1efeAtYx5_0;
	wire w_dff_A_iYRibRUl1_1;
	wire w_dff_A_DtfApZ644_0;
	wire w_dff_A_spBeFz7Q1_0;
	wire w_dff_A_zggI7YUb0_0;
	wire w_dff_A_uqnBezBm3_0;
	wire w_dff_A_4M7CeSQk3_0;
	wire w_dff_A_DJ6AhKP72_0;
	wire w_dff_A_BFztI4Bh1_0;
	wire w_dff_A_cqJA7KfR5_0;
	wire w_dff_A_zsGQi5M20_0;
	wire w_dff_A_UlVdO9237_0;
	wire w_dff_A_wUk8zebQ7_0;
	wire w_dff_A_pmgoKI551_0;
	wire w_dff_A_rM84gTKC2_0;
	wire w_dff_A_HrFf6mQx3_0;
	wire w_dff_A_YfYXewFo9_0;
	wire w_dff_A_r2MSjyaJ9_0;
	wire w_dff_A_jcBqriGy5_0;
	wire w_dff_A_jwfMJWPO3_0;
	wire w_dff_A_l0XUuEHd6_0;
	wire w_dff_A_TLmp5ND70_0;
	wire w_dff_A_CQbFnLfr6_0;
	wire w_dff_A_SKbKcetk1_0;
	wire w_dff_A_L6IqURT07_0;
	wire w_dff_A_1RlyPywy1_0;
	wire w_dff_A_YM7WnGRF9_0;
	wire w_dff_A_EIe6eaZE5_0;
	wire w_dff_A_lslajPSF1_0;
	wire w_dff_A_e8ZfvcSP1_0;
	wire w_dff_A_9SlHEK3L8_0;
	wire w_dff_A_CIp6Cpqx5_0;
	wire w_dff_A_c906w5Tr0_0;
	wire w_dff_A_KzHKDdGE1_0;
	wire w_dff_A_UBBuUfUc6_0;
	wire w_dff_A_6wW9gcSs6_0;
	wire w_dff_A_kJxTHZ8z4_0;
	wire w_dff_A_tsINoMcR6_1;
	wire w_dff_A_XIOyU0On8_0;
	wire w_dff_A_DKq3e43b4_0;
	wire w_dff_A_czLKlFlI1_0;
	wire w_dff_A_kneUDeSo9_0;
	wire w_dff_A_asRLFjFv8_0;
	wire w_dff_A_dmSL62r85_0;
	wire w_dff_A_WGYuRayh3_0;
	wire w_dff_A_t6Yo5nF36_0;
	wire w_dff_A_ff0bDvq20_0;
	wire w_dff_A_YprfJ5oT0_0;
	wire w_dff_A_joTFkHDa9_0;
	wire w_dff_A_e3zsG0NN4_0;
	wire w_dff_A_GiAcPx413_0;
	wire w_dff_A_dK4zzXzr1_0;
	wire w_dff_A_Ht2WsStZ1_0;
	wire w_dff_A_cQMboIm72_0;
	wire w_dff_A_8ON1Eriq9_0;
	wire w_dff_A_v8lLApdP1_0;
	wire w_dff_A_zuxOMWEg1_0;
	wire w_dff_A_XM4UcsAw0_0;
	wire w_dff_A_2hzFlrvq5_0;
	wire w_dff_A_MfntoeHo8_0;
	wire w_dff_A_sNo8GWjO7_0;
	wire w_dff_A_gQqToHrd4_0;
	wire w_dff_A_dmv0xlOx5_0;
	wire w_dff_A_Axk2z5rC2_0;
	wire w_dff_A_YnNXsQSi6_0;
	wire w_dff_A_HYgM8sFp3_0;
	wire w_dff_A_4jlBtAG66_0;
	wire w_dff_A_qu88kCpS4_0;
	wire w_dff_A_vZjIRnTp8_0;
	wire w_dff_A_YBpAlVzF8_0;
	wire w_dff_A_wUcfwBcW0_0;
	wire w_dff_A_97LBmKt26_0;
	wire w_dff_A_E8Kfagdu4_0;
	wire w_dff_A_qBosUjhi3_1;
	wire w_dff_A_XmgoDoCt4_0;
	wire w_dff_A_itObX5ox0_0;
	wire w_dff_A_Rpp4e2bC3_0;
	wire w_dff_A_lTkrdVcb8_0;
	wire w_dff_A_D5p6PecJ3_0;
	wire w_dff_A_JXSZ5SvE0_0;
	wire w_dff_A_3Z2f4XkW7_0;
	wire w_dff_A_A9OrukCD7_0;
	wire w_dff_A_NAYmCd8j7_0;
	wire w_dff_A_xupyWn3O3_0;
	wire w_dff_A_H4RuCvSp8_0;
	wire w_dff_A_zZ1EwvVA0_0;
	wire w_dff_A_czCWPgKP9_0;
	wire w_dff_A_xNdcvHzM6_0;
	wire w_dff_A_j87HSMIm3_0;
	wire w_dff_A_GmbMW3xD9_0;
	wire w_dff_A_C18XUQQa7_0;
	wire w_dff_A_naa32m2T6_0;
	wire w_dff_A_cOfx9NFv1_0;
	wire w_dff_A_4hpYc9fY4_0;
	wire w_dff_A_XsJpSv5p8_0;
	wire w_dff_A_fqUaLZyf4_0;
	wire w_dff_A_8RZ7vtGk9_0;
	wire w_dff_A_ODlXNWHL3_0;
	wire w_dff_A_4swP6WIa2_0;
	wire w_dff_A_d6Mo7nOM4_0;
	wire w_dff_A_KTfYlTgG4_0;
	wire w_dff_A_Zyw4Hh4c6_0;
	wire w_dff_A_n2kFEPZK1_0;
	wire w_dff_A_aJ1zcPEv6_0;
	wire w_dff_A_6irygS6R2_0;
	wire w_dff_A_bolcnoIS3_0;
	wire w_dff_A_uSEjDQWZ8_0;
	wire w_dff_A_KL8TYi5m6_0;
	wire w_dff_A_kQwDryEX1_0;
	wire w_dff_A_xbTcNRte5_0;
	wire w_dff_A_lAwUlNW61_0;
	wire w_dff_A_7CPkUKba1_1;
	wire w_dff_A_hFHRnq6W9_0;
	wire w_dff_A_cRkVY68A8_0;
	wire w_dff_A_IwjzF4j26_0;
	wire w_dff_A_JdS5G9fi0_0;
	wire w_dff_A_fOQ4OWmk6_0;
	wire w_dff_A_mLoOTjCq3_0;
	wire w_dff_A_HsuMZptG0_0;
	wire w_dff_A_ND3CZ08G8_0;
	wire w_dff_A_9BvbREtT2_0;
	wire w_dff_A_a4PKNzHV1_0;
	wire w_dff_A_5NBegsxh8_0;
	wire w_dff_A_dF4jaW3N3_0;
	wire w_dff_A_99JjSqbQ1_0;
	wire w_dff_A_p2BmPM2V6_0;
	wire w_dff_A_4ZozXwag7_0;
	wire w_dff_A_htkz3Bcv2_0;
	wire w_dff_A_btiXgu8q3_0;
	wire w_dff_A_FnFL6dh00_0;
	wire w_dff_A_afGZXWsr7_0;
	wire w_dff_A_v2n8Ng6n3_0;
	wire w_dff_A_d2BlWLgO1_0;
	wire w_dff_A_0Q0zobza8_0;
	wire w_dff_A_bgYQnZzi9_0;
	wire w_dff_A_5H3xuNUW5_0;
	wire w_dff_A_S7AHO3mo4_0;
	wire w_dff_A_jtWoDO2h5_0;
	wire w_dff_A_gBOFoBxy4_0;
	wire w_dff_A_RhFHycWi4_0;
	wire w_dff_A_DT78MEPQ2_0;
	wire w_dff_A_Oc6JN0xg0_0;
	wire w_dff_A_HdxBD7nt4_0;
	wire w_dff_A_bInwR5Tk5_0;
	wire w_dff_A_JFFF6dnL9_0;
	wire w_dff_A_xooZ55Ga8_0;
	wire w_dff_A_A4jbgDlv0_0;
	wire w_dff_A_GgnUw7223_0;
	wire w_dff_A_DK5nqAm15_0;
	wire w_dff_A_ssThCr5Y4_2;
	wire w_dff_A_M4P5kbJ74_0;
	wire w_dff_A_jl8WAa2z7_0;
	wire w_dff_A_5NHkHYdl1_0;
	wire w_dff_A_p1QNopHh9_0;
	wire w_dff_A_CKsYa0bN9_0;
	wire w_dff_A_fUcmldH32_0;
	wire w_dff_A_YXJAhgpv8_0;
	wire w_dff_A_bw2fKbEw5_0;
	wire w_dff_A_FJJLuoSa8_0;
	wire w_dff_A_o7Hz3tdQ5_0;
	wire w_dff_A_kzHlWNOg3_0;
	wire w_dff_A_PUqeC5lp1_0;
	wire w_dff_A_P07lZhrt0_0;
	wire w_dff_A_totwC3zQ5_0;
	wire w_dff_A_cMqDTa7Z0_0;
	wire w_dff_A_iBdouH5S5_0;
	wire w_dff_A_3VKFQcpz6_0;
	wire w_dff_A_T9P5G9uA4_0;
	wire w_dff_A_5rr3c4HZ8_0;
	wire w_dff_A_d8ncZiCq3_0;
	wire w_dff_A_KYIgKngs5_0;
	wire w_dff_A_qTx1po8g7_0;
	wire w_dff_A_0tW622NM2_0;
	wire w_dff_A_sdiKqK4P3_0;
	wire w_dff_A_gzziJXjC0_0;
	wire w_dff_A_USJhQbOg3_0;
	wire w_dff_A_LBF6doIT2_0;
	wire w_dff_A_fBpDS66K8_0;
	wire w_dff_A_icL07ajY8_0;
	wire w_dff_A_SS5zIw232_0;
	wire w_dff_A_qCEiOyxe6_0;
	wire w_dff_A_S4fqUD1W6_0;
	wire w_dff_A_VMd4BWbO7_0;
	wire w_dff_A_72TtIEga5_0;
	wire w_dff_A_GRCmtOQz2_0;
	wire w_dff_A_bM2a9uym8_0;
	wire w_dff_A_2CM4RefF3_1;
	wire w_dff_A_n5yoZDCf8_0;
	wire w_dff_A_bKF5IE3v5_0;
	wire w_dff_A_4zRKyYlP0_0;
	wire w_dff_A_VWD6FnwO0_0;
	wire w_dff_A_c7AkPyDO7_0;
	wire w_dff_A_NU8Yegop7_0;
	wire w_dff_A_FjyWPSxX2_0;
	wire w_dff_A_qX7D6fDA9_0;
	wire w_dff_A_jiIR7V6H0_0;
	wire w_dff_A_u69AqvrK0_0;
	wire w_dff_A_TSC8EBos4_0;
	wire w_dff_A_TMTyYm9x4_0;
	wire w_dff_A_iVmQubmu0_0;
	wire w_dff_A_4kYU3pSG2_0;
	wire w_dff_A_TOO6hyuv1_0;
	wire w_dff_A_pqZdBcaF9_0;
	wire w_dff_A_Fbjf0KqF1_0;
	wire w_dff_A_dB48OhgZ7_0;
	wire w_dff_A_zCkggYEu9_0;
	wire w_dff_A_XrWLbXV64_0;
	wire w_dff_A_nDeGW0gs1_0;
	wire w_dff_A_AWxxHpcb5_0;
	wire w_dff_A_KMlUbPeh0_0;
	wire w_dff_A_uLqjC8R84_0;
	wire w_dff_A_Wiwszthh8_0;
	wire w_dff_A_GQtNPTjH2_0;
	wire w_dff_A_ul6SvONu8_0;
	wire w_dff_A_3C3pdOhQ0_0;
	wire w_dff_A_gwXh8D4n5_0;
	wire w_dff_A_CwSzkxRm1_0;
	wire w_dff_A_N1pluRYG2_0;
	wire w_dff_A_Xa6DPwYr3_0;
	wire w_dff_A_GU7r6nvd5_0;
	wire w_dff_A_mrVNT3gD6_0;
	wire w_dff_A_coFlINwc6_0;
	wire w_dff_A_2i4GnoHT7_0;
	wire w_dff_A_GEUJn6gc6_0;
	wire w_dff_A_ZwTqURVo7_2;
	wire w_dff_A_plbNHkHT8_0;
	wire w_dff_A_62v67yL61_0;
	wire w_dff_A_lzLj9gwB7_0;
	wire w_dff_A_AMqU5Q7T1_0;
	wire w_dff_A_rKxjZvUk8_0;
	wire w_dff_A_IokWATAQ4_0;
	wire w_dff_A_BgZ99lLa4_0;
	wire w_dff_A_pJnvJxP37_0;
	wire w_dff_A_yxQp2DIN4_0;
	wire w_dff_A_ocwSjP7n9_0;
	wire w_dff_A_tgOR6fJn0_0;
	wire w_dff_A_h4ApIzZf9_0;
	wire w_dff_A_EKQhDHtQ6_0;
	wire w_dff_A_rTmEYGpL2_0;
	wire w_dff_A_Oh1EcsKi0_0;
	wire w_dff_A_QbVMJAyt6_0;
	wire w_dff_A_x38VK13U7_0;
	wire w_dff_A_Lf3y1ZlA5_0;
	wire w_dff_A_pkU8CXXw0_0;
	wire w_dff_A_yUQyUETs8_0;
	wire w_dff_A_kq3u3yqe7_0;
	wire w_dff_A_v9ZiQGw37_0;
	wire w_dff_A_4ryWWJ1Q2_0;
	wire w_dff_A_wzbqZFOy7_0;
	wire w_dff_A_j1ezqyNl7_0;
	wire w_dff_A_blHQsdka1_0;
	wire w_dff_A_5eU4ibM80_0;
	wire w_dff_A_AHgRfG8G2_0;
	wire w_dff_A_frXSsZH08_0;
	wire w_dff_A_0vJJS7Pc9_0;
	wire w_dff_A_EqH1qAAp1_0;
	wire w_dff_A_uUWmgIk26_0;
	wire w_dff_A_Xwr63UvT2_0;
	wire w_dff_A_aNtfbfzQ8_0;
	wire w_dff_A_n5p0vNWm1_0;
	wire w_dff_A_16veWjrJ2_0;
	wire w_dff_A_x6bwFvue0_2;
	wire w_dff_A_vJTDuolT8_0;
	wire w_dff_A_mVRE5PBb3_0;
	wire w_dff_A_j4HHhwUy1_0;
	wire w_dff_A_8ymnaPga4_0;
	wire w_dff_A_gMawEEuw6_0;
	wire w_dff_A_kkOSS41X7_0;
	wire w_dff_A_FokBI5dd4_0;
	wire w_dff_A_eKfA5OVK9_0;
	wire w_dff_A_oLhL8F5V8_0;
	wire w_dff_A_xm5UzF4w4_0;
	wire w_dff_A_xirkfDEl9_0;
	wire w_dff_A_VSyMBy6L9_0;
	wire w_dff_A_hwPy5vzu4_0;
	wire w_dff_A_bVZYnrVS2_0;
	wire w_dff_A_qKLwvFUP1_0;
	wire w_dff_A_PWdW3zAt4_0;
	wire w_dff_A_xPZrV0SC3_0;
	wire w_dff_A_fJaFXqRS8_0;
	wire w_dff_A_TPgnHYr46_0;
	wire w_dff_A_xAKLmj6O5_0;
	wire w_dff_A_QWWWZ0AH4_0;
	wire w_dff_A_s6o5VFmK0_0;
	wire w_dff_A_gXKFYeAi4_0;
	wire w_dff_A_KfUohfH77_0;
	wire w_dff_A_IxFXTg752_0;
	wire w_dff_A_fjgkxzkq0_0;
	wire w_dff_A_cR61TyC04_0;
	wire w_dff_A_lJS3UL8m0_0;
	wire w_dff_A_jzmgkfkQ5_0;
	wire w_dff_A_T7UAfG1r1_0;
	wire w_dff_A_PVcoIPhT0_0;
	wire w_dff_A_of390Vzo3_0;
	wire w_dff_A_GDUSIUm76_0;
	wire w_dff_A_hYnJaZzd3_0;
	wire w_dff_A_3SV0BPMb8_0;
	wire w_dff_A_0w6Csyvn8_1;
	wire w_dff_A_aJRzz02e8_0;
	wire w_dff_A_ySSvZSMX1_0;
	wire w_dff_A_817qS1Yx7_0;
	wire w_dff_A_vwTRdGvn7_0;
	wire w_dff_A_NmgrfalF8_0;
	wire w_dff_A_DMZsHzAL7_0;
	wire w_dff_A_wcMw7NWP6_0;
	wire w_dff_A_3gaDqzmV2_0;
	wire w_dff_A_WOxNUutk7_0;
	wire w_dff_A_Tpyuw7Lb4_0;
	wire w_dff_A_vGyNWZlW9_0;
	wire w_dff_A_vY89ozsT9_0;
	wire w_dff_A_W92VnVZr5_0;
	wire w_dff_A_1S4h1ec35_0;
	wire w_dff_A_nQYf6h6r3_0;
	wire w_dff_A_XFgQYpmq3_0;
	wire w_dff_A_dTAP4cXN1_0;
	wire w_dff_A_vCjQO0hF3_0;
	wire w_dff_A_32bftMGQ8_0;
	wire w_dff_A_T4hKSIS77_0;
	wire w_dff_A_REX2j62H4_0;
	wire w_dff_A_Gq3lznHz2_0;
	wire w_dff_A_QhEIEVDd9_0;
	wire w_dff_A_bHzDProK3_0;
	wire w_dff_A_ykyFEO5f6_0;
	wire w_dff_A_lNTfgc6s7_0;
	wire w_dff_A_oOdCMo2h3_0;
	wire w_dff_A_ZESI0Ss79_0;
	wire w_dff_A_EWfjLcQY6_0;
	wire w_dff_A_qmZVpdSi9_0;
	wire w_dff_A_2vQLWaaH3_0;
	wire w_dff_A_03PM1Ut50_0;
	wire w_dff_A_UhMHdjPL6_0;
	wire w_dff_A_uz1hkg592_0;
	wire w_dff_A_cCEHWIOR6_0;
	wire w_dff_A_9Pj9fEaC9_0;
	wire w_dff_A_vT7Mf1cx5_0;
	wire w_dff_A_UKxWtnJd8_2;
	wire w_dff_A_RuP9411f3_0;
	wire w_dff_A_ALhJE6hN7_0;
	wire w_dff_A_GbNS7SoF3_0;
	wire w_dff_A_cn5ShnvJ9_0;
	wire w_dff_A_qwTw1RaX2_0;
	wire w_dff_A_PNs8KCUb1_0;
	wire w_dff_A_93QzkCA82_0;
	wire w_dff_A_xglkL6wa8_0;
	wire w_dff_A_LXbpOo1Z0_0;
	wire w_dff_A_Xvh2uMQd3_0;
	wire w_dff_A_LRBna6GA3_0;
	wire w_dff_A_AESoj9m69_0;
	wire w_dff_A_SXECSwnZ7_0;
	wire w_dff_A_DKCrPw4f9_0;
	wire w_dff_A_eXmqM5jx6_0;
	wire w_dff_A_w4oSo3Yn8_0;
	wire w_dff_A_91V8v4Y38_0;
	wire w_dff_A_nULIvwbz1_0;
	wire w_dff_A_2c8d4vxf3_0;
	wire w_dff_A_rND2kL1W5_0;
	wire w_dff_A_vZpAs4mw8_0;
	wire w_dff_A_BZ0hxsoU0_0;
	wire w_dff_A_BDOGNpk46_0;
	wire w_dff_A_TZznJtTl5_0;
	wire w_dff_A_ZYFuPgoN6_0;
	wire w_dff_A_c1vNB3sB2_0;
	wire w_dff_A_tmxk6DYN5_0;
	wire w_dff_A_Flz6wzH57_0;
	wire w_dff_A_WzZOrcEQ3_0;
	wire w_dff_A_Pd7S7EJy4_0;
	wire w_dff_A_fVJNAEaJ9_0;
	wire w_dff_A_j7TRNiBv1_0;
	wire w_dff_A_jWybCdhP2_0;
	wire w_dff_A_RWyN0RFi0_0;
	wire w_dff_A_jQgGwhbs3_0;
	wire w_dff_A_M0HT7wKV8_1;
	wire w_dff_A_XEH1iaR35_0;
	wire w_dff_A_CqiTVAVZ2_0;
	wire w_dff_A_bsfuE8Sl1_0;
	wire w_dff_A_zWxyzn3l5_0;
	wire w_dff_A_WzuUtemE3_0;
	wire w_dff_A_paBSIU5t2_0;
	wire w_dff_A_nu7sBOC97_0;
	wire w_dff_A_HzvtWlB31_0;
	wire w_dff_A_kuGB9u1T4_0;
	wire w_dff_A_q0C6jZsZ7_0;
	wire w_dff_A_ATNOlEmw6_0;
	wire w_dff_A_l78yR6Lg3_0;
	wire w_dff_A_WeboNXlf9_0;
	wire w_dff_A_6Xgt1Nuk4_0;
	wire w_dff_A_BxZix9QQ3_0;
	wire w_dff_A_FwZWJJCL2_0;
	wire w_dff_A_lID18ov26_0;
	wire w_dff_A_AjzjY1pl6_0;
	wire w_dff_A_oNu8Qi0D7_0;
	wire w_dff_A_aZE4mLlt9_0;
	wire w_dff_A_bZMU7YKQ7_0;
	wire w_dff_A_RR9XyXBC3_0;
	wire w_dff_A_wrF4K1iO4_0;
	wire w_dff_A_x9NQhUqe8_0;
	wire w_dff_A_gOZDgZ043_0;
	wire w_dff_A_ZjsyHjk21_0;
	wire w_dff_A_S0Qy6RCn4_0;
	wire w_dff_A_d9rpGd3U9_0;
	wire w_dff_A_BUfKz0sK4_0;
	wire w_dff_A_xK4mRano6_0;
	wire w_dff_A_2RJVWX3P4_0;
	wire w_dff_A_KniBZR9T5_0;
	wire w_dff_A_sAHh03771_0;
	wire w_dff_A_iQckNP664_0;
	wire w_dff_A_v3a1Duhj4_0;
	wire w_dff_A_KWBqBybj2_0;
	wire w_dff_A_vcCgEMvk3_0;
	wire w_dff_A_EbglPHaX6_2;
	wire w_dff_A_swV84blL3_0;
	wire w_dff_A_MoTpyETq4_0;
	wire w_dff_A_befxaSdt5_0;
	wire w_dff_A_nj1S3wB41_0;
	wire w_dff_A_7C4MqCvJ4_0;
	wire w_dff_A_NJpT3PZq6_0;
	wire w_dff_A_rUUp3FX02_0;
	wire w_dff_A_fSutrgXe6_0;
	wire w_dff_A_VgcIlFzG8_0;
	wire w_dff_A_69izWaog9_0;
	wire w_dff_A_Cdzp4wZp7_0;
	wire w_dff_A_virqKLAN5_0;
	wire w_dff_A_5ENM3xos9_0;
	wire w_dff_A_V2tqs1vF0_0;
	wire w_dff_A_wk30Ygv81_0;
	wire w_dff_A_110pMlfj1_0;
	wire w_dff_A_hWdkipOI8_0;
	wire w_dff_A_GQm3qUCT1_0;
	wire w_dff_A_iIUXtAtb7_0;
	wire w_dff_A_ZsJAKTfe5_0;
	wire w_dff_A_qXeYCbkh8_0;
	wire w_dff_A_RFNpAnF93_0;
	wire w_dff_A_EjXHQbSF4_0;
	wire w_dff_A_40eeJVPZ1_0;
	wire w_dff_A_5QtKENZk9_0;
	wire w_dff_A_wkcGo9BV7_0;
	wire w_dff_A_Oit6hlsp3_0;
	wire w_dff_A_RmnDTltQ2_0;
	wire w_dff_A_EtNNyMz02_0;
	wire w_dff_A_rIrObztX0_0;
	wire w_dff_A_9dE3pU650_0;
	wire w_dff_A_6L9Z9La10_0;
	wire w_dff_A_rfwuTdbL8_0;
	wire w_dff_A_XcD2rOzf0_0;
	wire w_dff_A_siWTAYaz3_0;
	wire w_dff_A_POP02OC74_0;
	wire w_dff_A_rz4eBgoh6_0;
	wire w_dff_A_S8QuRzkE0_2;
	wire w_dff_A_dseyb2v74_0;
	wire w_dff_A_OUFirTFu9_0;
	wire w_dff_A_0TFd1sSJ4_0;
	wire w_dff_A_kXRCpNYU6_0;
	wire w_dff_A_YUdKZbFq6_0;
	wire w_dff_A_W5OsBaa58_0;
	wire w_dff_A_uu9vKEwQ8_0;
	wire w_dff_A_FMlwMk116_0;
	wire w_dff_A_XAK0UxfS4_0;
	wire w_dff_A_fvgllW6Q1_0;
	wire w_dff_A_XCi5mrWq6_0;
	wire w_dff_A_vMeoGz8n2_0;
	wire w_dff_A_0Bdpm1em9_0;
	wire w_dff_A_3nVUNd1z4_0;
	wire w_dff_A_q6yS1vd01_0;
	wire w_dff_A_VeUuPMa17_0;
	wire w_dff_A_XNT9SGAd2_0;
	wire w_dff_A_x7xCGkqj3_0;
	wire w_dff_A_T0wCi8o12_0;
	wire w_dff_A_Cely64dP6_0;
	wire w_dff_A_nrExZfeL0_0;
	wire w_dff_A_rQYLfaUN2_0;
	wire w_dff_A_12TaG0F05_0;
	wire w_dff_A_5a9NCTDT6_0;
	wire w_dff_A_aFXjbadQ2_0;
	wire w_dff_A_BBfr5o794_0;
	wire w_dff_A_B5YKQYA75_0;
	wire w_dff_A_tHYkYDFq7_0;
	wire w_dff_A_OxPfMyx55_0;
	wire w_dff_A_MvRVSvZU6_0;
	wire w_dff_A_T99Xbd8v0_0;
	wire w_dff_A_0ioXxkSG6_0;
	wire w_dff_A_C7Y9DVay5_2;
	wire w_dff_A_nzl4gXeX9_0;
	wire w_dff_A_H3VhH1vY2_0;
	wire w_dff_A_JZLqlW553_0;
	wire w_dff_A_kfVPIFvh6_0;
	wire w_dff_A_xZOhCyG66_0;
	wire w_dff_A_enRZMrRj2_0;
	wire w_dff_A_5ULdjhRT0_0;
	wire w_dff_A_ViaN4srH4_0;
	wire w_dff_A_9D32lsUc0_0;
	wire w_dff_A_xeF3ArdW7_0;
	wire w_dff_A_6veNz4KY3_2;
	wire w_dff_A_9HZvrbM50_0;
	wire w_dff_A_Iofqhzvn3_0;
	wire w_dff_A_Rpdsh7GX8_0;
	wire w_dff_A_ShHN4Y151_0;
	wire w_dff_A_KT01SSCm0_0;
	wire w_dff_A_jUpYjNDe8_0;
	wire w_dff_A_koFrxztT6_0;
	wire w_dff_A_Q3yJPoNu6_0;
	wire w_dff_A_jfYRn6PI6_0;
	wire w_dff_A_pJJ0Ihlt6_0;
	wire w_dff_A_oa0XxNvS3_2;
	wire w_dff_A_bB4avgpf0_0;
	wire w_dff_A_Nt3WlxA69_0;
	wire w_dff_A_IzCSaNRG4_0;
	wire w_dff_A_VqUfarth3_0;
	wire w_dff_A_CP0LNn3C8_0;
	wire w_dff_A_wBzVYZfD6_0;
	wire w_dff_A_Wko3XSpy7_0;
	wire w_dff_A_M0lcvcBX0_0;
	wire w_dff_A_yFOsYNUg9_0;
	wire w_dff_A_NED2kRvc1_0;
	wire w_dff_A_Y3lDAcRw4_0;
	wire w_dff_A_jOZt3TJ25_0;
	wire w_dff_A_JERUK1X57_0;
	wire w_dff_A_Ngvebk253_0;
	wire w_dff_A_w1ntX4QK4_0;
	wire w_dff_A_AYdDzrQq9_0;
	wire w_dff_A_hToYVN4Y9_0;
	wire w_dff_A_mcyC9mh01_0;
	wire w_dff_A_KuuqqpVz0_0;
	wire w_dff_A_cBOkQEx37_0;
	wire w_dff_A_NXSWMPmp2_0;
	wire w_dff_A_ftUV2bVH7_0;
	wire w_dff_A_sdKYZNvW4_0;
	wire w_dff_A_Ij8AChXO0_0;
	wire w_dff_A_NyvscHrC9_2;
	wire w_dff_A_x8uJ3uU14_0;
	wire w_dff_A_uWUq719U4_0;
	wire w_dff_A_Ra96J6TQ9_0;
	wire w_dff_A_oYmIiRKo1_0;
	wire w_dff_A_Ag0jBzgQ0_0;
	wire w_dff_A_6y2qeYlc9_0;
	wire w_dff_A_63ytucfX7_0;
	wire w_dff_A_DV8plbpk4_0;
	wire w_dff_A_D56M6mj31_0;
	wire w_dff_A_7vvA95Gx0_0;
	wire w_dff_A_7Pro7rEs1_0;
	wire w_dff_A_I7WGF6fh4_0;
	wire w_dff_A_QpadcRY80_0;
	wire w_dff_A_l7Pn9xLV6_0;
	wire w_dff_A_sdWqi4Go1_0;
	wire w_dff_A_oz2mxFWJ6_0;
	wire w_dff_A_UDnVxWWn3_0;
	wire w_dff_A_AldomAwp8_0;
	wire w_dff_A_8gjEDqU79_0;
	wire w_dff_A_F6GX7V5k7_0;
	wire w_dff_A_ylmtbOf76_0;
	wire w_dff_A_rXriJFTA6_0;
	wire w_dff_A_I33HmPdM2_0;
	wire w_dff_A_fjmmPZfX7_0;
	wire w_dff_A_rPh0qnnX6_0;
	wire w_dff_A_MLSieQRb5_0;
	wire w_dff_A_lPzfP2la9_2;
	wire w_dff_A_VEC37Kb97_0;
	wire w_dff_A_yKwTG61T1_0;
	wire w_dff_A_U29S5hfu4_0;
	wire w_dff_A_v6cvdGue5_0;
	wire w_dff_A_PgLsNzlD8_0;
	wire w_dff_A_IwHeJo6u7_0;
	wire w_dff_A_eepxyCLY5_0;
	wire w_dff_A_KoOHLsFp7_0;
	wire w_dff_A_GeuJQvZH1_0;
	wire w_dff_A_w9WqPI5b7_0;
	wire w_dff_A_h6KY3otM4_0;
	wire w_dff_A_pQXfIaEc7_0;
	wire w_dff_A_OGfNbo279_0;
	wire w_dff_A_OPysQK8j9_0;
	wire w_dff_A_YKfG7xbx4_0;
	wire w_dff_A_046HKjwD5_0;
	wire w_dff_A_nyu2S2zC0_0;
	wire w_dff_A_8ePTkFr49_0;
	wire w_dff_A_Efgp4oSm6_0;
	wire w_dff_A_6fJC1h071_0;
	wire w_dff_A_948eRYST5_0;
	wire w_dff_A_0Ee2ZB4q3_0;
	wire w_dff_A_s3R6TkFj3_0;
	wire w_dff_A_zKOEIkDr2_0;
	wire w_dff_A_2z1wE9Tr7_0;
	wire w_dff_A_CreCEGnX4_0;
	wire w_dff_A_ZVuNEt8t7_0;
	wire w_dff_A_IQkVbZHN5_0;
	wire w_dff_A_tL4B5Qt22_0;
	wire w_dff_A_JmJfu1Jx3_2;
	wire w_dff_A_prcnguFT9_0;
	wire w_dff_A_XKV3xiQI6_0;
	wire w_dff_A_sfGrFQKw2_0;
	wire w_dff_A_1TmbwBDk6_0;
	wire w_dff_A_GlJUvyaM9_0;
	wire w_dff_A_4vpgJdKb8_0;
	wire w_dff_A_E6RaSHGq9_0;
	wire w_dff_A_Z5vwzN8A5_0;
	wire w_dff_A_HaUUTyqT3_0;
	wire w_dff_A_Oqd4VR4j8_0;
	wire w_dff_A_XrCT66DO4_0;
	wire w_dff_A_fD6h7s5w5_0;
	wire w_dff_A_sBgo36vb4_0;
	wire w_dff_A_P6AVwomB9_0;
	wire w_dff_A_LGhfym0w3_0;
	wire w_dff_A_ismxpB1d4_0;
	wire w_dff_A_Qa4lUHWV6_0;
	wire w_dff_A_P5bnf5xA4_0;
	wire w_dff_A_TLWD8j7q8_0;
	wire w_dff_A_PmPFXRkm5_0;
	wire w_dff_A_1DEqSVSh8_0;
	wire w_dff_A_hvLRLS7Y4_0;
	wire w_dff_A_hBdyxDej5_0;
	wire w_dff_A_uVOIUjPU9_0;
	wire w_dff_A_LcmR00Rp7_0;
	wire w_dff_A_RLqxLHBO8_0;
	wire w_dff_A_nTjrgZKe8_0;
	wire w_dff_A_FFcBnvFW4_0;
	wire w_dff_A_TQEAN2BS3_0;
	wire w_dff_A_yAlJLw6x9_0;
	wire w_dff_A_SGZG573Y4_2;
	wire w_dff_A_9mPUOZh00_0;
	wire w_dff_A_Jnwu2Yhf4_0;
	wire w_dff_A_joi2S2HD0_0;
	wire w_dff_A_Jr2FxMJX9_0;
	wire w_dff_A_qzv6Kkxg3_0;
	wire w_dff_A_rov2lSPR2_0;
	wire w_dff_A_QmAp1mWZ8_0;
	wire w_dff_A_QZwkynxl6_0;
	wire w_dff_A_Iu7M7jYm4_0;
	wire w_dff_A_pOGcSKCK9_0;
	wire w_dff_A_mYyUNWY12_0;
	wire w_dff_A_dSTkFMBC4_0;
	wire w_dff_A_fJTZhBr26_0;
	wire w_dff_A_5JsqUKxw8_0;
	wire w_dff_A_3Rh7J9tu3_0;
	wire w_dff_A_bnz3u5M11_0;
	wire w_dff_A_xMdH4bvC6_0;
	wire w_dff_A_w14rmFCR8_0;
	wire w_dff_A_YIe0BZdp2_0;
	wire w_dff_A_1iQksQaM0_2;
	wire w_dff_A_hJfgijJH7_0;
	wire w_dff_A_ENMl7Ul43_0;
	wire w_dff_A_DExDC5NA7_0;
	wire w_dff_A_lvtQbmGm9_0;
	wire w_dff_A_Dn1W2jZo5_0;
	wire w_dff_A_oRVU4bwl0_0;
	wire w_dff_A_3EwZXQr04_0;
	wire w_dff_A_AdfZZQkV9_0;
	wire w_dff_A_cPHzPg2Q5_0;
	wire w_dff_A_Utf0xcYh7_0;
	wire w_dff_A_g5xImQhC7_0;
	wire w_dff_A_ASQRqqgS8_0;
	wire w_dff_A_npwC4EFi4_0;
	wire w_dff_A_TttgXi3p2_0;
	wire w_dff_A_xz1zoii98_0;
	wire w_dff_A_QZu0Vnbb5_0;
	wire w_dff_A_cuTUdWVQ7_0;
	wire w_dff_A_DmhPxgal5_0;
	wire w_dff_A_TU3bReNd5_0;
	wire w_dff_A_CtZh37QI7_0;
	wire w_dff_A_Pvsn6F9o5_0;
	wire w_dff_A_8hS9m2Y73_2;
	wire w_dff_A_81labtvY2_0;
	wire w_dff_A_akV4xtHz7_0;
	wire w_dff_A_nIGbZKFp1_0;
	wire w_dff_A_lUNlwOxw3_0;
	wire w_dff_A_gSSZ0jMX7_0;
	wire w_dff_A_rcRwI3k86_0;
	wire w_dff_A_4noCiurx9_0;
	wire w_dff_A_k94ta9Te0_0;
	wire w_dff_A_9ipDSy589_0;
	wire w_dff_A_uEyHgZvI9_0;
	wire w_dff_A_PSRTnObD1_0;
	wire w_dff_A_mvSPDdfY6_0;
	wire w_dff_A_QN6sim7e1_0;
	wire w_dff_A_JP63ReqE8_0;
	wire w_dff_A_y2sS8QCS1_0;
	wire w_dff_A_a5EPy4Eo6_0;
	wire w_dff_A_5o1x4bdg3_0;
	wire w_dff_A_3ICkKOD14_0;
	wire w_dff_A_C1hkKMUJ3_0;
	wire w_dff_A_JZvHAGLw5_0;
	wire w_dff_A_fyaugnMa2_0;
	wire w_dff_A_QdpmjzBx0_2;
	wire w_dff_A_iZEIChW01_0;
	wire w_dff_A_mn0c5MFP5_0;
	wire w_dff_A_Dj3tBW0L8_0;
	wire w_dff_A_7kaOGsd84_0;
	wire w_dff_A_0cWbSjBm6_0;
	wire w_dff_A_MIY5zbxi1_0;
	wire w_dff_A_wTQvmoWW0_0;
	wire w_dff_A_GAteg4uW2_0;
	wire w_dff_A_xVQkVIfh8_0;
	wire w_dff_A_HGnJh86x2_0;
	wire w_dff_A_OJvHaqSg2_0;
	wire w_dff_A_vxK1JuXe5_0;
	wire w_dff_A_lI7zYVwi0_0;
	wire w_dff_A_qgijVHmm8_0;
	wire w_dff_A_bQjDTPrO9_0;
	wire w_dff_A_vHHhn0rE8_0;
	wire w_dff_A_moKsCxe35_0;
	wire w_dff_A_fbVCFjhV8_0;
	wire w_dff_A_yxYhDQmB1_0;
	wire w_dff_A_VEG1LvX42_0;
	wire w_dff_A_DH8muabI7_0;
	wire w_dff_A_lvIBfCit0_0;
	wire w_dff_A_i6ELr4Gm8_0;
	wire w_dff_A_bjP8Gnko9_1;
	wire w_dff_A_JygE6xV54_0;
	wire w_dff_A_H4LIQZcz0_0;
	wire w_dff_A_9BdYvwWZ5_0;
	wire w_dff_A_xjFsUMIC1_0;
	wire w_dff_A_nBEVTmQl0_0;
	wire w_dff_A_ZTRW8m1r2_0;
	wire w_dff_A_vY0xZFyl9_0;
	wire w_dff_A_Mt9v6H714_0;
	wire w_dff_A_0YXCL5Ik2_0;
	wire w_dff_A_CBiBBm4n5_0;
	wire w_dff_A_iBsDKZqG6_0;
	wire w_dff_A_7WFgkYER7_0;
	wire w_dff_A_FsukPbtM5_0;
	wire w_dff_A_GugBEpix2_0;
	wire w_dff_A_V0skxr0F7_0;
	wire w_dff_A_XfMIXKrl8_0;
	wire w_dff_A_Ll27CUwy3_0;
	wire w_dff_A_NzGWomL06_0;
	wire w_dff_A_UUfhRLOj5_0;
	wire w_dff_A_o6KxQzLL7_0;
	wire w_dff_A_GfGoUerw9_0;
	wire w_dff_A_r2wZF0K61_0;
	wire w_dff_A_H9WEcLuX7_0;
	wire w_dff_A_cplgJl6L5_0;
	wire w_dff_A_kgzbzXtT2_0;
	wire w_dff_A_KY6aIAwW6_0;
	wire w_dff_A_vfpGiafr1_0;
	wire w_dff_A_I8w0B8AP8_1;
	wire w_dff_A_lvMnoDQb4_0;
	wire w_dff_A_quCktKZK7_0;
	wire w_dff_A_X2cIBIdp3_0;
	wire w_dff_A_t4blgWWg3_0;
	wire w_dff_A_Of6vaUcI3_0;
	wire w_dff_A_WCLfFFzk4_0;
	wire w_dff_A_hEk6ocyy6_0;
	wire w_dff_A_WBawVD2a9_0;
	wire w_dff_A_VycTajte5_0;
	wire w_dff_A_YhKGf7wL9_0;
	wire w_dff_A_Kz6Ru4PS6_0;
	wire w_dff_A_L0UlO98V6_0;
	wire w_dff_A_gR1jdJvZ9_0;
	wire w_dff_A_nExZUtR06_0;
	wire w_dff_A_5BU2K0yv5_0;
	wire w_dff_A_hT4K5FmC9_0;
	wire w_dff_A_5LoUhNRd9_0;
	wire w_dff_A_h0ewkhsh3_0;
	wire w_dff_A_btY6XhyT9_0;
	wire w_dff_A_A5zHOWMX2_0;
	wire w_dff_A_E7nqzzLD2_0;
	wire w_dff_A_aYNRGjsY9_0;
	wire w_dff_A_2uwE9oa72_0;
	wire w_dff_A_52KrNaZP3_0;
	wire w_dff_A_Udi0OLKP8_0;
	wire w_dff_A_pC563uJb1_0;
	wire w_dff_A_3jAjF1Gz6_0;
	wire w_dff_A_wwd0LvTI7_0;
	wire w_dff_A_fl9wfYSL3_0;
	wire w_dff_A_qkkR41lL2_1;
	wire w_dff_A_7ljZlT9V9_0;
	wire w_dff_A_shnOCCR11_0;
	wire w_dff_A_czG8FT767_0;
	wire w_dff_A_al6xBKIX6_0;
	wire w_dff_A_R7QPpjgf2_0;
	wire w_dff_A_pPRppIca7_0;
	wire w_dff_A_zO4s8VNy2_0;
	wire w_dff_A_NTX6bz143_0;
	wire w_dff_A_GhGmbBTX1_0;
	wire w_dff_A_uhyNS0uH7_0;
	wire w_dff_A_MKOz98611_0;
	wire w_dff_A_2LBlAj0V3_0;
	wire w_dff_A_S74WIrSZ4_0;
	wire w_dff_A_qBBnIvzr8_0;
	wire w_dff_A_6AmY8qAZ4_0;
	wire w_dff_A_Sr5tra2P7_0;
	wire w_dff_A_slxDaHWE6_0;
	wire w_dff_A_386anNwP6_0;
	wire w_dff_A_u4bbuj2R2_0;
	wire w_dff_A_BG3MG6e71_0;
	wire w_dff_A_XtDUCDlA7_0;
	wire w_dff_A_1P1c9G1b8_0;
	wire w_dff_A_M23WeA3w0_0;
	wire w_dff_A_y5ZnVpJd4_0;
	wire w_dff_A_kBitKUpS4_0;
	wire w_dff_A_mG0QgLiw8_0;
	wire w_dff_A_IMH9stej5_0;
	wire w_dff_A_ku4bgICf8_0;
	wire w_dff_A_ILSvZBEJ4_2;
	wire w_dff_A_OVLSzOC91_0;
	wire w_dff_A_ZyDKHbNT6_0;
	wire w_dff_A_01A7bkPs6_0;
	wire w_dff_A_SdsYbdir9_0;
	wire w_dff_A_yUIXDO435_0;
	wire w_dff_A_SFTo6Cfo7_0;
	wire w_dff_A_QK4jZoz99_0;
	wire w_dff_A_2krjyInS3_0;
	wire w_dff_A_P125zpNw4_0;
	wire w_dff_A_ediNWG1J7_0;
	wire w_dff_A_xfiKRwPP3_2;
	wire w_dff_A_aK0GLROY2_0;
	wire w_dff_A_36wbyAAn1_0;
	wire w_dff_A_i6rV34jg1_0;
	wire w_dff_A_vfccntIk7_0;
	wire w_dff_A_NZNHqxuW7_0;
	wire w_dff_A_fycggT6y2_0;
	wire w_dff_A_4o1FDuoc5_0;
	wire w_dff_A_FjvKrP1L7_0;
	wire w_dff_A_led1xBmg1_0;
	wire w_dff_A_X39QseWh6_0;
	wire w_dff_A_zrcXL1rl7_2;
	wire w_dff_A_V6rEcdFt9_0;
	wire w_dff_A_YVfZ5NnC0_0;
	wire w_dff_A_742KAgvO1_0;
	wire w_dff_A_qDtSjULd9_1;
	wire w_dff_A_ugdaHuIq3_0;
	wire w_dff_A_KsYWvMPz2_0;
	wire w_dff_A_pzKquxwd5_0;
	wire w_dff_A_xPDRx4bs8_0;
	wire w_dff_A_1XTG5deb9_0;
	wire w_dff_A_uDtlWOCu5_0;
	wire w_dff_A_VLrYmf5Z1_0;
	wire w_dff_A_spldhYxi7_0;
	wire w_dff_A_KhQG3VGM0_0;
	wire w_dff_A_n5Qvx2W22_0;
	wire w_dff_A_8S4rUr0x5_0;
	wire w_dff_A_PYLW6zl73_0;
	wire w_dff_A_mGLUpW3V3_0;
	wire w_dff_A_FIEAXlDu9_0;
	wire w_dff_A_1tJXCDZH5_0;
	wire w_dff_A_l5gMOBei4_0;
	wire w_dff_A_8qXkLzQl9_0;
	wire w_dff_A_5sNSkv1N1_0;
	wire w_dff_A_ASJ4J5SQ2_0;
	wire w_dff_A_w4VHtvYt5_0;
	wire w_dff_A_gwDlvvGS8_2;
	wire w_dff_A_pyMSuIju5_0;
	wire w_dff_A_HvPMqq5t9_0;
	wire w_dff_A_UGyAlJ6Y0_0;
	wire w_dff_A_XSrtizU08_0;
	wire w_dff_A_8lN7DabA1_0;
	wire w_dff_A_HM3MKpQL8_2;
	wire w_dff_A_R6jWaAUu3_0;
	wire w_dff_A_MBiSDkNg6_0;
	wire w_dff_A_TiLs4IDp0_0;
	wire w_dff_A_f2y4bC435_0;
	wire w_dff_A_90iJhh3S3_2;
	wire w_dff_A_wMVTovFG7_0;
	wire w_dff_A_sNDuGX0S8_0;
	wire w_dff_A_cNEKW8gF0_0;
	wire w_dff_A_uimQMgSQ5_0;
	wire w_dff_A_QhnLDcRO1_0;
	wire w_dff_A_QndRye4D9_0;
	wire w_dff_A_Qp3H3yc01_0;
	wire w_dff_A_eTQMF5Qy7_0;
	wire w_dff_A_3fDqDu737_2;
	wire w_dff_A_7KFerPuq5_0;
	wire w_dff_A_5Zm3OgNo7_0;
	wire w_dff_A_1rPRtXIg7_0;
	wire w_dff_A_LUjSBSBl2_0;
	wire w_dff_A_xgQlfr3r4_0;
	wire w_dff_A_CdS7RY2u4_0;
	wire w_dff_A_q2DaGNrb1_0;
	wire w_dff_A_eOEDl1WL5_0;
	wire w_dff_A_F5JBNVEW3_2;
	wire w_dff_A_Phw1tJnA6_0;
	wire w_dff_A_4qm3SZjK2_2;
	wire w_dff_A_WDRkfbAT3_0;
	wire w_dff_A_LuZMZecF1_2;
	wire w_dff_A_8FT8dgJl5_0;
	wire w_dff_A_DpK9MJgg0_2;
	wire w_dff_A_XmzPJ8Z65_0;
	wire w_dff_A_e8tpRDF93_0;
	wire w_dff_A_4bsi1gVk1_0;
	wire w_dff_A_RwTLNT8w2_0;
	wire w_dff_A_WfdH0IHe9_0;
	wire w_dff_A_0MxlA2ET8_0;
	wire w_dff_A_fkKoHX4M6_0;
	wire w_dff_A_tVu4vRE77_0;
	wire w_dff_A_sPJrOy6n7_0;
	wire w_dff_A_MSlCcuJr7_0;
	wire w_dff_A_5Faf9DTs9_0;
	wire w_dff_A_ZD0wqzCR0_0;
	wire w_dff_A_uN8TCNXs0_0;
	wire w_dff_A_OJOU4HGP3_0;
	wire w_dff_A_vrTN3nrh9_0;
	wire w_dff_A_Yu8avxCL4_0;
	wire w_dff_A_2dEyfsHJ7_0;
	wire w_dff_A_Ztvpptee8_0;
	wire w_dff_A_MexYlLuv6_0;
	wire w_dff_A_skz1TVNd4_0;
	wire w_dff_A_ja4VovS83_0;
	wire w_dff_A_cO5F2zJo7_0;
	wire w_dff_A_EvNvKbhg4_0;
	wire w_dff_A_7S3hWtba7_0;
	wire w_dff_A_66Kxv2s37_2;
	wire w_dff_A_5FuhfzB66_0;
	wire w_dff_A_9k1mbw330_0;
	wire w_dff_A_0o1hTSuY3_0;
	wire w_dff_A_u2QOunfA3_0;
	wire w_dff_A_5HB4DTtw9_0;
	wire w_dff_A_Zf5g3S756_2;
	wire w_dff_A_WL258vLB9_0;
	wire w_dff_A_nyc2roSQ8_0;
	wire w_dff_A_wgWE2OIF4_0;
	wire w_dff_A_EQdiu7Rs7_0;
	wire w_dff_A_7s1UEE4E9_0;
	wire w_dff_A_5ZJ7pWXu5_2;
	wire w_dff_A_B9hm0S602_0;
	wire w_dff_A_62ACiwer7_0;
	wire w_dff_A_33B314zn1_0;
	wire w_dff_A_1ORmC1Rr9_0;
	wire w_dff_A_UD0mHw0Y8_0;
	wire w_dff_A_xlZ8L1W07_2;
	wire w_dff_A_8RsmyaiI5_0;
	wire w_dff_A_t1a9Lv1z5_0;
	wire w_dff_A_1mvlSIxx1_0;
	wire w_dff_A_OPuVijkx7_0;
	wire w_dff_A_pN6rLBLl2_0;
	wire w_dff_A_Enrz0vw03_0;
	wire w_dff_A_ZNa2zk2F9_0;
	wire w_dff_A_NpO6pto17_2;
	wire w_dff_A_yGWClJHQ3_0;
	wire w_dff_A_KVuEHkkb2_0;
	wire w_dff_A_Tx2EeQEC5_0;
	wire w_dff_A_TRwoNDg73_0;
	wire w_dff_A_hikfPZ1u3_0;
	wire w_dff_A_7TrXXuFg1_0;
	wire w_dff_A_xNhO77ex5_0;
	wire w_dff_A_LNfNVx5v9_0;
	wire w_dff_A_lNXZEEmI6_0;
	wire w_dff_A_sxzLpbNr9_0;
	wire w_dff_A_QgfBEcCl0_0;
	wire w_dff_A_H4nuQuD29_0;
	wire w_dff_A_RmMNSInv4_0;
	wire w_dff_A_Cn0gG3nw8_0;
	wire w_dff_A_oEcxtlaH3_0;
	wire w_dff_A_kBA3nHEg5_0;
	wire w_dff_A_z4pndscK5_0;
	wire w_dff_A_zg3xNFJl1_0;
	wire w_dff_A_Izr64Mtx0_0;
	wire w_dff_A_5xWKymr18_2;
	wire w_dff_A_HlcRKYcW8_0;
	wire w_dff_A_TNQyhMuw3_2;
	wire w_dff_A_kyRgxR5R7_0;
	wire w_dff_A_gjRLzgIm3_2;
	wire w_dff_A_JXazmYKP2_0;
	wire w_dff_A_bEIjtywn2_0;
	wire w_dff_A_tPHdV3u70_0;
	wire w_dff_A_Lca0kmFz9_0;
	wire w_dff_A_X3BxciBC4_0;
	wire w_dff_A_VfdZ5erP6_0;
	wire w_dff_A_nvN9YVzL6_0;
	wire w_dff_A_Ng5PWTK74_0;
	wire w_dff_A_SRISsozN2_0;
	wire w_dff_A_zK39wwoO4_0;
	wire w_dff_A_n9IPYTyO1_0;
	wire w_dff_A_4k3rMu2f9_0;
	wire w_dff_A_MAHEbFBd1_0;
	wire w_dff_A_Bmfi1Pd85_0;
	wire w_dff_A_JWsvIb9c8_0;
	wire w_dff_A_fy6XihzP7_0;
	wire w_dff_A_6wJk8jyM6_0;
	wire w_dff_A_A4XOy4fh6_2;
	wire w_dff_A_gTN6iNlU9_0;
	wire w_dff_A_GCu76aiM2_0;
	wire w_dff_A_Vc4je3797_0;
	wire w_dff_A_LcOUrM4m3_0;
	wire w_dff_A_Wp5C6Slw5_0;
	wire w_dff_A_j7MCRLo46_0;
	wire w_dff_A_DBJGPkYD5_0;
	wire w_dff_A_13cYZlMt2_0;
	wire w_dff_A_zTHqLjhk6_0;
	wire w_dff_A_6L7oKnnq6_0;
	wire w_dff_A_XyI0mOA96_0;
	wire w_dff_A_CpHfLnY25_0;
	wire w_dff_A_ZqUBEiYz9_0;
	wire w_dff_A_8yoyiDDb7_0;
	wire w_dff_A_0RTInmma9_0;
	wire w_dff_A_OhYKUvWI1_0;
	wire w_dff_A_UPZ5k5Xb9_0;
	wire w_dff_A_aqO8jZ6A6_2;
	wire w_dff_A_AZzDua9b3_0;
	wire w_dff_A_6YO4tzXl6_0;
	wire w_dff_A_o0UazIW82_0;
	wire w_dff_A_YOBdtfMA2_0;
	wire w_dff_A_uCogFCmT3_0;
	wire w_dff_A_xWT3jQs29_0;
	wire w_dff_A_72h9EVtj2_0;
	wire w_dff_A_YzK76lN63_0;
	wire w_dff_A_TCxdCZHY1_0;
	wire w_dff_A_2UzDimiZ9_0;
	wire w_dff_A_7PP1sbCB6_0;
	wire w_dff_A_fQgQo2ye7_0;
	wire w_dff_A_5VkYQ8El0_0;
	wire w_dff_A_YGpfq2Jd9_0;
	wire w_dff_A_aOSDakV86_0;
	wire w_dff_A_Li7dGMDe5_0;
	wire w_dff_A_6NQCOJIc2_0;
	wire w_dff_A_7pKYbPVy4_2;
	wire w_dff_A_WBGl0WpB8_0;
	wire w_dff_A_WhsXkAvs8_0;
	wire w_dff_A_CDe5Np1a1_0;
	wire w_dff_A_akKupNvi7_0;
	wire w_dff_A_iWlaiOJf0_0;
	wire w_dff_A_eQUQsWTy3_0;
	wire w_dff_A_adO26Uvs3_0;
	wire w_dff_A_LgSqa9uP7_0;
	wire w_dff_A_eHYOdJuD0_0;
	wire w_dff_A_06QDEm150_0;
	wire w_dff_A_Uk1kWr2b3_0;
	wire w_dff_A_jphJM6sA5_0;
	wire w_dff_A_KZnSz4oG9_0;
	wire w_dff_A_FsiRgk9F2_0;
	wire w_dff_A_npPxXng34_0;
	wire w_dff_A_tggbj35D0_0;
	wire w_dff_A_f6zmQDRH2_0;
	wire w_dff_A_QExPo0Wj9_2;
	wire w_dff_A_zjSrlHje7_0;
	wire w_dff_A_64PeerYV0_0;
	wire w_dff_A_joX9QhWi4_0;
	wire w_dff_A_F4x6EZGn9_0;
	wire w_dff_A_I58el1FW9_0;
	wire w_dff_A_n7JEDQ8V9_0;
	wire w_dff_A_Muat5UCv8_0;
	wire w_dff_A_npOvNuPR5_0;
	wire w_dff_A_cigL26PG5_0;
	wire w_dff_A_v1AWzzSo9_0;
	wire w_dff_A_6D9PtInS1_0;
	wire w_dff_A_77ssRZCb2_0;
	wire w_dff_A_RRVhlcbP2_2;
	wire w_dff_A_Y3duYJiR3_0;
	wire w_dff_A_XZea749D9_0;
	wire w_dff_A_cd9govl93_0;
	wire w_dff_A_BiAC9qPC4_0;
	wire w_dff_A_SdAU7V2Q1_0;
	wire w_dff_A_tVFX3nj97_0;
	wire w_dff_A_Xy2JumR71_0;
	wire w_dff_A_eZlrCZqr9_0;
	wire w_dff_A_hvHvB2zE9_0;
	wire w_dff_A_fYKJRhen9_0;
	wire w_dff_A_lCZJMyYO7_0;
	wire w_dff_A_ko2P7GjQ4_0;
	wire w_dff_A_Dtcr2t8E9_0;
	wire w_dff_A_lnookEJx5_2;
	wire w_dff_A_hFSAKiyw3_0;
	wire w_dff_A_JEcEXyYJ5_0;
	wire w_dff_A_xGtgUL8o3_0;
	wire w_dff_A_nB9rpTsv6_0;
	wire w_dff_A_WQGQdT9K8_0;
	wire w_dff_A_pl2xJzib4_0;
	wire w_dff_A_wnqCkNDS2_0;
	wire w_dff_A_HwJX9iCr2_0;
	wire w_dff_A_z4uEjMGn0_0;
	wire w_dff_A_3WBHduyB5_0;
	wire w_dff_A_klBuYOAh1_0;
	wire w_dff_A_8Wg1UBbA2_0;
	wire w_dff_A_o2PvDGlQ1_0;
	wire w_dff_A_RrFeEEwF1_0;
	wire w_dff_A_wX30sGNI9_0;
	wire w_dff_A_fSEwKRmD3_2;
	wire w_dff_A_tdsQ6rES9_0;
	wire w_dff_A_hLvOlyGW9_0;
	wire w_dff_A_Hwn6ljTY8_0;
	wire w_dff_A_6oZDhHqT0_0;
	wire w_dff_A_LAsdIJpO2_0;
	wire w_dff_A_ZTTy8cRz9_0;
	wire w_dff_A_oaqnHzPb4_0;
	wire w_dff_A_asSJdhsN3_0;
	wire w_dff_A_icCUAyOh3_0;
	wire w_dff_A_zGpUNtdD2_0;
	wire w_dff_A_UpoGRkq93_0;
	wire w_dff_A_bK9inClz4_0;
	wire w_dff_A_557gcgzR0_0;
	wire w_dff_A_iFGbiI5M0_0;
	wire w_dff_A_CMGYIz2W0_0;
	wire w_dff_A_G4LGUiy17_0;
	wire w_dff_A_C2zreAzv5_0;
	wire w_dff_A_kjGGFBjr5_2;
	wire w_dff_A_mIhX1E8q9_0;
	wire w_dff_A_63iv9Lgt4_0;
	wire w_dff_A_syg62Qgg5_0;
	wire w_dff_A_XbNGlsgT6_0;
	wire w_dff_A_ocJ5WiQt8_0;
	wire w_dff_A_3AVLPWfs6_2;
	wire w_dff_A_oM4MwWtI5_2;
	wire w_dff_A_o8QafsO16_0;
	wire w_dff_A_Jqd4xWpb1_0;
	wire w_dff_A_Yo2qFoKU9_0;
	wire w_dff_A_pom0h5kE6_0;
	wire w_dff_A_OozD2UhM1_0;
	wire w_dff_A_BgCpmlhe9_0;
	wire w_dff_A_QBrIUpQs0_0;
	wire w_dff_A_NpIy8QxP0_0;
	wire w_dff_A_eRzlU6yE5_0;
	wire w_dff_A_bi5YO1QB7_0;
	wire w_dff_A_patlHC8c3_0;
	wire w_dff_A_HCOqsXlx4_0;
	wire w_dff_A_caS97pzf2_0;
	wire w_dff_A_5HZDyfup5_0;
	wire w_dff_A_04DFZzRO4_0;
	wire w_dff_A_iBbCuLEp4_0;
	wire w_dff_A_SZHKifOh5_2;
	wire w_dff_A_xrM9NinU7_0;
	wire w_dff_A_faxxTd5s3_0;
	wire w_dff_A_4ctQpcnd2_0;
	wire w_dff_A_iDNk4g734_0;
	wire w_dff_A_PSY8VEdo3_0;
	wire w_dff_A_eOFAMxXJ6_0;
	wire w_dff_A_QS29gxdM5_0;
	wire w_dff_A_UqQwMQpd0_0;
	wire w_dff_A_sNl1j9sY2_0;
	wire w_dff_A_eVXWxF4r8_0;
	wire w_dff_A_LVLxvjpj1_0;
	wire w_dff_A_utWrhI8o3_0;
	wire w_dff_A_j3c1f5To7_0;
	wire w_dff_A_EnSTdf7g6_0;
	wire w_dff_A_1vJFTEEo4_0;
	wire w_dff_A_Jt6aMDQ94_0;
	wire w_dff_A_9ZIm3fD33_0;
	wire w_dff_A_2MSuZMVk5_0;
	wire w_dff_A_Tm1UH8M69_0;
	wire w_dff_A_qp69ew1k3_0;
	jnot g0000(.din(w_G15_0[2]),.dout(w_dff_A_TnC3fYtR3_1),.clk(gclk));
	jor g0001(.dina(G57),.dinb(w_G5_1[1]),.dout(w_dff_A_158BVJfx5_2),.clk(gclk));
	jnot g0002(.din(G184),.dout(n317),.clk(gclk));
	jnot g0003(.din(G228),.dout(n318),.clk(gclk));
	jor g0004(.dina(n318),.dinb(n317),.dout(n319),.clk(gclk));
	jnot g0005(.din(G150),.dout(n320),.clk(gclk));
	jnot g0006(.din(G240),.dout(n321),.clk(gclk));
	jor g0007(.dina(n321),.dinb(n320),.dout(n322),.clk(gclk));
	jor g0008(.dina(n322),.dinb(n319),.dout(G404_fa_),.clk(gclk));
	jnot g0009(.din(G210),.dout(n324),.clk(gclk));
	jnot g0010(.din(G218),.dout(n325),.clk(gclk));
	jor g0011(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jnot g0012(.din(G152),.dout(n327),.clk(gclk));
	jnot g0013(.din(G230),.dout(n328),.clk(gclk));
	jor g0014(.dina(n328),.dinb(n327),.dout(n329),.clk(gclk));
	jor g0015(.dina(n329),.dinb(n326),.dout(G406_fa_),.clk(gclk));
	jnot g0016(.din(G183),.dout(n331),.clk(gclk));
	jnot g0017(.din(G185),.dout(n332),.clk(gclk));
	jor g0018(.dina(n332),.dinb(n331),.dout(n333),.clk(gclk));
	jnot g0019(.din(G182),.dout(n334),.clk(gclk));
	jnot g0020(.din(G186),.dout(n335),.clk(gclk));
	jor g0021(.dina(n335),.dinb(n334),.dout(n336),.clk(gclk));
	jor g0022(.dina(n336),.dinb(n333),.dout(G408_fa_),.clk(gclk));
	jnot g0023(.din(G172),.dout(n338),.clk(gclk));
	jnot g0024(.din(G188),.dout(n339),.clk(gclk));
	jor g0025(.dina(n339),.dinb(n338),.dout(n340),.clk(gclk));
	jnot g0026(.din(G162),.dout(n341),.clk(gclk));
	jnot g0027(.din(G199),.dout(n342),.clk(gclk));
	jor g0028(.dina(n342),.dinb(n341),.dout(n343),.clk(gclk));
	jor g0029(.dina(n343),.dinb(n340),.dout(G410_fa_),.clk(gclk));
	jnot g0030(.din(G1197),.dout(n345),.clk(gclk));
	jor g0031(.dina(w_n345_0[1]),.dinb(w_G5_1[0]),.dout(w_dff_A_ssThCr5Y4_2),.clk(gclk));
	jnot g0032(.din(G134),.dout(n347),.clk(gclk));
	jnot g0033(.din(G133),.dout(n348),.clk(gclk));
	jor g0034(.dina(n348),.dinb(w_G5_0[2]),.dout(n349),.clk(gclk));
	jor g0035(.dina(w_n349_0[1]),.dinb(w_n347_0[1]),.dout(w_dff_A_x6bwFvue0_2),.clk(gclk));
	jand g0036(.dina(G163),.dinb(w_G1_1[2]),.dout(w_dff_A_EbglPHaX6_2),.clk(gclk));
	jnot g0037(.din(w_G41_0[1]),.dout(n352),.clk(gclk));
	jor g0038(.dina(n352),.dinb(w_G18_49[2]),.dout(n353),.clk(gclk));
	jor g0039(.dina(w_n353_0[1]),.dinb(w_G3701_1[1]),.dout(n354),.clk(gclk));
	jnot g0040(.din(w_G18_49[1]),.dout(n355),.clk(gclk));
	jand g0041(.dina(w_G3701_1[0]),.dinb(w_n355_35[2]),.dout(n356),.clk(gclk));
	jand g0042(.dina(n356),.dinb(w_n353_0[0]),.dout(n357),.clk(gclk));
	jnot g0043(.din(w_n357_0[1]),.dout(n358),.clk(gclk));
	jand g0044(.dina(w_n358_0[1]),.dinb(w_n354_0[2]),.dout(n359),.clk(gclk));
	jxor g0045(.dina(w_n359_1[1]),.dinb(w_G4526_2[2]),.dout(w_dff_A_S8QuRzkE0_2),.clk(gclk));
	jnot g0046(.din(w_G38_2[2]),.dout(n361),.clk(gclk));
	jand g0047(.dina(w_G4528_0[2]),.dinb(w_G1492_1[1]),.dout(n362),.clk(gclk));
	jxor g0048(.dina(w_n362_0[2]),.dinb(w_n361_0[2]),.dout(n363),.clk(gclk));
	jand g0049(.dina(w_G4528_0[1]),.dinb(w_G1496_1[1]),.dout(n364),.clk(gclk));
	jor g0050(.dina(w_n364_0[2]),.dinb(w_n361_0[1]),.dout(n365),.clk(gclk));
	jnot g0051(.din(w_G1496_1[0]),.dout(n366),.clk(gclk));
	jnot g0052(.din(w_G4528_0[0]),.dout(n367),.clk(gclk));
	jor g0053(.dina(w_n367_0[1]),.dinb(w_G38_2[1]),.dout(n368),.clk(gclk));
	jor g0054(.dina(w_n368_0[1]),.dinb(w_n366_0[2]),.dout(n369),.clk(gclk));
	jand g0055(.dina(w_n369_0[1]),.dinb(w_dff_B_gPMZX7B71_1),.dout(n370),.clk(gclk));
	jnot g0056(.din(w_G1486_0[1]),.dout(n371),.clk(gclk));
	jand g0057(.dina(G12),.dinb(G9),.dout(n372),.clk(gclk));
	jnot g0058(.din(w_n372_0[1]),.dout(n373),.clk(gclk));
	jor g0059(.dina(w_dff_B_a909KlhV4_0),.dinb(w_n355_35[1]),.dout(n374),.clk(gclk));
	jand g0060(.dina(w_n374_0[1]),.dinb(w_n373_9[2]),.dout(n375),.clk(gclk));
	jand g0061(.dina(w_n375_0[2]),.dinb(w_n371_0[2]),.dout(n376),.clk(gclk));
	jxor g0062(.dina(w_n375_0[1]),.dinb(w_n371_0[1]),.dout(n377),.clk(gclk));
	jor g0063(.dina(w_dff_B_vxvT3Qbl3_0),.dinb(w_n355_35[0]),.dout(n378),.clk(gclk));
	jand g0064(.dina(w_n378_0[1]),.dinb(w_n373_9[1]),.dout(n379),.clk(gclk));
	jnot g0065(.din(w_n379_0[2]),.dout(n380),.clk(gclk));
	jand g0066(.dina(w_n380_0[1]),.dinb(w_G1480_0[2]),.dout(n381),.clk(gclk));
	jnot g0067(.din(n381),.dout(n382),.clk(gclk));
	jnot g0068(.din(w_G1480_0[1]),.dout(n383),.clk(gclk));
	jand g0069(.dina(w_n379_0[1]),.dinb(w_n383_0[2]),.dout(n384),.clk(gclk));
	jnot g0070(.din(w_G106_1[1]),.dout(n385),.clk(gclk));
	jor g0071(.dina(w_dff_B_ZagUfvbl0_0),.dinb(w_n355_34[2]),.dout(n386),.clk(gclk));
	jand g0072(.dina(w_n386_0[1]),.dinb(w_n373_9[0]),.dout(n387),.clk(gclk));
	jxor g0073(.dina(w_n387_1[1]),.dinb(w_n385_0[1]),.dout(n388),.clk(gclk));
	jnot g0074(.din(w_G1462_0[1]),.dout(n389),.clk(gclk));
	jor g0075(.dina(w_G209_0[1]),.dinb(w_n355_34[1]),.dout(n390),.clk(gclk));
	jand g0076(.dina(n390),.dinb(w_n373_8[2]),.dout(n391),.clk(gclk));
	jand g0077(.dina(w_n391_0[2]),.dinb(w_n389_1[1]),.dout(n392),.clk(gclk));
	jnot g0078(.din(w_G1469_0[1]),.dout(n393),.clk(gclk));
	jor g0079(.dina(w_dff_B_bZf3Y5AV4_0),.dinb(w_n355_34[0]),.dout(n394),.clk(gclk));
	jand g0080(.dina(w_n394_0[1]),.dinb(w_n373_8[1]),.dout(n395),.clk(gclk));
	jxor g0081(.dina(w_n395_1[1]),.dinb(w_n393_1[1]),.dout(n396),.clk(gclk));
	jand g0082(.dina(w_n396_1[2]),.dinb(w_n392_0[2]),.dout(n397),.clk(gclk));
	jand g0083(.dina(w_n397_0[1]),.dinb(w_n388_1[2]),.dout(n398),.clk(gclk));
	jnot g0084(.din(n398),.dout(n399),.clk(gclk));
	jand g0085(.dina(w_n387_1[0]),.dinb(w_n385_0[0]),.dout(n400),.clk(gclk));
	jnot g0086(.din(n400),.dout(n401),.clk(gclk));
	jnot g0087(.din(w_n387_0[2]),.dout(n402),.clk(gclk));
	jand g0088(.dina(n402),.dinb(w_G106_1[0]),.dout(n403),.clk(gclk));
	jand g0089(.dina(w_n395_1[0]),.dinb(w_n393_1[0]),.dout(n404),.clk(gclk));
	jnot g0090(.din(n404),.dout(n405),.clk(gclk));
	jor g0091(.dina(w_n405_0[2]),.dinb(n403),.dout(n406),.clk(gclk));
	jand g0092(.dina(n406),.dinb(w_dff_B_ip9tF0zH7_1),.dout(n407),.clk(gclk));
	jand g0093(.dina(w_n407_0[1]),.dinb(n399),.dout(n408),.clk(gclk));
	jnot g0094(.din(n408),.dout(n409),.clk(gclk));
	jor g0095(.dina(w_n409_1[1]),.dinb(w_dff_B_Cw6wK2kq0_1),.dout(n410),.clk(gclk));
	jand g0096(.dina(n410),.dinb(w_dff_B_9j5IoNto8_1),.dout(n411),.clk(gclk));
	jand g0097(.dina(w_n411_1[1]),.dinb(w_n377_1[2]),.dout(n412),.clk(gclk));
	jor g0098(.dina(n412),.dinb(w_dff_B_GP6CBlmT3_1),.dout(n413),.clk(gclk));
	jxor g0099(.dina(w_n391_0[1]),.dinb(w_n389_1[0]),.dout(n414),.clk(gclk));
	jand g0100(.dina(w_n414_1[1]),.dinb(w_n396_1[1]),.dout(n415),.clk(gclk));
	jxor g0101(.dina(w_n379_0[0]),.dinb(w_n383_0[1]),.dout(n416),.clk(gclk));
	jand g0102(.dina(w_n416_0[2]),.dinb(w_n388_1[1]),.dout(n417),.clk(gclk));
	jand g0103(.dina(n417),.dinb(w_n415_0[1]),.dout(n418),.clk(gclk));
	jand g0104(.dina(w_n418_0[1]),.dinb(w_n377_1[1]),.dout(n419),.clk(gclk));
	jor g0105(.dina(w_n419_0[1]),.dinb(w_n413_1[1]),.dout(n420),.clk(gclk));
	jnot g0106(.din(w_G2256_0[1]),.dout(n421),.clk(gclk));
	jor g0107(.dina(w_dff_B_KrwkUrhI8_0),.dinb(w_n355_33[2]),.dout(n422),.clk(gclk));
	jand g0108(.dina(w_n422_0[1]),.dinb(w_n373_8[0]),.dout(n423),.clk(gclk));
	jand g0109(.dina(w_n423_0[2]),.dinb(w_n421_0[2]),.dout(n424),.clk(gclk));
	jxor g0110(.dina(w_n423_0[1]),.dinb(w_n421_0[1]),.dout(n425),.clk(gclk));
	jnot g0111(.din(w_G2253_0[2]),.dout(n426),.clk(gclk));
	jor g0112(.dina(w_dff_B_8UG59Vca7_0),.dinb(w_n355_33[1]),.dout(n427),.clk(gclk));
	jand g0113(.dina(w_n427_0[1]),.dinb(w_n373_7[2]),.dout(n428),.clk(gclk));
	jxor g0114(.dina(w_n428_0[2]),.dinb(w_n426_0[2]),.dout(n429),.clk(gclk));
	jnot g0115(.din(w_G2247_0[2]),.dout(n430),.clk(gclk));
	jor g0116(.dina(w_dff_B_F1xHy1Kr0_0),.dinb(w_n355_33[0]),.dout(n431),.clk(gclk));
	jand g0117(.dina(w_n431_0[1]),.dinb(w_n373_7[1]),.dout(n432),.clk(gclk));
	jxor g0118(.dina(w_n432_0[2]),.dinb(w_n430_0[1]),.dout(n433),.clk(gclk));
	jnot g0119(.din(w_G2239_1[1]),.dout(n434),.clk(gclk));
	jor g0120(.dina(w_dff_B_wEA3Mhyp8_0),.dinb(w_n355_32[2]),.dout(n435),.clk(gclk));
	jand g0121(.dina(w_n435_0[1]),.dinb(w_n373_7[0]),.dout(n436),.clk(gclk));
	jxor g0122(.dina(w_n436_0[2]),.dinb(w_n434_0[1]),.dout(n437),.clk(gclk));
	jand g0123(.dina(w_n437_0[2]),.dinb(w_n433_1[2]),.dout(n438),.clk(gclk));
	jand g0124(.dina(w_n438_0[1]),.dinb(w_n429_0[2]),.dout(n439),.clk(gclk));
	jnot g0125(.din(w_n428_0[1]),.dout(n440),.clk(gclk));
	jand g0126(.dina(w_n440_0[1]),.dinb(w_G2253_0[1]),.dout(n441),.clk(gclk));
	jnot g0127(.din(n441),.dout(n442),.clk(gclk));
	jand g0128(.dina(w_n428_0[0]),.dinb(w_n426_0[1]),.dout(n443),.clk(gclk));
	jand g0129(.dina(w_n432_0[1]),.dinb(w_n430_0[0]),.dout(n444),.clk(gclk));
	jand g0130(.dina(w_n436_0[1]),.dinb(w_n434_0[0]),.dout(n445),.clk(gclk));
	jand g0131(.dina(w_n445_0[2]),.dinb(w_n433_1[1]),.dout(n446),.clk(gclk));
	jor g0132(.dina(n446),.dinb(w_n444_0[2]),.dout(n447),.clk(gclk));
	jor g0133(.dina(w_n447_0[2]),.dinb(w_dff_B_2P3d0CEE3_1),.dout(n448),.clk(gclk));
	jand g0134(.dina(n448),.dinb(w_dff_B_pVUVu6oE9_1),.dout(n449),.clk(gclk));
	jor g0135(.dina(w_n449_1[1]),.dinb(w_dff_B_BiI0ZTCU1_1),.dout(n450),.clk(gclk));
	jnot g0136(.din(w_G2236_0[2]),.dout(n451),.clk(gclk));
	jor g0137(.dina(w_dff_B_1NhAGwVz7_0),.dinb(w_n355_32[1]),.dout(n452),.clk(gclk));
	jand g0138(.dina(n452),.dinb(w_n373_6[2]),.dout(n453),.clk(gclk));
	jand g0139(.dina(w_n453_1[1]),.dinb(w_n451_0[2]),.dout(n454),.clk(gclk));
	jor g0140(.dina(w_n453_1[0]),.dinb(w_n451_0[1]),.dout(n455),.clk(gclk));
	jnot g0141(.din(w_G2230_0[2]),.dout(n456),.clk(gclk));
	jand g0142(.dina(w_dff_B_W1sljb7y0_0),.dinb(w_n355_32[0]),.dout(n457),.clk(gclk));
	jand g0143(.dina(G158),.dinb(w_G18_49[0]),.dout(n458),.clk(gclk));
	jor g0144(.dina(w_dff_B_4ktNGoya8_0),.dinb(w_n457_0[1]),.dout(n459),.clk(gclk));
	jand g0145(.dina(w_n459_0[2]),.dinb(w_n456_0[2]),.dout(n460),.clk(gclk));
	jand g0146(.dina(w_n460_1[2]),.dinb(n455),.dout(n461),.clk(gclk));
	jor g0147(.dina(n461),.dinb(w_dff_B_ROfqi5sd5_1),.dout(n462),.clk(gclk));
	jxor g0148(.dina(w_n453_0[2]),.dinb(w_n451_0[0]),.dout(n463),.clk(gclk));
	jxor g0149(.dina(w_n459_0[1]),.dinb(w_n456_0[1]),.dout(n464),.clk(gclk));
	jand g0150(.dina(w_n464_0[2]),.dinb(w_n463_1[1]),.dout(n465),.clk(gclk));
	jnot g0151(.din(w_G2224_1[1]),.dout(n466),.clk(gclk));
	jand g0152(.dina(w_dff_B_FXRdcySs7_0),.dinb(w_n355_31[2]),.dout(n467),.clk(gclk));
	jand g0153(.dina(G159),.dinb(w_G18_48[2]),.dout(n468),.clk(gclk));
	jor g0154(.dina(w_dff_B_s4eA4dZI1_0),.dinb(w_n467_0[1]),.dout(n469),.clk(gclk));
	jxor g0155(.dina(w_n469_1[1]),.dinb(w_n466_0[1]),.dout(n470),.clk(gclk));
	jnot g0156(.din(w_G2218_0[2]),.dout(n471),.clk(gclk));
	jand g0157(.dina(w_dff_B_i95EsnAB8_0),.dinb(w_n355_31[1]),.dout(n472),.clk(gclk));
	jand g0158(.dina(G160),.dinb(w_G18_48[1]),.dout(n473),.clk(gclk));
	jor g0159(.dina(w_dff_B_MQuA8mp51_0),.dinb(w_n472_0[1]),.dout(n474),.clk(gclk));
	jxor g0160(.dina(w_n474_0[2]),.dinb(w_n471_0[2]),.dout(n475),.clk(gclk));
	jnot g0161(.din(w_G2211_0[2]),.dout(n476),.clk(gclk));
	jand g0162(.dina(w_dff_B_0RG5tioS2_0),.dinb(w_n355_31[0]),.dout(n477),.clk(gclk));
	jand g0163(.dina(G151),.dinb(w_G18_48[0]),.dout(n478),.clk(gclk));
	jor g0164(.dina(w_dff_B_tvoDF4FO0_0),.dinb(w_n477_0[1]),.dout(n479),.clk(gclk));
	jxor g0165(.dina(w_n479_1[1]),.dinb(w_n476_0[2]),.dout(n480),.clk(gclk));
	jand g0166(.dina(w_n480_1[1]),.dinb(w_n475_0[2]),.dout(n481),.clk(gclk));
	jand g0167(.dina(w_n481_0[1]),.dinb(w_n470_0[2]),.dout(n482),.clk(gclk));
	jnot g0168(.din(w_n469_1[0]),.dout(n483),.clk(gclk));
	jand g0169(.dina(n483),.dinb(w_G2224_1[0]),.dout(n484),.clk(gclk));
	jnot g0170(.din(w_n474_0[1]),.dout(n485),.clk(gclk));
	jand g0171(.dina(w_n485_0[1]),.dinb(w_G2218_0[1]),.dout(n486),.clk(gclk));
	jand g0172(.dina(w_n479_1[0]),.dinb(w_n476_0[1]),.dout(n487),.clk(gclk));
	jnot g0173(.din(w_n487_0[2]),.dout(n488),.clk(gclk));
	jor g0174(.dina(n488),.dinb(w_n486_0[1]),.dout(n489),.clk(gclk));
	jand g0175(.dina(w_n469_0[2]),.dinb(w_n466_0[0]),.dout(n490),.clk(gclk));
	jand g0176(.dina(w_n474_0[0]),.dinb(w_n471_0[1]),.dout(n491),.clk(gclk));
	jor g0177(.dina(w_n491_1[1]),.dinb(n490),.dout(n492),.clk(gclk));
	jnot g0178(.din(n492),.dout(n493),.clk(gclk));
	jand g0179(.dina(n493),.dinb(w_n489_0[2]),.dout(n494),.clk(gclk));
	jor g0180(.dina(n494),.dinb(w_dff_B_GMRm2J0a2_1),.dout(n495),.clk(gclk));
	jnot g0181(.din(w_n495_1[1]),.dout(n496),.clk(gclk));
	jor g0182(.dina(w_n496_0[2]),.dinb(w_dff_B_gyQ2zbRa9_1),.dout(n497),.clk(gclk));
	jand g0183(.dina(w_n497_1[1]),.dinb(w_n465_0[1]),.dout(n498),.clk(gclk));
	jor g0184(.dina(n498),.dinb(w_n462_0[2]),.dout(n499),.clk(gclk));
	jand g0185(.dina(w_n496_0[1]),.dinb(w_n465_0[0]),.dout(n500),.clk(gclk));
	jnot g0186(.din(w_G4437_0[2]),.dout(n501),.clk(gclk));
	jand g0187(.dina(G219),.dinb(w_G18_47[2]),.dout(n502),.clk(gclk));
	jand g0188(.dina(w_dff_B_K91H5ioU1_0),.dinb(w_n355_30[2]),.dout(n503),.clk(gclk));
	jor g0189(.dina(w_n503_0[1]),.dinb(w_dff_B_Wb2jObOc6_1),.dout(n504),.clk(gclk));
	jand g0190(.dina(w_n504_1[1]),.dinb(w_n501_0[2]),.dout(n505),.clk(gclk));
	jnot g0191(.din(w_n504_1[0]),.dout(n506),.clk(gclk));
	jand g0192(.dina(n506),.dinb(w_G4437_0[1]),.dout(n507),.clk(gclk));
	jnot g0193(.din(w_n507_0[1]),.dout(n508),.clk(gclk));
	jnot g0194(.din(w_G4432_0[2]),.dout(n509),.clk(gclk));
	jand g0195(.dina(G220),.dinb(w_G18_47[1]),.dout(n510),.clk(gclk));
	jand g0196(.dina(w_dff_B_GlAauAlX5_0),.dinb(w_n355_30[1]),.dout(n511),.clk(gclk));
	jor g0197(.dina(w_n511_0[1]),.dinb(w_dff_B_S7QK8PnQ1_1),.dout(n512),.clk(gclk));
	jxor g0198(.dina(w_n512_0[2]),.dinb(w_n509_0[2]),.dout(n513),.clk(gclk));
	jnot g0199(.din(w_G4420_1[1]),.dout(n514),.clk(gclk));
	jand g0200(.dina(G222),.dinb(w_G18_47[0]),.dout(n515),.clk(gclk));
	jand g0201(.dina(w_dff_B_ZDKRkgen7_0),.dinb(w_n355_30[0]),.dout(n516),.clk(gclk));
	jor g0202(.dina(w_n516_0[1]),.dinb(w_dff_B_1BBgLLMX6_1),.dout(n517),.clk(gclk));
	jand g0203(.dina(w_n517_1[1]),.dinb(w_n514_0[1]),.dout(n518),.clk(gclk));
	jnot g0204(.din(w_n518_1[2]),.dout(n519),.clk(gclk));
	jnot g0205(.din(w_G4427_0[2]),.dout(n520),.clk(gclk));
	jand g0206(.dina(G221),.dinb(w_G18_46[2]),.dout(n521),.clk(gclk));
	jand g0207(.dina(w_dff_B_Tf4sktAQ5_0),.dinb(w_n355_29[2]),.dout(n522),.clk(gclk));
	jor g0208(.dina(w_n522_0[1]),.dinb(w_dff_B_hfhO92eX9_1),.dout(n523),.clk(gclk));
	jxor g0209(.dina(w_n523_0[2]),.dinb(w_n520_0[1]),.dout(n524),.clk(gclk));
	jnot g0210(.din(w_n517_1[0]),.dout(n525),.clk(gclk));
	jand g0211(.dina(n525),.dinb(w_G4420_1[0]),.dout(n526),.clk(gclk));
	jnot g0212(.din(w_n526_0[2]),.dout(n527),.clk(gclk));
	jnot g0213(.din(w_G4415_1[1]),.dout(n528),.clk(gclk));
	jand g0214(.dina(G223),.dinb(w_G18_46[1]),.dout(n529),.clk(gclk));
	jand g0215(.dina(w_dff_B_zO4tm7vU4_0),.dinb(w_n355_29[1]),.dout(n530),.clk(gclk));
	jor g0216(.dina(w_n530_0[1]),.dinb(w_dff_B_hpaCQnrD8_1),.dout(n531),.clk(gclk));
	jand g0217(.dina(w_n531_1[1]),.dinb(w_n528_0[1]),.dout(n532),.clk(gclk));
	jnot g0218(.din(w_n531_1[0]),.dout(n533),.clk(gclk));
	jand g0219(.dina(n533),.dinb(w_G4415_1[0]),.dout(n534),.clk(gclk));
	jnot g0220(.din(n534),.dout(n535),.clk(gclk));
	jnot g0221(.din(w_G4410_0[2]),.dout(n536),.clk(gclk));
	jand g0222(.dina(G224),.dinb(w_G18_46[0]),.dout(n537),.clk(gclk));
	jand g0223(.dina(w_dff_B_VTqLAKE61_0),.dinb(w_n355_29[0]),.dout(n538),.clk(gclk));
	jor g0224(.dina(w_n538_0[1]),.dinb(w_dff_B_eBTD6XLU8_1),.dout(n539),.clk(gclk));
	jand g0225(.dina(w_n539_1[1]),.dinb(w_n536_0[2]),.dout(n540),.clk(gclk));
	jnot g0226(.din(w_n539_1[0]),.dout(n541),.clk(gclk));
	jand g0227(.dina(n541),.dinb(w_G4410_0[1]),.dout(n542),.clk(gclk));
	jnot g0228(.din(n542),.dout(n543),.clk(gclk));
	jnot g0229(.din(w_G4405_1[1]),.dout(n544),.clk(gclk));
	jand g0230(.dina(G225),.dinb(w_G18_45[2]),.dout(n545),.clk(gclk));
	jand g0231(.dina(w_dff_B_NdacBAVQ8_0),.dinb(w_n355_28[2]),.dout(n546),.clk(gclk));
	jor g0232(.dina(w_n546_0[1]),.dinb(w_dff_B_lncsuzpc2_1),.dout(n547),.clk(gclk));
	jand g0233(.dina(w_n547_1[1]),.dinb(w_n544_0[1]),.dout(n548),.clk(gclk));
	jnot g0234(.din(w_n547_1[0]),.dout(n549),.clk(gclk));
	jand g0235(.dina(n549),.dinb(w_G4405_1[0]),.dout(n550),.clk(gclk));
	jnot g0236(.din(w_n550_0[1]),.dout(n551),.clk(gclk));
	jnot g0237(.din(w_G4400_1[1]),.dout(n552),.clk(gclk));
	jand g0238(.dina(G226),.dinb(w_G18_45[1]),.dout(n553),.clk(gclk));
	jand g0239(.dina(w_dff_B_d32fgfP58_0),.dinb(w_n355_28[1]),.dout(n554),.clk(gclk));
	jor g0240(.dina(w_n554_0[1]),.dinb(w_dff_B_Ay4BhMt72_1),.dout(n555),.clk(gclk));
	jand g0241(.dina(w_n555_1[1]),.dinb(w_n552_0[1]),.dout(n556),.clk(gclk));
	jnot g0242(.din(w_n555_1[0]),.dout(n557),.clk(gclk));
	jand g0243(.dina(n557),.dinb(w_G4400_1[0]),.dout(n558),.clk(gclk));
	jnot g0244(.din(w_n558_0[1]),.dout(n559),.clk(gclk));
	jnot g0245(.din(w_G4394_1[1]),.dout(n560),.clk(gclk));
	jand g0246(.dina(G217),.dinb(w_G18_45[0]),.dout(n561),.clk(gclk));
	jand g0247(.dina(w_dff_B_B9vMYkRe1_0),.dinb(w_n355_28[0]),.dout(n562),.clk(gclk));
	jor g0248(.dina(w_n562_0[1]),.dinb(w_dff_B_zfeiiKV59_1),.dout(n563),.clk(gclk));
	jand g0249(.dina(w_n563_1[1]),.dinb(w_n560_0[1]),.dout(n564),.clk(gclk));
	jand g0250(.dina(w_n564_0[2]),.dinb(n559),.dout(n565),.clk(gclk));
	jor g0251(.dina(w_n565_0[1]),.dinb(w_n556_0[2]),.dout(n566),.clk(gclk));
	jand g0252(.dina(w_n566_0[2]),.dinb(w_dff_B_Md0cH27z3_1),.dout(n567),.clk(gclk));
	jor g0253(.dina(n567),.dinb(w_n548_0[1]),.dout(n568),.clk(gclk));
	jand g0254(.dina(w_n568_0[2]),.dinb(w_dff_B_Hit352gK4_1),.dout(n569),.clk(gclk));
	jor g0255(.dina(n569),.dinb(w_dff_B_aKKKoBAO2_1),.dout(n570),.clk(gclk));
	jand g0256(.dina(w_n570_1[2]),.dinb(w_dff_B_o9pz9yqM5_1),.dout(n571),.clk(gclk));
	jor g0257(.dina(n571),.dinb(w_dff_B_w5dep8MM1_1),.dout(n572),.clk(gclk));
	jxor g0258(.dina(w_n531_0[2]),.dinb(w_n528_0[0]),.dout(n573),.clk(gclk));
	jxor g0259(.dina(w_n555_0[2]),.dinb(w_n552_0[0]),.dout(n574),.clk(gclk));
	jxor g0260(.dina(w_n563_1[0]),.dinb(w_n560_0[0]),.dout(n575),.clk(gclk));
	jand g0261(.dina(w_n575_1[1]),.dinb(w_n574_0[2]),.dout(n576),.clk(gclk));
	jxor g0262(.dina(w_n539_0[2]),.dinb(w_n536_0[1]),.dout(n577),.clk(gclk));
	jxor g0263(.dina(w_n547_0[2]),.dinb(w_n544_0[0]),.dout(n578),.clk(gclk));
	jand g0264(.dina(w_n578_0[2]),.dinb(w_n577_0[1]),.dout(n579),.clk(gclk));
	jand g0265(.dina(n579),.dinb(w_n576_0[2]),.dout(n580),.clk(gclk));
	jand g0266(.dina(w_n580_0[2]),.dinb(w_n573_1[1]),.dout(n581),.clk(gclk));
	jnot g0267(.din(w_G3749_0[2]),.dout(n582),.clk(gclk));
	jand g0268(.dina(G231),.dinb(w_G18_44[2]),.dout(n583),.clk(gclk));
	jand g0269(.dina(w_dff_B_pbQHyWMd6_0),.dinb(w_n355_27[2]),.dout(n584),.clk(gclk));
	jor g0270(.dina(w_n584_0[1]),.dinb(w_dff_B_izFmWNtm7_1),.dout(n585),.clk(gclk));
	jand g0271(.dina(w_n585_1[1]),.dinb(w_n582_0[2]),.dout(n586),.clk(gclk));
	jnot g0272(.din(w_n585_1[0]),.dout(n587),.clk(gclk));
	jand g0273(.dina(n587),.dinb(w_G3749_0[1]),.dout(n588),.clk(gclk));
	jnot g0274(.din(w_n588_0[1]),.dout(n589),.clk(gclk));
	jnot g0275(.din(w_G3743_0[2]),.dout(n590),.clk(gclk));
	jand g0276(.dina(G232),.dinb(w_G18_44[1]),.dout(n591),.clk(gclk));
	jand g0277(.dina(w_dff_B_Vz2Xni5H6_0),.dinb(w_n355_27[1]),.dout(n592),.clk(gclk));
	jor g0278(.dina(w_n592_0[1]),.dinb(w_dff_B_0Y1cWcdy6_1),.dout(n593),.clk(gclk));
	jxor g0279(.dina(w_n593_1[1]),.dinb(w_n590_0[2]),.dout(n594),.clk(gclk));
	jnot g0280(.din(w_G3737_0[2]),.dout(n595),.clk(gclk));
	jand g0281(.dina(G233),.dinb(w_G18_44[0]),.dout(n596),.clk(gclk));
	jand g0282(.dina(w_dff_B_XAFmI2px1_0),.dinb(w_n355_27[0]),.dout(n597),.clk(gclk));
	jor g0283(.dina(w_n597_0[1]),.dinb(w_dff_B_XueDhB7k7_1),.dout(n598),.clk(gclk));
	jxor g0284(.dina(w_n598_1[1]),.dinb(w_n595_0[2]),.dout(n599),.clk(gclk));
	jnot g0285(.din(w_G3729_1[1]),.dout(n600),.clk(gclk));
	jand g0286(.dina(G234),.dinb(w_G18_43[2]),.dout(n601),.clk(gclk));
	jand g0287(.dina(w_dff_B_0p2ojq8i8_0),.dinb(w_n355_26[2]),.dout(n602),.clk(gclk));
	jor g0288(.dina(w_n602_0[1]),.dinb(w_dff_B_lULSSn2v6_1),.dout(n603),.clk(gclk));
	jxor g0289(.dina(w_n603_1[1]),.dinb(w_n600_0[1]),.dout(n604),.clk(gclk));
	jand g0290(.dina(w_n604_0[1]),.dinb(w_n599_0[2]),.dout(n605),.clk(gclk));
	jand g0291(.dina(w_n605_0[2]),.dinb(w_n594_0[2]),.dout(n606),.clk(gclk));
	jnot g0292(.din(n606),.dout(n607),.clk(gclk));
	jnot g0293(.din(w_n593_1[0]),.dout(n608),.clk(gclk));
	jand g0294(.dina(n608),.dinb(w_G3743_0[1]),.dout(n609),.clk(gclk));
	jand g0295(.dina(w_n593_0[2]),.dinb(w_n590_0[1]),.dout(n610),.clk(gclk));
	jnot g0296(.din(w_n610_0[1]),.dout(n611),.clk(gclk));
	jand g0297(.dina(w_n598_1[0]),.dinb(w_n595_0[1]),.dout(n612),.clk(gclk));
	jand g0298(.dina(w_n603_1[0]),.dinb(w_n600_0[0]),.dout(n613),.clk(gclk));
	jand g0299(.dina(w_n613_0[2]),.dinb(w_n599_0[1]),.dout(n614),.clk(gclk));
	jor g0300(.dina(n614),.dinb(w_n612_0[1]),.dout(n615),.clk(gclk));
	jnot g0301(.din(w_n615_0[2]),.dout(n616),.clk(gclk));
	jand g0302(.dina(w_n616_0[1]),.dinb(w_dff_B_1aY1013Z9_1),.dout(n617),.clk(gclk));
	jor g0303(.dina(n617),.dinb(w_n609_0[1]),.dout(n618),.clk(gclk));
	jand g0304(.dina(w_n618_0[2]),.dinb(w_dff_B_Q8FR69JP3_1),.dout(n619),.clk(gclk));
	jnot g0305(.din(w_n619_0[2]),.dout(n620),.clk(gclk));
	jnot g0306(.din(w_n618_0[1]),.dout(n621),.clk(gclk));
	jnot g0307(.din(w_G3723_0[2]),.dout(n622),.clk(gclk));
	jand g0308(.dina(G235),.dinb(w_G18_43[1]),.dout(n623),.clk(gclk));
	jand g0309(.dina(w_dff_B_uNyvENmp2_0),.dinb(w_n355_26[1]),.dout(n624),.clk(gclk));
	jor g0310(.dina(w_n624_0[1]),.dinb(w_dff_B_A084MN4E7_1),.dout(n625),.clk(gclk));
	jxor g0311(.dina(w_n625_1[1]),.dinb(w_n622_0[2]),.dout(n626),.clk(gclk));
	jnot g0312(.din(w_G3717_0[2]),.dout(n627),.clk(gclk));
	jand g0313(.dina(G236),.dinb(w_G18_43[0]),.dout(n628),.clk(gclk));
	jand g0314(.dina(w_dff_B_qWV7iYu50_0),.dinb(w_n355_26[0]),.dout(n629),.clk(gclk));
	jor g0315(.dina(w_n629_0[1]),.dinb(w_dff_B_eSI8rUsk5_1),.dout(n630),.clk(gclk));
	jxor g0316(.dina(w_n630_0[2]),.dinb(w_n627_0[2]),.dout(n631),.clk(gclk));
	jnot g0317(.din(w_G3711_0[1]),.dout(n632),.clk(gclk));
	jand g0318(.dina(G237),.dinb(w_G18_42[2]),.dout(n633),.clk(gclk));
	jand g0319(.dina(w_dff_B_imc1wVcA6_0),.dinb(w_n355_25[2]),.dout(n634),.clk(gclk));
	jor g0320(.dina(w_n634_0[1]),.dinb(w_dff_B_C6xg2Z3Z4_1),.dout(n635),.clk(gclk));
	jxor g0321(.dina(w_n635_1[1]),.dinb(w_n632_1[1]),.dout(n636),.clk(gclk));
	jnot g0322(.din(w_G238_0[1]),.dout(n637),.clk(gclk));
	jor g0323(.dina(n637),.dinb(w_n355_25[1]),.dout(n638),.clk(gclk));
	jnot g0324(.din(w_G29_0[1]),.dout(n639),.clk(gclk));
	jor g0325(.dina(n639),.dinb(w_G18_42[1]),.dout(n640),.clk(gclk));
	jand g0326(.dina(n640),.dinb(n638),.dout(n641),.clk(gclk));
	jxor g0327(.dina(w_n641_0[2]),.dinb(w_G3705_1[2]),.dout(n642),.clk(gclk));
	jand g0328(.dina(w_n642_0[2]),.dinb(w_n359_1[0]),.dout(n643),.clk(gclk));
	jand g0329(.dina(n643),.dinb(w_n636_0[2]),.dout(n644),.clk(gclk));
	jand g0330(.dina(w_n644_0[1]),.dinb(w_n631_0[2]),.dout(n645),.clk(gclk));
	jand g0331(.dina(w_n645_0[1]),.dinb(w_n626_1[1]),.dout(n646),.clk(gclk));
	jand g0332(.dina(w_n625_1[0]),.dinb(w_n622_0[1]),.dout(n647),.clk(gclk));
	jnot g0333(.din(w_n625_0[2]),.dout(n648),.clk(gclk));
	jand g0334(.dina(n648),.dinb(w_G3723_0[1]),.dout(n649),.clk(gclk));
	jnot g0335(.din(w_n649_0[1]),.dout(n650),.clk(gclk));
	jnot g0336(.din(w_n630_0[1]),.dout(n651),.clk(gclk));
	jand g0337(.dina(w_n651_0[1]),.dinb(w_G3717_0[1]),.dout(n652),.clk(gclk));
	jnot g0338(.din(w_n652_0[1]),.dout(n653),.clk(gclk));
	jand g0339(.dina(w_n630_0[0]),.dinb(w_n627_0[1]),.dout(n654),.clk(gclk));
	jand g0340(.dina(w_n635_1[0]),.dinb(w_n632_1[0]),.dout(n655),.clk(gclk));
	jor g0341(.dina(w_n635_0[2]),.dinb(w_n632_0[2]),.dout(n656),.clk(gclk));
	jnot g0342(.din(w_G3705_1[1]),.dout(n657),.clk(gclk));
	jand g0343(.dina(w_G238_0[0]),.dinb(w_G18_42[0]),.dout(n658),.clk(gclk));
	jand g0344(.dina(w_G29_0[0]),.dinb(w_n355_25[0]),.dout(n659),.clk(gclk));
	jor g0345(.dina(w_n659_0[1]),.dinb(w_dff_B_pTaV3zpz2_1),.dout(n660),.clk(gclk));
	jor g0346(.dina(w_n660_0[2]),.dinb(w_n657_0[2]),.dout(n661),.clk(gclk));
	jnot g0347(.din(w_G3701_0[2]),.dout(n662),.clk(gclk));
	jand g0348(.dina(w_G41_0[0]),.dinb(w_n355_24[2]),.dout(n663),.clk(gclk));
	jand g0349(.dina(w_n663_1[1]),.dinb(w_n662_0[1]),.dout(n664),.clk(gclk));
	jand g0350(.dina(w_n660_0[1]),.dinb(w_n657_0[1]),.dout(n665),.clk(gclk));
	jor g0351(.dina(n665),.dinb(w_n664_0[1]),.dout(n666),.clk(gclk));
	jand g0352(.dina(w_n666_0[1]),.dinb(w_n661_0[2]),.dout(n667),.clk(gclk));
	jand g0353(.dina(n667),.dinb(w_n656_0[1]),.dout(n668),.clk(gclk));
	jor g0354(.dina(n668),.dinb(w_n655_0[1]),.dout(n669),.clk(gclk));
	jor g0355(.dina(w_n669_0[1]),.dinb(w_n654_0[2]),.dout(n670),.clk(gclk));
	jand g0356(.dina(n670),.dinb(w_n653_0[1]),.dout(n671),.clk(gclk));
	jand g0357(.dina(w_n671_0[1]),.dinb(w_dff_B_KOksx7kp3_1),.dout(n672),.clk(gclk));
	jor g0358(.dina(n672),.dinb(w_n647_0[1]),.dout(n673),.clk(gclk));
	jor g0359(.dina(w_n673_0[2]),.dinb(w_n646_0[1]),.dout(n674),.clk(gclk));
	jor g0360(.dina(w_n673_0[1]),.dinb(w_G4526_2[1]),.dout(n675),.clk(gclk));
	jand g0361(.dina(n675),.dinb(w_n674_0[1]),.dout(n676),.clk(gclk));
	jor g0362(.dina(w_n676_0[2]),.dinb(w_dff_B_arJKPxfw8_1),.dout(n677),.clk(gclk));
	jand g0363(.dina(n677),.dinb(w_dff_B_DN46X9li4_1),.dout(n678),.clk(gclk));
	jand g0364(.dina(w_n678_0[1]),.dinb(w_dff_B_VXnoGf3b7_1),.dout(n679),.clk(gclk));
	jor g0365(.dina(n679),.dinb(w_n586_0[2]),.dout(n680),.clk(gclk));
	jand g0366(.dina(w_n680_2[2]),.dinb(w_n581_0[2]),.dout(n681),.clk(gclk));
	jor g0367(.dina(n681),.dinb(w_n572_1[1]),.dout(n682),.clk(gclk));
	jand g0368(.dina(w_n682_0[1]),.dinb(w_dff_B_qToOmZvf7_1),.dout(n683),.clk(gclk));
	jand g0369(.dina(w_n683_0[1]),.dinb(w_n524_1[2]),.dout(n684),.clk(gclk));
	jand g0370(.dina(n684),.dinb(w_dff_B_pE2wBYNa4_1),.dout(n685),.clk(gclk));
	jand g0371(.dina(n685),.dinb(w_n513_1[1]),.dout(n686),.clk(gclk));
	jand g0372(.dina(w_n512_0[1]),.dinb(w_n509_0[1]),.dout(n687),.clk(gclk));
	jnot g0373(.din(w_n687_0[1]),.dout(n688),.clk(gclk));
	jnot g0374(.din(w_n512_0[0]),.dout(n689),.clk(gclk));
	jand g0375(.dina(w_n689_0[1]),.dinb(w_G4432_0[1]),.dout(n690),.clk(gclk));
	jand g0376(.dina(w_n523_0[1]),.dinb(w_n520_0[0]),.dout(n691),.clk(gclk));
	jand g0377(.dina(w_n524_1[1]),.dinb(w_n518_1[1]),.dout(n692),.clk(gclk));
	jor g0378(.dina(n692),.dinb(w_dff_B_0gubTSiJ7_1),.dout(n693),.clk(gclk));
	jnot g0379(.din(w_n693_0[1]),.dout(n694),.clk(gclk));
	jor g0380(.dina(w_n694_0[1]),.dinb(w_n690_0[1]),.dout(n695),.clk(gclk));
	jand g0381(.dina(w_n695_0[1]),.dinb(w_dff_B_2OvdcqoQ8_1),.dout(n696),.clk(gclk));
	jnot g0382(.din(w_n696_0[1]),.dout(n697),.clk(gclk));
	jor g0383(.dina(w_dff_B_pce0MwIA2_0),.dinb(n686),.dout(n698),.clk(gclk));
	jand g0384(.dina(w_n698_0[1]),.dinb(w_dff_B_ivJcWUpd4_1),.dout(n699),.clk(gclk));
	jor g0385(.dina(n699),.dinb(w_n505_0[1]),.dout(n700),.clk(gclk));
	jor g0386(.dina(w_n700_1[1]),.dinb(w_n462_0[1]),.dout(n701),.clk(gclk));
	jor g0387(.dina(n701),.dinb(w_n500_0[1]),.dout(n702),.clk(gclk));
	jand g0388(.dina(n702),.dinb(w_n499_0[1]),.dout(n703),.clk(gclk));
	jor g0389(.dina(w_n703_1[2]),.dinb(w_n449_1[0]),.dout(n704),.clk(gclk));
	jand g0390(.dina(n704),.dinb(w_n450_0[2]),.dout(n705),.clk(gclk));
	jand g0391(.dina(w_n705_0[1]),.dinb(w_n425_1[1]),.dout(n706),.clk(gclk));
	jor g0392(.dina(n706),.dinb(w_n424_0[1]),.dout(n707),.clk(gclk));
	jor g0393(.dina(w_n707_1[2]),.dinb(w_n413_1[0]),.dout(n708),.clk(gclk));
	jand g0394(.dina(n708),.dinb(w_n420_0[1]),.dout(n709),.clk(gclk));
	jand g0395(.dina(w_n709_1[1]),.dinb(w_n370_0[2]),.dout(n710),.clk(gclk));
	jand g0396(.dina(n710),.dinb(w_n363_0[2]),.dout(n711),.clk(gclk));
	jnot g0397(.din(w_n362_0[1]),.dout(n712),.clk(gclk));
	jand g0398(.dina(w_n712_0[2]),.dinb(w_G38_2[0]),.dout(n713),.clk(gclk));
	jand g0399(.dina(w_n366_0[1]),.dinb(w_G38_1[2]),.dout(n714),.clk(gclk));
	jor g0400(.dina(w_dff_B_ZQL03hyj8_0),.dinb(w_n713_0[1]),.dout(n715),.clk(gclk));
	jor g0401(.dina(w_n715_1[1]),.dinb(w_n711_1[1]),.dout(G246),.clk(gclk));
	jand g0402(.dina(w_G2204_0[2]),.dinb(w_G1455_0[2]),.dout(n717),.clk(gclk));
	jor g0403(.dina(w_dff_B_Xp7qq0Vb4_0),.dinb(w_n368_0[0]),.dout(n718),.clk(gclk));
	jor g0404(.dina(w_dff_B_LdDA1UfB9_0),.dinb(w_n355_24[1]),.dout(n719),.clk(gclk));
	jand g0405(.dina(w_n719_0[1]),.dinb(w_n373_6[1]),.dout(n720),.clk(gclk));
	jor g0406(.dina(w_n371_0[0]),.dinb(w_n355_24[0]),.dout(n721),.clk(gclk));
	jor g0407(.dina(G88),.dinb(w_G18_41[2]),.dout(n722),.clk(gclk));
	jand g0408(.dina(w_dff_B_suekqKZF4_0),.dinb(n721),.dout(n723),.clk(gclk));
	jxor g0409(.dina(w_n723_0[2]),.dinb(w_n720_0[2]),.dout(n724),.clk(gclk));
	jor g0410(.dina(w_dff_B_X6BYXpZV8_0),.dinb(w_n355_23[2]),.dout(n725),.clk(gclk));
	jand g0411(.dina(w_n725_0[1]),.dinb(w_n373_6[0]),.dout(n726),.clk(gclk));
	jor g0412(.dina(w_n383_0[0]),.dinb(w_n355_23[1]),.dout(n727),.clk(gclk));
	jor g0413(.dina(G112),.dinb(w_G18_41[1]),.dout(n728),.clk(gclk));
	jand g0414(.dina(w_dff_B_PknzMfj32_0),.dinb(n727),.dout(n729),.clk(gclk));
	jor g0415(.dina(w_n729_1[1]),.dinb(w_n726_1[1]),.dout(n730),.clk(gclk));
	jand g0416(.dina(w_n729_1[0]),.dinb(w_n726_1[0]),.dout(n731),.clk(gclk));
	jor g0417(.dina(w_n389_0[2]),.dinb(w_n355_23[0]),.dout(n732),.clk(gclk));
	jor g0418(.dina(G113),.dinb(w_G18_41[0]),.dout(n733),.clk(gclk));
	jand g0419(.dina(w_dff_B_U8wghQvY4_0),.dinb(n732),.dout(n734),.clk(gclk));
	jand g0420(.dina(w_n734_0[2]),.dinb(w_n373_5[2]),.dout(n735),.clk(gclk));
	jor g0421(.dina(w_dff_B_IC7aNWb99_0),.dinb(w_n355_22[2]),.dout(n736),.clk(gclk));
	jand g0422(.dina(w_n736_0[1]),.dinb(w_n373_5[1]),.dout(n737),.clk(gclk));
	jand g0423(.dina(w_G106_0[2]),.dinb(w_G18_40[2]),.dout(n738),.clk(gclk));
	jnot g0424(.din(n738),.dout(n739),.clk(gclk));
	jor g0425(.dina(G87),.dinb(w_G18_40[1]),.dout(n740),.clk(gclk));
	jand g0426(.dina(w_dff_B_oVCXBg7B5_0),.dinb(n739),.dout(n741),.clk(gclk));
	jxor g0427(.dina(w_n741_1[1]),.dinb(w_n737_1[1]),.dout(n742),.clk(gclk));
	jor g0428(.dina(w_dff_B_q4LyJ9mr1_0),.dinb(w_n355_22[1]),.dout(n743),.clk(gclk));
	jand g0429(.dina(w_n743_0[1]),.dinb(w_n373_5[0]),.dout(n744),.clk(gclk));
	jor g0430(.dina(w_n393_0[2]),.dinb(w_n355_22[0]),.dout(n745),.clk(gclk));
	jor g0431(.dina(G111),.dinb(w_G18_40[0]),.dout(n746),.clk(gclk));
	jand g0432(.dina(w_dff_B_KVIsyAul7_0),.dinb(n745),.dout(n747),.clk(gclk));
	jxor g0433(.dina(w_n747_0[2]),.dinb(w_n744_0[2]),.dout(n748),.clk(gclk));
	jand g0434(.dina(n748),.dinb(n742),.dout(n749),.clk(gclk));
	jand g0435(.dina(w_n749_0[1]),.dinb(w_dff_B_XLCg4Vxz6_1),.dout(n750),.clk(gclk));
	jor g0436(.dina(n750),.dinb(w_dff_B_m7N8lvTH8_1),.dout(n751),.clk(gclk));
	jand g0437(.dina(n751),.dinb(w_dff_B_TSRR2EAS2_1),.dout(n752),.clk(gclk));
	jand g0438(.dina(n752),.dinb(w_n724_0[1]),.dout(n753),.clk(gclk));
	jor g0439(.dina(w_dff_B_rilexsIN7_0),.dinb(w_n355_21[2]),.dout(n754),.clk(gclk));
	jand g0440(.dina(w_n754_0[1]),.dinb(w_n373_4[2]),.dout(n755),.clk(gclk));
	jor g0441(.dina(w_n421_0[0]),.dinb(w_n355_21[1]),.dout(n756),.clk(gclk));
	jor g0442(.dina(G110),.dinb(w_G18_39[2]),.dout(n757),.clk(gclk));
	jand g0443(.dina(w_dff_B_hZpeGKhD7_0),.dinb(n756),.dout(n758),.clk(gclk));
	jxor g0444(.dina(w_n758_1[1]),.dinb(w_n755_1[1]),.dout(n759),.clk(gclk));
	jor g0445(.dina(w_dff_B_xlnYYd9P9_0),.dinb(w_n355_21[0]),.dout(n760),.clk(gclk));
	jand g0446(.dina(w_n760_0[1]),.dinb(w_n373_4[1]),.dout(n761),.clk(gclk));
	jor g0447(.dina(w_n426_0[0]),.dinb(w_n355_20[2]),.dout(n762),.clk(gclk));
	jor g0448(.dina(G109),.dinb(w_G18_39[1]),.dout(n763),.clk(gclk));
	jand g0449(.dina(w_dff_B_6S4NPvSl2_0),.dinb(n762),.dout(n764),.clk(gclk));
	jxor g0450(.dina(w_n764_0[2]),.dinb(w_n761_0[2]),.dout(n765),.clk(gclk));
	jand g0451(.dina(n765),.dinb(n759),.dout(n766),.clk(gclk));
	jor g0452(.dina(w_dff_B_lVJBxmwj6_0),.dinb(w_n355_20[1]),.dout(n767),.clk(gclk));
	jand g0453(.dina(w_n767_0[1]),.dinb(w_n373_4[0]),.dout(n768),.clk(gclk));
	jand g0454(.dina(w_G2247_0[1]),.dinb(w_G18_39[0]),.dout(n769),.clk(gclk));
	jnot g0455(.din(n769),.dout(n770),.clk(gclk));
	jor g0456(.dina(G86),.dinb(w_G18_38[2]),.dout(n771),.clk(gclk));
	jand g0457(.dina(w_dff_B_rZiy9hkI1_0),.dinb(n770),.dout(n772),.clk(gclk));
	jand g0458(.dina(w_n772_0[2]),.dinb(w_n768_0[2]),.dout(n773),.clk(gclk));
	jor g0459(.dina(w_n772_0[1]),.dinb(w_n768_0[1]),.dout(n774),.clk(gclk));
	jor g0460(.dina(w_dff_B_ACptuE0V4_0),.dinb(w_n355_20[0]),.dout(n775),.clk(gclk));
	jand g0461(.dina(w_n775_0[1]),.dinb(w_n373_3[2]),.dout(n776),.clk(gclk));
	jand g0462(.dina(w_G2239_1[0]),.dinb(w_G18_38[1]),.dout(n777),.clk(gclk));
	jnot g0463(.din(n777),.dout(n778),.clk(gclk));
	jor g0464(.dina(G63),.dinb(w_G18_38[0]),.dout(n779),.clk(gclk));
	jand g0465(.dina(w_dff_B_MevoUuZj5_0),.dinb(n778),.dout(n780),.clk(gclk));
	jand g0466(.dina(w_n780_0[2]),.dinb(w_n776_0[2]),.dout(n781),.clk(gclk));
	jand g0467(.dina(w_n781_0[1]),.dinb(w_n774_0[1]),.dout(n782),.clk(gclk));
	jor g0468(.dina(n782),.dinb(w_n773_0[1]),.dout(n783),.clk(gclk));
	jand g0469(.dina(n783),.dinb(w_n766_0[1]),.dout(n784),.clk(gclk));
	jand g0470(.dina(w_n758_1[0]),.dinb(w_n755_1[0]),.dout(n785),.clk(gclk));
	jor g0471(.dina(w_n758_0[2]),.dinb(w_n755_0[2]),.dout(n786),.clk(gclk));
	jand g0472(.dina(w_n764_0[1]),.dinb(w_n761_0[1]),.dout(n787),.clk(gclk));
	jand g0473(.dina(n787),.dinb(n786),.dout(n788),.clk(gclk));
	jor g0474(.dina(n788),.dinb(w_dff_B_AysCa2sL2_1),.dout(n789),.clk(gclk));
	jor g0475(.dina(w_dff_B_7UnKPXbe2_0),.dinb(n784),.dout(n790),.clk(gclk));
	jnot g0476(.din(w_n773_0[0]),.dout(n791),.clk(gclk));
	jnot g0477(.din(w_n781_0[0]),.dout(n792),.clk(gclk));
	jand g0478(.dina(n792),.dinb(n791),.dout(n793),.clk(gclk));
	jand g0479(.dina(n793),.dinb(w_n766_0[0]),.dout(n794),.clk(gclk));
	jor g0480(.dina(w_dff_B_neYfZjv58_0),.dinb(w_n355_19[2]),.dout(n795),.clk(gclk));
	jand g0481(.dina(n795),.dinb(w_n373_3[1]),.dout(n796),.clk(gclk));
	jand g0482(.dina(w_G2236_0[1]),.dinb(w_G18_37[2]),.dout(n797),.clk(gclk));
	jnot g0483(.din(n797),.dout(n798),.clk(gclk));
	jor g0484(.dina(G64),.dinb(w_G18_37[1]),.dout(n799),.clk(gclk));
	jand g0485(.dina(w_dff_B_Q1fKgDge9_0),.dinb(n798),.dout(n800),.clk(gclk));
	jxor g0486(.dina(w_n800_1[1]),.dinb(w_n796_1[1]),.dout(n801),.clk(gclk));
	jand g0487(.dina(G178),.dinb(w_G18_37[0]),.dout(n802),.clk(gclk));
	jor g0488(.dina(w_dff_B_8afCptDr6_0),.dinb(w_n457_0[0]),.dout(n803),.clk(gclk));
	jor g0489(.dina(w_n456_0[0]),.dinb(w_n355_19[1]),.dout(n804),.clk(gclk));
	jor g0490(.dina(G85),.dinb(w_G18_36[2]),.dout(n805),.clk(gclk));
	jand g0491(.dina(w_dff_B_IHKWq1ZS2_0),.dinb(n804),.dout(n806),.clk(gclk));
	jxor g0492(.dina(w_n806_0[2]),.dinb(w_n803_0[2]),.dout(n807),.clk(gclk));
	jand g0493(.dina(n807),.dinb(n801),.dout(n808),.clk(gclk));
	jand g0494(.dina(G179),.dinb(w_G18_36[1]),.dout(n809),.clk(gclk));
	jor g0495(.dina(w_dff_B_HI17SWLs1_0),.dinb(w_n467_0[0]),.dout(n810),.clk(gclk));
	jand g0496(.dina(w_G2224_0[2]),.dinb(w_G18_36[0]),.dout(n811),.clk(gclk));
	jnot g0497(.din(n811),.dout(n812),.clk(gclk));
	jor g0498(.dina(G84),.dinb(w_G18_35[2]),.dout(n813),.clk(gclk));
	jand g0499(.dina(w_dff_B_aJMHWVVK0_0),.dinb(n812),.dout(n814),.clk(gclk));
	jxor g0500(.dina(w_n814_1[1]),.dinb(w_n810_1[1]),.dout(n815),.clk(gclk));
	jand g0501(.dina(G180),.dinb(w_G18_35[1]),.dout(n816),.clk(gclk));
	jor g0502(.dina(w_dff_B_VCPo7aj54_0),.dinb(w_n472_0[0]),.dout(n817),.clk(gclk));
	jor g0503(.dina(w_n471_0[0]),.dinb(w_n355_19[0]),.dout(n818),.clk(gclk));
	jor g0504(.dina(G83),.dinb(w_G18_35[0]),.dout(n819),.clk(gclk));
	jand g0505(.dina(w_dff_B_LlYTllIS2_0),.dinb(n818),.dout(n820),.clk(gclk));
	jxor g0506(.dina(w_n820_0[2]),.dinb(w_n817_0[2]),.dout(n821),.clk(gclk));
	jand g0507(.dina(n821),.dinb(n815),.dout(n822),.clk(gclk));
	jand g0508(.dina(G171),.dinb(w_G18_34[2]),.dout(n823),.clk(gclk));
	jor g0509(.dina(w_dff_B_XobirX4R6_0),.dinb(w_n477_0[0]),.dout(n824),.clk(gclk));
	jor g0510(.dina(w_n476_0[0]),.dinb(w_n355_18[2]),.dout(n825),.clk(gclk));
	jor g0511(.dina(G65),.dinb(w_G18_34[1]),.dout(n826),.clk(gclk));
	jand g0512(.dina(w_dff_B_NXZo4Vpb7_0),.dinb(n825),.dout(n827),.clk(gclk));
	jand g0513(.dina(w_n827_0[2]),.dinb(w_n824_0[2]),.dout(n828),.clk(gclk));
	jand g0514(.dina(w_dff_B_PkOzYPwq0_0),.dinb(w_n822_0[1]),.dout(n829),.clk(gclk));
	jand g0515(.dina(w_n814_1[0]),.dinb(w_n810_1[0]),.dout(n830),.clk(gclk));
	jor g0516(.dina(w_n814_0[2]),.dinb(w_n810_0[2]),.dout(n831),.clk(gclk));
	jand g0517(.dina(w_n820_0[1]),.dinb(w_n817_0[1]),.dout(n832),.clk(gclk));
	jand g0518(.dina(n832),.dinb(n831),.dout(n833),.clk(gclk));
	jor g0519(.dina(n833),.dinb(w_dff_B_fNbtVY718_1),.dout(n834),.clk(gclk));
	jor g0520(.dina(n834),.dinb(n829),.dout(n835),.clk(gclk));
	jand g0521(.dina(n835),.dinb(w_n808_0[1]),.dout(n836),.clk(gclk));
	jand g0522(.dina(w_n800_1[0]),.dinb(w_n796_1[0]),.dout(n837),.clk(gclk));
	jor g0523(.dina(w_n800_0[2]),.dinb(w_n796_0[2]),.dout(n838),.clk(gclk));
	jand g0524(.dina(w_n806_0[1]),.dinb(w_n803_0[1]),.dout(n839),.clk(gclk));
	jand g0525(.dina(n839),.dinb(n838),.dout(n840),.clk(gclk));
	jor g0526(.dina(n840),.dinb(w_dff_B_ZkmYrJx73_1),.dout(n841),.clk(gclk));
	jor g0527(.dina(w_dff_B_RuudyVQP2_0),.dinb(n836),.dout(n842),.clk(gclk));
	jand g0528(.dina(w_n822_0[0]),.dinb(w_n808_0[0]),.dout(n843),.clk(gclk));
	jand g0529(.dina(G189),.dinb(w_G18_34[0]),.dout(n844),.clk(gclk));
	jor g0530(.dina(w_dff_B_mTocefGd9_0),.dinb(w_n503_0[0]),.dout(n845),.clk(gclk));
	jor g0531(.dina(w_n501_0[1]),.dinb(w_n355_18[1]),.dout(n846),.clk(gclk));
	jor g0532(.dina(G62),.dinb(w_G18_33[2]),.dout(n847),.clk(gclk));
	jand g0533(.dina(w_dff_B_bTJoSfQD1_0),.dinb(n846),.dout(n848),.clk(gclk));
	jxor g0534(.dina(w_n848_1[1]),.dinb(w_n845_1[1]),.dout(n849),.clk(gclk));
	jand g0535(.dina(G190),.dinb(w_G18_33[1]),.dout(n850),.clk(gclk));
	jor g0536(.dina(w_dff_B_mVGGaIz23_0),.dinb(w_n511_0[0]),.dout(n851),.clk(gclk));
	jor g0537(.dina(w_n509_0[0]),.dinb(w_n355_18[0]),.dout(n852),.clk(gclk));
	jor g0538(.dina(G61),.dinb(w_G18_33[0]),.dout(n853),.clk(gclk));
	jand g0539(.dina(w_dff_B_VMN7qhTg7_0),.dinb(n852),.dout(n854),.clk(gclk));
	jxor g0540(.dina(w_n854_0[2]),.dinb(w_n851_0[2]),.dout(n855),.clk(gclk));
	jand g0541(.dina(n855),.dinb(n849),.dout(n856),.clk(gclk));
	jand g0542(.dina(G191),.dinb(w_G18_32[2]),.dout(n857),.clk(gclk));
	jor g0543(.dina(w_dff_B_fV89OfNc8_0),.dinb(w_n522_0[0]),.dout(n858),.clk(gclk));
	jand g0544(.dina(w_G4427_0[1]),.dinb(w_G18_32[1]),.dout(n859),.clk(gclk));
	jnot g0545(.din(n859),.dout(n860),.clk(gclk));
	jor g0546(.dina(G60),.dinb(w_G18_32[0]),.dout(n861),.clk(gclk));
	jand g0547(.dina(w_dff_B_sQF7XcW14_0),.dinb(n860),.dout(n862),.clk(gclk));
	jand g0548(.dina(w_n862_0[2]),.dinb(w_n858_0[2]),.dout(n863),.clk(gclk));
	jor g0549(.dina(w_n862_0[1]),.dinb(w_n858_0[1]),.dout(n864),.clk(gclk));
	jand g0550(.dina(G192),.dinb(w_G18_31[2]),.dout(n865),.clk(gclk));
	jor g0551(.dina(w_dff_B_dnkm3fBP6_0),.dinb(w_n516_0[0]),.dout(n866),.clk(gclk));
	jand g0552(.dina(w_G4420_0[2]),.dinb(w_G18_31[1]),.dout(n867),.clk(gclk));
	jnot g0553(.din(n867),.dout(n868),.clk(gclk));
	jor g0554(.dina(G79),.dinb(w_G18_31[0]),.dout(n869),.clk(gclk));
	jand g0555(.dina(w_dff_B_i1Wnk4No1_0),.dinb(n868),.dout(n870),.clk(gclk));
	jand g0556(.dina(w_n870_0[2]),.dinb(w_n866_0[2]),.dout(n871),.clk(gclk));
	jand g0557(.dina(w_n871_0[1]),.dinb(w_n864_0[1]),.dout(n872),.clk(gclk));
	jor g0558(.dina(n872),.dinb(w_n863_0[1]),.dout(n873),.clk(gclk));
	jand g0559(.dina(n873),.dinb(w_n856_0[1]),.dout(n874),.clk(gclk));
	jand g0560(.dina(w_n848_1[0]),.dinb(w_n845_1[0]),.dout(n875),.clk(gclk));
	jor g0561(.dina(w_n848_0[2]),.dinb(w_n845_0[2]),.dout(n876),.clk(gclk));
	jand g0562(.dina(w_n854_0[1]),.dinb(w_n851_0[1]),.dout(n877),.clk(gclk));
	jand g0563(.dina(n877),.dinb(n876),.dout(n878),.clk(gclk));
	jor g0564(.dina(n878),.dinb(w_dff_B_R2ssDfRx2_1),.dout(n879),.clk(gclk));
	jor g0565(.dina(w_dff_B_xCGAEQP75_0),.dinb(n874),.dout(n880),.clk(gclk));
	jor g0566(.dina(w_n870_0[1]),.dinb(w_n866_0[1]),.dout(n881),.clk(gclk));
	jand g0567(.dina(n881),.dinb(w_n864_0[0]),.dout(n882),.clk(gclk));
	jand g0568(.dina(n882),.dinb(w_n856_0[0]),.dout(n883),.clk(gclk));
	jand g0569(.dina(G205),.dinb(w_G18_30[2]),.dout(n884),.clk(gclk));
	jor g0570(.dina(w_dff_B_9SokRwpu0_0),.dinb(w_n629_0[0]),.dout(n885),.clk(gclk));
	jor g0571(.dina(w_n627_0[0]),.dinb(w_n355_17[2]),.dout(n886),.clk(gclk));
	jor g0572(.dina(G75),.dinb(w_G18_30[1]),.dout(n887),.clk(gclk));
	jand g0573(.dina(w_dff_B_LTj0zE0V5_0),.dinb(n886),.dout(n888),.clk(gclk));
	jor g0574(.dina(w_n888_0[2]),.dinb(w_n885_0[2]),.dout(n889),.clk(gclk));
	jand g0575(.dina(G206),.dinb(w_G18_30[0]),.dout(n890),.clk(gclk));
	jor g0576(.dina(w_dff_B_MxQHdMvy2_0),.dinb(w_n634_0[0]),.dout(n891),.clk(gclk));
	jor g0577(.dina(w_n632_0[1]),.dinb(w_n355_17[1]),.dout(n892),.clk(gclk));
	jor g0578(.dina(G76),.dinb(w_G18_29[2]),.dout(n893),.clk(gclk));
	jand g0579(.dina(w_dff_B_bEl0xenY5_0),.dinb(n892),.dout(n894),.clk(gclk));
	jand g0580(.dina(w_n894_0[2]),.dinb(w_n891_0[2]),.dout(n895),.clk(gclk));
	jor g0581(.dina(w_G89_0[1]),.dinb(w_G70_0[1]),.dout(n896),.clk(gclk));
	jand g0582(.dina(w_dff_B_BNFVeHPN2_0),.dinb(w_n663_1[0]),.dout(n897),.clk(gclk));
	jor g0583(.dina(w_dff_B_RnXkE3it4_0),.dinb(w_n895_0[1]),.dout(n898),.clk(gclk));
	jand g0584(.dina(G207),.dinb(w_G18_29[1]),.dout(n899),.clk(gclk));
	jor g0585(.dina(w_dff_B_bxk0bZM88_0),.dinb(w_n659_0[0]),.dout(n900),.clk(gclk));
	jor g0586(.dina(w_n657_0[0]),.dinb(w_n355_17[0]),.dout(n901),.clk(gclk));
	jor g0587(.dina(G74),.dinb(w_G18_29[0]),.dout(n902),.clk(gclk));
	jand g0588(.dina(w_dff_B_6S7kVID85_0),.dinb(n901),.dout(n903),.clk(gclk));
	jand g0589(.dina(w_n903_0[2]),.dinb(w_n900_0[2]),.dout(n904),.clk(gclk));
	jor g0590(.dina(w_G70_0[0]),.dinb(w_G18_28[2]),.dout(n905),.clk(gclk));
	jand g0591(.dina(w_n905_0[1]),.dinb(w_G89_0[0]),.dout(n906),.clk(gclk));
	jor g0592(.dina(w_dff_B_1SRk8rnZ7_0),.dinb(n904),.dout(n907),.clk(gclk));
	jor g0593(.dina(n907),.dinb(n898),.dout(n908),.clk(gclk));
	jor g0594(.dina(w_n903_0[1]),.dinb(w_n900_0[1]),.dout(n909),.clk(gclk));
	jor g0595(.dina(w_n894_0[1]),.dinb(w_n891_0[1]),.dout(n910),.clk(gclk));
	jand g0596(.dina(n910),.dinb(n909),.dout(n911),.clk(gclk));
	jor g0597(.dina(n911),.dinb(w_n895_0[0]),.dout(n912),.clk(gclk));
	jand g0598(.dina(n912),.dinb(n908),.dout(n913),.clk(gclk));
	jand g0599(.dina(n913),.dinb(w_dff_B_ZauRDTiH8_1),.dout(n914),.clk(gclk));
	jand g0600(.dina(G204),.dinb(w_G18_28[1]),.dout(n915),.clk(gclk));
	jor g0601(.dina(w_dff_B_ZKWIEJTp2_0),.dinb(w_n624_0[0]),.dout(n916),.clk(gclk));
	jor g0602(.dina(w_n622_0[0]),.dinb(w_n355_16[2]),.dout(n917),.clk(gclk));
	jor g0603(.dina(G73),.dinb(w_G18_28[0]),.dout(n918),.clk(gclk));
	jand g0604(.dina(w_dff_B_erXJUqiE4_0),.dinb(n917),.dout(n919),.clk(gclk));
	jand g0605(.dina(w_n919_0[2]),.dinb(w_n916_0[2]),.dout(n920),.clk(gclk));
	jand g0606(.dina(w_n888_0[1]),.dinb(w_n885_0[1]),.dout(n921),.clk(gclk));
	jor g0607(.dina(n921),.dinb(n920),.dout(n922),.clk(gclk));
	jor g0608(.dina(w_dff_B_nggOTCOy9_0),.dinb(n914),.dout(n923),.clk(gclk));
	jor g0609(.dina(w_n919_0[1]),.dinb(w_n916_0[1]),.dout(n924),.clk(gclk));
	jand g0610(.dina(G203),.dinb(w_G18_27[2]),.dout(n925),.clk(gclk));
	jor g0611(.dina(w_dff_B_4s9IArk87_0),.dinb(w_n602_0[0]),.dout(n926),.clk(gclk));
	jand g0612(.dina(w_G3729_1[0]),.dinb(w_G18_27[1]),.dout(n927),.clk(gclk));
	jnot g0613(.din(n927),.dout(n928),.clk(gclk));
	jor g0614(.dina(G53),.dinb(w_G18_27[0]),.dout(n929),.clk(gclk));
	jand g0615(.dina(w_dff_B_GVGkWjOU8_0),.dinb(n928),.dout(n930),.clk(gclk));
	jor g0616(.dina(w_n930_0[2]),.dinb(w_n926_0[2]),.dout(n931),.clk(gclk));
	jand g0617(.dina(n931),.dinb(n924),.dout(n932),.clk(gclk));
	jand g0618(.dina(w_dff_B_k180PTCX8_0),.dinb(n923),.dout(n933),.clk(gclk));
	jand g0619(.dina(G202),.dinb(w_G18_26[2]),.dout(n934),.clk(gclk));
	jor g0620(.dina(w_dff_B_q9i22s8O9_0),.dinb(w_n597_0[0]),.dout(n935),.clk(gclk));
	jor g0621(.dina(w_n595_0[0]),.dinb(w_n355_16[1]),.dout(n936),.clk(gclk));
	jor g0622(.dina(G54),.dinb(w_G18_26[1]),.dout(n937),.clk(gclk));
	jand g0623(.dina(w_dff_B_DjGqyaxc6_0),.dinb(n936),.dout(n938),.clk(gclk));
	jand g0624(.dina(w_n938_0[2]),.dinb(w_n935_0[2]),.dout(n939),.clk(gclk));
	jand g0625(.dina(w_n930_0[1]),.dinb(w_n926_0[1]),.dout(n940),.clk(gclk));
	jor g0626(.dina(n940),.dinb(n939),.dout(n941),.clk(gclk));
	jor g0627(.dina(w_dff_B_BppfZCnu1_0),.dinb(n933),.dout(n942),.clk(gclk));
	jand g0628(.dina(G201),.dinb(w_G18_26[0]),.dout(n943),.clk(gclk));
	jor g0629(.dina(w_dff_B_tC5oChiN6_0),.dinb(w_n592_0[0]),.dout(n944),.clk(gclk));
	jor g0630(.dina(w_n590_0[0]),.dinb(w_n355_16[0]),.dout(n945),.clk(gclk));
	jor g0631(.dina(G55),.dinb(w_G18_25[2]),.dout(n946),.clk(gclk));
	jand g0632(.dina(w_dff_B_kX1qkxWd0_0),.dinb(n945),.dout(n947),.clk(gclk));
	jxor g0633(.dina(w_n947_0[2]),.dinb(w_n944_0[2]),.dout(n948),.clk(gclk));
	jand g0634(.dina(G200),.dinb(w_G18_25[1]),.dout(n949),.clk(gclk));
	jor g0635(.dina(w_dff_B_4nTjbmam1_0),.dinb(w_n584_0[0]),.dout(n950),.clk(gclk));
	jor g0636(.dina(w_n582_0[1]),.dinb(w_n355_15[2]),.dout(n951),.clk(gclk));
	jor g0637(.dina(G56),.dinb(w_G18_25[0]),.dout(n952),.clk(gclk));
	jand g0638(.dina(w_dff_B_K8YkDxMJ7_0),.dinb(n951),.dout(n953),.clk(gclk));
	jxor g0639(.dina(w_n953_1[1]),.dinb(w_n950_1[1]),.dout(n954),.clk(gclk));
	jand g0640(.dina(n954),.dinb(n948),.dout(n955),.clk(gclk));
	jor g0641(.dina(w_n938_0[1]),.dinb(w_n935_0[1]),.dout(n956),.clk(gclk));
	jand g0642(.dina(w_dff_B_estVN0us2_0),.dinb(n955),.dout(n957),.clk(gclk));
	jand g0643(.dina(w_dff_B_3bJApQEN4_0),.dinb(n942),.dout(n958),.clk(gclk));
	jand g0644(.dina(w_n953_1[0]),.dinb(w_n950_1[0]),.dout(n959),.clk(gclk));
	jand g0645(.dina(w_n947_0[1]),.dinb(w_n944_0[1]),.dout(n960),.clk(gclk));
	jor g0646(.dina(w_n953_0[2]),.dinb(w_n950_0[2]),.dout(n961),.clk(gclk));
	jand g0647(.dina(n961),.dinb(n960),.dout(n962),.clk(gclk));
	jor g0648(.dina(n962),.dinb(w_dff_B_orv1wjnb3_1),.dout(n963),.clk(gclk));
	jor g0649(.dina(w_dff_B_uZ9L45DT7_0),.dinb(n958),.dout(n964),.clk(gclk));
	jand g0650(.dina(G187),.dinb(w_G18_24[2]),.dout(n965),.clk(gclk));
	jor g0651(.dina(w_dff_B_fT6cpS2r5_0),.dinb(w_n562_0[0]),.dout(n966),.clk(gclk));
	jand g0652(.dina(w_G4394_1[0]),.dinb(w_G18_24[1]),.dout(n967),.clk(gclk));
	jnot g0653(.din(n967),.dout(n968),.clk(gclk));
	jor g0654(.dina(G77),.dinb(w_G18_24[0]),.dout(n969),.clk(gclk));
	jand g0655(.dina(w_dff_B_8rIQAGib9_0),.dinb(n968),.dout(n970),.clk(gclk));
	jor g0656(.dina(w_n970_0[2]),.dinb(w_n966_0[2]),.dout(n971),.clk(gclk));
	jand g0657(.dina(G193),.dinb(w_G18_23[2]),.dout(n972),.clk(gclk));
	jor g0658(.dina(w_dff_B_fFR3xlQT2_0),.dinb(w_n530_0[0]),.dout(n973),.clk(gclk));
	jand g0659(.dina(w_G4415_0[2]),.dinb(w_G18_23[1]),.dout(n974),.clk(gclk));
	jnot g0660(.din(n974),.dout(n975),.clk(gclk));
	jor g0661(.dina(G80),.dinb(w_G18_23[0]),.dout(n976),.clk(gclk));
	jand g0662(.dina(w_dff_B_l3G4sekk1_0),.dinb(n975),.dout(n977),.clk(gclk));
	jxor g0663(.dina(w_n977_1[1]),.dinb(w_n973_1[1]),.dout(n978),.clk(gclk));
	jand g0664(.dina(G194),.dinb(w_G18_22[2]),.dout(n979),.clk(gclk));
	jor g0665(.dina(w_dff_B_NfZNRfxe8_0),.dinb(w_n538_0[0]),.dout(n980),.clk(gclk));
	jor g0666(.dina(w_n536_0[0]),.dinb(w_n355_15[1]),.dout(n981),.clk(gclk));
	jor g0667(.dina(G81),.dinb(w_G18_22[1]),.dout(n982),.clk(gclk));
	jand g0668(.dina(w_dff_B_UQfx4r7m6_0),.dinb(n981),.dout(n983),.clk(gclk));
	jxor g0669(.dina(w_n983_0[2]),.dinb(w_n980_0[2]),.dout(n984),.clk(gclk));
	jand g0670(.dina(n984),.dinb(n978),.dout(n985),.clk(gclk));
	jand g0671(.dina(G196),.dinb(w_G18_22[0]),.dout(n986),.clk(gclk));
	jor g0672(.dina(w_dff_B_cQLPEVoP8_0),.dinb(w_n554_0[0]),.dout(n987),.clk(gclk));
	jand g0673(.dina(w_G4400_0[2]),.dinb(w_G18_21[2]),.dout(n988),.clk(gclk));
	jnot g0674(.din(n988),.dout(n989),.clk(gclk));
	jor g0675(.dina(G78),.dinb(w_G18_21[1]),.dout(n990),.clk(gclk));
	jand g0676(.dina(w_dff_B_lmDZK8E89_0),.dinb(n989),.dout(n991),.clk(gclk));
	jand g0677(.dina(w_n991_0[2]),.dinb(w_n987_0[2]),.dout(n992),.clk(gclk));
	jnot g0678(.din(w_n992_0[1]),.dout(n993),.clk(gclk));
	jand g0679(.dina(G195),.dinb(w_G18_21[0]),.dout(n994),.clk(gclk));
	jor g0680(.dina(w_dff_B_XXe0m7kV4_0),.dinb(w_n546_0[0]),.dout(n995),.clk(gclk));
	jand g0681(.dina(w_G4405_0[2]),.dinb(w_G18_20[2]),.dout(n996),.clk(gclk));
	jnot g0682(.din(n996),.dout(n997),.clk(gclk));
	jor g0683(.dina(G59),.dinb(w_G18_20[1]),.dout(n998),.clk(gclk));
	jand g0684(.dina(w_dff_B_hIfhACI74_0),.dinb(n997),.dout(n999),.clk(gclk));
	jor g0685(.dina(w_n999_0[2]),.dinb(w_n995_0[2]),.dout(n1000),.clk(gclk));
	jand g0686(.dina(w_n1000_0[1]),.dinb(n993),.dout(n1001),.clk(gclk));
	jor g0687(.dina(w_n991_0[1]),.dinb(w_n987_0[1]),.dout(n1002),.clk(gclk));
	jand g0688(.dina(w_n999_0[1]),.dinb(w_n995_0[1]),.dout(n1003),.clk(gclk));
	jnot g0689(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jand g0690(.dina(n1004),.dinb(w_dff_B_Ah2aUiDQ3_1),.dout(n1005),.clk(gclk));
	jand g0691(.dina(n1005),.dinb(n1001),.dout(n1006),.clk(gclk));
	jand g0692(.dina(n1006),.dinb(w_n985_0[1]),.dout(n1007),.clk(gclk));
	jand g0693(.dina(w_n970_0[1]),.dinb(w_n966_0[1]),.dout(n1008),.clk(gclk));
	jnot g0694(.din(w_n1008_0[1]),.dout(n1009),.clk(gclk));
	jand g0695(.dina(w_dff_B_HgrYxgY77_0),.dinb(w_n1007_0[1]),.dout(n1010),.clk(gclk));
	jand g0696(.dina(n1010),.dinb(w_dff_B_iSDLFJwX9_1),.dout(n1011),.clk(gclk));
	jand g0697(.dina(w_dff_B_4bXAa7Qs8_0),.dinb(n964),.dout(n1012),.clk(gclk));
	jand g0698(.dina(w_n977_1[0]),.dinb(w_n973_1[0]),.dout(n1013),.clk(gclk));
	jor g0699(.dina(w_n977_0[2]),.dinb(w_n973_0[2]),.dout(n1014),.clk(gclk));
	jand g0700(.dina(w_n983_0[1]),.dinb(w_n980_0[1]),.dout(n1015),.clk(gclk));
	jand g0701(.dina(n1015),.dinb(n1014),.dout(n1016),.clk(gclk));
	jor g0702(.dina(n1016),.dinb(w_dff_B_bLFA0pqD5_1),.dout(n1017),.clk(gclk));
	jand g0703(.dina(w_n1008_0[0]),.dinb(w_n1007_0[0]),.dout(n1018),.clk(gclk));
	jand g0704(.dina(w_n1000_0[0]),.dinb(w_n992_0[0]),.dout(n1019),.clk(gclk));
	jor g0705(.dina(n1019),.dinb(w_n1003_0[0]),.dout(n1020),.clk(gclk));
	jand g0706(.dina(n1020),.dinb(w_n985_0[0]),.dout(n1021),.clk(gclk));
	jor g0707(.dina(w_dff_B_fKc0yDPw9_0),.dinb(n1018),.dout(n1022),.clk(gclk));
	jor g0708(.dina(n1022),.dinb(w_dff_B_jorYkMEJ4_1),.dout(n1023),.clk(gclk));
	jor g0709(.dina(w_dff_B_JQsr2JeB4_0),.dinb(n1012),.dout(n1024),.clk(gclk));
	jnot g0710(.din(w_n863_0[0]),.dout(n1025),.clk(gclk));
	jnot g0711(.din(w_n871_0[0]),.dout(n1026),.clk(gclk));
	jand g0712(.dina(n1026),.dinb(n1025),.dout(n1027),.clk(gclk));
	jand g0713(.dina(w_dff_B_23Ep1ycX0_0),.dinb(n1024),.dout(n1028),.clk(gclk));
	jand g0714(.dina(n1028),.dinb(w_dff_B_hoqQbiCM6_1),.dout(n1029),.clk(gclk));
	jor g0715(.dina(n1029),.dinb(w_dff_B_lx5nZqAc0_1),.dout(G252_fa_),.clk(gclk));
	jxor g0716(.dina(w_n827_0[1]),.dinb(w_n824_0[1]),.dout(n1031),.clk(gclk));
	jand g0717(.dina(w_dff_B_cuMzDEww9_0),.dinb(w_G252_0),.dout(n1032),.clk(gclk));
	jand g0718(.dina(n1032),.dinb(w_dff_B_6ZZMi8gg9_1),.dout(n1033),.clk(gclk));
	jor g0719(.dina(n1033),.dinb(w_dff_B_jilyhg740_1),.dout(n1034),.clk(gclk));
	jor g0720(.dina(w_n780_0[1]),.dinb(w_n776_0[1]),.dout(n1035),.clk(gclk));
	jand g0721(.dina(n1035),.dinb(w_n774_0[0]),.dout(n1036),.clk(gclk));
	jand g0722(.dina(w_dff_B_Wrw5Hqd19_0),.dinb(n1034),.dout(n1037),.clk(gclk));
	jand g0723(.dina(n1037),.dinb(w_dff_B_gbMbJoQG1_1),.dout(n1038),.clk(gclk));
	jor g0724(.dina(n1038),.dinb(w_dff_B_q2ed6MJC2_1),.dout(n1039),.clk(gclk));
	jxor g0725(.dina(w_n734_0[1]),.dinb(w_n373_3[0]),.dout(n1040),.clk(gclk));
	jxor g0726(.dina(w_n729_0[2]),.dinb(w_n726_0[2]),.dout(n1041),.clk(gclk));
	jand g0727(.dina(n1041),.dinb(w_n724_0[0]),.dout(n1042),.clk(gclk));
	jand g0728(.dina(w_n1042_0[1]),.dinb(w_n749_0[0]),.dout(n1043),.clk(gclk));
	jand g0729(.dina(n1043),.dinb(w_dff_B_akVBs4rW7_1),.dout(n1044),.clk(gclk));
	jand g0730(.dina(w_dff_B_g3X5V15h0_0),.dinb(n1039),.dout(n1045),.clk(gclk));
	jor g0731(.dina(w_G2204_0[1]),.dinb(w_G1455_0[1]),.dout(n1046),.clk(gclk));
	jor g0732(.dina(n1046),.dinb(w_n367_0[0]),.dout(n1047),.clk(gclk));
	jand g0733(.dina(n1047),.dinb(w_G38_1[1]),.dout(n1048),.clk(gclk));
	jand g0734(.dina(w_n723_0[1]),.dinb(w_n720_0[1]),.dout(n1049),.clk(gclk));
	jand g0735(.dina(w_n741_1[0]),.dinb(w_n737_1[0]),.dout(n1050),.clk(gclk));
	jor g0736(.dina(w_n741_0[2]),.dinb(w_n737_0[2]),.dout(n1051),.clk(gclk));
	jand g0737(.dina(w_n747_0[1]),.dinb(w_n744_0[1]),.dout(n1052),.clk(gclk));
	jand g0738(.dina(n1052),.dinb(n1051),.dout(n1053),.clk(gclk));
	jor g0739(.dina(n1053),.dinb(w_dff_B_gMtGkkf78_1),.dout(n1054),.clk(gclk));
	jand g0740(.dina(n1054),.dinb(w_n1042_0[0]),.dout(n1055),.clk(gclk));
	jor g0741(.dina(n1055),.dinb(w_dff_B_LOovrd8T7_1),.dout(n1056),.clk(gclk));
	jor g0742(.dina(n1056),.dinb(w_dff_B_aLZtl6TB0_1),.dout(n1057),.clk(gclk));
	jor g0743(.dina(w_dff_B_4OlEFcVr6_0),.dinb(n1045),.dout(n1058),.clk(gclk));
	jor g0744(.dina(n1058),.dinb(w_dff_B_BQCItuAB9_1),.dout(n1059),.clk(gclk));
	jand g0745(.dina(w_n1059_0[2]),.dinb(w_n718_0[2]),.dout(w_dff_A_C7Y9DVay5_2),.clk(gclk));
	jnot g0746(.din(w_n644_0[0]),.dout(n1061),.clk(gclk));
	jnot g0747(.din(w_n655_0[0]),.dout(n1062),.clk(gclk));
	jnot g0748(.din(w_n656_0[0]),.dout(n1063),.clk(gclk));
	jand g0749(.dina(w_n641_0[1]),.dinb(w_G3705_1[0]),.dout(n1064),.clk(gclk));
	jor g0750(.dina(w_n641_0[0]),.dinb(w_G3705_0[2]),.dout(n1065),.clk(gclk));
	jand g0751(.dina(n1065),.dinb(w_n354_0[1]),.dout(n1066),.clk(gclk));
	jor g0752(.dina(n1066),.dinb(w_dff_B_q4V9eCAW1_1),.dout(n1067),.clk(gclk));
	jor g0753(.dina(w_n1067_0[2]),.dinb(w_dff_B_8t3jpyCn9_1),.dout(n1068),.clk(gclk));
	jand g0754(.dina(n1068),.dinb(w_dff_B_Tjb98FfF9_1),.dout(n1069),.clk(gclk));
	jand g0755(.dina(w_n1069_0[2]),.dinb(n1061),.dout(n1070),.clk(gclk));
	jnot g0756(.din(w_n1070_0[1]),.dout(n1071),.clk(gclk));
	jor g0757(.dina(w_n669_0[0]),.dinb(w_G4526_2[0]),.dout(n1072),.clk(gclk));
	jand g0758(.dina(w_dff_B_QW2NFVLj0_0),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0759(.dina(w_n1073_0[1]),.dinb(w_n654_0[1]),.dout(n1074),.clk(gclk));
	jand g0760(.dina(n1074),.dinb(w_n653_0[0]),.dout(n1075),.clk(gclk));
	jxor g0761(.dina(n1075),.dinb(w_n626_1[0]),.dout(w_dff_A_oa0XxNvS3_2),.clk(gclk));
	jxor g0762(.dina(w_n1073_0[0]),.dinb(w_n631_0[1]),.dout(w_dff_A_NyvscHrC9_2),.clk(gclk));
	jand g0763(.dina(w_n359_0[2]),.dinb(w_G4526_1[2]),.dout(n1078),.clk(gclk));
	jor g0764(.dina(w_n666_0[0]),.dinb(w_n1078_0[1]),.dout(n1079),.clk(gclk));
	jand g0765(.dina(n1079),.dinb(w_n661_0[1]),.dout(n1080),.clk(gclk));
	jxor g0766(.dina(n1080),.dinb(w_n636_0[1]),.dout(w_dff_A_lPzfP2la9_2),.clk(gclk));
	jor g0767(.dina(w_n1078_0[0]),.dinb(w_n664_0[0]),.dout(n1082),.clk(gclk));
	jxor g0768(.dina(n1082),.dinb(w_n642_0[1]),.dout(w_dff_A_JmJfu1Jx3_2),.clk(gclk));
	jxor g0769(.dina(w_n585_0[2]),.dinb(w_n582_0[0]),.dout(n1084),.clk(gclk));
	jor g0770(.dina(w_n1084_0[2]),.dinb(w_n678_0[0]),.dout(n1085),.clk(gclk));
	jnot g0771(.din(w_n646_0[0]),.dout(n1086),.clk(gclk));
	jnot g0772(.din(w_n647_0[0]),.dout(n1087),.clk(gclk));
	jnot g0773(.din(w_n654_0[0]),.dout(n1088),.clk(gclk));
	jand g0774(.dina(w_n1069_0[1]),.dinb(w_dff_B_45VyFlQB5_1),.dout(n1089),.clk(gclk));
	jor g0775(.dina(n1089),.dinb(w_n652_0[0]),.dout(n1090),.clk(gclk));
	jor g0776(.dina(w_n1090_0[1]),.dinb(w_n649_0[0]),.dout(n1091),.clk(gclk));
	jand g0777(.dina(n1091),.dinb(w_dff_B_bqNfjuoh2_1),.dout(n1092),.clk(gclk));
	jand g0778(.dina(w_n1092_0[2]),.dinb(w_n1086_0[1]),.dout(n1093),.clk(gclk));
	jnot g0779(.din(w_G4526_1[1]),.dout(n1094),.clk(gclk));
	jand g0780(.dina(w_n1092_0[1]),.dinb(w_n1094_0[2]),.dout(n1095),.clk(gclk));
	jor g0781(.dina(n1095),.dinb(n1093),.dout(n1096),.clk(gclk));
	jand g0782(.dina(w_n1096_0[1]),.dinb(w_n618_0[0]),.dout(n1097),.clk(gclk));
	jor g0783(.dina(n1097),.dinb(w_n619_0[1]),.dout(n1098),.clk(gclk));
	jor g0784(.dina(n1098),.dinb(w_n588_0[0]),.dout(n1099),.clk(gclk));
	jor g0785(.dina(w_n1099_0[1]),.dinb(w_n586_0[1]),.dout(n1100),.clk(gclk));
	jand g0786(.dina(n1100),.dinb(w_dff_B_iv2qALu13_1),.dout(w_dff_A_SGZG573Y4_2),.clk(gclk));
	jand g0787(.dina(w_n676_0[1]),.dinb(w_n605_0[1]),.dout(n1102),.clk(gclk));
	jor g0788(.dina(n1102),.dinb(w_n615_0[1]),.dout(n1103),.clk(gclk));
	jxor g0789(.dina(n1103),.dinb(w_n594_0[1]),.dout(w_dff_A_1iQksQaM0_2),.clk(gclk));
	jnot g0790(.din(w_n599_0[0]),.dout(n1105),.clk(gclk));
	jnot g0791(.din(w_n613_0[1]),.dout(n1106),.clk(gclk));
	jnot g0792(.din(w_n603_0[2]),.dout(n1107),.clk(gclk));
	jand g0793(.dina(n1107),.dinb(w_G3729_0[2]),.dout(n1108),.clk(gclk));
	jor g0794(.dina(w_n1096_0[0]),.dinb(w_n1108_0[1]),.dout(n1109),.clk(gclk));
	jand g0795(.dina(n1109),.dinb(w_n1106_0[1]),.dout(n1110),.clk(gclk));
	jxor g0796(.dina(n1110),.dinb(w_n1105_0[1]),.dout(w_dff_A_8hS9m2Y73_2),.clk(gclk));
	jxor g0797(.dina(w_n676_0[0]),.dinb(w_n604_0[0]),.dout(w_dff_A_QdpmjzBx0_2),.clk(gclk));
	jnot g0798(.din(w_n436_0[0]),.dout(n1113),.clk(gclk));
	jor g0799(.dina(w_n1113_0[1]),.dinb(w_n431_0[0]),.dout(n1114),.clk(gclk));
	jnot g0800(.din(w_n432_0[0]),.dout(n1115),.clk(gclk));
	jor g0801(.dina(w_n435_0[0]),.dinb(n1115),.dout(n1116),.clk(gclk));
	jand g0802(.dina(n1116),.dinb(n1114),.dout(n1117),.clk(gclk));
	jnot g0803(.din(w_n459_0[0]),.dout(n1118),.clk(gclk));
	jxor g0804(.dina(w_n1118_0[1]),.dinb(w_n453_0[1]),.dout(n1119),.clk(gclk));
	jxor g0805(.dina(w_dff_B_gg1Pz5RC7_0),.dinb(n1117),.dout(n1120),.clk(gclk));
	jxor g0806(.dina(w_n485_0[0]),.dinb(w_n469_0[1]),.dout(n1121),.clk(gclk));
	jor g0807(.dina(w_n440_0[0]),.dinb(w_n422_0[0]),.dout(n1122),.clk(gclk));
	jnot g0808(.din(w_n423_0[0]),.dout(n1123),.clk(gclk));
	jor g0809(.dina(w_n427_0[0]),.dinb(n1123),.dout(n1124),.clk(gclk));
	jand g0810(.dina(n1124),.dinb(n1122),.dout(n1125),.clk(gclk));
	jnot g0811(.din(G141),.dout(n1126),.clk(gclk));
	jor g0812(.dina(n1126),.dinb(w_G18_20[0]),.dout(n1127),.clk(gclk));
	jnot g0813(.din(G161),.dout(n1128),.clk(gclk));
	jor g0814(.dina(n1128),.dinb(w_n355_15[0]),.dout(n1129),.clk(gclk));
	jand g0815(.dina(n1129),.dinb(w_n1127_0[1]),.dout(n1130),.clk(gclk));
	jxor g0816(.dina(n1130),.dinb(w_n479_0[2]),.dout(n1131),.clk(gclk));
	jxor g0817(.dina(w_dff_B_jXbhs1Ts2_0),.dinb(n1125),.dout(n1132),.clk(gclk));
	jxor g0818(.dina(n1132),.dinb(w_dff_B_31ztlG9W9_1),.dout(n1133),.clk(gclk));
	jxor g0819(.dina(n1133),.dinb(w_dff_B_oSRhgFo17_1),.dout(n1134),.clk(gclk));
	jxor g0820(.dina(w_n603_0[1]),.dinb(w_n598_0[2]),.dout(n1135),.clk(gclk));
	jand g0821(.dina(G239),.dinb(w_G18_19[2]),.dout(n1136),.clk(gclk));
	jand g0822(.dina(w_dff_B_1rrGnPMp2_0),.dinb(w_n355_14[2]),.dout(n1137),.clk(gclk));
	jor g0823(.dina(w_n1137_0[1]),.dinb(w_dff_B_8KC414ka4_1),.dout(n1138),.clk(gclk));
	jxor g0824(.dina(w_dff_B_gX7dCrmQ4_0),.dinb(w_n651_0[0]),.dout(n1139),.clk(gclk));
	jxor g0825(.dina(n1139),.dinb(w_dff_B_L7MDHylB8_1),.dout(n1140),.clk(gclk));
	jand g0826(.dina(G229),.dinb(w_G18_19[1]),.dout(n1141),.clk(gclk));
	jor g0827(.dina(w_dff_B_T8lypvRC0_0),.dinb(w_n663_0[2]),.dout(n1142),.clk(gclk));
	jxor g0828(.dina(n1142),.dinb(w_n660_0[0]),.dout(n1143),.clk(gclk));
	jxor g0829(.dina(w_n635_0[1]),.dinb(w_n625_0[1]),.dout(n1144),.clk(gclk));
	jxor g0830(.dina(n1144),.dinb(n1143),.dout(n1145),.clk(gclk));
	jxor g0831(.dina(w_n593_0[1]),.dinb(w_n585_0[1]),.dout(n1146),.clk(gclk));
	jxor g0832(.dina(w_dff_B_VqDCOUdL7_0),.dinb(n1145),.dout(n1147),.clk(gclk));
	jxor g0833(.dina(n1147),.dinb(n1140),.dout(n1148),.clk(gclk));
	jor g0834(.dina(w_dff_B_DruvH7gb4_0),.dinb(n1134),.dout(n1149),.clk(gclk));
	jor g0835(.dina(w_n372_0[0]),.dinb(w_n355_14[1]),.dout(n1150),.clk(gclk));
	jxor g0836(.dina(G212),.dinb(G211),.dout(n1151),.clk(gclk));
	jxor g0837(.dina(n1151),.dinb(w_G209_0[0]),.dout(n1152),.clk(gclk));
	jor g0838(.dina(n1152),.dinb(w_n1150_0[1]),.dout(n1153),.clk(gclk));
	jnot g0839(.din(w_n386_0[0]),.dout(n1154),.clk(gclk));
	jand g0840(.dina(w_n395_0[2]),.dinb(n1154),.dout(n1155),.clk(gclk));
	jnot g0841(.din(w_n394_0[0]),.dout(n1156),.clk(gclk));
	jand g0842(.dina(n1156),.dinb(w_n387_0[1]),.dout(n1157),.clk(gclk));
	jor g0843(.dina(n1157),.dinb(n1155),.dout(n1158),.clk(gclk));
	jor g0844(.dina(w_n380_0[0]),.dinb(w_n374_0[0]),.dout(n1159),.clk(gclk));
	jnot g0845(.din(w_n375_0[0]),.dout(n1160),.clk(gclk));
	jor g0846(.dina(w_n378_0[0]),.dinb(n1160),.dout(n1161),.clk(gclk));
	jand g0847(.dina(n1161),.dinb(n1159),.dout(n1162),.clk(gclk));
	jxor g0848(.dina(n1162),.dinb(w_dff_B_ElLWtjbo3_1),.dout(n1163),.clk(gclk));
	jxor g0849(.dina(n1163),.dinb(w_dff_B_r4wVXBmI4_1),.dout(n1164),.clk(gclk));
	jxor g0850(.dina(w_n689_0[0]),.dinb(w_n504_0[2]),.dout(n1165),.clk(gclk));
	jxor g0851(.dina(w_n523_0[0]),.dinb(w_n517_0[2]),.dout(n1166),.clk(gclk));
	jxor g0852(.dina(w_dff_B_hETOkRjX2_0),.dinb(n1165),.dout(n1167),.clk(gclk));
	jxor g0853(.dina(w_n555_0[1]),.dinb(w_n539_0[1]),.dout(n1168),.clk(gclk));
	jxor g0854(.dina(w_n547_0[1]),.dinb(w_n531_0[1]),.dout(n1169),.clk(gclk));
	jxor g0855(.dina(n1169),.dinb(n1168),.dout(n1170),.clk(gclk));
	jand g0856(.dina(G227),.dinb(w_G18_19[0]),.dout(n1171),.clk(gclk));
	jand g0857(.dina(w_dff_B_CwWHlkEl2_0),.dinb(w_n355_14[0]),.dout(n1172),.clk(gclk));
	jor g0858(.dina(w_n1172_0[1]),.dinb(w_dff_B_iO12gpId8_1),.dout(n1173),.clk(gclk));
	jxor g0859(.dina(n1173),.dinb(w_n563_0[2]),.dout(n1174),.clk(gclk));
	jxor g0860(.dina(w_dff_B_qZ37TkEr6_0),.dinb(n1170),.dout(n1175),.clk(gclk));
	jxor g0861(.dina(n1175),.dinb(n1167),.dout(n1176),.clk(gclk));
	jor g0862(.dina(w_dff_B_nYIWO4Zh3_0),.dinb(n1164),.dout(n1177),.clk(gclk));
	jor g0863(.dina(w_dff_B_rfMi1FXX7_0),.dinb(n1149),.dout(G412_fa_),.clk(gclk));
	jnot g0864(.din(w_n772_0[0]),.dout(n1179),.clk(gclk));
	jxor g0865(.dina(w_n780_0[0]),.dinb(n1179),.dout(n1180),.clk(gclk));
	jnot g0866(.din(w_G2208_0[1]),.dout(n1181),.clk(gclk));
	jor g0867(.dina(n1181),.dinb(w_n355_13[2]),.dout(n1182),.clk(gclk));
	jor g0868(.dina(G82),.dinb(w_G18_18[2]),.dout(n1183),.clk(gclk));
	jand g0869(.dina(w_dff_B_motdm5k38_0),.dinb(n1182),.dout(n1184),.clk(gclk));
	jxor g0870(.dina(n1184),.dinb(w_n827_0[0]),.dout(n1185),.clk(gclk));
	jxor g0871(.dina(w_dff_B_eweljXyV3_0),.dinb(n1180),.dout(n1186),.clk(gclk));
	jxor g0872(.dina(w_n806_0[0]),.dinb(w_n800_0[1]),.dout(n1187),.clk(gclk));
	jxor g0873(.dina(w_n820_0[0]),.dinb(w_n814_0[1]),.dout(n1188),.clk(gclk));
	jxor g0874(.dina(n1188),.dinb(n1187),.dout(n1189),.clk(gclk));
	jxor g0875(.dina(w_n764_0[0]),.dinb(w_n758_0[1]),.dout(n1190),.clk(gclk));
	jxor g0876(.dina(w_dff_B_ZDQVdoiT8_0),.dinb(n1189),.dout(n1191),.clk(gclk));
	jxor g0877(.dina(n1191),.dinb(n1186),.dout(n1192),.clk(gclk));
	jxor g0878(.dina(w_n953_0[1]),.dinb(w_n947_0[0]),.dout(n1193),.clk(gclk));
	jxor g0879(.dina(w_n903_0[0]),.dinb(w_n894_0[0]),.dout(n1194),.clk(gclk));
	jxor g0880(.dina(n1194),.dinb(n1193),.dout(n1195),.clk(gclk));
	jnot g0881(.din(w_G3698_0[1]),.dout(n1196),.clk(gclk));
	jor g0882(.dina(n1196),.dinb(w_n355_13[1]),.dout(n1197),.clk(gclk));
	jor g0883(.dina(G69),.dinb(w_G18_18[1]),.dout(n1198),.clk(gclk));
	jand g0884(.dina(w_dff_B_jCyB9P0P2_0),.dinb(n1197),.dout(n1199),.clk(gclk));
	jxor g0885(.dina(n1199),.dinb(w_n888_0[0]),.dout(n1200),.clk(gclk));
	jor g0886(.dina(w_n662_0[0]),.dinb(w_n355_13[0]),.dout(n1201),.clk(gclk));
	jand g0887(.dina(n1201),.dinb(w_n905_0[0]),.dout(n1202),.clk(gclk));
	jxor g0888(.dina(n1202),.dinb(w_n919_0[0]),.dout(n1203),.clk(gclk));
	jxor g0889(.dina(n1203),.dinb(n1200),.dout(n1204),.clk(gclk));
	jnot g0890(.din(w_n930_0[0]),.dout(n1205),.clk(gclk));
	jxor g0891(.dina(w_n938_0[0]),.dinb(n1205),.dout(n1206),.clk(gclk));
	jxor g0892(.dina(n1206),.dinb(n1204),.dout(n1207),.clk(gclk));
	jxor g0893(.dina(n1207),.dinb(w_dff_B_LWRHO66N8_1),.dout(n1208),.clk(gclk));
	jor g0894(.dina(n1208),.dinb(n1192),.dout(n1209),.clk(gclk));
	jxor g0895(.dina(w_n854_0[0]),.dinb(w_n848_0[1]),.dout(n1210),.clk(gclk));
	jxor g0896(.dina(w_n870_0[0]),.dinb(w_n862_0[0]),.dout(n1211),.clk(gclk));
	jxor g0897(.dina(n1211),.dinb(n1210),.dout(n1212),.clk(gclk));
	jxor g0898(.dina(w_n983_0[0]),.dinb(w_n977_0[1]),.dout(n1213),.clk(gclk));
	jand g0899(.dina(w_G4393_0[1]),.dinb(w_G18_18[0]),.dout(n1214),.clk(gclk));
	jnot g0900(.din(G58),.dout(n1215),.clk(gclk));
	jand g0901(.dina(n1215),.dinb(w_n355_12[2]),.dout(n1216),.clk(gclk));
	jor g0902(.dina(n1216),.dinb(w_dff_B_VAnidCBK9_1),.dout(n1217),.clk(gclk));
	jxor g0903(.dina(n1217),.dinb(w_n970_0[0]),.dout(n1218),.clk(gclk));
	jxor g0904(.dina(w_n999_0[0]),.dinb(w_n991_0[0]),.dout(n1219),.clk(gclk));
	jxor g0905(.dina(n1219),.dinb(n1218),.dout(n1220),.clk(gclk));
	jxor g0906(.dina(n1220),.dinb(w_dff_B_mmKU2qf88_1),.dout(n1221),.clk(gclk));
	jxor g0907(.dina(n1221),.dinb(w_dff_B_UT7DX8AU3_1),.dout(n1222),.clk(gclk));
	jxor g0908(.dina(w_n366_0[0]),.dinb(w_G1492_1[0]),.dout(n1223),.clk(gclk));
	jor g0909(.dina(n1223),.dinb(w_n355_12[1]),.dout(n1224),.clk(gclk));
	jnot g0910(.din(w_G1455_0[0]),.dout(n1225),.clk(gclk));
	jxor g0911(.dina(w_G2204_0[0]),.dinb(n1225),.dout(n1226),.clk(gclk));
	jor g0912(.dina(n1226),.dinb(w_G18_17[2]),.dout(n1227),.clk(gclk));
	jand g0913(.dina(n1227),.dinb(n1224),.dout(n1228),.clk(gclk));
	jxor g0914(.dina(w_n729_0[1]),.dinb(w_n723_0[0]),.dout(n1229),.clk(gclk));
	jxor g0915(.dina(w_n747_0[0]),.dinb(w_n741_0[1]),.dout(n1230),.clk(gclk));
	jxor g0916(.dina(n1230),.dinb(n1229),.dout(n1231),.clk(gclk));
	jnot g0917(.din(w_G1459_0[1]),.dout(n1232),.clk(gclk));
	jor g0918(.dina(n1232),.dinb(w_n355_12[0]),.dout(n1233),.clk(gclk));
	jor g0919(.dina(G114),.dinb(w_G18_17[1]),.dout(n1234),.clk(gclk));
	jand g0920(.dina(w_dff_B_FIx2mURg1_0),.dinb(n1233),.dout(n1235),.clk(gclk));
	jxor g0921(.dina(n1235),.dinb(w_n734_0[0]),.dout(n1236),.clk(gclk));
	jxor g0922(.dina(w_dff_B_VaOgOo7R7_0),.dinb(n1231),.dout(n1237),.clk(gclk));
	jxor g0923(.dina(n1237),.dinb(w_dff_B_Y00uvtA76_1),.dout(n1238),.clk(gclk));
	jor g0924(.dina(n1238),.dinb(n1222),.dout(n1239),.clk(gclk));
	jor g0925(.dina(n1239),.dinb(n1209),.dout(G414_fa_),.clk(gclk));
	jnot g0926(.din(w_n935_0[0]),.dout(n1241),.clk(gclk));
	jxor g0927(.dina(n1241),.dinb(w_n926_0[0]),.dout(n1242),.clk(gclk));
	jxor g0928(.dina(w_n950_0[1]),.dinb(w_n944_0[0]),.dout(n1243),.clk(gclk));
	jxor g0929(.dina(w_dff_B_5YrEWmCa8_0),.dinb(n1242),.dout(n1244),.clk(gclk));
	jand g0930(.dina(G208),.dinb(w_G18_17[0]),.dout(n1245),.clk(gclk));
	jor g0931(.dina(w_dff_B_Jrk5eOK59_0),.dinb(w_n1137_0[0]),.dout(n1246),.clk(gclk));
	jand g0932(.dina(G198),.dinb(w_G18_16[2]),.dout(n1247),.clk(gclk));
	jor g0933(.dina(w_dff_B_9bgLBXQJ9_0),.dinb(w_n663_0[1]),.dout(n1248),.clk(gclk));
	jxor g0934(.dina(n1248),.dinb(n1246),.dout(n1249),.clk(gclk));
	jxor g0935(.dina(w_n916_0[0]),.dinb(w_n885_0[0]),.dout(n1250),.clk(gclk));
	jxor g0936(.dina(n1250),.dinb(n1249),.dout(n1251),.clk(gclk));
	jxor g0937(.dina(w_n900_0[0]),.dinb(w_n891_0[0]),.dout(n1252),.clk(gclk));
	jxor g0938(.dina(w_dff_B_g6xz6nVJ6_0),.dinb(n1251),.dout(n1253),.clk(gclk));
	jxor g0939(.dina(n1253),.dinb(n1244),.dout(n1254),.clk(gclk));
	jxor g0940(.dina(w_n866_0[0]),.dinb(w_n858_0[0]),.dout(n1255),.clk(gclk));
	jxor g0941(.dina(w_n995_0[0]),.dinb(w_n987_0[0]),.dout(n1256),.clk(gclk));
	jxor g0942(.dina(n1256),.dinb(n1255),.dout(n1257),.clk(gclk));
	jxor g0943(.dina(w_n980_0[0]),.dinb(w_n973_0[1]),.dout(n1258),.clk(gclk));
	jand g0944(.dina(G197),.dinb(w_G18_16[1]),.dout(n1259),.clk(gclk));
	jor g0945(.dina(w_dff_B_lnZwKp530_0),.dinb(w_n1172_0[0]),.dout(n1260),.clk(gclk));
	jxor g0946(.dina(n1260),.dinb(w_n966_0[0]),.dout(n1261),.clk(gclk));
	jxor g0947(.dina(n1261),.dinb(n1258),.dout(n1262),.clk(gclk));
	jnot g0948(.din(w_n851_0[0]),.dout(n1263),.clk(gclk));
	jxor g0949(.dina(n1263),.dinb(w_n845_0[1]),.dout(n1264),.clk(gclk));
	jxor g0950(.dina(n1264),.dinb(n1262),.dout(n1265),.clk(gclk));
	jxor g0951(.dina(n1265),.dinb(w_dff_B_9v9MOOrH2_1),.dout(n1266),.clk(gclk));
	jor g0952(.dina(n1266),.dinb(n1254),.dout(n1267),.clk(gclk));
	jxor g0953(.dina(G165),.dinb(G164),.dout(n1268),.clk(gclk));
	jxor g0954(.dina(n1268),.dinb(w_dff_B_4OUwLuKY1_1),.dout(n1269),.clk(gclk));
	jor g0955(.dina(n1269),.dinb(w_n1150_0[0]),.dout(n1270),.clk(gclk));
	jnot g0956(.din(w_n736_0[0]),.dout(n1271),.clk(gclk));
	jand g0957(.dina(w_n744_0[0]),.dinb(n1271),.dout(n1272),.clk(gclk));
	jnot g0958(.din(w_n743_0[0]),.dout(n1273),.clk(gclk));
	jand g0959(.dina(n1273),.dinb(w_n737_0[1]),.dout(n1274),.clk(gclk));
	jor g0960(.dina(n1274),.dinb(n1272),.dout(n1275),.clk(gclk));
	jnot g0961(.din(w_n726_0[1]),.dout(n1276),.clk(gclk));
	jor g0962(.dina(n1276),.dinb(w_n719_0[0]),.dout(n1277),.clk(gclk));
	jnot g0963(.din(w_n720_0[0]),.dout(n1278),.clk(gclk));
	jor g0964(.dina(w_n725_0[0]),.dinb(n1278),.dout(n1279),.clk(gclk));
	jand g0965(.dina(n1279),.dinb(n1277),.dout(n1280),.clk(gclk));
	jxor g0966(.dina(n1280),.dinb(w_dff_B_9B07w0IG3_1),.dout(n1281),.clk(gclk));
	jxor g0967(.dina(n1281),.dinb(w_dff_B_yr36TW4i6_1),.dout(n1282),.clk(gclk));
	jor g0968(.dina(n1282),.dinb(n1267),.dout(n1283),.clk(gclk));
	jnot g0969(.din(G181),.dout(n1284),.clk(gclk));
	jor g0970(.dina(n1284),.dinb(w_n355_11[2]),.dout(n1285),.clk(gclk));
	jand g0971(.dina(n1285),.dinb(w_n1127_0[0]),.dout(n1286),.clk(gclk));
	jxor g0972(.dina(n1286),.dinb(w_n824_0[0]),.dout(n1287),.clk(gclk));
	jxor g0973(.dina(w_n803_0[0]),.dinb(w_n796_0[1]),.dout(n1288),.clk(gclk));
	jxor g0974(.dina(n1288),.dinb(n1287),.dout(n1289),.clk(gclk));
	jnot g0975(.din(w_n767_0[0]),.dout(n1290),.clk(gclk));
	jand g0976(.dina(w_n776_0[0]),.dinb(n1290),.dout(n1291),.clk(gclk));
	jnot g0977(.din(w_n775_0[0]),.dout(n1292),.clk(gclk));
	jand g0978(.dina(n1292),.dinb(w_n768_0[0]),.dout(n1293),.clk(gclk));
	jor g0979(.dina(n1293),.dinb(n1291),.dout(n1294),.clk(gclk));
	jnot g0980(.din(w_n754_0[0]),.dout(n1295),.clk(gclk));
	jand g0981(.dina(w_n761_0[0]),.dinb(n1295),.dout(n1296),.clk(gclk));
	jnot g0982(.din(w_n760_0[0]),.dout(n1297),.clk(gclk));
	jand g0983(.dina(n1297),.dinb(w_n755_0[1]),.dout(n1298),.clk(gclk));
	jor g0984(.dina(n1298),.dinb(n1296),.dout(n1299),.clk(gclk));
	jxor g0985(.dina(n1299),.dinb(n1294),.dout(n1300),.clk(gclk));
	jxor g0986(.dina(w_n817_0[0]),.dinb(w_n810_0[1]),.dout(n1301),.clk(gclk));
	jxor g0987(.dina(w_dff_B_78xqVym44_0),.dinb(n1300),.dout(n1302),.clk(gclk));
	jxor g0988(.dina(n1302),.dinb(w_dff_B_pwJz712V9_1),.dout(n1303),.clk(gclk));
	jor g0989(.dina(w_dff_B_dxTagTcf8_0),.dinb(n1283),.dout(G416_fa_),.clk(gclk));
	jnot g0990(.din(w_n480_1[0]),.dout(n1305),.clk(gclk));
	jnot g0991(.din(w_n505_0[0]),.dout(n1306),.clk(gclk));
	jnot g0992(.din(w_n513_1[0]),.dout(n1307),.clk(gclk));
	jnot g0993(.din(w_n524_1[0]),.dout(n1308),.clk(gclk));
	jnot g0994(.din(w_n572_1[0]),.dout(n1309),.clk(gclk));
	jnot g0995(.din(w_n581_0[1]),.dout(n1310),.clk(gclk));
	jnot g0996(.din(w_n586_0[0]),.dout(n1311),.clk(gclk));
	jand g0997(.dina(w_n1099_0[0]),.dinb(w_dff_B_R7AEYJd50_1),.dout(n1312),.clk(gclk));
	jor g0998(.dina(w_n1312_1[1]),.dinb(w_n1310_0[1]),.dout(n1313),.clk(gclk));
	jand g0999(.dina(n1313),.dinb(w_n1309_0[1]),.dout(n1314),.clk(gclk));
	jor g1000(.dina(n1314),.dinb(w_n526_0[1]),.dout(n1315),.clk(gclk));
	jor g1001(.dina(n1315),.dinb(w_n1308_0[1]),.dout(n1316),.clk(gclk));
	jor g1002(.dina(w_n1316_0[1]),.dinb(w_n518_1[0]),.dout(n1317),.clk(gclk));
	jor g1003(.dina(w_n1317_0[1]),.dinb(w_n1307_0[1]),.dout(n1318),.clk(gclk));
	jand g1004(.dina(w_n696_0[0]),.dinb(n1318),.dout(n1319),.clk(gclk));
	jor g1005(.dina(n1319),.dinb(w_n507_0[0]),.dout(n1320),.clk(gclk));
	jand g1006(.dina(n1320),.dinb(w_dff_B_ikio3lpP7_1),.dout(n1321),.clk(gclk));
	jxor g1007(.dina(w_n1321_1[1]),.dinb(w_dff_B_ypHWpTQ32_1),.dout(w_dff_A_xfiKRwPP3_2),.clk(gclk));
	jnot g1008(.din(w_n414_1[0]),.dout(n1323),.clk(gclk));
	jnot g1009(.din(w_n424_0[0]),.dout(n1324),.clk(gclk));
	jnot g1010(.din(w_n425_1[0]),.dout(n1325),.clk(gclk));
	jnot g1011(.din(w_n450_0[1]),.dout(n1326),.clk(gclk));
	jnot g1012(.din(w_n449_0[2]),.dout(n1327),.clk(gclk));
	jnot g1013(.din(w_n499_0[0]),.dout(n1328),.clk(gclk));
	jnot g1014(.din(w_n500_0[0]),.dout(n1329),.clk(gclk));
	jnot g1015(.din(w_n462_0[0]),.dout(n1330),.clk(gclk));
	jand g1016(.dina(w_n1321_1[0]),.dinb(w_dff_B_luDCltd93_1),.dout(n1331),.clk(gclk));
	jand g1017(.dina(n1331),.dinb(w_dff_B_rHabs0Ds3_1),.dout(n1332),.clk(gclk));
	jor g1018(.dina(n1332),.dinb(w_dff_B_NAgtVxZD0_1),.dout(n1333),.clk(gclk));
	jand g1019(.dina(w_n1333_0[1]),.dinb(w_dff_B_nd1RsLIr9_1),.dout(n1334),.clk(gclk));
	jor g1020(.dina(n1334),.dinb(w_dff_B_rnCe3Ork8_1),.dout(n1335),.clk(gclk));
	jor g1021(.dina(n1335),.dinb(w_dff_B_vp9A2Y2X7_1),.dout(n1336),.clk(gclk));
	jand g1022(.dina(n1336),.dinb(w_dff_B_zmbOQOvP3_1),.dout(n1337),.clk(gclk));
	jxor g1023(.dina(w_n1337_1[1]),.dinb(w_n1323_0[1]),.dout(w_dff_A_zrcXL1rl7_2),.clk(gclk));
	jand g1024(.dina(w_n1118_0[0]),.dinb(w_G2230_0[1]),.dout(n1339),.clk(gclk));
	jnot g1025(.din(n1339),.dout(n1340),.clk(gclk));
	jand g1026(.dina(w_n1321_0[2]),.dinb(w_n495_1[0]),.dout(n1341),.clk(gclk));
	jnot g1027(.din(n1341),.dout(n1342),.clk(gclk));
	jand g1028(.dina(n1342),.dinb(w_n497_1[0]),.dout(n1343),.clk(gclk));
	jand g1029(.dina(w_n1343_0[1]),.dinb(w_n1340_0[2]),.dout(n1344),.clk(gclk));
	jor g1030(.dina(w_n1344_0[1]),.dinb(w_n460_1[1]),.dout(n1345),.clk(gclk));
	jxor g1031(.dina(n1345),.dinb(w_n463_1[0]),.dout(w_dff_A_gwDlvvGS8_2),.clk(gclk));
	jor g1032(.dina(w_n1343_0[0]),.dinb(w_n464_0[1]),.dout(n1347),.clk(gclk));
	jnot g1033(.din(w_n1344_0[0]),.dout(n1348),.clk(gclk));
	jor g1034(.dina(n1348),.dinb(w_n460_1[0]),.dout(n1349),.clk(gclk));
	jand g1035(.dina(n1349),.dinb(w_dff_B_y6tAviAl7_1),.dout(w_dff_A_HM3MKpQL8_2),.clk(gclk));
	jnot g1036(.din(w_n489_0[1]),.dout(n1351),.clk(gclk));
	jor g1037(.dina(n1351),.dinb(w_n491_1[0]),.dout(n1352),.clk(gclk));
	jand g1038(.dina(w_n700_1[0]),.dinb(w_n481_0[0]),.dout(n1353),.clk(gclk));
	jor g1039(.dina(n1353),.dinb(w_dff_B_Yyae2c6K8_1),.dout(n1354),.clk(gclk));
	jxor g1040(.dina(n1354),.dinb(w_n470_0[1]),.dout(w_dff_A_90iJhh3S3_2),.clk(gclk));
	jand g1041(.dina(w_n700_0[2]),.dinb(w_n480_0[2]),.dout(n1356),.clk(gclk));
	jor g1042(.dina(n1356),.dinb(w_n487_0[1]),.dout(n1357),.clk(gclk));
	jxor g1043(.dina(n1357),.dinb(w_n475_0[1]),.dout(w_dff_A_3fDqDu737_2),.clk(gclk));
	jor g1044(.dina(w_n418_0[0]),.dinb(w_n411_1[0]),.dout(n1359),.clk(gclk));
	jor g1045(.dina(w_n707_1[1]),.dinb(w_n411_0[2]),.dout(n1360),.clk(gclk));
	jand g1046(.dina(n1360),.dinb(w_n1359_0[1]),.dout(n1361),.clk(gclk));
	jxor g1047(.dina(n1361),.dinb(w_n377_1[0]),.dout(w_dff_A_F5JBNVEW3_2),.clk(gclk));
	jand g1048(.dina(w_n415_0[0]),.dinb(w_n388_1[0]),.dout(n1363),.clk(gclk));
	jor g1049(.dina(w_dff_B_6Xm9GNkp1_0),.dinb(w_n409_1[0]),.dout(n1364),.clk(gclk));
	jor g1050(.dina(w_n707_1[0]),.dinb(w_n409_0[2]),.dout(n1365),.clk(gclk));
	jand g1051(.dina(n1365),.dinb(w_n1364_0[1]),.dout(n1366),.clk(gclk));
	jxor g1052(.dina(n1366),.dinb(w_n416_0[1]),.dout(w_dff_A_4qm3SZjK2_2),.clk(gclk));
	jnot g1053(.din(w_n388_0[2]),.dout(n1368),.clk(gclk));
	jnot g1054(.din(w_n396_1[0]),.dout(n1369),.clk(gclk));
	jnot g1055(.din(w_n392_0[1]),.dout(n1370),.clk(gclk));
	jor g1056(.dina(w_n1337_1[0]),.dinb(w_n1323_0[0]),.dout(n1371),.clk(gclk));
	jand g1057(.dina(n1371),.dinb(w_n1370_0[1]),.dout(n1372),.clk(gclk));
	jor g1058(.dina(w_n1372_0[1]),.dinb(w_n1369_0[1]),.dout(n1373),.clk(gclk));
	jand g1059(.dina(n1373),.dinb(w_n405_0[1]),.dout(n1374),.clk(gclk));
	jxor g1060(.dina(n1374),.dinb(w_dff_B_Vk81izGt4_1),.dout(G333),.clk(gclk));
	jxor g1061(.dina(w_n1372_0[0]),.dinb(w_n1369_0[0]),.dout(w_dff_A_LuZMZecF1_2),.clk(gclk));
	jor g1062(.dina(w_G416_0),.dinb(w_G414_0),.dout(n1377),.clk(gclk));
	jor g1063(.dina(w_G408_0),.dinb(w_G404_0),.dout(n1378),.clk(gclk));
	jor g1064(.dina(w_G410_0),.dinb(w_G406_0),.dout(n1379),.clk(gclk));
	jor g1065(.dina(w_dff_B_hU40mBNJ5_0),.dinb(w_G412_0),.dout(n1380),.clk(gclk));
	jor g1066(.dina(n1380),.dinb(w_dff_B_D3ju29x52_1),.dout(n1381),.clk(gclk));
	jor g1067(.dina(n1381),.dinb(w_dff_B_oJ3uk5Yu9_1),.dout(w_dff_A_DpK9MJgg0_2),.clk(gclk));
	jxor g1068(.dina(w_n705_0[0]),.dinb(w_n425_0[2]),.dout(w_dff_A_66Kxv2s37_2),.clk(gclk));
	jand g1069(.dina(w_n703_1[1]),.dinb(w_n438_0[0]),.dout(n1384),.clk(gclk));
	jor g1070(.dina(n1384),.dinb(w_n447_0[1]),.dout(n1385),.clk(gclk));
	jxor g1071(.dina(n1385),.dinb(w_n429_0[1]),.dout(w_dff_A_Zf5g3S756_2),.clk(gclk));
	jand g1072(.dina(w_n1113_0[0]),.dinb(w_G2239_0[2]),.dout(n1387),.clk(gclk));
	jnot g1073(.din(w_n1387_0[1]),.dout(n1388),.clk(gclk));
	jor g1074(.dina(w_n703_1[0]),.dinb(w_n445_0[1]),.dout(n1389),.clk(gclk));
	jand g1075(.dina(n1389),.dinb(w_n1388_0[1]),.dout(n1390),.clk(gclk));
	jxor g1076(.dina(n1390),.dinb(w_n433_1[0]),.dout(w_dff_A_5ZJ7pWXu5_2),.clk(gclk));
	jxor g1077(.dina(w_n703_0[2]),.dinb(w_n437_0[1]),.dout(w_dff_A_xlZ8L1W07_2),.clk(gclk));
	jxor g1078(.dina(w_n680_2[1]),.dinb(w_n575_1[0]),.dout(w_dff_A_NpO6pto17_2),.clk(gclk));
	jor g1079(.dina(w_n712_0[1]),.dinb(w_G38_1[0]),.dout(n1394),.clk(gclk));
	jor g1080(.dina(w_n713_0[0]),.dinb(w_n709_1[0]),.dout(n1395),.clk(gclk));
	jand g1081(.dina(n1395),.dinb(w_dff_B_5a4TbPj14_1),.dout(n1396),.clk(gclk));
	jxor g1082(.dina(w_n1396_0[1]),.dinb(w_n370_0[1]),.dout(G422),.clk(gclk));
	jxor g1083(.dina(w_n709_0[2]),.dinb(w_n363_0[1]),.dout(w_dff_A_5xWKymr18_2),.clk(gclk));
	jand g1084(.dina(w_n680_2[0]),.dinb(w_n580_0[1]),.dout(n1399),.clk(gclk));
	jor g1085(.dina(n1399),.dinb(w_n570_1[1]),.dout(n1400),.clk(gclk));
	jxor g1086(.dina(n1400),.dinb(w_n573_1[0]),.dout(w_dff_A_gjRLzgIm3_2),.clk(gclk));
	jnot g1087(.din(w_n577_0[0]),.dout(n1402),.clk(gclk));
	jnot g1088(.din(w_n548_0[0]),.dout(n1403),.clk(gclk));
	jnot g1089(.din(w_n566_0[1]),.dout(n1404),.clk(gclk));
	jnot g1090(.din(w_n576_0[1]),.dout(n1405),.clk(gclk));
	jand g1091(.dina(w_dff_B_CnVb1Lwf1_0),.dinb(n1404),.dout(n1406),.clk(gclk));
	jor g1092(.dina(n1406),.dinb(w_n550_0[0]),.dout(n1407),.clk(gclk));
	jand g1093(.dina(n1407),.dinb(w_dff_B_rqgIY5ES8_1),.dout(n1408),.clk(gclk));
	jnot g1094(.din(w_n568_0[1]),.dout(n1409),.clk(gclk));
	jand g1095(.dina(w_n1312_1[0]),.dinb(w_dff_B_LQia12gc9_1),.dout(n1410),.clk(gclk));
	jor g1096(.dina(n1410),.dinb(w_n1408_0[1]),.dout(n1411),.clk(gclk));
	jxor g1097(.dina(n1411),.dinb(w_n1402_0[1]),.dout(w_dff_A_A4XOy4fh6_2),.clk(gclk));
	jand g1098(.dina(w_n680_1[2]),.dinb(w_n576_0[0]),.dout(n1413),.clk(gclk));
	jor g1099(.dina(n1413),.dinb(w_n566_0[0]),.dout(n1414),.clk(gclk));
	jxor g1100(.dina(n1414),.dinb(w_n578_0[1]),.dout(w_dff_A_aqO8jZ6A6_2),.clk(gclk));
	jand g1101(.dina(w_n680_1[1]),.dinb(w_n575_0[2]),.dout(n1416),.clk(gclk));
	jor g1102(.dina(n1416),.dinb(w_n564_0[1]),.dout(n1417),.clk(gclk));
	jxor g1103(.dina(n1417),.dinb(w_n574_0[1]),.dout(w_dff_A_7pKYbPVy4_2),.clk(gclk));
	jxor g1104(.dina(w_n504_0[1]),.dinb(w_n501_0[0]),.dout(n1419),.clk(gclk));
	jxor g1105(.dina(w_n1419_0[1]),.dinb(w_n698_0[0]),.dout(w_dff_A_QExPo0Wj9_2),.clk(gclk));
	jand g1106(.dina(w_n694_0[0]),.dinb(w_n1317_0[0]),.dout(n1421),.clk(gclk));
	jxor g1107(.dina(n1421),.dinb(w_n1307_0[0]),.dout(w_dff_A_RRVhlcbP2_2),.clk(gclk));
	jxor g1108(.dina(w_n524_0[2]),.dinb(w_n518_0[2]),.dout(n1423),.clk(gclk));
	jor g1109(.dina(w_dff_B_9Ijh9dG00_0),.dinb(w_n683_0[0]),.dout(n1424),.clk(gclk));
	jand g1110(.dina(n1424),.dinb(w_n1316_0[0]),.dout(w_dff_A_lnookEJx5_2),.clk(gclk));
	jxor g1111(.dina(w_n517_0[1]),.dinb(w_n514_0[0]),.dout(n1426),.clk(gclk));
	jxor g1112(.dina(w_n1426_0[1]),.dinb(w_n682_0[0]),.dout(w_dff_A_fSEwKRmD3_2),.clk(gclk));
	jxor g1113(.dina(w_n429_0[0]),.dinb(w_n425_0[1]),.dout(n1431),.clk(gclk));
	jor g1114(.dina(w_n1388_0[0]),.dinb(w_n444_0[1]),.dout(n1432),.clk(gclk));
	jnot g1115(.din(w_n447_0[0]),.dout(n1433),.clk(gclk));
	jor g1116(.dina(w_n1433_0[1]),.dinb(w_n1387_0[0]),.dout(n1434),.clk(gclk));
	jand g1117(.dina(n1434),.dinb(w_dff_B_Jyi5VW8h0_1),.dout(n1435),.clk(gclk));
	jxor g1118(.dina(n1435),.dinb(w_n1431_0[1]),.dout(n1436),.clk(gclk));
	jxor g1119(.dina(w_n449_0[1]),.dinb(w_n433_0[2]),.dout(n1437),.clk(gclk));
	jxor g1120(.dina(w_dff_B_bZewYbaQ4_0),.dinb(n1436),.dout(n1438),.clk(gclk));
	jand g1121(.dina(w_dff_B_kGTsVbyO2_0),.dinb(w_n1333_0[0]),.dout(n1439),.clk(gclk));
	jxor g1122(.dina(w_n445_0[0]),.dinb(w_n433_0[1]),.dout(n1440),.clk(gclk));
	jnot g1123(.din(w_n1440_0[1]),.dout(n1441),.clk(gclk));
	jand g1124(.dina(w_dff_B_pUYv3kJb8_0),.dinb(w_n1433_0[0]),.dout(n1442),.clk(gclk));
	jor g1125(.dina(w_n437_0[0]),.dinb(w_n444_0[0]),.dout(n1443),.clk(gclk));
	jand g1126(.dina(n1443),.dinb(w_n1440_0[0]),.dout(n1444),.clk(gclk));
	jor g1127(.dina(w_dff_B_V51AO53A2_0),.dinb(n1442),.dout(n1445),.clk(gclk));
	jxor g1128(.dina(w_n1431_0[0]),.dinb(w_n450_0[0]),.dout(n1446),.clk(gclk));
	jxor g1129(.dina(n1446),.dinb(w_dff_B_4HAgZNzg2_1),.dout(n1447),.clk(gclk));
	jand g1130(.dina(w_dff_B_NGsbwMpe2_0),.dinb(w_n703_0[1]),.dout(n1448),.clk(gclk));
	jor g1131(.dina(n1448),.dinb(n1439),.dout(n1449),.clk(gclk));
	jand g1132(.dina(w_n497_0[2]),.dinb(w_n1340_0[1]),.dout(n1450),.clk(gclk));
	jor g1133(.dina(n1450),.dinb(w_n460_0[2]),.dout(n1451),.clk(gclk));
	jxor g1134(.dina(w_n480_0[1]),.dinb(w_n475_0[0]),.dout(n1452),.clk(gclk));
	jand g1135(.dina(w_n1452_0[2]),.dinb(w_n495_0[2]),.dout(n1453),.clk(gclk));
	jnot g1136(.din(w_n1452_0[1]),.dout(n1454),.clk(gclk));
	jand g1137(.dina(w_dff_B_lc2rTYBf5_0),.dinb(w_n497_0[1]),.dout(n1455),.clk(gclk));
	jor g1138(.dina(n1455),.dinb(w_dff_B_8MmWqEbC1_1),.dout(n1456),.clk(gclk));
	jnot g1139(.din(w_n479_0[1]),.dout(n1457),.clk(gclk));
	jand g1140(.dina(n1457),.dinb(w_G2211_0[1]),.dout(n1458),.clk(gclk));
	jnot g1141(.din(w_n1458_0[1]),.dout(n1459),.clk(gclk));
	jor g1142(.dina(n1459),.dinb(w_n491_0[2]),.dout(n1460),.clk(gclk));
	jor g1143(.dina(w_n1458_0[0]),.dinb(w_n486_0[0]),.dout(n1461),.clk(gclk));
	jand g1144(.dina(w_dff_B_KYND4Y7A2_0),.dinb(n1460),.dout(n1462),.clk(gclk));
	jxor g1145(.dina(n1462),.dinb(w_n463_0[2]),.dout(n1463),.clk(gclk));
	jxor g1146(.dina(w_dff_B_b9b3rXR82_0),.dinb(n1456),.dout(n1464),.clk(gclk));
	jxor g1147(.dina(n1464),.dinb(w_dff_B_PL1JEJ9U9_1),.dout(n1465),.clk(gclk));
	jand g1148(.dina(w_dff_B_INOpmN2v9_0),.dinb(w_n700_0[1]),.dout(n1466),.clk(gclk));
	jand g1149(.dina(w_n496_0[0]),.dinb(w_n1340_0[0]),.dout(n1467),.clk(gclk));
	jor g1150(.dina(n1467),.dinb(w_n460_0[1]),.dout(n1468),.clk(gclk));
	jor g1151(.dina(w_n487_0[0]),.dinb(w_n491_0[1]),.dout(n1469),.clk(gclk));
	jand g1152(.dina(w_dff_B_mxWw4cXU4_0),.dinb(w_n489_0[0]),.dout(n1470),.clk(gclk));
	jxor g1153(.dina(n1470),.dinb(w_n463_0[1]),.dout(n1471),.clk(gclk));
	jxor g1154(.dina(n1471),.dinb(w_n495_0[1]),.dout(n1472),.clk(gclk));
	jxor g1155(.dina(n1472),.dinb(w_n1452_0[0]),.dout(n1473),.clk(gclk));
	jxor g1156(.dina(w_dff_B_hephm8TV5_0),.dinb(n1468),.dout(n1474),.clk(gclk));
	jand g1157(.dina(w_dff_B_GfyjoT731_0),.dinb(w_n1321_0[1]),.dout(n1475),.clk(gclk));
	jor g1158(.dina(n1475),.dinb(n1466),.dout(n1476),.clk(gclk));
	jxor g1159(.dina(w_n470_0[0]),.dinb(w_n464_0[0]),.dout(n1477),.clk(gclk));
	jxor g1160(.dina(w_dff_B_AXN5zYGA4_0),.dinb(n1476),.dout(n1478),.clk(gclk));
	jxor g1161(.dina(w_dff_B_12HAZl668_0),.dinb(n1449),.dout(w_dff_A_kjGGFBjr5_2),.clk(gclk));
	jxor g1162(.dina(w_n416_0[0]),.dinb(w_n388_0[1]),.dout(n1480),.clk(gclk));
	jxor g1163(.dina(w_n411_0[1]),.dinb(w_n377_0[2]),.dout(n1481),.clk(gclk));
	jand g1164(.dina(w_n407_0[0]),.dinb(w_n1370_0[0]),.dout(n1482),.clk(gclk));
	jand g1165(.dina(w_n409_0[1]),.dinb(w_n392_0[0]),.dout(n1483),.clk(gclk));
	jor g1166(.dina(n1483),.dinb(w_dff_B_0FngQeLD3_1),.dout(n1484),.clk(gclk));
	jnot g1167(.din(w_n397_0[0]),.dout(n1485),.clk(gclk));
	jand g1168(.dina(n1485),.dinb(w_n405_0[0]),.dout(n1486),.clk(gclk));
	jxor g1169(.dina(w_n414_0[2]),.dinb(w_n396_0[2]),.dout(n1487),.clk(gclk));
	jxor g1170(.dina(w_dff_B_nODN7bvz1_0),.dinb(w_n1486_0[1]),.dout(n1488),.clk(gclk));
	jxor g1171(.dina(w_dff_B_4T9BR8210_0),.dinb(n1484),.dout(n1489),.clk(gclk));
	jxor g1172(.dina(n1489),.dinb(n1481),.dout(n1490),.clk(gclk));
	jor g1173(.dina(w_dff_B_QktJqICt2_0),.dinb(w_n707_0[2]),.dout(n1491),.clk(gclk));
	jor g1174(.dina(w_n391_0[0]),.dinb(w_n389_0[1]),.dout(n1492),.clk(gclk));
	jor g1175(.dina(w_n395_0[1]),.dinb(w_n393_0[1]),.dout(n1493),.clk(gclk));
	jand g1176(.dina(n1493),.dinb(w_n1492_0[1]),.dout(n1494),.clk(gclk));
	jnot g1177(.din(w_n1492_0[0]),.dout(n1495),.clk(gclk));
	jand g1178(.dina(w_n1486_0[0]),.dinb(w_dff_B_zpFoqYh97_1),.dout(n1496),.clk(gclk));
	jor g1179(.dina(n1496),.dinb(w_dff_B_SFXMS2uJ4_1),.dout(n1497),.clk(gclk));
	jxor g1180(.dina(w_n396_0[1]),.dinb(w_n377_0[1]),.dout(n1498),.clk(gclk));
	jxor g1181(.dina(w_dff_B_7TJ07BqD6_0),.dinb(w_n1364_0[0]),.dout(n1499),.clk(gclk));
	jxor g1182(.dina(n1499),.dinb(w_dff_B_Wz9LiyGS3_1),.dout(n1500),.clk(gclk));
	jxor g1183(.dina(n1500),.dinb(w_n414_0[1]),.dout(n1501),.clk(gclk));
	jxor g1184(.dina(n1501),.dinb(w_n1359_0[0]),.dout(n1502),.clk(gclk));
	jor g1185(.dina(w_dff_B_AHUCtzZZ4_0),.dinb(w_n1337_0[2]),.dout(n1503),.clk(gclk));
	jand g1186(.dina(n1503),.dinb(n1491),.dout(n1504),.clk(gclk));
	jxor g1187(.dina(n1504),.dinb(w_dff_B_QwCIe8H74_1),.dout(n1505),.clk(gclk));
	jand g1188(.dina(w_n362_0[0]),.dinb(w_G38_0[2]),.dout(n1506),.clk(gclk));
	jnot g1189(.din(w_n364_0[1]),.dout(n1507),.clk(gclk));
	jor g1190(.dina(n1507),.dinb(w_n1506_0[1]),.dout(n1508),.clk(gclk));
	jnot g1191(.din(w_n1506_0[0]),.dout(n1509),.clk(gclk));
	jor g1192(.dina(n1509),.dinb(w_G1496_0[2]),.dout(n1510),.clk(gclk));
	jand g1193(.dina(n1510),.dinb(w_dff_B_GB5UhtBF0_1),.dout(n1511),.clk(gclk));
	jand g1194(.dina(w_n1511_0[1]),.dinb(w_n413_0[2]),.dout(n1512),.clk(gclk));
	jnot g1195(.din(w_n413_0[1]),.dout(n1513),.clk(gclk));
	jand g1196(.dina(w_n712_0[0]),.dinb(w_n361_0[0]),.dout(n1514),.clk(gclk));
	jor g1197(.dina(w_n364_0[0]),.dinb(n1514),.dout(n1515),.clk(gclk));
	jor g1198(.dina(w_n369_0[0]),.dinb(w_G1492_0[2]),.dout(n1516),.clk(gclk));
	jand g1199(.dina(n1516),.dinb(n1515),.dout(n1517),.clk(gclk));
	jand g1200(.dina(w_dff_B_myCTkUXi8_0),.dinb(n1513),.dout(n1518),.clk(gclk));
	jor g1201(.dina(w_n1518_0[1]),.dinb(w_dff_B_iVnIzRsb0_1),.dout(n1519),.clk(gclk));
	jor g1202(.dina(w_dff_B_Nrh579qe2_0),.dinb(w_n707_0[1]),.dout(n1520),.clk(gclk));
	jnot g1203(.din(w_n419_0[0]),.dout(n1521),.clk(gclk));
	jand g1204(.dina(w_n1518_0[0]),.dinb(w_dff_B_28qkGFQB2_1),.dout(n1522),.clk(gclk));
	jand g1205(.dina(w_n1511_0[0]),.dinb(w_n420_0[0]),.dout(n1523),.clk(gclk));
	jor g1206(.dina(w_dff_B_JwRnG0pd9_0),.dinb(n1522),.dout(n1524),.clk(gclk));
	jor g1207(.dina(w_dff_B_JykNhceB1_0),.dinb(w_n1337_0[1]),.dout(n1525),.clk(gclk));
	jand g1208(.dina(n1525),.dinb(n1520),.dout(n1526),.clk(gclk));
	jxor g1209(.dina(w_dff_B_7Lz0IC683_0),.dinb(n1505),.dout(w_dff_A_3AVLPWfs6_2),.clk(gclk));
	jor g1210(.dina(w_n693_0[0]),.dinb(w_n687_0[0]),.dout(n1528),.clk(gclk));
	jand g1211(.dina(w_dff_B_X5UPQFDB0_0),.dinb(w_n695_0[0]),.dout(n1529),.clk(gclk));
	jor g1212(.dina(w_n1529_0[1]),.dinb(w_n513_0[2]),.dout(n1530),.clk(gclk));
	jxor g1213(.dina(w_n1419_0[0]),.dinb(w_n1308_0[0]),.dout(n1531),.clk(gclk));
	jxor g1214(.dina(w_n1531_0[1]),.dinb(w_n526_0[0]),.dout(n1532),.clk(gclk));
	jxor g1215(.dina(w_dff_B_qoeLEU5k2_0),.dinb(n1530),.dout(n1533),.clk(gclk));
	jand g1216(.dina(w_dff_B_mrMzToCv7_0),.dinb(w_n1309_0[0]),.dout(n1534),.clk(gclk));
	jand g1217(.dina(w_n1534_0[1]),.dinb(w_n1310_0[0]),.dout(n1535),.clk(gclk));
	jand g1218(.dina(w_n1426_0[0]),.dinb(w_n524_0[1]),.dout(n1536),.clk(gclk));
	jnot g1219(.din(w_n1536_0[1]),.dout(n1537),.clk(gclk));
	jor g1220(.dina(n1537),.dinb(w_n690_0[0]),.dout(n1538),.clk(gclk));
	jor g1221(.dina(w_n1536_0[0]),.dinb(w_n1529_0[0]),.dout(n1539),.clk(gclk));
	jand g1222(.dina(n1539),.dinb(w_dff_B_EU2ykJhL3_1),.dout(n1540),.clk(gclk));
	jxor g1223(.dina(w_n518_0[1]),.dinb(w_n513_0[1]),.dout(n1541),.clk(gclk));
	jxor g1224(.dina(w_dff_B_FkQP94Gv6_0),.dinb(w_n1531_0[0]),.dout(n1542),.clk(gclk));
	jxor g1225(.dina(w_dff_B_4xMheUue8_0),.dinb(n1540),.dout(n1543),.clk(gclk));
	jor g1226(.dina(w_n581_0[0]),.dinb(w_n572_0[2]),.dout(n1544),.clk(gclk));
	jand g1227(.dina(n1544),.dinb(w_n1543_0[1]),.dout(n1545),.clk(gclk));
	jor g1228(.dina(w_dff_B_eZ81QOBf4_0),.dinb(n1535),.dout(n1546),.clk(gclk));
	jand g1229(.dina(n1546),.dinb(w_n680_1[0]),.dout(n1547),.clk(gclk));
	jand g1230(.dina(w_n1543_0[0]),.dinb(w_n572_0[1]),.dout(n1548),.clk(gclk));
	jor g1231(.dina(w_dff_B_JC4Q6jwA2_0),.dinb(w_n1534_0[0]),.dout(n1549),.clk(gclk));
	jand g1232(.dina(w_dff_B_1eGYARXL9_0),.dinb(w_n1312_0[2]),.dout(n1550),.clk(gclk));
	jor g1233(.dina(n1550),.dinb(n1547),.dout(n1551),.clk(gclk));
	jxor g1234(.dina(w_n578_0[0]),.dinb(w_n1402_0[0]),.dout(n1552),.clk(gclk));
	jnot g1235(.din(w_n563_0[1]),.dout(n1553),.clk(gclk));
	jand g1236(.dina(n1553),.dinb(w_G4394_0[2]),.dout(n1554),.clk(gclk));
	jnot g1237(.din(w_n1554_0[1]),.dout(n1555),.clk(gclk));
	jand g1238(.dina(n1555),.dinb(w_n558_0[0]),.dout(n1556),.clk(gclk));
	jand g1239(.dina(w_n1554_0[0]),.dinb(w_n556_0[1]),.dout(n1557),.clk(gclk));
	jor g1240(.dina(w_dff_B_FFuF2WM68_0),.dinb(n1556),.dout(n1558),.clk(gclk));
	jxor g1241(.dina(n1558),.dinb(w_n573_0[2]),.dout(n1559),.clk(gclk));
	jxor g1242(.dina(w_dff_B_I4GYQyWz0_0),.dinb(w_n1408_0[0]),.dout(n1560),.clk(gclk));
	jnot g1243(.din(w_n570_1[0]),.dout(n1561),.clk(gclk));
	jxor g1244(.dina(w_n575_0[1]),.dinb(w_n574_0[0]),.dout(n1562),.clk(gclk));
	jnot g1245(.din(w_n1562_0[2]),.dout(n1563),.clk(gclk));
	jor g1246(.dina(w_dff_B_zwd4YUXK8_0),.dinb(n1561),.dout(n1564),.clk(gclk));
	jor g1247(.dina(w_n1562_0[1]),.dinb(w_n570_0[2]),.dout(n1565),.clk(gclk));
	jor g1248(.dina(n1565),.dinb(w_n580_0[0]),.dout(n1566),.clk(gclk));
	jand g1249(.dina(n1566),.dinb(n1564),.dout(n1567),.clk(gclk));
	jxor g1250(.dina(n1567),.dinb(w_dff_B_USdYKckw6_1),.dout(n1568),.clk(gclk));
	jor g1251(.dina(w_dff_B_qgka1V8r4_0),.dinb(w_n1312_0[1]),.dout(n1569),.clk(gclk));
	jxor g1252(.dina(w_n1562_0[0]),.dinb(w_n570_0[1]),.dout(n1570),.clk(gclk));
	jnot g1253(.din(w_n565_0[0]),.dout(n1571),.clk(gclk));
	jor g1254(.dina(w_n564_0[0]),.dinb(w_n556_0[0]),.dout(n1572),.clk(gclk));
	jand g1255(.dina(w_dff_B_23s7cY9T8_0),.dinb(n1571),.dout(n1573),.clk(gclk));
	jxor g1256(.dina(n1573),.dinb(w_n573_0[1]),.dout(n1574),.clk(gclk));
	jxor g1257(.dina(n1574),.dinb(w_n568_0[0]),.dout(n1575),.clk(gclk));
	jxor g1258(.dina(w_dff_B_iiTVZbst1_0),.dinb(n1570),.dout(n1576),.clk(gclk));
	jor g1259(.dina(w_dff_B_zXwjkqDF0_0),.dinb(w_n680_0[2]),.dout(n1577),.clk(gclk));
	jand g1260(.dina(n1577),.dinb(n1569),.dout(n1578),.clk(gclk));
	jxor g1261(.dina(n1578),.dinb(w_dff_B_c6sAlVSH7_1),.dout(n1579),.clk(gclk));
	jxor g1262(.dina(n1579),.dinb(w_dff_B_03bsOFBl3_1),.dout(w_dff_A_oM4MwWtI5_2),.clk(gclk));
	jxor g1263(.dina(w_n1084_0[1]),.dinb(w_n1108_0[0]),.dout(n1581),.clk(gclk));
	jxor g1264(.dina(n1581),.dinb(w_n1105_0[0]),.dout(n1582),.clk(gclk));
	jand g1265(.dina(w_n616_0[0]),.dinb(w_n609_0[0]),.dout(n1583),.clk(gclk));
	jand g1266(.dina(w_n615_0[0]),.dinb(w_n610_0[0]),.dout(n1584),.clk(gclk));
	jor g1267(.dina(w_dff_B_JV2A6PtL3_0),.dinb(n1583),.dout(n1585),.clk(gclk));
	jxor g1268(.dina(n1585),.dinb(w_dff_B_mGxIXwGq5_1),.dout(n1586),.clk(gclk));
	jand g1269(.dina(w_dff_B_ivaSIiH18_0),.dinb(w_n1092_0[0]),.dout(n1587),.clk(gclk));
	jand g1270(.dina(w_n1587_0[1]),.dinb(w_n1086_0[0]),.dout(n1588),.clk(gclk));
	jnot g1271(.din(w_n598_0[1]),.dout(n1589),.clk(gclk));
	jand g1272(.dina(n1589),.dinb(w_G3737_0[1]),.dout(n1590),.clk(gclk));
	jand g1273(.dina(w_n1106_0[0]),.dinb(n1590),.dout(n1591),.clk(gclk));
	jand g1274(.dina(w_n613_0[0]),.dinb(w_n612_0[0]),.dout(n1592),.clk(gclk));
	jor g1275(.dina(w_dff_B_0XqqsElB1_0),.dinb(n1591),.dout(n1593),.clk(gclk));
	jor g1276(.dina(n1593),.dinb(w_n605_0[0]),.dout(n1594),.clk(gclk));
	jxor g1277(.dina(w_n1084_0[0]),.dinb(w_n594_0[0]),.dout(n1595),.clk(gclk));
	jxor g1278(.dina(w_dff_B_ZmV7R1xK6_0),.dinb(n1594),.dout(n1596),.clk(gclk));
	jxor g1279(.dina(w_dff_B_3XopZPmy5_0),.dinb(w_n619_0[0]),.dout(n1597),.clk(gclk));
	jand g1280(.dina(w_n1597_0[1]),.dinb(w_n674_0[0]),.dout(n1598),.clk(gclk));
	jor g1281(.dina(n1598),.dinb(w_n1094_0[1]),.dout(n1599),.clk(gclk));
	jor g1282(.dina(n1599),.dinb(w_dff_B_YtMXNCep7_1),.dout(n1600),.clk(gclk));
	jand g1283(.dina(w_n1597_0[0]),.dinb(w_n673_0[0]),.dout(n1601),.clk(gclk));
	jor g1284(.dina(n1601),.dinb(w_n1587_0[0]),.dout(n1602),.clk(gclk));
	jor g1285(.dina(n1602),.dinb(w_G4526_1[0]),.dout(n1603),.clk(gclk));
	jand g1286(.dina(w_dff_B_NWmQF8Ab9_0),.dinb(n1600),.dout(n1604),.clk(gclk));
	jxor g1287(.dina(w_n642_0[0]),.dinb(w_n359_0[1]),.dout(n1605),.clk(gclk));
	jxor g1288(.dina(w_n1605_0[1]),.dinb(w_n1067_0[1]),.dout(n1606),.clk(gclk));
	jxor g1289(.dina(w_dff_B_5Ifwxcif7_0),.dinb(w_n1069_0[0]),.dout(n1607),.clk(gclk));
	jnot g1290(.din(w_n1607_0[1]),.dout(n1608),.clk(gclk));
	jxor g1291(.dina(w_n626_0[2]),.dinb(w_n354_0[0]),.dout(n1609),.clk(gclk));
	jxor g1292(.dina(w_dff_B_fEle8DqW2_0),.dinb(w_n671_0[0]),.dout(n1610),.clk(gclk));
	jor g1293(.dina(w_n1610_0[1]),.dinb(w_dff_B_pGs50NTd7_1),.dout(n1611),.clk(gclk));
	jnot g1294(.din(w_n1610_0[0]),.dout(n1612),.clk(gclk));
	jor g1295(.dina(n1612),.dinb(w_n1607_0[0]),.dout(n1613),.clk(gclk));
	jand g1296(.dina(n1613),.dinb(w_n1094_0[0]),.dout(n1614),.clk(gclk));
	jand g1297(.dina(n1614),.dinb(w_dff_B_9hQjcZU16_1),.dout(n1615),.clk(gclk));
	jand g1298(.dina(w_n1067_0[0]),.dinb(w_n357_0[0]),.dout(n1616),.clk(gclk));
	jand g1299(.dina(w_n661_0[0]),.dinb(w_n358_0[0]),.dout(n1617),.clk(gclk));
	jor g1300(.dina(w_dff_B_r2mzG9rG0_0),.dinb(n1616),.dout(n1618),.clk(gclk));
	jxor g1301(.dina(n1618),.dinb(w_n626_0[1]),.dout(n1619),.clk(gclk));
	jxor g1302(.dina(n1619),.dinb(w_n1070_0[0]),.dout(n1620),.clk(gclk));
	jnot g1303(.din(w_n1620_0[1]),.dout(n1621),.clk(gclk));
	jnot g1304(.din(w_n645_0[0]),.dout(n1622),.clk(gclk));
	jand g1305(.dina(w_n1090_0[0]),.dinb(w_dff_B_qI4S16l17_1),.dout(n1623),.clk(gclk));
	jxor g1306(.dina(n1623),.dinb(w_n1605_0[0]),.dout(n1624),.clk(gclk));
	jnot g1307(.din(w_n1624_0[1]),.dout(n1625),.clk(gclk));
	jor g1308(.dina(n1625),.dinb(w_dff_B_NIqczoov3_1),.dout(n1626),.clk(gclk));
	jor g1309(.dina(w_n1624_0[0]),.dinb(w_n1620_0[0]),.dout(n1627),.clk(gclk));
	jand g1310(.dina(n1627),.dinb(w_G4526_0[2]),.dout(n1628),.clk(gclk));
	jand g1311(.dina(n1628),.dinb(n1626),.dout(n1629),.clk(gclk));
	jor g1312(.dina(n1629),.dinb(n1615),.dout(n1630),.clk(gclk));
	jxor g1313(.dina(w_n636_0[0]),.dinb(w_n631_0[0]),.dout(n1631),.clk(gclk));
	jxor g1314(.dina(w_dff_B_dE3sVdpW8_0),.dinb(n1630),.dout(n1632),.clk(gclk));
	jxor g1315(.dina(n1632),.dinb(n1604),.dout(w_dff_A_SZHKifOh5_2),.clk(gclk));
	jdff g1316(.din(w_G1_1[1]),.dout(w_dff_A_StDwqhMe5_1),.clk(gclk));
	jdff g1317(.din(w_G1_1[0]),.dout(w_dff_A_lnaQpt5X0_1),.clk(gclk));
	jdff g1318(.din(w_G1459_0[0]),.dout(w_dff_A_nByzfYml7_1),.clk(gclk));
	jdff g1319(.din(w_G1469_0[0]),.dout(w_dff_A_X1gH7vPc7_1),.clk(gclk));
	jdff g1320(.din(w_G1480_0[0]),.dout(w_dff_A_uLsdXGj77_1),.clk(gclk));
	jdff g1321(.din(w_G1486_0[0]),.dout(w_dff_A_2l1hqVy46_1),.clk(gclk));
	jdff g1322(.din(w_G1492_0[1]),.dout(w_dff_A_HiWLfWKP7_1),.clk(gclk));
	jdff g1323(.din(w_G1496_0[1]),.dout(w_dff_A_kvGxlUzO4_1),.clk(gclk));
	jdff g1324(.din(w_G2208_0[0]),.dout(w_dff_A_fKxVyEvG8_1),.clk(gclk));
	jdff g1325(.din(w_G2218_0[0]),.dout(w_dff_A_AcwEvtBl8_1),.clk(gclk));
	jdff g1326(.din(w_G2224_0[1]),.dout(w_dff_A_z4lHrBEn5_1),.clk(gclk));
	jdff g1327(.din(w_G2230_0[0]),.dout(w_dff_A_36IIFIIA7_1),.clk(gclk));
	jdff g1328(.din(w_G2236_0[0]),.dout(w_dff_A_DXzas7OV3_1),.clk(gclk));
	jdff g1329(.din(w_G2239_0[1]),.dout(w_dff_A_8wLrcBEf7_1),.clk(gclk));
	jdff g1330(.din(w_G2247_0[0]),.dout(w_dff_A_0XQfGMjy7_1),.clk(gclk));
	jdff g1331(.din(w_G2253_0[0]),.dout(w_dff_A_azIhLlon4_1),.clk(gclk));
	jdff g1332(.din(w_G2256_0[0]),.dout(w_dff_A_OfRm1bFs5_1),.clk(gclk));
	jdff g1333(.din(w_G3698_0[0]),.dout(w_dff_A_4CAs5RJf1_1),.clk(gclk));
	jdff g1334(.din(w_G3701_0[1]),.dout(w_dff_A_C0h2PJSo2_1),.clk(gclk));
	jdff g1335(.din(w_G3705_0[1]),.dout(w_dff_A_pxhHMs847_1),.clk(gclk));
	jdff g1336(.din(w_G3711_0[0]),.dout(w_dff_A_PaiAskYr6_1),.clk(gclk));
	jdff g1337(.din(w_G3717_0[0]),.dout(w_dff_A_Nu4uyITW4_1),.clk(gclk));
	jdff g1338(.din(w_G3723_0[0]),.dout(w_dff_A_Ol3YBVCw1_1),.clk(gclk));
	jdff g1339(.din(w_G3729_0[1]),.dout(w_dff_A_vskJrkeb7_1),.clk(gclk));
	jdff g1340(.din(w_G3737_0[0]),.dout(w_dff_A_RaK8syet9_1),.clk(gclk));
	jdff g1341(.din(w_G3743_0[0]),.dout(w_dff_A_rcmF46MD0_1),.clk(gclk));
	jdff g1342(.din(w_G3749_0[0]),.dout(w_dff_A_dxxPtiY89_1),.clk(gclk));
	jdff g1343(.din(w_G4393_0[0]),.dout(w_dff_A_k9lEreo95_1),.clk(gclk));
	jdff g1344(.din(w_G4400_0[1]),.dout(w_dff_A_OvoAegEm6_1),.clk(gclk));
	jdff g1345(.din(w_G4405_0[1]),.dout(w_dff_A_tWFx69fK7_1),.clk(gclk));
	jdff g1346(.din(w_G4410_0[0]),.dout(w_dff_A_WpSOD8rp3_1),.clk(gclk));
	jdff g1347(.din(w_G4415_0[1]),.dout(w_dff_A_0Bt12MFX2_1),.clk(gclk));
	jdff g1348(.din(w_G4420_0[1]),.dout(w_dff_A_Btoykzj63_1),.clk(gclk));
	jdff g1349(.din(w_G4427_0[0]),.dout(w_dff_A_Mp0c0e9T0_1),.clk(gclk));
	jdff g1350(.din(w_G4432_0[0]),.dout(w_dff_A_ReeCzHam0_1),.clk(gclk));
	jdff g1351(.din(w_G4437_0[0]),.dout(w_dff_A_wNDkqV9X6_1),.clk(gclk));
	jdff g1352(.din(w_G1462_0[0]),.dout(w_dff_A_3rxkWg5S9_1),.clk(gclk));
	jdff g1353(.din(w_G2211_0[0]),.dout(w_dff_A_VGhsnYzH9_1),.clk(gclk));
	jdff g1354(.din(w_G4394_0[1]),.dout(w_dff_A_JFXSKKkp5_1),.clk(gclk));
	jdff g1355(.din(w_G1_0[2]),.dout(w_dff_A_qBosUjhi3_1),.clk(gclk));
	jdff g1356(.din(w_G106_0[1]),.dout(w_dff_A_7CPkUKba1_1),.clk(gclk));
	jnot g1357(.din(w_G15_0[1]),.dout(w_dff_A_2CM4RefF3_1),.clk(gclk));
	jor g1358(.dina(w_n345_0[0]),.dinb(w_G5_0[1]),.dout(w_dff_A_ZwTqURVo7_2),.clk(gclk));
	jnot g1359(.din(w_G15_0[0]),.dout(w_dff_A_0w6Csyvn8_1),.clk(gclk));
	jor g1360(.dina(w_n349_0[0]),.dinb(w_n347_0[0]),.dout(w_dff_A_UKxWtnJd8_2),.clk(gclk));
	jdff g1361(.din(w_G1_0[1]),.dout(w_dff_A_M0HT7wKV8_1),.clk(gclk));
	jand g1362(.dina(w_n1059_0[1]),.dinb(w_n718_0[1]),.dout(w_dff_A_6veNz4KY3_2),.clk(gclk));
	jor g1363(.dina(w_n715_1[0]),.dinb(w_n711_1[0]),.dout(G270),.clk(gclk));
	jand g1364(.dina(w_n1059_0[0]),.dinb(w_n718_0[0]),.dout(w_dff_A_ILSvZBEJ4_2),.clk(gclk));
	jor g1365(.dina(w_n715_0[2]),.dinb(w_n711_0[2]),.dout(G276),.clk(gclk));
	jor g1366(.dina(w_n715_0[1]),.dinb(w_n711_0[1]),.dout(G273),.clk(gclk));
	jxor g1367(.dina(w_n1396_0[0]),.dinb(w_n370_0[0]),.dout(G469),.clk(gclk));
	jxor g1368(.dina(w_n709_0[1]),.dinb(w_n363_0[0]),.dout(w_dff_A_TNQyhMuw3_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G5_0(.douta(w_G5_0[0]),.doutb(w_dff_A_7au7tv7s7_1),.doutc(w_dff_A_QQzWuTYo3_2),.din(G5));
	jspl jspl_w_G5_1(.douta(w_dff_A_n9g5SFgC7_0),.doutb(w_G5_1[1]),.din(w_G5_0[0]));
	jspl3 jspl3_w_G15_0(.douta(w_G15_0[0]),.doutb(w_G15_0[1]),.doutc(w_G15_0[2]),.din(G15));
	jspl3 jspl3_w_G18_0(.douta(w_G18_0[0]),.doutb(w_G18_0[1]),.doutc(w_G18_0[2]),.din(G18));
	jspl3 jspl3_w_G18_1(.douta(w_G18_1[0]),.doutb(w_G18_1[1]),.doutc(w_G18_1[2]),.din(w_G18_0[0]));
	jspl3 jspl3_w_G18_2(.douta(w_G18_2[0]),.doutb(w_G18_2[1]),.doutc(w_G18_2[2]),.din(w_G18_0[1]));
	jspl3 jspl3_w_G18_3(.douta(w_G18_3[0]),.doutb(w_G18_3[1]),.doutc(w_G18_3[2]),.din(w_G18_0[2]));
	jspl3 jspl3_w_G18_4(.douta(w_G18_4[0]),.doutb(w_G18_4[1]),.doutc(w_G18_4[2]),.din(w_G18_1[0]));
	jspl3 jspl3_w_G18_5(.douta(w_G18_5[0]),.doutb(w_G18_5[1]),.doutc(w_G18_5[2]),.din(w_G18_1[1]));
	jspl3 jspl3_w_G18_6(.douta(w_G18_6[0]),.doutb(w_G18_6[1]),.doutc(w_G18_6[2]),.din(w_G18_1[2]));
	jspl3 jspl3_w_G18_7(.douta(w_G18_7[0]),.doutb(w_G18_7[1]),.doutc(w_G18_7[2]),.din(w_G18_2[0]));
	jspl3 jspl3_w_G18_8(.douta(w_G18_8[0]),.doutb(w_G18_8[1]),.doutc(w_G18_8[2]),.din(w_G18_2[1]));
	jspl3 jspl3_w_G18_9(.douta(w_G18_9[0]),.doutb(w_G18_9[1]),.doutc(w_G18_9[2]),.din(w_G18_2[2]));
	jspl3 jspl3_w_G18_10(.douta(w_G18_10[0]),.doutb(w_G18_10[1]),.doutc(w_G18_10[2]),.din(w_G18_3[0]));
	jspl3 jspl3_w_G18_11(.douta(w_G18_11[0]),.doutb(w_G18_11[1]),.doutc(w_G18_11[2]),.din(w_G18_3[1]));
	jspl3 jspl3_w_G18_12(.douta(w_G18_12[0]),.doutb(w_G18_12[1]),.doutc(w_G18_12[2]),.din(w_G18_3[2]));
	jspl3 jspl3_w_G18_13(.douta(w_G18_13[0]),.doutb(w_G18_13[1]),.doutc(w_G18_13[2]),.din(w_G18_4[0]));
	jspl3 jspl3_w_G18_14(.douta(w_G18_14[0]),.doutb(w_G18_14[1]),.doutc(w_G18_14[2]),.din(w_G18_4[1]));
	jspl3 jspl3_w_G18_15(.douta(w_G18_15[0]),.doutb(w_G18_15[1]),.doutc(w_G18_15[2]),.din(w_G18_4[2]));
	jspl3 jspl3_w_G18_16(.douta(w_G18_16[0]),.doutb(w_G18_16[1]),.doutc(w_G18_16[2]),.din(w_G18_5[0]));
	jspl3 jspl3_w_G18_17(.douta(w_G18_17[0]),.doutb(w_G18_17[1]),.doutc(w_dff_A_1ikDeAhx6_2),.din(w_G18_5[1]));
	jspl3 jspl3_w_G18_18(.douta(w_G18_18[0]),.doutb(w_G18_18[1]),.doutc(w_G18_18[2]),.din(w_G18_5[2]));
	jspl3 jspl3_w_G18_19(.douta(w_G18_19[0]),.doutb(w_G18_19[1]),.doutc(w_G18_19[2]),.din(w_G18_6[0]));
	jspl3 jspl3_w_G18_20(.douta(w_dff_A_HQPL7rNf1_0),.doutb(w_G18_20[1]),.doutc(w_G18_20[2]),.din(w_G18_6[1]));
	jspl3 jspl3_w_G18_21(.douta(w_G18_21[0]),.doutb(w_G18_21[1]),.doutc(w_G18_21[2]),.din(w_G18_6[2]));
	jspl3 jspl3_w_G18_22(.douta(w_G18_22[0]),.doutb(w_G18_22[1]),.doutc(w_G18_22[2]),.din(w_G18_7[0]));
	jspl3 jspl3_w_G18_23(.douta(w_G18_23[0]),.doutb(w_G18_23[1]),.doutc(w_G18_23[2]),.din(w_G18_7[1]));
	jspl3 jspl3_w_G18_24(.douta(w_G18_24[0]),.doutb(w_G18_24[1]),.doutc(w_G18_24[2]),.din(w_G18_7[2]));
	jspl3 jspl3_w_G18_25(.douta(w_G18_25[0]),.doutb(w_G18_25[1]),.doutc(w_G18_25[2]),.din(w_G18_8[0]));
	jspl3 jspl3_w_G18_26(.douta(w_G18_26[0]),.doutb(w_G18_26[1]),.doutc(w_G18_26[2]),.din(w_G18_8[1]));
	jspl3 jspl3_w_G18_27(.douta(w_G18_27[0]),.doutb(w_G18_27[1]),.doutc(w_G18_27[2]),.din(w_G18_8[2]));
	jspl3 jspl3_w_G18_28(.douta(w_G18_28[0]),.doutb(w_G18_28[1]),.doutc(w_G18_28[2]),.din(w_G18_9[0]));
	jspl3 jspl3_w_G18_29(.douta(w_G18_29[0]),.doutb(w_G18_29[1]),.doutc(w_G18_29[2]),.din(w_G18_9[1]));
	jspl3 jspl3_w_G18_30(.douta(w_G18_30[0]),.doutb(w_G18_30[1]),.doutc(w_G18_30[2]),.din(w_G18_9[2]));
	jspl3 jspl3_w_G18_31(.douta(w_G18_31[0]),.doutb(w_G18_31[1]),.doutc(w_G18_31[2]),.din(w_G18_10[0]));
	jspl3 jspl3_w_G18_32(.douta(w_G18_32[0]),.doutb(w_G18_32[1]),.doutc(w_G18_32[2]),.din(w_G18_10[1]));
	jspl3 jspl3_w_G18_33(.douta(w_G18_33[0]),.doutb(w_G18_33[1]),.doutc(w_G18_33[2]),.din(w_G18_10[2]));
	jspl3 jspl3_w_G18_34(.douta(w_G18_34[0]),.doutb(w_G18_34[1]),.doutc(w_G18_34[2]),.din(w_G18_11[0]));
	jspl3 jspl3_w_G18_35(.douta(w_G18_35[0]),.doutb(w_G18_35[1]),.doutc(w_G18_35[2]),.din(w_G18_11[1]));
	jspl3 jspl3_w_G18_36(.douta(w_G18_36[0]),.doutb(w_G18_36[1]),.doutc(w_G18_36[2]),.din(w_G18_11[2]));
	jspl3 jspl3_w_G18_37(.douta(w_G18_37[0]),.doutb(w_G18_37[1]),.doutc(w_G18_37[2]),.din(w_G18_12[0]));
	jspl3 jspl3_w_G18_38(.douta(w_G18_38[0]),.doutb(w_G18_38[1]),.doutc(w_G18_38[2]),.din(w_G18_12[1]));
	jspl3 jspl3_w_G18_39(.douta(w_G18_39[0]),.doutb(w_G18_39[1]),.doutc(w_G18_39[2]),.din(w_G18_12[2]));
	jspl3 jspl3_w_G18_40(.douta(w_G18_40[0]),.doutb(w_G18_40[1]),.doutc(w_G18_40[2]),.din(w_G18_13[0]));
	jspl3 jspl3_w_G18_41(.douta(w_G18_41[0]),.doutb(w_G18_41[1]),.doutc(w_G18_41[2]),.din(w_G18_13[1]));
	jspl3 jspl3_w_G18_42(.douta(w_G18_42[0]),.doutb(w_dff_A_h8yjWpDz5_1),.doutc(w_G18_42[2]),.din(w_G18_13[2]));
	jspl3 jspl3_w_G18_43(.douta(w_G18_43[0]),.doutb(w_G18_43[1]),.doutc(w_G18_43[2]),.din(w_G18_14[0]));
	jspl3 jspl3_w_G18_44(.douta(w_G18_44[0]),.doutb(w_G18_44[1]),.doutc(w_G18_44[2]),.din(w_G18_14[1]));
	jspl3 jspl3_w_G18_45(.douta(w_G18_45[0]),.doutb(w_G18_45[1]),.doutc(w_G18_45[2]),.din(w_G18_14[2]));
	jspl3 jspl3_w_G18_46(.douta(w_G18_46[0]),.doutb(w_G18_46[1]),.doutc(w_G18_46[2]),.din(w_G18_15[0]));
	jspl3 jspl3_w_G18_47(.douta(w_G18_47[0]),.doutb(w_G18_47[1]),.doutc(w_G18_47[2]),.din(w_G18_15[1]));
	jspl3 jspl3_w_G18_48(.douta(w_G18_48[0]),.doutb(w_G18_48[1]),.doutc(w_G18_48[2]),.din(w_G18_15[2]));
	jspl3 jspl3_w_G18_49(.douta(w_G18_49[0]),.doutb(w_G18_49[1]),.doutc(w_dff_A_sd1wNqVa8_2),.din(w_G18_16[0]));
	jspl jspl_w_G29_0(.douta(w_dff_A_tj16hwk92_0),.doutb(w_G29_0[1]),.din(G29));
	jspl3 jspl3_w_G38_0(.douta(w_dff_A_FQOPaHzv0_0),.doutb(w_G38_0[1]),.doutc(w_dff_A_sWXvFQX26_2),.din(G38));
	jspl3 jspl3_w_G38_1(.douta(w_dff_A_wVLQgSOY1_0),.doutb(w_dff_A_ihZcVA6G5_1),.doutc(w_G38_1[2]),.din(w_G38_0[0]));
	jspl3 jspl3_w_G38_2(.douta(w_dff_A_0RqgLhFE7_0),.doutb(w_dff_A_AV8fO8in9_1),.doutc(w_G38_2[2]),.din(w_G38_0[1]));
	jspl jspl_w_G41_0(.douta(w_dff_A_ox4zSsWX7_0),.doutb(w_G41_0[1]),.din(G41));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(G70));
	jspl jspl_w_G89_0(.douta(w_dff_A_ZZDYvtpd2_0),.doutb(w_G89_0[1]),.din(G89));
	jspl3 jspl3_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.doutc(w_G106_0[2]),.din(G106));
	jspl jspl_w_G106_1(.douta(w_dff_A_Ooh0LBXd5_0),.doutb(w_G106_1[1]),.din(w_G106_0[0]));
	jspl jspl_w_G209_0(.douta(w_G209_0[0]),.doutb(w_G209_0[1]),.din(w_dff_B_SYp4AUKk5_2));
	jspl jspl_w_G238_0(.douta(w_G238_0[0]),.doutb(w_G238_0[1]),.din(G238));
	jspl3 jspl3_w_G1455_0(.douta(w_G1455_0[0]),.doutb(w_G1455_0[1]),.doutc(w_G1455_0[2]),.din(G1455));
	jspl jspl_w_G1459_0(.douta(w_G1459_0[0]),.doutb(w_G1459_0[1]),.din(G1459));
	jspl jspl_w_G1462_0(.douta(w_G1462_0[0]),.doutb(w_G1462_0[1]),.din(G1462));
	jspl jspl_w_G1469_0(.douta(w_G1469_0[0]),.doutb(w_G1469_0[1]),.din(G1469));
	jspl3 jspl3_w_G1480_0(.douta(w_G1480_0[0]),.doutb(w_G1480_0[1]),.doutc(w_dff_A_lACnqkSy8_2),.din(G1480));
	jspl jspl_w_G1486_0(.douta(w_G1486_0[0]),.doutb(w_G1486_0[1]),.din(G1486));
	jspl3 jspl3_w_G1492_0(.douta(w_G1492_0[0]),.doutb(w_G1492_0[1]),.doutc(w_dff_A_0Ti9dv7b3_2),.din(G1492));
	jspl jspl_w_G1492_1(.douta(w_dff_A_jj8FWGRv1_0),.doutb(w_G1492_1[1]),.din(w_G1492_0[0]));
	jspl3 jspl3_w_G1496_0(.douta(w_G1496_0[0]),.doutb(w_G1496_0[1]),.doutc(w_dff_A_om8WZW3x7_2),.din(G1496));
	jspl jspl_w_G1496_1(.douta(w_G1496_1[0]),.doutb(w_G1496_1[1]),.din(w_G1496_0[0]));
	jspl3 jspl3_w_G2204_0(.douta(w_dff_A_Cid0r0AO1_0),.doutb(w_G2204_0[1]),.doutc(w_G2204_0[2]),.din(G2204));
	jspl jspl_w_G2208_0(.douta(w_G2208_0[0]),.doutb(w_G2208_0[1]),.din(G2208));
	jspl3 jspl3_w_G2211_0(.douta(w_G2211_0[0]),.doutb(w_dff_A_SR3YcPDr8_1),.doutc(w_G2211_0[2]),.din(G2211));
	jspl3 jspl3_w_G2218_0(.douta(w_G2218_0[0]),.doutb(w_dff_A_MCNX1YCM4_1),.doutc(w_G2218_0[2]),.din(G2218));
	jspl3 jspl3_w_G2224_0(.douta(w_G2224_0[0]),.doutb(w_G2224_0[1]),.doutc(w_G2224_0[2]),.din(G2224));
	jspl jspl_w_G2224_1(.douta(w_dff_A_hBAC02z23_0),.doutb(w_G2224_1[1]),.din(w_G2224_0[0]));
	jspl3 jspl3_w_G2230_0(.douta(w_G2230_0[0]),.doutb(w_dff_A_cqRjat6f7_1),.doutc(w_G2230_0[2]),.din(G2230));
	jspl3 jspl3_w_G2236_0(.douta(w_G2236_0[0]),.doutb(w_G2236_0[1]),.doutc(w_G2236_0[2]),.din(G2236));
	jspl3 jspl3_w_G2239_0(.douta(w_G2239_0[0]),.doutb(w_G2239_0[1]),.doutc(w_dff_A_LcmCCn9p0_2),.din(G2239));
	jspl jspl_w_G2239_1(.douta(w_G2239_1[0]),.doutb(w_G2239_1[1]),.din(w_G2239_0[0]));
	jspl3 jspl3_w_G2247_0(.douta(w_G2247_0[0]),.doutb(w_G2247_0[1]),.doutc(w_G2247_0[2]),.din(G2247));
	jspl3 jspl3_w_G2253_0(.douta(w_G2253_0[0]),.doutb(w_dff_A_Pn0AJcb18_1),.doutc(w_G2253_0[2]),.din(G2253));
	jspl jspl_w_G2256_0(.douta(w_G2256_0[0]),.doutb(w_G2256_0[1]),.din(G2256));
	jspl jspl_w_G3698_0(.douta(w_G3698_0[0]),.doutb(w_G3698_0[1]),.din(G3698));
	jspl3 jspl3_w_G3701_0(.douta(w_dff_A_Pqsjnv4v5_0),.doutb(w_G3701_0[1]),.doutc(w_G3701_0[2]),.din(G3701));
	jspl jspl_w_G3701_1(.douta(w_G3701_1[0]),.doutb(w_dff_A_8S7dEa0i4_1),.din(w_G3701_0[0]));
	jspl3 jspl3_w_G3705_0(.douta(w_G3705_0[0]),.doutb(w_G3705_0[1]),.doutc(w_dff_A_w8ug4njh8_2),.din(G3705));
	jspl3 jspl3_w_G3705_1(.douta(w_dff_A_4z0juuWj9_0),.doutb(w_G3705_1[1]),.doutc(w_dff_A_YPFFoyh43_2),.din(w_G3705_0[0]));
	jspl jspl_w_G3711_0(.douta(w_G3711_0[0]),.doutb(w_G3711_0[1]),.din(G3711));
	jspl3 jspl3_w_G3717_0(.douta(w_G3717_0[0]),.doutb(w_dff_A_x0EMkzxd8_1),.doutc(w_G3717_0[2]),.din(G3717));
	jspl3 jspl3_w_G3723_0(.douta(w_G3723_0[0]),.doutb(w_dff_A_RgggCuSl6_1),.doutc(w_G3723_0[2]),.din(G3723));
	jspl3 jspl3_w_G3729_0(.douta(w_G3729_0[0]),.doutb(w_G3729_0[1]),.doutc(w_dff_A_Uq2Gp1T96_2),.din(G3729));
	jspl jspl_w_G3729_1(.douta(w_G3729_1[0]),.doutb(w_G3729_1[1]),.din(w_G3729_0[0]));
	jspl3 jspl3_w_G3737_0(.douta(w_G3737_0[0]),.doutb(w_dff_A_wq8328gB9_1),.doutc(w_G3737_0[2]),.din(G3737));
	jspl3 jspl3_w_G3743_0(.douta(w_G3743_0[0]),.doutb(w_dff_A_ggo8CN6V0_1),.doutc(w_G3743_0[2]),.din(G3743));
	jspl3 jspl3_w_G3749_0(.douta(w_G3749_0[0]),.doutb(w_dff_A_zBnmxytd5_1),.doutc(w_G3749_0[2]),.din(G3749));
	jspl jspl_w_G4393_0(.douta(w_G4393_0[0]),.doutb(w_G4393_0[1]),.din(G4393));
	jspl3 jspl3_w_G4394_0(.douta(w_G4394_0[0]),.doutb(w_G4394_0[1]),.doutc(w_dff_A_E5eUml0l6_2),.din(G4394));
	jspl jspl_w_G4394_1(.douta(w_G4394_1[0]),.doutb(w_G4394_1[1]),.din(w_G4394_0[0]));
	jspl3 jspl3_w_G4400_0(.douta(w_G4400_0[0]),.doutb(w_G4400_0[1]),.doutc(w_G4400_0[2]),.din(G4400));
	jspl jspl_w_G4400_1(.douta(w_dff_A_pTOs2fBc6_0),.doutb(w_G4400_1[1]),.din(w_G4400_0[0]));
	jspl3 jspl3_w_G4405_0(.douta(w_G4405_0[0]),.doutb(w_G4405_0[1]),.doutc(w_G4405_0[2]),.din(G4405));
	jspl jspl_w_G4405_1(.douta(w_dff_A_KsBxcwTl2_0),.doutb(w_G4405_1[1]),.din(w_G4405_0[0]));
	jspl3 jspl3_w_G4410_0(.douta(w_G4410_0[0]),.doutb(w_dff_A_RQNKq2ED1_1),.doutc(w_G4410_0[2]),.din(G4410));
	jspl3 jspl3_w_G4415_0(.douta(w_G4415_0[0]),.doutb(w_G4415_0[1]),.doutc(w_G4415_0[2]),.din(G4415));
	jspl jspl_w_G4415_1(.douta(w_dff_A_9AKXfkfi4_0),.doutb(w_G4415_1[1]),.din(w_G4415_0[0]));
	jspl3 jspl3_w_G4420_0(.douta(w_G4420_0[0]),.doutb(w_G4420_0[1]),.doutc(w_G4420_0[2]),.din(G4420));
	jspl jspl_w_G4420_1(.douta(w_dff_A_QOT75w8e3_0),.doutb(w_G4420_1[1]),.din(w_G4420_0[0]));
	jspl3 jspl3_w_G4427_0(.douta(w_G4427_0[0]),.doutb(w_G4427_0[1]),.doutc(w_G4427_0[2]),.din(G4427));
	jspl3 jspl3_w_G4432_0(.douta(w_G4432_0[0]),.doutb(w_dff_A_ttAswpf56_1),.doutc(w_G4432_0[2]),.din(G4432));
	jspl3 jspl3_w_G4437_0(.douta(w_G4437_0[0]),.doutb(w_dff_A_bdb0wrOh4_1),.doutc(w_G4437_0[2]),.din(G4437));
	jspl3 jspl3_w_G4526_0(.douta(w_G4526_0[0]),.doutb(w_dff_A_AAVX09nF5_1),.doutc(w_dff_A_M4E1PaT90_2),.din(G4526));
	jspl3 jspl3_w_G4526_1(.douta(w_dff_A_WgW83LfH5_0),.doutb(w_G4526_1[1]),.doutc(w_dff_A_vIdPQ6qN6_2),.din(w_G4526_0[0]));
	jspl3 jspl3_w_G4526_2(.douta(w_dff_A_eGfvfQ5k5_0),.doutb(w_dff_A_dzxADrtF4_1),.doutc(w_G4526_2[2]),.din(w_G4526_0[1]));
	jspl3 jspl3_w_G4528_0(.douta(w_G4528_0[0]),.doutb(w_G4528_0[1]),.doutc(w_G4528_0[2]),.din(G4528));
	jspl jspl_w_G404_0(.douta(w_G404_0),.doutb(w_dff_A_GynMmCSi4_1),.din(G404_fa_));
	jspl jspl_w_G406_0(.douta(w_G406_0),.doutb(w_dff_A_QtSapZun2_1),.din(G406_fa_));
	jspl jspl_w_G408_0(.douta(w_G408_0),.doutb(w_dff_A_iYRibRUl1_1),.din(G408_fa_));
	jspl jspl_w_G410_0(.douta(w_G410_0),.doutb(w_dff_A_tsINoMcR6_1),.din(G410_fa_));
	jspl jspl_w_G412_0(.douta(w_G412_0),.doutb(w_dff_A_bjP8Gnko9_1),.din(G412_fa_));
	jspl jspl_w_G414_0(.douta(w_dff_A_ERBY7ag16_0),.doutb(w_dff_A_I8w0B8AP8_1),.din(G414_fa_));
	jspl jspl_w_G416_0(.douta(w_G416_0),.doutb(w_dff_A_qkkR41lL2_1),.din(G416_fa_));
	jspl jspl_w_G252_0(.douta(w_G252_0),.doutb(w_dff_A_qDtSjULd9_1),.din(G252_fa_));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(n345));
	jspl jspl_w_n347_0(.douta(w_n347_0[0]),.doutb(w_n347_0[1]),.din(w_dff_B_eVb1uE7h3_2));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl jspl_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.din(n353));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_n354_0[2]),.din(w_dff_B_bRLAOsI35_3));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl3 jspl3_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.doutc(w_n355_1[2]),.din(w_n355_0[0]));
	jspl3 jspl3_w_n355_2(.douta(w_n355_2[0]),.doutb(w_n355_2[1]),.doutc(w_n355_2[2]),.din(w_n355_0[1]));
	jspl3 jspl3_w_n355_3(.douta(w_n355_3[0]),.doutb(w_n355_3[1]),.doutc(w_n355_3[2]),.din(w_n355_0[2]));
	jspl3 jspl3_w_n355_4(.douta(w_n355_4[0]),.doutb(w_n355_4[1]),.doutc(w_n355_4[2]),.din(w_n355_1[0]));
	jspl3 jspl3_w_n355_5(.douta(w_n355_5[0]),.doutb(w_n355_5[1]),.doutc(w_n355_5[2]),.din(w_n355_1[1]));
	jspl3 jspl3_w_n355_6(.douta(w_n355_6[0]),.doutb(w_n355_6[1]),.doutc(w_n355_6[2]),.din(w_n355_1[2]));
	jspl3 jspl3_w_n355_7(.douta(w_n355_7[0]),.doutb(w_n355_7[1]),.doutc(w_n355_7[2]),.din(w_n355_2[0]));
	jspl3 jspl3_w_n355_8(.douta(w_n355_8[0]),.doutb(w_n355_8[1]),.doutc(w_n355_8[2]),.din(w_n355_2[1]));
	jspl3 jspl3_w_n355_9(.douta(w_n355_9[0]),.doutb(w_n355_9[1]),.doutc(w_n355_9[2]),.din(w_n355_2[2]));
	jspl3 jspl3_w_n355_10(.douta(w_n355_10[0]),.doutb(w_n355_10[1]),.doutc(w_n355_10[2]),.din(w_n355_3[0]));
	jspl3 jspl3_w_n355_11(.douta(w_n355_11[0]),.doutb(w_n355_11[1]),.doutc(w_n355_11[2]),.din(w_n355_3[1]));
	jspl3 jspl3_w_n355_12(.douta(w_n355_12[0]),.doutb(w_dff_A_t7Tf8XrA0_1),.doutc(w_n355_12[2]),.din(w_n355_3[2]));
	jspl3 jspl3_w_n355_13(.douta(w_n355_13[0]),.doutb(w_n355_13[1]),.doutc(w_n355_13[2]),.din(w_n355_4[0]));
	jspl3 jspl3_w_n355_14(.douta(w_n355_14[0]),.doutb(w_n355_14[1]),.doutc(w_n355_14[2]),.din(w_n355_4[1]));
	jspl3 jspl3_w_n355_15(.douta(w_n355_15[0]),.doutb(w_n355_15[1]),.doutc(w_n355_15[2]),.din(w_n355_4[2]));
	jspl3 jspl3_w_n355_16(.douta(w_n355_16[0]),.doutb(w_n355_16[1]),.doutc(w_n355_16[2]),.din(w_n355_5[0]));
	jspl3 jspl3_w_n355_17(.douta(w_n355_17[0]),.doutb(w_n355_17[1]),.doutc(w_n355_17[2]),.din(w_n355_5[1]));
	jspl3 jspl3_w_n355_18(.douta(w_n355_18[0]),.doutb(w_n355_18[1]),.doutc(w_n355_18[2]),.din(w_n355_5[2]));
	jspl3 jspl3_w_n355_19(.douta(w_n355_19[0]),.doutb(w_n355_19[1]),.doutc(w_n355_19[2]),.din(w_n355_6[0]));
	jspl3 jspl3_w_n355_20(.douta(w_n355_20[0]),.doutb(w_n355_20[1]),.doutc(w_n355_20[2]),.din(w_n355_6[1]));
	jspl3 jspl3_w_n355_21(.douta(w_n355_21[0]),.doutb(w_n355_21[1]),.doutc(w_n355_21[2]),.din(w_n355_6[2]));
	jspl3 jspl3_w_n355_22(.douta(w_n355_22[0]),.doutb(w_n355_22[1]),.doutc(w_n355_22[2]),.din(w_n355_7[0]));
	jspl3 jspl3_w_n355_23(.douta(w_n355_23[0]),.doutb(w_n355_23[1]),.doutc(w_n355_23[2]),.din(w_n355_7[1]));
	jspl3 jspl3_w_n355_24(.douta(w_n355_24[0]),.doutb(w_n355_24[1]),.doutc(w_n355_24[2]),.din(w_n355_7[2]));
	jspl3 jspl3_w_n355_25(.douta(w_n355_25[0]),.doutb(w_n355_25[1]),.doutc(w_n355_25[2]),.din(w_n355_8[0]));
	jspl3 jspl3_w_n355_26(.douta(w_n355_26[0]),.doutb(w_n355_26[1]),.doutc(w_n355_26[2]),.din(w_n355_8[1]));
	jspl3 jspl3_w_n355_27(.douta(w_n355_27[0]),.doutb(w_n355_27[1]),.doutc(w_n355_27[2]),.din(w_n355_8[2]));
	jspl3 jspl3_w_n355_28(.douta(w_n355_28[0]),.doutb(w_n355_28[1]),.doutc(w_n355_28[2]),.din(w_n355_9[0]));
	jspl3 jspl3_w_n355_29(.douta(w_n355_29[0]),.doutb(w_n355_29[1]),.doutc(w_n355_29[2]),.din(w_n355_9[1]));
	jspl3 jspl3_w_n355_30(.douta(w_n355_30[0]),.doutb(w_n355_30[1]),.doutc(w_n355_30[2]),.din(w_n355_9[2]));
	jspl3 jspl3_w_n355_31(.douta(w_n355_31[0]),.doutb(w_n355_31[1]),.doutc(w_n355_31[2]),.din(w_n355_10[0]));
	jspl3 jspl3_w_n355_32(.douta(w_n355_32[0]),.doutb(w_n355_32[1]),.doutc(w_n355_32[2]),.din(w_n355_10[1]));
	jspl3 jspl3_w_n355_33(.douta(w_n355_33[0]),.doutb(w_n355_33[1]),.doutc(w_n355_33[2]),.din(w_n355_10[2]));
	jspl3 jspl3_w_n355_34(.douta(w_n355_34[0]),.doutb(w_n355_34[1]),.doutc(w_n355_34[2]),.din(w_n355_11[0]));
	jspl3 jspl3_w_n355_35(.douta(w_n355_35[0]),.doutb(w_n355_35[1]),.doutc(w_n355_35[2]),.din(w_n355_11[1]));
	jspl jspl_w_n357_0(.douta(w_dff_A_8u8zz0hI7_0),.doutb(w_n357_0[1]),.din(n357));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(n358));
	jspl3 jspl3_w_n359_0(.douta(w_n359_0[0]),.doutb(w_n359_0[1]),.doutc(w_n359_0[2]),.din(n359));
	jspl jspl_w_n359_1(.douta(w_n359_1[0]),.doutb(w_n359_1[1]),.din(w_n359_0[0]));
	jspl3 jspl3_w_n361_0(.douta(w_dff_A_4pDBzIkj8_0),.doutb(w_n361_0[1]),.doutc(w_n361_0[2]),.din(n361));
	jspl3 jspl3_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.doutc(w_n362_0[2]),.din(n362));
	jspl3 jspl3_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.doutc(w_dff_A_DpxLS1m19_2),.din(w_dff_B_ICQHecuV9_3));
	jspl3 jspl3_w_n364_0(.douta(w_dff_A_XrVfKjOm6_0),.doutb(w_n364_0[1]),.doutc(w_n364_0[2]),.din(n364));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_dff_A_QNIvOtTH5_2),.din(n366));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(n368));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl3 jspl3_w_n370_0(.douta(w_dff_A_2FSUKeD00_0),.doutb(w_dff_A_ehSBP0Yb4_1),.doutc(w_n370_0[2]),.din(w_dff_B_nxbVmBxn9_3));
	jspl3 jspl3_w_n371_0(.douta(w_n371_0[0]),.doutb(w_dff_A_nuxPCBOz4_1),.doutc(w_dff_A_fWSAdVKo6_2),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl3 jspl3_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.doutc(w_n373_0[2]),.din(n373));
	jspl3 jspl3_w_n373_1(.douta(w_n373_1[0]),.doutb(w_n373_1[1]),.doutc(w_n373_1[2]),.din(w_n373_0[0]));
	jspl3 jspl3_w_n373_2(.douta(w_n373_2[0]),.doutb(w_n373_2[1]),.doutc(w_n373_2[2]),.din(w_n373_0[1]));
	jspl3 jspl3_w_n373_3(.douta(w_dff_A_dvAMxUoN8_0),.doutb(w_n373_3[1]),.doutc(w_n373_3[2]),.din(w_n373_0[2]));
	jspl3 jspl3_w_n373_4(.douta(w_n373_4[0]),.doutb(w_n373_4[1]),.doutc(w_n373_4[2]),.din(w_n373_1[0]));
	jspl3 jspl3_w_n373_5(.douta(w_n373_5[0]),.doutb(w_n373_5[1]),.doutc(w_dff_A_8Cb6vKBt0_2),.din(w_n373_1[1]));
	jspl3 jspl3_w_n373_6(.douta(w_n373_6[0]),.doutb(w_n373_6[1]),.doutc(w_n373_6[2]),.din(w_n373_1[2]));
	jspl3 jspl3_w_n373_7(.douta(w_n373_7[0]),.doutb(w_n373_7[1]),.doutc(w_n373_7[2]),.din(w_n373_2[0]));
	jspl3 jspl3_w_n373_8(.douta(w_n373_8[0]),.doutb(w_n373_8[1]),.doutc(w_n373_8[2]),.din(w_n373_2[1]));
	jspl3 jspl3_w_n373_9(.douta(w_n373_9[0]),.doutb(w_n373_9[1]),.doutc(w_n373_9[2]),.din(w_n373_2[2]));
	jspl jspl_w_n374_0(.douta(w_dff_A_tkqNoS2v5_0),.doutb(w_n374_0[1]),.din(n374));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl3 jspl3_w_n377_0(.douta(w_dff_A_t6sCCjTH2_0),.doutb(w_n377_0[1]),.doutc(w_dff_A_idthlT9g4_2),.din(n377));
	jspl3 jspl3_w_n377_1(.douta(w_dff_A_9QatQ9tk9_0),.doutb(w_n377_1[1]),.doutc(w_dff_A_khjwgLvX2_2),.din(w_n377_0[0]));
	jspl jspl_w_n378_0(.douta(w_dff_A_zj7Wtcb85_0),.doutb(w_n378_0[1]),.din(n378));
	jspl3 jspl3_w_n379_0(.douta(w_n379_0[0]),.doutb(w_n379_0[1]),.doutc(w_n379_0[2]),.din(n379));
	jspl jspl_w_n380_0(.douta(w_n380_0[0]),.doutb(w_n380_0[1]),.din(n380));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_dff_A_DY0VH9bL9_1),.doutc(w_dff_A_4u7xADtA8_2),.din(n383));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(w_dff_B_8TkpM3NK2_2));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_n388_0[2]),.din(n388));
	jspl3 jspl3_w_n388_1(.douta(w_dff_A_j3rjMdM79_0),.doutb(w_n388_1[1]),.doutc(w_dff_A_SRJSWJeu4_2),.din(w_n388_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_dff_A_qqy3ED7z2_0),.doutb(w_dff_A_JXnlarNW9_1),.doutc(w_n389_0[2]),.din(n389));
	jspl jspl_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.din(w_n389_0[0]));
	jspl3 jspl3_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.doutc(w_n391_0[2]),.din(n391));
	jspl3 jspl3_w_n392_0(.douta(w_dff_A_wx8BE9BM7_0),.doutb(w_n392_0[1]),.doutc(w_n392_0[2]),.din(n392));
	jspl3 jspl3_w_n393_0(.douta(w_dff_A_BBzGkKiJ5_0),.doutb(w_dff_A_oj1IjktD9_1),.doutc(w_n393_0[2]),.din(n393));
	jspl jspl_w_n393_1(.douta(w_n393_1[0]),.doutb(w_n393_1[1]),.din(w_n393_0[0]));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl3 jspl3_w_n395_0(.douta(w_n395_0[0]),.doutb(w_n395_0[1]),.doutc(w_n395_0[2]),.din(n395));
	jspl jspl_w_n395_1(.douta(w_n395_1[0]),.doutb(w_n395_1[1]),.din(w_n395_0[0]));
	jspl3 jspl3_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.doutc(w_n396_0[2]),.din(n396));
	jspl3 jspl3_w_n396_1(.douta(w_n396_1[0]),.doutb(w_n396_1[1]),.doutc(w_n396_1[2]),.din(w_n396_0[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl3 jspl3_w_n405_0(.douta(w_dff_A_0KsNRUZ00_0),.doutb(w_dff_A_nsaHze9V0_1),.doutc(w_n405_0[2]),.din(n405));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl3 jspl3_w_n409_0(.douta(w_n409_0[0]),.doutb(w_n409_0[1]),.doutc(w_dff_A_Amuwpa848_2),.din(n409));
	jspl jspl_w_n409_1(.douta(w_n409_1[0]),.doutb(w_n409_1[1]),.din(w_n409_0[0]));
	jspl3 jspl3_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.doutc(w_dff_A_C5SgrmPL0_2),.din(n411));
	jspl jspl_w_n411_1(.douta(w_n411_1[0]),.doutb(w_n411_1[1]),.din(w_n411_0[0]));
	jspl3 jspl3_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.doutc(w_n413_0[2]),.din(n413));
	jspl jspl_w_n413_1(.douta(w_dff_A_msS3zn0b7_0),.doutb(w_n413_1[1]),.din(w_n413_0[0]));
	jspl3 jspl3_w_n414_0(.douta(w_n414_0[0]),.doutb(w_dff_A_qWKx2dOq8_1),.doutc(w_n414_0[2]),.din(n414));
	jspl jspl_w_n414_1(.douta(w_n414_1[0]),.doutb(w_n414_1[1]),.din(w_n414_0[0]));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl3 jspl3_w_n416_0(.douta(w_n416_0[0]),.doutb(w_dff_A_1zVdYsML7_1),.doutc(w_n416_0[2]),.din(n416));
	jspl jspl_w_n418_0(.douta(w_dff_A_iWAGMO7h6_0),.doutb(w_n418_0[1]),.din(n418));
	jspl jspl_w_n419_0(.douta(w_n419_0[0]),.doutb(w_dff_A_StSoeVLD8_1),.din(n419));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_dff_A_keEUnYQ00_1),.din(n420));
	jspl3 jspl3_w_n421_0(.douta(w_n421_0[0]),.doutb(w_dff_A_J5y6YU0r4_1),.doutc(w_dff_A_fzPZDmtX3_2),.din(n421));
	jspl jspl_w_n422_0(.douta(w_dff_A_3oLcbMUW2_0),.doutb(w_n422_0[1]),.din(n422));
	jspl3 jspl3_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.doutc(w_n423_0[2]),.din(n423));
	jspl jspl_w_n424_0(.douta(w_n424_0[0]),.doutb(w_dff_A_6GHje0Ez4_1),.din(n424));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_dff_A_wqPvJ2r96_2),.din(n425));
	jspl jspl_w_n425_1(.douta(w_n425_1[0]),.doutb(w_dff_A_fHouZqGt3_1),.din(w_n425_0[0]));
	jspl3 jspl3_w_n426_0(.douta(w_n426_0[0]),.doutb(w_dff_A_Ggj1yM443_1),.doutc(w_dff_A_K5ZBCKeC9_2),.din(n426));
	jspl jspl_w_n427_0(.douta(w_dff_A_Etqypq3F7_0),.doutb(w_n427_0[1]),.din(n427));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.doutc(w_n428_0[2]),.din(n428));
	jspl3 jspl3_w_n429_0(.douta(w_n429_0[0]),.doutb(w_dff_A_YUTW2DAO3_1),.doutc(w_dff_A_9gVNd9nX7_2),.din(n429));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(w_dff_B_qfxNow3q4_2));
	jspl jspl_w_n431_0(.douta(w_dff_A_rZYiXbkz5_0),.doutb(w_n431_0[1]),.din(n431));
	jspl3 jspl3_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.doutc(w_n432_0[2]),.din(n432));
	jspl3 jspl3_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.doutc(w_dff_A_ky3EWdLW5_2),.din(n433));
	jspl3 jspl3_w_n433_1(.douta(w_dff_A_OuOmfGs39_0),.doutb(w_n433_1[1]),.doutc(w_n433_1[2]),.din(w_n433_0[0]));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(w_dff_B_59IVopTg7_2));
	jspl jspl_w_n435_0(.douta(w_dff_A_Dxy3LhG70_0),.doutb(w_n435_0[1]),.din(n435));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n437_0(.douta(w_n437_0[0]),.doutb(w_dff_A_R1lrvgxA0_1),.doutc(w_n437_0[2]),.din(n437));
	jspl jspl_w_n438_0(.douta(w_dff_A_b9i0mVPX4_0),.doutb(w_n438_0[1]),.din(n438));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl3 jspl3_w_n444_0(.douta(w_n444_0[0]),.doutb(w_dff_A_mfUBjL8h2_1),.doutc(w_dff_A_jGvha8wF0_2),.din(n444));
	jspl3 jspl3_w_n445_0(.douta(w_n445_0[0]),.doutb(w_dff_A_nRvZGQid1_1),.doutc(w_n445_0[2]),.din(n445));
	jspl3 jspl3_w_n447_0(.douta(w_n447_0[0]),.doutb(w_dff_A_DBXmQNFG7_1),.doutc(w_n447_0[2]),.din(n447));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl jspl_w_n449_1(.douta(w_dff_A_YDSTlRFl9_0),.doutb(w_n449_1[1]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n450_0(.douta(w_n450_0[0]),.doutb(w_n450_0[1]),.doutc(w_dff_A_yOGMEFVi3_2),.din(n450));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_n451_0[1]),.doutc(w_n451_0[2]),.din(w_dff_B_ZTy8EqPV4_3));
	jspl3 jspl3_w_n453_0(.douta(w_n453_0[0]),.doutb(w_dff_A_tqesnuAW6_1),.doutc(w_n453_0[2]),.din(n453));
	jspl jspl_w_n453_1(.douta(w_n453_1[0]),.doutb(w_n453_1[1]),.din(w_n453_0[0]));
	jspl3 jspl3_w_n456_0(.douta(w_n456_0[0]),.doutb(w_dff_A_JnxynNQZ7_1),.doutc(w_dff_A_fzA0RuAB8_2),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.doutc(w_n459_0[2]),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_dff_A_ELfZLHUX2_1),.doutc(w_dff_A_9WxyhcV15_2),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_dff_A_wPtHeeCc1_0),.doutb(w_dff_A_6Hqpq9og1_1),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_X9cBIOx54_1),.doutc(w_dff_A_l6iDbYvx2_2),.din(n462));
	jspl3 jspl3_w_n463_0(.douta(w_n463_0[0]),.doutb(w_dff_A_QVBtoqvc1_1),.doutc(w_dff_A_iJUqX09N6_2),.din(n463));
	jspl jspl_w_n463_1(.douta(w_dff_A_NO57E4si4_0),.doutb(w_n463_1[1]),.din(w_n463_0[0]));
	jspl3 jspl3_w_n464_0(.douta(w_n464_0[0]),.doutb(w_dff_A_4UQNzWyN7_1),.doutc(w_n464_0[2]),.din(n464));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_dff_A_cjpTw9ug5_1),.din(w_dff_B_La6GKKE27_2));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(w_dff_B_JpelzHeC9_2));
	jspl jspl_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.din(n467));
	jspl3 jspl3_w_n469_0(.douta(w_n469_0[0]),.doutb(w_dff_A_u8HoK95L0_1),.doutc(w_n469_0[2]),.din(n469));
	jspl jspl_w_n469_1(.douta(w_n469_1[0]),.doutb(w_n469_1[1]),.din(w_n469_0[0]));
	jspl3 jspl3_w_n470_0(.douta(w_n470_0[0]),.doutb(w_dff_A_5A8AnfSW3_1),.doutc(w_dff_A_PvTO2xKm6_2),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_dff_A_KfIMhN2W7_1),.doutc(w_dff_A_vtutKMai1_2),.din(n471));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl3 jspl3_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.doutc(w_n474_0[2]),.din(n474));
	jspl3 jspl3_w_n475_0(.douta(w_n475_0[0]),.doutb(w_dff_A_mti1uzGy6_1),.doutc(w_n475_0[2]),.din(n475));
	jspl3 jspl3_w_n476_0(.douta(w_n476_0[0]),.doutb(w_dff_A_kyLWR7fF2_1),.doutc(w_dff_A_O9ZEuD0F3_2),.din(n476));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl3 jspl3_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.doutc(w_n479_0[2]),.din(n479));
	jspl jspl_w_n479_1(.douta(w_n479_1[0]),.doutb(w_n479_1[1]),.din(w_n479_0[0]));
	jspl3 jspl3_w_n480_0(.douta(w_n480_0[0]),.doutb(w_n480_0[1]),.doutc(w_dff_A_oyn8YtEy2_2),.din(n480));
	jspl jspl_w_n480_1(.douta(w_n480_1[0]),.doutb(w_n480_1[1]),.din(w_n480_0[0]));
	jspl jspl_w_n481_0(.douta(w_dff_A_NTePZsvj2_0),.doutb(w_n481_0[1]),.din(n481));
	jspl jspl_w_n485_0(.douta(w_n485_0[0]),.doutb(w_n485_0[1]),.din(n485));
	jspl jspl_w_n486_0(.douta(w_n486_0[0]),.doutb(w_n486_0[1]),.din(n486));
	jspl3 jspl3_w_n487_0(.douta(w_n487_0[0]),.doutb(w_dff_A_JIc1SOCK2_1),.doutc(w_n487_0[2]),.din(n487));
	jspl3 jspl3_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.doutc(w_n489_0[2]),.din(n489));
	jspl3 jspl3_w_n491_0(.douta(w_n491_0[0]),.doutb(w_n491_0[1]),.doutc(w_dff_A_8J2edwd05_2),.din(n491));
	jspl jspl_w_n491_1(.douta(w_dff_A_heQPLmxD8_0),.doutb(w_n491_1[1]),.din(w_n491_0[0]));
	jspl3 jspl3_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.doutc(w_n495_0[2]),.din(n495));
	jspl jspl_w_n495_1(.douta(w_dff_A_U03xe2o77_0),.doutb(w_n495_1[1]),.din(w_n495_0[0]));
	jspl3 jspl3_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.doutc(w_n496_0[2]),.din(n496));
	jspl3 jspl3_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.doutc(w_n497_0[2]),.din(n497));
	jspl jspl_w_n497_1(.douta(w_dff_A_IHcVICTS5_0),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_dff_A_YKcXgaSB9_1),.din(n499));
	jspl jspl_w_n500_0(.douta(w_n500_0[0]),.doutb(w_dff_A_AJ2RaLHq2_1),.din(n500));
	jspl3 jspl3_w_n501_0(.douta(w_dff_A_KG5akhGz9_0),.doutb(w_n501_0[1]),.doutc(w_dff_A_qIxN32vE1_2),.din(n501));
	jspl jspl_w_n503_0(.douta(w_n503_0[0]),.doutb(w_n503_0[1]),.din(n503));
	jspl3 jspl3_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.doutc(w_dff_A_FmgsxsHO6_2),.din(n504));
	jspl jspl_w_n504_1(.douta(w_n504_1[0]),.doutb(w_n504_1[1]),.din(w_n504_0[0]));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_dff_A_RxW72wH48_1),.din(n505));
	jspl jspl_w_n507_0(.douta(w_dff_A_nQGtR75U2_0),.doutb(w_n507_0[1]),.din(n507));
	jspl3 jspl3_w_n509_0(.douta(w_n509_0[0]),.doutb(w_dff_A_ze2TbJmO2_1),.doutc(w_dff_A_DSMLlou83_2),.din(n509));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl3 jspl3_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.doutc(w_n512_0[2]),.din(n512));
	jspl3 jspl3_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.doutc(w_dff_A_VgXoLfYa4_2),.din(n513));
	jspl jspl_w_n513_1(.douta(w_n513_1[0]),.doutb(w_dff_A_6rMMNjas3_1),.din(w_n513_0[0]));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(w_dff_B_o50higMX4_2));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl3 jspl3_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.doutc(w_n517_0[2]),.din(n517));
	jspl jspl_w_n517_1(.douta(w_n517_1[0]),.doutb(w_n517_1[1]),.din(w_n517_0[0]));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl3 jspl3_w_n518_1(.douta(w_dff_A_lCny2K5N7_0),.doutb(w_n518_1[1]),.doutc(w_n518_1[2]),.din(w_n518_0[0]));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(w_dff_B_s3BtrIMB0_2));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.doutc(w_n523_0[2]),.din(n523));
	jspl3 jspl3_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.doutc(w_n524_0[2]),.din(n524));
	jspl3 jspl3_w_n524_1(.douta(w_n524_1[0]),.doutb(w_n524_1[1]),.doutc(w_dff_A_rPeFpmjZ9_2),.din(w_n524_0[0]));
	jspl3 jspl3_w_n526_0(.douta(w_dff_A_gcnzPzKn1_0),.doutb(w_dff_A_xxYf9NAS1_1),.doutc(w_n526_0[2]),.din(n526));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(w_dff_B_6kXN9UvO1_2));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(n530));
	jspl3 jspl3_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.doutc(w_n531_0[2]),.din(n531));
	jspl jspl_w_n531_1(.douta(w_n531_1[0]),.doutb(w_n531_1[1]),.din(w_n531_0[0]));
	jspl3 jspl3_w_n536_0(.douta(w_n536_0[0]),.doutb(w_dff_A_hOgeOUPF7_1),.doutc(w_dff_A_iC5C8OjB4_2),.din(n536));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl3 jspl3_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.doutc(w_n539_0[2]),.din(n539));
	jspl jspl_w_n539_1(.douta(w_n539_1[0]),.doutb(w_n539_1[1]),.din(w_n539_0[0]));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(w_dff_B_JLLYtHSi6_2));
	jspl jspl_w_n546_0(.douta(w_n546_0[0]),.doutb(w_n546_0[1]),.din(n546));
	jspl3 jspl3_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.doutc(w_n547_0[2]),.din(n547));
	jspl jspl_w_n547_1(.douta(w_n547_1[0]),.doutb(w_n547_1[1]),.din(w_n547_0[0]));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_dff_A_3WoZ6Qs11_1),.din(n548));
	jspl jspl_w_n550_0(.douta(w_dff_A_HAQrLaVw1_0),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(w_dff_B_o3YYZP3c6_2));
	jspl jspl_w_n554_0(.douta(w_n554_0[0]),.doutb(w_n554_0[1]),.din(n554));
	jspl3 jspl3_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.doutc(w_n555_0[2]),.din(n555));
	jspl jspl_w_n555_1(.douta(w_n555_1[0]),.doutb(w_n555_1[1]),.din(w_n555_0[0]));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_dff_A_oQuHNRS80_1),.doutc(w_dff_A_dGv0HnBV7_2),.din(n556));
	jspl jspl_w_n558_0(.douta(w_dff_A_9H7CSzP19_0),.doutb(w_n558_0[1]),.din(n558));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(w_dff_B_mbNgPm2M9_2));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.doutc(w_n563_0[2]),.din(n563));
	jspl jspl_w_n563_1(.douta(w_n563_1[0]),.doutb(w_n563_1[1]),.din(w_n563_0[0]));
	jspl3 jspl3_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_hFM6fXmV7_1),.doutc(w_dff_A_md8RtMPF9_2),.din(n564));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl3 jspl3_w_n566_0(.douta(w_dff_A_TRgHmW7P3_0),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.doutc(w_n568_0[2]),.din(n568));
	jspl3 jspl3_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.doutc(w_n570_0[2]),.din(n570));
	jspl3 jspl3_w_n570_1(.douta(w_n570_1[0]),.doutb(w_dff_A_a2DMK6Mh4_1),.doutc(w_n570_1[2]),.din(w_n570_0[0]));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl jspl_w_n572_1(.douta(w_n572_1[0]),.doutb(w_dff_A_qmdxOz5k3_1),.din(w_n572_0[0]));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_dff_A_zkIvd3R72_1),.doutc(w_dff_A_Pvhb6ZV98_2),.din(w_dff_B_w0b9mGea6_3));
	jspl jspl_w_n573_1(.douta(w_dff_A_hguD7QRp5_0),.doutb(w_n573_1[1]),.din(w_n573_0[0]));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_dff_A_XafuP8tA7_1),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.doutc(w_dff_A_vgM6wKl89_2),.din(n575));
	jspl jspl_w_n575_1(.douta(w_dff_A_834GmKxn6_0),.doutb(w_n575_1[1]),.din(w_n575_0[0]));
	jspl3 jspl3_w_n576_0(.douta(w_dff_A_LqCO2wEt1_0),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_dff_A_m1xlhcAx1_0),.doutb(w_dff_A_Jy21ZVUD4_1),.doutc(w_n578_0[2]),.din(n578));
	jspl3 jspl3_w_n580_0(.douta(w_dff_A_IYP4Qtpr2_0),.doutb(w_dff_A_nSimRdzg0_1),.doutc(w_n580_0[2]),.din(n580));
	jspl3 jspl3_w_n581_0(.douta(w_dff_A_ljIFcQ6O6_0),.doutb(w_n581_0[1]),.doutc(w_dff_A_2EevMicO9_2),.din(n581));
	jspl3 jspl3_w_n582_0(.douta(w_dff_A_bSEYi0OK8_0),.doutb(w_n582_0[1]),.doutc(w_dff_A_ouNZOQcj1_2),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl3 jspl3_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.doutc(w_n585_0[2]),.din(n585));
	jspl jspl_w_n585_1(.douta(w_n585_1[0]),.doutb(w_n585_1[1]),.din(w_n585_0[0]));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_dff_A_UOjkKZjf8_1),.doutc(w_dff_A_Jif3DlyP9_2),.din(n586));
	jspl jspl_w_n588_0(.douta(w_dff_A_I8ZCmTMw6_0),.doutb(w_n588_0[1]),.din(n588));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_dff_A_9ZEcId8N2_1),.doutc(w_dff_A_agWuWEKK0_2),.din(n590));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(n592));
	jspl3 jspl3_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.doutc(w_n593_0[2]),.din(n593));
	jspl jspl_w_n593_1(.douta(w_n593_1[0]),.doutb(w_n593_1[1]),.din(w_n593_0[0]));
	jspl3 jspl3_w_n594_0(.douta(w_n594_0[0]),.doutb(w_dff_A_kmmA1FoC8_1),.doutc(w_dff_A_R7HIKgfX4_2),.din(n594));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_dff_A_hKABPv192_1),.doutc(w_dff_A_OtRZhWkL0_2),.din(n595));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl3 jspl3_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.doutc(w_n598_0[2]),.din(n598));
	jspl jspl_w_n598_1(.douta(w_n598_1[0]),.doutb(w_n598_1[1]),.din(w_n598_0[0]));
	jspl3 jspl3_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.doutc(w_n599_0[2]),.din(n599));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(w_dff_B_BXVAVGHI5_2));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.doutc(w_n603_0[2]),.din(n603));
	jspl jspl_w_n603_1(.douta(w_n603_1[0]),.doutb(w_n603_1[1]),.din(w_n603_0[0]));
	jspl jspl_w_n604_0(.douta(w_dff_A_eybIkGQx0_0),.doutb(w_n604_0[1]),.din(n604));
	jspl3 jspl3_w_n605_0(.douta(w_dff_A_tPE7GcZP7_0),.doutb(w_dff_A_0KXMix2R7_1),.doutc(w_n605_0[2]),.din(n605));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_dff_A_PWYghY9h1_1),.din(w_dff_B_tJHYdyLG7_2));
	jspl jspl_w_n610_0(.douta(w_dff_A_iag1hkad3_0),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_dff_A_NJ16sLVB1_1),.din(n612));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n615_0(.douta(w_n615_0[0]),.doutb(w_dff_A_6QjljWL94_1),.doutc(w_n615_0[2]),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl3 jspl3_w_n618_0(.douta(w_dff_A_4HO5pGpq3_0),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_dff_A_9j1YVS9y4_1),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_dff_A_Ovq9bdPh2_1),.doutc(w_dff_A_erNsfYQU8_2),.din(n622));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n625_1(.douta(w_n625_1[0]),.doutb(w_n625_1[1]),.din(w_n625_0[0]));
	jspl3 jspl3_w_n626_0(.douta(w_dff_A_3kVY6l0E9_0),.doutb(w_dff_A_wND6vBd05_1),.doutc(w_n626_0[2]),.din(n626));
	jspl jspl_w_n626_1(.douta(w_dff_A_Gs5W5Cso5_0),.doutb(w_n626_1[1]),.din(w_n626_0[0]));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_dff_A_imEWMNjW5_1),.doutc(w_dff_A_woTKomL55_2),.din(n627));
	jspl jspl_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.din(n629));
	jspl3 jspl3_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.doutc(w_n630_0[2]),.din(n630));
	jspl3 jspl3_w_n631_0(.douta(w_n631_0[0]),.doutb(w_dff_A_tikeZxdx1_1),.doutc(w_dff_A_FSv2gqVb9_2),.din(n631));
	jspl3 jspl3_w_n632_0(.douta(w_dff_A_oKX0JHAy5_0),.doutb(w_n632_0[1]),.doutc(w_dff_A_nAx8PBdD7_2),.din(n632));
	jspl jspl_w_n632_1(.douta(w_n632_1[0]),.doutb(w_n632_1[1]),.din(w_n632_0[0]));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n635_1(.douta(w_n635_1[0]),.doutb(w_n635_1[1]),.din(w_n635_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_dff_A_gg61SxAS4_1),.doutc(w_dff_A_fEUrzPyw6_2),.din(n636));
	jspl3 jspl3_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.doutc(w_n641_0[2]),.din(n641));
	jspl3 jspl3_w_n642_0(.douta(w_n642_0[0]),.doutb(w_dff_A_VjQZaMGs4_1),.doutc(w_n642_0[2]),.din(w_dff_B_NUMZYu669_3));
	jspl jspl_w_n644_0(.douta(w_n644_0[0]),.doutb(w_n644_0[1]),.din(n644));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n646_0(.douta(w_n646_0[0]),.doutb(w_dff_A_Xub83BwO5_1),.din(n646));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_dff_A_wGTAaL9u6_1),.din(n647));
	jspl jspl_w_n649_0(.douta(w_dff_A_9aQUFTwP0_0),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.din(n651));
	jspl jspl_w_n652_0(.douta(w_dff_A_nJFI4ewU7_0),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n653_0(.douta(w_dff_A_UjSvI0Ny8_0),.doutb(w_n653_0[1]),.din(w_dff_B_aEhxahxj8_2));
	jspl3 jspl3_w_n654_0(.douta(w_n654_0[0]),.doutb(w_dff_A_ce8Cg8FA8_1),.doutc(w_dff_A_zA6O4Agt9_2),.din(n654));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_dff_A_PDijplF23_1),.din(n655));
	jspl jspl_w_n656_0(.douta(w_n656_0[0]),.doutb(w_dff_A_bU3HxgH34_1),.din(n656));
	jspl3 jspl3_w_n657_0(.douta(w_n657_0[0]),.doutb(w_dff_A_A1OPI00p8_1),.doutc(w_dff_A_2GrllwjR3_2),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_n660_0[2]),.din(n660));
	jspl3 jspl3_w_n661_0(.douta(w_n661_0[0]),.doutb(w_dff_A_kXj7iwpq7_1),.doutc(w_dff_A_yUGoHWWg2_2),.din(n661));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_dff_A_UqyDJu4D5_1),.din(n662));
	jspl3 jspl3_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.doutc(w_n663_0[2]),.din(n663));
	jspl jspl_w_n663_1(.douta(w_n663_1[0]),.doutb(w_n663_1[1]),.din(w_n663_0[0]));
	jspl jspl_w_n664_0(.douta(w_dff_A_nBMtiG5B5_0),.doutb(w_n664_0[1]),.din(w_dff_B_eLWVEYyq7_2));
	jspl jspl_w_n666_0(.douta(w_dff_A_Bwoqm0jQ7_0),.doutb(w_n666_0[1]),.din(n666));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(n669));
	jspl jspl_w_n671_0(.douta(w_n671_0[0]),.doutb(w_n671_0[1]),.din(n671));
	jspl3 jspl3_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.doutc(w_n673_0[2]),.din(n673));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(n674));
	jspl3 jspl3_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.doutc(w_n676_0[2]),.din(n676));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl3 jspl3_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.doutc(w_n680_0[2]),.din(n680));
	jspl3 jspl3_w_n680_1(.douta(w_n680_1[0]),.doutb(w_n680_1[1]),.doutc(w_n680_1[2]),.din(w_n680_0[0]));
	jspl3 jspl3_w_n680_2(.douta(w_n680_2[0]),.doutb(w_n680_2[1]),.doutc(w_n680_2[2]),.din(w_n680_0[1]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n687_0(.douta(w_dff_A_Sv7nSz9l8_0),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_dff_A_9ccwibTO2_1),.din(w_dff_B_xsOrJPyQ6_2));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_dff_A_RF0FdYnX6_0),.doutb(w_n694_0[1]),.din(n694));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n696_0(.douta(w_dff_A_b1VtYyyq2_0),.doutb(w_n696_0[1]),.din(n696));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(n698));
	jspl3 jspl3_w_n700_0(.douta(w_n700_0[0]),.doutb(w_n700_0[1]),.doutc(w_n700_0[2]),.din(n700));
	jspl jspl_w_n700_1(.douta(w_n700_1[0]),.doutb(w_n700_1[1]),.din(w_n700_0[0]));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl3 jspl3_w_n703_1(.douta(w_n703_1[0]),.doutb(w_n703_1[1]),.doutc(w_n703_1[2]),.din(w_n703_0[0]));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.doutc(w_n707_0[2]),.din(n707));
	jspl3 jspl3_w_n707_1(.douta(w_n707_1[0]),.doutb(w_n707_1[1]),.doutc(w_n707_1[2]),.din(w_n707_0[0]));
	jspl3 jspl3_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.doutc(w_n709_0[2]),.din(n709));
	jspl jspl_w_n709_1(.douta(w_n709_1[0]),.doutb(w_n709_1[1]),.din(w_n709_0[0]));
	jspl3 jspl3_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.doutc(w_n711_0[2]),.din(n711));
	jspl jspl_w_n711_1(.douta(w_n711_1[0]),.doutb(w_n711_1[1]),.din(w_n711_0[0]));
	jspl3 jspl3_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.doutc(w_n712_0[2]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_dff_A_1NxDNOAD3_0),.doutb(w_n713_0[1]),.din(n713));
	jspl3 jspl3_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.doutc(w_n715_0[2]),.din(w_dff_B_jHOlOr462_3));
	jspl jspl_w_n715_1(.douta(w_n715_1[0]),.doutb(w_n715_1[1]),.din(w_n715_0[0]));
	jspl3 jspl3_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.doutc(w_n718_0[2]),.din(w_dff_B_47SaYpgW2_3));
	jspl jspl_w_n719_0(.douta(w_dff_A_2hx7wOQO9_0),.doutb(w_n719_0[1]),.din(n719));
	jspl3 jspl3_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.doutc(w_n720_0[2]),.din(n720));
	jspl3 jspl3_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.doutc(w_n723_0[2]),.din(n723));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_dff_A_lttAXzVh7_1),.din(n724));
	jspl jspl_w_n725_0(.douta(w_dff_A_PpFG70SJ1_0),.doutb(w_n725_0[1]),.din(n725));
	jspl3 jspl3_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.doutc(w_n726_0[2]),.din(n726));
	jspl jspl_w_n726_1(.douta(w_n726_1[0]),.doutb(w_n726_1[1]),.din(w_n726_0[0]));
	jspl3 jspl3_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.doutc(w_n729_0[2]),.din(n729));
	jspl jspl_w_n729_1(.douta(w_n729_1[0]),.doutb(w_n729_1[1]),.din(w_n729_0[0]));
	jspl3 jspl3_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.doutc(w_n734_0[2]),.din(n734));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl3 jspl3_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl jspl_w_n737_1(.douta(w_n737_1[0]),.doutb(w_n737_1[1]),.din(w_n737_0[0]));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n741_1(.douta(w_n741_1[0]),.doutb(w_n741_1[1]),.din(w_n741_0[0]));
	jspl jspl_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.din(n743));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_n744_0[2]),.din(n744));
	jspl3 jspl3_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.doutc(w_n747_0[2]),.din(n747));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(n749));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl3 jspl3_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.doutc(w_n755_0[2]),.din(n755));
	jspl jspl_w_n755_1(.douta(w_n755_1[0]),.doutb(w_n755_1[1]),.din(w_n755_0[0]));
	jspl3 jspl3_w_n758_0(.douta(w_n758_0[0]),.doutb(w_n758_0[1]),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n758_1(.douta(w_n758_1[0]),.doutb(w_n758_1[1]),.din(w_n758_0[0]));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl3 jspl3_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.doutc(w_n761_0[2]),.din(n761));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_n764_0[2]),.din(n764));
	jspl jspl_w_n766_0(.douta(w_n766_0[0]),.doutb(w_n766_0[1]),.din(w_dff_B_9uMlF7Ay0_2));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl3 jspl3_w_n768_0(.douta(w_n768_0[0]),.doutb(w_n768_0[1]),.doutc(w_n768_0[2]),.din(n768));
	jspl3 jspl3_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.doutc(w_n772_0[2]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_dff_A_hL4QtHdo2_1),.din(n773));
	jspl jspl_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.din(n774));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl3 jspl3_w_n776_0(.douta(w_n776_0[0]),.doutb(w_n776_0[1]),.doutc(w_n776_0[2]),.din(n776));
	jspl3 jspl3_w_n780_0(.douta(w_dff_A_RwjGpHMx3_0),.doutb(w_n780_0[1]),.doutc(w_n780_0[2]),.din(n780));
	jspl jspl_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.din(n781));
	jspl3 jspl3_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.doutc(w_n796_0[2]),.din(n796));
	jspl jspl_w_n796_1(.douta(w_n796_1[0]),.doutb(w_n796_1[1]),.din(w_n796_0[0]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.doutc(w_n800_0[2]),.din(n800));
	jspl jspl_w_n800_1(.douta(w_n800_1[0]),.doutb(w_n800_1[1]),.din(w_n800_0[0]));
	jspl3 jspl3_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.doutc(w_n803_0[2]),.din(n803));
	jspl3 jspl3_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.doutc(w_n806_0[2]),.din(n806));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_dff_A_K0UyC9ij2_1),.din(n808));
	jspl3 jspl3_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.doutc(w_n810_0[2]),.din(n810));
	jspl jspl_w_n810_1(.douta(w_n810_1[0]),.doutb(w_n810_1[1]),.din(w_n810_0[0]));
	jspl3 jspl3_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.doutc(w_n814_0[2]),.din(n814));
	jspl jspl_w_n814_1(.douta(w_n814_1[0]),.doutb(w_n814_1[1]),.din(w_n814_0[0]));
	jspl3 jspl3_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.doutc(w_n817_0[2]),.din(n817));
	jspl3 jspl3_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.doutc(w_n820_0[2]),.din(n820));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(n822));
	jspl3 jspl3_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.doutc(w_n824_0[2]),.din(n824));
	jspl3 jspl3_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.doutc(w_n827_0[2]),.din(n827));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_dff_A_9BgNPRCU5_1),.doutc(w_n845_0[2]),.din(n845));
	jspl jspl_w_n845_1(.douta(w_n845_1[0]),.doutb(w_n845_1[1]),.din(w_n845_0[0]));
	jspl3 jspl3_w_n848_0(.douta(w_n848_0[0]),.doutb(w_n848_0[1]),.doutc(w_n848_0[2]),.din(n848));
	jspl jspl_w_n848_1(.douta(w_n848_1[0]),.doutb(w_n848_1[1]),.din(w_n848_0[0]));
	jspl3 jspl3_w_n851_0(.douta(w_n851_0[0]),.doutb(w_n851_0[1]),.doutc(w_n851_0[2]),.din(n851));
	jspl3 jspl3_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.doutc(w_n854_0[2]),.din(n854));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_dff_A_RuXzwzZo6_1),.din(n856));
	jspl3 jspl3_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.doutc(w_n858_0[2]),.din(n858));
	jspl3 jspl3_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.doutc(w_n862_0[2]),.din(n862));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_dff_A_Ig6Jd2UU0_1),.din(n863));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl3 jspl3_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.doutc(w_n866_0[2]),.din(n866));
	jspl3 jspl3_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.doutc(w_n870_0[2]),.din(n870));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl3 jspl3_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.doutc(w_n885_0[2]),.din(n885));
	jspl3 jspl3_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.doutc(w_n888_0[2]),.din(n888));
	jspl3 jspl3_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.doutc(w_n891_0[2]),.din(n891));
	jspl3 jspl3_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.doutc(w_n894_0[2]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_dff_A_fwEvooYQ0_0),.doutb(w_n895_0[1]),.din(n895));
	jspl3 jspl3_w_n900_0(.douta(w_n900_0[0]),.doutb(w_n900_0[1]),.doutc(w_n900_0[2]),.din(n900));
	jspl3 jspl3_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.doutc(w_n903_0[2]),.din(n903));
	jspl jspl_w_n905_0(.douta(w_dff_A_rNjZUdEz4_0),.doutb(w_n905_0[1]),.din(n905));
	jspl3 jspl3_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.doutc(w_n916_0[2]),.din(n916));
	jspl3 jspl3_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.doutc(w_n919_0[2]),.din(n919));
	jspl3 jspl3_w_n926_0(.douta(w_dff_A_ZFgUO11s5_0),.doutb(w_n926_0[1]),.doutc(w_n926_0[2]),.din(n926));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_n930_0[2]),.din(n930));
	jspl3 jspl3_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.doutc(w_n935_0[2]),.din(n935));
	jspl3 jspl3_w_n938_0(.douta(w_dff_A_6HllCUn99_0),.doutb(w_n938_0[1]),.doutc(w_n938_0[2]),.din(n938));
	jspl3 jspl3_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.doutc(w_n944_0[2]),.din(n944));
	jspl3 jspl3_w_n947_0(.douta(w_n947_0[0]),.doutb(w_n947_0[1]),.doutc(w_n947_0[2]),.din(n947));
	jspl3 jspl3_w_n950_0(.douta(w_n950_0[0]),.doutb(w_n950_0[1]),.doutc(w_n950_0[2]),.din(n950));
	jspl jspl_w_n950_1(.douta(w_n950_1[0]),.doutb(w_n950_1[1]),.din(w_n950_0[0]));
	jspl3 jspl3_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.doutc(w_n953_0[2]),.din(n953));
	jspl jspl_w_n953_1(.douta(w_n953_1[0]),.doutb(w_n953_1[1]),.din(w_n953_0[0]));
	jspl3 jspl3_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.doutc(w_n966_0[2]),.din(n966));
	jspl3 jspl3_w_n970_0(.douta(w_n970_0[0]),.doutb(w_n970_0[1]),.doutc(w_n970_0[2]),.din(n970));
	jspl3 jspl3_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.doutc(w_n973_0[2]),.din(n973));
	jspl jspl_w_n973_1(.douta(w_n973_1[0]),.doutb(w_n973_1[1]),.din(w_n973_0[0]));
	jspl3 jspl3_w_n977_0(.douta(w_n977_0[0]),.doutb(w_n977_0[1]),.doutc(w_n977_0[2]),.din(n977));
	jspl jspl_w_n977_1(.douta(w_n977_1[0]),.doutb(w_n977_1[1]),.din(w_n977_0[0]));
	jspl3 jspl3_w_n980_0(.douta(w_n980_0[0]),.doutb(w_n980_0[1]),.doutc(w_n980_0[2]),.din(n980));
	jspl3 jspl3_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.doutc(w_n983_0[2]),.din(n983));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_dff_A_RhqxIhuS9_1),.din(w_dff_B_83cBPOSs0_2));
	jspl3 jspl3_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.doutc(w_n987_0[2]),.din(n987));
	jspl3 jspl3_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.doutc(w_n991_0[2]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl3 jspl3_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.doutc(w_n995_0[2]),.din(n995));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.doutc(w_n999_0[2]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_dff_A_N3BsIWX12_1),.din(n1000));
	jspl jspl_w_n1003_0(.douta(w_dff_A_ezWMIB7q9_0),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_dff_A_A4sJ5E0u2_0),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1042_0(.douta(w_dff_A_etnL63KJ2_0),.doutb(w_n1042_0[1]),.din(n1042));
	jspl3 jspl3_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.doutc(w_n1059_0[2]),.din(n1059));
	jspl3 jspl3_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.doutc(w_n1067_0[2]),.din(n1067));
	jspl3 jspl3_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.doutc(w_n1069_0[2]),.din(n1069));
	jspl jspl_w_n1070_0(.douta(w_n1070_0[0]),.doutb(w_n1070_0[1]),.din(n1070));
	jspl jspl_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.din(n1073));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(n1078));
	jspl3 jspl3_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_dff_A_689w9I3n8_1),.doutc(w_dff_A_zIaVZtZh8_2),.din(n1084));
	jspl jspl_w_n1086_0(.douta(w_dff_A_5np9xzlW8_0),.doutb(w_n1086_0[1]),.din(w_dff_B_IrzrFxNw3_2));
	jspl jspl_w_n1090_0(.douta(w_n1090_0[0]),.doutb(w_n1090_0[1]),.din(n1090));
	jspl3 jspl3_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.doutc(w_n1092_0[2]),.din(n1092));
	jspl3 jspl3_w_n1094_0(.douta(w_dff_A_Rkv4QTmw4_0),.doutb(w_dff_A_dlGEQ5aM2_1),.doutc(w_n1094_0[2]),.din(w_dff_B_18wAMXjE5_3));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_dff_A_eNTiblVA7_1),.din(w_dff_B_dqPP4jvQ7_2));
	jspl jspl_w_n1106_0(.douta(w_n1106_0[0]),.doutb(w_dff_A_Da3PXiuw3_1),.din(n1106));
	jspl jspl_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_dff_A_ym1Eibhz7_1),.din(n1108));
	jspl jspl_w_n1113_0(.douta(w_n1113_0[0]),.doutb(w_n1113_0[1]),.din(n1113));
	jspl jspl_w_n1118_0(.douta(w_n1118_0[0]),.doutb(w_n1118_0[1]),.din(n1118));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(n1127));
	jspl jspl_w_n1137_0(.douta(w_n1137_0[0]),.doutb(w_n1137_0[1]),.din(n1137));
	jspl jspl_w_n1150_0(.douta(w_n1150_0[0]),.doutb(w_n1150_0[1]),.din(n1150));
	jspl jspl_w_n1172_0(.douta(w_n1172_0[0]),.doutb(w_n1172_0[1]),.din(n1172));
	jspl jspl_w_n1307_0(.douta(w_dff_A_IuxooMrp3_0),.doutb(w_n1307_0[1]),.din(w_dff_B_Y5woxDGt8_2));
	jspl jspl_w_n1308_0(.douta(w_n1308_0[0]),.doutb(w_dff_A_sEhCQmEg5_1),.din(n1308));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_dff_A_Uy6kw2GG4_1),.din(n1309));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_dff_A_oKs18H4K4_1),.din(w_dff_B_jm3SBMPv0_2));
	jspl3 jspl3_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.doutc(w_n1312_0[2]),.din(n1312));
	jspl jspl_w_n1312_1(.douta(w_n1312_1[0]),.doutb(w_n1312_1[1]),.din(w_n1312_0[0]));
	jspl jspl_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.din(n1316));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl3 jspl3_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.doutc(w_n1321_0[2]),.din(n1321));
	jspl jspl_w_n1321_1(.douta(w_n1321_1[0]),.doutb(w_n1321_1[1]),.din(w_n1321_0[0]));
	jspl jspl_w_n1323_0(.douta(w_n1323_0[0]),.doutb(w_n1323_0[1]),.din(w_dff_B_eapPgTTJ3_2));
	jspl jspl_w_n1333_0(.douta(w_n1333_0[0]),.doutb(w_n1333_0[1]),.din(n1333));
	jspl3 jspl3_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.doutc(w_n1337_0[2]),.din(n1337));
	jspl jspl_w_n1337_1(.douta(w_n1337_1[0]),.doutb(w_n1337_1[1]),.din(w_n1337_0[0]));
	jspl3 jspl3_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_dff_A_krkk7XAh3_1),.doutc(w_dff_A_jJI5G6gM5_2),.din(w_dff_B_tof5vAxJ8_3));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(n1343));
	jspl jspl_w_n1344_0(.douta(w_n1344_0[0]),.doutb(w_n1344_0[1]),.din(n1344));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_dff_A_OQiWABd12_1),.din(w_dff_B_H8oXmmA94_2));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_dff_A_xuCJl1nq8_1),.din(n1364));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(w_dff_B_rYSpOFRW4_2));
	jspl jspl_w_n1370_0(.douta(w_n1370_0[0]),.doutb(w_dff_A_Mo5ZWezW7_1),.din(w_dff_B_lJ5QNjnV4_2));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl jspl_w_n1387_0(.douta(w_dff_A_aqmJyNgr3_0),.doutb(w_n1387_0[1]),.din(n1387));
	jspl jspl_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_dff_A_LPFnN2Nq5_1),.din(n1388));
	jspl jspl_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.din(n1396));
	jspl jspl_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_dff_A_07VbPBFq4_1),.din(n1402));
	jspl jspl_w_n1408_0(.douta(w_n1408_0[0]),.doutb(w_dff_A_H227V6P77_1),.din(n1408));
	jspl jspl_w_n1419_0(.douta(w_n1419_0[0]),.doutb(w_dff_A_NRvr2xNV3_1),.din(w_dff_B_XkcTUA521_2));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_dff_A_mdctKRx36_1),.din(n1426));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(w_dff_B_34c1KuyF5_2));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.din(n1440));
	jspl3 jspl3_w_n1452_0(.douta(w_dff_A_TtsvZyKe2_0),.doutb(w_n1452_0[1]),.doutc(w_dff_A_7oZDXmlx4_2),.din(n1452));
	jspl jspl_w_n1458_0(.douta(w_n1458_0[0]),.doutb(w_n1458_0[1]),.din(n1458));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(n1486));
	jspl jspl_w_n1492_0(.douta(w_n1492_0[0]),.doutb(w_n1492_0[1]),.din(n1492));
	jspl jspl_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.din(n1506));
	jspl jspl_w_n1511_0(.douta(w_dff_A_GEC2RqG04_0),.doutb(w_n1511_0[1]),.din(w_dff_B_n59tdYKQ9_2));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.din(n1529));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(n1531));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(n1534));
	jspl jspl_w_n1536_0(.douta(w_dff_A_W85UgazU7_0),.doutb(w_n1536_0[1]),.din(n1536));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_dff_A_3BncMQJW6_1),.din(w_dff_B_24mtxUlb8_2));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl3 jspl3_w_n1562_0(.douta(w_dff_A_uzD2hOmg0_0),.doutb(w_dff_A_BGKrLFec7_1),.doutc(w_n1562_0[2]),.din(n1562));
	jspl jspl_w_n1587_0(.douta(w_n1587_0[0]),.doutb(w_n1587_0[1]),.din(n1587));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_dff_A_cU7m0Lw71_1),.din(w_dff_B_w8rOjI4n1_2));
	jspl jspl_w_n1605_0(.douta(w_dff_A_dOaRQNjy6_0),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1607_0(.douta(w_dff_A_6NPsbDMG0_0),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1620_0(.douta(w_dff_A_o1ibeUd56_0),.doutb(w_n1620_0[1]),.din(n1620));
	jspl jspl_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.din(n1624));
	jdff dff_A_n9g5SFgC7_0(.dout(w_G5_1[0]),.din(w_dff_A_n9g5SFgC7_0),.clk(gclk));
	jdff dff_A_7au7tv7s7_1(.dout(w_G5_0[1]),.din(w_dff_A_7au7tv7s7_1),.clk(gclk));
	jdff dff_A_QQzWuTYo3_2(.dout(w_G5_0[2]),.din(w_dff_A_QQzWuTYo3_2),.clk(gclk));
	jdff dff_B_eVb1uE7h3_2(.din(n347),.dout(w_dff_B_eVb1uE7h3_2),.clk(gclk));
	jdff dff_B_QW2NFVLj0_0(.din(n1072),.dout(w_dff_B_QW2NFVLj0_0),.clk(gclk));
	jdff dff_B_iv2qALu13_1(.din(n1085),.dout(w_dff_B_iv2qALu13_1),.clk(gclk));
	jdff dff_B_JL3Uxk8f4_1(.din(n753),.dout(w_dff_B_JL3Uxk8f4_1),.clk(gclk));
	jdff dff_B_nVkUxcQh2_1(.din(w_dff_B_JL3Uxk8f4_1),.dout(w_dff_B_nVkUxcQh2_1),.clk(gclk));
	jdff dff_B_dZFVaLSq9_1(.din(w_dff_B_nVkUxcQh2_1),.dout(w_dff_B_dZFVaLSq9_1),.clk(gclk));
	jdff dff_B_bxUYwUlW2_1(.din(w_dff_B_dZFVaLSq9_1),.dout(w_dff_B_bxUYwUlW2_1),.clk(gclk));
	jdff dff_B_rFvENq0u8_1(.din(w_dff_B_bxUYwUlW2_1),.dout(w_dff_B_rFvENq0u8_1),.clk(gclk));
	jdff dff_B_hlzU7xKp9_1(.din(w_dff_B_rFvENq0u8_1),.dout(w_dff_B_hlzU7xKp9_1),.clk(gclk));
	jdff dff_B_crLpbJdd3_1(.din(w_dff_B_hlzU7xKp9_1),.dout(w_dff_B_crLpbJdd3_1),.clk(gclk));
	jdff dff_B_7ugGyDHY8_1(.din(w_dff_B_crLpbJdd3_1),.dout(w_dff_B_7ugGyDHY8_1),.clk(gclk));
	jdff dff_B_aM0y4fTl0_1(.din(w_dff_B_7ugGyDHY8_1),.dout(w_dff_B_aM0y4fTl0_1),.clk(gclk));
	jdff dff_B_oKopyVDu0_1(.din(w_dff_B_aM0y4fTl0_1),.dout(w_dff_B_oKopyVDu0_1),.clk(gclk));
	jdff dff_B_VzZUjfJJ3_1(.din(w_dff_B_oKopyVDu0_1),.dout(w_dff_B_VzZUjfJJ3_1),.clk(gclk));
	jdff dff_B_LysNLlf65_1(.din(w_dff_B_VzZUjfJJ3_1),.dout(w_dff_B_LysNLlf65_1),.clk(gclk));
	jdff dff_B_ZSK9EZ2f6_1(.din(w_dff_B_LysNLlf65_1),.dout(w_dff_B_ZSK9EZ2f6_1),.clk(gclk));
	jdff dff_B_w359KRXJ1_1(.din(w_dff_B_ZSK9EZ2f6_1),.dout(w_dff_B_w359KRXJ1_1),.clk(gclk));
	jdff dff_B_QDqV3Viq0_1(.din(w_dff_B_w359KRXJ1_1),.dout(w_dff_B_QDqV3Viq0_1),.clk(gclk));
	jdff dff_B_izIiGylm2_1(.din(w_dff_B_QDqV3Viq0_1),.dout(w_dff_B_izIiGylm2_1),.clk(gclk));
	jdff dff_B_BQCItuAB9_1(.din(w_dff_B_izIiGylm2_1),.dout(w_dff_B_BQCItuAB9_1),.clk(gclk));
	jdff dff_B_8HFHMBLa2_0(.din(n1057),.dout(w_dff_B_8HFHMBLa2_0),.clk(gclk));
	jdff dff_B_Fh2BoDEf2_0(.din(w_dff_B_8HFHMBLa2_0),.dout(w_dff_B_Fh2BoDEf2_0),.clk(gclk));
	jdff dff_B_LVM4weCC0_0(.din(w_dff_B_Fh2BoDEf2_0),.dout(w_dff_B_LVM4weCC0_0),.clk(gclk));
	jdff dff_B_gW8CMy1h9_0(.din(w_dff_B_LVM4weCC0_0),.dout(w_dff_B_gW8CMy1h9_0),.clk(gclk));
	jdff dff_B_cxf56XXI2_0(.din(w_dff_B_gW8CMy1h9_0),.dout(w_dff_B_cxf56XXI2_0),.clk(gclk));
	jdff dff_B_EALYBs6j4_0(.din(w_dff_B_cxf56XXI2_0),.dout(w_dff_B_EALYBs6j4_0),.clk(gclk));
	jdff dff_B_RfPtmtFx6_0(.din(w_dff_B_EALYBs6j4_0),.dout(w_dff_B_RfPtmtFx6_0),.clk(gclk));
	jdff dff_B_HNUnMUZf5_0(.din(w_dff_B_RfPtmtFx6_0),.dout(w_dff_B_HNUnMUZf5_0),.clk(gclk));
	jdff dff_B_3yh1LDUD9_0(.din(w_dff_B_HNUnMUZf5_0),.dout(w_dff_B_3yh1LDUD9_0),.clk(gclk));
	jdff dff_B_rPsERgDg4_0(.din(w_dff_B_3yh1LDUD9_0),.dout(w_dff_B_rPsERgDg4_0),.clk(gclk));
	jdff dff_B_6aWEYUU27_0(.din(w_dff_B_rPsERgDg4_0),.dout(w_dff_B_6aWEYUU27_0),.clk(gclk));
	jdff dff_B_2gyqvWcx3_0(.din(w_dff_B_6aWEYUU27_0),.dout(w_dff_B_2gyqvWcx3_0),.clk(gclk));
	jdff dff_B_OJFaf4C45_0(.din(w_dff_B_2gyqvWcx3_0),.dout(w_dff_B_OJFaf4C45_0),.clk(gclk));
	jdff dff_B_agc9kbSX2_0(.din(w_dff_B_OJFaf4C45_0),.dout(w_dff_B_agc9kbSX2_0),.clk(gclk));
	jdff dff_B_QhklNHYJ1_0(.din(w_dff_B_agc9kbSX2_0),.dout(w_dff_B_QhklNHYJ1_0),.clk(gclk));
	jdff dff_B_4OlEFcVr6_0(.din(w_dff_B_QhklNHYJ1_0),.dout(w_dff_B_4OlEFcVr6_0),.clk(gclk));
	jdff dff_B_UWyCibH59_1(.din(n1048),.dout(w_dff_B_UWyCibH59_1),.clk(gclk));
	jdff dff_B_8JBo7MtE0_1(.din(w_dff_B_UWyCibH59_1),.dout(w_dff_B_8JBo7MtE0_1),.clk(gclk));
	jdff dff_B_2JDqAnWF6_1(.din(w_dff_B_8JBo7MtE0_1),.dout(w_dff_B_2JDqAnWF6_1),.clk(gclk));
	jdff dff_B_PNmrDce39_1(.din(w_dff_B_2JDqAnWF6_1),.dout(w_dff_B_PNmrDce39_1),.clk(gclk));
	jdff dff_B_aLZtl6TB0_1(.din(w_dff_B_PNmrDce39_1),.dout(w_dff_B_aLZtl6TB0_1),.clk(gclk));
	jdff dff_B_PVYmZCkK3_1(.din(n1049),.dout(w_dff_B_PVYmZCkK3_1),.clk(gclk));
	jdff dff_B_rhWpG1sa2_1(.din(w_dff_B_PVYmZCkK3_1),.dout(w_dff_B_rhWpG1sa2_1),.clk(gclk));
	jdff dff_B_LOovrd8T7_1(.din(w_dff_B_rhWpG1sa2_1),.dout(w_dff_B_LOovrd8T7_1),.clk(gclk));
	jdff dff_B_gMtGkkf78_1(.din(n1050),.dout(w_dff_B_gMtGkkf78_1),.clk(gclk));
	jdff dff_B_Xgr1Rhsw9_0(.din(n1044),.dout(w_dff_B_Xgr1Rhsw9_0),.clk(gclk));
	jdff dff_B_QB02PcLq1_0(.din(w_dff_B_Xgr1Rhsw9_0),.dout(w_dff_B_QB02PcLq1_0),.clk(gclk));
	jdff dff_B_oatz0fpB2_0(.din(w_dff_B_QB02PcLq1_0),.dout(w_dff_B_oatz0fpB2_0),.clk(gclk));
	jdff dff_B_XQf3rFE19_0(.din(w_dff_B_oatz0fpB2_0),.dout(w_dff_B_XQf3rFE19_0),.clk(gclk));
	jdff dff_B_vxvH3OFK4_0(.din(w_dff_B_XQf3rFE19_0),.dout(w_dff_B_vxvH3OFK4_0),.clk(gclk));
	jdff dff_B_GrPooNUC1_0(.din(w_dff_B_vxvH3OFK4_0),.dout(w_dff_B_GrPooNUC1_0),.clk(gclk));
	jdff dff_B_OfgiU85C0_0(.din(w_dff_B_GrPooNUC1_0),.dout(w_dff_B_OfgiU85C0_0),.clk(gclk));
	jdff dff_B_qPumAjg09_0(.din(w_dff_B_OfgiU85C0_0),.dout(w_dff_B_qPumAjg09_0),.clk(gclk));
	jdff dff_B_V0LyciSs5_0(.din(w_dff_B_qPumAjg09_0),.dout(w_dff_B_V0LyciSs5_0),.clk(gclk));
	jdff dff_B_Ka3Cw3Gj3_0(.din(w_dff_B_V0LyciSs5_0),.dout(w_dff_B_Ka3Cw3Gj3_0),.clk(gclk));
	jdff dff_B_BJYVUQtv6_0(.din(w_dff_B_Ka3Cw3Gj3_0),.dout(w_dff_B_BJYVUQtv6_0),.clk(gclk));
	jdff dff_B_GSjd4Lz08_0(.din(w_dff_B_BJYVUQtv6_0),.dout(w_dff_B_GSjd4Lz08_0),.clk(gclk));
	jdff dff_B_OQGKkDLd6_0(.din(w_dff_B_GSjd4Lz08_0),.dout(w_dff_B_OQGKkDLd6_0),.clk(gclk));
	jdff dff_B_uRaaM5jN4_0(.din(w_dff_B_OQGKkDLd6_0),.dout(w_dff_B_uRaaM5jN4_0),.clk(gclk));
	jdff dff_B_Q0RK8VJb7_0(.din(w_dff_B_uRaaM5jN4_0),.dout(w_dff_B_Q0RK8VJb7_0),.clk(gclk));
	jdff dff_B_RtWilZ243_0(.din(w_dff_B_Q0RK8VJb7_0),.dout(w_dff_B_RtWilZ243_0),.clk(gclk));
	jdff dff_B_g3X5V15h0_0(.din(w_dff_B_RtWilZ243_0),.dout(w_dff_B_g3X5V15h0_0),.clk(gclk));
	jdff dff_B_nKOYJWaS6_1(.din(n1040),.dout(w_dff_B_nKOYJWaS6_1),.clk(gclk));
	jdff dff_B_akVBs4rW7_1(.din(w_dff_B_nKOYJWaS6_1),.dout(w_dff_B_akVBs4rW7_1),.clk(gclk));
	jdff dff_A_etnL63KJ2_0(.dout(w_n1042_0[0]),.din(w_dff_A_etnL63KJ2_0),.clk(gclk));
	jdff dff_B_2PwnoF0C9_1(.din(n790),.dout(w_dff_B_2PwnoF0C9_1),.clk(gclk));
	jdff dff_B_BGoAAQot9_1(.din(w_dff_B_2PwnoF0C9_1),.dout(w_dff_B_BGoAAQot9_1),.clk(gclk));
	jdff dff_B_mjwidCI77_1(.din(w_dff_B_BGoAAQot9_1),.dout(w_dff_B_mjwidCI77_1),.clk(gclk));
	jdff dff_B_V9nMdID11_1(.din(w_dff_B_mjwidCI77_1),.dout(w_dff_B_V9nMdID11_1),.clk(gclk));
	jdff dff_B_tYdbC80R0_1(.din(w_dff_B_V9nMdID11_1),.dout(w_dff_B_tYdbC80R0_1),.clk(gclk));
	jdff dff_B_TH4u9rLa8_1(.din(w_dff_B_tYdbC80R0_1),.dout(w_dff_B_TH4u9rLa8_1),.clk(gclk));
	jdff dff_B_lAxSjQ1s9_1(.din(w_dff_B_TH4u9rLa8_1),.dout(w_dff_B_lAxSjQ1s9_1),.clk(gclk));
	jdff dff_B_5FUHYWFc4_1(.din(w_dff_B_lAxSjQ1s9_1),.dout(w_dff_B_5FUHYWFc4_1),.clk(gclk));
	jdff dff_B_En9U1VzK2_1(.din(w_dff_B_5FUHYWFc4_1),.dout(w_dff_B_En9U1VzK2_1),.clk(gclk));
	jdff dff_B_N2JrJOuG9_1(.din(w_dff_B_En9U1VzK2_1),.dout(w_dff_B_N2JrJOuG9_1),.clk(gclk));
	jdff dff_B_BlWityMK6_1(.din(w_dff_B_N2JrJOuG9_1),.dout(w_dff_B_BlWityMK6_1),.clk(gclk));
	jdff dff_B_jwk2BptA6_1(.din(w_dff_B_BlWityMK6_1),.dout(w_dff_B_jwk2BptA6_1),.clk(gclk));
	jdff dff_B_zPqGfzw23_1(.din(w_dff_B_jwk2BptA6_1),.dout(w_dff_B_zPqGfzw23_1),.clk(gclk));
	jdff dff_B_RbCkI6so9_1(.din(w_dff_B_zPqGfzw23_1),.dout(w_dff_B_RbCkI6so9_1),.clk(gclk));
	jdff dff_B_q2ed6MJC2_1(.din(w_dff_B_RbCkI6so9_1),.dout(w_dff_B_q2ed6MJC2_1),.clk(gclk));
	jdff dff_B_3dj0ESMk7_1(.din(n794),.dout(w_dff_B_3dj0ESMk7_1),.clk(gclk));
	jdff dff_B_Ly1Pwmrj8_1(.din(w_dff_B_3dj0ESMk7_1),.dout(w_dff_B_Ly1Pwmrj8_1),.clk(gclk));
	jdff dff_B_b8V7jSAR0_1(.din(w_dff_B_Ly1Pwmrj8_1),.dout(w_dff_B_b8V7jSAR0_1),.clk(gclk));
	jdff dff_B_ISYftX5M2_1(.din(w_dff_B_b8V7jSAR0_1),.dout(w_dff_B_ISYftX5M2_1),.clk(gclk));
	jdff dff_B_OJlOckdU6_1(.din(w_dff_B_ISYftX5M2_1),.dout(w_dff_B_OJlOckdU6_1),.clk(gclk));
	jdff dff_B_3UocEI9x1_1(.din(w_dff_B_OJlOckdU6_1),.dout(w_dff_B_3UocEI9x1_1),.clk(gclk));
	jdff dff_B_Zltogmk66_1(.din(w_dff_B_3UocEI9x1_1),.dout(w_dff_B_Zltogmk66_1),.clk(gclk));
	jdff dff_B_aGNbQitz5_1(.din(w_dff_B_Zltogmk66_1),.dout(w_dff_B_aGNbQitz5_1),.clk(gclk));
	jdff dff_B_tGTEbQFu9_1(.din(w_dff_B_aGNbQitz5_1),.dout(w_dff_B_tGTEbQFu9_1),.clk(gclk));
	jdff dff_B_t4PbNbjN9_1(.din(w_dff_B_tGTEbQFu9_1),.dout(w_dff_B_t4PbNbjN9_1),.clk(gclk));
	jdff dff_B_k4zYkSZL1_1(.din(w_dff_B_t4PbNbjN9_1),.dout(w_dff_B_k4zYkSZL1_1),.clk(gclk));
	jdff dff_B_pQAnTvFN7_1(.din(w_dff_B_k4zYkSZL1_1),.dout(w_dff_B_pQAnTvFN7_1),.clk(gclk));
	jdff dff_B_o6SHvsb31_1(.din(w_dff_B_pQAnTvFN7_1),.dout(w_dff_B_o6SHvsb31_1),.clk(gclk));
	jdff dff_B_17DmmvCM8_1(.din(w_dff_B_o6SHvsb31_1),.dout(w_dff_B_17DmmvCM8_1),.clk(gclk));
	jdff dff_B_gbMbJoQG1_1(.din(w_dff_B_17DmmvCM8_1),.dout(w_dff_B_gbMbJoQG1_1),.clk(gclk));
	jdff dff_B_CFcAvKLj6_0(.din(n1036),.dout(w_dff_B_CFcAvKLj6_0),.clk(gclk));
	jdff dff_B_rQbrq56t8_0(.din(w_dff_B_CFcAvKLj6_0),.dout(w_dff_B_rQbrq56t8_0),.clk(gclk));
	jdff dff_B_HmzUSUyA1_0(.din(w_dff_B_rQbrq56t8_0),.dout(w_dff_B_HmzUSUyA1_0),.clk(gclk));
	jdff dff_B_QXc6b5cQ2_0(.din(w_dff_B_HmzUSUyA1_0),.dout(w_dff_B_QXc6b5cQ2_0),.clk(gclk));
	jdff dff_B_X0FCGtHk4_0(.din(w_dff_B_QXc6b5cQ2_0),.dout(w_dff_B_X0FCGtHk4_0),.clk(gclk));
	jdff dff_B_PRKVWczS3_0(.din(w_dff_B_X0FCGtHk4_0),.dout(w_dff_B_PRKVWczS3_0),.clk(gclk));
	jdff dff_B_FDHQqxPH7_0(.din(w_dff_B_PRKVWczS3_0),.dout(w_dff_B_FDHQqxPH7_0),.clk(gclk));
	jdff dff_B_CdpEen625_0(.din(w_dff_B_FDHQqxPH7_0),.dout(w_dff_B_CdpEen625_0),.clk(gclk));
	jdff dff_B_h5sEIVQ94_0(.din(w_dff_B_CdpEen625_0),.dout(w_dff_B_h5sEIVQ94_0),.clk(gclk));
	jdff dff_B_hIYWDFIz8_0(.din(w_dff_B_h5sEIVQ94_0),.dout(w_dff_B_hIYWDFIz8_0),.clk(gclk));
	jdff dff_B_JQlIRtgm7_0(.din(w_dff_B_hIYWDFIz8_0),.dout(w_dff_B_JQlIRtgm7_0),.clk(gclk));
	jdff dff_B_dHo87xgk2_0(.din(w_dff_B_JQlIRtgm7_0),.dout(w_dff_B_dHo87xgk2_0),.clk(gclk));
	jdff dff_B_1QSc33RG0_0(.din(w_dff_B_dHo87xgk2_0),.dout(w_dff_B_1QSc33RG0_0),.clk(gclk));
	jdff dff_B_DWOeTdVH9_0(.din(w_dff_B_1QSc33RG0_0),.dout(w_dff_B_DWOeTdVH9_0),.clk(gclk));
	jdff dff_B_A988JWCx6_0(.din(w_dff_B_DWOeTdVH9_0),.dout(w_dff_B_A988JWCx6_0),.clk(gclk));
	jdff dff_B_Wrw5Hqd19_0(.din(w_dff_B_A988JWCx6_0),.dout(w_dff_B_Wrw5Hqd19_0),.clk(gclk));
	jdff dff_B_udaqWIxX2_1(.din(n842),.dout(w_dff_B_udaqWIxX2_1),.clk(gclk));
	jdff dff_B_UtZYf41y7_1(.din(w_dff_B_udaqWIxX2_1),.dout(w_dff_B_UtZYf41y7_1),.clk(gclk));
	jdff dff_B_SnWwyTbr1_1(.din(w_dff_B_UtZYf41y7_1),.dout(w_dff_B_SnWwyTbr1_1),.clk(gclk));
	jdff dff_B_DeBSnkJO1_1(.din(w_dff_B_SnWwyTbr1_1),.dout(w_dff_B_DeBSnkJO1_1),.clk(gclk));
	jdff dff_B_Ibq7IEn14_1(.din(w_dff_B_DeBSnkJO1_1),.dout(w_dff_B_Ibq7IEn14_1),.clk(gclk));
	jdff dff_B_V5letM908_1(.din(w_dff_B_Ibq7IEn14_1),.dout(w_dff_B_V5letM908_1),.clk(gclk));
	jdff dff_B_xZ4Xqwaj8_1(.din(w_dff_B_V5letM908_1),.dout(w_dff_B_xZ4Xqwaj8_1),.clk(gclk));
	jdff dff_B_DR71AT8P1_1(.din(w_dff_B_xZ4Xqwaj8_1),.dout(w_dff_B_DR71AT8P1_1),.clk(gclk));
	jdff dff_B_1HW4sbfE6_1(.din(w_dff_B_DR71AT8P1_1),.dout(w_dff_B_1HW4sbfE6_1),.clk(gclk));
	jdff dff_B_hqillBlo1_1(.din(w_dff_B_1HW4sbfE6_1),.dout(w_dff_B_hqillBlo1_1),.clk(gclk));
	jdff dff_B_jilyhg740_1(.din(w_dff_B_hqillBlo1_1),.dout(w_dff_B_jilyhg740_1),.clk(gclk));
	jdff dff_B_kU0byQFR8_1(.din(n843),.dout(w_dff_B_kU0byQFR8_1),.clk(gclk));
	jdff dff_B_Sx1uNu5a3_1(.din(w_dff_B_kU0byQFR8_1),.dout(w_dff_B_Sx1uNu5a3_1),.clk(gclk));
	jdff dff_B_dZGAQpab0_1(.din(w_dff_B_Sx1uNu5a3_1),.dout(w_dff_B_dZGAQpab0_1),.clk(gclk));
	jdff dff_B_xLdrZaIi8_1(.din(w_dff_B_dZGAQpab0_1),.dout(w_dff_B_xLdrZaIi8_1),.clk(gclk));
	jdff dff_B_JqCmj6pN7_1(.din(w_dff_B_xLdrZaIi8_1),.dout(w_dff_B_JqCmj6pN7_1),.clk(gclk));
	jdff dff_B_4Wuzp8db7_1(.din(w_dff_B_JqCmj6pN7_1),.dout(w_dff_B_4Wuzp8db7_1),.clk(gclk));
	jdff dff_B_wZtY4F0h6_1(.din(w_dff_B_4Wuzp8db7_1),.dout(w_dff_B_wZtY4F0h6_1),.clk(gclk));
	jdff dff_B_LWD6H3D95_1(.din(w_dff_B_wZtY4F0h6_1),.dout(w_dff_B_LWD6H3D95_1),.clk(gclk));
	jdff dff_B_FyyDFzm21_1(.din(w_dff_B_LWD6H3D95_1),.dout(w_dff_B_FyyDFzm21_1),.clk(gclk));
	jdff dff_B_hSbRrYUw8_1(.din(w_dff_B_FyyDFzm21_1),.dout(w_dff_B_hSbRrYUw8_1),.clk(gclk));
	jdff dff_B_UAu2N2p05_1(.din(w_dff_B_hSbRrYUw8_1),.dout(w_dff_B_UAu2N2p05_1),.clk(gclk));
	jdff dff_B_hDBXXTch2_1(.din(w_dff_B_UAu2N2p05_1),.dout(w_dff_B_hDBXXTch2_1),.clk(gclk));
	jdff dff_B_6ZZMi8gg9_1(.din(w_dff_B_hDBXXTch2_1),.dout(w_dff_B_6ZZMi8gg9_1),.clk(gclk));
	jdff dff_B_bp3JTHAO6_0(.din(n1031),.dout(w_dff_B_bp3JTHAO6_0),.clk(gclk));
	jdff dff_B_VOa6mjkz4_0(.din(w_dff_B_bp3JTHAO6_0),.dout(w_dff_B_VOa6mjkz4_0),.clk(gclk));
	jdff dff_B_obl5F4as6_0(.din(w_dff_B_VOa6mjkz4_0),.dout(w_dff_B_obl5F4as6_0),.clk(gclk));
	jdff dff_B_gcpaaMQq6_0(.din(w_dff_B_obl5F4as6_0),.dout(w_dff_B_gcpaaMQq6_0),.clk(gclk));
	jdff dff_B_C5z9MrMH0_0(.din(w_dff_B_gcpaaMQq6_0),.dout(w_dff_B_C5z9MrMH0_0),.clk(gclk));
	jdff dff_B_F25zxsnW1_0(.din(w_dff_B_C5z9MrMH0_0),.dout(w_dff_B_F25zxsnW1_0),.clk(gclk));
	jdff dff_B_xfLNtrgX0_0(.din(w_dff_B_F25zxsnW1_0),.dout(w_dff_B_xfLNtrgX0_0),.clk(gclk));
	jdff dff_B_hNdKFqWY8_0(.din(w_dff_B_xfLNtrgX0_0),.dout(w_dff_B_hNdKFqWY8_0),.clk(gclk));
	jdff dff_B_w78BfbYk0_0(.din(w_dff_B_hNdKFqWY8_0),.dout(w_dff_B_w78BfbYk0_0),.clk(gclk));
	jdff dff_B_IN28J2OI0_0(.din(w_dff_B_w78BfbYk0_0),.dout(w_dff_B_IN28J2OI0_0),.clk(gclk));
	jdff dff_B_g0IXKYU45_0(.din(w_dff_B_IN28J2OI0_0),.dout(w_dff_B_g0IXKYU45_0),.clk(gclk));
	jdff dff_B_4iCGeQns8_0(.din(w_dff_B_g0IXKYU45_0),.dout(w_dff_B_4iCGeQns8_0),.clk(gclk));
	jdff dff_B_Cz8YghvD9_0(.din(w_dff_B_4iCGeQns8_0),.dout(w_dff_B_Cz8YghvD9_0),.clk(gclk));
	jdff dff_B_cuMzDEww9_0(.din(w_dff_B_Cz8YghvD9_0),.dout(w_dff_B_cuMzDEww9_0),.clk(gclk));
	jdff dff_B_1fYsCXVZ7_0(.din(n841),.dout(w_dff_B_1fYsCXVZ7_0),.clk(gclk));
	jdff dff_B_RuudyVQP2_0(.din(w_dff_B_1fYsCXVZ7_0),.dout(w_dff_B_RuudyVQP2_0),.clk(gclk));
	jdff dff_B_ZkmYrJx73_1(.din(n837),.dout(w_dff_B_ZkmYrJx73_1),.clk(gclk));
	jdff dff_B_fNbtVY718_1(.din(n830),.dout(w_dff_B_fNbtVY718_1),.clk(gclk));
	jdff dff_B_PkOzYPwq0_0(.din(n828),.dout(w_dff_B_PkOzYPwq0_0),.clk(gclk));
	jdff dff_A_ZGaBYqMV5_1(.dout(w_n808_0[1]),.din(w_dff_A_ZGaBYqMV5_1),.clk(gclk));
	jdff dff_A_K0UyC9ij2_1(.dout(w_dff_A_ZGaBYqMV5_1),.din(w_dff_A_K0UyC9ij2_1),.clk(gclk));
	jdff dff_B_7UnKPXbe2_0(.din(n789),.dout(w_dff_B_7UnKPXbe2_0),.clk(gclk));
	jdff dff_B_AysCa2sL2_1(.din(n785),.dout(w_dff_B_AysCa2sL2_1),.clk(gclk));
	jdff dff_A_hL4QtHdo2_1(.dout(w_n773_0[1]),.din(w_dff_A_hL4QtHdo2_1),.clk(gclk));
	jdff dff_B_9uMlF7Ay0_2(.din(n766),.dout(w_dff_B_9uMlF7Ay0_2),.clk(gclk));
	jdff dff_B_tsEoyIJd7_1(.din(n730),.dout(w_dff_B_tsEoyIJd7_1),.clk(gclk));
	jdff dff_B_dobygOqp2_1(.din(w_dff_B_tsEoyIJd7_1),.dout(w_dff_B_dobygOqp2_1),.clk(gclk));
	jdff dff_B_TSRR2EAS2_1(.din(w_dff_B_dobygOqp2_1),.dout(w_dff_B_TSRR2EAS2_1),.clk(gclk));
	jdff dff_B_br1cFjSc2_1(.din(n731),.dout(w_dff_B_br1cFjSc2_1),.clk(gclk));
	jdff dff_B_m7N8lvTH8_1(.din(w_dff_B_br1cFjSc2_1),.dout(w_dff_B_m7N8lvTH8_1),.clk(gclk));
	jdff dff_B_XLCg4Vxz6_1(.din(n735),.dout(w_dff_B_XLCg4Vxz6_1),.clk(gclk));
	jdff dff_A_Jl51lhWb4_1(.dout(w_n724_0[1]),.din(w_dff_A_Jl51lhWb4_1),.clk(gclk));
	jdff dff_A_YFJq84cV2_1(.dout(w_dff_A_Jl51lhWb4_1),.din(w_dff_A_YFJq84cV2_1),.clk(gclk));
	jdff dff_A_UCuGhZcJ5_1(.dout(w_dff_A_YFJq84cV2_1),.din(w_dff_A_UCuGhZcJ5_1),.clk(gclk));
	jdff dff_A_lttAXzVh7_1(.dout(w_dff_A_UCuGhZcJ5_1),.din(w_dff_A_lttAXzVh7_1),.clk(gclk));
	jdff dff_B_wyZkRwqg1_3(.din(n718),.dout(w_dff_B_wyZkRwqg1_3),.clk(gclk));
	jdff dff_B_WFFcg9b19_3(.din(w_dff_B_wyZkRwqg1_3),.dout(w_dff_B_WFFcg9b19_3),.clk(gclk));
	jdff dff_B_GjJNepL59_3(.din(w_dff_B_WFFcg9b19_3),.dout(w_dff_B_GjJNepL59_3),.clk(gclk));
	jdff dff_B_3Y7CzIhi9_3(.din(w_dff_B_GjJNepL59_3),.dout(w_dff_B_3Y7CzIhi9_3),.clk(gclk));
	jdff dff_B_5FjumPSY2_3(.din(w_dff_B_3Y7CzIhi9_3),.dout(w_dff_B_5FjumPSY2_3),.clk(gclk));
	jdff dff_B_lnJSQtNq1_3(.din(w_dff_B_5FjumPSY2_3),.dout(w_dff_B_lnJSQtNq1_3),.clk(gclk));
	jdff dff_B_VYBVRL0s7_3(.din(w_dff_B_lnJSQtNq1_3),.dout(w_dff_B_VYBVRL0s7_3),.clk(gclk));
	jdff dff_B_cshPhwWY7_3(.din(w_dff_B_VYBVRL0s7_3),.dout(w_dff_B_cshPhwWY7_3),.clk(gclk));
	jdff dff_B_fAR5PAi63_3(.din(w_dff_B_cshPhwWY7_3),.dout(w_dff_B_fAR5PAi63_3),.clk(gclk));
	jdff dff_B_Tstrbp4H5_3(.din(w_dff_B_fAR5PAi63_3),.dout(w_dff_B_Tstrbp4H5_3),.clk(gclk));
	jdff dff_B_gwZrCtHh3_3(.din(w_dff_B_Tstrbp4H5_3),.dout(w_dff_B_gwZrCtHh3_3),.clk(gclk));
	jdff dff_B_ecySOCm87_3(.din(w_dff_B_gwZrCtHh3_3),.dout(w_dff_B_ecySOCm87_3),.clk(gclk));
	jdff dff_B_rYNRIiR07_3(.din(w_dff_B_ecySOCm87_3),.dout(w_dff_B_rYNRIiR07_3),.clk(gclk));
	jdff dff_B_KfHtvRn50_3(.din(w_dff_B_rYNRIiR07_3),.dout(w_dff_B_KfHtvRn50_3),.clk(gclk));
	jdff dff_B_AnFO0cLV7_3(.din(w_dff_B_KfHtvRn50_3),.dout(w_dff_B_AnFO0cLV7_3),.clk(gclk));
	jdff dff_B_qLiOIZ6E7_3(.din(w_dff_B_AnFO0cLV7_3),.dout(w_dff_B_qLiOIZ6E7_3),.clk(gclk));
	jdff dff_B_36q99d5L1_3(.din(w_dff_B_qLiOIZ6E7_3),.dout(w_dff_B_36q99d5L1_3),.clk(gclk));
	jdff dff_B_jN5ZtIgq2_3(.din(w_dff_B_36q99d5L1_3),.dout(w_dff_B_jN5ZtIgq2_3),.clk(gclk));
	jdff dff_B_Z4txTq0q7_3(.din(w_dff_B_jN5ZtIgq2_3),.dout(w_dff_B_Z4txTq0q7_3),.clk(gclk));
	jdff dff_B_CNLUHhKi7_3(.din(w_dff_B_Z4txTq0q7_3),.dout(w_dff_B_CNLUHhKi7_3),.clk(gclk));
	jdff dff_B_iTjKjlLP6_3(.din(w_dff_B_CNLUHhKi7_3),.dout(w_dff_B_iTjKjlLP6_3),.clk(gclk));
	jdff dff_B_NWmhIE741_3(.din(w_dff_B_iTjKjlLP6_3),.dout(w_dff_B_NWmhIE741_3),.clk(gclk));
	jdff dff_B_moekdsPF3_3(.din(w_dff_B_NWmhIE741_3),.dout(w_dff_B_moekdsPF3_3),.clk(gclk));
	jdff dff_B_47SaYpgW2_3(.din(w_dff_B_moekdsPF3_3),.dout(w_dff_B_47SaYpgW2_3),.clk(gclk));
	jdff dff_B_Xp7qq0Vb4_0(.din(n717),.dout(w_dff_B_Xp7qq0Vb4_0),.clk(gclk));
	jdff dff_B_XwvYcmZv1_1(.din(n1305),.dout(w_dff_B_XwvYcmZv1_1),.clk(gclk));
	jdff dff_B_1KBvtN5y0_1(.din(w_dff_B_XwvYcmZv1_1),.dout(w_dff_B_1KBvtN5y0_1),.clk(gclk));
	jdff dff_B_Z1MCnMhS5_1(.din(w_dff_B_1KBvtN5y0_1),.dout(w_dff_B_Z1MCnMhS5_1),.clk(gclk));
	jdff dff_B_8p0wyfGX5_1(.din(w_dff_B_Z1MCnMhS5_1),.dout(w_dff_B_8p0wyfGX5_1),.clk(gclk));
	jdff dff_B_BTItQeXr3_1(.din(w_dff_B_8p0wyfGX5_1),.dout(w_dff_B_BTItQeXr3_1),.clk(gclk));
	jdff dff_B_GcJ6Qs3N9_1(.din(w_dff_B_BTItQeXr3_1),.dout(w_dff_B_GcJ6Qs3N9_1),.clk(gclk));
	jdff dff_B_F2Ipz71k2_1(.din(w_dff_B_GcJ6Qs3N9_1),.dout(w_dff_B_F2Ipz71k2_1),.clk(gclk));
	jdff dff_B_Dnilearv7_1(.din(w_dff_B_F2Ipz71k2_1),.dout(w_dff_B_Dnilearv7_1),.clk(gclk));
	jdff dff_B_GanduZdd6_1(.din(w_dff_B_Dnilearv7_1),.dout(w_dff_B_GanduZdd6_1),.clk(gclk));
	jdff dff_B_OL0A4bTl4_1(.din(w_dff_B_GanduZdd6_1),.dout(w_dff_B_OL0A4bTl4_1),.clk(gclk));
	jdff dff_B_vEEIB46e3_1(.din(w_dff_B_OL0A4bTl4_1),.dout(w_dff_B_vEEIB46e3_1),.clk(gclk));
	jdff dff_B_lxQHE9iJ3_1(.din(w_dff_B_vEEIB46e3_1),.dout(w_dff_B_lxQHE9iJ3_1),.clk(gclk));
	jdff dff_B_YGEwG3Zv8_1(.din(w_dff_B_lxQHE9iJ3_1),.dout(w_dff_B_YGEwG3Zv8_1),.clk(gclk));
	jdff dff_B_oZNzsOXp5_1(.din(w_dff_B_YGEwG3Zv8_1),.dout(w_dff_B_oZNzsOXp5_1),.clk(gclk));
	jdff dff_B_PzZ9sjmD6_1(.din(w_dff_B_oZNzsOXp5_1),.dout(w_dff_B_PzZ9sjmD6_1),.clk(gclk));
	jdff dff_B_jDmQfozV5_1(.din(w_dff_B_PzZ9sjmD6_1),.dout(w_dff_B_jDmQfozV5_1),.clk(gclk));
	jdff dff_B_OQxyPvgY5_1(.din(w_dff_B_jDmQfozV5_1),.dout(w_dff_B_OQxyPvgY5_1),.clk(gclk));
	jdff dff_B_HZJ6luck2_1(.din(w_dff_B_OQxyPvgY5_1),.dout(w_dff_B_HZJ6luck2_1),.clk(gclk));
	jdff dff_B_iu6b9rUm6_1(.din(w_dff_B_HZJ6luck2_1),.dout(w_dff_B_iu6b9rUm6_1),.clk(gclk));
	jdff dff_B_kEcfKRZY5_1(.din(w_dff_B_iu6b9rUm6_1),.dout(w_dff_B_kEcfKRZY5_1),.clk(gclk));
	jdff dff_B_nnbLFFhQ7_1(.din(w_dff_B_kEcfKRZY5_1),.dout(w_dff_B_nnbLFFhQ7_1),.clk(gclk));
	jdff dff_B_ypHWpTQ32_1(.din(w_dff_B_nnbLFFhQ7_1),.dout(w_dff_B_ypHWpTQ32_1),.clk(gclk));
	jdff dff_B_LxQ2xTZx8_1(.din(n880),.dout(w_dff_B_LxQ2xTZx8_1),.clk(gclk));
	jdff dff_B_6sAumDgf3_1(.din(w_dff_B_LxQ2xTZx8_1),.dout(w_dff_B_6sAumDgf3_1),.clk(gclk));
	jdff dff_B_kfwgKews0_1(.din(w_dff_B_6sAumDgf3_1),.dout(w_dff_B_kfwgKews0_1),.clk(gclk));
	jdff dff_B_7Dn82H1x6_1(.din(w_dff_B_kfwgKews0_1),.dout(w_dff_B_7Dn82H1x6_1),.clk(gclk));
	jdff dff_B_jStP1M7t8_1(.din(w_dff_B_7Dn82H1x6_1),.dout(w_dff_B_jStP1M7t8_1),.clk(gclk));
	jdff dff_B_tOhu7D1u7_1(.din(w_dff_B_jStP1M7t8_1),.dout(w_dff_B_tOhu7D1u7_1),.clk(gclk));
	jdff dff_B_Mag9w8OI4_1(.din(w_dff_B_tOhu7D1u7_1),.dout(w_dff_B_Mag9w8OI4_1),.clk(gclk));
	jdff dff_B_ZdJKHoFX8_1(.din(w_dff_B_Mag9w8OI4_1),.dout(w_dff_B_ZdJKHoFX8_1),.clk(gclk));
	jdff dff_B_lx5nZqAc0_1(.din(w_dff_B_ZdJKHoFX8_1),.dout(w_dff_B_lx5nZqAc0_1),.clk(gclk));
	jdff dff_B_Oo0QY9Ih6_1(.din(n883),.dout(w_dff_B_Oo0QY9Ih6_1),.clk(gclk));
	jdff dff_B_QJBBCxc72_1(.din(w_dff_B_Oo0QY9Ih6_1),.dout(w_dff_B_QJBBCxc72_1),.clk(gclk));
	jdff dff_B_ttWn3OQ39_1(.din(w_dff_B_QJBBCxc72_1),.dout(w_dff_B_ttWn3OQ39_1),.clk(gclk));
	jdff dff_B_7TZ60Xwn9_1(.din(w_dff_B_ttWn3OQ39_1),.dout(w_dff_B_7TZ60Xwn9_1),.clk(gclk));
	jdff dff_B_ZgiK9XAF4_1(.din(w_dff_B_7TZ60Xwn9_1),.dout(w_dff_B_ZgiK9XAF4_1),.clk(gclk));
	jdff dff_B_Plyq66uC2_1(.din(w_dff_B_ZgiK9XAF4_1),.dout(w_dff_B_Plyq66uC2_1),.clk(gclk));
	jdff dff_B_uNYCFD427_1(.din(w_dff_B_Plyq66uC2_1),.dout(w_dff_B_uNYCFD427_1),.clk(gclk));
	jdff dff_B_P2UJUTcZ8_1(.din(w_dff_B_uNYCFD427_1),.dout(w_dff_B_P2UJUTcZ8_1),.clk(gclk));
	jdff dff_B_YTkSdiyG8_1(.din(w_dff_B_P2UJUTcZ8_1),.dout(w_dff_B_YTkSdiyG8_1),.clk(gclk));
	jdff dff_B_hoqQbiCM6_1(.din(w_dff_B_YTkSdiyG8_1),.dout(w_dff_B_hoqQbiCM6_1),.clk(gclk));
	jdff dff_B_8Nz34Ps88_0(.din(n1027),.dout(w_dff_B_8Nz34Ps88_0),.clk(gclk));
	jdff dff_B_RF3upjcN2_0(.din(w_dff_B_8Nz34Ps88_0),.dout(w_dff_B_RF3upjcN2_0),.clk(gclk));
	jdff dff_B_JB2wzUzL0_0(.din(w_dff_B_RF3upjcN2_0),.dout(w_dff_B_JB2wzUzL0_0),.clk(gclk));
	jdff dff_B_sQ5WW1bI7_0(.din(w_dff_B_JB2wzUzL0_0),.dout(w_dff_B_sQ5WW1bI7_0),.clk(gclk));
	jdff dff_B_Cwm1zvf69_0(.din(w_dff_B_sQ5WW1bI7_0),.dout(w_dff_B_Cwm1zvf69_0),.clk(gclk));
	jdff dff_B_kKSLLmd88_0(.din(w_dff_B_Cwm1zvf69_0),.dout(w_dff_B_kKSLLmd88_0),.clk(gclk));
	jdff dff_B_lh8VyK5u1_0(.din(w_dff_B_kKSLLmd88_0),.dout(w_dff_B_lh8VyK5u1_0),.clk(gclk));
	jdff dff_B_B2omcMka9_0(.din(w_dff_B_lh8VyK5u1_0),.dout(w_dff_B_B2omcMka9_0),.clk(gclk));
	jdff dff_B_23Ep1ycX0_0(.din(w_dff_B_B2omcMka9_0),.dout(w_dff_B_23Ep1ycX0_0),.clk(gclk));
	jdff dff_B_otYfyN7k6_0(.din(n1023),.dout(w_dff_B_otYfyN7k6_0),.clk(gclk));
	jdff dff_B_mFzj0fnV1_0(.din(w_dff_B_otYfyN7k6_0),.dout(w_dff_B_mFzj0fnV1_0),.clk(gclk));
	jdff dff_B_JQsr2JeB4_0(.din(w_dff_B_mFzj0fnV1_0),.dout(w_dff_B_JQsr2JeB4_0),.clk(gclk));
	jdff dff_B_QNMsegxi0_1(.din(n1017),.dout(w_dff_B_QNMsegxi0_1),.clk(gclk));
	jdff dff_B_PNhe6DRF0_1(.din(w_dff_B_QNMsegxi0_1),.dout(w_dff_B_PNhe6DRF0_1),.clk(gclk));
	jdff dff_B_AwPlcsak5_1(.din(w_dff_B_PNhe6DRF0_1),.dout(w_dff_B_AwPlcsak5_1),.clk(gclk));
	jdff dff_B_jorYkMEJ4_1(.din(w_dff_B_AwPlcsak5_1),.dout(w_dff_B_jorYkMEJ4_1),.clk(gclk));
	jdff dff_B_Hhr9qj9p0_0(.din(n1021),.dout(w_dff_B_Hhr9qj9p0_0),.clk(gclk));
	jdff dff_B_fKc0yDPw9_0(.din(w_dff_B_Hhr9qj9p0_0),.dout(w_dff_B_fKc0yDPw9_0),.clk(gclk));
	jdff dff_B_bLFA0pqD5_1(.din(n1013),.dout(w_dff_B_bLFA0pqD5_1),.clk(gclk));
	jdff dff_B_vETxS4Ly4_0(.din(n1011),.dout(w_dff_B_vETxS4Ly4_0),.clk(gclk));
	jdff dff_B_1vllwRkt2_0(.din(w_dff_B_vETxS4Ly4_0),.dout(w_dff_B_1vllwRkt2_0),.clk(gclk));
	jdff dff_B_4bXAa7Qs8_0(.din(w_dff_B_1vllwRkt2_0),.dout(w_dff_B_4bXAa7Qs8_0),.clk(gclk));
	jdff dff_B_Z2MGMkkr8_1(.din(n971),.dout(w_dff_B_Z2MGMkkr8_1),.clk(gclk));
	jdff dff_B_e3nt4qMF6_1(.din(w_dff_B_Z2MGMkkr8_1),.dout(w_dff_B_e3nt4qMF6_1),.clk(gclk));
	jdff dff_B_34isNXdR2_1(.din(w_dff_B_e3nt4qMF6_1),.dout(w_dff_B_34isNXdR2_1),.clk(gclk));
	jdff dff_B_3JTNGUfp6_1(.din(w_dff_B_34isNXdR2_1),.dout(w_dff_B_3JTNGUfp6_1),.clk(gclk));
	jdff dff_B_iSDLFJwX9_1(.din(w_dff_B_3JTNGUfp6_1),.dout(w_dff_B_iSDLFJwX9_1),.clk(gclk));
	jdff dff_B_ge5PWEz40_0(.din(n1009),.dout(w_dff_B_ge5PWEz40_0),.clk(gclk));
	jdff dff_B_ZDcraaM70_0(.din(w_dff_B_ge5PWEz40_0),.dout(w_dff_B_ZDcraaM70_0),.clk(gclk));
	jdff dff_B_HgrYxgY77_0(.din(w_dff_B_ZDcraaM70_0),.dout(w_dff_B_HgrYxgY77_0),.clk(gclk));
	jdff dff_A_wbodIdqm6_0(.dout(w_n1008_0[0]),.din(w_dff_A_wbodIdqm6_0),.clk(gclk));
	jdff dff_A_EAfLFRDE2_0(.dout(w_dff_A_wbodIdqm6_0),.din(w_dff_A_EAfLFRDE2_0),.clk(gclk));
	jdff dff_A_ZZF8lVze4_0(.dout(w_dff_A_EAfLFRDE2_0),.din(w_dff_A_ZZF8lVze4_0),.clk(gclk));
	jdff dff_A_A4sJ5E0u2_0(.dout(w_dff_A_ZZF8lVze4_0),.din(w_dff_A_A4sJ5E0u2_0),.clk(gclk));
	jdff dff_B_Ah2aUiDQ3_1(.din(n1002),.dout(w_dff_B_Ah2aUiDQ3_1),.clk(gclk));
	jdff dff_A_ezWMIB7q9_0(.dout(w_n1003_0[0]),.din(w_dff_A_ezWMIB7q9_0),.clk(gclk));
	jdff dff_A_N3BsIWX12_1(.dout(w_n1000_0[1]),.din(w_dff_A_N3BsIWX12_1),.clk(gclk));
	jdff dff_A_RhqxIhuS9_1(.dout(w_n985_0[1]),.din(w_dff_A_RhqxIhuS9_1),.clk(gclk));
	jdff dff_B_83cBPOSs0_2(.din(n985),.dout(w_dff_B_83cBPOSs0_2),.clk(gclk));
	jdff dff_B_sdDMOuXZ9_0(.din(n963),.dout(w_dff_B_sdDMOuXZ9_0),.clk(gclk));
	jdff dff_B_LEgRd1n37_0(.din(w_dff_B_sdDMOuXZ9_0),.dout(w_dff_B_LEgRd1n37_0),.clk(gclk));
	jdff dff_B_P0OTCDOI4_0(.din(w_dff_B_LEgRd1n37_0),.dout(w_dff_B_P0OTCDOI4_0),.clk(gclk));
	jdff dff_B_zkNYjj430_0(.din(w_dff_B_P0OTCDOI4_0),.dout(w_dff_B_zkNYjj430_0),.clk(gclk));
	jdff dff_B_tnYWgAfx1_0(.din(w_dff_B_zkNYjj430_0),.dout(w_dff_B_tnYWgAfx1_0),.clk(gclk));
	jdff dff_B_uZ9L45DT7_0(.din(w_dff_B_tnYWgAfx1_0),.dout(w_dff_B_uZ9L45DT7_0),.clk(gclk));
	jdff dff_B_orv1wjnb3_1(.din(n959),.dout(w_dff_B_orv1wjnb3_1),.clk(gclk));
	jdff dff_B_CNN3Tmiw0_0(.din(n957),.dout(w_dff_B_CNN3Tmiw0_0),.clk(gclk));
	jdff dff_B_4kWLMhoZ9_0(.din(w_dff_B_CNN3Tmiw0_0),.dout(w_dff_B_4kWLMhoZ9_0),.clk(gclk));
	jdff dff_B_xFBDYDCS7_0(.din(w_dff_B_4kWLMhoZ9_0),.dout(w_dff_B_xFBDYDCS7_0),.clk(gclk));
	jdff dff_B_JdUiZGCi0_0(.din(w_dff_B_xFBDYDCS7_0),.dout(w_dff_B_JdUiZGCi0_0),.clk(gclk));
	jdff dff_B_3bJApQEN4_0(.din(w_dff_B_JdUiZGCi0_0),.dout(w_dff_B_3bJApQEN4_0),.clk(gclk));
	jdff dff_B_estVN0us2_0(.din(n956),.dout(w_dff_B_estVN0us2_0),.clk(gclk));
	jdff dff_B_NehKFbxp0_0(.din(n941),.dout(w_dff_B_NehKFbxp0_0),.clk(gclk));
	jdff dff_B_9iZzCCub3_0(.din(w_dff_B_NehKFbxp0_0),.dout(w_dff_B_9iZzCCub3_0),.clk(gclk));
	jdff dff_B_CidzbUxa3_0(.din(w_dff_B_9iZzCCub3_0),.dout(w_dff_B_CidzbUxa3_0),.clk(gclk));
	jdff dff_B_MapM6INs9_0(.din(w_dff_B_CidzbUxa3_0),.dout(w_dff_B_MapM6INs9_0),.clk(gclk));
	jdff dff_B_BppfZCnu1_0(.din(w_dff_B_MapM6INs9_0),.dout(w_dff_B_BppfZCnu1_0),.clk(gclk));
	jdff dff_B_Nz54HwJD5_0(.din(n932),.dout(w_dff_B_Nz54HwJD5_0),.clk(gclk));
	jdff dff_B_ID7XDYqu7_0(.din(w_dff_B_Nz54HwJD5_0),.dout(w_dff_B_ID7XDYqu7_0),.clk(gclk));
	jdff dff_B_DwOjqOiE3_0(.din(w_dff_B_ID7XDYqu7_0),.dout(w_dff_B_DwOjqOiE3_0),.clk(gclk));
	jdff dff_B_k180PTCX8_0(.din(w_dff_B_DwOjqOiE3_0),.dout(w_dff_B_k180PTCX8_0),.clk(gclk));
	jdff dff_B_gxkXCOrE5_0(.din(n922),.dout(w_dff_B_gxkXCOrE5_0),.clk(gclk));
	jdff dff_B_zxf4LBxI1_0(.din(w_dff_B_gxkXCOrE5_0),.dout(w_dff_B_zxf4LBxI1_0),.clk(gclk));
	jdff dff_B_nggOTCOy9_0(.din(w_dff_B_zxf4LBxI1_0),.dout(w_dff_B_nggOTCOy9_0),.clk(gclk));
	jdff dff_B_bo2wYj5S3_1(.din(n889),.dout(w_dff_B_bo2wYj5S3_1),.clk(gclk));
	jdff dff_B_q6EnlDxl3_1(.din(w_dff_B_bo2wYj5S3_1),.dout(w_dff_B_q6EnlDxl3_1),.clk(gclk));
	jdff dff_B_ZauRDTiH8_1(.din(w_dff_B_q6EnlDxl3_1),.dout(w_dff_B_ZauRDTiH8_1),.clk(gclk));
	jdff dff_B_wRFYCBmU5_0(.din(n906),.dout(w_dff_B_wRFYCBmU5_0),.clk(gclk));
	jdff dff_B_1SRk8rnZ7_0(.din(w_dff_B_wRFYCBmU5_0),.dout(w_dff_B_1SRk8rnZ7_0),.clk(gclk));
	jdff dff_B_RnXkE3it4_0(.din(n897),.dout(w_dff_B_RnXkE3it4_0),.clk(gclk));
	jdff dff_B_BNFVeHPN2_0(.din(n896),.dout(w_dff_B_BNFVeHPN2_0),.clk(gclk));
	jdff dff_A_ZZDYvtpd2_0(.dout(w_G89_0[0]),.din(w_dff_A_ZZDYvtpd2_0),.clk(gclk));
	jdff dff_A_fwEvooYQ0_0(.dout(w_n895_0[0]),.din(w_dff_A_fwEvooYQ0_0),.clk(gclk));
	jdff dff_B_xCGAEQP75_0(.din(n879),.dout(w_dff_B_xCGAEQP75_0),.clk(gclk));
	jdff dff_B_R2ssDfRx2_1(.din(n875),.dout(w_dff_B_R2ssDfRx2_1),.clk(gclk));
	jdff dff_A_Ig6Jd2UU0_1(.dout(w_n863_0[1]),.din(w_dff_A_Ig6Jd2UU0_1),.clk(gclk));
	jdff dff_A_RuXzwzZo6_1(.dout(w_n856_0[1]),.din(w_dff_A_RuXzwzZo6_1),.clk(gclk));
	jdff dff_B_s5Hp0cC17_1(.din(n1347),.dout(w_dff_B_s5Hp0cC17_1),.clk(gclk));
	jdff dff_B_y6tAviAl7_1(.din(w_dff_B_s5Hp0cC17_1),.dout(w_dff_B_y6tAviAl7_1),.clk(gclk));
	jdff dff_B_eQadKVK99_1(.din(n1352),.dout(w_dff_B_eQadKVK99_1),.clk(gclk));
	jdff dff_B_QOmj15Uf4_1(.din(w_dff_B_eQadKVK99_1),.dout(w_dff_B_QOmj15Uf4_1),.clk(gclk));
	jdff dff_B_c06RZygx3_1(.din(w_dff_B_QOmj15Uf4_1),.dout(w_dff_B_c06RZygx3_1),.clk(gclk));
	jdff dff_B_sjOvuJzq8_1(.din(w_dff_B_c06RZygx3_1),.dout(w_dff_B_sjOvuJzq8_1),.clk(gclk));
	jdff dff_B_OaYYyJIi8_1(.din(w_dff_B_sjOvuJzq8_1),.dout(w_dff_B_OaYYyJIi8_1),.clk(gclk));
	jdff dff_B_YYagu3qC3_1(.din(w_dff_B_OaYYyJIi8_1),.dout(w_dff_B_YYagu3qC3_1),.clk(gclk));
	jdff dff_B_PNEekTyH5_1(.din(w_dff_B_YYagu3qC3_1),.dout(w_dff_B_PNEekTyH5_1),.clk(gclk));
	jdff dff_B_fUtICkG03_1(.din(w_dff_B_PNEekTyH5_1),.dout(w_dff_B_fUtICkG03_1),.clk(gclk));
	jdff dff_B_NQhm448A5_1(.din(w_dff_B_fUtICkG03_1),.dout(w_dff_B_NQhm448A5_1),.clk(gclk));
	jdff dff_B_26CUA39Z9_1(.din(w_dff_B_NQhm448A5_1),.dout(w_dff_B_26CUA39Z9_1),.clk(gclk));
	jdff dff_B_tnretszl7_1(.din(w_dff_B_26CUA39Z9_1),.dout(w_dff_B_tnretszl7_1),.clk(gclk));
	jdff dff_B_YnwHMZT42_1(.din(w_dff_B_tnretszl7_1),.dout(w_dff_B_YnwHMZT42_1),.clk(gclk));
	jdff dff_B_sfp0FJc35_1(.din(w_dff_B_YnwHMZT42_1),.dout(w_dff_B_sfp0FJc35_1),.clk(gclk));
	jdff dff_B_j8VXcBKN6_1(.din(w_dff_B_sfp0FJc35_1),.dout(w_dff_B_j8VXcBKN6_1),.clk(gclk));
	jdff dff_B_b2IvIusC6_1(.din(w_dff_B_j8VXcBKN6_1),.dout(w_dff_B_b2IvIusC6_1),.clk(gclk));
	jdff dff_B_PAWkJtJY9_1(.din(w_dff_B_b2IvIusC6_1),.dout(w_dff_B_PAWkJtJY9_1),.clk(gclk));
	jdff dff_B_v8NiatIJ7_1(.din(w_dff_B_PAWkJtJY9_1),.dout(w_dff_B_v8NiatIJ7_1),.clk(gclk));
	jdff dff_B_j67HeSxg9_1(.din(w_dff_B_v8NiatIJ7_1),.dout(w_dff_B_j67HeSxg9_1),.clk(gclk));
	jdff dff_B_rk62XQu75_1(.din(w_dff_B_j67HeSxg9_1),.dout(w_dff_B_rk62XQu75_1),.clk(gclk));
	jdff dff_B_Yyae2c6K8_1(.din(w_dff_B_rk62XQu75_1),.dout(w_dff_B_Yyae2c6K8_1),.clk(gclk));
	jdff dff_B_PzBMoEd49_1(.din(n1368),.dout(w_dff_B_PzBMoEd49_1),.clk(gclk));
	jdff dff_B_IPsu51sy8_1(.din(w_dff_B_PzBMoEd49_1),.dout(w_dff_B_IPsu51sy8_1),.clk(gclk));
	jdff dff_B_YCx18kfC2_1(.din(w_dff_B_IPsu51sy8_1),.dout(w_dff_B_YCx18kfC2_1),.clk(gclk));
	jdff dff_B_EBsTKoK00_1(.din(w_dff_B_YCx18kfC2_1),.dout(w_dff_B_EBsTKoK00_1),.clk(gclk));
	jdff dff_B_Biz1UDPJ3_1(.din(w_dff_B_EBsTKoK00_1),.dout(w_dff_B_Biz1UDPJ3_1),.clk(gclk));
	jdff dff_B_5rz7YNcP1_1(.din(w_dff_B_Biz1UDPJ3_1),.dout(w_dff_B_5rz7YNcP1_1),.clk(gclk));
	jdff dff_B_veDgjCRN8_1(.din(w_dff_B_5rz7YNcP1_1),.dout(w_dff_B_veDgjCRN8_1),.clk(gclk));
	jdff dff_B_LlzMOLUu9_1(.din(w_dff_B_veDgjCRN8_1),.dout(w_dff_B_LlzMOLUu9_1),.clk(gclk));
	jdff dff_B_jKGlioYE1_1(.din(w_dff_B_LlzMOLUu9_1),.dout(w_dff_B_jKGlioYE1_1),.clk(gclk));
	jdff dff_B_r3vDdZ8X0_1(.din(w_dff_B_jKGlioYE1_1),.dout(w_dff_B_r3vDdZ8X0_1),.clk(gclk));
	jdff dff_B_3AZH8EsJ1_1(.din(w_dff_B_r3vDdZ8X0_1),.dout(w_dff_B_3AZH8EsJ1_1),.clk(gclk));
	jdff dff_B_TIhj8ilP0_1(.din(w_dff_B_3AZH8EsJ1_1),.dout(w_dff_B_TIhj8ilP0_1),.clk(gclk));
	jdff dff_B_zAuZVIdH9_1(.din(w_dff_B_TIhj8ilP0_1),.dout(w_dff_B_zAuZVIdH9_1),.clk(gclk));
	jdff dff_B_mHSbwIWC5_1(.din(w_dff_B_zAuZVIdH9_1),.dout(w_dff_B_mHSbwIWC5_1),.clk(gclk));
	jdff dff_B_r0Yh98b39_1(.din(w_dff_B_mHSbwIWC5_1),.dout(w_dff_B_r0Yh98b39_1),.clk(gclk));
	jdff dff_B_lEZTA7sg4_1(.din(w_dff_B_r0Yh98b39_1),.dout(w_dff_B_lEZTA7sg4_1),.clk(gclk));
	jdff dff_B_Ib8tCxxr1_1(.din(w_dff_B_lEZTA7sg4_1),.dout(w_dff_B_Ib8tCxxr1_1),.clk(gclk));
	jdff dff_B_YW26d8oN5_1(.din(w_dff_B_Ib8tCxxr1_1),.dout(w_dff_B_YW26d8oN5_1),.clk(gclk));
	jdff dff_B_gtvralSJ4_1(.din(w_dff_B_YW26d8oN5_1),.dout(w_dff_B_gtvralSJ4_1),.clk(gclk));
	jdff dff_B_50cW6R5h5_1(.din(w_dff_B_gtvralSJ4_1),.dout(w_dff_B_50cW6R5h5_1),.clk(gclk));
	jdff dff_B_9vv4BaAl1_1(.din(w_dff_B_50cW6R5h5_1),.dout(w_dff_B_9vv4BaAl1_1),.clk(gclk));
	jdff dff_B_lT7YcpLB1_1(.din(w_dff_B_9vv4BaAl1_1),.dout(w_dff_B_lT7YcpLB1_1),.clk(gclk));
	jdff dff_B_RDORgMqD4_1(.din(w_dff_B_lT7YcpLB1_1),.dout(w_dff_B_RDORgMqD4_1),.clk(gclk));
	jdff dff_B_ALJ4lXBz2_1(.din(w_dff_B_RDORgMqD4_1),.dout(w_dff_B_ALJ4lXBz2_1),.clk(gclk));
	jdff dff_B_LX7CG5Qt4_1(.din(w_dff_B_ALJ4lXBz2_1),.dout(w_dff_B_LX7CG5Qt4_1),.clk(gclk));
	jdff dff_B_LZwkqAo59_1(.din(w_dff_B_LX7CG5Qt4_1),.dout(w_dff_B_LZwkqAo59_1),.clk(gclk));
	jdff dff_B_1DLfnPfQ1_1(.din(w_dff_B_LZwkqAo59_1),.dout(w_dff_B_1DLfnPfQ1_1),.clk(gclk));
	jdff dff_B_EcLzNYaP2_1(.din(w_dff_B_1DLfnPfQ1_1),.dout(w_dff_B_EcLzNYaP2_1),.clk(gclk));
	jdff dff_B_5DVjiJ859_1(.din(w_dff_B_EcLzNYaP2_1),.dout(w_dff_B_5DVjiJ859_1),.clk(gclk));
	jdff dff_B_97LKRyJs4_1(.din(w_dff_B_5DVjiJ859_1),.dout(w_dff_B_97LKRyJs4_1),.clk(gclk));
	jdff dff_B_hy9CQt7z0_1(.din(w_dff_B_97LKRyJs4_1),.dout(w_dff_B_hy9CQt7z0_1),.clk(gclk));
	jdff dff_B_JDntq90E5_1(.din(w_dff_B_hy9CQt7z0_1),.dout(w_dff_B_JDntq90E5_1),.clk(gclk));
	jdff dff_B_Vk81izGt4_1(.din(w_dff_B_JDntq90E5_1),.dout(w_dff_B_Vk81izGt4_1),.clk(gclk));
	jdff dff_B_ahLpG0yz2_2(.din(n1323),.dout(w_dff_B_ahLpG0yz2_2),.clk(gclk));
	jdff dff_B_A8Ubha8d9_2(.din(w_dff_B_ahLpG0yz2_2),.dout(w_dff_B_A8Ubha8d9_2),.clk(gclk));
	jdff dff_B_Pfp9khLw3_2(.din(w_dff_B_A8Ubha8d9_2),.dout(w_dff_B_Pfp9khLw3_2),.clk(gclk));
	jdff dff_B_JRXQ9fNn1_2(.din(w_dff_B_Pfp9khLw3_2),.dout(w_dff_B_JRXQ9fNn1_2),.clk(gclk));
	jdff dff_B_IIjiu3Bv2_2(.din(w_dff_B_JRXQ9fNn1_2),.dout(w_dff_B_IIjiu3Bv2_2),.clk(gclk));
	jdff dff_B_oLXc25eD2_2(.din(w_dff_B_IIjiu3Bv2_2),.dout(w_dff_B_oLXc25eD2_2),.clk(gclk));
	jdff dff_B_HiNlUkE01_2(.din(w_dff_B_oLXc25eD2_2),.dout(w_dff_B_HiNlUkE01_2),.clk(gclk));
	jdff dff_B_wsUnivT46_2(.din(w_dff_B_HiNlUkE01_2),.dout(w_dff_B_wsUnivT46_2),.clk(gclk));
	jdff dff_B_fsDYXqJj3_2(.din(w_dff_B_wsUnivT46_2),.dout(w_dff_B_fsDYXqJj3_2),.clk(gclk));
	jdff dff_B_cLBQPQYd8_2(.din(w_dff_B_fsDYXqJj3_2),.dout(w_dff_B_cLBQPQYd8_2),.clk(gclk));
	jdff dff_B_6NYEkpyw4_2(.din(w_dff_B_cLBQPQYd8_2),.dout(w_dff_B_6NYEkpyw4_2),.clk(gclk));
	jdff dff_B_Xzmf6IqD8_2(.din(w_dff_B_6NYEkpyw4_2),.dout(w_dff_B_Xzmf6IqD8_2),.clk(gclk));
	jdff dff_B_YNLKOk187_2(.din(w_dff_B_Xzmf6IqD8_2),.dout(w_dff_B_YNLKOk187_2),.clk(gclk));
	jdff dff_B_eQvRwRHh1_2(.din(w_dff_B_YNLKOk187_2),.dout(w_dff_B_eQvRwRHh1_2),.clk(gclk));
	jdff dff_B_LlkwaQ854_2(.din(w_dff_B_eQvRwRHh1_2),.dout(w_dff_B_LlkwaQ854_2),.clk(gclk));
	jdff dff_B_ofEo3QIb5_2(.din(w_dff_B_LlkwaQ854_2),.dout(w_dff_B_ofEo3QIb5_2),.clk(gclk));
	jdff dff_B_sOpolSFo4_2(.din(w_dff_B_ofEo3QIb5_2),.dout(w_dff_B_sOpolSFo4_2),.clk(gclk));
	jdff dff_B_sqbqov2b6_2(.din(w_dff_B_sOpolSFo4_2),.dout(w_dff_B_sqbqov2b6_2),.clk(gclk));
	jdff dff_B_zQFllWNM0_2(.din(w_dff_B_sqbqov2b6_2),.dout(w_dff_B_zQFllWNM0_2),.clk(gclk));
	jdff dff_B_cRySGfZj1_2(.din(w_dff_B_zQFllWNM0_2),.dout(w_dff_B_cRySGfZj1_2),.clk(gclk));
	jdff dff_B_x3F9zCXM5_2(.din(w_dff_B_cRySGfZj1_2),.dout(w_dff_B_x3F9zCXM5_2),.clk(gclk));
	jdff dff_B_Iwz6rXXn2_2(.din(w_dff_B_x3F9zCXM5_2),.dout(w_dff_B_Iwz6rXXn2_2),.clk(gclk));
	jdff dff_B_2wAmErmz5_2(.din(w_dff_B_Iwz6rXXn2_2),.dout(w_dff_B_2wAmErmz5_2),.clk(gclk));
	jdff dff_B_nPlACwd95_2(.din(w_dff_B_2wAmErmz5_2),.dout(w_dff_B_nPlACwd95_2),.clk(gclk));
	jdff dff_B_FfWgKOYy4_2(.din(w_dff_B_nPlACwd95_2),.dout(w_dff_B_FfWgKOYy4_2),.clk(gclk));
	jdff dff_B_1ul6ytrd7_2(.din(w_dff_B_FfWgKOYy4_2),.dout(w_dff_B_1ul6ytrd7_2),.clk(gclk));
	jdff dff_B_C7pro73t8_2(.din(w_dff_B_1ul6ytrd7_2),.dout(w_dff_B_C7pro73t8_2),.clk(gclk));
	jdff dff_B_xetpYuPs7_2(.din(w_dff_B_C7pro73t8_2),.dout(w_dff_B_xetpYuPs7_2),.clk(gclk));
	jdff dff_B_eapPgTTJ3_2(.din(w_dff_B_xetpYuPs7_2),.dout(w_dff_B_eapPgTTJ3_2),.clk(gclk));
	jdff dff_B_Nsi5X4a68_2(.din(n1369),.dout(w_dff_B_Nsi5X4a68_2),.clk(gclk));
	jdff dff_B_Bh2we42W7_2(.din(w_dff_B_Nsi5X4a68_2),.dout(w_dff_B_Bh2we42W7_2),.clk(gclk));
	jdff dff_B_ZQeZ26oA8_2(.din(w_dff_B_Bh2we42W7_2),.dout(w_dff_B_ZQeZ26oA8_2),.clk(gclk));
	jdff dff_B_XFy51k1n4_2(.din(w_dff_B_ZQeZ26oA8_2),.dout(w_dff_B_XFy51k1n4_2),.clk(gclk));
	jdff dff_B_0Ktn2SDL8_2(.din(w_dff_B_XFy51k1n4_2),.dout(w_dff_B_0Ktn2SDL8_2),.clk(gclk));
	jdff dff_B_V0recqrJ1_2(.din(w_dff_B_0Ktn2SDL8_2),.dout(w_dff_B_V0recqrJ1_2),.clk(gclk));
	jdff dff_B_3cYDWd4q5_2(.din(w_dff_B_V0recqrJ1_2),.dout(w_dff_B_3cYDWd4q5_2),.clk(gclk));
	jdff dff_B_cCwouaHD3_2(.din(w_dff_B_3cYDWd4q5_2),.dout(w_dff_B_cCwouaHD3_2),.clk(gclk));
	jdff dff_B_zOLsnwPo4_2(.din(w_dff_B_cCwouaHD3_2),.dout(w_dff_B_zOLsnwPo4_2),.clk(gclk));
	jdff dff_B_TW8d3bdG2_2(.din(w_dff_B_zOLsnwPo4_2),.dout(w_dff_B_TW8d3bdG2_2),.clk(gclk));
	jdff dff_B_ZAW1SaQB6_2(.din(w_dff_B_TW8d3bdG2_2),.dout(w_dff_B_ZAW1SaQB6_2),.clk(gclk));
	jdff dff_B_XL2DLYm64_2(.din(w_dff_B_ZAW1SaQB6_2),.dout(w_dff_B_XL2DLYm64_2),.clk(gclk));
	jdff dff_B_vOkVqBPd0_2(.din(w_dff_B_XL2DLYm64_2),.dout(w_dff_B_vOkVqBPd0_2),.clk(gclk));
	jdff dff_B_N2PZ3a1Q0_2(.din(w_dff_B_vOkVqBPd0_2),.dout(w_dff_B_N2PZ3a1Q0_2),.clk(gclk));
	jdff dff_B_SH94kbda1_2(.din(w_dff_B_N2PZ3a1Q0_2),.dout(w_dff_B_SH94kbda1_2),.clk(gclk));
	jdff dff_B_4a0rIBNL6_2(.din(w_dff_B_SH94kbda1_2),.dout(w_dff_B_4a0rIBNL6_2),.clk(gclk));
	jdff dff_B_Gor3mNL25_2(.din(w_dff_B_4a0rIBNL6_2),.dout(w_dff_B_Gor3mNL25_2),.clk(gclk));
	jdff dff_B_7vaA25NE1_2(.din(w_dff_B_Gor3mNL25_2),.dout(w_dff_B_7vaA25NE1_2),.clk(gclk));
	jdff dff_B_0YPyJ8Uc4_2(.din(w_dff_B_7vaA25NE1_2),.dout(w_dff_B_0YPyJ8Uc4_2),.clk(gclk));
	jdff dff_B_aXUwLWky9_2(.din(w_dff_B_0YPyJ8Uc4_2),.dout(w_dff_B_aXUwLWky9_2),.clk(gclk));
	jdff dff_B_2eIhZ2w12_2(.din(w_dff_B_aXUwLWky9_2),.dout(w_dff_B_2eIhZ2w12_2),.clk(gclk));
	jdff dff_B_C4w7ZstR7_2(.din(w_dff_B_2eIhZ2w12_2),.dout(w_dff_B_C4w7ZstR7_2),.clk(gclk));
	jdff dff_B_JjtbViYg2_2(.din(w_dff_B_C4w7ZstR7_2),.dout(w_dff_B_JjtbViYg2_2),.clk(gclk));
	jdff dff_B_vGWTtvqL1_2(.din(w_dff_B_JjtbViYg2_2),.dout(w_dff_B_vGWTtvqL1_2),.clk(gclk));
	jdff dff_B_7ZadreeO3_2(.din(w_dff_B_vGWTtvqL1_2),.dout(w_dff_B_7ZadreeO3_2),.clk(gclk));
	jdff dff_B_agoTf6pK2_2(.din(w_dff_B_7ZadreeO3_2),.dout(w_dff_B_agoTf6pK2_2),.clk(gclk));
	jdff dff_B_lCJ7p6YX6_2(.din(w_dff_B_agoTf6pK2_2),.dout(w_dff_B_lCJ7p6YX6_2),.clk(gclk));
	jdff dff_B_rqPDnjiC8_2(.din(w_dff_B_lCJ7p6YX6_2),.dout(w_dff_B_rqPDnjiC8_2),.clk(gclk));
	jdff dff_B_vuxAlKJW3_2(.din(w_dff_B_rqPDnjiC8_2),.dout(w_dff_B_vuxAlKJW3_2),.clk(gclk));
	jdff dff_B_gm6zH1U62_2(.din(w_dff_B_vuxAlKJW3_2),.dout(w_dff_B_gm6zH1U62_2),.clk(gclk));
	jdff dff_B_rYSpOFRW4_2(.din(w_dff_B_gm6zH1U62_2),.dout(w_dff_B_rYSpOFRW4_2),.clk(gclk));
	jdff dff_B_nnIPsxnx3_1(.din(n1377),.dout(w_dff_B_nnIPsxnx3_1),.clk(gclk));
	jdff dff_B_oJ3uk5Yu9_1(.din(w_dff_B_nnIPsxnx3_1),.dout(w_dff_B_oJ3uk5Yu9_1),.clk(gclk));
	jdff dff_B_5GBMW2tW7_1(.din(n1378),.dout(w_dff_B_5GBMW2tW7_1),.clk(gclk));
	jdff dff_B_SQrA1Ldx3_1(.din(w_dff_B_5GBMW2tW7_1),.dout(w_dff_B_SQrA1Ldx3_1),.clk(gclk));
	jdff dff_B_QfoNWJZa1_1(.din(w_dff_B_SQrA1Ldx3_1),.dout(w_dff_B_QfoNWJZa1_1),.clk(gclk));
	jdff dff_B_jZ1VNd3j9_1(.din(w_dff_B_QfoNWJZa1_1),.dout(w_dff_B_jZ1VNd3j9_1),.clk(gclk));
	jdff dff_B_zbpEuFZc3_1(.din(w_dff_B_jZ1VNd3j9_1),.dout(w_dff_B_zbpEuFZc3_1),.clk(gclk));
	jdff dff_B_6neiXGcZ2_1(.din(w_dff_B_zbpEuFZc3_1),.dout(w_dff_B_6neiXGcZ2_1),.clk(gclk));
	jdff dff_B_WsznJuhN4_1(.din(w_dff_B_6neiXGcZ2_1),.dout(w_dff_B_WsznJuhN4_1),.clk(gclk));
	jdff dff_B_D3ju29x52_1(.din(w_dff_B_WsznJuhN4_1),.dout(w_dff_B_D3ju29x52_1),.clk(gclk));
	jdff dff_B_NRiDnaVs1_0(.din(n1379),.dout(w_dff_B_NRiDnaVs1_0),.clk(gclk));
	jdff dff_B_xYAtRbtz9_0(.din(w_dff_B_NRiDnaVs1_0),.dout(w_dff_B_xYAtRbtz9_0),.clk(gclk));
	jdff dff_B_0P283q1G0_0(.din(w_dff_B_xYAtRbtz9_0),.dout(w_dff_B_0P283q1G0_0),.clk(gclk));
	jdff dff_B_DwLSuusb8_0(.din(w_dff_B_0P283q1G0_0),.dout(w_dff_B_DwLSuusb8_0),.clk(gclk));
	jdff dff_B_e5eFDp330_0(.din(w_dff_B_DwLSuusb8_0),.dout(w_dff_B_e5eFDp330_0),.clk(gclk));
	jdff dff_B_qNU6KT989_0(.din(w_dff_B_e5eFDp330_0),.dout(w_dff_B_qNU6KT989_0),.clk(gclk));
	jdff dff_B_hU40mBNJ5_0(.din(w_dff_B_qNU6KT989_0),.dout(w_dff_B_hU40mBNJ5_0),.clk(gclk));
	jdff dff_B_rfMi1FXX7_0(.din(n1177),.dout(w_dff_B_rfMi1FXX7_0),.clk(gclk));
	jdff dff_B_nYIWO4Zh3_0(.din(n1176),.dout(w_dff_B_nYIWO4Zh3_0),.clk(gclk));
	jdff dff_B_qZ37TkEr6_0(.din(n1174),.dout(w_dff_B_qZ37TkEr6_0),.clk(gclk));
	jdff dff_B_iO12gpId8_1(.din(n1171),.dout(w_dff_B_iO12gpId8_1),.clk(gclk));
	jdff dff_B_hETOkRjX2_0(.din(n1166),.dout(w_dff_B_hETOkRjX2_0),.clk(gclk));
	jdff dff_B_7CjXRu199_1(.din(n1153),.dout(w_dff_B_7CjXRu199_1),.clk(gclk));
	jdff dff_B_MEpDpiEk0_1(.din(w_dff_B_7CjXRu199_1),.dout(w_dff_B_MEpDpiEk0_1),.clk(gclk));
	jdff dff_B_jhQ9ZwHH8_1(.din(w_dff_B_MEpDpiEk0_1),.dout(w_dff_B_jhQ9ZwHH8_1),.clk(gclk));
	jdff dff_B_r4wVXBmI4_1(.din(w_dff_B_jhQ9ZwHH8_1),.dout(w_dff_B_r4wVXBmI4_1),.clk(gclk));
	jdff dff_B_ElLWtjbo3_1(.din(n1158),.dout(w_dff_B_ElLWtjbo3_1),.clk(gclk));
	jdff dff_B_yxh4zwZu0_0(.din(n1148),.dout(w_dff_B_yxh4zwZu0_0),.clk(gclk));
	jdff dff_B_DruvH7gb4_0(.din(w_dff_B_yxh4zwZu0_0),.dout(w_dff_B_DruvH7gb4_0),.clk(gclk));
	jdff dff_B_VqDCOUdL7_0(.din(n1146),.dout(w_dff_B_VqDCOUdL7_0),.clk(gclk));
	jdff dff_B_T8lypvRC0_0(.din(n1141),.dout(w_dff_B_T8lypvRC0_0),.clk(gclk));
	jdff dff_B_L7MDHylB8_1(.din(n1135),.dout(w_dff_B_L7MDHylB8_1),.clk(gclk));
	jdff dff_B_gX7dCrmQ4_0(.din(n1138),.dout(w_dff_B_gX7dCrmQ4_0),.clk(gclk));
	jdff dff_B_8KC414ka4_1(.din(n1136),.dout(w_dff_B_8KC414ka4_1),.clk(gclk));
	jdff dff_B_oSRhgFo17_1(.din(n1120),.dout(w_dff_B_oSRhgFo17_1),.clk(gclk));
	jdff dff_B_cxn5ESvY5_1(.din(n1121),.dout(w_dff_B_cxn5ESvY5_1),.clk(gclk));
	jdff dff_B_31ztlG9W9_1(.din(w_dff_B_cxn5ESvY5_1),.dout(w_dff_B_31ztlG9W9_1),.clk(gclk));
	jdff dff_B_LCvwGGe99_0(.din(n1131),.dout(w_dff_B_LCvwGGe99_0),.clk(gclk));
	jdff dff_B_jXbhs1Ts2_0(.din(w_dff_B_LCvwGGe99_0),.dout(w_dff_B_jXbhs1Ts2_0),.clk(gclk));
	jdff dff_B_gg1Pz5RC7_0(.din(n1119),.dout(w_dff_B_gg1Pz5RC7_0),.clk(gclk));
	jdff dff_B_dxTagTcf8_0(.din(n1303),.dout(w_dff_B_dxTagTcf8_0),.clk(gclk));
	jdff dff_B_8NSQiVkX4_1(.din(n1289),.dout(w_dff_B_8NSQiVkX4_1),.clk(gclk));
	jdff dff_B_pwJz712V9_1(.din(w_dff_B_8NSQiVkX4_1),.dout(w_dff_B_pwJz712V9_1),.clk(gclk));
	jdff dff_B_9OoVwt040_0(.din(n1301),.dout(w_dff_B_9OoVwt040_0),.clk(gclk));
	jdff dff_B_78xqVym44_0(.din(w_dff_B_9OoVwt040_0),.dout(w_dff_B_78xqVym44_0),.clk(gclk));
	jdff dff_B_VCPo7aj54_0(.din(n816),.dout(w_dff_B_VCPo7aj54_0),.clk(gclk));
	jdff dff_B_HI17SWLs1_0(.din(n809),.dout(w_dff_B_HI17SWLs1_0),.clk(gclk));
	jdff dff_B_xlnYYd9P9_0(.din(G174),.dout(w_dff_B_xlnYYd9P9_0),.clk(gclk));
	jdff dff_B_rilexsIN7_0(.din(G173),.dout(w_dff_B_rilexsIN7_0),.clk(gclk));
	jdff dff_B_ACptuE0V4_0(.din(G176),.dout(w_dff_B_ACptuE0V4_0),.clk(gclk));
	jdff dff_B_lVJBxmwj6_0(.din(G175),.dout(w_dff_B_lVJBxmwj6_0),.clk(gclk));
	jdff dff_B_8afCptDr6_0(.din(n802),.dout(w_dff_B_8afCptDr6_0),.clk(gclk));
	jdff dff_B_neYfZjv58_0(.din(G177),.dout(w_dff_B_neYfZjv58_0),.clk(gclk));
	jdff dff_A_dvAMxUoN8_0(.dout(w_n373_3[0]),.din(w_dff_A_dvAMxUoN8_0),.clk(gclk));
	jdff dff_B_XobirX4R6_0(.din(n823),.dout(w_dff_B_XobirX4R6_0),.clk(gclk));
	jdff dff_B_bqA7wn954_1(.din(n1270),.dout(w_dff_B_bqA7wn954_1),.clk(gclk));
	jdff dff_B_wiIQHOaU6_1(.din(w_dff_B_bqA7wn954_1),.dout(w_dff_B_wiIQHOaU6_1),.clk(gclk));
	jdff dff_B_bWgIHx2K6_1(.din(w_dff_B_wiIQHOaU6_1),.dout(w_dff_B_bWgIHx2K6_1),.clk(gclk));
	jdff dff_B_yr36TW4i6_1(.din(w_dff_B_bWgIHx2K6_1),.dout(w_dff_B_yr36TW4i6_1),.clk(gclk));
	jdff dff_B_9B07w0IG3_1(.din(n1275),.dout(w_dff_B_9B07w0IG3_1),.clk(gclk));
	jdff dff_A_kPtUaf2H8_0(.dout(w_n725_0[0]),.din(w_dff_A_kPtUaf2H8_0),.clk(gclk));
	jdff dff_A_PpFG70SJ1_0(.dout(w_dff_A_kPtUaf2H8_0),.din(w_dff_A_PpFG70SJ1_0),.clk(gclk));
	jdff dff_B_X6BYXpZV8_0(.din(G167),.dout(w_dff_B_X6BYXpZV8_0),.clk(gclk));
	jdff dff_A_kCiJr1094_0(.dout(w_n719_0[0]),.din(w_dff_A_kCiJr1094_0),.clk(gclk));
	jdff dff_A_2hx7wOQO9_0(.dout(w_dff_A_kCiJr1094_0),.din(w_dff_A_2hx7wOQO9_0),.clk(gclk));
	jdff dff_B_LdDA1UfB9_0(.din(G166),.dout(w_dff_B_LdDA1UfB9_0),.clk(gclk));
	jdff dff_B_q4LyJ9mr1_0(.din(G169),.dout(w_dff_B_q4LyJ9mr1_0),.clk(gclk));
	jdff dff_A_8Cb6vKBt0_2(.dout(w_n373_5[2]),.din(w_dff_A_8Cb6vKBt0_2),.clk(gclk));
	jdff dff_B_IC7aNWb99_0(.din(G168),.dout(w_dff_B_IC7aNWb99_0),.clk(gclk));
	jdff dff_B_4OUwLuKY1_1(.din(G170),.dout(w_dff_B_4OUwLuKY1_1),.clk(gclk));
	jdff dff_B_9v9MOOrH2_1(.din(n1257),.dout(w_dff_B_9v9MOOrH2_1),.clk(gclk));
	jdff dff_B_mVGGaIz23_0(.din(n850),.dout(w_dff_B_mVGGaIz23_0),.clk(gclk));
	jdff dff_A_9BgNPRCU5_1(.dout(w_n845_0[1]),.din(w_dff_A_9BgNPRCU5_1),.clk(gclk));
	jdff dff_B_mTocefGd9_0(.din(n844),.dout(w_dff_B_mTocefGd9_0),.clk(gclk));
	jdff dff_B_lnZwKp530_0(.din(n1259),.dout(w_dff_B_lnZwKp530_0),.clk(gclk));
	jdff dff_B_CwWHlkEl2_0(.din(G115),.dout(w_dff_B_CwWHlkEl2_0),.clk(gclk));
	jdff dff_B_fT6cpS2r5_0(.din(n965),.dout(w_dff_B_fT6cpS2r5_0),.clk(gclk));
	jdff dff_B_NfZNRfxe8_0(.din(n979),.dout(w_dff_B_NfZNRfxe8_0),.clk(gclk));
	jdff dff_B_fFR3xlQT2_0(.din(n972),.dout(w_dff_B_fFR3xlQT2_0),.clk(gclk));
	jdff dff_B_XXe0m7kV4_0(.din(n994),.dout(w_dff_B_XXe0m7kV4_0),.clk(gclk));
	jdff dff_B_cQLPEVoP8_0(.din(n986),.dout(w_dff_B_cQLPEVoP8_0),.clk(gclk));
	jdff dff_B_dnkm3fBP6_0(.din(n865),.dout(w_dff_B_dnkm3fBP6_0),.clk(gclk));
	jdff dff_B_fV89OfNc8_0(.din(n857),.dout(w_dff_B_fV89OfNc8_0),.clk(gclk));
	jdff dff_B_g6xz6nVJ6_0(.din(n1252),.dout(w_dff_B_g6xz6nVJ6_0),.clk(gclk));
	jdff dff_B_bxk0bZM88_0(.din(n899),.dout(w_dff_B_bxk0bZM88_0),.clk(gclk));
	jdff dff_B_MxQHdMvy2_0(.din(n890),.dout(w_dff_B_MxQHdMvy2_0),.clk(gclk));
	jdff dff_B_ZKWIEJTp2_0(.din(n915),.dout(w_dff_B_ZKWIEJTp2_0),.clk(gclk));
	jdff dff_B_9SokRwpu0_0(.din(n884),.dout(w_dff_B_9SokRwpu0_0),.clk(gclk));
	jdff dff_B_9bgLBXQJ9_0(.din(n1247),.dout(w_dff_B_9bgLBXQJ9_0),.clk(gclk));
	jdff dff_B_Jrk5eOK59_0(.din(n1245),.dout(w_dff_B_Jrk5eOK59_0),.clk(gclk));
	jdff dff_B_1rrGnPMp2_0(.din(G44),.dout(w_dff_B_1rrGnPMp2_0),.clk(gclk));
	jdff dff_B_5YrEWmCa8_0(.din(n1243),.dout(w_dff_B_5YrEWmCa8_0),.clk(gclk));
	jdff dff_B_4nTjbmam1_0(.din(n949),.dout(w_dff_B_4nTjbmam1_0),.clk(gclk));
	jdff dff_B_tC5oChiN6_0(.din(n943),.dout(w_dff_B_tC5oChiN6_0),.clk(gclk));
	jdff dff_B_q9i22s8O9_0(.din(n934),.dout(w_dff_B_q9i22s8O9_0),.clk(gclk));
	jdff dff_A_ZFgUO11s5_0(.dout(w_n926_0[0]),.din(w_dff_A_ZFgUO11s5_0),.clk(gclk));
	jdff dff_B_4s9IArk87_0(.din(n925),.dout(w_dff_B_4s9IArk87_0),.clk(gclk));
	jdff dff_A_ERBY7ag16_0(.dout(w_G414_0),.din(w_dff_A_ERBY7ag16_0),.clk(gclk));
	jdff dff_B_gRr2QMWX6_1(.din(n1228),.dout(w_dff_B_gRr2QMWX6_1),.clk(gclk));
	jdff dff_B_Y00uvtA76_1(.din(w_dff_B_gRr2QMWX6_1),.dout(w_dff_B_Y00uvtA76_1),.clk(gclk));
	jdff dff_B_VaOgOo7R7_0(.din(n1236),.dout(w_dff_B_VaOgOo7R7_0),.clk(gclk));
	jdff dff_B_FIx2mURg1_0(.din(n1234),.dout(w_dff_B_FIx2mURg1_0),.clk(gclk));
	jdff dff_B_U8wghQvY4_0(.din(n733),.dout(w_dff_B_U8wghQvY4_0),.clk(gclk));
	jdff dff_B_KVIsyAul7_0(.din(n746),.dout(w_dff_B_KVIsyAul7_0),.clk(gclk));
	jdff dff_B_oVCXBg7B5_0(.din(n740),.dout(w_dff_B_oVCXBg7B5_0),.clk(gclk));
	jdff dff_B_PknzMfj32_0(.din(n728),.dout(w_dff_B_PknzMfj32_0),.clk(gclk));
	jdff dff_B_suekqKZF4_0(.din(n722),.dout(w_dff_B_suekqKZF4_0),.clk(gclk));
	jdff dff_A_Cid0r0AO1_0(.dout(w_G2204_0[0]),.din(w_dff_A_Cid0r0AO1_0),.clk(gclk));
	jdff dff_A_RIAEFIVh8_2(.dout(w_G18_17[2]),.din(w_dff_A_RIAEFIVh8_2),.clk(gclk));
	jdff dff_A_1ikDeAhx6_2(.dout(w_dff_A_RIAEFIVh8_2),.din(w_dff_A_1ikDeAhx6_2),.clk(gclk));
	jdff dff_B_UT7DX8AU3_1(.din(n1212),.dout(w_dff_B_UT7DX8AU3_1),.clk(gclk));
	jdff dff_B_mmKU2qf88_1(.din(n1213),.dout(w_dff_B_mmKU2qf88_1),.clk(gclk));
	jdff dff_B_hIfhACI74_0(.din(n998),.dout(w_dff_B_hIfhACI74_0),.clk(gclk));
	jdff dff_A_HQPL7rNf1_0(.dout(w_G18_20[0]),.din(w_dff_A_HQPL7rNf1_0),.clk(gclk));
	jdff dff_B_lmDZK8E89_0(.din(n990),.dout(w_dff_B_lmDZK8E89_0),.clk(gclk));
	jdff dff_B_VAnidCBK9_1(.din(n1214),.dout(w_dff_B_VAnidCBK9_1),.clk(gclk));
	jdff dff_A_t7Tf8XrA0_1(.dout(w_n355_12[1]),.din(w_dff_A_t7Tf8XrA0_1),.clk(gclk));
	jdff dff_B_8rIQAGib9_0(.din(n969),.dout(w_dff_B_8rIQAGib9_0),.clk(gclk));
	jdff dff_B_UQfx4r7m6_0(.din(n982),.dout(w_dff_B_UQfx4r7m6_0),.clk(gclk));
	jdff dff_B_l3G4sekk1_0(.din(n976),.dout(w_dff_B_l3G4sekk1_0),.clk(gclk));
	jdff dff_B_i1Wnk4No1_0(.din(n869),.dout(w_dff_B_i1Wnk4No1_0),.clk(gclk));
	jdff dff_B_sQF7XcW14_0(.din(n861),.dout(w_dff_B_sQF7XcW14_0),.clk(gclk));
	jdff dff_B_VMN7qhTg7_0(.din(n853),.dout(w_dff_B_VMN7qhTg7_0),.clk(gclk));
	jdff dff_B_bTJoSfQD1_0(.din(n847),.dout(w_dff_B_bTJoSfQD1_0),.clk(gclk));
	jdff dff_B_LWRHO66N8_1(.din(n1195),.dout(w_dff_B_LWRHO66N8_1),.clk(gclk));
	jdff dff_A_6HllCUn99_0(.dout(w_n938_0[0]),.din(w_dff_A_6HllCUn99_0),.clk(gclk));
	jdff dff_B_DjGqyaxc6_0(.din(n937),.dout(w_dff_B_DjGqyaxc6_0),.clk(gclk));
	jdff dff_B_GVGkWjOU8_0(.din(n929),.dout(w_dff_B_GVGkWjOU8_0),.clk(gclk));
	jdff dff_A_rNjZUdEz4_0(.dout(w_n905_0[0]),.din(w_dff_A_rNjZUdEz4_0),.clk(gclk));
	jdff dff_B_erXJUqiE4_0(.din(n918),.dout(w_dff_B_erXJUqiE4_0),.clk(gclk));
	jdff dff_B_jCyB9P0P2_0(.din(n1198),.dout(w_dff_B_jCyB9P0P2_0),.clk(gclk));
	jdff dff_B_LTj0zE0V5_0(.din(n887),.dout(w_dff_B_LTj0zE0V5_0),.clk(gclk));
	jdff dff_B_6S7kVID85_0(.din(n902),.dout(w_dff_B_6S7kVID85_0),.clk(gclk));
	jdff dff_B_bEl0xenY5_0(.din(n893),.dout(w_dff_B_bEl0xenY5_0),.clk(gclk));
	jdff dff_B_K8YkDxMJ7_0(.din(n952),.dout(w_dff_B_K8YkDxMJ7_0),.clk(gclk));
	jdff dff_B_kX1qkxWd0_0(.din(n946),.dout(w_dff_B_kX1qkxWd0_0),.clk(gclk));
	jdff dff_B_ZDQVdoiT8_0(.din(n1190),.dout(w_dff_B_ZDQVdoiT8_0),.clk(gclk));
	jdff dff_B_6S4NPvSl2_0(.din(n763),.dout(w_dff_B_6S4NPvSl2_0),.clk(gclk));
	jdff dff_B_hZpeGKhD7_0(.din(n757),.dout(w_dff_B_hZpeGKhD7_0),.clk(gclk));
	jdff dff_B_LlYTllIS2_0(.din(n819),.dout(w_dff_B_LlYTllIS2_0),.clk(gclk));
	jdff dff_B_aJMHWVVK0_0(.din(n813),.dout(w_dff_B_aJMHWVVK0_0),.clk(gclk));
	jdff dff_B_IHKWq1ZS2_0(.din(n805),.dout(w_dff_B_IHKWq1ZS2_0),.clk(gclk));
	jdff dff_B_Q1fKgDge9_0(.din(n799),.dout(w_dff_B_Q1fKgDge9_0),.clk(gclk));
	jdff dff_B_eweljXyV3_0(.din(n1185),.dout(w_dff_B_eweljXyV3_0),.clk(gclk));
	jdff dff_B_motdm5k38_0(.din(n1183),.dout(w_dff_B_motdm5k38_0),.clk(gclk));
	jdff dff_B_NXZo4Vpb7_0(.din(n826),.dout(w_dff_B_NXZo4Vpb7_0),.clk(gclk));
	jdff dff_A_RwjGpHMx3_0(.dout(w_n780_0[0]),.din(w_dff_A_RwjGpHMx3_0),.clk(gclk));
	jdff dff_B_MevoUuZj5_0(.din(n779),.dout(w_dff_B_MevoUuZj5_0),.clk(gclk));
	jdff dff_B_rZiy9hkI1_0(.din(n771),.dout(w_dff_B_rZiy9hkI1_0),.clk(gclk));
	jdff dff_B_7harNJMF0_3(.din(n715),.dout(w_dff_B_7harNJMF0_3),.clk(gclk));
	jdff dff_B_8OB2MLuA2_3(.din(w_dff_B_7harNJMF0_3),.dout(w_dff_B_8OB2MLuA2_3),.clk(gclk));
	jdff dff_B_YnPVhjWc0_3(.din(w_dff_B_8OB2MLuA2_3),.dout(w_dff_B_YnPVhjWc0_3),.clk(gclk));
	jdff dff_B_eu4nILTo8_3(.din(w_dff_B_YnPVhjWc0_3),.dout(w_dff_B_eu4nILTo8_3),.clk(gclk));
	jdff dff_B_Vk2AVHSq9_3(.din(w_dff_B_eu4nILTo8_3),.dout(w_dff_B_Vk2AVHSq9_3),.clk(gclk));
	jdff dff_B_LJJj8OGw5_3(.din(w_dff_B_Vk2AVHSq9_3),.dout(w_dff_B_LJJj8OGw5_3),.clk(gclk));
	jdff dff_B_HIa3BgOe6_3(.din(w_dff_B_LJJj8OGw5_3),.dout(w_dff_B_HIa3BgOe6_3),.clk(gclk));
	jdff dff_B_JgJYS9W98_3(.din(w_dff_B_HIa3BgOe6_3),.dout(w_dff_B_JgJYS9W98_3),.clk(gclk));
	jdff dff_B_ESPycNKz5_3(.din(w_dff_B_JgJYS9W98_3),.dout(w_dff_B_ESPycNKz5_3),.clk(gclk));
	jdff dff_B_yWHsUTY29_3(.din(w_dff_B_ESPycNKz5_3),.dout(w_dff_B_yWHsUTY29_3),.clk(gclk));
	jdff dff_B_0gzNXEkO3_3(.din(w_dff_B_yWHsUTY29_3),.dout(w_dff_B_0gzNXEkO3_3),.clk(gclk));
	jdff dff_B_VvcJRpKe3_3(.din(w_dff_B_0gzNXEkO3_3),.dout(w_dff_B_VvcJRpKe3_3),.clk(gclk));
	jdff dff_B_Pf0PwEVi3_3(.din(w_dff_B_VvcJRpKe3_3),.dout(w_dff_B_Pf0PwEVi3_3),.clk(gclk));
	jdff dff_B_WPCQJIqE3_3(.din(w_dff_B_Pf0PwEVi3_3),.dout(w_dff_B_WPCQJIqE3_3),.clk(gclk));
	jdff dff_B_58YVGJTN1_3(.din(w_dff_B_WPCQJIqE3_3),.dout(w_dff_B_58YVGJTN1_3),.clk(gclk));
	jdff dff_B_MdRPCVhl7_3(.din(w_dff_B_58YVGJTN1_3),.dout(w_dff_B_MdRPCVhl7_3),.clk(gclk));
	jdff dff_B_Oew8zBW70_3(.din(w_dff_B_MdRPCVhl7_3),.dout(w_dff_B_Oew8zBW70_3),.clk(gclk));
	jdff dff_B_w0Mvhv1d9_3(.din(w_dff_B_Oew8zBW70_3),.dout(w_dff_B_w0Mvhv1d9_3),.clk(gclk));
	jdff dff_B_c8js4H3A1_3(.din(w_dff_B_w0Mvhv1d9_3),.dout(w_dff_B_c8js4H3A1_3),.clk(gclk));
	jdff dff_B_MBpvApYr2_3(.din(w_dff_B_c8js4H3A1_3),.dout(w_dff_B_MBpvApYr2_3),.clk(gclk));
	jdff dff_B_6rziHhf50_3(.din(w_dff_B_MBpvApYr2_3),.dout(w_dff_B_6rziHhf50_3),.clk(gclk));
	jdff dff_B_YeNXfyw63_3(.din(w_dff_B_6rziHhf50_3),.dout(w_dff_B_YeNXfyw63_3),.clk(gclk));
	jdff dff_B_yOSJnDMg0_3(.din(w_dff_B_YeNXfyw63_3),.dout(w_dff_B_yOSJnDMg0_3),.clk(gclk));
	jdff dff_B_U4aXV4h35_3(.din(w_dff_B_yOSJnDMg0_3),.dout(w_dff_B_U4aXV4h35_3),.clk(gclk));
	jdff dff_B_qEa75UDU2_3(.din(w_dff_B_U4aXV4h35_3),.dout(w_dff_B_qEa75UDU2_3),.clk(gclk));
	jdff dff_B_GVWJ8yq63_3(.din(w_dff_B_qEa75UDU2_3),.dout(w_dff_B_GVWJ8yq63_3),.clk(gclk));
	jdff dff_B_zSMpWHB00_3(.din(w_dff_B_GVWJ8yq63_3),.dout(w_dff_B_zSMpWHB00_3),.clk(gclk));
	jdff dff_B_v4tQL05P7_3(.din(w_dff_B_zSMpWHB00_3),.dout(w_dff_B_v4tQL05P7_3),.clk(gclk));
	jdff dff_B_Jl9eAITO4_3(.din(w_dff_B_v4tQL05P7_3),.dout(w_dff_B_Jl9eAITO4_3),.clk(gclk));
	jdff dff_B_E0sjvPnC4_3(.din(w_dff_B_Jl9eAITO4_3),.dout(w_dff_B_E0sjvPnC4_3),.clk(gclk));
	jdff dff_B_jz4mq0wf2_3(.din(w_dff_B_E0sjvPnC4_3),.dout(w_dff_B_jz4mq0wf2_3),.clk(gclk));
	jdff dff_B_htuktq9e4_3(.din(w_dff_B_jz4mq0wf2_3),.dout(w_dff_B_htuktq9e4_3),.clk(gclk));
	jdff dff_B_cHzQtCIR4_3(.din(w_dff_B_htuktq9e4_3),.dout(w_dff_B_cHzQtCIR4_3),.clk(gclk));
	jdff dff_B_jHOlOr462_3(.din(w_dff_B_cHzQtCIR4_3),.dout(w_dff_B_jHOlOr462_3),.clk(gclk));
	jdff dff_B_ZQL03hyj8_0(.din(n714),.dout(w_dff_B_ZQL03hyj8_0),.clk(gclk));
	jdff dff_B_twlXeJ7q4_1(.din(n1394),.dout(w_dff_B_twlXeJ7q4_1),.clk(gclk));
	jdff dff_B_XtVTCOOT6_1(.din(w_dff_B_twlXeJ7q4_1),.dout(w_dff_B_XtVTCOOT6_1),.clk(gclk));
	jdff dff_B_0ajKQru93_1(.din(w_dff_B_XtVTCOOT6_1),.dout(w_dff_B_0ajKQru93_1),.clk(gclk));
	jdff dff_B_mObBsoMl9_1(.din(w_dff_B_0ajKQru93_1),.dout(w_dff_B_mObBsoMl9_1),.clk(gclk));
	jdff dff_B_5NRuV43X0_1(.din(w_dff_B_mObBsoMl9_1),.dout(w_dff_B_5NRuV43X0_1),.clk(gclk));
	jdff dff_B_T6QZYIjE6_1(.din(w_dff_B_5NRuV43X0_1),.dout(w_dff_B_T6QZYIjE6_1),.clk(gclk));
	jdff dff_B_z2e1mNPa3_1(.din(w_dff_B_T6QZYIjE6_1),.dout(w_dff_B_z2e1mNPa3_1),.clk(gclk));
	jdff dff_B_JDGzKElI0_1(.din(w_dff_B_z2e1mNPa3_1),.dout(w_dff_B_JDGzKElI0_1),.clk(gclk));
	jdff dff_B_jZweMMIS4_1(.din(w_dff_B_JDGzKElI0_1),.dout(w_dff_B_jZweMMIS4_1),.clk(gclk));
	jdff dff_B_rmHqHeNi5_1(.din(w_dff_B_jZweMMIS4_1),.dout(w_dff_B_rmHqHeNi5_1),.clk(gclk));
	jdff dff_B_tkqYSXQp0_1(.din(w_dff_B_rmHqHeNi5_1),.dout(w_dff_B_tkqYSXQp0_1),.clk(gclk));
	jdff dff_B_JyJLMoj38_1(.din(w_dff_B_tkqYSXQp0_1),.dout(w_dff_B_JyJLMoj38_1),.clk(gclk));
	jdff dff_B_NOccPzQb0_1(.din(w_dff_B_JyJLMoj38_1),.dout(w_dff_B_NOccPzQb0_1),.clk(gclk));
	jdff dff_B_h6faLEoc9_1(.din(w_dff_B_NOccPzQb0_1),.dout(w_dff_B_h6faLEoc9_1),.clk(gclk));
	jdff dff_B_DpojqN0o5_1(.din(w_dff_B_h6faLEoc9_1),.dout(w_dff_B_DpojqN0o5_1),.clk(gclk));
	jdff dff_B_PERSpz908_1(.din(w_dff_B_DpojqN0o5_1),.dout(w_dff_B_PERSpz908_1),.clk(gclk));
	jdff dff_B_Lpz9wFYH3_1(.din(w_dff_B_PERSpz908_1),.dout(w_dff_B_Lpz9wFYH3_1),.clk(gclk));
	jdff dff_B_iBF0zSIX9_1(.din(w_dff_B_Lpz9wFYH3_1),.dout(w_dff_B_iBF0zSIX9_1),.clk(gclk));
	jdff dff_B_yEufKW7X7_1(.din(w_dff_B_iBF0zSIX9_1),.dout(w_dff_B_yEufKW7X7_1),.clk(gclk));
	jdff dff_B_fq0e9X9X7_1(.din(w_dff_B_yEufKW7X7_1),.dout(w_dff_B_fq0e9X9X7_1),.clk(gclk));
	jdff dff_B_FJr2wMqf2_1(.din(w_dff_B_fq0e9X9X7_1),.dout(w_dff_B_FJr2wMqf2_1),.clk(gclk));
	jdff dff_B_03xCJqGp8_1(.din(w_dff_B_FJr2wMqf2_1),.dout(w_dff_B_03xCJqGp8_1),.clk(gclk));
	jdff dff_B_sVVjQfj48_1(.din(w_dff_B_03xCJqGp8_1),.dout(w_dff_B_sVVjQfj48_1),.clk(gclk));
	jdff dff_B_BKunGsue7_1(.din(w_dff_B_sVVjQfj48_1),.dout(w_dff_B_BKunGsue7_1),.clk(gclk));
	jdff dff_B_8R73yoEh1_1(.din(w_dff_B_BKunGsue7_1),.dout(w_dff_B_8R73yoEh1_1),.clk(gclk));
	jdff dff_B_qjyl5HXG2_1(.din(w_dff_B_8R73yoEh1_1),.dout(w_dff_B_qjyl5HXG2_1),.clk(gclk));
	jdff dff_B_7EXr7k8h9_1(.din(w_dff_B_qjyl5HXG2_1),.dout(w_dff_B_7EXr7k8h9_1),.clk(gclk));
	jdff dff_B_0IJlOyoJ7_1(.din(w_dff_B_7EXr7k8h9_1),.dout(w_dff_B_0IJlOyoJ7_1),.clk(gclk));
	jdff dff_B_sUkka6jM2_1(.din(w_dff_B_0IJlOyoJ7_1),.dout(w_dff_B_sUkka6jM2_1),.clk(gclk));
	jdff dff_B_RSrplJz97_1(.din(w_dff_B_sUkka6jM2_1),.dout(w_dff_B_RSrplJz97_1),.clk(gclk));
	jdff dff_B_q3iB6P8T0_1(.din(w_dff_B_RSrplJz97_1),.dout(w_dff_B_q3iB6P8T0_1),.clk(gclk));
	jdff dff_B_gBVPGCjC2_1(.din(w_dff_B_q3iB6P8T0_1),.dout(w_dff_B_gBVPGCjC2_1),.clk(gclk));
	jdff dff_B_PO5zx7vC7_1(.din(w_dff_B_gBVPGCjC2_1),.dout(w_dff_B_PO5zx7vC7_1),.clk(gclk));
	jdff dff_B_5a4TbPj14_1(.din(w_dff_B_PO5zx7vC7_1),.dout(w_dff_B_5a4TbPj14_1),.clk(gclk));
	jdff dff_A_HBTyAc6I7_0(.dout(w_n713_0[0]),.din(w_dff_A_HBTyAc6I7_0),.clk(gclk));
	jdff dff_A_eMHmEffM2_0(.dout(w_dff_A_HBTyAc6I7_0),.din(w_dff_A_eMHmEffM2_0),.clk(gclk));
	jdff dff_A_5RNSaOsB4_0(.dout(w_dff_A_eMHmEffM2_0),.din(w_dff_A_5RNSaOsB4_0),.clk(gclk));
	jdff dff_A_7QrLGILF0_0(.dout(w_dff_A_5RNSaOsB4_0),.din(w_dff_A_7QrLGILF0_0),.clk(gclk));
	jdff dff_A_UqDAvpNu7_0(.dout(w_dff_A_7QrLGILF0_0),.din(w_dff_A_UqDAvpNu7_0),.clk(gclk));
	jdff dff_A_08piZveL4_0(.dout(w_dff_A_UqDAvpNu7_0),.din(w_dff_A_08piZveL4_0),.clk(gclk));
	jdff dff_A_GLjZCPGx4_0(.dout(w_dff_A_08piZveL4_0),.din(w_dff_A_GLjZCPGx4_0),.clk(gclk));
	jdff dff_A_dGsttuS78_0(.dout(w_dff_A_GLjZCPGx4_0),.din(w_dff_A_dGsttuS78_0),.clk(gclk));
	jdff dff_A_R3LwgNdi5_0(.dout(w_dff_A_dGsttuS78_0),.din(w_dff_A_R3LwgNdi5_0),.clk(gclk));
	jdff dff_A_z2ZIgc8r4_0(.dout(w_dff_A_R3LwgNdi5_0),.din(w_dff_A_z2ZIgc8r4_0),.clk(gclk));
	jdff dff_A_DYkcfs9h4_0(.dout(w_dff_A_z2ZIgc8r4_0),.din(w_dff_A_DYkcfs9h4_0),.clk(gclk));
	jdff dff_A_9ULzOk1L2_0(.dout(w_dff_A_DYkcfs9h4_0),.din(w_dff_A_9ULzOk1L2_0),.clk(gclk));
	jdff dff_A_a9dCG73h6_0(.dout(w_dff_A_9ULzOk1L2_0),.din(w_dff_A_a9dCG73h6_0),.clk(gclk));
	jdff dff_A_V3cVFiR18_0(.dout(w_dff_A_a9dCG73h6_0),.din(w_dff_A_V3cVFiR18_0),.clk(gclk));
	jdff dff_A_xwI6hixk2_0(.dout(w_dff_A_V3cVFiR18_0),.din(w_dff_A_xwI6hixk2_0),.clk(gclk));
	jdff dff_A_83rLeqmB9_0(.dout(w_dff_A_xwI6hixk2_0),.din(w_dff_A_83rLeqmB9_0),.clk(gclk));
	jdff dff_A_XXUM6CNb9_0(.dout(w_dff_A_83rLeqmB9_0),.din(w_dff_A_XXUM6CNb9_0),.clk(gclk));
	jdff dff_A_5zaQv1Fu1_0(.dout(w_dff_A_XXUM6CNb9_0),.din(w_dff_A_5zaQv1Fu1_0),.clk(gclk));
	jdff dff_A_migGWQ6K0_0(.dout(w_dff_A_5zaQv1Fu1_0),.din(w_dff_A_migGWQ6K0_0),.clk(gclk));
	jdff dff_A_lbXWVGxB4_0(.dout(w_dff_A_migGWQ6K0_0),.din(w_dff_A_lbXWVGxB4_0),.clk(gclk));
	jdff dff_A_uo4fPLGn1_0(.dout(w_dff_A_lbXWVGxB4_0),.din(w_dff_A_uo4fPLGn1_0),.clk(gclk));
	jdff dff_A_9v7X2MgY2_0(.dout(w_dff_A_uo4fPLGn1_0),.din(w_dff_A_9v7X2MgY2_0),.clk(gclk));
	jdff dff_A_zh8uifpR5_0(.dout(w_dff_A_9v7X2MgY2_0),.din(w_dff_A_zh8uifpR5_0),.clk(gclk));
	jdff dff_A_XDFsk4m49_0(.dout(w_dff_A_zh8uifpR5_0),.din(w_dff_A_XDFsk4m49_0),.clk(gclk));
	jdff dff_A_t8tGgAvN9_0(.dout(w_dff_A_XDFsk4m49_0),.din(w_dff_A_t8tGgAvN9_0),.clk(gclk));
	jdff dff_A_IvULAnd04_0(.dout(w_dff_A_t8tGgAvN9_0),.din(w_dff_A_IvULAnd04_0),.clk(gclk));
	jdff dff_A_5inUDP0s4_0(.dout(w_dff_A_IvULAnd04_0),.din(w_dff_A_5inUDP0s4_0),.clk(gclk));
	jdff dff_A_lDbIQf1M1_0(.dout(w_dff_A_5inUDP0s4_0),.din(w_dff_A_lDbIQf1M1_0),.clk(gclk));
	jdff dff_A_TLi6Ey8p3_0(.dout(w_dff_A_lDbIQf1M1_0),.din(w_dff_A_TLi6Ey8p3_0),.clk(gclk));
	jdff dff_A_C4WFfANq9_0(.dout(w_dff_A_TLi6Ey8p3_0),.din(w_dff_A_C4WFfANq9_0),.clk(gclk));
	jdff dff_A_UID0nzDd2_0(.dout(w_dff_A_C4WFfANq9_0),.din(w_dff_A_UID0nzDd2_0),.clk(gclk));
	jdff dff_A_brOidayp1_0(.dout(w_dff_A_UID0nzDd2_0),.din(w_dff_A_brOidayp1_0),.clk(gclk));
	jdff dff_A_1NxDNOAD3_0(.dout(w_dff_A_brOidayp1_0),.din(w_dff_A_1NxDNOAD3_0),.clk(gclk));
	jdff dff_A_wVLQgSOY1_0(.dout(w_G38_1[0]),.din(w_dff_A_wVLQgSOY1_0),.clk(gclk));
	jdff dff_A_ihZcVA6G5_1(.dout(w_G38_1[1]),.din(w_dff_A_ihZcVA6G5_1),.clk(gclk));
	jdff dff_A_BHKCSiIk4_0(.dout(w_n370_0[0]),.din(w_dff_A_BHKCSiIk4_0),.clk(gclk));
	jdff dff_A_2FSUKeD00_0(.dout(w_dff_A_BHKCSiIk4_0),.din(w_dff_A_2FSUKeD00_0),.clk(gclk));
	jdff dff_A_cEOHc9J08_1(.dout(w_n370_0[1]),.din(w_dff_A_cEOHc9J08_1),.clk(gclk));
	jdff dff_A_ehSBP0Yb4_1(.dout(w_dff_A_cEOHc9J08_1),.din(w_dff_A_ehSBP0Yb4_1),.clk(gclk));
	jdff dff_B_q0LQ1LIh0_3(.din(n370),.dout(w_dff_B_q0LQ1LIh0_3),.clk(gclk));
	jdff dff_B_E7JCIvke2_3(.din(w_dff_B_q0LQ1LIh0_3),.dout(w_dff_B_E7JCIvke2_3),.clk(gclk));
	jdff dff_B_wMLwoEFJ5_3(.din(w_dff_B_E7JCIvke2_3),.dout(w_dff_B_wMLwoEFJ5_3),.clk(gclk));
	jdff dff_B_FFS9hwVn0_3(.din(w_dff_B_wMLwoEFJ5_3),.dout(w_dff_B_FFS9hwVn0_3),.clk(gclk));
	jdff dff_B_Gj4y2JOc4_3(.din(w_dff_B_FFS9hwVn0_3),.dout(w_dff_B_Gj4y2JOc4_3),.clk(gclk));
	jdff dff_B_6PjPud009_3(.din(w_dff_B_Gj4y2JOc4_3),.dout(w_dff_B_6PjPud009_3),.clk(gclk));
	jdff dff_B_0Zy8qH1L9_3(.din(w_dff_B_6PjPud009_3),.dout(w_dff_B_0Zy8qH1L9_3),.clk(gclk));
	jdff dff_B_mHJbPJ679_3(.din(w_dff_B_0Zy8qH1L9_3),.dout(w_dff_B_mHJbPJ679_3),.clk(gclk));
	jdff dff_B_tBka5SwJ4_3(.din(w_dff_B_mHJbPJ679_3),.dout(w_dff_B_tBka5SwJ4_3),.clk(gclk));
	jdff dff_B_DdEpOIuM5_3(.din(w_dff_B_tBka5SwJ4_3),.dout(w_dff_B_DdEpOIuM5_3),.clk(gclk));
	jdff dff_B_RerjznoS2_3(.din(w_dff_B_DdEpOIuM5_3),.dout(w_dff_B_RerjznoS2_3),.clk(gclk));
	jdff dff_B_6iBaV3qT7_3(.din(w_dff_B_RerjznoS2_3),.dout(w_dff_B_6iBaV3qT7_3),.clk(gclk));
	jdff dff_B_y2IhB3Wx2_3(.din(w_dff_B_6iBaV3qT7_3),.dout(w_dff_B_y2IhB3Wx2_3),.clk(gclk));
	jdff dff_B_JFyCRsdG0_3(.din(w_dff_B_y2IhB3Wx2_3),.dout(w_dff_B_JFyCRsdG0_3),.clk(gclk));
	jdff dff_B_KuS2jGWu0_3(.din(w_dff_B_JFyCRsdG0_3),.dout(w_dff_B_KuS2jGWu0_3),.clk(gclk));
	jdff dff_B_xuvGn3c46_3(.din(w_dff_B_KuS2jGWu0_3),.dout(w_dff_B_xuvGn3c46_3),.clk(gclk));
	jdff dff_B_pc5SgHtI1_3(.din(w_dff_B_xuvGn3c46_3),.dout(w_dff_B_pc5SgHtI1_3),.clk(gclk));
	jdff dff_B_xUOIYxBN4_3(.din(w_dff_B_pc5SgHtI1_3),.dout(w_dff_B_xUOIYxBN4_3),.clk(gclk));
	jdff dff_B_DVHmYXEY2_3(.din(w_dff_B_xUOIYxBN4_3),.dout(w_dff_B_DVHmYXEY2_3),.clk(gclk));
	jdff dff_B_vEQQW6vH5_3(.din(w_dff_B_DVHmYXEY2_3),.dout(w_dff_B_vEQQW6vH5_3),.clk(gclk));
	jdff dff_B_0TcigI3U1_3(.din(w_dff_B_vEQQW6vH5_3),.dout(w_dff_B_0TcigI3U1_3),.clk(gclk));
	jdff dff_B_AlUWaXrM6_3(.din(w_dff_B_0TcigI3U1_3),.dout(w_dff_B_AlUWaXrM6_3),.clk(gclk));
	jdff dff_B_UJ55DKDV2_3(.din(w_dff_B_AlUWaXrM6_3),.dout(w_dff_B_UJ55DKDV2_3),.clk(gclk));
	jdff dff_B_adZOlTAc3_3(.din(w_dff_B_UJ55DKDV2_3),.dout(w_dff_B_adZOlTAc3_3),.clk(gclk));
	jdff dff_B_ZtTqyoaC8_3(.din(w_dff_B_adZOlTAc3_3),.dout(w_dff_B_ZtTqyoaC8_3),.clk(gclk));
	jdff dff_B_IIYzzFNh4_3(.din(w_dff_B_ZtTqyoaC8_3),.dout(w_dff_B_IIYzzFNh4_3),.clk(gclk));
	jdff dff_B_XKCGeKdu6_3(.din(w_dff_B_IIYzzFNh4_3),.dout(w_dff_B_XKCGeKdu6_3),.clk(gclk));
	jdff dff_B_xIIADPOF8_3(.din(w_dff_B_XKCGeKdu6_3),.dout(w_dff_B_xIIADPOF8_3),.clk(gclk));
	jdff dff_B_pKKk1fqI5_3(.din(w_dff_B_xIIADPOF8_3),.dout(w_dff_B_pKKk1fqI5_3),.clk(gclk));
	jdff dff_B_3UxzEWLV4_3(.din(w_dff_B_pKKk1fqI5_3),.dout(w_dff_B_3UxzEWLV4_3),.clk(gclk));
	jdff dff_B_otunNgPD3_3(.din(w_dff_B_3UxzEWLV4_3),.dout(w_dff_B_otunNgPD3_3),.clk(gclk));
	jdff dff_B_nxbVmBxn9_3(.din(w_dff_B_otunNgPD3_3),.dout(w_dff_B_nxbVmBxn9_3),.clk(gclk));
	jdff dff_B_gPMZX7B71_1(.din(n365),.dout(w_dff_B_gPMZX7B71_1),.clk(gclk));
	jdff dff_A_DpxLS1m19_2(.dout(w_n363_0[2]),.din(w_dff_A_DpxLS1m19_2),.clk(gclk));
	jdff dff_B_Uq11c23E3_3(.din(n363),.dout(w_dff_B_Uq11c23E3_3),.clk(gclk));
	jdff dff_B_QhcL4qzt4_3(.din(w_dff_B_Uq11c23E3_3),.dout(w_dff_B_QhcL4qzt4_3),.clk(gclk));
	jdff dff_B_1mfOWhPf0_3(.din(w_dff_B_QhcL4qzt4_3),.dout(w_dff_B_1mfOWhPf0_3),.clk(gclk));
	jdff dff_B_Rosh9z2W5_3(.din(w_dff_B_1mfOWhPf0_3),.dout(w_dff_B_Rosh9z2W5_3),.clk(gclk));
	jdff dff_B_LvtAVJsN0_3(.din(w_dff_B_Rosh9z2W5_3),.dout(w_dff_B_LvtAVJsN0_3),.clk(gclk));
	jdff dff_B_3RjnZiL48_3(.din(w_dff_B_LvtAVJsN0_3),.dout(w_dff_B_3RjnZiL48_3),.clk(gclk));
	jdff dff_B_rPE1qjcr5_3(.din(w_dff_B_3RjnZiL48_3),.dout(w_dff_B_rPE1qjcr5_3),.clk(gclk));
	jdff dff_B_a8fbWRL04_3(.din(w_dff_B_rPE1qjcr5_3),.dout(w_dff_B_a8fbWRL04_3),.clk(gclk));
	jdff dff_B_epQU5li38_3(.din(w_dff_B_a8fbWRL04_3),.dout(w_dff_B_epQU5li38_3),.clk(gclk));
	jdff dff_B_FeAzPCQL2_3(.din(w_dff_B_epQU5li38_3),.dout(w_dff_B_FeAzPCQL2_3),.clk(gclk));
	jdff dff_B_ZLhaZyTj5_3(.din(w_dff_B_FeAzPCQL2_3),.dout(w_dff_B_ZLhaZyTj5_3),.clk(gclk));
	jdff dff_B_UOMizGQl3_3(.din(w_dff_B_ZLhaZyTj5_3),.dout(w_dff_B_UOMizGQl3_3),.clk(gclk));
	jdff dff_B_Zf7VFlvj9_3(.din(w_dff_B_UOMizGQl3_3),.dout(w_dff_B_Zf7VFlvj9_3),.clk(gclk));
	jdff dff_B_PlUhUOXm0_3(.din(w_dff_B_Zf7VFlvj9_3),.dout(w_dff_B_PlUhUOXm0_3),.clk(gclk));
	jdff dff_B_7fTbE3Qs0_3(.din(w_dff_B_PlUhUOXm0_3),.dout(w_dff_B_7fTbE3Qs0_3),.clk(gclk));
	jdff dff_B_140LrTg14_3(.din(w_dff_B_7fTbE3Qs0_3),.dout(w_dff_B_140LrTg14_3),.clk(gclk));
	jdff dff_B_meu9KNNh7_3(.din(w_dff_B_140LrTg14_3),.dout(w_dff_B_meu9KNNh7_3),.clk(gclk));
	jdff dff_B_MlF8rQDI4_3(.din(w_dff_B_meu9KNNh7_3),.dout(w_dff_B_MlF8rQDI4_3),.clk(gclk));
	jdff dff_B_p1VP9w0V4_3(.din(w_dff_B_MlF8rQDI4_3),.dout(w_dff_B_p1VP9w0V4_3),.clk(gclk));
	jdff dff_B_laQWJH2k2_3(.din(w_dff_B_p1VP9w0V4_3),.dout(w_dff_B_laQWJH2k2_3),.clk(gclk));
	jdff dff_B_nh8BRbDh6_3(.din(w_dff_B_laQWJH2k2_3),.dout(w_dff_B_nh8BRbDh6_3),.clk(gclk));
	jdff dff_B_VLp3duVg2_3(.din(w_dff_B_nh8BRbDh6_3),.dout(w_dff_B_VLp3duVg2_3),.clk(gclk));
	jdff dff_B_jIgyEFNl8_3(.din(w_dff_B_VLp3duVg2_3),.dout(w_dff_B_jIgyEFNl8_3),.clk(gclk));
	jdff dff_B_LO4dsblm8_3(.din(w_dff_B_jIgyEFNl8_3),.dout(w_dff_B_LO4dsblm8_3),.clk(gclk));
	jdff dff_B_ofiOtxJx9_3(.din(w_dff_B_LO4dsblm8_3),.dout(w_dff_B_ofiOtxJx9_3),.clk(gclk));
	jdff dff_B_12GJp60D6_3(.din(w_dff_B_ofiOtxJx9_3),.dout(w_dff_B_12GJp60D6_3),.clk(gclk));
	jdff dff_B_tCs5qjH55_3(.din(w_dff_B_12GJp60D6_3),.dout(w_dff_B_tCs5qjH55_3),.clk(gclk));
	jdff dff_B_FlfoBxZO6_3(.din(w_dff_B_tCs5qjH55_3),.dout(w_dff_B_FlfoBxZO6_3),.clk(gclk));
	jdff dff_B_et4NPvVk8_3(.din(w_dff_B_FlfoBxZO6_3),.dout(w_dff_B_et4NPvVk8_3),.clk(gclk));
	jdff dff_B_85JHcCmn5_3(.din(w_dff_B_et4NPvVk8_3),.dout(w_dff_B_85JHcCmn5_3),.clk(gclk));
	jdff dff_B_8iLpfF7G6_3(.din(w_dff_B_85JHcCmn5_3),.dout(w_dff_B_8iLpfF7G6_3),.clk(gclk));
	jdff dff_B_93hIVo6c5_3(.din(w_dff_B_8iLpfF7G6_3),.dout(w_dff_B_93hIVo6c5_3),.clk(gclk));
	jdff dff_B_GwLzA4Vi2_3(.din(w_dff_B_93hIVo6c5_3),.dout(w_dff_B_GwLzA4Vi2_3),.clk(gclk));
	jdff dff_B_ICQHecuV9_3(.din(w_dff_B_GwLzA4Vi2_3),.dout(w_dff_B_ICQHecuV9_3),.clk(gclk));
	jdff dff_B_wWZk4Lds0_1(.din(n1409),.dout(w_dff_B_wWZk4Lds0_1),.clk(gclk));
	jdff dff_B_wJv8Z09L0_1(.din(w_dff_B_wWZk4Lds0_1),.dout(w_dff_B_wJv8Z09L0_1),.clk(gclk));
	jdff dff_B_KGtdqV2A3_1(.din(w_dff_B_wJv8Z09L0_1),.dout(w_dff_B_KGtdqV2A3_1),.clk(gclk));
	jdff dff_B_5tREL57K7_1(.din(w_dff_B_KGtdqV2A3_1),.dout(w_dff_B_5tREL57K7_1),.clk(gclk));
	jdff dff_B_RF5t2aVj9_1(.din(w_dff_B_5tREL57K7_1),.dout(w_dff_B_RF5t2aVj9_1),.clk(gclk));
	jdff dff_B_WcJaMcar2_1(.din(w_dff_B_RF5t2aVj9_1),.dout(w_dff_B_WcJaMcar2_1),.clk(gclk));
	jdff dff_B_LQia12gc9_1(.din(w_dff_B_WcJaMcar2_1),.dout(w_dff_B_LQia12gc9_1),.clk(gclk));
	jdff dff_B_feOQWGXI5_0(.din(n1423),.dout(w_dff_B_feOQWGXI5_0),.clk(gclk));
	jdff dff_B_9nxREcP01_0(.din(w_dff_B_feOQWGXI5_0),.dout(w_dff_B_9nxREcP01_0),.clk(gclk));
	jdff dff_B_GBOVEWZc9_0(.din(w_dff_B_9nxREcP01_0),.dout(w_dff_B_GBOVEWZc9_0),.clk(gclk));
	jdff dff_B_yZhpUOE74_0(.din(w_dff_B_GBOVEWZc9_0),.dout(w_dff_B_yZhpUOE74_0),.clk(gclk));
	jdff dff_B_q5H8wVDo8_0(.din(w_dff_B_yZhpUOE74_0),.dout(w_dff_B_q5H8wVDo8_0),.clk(gclk));
	jdff dff_B_4SapPi330_0(.din(w_dff_B_q5H8wVDo8_0),.dout(w_dff_B_4SapPi330_0),.clk(gclk));
	jdff dff_B_qSPEZmw36_0(.din(w_dff_B_4SapPi330_0),.dout(w_dff_B_qSPEZmw36_0),.clk(gclk));
	jdff dff_B_PKJyVjaC7_0(.din(w_dff_B_qSPEZmw36_0),.dout(w_dff_B_PKJyVjaC7_0),.clk(gclk));
	jdff dff_B_1pLUySZd3_0(.din(w_dff_B_PKJyVjaC7_0),.dout(w_dff_B_1pLUySZd3_0),.clk(gclk));
	jdff dff_B_qZd0qqtg9_0(.din(w_dff_B_1pLUySZd3_0),.dout(w_dff_B_qZd0qqtg9_0),.clk(gclk));
	jdff dff_B_zb3Fl8IE9_0(.din(w_dff_B_qZd0qqtg9_0),.dout(w_dff_B_zb3Fl8IE9_0),.clk(gclk));
	jdff dff_B_nBniW0zQ0_0(.din(w_dff_B_zb3Fl8IE9_0),.dout(w_dff_B_nBniW0zQ0_0),.clk(gclk));
	jdff dff_B_oQY7Vf4N0_0(.din(w_dff_B_nBniW0zQ0_0),.dout(w_dff_B_oQY7Vf4N0_0),.clk(gclk));
	jdff dff_B_hvJq30dk8_0(.din(w_dff_B_oQY7Vf4N0_0),.dout(w_dff_B_hvJq30dk8_0),.clk(gclk));
	jdff dff_B_NDmSaG2h9_0(.din(w_dff_B_hvJq30dk8_0),.dout(w_dff_B_NDmSaG2h9_0),.clk(gclk));
	jdff dff_B_9Ijh9dG00_0(.din(w_dff_B_NDmSaG2h9_0),.dout(w_dff_B_9Ijh9dG00_0),.clk(gclk));
	jdff dff_B_TK2VkFiS0_0(.din(n1478),.dout(w_dff_B_TK2VkFiS0_0),.clk(gclk));
	jdff dff_B_12HAZl668_0(.din(w_dff_B_TK2VkFiS0_0),.dout(w_dff_B_12HAZl668_0),.clk(gclk));
	jdff dff_B_oSPfDfeT1_0(.din(n1477),.dout(w_dff_B_oSPfDfeT1_0),.clk(gclk));
	jdff dff_B_3A12Cw1k7_0(.din(w_dff_B_oSPfDfeT1_0),.dout(w_dff_B_3A12Cw1k7_0),.clk(gclk));
	jdff dff_B_1NZYUUDW3_0(.din(w_dff_B_3A12Cw1k7_0),.dout(w_dff_B_1NZYUUDW3_0),.clk(gclk));
	jdff dff_B_DxnJ7JMd7_0(.din(w_dff_B_1NZYUUDW3_0),.dout(w_dff_B_DxnJ7JMd7_0),.clk(gclk));
	jdff dff_B_ruU84gPK4_0(.din(w_dff_B_DxnJ7JMd7_0),.dout(w_dff_B_ruU84gPK4_0),.clk(gclk));
	jdff dff_B_D5dEVWu88_0(.din(w_dff_B_ruU84gPK4_0),.dout(w_dff_B_D5dEVWu88_0),.clk(gclk));
	jdff dff_B_8vozDF7V2_0(.din(w_dff_B_D5dEVWu88_0),.dout(w_dff_B_8vozDF7V2_0),.clk(gclk));
	jdff dff_B_5qcoIMpU2_0(.din(w_dff_B_8vozDF7V2_0),.dout(w_dff_B_5qcoIMpU2_0),.clk(gclk));
	jdff dff_B_Ca4LTnJZ4_0(.din(w_dff_B_5qcoIMpU2_0),.dout(w_dff_B_Ca4LTnJZ4_0),.clk(gclk));
	jdff dff_B_gIhRgRjM1_0(.din(w_dff_B_Ca4LTnJZ4_0),.dout(w_dff_B_gIhRgRjM1_0),.clk(gclk));
	jdff dff_B_Zt8ILZVx8_0(.din(w_dff_B_gIhRgRjM1_0),.dout(w_dff_B_Zt8ILZVx8_0),.clk(gclk));
	jdff dff_B_gUUhPHdx0_0(.din(w_dff_B_Zt8ILZVx8_0),.dout(w_dff_B_gUUhPHdx0_0),.clk(gclk));
	jdff dff_B_mhhPRSfj5_0(.din(w_dff_B_gUUhPHdx0_0),.dout(w_dff_B_mhhPRSfj5_0),.clk(gclk));
	jdff dff_B_x2Z9RvSJ7_0(.din(w_dff_B_mhhPRSfj5_0),.dout(w_dff_B_x2Z9RvSJ7_0),.clk(gclk));
	jdff dff_B_ElOjTrJk8_0(.din(w_dff_B_x2Z9RvSJ7_0),.dout(w_dff_B_ElOjTrJk8_0),.clk(gclk));
	jdff dff_B_6a3XpskK7_0(.din(w_dff_B_ElOjTrJk8_0),.dout(w_dff_B_6a3XpskK7_0),.clk(gclk));
	jdff dff_B_bLwZTJWi7_0(.din(w_dff_B_6a3XpskK7_0),.dout(w_dff_B_bLwZTJWi7_0),.clk(gclk));
	jdff dff_B_OUDgAJoO4_0(.din(w_dff_B_bLwZTJWi7_0),.dout(w_dff_B_OUDgAJoO4_0),.clk(gclk));
	jdff dff_B_rwukpntz1_0(.din(w_dff_B_OUDgAJoO4_0),.dout(w_dff_B_rwukpntz1_0),.clk(gclk));
	jdff dff_B_9FbwB4DN9_0(.din(w_dff_B_rwukpntz1_0),.dout(w_dff_B_9FbwB4DN9_0),.clk(gclk));
	jdff dff_B_4EJ33MHl7_0(.din(w_dff_B_9FbwB4DN9_0),.dout(w_dff_B_4EJ33MHl7_0),.clk(gclk));
	jdff dff_B_reTKQ3Mt8_0(.din(w_dff_B_4EJ33MHl7_0),.dout(w_dff_B_reTKQ3Mt8_0),.clk(gclk));
	jdff dff_B_GQZn4cF11_0(.din(w_dff_B_reTKQ3Mt8_0),.dout(w_dff_B_GQZn4cF11_0),.clk(gclk));
	jdff dff_B_AXN5zYGA4_0(.din(w_dff_B_GQZn4cF11_0),.dout(w_dff_B_AXN5zYGA4_0),.clk(gclk));
	jdff dff_B_2738FR838_0(.din(n1474),.dout(w_dff_B_2738FR838_0),.clk(gclk));
	jdff dff_B_mQA7HCfO5_0(.din(w_dff_B_2738FR838_0),.dout(w_dff_B_mQA7HCfO5_0),.clk(gclk));
	jdff dff_B_8fkx1HXv7_0(.din(w_dff_B_mQA7HCfO5_0),.dout(w_dff_B_8fkx1HXv7_0),.clk(gclk));
	jdff dff_B_HGeN4flO9_0(.din(w_dff_B_8fkx1HXv7_0),.dout(w_dff_B_HGeN4flO9_0),.clk(gclk));
	jdff dff_B_u2t1JI6M1_0(.din(w_dff_B_HGeN4flO9_0),.dout(w_dff_B_u2t1JI6M1_0),.clk(gclk));
	jdff dff_B_Jbq6DmhX3_0(.din(w_dff_B_u2t1JI6M1_0),.dout(w_dff_B_Jbq6DmhX3_0),.clk(gclk));
	jdff dff_B_rqNvkiyT5_0(.din(w_dff_B_Jbq6DmhX3_0),.dout(w_dff_B_rqNvkiyT5_0),.clk(gclk));
	jdff dff_B_80hPncZ95_0(.din(w_dff_B_rqNvkiyT5_0),.dout(w_dff_B_80hPncZ95_0),.clk(gclk));
	jdff dff_B_S7F6LStF1_0(.din(w_dff_B_80hPncZ95_0),.dout(w_dff_B_S7F6LStF1_0),.clk(gclk));
	jdff dff_B_BRMmmpfL0_0(.din(w_dff_B_S7F6LStF1_0),.dout(w_dff_B_BRMmmpfL0_0),.clk(gclk));
	jdff dff_B_nRPVgKWW5_0(.din(w_dff_B_BRMmmpfL0_0),.dout(w_dff_B_nRPVgKWW5_0),.clk(gclk));
	jdff dff_B_8kAVW8gB0_0(.din(w_dff_B_nRPVgKWW5_0),.dout(w_dff_B_8kAVW8gB0_0),.clk(gclk));
	jdff dff_B_GmWRTMoa6_0(.din(w_dff_B_8kAVW8gB0_0),.dout(w_dff_B_GmWRTMoa6_0),.clk(gclk));
	jdff dff_B_d4kiu3Y44_0(.din(w_dff_B_GmWRTMoa6_0),.dout(w_dff_B_d4kiu3Y44_0),.clk(gclk));
	jdff dff_B_GfyjoT731_0(.din(w_dff_B_d4kiu3Y44_0),.dout(w_dff_B_GfyjoT731_0),.clk(gclk));
	jdff dff_B_hephm8TV5_0(.din(n1473),.dout(w_dff_B_hephm8TV5_0),.clk(gclk));
	jdff dff_B_mxWw4cXU4_0(.din(n1469),.dout(w_dff_B_mxWw4cXU4_0),.clk(gclk));
	jdff dff_B_JFGY0C2l5_0(.din(n1465),.dout(w_dff_B_JFGY0C2l5_0),.clk(gclk));
	jdff dff_B_ACIfsFgv6_0(.din(w_dff_B_JFGY0C2l5_0),.dout(w_dff_B_ACIfsFgv6_0),.clk(gclk));
	jdff dff_B_oAbW667H2_0(.din(w_dff_B_ACIfsFgv6_0),.dout(w_dff_B_oAbW667H2_0),.clk(gclk));
	jdff dff_B_Rsfrln7j2_0(.din(w_dff_B_oAbW667H2_0),.dout(w_dff_B_Rsfrln7j2_0),.clk(gclk));
	jdff dff_B_8IkfZdUQ2_0(.din(w_dff_B_Rsfrln7j2_0),.dout(w_dff_B_8IkfZdUQ2_0),.clk(gclk));
	jdff dff_B_jZ7TKH3V2_0(.din(w_dff_B_8IkfZdUQ2_0),.dout(w_dff_B_jZ7TKH3V2_0),.clk(gclk));
	jdff dff_B_ICu2GORB2_0(.din(w_dff_B_jZ7TKH3V2_0),.dout(w_dff_B_ICu2GORB2_0),.clk(gclk));
	jdff dff_B_dNevHoGM4_0(.din(w_dff_B_ICu2GORB2_0),.dout(w_dff_B_dNevHoGM4_0),.clk(gclk));
	jdff dff_B_W25aDOCw2_0(.din(w_dff_B_dNevHoGM4_0),.dout(w_dff_B_W25aDOCw2_0),.clk(gclk));
	jdff dff_B_uJpGYrPR3_0(.din(w_dff_B_W25aDOCw2_0),.dout(w_dff_B_uJpGYrPR3_0),.clk(gclk));
	jdff dff_B_7mnuJ1KH0_0(.din(w_dff_B_uJpGYrPR3_0),.dout(w_dff_B_7mnuJ1KH0_0),.clk(gclk));
	jdff dff_B_s4mshVr45_0(.din(w_dff_B_7mnuJ1KH0_0),.dout(w_dff_B_s4mshVr45_0),.clk(gclk));
	jdff dff_B_INOpmN2v9_0(.din(w_dff_B_s4mshVr45_0),.dout(w_dff_B_INOpmN2v9_0),.clk(gclk));
	jdff dff_B_PL1JEJ9U9_1(.din(n1451),.dout(w_dff_B_PL1JEJ9U9_1),.clk(gclk));
	jdff dff_B_1FyWNS501_0(.din(n1463),.dout(w_dff_B_1FyWNS501_0),.clk(gclk));
	jdff dff_B_NozrAiAC0_0(.din(w_dff_B_1FyWNS501_0),.dout(w_dff_B_NozrAiAC0_0),.clk(gclk));
	jdff dff_B_b9b3rXR82_0(.din(w_dff_B_NozrAiAC0_0),.dout(w_dff_B_b9b3rXR82_0),.clk(gclk));
	jdff dff_B_KYND4Y7A2_0(.din(n1461),.dout(w_dff_B_KYND4Y7A2_0),.clk(gclk));
	jdff dff_B_ew9BjGEv2_1(.din(n1453),.dout(w_dff_B_ew9BjGEv2_1),.clk(gclk));
	jdff dff_B_8MmWqEbC1_1(.din(w_dff_B_ew9BjGEv2_1),.dout(w_dff_B_8MmWqEbC1_1),.clk(gclk));
	jdff dff_B_yv0IKcgm6_0(.din(n1454),.dout(w_dff_B_yv0IKcgm6_0),.clk(gclk));
	jdff dff_B_N2OCdIRW9_0(.din(w_dff_B_yv0IKcgm6_0),.dout(w_dff_B_N2OCdIRW9_0),.clk(gclk));
	jdff dff_B_xpKKAL3M3_0(.din(w_dff_B_N2OCdIRW9_0),.dout(w_dff_B_xpKKAL3M3_0),.clk(gclk));
	jdff dff_B_lc2rTYBf5_0(.din(w_dff_B_xpKKAL3M3_0),.dout(w_dff_B_lc2rTYBf5_0),.clk(gclk));
	jdff dff_A_719EER1D0_0(.dout(w_n1452_0[0]),.din(w_dff_A_719EER1D0_0),.clk(gclk));
	jdff dff_A_OjBgAxHs3_0(.dout(w_dff_A_719EER1D0_0),.din(w_dff_A_OjBgAxHs3_0),.clk(gclk));
	jdff dff_A_W0PFkf9e6_0(.dout(w_dff_A_OjBgAxHs3_0),.din(w_dff_A_W0PFkf9e6_0),.clk(gclk));
	jdff dff_A_TtsvZyKe2_0(.dout(w_dff_A_W0PFkf9e6_0),.din(w_dff_A_TtsvZyKe2_0),.clk(gclk));
	jdff dff_A_gbJB54ha2_2(.dout(w_n1452_0[2]),.din(w_dff_A_gbJB54ha2_2),.clk(gclk));
	jdff dff_A_PzrwB98c9_2(.dout(w_dff_A_gbJB54ha2_2),.din(w_dff_A_PzrwB98c9_2),.clk(gclk));
	jdff dff_A_7oZDXmlx4_2(.dout(w_dff_A_PzrwB98c9_2),.din(w_dff_A_7oZDXmlx4_2),.clk(gclk));
	jdff dff_A_krkk7XAh3_1(.dout(w_n1340_0[1]),.din(w_dff_A_krkk7XAh3_1),.clk(gclk));
	jdff dff_A_aBj6fkYF0_2(.dout(w_n1340_0[2]),.din(w_dff_A_aBj6fkYF0_2),.clk(gclk));
	jdff dff_A_2zKwrxka1_2(.dout(w_dff_A_aBj6fkYF0_2),.din(w_dff_A_2zKwrxka1_2),.clk(gclk));
	jdff dff_A_HUrhjDSj0_2(.dout(w_dff_A_2zKwrxka1_2),.din(w_dff_A_HUrhjDSj0_2),.clk(gclk));
	jdff dff_A_beI3AcAP1_2(.dout(w_dff_A_HUrhjDSj0_2),.din(w_dff_A_beI3AcAP1_2),.clk(gclk));
	jdff dff_A_QhrjhUhk6_2(.dout(w_dff_A_beI3AcAP1_2),.din(w_dff_A_QhrjhUhk6_2),.clk(gclk));
	jdff dff_A_5r8eP85j4_2(.dout(w_dff_A_QhrjhUhk6_2),.din(w_dff_A_5r8eP85j4_2),.clk(gclk));
	jdff dff_A_WEP0MKFF0_2(.dout(w_dff_A_5r8eP85j4_2),.din(w_dff_A_WEP0MKFF0_2),.clk(gclk));
	jdff dff_A_YrUKhixG1_2(.dout(w_dff_A_WEP0MKFF0_2),.din(w_dff_A_YrUKhixG1_2),.clk(gclk));
	jdff dff_A_eIOkxsDs3_2(.dout(w_dff_A_YrUKhixG1_2),.din(w_dff_A_eIOkxsDs3_2),.clk(gclk));
	jdff dff_A_q5O3GhCj0_2(.dout(w_dff_A_eIOkxsDs3_2),.din(w_dff_A_q5O3GhCj0_2),.clk(gclk));
	jdff dff_A_LsF4A0HY3_2(.dout(w_dff_A_q5O3GhCj0_2),.din(w_dff_A_LsF4A0HY3_2),.clk(gclk));
	jdff dff_A_jtg43NQK5_2(.dout(w_dff_A_LsF4A0HY3_2),.din(w_dff_A_jtg43NQK5_2),.clk(gclk));
	jdff dff_A_7yNIHFGd2_2(.dout(w_dff_A_jtg43NQK5_2),.din(w_dff_A_7yNIHFGd2_2),.clk(gclk));
	jdff dff_A_QcorbPoi1_2(.dout(w_dff_A_7yNIHFGd2_2),.din(w_dff_A_QcorbPoi1_2),.clk(gclk));
	jdff dff_A_ePWatc187_2(.dout(w_dff_A_QcorbPoi1_2),.din(w_dff_A_ePWatc187_2),.clk(gclk));
	jdff dff_A_XQE8hrzm9_2(.dout(w_dff_A_ePWatc187_2),.din(w_dff_A_XQE8hrzm9_2),.clk(gclk));
	jdff dff_A_gUPboYWa9_2(.dout(w_dff_A_XQE8hrzm9_2),.din(w_dff_A_gUPboYWa9_2),.clk(gclk));
	jdff dff_A_t7SZ7ibq3_2(.dout(w_dff_A_gUPboYWa9_2),.din(w_dff_A_t7SZ7ibq3_2),.clk(gclk));
	jdff dff_A_i00KGOL32_2(.dout(w_dff_A_t7SZ7ibq3_2),.din(w_dff_A_i00KGOL32_2),.clk(gclk));
	jdff dff_A_HvtO3RM12_2(.dout(w_dff_A_i00KGOL32_2),.din(w_dff_A_HvtO3RM12_2),.clk(gclk));
	jdff dff_A_jJI5G6gM5_2(.dout(w_dff_A_HvtO3RM12_2),.din(w_dff_A_jJI5G6gM5_2),.clk(gclk));
	jdff dff_B_VayDGo799_3(.din(n1340),.dout(w_dff_B_VayDGo799_3),.clk(gclk));
	jdff dff_B_rDo5NBVx2_3(.din(w_dff_B_VayDGo799_3),.dout(w_dff_B_rDo5NBVx2_3),.clk(gclk));
	jdff dff_B_tof5vAxJ8_3(.din(w_dff_B_rDo5NBVx2_3),.dout(w_dff_B_tof5vAxJ8_3),.clk(gclk));
	jdff dff_B_ijaMgSks0_0(.din(n1447),.dout(w_dff_B_ijaMgSks0_0),.clk(gclk));
	jdff dff_B_3rEMfBpF3_0(.din(w_dff_B_ijaMgSks0_0),.dout(w_dff_B_3rEMfBpF3_0),.clk(gclk));
	jdff dff_B_hK5XbLPc3_0(.din(w_dff_B_3rEMfBpF3_0),.dout(w_dff_B_hK5XbLPc3_0),.clk(gclk));
	jdff dff_B_bzBj97qH0_0(.din(w_dff_B_hK5XbLPc3_0),.dout(w_dff_B_bzBj97qH0_0),.clk(gclk));
	jdff dff_B_GAaUEI6x9_0(.din(w_dff_B_bzBj97qH0_0),.dout(w_dff_B_GAaUEI6x9_0),.clk(gclk));
	jdff dff_B_Mv1xrPiQ3_0(.din(w_dff_B_GAaUEI6x9_0),.dout(w_dff_B_Mv1xrPiQ3_0),.clk(gclk));
	jdff dff_B_r8l9RA577_0(.din(w_dff_B_Mv1xrPiQ3_0),.dout(w_dff_B_r8l9RA577_0),.clk(gclk));
	jdff dff_B_ChH0EEBX8_0(.din(w_dff_B_r8l9RA577_0),.dout(w_dff_B_ChH0EEBX8_0),.clk(gclk));
	jdff dff_B_BSKntXx67_0(.din(w_dff_B_ChH0EEBX8_0),.dout(w_dff_B_BSKntXx67_0),.clk(gclk));
	jdff dff_B_77aDa9LM9_0(.din(w_dff_B_BSKntXx67_0),.dout(w_dff_B_77aDa9LM9_0),.clk(gclk));
	jdff dff_B_UtGWPSW14_0(.din(w_dff_B_77aDa9LM9_0),.dout(w_dff_B_UtGWPSW14_0),.clk(gclk));
	jdff dff_B_B4SL31yq2_0(.din(w_dff_B_UtGWPSW14_0),.dout(w_dff_B_B4SL31yq2_0),.clk(gclk));
	jdff dff_B_zfRgEin34_0(.din(w_dff_B_B4SL31yq2_0),.dout(w_dff_B_zfRgEin34_0),.clk(gclk));
	jdff dff_B_86m7VksF8_0(.din(w_dff_B_zfRgEin34_0),.dout(w_dff_B_86m7VksF8_0),.clk(gclk));
	jdff dff_B_5avHTFlS5_0(.din(w_dff_B_86m7VksF8_0),.dout(w_dff_B_5avHTFlS5_0),.clk(gclk));
	jdff dff_B_UAJSjZ4p4_0(.din(w_dff_B_5avHTFlS5_0),.dout(w_dff_B_UAJSjZ4p4_0),.clk(gclk));
	jdff dff_B_xP21tEYM0_0(.din(w_dff_B_UAJSjZ4p4_0),.dout(w_dff_B_xP21tEYM0_0),.clk(gclk));
	jdff dff_B_fYPvapMd8_0(.din(w_dff_B_xP21tEYM0_0),.dout(w_dff_B_fYPvapMd8_0),.clk(gclk));
	jdff dff_B_NGsbwMpe2_0(.din(w_dff_B_fYPvapMd8_0),.dout(w_dff_B_NGsbwMpe2_0),.clk(gclk));
	jdff dff_B_4HAgZNzg2_1(.din(n1445),.dout(w_dff_B_4HAgZNzg2_1),.clk(gclk));
	jdff dff_B_nuGxlRcY6_0(.din(n1444),.dout(w_dff_B_nuGxlRcY6_0),.clk(gclk));
	jdff dff_B_V51AO53A2_0(.din(w_dff_B_nuGxlRcY6_0),.dout(w_dff_B_V51AO53A2_0),.clk(gclk));
	jdff dff_B_pUYv3kJb8_0(.din(n1441),.dout(w_dff_B_pUYv3kJb8_0),.clk(gclk));
	jdff dff_B_8p8f9pN02_0(.din(n1438),.dout(w_dff_B_8p8f9pN02_0),.clk(gclk));
	jdff dff_B_eDA1cr683_0(.din(w_dff_B_8p8f9pN02_0),.dout(w_dff_B_eDA1cr683_0),.clk(gclk));
	jdff dff_B_2NVuRVOw5_0(.din(w_dff_B_eDA1cr683_0),.dout(w_dff_B_2NVuRVOw5_0),.clk(gclk));
	jdff dff_B_Hr4UWyl12_0(.din(w_dff_B_2NVuRVOw5_0),.dout(w_dff_B_Hr4UWyl12_0),.clk(gclk));
	jdff dff_B_CXgMz9647_0(.din(w_dff_B_Hr4UWyl12_0),.dout(w_dff_B_CXgMz9647_0),.clk(gclk));
	jdff dff_B_OERe5ODg6_0(.din(w_dff_B_CXgMz9647_0),.dout(w_dff_B_OERe5ODg6_0),.clk(gclk));
	jdff dff_B_ImMSh5TZ2_0(.din(w_dff_B_OERe5ODg6_0),.dout(w_dff_B_ImMSh5TZ2_0),.clk(gclk));
	jdff dff_B_QaXdQIWl1_0(.din(w_dff_B_ImMSh5TZ2_0),.dout(w_dff_B_QaXdQIWl1_0),.clk(gclk));
	jdff dff_B_1YZVfkZN3_0(.din(w_dff_B_QaXdQIWl1_0),.dout(w_dff_B_1YZVfkZN3_0),.clk(gclk));
	jdff dff_B_6rUDTuxD3_0(.din(w_dff_B_1YZVfkZN3_0),.dout(w_dff_B_6rUDTuxD3_0),.clk(gclk));
	jdff dff_B_6lcabkyl5_0(.din(w_dff_B_6rUDTuxD3_0),.dout(w_dff_B_6lcabkyl5_0),.clk(gclk));
	jdff dff_B_YhVmrNL97_0(.din(w_dff_B_6lcabkyl5_0),.dout(w_dff_B_YhVmrNL97_0),.clk(gclk));
	jdff dff_B_mSlToNXx6_0(.din(w_dff_B_YhVmrNL97_0),.dout(w_dff_B_mSlToNXx6_0),.clk(gclk));
	jdff dff_B_MefwuRR94_0(.din(w_dff_B_mSlToNXx6_0),.dout(w_dff_B_MefwuRR94_0),.clk(gclk));
	jdff dff_B_3xR3Qjsu8_0(.din(w_dff_B_MefwuRR94_0),.dout(w_dff_B_3xR3Qjsu8_0),.clk(gclk));
	jdff dff_B_wgTQbKLv9_0(.din(w_dff_B_3xR3Qjsu8_0),.dout(w_dff_B_wgTQbKLv9_0),.clk(gclk));
	jdff dff_B_MG03m1yT9_0(.din(w_dff_B_wgTQbKLv9_0),.dout(w_dff_B_MG03m1yT9_0),.clk(gclk));
	jdff dff_B_hYjjC3xx1_0(.din(w_dff_B_MG03m1yT9_0),.dout(w_dff_B_hYjjC3xx1_0),.clk(gclk));
	jdff dff_B_kGTsVbyO2_0(.din(w_dff_B_hYjjC3xx1_0),.dout(w_dff_B_kGTsVbyO2_0),.clk(gclk));
	jdff dff_B_bZewYbaQ4_0(.din(n1437),.dout(w_dff_B_bZewYbaQ4_0),.clk(gclk));
	jdff dff_B_Jyi5VW8h0_1(.din(n1432),.dout(w_dff_B_Jyi5VW8h0_1),.clk(gclk));
	jdff dff_A_ND9Xw4v67_1(.dout(w_n1388_0[1]),.din(w_dff_A_ND9Xw4v67_1),.clk(gclk));
	jdff dff_A_x46G1Kg41_1(.dout(w_dff_A_ND9Xw4v67_1),.din(w_dff_A_x46G1Kg41_1),.clk(gclk));
	jdff dff_A_mBJj3KzO0_1(.dout(w_dff_A_x46G1Kg41_1),.din(w_dff_A_mBJj3KzO0_1),.clk(gclk));
	jdff dff_A_YbNCaeJ37_1(.dout(w_dff_A_mBJj3KzO0_1),.din(w_dff_A_YbNCaeJ37_1),.clk(gclk));
	jdff dff_A_oTD6dlzB2_1(.dout(w_dff_A_YbNCaeJ37_1),.din(w_dff_A_oTD6dlzB2_1),.clk(gclk));
	jdff dff_A_OgqFqi3b7_1(.dout(w_dff_A_oTD6dlzB2_1),.din(w_dff_A_OgqFqi3b7_1),.clk(gclk));
	jdff dff_A_Ou7NyWKl8_1(.dout(w_dff_A_OgqFqi3b7_1),.din(w_dff_A_Ou7NyWKl8_1),.clk(gclk));
	jdff dff_A_Y6s8OPQO9_1(.dout(w_dff_A_Ou7NyWKl8_1),.din(w_dff_A_Y6s8OPQO9_1),.clk(gclk));
	jdff dff_A_2VYW4K1v6_1(.dout(w_dff_A_Y6s8OPQO9_1),.din(w_dff_A_2VYW4K1v6_1),.clk(gclk));
	jdff dff_A_7fH6kUON8_1(.dout(w_dff_A_2VYW4K1v6_1),.din(w_dff_A_7fH6kUON8_1),.clk(gclk));
	jdff dff_A_cevX7o0u9_1(.dout(w_dff_A_7fH6kUON8_1),.din(w_dff_A_cevX7o0u9_1),.clk(gclk));
	jdff dff_A_b4P4GOG36_1(.dout(w_dff_A_cevX7o0u9_1),.din(w_dff_A_b4P4GOG36_1),.clk(gclk));
	jdff dff_A_tEyVDrMj6_1(.dout(w_dff_A_b4P4GOG36_1),.din(w_dff_A_tEyVDrMj6_1),.clk(gclk));
	jdff dff_A_zVfKWdjQ9_1(.dout(w_dff_A_tEyVDrMj6_1),.din(w_dff_A_zVfKWdjQ9_1),.clk(gclk));
	jdff dff_A_CAAk2uRn9_1(.dout(w_dff_A_zVfKWdjQ9_1),.din(w_dff_A_CAAk2uRn9_1),.clk(gclk));
	jdff dff_A_PIqAJi5a8_1(.dout(w_dff_A_CAAk2uRn9_1),.din(w_dff_A_PIqAJi5a8_1),.clk(gclk));
	jdff dff_A_3NmO94mg2_1(.dout(w_dff_A_PIqAJi5a8_1),.din(w_dff_A_3NmO94mg2_1),.clk(gclk));
	jdff dff_A_3IP9oUZD1_1(.dout(w_dff_A_3NmO94mg2_1),.din(w_dff_A_3IP9oUZD1_1),.clk(gclk));
	jdff dff_A_qc6uFhI29_1(.dout(w_dff_A_3IP9oUZD1_1),.din(w_dff_A_qc6uFhI29_1),.clk(gclk));
	jdff dff_A_fQOs5RJI0_1(.dout(w_dff_A_qc6uFhI29_1),.din(w_dff_A_fQOs5RJI0_1),.clk(gclk));
	jdff dff_A_cHkkuZrw5_1(.dout(w_dff_A_fQOs5RJI0_1),.din(w_dff_A_cHkkuZrw5_1),.clk(gclk));
	jdff dff_A_yBrlKAMT0_1(.dout(w_dff_A_cHkkuZrw5_1),.din(w_dff_A_yBrlKAMT0_1),.clk(gclk));
	jdff dff_A_L37J9nCp5_1(.dout(w_dff_A_yBrlKAMT0_1),.din(w_dff_A_L37J9nCp5_1),.clk(gclk));
	jdff dff_A_Xlj8jfvv7_1(.dout(w_dff_A_L37J9nCp5_1),.din(w_dff_A_Xlj8jfvv7_1),.clk(gclk));
	jdff dff_A_LPFnN2Nq5_1(.dout(w_dff_A_Xlj8jfvv7_1),.din(w_dff_A_LPFnN2Nq5_1),.clk(gclk));
	jdff dff_A_UTUX7qT57_0(.dout(w_n1387_0[0]),.din(w_dff_A_UTUX7qT57_0),.clk(gclk));
	jdff dff_A_aqmJyNgr3_0(.dout(w_dff_A_UTUX7qT57_0),.din(w_dff_A_aqmJyNgr3_0),.clk(gclk));
	jdff dff_B_M4BynVLC9_2(.din(n1431),.dout(w_dff_B_M4BynVLC9_2),.clk(gclk));
	jdff dff_B_cUsg1qKh9_2(.din(w_dff_B_M4BynVLC9_2),.dout(w_dff_B_cUsg1qKh9_2),.clk(gclk));
	jdff dff_B_0E7z0d090_2(.din(w_dff_B_cUsg1qKh9_2),.dout(w_dff_B_0E7z0d090_2),.clk(gclk));
	jdff dff_B_34c1KuyF5_2(.din(w_dff_B_0E7z0d090_2),.dout(w_dff_B_34c1KuyF5_2),.clk(gclk));
	jdff dff_B_7Lz0IC683_0(.din(n1526),.dout(w_dff_B_7Lz0IC683_0),.clk(gclk));
	jdff dff_B_Tq42sKlL7_0(.din(n1524),.dout(w_dff_B_Tq42sKlL7_0),.clk(gclk));
	jdff dff_B_QJJewbSj4_0(.din(w_dff_B_Tq42sKlL7_0),.dout(w_dff_B_QJJewbSj4_0),.clk(gclk));
	jdff dff_B_1AgZ3Bjn8_0(.din(w_dff_B_QJJewbSj4_0),.dout(w_dff_B_1AgZ3Bjn8_0),.clk(gclk));
	jdff dff_B_whGa9iPH5_0(.din(w_dff_B_1AgZ3Bjn8_0),.dout(w_dff_B_whGa9iPH5_0),.clk(gclk));
	jdff dff_B_1AnSKQfI2_0(.din(w_dff_B_whGa9iPH5_0),.dout(w_dff_B_1AnSKQfI2_0),.clk(gclk));
	jdff dff_B_REgLsSAk6_0(.din(w_dff_B_1AnSKQfI2_0),.dout(w_dff_B_REgLsSAk6_0),.clk(gclk));
	jdff dff_B_yoFNMVqF6_0(.din(w_dff_B_REgLsSAk6_0),.dout(w_dff_B_yoFNMVqF6_0),.clk(gclk));
	jdff dff_B_LO8MsGPn6_0(.din(w_dff_B_yoFNMVqF6_0),.dout(w_dff_B_LO8MsGPn6_0),.clk(gclk));
	jdff dff_B_MPZomksl0_0(.din(w_dff_B_LO8MsGPn6_0),.dout(w_dff_B_MPZomksl0_0),.clk(gclk));
	jdff dff_B_qPloL37m9_0(.din(w_dff_B_MPZomksl0_0),.dout(w_dff_B_qPloL37m9_0),.clk(gclk));
	jdff dff_B_EQRiOYtZ7_0(.din(w_dff_B_qPloL37m9_0),.dout(w_dff_B_EQRiOYtZ7_0),.clk(gclk));
	jdff dff_B_5qvJ2mKi1_0(.din(w_dff_B_EQRiOYtZ7_0),.dout(w_dff_B_5qvJ2mKi1_0),.clk(gclk));
	jdff dff_B_VEzlivPG9_0(.din(w_dff_B_5qvJ2mKi1_0),.dout(w_dff_B_VEzlivPG9_0),.clk(gclk));
	jdff dff_B_luoQV8yu9_0(.din(w_dff_B_VEzlivPG9_0),.dout(w_dff_B_luoQV8yu9_0),.clk(gclk));
	jdff dff_B_l96kWJPL1_0(.din(w_dff_B_luoQV8yu9_0),.dout(w_dff_B_l96kWJPL1_0),.clk(gclk));
	jdff dff_B_lT3Pp4zg7_0(.din(w_dff_B_l96kWJPL1_0),.dout(w_dff_B_lT3Pp4zg7_0),.clk(gclk));
	jdff dff_B_JykNhceB1_0(.din(w_dff_B_lT3Pp4zg7_0),.dout(w_dff_B_JykNhceB1_0),.clk(gclk));
	jdff dff_B_JwRnG0pd9_0(.din(n1523),.dout(w_dff_B_JwRnG0pd9_0),.clk(gclk));
	jdff dff_A_8AxGSzgb4_1(.dout(w_n420_0[1]),.din(w_dff_A_8AxGSzgb4_1),.clk(gclk));
	jdff dff_A_GAnxm2I85_1(.dout(w_dff_A_8AxGSzgb4_1),.din(w_dff_A_GAnxm2I85_1),.clk(gclk));
	jdff dff_A_t9iASt3X5_1(.dout(w_dff_A_GAnxm2I85_1),.din(w_dff_A_t9iASt3X5_1),.clk(gclk));
	jdff dff_A_zV6UWLfI6_1(.dout(w_dff_A_t9iASt3X5_1),.din(w_dff_A_zV6UWLfI6_1),.clk(gclk));
	jdff dff_A_7y77P9SC0_1(.dout(w_dff_A_zV6UWLfI6_1),.din(w_dff_A_7y77P9SC0_1),.clk(gclk));
	jdff dff_A_2RVeAT833_1(.dout(w_dff_A_7y77P9SC0_1),.din(w_dff_A_2RVeAT833_1),.clk(gclk));
	jdff dff_A_e9Go8sPr9_1(.dout(w_dff_A_2RVeAT833_1),.din(w_dff_A_e9Go8sPr9_1),.clk(gclk));
	jdff dff_A_HxTrJinE0_1(.dout(w_dff_A_e9Go8sPr9_1),.din(w_dff_A_HxTrJinE0_1),.clk(gclk));
	jdff dff_A_nYkfMcrM3_1(.dout(w_dff_A_HxTrJinE0_1),.din(w_dff_A_nYkfMcrM3_1),.clk(gclk));
	jdff dff_A_hbPUZvC87_1(.dout(w_dff_A_nYkfMcrM3_1),.din(w_dff_A_hbPUZvC87_1),.clk(gclk));
	jdff dff_A_OZqdLF5D0_1(.dout(w_dff_A_hbPUZvC87_1),.din(w_dff_A_OZqdLF5D0_1),.clk(gclk));
	jdff dff_A_dEH2fRdO4_1(.dout(w_dff_A_OZqdLF5D0_1),.din(w_dff_A_dEH2fRdO4_1),.clk(gclk));
	jdff dff_A_aspEWJ8J4_1(.dout(w_dff_A_dEH2fRdO4_1),.din(w_dff_A_aspEWJ8J4_1),.clk(gclk));
	jdff dff_A_UPBiKVTm1_1(.dout(w_dff_A_aspEWJ8J4_1),.din(w_dff_A_UPBiKVTm1_1),.clk(gclk));
	jdff dff_A_mxFMN0K67_1(.dout(w_dff_A_UPBiKVTm1_1),.din(w_dff_A_mxFMN0K67_1),.clk(gclk));
	jdff dff_A_r997vqh18_1(.dout(w_dff_A_mxFMN0K67_1),.din(w_dff_A_r997vqh18_1),.clk(gclk));
	jdff dff_A_en48fLNx7_1(.dout(w_dff_A_r997vqh18_1),.din(w_dff_A_en48fLNx7_1),.clk(gclk));
	jdff dff_A_eIgdf5oS8_1(.dout(w_dff_A_en48fLNx7_1),.din(w_dff_A_eIgdf5oS8_1),.clk(gclk));
	jdff dff_A_b6NpkqnL3_1(.dout(w_dff_A_eIgdf5oS8_1),.din(w_dff_A_b6NpkqnL3_1),.clk(gclk));
	jdff dff_A_l9fYWk477_1(.dout(w_dff_A_b6NpkqnL3_1),.din(w_dff_A_l9fYWk477_1),.clk(gclk));
	jdff dff_A_keEUnYQ00_1(.dout(w_dff_A_l9fYWk477_1),.din(w_dff_A_keEUnYQ00_1),.clk(gclk));
	jdff dff_A_M7KmyMdH9_0(.dout(w_n413_1[0]),.din(w_dff_A_M7KmyMdH9_0),.clk(gclk));
	jdff dff_A_tpY9nJRG5_0(.dout(w_dff_A_M7KmyMdH9_0),.din(w_dff_A_tpY9nJRG5_0),.clk(gclk));
	jdff dff_A_FNA0fCSX4_0(.dout(w_dff_A_tpY9nJRG5_0),.din(w_dff_A_FNA0fCSX4_0),.clk(gclk));
	jdff dff_A_cnEMWUXq2_0(.dout(w_dff_A_FNA0fCSX4_0),.din(w_dff_A_cnEMWUXq2_0),.clk(gclk));
	jdff dff_A_JkaivZjF0_0(.dout(w_dff_A_cnEMWUXq2_0),.din(w_dff_A_JkaivZjF0_0),.clk(gclk));
	jdff dff_A_OEgsPleW8_0(.dout(w_dff_A_JkaivZjF0_0),.din(w_dff_A_OEgsPleW8_0),.clk(gclk));
	jdff dff_A_l1KiWBJ80_0(.dout(w_dff_A_OEgsPleW8_0),.din(w_dff_A_l1KiWBJ80_0),.clk(gclk));
	jdff dff_A_7L673EWa7_0(.dout(w_dff_A_l1KiWBJ80_0),.din(w_dff_A_7L673EWa7_0),.clk(gclk));
	jdff dff_A_QgYzijuN2_0(.dout(w_dff_A_7L673EWa7_0),.din(w_dff_A_QgYzijuN2_0),.clk(gclk));
	jdff dff_A_Edtt8bzm2_0(.dout(w_dff_A_QgYzijuN2_0),.din(w_dff_A_Edtt8bzm2_0),.clk(gclk));
	jdff dff_A_bcSouc1D2_0(.dout(w_dff_A_Edtt8bzm2_0),.din(w_dff_A_bcSouc1D2_0),.clk(gclk));
	jdff dff_A_36YJjSOi8_0(.dout(w_dff_A_bcSouc1D2_0),.din(w_dff_A_36YJjSOi8_0),.clk(gclk));
	jdff dff_A_cC7PaEWc9_0(.dout(w_dff_A_36YJjSOi8_0),.din(w_dff_A_cC7PaEWc9_0),.clk(gclk));
	jdff dff_A_CaRJ8C2P2_0(.dout(w_dff_A_cC7PaEWc9_0),.din(w_dff_A_CaRJ8C2P2_0),.clk(gclk));
	jdff dff_A_AR8wxLEs0_0(.dout(w_dff_A_CaRJ8C2P2_0),.din(w_dff_A_AR8wxLEs0_0),.clk(gclk));
	jdff dff_A_Uv5lnRWA8_0(.dout(w_dff_A_AR8wxLEs0_0),.din(w_dff_A_Uv5lnRWA8_0),.clk(gclk));
	jdff dff_A_iMxzCyTs2_0(.dout(w_dff_A_Uv5lnRWA8_0),.din(w_dff_A_iMxzCyTs2_0),.clk(gclk));
	jdff dff_A_xpiY8Ufd5_0(.dout(w_dff_A_iMxzCyTs2_0),.din(w_dff_A_xpiY8Ufd5_0),.clk(gclk));
	jdff dff_A_liH9GRf56_0(.dout(w_dff_A_xpiY8Ufd5_0),.din(w_dff_A_liH9GRf56_0),.clk(gclk));
	jdff dff_A_9gO6g7tX7_0(.dout(w_dff_A_liH9GRf56_0),.din(w_dff_A_9gO6g7tX7_0),.clk(gclk));
	jdff dff_A_msS3zn0b7_0(.dout(w_dff_A_9gO6g7tX7_0),.din(w_dff_A_msS3zn0b7_0),.clk(gclk));
	jdff dff_B_OnYKiijy7_1(.din(n1521),.dout(w_dff_B_OnYKiijy7_1),.clk(gclk));
	jdff dff_B_BwhpK7Re8_1(.din(w_dff_B_OnYKiijy7_1),.dout(w_dff_B_BwhpK7Re8_1),.clk(gclk));
	jdff dff_B_u7raKxTd3_1(.din(w_dff_B_BwhpK7Re8_1),.dout(w_dff_B_u7raKxTd3_1),.clk(gclk));
	jdff dff_B_p95jurqh9_1(.din(w_dff_B_u7raKxTd3_1),.dout(w_dff_B_p95jurqh9_1),.clk(gclk));
	jdff dff_B_rIxcZSoR5_1(.din(w_dff_B_p95jurqh9_1),.dout(w_dff_B_rIxcZSoR5_1),.clk(gclk));
	jdff dff_B_i4G7rVJD8_1(.din(w_dff_B_rIxcZSoR5_1),.dout(w_dff_B_i4G7rVJD8_1),.clk(gclk));
	jdff dff_B_28qkGFQB2_1(.din(w_dff_B_i4G7rVJD8_1),.dout(w_dff_B_28qkGFQB2_1),.clk(gclk));
	jdff dff_A_UHdhm1WF6_1(.dout(w_n419_0[1]),.din(w_dff_A_UHdhm1WF6_1),.clk(gclk));
	jdff dff_A_ThXDYTK74_1(.dout(w_dff_A_UHdhm1WF6_1),.din(w_dff_A_ThXDYTK74_1),.clk(gclk));
	jdff dff_A_wahFABi94_1(.dout(w_dff_A_ThXDYTK74_1),.din(w_dff_A_wahFABi94_1),.clk(gclk));
	jdff dff_A_qhGdko7W8_1(.dout(w_dff_A_wahFABi94_1),.din(w_dff_A_qhGdko7W8_1),.clk(gclk));
	jdff dff_A_oh1B2yho0_1(.dout(w_dff_A_qhGdko7W8_1),.din(w_dff_A_oh1B2yho0_1),.clk(gclk));
	jdff dff_A_StSoeVLD8_1(.dout(w_dff_A_oh1B2yho0_1),.din(w_dff_A_StSoeVLD8_1),.clk(gclk));
	jdff dff_B_oiF3CoFo6_0(.din(n1519),.dout(w_dff_B_oiF3CoFo6_0),.clk(gclk));
	jdff dff_B_K5OSU1ID5_0(.din(w_dff_B_oiF3CoFo6_0),.dout(w_dff_B_K5OSU1ID5_0),.clk(gclk));
	jdff dff_B_uYuGoqJ38_0(.din(w_dff_B_K5OSU1ID5_0),.dout(w_dff_B_uYuGoqJ38_0),.clk(gclk));
	jdff dff_B_5A1JMwbV0_0(.din(w_dff_B_uYuGoqJ38_0),.dout(w_dff_B_5A1JMwbV0_0),.clk(gclk));
	jdff dff_B_Bib73DXc3_0(.din(w_dff_B_5A1JMwbV0_0),.dout(w_dff_B_Bib73DXc3_0),.clk(gclk));
	jdff dff_B_gxFZF1cC6_0(.din(w_dff_B_Bib73DXc3_0),.dout(w_dff_B_gxFZF1cC6_0),.clk(gclk));
	jdff dff_B_T1a1nCr90_0(.din(w_dff_B_gxFZF1cC6_0),.dout(w_dff_B_T1a1nCr90_0),.clk(gclk));
	jdff dff_B_cmmUvgXQ2_0(.din(w_dff_B_T1a1nCr90_0),.dout(w_dff_B_cmmUvgXQ2_0),.clk(gclk));
	jdff dff_B_VcA1N3op7_0(.din(w_dff_B_cmmUvgXQ2_0),.dout(w_dff_B_VcA1N3op7_0),.clk(gclk));
	jdff dff_B_DpD6zRwG4_0(.din(w_dff_B_VcA1N3op7_0),.dout(w_dff_B_DpD6zRwG4_0),.clk(gclk));
	jdff dff_B_9EtzbZrf0_0(.din(w_dff_B_DpD6zRwG4_0),.dout(w_dff_B_9EtzbZrf0_0),.clk(gclk));
	jdff dff_B_shyeRnQy5_0(.din(w_dff_B_9EtzbZrf0_0),.dout(w_dff_B_shyeRnQy5_0),.clk(gclk));
	jdff dff_B_SzAEIMD45_0(.din(w_dff_B_shyeRnQy5_0),.dout(w_dff_B_SzAEIMD45_0),.clk(gclk));
	jdff dff_B_Dkxpceow1_0(.din(w_dff_B_SzAEIMD45_0),.dout(w_dff_B_Dkxpceow1_0),.clk(gclk));
	jdff dff_B_ir71D0UF7_0(.din(w_dff_B_Dkxpceow1_0),.dout(w_dff_B_ir71D0UF7_0),.clk(gclk));
	jdff dff_B_6iJ4ZQlC5_0(.din(w_dff_B_ir71D0UF7_0),.dout(w_dff_B_6iJ4ZQlC5_0),.clk(gclk));
	jdff dff_B_R6auYvqy2_0(.din(w_dff_B_6iJ4ZQlC5_0),.dout(w_dff_B_R6auYvqy2_0),.clk(gclk));
	jdff dff_B_Nrh579qe2_0(.din(w_dff_B_R6auYvqy2_0),.dout(w_dff_B_Nrh579qe2_0),.clk(gclk));
	jdff dff_B_iVnIzRsb0_1(.din(n1512),.dout(w_dff_B_iVnIzRsb0_1),.clk(gclk));
	jdff dff_B_rUCszkdl1_0(.din(n1517),.dout(w_dff_B_rUCszkdl1_0),.clk(gclk));
	jdff dff_B_IKQhlY9y6_0(.din(w_dff_B_rUCszkdl1_0),.dout(w_dff_B_IKQhlY9y6_0),.clk(gclk));
	jdff dff_B_RGnY6viN6_0(.din(w_dff_B_IKQhlY9y6_0),.dout(w_dff_B_RGnY6viN6_0),.clk(gclk));
	jdff dff_B_sJYrScQ83_0(.din(w_dff_B_RGnY6viN6_0),.dout(w_dff_B_sJYrScQ83_0),.clk(gclk));
	jdff dff_B_YpX15TpO5_0(.din(w_dff_B_sJYrScQ83_0),.dout(w_dff_B_YpX15TpO5_0),.clk(gclk));
	jdff dff_B_1MTnPnjM5_0(.din(w_dff_B_YpX15TpO5_0),.dout(w_dff_B_1MTnPnjM5_0),.clk(gclk));
	jdff dff_B_9wr4v2i46_0(.din(w_dff_B_1MTnPnjM5_0),.dout(w_dff_B_9wr4v2i46_0),.clk(gclk));
	jdff dff_B_7M0PEGo79_0(.din(w_dff_B_9wr4v2i46_0),.dout(w_dff_B_7M0PEGo79_0),.clk(gclk));
	jdff dff_B_myCTkUXi8_0(.din(w_dff_B_7M0PEGo79_0),.dout(w_dff_B_myCTkUXi8_0),.clk(gclk));
	jdff dff_A_QNIvOtTH5_2(.dout(w_n366_0[2]),.din(w_dff_A_QNIvOtTH5_2),.clk(gclk));
	jdff dff_A_4pDBzIkj8_0(.dout(w_n361_0[0]),.din(w_dff_A_4pDBzIkj8_0),.clk(gclk));
	jdff dff_A_AoXjLKEa2_0(.dout(w_G38_2[0]),.din(w_dff_A_AoXjLKEa2_0),.clk(gclk));
	jdff dff_A_0RqgLhFE7_0(.dout(w_dff_A_AoXjLKEa2_0),.din(w_dff_A_0RqgLhFE7_0),.clk(gclk));
	jdff dff_A_AV8fO8in9_1(.dout(w_G38_2[1]),.din(w_dff_A_AV8fO8in9_1),.clk(gclk));
	jdff dff_A_GEC2RqG04_0(.dout(w_n1511_0[0]),.din(w_dff_A_GEC2RqG04_0),.clk(gclk));
	jdff dff_B_k6xiZitH3_2(.din(n1511),.dout(w_dff_B_k6xiZitH3_2),.clk(gclk));
	jdff dff_B_h91Oegy59_2(.din(w_dff_B_k6xiZitH3_2),.dout(w_dff_B_h91Oegy59_2),.clk(gclk));
	jdff dff_B_ceZN13d44_2(.din(w_dff_B_h91Oegy59_2),.dout(w_dff_B_ceZN13d44_2),.clk(gclk));
	jdff dff_B_gItFd5wj3_2(.din(w_dff_B_ceZN13d44_2),.dout(w_dff_B_gItFd5wj3_2),.clk(gclk));
	jdff dff_B_UaCCBgEI4_2(.din(w_dff_B_gItFd5wj3_2),.dout(w_dff_B_UaCCBgEI4_2),.clk(gclk));
	jdff dff_B_6cX0yVnW7_2(.din(w_dff_B_UaCCBgEI4_2),.dout(w_dff_B_6cX0yVnW7_2),.clk(gclk));
	jdff dff_B_yeZl5t8Z9_2(.din(w_dff_B_6cX0yVnW7_2),.dout(w_dff_B_yeZl5t8Z9_2),.clk(gclk));
	jdff dff_B_n59tdYKQ9_2(.din(w_dff_B_yeZl5t8Z9_2),.dout(w_dff_B_n59tdYKQ9_2),.clk(gclk));
	jdff dff_B_GB5UhtBF0_1(.din(n1508),.dout(w_dff_B_GB5UhtBF0_1),.clk(gclk));
	jdff dff_A_JsrNYtsM8_0(.dout(w_n364_0[0]),.din(w_dff_A_JsrNYtsM8_0),.clk(gclk));
	jdff dff_A_XrVfKjOm6_0(.dout(w_dff_A_JsrNYtsM8_0),.din(w_dff_A_XrVfKjOm6_0),.clk(gclk));
	jdff dff_A_HXEhRKtJ6_2(.dout(w_G1496_0[2]),.din(w_dff_A_HXEhRKtJ6_2),.clk(gclk));
	jdff dff_A_TygEWVQm6_2(.dout(w_dff_A_HXEhRKtJ6_2),.din(w_dff_A_TygEWVQm6_2),.clk(gclk));
	jdff dff_A_om8WZW3x7_2(.dout(w_dff_A_TygEWVQm6_2),.din(w_dff_A_om8WZW3x7_2),.clk(gclk));
	jdff dff_A_jj8FWGRv1_0(.dout(w_G1492_1[0]),.din(w_dff_A_jj8FWGRv1_0),.clk(gclk));
	jdff dff_A_5EyIJLb49_2(.dout(w_G1492_0[2]),.din(w_dff_A_5EyIJLb49_2),.clk(gclk));
	jdff dff_A_z84Sivjb7_2(.dout(w_dff_A_5EyIJLb49_2),.din(w_dff_A_z84Sivjb7_2),.clk(gclk));
	jdff dff_A_0Ti9dv7b3_2(.dout(w_dff_A_z84Sivjb7_2),.din(w_dff_A_0Ti9dv7b3_2),.clk(gclk));
	jdff dff_A_FQOPaHzv0_0(.dout(w_G38_0[0]),.din(w_dff_A_FQOPaHzv0_0),.clk(gclk));
	jdff dff_A_sWXvFQX26_2(.dout(w_G38_0[2]),.din(w_dff_A_sWXvFQX26_2),.clk(gclk));
	jdff dff_B_kXl7AKD53_1(.din(n376),.dout(w_dff_B_kXl7AKD53_1),.clk(gclk));
	jdff dff_B_gXPd4Jwn9_1(.din(w_dff_B_kXl7AKD53_1),.dout(w_dff_B_gXPd4Jwn9_1),.clk(gclk));
	jdff dff_B_skhcZKns8_1(.din(w_dff_B_gXPd4Jwn9_1),.dout(w_dff_B_skhcZKns8_1),.clk(gclk));
	jdff dff_B_3MxGaw4F7_1(.din(w_dff_B_skhcZKns8_1),.dout(w_dff_B_3MxGaw4F7_1),.clk(gclk));
	jdff dff_B_1leuiOL64_1(.din(w_dff_B_3MxGaw4F7_1),.dout(w_dff_B_1leuiOL64_1),.clk(gclk));
	jdff dff_B_6za001C86_1(.din(w_dff_B_1leuiOL64_1),.dout(w_dff_B_6za001C86_1),.clk(gclk));
	jdff dff_B_1VpL3ITN8_1(.din(w_dff_B_6za001C86_1),.dout(w_dff_B_1VpL3ITN8_1),.clk(gclk));
	jdff dff_B_GP6CBlmT3_1(.din(w_dff_B_1VpL3ITN8_1),.dout(w_dff_B_GP6CBlmT3_1),.clk(gclk));
	jdff dff_A_2scM1JL69_0(.dout(w_n377_1[0]),.din(w_dff_A_2scM1JL69_0),.clk(gclk));
	jdff dff_A_HT7AMlND8_0(.dout(w_dff_A_2scM1JL69_0),.din(w_dff_A_HT7AMlND8_0),.clk(gclk));
	jdff dff_A_3ny3aAEH1_0(.dout(w_dff_A_HT7AMlND8_0),.din(w_dff_A_3ny3aAEH1_0),.clk(gclk));
	jdff dff_A_Wp3jAbI40_0(.dout(w_dff_A_3ny3aAEH1_0),.din(w_dff_A_Wp3jAbI40_0),.clk(gclk));
	jdff dff_A_5spAxOzI6_0(.dout(w_dff_A_Wp3jAbI40_0),.din(w_dff_A_5spAxOzI6_0),.clk(gclk));
	jdff dff_A_19uBMY4k7_0(.dout(w_dff_A_5spAxOzI6_0),.din(w_dff_A_19uBMY4k7_0),.clk(gclk));
	jdff dff_A_7ylir7V19_0(.dout(w_dff_A_19uBMY4k7_0),.din(w_dff_A_7ylir7V19_0),.clk(gclk));
	jdff dff_A_clLEDIGw9_0(.dout(w_dff_A_7ylir7V19_0),.din(w_dff_A_clLEDIGw9_0),.clk(gclk));
	jdff dff_A_ePeB584u3_0(.dout(w_dff_A_clLEDIGw9_0),.din(w_dff_A_ePeB584u3_0),.clk(gclk));
	jdff dff_A_CT1Zwr7E6_0(.dout(w_dff_A_ePeB584u3_0),.din(w_dff_A_CT1Zwr7E6_0),.clk(gclk));
	jdff dff_A_NA3emlrz5_0(.dout(w_dff_A_CT1Zwr7E6_0),.din(w_dff_A_NA3emlrz5_0),.clk(gclk));
	jdff dff_A_1tUvtlUT3_0(.dout(w_dff_A_NA3emlrz5_0),.din(w_dff_A_1tUvtlUT3_0),.clk(gclk));
	jdff dff_A_7EcG6Nh41_0(.dout(w_dff_A_1tUvtlUT3_0),.din(w_dff_A_7EcG6Nh41_0),.clk(gclk));
	jdff dff_A_4n9Cq2BZ1_0(.dout(w_dff_A_7EcG6Nh41_0),.din(w_dff_A_4n9Cq2BZ1_0),.clk(gclk));
	jdff dff_A_xbcpzsOe3_0(.dout(w_dff_A_4n9Cq2BZ1_0),.din(w_dff_A_xbcpzsOe3_0),.clk(gclk));
	jdff dff_A_pWnRGosz6_0(.dout(w_dff_A_xbcpzsOe3_0),.din(w_dff_A_pWnRGosz6_0),.clk(gclk));
	jdff dff_A_Nfs8BZD57_0(.dout(w_dff_A_pWnRGosz6_0),.din(w_dff_A_Nfs8BZD57_0),.clk(gclk));
	jdff dff_A_fVC9dVDB5_0(.dout(w_dff_A_Nfs8BZD57_0),.din(w_dff_A_fVC9dVDB5_0),.clk(gclk));
	jdff dff_A_9jIclCX84_0(.dout(w_dff_A_fVC9dVDB5_0),.din(w_dff_A_9jIclCX84_0),.clk(gclk));
	jdff dff_A_G9eBYFVB8_0(.dout(w_dff_A_9jIclCX84_0),.din(w_dff_A_G9eBYFVB8_0),.clk(gclk));
	jdff dff_A_73VINfOf7_0(.dout(w_dff_A_G9eBYFVB8_0),.din(w_dff_A_73VINfOf7_0),.clk(gclk));
	jdff dff_A_q4Rcgtd79_0(.dout(w_dff_A_73VINfOf7_0),.din(w_dff_A_q4Rcgtd79_0),.clk(gclk));
	jdff dff_A_VuJDRYHz4_0(.dout(w_dff_A_q4Rcgtd79_0),.din(w_dff_A_VuJDRYHz4_0),.clk(gclk));
	jdff dff_A_PFxXQQEF3_0(.dout(w_dff_A_VuJDRYHz4_0),.din(w_dff_A_PFxXQQEF3_0),.clk(gclk));
	jdff dff_A_biG1YBpe4_0(.dout(w_dff_A_PFxXQQEF3_0),.din(w_dff_A_biG1YBpe4_0),.clk(gclk));
	jdff dff_A_UOo25iMB9_0(.dout(w_dff_A_biG1YBpe4_0),.din(w_dff_A_UOo25iMB9_0),.clk(gclk));
	jdff dff_A_2DWOwWGn1_0(.dout(w_dff_A_UOo25iMB9_0),.din(w_dff_A_2DWOwWGn1_0),.clk(gclk));
	jdff dff_A_otJcy7zp3_0(.dout(w_dff_A_2DWOwWGn1_0),.din(w_dff_A_otJcy7zp3_0),.clk(gclk));
	jdff dff_A_P3Kbsd9q8_0(.dout(w_dff_A_otJcy7zp3_0),.din(w_dff_A_P3Kbsd9q8_0),.clk(gclk));
	jdff dff_A_9QatQ9tk9_0(.dout(w_dff_A_P3Kbsd9q8_0),.din(w_dff_A_9QatQ9tk9_0),.clk(gclk));
	jdff dff_A_SiChp53D2_2(.dout(w_n377_1[2]),.din(w_dff_A_SiChp53D2_2),.clk(gclk));
	jdff dff_A_OpQKdVDa4_2(.dout(w_dff_A_SiChp53D2_2),.din(w_dff_A_OpQKdVDa4_2),.clk(gclk));
	jdff dff_A_CsClAuT21_2(.dout(w_dff_A_OpQKdVDa4_2),.din(w_dff_A_CsClAuT21_2),.clk(gclk));
	jdff dff_A_iNggLAeh1_2(.dout(w_dff_A_CsClAuT21_2),.din(w_dff_A_iNggLAeh1_2),.clk(gclk));
	jdff dff_A_khjwgLvX2_2(.dout(w_dff_A_iNggLAeh1_2),.din(w_dff_A_khjwgLvX2_2),.clk(gclk));
	jdff dff_B_4URZCTKT2_1(.din(n1480),.dout(w_dff_B_4URZCTKT2_1),.clk(gclk));
	jdff dff_B_IIRAvDTi4_1(.din(w_dff_B_4URZCTKT2_1),.dout(w_dff_B_IIRAvDTi4_1),.clk(gclk));
	jdff dff_B_H9669h9Z1_1(.din(w_dff_B_IIRAvDTi4_1),.dout(w_dff_B_H9669h9Z1_1),.clk(gclk));
	jdff dff_B_XCrdcWAr7_1(.din(w_dff_B_H9669h9Z1_1),.dout(w_dff_B_XCrdcWAr7_1),.clk(gclk));
	jdff dff_B_MScwB68L7_1(.din(w_dff_B_XCrdcWAr7_1),.dout(w_dff_B_MScwB68L7_1),.clk(gclk));
	jdff dff_B_n5I8J8zb3_1(.din(w_dff_B_MScwB68L7_1),.dout(w_dff_B_n5I8J8zb3_1),.clk(gclk));
	jdff dff_B_VecfdJva2_1(.din(w_dff_B_n5I8J8zb3_1),.dout(w_dff_B_VecfdJva2_1),.clk(gclk));
	jdff dff_B_lmdSCRQa8_1(.din(w_dff_B_VecfdJva2_1),.dout(w_dff_B_lmdSCRQa8_1),.clk(gclk));
	jdff dff_B_dQLeCAFX5_1(.din(w_dff_B_lmdSCRQa8_1),.dout(w_dff_B_dQLeCAFX5_1),.clk(gclk));
	jdff dff_B_52g9Ls848_1(.din(w_dff_B_dQLeCAFX5_1),.dout(w_dff_B_52g9Ls848_1),.clk(gclk));
	jdff dff_B_NATieFFa3_1(.din(w_dff_B_52g9Ls848_1),.dout(w_dff_B_NATieFFa3_1),.clk(gclk));
	jdff dff_B_2ZjSOoZk1_1(.din(w_dff_B_NATieFFa3_1),.dout(w_dff_B_2ZjSOoZk1_1),.clk(gclk));
	jdff dff_B_K565x8eR5_1(.din(w_dff_B_2ZjSOoZk1_1),.dout(w_dff_B_K565x8eR5_1),.clk(gclk));
	jdff dff_B_jJYMotSy6_1(.din(w_dff_B_K565x8eR5_1),.dout(w_dff_B_jJYMotSy6_1),.clk(gclk));
	jdff dff_B_DPT6iVDN3_1(.din(w_dff_B_jJYMotSy6_1),.dout(w_dff_B_DPT6iVDN3_1),.clk(gclk));
	jdff dff_B_2Rq562tP6_1(.din(w_dff_B_DPT6iVDN3_1),.dout(w_dff_B_2Rq562tP6_1),.clk(gclk));
	jdff dff_B_v5OaJ4Ow5_1(.din(w_dff_B_2Rq562tP6_1),.dout(w_dff_B_v5OaJ4Ow5_1),.clk(gclk));
	jdff dff_B_1eXPyZuP0_1(.din(w_dff_B_v5OaJ4Ow5_1),.dout(w_dff_B_1eXPyZuP0_1),.clk(gclk));
	jdff dff_B_2yN8lW562_1(.din(w_dff_B_1eXPyZuP0_1),.dout(w_dff_B_2yN8lW562_1),.clk(gclk));
	jdff dff_B_4bfEc6Q59_1(.din(w_dff_B_2yN8lW562_1),.dout(w_dff_B_4bfEc6Q59_1),.clk(gclk));
	jdff dff_B_iKOJSfaE1_1(.din(w_dff_B_4bfEc6Q59_1),.dout(w_dff_B_iKOJSfaE1_1),.clk(gclk));
	jdff dff_B_OBsVua4Z4_1(.din(w_dff_B_iKOJSfaE1_1),.dout(w_dff_B_OBsVua4Z4_1),.clk(gclk));
	jdff dff_B_dUJDzBcM6_1(.din(w_dff_B_OBsVua4Z4_1),.dout(w_dff_B_dUJDzBcM6_1),.clk(gclk));
	jdff dff_B_YoHRC7kQ1_1(.din(w_dff_B_dUJDzBcM6_1),.dout(w_dff_B_YoHRC7kQ1_1),.clk(gclk));
	jdff dff_B_KUJFyn363_1(.din(w_dff_B_YoHRC7kQ1_1),.dout(w_dff_B_KUJFyn363_1),.clk(gclk));
	jdff dff_B_a0A0R9iS4_1(.din(w_dff_B_KUJFyn363_1),.dout(w_dff_B_a0A0R9iS4_1),.clk(gclk));
	jdff dff_B_iBqu3Y7d7_1(.din(w_dff_B_a0A0R9iS4_1),.dout(w_dff_B_iBqu3Y7d7_1),.clk(gclk));
	jdff dff_B_57n7TXKg3_1(.din(w_dff_B_iBqu3Y7d7_1),.dout(w_dff_B_57n7TXKg3_1),.clk(gclk));
	jdff dff_B_EzkNbk9Z3_1(.din(w_dff_B_57n7TXKg3_1),.dout(w_dff_B_EzkNbk9Z3_1),.clk(gclk));
	jdff dff_B_YaANBgLp9_1(.din(w_dff_B_EzkNbk9Z3_1),.dout(w_dff_B_YaANBgLp9_1),.clk(gclk));
	jdff dff_B_QwCIe8H74_1(.din(w_dff_B_YaANBgLp9_1),.dout(w_dff_B_QwCIe8H74_1),.clk(gclk));
	jdff dff_B_zAPGi7sQ9_0(.din(n1502),.dout(w_dff_B_zAPGi7sQ9_0),.clk(gclk));
	jdff dff_B_kpcEDEf08_0(.din(w_dff_B_zAPGi7sQ9_0),.dout(w_dff_B_kpcEDEf08_0),.clk(gclk));
	jdff dff_B_cxTFnbYF4_0(.din(w_dff_B_kpcEDEf08_0),.dout(w_dff_B_cxTFnbYF4_0),.clk(gclk));
	jdff dff_B_uPPHhfSG4_0(.din(w_dff_B_cxTFnbYF4_0),.dout(w_dff_B_uPPHhfSG4_0),.clk(gclk));
	jdff dff_B_XK8ll53l8_0(.din(w_dff_B_uPPHhfSG4_0),.dout(w_dff_B_XK8ll53l8_0),.clk(gclk));
	jdff dff_B_azRK4Jwg0_0(.din(w_dff_B_XK8ll53l8_0),.dout(w_dff_B_azRK4Jwg0_0),.clk(gclk));
	jdff dff_B_QVinhlI20_0(.din(w_dff_B_azRK4Jwg0_0),.dout(w_dff_B_QVinhlI20_0),.clk(gclk));
	jdff dff_B_rawBPdkp5_0(.din(w_dff_B_QVinhlI20_0),.dout(w_dff_B_rawBPdkp5_0),.clk(gclk));
	jdff dff_B_fexPNuMS8_0(.din(w_dff_B_rawBPdkp5_0),.dout(w_dff_B_fexPNuMS8_0),.clk(gclk));
	jdff dff_B_MaMLRemh2_0(.din(w_dff_B_fexPNuMS8_0),.dout(w_dff_B_MaMLRemh2_0),.clk(gclk));
	jdff dff_B_A901igYJ6_0(.din(w_dff_B_MaMLRemh2_0),.dout(w_dff_B_A901igYJ6_0),.clk(gclk));
	jdff dff_B_dxs6qdP81_0(.din(w_dff_B_A901igYJ6_0),.dout(w_dff_B_dxs6qdP81_0),.clk(gclk));
	jdff dff_B_LVMcigG42_0(.din(w_dff_B_dxs6qdP81_0),.dout(w_dff_B_LVMcigG42_0),.clk(gclk));
	jdff dff_B_EOpICpsq9_0(.din(w_dff_B_LVMcigG42_0),.dout(w_dff_B_EOpICpsq9_0),.clk(gclk));
	jdff dff_B_sA3whaAc2_0(.din(w_dff_B_EOpICpsq9_0),.dout(w_dff_B_sA3whaAc2_0),.clk(gclk));
	jdff dff_B_gvLAsJf49_0(.din(w_dff_B_sA3whaAc2_0),.dout(w_dff_B_gvLAsJf49_0),.clk(gclk));
	jdff dff_B_vfS4H3GJ8_0(.din(w_dff_B_gvLAsJf49_0),.dout(w_dff_B_vfS4H3GJ8_0),.clk(gclk));
	jdff dff_B_IU8FPb0D3_0(.din(w_dff_B_vfS4H3GJ8_0),.dout(w_dff_B_IU8FPb0D3_0),.clk(gclk));
	jdff dff_B_3IfdK66J1_0(.din(w_dff_B_IU8FPb0D3_0),.dout(w_dff_B_3IfdK66J1_0),.clk(gclk));
	jdff dff_B_AHUCtzZZ4_0(.din(w_dff_B_3IfdK66J1_0),.dout(w_dff_B_AHUCtzZZ4_0),.clk(gclk));
	jdff dff_B_VG3jWbMU3_1(.din(n1497),.dout(w_dff_B_VG3jWbMU3_1),.clk(gclk));
	jdff dff_B_Wz9LiyGS3_1(.din(w_dff_B_VG3jWbMU3_1),.dout(w_dff_B_Wz9LiyGS3_1),.clk(gclk));
	jdff dff_B_xStXXyDX5_0(.din(n1498),.dout(w_dff_B_xStXXyDX5_0),.clk(gclk));
	jdff dff_B_8C6OP5B58_0(.din(w_dff_B_xStXXyDX5_0),.dout(w_dff_B_8C6OP5B58_0),.clk(gclk));
	jdff dff_B_EkJW2d739_0(.din(w_dff_B_8C6OP5B58_0),.dout(w_dff_B_EkJW2d739_0),.clk(gclk));
	jdff dff_B_GfHZKRgn0_0(.din(w_dff_B_EkJW2d739_0),.dout(w_dff_B_GfHZKRgn0_0),.clk(gclk));
	jdff dff_B_7TJ07BqD6_0(.din(w_dff_B_GfHZKRgn0_0),.dout(w_dff_B_7TJ07BqD6_0),.clk(gclk));
	jdff dff_A_FGO3VwDe7_1(.dout(w_n1364_0[1]),.din(w_dff_A_FGO3VwDe7_1),.clk(gclk));
	jdff dff_A_4GxBDFuK5_1(.dout(w_dff_A_FGO3VwDe7_1),.din(w_dff_A_4GxBDFuK5_1),.clk(gclk));
	jdff dff_A_9Dandry36_1(.dout(w_dff_A_4GxBDFuK5_1),.din(w_dff_A_9Dandry36_1),.clk(gclk));
	jdff dff_A_WsZgq4ld1_1(.dout(w_dff_A_9Dandry36_1),.din(w_dff_A_WsZgq4ld1_1),.clk(gclk));
	jdff dff_A_62agWQZ76_1(.dout(w_dff_A_WsZgq4ld1_1),.din(w_dff_A_62agWQZ76_1),.clk(gclk));
	jdff dff_A_AquFdCbi3_1(.dout(w_dff_A_62agWQZ76_1),.din(w_dff_A_AquFdCbi3_1),.clk(gclk));
	jdff dff_A_FE4fiykW8_1(.dout(w_dff_A_AquFdCbi3_1),.din(w_dff_A_FE4fiykW8_1),.clk(gclk));
	jdff dff_A_pOPNpuih6_1(.dout(w_dff_A_FE4fiykW8_1),.din(w_dff_A_pOPNpuih6_1),.clk(gclk));
	jdff dff_A_A4OjkDoC9_1(.dout(w_dff_A_pOPNpuih6_1),.din(w_dff_A_A4OjkDoC9_1),.clk(gclk));
	jdff dff_A_96IQSY3P0_1(.dout(w_dff_A_A4OjkDoC9_1),.din(w_dff_A_96IQSY3P0_1),.clk(gclk));
	jdff dff_A_rcEpXCLT9_1(.dout(w_dff_A_96IQSY3P0_1),.din(w_dff_A_rcEpXCLT9_1),.clk(gclk));
	jdff dff_A_FueC69Vb4_1(.dout(w_dff_A_rcEpXCLT9_1),.din(w_dff_A_FueC69Vb4_1),.clk(gclk));
	jdff dff_A_VZSUXcJR1_1(.dout(w_dff_A_FueC69Vb4_1),.din(w_dff_A_VZSUXcJR1_1),.clk(gclk));
	jdff dff_A_XdQMZGYT8_1(.dout(w_dff_A_VZSUXcJR1_1),.din(w_dff_A_XdQMZGYT8_1),.clk(gclk));
	jdff dff_A_KKXS9DGc4_1(.dout(w_dff_A_XdQMZGYT8_1),.din(w_dff_A_KKXS9DGc4_1),.clk(gclk));
	jdff dff_A_iEOT29u52_1(.dout(w_dff_A_KKXS9DGc4_1),.din(w_dff_A_iEOT29u52_1),.clk(gclk));
	jdff dff_A_xhJreGxM4_1(.dout(w_dff_A_iEOT29u52_1),.din(w_dff_A_xhJreGxM4_1),.clk(gclk));
	jdff dff_A_5rZqYOZF2_1(.dout(w_dff_A_xhJreGxM4_1),.din(w_dff_A_5rZqYOZF2_1),.clk(gclk));
	jdff dff_A_JMGaejtI5_1(.dout(w_dff_A_5rZqYOZF2_1),.din(w_dff_A_JMGaejtI5_1),.clk(gclk));
	jdff dff_A_6kHtavVd7_1(.dout(w_dff_A_JMGaejtI5_1),.din(w_dff_A_6kHtavVd7_1),.clk(gclk));
	jdff dff_A_BtTuPcIS1_1(.dout(w_dff_A_6kHtavVd7_1),.din(w_dff_A_BtTuPcIS1_1),.clk(gclk));
	jdff dff_A_VTtE4p5y2_1(.dout(w_dff_A_BtTuPcIS1_1),.din(w_dff_A_VTtE4p5y2_1),.clk(gclk));
	jdff dff_A_aMUHQ7Iu9_1(.dout(w_dff_A_VTtE4p5y2_1),.din(w_dff_A_aMUHQ7Iu9_1),.clk(gclk));
	jdff dff_A_G14UZ7Ts8_1(.dout(w_dff_A_aMUHQ7Iu9_1),.din(w_dff_A_G14UZ7Ts8_1),.clk(gclk));
	jdff dff_A_xuCJl1nq8_1(.dout(w_dff_A_G14UZ7Ts8_1),.din(w_dff_A_xuCJl1nq8_1),.clk(gclk));
	jdff dff_B_6dr2HROu8_0(.din(n1363),.dout(w_dff_B_6dr2HROu8_0),.clk(gclk));
	jdff dff_B_CJN2F4J86_0(.din(w_dff_B_6dr2HROu8_0),.dout(w_dff_B_CJN2F4J86_0),.clk(gclk));
	jdff dff_B_6Xm9GNkp1_0(.din(w_dff_B_CJN2F4J86_0),.dout(w_dff_B_6Xm9GNkp1_0),.clk(gclk));
	jdff dff_B_jvy3VoAt6_1(.din(n1494),.dout(w_dff_B_jvy3VoAt6_1),.clk(gclk));
	jdff dff_B_iTP5sQCM5_1(.din(w_dff_B_jvy3VoAt6_1),.dout(w_dff_B_iTP5sQCM5_1),.clk(gclk));
	jdff dff_B_SFXMS2uJ4_1(.din(w_dff_B_iTP5sQCM5_1),.dout(w_dff_B_SFXMS2uJ4_1),.clk(gclk));
	jdff dff_B_qVejruuc3_1(.din(n1495),.dout(w_dff_B_qVejruuc3_1),.clk(gclk));
	jdff dff_B_zpFoqYh97_1(.din(w_dff_B_qVejruuc3_1),.dout(w_dff_B_zpFoqYh97_1),.clk(gclk));
	jdff dff_A_qQNwmH5o6_1(.dout(w_n1359_0[1]),.din(w_dff_A_qQNwmH5o6_1),.clk(gclk));
	jdff dff_A_nVFKisTE2_1(.dout(w_dff_A_qQNwmH5o6_1),.din(w_dff_A_nVFKisTE2_1),.clk(gclk));
	jdff dff_A_ktLMMZcL7_1(.dout(w_dff_A_nVFKisTE2_1),.din(w_dff_A_ktLMMZcL7_1),.clk(gclk));
	jdff dff_A_SLotKsRL8_1(.dout(w_dff_A_ktLMMZcL7_1),.din(w_dff_A_SLotKsRL8_1),.clk(gclk));
	jdff dff_A_EzpjlKyO6_1(.dout(w_dff_A_SLotKsRL8_1),.din(w_dff_A_EzpjlKyO6_1),.clk(gclk));
	jdff dff_A_HfGWA7UL9_1(.dout(w_dff_A_EzpjlKyO6_1),.din(w_dff_A_HfGWA7UL9_1),.clk(gclk));
	jdff dff_A_hKV06LHL6_1(.dout(w_dff_A_HfGWA7UL9_1),.din(w_dff_A_hKV06LHL6_1),.clk(gclk));
	jdff dff_A_7nE0DL139_1(.dout(w_dff_A_hKV06LHL6_1),.din(w_dff_A_7nE0DL139_1),.clk(gclk));
	jdff dff_A_YmS8dCMC5_1(.dout(w_dff_A_7nE0DL139_1),.din(w_dff_A_YmS8dCMC5_1),.clk(gclk));
	jdff dff_A_UbIBYy1D3_1(.dout(w_dff_A_YmS8dCMC5_1),.din(w_dff_A_UbIBYy1D3_1),.clk(gclk));
	jdff dff_A_k0dx8DWQ3_1(.dout(w_dff_A_UbIBYy1D3_1),.din(w_dff_A_k0dx8DWQ3_1),.clk(gclk));
	jdff dff_A_0m2DTqYc6_1(.dout(w_dff_A_k0dx8DWQ3_1),.din(w_dff_A_0m2DTqYc6_1),.clk(gclk));
	jdff dff_A_TCvrdDZE9_1(.dout(w_dff_A_0m2DTqYc6_1),.din(w_dff_A_TCvrdDZE9_1),.clk(gclk));
	jdff dff_A_7Ayixigf7_1(.dout(w_dff_A_TCvrdDZE9_1),.din(w_dff_A_7Ayixigf7_1),.clk(gclk));
	jdff dff_A_Iq0hghM34_1(.dout(w_dff_A_7Ayixigf7_1),.din(w_dff_A_Iq0hghM34_1),.clk(gclk));
	jdff dff_A_nYKAr1b15_1(.dout(w_dff_A_Iq0hghM34_1),.din(w_dff_A_nYKAr1b15_1),.clk(gclk));
	jdff dff_A_ARd6ITmS7_1(.dout(w_dff_A_nYKAr1b15_1),.din(w_dff_A_ARd6ITmS7_1),.clk(gclk));
	jdff dff_A_GXlCHxSq3_1(.dout(w_dff_A_ARd6ITmS7_1),.din(w_dff_A_GXlCHxSq3_1),.clk(gclk));
	jdff dff_A_1i44VYq57_1(.dout(w_dff_A_GXlCHxSq3_1),.din(w_dff_A_1i44VYq57_1),.clk(gclk));
	jdff dff_A_xdS4xNOl2_1(.dout(w_dff_A_1i44VYq57_1),.din(w_dff_A_xdS4xNOl2_1),.clk(gclk));
	jdff dff_A_6GealkN51_1(.dout(w_dff_A_xdS4xNOl2_1),.din(w_dff_A_6GealkN51_1),.clk(gclk));
	jdff dff_A_OQiWABd12_1(.dout(w_dff_A_6GealkN51_1),.din(w_dff_A_OQiWABd12_1),.clk(gclk));
	jdff dff_B_H8oXmmA94_2(.din(n1359),.dout(w_dff_B_H8oXmmA94_2),.clk(gclk));
	jdff dff_A_nfikk4AQ6_0(.dout(w_n418_0[0]),.din(w_dff_A_nfikk4AQ6_0),.clk(gclk));
	jdff dff_A_lkcE2c0P4_0(.dout(w_dff_A_nfikk4AQ6_0),.din(w_dff_A_lkcE2c0P4_0),.clk(gclk));
	jdff dff_A_qxMPcfHI4_0(.dout(w_dff_A_lkcE2c0P4_0),.din(w_dff_A_qxMPcfHI4_0),.clk(gclk));
	jdff dff_A_h4etcT9V1_0(.dout(w_dff_A_qxMPcfHI4_0),.din(w_dff_A_h4etcT9V1_0),.clk(gclk));
	jdff dff_A_iWAGMO7h6_0(.dout(w_dff_A_h4etcT9V1_0),.din(w_dff_A_iWAGMO7h6_0),.clk(gclk));
	jdff dff_B_bFGdTcFl7_1(.din(n1324),.dout(w_dff_B_bFGdTcFl7_1),.clk(gclk));
	jdff dff_B_uktRUa4U6_1(.din(w_dff_B_bFGdTcFl7_1),.dout(w_dff_B_uktRUa4U6_1),.clk(gclk));
	jdff dff_B_yPB3bYIt8_1(.din(w_dff_B_uktRUa4U6_1),.dout(w_dff_B_yPB3bYIt8_1),.clk(gclk));
	jdff dff_B_SnoR0ISc2_1(.din(w_dff_B_yPB3bYIt8_1),.dout(w_dff_B_SnoR0ISc2_1),.clk(gclk));
	jdff dff_B_a6kOW1KS8_1(.din(w_dff_B_SnoR0ISc2_1),.dout(w_dff_B_a6kOW1KS8_1),.clk(gclk));
	jdff dff_B_mZtiIKQf2_1(.din(w_dff_B_a6kOW1KS8_1),.dout(w_dff_B_mZtiIKQf2_1),.clk(gclk));
	jdff dff_B_pZ9D4wAW0_1(.din(w_dff_B_mZtiIKQf2_1),.dout(w_dff_B_pZ9D4wAW0_1),.clk(gclk));
	jdff dff_B_GclWk9i40_1(.din(w_dff_B_pZ9D4wAW0_1),.dout(w_dff_B_GclWk9i40_1),.clk(gclk));
	jdff dff_B_NEiHFAHC2_1(.din(w_dff_B_GclWk9i40_1),.dout(w_dff_B_NEiHFAHC2_1),.clk(gclk));
	jdff dff_B_aR29EeWm8_1(.din(w_dff_B_NEiHFAHC2_1),.dout(w_dff_B_aR29EeWm8_1),.clk(gclk));
	jdff dff_B_URtq9owT4_1(.din(w_dff_B_aR29EeWm8_1),.dout(w_dff_B_URtq9owT4_1),.clk(gclk));
	jdff dff_B_4g3291wX8_1(.din(w_dff_B_URtq9owT4_1),.dout(w_dff_B_4g3291wX8_1),.clk(gclk));
	jdff dff_B_X2fhvDj11_1(.din(w_dff_B_4g3291wX8_1),.dout(w_dff_B_X2fhvDj11_1),.clk(gclk));
	jdff dff_B_JJ2mHynC8_1(.din(w_dff_B_X2fhvDj11_1),.dout(w_dff_B_JJ2mHynC8_1),.clk(gclk));
	jdff dff_B_gUZoFocb4_1(.din(w_dff_B_JJ2mHynC8_1),.dout(w_dff_B_gUZoFocb4_1),.clk(gclk));
	jdff dff_B_GFxji9EJ8_1(.din(w_dff_B_gUZoFocb4_1),.dout(w_dff_B_GFxji9EJ8_1),.clk(gclk));
	jdff dff_B_HE4ZSF592_1(.din(w_dff_B_GFxji9EJ8_1),.dout(w_dff_B_HE4ZSF592_1),.clk(gclk));
	jdff dff_B_48tK7MUN0_1(.din(w_dff_B_HE4ZSF592_1),.dout(w_dff_B_48tK7MUN0_1),.clk(gclk));
	jdff dff_B_Su3kwOrT5_1(.din(w_dff_B_48tK7MUN0_1),.dout(w_dff_B_Su3kwOrT5_1),.clk(gclk));
	jdff dff_B_DkS7F9ki1_1(.din(w_dff_B_Su3kwOrT5_1),.dout(w_dff_B_DkS7F9ki1_1),.clk(gclk));
	jdff dff_B_OiLJXAWd0_1(.din(w_dff_B_DkS7F9ki1_1),.dout(w_dff_B_OiLJXAWd0_1),.clk(gclk));
	jdff dff_B_jet4qFZK3_1(.din(w_dff_B_OiLJXAWd0_1),.dout(w_dff_B_jet4qFZK3_1),.clk(gclk));
	jdff dff_B_0LPA7P8j1_1(.din(w_dff_B_jet4qFZK3_1),.dout(w_dff_B_0LPA7P8j1_1),.clk(gclk));
	jdff dff_B_lInV46iW7_1(.din(w_dff_B_0LPA7P8j1_1),.dout(w_dff_B_lInV46iW7_1),.clk(gclk));
	jdff dff_B_8xwmUzaQ2_1(.din(w_dff_B_lInV46iW7_1),.dout(w_dff_B_8xwmUzaQ2_1),.clk(gclk));
	jdff dff_B_sn5wKndL8_1(.din(w_dff_B_8xwmUzaQ2_1),.dout(w_dff_B_sn5wKndL8_1),.clk(gclk));
	jdff dff_B_k4OnJtg44_1(.din(w_dff_B_sn5wKndL8_1),.dout(w_dff_B_k4OnJtg44_1),.clk(gclk));
	jdff dff_B_zmbOQOvP3_1(.din(w_dff_B_k4OnJtg44_1),.dout(w_dff_B_zmbOQOvP3_1),.clk(gclk));
	jdff dff_B_U3fnmt7e9_1(.din(n1325),.dout(w_dff_B_U3fnmt7e9_1),.clk(gclk));
	jdff dff_B_PXcm5kGH7_1(.din(w_dff_B_U3fnmt7e9_1),.dout(w_dff_B_PXcm5kGH7_1),.clk(gclk));
	jdff dff_B_Du06je7b1_1(.din(w_dff_B_PXcm5kGH7_1),.dout(w_dff_B_Du06je7b1_1),.clk(gclk));
	jdff dff_B_4e5OsMwi1_1(.din(w_dff_B_Du06je7b1_1),.dout(w_dff_B_4e5OsMwi1_1),.clk(gclk));
	jdff dff_B_Nt7kok2D2_1(.din(w_dff_B_4e5OsMwi1_1),.dout(w_dff_B_Nt7kok2D2_1),.clk(gclk));
	jdff dff_B_LHcp6NtL3_1(.din(w_dff_B_Nt7kok2D2_1),.dout(w_dff_B_LHcp6NtL3_1),.clk(gclk));
	jdff dff_B_s0BKhxcC7_1(.din(w_dff_B_LHcp6NtL3_1),.dout(w_dff_B_s0BKhxcC7_1),.clk(gclk));
	jdff dff_B_uXUOpUnp0_1(.din(w_dff_B_s0BKhxcC7_1),.dout(w_dff_B_uXUOpUnp0_1),.clk(gclk));
	jdff dff_B_IuDRgzOw6_1(.din(w_dff_B_uXUOpUnp0_1),.dout(w_dff_B_IuDRgzOw6_1),.clk(gclk));
	jdff dff_B_iX6HCfrX8_1(.din(w_dff_B_IuDRgzOw6_1),.dout(w_dff_B_iX6HCfrX8_1),.clk(gclk));
	jdff dff_B_TkAQmy2F6_1(.din(w_dff_B_iX6HCfrX8_1),.dout(w_dff_B_TkAQmy2F6_1),.clk(gclk));
	jdff dff_B_HZP9cHmN3_1(.din(w_dff_B_TkAQmy2F6_1),.dout(w_dff_B_HZP9cHmN3_1),.clk(gclk));
	jdff dff_B_SErHn3Co3_1(.din(w_dff_B_HZP9cHmN3_1),.dout(w_dff_B_SErHn3Co3_1),.clk(gclk));
	jdff dff_B_a5KWdw619_1(.din(w_dff_B_SErHn3Co3_1),.dout(w_dff_B_a5KWdw619_1),.clk(gclk));
	jdff dff_B_6nfR4x0N9_1(.din(w_dff_B_a5KWdw619_1),.dout(w_dff_B_6nfR4x0N9_1),.clk(gclk));
	jdff dff_B_oqP1e4z64_1(.din(w_dff_B_6nfR4x0N9_1),.dout(w_dff_B_oqP1e4z64_1),.clk(gclk));
	jdff dff_B_HrBH1RxL0_1(.din(w_dff_B_oqP1e4z64_1),.dout(w_dff_B_HrBH1RxL0_1),.clk(gclk));
	jdff dff_B_yxSWqYma7_1(.din(w_dff_B_HrBH1RxL0_1),.dout(w_dff_B_yxSWqYma7_1),.clk(gclk));
	jdff dff_B_o8Emg5SK9_1(.din(w_dff_B_yxSWqYma7_1),.dout(w_dff_B_o8Emg5SK9_1),.clk(gclk));
	jdff dff_B_Rktz6AM47_1(.din(w_dff_B_o8Emg5SK9_1),.dout(w_dff_B_Rktz6AM47_1),.clk(gclk));
	jdff dff_B_0QIdrxkI4_1(.din(w_dff_B_Rktz6AM47_1),.dout(w_dff_B_0QIdrxkI4_1),.clk(gclk));
	jdff dff_B_Cf7HDrTi8_1(.din(w_dff_B_0QIdrxkI4_1),.dout(w_dff_B_Cf7HDrTi8_1),.clk(gclk));
	jdff dff_B_ZsIJhXav8_1(.din(w_dff_B_Cf7HDrTi8_1),.dout(w_dff_B_ZsIJhXav8_1),.clk(gclk));
	jdff dff_B_MpGPcPli1_1(.din(w_dff_B_ZsIJhXav8_1),.dout(w_dff_B_MpGPcPli1_1),.clk(gclk));
	jdff dff_B_QxqAoEww1_1(.din(w_dff_B_MpGPcPli1_1),.dout(w_dff_B_QxqAoEww1_1),.clk(gclk));
	jdff dff_B_usKxzaUL4_1(.din(w_dff_B_QxqAoEww1_1),.dout(w_dff_B_usKxzaUL4_1),.clk(gclk));
	jdff dff_B_vp9A2Y2X7_1(.din(w_dff_B_usKxzaUL4_1),.dout(w_dff_B_vp9A2Y2X7_1),.clk(gclk));
	jdff dff_B_cESwo7Oj0_1(.din(n1326),.dout(w_dff_B_cESwo7Oj0_1),.clk(gclk));
	jdff dff_B_R69Topu95_1(.din(w_dff_B_cESwo7Oj0_1),.dout(w_dff_B_R69Topu95_1),.clk(gclk));
	jdff dff_B_67skyuQZ3_1(.din(w_dff_B_R69Topu95_1),.dout(w_dff_B_67skyuQZ3_1),.clk(gclk));
	jdff dff_B_AxBhauOz4_1(.din(w_dff_B_67skyuQZ3_1),.dout(w_dff_B_AxBhauOz4_1),.clk(gclk));
	jdff dff_B_KEgrpVWj1_1(.din(w_dff_B_AxBhauOz4_1),.dout(w_dff_B_KEgrpVWj1_1),.clk(gclk));
	jdff dff_B_8zSm99nB1_1(.din(w_dff_B_KEgrpVWj1_1),.dout(w_dff_B_8zSm99nB1_1),.clk(gclk));
	jdff dff_B_gPFETUWy8_1(.din(w_dff_B_8zSm99nB1_1),.dout(w_dff_B_gPFETUWy8_1),.clk(gclk));
	jdff dff_B_BQXFmObV5_1(.din(w_dff_B_gPFETUWy8_1),.dout(w_dff_B_BQXFmObV5_1),.clk(gclk));
	jdff dff_B_pKtYLJ7Z5_1(.din(w_dff_B_BQXFmObV5_1),.dout(w_dff_B_pKtYLJ7Z5_1),.clk(gclk));
	jdff dff_B_wV0BdER56_1(.din(w_dff_B_pKtYLJ7Z5_1),.dout(w_dff_B_wV0BdER56_1),.clk(gclk));
	jdff dff_B_JPv22FWC9_1(.din(w_dff_B_wV0BdER56_1),.dout(w_dff_B_JPv22FWC9_1),.clk(gclk));
	jdff dff_B_XnJiykrU9_1(.din(w_dff_B_JPv22FWC9_1),.dout(w_dff_B_XnJiykrU9_1),.clk(gclk));
	jdff dff_B_FL6Sb9Lk6_1(.din(w_dff_B_XnJiykrU9_1),.dout(w_dff_B_FL6Sb9Lk6_1),.clk(gclk));
	jdff dff_B_T0wtvQYU4_1(.din(w_dff_B_FL6Sb9Lk6_1),.dout(w_dff_B_T0wtvQYU4_1),.clk(gclk));
	jdff dff_B_cCF5SyOg4_1(.din(w_dff_B_T0wtvQYU4_1),.dout(w_dff_B_cCF5SyOg4_1),.clk(gclk));
	jdff dff_B_KX9axuSC7_1(.din(w_dff_B_cCF5SyOg4_1),.dout(w_dff_B_KX9axuSC7_1),.clk(gclk));
	jdff dff_B_NOkpmACW8_1(.din(w_dff_B_KX9axuSC7_1),.dout(w_dff_B_NOkpmACW8_1),.clk(gclk));
	jdff dff_B_Jb6RIUga0_1(.din(w_dff_B_NOkpmACW8_1),.dout(w_dff_B_Jb6RIUga0_1),.clk(gclk));
	jdff dff_B_vdkrFCYN1_1(.din(w_dff_B_Jb6RIUga0_1),.dout(w_dff_B_vdkrFCYN1_1),.clk(gclk));
	jdff dff_B_ZsqlCYh01_1(.din(w_dff_B_vdkrFCYN1_1),.dout(w_dff_B_ZsqlCYh01_1),.clk(gclk));
	jdff dff_B_rnCe3Ork8_1(.din(w_dff_B_ZsqlCYh01_1),.dout(w_dff_B_rnCe3Ork8_1),.clk(gclk));
	jdff dff_B_k128GXOQ4_1(.din(n1327),.dout(w_dff_B_k128GXOQ4_1),.clk(gclk));
	jdff dff_B_8v1f5lu64_1(.din(w_dff_B_k128GXOQ4_1),.dout(w_dff_B_8v1f5lu64_1),.clk(gclk));
	jdff dff_B_qDMTBvTM4_1(.din(w_dff_B_8v1f5lu64_1),.dout(w_dff_B_qDMTBvTM4_1),.clk(gclk));
	jdff dff_B_RpTJ8ne29_1(.din(w_dff_B_qDMTBvTM4_1),.dout(w_dff_B_RpTJ8ne29_1),.clk(gclk));
	jdff dff_B_AshLw6qE3_1(.din(w_dff_B_RpTJ8ne29_1),.dout(w_dff_B_AshLw6qE3_1),.clk(gclk));
	jdff dff_B_Tc9xDrxg9_1(.din(w_dff_B_AshLw6qE3_1),.dout(w_dff_B_Tc9xDrxg9_1),.clk(gclk));
	jdff dff_B_5mxyAtXC7_1(.din(w_dff_B_Tc9xDrxg9_1),.dout(w_dff_B_5mxyAtXC7_1),.clk(gclk));
	jdff dff_B_nrRkeC0n1_1(.din(w_dff_B_5mxyAtXC7_1),.dout(w_dff_B_nrRkeC0n1_1),.clk(gclk));
	jdff dff_B_sJ1BlAHw3_1(.din(w_dff_B_nrRkeC0n1_1),.dout(w_dff_B_sJ1BlAHw3_1),.clk(gclk));
	jdff dff_B_NgtP7nAb7_1(.din(w_dff_B_sJ1BlAHw3_1),.dout(w_dff_B_NgtP7nAb7_1),.clk(gclk));
	jdff dff_B_rae1xR3N7_1(.din(w_dff_B_NgtP7nAb7_1),.dout(w_dff_B_rae1xR3N7_1),.clk(gclk));
	jdff dff_B_IK8yuc0C4_1(.din(w_dff_B_rae1xR3N7_1),.dout(w_dff_B_IK8yuc0C4_1),.clk(gclk));
	jdff dff_B_3kuzFPr53_1(.din(w_dff_B_IK8yuc0C4_1),.dout(w_dff_B_3kuzFPr53_1),.clk(gclk));
	jdff dff_B_CyWgGN208_1(.din(w_dff_B_3kuzFPr53_1),.dout(w_dff_B_CyWgGN208_1),.clk(gclk));
	jdff dff_B_NNvIj3sz2_1(.din(w_dff_B_CyWgGN208_1),.dout(w_dff_B_NNvIj3sz2_1),.clk(gclk));
	jdff dff_B_qnAH5L7I0_1(.din(w_dff_B_NNvIj3sz2_1),.dout(w_dff_B_qnAH5L7I0_1),.clk(gclk));
	jdff dff_B_RgWgAMLJ0_1(.din(w_dff_B_qnAH5L7I0_1),.dout(w_dff_B_RgWgAMLJ0_1),.clk(gclk));
	jdff dff_B_Jrt6afgO4_1(.din(w_dff_B_RgWgAMLJ0_1),.dout(w_dff_B_Jrt6afgO4_1),.clk(gclk));
	jdff dff_B_4gExAVhN2_1(.din(w_dff_B_Jrt6afgO4_1),.dout(w_dff_B_4gExAVhN2_1),.clk(gclk));
	jdff dff_B_lwVZCQWe7_1(.din(w_dff_B_4gExAVhN2_1),.dout(w_dff_B_lwVZCQWe7_1),.clk(gclk));
	jdff dff_B_nd1RsLIr9_1(.din(w_dff_B_lwVZCQWe7_1),.dout(w_dff_B_nd1RsLIr9_1),.clk(gclk));
	jdff dff_B_HCXKnUV56_1(.din(n1328),.dout(w_dff_B_HCXKnUV56_1),.clk(gclk));
	jdff dff_B_44gYAvYT5_1(.din(w_dff_B_HCXKnUV56_1),.dout(w_dff_B_44gYAvYT5_1),.clk(gclk));
	jdff dff_B_ODsjwKZU9_1(.din(w_dff_B_44gYAvYT5_1),.dout(w_dff_B_ODsjwKZU9_1),.clk(gclk));
	jdff dff_B_ohRFURxK8_1(.din(w_dff_B_ODsjwKZU9_1),.dout(w_dff_B_ohRFURxK8_1),.clk(gclk));
	jdff dff_B_hw8qqWUl6_1(.din(w_dff_B_ohRFURxK8_1),.dout(w_dff_B_hw8qqWUl6_1),.clk(gclk));
	jdff dff_B_ZFrDDfpJ6_1(.din(w_dff_B_hw8qqWUl6_1),.dout(w_dff_B_ZFrDDfpJ6_1),.clk(gclk));
	jdff dff_B_D5IQZtkR1_1(.din(w_dff_B_ZFrDDfpJ6_1),.dout(w_dff_B_D5IQZtkR1_1),.clk(gclk));
	jdff dff_B_UPCU2CmB6_1(.din(w_dff_B_D5IQZtkR1_1),.dout(w_dff_B_UPCU2CmB6_1),.clk(gclk));
	jdff dff_B_u6yzwprT5_1(.din(w_dff_B_UPCU2CmB6_1),.dout(w_dff_B_u6yzwprT5_1),.clk(gclk));
	jdff dff_B_BonRRWPv8_1(.din(w_dff_B_u6yzwprT5_1),.dout(w_dff_B_BonRRWPv8_1),.clk(gclk));
	jdff dff_B_77XlgZEc1_1(.din(w_dff_B_BonRRWPv8_1),.dout(w_dff_B_77XlgZEc1_1),.clk(gclk));
	jdff dff_B_Akr6oeE66_1(.din(w_dff_B_77XlgZEc1_1),.dout(w_dff_B_Akr6oeE66_1),.clk(gclk));
	jdff dff_B_D03abrMJ9_1(.din(w_dff_B_Akr6oeE66_1),.dout(w_dff_B_D03abrMJ9_1),.clk(gclk));
	jdff dff_B_8lvX44m70_1(.din(w_dff_B_D03abrMJ9_1),.dout(w_dff_B_8lvX44m70_1),.clk(gclk));
	jdff dff_B_MQlJAE9M7_1(.din(w_dff_B_8lvX44m70_1),.dout(w_dff_B_MQlJAE9M7_1),.clk(gclk));
	jdff dff_B_NAgtVxZD0_1(.din(w_dff_B_MQlJAE9M7_1),.dout(w_dff_B_NAgtVxZD0_1),.clk(gclk));
	jdff dff_B_Y5YldpcH8_1(.din(n1329),.dout(w_dff_B_Y5YldpcH8_1),.clk(gclk));
	jdff dff_B_DP4CX1mM1_1(.din(w_dff_B_Y5YldpcH8_1),.dout(w_dff_B_DP4CX1mM1_1),.clk(gclk));
	jdff dff_B_5tklbAaM3_1(.din(w_dff_B_DP4CX1mM1_1),.dout(w_dff_B_5tklbAaM3_1),.clk(gclk));
	jdff dff_B_Byl5Z62t8_1(.din(w_dff_B_5tklbAaM3_1),.dout(w_dff_B_Byl5Z62t8_1),.clk(gclk));
	jdff dff_B_ytgcOuN60_1(.din(w_dff_B_Byl5Z62t8_1),.dout(w_dff_B_ytgcOuN60_1),.clk(gclk));
	jdff dff_B_0kADtmeq4_1(.din(w_dff_B_ytgcOuN60_1),.dout(w_dff_B_0kADtmeq4_1),.clk(gclk));
	jdff dff_B_u6FH1tbz5_1(.din(w_dff_B_0kADtmeq4_1),.dout(w_dff_B_u6FH1tbz5_1),.clk(gclk));
	jdff dff_B_jW935lNA8_1(.din(w_dff_B_u6FH1tbz5_1),.dout(w_dff_B_jW935lNA8_1),.clk(gclk));
	jdff dff_B_rLGvwbtD6_1(.din(w_dff_B_jW935lNA8_1),.dout(w_dff_B_rLGvwbtD6_1),.clk(gclk));
	jdff dff_B_nlH3rkY76_1(.din(w_dff_B_rLGvwbtD6_1),.dout(w_dff_B_nlH3rkY76_1),.clk(gclk));
	jdff dff_B_i7s5kYnd1_1(.din(w_dff_B_nlH3rkY76_1),.dout(w_dff_B_i7s5kYnd1_1),.clk(gclk));
	jdff dff_B_wYoPpZ6N7_1(.din(w_dff_B_i7s5kYnd1_1),.dout(w_dff_B_wYoPpZ6N7_1),.clk(gclk));
	jdff dff_B_YTdOoUHr3_1(.din(w_dff_B_wYoPpZ6N7_1),.dout(w_dff_B_YTdOoUHr3_1),.clk(gclk));
	jdff dff_B_e52IBdTD4_1(.din(w_dff_B_YTdOoUHr3_1),.dout(w_dff_B_e52IBdTD4_1),.clk(gclk));
	jdff dff_B_j0QpTQHF5_1(.din(w_dff_B_e52IBdTD4_1),.dout(w_dff_B_j0QpTQHF5_1),.clk(gclk));
	jdff dff_B_TOdfTB2l7_1(.din(w_dff_B_j0QpTQHF5_1),.dout(w_dff_B_TOdfTB2l7_1),.clk(gclk));
	jdff dff_B_rHabs0Ds3_1(.din(w_dff_B_TOdfTB2l7_1),.dout(w_dff_B_rHabs0Ds3_1),.clk(gclk));
	jdff dff_B_xlnIwjUB5_1(.din(n1330),.dout(w_dff_B_xlnIwjUB5_1),.clk(gclk));
	jdff dff_B_epeUJmat6_1(.din(w_dff_B_xlnIwjUB5_1),.dout(w_dff_B_epeUJmat6_1),.clk(gclk));
	jdff dff_B_3bOwUSDR6_1(.din(w_dff_B_epeUJmat6_1),.dout(w_dff_B_3bOwUSDR6_1),.clk(gclk));
	jdff dff_B_7oCASZGe3_1(.din(w_dff_B_3bOwUSDR6_1),.dout(w_dff_B_7oCASZGe3_1),.clk(gclk));
	jdff dff_B_4VyW49zX9_1(.din(w_dff_B_7oCASZGe3_1),.dout(w_dff_B_4VyW49zX9_1),.clk(gclk));
	jdff dff_B_pk97WiTA1_1(.din(w_dff_B_4VyW49zX9_1),.dout(w_dff_B_pk97WiTA1_1),.clk(gclk));
	jdff dff_B_xZKYKqV27_1(.din(w_dff_B_pk97WiTA1_1),.dout(w_dff_B_xZKYKqV27_1),.clk(gclk));
	jdff dff_B_Mz1q1YI47_1(.din(w_dff_B_xZKYKqV27_1),.dout(w_dff_B_Mz1q1YI47_1),.clk(gclk));
	jdff dff_B_o1XJSCTh3_1(.din(w_dff_B_Mz1q1YI47_1),.dout(w_dff_B_o1XJSCTh3_1),.clk(gclk));
	jdff dff_B_IGC0S6jD6_1(.din(w_dff_B_o1XJSCTh3_1),.dout(w_dff_B_IGC0S6jD6_1),.clk(gclk));
	jdff dff_B_aTPdqReg6_1(.din(w_dff_B_IGC0S6jD6_1),.dout(w_dff_B_aTPdqReg6_1),.clk(gclk));
	jdff dff_B_vxIYgitq5_1(.din(w_dff_B_aTPdqReg6_1),.dout(w_dff_B_vxIYgitq5_1),.clk(gclk));
	jdff dff_B_ZXtwGK773_1(.din(w_dff_B_vxIYgitq5_1),.dout(w_dff_B_ZXtwGK773_1),.clk(gclk));
	jdff dff_B_2iFnCUuU8_1(.din(w_dff_B_ZXtwGK773_1),.dout(w_dff_B_2iFnCUuU8_1),.clk(gclk));
	jdff dff_B_RsyCdviq3_1(.din(w_dff_B_2iFnCUuU8_1),.dout(w_dff_B_RsyCdviq3_1),.clk(gclk));
	jdff dff_B_nfriTmIm4_1(.din(w_dff_B_RsyCdviq3_1),.dout(w_dff_B_nfriTmIm4_1),.clk(gclk));
	jdff dff_B_oO0jZObY5_1(.din(w_dff_B_nfriTmIm4_1),.dout(w_dff_B_oO0jZObY5_1),.clk(gclk));
	jdff dff_B_BrvrR8gC2_1(.din(w_dff_B_oO0jZObY5_1),.dout(w_dff_B_BrvrR8gC2_1),.clk(gclk));
	jdff dff_B_LJxHPsYZ4_1(.din(w_dff_B_BrvrR8gC2_1),.dout(w_dff_B_LJxHPsYZ4_1),.clk(gclk));
	jdff dff_B_luDCltd93_1(.din(w_dff_B_LJxHPsYZ4_1),.dout(w_dff_B_luDCltd93_1),.clk(gclk));
	jdff dff_B_jDfHQxtX6_1(.din(n1306),.dout(w_dff_B_jDfHQxtX6_1),.clk(gclk));
	jdff dff_B_padfVtME6_1(.din(w_dff_B_jDfHQxtX6_1),.dout(w_dff_B_padfVtME6_1),.clk(gclk));
	jdff dff_B_YNsgfuEa4_1(.din(w_dff_B_padfVtME6_1),.dout(w_dff_B_YNsgfuEa4_1),.clk(gclk));
	jdff dff_B_ySbCi0UA4_1(.din(w_dff_B_YNsgfuEa4_1),.dout(w_dff_B_ySbCi0UA4_1),.clk(gclk));
	jdff dff_B_sT2LG1VA4_1(.din(w_dff_B_ySbCi0UA4_1),.dout(w_dff_B_sT2LG1VA4_1),.clk(gclk));
	jdff dff_B_VkuhmvWQ4_1(.din(w_dff_B_sT2LG1VA4_1),.dout(w_dff_B_VkuhmvWQ4_1),.clk(gclk));
	jdff dff_B_weELPwBH8_1(.din(w_dff_B_VkuhmvWQ4_1),.dout(w_dff_B_weELPwBH8_1),.clk(gclk));
	jdff dff_B_MoK8K3V77_1(.din(w_dff_B_weELPwBH8_1),.dout(w_dff_B_MoK8K3V77_1),.clk(gclk));
	jdff dff_B_aFiCM8Xa7_1(.din(w_dff_B_MoK8K3V77_1),.dout(w_dff_B_aFiCM8Xa7_1),.clk(gclk));
	jdff dff_B_RmXhfKrA5_1(.din(w_dff_B_aFiCM8Xa7_1),.dout(w_dff_B_RmXhfKrA5_1),.clk(gclk));
	jdff dff_B_A9342yTM3_1(.din(w_dff_B_RmXhfKrA5_1),.dout(w_dff_B_A9342yTM3_1),.clk(gclk));
	jdff dff_B_DuUQPFvb7_1(.din(w_dff_B_A9342yTM3_1),.dout(w_dff_B_DuUQPFvb7_1),.clk(gclk));
	jdff dff_B_uo74DPz82_1(.din(w_dff_B_DuUQPFvb7_1),.dout(w_dff_B_uo74DPz82_1),.clk(gclk));
	jdff dff_B_PncgLYtv6_1(.din(w_dff_B_uo74DPz82_1),.dout(w_dff_B_PncgLYtv6_1),.clk(gclk));
	jdff dff_B_1oMPnq7s8_1(.din(w_dff_B_PncgLYtv6_1),.dout(w_dff_B_1oMPnq7s8_1),.clk(gclk));
	jdff dff_B_Y4voQsKt4_1(.din(w_dff_B_1oMPnq7s8_1),.dout(w_dff_B_Y4voQsKt4_1),.clk(gclk));
	jdff dff_B_6ZOy3w3J2_1(.din(w_dff_B_Y4voQsKt4_1),.dout(w_dff_B_6ZOy3w3J2_1),.clk(gclk));
	jdff dff_B_OcKKJx5L0_1(.din(w_dff_B_6ZOy3w3J2_1),.dout(w_dff_B_OcKKJx5L0_1),.clk(gclk));
	jdff dff_B_MLZPxglE7_1(.din(w_dff_B_OcKKJx5L0_1),.dout(w_dff_B_MLZPxglE7_1),.clk(gclk));
	jdff dff_B_1H8NVeIm3_1(.din(w_dff_B_MLZPxglE7_1),.dout(w_dff_B_1H8NVeIm3_1),.clk(gclk));
	jdff dff_B_ikio3lpP7_1(.din(w_dff_B_1H8NVeIm3_1),.dout(w_dff_B_ikio3lpP7_1),.clk(gclk));
	jdff dff_A_IuxooMrp3_0(.dout(w_n1307_0[0]),.din(w_dff_A_IuxooMrp3_0),.clk(gclk));
	jdff dff_B_g5yGYdSh2_2(.din(n1307),.dout(w_dff_B_g5yGYdSh2_2),.clk(gclk));
	jdff dff_B_roBgkliS7_2(.din(w_dff_B_g5yGYdSh2_2),.dout(w_dff_B_roBgkliS7_2),.clk(gclk));
	jdff dff_B_5yXtPHCI4_2(.din(w_dff_B_roBgkliS7_2),.dout(w_dff_B_5yXtPHCI4_2),.clk(gclk));
	jdff dff_B_czORjX8i6_2(.din(w_dff_B_5yXtPHCI4_2),.dout(w_dff_B_czORjX8i6_2),.clk(gclk));
	jdff dff_B_vkNiYCuI6_2(.din(w_dff_B_czORjX8i6_2),.dout(w_dff_B_vkNiYCuI6_2),.clk(gclk));
	jdff dff_B_AamhJqBS7_2(.din(w_dff_B_vkNiYCuI6_2),.dout(w_dff_B_AamhJqBS7_2),.clk(gclk));
	jdff dff_B_omN9lnRC1_2(.din(w_dff_B_AamhJqBS7_2),.dout(w_dff_B_omN9lnRC1_2),.clk(gclk));
	jdff dff_B_BvWSSrzu4_2(.din(w_dff_B_omN9lnRC1_2),.dout(w_dff_B_BvWSSrzu4_2),.clk(gclk));
	jdff dff_B_V4gj3nKw4_2(.din(w_dff_B_BvWSSrzu4_2),.dout(w_dff_B_V4gj3nKw4_2),.clk(gclk));
	jdff dff_B_SMP7N7Ck0_2(.din(w_dff_B_V4gj3nKw4_2),.dout(w_dff_B_SMP7N7Ck0_2),.clk(gclk));
	jdff dff_B_Up4m6slZ1_2(.din(w_dff_B_SMP7N7Ck0_2),.dout(w_dff_B_Up4m6slZ1_2),.clk(gclk));
	jdff dff_B_UrTGNWhK7_2(.din(w_dff_B_Up4m6slZ1_2),.dout(w_dff_B_UrTGNWhK7_2),.clk(gclk));
	jdff dff_B_mBdl030i6_2(.din(w_dff_B_UrTGNWhK7_2),.dout(w_dff_B_mBdl030i6_2),.clk(gclk));
	jdff dff_B_8pQKnd758_2(.din(w_dff_B_mBdl030i6_2),.dout(w_dff_B_8pQKnd758_2),.clk(gclk));
	jdff dff_B_6ObSEDAw4_2(.din(w_dff_B_8pQKnd758_2),.dout(w_dff_B_6ObSEDAw4_2),.clk(gclk));
	jdff dff_B_KGY4CxUr5_2(.din(w_dff_B_6ObSEDAw4_2),.dout(w_dff_B_KGY4CxUr5_2),.clk(gclk));
	jdff dff_B_qXfQcp5F7_2(.din(w_dff_B_KGY4CxUr5_2),.dout(w_dff_B_qXfQcp5F7_2),.clk(gclk));
	jdff dff_B_Y5woxDGt8_2(.din(w_dff_B_qXfQcp5F7_2),.dout(w_dff_B_Y5woxDGt8_2),.clk(gclk));
	jdff dff_B_AGhvN9KA2_0(.din(n1490),.dout(w_dff_B_AGhvN9KA2_0),.clk(gclk));
	jdff dff_B_0gJncxEk9_0(.din(w_dff_B_AGhvN9KA2_0),.dout(w_dff_B_0gJncxEk9_0),.clk(gclk));
	jdff dff_B_AdBgfhpW3_0(.din(w_dff_B_0gJncxEk9_0),.dout(w_dff_B_AdBgfhpW3_0),.clk(gclk));
	jdff dff_B_0TCVwuZs8_0(.din(w_dff_B_AdBgfhpW3_0),.dout(w_dff_B_0TCVwuZs8_0),.clk(gclk));
	jdff dff_B_rfKLOvf55_0(.din(w_dff_B_0TCVwuZs8_0),.dout(w_dff_B_rfKLOvf55_0),.clk(gclk));
	jdff dff_B_05v4G4EF4_0(.din(w_dff_B_rfKLOvf55_0),.dout(w_dff_B_05v4G4EF4_0),.clk(gclk));
	jdff dff_B_FOqQI0gV0_0(.din(w_dff_B_05v4G4EF4_0),.dout(w_dff_B_FOqQI0gV0_0),.clk(gclk));
	jdff dff_B_8ImvVHjO3_0(.din(w_dff_B_FOqQI0gV0_0),.dout(w_dff_B_8ImvVHjO3_0),.clk(gclk));
	jdff dff_B_X2YReIlf9_0(.din(w_dff_B_8ImvVHjO3_0),.dout(w_dff_B_X2YReIlf9_0),.clk(gclk));
	jdff dff_B_LZXWKBZ50_0(.din(w_dff_B_X2YReIlf9_0),.dout(w_dff_B_LZXWKBZ50_0),.clk(gclk));
	jdff dff_B_9xnFQAWl5_0(.din(w_dff_B_LZXWKBZ50_0),.dout(w_dff_B_9xnFQAWl5_0),.clk(gclk));
	jdff dff_B_98YENKx82_0(.din(w_dff_B_9xnFQAWl5_0),.dout(w_dff_B_98YENKx82_0),.clk(gclk));
	jdff dff_B_E4vM521R1_0(.din(w_dff_B_98YENKx82_0),.dout(w_dff_B_E4vM521R1_0),.clk(gclk));
	jdff dff_B_L07YgFGf5_0(.din(w_dff_B_E4vM521R1_0),.dout(w_dff_B_L07YgFGf5_0),.clk(gclk));
	jdff dff_B_svOPQ0IX8_0(.din(w_dff_B_L07YgFGf5_0),.dout(w_dff_B_svOPQ0IX8_0),.clk(gclk));
	jdff dff_B_XoqK1Qrf7_0(.din(w_dff_B_svOPQ0IX8_0),.dout(w_dff_B_XoqK1Qrf7_0),.clk(gclk));
	jdff dff_B_mNVELAZ65_0(.din(w_dff_B_XoqK1Qrf7_0),.dout(w_dff_B_mNVELAZ65_0),.clk(gclk));
	jdff dff_B_wNjScP6a2_0(.din(w_dff_B_mNVELAZ65_0),.dout(w_dff_B_wNjScP6a2_0),.clk(gclk));
	jdff dff_B_F1pYMPkp7_0(.din(w_dff_B_wNjScP6a2_0),.dout(w_dff_B_F1pYMPkp7_0),.clk(gclk));
	jdff dff_B_f6SH1Swa5_0(.din(w_dff_B_F1pYMPkp7_0),.dout(w_dff_B_f6SH1Swa5_0),.clk(gclk));
	jdff dff_B_QktJqICt2_0(.din(w_dff_B_f6SH1Swa5_0),.dout(w_dff_B_QktJqICt2_0),.clk(gclk));
	jdff dff_B_sF6oPbsM6_0(.din(n1488),.dout(w_dff_B_sF6oPbsM6_0),.clk(gclk));
	jdff dff_B_5kIPSHbN4_0(.din(w_dff_B_sF6oPbsM6_0),.dout(w_dff_B_5kIPSHbN4_0),.clk(gclk));
	jdff dff_B_4T9BR8210_0(.din(w_dff_B_5kIPSHbN4_0),.dout(w_dff_B_4T9BR8210_0),.clk(gclk));
	jdff dff_B_Kzz4PDiU8_0(.din(n1487),.dout(w_dff_B_Kzz4PDiU8_0),.clk(gclk));
	jdff dff_B_nODN7bvz1_0(.din(w_dff_B_Kzz4PDiU8_0),.dout(w_dff_B_nODN7bvz1_0),.clk(gclk));
	jdff dff_A_gwZYhnKO5_1(.dout(w_n414_0[1]),.din(w_dff_A_gwZYhnKO5_1),.clk(gclk));
	jdff dff_A_RvPdg9DA4_1(.dout(w_dff_A_gwZYhnKO5_1),.din(w_dff_A_RvPdg9DA4_1),.clk(gclk));
	jdff dff_A_r5vwT7TT8_1(.dout(w_dff_A_RvPdg9DA4_1),.din(w_dff_A_r5vwT7TT8_1),.clk(gclk));
	jdff dff_A_0EY8Gc0Y3_1(.dout(w_dff_A_r5vwT7TT8_1),.din(w_dff_A_0EY8Gc0Y3_1),.clk(gclk));
	jdff dff_A_L9KEOYBB9_1(.dout(w_dff_A_0EY8Gc0Y3_1),.din(w_dff_A_L9KEOYBB9_1),.clk(gclk));
	jdff dff_A_m5ViydYv5_1(.dout(w_dff_A_L9KEOYBB9_1),.din(w_dff_A_m5ViydYv5_1),.clk(gclk));
	jdff dff_A_yoPZSWl13_1(.dout(w_dff_A_m5ViydYv5_1),.din(w_dff_A_yoPZSWl13_1),.clk(gclk));
	jdff dff_A_qWKx2dOq8_1(.dout(w_dff_A_yoPZSWl13_1),.din(w_dff_A_qWKx2dOq8_1),.clk(gclk));
	jdff dff_B_eFgGSVwm2_1(.din(n1482),.dout(w_dff_B_eFgGSVwm2_1),.clk(gclk));
	jdff dff_B_0FngQeLD3_1(.din(w_dff_B_eFgGSVwm2_1),.dout(w_dff_B_0FngQeLD3_1),.clk(gclk));
	jdff dff_A_eZXnlpvS8_1(.dout(w_n1370_0[1]),.din(w_dff_A_eZXnlpvS8_1),.clk(gclk));
	jdff dff_A_6h3bIYF37_1(.dout(w_dff_A_eZXnlpvS8_1),.din(w_dff_A_6h3bIYF37_1),.clk(gclk));
	jdff dff_A_7VYmYoYr9_1(.dout(w_dff_A_6h3bIYF37_1),.din(w_dff_A_7VYmYoYr9_1),.clk(gclk));
	jdff dff_A_2poalKMA2_1(.dout(w_dff_A_7VYmYoYr9_1),.din(w_dff_A_2poalKMA2_1),.clk(gclk));
	jdff dff_A_KIx2VHi19_1(.dout(w_dff_A_2poalKMA2_1),.din(w_dff_A_KIx2VHi19_1),.clk(gclk));
	jdff dff_A_5cO6ktaw9_1(.dout(w_dff_A_KIx2VHi19_1),.din(w_dff_A_5cO6ktaw9_1),.clk(gclk));
	jdff dff_A_JejYPRDo3_1(.dout(w_dff_A_5cO6ktaw9_1),.din(w_dff_A_JejYPRDo3_1),.clk(gclk));
	jdff dff_A_wCJ2uaZ43_1(.dout(w_dff_A_JejYPRDo3_1),.din(w_dff_A_wCJ2uaZ43_1),.clk(gclk));
	jdff dff_A_6xxYKv2a0_1(.dout(w_dff_A_wCJ2uaZ43_1),.din(w_dff_A_6xxYKv2a0_1),.clk(gclk));
	jdff dff_A_tylyX5up8_1(.dout(w_dff_A_6xxYKv2a0_1),.din(w_dff_A_tylyX5up8_1),.clk(gclk));
	jdff dff_A_EZadv2aC4_1(.dout(w_dff_A_tylyX5up8_1),.din(w_dff_A_EZadv2aC4_1),.clk(gclk));
	jdff dff_A_K311HNM89_1(.dout(w_dff_A_EZadv2aC4_1),.din(w_dff_A_K311HNM89_1),.clk(gclk));
	jdff dff_A_3pwP2hv86_1(.dout(w_dff_A_K311HNM89_1),.din(w_dff_A_3pwP2hv86_1),.clk(gclk));
	jdff dff_A_4NJksY3z7_1(.dout(w_dff_A_3pwP2hv86_1),.din(w_dff_A_4NJksY3z7_1),.clk(gclk));
	jdff dff_A_1Mj12XJM8_1(.dout(w_dff_A_4NJksY3z7_1),.din(w_dff_A_1Mj12XJM8_1),.clk(gclk));
	jdff dff_A_fEZDBPaJ9_1(.dout(w_dff_A_1Mj12XJM8_1),.din(w_dff_A_fEZDBPaJ9_1),.clk(gclk));
	jdff dff_A_9ZwlWKzu7_1(.dout(w_dff_A_fEZDBPaJ9_1),.din(w_dff_A_9ZwlWKzu7_1),.clk(gclk));
	jdff dff_A_BZTD7tpw2_1(.dout(w_dff_A_9ZwlWKzu7_1),.din(w_dff_A_BZTD7tpw2_1),.clk(gclk));
	jdff dff_A_qjjDobR02_1(.dout(w_dff_A_BZTD7tpw2_1),.din(w_dff_A_qjjDobR02_1),.clk(gclk));
	jdff dff_A_OjhF358c0_1(.dout(w_dff_A_qjjDobR02_1),.din(w_dff_A_OjhF358c0_1),.clk(gclk));
	jdff dff_A_Tz7kdlG23_1(.dout(w_dff_A_OjhF358c0_1),.din(w_dff_A_Tz7kdlG23_1),.clk(gclk));
	jdff dff_A_9McRTXCu6_1(.dout(w_dff_A_Tz7kdlG23_1),.din(w_dff_A_9McRTXCu6_1),.clk(gclk));
	jdff dff_A_XBoqCcEx7_1(.dout(w_dff_A_9McRTXCu6_1),.din(w_dff_A_XBoqCcEx7_1),.clk(gclk));
	jdff dff_A_fdzOriLl1_1(.dout(w_dff_A_XBoqCcEx7_1),.din(w_dff_A_fdzOriLl1_1),.clk(gclk));
	jdff dff_A_vYHgwxc30_1(.dout(w_dff_A_fdzOriLl1_1),.din(w_dff_A_vYHgwxc30_1),.clk(gclk));
	jdff dff_A_PZw6Hh9P7_1(.dout(w_dff_A_vYHgwxc30_1),.din(w_dff_A_PZw6Hh9P7_1),.clk(gclk));
	jdff dff_A_jarPTf8q0_1(.dout(w_dff_A_PZw6Hh9P7_1),.din(w_dff_A_jarPTf8q0_1),.clk(gclk));
	jdff dff_A_Mo5ZWezW7_1(.dout(w_dff_A_jarPTf8q0_1),.din(w_dff_A_Mo5ZWezW7_1),.clk(gclk));
	jdff dff_B_AnofVKPO2_2(.din(n1370),.dout(w_dff_B_AnofVKPO2_2),.clk(gclk));
	jdff dff_B_lJ5QNjnV4_2(.din(w_dff_B_AnofVKPO2_2),.dout(w_dff_B_lJ5QNjnV4_2),.clk(gclk));
	jdff dff_A_g92e85O21_2(.dout(w_n411_0[2]),.din(w_dff_A_g92e85O21_2),.clk(gclk));
	jdff dff_A_aglXCVb96_2(.dout(w_dff_A_g92e85O21_2),.din(w_dff_A_aglXCVb96_2),.clk(gclk));
	jdff dff_A_YWRAjuvE8_2(.dout(w_dff_A_aglXCVb96_2),.din(w_dff_A_YWRAjuvE8_2),.clk(gclk));
	jdff dff_A_i34odZJ98_2(.dout(w_dff_A_YWRAjuvE8_2),.din(w_dff_A_i34odZJ98_2),.clk(gclk));
	jdff dff_A_3uf1oS8C3_2(.dout(w_dff_A_i34odZJ98_2),.din(w_dff_A_3uf1oS8C3_2),.clk(gclk));
	jdff dff_A_fYTI9cJ48_2(.dout(w_dff_A_3uf1oS8C3_2),.din(w_dff_A_fYTI9cJ48_2),.clk(gclk));
	jdff dff_A_AevRGeN78_2(.dout(w_dff_A_fYTI9cJ48_2),.din(w_dff_A_AevRGeN78_2),.clk(gclk));
	jdff dff_A_3J8NWZDi6_2(.dout(w_dff_A_AevRGeN78_2),.din(w_dff_A_3J8NWZDi6_2),.clk(gclk));
	jdff dff_A_TnqrOvdt0_2(.dout(w_dff_A_3J8NWZDi6_2),.din(w_dff_A_TnqrOvdt0_2),.clk(gclk));
	jdff dff_A_51aRyeB72_2(.dout(w_dff_A_TnqrOvdt0_2),.din(w_dff_A_51aRyeB72_2),.clk(gclk));
	jdff dff_A_woUc07xg0_2(.dout(w_dff_A_51aRyeB72_2),.din(w_dff_A_woUc07xg0_2),.clk(gclk));
	jdff dff_A_IjzyheDb7_2(.dout(w_dff_A_woUc07xg0_2),.din(w_dff_A_IjzyheDb7_2),.clk(gclk));
	jdff dff_A_CxhTikps9_2(.dout(w_dff_A_IjzyheDb7_2),.din(w_dff_A_CxhTikps9_2),.clk(gclk));
	jdff dff_A_MQNbCX390_2(.dout(w_dff_A_CxhTikps9_2),.din(w_dff_A_MQNbCX390_2),.clk(gclk));
	jdff dff_A_UE8spiDH8_2(.dout(w_dff_A_MQNbCX390_2),.din(w_dff_A_UE8spiDH8_2),.clk(gclk));
	jdff dff_A_qrthNcPY3_2(.dout(w_dff_A_UE8spiDH8_2),.din(w_dff_A_qrthNcPY3_2),.clk(gclk));
	jdff dff_A_nXS0nba76_2(.dout(w_dff_A_qrthNcPY3_2),.din(w_dff_A_nXS0nba76_2),.clk(gclk));
	jdff dff_A_W52wLRxE4_2(.dout(w_dff_A_nXS0nba76_2),.din(w_dff_A_W52wLRxE4_2),.clk(gclk));
	jdff dff_A_jRNRbCtR5_2(.dout(w_dff_A_W52wLRxE4_2),.din(w_dff_A_jRNRbCtR5_2),.clk(gclk));
	jdff dff_A_v90dEzJ47_2(.dout(w_dff_A_jRNRbCtR5_2),.din(w_dff_A_v90dEzJ47_2),.clk(gclk));
	jdff dff_A_DvqT2GfO2_2(.dout(w_dff_A_v90dEzJ47_2),.din(w_dff_A_DvqT2GfO2_2),.clk(gclk));
	jdff dff_A_gAZ44v0g8_2(.dout(w_dff_A_DvqT2GfO2_2),.din(w_dff_A_gAZ44v0g8_2),.clk(gclk));
	jdff dff_A_C5SgrmPL0_2(.dout(w_dff_A_gAZ44v0g8_2),.din(w_dff_A_C5SgrmPL0_2),.clk(gclk));
	jdff dff_B_Xzk5kxbQ0_1(.din(n382),.dout(w_dff_B_Xzk5kxbQ0_1),.clk(gclk));
	jdff dff_B_EDueLPXN5_1(.din(w_dff_B_Xzk5kxbQ0_1),.dout(w_dff_B_EDueLPXN5_1),.clk(gclk));
	jdff dff_B_pYGNNO9i9_1(.din(w_dff_B_EDueLPXN5_1),.dout(w_dff_B_pYGNNO9i9_1),.clk(gclk));
	jdff dff_B_9j5IoNto8_1(.din(w_dff_B_pYGNNO9i9_1),.dout(w_dff_B_9j5IoNto8_1),.clk(gclk));
	jdff dff_B_RWZ0nrv75_1(.din(n384),.dout(w_dff_B_RWZ0nrv75_1),.clk(gclk));
	jdff dff_B_erbnnowH2_1(.din(w_dff_B_RWZ0nrv75_1),.dout(w_dff_B_erbnnowH2_1),.clk(gclk));
	jdff dff_B_R04qSkmn0_1(.din(w_dff_B_erbnnowH2_1),.dout(w_dff_B_R04qSkmn0_1),.clk(gclk));
	jdff dff_B_ZQDWXIqq6_1(.din(w_dff_B_R04qSkmn0_1),.dout(w_dff_B_ZQDWXIqq6_1),.clk(gclk));
	jdff dff_B_Cw6wK2kq0_1(.din(w_dff_B_ZQDWXIqq6_1),.dout(w_dff_B_Cw6wK2kq0_1),.clk(gclk));
	jdff dff_A_BrJEZedj3_2(.dout(w_n409_0[2]),.din(w_dff_A_BrJEZedj3_2),.clk(gclk));
	jdff dff_A_HHPEyq3M9_2(.dout(w_dff_A_BrJEZedj3_2),.din(w_dff_A_HHPEyq3M9_2),.clk(gclk));
	jdff dff_A_CJL8xyZz6_2(.dout(w_dff_A_HHPEyq3M9_2),.din(w_dff_A_CJL8xyZz6_2),.clk(gclk));
	jdff dff_A_dVODatoS0_2(.dout(w_dff_A_CJL8xyZz6_2),.din(w_dff_A_dVODatoS0_2),.clk(gclk));
	jdff dff_A_oU1ZM55K8_2(.dout(w_dff_A_dVODatoS0_2),.din(w_dff_A_oU1ZM55K8_2),.clk(gclk));
	jdff dff_A_sGjIIncj7_2(.dout(w_dff_A_oU1ZM55K8_2),.din(w_dff_A_sGjIIncj7_2),.clk(gclk));
	jdff dff_A_6llkRCZ02_2(.dout(w_dff_A_sGjIIncj7_2),.din(w_dff_A_6llkRCZ02_2),.clk(gclk));
	jdff dff_A_SIOtIOml7_2(.dout(w_dff_A_6llkRCZ02_2),.din(w_dff_A_SIOtIOml7_2),.clk(gclk));
	jdff dff_A_glWGlEd73_2(.dout(w_dff_A_SIOtIOml7_2),.din(w_dff_A_glWGlEd73_2),.clk(gclk));
	jdff dff_A_Cgz9fZJ48_2(.dout(w_dff_A_glWGlEd73_2),.din(w_dff_A_Cgz9fZJ48_2),.clk(gclk));
	jdff dff_A_OILiBMmN9_2(.dout(w_dff_A_Cgz9fZJ48_2),.din(w_dff_A_OILiBMmN9_2),.clk(gclk));
	jdff dff_A_XSWRAldS2_2(.dout(w_dff_A_OILiBMmN9_2),.din(w_dff_A_XSWRAldS2_2),.clk(gclk));
	jdff dff_A_9HBIlFH77_2(.dout(w_dff_A_XSWRAldS2_2),.din(w_dff_A_9HBIlFH77_2),.clk(gclk));
	jdff dff_A_skJRAPsS0_2(.dout(w_dff_A_9HBIlFH77_2),.din(w_dff_A_skJRAPsS0_2),.clk(gclk));
	jdff dff_A_SPi4HDhp5_2(.dout(w_dff_A_skJRAPsS0_2),.din(w_dff_A_SPi4HDhp5_2),.clk(gclk));
	jdff dff_A_LoqPWNol5_2(.dout(w_dff_A_SPi4HDhp5_2),.din(w_dff_A_LoqPWNol5_2),.clk(gclk));
	jdff dff_A_UUzoMG4o9_2(.dout(w_dff_A_LoqPWNol5_2),.din(w_dff_A_UUzoMG4o9_2),.clk(gclk));
	jdff dff_A_lhgEor1P6_2(.dout(w_dff_A_UUzoMG4o9_2),.din(w_dff_A_lhgEor1P6_2),.clk(gclk));
	jdff dff_A_zMNFwiqL0_2(.dout(w_dff_A_lhgEor1P6_2),.din(w_dff_A_zMNFwiqL0_2),.clk(gclk));
	jdff dff_A_jYck3y3b9_2(.dout(w_dff_A_zMNFwiqL0_2),.din(w_dff_A_jYck3y3b9_2),.clk(gclk));
	jdff dff_A_2NPYQQ0K2_2(.dout(w_dff_A_jYck3y3b9_2),.din(w_dff_A_2NPYQQ0K2_2),.clk(gclk));
	jdff dff_A_BzExDJok8_2(.dout(w_dff_A_2NPYQQ0K2_2),.din(w_dff_A_BzExDJok8_2),.clk(gclk));
	jdff dff_A_lXNnTDcK2_2(.dout(w_dff_A_BzExDJok8_2),.din(w_dff_A_lXNnTDcK2_2),.clk(gclk));
	jdff dff_A_r0jkB8Pt3_2(.dout(w_dff_A_lXNnTDcK2_2),.din(w_dff_A_r0jkB8Pt3_2),.clk(gclk));
	jdff dff_A_Amuwpa848_2(.dout(w_dff_A_r0jkB8Pt3_2),.din(w_dff_A_Amuwpa848_2),.clk(gclk));
	jdff dff_B_ip9tF0zH7_1(.din(n401),.dout(w_dff_B_ip9tF0zH7_1),.clk(gclk));
	jdff dff_A_0KsNRUZ00_0(.dout(w_n405_0[0]),.din(w_dff_A_0KsNRUZ00_0),.clk(gclk));
	jdff dff_A_Vzst1tsa8_1(.dout(w_n405_0[1]),.din(w_dff_A_Vzst1tsa8_1),.clk(gclk));
	jdff dff_A_HW0CNNaM1_1(.dout(w_dff_A_Vzst1tsa8_1),.din(w_dff_A_HW0CNNaM1_1),.clk(gclk));
	jdff dff_A_LiijGa0q0_1(.dout(w_dff_A_HW0CNNaM1_1),.din(w_dff_A_LiijGa0q0_1),.clk(gclk));
	jdff dff_A_Rk8SrjUc5_1(.dout(w_dff_A_LiijGa0q0_1),.din(w_dff_A_Rk8SrjUc5_1),.clk(gclk));
	jdff dff_A_DSp4yWnr1_1(.dout(w_dff_A_Rk8SrjUc5_1),.din(w_dff_A_DSp4yWnr1_1),.clk(gclk));
	jdff dff_A_LmdZapYT8_1(.dout(w_dff_A_DSp4yWnr1_1),.din(w_dff_A_LmdZapYT8_1),.clk(gclk));
	jdff dff_A_Q4snMDE10_1(.dout(w_dff_A_LmdZapYT8_1),.din(w_dff_A_Q4snMDE10_1),.clk(gclk));
	jdff dff_A_nczq2ASh7_1(.dout(w_dff_A_Q4snMDE10_1),.din(w_dff_A_nczq2ASh7_1),.clk(gclk));
	jdff dff_A_rqdMaNH98_1(.dout(w_dff_A_nczq2ASh7_1),.din(w_dff_A_rqdMaNH98_1),.clk(gclk));
	jdff dff_A_K1SvHrs10_1(.dout(w_dff_A_rqdMaNH98_1),.din(w_dff_A_K1SvHrs10_1),.clk(gclk));
	jdff dff_A_Z4gY4QN91_1(.dout(w_dff_A_K1SvHrs10_1),.din(w_dff_A_Z4gY4QN91_1),.clk(gclk));
	jdff dff_A_v3e3znSJ6_1(.dout(w_dff_A_Z4gY4QN91_1),.din(w_dff_A_v3e3znSJ6_1),.clk(gclk));
	jdff dff_A_986pFOJR1_1(.dout(w_dff_A_v3e3znSJ6_1),.din(w_dff_A_986pFOJR1_1),.clk(gclk));
	jdff dff_A_5DzojULb4_1(.dout(w_dff_A_986pFOJR1_1),.din(w_dff_A_5DzojULb4_1),.clk(gclk));
	jdff dff_A_Wrp4ADXB5_1(.dout(w_dff_A_5DzojULb4_1),.din(w_dff_A_Wrp4ADXB5_1),.clk(gclk));
	jdff dff_A_EKEE6Tlo2_1(.dout(w_dff_A_Wrp4ADXB5_1),.din(w_dff_A_EKEE6Tlo2_1),.clk(gclk));
	jdff dff_A_b7NjEgFW8_1(.dout(w_dff_A_EKEE6Tlo2_1),.din(w_dff_A_b7NjEgFW8_1),.clk(gclk));
	jdff dff_A_A9wfmooN6_1(.dout(w_dff_A_b7NjEgFW8_1),.din(w_dff_A_A9wfmooN6_1),.clk(gclk));
	jdff dff_A_mTKAX2b75_1(.dout(w_dff_A_A9wfmooN6_1),.din(w_dff_A_mTKAX2b75_1),.clk(gclk));
	jdff dff_A_Z0DGIgll9_1(.dout(w_dff_A_mTKAX2b75_1),.din(w_dff_A_Z0DGIgll9_1),.clk(gclk));
	jdff dff_A_Xxub7PmQ3_1(.dout(w_dff_A_Z0DGIgll9_1),.din(w_dff_A_Xxub7PmQ3_1),.clk(gclk));
	jdff dff_A_Pq2XUUwU2_1(.dout(w_dff_A_Xxub7PmQ3_1),.din(w_dff_A_Pq2XUUwU2_1),.clk(gclk));
	jdff dff_A_jcUCBrq45_1(.dout(w_dff_A_Pq2XUUwU2_1),.din(w_dff_A_jcUCBrq45_1),.clk(gclk));
	jdff dff_A_dkolpX118_1(.dout(w_dff_A_jcUCBrq45_1),.din(w_dff_A_dkolpX118_1),.clk(gclk));
	jdff dff_A_njsPvHKF3_1(.dout(w_dff_A_dkolpX118_1),.din(w_dff_A_njsPvHKF3_1),.clk(gclk));
	jdff dff_A_hbAV5I5r2_1(.dout(w_dff_A_njsPvHKF3_1),.din(w_dff_A_hbAV5I5r2_1),.clk(gclk));
	jdff dff_A_RhSNtQ7o7_1(.dout(w_dff_A_hbAV5I5r2_1),.din(w_dff_A_RhSNtQ7o7_1),.clk(gclk));
	jdff dff_A_vHpQMJM47_1(.dout(w_dff_A_RhSNtQ7o7_1),.din(w_dff_A_vHpQMJM47_1),.clk(gclk));
	jdff dff_A_Apmk8SeQ1_1(.dout(w_dff_A_vHpQMJM47_1),.din(w_dff_A_Apmk8SeQ1_1),.clk(gclk));
	jdff dff_A_BhdubKHE1_1(.dout(w_dff_A_Apmk8SeQ1_1),.din(w_dff_A_BhdubKHE1_1),.clk(gclk));
	jdff dff_A_5xjHTlCY6_1(.dout(w_dff_A_BhdubKHE1_1),.din(w_dff_A_5xjHTlCY6_1),.clk(gclk));
	jdff dff_A_nsaHze9V0_1(.dout(w_dff_A_5xjHTlCY6_1),.din(w_dff_A_nsaHze9V0_1),.clk(gclk));
	jdff dff_B_bZf3Y5AV4_0(.din(G216),.dout(w_dff_B_bZf3Y5AV4_0),.clk(gclk));
	jdff dff_A_rOTyxRsQ1_0(.dout(w_n393_0[0]),.din(w_dff_A_rOTyxRsQ1_0),.clk(gclk));
	jdff dff_A_BBzGkKiJ5_0(.dout(w_dff_A_rOTyxRsQ1_0),.din(w_dff_A_BBzGkKiJ5_0),.clk(gclk));
	jdff dff_A_ueWiOO963_1(.dout(w_n393_0[1]),.din(w_dff_A_ueWiOO963_1),.clk(gclk));
	jdff dff_A_oj1IjktD9_1(.dout(w_dff_A_ueWiOO963_1),.din(w_dff_A_oj1IjktD9_1),.clk(gclk));
	jdff dff_A_MChL85tW9_0(.dout(w_n392_0[0]),.din(w_dff_A_MChL85tW9_0),.clk(gclk));
	jdff dff_A_XMXSjf4L9_0(.dout(w_dff_A_MChL85tW9_0),.din(w_dff_A_XMXSjf4L9_0),.clk(gclk));
	jdff dff_A_UyLnJLpV5_0(.dout(w_dff_A_XMXSjf4L9_0),.din(w_dff_A_UyLnJLpV5_0),.clk(gclk));
	jdff dff_A_XvxZdTNf7_0(.dout(w_dff_A_UyLnJLpV5_0),.din(w_dff_A_XvxZdTNf7_0),.clk(gclk));
	jdff dff_A_wx8BE9BM7_0(.dout(w_dff_A_XvxZdTNf7_0),.din(w_dff_A_wx8BE9BM7_0),.clk(gclk));
	jdff dff_B_SYp4AUKk5_2(.din(G209),.dout(w_dff_B_SYp4AUKk5_2),.clk(gclk));
	jdff dff_A_5XFw2BK36_0(.dout(w_n389_0[0]),.din(w_dff_A_5XFw2BK36_0),.clk(gclk));
	jdff dff_A_qqy3ED7z2_0(.dout(w_dff_A_5XFw2BK36_0),.din(w_dff_A_qqy3ED7z2_0),.clk(gclk));
	jdff dff_A_GpfuqmSP6_1(.dout(w_n389_0[1]),.din(w_dff_A_GpfuqmSP6_1),.clk(gclk));
	jdff dff_A_JXnlarNW9_1(.dout(w_dff_A_GpfuqmSP6_1),.din(w_dff_A_JXnlarNW9_1),.clk(gclk));
	jdff dff_A_j3rjMdM79_0(.dout(w_n388_1[0]),.din(w_dff_A_j3rjMdM79_0),.clk(gclk));
	jdff dff_A_SRJSWJeu4_2(.dout(w_n388_1[2]),.din(w_dff_A_SRJSWJeu4_2),.clk(gclk));
	jdff dff_A_vKP5qq0L8_0(.dout(w_n377_0[0]),.din(w_dff_A_vKP5qq0L8_0),.clk(gclk));
	jdff dff_A_t6sCCjTH2_0(.dout(w_dff_A_vKP5qq0L8_0),.din(w_dff_A_t6sCCjTH2_0),.clk(gclk));
	jdff dff_A_p5p2AGaa0_2(.dout(w_n377_0[2]),.din(w_dff_A_p5p2AGaa0_2),.clk(gclk));
	jdff dff_A_zbGCICaN3_2(.dout(w_dff_A_p5p2AGaa0_2),.din(w_dff_A_zbGCICaN3_2),.clk(gclk));
	jdff dff_A_eO1qbKxK0_2(.dout(w_dff_A_zbGCICaN3_2),.din(w_dff_A_eO1qbKxK0_2),.clk(gclk));
	jdff dff_A_bSvOCi7B0_2(.dout(w_dff_A_eO1qbKxK0_2),.din(w_dff_A_bSvOCi7B0_2),.clk(gclk));
	jdff dff_A_TP1DRJpF5_2(.dout(w_dff_A_bSvOCi7B0_2),.din(w_dff_A_TP1DRJpF5_2),.clk(gclk));
	jdff dff_A_zxZQCvQJ6_2(.dout(w_dff_A_TP1DRJpF5_2),.din(w_dff_A_zxZQCvQJ6_2),.clk(gclk));
	jdff dff_A_idthlT9g4_2(.dout(w_dff_A_zxZQCvQJ6_2),.din(w_dff_A_idthlT9g4_2),.clk(gclk));
	jdff dff_A_kjpjMtHF4_0(.dout(w_n374_0[0]),.din(w_dff_A_kjpjMtHF4_0),.clk(gclk));
	jdff dff_A_tkqNoS2v5_0(.dout(w_dff_A_kjpjMtHF4_0),.din(w_dff_A_tkqNoS2v5_0),.clk(gclk));
	jdff dff_B_a909KlhV4_0(.din(G213),.dout(w_dff_B_a909KlhV4_0),.clk(gclk));
	jdff dff_A_X1TuwsZf3_1(.dout(w_n371_0[1]),.din(w_dff_A_X1TuwsZf3_1),.clk(gclk));
	jdff dff_A_nuxPCBOz4_1(.dout(w_dff_A_X1TuwsZf3_1),.din(w_dff_A_nuxPCBOz4_1),.clk(gclk));
	jdff dff_A_FM3mH6a44_2(.dout(w_n371_0[2]),.din(w_dff_A_FM3mH6a44_2),.clk(gclk));
	jdff dff_A_fWSAdVKo6_2(.dout(w_dff_A_FM3mH6a44_2),.din(w_dff_A_fWSAdVKo6_2),.clk(gclk));
	jdff dff_B_dxI4Drpe8_1(.din(n508),.dout(w_dff_B_dxI4Drpe8_1),.clk(gclk));
	jdff dff_B_pmThCi3D0_1(.din(w_dff_B_dxI4Drpe8_1),.dout(w_dff_B_pmThCi3D0_1),.clk(gclk));
	jdff dff_B_iAKDS9Hl0_1(.din(w_dff_B_pmThCi3D0_1),.dout(w_dff_B_iAKDS9Hl0_1),.clk(gclk));
	jdff dff_B_fLkGQpSK7_1(.din(w_dff_B_iAKDS9Hl0_1),.dout(w_dff_B_fLkGQpSK7_1),.clk(gclk));
	jdff dff_B_ouyj905a4_1(.din(w_dff_B_fLkGQpSK7_1),.dout(w_dff_B_ouyj905a4_1),.clk(gclk));
	jdff dff_B_wsYh0W1j6_1(.din(w_dff_B_ouyj905a4_1),.dout(w_dff_B_wsYh0W1j6_1),.clk(gclk));
	jdff dff_B_s7kfYvyR7_1(.din(w_dff_B_wsYh0W1j6_1),.dout(w_dff_B_s7kfYvyR7_1),.clk(gclk));
	jdff dff_B_djipIL9X3_1(.din(w_dff_B_s7kfYvyR7_1),.dout(w_dff_B_djipIL9X3_1),.clk(gclk));
	jdff dff_B_HaqvBl8E4_1(.din(w_dff_B_djipIL9X3_1),.dout(w_dff_B_HaqvBl8E4_1),.clk(gclk));
	jdff dff_B_3wgKmfbH2_1(.din(w_dff_B_HaqvBl8E4_1),.dout(w_dff_B_3wgKmfbH2_1),.clk(gclk));
	jdff dff_B_g1HA1iMZ8_1(.din(w_dff_B_3wgKmfbH2_1),.dout(w_dff_B_g1HA1iMZ8_1),.clk(gclk));
	jdff dff_B_hV6BjzUi4_1(.din(w_dff_B_g1HA1iMZ8_1),.dout(w_dff_B_hV6BjzUi4_1),.clk(gclk));
	jdff dff_B_gLD3NANP0_1(.din(w_dff_B_hV6BjzUi4_1),.dout(w_dff_B_gLD3NANP0_1),.clk(gclk));
	jdff dff_B_6uYLmdzp6_1(.din(w_dff_B_gLD3NANP0_1),.dout(w_dff_B_6uYLmdzp6_1),.clk(gclk));
	jdff dff_B_1XOwPlP90_1(.din(w_dff_B_6uYLmdzp6_1),.dout(w_dff_B_1XOwPlP90_1),.clk(gclk));
	jdff dff_B_jhN7ONri7_1(.din(w_dff_B_1XOwPlP90_1),.dout(w_dff_B_jhN7ONri7_1),.clk(gclk));
	jdff dff_B_jQqlgt9b9_1(.din(w_dff_B_jhN7ONri7_1),.dout(w_dff_B_jQqlgt9b9_1),.clk(gclk));
	jdff dff_B_eOrW3sMd4_1(.din(w_dff_B_jQqlgt9b9_1),.dout(w_dff_B_eOrW3sMd4_1),.clk(gclk));
	jdff dff_B_ivJcWUpd4_1(.din(w_dff_B_eOrW3sMd4_1),.dout(w_dff_B_ivJcWUpd4_1),.clk(gclk));
	jdff dff_B_A9ljM3pL5_0(.din(n697),.dout(w_dff_B_A9ljM3pL5_0),.clk(gclk));
	jdff dff_B_vWTXuyzV1_0(.din(w_dff_B_A9ljM3pL5_0),.dout(w_dff_B_vWTXuyzV1_0),.clk(gclk));
	jdff dff_B_gFmnUpz72_0(.din(w_dff_B_vWTXuyzV1_0),.dout(w_dff_B_gFmnUpz72_0),.clk(gclk));
	jdff dff_B_5hs3d9dS8_0(.din(w_dff_B_gFmnUpz72_0),.dout(w_dff_B_5hs3d9dS8_0),.clk(gclk));
	jdff dff_B_glKRk3gR5_0(.din(w_dff_B_5hs3d9dS8_0),.dout(w_dff_B_glKRk3gR5_0),.clk(gclk));
	jdff dff_B_9rtOB0Lq3_0(.din(w_dff_B_glKRk3gR5_0),.dout(w_dff_B_9rtOB0Lq3_0),.clk(gclk));
	jdff dff_B_3yjIZrto9_0(.din(w_dff_B_9rtOB0Lq3_0),.dout(w_dff_B_3yjIZrto9_0),.clk(gclk));
	jdff dff_B_O2veVFGl5_0(.din(w_dff_B_3yjIZrto9_0),.dout(w_dff_B_O2veVFGl5_0),.clk(gclk));
	jdff dff_B_7TVa7QrY6_0(.din(w_dff_B_O2veVFGl5_0),.dout(w_dff_B_7TVa7QrY6_0),.clk(gclk));
	jdff dff_B_sagEw58q7_0(.din(w_dff_B_7TVa7QrY6_0),.dout(w_dff_B_sagEw58q7_0),.clk(gclk));
	jdff dff_B_c6HAdUaN2_0(.din(w_dff_B_sagEw58q7_0),.dout(w_dff_B_c6HAdUaN2_0),.clk(gclk));
	jdff dff_B_lAEfoLb51_0(.din(w_dff_B_c6HAdUaN2_0),.dout(w_dff_B_lAEfoLb51_0),.clk(gclk));
	jdff dff_B_n6A6nBpW3_0(.din(w_dff_B_lAEfoLb51_0),.dout(w_dff_B_n6A6nBpW3_0),.clk(gclk));
	jdff dff_B_pce0MwIA2_0(.din(w_dff_B_n6A6nBpW3_0),.dout(w_dff_B_pce0MwIA2_0),.clk(gclk));
	jdff dff_A_I7xDzB0S6_0(.dout(w_n696_0[0]),.din(w_dff_A_I7xDzB0S6_0),.clk(gclk));
	jdff dff_A_cNv0txgm3_0(.dout(w_dff_A_I7xDzB0S6_0),.din(w_dff_A_cNv0txgm3_0),.clk(gclk));
	jdff dff_A_aoVUsHNH4_0(.dout(w_dff_A_cNv0txgm3_0),.din(w_dff_A_aoVUsHNH4_0),.clk(gclk));
	jdff dff_A_uMMjXF7A7_0(.dout(w_dff_A_aoVUsHNH4_0),.din(w_dff_A_uMMjXF7A7_0),.clk(gclk));
	jdff dff_A_jRglSfii3_0(.dout(w_dff_A_uMMjXF7A7_0),.din(w_dff_A_jRglSfii3_0),.clk(gclk));
	jdff dff_A_5hsSyzRu8_0(.dout(w_dff_A_jRglSfii3_0),.din(w_dff_A_5hsSyzRu8_0),.clk(gclk));
	jdff dff_A_aXu3DKeP5_0(.dout(w_dff_A_5hsSyzRu8_0),.din(w_dff_A_aXu3DKeP5_0),.clk(gclk));
	jdff dff_A_nmfzxFhA3_0(.dout(w_dff_A_aXu3DKeP5_0),.din(w_dff_A_nmfzxFhA3_0),.clk(gclk));
	jdff dff_A_USPKJ8132_0(.dout(w_dff_A_nmfzxFhA3_0),.din(w_dff_A_USPKJ8132_0),.clk(gclk));
	jdff dff_A_X2pZoTDj5_0(.dout(w_dff_A_USPKJ8132_0),.din(w_dff_A_X2pZoTDj5_0),.clk(gclk));
	jdff dff_A_f4xdTZ1k0_0(.dout(w_dff_A_X2pZoTDj5_0),.din(w_dff_A_f4xdTZ1k0_0),.clk(gclk));
	jdff dff_A_Rszs5hxt9_0(.dout(w_dff_A_f4xdTZ1k0_0),.din(w_dff_A_Rszs5hxt9_0),.clk(gclk));
	jdff dff_A_0C7stwN52_0(.dout(w_dff_A_Rszs5hxt9_0),.din(w_dff_A_0C7stwN52_0),.clk(gclk));
	jdff dff_A_JicpSNRF3_0(.dout(w_dff_A_0C7stwN52_0),.din(w_dff_A_JicpSNRF3_0),.clk(gclk));
	jdff dff_A_b1VtYyyq2_0(.dout(w_dff_A_JicpSNRF3_0),.din(w_dff_A_b1VtYyyq2_0),.clk(gclk));
	jdff dff_B_4l6EjjZ92_1(.din(n688),.dout(w_dff_B_4l6EjjZ92_1),.clk(gclk));
	jdff dff_B_4mONRwjK5_1(.din(w_dff_B_4l6EjjZ92_1),.dout(w_dff_B_4mONRwjK5_1),.clk(gclk));
	jdff dff_B_2OvdcqoQ8_1(.din(w_dff_B_4mONRwjK5_1),.dout(w_dff_B_2OvdcqoQ8_1),.clk(gclk));
	jdff dff_B_tWHvgilG5_1(.din(n519),.dout(w_dff_B_tWHvgilG5_1),.clk(gclk));
	jdff dff_B_j3c8LBmL0_1(.din(w_dff_B_tWHvgilG5_1),.dout(w_dff_B_j3c8LBmL0_1),.clk(gclk));
	jdff dff_B_NRkqAHc08_1(.din(w_dff_B_j3c8LBmL0_1),.dout(w_dff_B_NRkqAHc08_1),.clk(gclk));
	jdff dff_B_UU5OWMm29_1(.din(w_dff_B_NRkqAHc08_1),.dout(w_dff_B_UU5OWMm29_1),.clk(gclk));
	jdff dff_B_FF9BiwNp5_1(.din(w_dff_B_UU5OWMm29_1),.dout(w_dff_B_FF9BiwNp5_1),.clk(gclk));
	jdff dff_B_ydLvFe607_1(.din(w_dff_B_FF9BiwNp5_1),.dout(w_dff_B_ydLvFe607_1),.clk(gclk));
	jdff dff_B_OaK0ATQs6_1(.din(w_dff_B_ydLvFe607_1),.dout(w_dff_B_OaK0ATQs6_1),.clk(gclk));
	jdff dff_B_BkLkavyk7_1(.din(w_dff_B_OaK0ATQs6_1),.dout(w_dff_B_BkLkavyk7_1),.clk(gclk));
	jdff dff_B_xt3rlacS3_1(.din(w_dff_B_BkLkavyk7_1),.dout(w_dff_B_xt3rlacS3_1),.clk(gclk));
	jdff dff_B_Nb90LzJ29_1(.din(w_dff_B_xt3rlacS3_1),.dout(w_dff_B_Nb90LzJ29_1),.clk(gclk));
	jdff dff_B_xEI4AJRJ0_1(.din(w_dff_B_Nb90LzJ29_1),.dout(w_dff_B_xEI4AJRJ0_1),.clk(gclk));
	jdff dff_B_BuNIFx2m3_1(.din(w_dff_B_xEI4AJRJ0_1),.dout(w_dff_B_BuNIFx2m3_1),.clk(gclk));
	jdff dff_B_uwJGeuQo2_1(.din(w_dff_B_BuNIFx2m3_1),.dout(w_dff_B_uwJGeuQo2_1),.clk(gclk));
	jdff dff_B_fLrw1hNJ4_1(.din(w_dff_B_uwJGeuQo2_1),.dout(w_dff_B_fLrw1hNJ4_1),.clk(gclk));
	jdff dff_B_KpiQnyyo5_1(.din(w_dff_B_fLrw1hNJ4_1),.dout(w_dff_B_KpiQnyyo5_1),.clk(gclk));
	jdff dff_B_4YOywbhc6_1(.din(w_dff_B_KpiQnyyo5_1),.dout(w_dff_B_4YOywbhc6_1),.clk(gclk));
	jdff dff_B_pE2wBYNa4_1(.din(w_dff_B_4YOywbhc6_1),.dout(w_dff_B_pE2wBYNa4_1),.clk(gclk));
	jdff dff_B_ZCvoo7Hx9_1(.din(n527),.dout(w_dff_B_ZCvoo7Hx9_1),.clk(gclk));
	jdff dff_B_pW0r1VbN2_1(.din(w_dff_B_ZCvoo7Hx9_1),.dout(w_dff_B_pW0r1VbN2_1),.clk(gclk));
	jdff dff_B_ZnnPsRxJ0_1(.din(w_dff_B_pW0r1VbN2_1),.dout(w_dff_B_ZnnPsRxJ0_1),.clk(gclk));
	jdff dff_B_MQNi7O0W7_1(.din(w_dff_B_ZnnPsRxJ0_1),.dout(w_dff_B_MQNi7O0W7_1),.clk(gclk));
	jdff dff_B_aoeJBiiz8_1(.din(w_dff_B_MQNi7O0W7_1),.dout(w_dff_B_aoeJBiiz8_1),.clk(gclk));
	jdff dff_B_P0hiPupE3_1(.din(w_dff_B_aoeJBiiz8_1),.dout(w_dff_B_P0hiPupE3_1),.clk(gclk));
	jdff dff_B_HR0JZQQm7_1(.din(w_dff_B_P0hiPupE3_1),.dout(w_dff_B_HR0JZQQm7_1),.clk(gclk));
	jdff dff_B_BPWMRp4e6_1(.din(w_dff_B_HR0JZQQm7_1),.dout(w_dff_B_BPWMRp4e6_1),.clk(gclk));
	jdff dff_B_hD6mkblq0_1(.din(w_dff_B_BPWMRp4e6_1),.dout(w_dff_B_hD6mkblq0_1),.clk(gclk));
	jdff dff_B_bOk8bYvH9_1(.din(w_dff_B_hD6mkblq0_1),.dout(w_dff_B_bOk8bYvH9_1),.clk(gclk));
	jdff dff_B_sBFOXOMN7_1(.din(w_dff_B_bOk8bYvH9_1),.dout(w_dff_B_sBFOXOMN7_1),.clk(gclk));
	jdff dff_B_vvQeQ9IZ6_1(.din(w_dff_B_sBFOXOMN7_1),.dout(w_dff_B_vvQeQ9IZ6_1),.clk(gclk));
	jdff dff_B_KrkYt20q1_1(.din(w_dff_B_vvQeQ9IZ6_1),.dout(w_dff_B_KrkYt20q1_1),.clk(gclk));
	jdff dff_B_qToOmZvf7_1(.din(w_dff_B_KrkYt20q1_1),.dout(w_dff_B_qToOmZvf7_1),.clk(gclk));
	jdff dff_A_4AY1VK1h7_1(.dout(w_n513_1[1]),.din(w_dff_A_4AY1VK1h7_1),.clk(gclk));
	jdff dff_A_OiCKnY8w5_1(.dout(w_dff_A_4AY1VK1h7_1),.din(w_dff_A_OiCKnY8w5_1),.clk(gclk));
	jdff dff_A_e0Ejqhux7_1(.dout(w_dff_A_OiCKnY8w5_1),.din(w_dff_A_e0Ejqhux7_1),.clk(gclk));
	jdff dff_A_5h6Q7F6G2_1(.dout(w_dff_A_e0Ejqhux7_1),.din(w_dff_A_5h6Q7F6G2_1),.clk(gclk));
	jdff dff_A_kBBqhWdO2_1(.dout(w_dff_A_5h6Q7F6G2_1),.din(w_dff_A_kBBqhWdO2_1),.clk(gclk));
	jdff dff_A_A1dL6dWk5_1(.dout(w_dff_A_kBBqhWdO2_1),.din(w_dff_A_A1dL6dWk5_1),.clk(gclk));
	jdff dff_A_n0BAAhXE8_1(.dout(w_dff_A_A1dL6dWk5_1),.din(w_dff_A_n0BAAhXE8_1),.clk(gclk));
	jdff dff_A_8vjMpDMc9_1(.dout(w_dff_A_n0BAAhXE8_1),.din(w_dff_A_8vjMpDMc9_1),.clk(gclk));
	jdff dff_A_F3FI9HFu1_1(.dout(w_dff_A_8vjMpDMc9_1),.din(w_dff_A_F3FI9HFu1_1),.clk(gclk));
	jdff dff_A_bUTvmJwf9_1(.dout(w_dff_A_F3FI9HFu1_1),.din(w_dff_A_bUTvmJwf9_1),.clk(gclk));
	jdff dff_A_W6Q6hwAB4_1(.dout(w_dff_A_bUTvmJwf9_1),.din(w_dff_A_W6Q6hwAB4_1),.clk(gclk));
	jdff dff_A_CcYGYwLY7_1(.dout(w_dff_A_W6Q6hwAB4_1),.din(w_dff_A_CcYGYwLY7_1),.clk(gclk));
	jdff dff_A_UGw49bNO0_1(.dout(w_dff_A_CcYGYwLY7_1),.din(w_dff_A_UGw49bNO0_1),.clk(gclk));
	jdff dff_A_elMZDeJw5_1(.dout(w_dff_A_UGw49bNO0_1),.din(w_dff_A_elMZDeJw5_1),.clk(gclk));
	jdff dff_A_IATSXNEX0_1(.dout(w_dff_A_elMZDeJw5_1),.din(w_dff_A_IATSXNEX0_1),.clk(gclk));
	jdff dff_A_7TcVFsax4_1(.dout(w_dff_A_IATSXNEX0_1),.din(w_dff_A_7TcVFsax4_1),.clk(gclk));
	jdff dff_A_YY9Wa9DR3_1(.dout(w_dff_A_7TcVFsax4_1),.din(w_dff_A_YY9Wa9DR3_1),.clk(gclk));
	jdff dff_A_wAQ3i3Jc9_1(.dout(w_dff_A_YY9Wa9DR3_1),.din(w_dff_A_wAQ3i3Jc9_1),.clk(gclk));
	jdff dff_A_6rMMNjas3_1(.dout(w_dff_A_wAQ3i3Jc9_1),.din(w_dff_A_6rMMNjas3_1),.clk(gclk));
	jdff dff_A_mysvAp8W3_0(.dout(w_n507_0[0]),.din(w_dff_A_mysvAp8W3_0),.clk(gclk));
	jdff dff_A_W2jLkjl70_0(.dout(w_dff_A_mysvAp8W3_0),.din(w_dff_A_W2jLkjl70_0),.clk(gclk));
	jdff dff_A_wBl7ND0M6_0(.dout(w_dff_A_W2jLkjl70_0),.din(w_dff_A_wBl7ND0M6_0),.clk(gclk));
	jdff dff_A_1kHYwltR7_0(.dout(w_dff_A_wBl7ND0M6_0),.din(w_dff_A_1kHYwltR7_0),.clk(gclk));
	jdff dff_A_wVENETGK6_0(.dout(w_dff_A_1kHYwltR7_0),.din(w_dff_A_wVENETGK6_0),.clk(gclk));
	jdff dff_A_9T32hcbM6_0(.dout(w_dff_A_wVENETGK6_0),.din(w_dff_A_9T32hcbM6_0),.clk(gclk));
	jdff dff_A_cIucq7oY5_0(.dout(w_dff_A_9T32hcbM6_0),.din(w_dff_A_cIucq7oY5_0),.clk(gclk));
	jdff dff_A_DIfLTP544_0(.dout(w_dff_A_cIucq7oY5_0),.din(w_dff_A_DIfLTP544_0),.clk(gclk));
	jdff dff_A_FEqIZsnq9_0(.dout(w_dff_A_DIfLTP544_0),.din(w_dff_A_FEqIZsnq9_0),.clk(gclk));
	jdff dff_A_EurOJcZ53_0(.dout(w_dff_A_FEqIZsnq9_0),.din(w_dff_A_EurOJcZ53_0),.clk(gclk));
	jdff dff_A_8oSIy0W82_0(.dout(w_dff_A_EurOJcZ53_0),.din(w_dff_A_8oSIy0W82_0),.clk(gclk));
	jdff dff_A_4nbLLgR66_0(.dout(w_dff_A_8oSIy0W82_0),.din(w_dff_A_4nbLLgR66_0),.clk(gclk));
	jdff dff_A_N0awK1a70_0(.dout(w_dff_A_4nbLLgR66_0),.din(w_dff_A_N0awK1a70_0),.clk(gclk));
	jdff dff_A_hY21ZafV7_0(.dout(w_dff_A_N0awK1a70_0),.din(w_dff_A_hY21ZafV7_0),.clk(gclk));
	jdff dff_A_4jEY70Uv7_0(.dout(w_dff_A_hY21ZafV7_0),.din(w_dff_A_4jEY70Uv7_0),.clk(gclk));
	jdff dff_A_hVdWN37r8_0(.dout(w_dff_A_4jEY70Uv7_0),.din(w_dff_A_hVdWN37r8_0),.clk(gclk));
	jdff dff_A_bZG6rCt02_0(.dout(w_dff_A_hVdWN37r8_0),.din(w_dff_A_bZG6rCt02_0),.clk(gclk));
	jdff dff_A_j8Yyd3C18_0(.dout(w_dff_A_bZG6rCt02_0),.din(w_dff_A_j8Yyd3C18_0),.clk(gclk));
	jdff dff_A_TytrfGEn0_0(.dout(w_dff_A_j8Yyd3C18_0),.din(w_dff_A_TytrfGEn0_0),.clk(gclk));
	jdff dff_A_nQGtR75U2_0(.dout(w_dff_A_TytrfGEn0_0),.din(w_dff_A_nQGtR75U2_0),.clk(gclk));
	jdff dff_A_wXmX0e7m5_1(.dout(w_n505_0[1]),.din(w_dff_A_wXmX0e7m5_1),.clk(gclk));
	jdff dff_A_dhNvzuby7_1(.dout(w_dff_A_wXmX0e7m5_1),.din(w_dff_A_dhNvzuby7_1),.clk(gclk));
	jdff dff_A_DJqP3u7M2_1(.dout(w_dff_A_dhNvzuby7_1),.din(w_dff_A_DJqP3u7M2_1),.clk(gclk));
	jdff dff_A_7Fqir6Uc3_1(.dout(w_dff_A_DJqP3u7M2_1),.din(w_dff_A_7Fqir6Uc3_1),.clk(gclk));
	jdff dff_A_lRaNFEFP2_1(.dout(w_dff_A_7Fqir6Uc3_1),.din(w_dff_A_lRaNFEFP2_1),.clk(gclk));
	jdff dff_A_4lf6tUkl5_1(.dout(w_dff_A_lRaNFEFP2_1),.din(w_dff_A_4lf6tUkl5_1),.clk(gclk));
	jdff dff_A_xVpNistd5_1(.dout(w_dff_A_4lf6tUkl5_1),.din(w_dff_A_xVpNistd5_1),.clk(gclk));
	jdff dff_A_4Q0HkovC8_1(.dout(w_dff_A_xVpNistd5_1),.din(w_dff_A_4Q0HkovC8_1),.clk(gclk));
	jdff dff_A_05cVpLKY5_1(.dout(w_dff_A_4Q0HkovC8_1),.din(w_dff_A_05cVpLKY5_1),.clk(gclk));
	jdff dff_A_I3EHgkKR5_1(.dout(w_dff_A_05cVpLKY5_1),.din(w_dff_A_I3EHgkKR5_1),.clk(gclk));
	jdff dff_A_TDuqIGv35_1(.dout(w_dff_A_I3EHgkKR5_1),.din(w_dff_A_TDuqIGv35_1),.clk(gclk));
	jdff dff_A_H5Du67Uf9_1(.dout(w_dff_A_TDuqIGv35_1),.din(w_dff_A_H5Du67Uf9_1),.clk(gclk));
	jdff dff_A_4FXWiXsM1_1(.dout(w_dff_A_H5Du67Uf9_1),.din(w_dff_A_4FXWiXsM1_1),.clk(gclk));
	jdff dff_A_DavtVEpX0_1(.dout(w_dff_A_4FXWiXsM1_1),.din(w_dff_A_DavtVEpX0_1),.clk(gclk));
	jdff dff_A_Cfo0Ft2p4_1(.dout(w_dff_A_DavtVEpX0_1),.din(w_dff_A_Cfo0Ft2p4_1),.clk(gclk));
	jdff dff_A_92OGamdW0_1(.dout(w_dff_A_Cfo0Ft2p4_1),.din(w_dff_A_92OGamdW0_1),.clk(gclk));
	jdff dff_A_lUlKWWju8_1(.dout(w_dff_A_92OGamdW0_1),.din(w_dff_A_lUlKWWju8_1),.clk(gclk));
	jdff dff_A_IsUwWonB5_1(.dout(w_dff_A_lUlKWWju8_1),.din(w_dff_A_IsUwWonB5_1),.clk(gclk));
	jdff dff_A_ZAjNNJfD7_1(.dout(w_dff_A_IsUwWonB5_1),.din(w_dff_A_ZAjNNJfD7_1),.clk(gclk));
	jdff dff_A_1VSTvnbX6_1(.dout(w_dff_A_ZAjNNJfD7_1),.din(w_dff_A_1VSTvnbX6_1),.clk(gclk));
	jdff dff_A_gHh1LAwz8_1(.dout(w_dff_A_1VSTvnbX6_1),.din(w_dff_A_gHh1LAwz8_1),.clk(gclk));
	jdff dff_A_RxW72wH48_1(.dout(w_dff_A_gHh1LAwz8_1),.din(w_dff_A_RxW72wH48_1),.clk(gclk));
	jdff dff_A_pV3i2Oqw1_1(.dout(w_n500_0[1]),.din(w_dff_A_pV3i2Oqw1_1),.clk(gclk));
	jdff dff_A_rZ0hgTC95_1(.dout(w_dff_A_pV3i2Oqw1_1),.din(w_dff_A_rZ0hgTC95_1),.clk(gclk));
	jdff dff_A_hQTC4fE15_1(.dout(w_dff_A_rZ0hgTC95_1),.din(w_dff_A_hQTC4fE15_1),.clk(gclk));
	jdff dff_A_mslwNtHw0_1(.dout(w_dff_A_hQTC4fE15_1),.din(w_dff_A_mslwNtHw0_1),.clk(gclk));
	jdff dff_A_ijRyzMBZ9_1(.dout(w_dff_A_mslwNtHw0_1),.din(w_dff_A_ijRyzMBZ9_1),.clk(gclk));
	jdff dff_A_wlVkLV6h4_1(.dout(w_dff_A_ijRyzMBZ9_1),.din(w_dff_A_wlVkLV6h4_1),.clk(gclk));
	jdff dff_A_yWUIeNXJ3_1(.dout(w_dff_A_wlVkLV6h4_1),.din(w_dff_A_yWUIeNXJ3_1),.clk(gclk));
	jdff dff_A_pQb2xkDp4_1(.dout(w_dff_A_yWUIeNXJ3_1),.din(w_dff_A_pQb2xkDp4_1),.clk(gclk));
	jdff dff_A_8yZtTeNR1_1(.dout(w_dff_A_pQb2xkDp4_1),.din(w_dff_A_8yZtTeNR1_1),.clk(gclk));
	jdff dff_A_HSRsi5bl1_1(.dout(w_dff_A_8yZtTeNR1_1),.din(w_dff_A_HSRsi5bl1_1),.clk(gclk));
	jdff dff_A_cFUZ2Tor7_1(.dout(w_dff_A_HSRsi5bl1_1),.din(w_dff_A_cFUZ2Tor7_1),.clk(gclk));
	jdff dff_A_3YjeGyEk6_1(.dout(w_dff_A_cFUZ2Tor7_1),.din(w_dff_A_3YjeGyEk6_1),.clk(gclk));
	jdff dff_A_kodrTzqj5_1(.dout(w_dff_A_3YjeGyEk6_1),.din(w_dff_A_kodrTzqj5_1),.clk(gclk));
	jdff dff_A_lMCx3fHi1_1(.dout(w_dff_A_kodrTzqj5_1),.din(w_dff_A_lMCx3fHi1_1),.clk(gclk));
	jdff dff_A_ySDlUllu3_1(.dout(w_dff_A_lMCx3fHi1_1),.din(w_dff_A_ySDlUllu3_1),.clk(gclk));
	jdff dff_A_fNRZdPWU1_1(.dout(w_dff_A_ySDlUllu3_1),.din(w_dff_A_fNRZdPWU1_1),.clk(gclk));
	jdff dff_A_wmgdaXR69_1(.dout(w_dff_A_fNRZdPWU1_1),.din(w_dff_A_wmgdaXR69_1),.clk(gclk));
	jdff dff_A_AJ2RaLHq2_1(.dout(w_dff_A_wmgdaXR69_1),.din(w_dff_A_AJ2RaLHq2_1),.clk(gclk));
	jdff dff_A_ZHrf0Wum6_1(.dout(w_n499_0[1]),.din(w_dff_A_ZHrf0Wum6_1),.clk(gclk));
	jdff dff_A_tIa5nNvV2_1(.dout(w_dff_A_ZHrf0Wum6_1),.din(w_dff_A_tIa5nNvV2_1),.clk(gclk));
	jdff dff_A_g1XOuA2k6_1(.dout(w_dff_A_tIa5nNvV2_1),.din(w_dff_A_g1XOuA2k6_1),.clk(gclk));
	jdff dff_A_5RRLB7Y64_1(.dout(w_dff_A_g1XOuA2k6_1),.din(w_dff_A_5RRLB7Y64_1),.clk(gclk));
	jdff dff_A_CpQPaSC28_1(.dout(w_dff_A_5RRLB7Y64_1),.din(w_dff_A_CpQPaSC28_1),.clk(gclk));
	jdff dff_A_BTgskNrm5_1(.dout(w_dff_A_CpQPaSC28_1),.din(w_dff_A_BTgskNrm5_1),.clk(gclk));
	jdff dff_A_4IMIwSgI0_1(.dout(w_dff_A_BTgskNrm5_1),.din(w_dff_A_4IMIwSgI0_1),.clk(gclk));
	jdff dff_A_8XtrJMHW8_1(.dout(w_dff_A_4IMIwSgI0_1),.din(w_dff_A_8XtrJMHW8_1),.clk(gclk));
	jdff dff_A_FXU8MAlH3_1(.dout(w_dff_A_8XtrJMHW8_1),.din(w_dff_A_FXU8MAlH3_1),.clk(gclk));
	jdff dff_A_pfxgqJCX4_1(.dout(w_dff_A_FXU8MAlH3_1),.din(w_dff_A_pfxgqJCX4_1),.clk(gclk));
	jdff dff_A_nNkPY3zj6_1(.dout(w_dff_A_pfxgqJCX4_1),.din(w_dff_A_nNkPY3zj6_1),.clk(gclk));
	jdff dff_A_2CeUZ8G02_1(.dout(w_dff_A_nNkPY3zj6_1),.din(w_dff_A_2CeUZ8G02_1),.clk(gclk));
	jdff dff_A_mRi2UOy46_1(.dout(w_dff_A_2CeUZ8G02_1),.din(w_dff_A_mRi2UOy46_1),.clk(gclk));
	jdff dff_A_bxcvZCMb8_1(.dout(w_dff_A_mRi2UOy46_1),.din(w_dff_A_bxcvZCMb8_1),.clk(gclk));
	jdff dff_A_ELfkE1sR4_1(.dout(w_dff_A_bxcvZCMb8_1),.din(w_dff_A_ELfkE1sR4_1),.clk(gclk));
	jdff dff_A_SzNhROO54_1(.dout(w_dff_A_ELfkE1sR4_1),.din(w_dff_A_SzNhROO54_1),.clk(gclk));
	jdff dff_A_YKcXgaSB9_1(.dout(w_dff_A_SzNhROO54_1),.din(w_dff_A_YKcXgaSB9_1),.clk(gclk));
	jdff dff_A_2h3sDGq20_0(.dout(w_n497_1[0]),.din(w_dff_A_2h3sDGq20_0),.clk(gclk));
	jdff dff_A_xQp4L2oT1_0(.dout(w_dff_A_2h3sDGq20_0),.din(w_dff_A_xQp4L2oT1_0),.clk(gclk));
	jdff dff_A_lP7LBitw2_0(.dout(w_dff_A_xQp4L2oT1_0),.din(w_dff_A_lP7LBitw2_0),.clk(gclk));
	jdff dff_A_NeiOiegw4_0(.dout(w_dff_A_lP7LBitw2_0),.din(w_dff_A_NeiOiegw4_0),.clk(gclk));
	jdff dff_A_YCAS7qFR3_0(.dout(w_dff_A_NeiOiegw4_0),.din(w_dff_A_YCAS7qFR3_0),.clk(gclk));
	jdff dff_A_aVVmcqqy9_0(.dout(w_dff_A_YCAS7qFR3_0),.din(w_dff_A_aVVmcqqy9_0),.clk(gclk));
	jdff dff_A_xqJnR9AY2_0(.dout(w_dff_A_aVVmcqqy9_0),.din(w_dff_A_xqJnR9AY2_0),.clk(gclk));
	jdff dff_A_5pBWwoNE3_0(.dout(w_dff_A_xqJnR9AY2_0),.din(w_dff_A_5pBWwoNE3_0),.clk(gclk));
	jdff dff_A_3Y0zYfS50_0(.dout(w_dff_A_5pBWwoNE3_0),.din(w_dff_A_3Y0zYfS50_0),.clk(gclk));
	jdff dff_A_QA8uoGzG6_0(.dout(w_dff_A_3Y0zYfS50_0),.din(w_dff_A_QA8uoGzG6_0),.clk(gclk));
	jdff dff_A_Ei0Pduxf5_0(.dout(w_dff_A_QA8uoGzG6_0),.din(w_dff_A_Ei0Pduxf5_0),.clk(gclk));
	jdff dff_A_AzQzgRyV6_0(.dout(w_dff_A_Ei0Pduxf5_0),.din(w_dff_A_AzQzgRyV6_0),.clk(gclk));
	jdff dff_A_tVVeXCWX9_0(.dout(w_dff_A_AzQzgRyV6_0),.din(w_dff_A_tVVeXCWX9_0),.clk(gclk));
	jdff dff_A_M04ERNrn8_0(.dout(w_dff_A_tVVeXCWX9_0),.din(w_dff_A_M04ERNrn8_0),.clk(gclk));
	jdff dff_A_DURmX0lG4_0(.dout(w_dff_A_M04ERNrn8_0),.din(w_dff_A_DURmX0lG4_0),.clk(gclk));
	jdff dff_A_HshRxNag0_0(.dout(w_dff_A_DURmX0lG4_0),.din(w_dff_A_HshRxNag0_0),.clk(gclk));
	jdff dff_A_qnv7e2B19_0(.dout(w_dff_A_HshRxNag0_0),.din(w_dff_A_qnv7e2B19_0),.clk(gclk));
	jdff dff_A_M68AdHPb8_0(.dout(w_dff_A_qnv7e2B19_0),.din(w_dff_A_M68AdHPb8_0),.clk(gclk));
	jdff dff_A_IHcVICTS5_0(.dout(w_dff_A_M68AdHPb8_0),.din(w_dff_A_IHcVICTS5_0),.clk(gclk));
	jdff dff_B_tus5eRkm1_1(.din(n482),.dout(w_dff_B_tus5eRkm1_1),.clk(gclk));
	jdff dff_B_eAXF9DqD6_1(.din(w_dff_B_tus5eRkm1_1),.dout(w_dff_B_eAXF9DqD6_1),.clk(gclk));
	jdff dff_B_gyQ2zbRa9_1(.din(w_dff_B_eAXF9DqD6_1),.dout(w_dff_B_gyQ2zbRa9_1),.clk(gclk));
	jdff dff_A_tuc5fw9a7_0(.dout(w_n495_1[0]),.din(w_dff_A_tuc5fw9a7_0),.clk(gclk));
	jdff dff_A_IS805HAQ7_0(.dout(w_dff_A_tuc5fw9a7_0),.din(w_dff_A_IS805HAQ7_0),.clk(gclk));
	jdff dff_A_UFxIPcbP1_0(.dout(w_dff_A_IS805HAQ7_0),.din(w_dff_A_UFxIPcbP1_0),.clk(gclk));
	jdff dff_A_yetBByJb6_0(.dout(w_dff_A_UFxIPcbP1_0),.din(w_dff_A_yetBByJb6_0),.clk(gclk));
	jdff dff_A_ZQPQV9Ht5_0(.dout(w_dff_A_yetBByJb6_0),.din(w_dff_A_ZQPQV9Ht5_0),.clk(gclk));
	jdff dff_A_fDVTvTrs4_0(.dout(w_dff_A_ZQPQV9Ht5_0),.din(w_dff_A_fDVTvTrs4_0),.clk(gclk));
	jdff dff_A_LR0mbwcR8_0(.dout(w_dff_A_fDVTvTrs4_0),.din(w_dff_A_LR0mbwcR8_0),.clk(gclk));
	jdff dff_A_WnKG3TWf8_0(.dout(w_dff_A_LR0mbwcR8_0),.din(w_dff_A_WnKG3TWf8_0),.clk(gclk));
	jdff dff_A_x4xG804r2_0(.dout(w_dff_A_WnKG3TWf8_0),.din(w_dff_A_x4xG804r2_0),.clk(gclk));
	jdff dff_A_rXbJPyvP6_0(.dout(w_dff_A_x4xG804r2_0),.din(w_dff_A_rXbJPyvP6_0),.clk(gclk));
	jdff dff_A_YUovUFfc3_0(.dout(w_dff_A_rXbJPyvP6_0),.din(w_dff_A_YUovUFfc3_0),.clk(gclk));
	jdff dff_A_oDpyawyB1_0(.dout(w_dff_A_YUovUFfc3_0),.din(w_dff_A_oDpyawyB1_0),.clk(gclk));
	jdff dff_A_J66xRmJJ2_0(.dout(w_dff_A_oDpyawyB1_0),.din(w_dff_A_J66xRmJJ2_0),.clk(gclk));
	jdff dff_A_bvfMJeKd6_0(.dout(w_dff_A_J66xRmJJ2_0),.din(w_dff_A_bvfMJeKd6_0),.clk(gclk));
	jdff dff_A_qbs6oP5o0_0(.dout(w_dff_A_bvfMJeKd6_0),.din(w_dff_A_qbs6oP5o0_0),.clk(gclk));
	jdff dff_A_mMtwPRWV7_0(.dout(w_dff_A_qbs6oP5o0_0),.din(w_dff_A_mMtwPRWV7_0),.clk(gclk));
	jdff dff_A_9hRxczGh1_0(.dout(w_dff_A_mMtwPRWV7_0),.din(w_dff_A_9hRxczGh1_0),.clk(gclk));
	jdff dff_A_2OlbOgEd7_0(.dout(w_dff_A_9hRxczGh1_0),.din(w_dff_A_2OlbOgEd7_0),.clk(gclk));
	jdff dff_A_U03xe2o77_0(.dout(w_dff_A_2OlbOgEd7_0),.din(w_dff_A_U03xe2o77_0),.clk(gclk));
	jdff dff_B_Yv1yDio26_1(.din(n484),.dout(w_dff_B_Yv1yDio26_1),.clk(gclk));
	jdff dff_B_GMRm2J0a2_1(.din(w_dff_B_Yv1yDio26_1),.dout(w_dff_B_GMRm2J0a2_1),.clk(gclk));
	jdff dff_A_DgLoT3Cl6_0(.dout(w_n491_1[0]),.din(w_dff_A_DgLoT3Cl6_0),.clk(gclk));
	jdff dff_A_EeUnnpzw5_0(.dout(w_dff_A_DgLoT3Cl6_0),.din(w_dff_A_EeUnnpzw5_0),.clk(gclk));
	jdff dff_A_heQPLmxD8_0(.dout(w_dff_A_EeUnnpzw5_0),.din(w_dff_A_heQPLmxD8_0),.clk(gclk));
	jdff dff_A_HhlvpK5i5_2(.dout(w_n491_0[2]),.din(w_dff_A_HhlvpK5i5_2),.clk(gclk));
	jdff dff_A_8J2edwd05_2(.dout(w_dff_A_HhlvpK5i5_2),.din(w_dff_A_8J2edwd05_2),.clk(gclk));
	jdff dff_A_wEhkXbVQ8_1(.dout(w_n487_0[1]),.din(w_dff_A_wEhkXbVQ8_1),.clk(gclk));
	jdff dff_A_hoEmSdRR5_1(.dout(w_dff_A_wEhkXbVQ8_1),.din(w_dff_A_hoEmSdRR5_1),.clk(gclk));
	jdff dff_A_Yqac6JF91_1(.dout(w_dff_A_hoEmSdRR5_1),.din(w_dff_A_Yqac6JF91_1),.clk(gclk));
	jdff dff_A_cQq5FWtM1_1(.dout(w_dff_A_Yqac6JF91_1),.din(w_dff_A_cQq5FWtM1_1),.clk(gclk));
	jdff dff_A_kkyJwqUr4_1(.dout(w_dff_A_cQq5FWtM1_1),.din(w_dff_A_kkyJwqUr4_1),.clk(gclk));
	jdff dff_A_MVluvxhh8_1(.dout(w_dff_A_kkyJwqUr4_1),.din(w_dff_A_MVluvxhh8_1),.clk(gclk));
	jdff dff_A_JqRgh5A39_1(.dout(w_dff_A_MVluvxhh8_1),.din(w_dff_A_JqRgh5A39_1),.clk(gclk));
	jdff dff_A_XAPlT4QL3_1(.dout(w_dff_A_JqRgh5A39_1),.din(w_dff_A_XAPlT4QL3_1),.clk(gclk));
	jdff dff_A_uH5x4HXz4_1(.dout(w_dff_A_XAPlT4QL3_1),.din(w_dff_A_uH5x4HXz4_1),.clk(gclk));
	jdff dff_A_JDkxCPk02_1(.dout(w_dff_A_uH5x4HXz4_1),.din(w_dff_A_JDkxCPk02_1),.clk(gclk));
	jdff dff_A_EU9PD6dJ6_1(.dout(w_dff_A_JDkxCPk02_1),.din(w_dff_A_EU9PD6dJ6_1),.clk(gclk));
	jdff dff_A_nlTJAkyk4_1(.dout(w_dff_A_EU9PD6dJ6_1),.din(w_dff_A_nlTJAkyk4_1),.clk(gclk));
	jdff dff_A_ihrt3K1E9_1(.dout(w_dff_A_nlTJAkyk4_1),.din(w_dff_A_ihrt3K1E9_1),.clk(gclk));
	jdff dff_A_Xijo1cgG4_1(.dout(w_dff_A_ihrt3K1E9_1),.din(w_dff_A_Xijo1cgG4_1),.clk(gclk));
	jdff dff_A_dkJWDnAp9_1(.dout(w_dff_A_Xijo1cgG4_1),.din(w_dff_A_dkJWDnAp9_1),.clk(gclk));
	jdff dff_A_28sMcNK85_1(.dout(w_dff_A_dkJWDnAp9_1),.din(w_dff_A_28sMcNK85_1),.clk(gclk));
	jdff dff_A_OMaqpi0d6_1(.dout(w_dff_A_28sMcNK85_1),.din(w_dff_A_OMaqpi0d6_1),.clk(gclk));
	jdff dff_A_j1cVR0RX7_1(.dout(w_dff_A_OMaqpi0d6_1),.din(w_dff_A_j1cVR0RX7_1),.clk(gclk));
	jdff dff_A_ks5Qe54q5_1(.dout(w_dff_A_j1cVR0RX7_1),.din(w_dff_A_ks5Qe54q5_1),.clk(gclk));
	jdff dff_A_4dWtdapo3_1(.dout(w_dff_A_ks5Qe54q5_1),.din(w_dff_A_4dWtdapo3_1),.clk(gclk));
	jdff dff_A_zpqqx4lL9_1(.dout(w_dff_A_4dWtdapo3_1),.din(w_dff_A_zpqqx4lL9_1),.clk(gclk));
	jdff dff_A_xLymxBEh4_1(.dout(w_dff_A_zpqqx4lL9_1),.din(w_dff_A_xLymxBEh4_1),.clk(gclk));
	jdff dff_A_FquwOoCd0_1(.dout(w_dff_A_xLymxBEh4_1),.din(w_dff_A_FquwOoCd0_1),.clk(gclk));
	jdff dff_A_JIc1SOCK2_1(.dout(w_dff_A_FquwOoCd0_1),.din(w_dff_A_JIc1SOCK2_1),.clk(gclk));
	jdff dff_A_GqDk9loR0_0(.dout(w_n481_0[0]),.din(w_dff_A_GqDk9loR0_0),.clk(gclk));
	jdff dff_A_4Le9nGDZ9_0(.dout(w_dff_A_GqDk9loR0_0),.din(w_dff_A_4Le9nGDZ9_0),.clk(gclk));
	jdff dff_A_OS89iIST8_0(.dout(w_dff_A_4Le9nGDZ9_0),.din(w_dff_A_OS89iIST8_0),.clk(gclk));
	jdff dff_A_MBUxQrmc6_0(.dout(w_dff_A_OS89iIST8_0),.din(w_dff_A_MBUxQrmc6_0),.clk(gclk));
	jdff dff_A_oFywIdMs1_0(.dout(w_dff_A_MBUxQrmc6_0),.din(w_dff_A_oFywIdMs1_0),.clk(gclk));
	jdff dff_A_GRSvb2ma3_0(.dout(w_dff_A_oFywIdMs1_0),.din(w_dff_A_GRSvb2ma3_0),.clk(gclk));
	jdff dff_A_VLOtDGPW1_0(.dout(w_dff_A_GRSvb2ma3_0),.din(w_dff_A_VLOtDGPW1_0),.clk(gclk));
	jdff dff_A_5ucflLL96_0(.dout(w_dff_A_VLOtDGPW1_0),.din(w_dff_A_5ucflLL96_0),.clk(gclk));
	jdff dff_A_zZEu0zwH3_0(.dout(w_dff_A_5ucflLL96_0),.din(w_dff_A_zZEu0zwH3_0),.clk(gclk));
	jdff dff_A_s0PqEE7h4_0(.dout(w_dff_A_zZEu0zwH3_0),.din(w_dff_A_s0PqEE7h4_0),.clk(gclk));
	jdff dff_A_bsGkyXTe7_0(.dout(w_dff_A_s0PqEE7h4_0),.din(w_dff_A_bsGkyXTe7_0),.clk(gclk));
	jdff dff_A_3b34rWmF2_0(.dout(w_dff_A_bsGkyXTe7_0),.din(w_dff_A_3b34rWmF2_0),.clk(gclk));
	jdff dff_A_zJq1VtZc4_0(.dout(w_dff_A_3b34rWmF2_0),.din(w_dff_A_zJq1VtZc4_0),.clk(gclk));
	jdff dff_A_66Rg3Y1y9_0(.dout(w_dff_A_zJq1VtZc4_0),.din(w_dff_A_66Rg3Y1y9_0),.clk(gclk));
	jdff dff_A_ScUGOy2X8_0(.dout(w_dff_A_66Rg3Y1y9_0),.din(w_dff_A_ScUGOy2X8_0),.clk(gclk));
	jdff dff_A_dKUNbawA1_0(.dout(w_dff_A_ScUGOy2X8_0),.din(w_dff_A_dKUNbawA1_0),.clk(gclk));
	jdff dff_A_a5IIealN0_0(.dout(w_dff_A_dKUNbawA1_0),.din(w_dff_A_a5IIealN0_0),.clk(gclk));
	jdff dff_A_uNdcLaJw2_0(.dout(w_dff_A_a5IIealN0_0),.din(w_dff_A_uNdcLaJw2_0),.clk(gclk));
	jdff dff_A_Nm6jfFKM7_0(.dout(w_dff_A_uNdcLaJw2_0),.din(w_dff_A_Nm6jfFKM7_0),.clk(gclk));
	jdff dff_A_ONH35l2Y7_0(.dout(w_dff_A_Nm6jfFKM7_0),.din(w_dff_A_ONH35l2Y7_0),.clk(gclk));
	jdff dff_A_99OCfEXo9_0(.dout(w_dff_A_ONH35l2Y7_0),.din(w_dff_A_99OCfEXo9_0),.clk(gclk));
	jdff dff_A_NTePZsvj2_0(.dout(w_dff_A_99OCfEXo9_0),.din(w_dff_A_NTePZsvj2_0),.clk(gclk));
	jdff dff_A_7x6e1Cwz1_2(.dout(w_n480_0[2]),.din(w_dff_A_7x6e1Cwz1_2),.clk(gclk));
	jdff dff_A_h0mCwTHF4_2(.dout(w_dff_A_7x6e1Cwz1_2),.din(w_dff_A_h0mCwTHF4_2),.clk(gclk));
	jdff dff_A_a2L6b9wV5_2(.dout(w_dff_A_h0mCwTHF4_2),.din(w_dff_A_a2L6b9wV5_2),.clk(gclk));
	jdff dff_A_RIidhpSp9_2(.dout(w_dff_A_a2L6b9wV5_2),.din(w_dff_A_RIidhpSp9_2),.clk(gclk));
	jdff dff_A_FUPkHfDt6_2(.dout(w_dff_A_RIidhpSp9_2),.din(w_dff_A_FUPkHfDt6_2),.clk(gclk));
	jdff dff_A_Z8wG2pGa3_2(.dout(w_dff_A_FUPkHfDt6_2),.din(w_dff_A_Z8wG2pGa3_2),.clk(gclk));
	jdff dff_A_3nBVnkpo2_2(.dout(w_dff_A_Z8wG2pGa3_2),.din(w_dff_A_3nBVnkpo2_2),.clk(gclk));
	jdff dff_A_y1aQQWlZ6_2(.dout(w_dff_A_3nBVnkpo2_2),.din(w_dff_A_y1aQQWlZ6_2),.clk(gclk));
	jdff dff_A_1vWIW1Rv9_2(.dout(w_dff_A_y1aQQWlZ6_2),.din(w_dff_A_1vWIW1Rv9_2),.clk(gclk));
	jdff dff_A_UpnmtUR61_2(.dout(w_dff_A_1vWIW1Rv9_2),.din(w_dff_A_UpnmtUR61_2),.clk(gclk));
	jdff dff_A_99gaBX5H7_2(.dout(w_dff_A_UpnmtUR61_2),.din(w_dff_A_99gaBX5H7_2),.clk(gclk));
	jdff dff_A_SJJq44Bw8_2(.dout(w_dff_A_99gaBX5H7_2),.din(w_dff_A_SJJq44Bw8_2),.clk(gclk));
	jdff dff_A_uc3cELp54_2(.dout(w_dff_A_SJJq44Bw8_2),.din(w_dff_A_uc3cELp54_2),.clk(gclk));
	jdff dff_A_s8lCTllk8_2(.dout(w_dff_A_uc3cELp54_2),.din(w_dff_A_s8lCTllk8_2),.clk(gclk));
	jdff dff_A_17Tjddwp7_2(.dout(w_dff_A_s8lCTllk8_2),.din(w_dff_A_17Tjddwp7_2),.clk(gclk));
	jdff dff_A_tNy0GlAU6_2(.dout(w_dff_A_17Tjddwp7_2),.din(w_dff_A_tNy0GlAU6_2),.clk(gclk));
	jdff dff_A_zr4HOGbH2_2(.dout(w_dff_A_tNy0GlAU6_2),.din(w_dff_A_zr4HOGbH2_2),.clk(gclk));
	jdff dff_A_zVRQU6PJ5_2(.dout(w_dff_A_zr4HOGbH2_2),.din(w_dff_A_zVRQU6PJ5_2),.clk(gclk));
	jdff dff_A_t0EtXzjT4_2(.dout(w_dff_A_zVRQU6PJ5_2),.din(w_dff_A_t0EtXzjT4_2),.clk(gclk));
	jdff dff_A_dymjYP6Y2_2(.dout(w_dff_A_t0EtXzjT4_2),.din(w_dff_A_dymjYP6Y2_2),.clk(gclk));
	jdff dff_A_E2nBjFEw2_2(.dout(w_dff_A_dymjYP6Y2_2),.din(w_dff_A_E2nBjFEw2_2),.clk(gclk));
	jdff dff_A_SKdSkvRK0_2(.dout(w_dff_A_E2nBjFEw2_2),.din(w_dff_A_SKdSkvRK0_2),.clk(gclk));
	jdff dff_A_oyn8YtEy2_2(.dout(w_dff_A_SKdSkvRK0_2),.din(w_dff_A_oyn8YtEy2_2),.clk(gclk));
	jdff dff_B_tvoDF4FO0_0(.din(n478),.dout(w_dff_B_tvoDF4FO0_0),.clk(gclk));
	jdff dff_B_0RG5tioS2_0(.din(G147),.dout(w_dff_B_0RG5tioS2_0),.clk(gclk));
	jdff dff_A_tpcB4Xpz7_1(.dout(w_n476_0[1]),.din(w_dff_A_tpcB4Xpz7_1),.clk(gclk));
	jdff dff_A_kyLWR7fF2_1(.dout(w_dff_A_tpcB4Xpz7_1),.din(w_dff_A_kyLWR7fF2_1),.clk(gclk));
	jdff dff_A_WCVFLqku1_2(.dout(w_n476_0[2]),.din(w_dff_A_WCVFLqku1_2),.clk(gclk));
	jdff dff_A_O9ZEuD0F3_2(.dout(w_dff_A_WCVFLqku1_2),.din(w_dff_A_O9ZEuD0F3_2),.clk(gclk));
	jdff dff_A_cxp9Ss3B8_1(.dout(w_G2211_0[1]),.din(w_dff_A_cxp9Ss3B8_1),.clk(gclk));
	jdff dff_A_M4kje5Xf9_1(.dout(w_dff_A_cxp9Ss3B8_1),.din(w_dff_A_M4kje5Xf9_1),.clk(gclk));
	jdff dff_A_6v2Rtka73_1(.dout(w_dff_A_M4kje5Xf9_1),.din(w_dff_A_6v2Rtka73_1),.clk(gclk));
	jdff dff_A_SR3YcPDr8_1(.dout(w_dff_A_6v2Rtka73_1),.din(w_dff_A_SR3YcPDr8_1),.clk(gclk));
	jdff dff_A_PFQbUgFH1_1(.dout(w_n475_0[1]),.din(w_dff_A_PFQbUgFH1_1),.clk(gclk));
	jdff dff_A_Th03vIP36_1(.dout(w_dff_A_PFQbUgFH1_1),.din(w_dff_A_Th03vIP36_1),.clk(gclk));
	jdff dff_A_ZKmtSBG20_1(.dout(w_dff_A_Th03vIP36_1),.din(w_dff_A_ZKmtSBG20_1),.clk(gclk));
	jdff dff_A_RkLwn8DP2_1(.dout(w_dff_A_ZKmtSBG20_1),.din(w_dff_A_RkLwn8DP2_1),.clk(gclk));
	jdff dff_A_TTpxHY2E4_1(.dout(w_dff_A_RkLwn8DP2_1),.din(w_dff_A_TTpxHY2E4_1),.clk(gclk));
	jdff dff_A_C2fZkQEP0_1(.dout(w_dff_A_TTpxHY2E4_1),.din(w_dff_A_C2fZkQEP0_1),.clk(gclk));
	jdff dff_A_0xmRz43N0_1(.dout(w_dff_A_C2fZkQEP0_1),.din(w_dff_A_0xmRz43N0_1),.clk(gclk));
	jdff dff_A_2RU396mk8_1(.dout(w_dff_A_0xmRz43N0_1),.din(w_dff_A_2RU396mk8_1),.clk(gclk));
	jdff dff_A_jNqaqBZC6_1(.dout(w_dff_A_2RU396mk8_1),.din(w_dff_A_jNqaqBZC6_1),.clk(gclk));
	jdff dff_A_jJlfJYnV6_1(.dout(w_dff_A_jNqaqBZC6_1),.din(w_dff_A_jJlfJYnV6_1),.clk(gclk));
	jdff dff_A_jN5FDuS95_1(.dout(w_dff_A_jJlfJYnV6_1),.din(w_dff_A_jN5FDuS95_1),.clk(gclk));
	jdff dff_A_nyXxN85x1_1(.dout(w_dff_A_jN5FDuS95_1),.din(w_dff_A_nyXxN85x1_1),.clk(gclk));
	jdff dff_A_EZt5qb8B7_1(.dout(w_dff_A_nyXxN85x1_1),.din(w_dff_A_EZt5qb8B7_1),.clk(gclk));
	jdff dff_A_7X9AVkNe8_1(.dout(w_dff_A_EZt5qb8B7_1),.din(w_dff_A_7X9AVkNe8_1),.clk(gclk));
	jdff dff_A_iQ8Yl5Ej1_1(.dout(w_dff_A_7X9AVkNe8_1),.din(w_dff_A_iQ8Yl5Ej1_1),.clk(gclk));
	jdff dff_A_ROcfoLcr4_1(.dout(w_dff_A_iQ8Yl5Ej1_1),.din(w_dff_A_ROcfoLcr4_1),.clk(gclk));
	jdff dff_A_vSmminsJ0_1(.dout(w_dff_A_ROcfoLcr4_1),.din(w_dff_A_vSmminsJ0_1),.clk(gclk));
	jdff dff_A_NUDMmJ1L5_1(.dout(w_dff_A_vSmminsJ0_1),.din(w_dff_A_NUDMmJ1L5_1),.clk(gclk));
	jdff dff_A_a5HHw5Zd5_1(.dout(w_dff_A_NUDMmJ1L5_1),.din(w_dff_A_a5HHw5Zd5_1),.clk(gclk));
	jdff dff_A_o38x5oMh6_1(.dout(w_dff_A_a5HHw5Zd5_1),.din(w_dff_A_o38x5oMh6_1),.clk(gclk));
	jdff dff_A_VmET2hKb8_1(.dout(w_dff_A_o38x5oMh6_1),.din(w_dff_A_VmET2hKb8_1),.clk(gclk));
	jdff dff_A_YNAHWE8k5_1(.dout(w_dff_A_VmET2hKb8_1),.din(w_dff_A_YNAHWE8k5_1),.clk(gclk));
	jdff dff_A_y5Wqknl02_1(.dout(w_dff_A_YNAHWE8k5_1),.din(w_dff_A_y5Wqknl02_1),.clk(gclk));
	jdff dff_A_UgbKSko40_1(.dout(w_dff_A_y5Wqknl02_1),.din(w_dff_A_UgbKSko40_1),.clk(gclk));
	jdff dff_A_mti1uzGy6_1(.dout(w_dff_A_UgbKSko40_1),.din(w_dff_A_mti1uzGy6_1),.clk(gclk));
	jdff dff_B_MQuA8mp51_0(.din(n473),.dout(w_dff_B_MQuA8mp51_0),.clk(gclk));
	jdff dff_B_i95EsnAB8_0(.din(G138),.dout(w_dff_B_i95EsnAB8_0),.clk(gclk));
	jdff dff_A_J2I59kpR2_1(.dout(w_n471_0[1]),.din(w_dff_A_J2I59kpR2_1),.clk(gclk));
	jdff dff_A_KfIMhN2W7_1(.dout(w_dff_A_J2I59kpR2_1),.din(w_dff_A_KfIMhN2W7_1),.clk(gclk));
	jdff dff_A_ZJQ3nsOw6_2(.dout(w_n471_0[2]),.din(w_dff_A_ZJQ3nsOw6_2),.clk(gclk));
	jdff dff_A_vtutKMai1_2(.dout(w_dff_A_ZJQ3nsOw6_2),.din(w_dff_A_vtutKMai1_2),.clk(gclk));
	jdff dff_A_sRfhcl926_1(.dout(w_G2218_0[1]),.din(w_dff_A_sRfhcl926_1),.clk(gclk));
	jdff dff_A_ihW1BRz73_1(.dout(w_dff_A_sRfhcl926_1),.din(w_dff_A_ihW1BRz73_1),.clk(gclk));
	jdff dff_A_XHsNrMzL4_1(.dout(w_dff_A_ihW1BRz73_1),.din(w_dff_A_XHsNrMzL4_1),.clk(gclk));
	jdff dff_A_MCNX1YCM4_1(.dout(w_dff_A_XHsNrMzL4_1),.din(w_dff_A_MCNX1YCM4_1),.clk(gclk));
	jdff dff_A_K2FeAn602_1(.dout(w_n470_0[1]),.din(w_dff_A_K2FeAn602_1),.clk(gclk));
	jdff dff_A_lkVNIif41_1(.dout(w_dff_A_K2FeAn602_1),.din(w_dff_A_lkVNIif41_1),.clk(gclk));
	jdff dff_A_5OAbYRuu6_1(.dout(w_dff_A_lkVNIif41_1),.din(w_dff_A_5OAbYRuu6_1),.clk(gclk));
	jdff dff_A_m59Tvl0e4_1(.dout(w_dff_A_5OAbYRuu6_1),.din(w_dff_A_m59Tvl0e4_1),.clk(gclk));
	jdff dff_A_3B1BqbPB2_1(.dout(w_dff_A_m59Tvl0e4_1),.din(w_dff_A_3B1BqbPB2_1),.clk(gclk));
	jdff dff_A_KcalhAAw7_1(.dout(w_dff_A_3B1BqbPB2_1),.din(w_dff_A_KcalhAAw7_1),.clk(gclk));
	jdff dff_A_126Nwlt32_1(.dout(w_dff_A_KcalhAAw7_1),.din(w_dff_A_126Nwlt32_1),.clk(gclk));
	jdff dff_A_8gbLF7Hy3_1(.dout(w_dff_A_126Nwlt32_1),.din(w_dff_A_8gbLF7Hy3_1),.clk(gclk));
	jdff dff_A_8R3nUI8J7_1(.dout(w_dff_A_8gbLF7Hy3_1),.din(w_dff_A_8R3nUI8J7_1),.clk(gclk));
	jdff dff_A_XbsvL4823_1(.dout(w_dff_A_8R3nUI8J7_1),.din(w_dff_A_XbsvL4823_1),.clk(gclk));
	jdff dff_A_9xyuKzU62_1(.dout(w_dff_A_XbsvL4823_1),.din(w_dff_A_9xyuKzU62_1),.clk(gclk));
	jdff dff_A_sqdGKtFa8_1(.dout(w_dff_A_9xyuKzU62_1),.din(w_dff_A_sqdGKtFa8_1),.clk(gclk));
	jdff dff_A_1KBnA3xU1_1(.dout(w_dff_A_sqdGKtFa8_1),.din(w_dff_A_1KBnA3xU1_1),.clk(gclk));
	jdff dff_A_JrGpFuJX4_1(.dout(w_dff_A_1KBnA3xU1_1),.din(w_dff_A_JrGpFuJX4_1),.clk(gclk));
	jdff dff_A_vkXhnAcW9_1(.dout(w_dff_A_JrGpFuJX4_1),.din(w_dff_A_vkXhnAcW9_1),.clk(gclk));
	jdff dff_A_oxU45Yxl4_1(.dout(w_dff_A_vkXhnAcW9_1),.din(w_dff_A_oxU45Yxl4_1),.clk(gclk));
	jdff dff_A_XhlpIIz80_1(.dout(w_dff_A_oxU45Yxl4_1),.din(w_dff_A_XhlpIIz80_1),.clk(gclk));
	jdff dff_A_EKDNYNzA3_1(.dout(w_dff_A_XhlpIIz80_1),.din(w_dff_A_EKDNYNzA3_1),.clk(gclk));
	jdff dff_A_S6jx6gYA3_1(.dout(w_dff_A_EKDNYNzA3_1),.din(w_dff_A_S6jx6gYA3_1),.clk(gclk));
	jdff dff_A_Z31eQSZF6_1(.dout(w_dff_A_S6jx6gYA3_1),.din(w_dff_A_Z31eQSZF6_1),.clk(gclk));
	jdff dff_A_DZZnkvIi2_1(.dout(w_dff_A_Z31eQSZF6_1),.din(w_dff_A_DZZnkvIi2_1),.clk(gclk));
	jdff dff_A_9cFfsQxC2_1(.dout(w_dff_A_DZZnkvIi2_1),.din(w_dff_A_9cFfsQxC2_1),.clk(gclk));
	jdff dff_A_qogrGZcT3_1(.dout(w_dff_A_9cFfsQxC2_1),.din(w_dff_A_qogrGZcT3_1),.clk(gclk));
	jdff dff_A_O3raPL9z5_1(.dout(w_dff_A_qogrGZcT3_1),.din(w_dff_A_O3raPL9z5_1),.clk(gclk));
	jdff dff_A_5A8AnfSW3_1(.dout(w_dff_A_O3raPL9z5_1),.din(w_dff_A_5A8AnfSW3_1),.clk(gclk));
	jdff dff_A_PvTO2xKm6_2(.dout(w_n470_0[2]),.din(w_dff_A_PvTO2xKm6_2),.clk(gclk));
	jdff dff_A_u8HoK95L0_1(.dout(w_n469_0[1]),.din(w_dff_A_u8HoK95L0_1),.clk(gclk));
	jdff dff_B_s4eA4dZI1_0(.din(n468),.dout(w_dff_B_s4eA4dZI1_0),.clk(gclk));
	jdff dff_B_FXRdcySs7_0(.din(G144),.dout(w_dff_B_FXRdcySs7_0),.clk(gclk));
	jdff dff_B_1p7mmdux0_2(.din(n466),.dout(w_dff_B_1p7mmdux0_2),.clk(gclk));
	jdff dff_B_JpelzHeC9_2(.din(w_dff_B_1p7mmdux0_2),.dout(w_dff_B_JpelzHeC9_2),.clk(gclk));
	jdff dff_A_M8I6GfXi6_0(.dout(w_G2224_1[0]),.din(w_dff_A_M8I6GfXi6_0),.clk(gclk));
	jdff dff_A_NQpzEZHc9_0(.dout(w_dff_A_M8I6GfXi6_0),.din(w_dff_A_NQpzEZHc9_0),.clk(gclk));
	jdff dff_A_ihlNcuCP0_0(.dout(w_dff_A_NQpzEZHc9_0),.din(w_dff_A_ihlNcuCP0_0),.clk(gclk));
	jdff dff_A_hBAC02z23_0(.dout(w_dff_A_ihlNcuCP0_0),.din(w_dff_A_hBAC02z23_0),.clk(gclk));
	jdff dff_A_cjpTw9ug5_1(.dout(w_n465_0[1]),.din(w_dff_A_cjpTw9ug5_1),.clk(gclk));
	jdff dff_B_VNDBVOTU3_2(.din(n465),.dout(w_dff_B_VNDBVOTU3_2),.clk(gclk));
	jdff dff_B_RtRPpRmP0_2(.din(w_dff_B_VNDBVOTU3_2),.dout(w_dff_B_RtRPpRmP0_2),.clk(gclk));
	jdff dff_B_VqLeReC87_2(.din(w_dff_B_RtRPpRmP0_2),.dout(w_dff_B_VqLeReC87_2),.clk(gclk));
	jdff dff_B_La6GKKE27_2(.din(w_dff_B_VqLeReC87_2),.dout(w_dff_B_La6GKKE27_2),.clk(gclk));
	jdff dff_A_HnBWU2jf4_1(.dout(w_n464_0[1]),.din(w_dff_A_HnBWU2jf4_1),.clk(gclk));
	jdff dff_A_1Vt5rRGr6_1(.dout(w_dff_A_HnBWU2jf4_1),.din(w_dff_A_1Vt5rRGr6_1),.clk(gclk));
	jdff dff_A_Dgt347V98_1(.dout(w_dff_A_1Vt5rRGr6_1),.din(w_dff_A_Dgt347V98_1),.clk(gclk));
	jdff dff_A_aLjvMWy45_1(.dout(w_dff_A_Dgt347V98_1),.din(w_dff_A_aLjvMWy45_1),.clk(gclk));
	jdff dff_A_nwifDyRU6_1(.dout(w_dff_A_aLjvMWy45_1),.din(w_dff_A_nwifDyRU6_1),.clk(gclk));
	jdff dff_A_M8CUetKr4_1(.dout(w_dff_A_nwifDyRU6_1),.din(w_dff_A_M8CUetKr4_1),.clk(gclk));
	jdff dff_A_UffxN78d5_1(.dout(w_dff_A_M8CUetKr4_1),.din(w_dff_A_UffxN78d5_1),.clk(gclk));
	jdff dff_A_p7TklzM11_1(.dout(w_dff_A_UffxN78d5_1),.din(w_dff_A_p7TklzM11_1),.clk(gclk));
	jdff dff_A_lu1XPUva1_1(.dout(w_dff_A_p7TklzM11_1),.din(w_dff_A_lu1XPUva1_1),.clk(gclk));
	jdff dff_A_xUke9Sjr9_1(.dout(w_dff_A_lu1XPUva1_1),.din(w_dff_A_xUke9Sjr9_1),.clk(gclk));
	jdff dff_A_N7g21i1s1_1(.dout(w_dff_A_xUke9Sjr9_1),.din(w_dff_A_N7g21i1s1_1),.clk(gclk));
	jdff dff_A_ZS28p3fN6_1(.dout(w_dff_A_N7g21i1s1_1),.din(w_dff_A_ZS28p3fN6_1),.clk(gclk));
	jdff dff_A_76zefZ4f4_1(.dout(w_dff_A_ZS28p3fN6_1),.din(w_dff_A_76zefZ4f4_1),.clk(gclk));
	jdff dff_A_hVXxn5s43_1(.dout(w_dff_A_76zefZ4f4_1),.din(w_dff_A_hVXxn5s43_1),.clk(gclk));
	jdff dff_A_vvj5LD029_1(.dout(w_dff_A_hVXxn5s43_1),.din(w_dff_A_vvj5LD029_1),.clk(gclk));
	jdff dff_A_FR1jVPtN9_1(.dout(w_dff_A_vvj5LD029_1),.din(w_dff_A_FR1jVPtN9_1),.clk(gclk));
	jdff dff_A_6A0JHep92_1(.dout(w_dff_A_FR1jVPtN9_1),.din(w_dff_A_6A0JHep92_1),.clk(gclk));
	jdff dff_A_0VlJsJY14_1(.dout(w_dff_A_6A0JHep92_1),.din(w_dff_A_0VlJsJY14_1),.clk(gclk));
	jdff dff_A_IBc3Xsp34_1(.dout(w_dff_A_0VlJsJY14_1),.din(w_dff_A_IBc3Xsp34_1),.clk(gclk));
	jdff dff_A_VlQXuF739_1(.dout(w_dff_A_IBc3Xsp34_1),.din(w_dff_A_VlQXuF739_1),.clk(gclk));
	jdff dff_A_zq2jNuoz6_1(.dout(w_dff_A_VlQXuF739_1),.din(w_dff_A_zq2jNuoz6_1),.clk(gclk));
	jdff dff_A_BWZ39dDq9_1(.dout(w_dff_A_zq2jNuoz6_1),.din(w_dff_A_BWZ39dDq9_1),.clk(gclk));
	jdff dff_A_xPtfVNsz4_1(.dout(w_dff_A_BWZ39dDq9_1),.din(w_dff_A_xPtfVNsz4_1),.clk(gclk));
	jdff dff_A_Bu5drJXT4_1(.dout(w_dff_A_xPtfVNsz4_1),.din(w_dff_A_Bu5drJXT4_1),.clk(gclk));
	jdff dff_A_z48JbY1H5_1(.dout(w_dff_A_Bu5drJXT4_1),.din(w_dff_A_z48JbY1H5_1),.clk(gclk));
	jdff dff_A_4UQNzWyN7_1(.dout(w_dff_A_z48JbY1H5_1),.din(w_dff_A_4UQNzWyN7_1),.clk(gclk));
	jdff dff_A_TYg8Tdpr4_0(.dout(w_n463_1[0]),.din(w_dff_A_TYg8Tdpr4_0),.clk(gclk));
	jdff dff_A_jMkhOUGu5_0(.dout(w_dff_A_TYg8Tdpr4_0),.din(w_dff_A_jMkhOUGu5_0),.clk(gclk));
	jdff dff_A_9ygve7a99_0(.dout(w_dff_A_jMkhOUGu5_0),.din(w_dff_A_9ygve7a99_0),.clk(gclk));
	jdff dff_A_bDWqOgy68_0(.dout(w_dff_A_9ygve7a99_0),.din(w_dff_A_bDWqOgy68_0),.clk(gclk));
	jdff dff_A_4wlQ1R3V9_0(.dout(w_dff_A_bDWqOgy68_0),.din(w_dff_A_4wlQ1R3V9_0),.clk(gclk));
	jdff dff_A_h1X0O4xv7_0(.dout(w_dff_A_4wlQ1R3V9_0),.din(w_dff_A_h1X0O4xv7_0),.clk(gclk));
	jdff dff_A_3zzVk0uX3_0(.dout(w_dff_A_h1X0O4xv7_0),.din(w_dff_A_3zzVk0uX3_0),.clk(gclk));
	jdff dff_A_RI2R0slG6_0(.dout(w_dff_A_3zzVk0uX3_0),.din(w_dff_A_RI2R0slG6_0),.clk(gclk));
	jdff dff_A_aZaxS6Bx2_0(.dout(w_dff_A_RI2R0slG6_0),.din(w_dff_A_aZaxS6Bx2_0),.clk(gclk));
	jdff dff_A_H1S0Lj2M4_0(.dout(w_dff_A_aZaxS6Bx2_0),.din(w_dff_A_H1S0Lj2M4_0),.clk(gclk));
	jdff dff_A_GRgmCoC55_0(.dout(w_dff_A_H1S0Lj2M4_0),.din(w_dff_A_GRgmCoC55_0),.clk(gclk));
	jdff dff_A_qQkC2sPC0_0(.dout(w_dff_A_GRgmCoC55_0),.din(w_dff_A_qQkC2sPC0_0),.clk(gclk));
	jdff dff_A_hEXqIV035_0(.dout(w_dff_A_qQkC2sPC0_0),.din(w_dff_A_hEXqIV035_0),.clk(gclk));
	jdff dff_A_CAsVwaVG4_0(.dout(w_dff_A_hEXqIV035_0),.din(w_dff_A_CAsVwaVG4_0),.clk(gclk));
	jdff dff_A_ntPRJ1Yt2_0(.dout(w_dff_A_CAsVwaVG4_0),.din(w_dff_A_ntPRJ1Yt2_0),.clk(gclk));
	jdff dff_A_UfHD95A03_0(.dout(w_dff_A_ntPRJ1Yt2_0),.din(w_dff_A_UfHD95A03_0),.clk(gclk));
	jdff dff_A_xwjjFYpY0_0(.dout(w_dff_A_UfHD95A03_0),.din(w_dff_A_xwjjFYpY0_0),.clk(gclk));
	jdff dff_A_HY38IcR00_0(.dout(w_dff_A_xwjjFYpY0_0),.din(w_dff_A_HY38IcR00_0),.clk(gclk));
	jdff dff_A_lgy4JPt34_0(.dout(w_dff_A_HY38IcR00_0),.din(w_dff_A_lgy4JPt34_0),.clk(gclk));
	jdff dff_A_vL5RymjX7_0(.dout(w_dff_A_lgy4JPt34_0),.din(w_dff_A_vL5RymjX7_0),.clk(gclk));
	jdff dff_A_dhVN3lCB6_0(.dout(w_dff_A_vL5RymjX7_0),.din(w_dff_A_dhVN3lCB6_0),.clk(gclk));
	jdff dff_A_prACCyXJ7_0(.dout(w_dff_A_dhVN3lCB6_0),.din(w_dff_A_prACCyXJ7_0),.clk(gclk));
	jdff dff_A_rz6XL2OO5_0(.dout(w_dff_A_prACCyXJ7_0),.din(w_dff_A_rz6XL2OO5_0),.clk(gclk));
	jdff dff_A_u4ZDMtqK4_0(.dout(w_dff_A_rz6XL2OO5_0),.din(w_dff_A_u4ZDMtqK4_0),.clk(gclk));
	jdff dff_A_28w2Jigz5_0(.dout(w_dff_A_u4ZDMtqK4_0),.din(w_dff_A_28w2Jigz5_0),.clk(gclk));
	jdff dff_A_cP91ZrdY0_0(.dout(w_dff_A_28w2Jigz5_0),.din(w_dff_A_cP91ZrdY0_0),.clk(gclk));
	jdff dff_A_ADIvEDMc5_0(.dout(w_dff_A_cP91ZrdY0_0),.din(w_dff_A_ADIvEDMc5_0),.clk(gclk));
	jdff dff_A_NO57E4si4_0(.dout(w_dff_A_ADIvEDMc5_0),.din(w_dff_A_NO57E4si4_0),.clk(gclk));
	jdff dff_A_31WWWRHU3_1(.dout(w_n463_0[1]),.din(w_dff_A_31WWWRHU3_1),.clk(gclk));
	jdff dff_A_1aLQFsMz9_1(.dout(w_dff_A_31WWWRHU3_1),.din(w_dff_A_1aLQFsMz9_1),.clk(gclk));
	jdff dff_A_QVBtoqvc1_1(.dout(w_dff_A_1aLQFsMz9_1),.din(w_dff_A_QVBtoqvc1_1),.clk(gclk));
	jdff dff_A_xC4ZM0WA6_2(.dout(w_n463_0[2]),.din(w_dff_A_xC4ZM0WA6_2),.clk(gclk));
	jdff dff_A_QF1WnZsW7_2(.dout(w_dff_A_xC4ZM0WA6_2),.din(w_dff_A_QF1WnZsW7_2),.clk(gclk));
	jdff dff_A_Dujt7ChK9_2(.dout(w_dff_A_QF1WnZsW7_2),.din(w_dff_A_Dujt7ChK9_2),.clk(gclk));
	jdff dff_A_iJUqX09N6_2(.dout(w_dff_A_Dujt7ChK9_2),.din(w_dff_A_iJUqX09N6_2),.clk(gclk));
	jdff dff_A_g2m1xBFl8_1(.dout(w_n462_0[1]),.din(w_dff_A_g2m1xBFl8_1),.clk(gclk));
	jdff dff_A_B0oME9l07_1(.dout(w_dff_A_g2m1xBFl8_1),.din(w_dff_A_B0oME9l07_1),.clk(gclk));
	jdff dff_A_9jqs9Xlx5_1(.dout(w_dff_A_B0oME9l07_1),.din(w_dff_A_9jqs9Xlx5_1),.clk(gclk));
	jdff dff_A_uaDqfkQw2_1(.dout(w_dff_A_9jqs9Xlx5_1),.din(w_dff_A_uaDqfkQw2_1),.clk(gclk));
	jdff dff_A_IvlrDlFz0_1(.dout(w_dff_A_uaDqfkQw2_1),.din(w_dff_A_IvlrDlFz0_1),.clk(gclk));
	jdff dff_A_vWMoivkc3_1(.dout(w_dff_A_IvlrDlFz0_1),.din(w_dff_A_vWMoivkc3_1),.clk(gclk));
	jdff dff_A_OU0AZkxh6_1(.dout(w_dff_A_vWMoivkc3_1),.din(w_dff_A_OU0AZkxh6_1),.clk(gclk));
	jdff dff_A_hOFzT9tM4_1(.dout(w_dff_A_OU0AZkxh6_1),.din(w_dff_A_hOFzT9tM4_1),.clk(gclk));
	jdff dff_A_kXitvI2w6_1(.dout(w_dff_A_hOFzT9tM4_1),.din(w_dff_A_kXitvI2w6_1),.clk(gclk));
	jdff dff_A_kEHsHiiy8_1(.dout(w_dff_A_kXitvI2w6_1),.din(w_dff_A_kEHsHiiy8_1),.clk(gclk));
	jdff dff_A_igPE98EO4_1(.dout(w_dff_A_kEHsHiiy8_1),.din(w_dff_A_igPE98EO4_1),.clk(gclk));
	jdff dff_A_MdzvNzrV6_1(.dout(w_dff_A_igPE98EO4_1),.din(w_dff_A_MdzvNzrV6_1),.clk(gclk));
	jdff dff_A_FhSiNrK38_1(.dout(w_dff_A_MdzvNzrV6_1),.din(w_dff_A_FhSiNrK38_1),.clk(gclk));
	jdff dff_A_aH8OxooQ2_1(.dout(w_dff_A_FhSiNrK38_1),.din(w_dff_A_aH8OxooQ2_1),.clk(gclk));
	jdff dff_A_Qu7i0AOX5_1(.dout(w_dff_A_aH8OxooQ2_1),.din(w_dff_A_Qu7i0AOX5_1),.clk(gclk));
	jdff dff_A_KUTh1DLr8_1(.dout(w_dff_A_Qu7i0AOX5_1),.din(w_dff_A_KUTh1DLr8_1),.clk(gclk));
	jdff dff_A_Ua2Ycfdy6_1(.dout(w_dff_A_KUTh1DLr8_1),.din(w_dff_A_Ua2Ycfdy6_1),.clk(gclk));
	jdff dff_A_gHT68AVI8_1(.dout(w_dff_A_Ua2Ycfdy6_1),.din(w_dff_A_gHT68AVI8_1),.clk(gclk));
	jdff dff_A_qNbB8PSW1_1(.dout(w_dff_A_gHT68AVI8_1),.din(w_dff_A_qNbB8PSW1_1),.clk(gclk));
	jdff dff_A_pmqbbcJL1_1(.dout(w_dff_A_qNbB8PSW1_1),.din(w_dff_A_pmqbbcJL1_1),.clk(gclk));
	jdff dff_A_X9cBIOx54_1(.dout(w_dff_A_pmqbbcJL1_1),.din(w_dff_A_X9cBIOx54_1),.clk(gclk));
	jdff dff_A_5Z81xz2U1_2(.dout(w_n462_0[2]),.din(w_dff_A_5Z81xz2U1_2),.clk(gclk));
	jdff dff_A_LnyJASmM1_2(.dout(w_dff_A_5Z81xz2U1_2),.din(w_dff_A_LnyJASmM1_2),.clk(gclk));
	jdff dff_A_j0ldxZUh0_2(.dout(w_dff_A_LnyJASmM1_2),.din(w_dff_A_j0ldxZUh0_2),.clk(gclk));
	jdff dff_A_HIduge0I7_2(.dout(w_dff_A_j0ldxZUh0_2),.din(w_dff_A_HIduge0I7_2),.clk(gclk));
	jdff dff_A_l6iDbYvx2_2(.dout(w_dff_A_HIduge0I7_2),.din(w_dff_A_l6iDbYvx2_2),.clk(gclk));
	jdff dff_B_ROfqi5sd5_1(.din(n454),.dout(w_dff_B_ROfqi5sd5_1),.clk(gclk));
	jdff dff_A_r9uNt09E4_0(.dout(w_n460_1[0]),.din(w_dff_A_r9uNt09E4_0),.clk(gclk));
	jdff dff_A_rkdl9ovW0_0(.dout(w_dff_A_r9uNt09E4_0),.din(w_dff_A_rkdl9ovW0_0),.clk(gclk));
	jdff dff_A_RK9WZi2Q1_0(.dout(w_dff_A_rkdl9ovW0_0),.din(w_dff_A_RK9WZi2Q1_0),.clk(gclk));
	jdff dff_A_43ymp5HH0_0(.dout(w_dff_A_RK9WZi2Q1_0),.din(w_dff_A_43ymp5HH0_0),.clk(gclk));
	jdff dff_A_PlUjBCk18_0(.dout(w_dff_A_43ymp5HH0_0),.din(w_dff_A_PlUjBCk18_0),.clk(gclk));
	jdff dff_A_nalhsrNs8_0(.dout(w_dff_A_PlUjBCk18_0),.din(w_dff_A_nalhsrNs8_0),.clk(gclk));
	jdff dff_A_gTodIcZt1_0(.dout(w_dff_A_nalhsrNs8_0),.din(w_dff_A_gTodIcZt1_0),.clk(gclk));
	jdff dff_A_0c4x3L2H1_0(.dout(w_dff_A_gTodIcZt1_0),.din(w_dff_A_0c4x3L2H1_0),.clk(gclk));
	jdff dff_A_8Wunz3Gz6_0(.dout(w_dff_A_0c4x3L2H1_0),.din(w_dff_A_8Wunz3Gz6_0),.clk(gclk));
	jdff dff_A_F96IB2Yj5_0(.dout(w_dff_A_8Wunz3Gz6_0),.din(w_dff_A_F96IB2Yj5_0),.clk(gclk));
	jdff dff_A_cVlb8Lai2_0(.dout(w_dff_A_F96IB2Yj5_0),.din(w_dff_A_cVlb8Lai2_0),.clk(gclk));
	jdff dff_A_q4kPMBVf3_0(.dout(w_dff_A_cVlb8Lai2_0),.din(w_dff_A_q4kPMBVf3_0),.clk(gclk));
	jdff dff_A_7ecolecs9_0(.dout(w_dff_A_q4kPMBVf3_0),.din(w_dff_A_7ecolecs9_0),.clk(gclk));
	jdff dff_A_dLJrDbS01_0(.dout(w_dff_A_7ecolecs9_0),.din(w_dff_A_dLJrDbS01_0),.clk(gclk));
	jdff dff_A_YNLs3Fpt1_0(.dout(w_dff_A_dLJrDbS01_0),.din(w_dff_A_YNLs3Fpt1_0),.clk(gclk));
	jdff dff_A_nWYj38gu5_0(.dout(w_dff_A_YNLs3Fpt1_0),.din(w_dff_A_nWYj38gu5_0),.clk(gclk));
	jdff dff_A_fjHQlS0k7_0(.dout(w_dff_A_nWYj38gu5_0),.din(w_dff_A_fjHQlS0k7_0),.clk(gclk));
	jdff dff_A_FmFN1t1E6_0(.dout(w_dff_A_fjHQlS0k7_0),.din(w_dff_A_FmFN1t1E6_0),.clk(gclk));
	jdff dff_A_07zxERxa6_0(.dout(w_dff_A_FmFN1t1E6_0),.din(w_dff_A_07zxERxa6_0),.clk(gclk));
	jdff dff_A_hE3TMeAi0_0(.dout(w_dff_A_07zxERxa6_0),.din(w_dff_A_hE3TMeAi0_0),.clk(gclk));
	jdff dff_A_vf7Phuzu2_0(.dout(w_dff_A_hE3TMeAi0_0),.din(w_dff_A_vf7Phuzu2_0),.clk(gclk));
	jdff dff_A_1k4KbDb68_0(.dout(w_dff_A_vf7Phuzu2_0),.din(w_dff_A_1k4KbDb68_0),.clk(gclk));
	jdff dff_A_wAN75iSl7_0(.dout(w_dff_A_1k4KbDb68_0),.din(w_dff_A_wAN75iSl7_0),.clk(gclk));
	jdff dff_A_YRBUIWw11_0(.dout(w_dff_A_wAN75iSl7_0),.din(w_dff_A_YRBUIWw11_0),.clk(gclk));
	jdff dff_A_9lgaDUz22_0(.dout(w_dff_A_YRBUIWw11_0),.din(w_dff_A_9lgaDUz22_0),.clk(gclk));
	jdff dff_A_HkY0Ozwo5_0(.dout(w_dff_A_9lgaDUz22_0),.din(w_dff_A_HkY0Ozwo5_0),.clk(gclk));
	jdff dff_A_pC9SxTcg1_0(.dout(w_dff_A_HkY0Ozwo5_0),.din(w_dff_A_pC9SxTcg1_0),.clk(gclk));
	jdff dff_A_wPtHeeCc1_0(.dout(w_dff_A_pC9SxTcg1_0),.din(w_dff_A_wPtHeeCc1_0),.clk(gclk));
	jdff dff_A_3ZpI47qr9_1(.dout(w_n460_1[1]),.din(w_dff_A_3ZpI47qr9_1),.clk(gclk));
	jdff dff_A_bFQNGcgB9_1(.dout(w_dff_A_3ZpI47qr9_1),.din(w_dff_A_bFQNGcgB9_1),.clk(gclk));
	jdff dff_A_MZshv5gh3_1(.dout(w_dff_A_bFQNGcgB9_1),.din(w_dff_A_MZshv5gh3_1),.clk(gclk));
	jdff dff_A_TwH1swP31_1(.dout(w_dff_A_MZshv5gh3_1),.din(w_dff_A_TwH1swP31_1),.clk(gclk));
	jdff dff_A_8HORNGw25_1(.dout(w_dff_A_TwH1swP31_1),.din(w_dff_A_8HORNGw25_1),.clk(gclk));
	jdff dff_A_xFMB9gpv5_1(.dout(w_dff_A_8HORNGw25_1),.din(w_dff_A_xFMB9gpv5_1),.clk(gclk));
	jdff dff_A_5NdSYsBJ7_1(.dout(w_dff_A_xFMB9gpv5_1),.din(w_dff_A_5NdSYsBJ7_1),.clk(gclk));
	jdff dff_A_vcR82Vn03_1(.dout(w_dff_A_5NdSYsBJ7_1),.din(w_dff_A_vcR82Vn03_1),.clk(gclk));
	jdff dff_A_reVZ7qnZ6_1(.dout(w_dff_A_vcR82Vn03_1),.din(w_dff_A_reVZ7qnZ6_1),.clk(gclk));
	jdff dff_A_DrHrwRI04_1(.dout(w_dff_A_reVZ7qnZ6_1),.din(w_dff_A_DrHrwRI04_1),.clk(gclk));
	jdff dff_A_tbLMEGHm9_1(.dout(w_dff_A_DrHrwRI04_1),.din(w_dff_A_tbLMEGHm9_1),.clk(gclk));
	jdff dff_A_0u21JPMa1_1(.dout(w_dff_A_tbLMEGHm9_1),.din(w_dff_A_0u21JPMa1_1),.clk(gclk));
	jdff dff_A_9W78x3VH4_1(.dout(w_dff_A_0u21JPMa1_1),.din(w_dff_A_9W78x3VH4_1),.clk(gclk));
	jdff dff_A_oHtssPdj0_1(.dout(w_dff_A_9W78x3VH4_1),.din(w_dff_A_oHtssPdj0_1),.clk(gclk));
	jdff dff_A_C2oswGKJ7_1(.dout(w_dff_A_oHtssPdj0_1),.din(w_dff_A_C2oswGKJ7_1),.clk(gclk));
	jdff dff_A_ez8dfd7Z7_1(.dout(w_dff_A_C2oswGKJ7_1),.din(w_dff_A_ez8dfd7Z7_1),.clk(gclk));
	jdff dff_A_V8dlpBUk4_1(.dout(w_dff_A_ez8dfd7Z7_1),.din(w_dff_A_V8dlpBUk4_1),.clk(gclk));
	jdff dff_A_y6e35GZE3_1(.dout(w_dff_A_V8dlpBUk4_1),.din(w_dff_A_y6e35GZE3_1),.clk(gclk));
	jdff dff_A_YErLJ0Y63_1(.dout(w_dff_A_y6e35GZE3_1),.din(w_dff_A_YErLJ0Y63_1),.clk(gclk));
	jdff dff_A_JWPlhfRX4_1(.dout(w_dff_A_YErLJ0Y63_1),.din(w_dff_A_JWPlhfRX4_1),.clk(gclk));
	jdff dff_A_oghk7Wwo4_1(.dout(w_dff_A_JWPlhfRX4_1),.din(w_dff_A_oghk7Wwo4_1),.clk(gclk));
	jdff dff_A_ZE5QrrRW7_1(.dout(w_dff_A_oghk7Wwo4_1),.din(w_dff_A_ZE5QrrRW7_1),.clk(gclk));
	jdff dff_A_jiaZanyy9_1(.dout(w_dff_A_ZE5QrrRW7_1),.din(w_dff_A_jiaZanyy9_1),.clk(gclk));
	jdff dff_A_qTxX4T0S2_1(.dout(w_dff_A_jiaZanyy9_1),.din(w_dff_A_qTxX4T0S2_1),.clk(gclk));
	jdff dff_A_Ni3xbxCS0_1(.dout(w_dff_A_qTxX4T0S2_1),.din(w_dff_A_Ni3xbxCS0_1),.clk(gclk));
	jdff dff_A_D5Uy5jKu4_1(.dout(w_dff_A_Ni3xbxCS0_1),.din(w_dff_A_D5Uy5jKu4_1),.clk(gclk));
	jdff dff_A_6Hqpq9og1_1(.dout(w_dff_A_D5Uy5jKu4_1),.din(w_dff_A_6Hqpq9og1_1),.clk(gclk));
	jdff dff_A_hi7zk1CR7_1(.dout(w_n460_0[1]),.din(w_dff_A_hi7zk1CR7_1),.clk(gclk));
	jdff dff_A_LF35YLmI6_1(.dout(w_dff_A_hi7zk1CR7_1),.din(w_dff_A_LF35YLmI6_1),.clk(gclk));
	jdff dff_A_zcRclED08_1(.dout(w_dff_A_LF35YLmI6_1),.din(w_dff_A_zcRclED08_1),.clk(gclk));
	jdff dff_A_fJ6Z2Fym0_1(.dout(w_dff_A_zcRclED08_1),.din(w_dff_A_fJ6Z2Fym0_1),.clk(gclk));
	jdff dff_A_H6YW1Fir0_1(.dout(w_dff_A_fJ6Z2Fym0_1),.din(w_dff_A_H6YW1Fir0_1),.clk(gclk));
	jdff dff_A_ELfZLHUX2_1(.dout(w_dff_A_H6YW1Fir0_1),.din(w_dff_A_ELfZLHUX2_1),.clk(gclk));
	jdff dff_A_tbc2fNk24_2(.dout(w_n460_0[2]),.din(w_dff_A_tbc2fNk24_2),.clk(gclk));
	jdff dff_A_ZO8xir4g0_2(.dout(w_dff_A_tbc2fNk24_2),.din(w_dff_A_ZO8xir4g0_2),.clk(gclk));
	jdff dff_A_llcSN2BG4_2(.dout(w_dff_A_ZO8xir4g0_2),.din(w_dff_A_llcSN2BG4_2),.clk(gclk));
	jdff dff_A_pUa3w54x3_2(.dout(w_dff_A_llcSN2BG4_2),.din(w_dff_A_pUa3w54x3_2),.clk(gclk));
	jdff dff_A_g3dRlHVv4_2(.dout(w_dff_A_pUa3w54x3_2),.din(w_dff_A_g3dRlHVv4_2),.clk(gclk));
	jdff dff_A_4iMejImJ9_2(.dout(w_dff_A_g3dRlHVv4_2),.din(w_dff_A_4iMejImJ9_2),.clk(gclk));
	jdff dff_A_9WxyhcV15_2(.dout(w_dff_A_4iMejImJ9_2),.din(w_dff_A_9WxyhcV15_2),.clk(gclk));
	jdff dff_B_4ktNGoya8_0(.din(n458),.dout(w_dff_B_4ktNGoya8_0),.clk(gclk));
	jdff dff_B_W1sljb7y0_0(.din(G135),.dout(w_dff_B_W1sljb7y0_0),.clk(gclk));
	jdff dff_A_K55uznzv1_1(.dout(w_n456_0[1]),.din(w_dff_A_K55uznzv1_1),.clk(gclk));
	jdff dff_A_JnxynNQZ7_1(.dout(w_dff_A_K55uznzv1_1),.din(w_dff_A_JnxynNQZ7_1),.clk(gclk));
	jdff dff_A_iSt3pmoL4_2(.dout(w_n456_0[2]),.din(w_dff_A_iSt3pmoL4_2),.clk(gclk));
	jdff dff_A_fzA0RuAB8_2(.dout(w_dff_A_iSt3pmoL4_2),.din(w_dff_A_fzA0RuAB8_2),.clk(gclk));
	jdff dff_A_62mwjYD83_1(.dout(w_G2230_0[1]),.din(w_dff_A_62mwjYD83_1),.clk(gclk));
	jdff dff_A_KHSdDUvG7_1(.dout(w_dff_A_62mwjYD83_1),.din(w_dff_A_KHSdDUvG7_1),.clk(gclk));
	jdff dff_A_WpstJHKE4_1(.dout(w_dff_A_KHSdDUvG7_1),.din(w_dff_A_WpstJHKE4_1),.clk(gclk));
	jdff dff_A_cqRjat6f7_1(.dout(w_dff_A_WpstJHKE4_1),.din(w_dff_A_cqRjat6f7_1),.clk(gclk));
	jdff dff_A_tqesnuAW6_1(.dout(w_n453_0[1]),.din(w_dff_A_tqesnuAW6_1),.clk(gclk));
	jdff dff_B_1NhAGwVz7_0(.din(G157),.dout(w_dff_B_1NhAGwVz7_0),.clk(gclk));
	jdff dff_B_K5txonfB4_3(.din(n451),.dout(w_dff_B_K5txonfB4_3),.clk(gclk));
	jdff dff_B_ZTy8EqPV4_3(.din(w_dff_B_K5txonfB4_3),.dout(w_dff_B_ZTy8EqPV4_3),.clk(gclk));
	jdff dff_A_MbeNTaRo8_2(.dout(w_n450_0[2]),.din(w_dff_A_MbeNTaRo8_2),.clk(gclk));
	jdff dff_A_VqFYbCB53_2(.dout(w_dff_A_MbeNTaRo8_2),.din(w_dff_A_VqFYbCB53_2),.clk(gclk));
	jdff dff_A_tg13M2sT7_2(.dout(w_dff_A_VqFYbCB53_2),.din(w_dff_A_tg13M2sT7_2),.clk(gclk));
	jdff dff_A_6XrtcXTY6_2(.dout(w_dff_A_tg13M2sT7_2),.din(w_dff_A_6XrtcXTY6_2),.clk(gclk));
	jdff dff_A_jPNMqTsu8_2(.dout(w_dff_A_6XrtcXTY6_2),.din(w_dff_A_jPNMqTsu8_2),.clk(gclk));
	jdff dff_A_iMez3pks7_2(.dout(w_dff_A_jPNMqTsu8_2),.din(w_dff_A_iMez3pks7_2),.clk(gclk));
	jdff dff_A_ZwyOmiDg8_2(.dout(w_dff_A_iMez3pks7_2),.din(w_dff_A_ZwyOmiDg8_2),.clk(gclk));
	jdff dff_A_1pWxHSlY1_2(.dout(w_dff_A_ZwyOmiDg8_2),.din(w_dff_A_1pWxHSlY1_2),.clk(gclk));
	jdff dff_A_JDyQ9ai18_2(.dout(w_dff_A_1pWxHSlY1_2),.din(w_dff_A_JDyQ9ai18_2),.clk(gclk));
	jdff dff_A_iR6B7duH2_2(.dout(w_dff_A_JDyQ9ai18_2),.din(w_dff_A_iR6B7duH2_2),.clk(gclk));
	jdff dff_A_OaDpa0iQ4_2(.dout(w_dff_A_iR6B7duH2_2),.din(w_dff_A_OaDpa0iQ4_2),.clk(gclk));
	jdff dff_A_dyS1aMqS3_2(.dout(w_dff_A_OaDpa0iQ4_2),.din(w_dff_A_dyS1aMqS3_2),.clk(gclk));
	jdff dff_A_6pCGcHdt6_2(.dout(w_dff_A_dyS1aMqS3_2),.din(w_dff_A_6pCGcHdt6_2),.clk(gclk));
	jdff dff_A_yYbDhjX34_2(.dout(w_dff_A_6pCGcHdt6_2),.din(w_dff_A_yYbDhjX34_2),.clk(gclk));
	jdff dff_A_hQ8yQrNP2_2(.dout(w_dff_A_yYbDhjX34_2),.din(w_dff_A_hQ8yQrNP2_2),.clk(gclk));
	jdff dff_A_41mxgmIB7_2(.dout(w_dff_A_hQ8yQrNP2_2),.din(w_dff_A_41mxgmIB7_2),.clk(gclk));
	jdff dff_A_pYHGwCkf2_2(.dout(w_dff_A_41mxgmIB7_2),.din(w_dff_A_pYHGwCkf2_2),.clk(gclk));
	jdff dff_A_2D8usgXT5_2(.dout(w_dff_A_pYHGwCkf2_2),.din(w_dff_A_2D8usgXT5_2),.clk(gclk));
	jdff dff_A_hYOCOZMz8_2(.dout(w_dff_A_2D8usgXT5_2),.din(w_dff_A_hYOCOZMz8_2),.clk(gclk));
	jdff dff_A_FQOKUYsv5_2(.dout(w_dff_A_hYOCOZMz8_2),.din(w_dff_A_FQOKUYsv5_2),.clk(gclk));
	jdff dff_A_BfJp3bsu6_2(.dout(w_dff_A_FQOKUYsv5_2),.din(w_dff_A_BfJp3bsu6_2),.clk(gclk));
	jdff dff_A_yOGMEFVi3_2(.dout(w_dff_A_BfJp3bsu6_2),.din(w_dff_A_yOGMEFVi3_2),.clk(gclk));
	jdff dff_B_bEDm3zYn1_1(.din(n439),.dout(w_dff_B_bEDm3zYn1_1),.clk(gclk));
	jdff dff_B_BiI0ZTCU1_1(.din(w_dff_B_bEDm3zYn1_1),.dout(w_dff_B_BiI0ZTCU1_1),.clk(gclk));
	jdff dff_A_wjKWvZBb3_0(.dout(w_n449_1[0]),.din(w_dff_A_wjKWvZBb3_0),.clk(gclk));
	jdff dff_A_dJgKxRIC5_0(.dout(w_dff_A_wjKWvZBb3_0),.din(w_dff_A_dJgKxRIC5_0),.clk(gclk));
	jdff dff_A_1ZBRyKC30_0(.dout(w_dff_A_dJgKxRIC5_0),.din(w_dff_A_1ZBRyKC30_0),.clk(gclk));
	jdff dff_A_cVv02Nlj1_0(.dout(w_dff_A_1ZBRyKC30_0),.din(w_dff_A_cVv02Nlj1_0),.clk(gclk));
	jdff dff_A_rRkeo3GP2_0(.dout(w_dff_A_cVv02Nlj1_0),.din(w_dff_A_rRkeo3GP2_0),.clk(gclk));
	jdff dff_A_bldm7o9G6_0(.dout(w_dff_A_rRkeo3GP2_0),.din(w_dff_A_bldm7o9G6_0),.clk(gclk));
	jdff dff_A_sBerXbpX6_0(.dout(w_dff_A_bldm7o9G6_0),.din(w_dff_A_sBerXbpX6_0),.clk(gclk));
	jdff dff_A_kEVfi8W48_0(.dout(w_dff_A_sBerXbpX6_0),.din(w_dff_A_kEVfi8W48_0),.clk(gclk));
	jdff dff_A_itbCi6411_0(.dout(w_dff_A_kEVfi8W48_0),.din(w_dff_A_itbCi6411_0),.clk(gclk));
	jdff dff_A_ePQy4ze88_0(.dout(w_dff_A_itbCi6411_0),.din(w_dff_A_ePQy4ze88_0),.clk(gclk));
	jdff dff_A_gpQCK13v9_0(.dout(w_dff_A_ePQy4ze88_0),.din(w_dff_A_gpQCK13v9_0),.clk(gclk));
	jdff dff_A_VgxrRdz78_0(.dout(w_dff_A_gpQCK13v9_0),.din(w_dff_A_VgxrRdz78_0),.clk(gclk));
	jdff dff_A_2ObhRrl09_0(.dout(w_dff_A_VgxrRdz78_0),.din(w_dff_A_2ObhRrl09_0),.clk(gclk));
	jdff dff_A_2D63Mkir0_0(.dout(w_dff_A_2ObhRrl09_0),.din(w_dff_A_2D63Mkir0_0),.clk(gclk));
	jdff dff_A_ssscaKOB5_0(.dout(w_dff_A_2D63Mkir0_0),.din(w_dff_A_ssscaKOB5_0),.clk(gclk));
	jdff dff_A_YYVbMTHo0_0(.dout(w_dff_A_ssscaKOB5_0),.din(w_dff_A_YYVbMTHo0_0),.clk(gclk));
	jdff dff_A_YoUP7csR4_0(.dout(w_dff_A_YYVbMTHo0_0),.din(w_dff_A_YoUP7csR4_0),.clk(gclk));
	jdff dff_A_RHxQU68j4_0(.dout(w_dff_A_YoUP7csR4_0),.din(w_dff_A_RHxQU68j4_0),.clk(gclk));
	jdff dff_A_Ol441Uz21_0(.dout(w_dff_A_RHxQU68j4_0),.din(w_dff_A_Ol441Uz21_0),.clk(gclk));
	jdff dff_A_bxayRSXS9_0(.dout(w_dff_A_Ol441Uz21_0),.din(w_dff_A_bxayRSXS9_0),.clk(gclk));
	jdff dff_A_KChkSnBZ2_0(.dout(w_dff_A_bxayRSXS9_0),.din(w_dff_A_KChkSnBZ2_0),.clk(gclk));
	jdff dff_A_YDSTlRFl9_0(.dout(w_dff_A_KChkSnBZ2_0),.din(w_dff_A_YDSTlRFl9_0),.clk(gclk));
	jdff dff_B_pVUVu6oE9_1(.din(n442),.dout(w_dff_B_pVUVu6oE9_1),.clk(gclk));
	jdff dff_B_VEsaFXyh2_1(.din(n443),.dout(w_dff_B_VEsaFXyh2_1),.clk(gclk));
	jdff dff_B_2P3d0CEE3_1(.din(w_dff_B_VEsaFXyh2_1),.dout(w_dff_B_2P3d0CEE3_1),.clk(gclk));
	jdff dff_A_Yx4risHu8_1(.dout(w_n447_0[1]),.din(w_dff_A_Yx4risHu8_1),.clk(gclk));
	jdff dff_A_LPyXdJn96_1(.dout(w_dff_A_Yx4risHu8_1),.din(w_dff_A_LPyXdJn96_1),.clk(gclk));
	jdff dff_A_YRV2LOo14_1(.dout(w_dff_A_LPyXdJn96_1),.din(w_dff_A_YRV2LOo14_1),.clk(gclk));
	jdff dff_A_jPrX1cbm8_1(.dout(w_dff_A_YRV2LOo14_1),.din(w_dff_A_jPrX1cbm8_1),.clk(gclk));
	jdff dff_A_BQ09mqDV6_1(.dout(w_dff_A_jPrX1cbm8_1),.din(w_dff_A_BQ09mqDV6_1),.clk(gclk));
	jdff dff_A_hnGbZB4c2_1(.dout(w_dff_A_BQ09mqDV6_1),.din(w_dff_A_hnGbZB4c2_1),.clk(gclk));
	jdff dff_A_LoWAeYgW8_1(.dout(w_dff_A_hnGbZB4c2_1),.din(w_dff_A_LoWAeYgW8_1),.clk(gclk));
	jdff dff_A_aga1Qr7U6_1(.dout(w_dff_A_LoWAeYgW8_1),.din(w_dff_A_aga1Qr7U6_1),.clk(gclk));
	jdff dff_A_E6b3rdbL2_1(.dout(w_dff_A_aga1Qr7U6_1),.din(w_dff_A_E6b3rdbL2_1),.clk(gclk));
	jdff dff_A_H2JKbEBc0_1(.dout(w_dff_A_E6b3rdbL2_1),.din(w_dff_A_H2JKbEBc0_1),.clk(gclk));
	jdff dff_A_tHGxxEfW7_1(.dout(w_dff_A_H2JKbEBc0_1),.din(w_dff_A_tHGxxEfW7_1),.clk(gclk));
	jdff dff_A_SV50TXc59_1(.dout(w_dff_A_tHGxxEfW7_1),.din(w_dff_A_SV50TXc59_1),.clk(gclk));
	jdff dff_A_ZCa0qgEb5_1(.dout(w_dff_A_SV50TXc59_1),.din(w_dff_A_ZCa0qgEb5_1),.clk(gclk));
	jdff dff_A_seWYdYZu5_1(.dout(w_dff_A_ZCa0qgEb5_1),.din(w_dff_A_seWYdYZu5_1),.clk(gclk));
	jdff dff_A_esdau1Ez5_1(.dout(w_dff_A_seWYdYZu5_1),.din(w_dff_A_esdau1Ez5_1),.clk(gclk));
	jdff dff_A_88KGpDJV7_1(.dout(w_dff_A_esdau1Ez5_1),.din(w_dff_A_88KGpDJV7_1),.clk(gclk));
	jdff dff_A_sKYU1zDx5_1(.dout(w_dff_A_88KGpDJV7_1),.din(w_dff_A_sKYU1zDx5_1),.clk(gclk));
	jdff dff_A_o83YnuwY8_1(.dout(w_dff_A_sKYU1zDx5_1),.din(w_dff_A_o83YnuwY8_1),.clk(gclk));
	jdff dff_A_Tp2bWoNb3_1(.dout(w_dff_A_o83YnuwY8_1),.din(w_dff_A_Tp2bWoNb3_1),.clk(gclk));
	jdff dff_A_hXMuAwq23_1(.dout(w_dff_A_Tp2bWoNb3_1),.din(w_dff_A_hXMuAwq23_1),.clk(gclk));
	jdff dff_A_aNHrWs2m3_1(.dout(w_dff_A_hXMuAwq23_1),.din(w_dff_A_aNHrWs2m3_1),.clk(gclk));
	jdff dff_A_DCRuM31d7_1(.dout(w_dff_A_aNHrWs2m3_1),.din(w_dff_A_DCRuM31d7_1),.clk(gclk));
	jdff dff_A_cYntFtSi4_1(.dout(w_dff_A_DCRuM31d7_1),.din(w_dff_A_cYntFtSi4_1),.clk(gclk));
	jdff dff_A_kiwYSKer5_1(.dout(w_dff_A_cYntFtSi4_1),.din(w_dff_A_kiwYSKer5_1),.clk(gclk));
	jdff dff_A_DBXmQNFG7_1(.dout(w_dff_A_kiwYSKer5_1),.din(w_dff_A_DBXmQNFG7_1),.clk(gclk));
	jdff dff_A_7PWrwykw5_1(.dout(w_n445_0[1]),.din(w_dff_A_7PWrwykw5_1),.clk(gclk));
	jdff dff_A_tVTt4gd04_1(.dout(w_dff_A_7PWrwykw5_1),.din(w_dff_A_tVTt4gd04_1),.clk(gclk));
	jdff dff_A_gLGe0Teh8_1(.dout(w_dff_A_tVTt4gd04_1),.din(w_dff_A_gLGe0Teh8_1),.clk(gclk));
	jdff dff_A_9zluSdTd1_1(.dout(w_dff_A_gLGe0Teh8_1),.din(w_dff_A_9zluSdTd1_1),.clk(gclk));
	jdff dff_A_tlvcJgdQ4_1(.dout(w_dff_A_9zluSdTd1_1),.din(w_dff_A_tlvcJgdQ4_1),.clk(gclk));
	jdff dff_A_SJerHwCp5_1(.dout(w_dff_A_tlvcJgdQ4_1),.din(w_dff_A_SJerHwCp5_1),.clk(gclk));
	jdff dff_A_O0RnGL9Z6_1(.dout(w_dff_A_SJerHwCp5_1),.din(w_dff_A_O0RnGL9Z6_1),.clk(gclk));
	jdff dff_A_8c5mLC0Q5_1(.dout(w_dff_A_O0RnGL9Z6_1),.din(w_dff_A_8c5mLC0Q5_1),.clk(gclk));
	jdff dff_A_iUP3jbLH0_1(.dout(w_dff_A_8c5mLC0Q5_1),.din(w_dff_A_iUP3jbLH0_1),.clk(gclk));
	jdff dff_A_iLH3P6Ny7_1(.dout(w_dff_A_iUP3jbLH0_1),.din(w_dff_A_iLH3P6Ny7_1),.clk(gclk));
	jdff dff_A_iraFo22z3_1(.dout(w_dff_A_iLH3P6Ny7_1),.din(w_dff_A_iraFo22z3_1),.clk(gclk));
	jdff dff_A_BIz3xtaL1_1(.dout(w_dff_A_iraFo22z3_1),.din(w_dff_A_BIz3xtaL1_1),.clk(gclk));
	jdff dff_A_9wo9M0UM2_1(.dout(w_dff_A_BIz3xtaL1_1),.din(w_dff_A_9wo9M0UM2_1),.clk(gclk));
	jdff dff_A_ZlWK9vG67_1(.dout(w_dff_A_9wo9M0UM2_1),.din(w_dff_A_ZlWK9vG67_1),.clk(gclk));
	jdff dff_A_mrAwvEfd2_1(.dout(w_dff_A_ZlWK9vG67_1),.din(w_dff_A_mrAwvEfd2_1),.clk(gclk));
	jdff dff_A_RW5hLxVc4_1(.dout(w_dff_A_mrAwvEfd2_1),.din(w_dff_A_RW5hLxVc4_1),.clk(gclk));
	jdff dff_A_5WviFnyq4_1(.dout(w_dff_A_RW5hLxVc4_1),.din(w_dff_A_5WviFnyq4_1),.clk(gclk));
	jdff dff_A_Pmjqmfgp6_1(.dout(w_dff_A_5WviFnyq4_1),.din(w_dff_A_Pmjqmfgp6_1),.clk(gclk));
	jdff dff_A_cW8swT584_1(.dout(w_dff_A_Pmjqmfgp6_1),.din(w_dff_A_cW8swT584_1),.clk(gclk));
	jdff dff_A_yiEcr5Fi0_1(.dout(w_dff_A_cW8swT584_1),.din(w_dff_A_yiEcr5Fi0_1),.clk(gclk));
	jdff dff_A_7fMavj4h1_1(.dout(w_dff_A_yiEcr5Fi0_1),.din(w_dff_A_7fMavj4h1_1),.clk(gclk));
	jdff dff_A_kMawKvbe0_1(.dout(w_dff_A_7fMavj4h1_1),.din(w_dff_A_kMawKvbe0_1),.clk(gclk));
	jdff dff_A_Wj9KDVlV5_1(.dout(w_dff_A_kMawKvbe0_1),.din(w_dff_A_Wj9KDVlV5_1),.clk(gclk));
	jdff dff_A_GxaZnX183_1(.dout(w_dff_A_Wj9KDVlV5_1),.din(w_dff_A_GxaZnX183_1),.clk(gclk));
	jdff dff_A_Wdxvnsr97_1(.dout(w_dff_A_GxaZnX183_1),.din(w_dff_A_Wdxvnsr97_1),.clk(gclk));
	jdff dff_A_nRvZGQid1_1(.dout(w_dff_A_Wdxvnsr97_1),.din(w_dff_A_nRvZGQid1_1),.clk(gclk));
	jdff dff_A_vlI9QMAP8_1(.dout(w_n444_0[1]),.din(w_dff_A_vlI9QMAP8_1),.clk(gclk));
	jdff dff_A_mfUBjL8h2_1(.dout(w_dff_A_vlI9QMAP8_1),.din(w_dff_A_mfUBjL8h2_1),.clk(gclk));
	jdff dff_A_jGvha8wF0_2(.dout(w_n444_0[2]),.din(w_dff_A_jGvha8wF0_2),.clk(gclk));
	jdff dff_A_kggdpM1j0_0(.dout(w_n438_0[0]),.din(w_dff_A_kggdpM1j0_0),.clk(gclk));
	jdff dff_A_0oJUP1386_0(.dout(w_dff_A_kggdpM1j0_0),.din(w_dff_A_0oJUP1386_0),.clk(gclk));
	jdff dff_A_k5pLKUhv3_0(.dout(w_dff_A_0oJUP1386_0),.din(w_dff_A_k5pLKUhv3_0),.clk(gclk));
	jdff dff_A_mJqz6rnL6_0(.dout(w_dff_A_k5pLKUhv3_0),.din(w_dff_A_mJqz6rnL6_0),.clk(gclk));
	jdff dff_A_PDW4LpkL6_0(.dout(w_dff_A_mJqz6rnL6_0),.din(w_dff_A_PDW4LpkL6_0),.clk(gclk));
	jdff dff_A_OmW5Xfae5_0(.dout(w_dff_A_PDW4LpkL6_0),.din(w_dff_A_OmW5Xfae5_0),.clk(gclk));
	jdff dff_A_EA2hOLsY0_0(.dout(w_dff_A_OmW5Xfae5_0),.din(w_dff_A_EA2hOLsY0_0),.clk(gclk));
	jdff dff_A_WbU7slYa3_0(.dout(w_dff_A_EA2hOLsY0_0),.din(w_dff_A_WbU7slYa3_0),.clk(gclk));
	jdff dff_A_d7qouoRC9_0(.dout(w_dff_A_WbU7slYa3_0),.din(w_dff_A_d7qouoRC9_0),.clk(gclk));
	jdff dff_A_1P1smI3R2_0(.dout(w_dff_A_d7qouoRC9_0),.din(w_dff_A_1P1smI3R2_0),.clk(gclk));
	jdff dff_A_Fg6V4p2y1_0(.dout(w_dff_A_1P1smI3R2_0),.din(w_dff_A_Fg6V4p2y1_0),.clk(gclk));
	jdff dff_A_ydOLMp6N6_0(.dout(w_dff_A_Fg6V4p2y1_0),.din(w_dff_A_ydOLMp6N6_0),.clk(gclk));
	jdff dff_A_EmUjLuic3_0(.dout(w_dff_A_ydOLMp6N6_0),.din(w_dff_A_EmUjLuic3_0),.clk(gclk));
	jdff dff_A_LUvcrnHy4_0(.dout(w_dff_A_EmUjLuic3_0),.din(w_dff_A_LUvcrnHy4_0),.clk(gclk));
	jdff dff_A_QTbTcMfe2_0(.dout(w_dff_A_LUvcrnHy4_0),.din(w_dff_A_QTbTcMfe2_0),.clk(gclk));
	jdff dff_A_xjM7abYy4_0(.dout(w_dff_A_QTbTcMfe2_0),.din(w_dff_A_xjM7abYy4_0),.clk(gclk));
	jdff dff_A_g46lyfAZ5_0(.dout(w_dff_A_xjM7abYy4_0),.din(w_dff_A_g46lyfAZ5_0),.clk(gclk));
	jdff dff_A_AiEyQROX8_0(.dout(w_dff_A_g46lyfAZ5_0),.din(w_dff_A_AiEyQROX8_0),.clk(gclk));
	jdff dff_A_XEDLWGuX6_0(.dout(w_dff_A_AiEyQROX8_0),.din(w_dff_A_XEDLWGuX6_0),.clk(gclk));
	jdff dff_A_S0iiNFFp4_0(.dout(w_dff_A_XEDLWGuX6_0),.din(w_dff_A_S0iiNFFp4_0),.clk(gclk));
	jdff dff_A_sXogL2F34_0(.dout(w_dff_A_S0iiNFFp4_0),.din(w_dff_A_sXogL2F34_0),.clk(gclk));
	jdff dff_A_Hf4XiKpk9_0(.dout(w_dff_A_sXogL2F34_0),.din(w_dff_A_Hf4XiKpk9_0),.clk(gclk));
	jdff dff_A_gl02tlid9_0(.dout(w_dff_A_Hf4XiKpk9_0),.din(w_dff_A_gl02tlid9_0),.clk(gclk));
	jdff dff_A_2G7fOMRi7_0(.dout(w_dff_A_gl02tlid9_0),.din(w_dff_A_2G7fOMRi7_0),.clk(gclk));
	jdff dff_A_b9i0mVPX4_0(.dout(w_dff_A_2G7fOMRi7_0),.din(w_dff_A_b9i0mVPX4_0),.clk(gclk));
	jdff dff_A_387xNCBw7_1(.dout(w_n437_0[1]),.din(w_dff_A_387xNCBw7_1),.clk(gclk));
	jdff dff_A_mTJizaas6_1(.dout(w_dff_A_387xNCBw7_1),.din(w_dff_A_mTJizaas6_1),.clk(gclk));
	jdff dff_A_eBFFZHSR0_1(.dout(w_dff_A_mTJizaas6_1),.din(w_dff_A_eBFFZHSR0_1),.clk(gclk));
	jdff dff_A_m7l1VNKy0_1(.dout(w_dff_A_eBFFZHSR0_1),.din(w_dff_A_m7l1VNKy0_1),.clk(gclk));
	jdff dff_A_lbqrYRH56_1(.dout(w_dff_A_m7l1VNKy0_1),.din(w_dff_A_lbqrYRH56_1),.clk(gclk));
	jdff dff_A_2RPepJyl2_1(.dout(w_dff_A_lbqrYRH56_1),.din(w_dff_A_2RPepJyl2_1),.clk(gclk));
	jdff dff_A_vsDihIaw3_1(.dout(w_dff_A_2RPepJyl2_1),.din(w_dff_A_vsDihIaw3_1),.clk(gclk));
	jdff dff_A_HR0oxJQG8_1(.dout(w_dff_A_vsDihIaw3_1),.din(w_dff_A_HR0oxJQG8_1),.clk(gclk));
	jdff dff_A_euFO73gY0_1(.dout(w_dff_A_HR0oxJQG8_1),.din(w_dff_A_euFO73gY0_1),.clk(gclk));
	jdff dff_A_y5wHyyBy4_1(.dout(w_dff_A_euFO73gY0_1),.din(w_dff_A_y5wHyyBy4_1),.clk(gclk));
	jdff dff_A_bTwg9hed6_1(.dout(w_dff_A_y5wHyyBy4_1),.din(w_dff_A_bTwg9hed6_1),.clk(gclk));
	jdff dff_A_PUmlXlX87_1(.dout(w_dff_A_bTwg9hed6_1),.din(w_dff_A_PUmlXlX87_1),.clk(gclk));
	jdff dff_A_Tmg5YTKb6_1(.dout(w_dff_A_PUmlXlX87_1),.din(w_dff_A_Tmg5YTKb6_1),.clk(gclk));
	jdff dff_A_z8vE3lil5_1(.dout(w_dff_A_Tmg5YTKb6_1),.din(w_dff_A_z8vE3lil5_1),.clk(gclk));
	jdff dff_A_Uu017SPj2_1(.dout(w_dff_A_z8vE3lil5_1),.din(w_dff_A_Uu017SPj2_1),.clk(gclk));
	jdff dff_A_SMs7wOsT4_1(.dout(w_dff_A_Uu017SPj2_1),.din(w_dff_A_SMs7wOsT4_1),.clk(gclk));
	jdff dff_A_ozyoaQiE6_1(.dout(w_dff_A_SMs7wOsT4_1),.din(w_dff_A_ozyoaQiE6_1),.clk(gclk));
	jdff dff_A_ItrCI28u1_1(.dout(w_dff_A_ozyoaQiE6_1),.din(w_dff_A_ItrCI28u1_1),.clk(gclk));
	jdff dff_A_LY8xMpdE4_1(.dout(w_dff_A_ItrCI28u1_1),.din(w_dff_A_LY8xMpdE4_1),.clk(gclk));
	jdff dff_A_w6LFbHZM6_1(.dout(w_dff_A_LY8xMpdE4_1),.din(w_dff_A_w6LFbHZM6_1),.clk(gclk));
	jdff dff_A_ydoMcFHd3_1(.dout(w_dff_A_w6LFbHZM6_1),.din(w_dff_A_ydoMcFHd3_1),.clk(gclk));
	jdff dff_A_zMW1l7rV8_1(.dout(w_dff_A_ydoMcFHd3_1),.din(w_dff_A_zMW1l7rV8_1),.clk(gclk));
	jdff dff_A_pWMSAPij5_1(.dout(w_dff_A_zMW1l7rV8_1),.din(w_dff_A_pWMSAPij5_1),.clk(gclk));
	jdff dff_A_ERRnKHiM3_1(.dout(w_dff_A_pWMSAPij5_1),.din(w_dff_A_ERRnKHiM3_1),.clk(gclk));
	jdff dff_A_GVpSceM11_1(.dout(w_dff_A_ERRnKHiM3_1),.din(w_dff_A_GVpSceM11_1),.clk(gclk));
	jdff dff_A_R1lrvgxA0_1(.dout(w_dff_A_GVpSceM11_1),.din(w_dff_A_R1lrvgxA0_1),.clk(gclk));
	jdff dff_A_ixPLp55g3_0(.dout(w_n435_0[0]),.din(w_dff_A_ixPLp55g3_0),.clk(gclk));
	jdff dff_A_Dxy3LhG70_0(.dout(w_dff_A_ixPLp55g3_0),.din(w_dff_A_Dxy3LhG70_0),.clk(gclk));
	jdff dff_B_wEA3Mhyp8_0(.din(G156),.dout(w_dff_B_wEA3Mhyp8_0),.clk(gclk));
	jdff dff_B_q2wugx5I4_2(.din(n434),.dout(w_dff_B_q2wugx5I4_2),.clk(gclk));
	jdff dff_B_59IVopTg7_2(.din(w_dff_B_q2wugx5I4_2),.dout(w_dff_B_59IVopTg7_2),.clk(gclk));
	jdff dff_A_3wBuw7q61_2(.dout(w_G2239_0[2]),.din(w_dff_A_3wBuw7q61_2),.clk(gclk));
	jdff dff_A_nKOwR62T0_2(.dout(w_dff_A_3wBuw7q61_2),.din(w_dff_A_nKOwR62T0_2),.clk(gclk));
	jdff dff_A_AUMhxIV25_2(.dout(w_dff_A_nKOwR62T0_2),.din(w_dff_A_AUMhxIV25_2),.clk(gclk));
	jdff dff_A_LcmCCn9p0_2(.dout(w_dff_A_AUMhxIV25_2),.din(w_dff_A_LcmCCn9p0_2),.clk(gclk));
	jdff dff_A_pAmu6KRT6_0(.dout(w_n433_1[0]),.din(w_dff_A_pAmu6KRT6_0),.clk(gclk));
	jdff dff_A_BdNNkt7t5_0(.dout(w_dff_A_pAmu6KRT6_0),.din(w_dff_A_BdNNkt7t5_0),.clk(gclk));
	jdff dff_A_GVtHqrqw2_0(.dout(w_dff_A_BdNNkt7t5_0),.din(w_dff_A_GVtHqrqw2_0),.clk(gclk));
	jdff dff_A_zema3Pci6_0(.dout(w_dff_A_GVtHqrqw2_0),.din(w_dff_A_zema3Pci6_0),.clk(gclk));
	jdff dff_A_pbkPyzqZ3_0(.dout(w_dff_A_zema3Pci6_0),.din(w_dff_A_pbkPyzqZ3_0),.clk(gclk));
	jdff dff_A_1snCvRQM9_0(.dout(w_dff_A_pbkPyzqZ3_0),.din(w_dff_A_1snCvRQM9_0),.clk(gclk));
	jdff dff_A_fvnDjC625_0(.dout(w_dff_A_1snCvRQM9_0),.din(w_dff_A_fvnDjC625_0),.clk(gclk));
	jdff dff_A_u8A8dzar6_0(.dout(w_dff_A_fvnDjC625_0),.din(w_dff_A_u8A8dzar6_0),.clk(gclk));
	jdff dff_A_xPZ30kMI6_0(.dout(w_dff_A_u8A8dzar6_0),.din(w_dff_A_xPZ30kMI6_0),.clk(gclk));
	jdff dff_A_igY3nnvL2_0(.dout(w_dff_A_xPZ30kMI6_0),.din(w_dff_A_igY3nnvL2_0),.clk(gclk));
	jdff dff_A_F5ZTxqAJ1_0(.dout(w_dff_A_igY3nnvL2_0),.din(w_dff_A_F5ZTxqAJ1_0),.clk(gclk));
	jdff dff_A_MTgprWJy7_0(.dout(w_dff_A_F5ZTxqAJ1_0),.din(w_dff_A_MTgprWJy7_0),.clk(gclk));
	jdff dff_A_G0bKuq5s8_0(.dout(w_dff_A_MTgprWJy7_0),.din(w_dff_A_G0bKuq5s8_0),.clk(gclk));
	jdff dff_A_RYW8Liwf4_0(.dout(w_dff_A_G0bKuq5s8_0),.din(w_dff_A_RYW8Liwf4_0),.clk(gclk));
	jdff dff_A_NOoDreEn2_0(.dout(w_dff_A_RYW8Liwf4_0),.din(w_dff_A_NOoDreEn2_0),.clk(gclk));
	jdff dff_A_jnJX9vzc5_0(.dout(w_dff_A_NOoDreEn2_0),.din(w_dff_A_jnJX9vzc5_0),.clk(gclk));
	jdff dff_A_sH9JF1vV8_0(.dout(w_dff_A_jnJX9vzc5_0),.din(w_dff_A_sH9JF1vV8_0),.clk(gclk));
	jdff dff_A_NrXAo8iN2_0(.dout(w_dff_A_sH9JF1vV8_0),.din(w_dff_A_NrXAo8iN2_0),.clk(gclk));
	jdff dff_A_KCGuJm2B2_0(.dout(w_dff_A_NrXAo8iN2_0),.din(w_dff_A_KCGuJm2B2_0),.clk(gclk));
	jdff dff_A_kfLL1v7W8_0(.dout(w_dff_A_KCGuJm2B2_0),.din(w_dff_A_kfLL1v7W8_0),.clk(gclk));
	jdff dff_A_GgfWM8fP3_0(.dout(w_dff_A_kfLL1v7W8_0),.din(w_dff_A_GgfWM8fP3_0),.clk(gclk));
	jdff dff_A_Qqjm0Ki83_0(.dout(w_dff_A_GgfWM8fP3_0),.din(w_dff_A_Qqjm0Ki83_0),.clk(gclk));
	jdff dff_A_2aihjCnZ1_0(.dout(w_dff_A_Qqjm0Ki83_0),.din(w_dff_A_2aihjCnZ1_0),.clk(gclk));
	jdff dff_A_elxtFNZ21_0(.dout(w_dff_A_2aihjCnZ1_0),.din(w_dff_A_elxtFNZ21_0),.clk(gclk));
	jdff dff_A_c7ZQRUbS3_0(.dout(w_dff_A_elxtFNZ21_0),.din(w_dff_A_c7ZQRUbS3_0),.clk(gclk));
	jdff dff_A_Ar18Dr8B6_0(.dout(w_dff_A_c7ZQRUbS3_0),.din(w_dff_A_Ar18Dr8B6_0),.clk(gclk));
	jdff dff_A_cd83q31D9_0(.dout(w_dff_A_Ar18Dr8B6_0),.din(w_dff_A_cd83q31D9_0),.clk(gclk));
	jdff dff_A_OuOmfGs39_0(.dout(w_dff_A_cd83q31D9_0),.din(w_dff_A_OuOmfGs39_0),.clk(gclk));
	jdff dff_A_UYjlfQK17_2(.dout(w_n433_0[2]),.din(w_dff_A_UYjlfQK17_2),.clk(gclk));
	jdff dff_A_YLcjpomc1_2(.dout(w_dff_A_UYjlfQK17_2),.din(w_dff_A_YLcjpomc1_2),.clk(gclk));
	jdff dff_A_yvXqhH371_2(.dout(w_dff_A_YLcjpomc1_2),.din(w_dff_A_yvXqhH371_2),.clk(gclk));
	jdff dff_A_ky3EWdLW5_2(.dout(w_dff_A_yvXqhH371_2),.din(w_dff_A_ky3EWdLW5_2),.clk(gclk));
	jdff dff_A_9FBXsJ5D7_0(.dout(w_n431_0[0]),.din(w_dff_A_9FBXsJ5D7_0),.clk(gclk));
	jdff dff_A_rZYiXbkz5_0(.dout(w_dff_A_9FBXsJ5D7_0),.din(w_dff_A_rZYiXbkz5_0),.clk(gclk));
	jdff dff_B_F1xHy1Kr0_0(.din(G155),.dout(w_dff_B_F1xHy1Kr0_0),.clk(gclk));
	jdff dff_B_aLOuqT6y1_2(.din(n430),.dout(w_dff_B_aLOuqT6y1_2),.clk(gclk));
	jdff dff_B_qfxNow3q4_2(.din(w_dff_B_aLOuqT6y1_2),.dout(w_dff_B_qfxNow3q4_2),.clk(gclk));
	jdff dff_A_09Rzbv0n9_1(.dout(w_n429_0[1]),.din(w_dff_A_09Rzbv0n9_1),.clk(gclk));
	jdff dff_A_zEQnSkvr7_1(.dout(w_dff_A_09Rzbv0n9_1),.din(w_dff_A_zEQnSkvr7_1),.clk(gclk));
	jdff dff_A_xGnoXxZc2_1(.dout(w_dff_A_zEQnSkvr7_1),.din(w_dff_A_xGnoXxZc2_1),.clk(gclk));
	jdff dff_A_sg9lbXIo8_1(.dout(w_dff_A_xGnoXxZc2_1),.din(w_dff_A_sg9lbXIo8_1),.clk(gclk));
	jdff dff_A_H6LTrRNq3_1(.dout(w_dff_A_sg9lbXIo8_1),.din(w_dff_A_H6LTrRNq3_1),.clk(gclk));
	jdff dff_A_suG4h3MQ2_1(.dout(w_dff_A_H6LTrRNq3_1),.din(w_dff_A_suG4h3MQ2_1),.clk(gclk));
	jdff dff_A_XwqpMb7r3_1(.dout(w_dff_A_suG4h3MQ2_1),.din(w_dff_A_XwqpMb7r3_1),.clk(gclk));
	jdff dff_A_gr4pZuZk5_1(.dout(w_dff_A_XwqpMb7r3_1),.din(w_dff_A_gr4pZuZk5_1),.clk(gclk));
	jdff dff_A_Zezn3gTG3_1(.dout(w_dff_A_gr4pZuZk5_1),.din(w_dff_A_Zezn3gTG3_1),.clk(gclk));
	jdff dff_A_79D3nSYZ5_1(.dout(w_dff_A_Zezn3gTG3_1),.din(w_dff_A_79D3nSYZ5_1),.clk(gclk));
	jdff dff_A_0m4mJ7o25_1(.dout(w_dff_A_79D3nSYZ5_1),.din(w_dff_A_0m4mJ7o25_1),.clk(gclk));
	jdff dff_A_RMSrkFxh6_1(.dout(w_dff_A_0m4mJ7o25_1),.din(w_dff_A_RMSrkFxh6_1),.clk(gclk));
	jdff dff_A_CmqjsdPN6_1(.dout(w_dff_A_RMSrkFxh6_1),.din(w_dff_A_CmqjsdPN6_1),.clk(gclk));
	jdff dff_A_fll1kGTT8_1(.dout(w_dff_A_CmqjsdPN6_1),.din(w_dff_A_fll1kGTT8_1),.clk(gclk));
	jdff dff_A_4E0of3rE9_1(.dout(w_dff_A_fll1kGTT8_1),.din(w_dff_A_4E0of3rE9_1),.clk(gclk));
	jdff dff_A_moFGrM1t2_1(.dout(w_dff_A_4E0of3rE9_1),.din(w_dff_A_moFGrM1t2_1),.clk(gclk));
	jdff dff_A_Mjxs4LXI1_1(.dout(w_dff_A_moFGrM1t2_1),.din(w_dff_A_Mjxs4LXI1_1),.clk(gclk));
	jdff dff_A_36A6DOYl2_1(.dout(w_dff_A_Mjxs4LXI1_1),.din(w_dff_A_36A6DOYl2_1),.clk(gclk));
	jdff dff_A_zF5Nd7pD3_1(.dout(w_dff_A_36A6DOYl2_1),.din(w_dff_A_zF5Nd7pD3_1),.clk(gclk));
	jdff dff_A_RwvSeBfy3_1(.dout(w_dff_A_zF5Nd7pD3_1),.din(w_dff_A_RwvSeBfy3_1),.clk(gclk));
	jdff dff_A_5gnAqyom9_1(.dout(w_dff_A_RwvSeBfy3_1),.din(w_dff_A_5gnAqyom9_1),.clk(gclk));
	jdff dff_A_DhltJnR27_1(.dout(w_dff_A_5gnAqyom9_1),.din(w_dff_A_DhltJnR27_1),.clk(gclk));
	jdff dff_A_cPYjnrig9_1(.dout(w_dff_A_DhltJnR27_1),.din(w_dff_A_cPYjnrig9_1),.clk(gclk));
	jdff dff_A_hrEXM8FB1_1(.dout(w_dff_A_cPYjnrig9_1),.din(w_dff_A_hrEXM8FB1_1),.clk(gclk));
	jdff dff_A_xddUA2Jw4_1(.dout(w_dff_A_hrEXM8FB1_1),.din(w_dff_A_xddUA2Jw4_1),.clk(gclk));
	jdff dff_A_cXhmlniw5_1(.dout(w_dff_A_xddUA2Jw4_1),.din(w_dff_A_cXhmlniw5_1),.clk(gclk));
	jdff dff_A_1Ymh6j8A3_1(.dout(w_dff_A_cXhmlniw5_1),.din(w_dff_A_1Ymh6j8A3_1),.clk(gclk));
	jdff dff_A_YUTW2DAO3_1(.dout(w_dff_A_1Ymh6j8A3_1),.din(w_dff_A_YUTW2DAO3_1),.clk(gclk));
	jdff dff_A_9gVNd9nX7_2(.dout(w_n429_0[2]),.din(w_dff_A_9gVNd9nX7_2),.clk(gclk));
	jdff dff_A_4arLlfmD9_0(.dout(w_n427_0[0]),.din(w_dff_A_4arLlfmD9_0),.clk(gclk));
	jdff dff_A_Etqypq3F7_0(.dout(w_dff_A_4arLlfmD9_0),.din(w_dff_A_Etqypq3F7_0),.clk(gclk));
	jdff dff_B_8UG59Vca7_0(.din(G154),.dout(w_dff_B_8UG59Vca7_0),.clk(gclk));
	jdff dff_A_QX1Bx6I01_1(.dout(w_n426_0[1]),.din(w_dff_A_QX1Bx6I01_1),.clk(gclk));
	jdff dff_A_Ggj1yM443_1(.dout(w_dff_A_QX1Bx6I01_1),.din(w_dff_A_Ggj1yM443_1),.clk(gclk));
	jdff dff_A_HTMGDVHZ1_2(.dout(w_n426_0[2]),.din(w_dff_A_HTMGDVHZ1_2),.clk(gclk));
	jdff dff_A_K5ZBCKeC9_2(.dout(w_dff_A_HTMGDVHZ1_2),.din(w_dff_A_K5ZBCKeC9_2),.clk(gclk));
	jdff dff_A_DY0byoKN3_1(.dout(w_G2253_0[1]),.din(w_dff_A_DY0byoKN3_1),.clk(gclk));
	jdff dff_A_poaqWqFO4_1(.dout(w_dff_A_DY0byoKN3_1),.din(w_dff_A_poaqWqFO4_1),.clk(gclk));
	jdff dff_A_otUmM6eA6_1(.dout(w_dff_A_poaqWqFO4_1),.din(w_dff_A_otUmM6eA6_1),.clk(gclk));
	jdff dff_A_Pn0AJcb18_1(.dout(w_dff_A_otUmM6eA6_1),.din(w_dff_A_Pn0AJcb18_1),.clk(gclk));
	jdff dff_A_baD3Q3CB8_1(.dout(w_n425_1[1]),.din(w_dff_A_baD3Q3CB8_1),.clk(gclk));
	jdff dff_A_1R9bhMXu3_1(.dout(w_dff_A_baD3Q3CB8_1),.din(w_dff_A_1R9bhMXu3_1),.clk(gclk));
	jdff dff_A_wWKFtqNt8_1(.dout(w_dff_A_1R9bhMXu3_1),.din(w_dff_A_wWKFtqNt8_1),.clk(gclk));
	jdff dff_A_71pj1lpB6_1(.dout(w_dff_A_wWKFtqNt8_1),.din(w_dff_A_71pj1lpB6_1),.clk(gclk));
	jdff dff_A_ryRSPHHA3_1(.dout(w_dff_A_71pj1lpB6_1),.din(w_dff_A_ryRSPHHA3_1),.clk(gclk));
	jdff dff_A_KavIGZoi1_1(.dout(w_dff_A_ryRSPHHA3_1),.din(w_dff_A_KavIGZoi1_1),.clk(gclk));
	jdff dff_A_OjjPaYin5_1(.dout(w_dff_A_KavIGZoi1_1),.din(w_dff_A_OjjPaYin5_1),.clk(gclk));
	jdff dff_A_49iVaXPm4_1(.dout(w_dff_A_OjjPaYin5_1),.din(w_dff_A_49iVaXPm4_1),.clk(gclk));
	jdff dff_A_uL3r89oo2_1(.dout(w_dff_A_49iVaXPm4_1),.din(w_dff_A_uL3r89oo2_1),.clk(gclk));
	jdff dff_A_K5wvCeqg4_1(.dout(w_dff_A_uL3r89oo2_1),.din(w_dff_A_K5wvCeqg4_1),.clk(gclk));
	jdff dff_A_8GZUAg3f1_1(.dout(w_dff_A_K5wvCeqg4_1),.din(w_dff_A_8GZUAg3f1_1),.clk(gclk));
	jdff dff_A_y6Lu6vUt2_1(.dout(w_dff_A_8GZUAg3f1_1),.din(w_dff_A_y6Lu6vUt2_1),.clk(gclk));
	jdff dff_A_yWVwfS0b3_1(.dout(w_dff_A_y6Lu6vUt2_1),.din(w_dff_A_yWVwfS0b3_1),.clk(gclk));
	jdff dff_A_uSkAOhDH6_1(.dout(w_dff_A_yWVwfS0b3_1),.din(w_dff_A_uSkAOhDH6_1),.clk(gclk));
	jdff dff_A_yh9jPnZQ7_1(.dout(w_dff_A_uSkAOhDH6_1),.din(w_dff_A_yh9jPnZQ7_1),.clk(gclk));
	jdff dff_A_CAjnkr406_1(.dout(w_dff_A_yh9jPnZQ7_1),.din(w_dff_A_CAjnkr406_1),.clk(gclk));
	jdff dff_A_bZpG9w7x0_1(.dout(w_dff_A_CAjnkr406_1),.din(w_dff_A_bZpG9w7x0_1),.clk(gclk));
	jdff dff_A_3nTGLdvQ8_1(.dout(w_dff_A_bZpG9w7x0_1),.din(w_dff_A_3nTGLdvQ8_1),.clk(gclk));
	jdff dff_A_Tqr5ye7V0_1(.dout(w_dff_A_3nTGLdvQ8_1),.din(w_dff_A_Tqr5ye7V0_1),.clk(gclk));
	jdff dff_A_MrxSu1Kd1_1(.dout(w_dff_A_Tqr5ye7V0_1),.din(w_dff_A_MrxSu1Kd1_1),.clk(gclk));
	jdff dff_A_z8TgFc517_1(.dout(w_dff_A_MrxSu1Kd1_1),.din(w_dff_A_z8TgFc517_1),.clk(gclk));
	jdff dff_A_iYFIVBXd1_1(.dout(w_dff_A_z8TgFc517_1),.din(w_dff_A_iYFIVBXd1_1),.clk(gclk));
	jdff dff_A_CKmlYBeT8_1(.dout(w_dff_A_iYFIVBXd1_1),.din(w_dff_A_CKmlYBeT8_1),.clk(gclk));
	jdff dff_A_Lq8qeYY98_1(.dout(w_dff_A_CKmlYBeT8_1),.din(w_dff_A_Lq8qeYY98_1),.clk(gclk));
	jdff dff_A_AY0Ygbpn0_1(.dout(w_dff_A_Lq8qeYY98_1),.din(w_dff_A_AY0Ygbpn0_1),.clk(gclk));
	jdff dff_A_tR2DfjdY3_1(.dout(w_dff_A_AY0Ygbpn0_1),.din(w_dff_A_tR2DfjdY3_1),.clk(gclk));
	jdff dff_A_udk0DvfK8_1(.dout(w_dff_A_tR2DfjdY3_1),.din(w_dff_A_udk0DvfK8_1),.clk(gclk));
	jdff dff_A_fHouZqGt3_1(.dout(w_dff_A_udk0DvfK8_1),.din(w_dff_A_fHouZqGt3_1),.clk(gclk));
	jdff dff_A_C5gFqW8C7_2(.dout(w_n425_0[2]),.din(w_dff_A_C5gFqW8C7_2),.clk(gclk));
	jdff dff_A_AzhajSGA9_2(.dout(w_dff_A_C5gFqW8C7_2),.din(w_dff_A_AzhajSGA9_2),.clk(gclk));
	jdff dff_A_anWRxKrp5_2(.dout(w_dff_A_AzhajSGA9_2),.din(w_dff_A_anWRxKrp5_2),.clk(gclk));
	jdff dff_A_CEBS9loZ4_2(.dout(w_dff_A_anWRxKrp5_2),.din(w_dff_A_CEBS9loZ4_2),.clk(gclk));
	jdff dff_A_zWpz9K373_2(.dout(w_dff_A_CEBS9loZ4_2),.din(w_dff_A_zWpz9K373_2),.clk(gclk));
	jdff dff_A_tS34ImiE8_2(.dout(w_dff_A_zWpz9K373_2),.din(w_dff_A_tS34ImiE8_2),.clk(gclk));
	jdff dff_A_i9BEr20I3_2(.dout(w_dff_A_tS34ImiE8_2),.din(w_dff_A_i9BEr20I3_2),.clk(gclk));
	jdff dff_A_6BNDKbQJ5_2(.dout(w_dff_A_i9BEr20I3_2),.din(w_dff_A_6BNDKbQJ5_2),.clk(gclk));
	jdff dff_A_wHvaS5eP5_2(.dout(w_dff_A_6BNDKbQJ5_2),.din(w_dff_A_wHvaS5eP5_2),.clk(gclk));
	jdff dff_A_2UJBnGw15_2(.dout(w_dff_A_wHvaS5eP5_2),.din(w_dff_A_2UJBnGw15_2),.clk(gclk));
	jdff dff_A_YHYPlSnV9_2(.dout(w_dff_A_2UJBnGw15_2),.din(w_dff_A_YHYPlSnV9_2),.clk(gclk));
	jdff dff_A_NmpRpQDc7_2(.dout(w_dff_A_YHYPlSnV9_2),.din(w_dff_A_NmpRpQDc7_2),.clk(gclk));
	jdff dff_A_IIb8Gdv16_2(.dout(w_dff_A_NmpRpQDc7_2),.din(w_dff_A_IIb8Gdv16_2),.clk(gclk));
	jdff dff_A_QwKkJGS42_2(.dout(w_dff_A_IIb8Gdv16_2),.din(w_dff_A_QwKkJGS42_2),.clk(gclk));
	jdff dff_A_FpE1NfNw5_2(.dout(w_dff_A_QwKkJGS42_2),.din(w_dff_A_FpE1NfNw5_2),.clk(gclk));
	jdff dff_A_ZAXYdkzJ8_2(.dout(w_dff_A_FpE1NfNw5_2),.din(w_dff_A_ZAXYdkzJ8_2),.clk(gclk));
	jdff dff_A_b3I5VCR79_2(.dout(w_dff_A_ZAXYdkzJ8_2),.din(w_dff_A_b3I5VCR79_2),.clk(gclk));
	jdff dff_A_M8tnH8qC1_2(.dout(w_dff_A_b3I5VCR79_2),.din(w_dff_A_M8tnH8qC1_2),.clk(gclk));
	jdff dff_A_TzFzFNrV6_2(.dout(w_dff_A_M8tnH8qC1_2),.din(w_dff_A_TzFzFNrV6_2),.clk(gclk));
	jdff dff_A_xkqkMJMN6_2(.dout(w_dff_A_TzFzFNrV6_2),.din(w_dff_A_xkqkMJMN6_2),.clk(gclk));
	jdff dff_A_jvauE3K24_2(.dout(w_dff_A_xkqkMJMN6_2),.din(w_dff_A_jvauE3K24_2),.clk(gclk));
	jdff dff_A_QQKBQqh65_2(.dout(w_dff_A_jvauE3K24_2),.din(w_dff_A_QQKBQqh65_2),.clk(gclk));
	jdff dff_A_tUUVP2Vy9_2(.dout(w_dff_A_QQKBQqh65_2),.din(w_dff_A_tUUVP2Vy9_2),.clk(gclk));
	jdff dff_A_BHs6HxvU7_2(.dout(w_dff_A_tUUVP2Vy9_2),.din(w_dff_A_BHs6HxvU7_2),.clk(gclk));
	jdff dff_A_VmcHDvd72_2(.dout(w_dff_A_BHs6HxvU7_2),.din(w_dff_A_VmcHDvd72_2),.clk(gclk));
	jdff dff_A_U6iUWgwA8_2(.dout(w_dff_A_VmcHDvd72_2),.din(w_dff_A_U6iUWgwA8_2),.clk(gclk));
	jdff dff_A_FNcJlQLL3_2(.dout(w_dff_A_U6iUWgwA8_2),.din(w_dff_A_FNcJlQLL3_2),.clk(gclk));
	jdff dff_A_wqPvJ2r96_2(.dout(w_dff_A_FNcJlQLL3_2),.din(w_dff_A_wqPvJ2r96_2),.clk(gclk));
	jdff dff_A_JPCot2ZB7_1(.dout(w_n424_0[1]),.din(w_dff_A_JPCot2ZB7_1),.clk(gclk));
	jdff dff_A_L7qavIXQ2_1(.dout(w_dff_A_JPCot2ZB7_1),.din(w_dff_A_L7qavIXQ2_1),.clk(gclk));
	jdff dff_A_AbUAfjVv8_1(.dout(w_dff_A_L7qavIXQ2_1),.din(w_dff_A_AbUAfjVv8_1),.clk(gclk));
	jdff dff_A_0vjlAh087_1(.dout(w_dff_A_AbUAfjVv8_1),.din(w_dff_A_0vjlAh087_1),.clk(gclk));
	jdff dff_A_rbzNotZQ9_1(.dout(w_dff_A_0vjlAh087_1),.din(w_dff_A_rbzNotZQ9_1),.clk(gclk));
	jdff dff_A_LIx7qTrD6_1(.dout(w_dff_A_rbzNotZQ9_1),.din(w_dff_A_LIx7qTrD6_1),.clk(gclk));
	jdff dff_A_TH2h2Jyo1_1(.dout(w_dff_A_LIx7qTrD6_1),.din(w_dff_A_TH2h2Jyo1_1),.clk(gclk));
	jdff dff_A_63KIUd6P4_1(.dout(w_dff_A_TH2h2Jyo1_1),.din(w_dff_A_63KIUd6P4_1),.clk(gclk));
	jdff dff_A_LytSijHB7_1(.dout(w_dff_A_63KIUd6P4_1),.din(w_dff_A_LytSijHB7_1),.clk(gclk));
	jdff dff_A_T6Pw4CQE5_1(.dout(w_dff_A_LytSijHB7_1),.din(w_dff_A_T6Pw4CQE5_1),.clk(gclk));
	jdff dff_A_FecUEcXq0_1(.dout(w_dff_A_T6Pw4CQE5_1),.din(w_dff_A_FecUEcXq0_1),.clk(gclk));
	jdff dff_A_jfqI3rik3_1(.dout(w_dff_A_FecUEcXq0_1),.din(w_dff_A_jfqI3rik3_1),.clk(gclk));
	jdff dff_A_2VydCtZr7_1(.dout(w_dff_A_jfqI3rik3_1),.din(w_dff_A_2VydCtZr7_1),.clk(gclk));
	jdff dff_A_RwDE5Bnv0_1(.dout(w_dff_A_2VydCtZr7_1),.din(w_dff_A_RwDE5Bnv0_1),.clk(gclk));
	jdff dff_A_3wkFOEgy6_1(.dout(w_dff_A_RwDE5Bnv0_1),.din(w_dff_A_3wkFOEgy6_1),.clk(gclk));
	jdff dff_A_r1jNPOol5_1(.dout(w_dff_A_3wkFOEgy6_1),.din(w_dff_A_r1jNPOol5_1),.clk(gclk));
	jdff dff_A_qv6uDbQW6_1(.dout(w_dff_A_r1jNPOol5_1),.din(w_dff_A_qv6uDbQW6_1),.clk(gclk));
	jdff dff_A_IxbBvkpg9_1(.dout(w_dff_A_qv6uDbQW6_1),.din(w_dff_A_IxbBvkpg9_1),.clk(gclk));
	jdff dff_A_nM5uXi1V4_1(.dout(w_dff_A_IxbBvkpg9_1),.din(w_dff_A_nM5uXi1V4_1),.clk(gclk));
	jdff dff_A_xs1WsFzi4_1(.dout(w_dff_A_nM5uXi1V4_1),.din(w_dff_A_xs1WsFzi4_1),.clk(gclk));
	jdff dff_A_h2OQWkcC5_1(.dout(w_dff_A_xs1WsFzi4_1),.din(w_dff_A_h2OQWkcC5_1),.clk(gclk));
	jdff dff_A_ZW4vS40h0_1(.dout(w_dff_A_h2OQWkcC5_1),.din(w_dff_A_ZW4vS40h0_1),.clk(gclk));
	jdff dff_A_BrYgqhBT2_1(.dout(w_dff_A_ZW4vS40h0_1),.din(w_dff_A_BrYgqhBT2_1),.clk(gclk));
	jdff dff_A_WVcPQJbm0_1(.dout(w_dff_A_BrYgqhBT2_1),.din(w_dff_A_WVcPQJbm0_1),.clk(gclk));
	jdff dff_A_lFLkfp0b5_1(.dout(w_dff_A_WVcPQJbm0_1),.din(w_dff_A_lFLkfp0b5_1),.clk(gclk));
	jdff dff_A_y8sCxpDE5_1(.dout(w_dff_A_lFLkfp0b5_1),.din(w_dff_A_y8sCxpDE5_1),.clk(gclk));
	jdff dff_A_vKkxQUhC6_1(.dout(w_dff_A_y8sCxpDE5_1),.din(w_dff_A_vKkxQUhC6_1),.clk(gclk));
	jdff dff_A_mXJSl3Zk9_1(.dout(w_dff_A_vKkxQUhC6_1),.din(w_dff_A_mXJSl3Zk9_1),.clk(gclk));
	jdff dff_A_6GHje0Ez4_1(.dout(w_dff_A_mXJSl3Zk9_1),.din(w_dff_A_6GHje0Ez4_1),.clk(gclk));
	jdff dff_A_HvRZD6YI7_0(.dout(w_n422_0[0]),.din(w_dff_A_HvRZD6YI7_0),.clk(gclk));
	jdff dff_A_3oLcbMUW2_0(.dout(w_dff_A_HvRZD6YI7_0),.din(w_dff_A_3oLcbMUW2_0),.clk(gclk));
	jdff dff_B_KrwkUrhI8_0(.din(G153),.dout(w_dff_B_KrwkUrhI8_0),.clk(gclk));
	jdff dff_A_GKk1bp1A7_1(.dout(w_n421_0[1]),.din(w_dff_A_GKk1bp1A7_1),.clk(gclk));
	jdff dff_A_J5y6YU0r4_1(.dout(w_dff_A_GKk1bp1A7_1),.din(w_dff_A_J5y6YU0r4_1),.clk(gclk));
	jdff dff_A_dIpyqVQs2_2(.dout(w_n421_0[2]),.din(w_dff_A_dIpyqVQs2_2),.clk(gclk));
	jdff dff_A_fzPZDmtX3_2(.dout(w_dff_A_dIpyqVQs2_2),.din(w_dff_A_fzPZDmtX3_2),.clk(gclk));
	jdff dff_A_bUrptudo5_1(.dout(w_n416_0[1]),.din(w_dff_A_bUrptudo5_1),.clk(gclk));
	jdff dff_A_aAH0WpaF9_1(.dout(w_dff_A_bUrptudo5_1),.din(w_dff_A_aAH0WpaF9_1),.clk(gclk));
	jdff dff_A_lNPuLJKy0_1(.dout(w_dff_A_aAH0WpaF9_1),.din(w_dff_A_lNPuLJKy0_1),.clk(gclk));
	jdff dff_A_8RIx3fbU2_1(.dout(w_dff_A_lNPuLJKy0_1),.din(w_dff_A_8RIx3fbU2_1),.clk(gclk));
	jdff dff_A_40hxMOXx5_1(.dout(w_dff_A_8RIx3fbU2_1),.din(w_dff_A_40hxMOXx5_1),.clk(gclk));
	jdff dff_A_Tfq0k3aS0_1(.dout(w_dff_A_40hxMOXx5_1),.din(w_dff_A_Tfq0k3aS0_1),.clk(gclk));
	jdff dff_A_rLdU8sJG5_1(.dout(w_dff_A_Tfq0k3aS0_1),.din(w_dff_A_rLdU8sJG5_1),.clk(gclk));
	jdff dff_A_GsibDraX6_1(.dout(w_dff_A_rLdU8sJG5_1),.din(w_dff_A_GsibDraX6_1),.clk(gclk));
	jdff dff_A_QlKpmL7l1_1(.dout(w_dff_A_GsibDraX6_1),.din(w_dff_A_QlKpmL7l1_1),.clk(gclk));
	jdff dff_A_idxDFid54_1(.dout(w_dff_A_QlKpmL7l1_1),.din(w_dff_A_idxDFid54_1),.clk(gclk));
	jdff dff_A_pFynIBHc3_1(.dout(w_dff_A_idxDFid54_1),.din(w_dff_A_pFynIBHc3_1),.clk(gclk));
	jdff dff_A_KylSvzqG0_1(.dout(w_dff_A_pFynIBHc3_1),.din(w_dff_A_KylSvzqG0_1),.clk(gclk));
	jdff dff_A_JRn941Bw9_1(.dout(w_dff_A_KylSvzqG0_1),.din(w_dff_A_JRn941Bw9_1),.clk(gclk));
	jdff dff_A_hnYhUgvT6_1(.dout(w_dff_A_JRn941Bw9_1),.din(w_dff_A_hnYhUgvT6_1),.clk(gclk));
	jdff dff_A_bKtJ0jLs3_1(.dout(w_dff_A_hnYhUgvT6_1),.din(w_dff_A_bKtJ0jLs3_1),.clk(gclk));
	jdff dff_A_Lf6bnXpT7_1(.dout(w_dff_A_bKtJ0jLs3_1),.din(w_dff_A_Lf6bnXpT7_1),.clk(gclk));
	jdff dff_A_EsfkNbea7_1(.dout(w_dff_A_Lf6bnXpT7_1),.din(w_dff_A_EsfkNbea7_1),.clk(gclk));
	jdff dff_A_eRFKiswX8_1(.dout(w_dff_A_EsfkNbea7_1),.din(w_dff_A_eRFKiswX8_1),.clk(gclk));
	jdff dff_A_sHTJBg2x2_1(.dout(w_dff_A_eRFKiswX8_1),.din(w_dff_A_sHTJBg2x2_1),.clk(gclk));
	jdff dff_A_zBdsHkwr0_1(.dout(w_dff_A_sHTJBg2x2_1),.din(w_dff_A_zBdsHkwr0_1),.clk(gclk));
	jdff dff_A_24gcnJs55_1(.dout(w_dff_A_zBdsHkwr0_1),.din(w_dff_A_24gcnJs55_1),.clk(gclk));
	jdff dff_A_2yoa0Xmg3_1(.dout(w_dff_A_24gcnJs55_1),.din(w_dff_A_2yoa0Xmg3_1),.clk(gclk));
	jdff dff_A_I5NxoADI0_1(.dout(w_dff_A_2yoa0Xmg3_1),.din(w_dff_A_I5NxoADI0_1),.clk(gclk));
	jdff dff_A_dWsgIMZl3_1(.dout(w_dff_A_I5NxoADI0_1),.din(w_dff_A_dWsgIMZl3_1),.clk(gclk));
	jdff dff_A_W9XIvgWl1_1(.dout(w_dff_A_dWsgIMZl3_1),.din(w_dff_A_W9XIvgWl1_1),.clk(gclk));
	jdff dff_A_5avsFQRR6_1(.dout(w_dff_A_W9XIvgWl1_1),.din(w_dff_A_5avsFQRR6_1),.clk(gclk));
	jdff dff_A_huoydXMQ2_1(.dout(w_dff_A_5avsFQRR6_1),.din(w_dff_A_huoydXMQ2_1),.clk(gclk));
	jdff dff_A_hYt7MMz02_1(.dout(w_dff_A_huoydXMQ2_1),.din(w_dff_A_hYt7MMz02_1),.clk(gclk));
	jdff dff_A_NlVCp1mj4_1(.dout(w_dff_A_hYt7MMz02_1),.din(w_dff_A_NlVCp1mj4_1),.clk(gclk));
	jdff dff_A_O4cQ5JZr6_1(.dout(w_dff_A_NlVCp1mj4_1),.din(w_dff_A_O4cQ5JZr6_1),.clk(gclk));
	jdff dff_A_SKbTFCZj2_1(.dout(w_dff_A_O4cQ5JZr6_1),.din(w_dff_A_SKbTFCZj2_1),.clk(gclk));
	jdff dff_A_1zVdYsML7_1(.dout(w_dff_A_SKbTFCZj2_1),.din(w_dff_A_1zVdYsML7_1),.clk(gclk));
	jdff dff_A_rGde2L1r5_0(.dout(w_n378_0[0]),.din(w_dff_A_rGde2L1r5_0),.clk(gclk));
	jdff dff_A_zj7Wtcb85_0(.dout(w_dff_A_rGde2L1r5_0),.din(w_dff_A_zj7Wtcb85_0),.clk(gclk));
	jdff dff_B_vxvT3Qbl3_0(.din(G214),.dout(w_dff_B_vxvT3Qbl3_0),.clk(gclk));
	jdff dff_A_ZmpSsmGr0_1(.dout(w_n383_0[1]),.din(w_dff_A_ZmpSsmGr0_1),.clk(gclk));
	jdff dff_A_DY0VH9bL9_1(.dout(w_dff_A_ZmpSsmGr0_1),.din(w_dff_A_DY0VH9bL9_1),.clk(gclk));
	jdff dff_A_w1WJmkCq5_2(.dout(w_n383_0[2]),.din(w_dff_A_w1WJmkCq5_2),.clk(gclk));
	jdff dff_A_4u7xADtA8_2(.dout(w_dff_A_w1WJmkCq5_2),.din(w_dff_A_4u7xADtA8_2),.clk(gclk));
	jdff dff_A_ob5eTzHp9_2(.dout(w_G1480_0[2]),.din(w_dff_A_ob5eTzHp9_2),.clk(gclk));
	jdff dff_A_3RoiRSzn7_2(.dout(w_dff_A_ob5eTzHp9_2),.din(w_dff_A_3RoiRSzn7_2),.clk(gclk));
	jdff dff_A_1guXg5S94_2(.dout(w_dff_A_3RoiRSzn7_2),.din(w_dff_A_1guXg5S94_2),.clk(gclk));
	jdff dff_A_lACnqkSy8_2(.dout(w_dff_A_1guXg5S94_2),.din(w_dff_A_lACnqkSy8_2),.clk(gclk));
	jdff dff_B_ZagUfvbl0_0(.din(G215),.dout(w_dff_B_ZagUfvbl0_0),.clk(gclk));
	jdff dff_B_wPxDIRJ71_2(.din(n385),.dout(w_dff_B_wPxDIRJ71_2),.clk(gclk));
	jdff dff_B_8TkpM3NK2_2(.din(w_dff_B_wPxDIRJ71_2),.dout(w_dff_B_8TkpM3NK2_2),.clk(gclk));
	jdff dff_A_hV1GeVxG4_0(.dout(w_G106_1[0]),.din(w_dff_A_hV1GeVxG4_0),.clk(gclk));
	jdff dff_A_B1dGCImi7_0(.dout(w_dff_A_hV1GeVxG4_0),.din(w_dff_A_B1dGCImi7_0),.clk(gclk));
	jdff dff_A_jwPzA63V8_0(.dout(w_dff_A_B1dGCImi7_0),.din(w_dff_A_jwPzA63V8_0),.clk(gclk));
	jdff dff_A_Ooh0LBXd5_0(.dout(w_dff_A_jwPzA63V8_0),.din(w_dff_A_Ooh0LBXd5_0),.clk(gclk));
	jdff dff_B_03bsOFBl3_1(.din(n1551),.dout(w_dff_B_03bsOFBl3_1),.clk(gclk));
	jdff dff_B_65zW7JSU8_1(.din(n1552),.dout(w_dff_B_65zW7JSU8_1),.clk(gclk));
	jdff dff_B_dDmxprc12_1(.din(w_dff_B_65zW7JSU8_1),.dout(w_dff_B_dDmxprc12_1),.clk(gclk));
	jdff dff_B_3SWdjrQz8_1(.din(w_dff_B_dDmxprc12_1),.dout(w_dff_B_3SWdjrQz8_1),.clk(gclk));
	jdff dff_B_lEXq7Dmk5_1(.din(w_dff_B_3SWdjrQz8_1),.dout(w_dff_B_lEXq7Dmk5_1),.clk(gclk));
	jdff dff_B_q2YQNKPl0_1(.din(w_dff_B_lEXq7Dmk5_1),.dout(w_dff_B_q2YQNKPl0_1),.clk(gclk));
	jdff dff_B_84g7pzSx1_1(.din(w_dff_B_q2YQNKPl0_1),.dout(w_dff_B_84g7pzSx1_1),.clk(gclk));
	jdff dff_B_UsAZKtNS6_1(.din(w_dff_B_84g7pzSx1_1),.dout(w_dff_B_UsAZKtNS6_1),.clk(gclk));
	jdff dff_B_7H7EWBKK6_1(.din(w_dff_B_UsAZKtNS6_1),.dout(w_dff_B_7H7EWBKK6_1),.clk(gclk));
	jdff dff_B_C6KzTMwc7_1(.din(w_dff_B_7H7EWBKK6_1),.dout(w_dff_B_C6KzTMwc7_1),.clk(gclk));
	jdff dff_B_r0ROCC9s4_1(.din(w_dff_B_C6KzTMwc7_1),.dout(w_dff_B_r0ROCC9s4_1),.clk(gclk));
	jdff dff_B_IjIqbyHH4_1(.din(w_dff_B_r0ROCC9s4_1),.dout(w_dff_B_IjIqbyHH4_1),.clk(gclk));
	jdff dff_B_flmF78nX9_1(.din(w_dff_B_IjIqbyHH4_1),.dout(w_dff_B_flmF78nX9_1),.clk(gclk));
	jdff dff_B_aofrh8mi9_1(.din(w_dff_B_flmF78nX9_1),.dout(w_dff_B_aofrh8mi9_1),.clk(gclk));
	jdff dff_B_c6sAlVSH7_1(.din(w_dff_B_aofrh8mi9_1),.dout(w_dff_B_c6sAlVSH7_1),.clk(gclk));
	jdff dff_B_sqaBfIcu0_0(.din(n1576),.dout(w_dff_B_sqaBfIcu0_0),.clk(gclk));
	jdff dff_B_Ao6mYGi31_0(.din(w_dff_B_sqaBfIcu0_0),.dout(w_dff_B_Ao6mYGi31_0),.clk(gclk));
	jdff dff_B_UuW7iBjA1_0(.din(w_dff_B_Ao6mYGi31_0),.dout(w_dff_B_UuW7iBjA1_0),.clk(gclk));
	jdff dff_B_zXwjkqDF0_0(.din(w_dff_B_UuW7iBjA1_0),.dout(w_dff_B_zXwjkqDF0_0),.clk(gclk));
	jdff dff_B_WYToY6Qz7_0(.din(n1575),.dout(w_dff_B_WYToY6Qz7_0),.clk(gclk));
	jdff dff_B_iiTVZbst1_0(.din(w_dff_B_WYToY6Qz7_0),.dout(w_dff_B_iiTVZbst1_0),.clk(gclk));
	jdff dff_B_dWg3EtNZ9_0(.din(n1572),.dout(w_dff_B_dWg3EtNZ9_0),.clk(gclk));
	jdff dff_B_2ddakiyz8_0(.din(w_dff_B_dWg3EtNZ9_0),.dout(w_dff_B_2ddakiyz8_0),.clk(gclk));
	jdff dff_B_23s7cY9T8_0(.din(w_dff_B_2ddakiyz8_0),.dout(w_dff_B_23s7cY9T8_0),.clk(gclk));
	jdff dff_B_v0dM5hOn8_0(.din(n1568),.dout(w_dff_B_v0dM5hOn8_0),.clk(gclk));
	jdff dff_B_qgka1V8r4_0(.din(w_dff_B_v0dM5hOn8_0),.dout(w_dff_B_qgka1V8r4_0),.clk(gclk));
	jdff dff_B_cVuH9BZP5_1(.din(n1560),.dout(w_dff_B_cVuH9BZP5_1),.clk(gclk));
	jdff dff_B_USdYKckw6_1(.din(w_dff_B_cVuH9BZP5_1),.dout(w_dff_B_USdYKckw6_1),.clk(gclk));
	jdff dff_B_uWWG181A2_0(.din(n1563),.dout(w_dff_B_uWWG181A2_0),.clk(gclk));
	jdff dff_B_rnq9dnf40_0(.din(w_dff_B_uWWG181A2_0),.dout(w_dff_B_rnq9dnf40_0),.clk(gclk));
	jdff dff_B_aqxciPkK8_0(.din(w_dff_B_rnq9dnf40_0),.dout(w_dff_B_aqxciPkK8_0),.clk(gclk));
	jdff dff_B_zcygb30n6_0(.din(w_dff_B_aqxciPkK8_0),.dout(w_dff_B_zcygb30n6_0),.clk(gclk));
	jdff dff_B_jjk4JYtM5_0(.din(w_dff_B_zcygb30n6_0),.dout(w_dff_B_jjk4JYtM5_0),.clk(gclk));
	jdff dff_B_mORKMFCh6_0(.din(w_dff_B_jjk4JYtM5_0),.dout(w_dff_B_mORKMFCh6_0),.clk(gclk));
	jdff dff_B_zwd4YUXK8_0(.din(w_dff_B_mORKMFCh6_0),.dout(w_dff_B_zwd4YUXK8_0),.clk(gclk));
	jdff dff_A_PAVCvIjB5_0(.dout(w_n1562_0[0]),.din(w_dff_A_PAVCvIjB5_0),.clk(gclk));
	jdff dff_A_OgBIZFUB7_0(.dout(w_dff_A_PAVCvIjB5_0),.din(w_dff_A_OgBIZFUB7_0),.clk(gclk));
	jdff dff_A_mN0ce6hD7_0(.dout(w_dff_A_OgBIZFUB7_0),.din(w_dff_A_mN0ce6hD7_0),.clk(gclk));
	jdff dff_A_jWx3Jy360_0(.dout(w_dff_A_mN0ce6hD7_0),.din(w_dff_A_jWx3Jy360_0),.clk(gclk));
	jdff dff_A_sNwyBztz9_0(.dout(w_dff_A_jWx3Jy360_0),.din(w_dff_A_sNwyBztz9_0),.clk(gclk));
	jdff dff_A_mwdLIJc12_0(.dout(w_dff_A_sNwyBztz9_0),.din(w_dff_A_mwdLIJc12_0),.clk(gclk));
	jdff dff_A_uzD2hOmg0_0(.dout(w_dff_A_mwdLIJc12_0),.din(w_dff_A_uzD2hOmg0_0),.clk(gclk));
	jdff dff_A_CNVqdke96_1(.dout(w_n1562_0[1]),.din(w_dff_A_CNVqdke96_1),.clk(gclk));
	jdff dff_A_XjAjlG513_1(.dout(w_dff_A_CNVqdke96_1),.din(w_dff_A_XjAjlG513_1),.clk(gclk));
	jdff dff_A_whqrPRhn5_1(.dout(w_dff_A_XjAjlG513_1),.din(w_dff_A_whqrPRhn5_1),.clk(gclk));
	jdff dff_A_hZU2Twyh5_1(.dout(w_dff_A_whqrPRhn5_1),.din(w_dff_A_hZU2Twyh5_1),.clk(gclk));
	jdff dff_A_4UNpTZPn2_1(.dout(w_dff_A_hZU2Twyh5_1),.din(w_dff_A_4UNpTZPn2_1),.clk(gclk));
	jdff dff_A_bqsqtYaC7_1(.dout(w_dff_A_4UNpTZPn2_1),.din(w_dff_A_bqsqtYaC7_1),.clk(gclk));
	jdff dff_A_BGKrLFec7_1(.dout(w_dff_A_bqsqtYaC7_1),.din(w_dff_A_BGKrLFec7_1),.clk(gclk));
	jdff dff_B_uLmvtIRD8_0(.din(n1559),.dout(w_dff_B_uLmvtIRD8_0),.clk(gclk));
	jdff dff_B_Rvwz1Ntt5_0(.din(w_dff_B_uLmvtIRD8_0),.dout(w_dff_B_Rvwz1Ntt5_0),.clk(gclk));
	jdff dff_B_I4GYQyWz0_0(.din(w_dff_B_Rvwz1Ntt5_0),.dout(w_dff_B_I4GYQyWz0_0),.clk(gclk));
	jdff dff_B_FFuF2WM68_0(.din(n1557),.dout(w_dff_B_FFuF2WM68_0),.clk(gclk));
	jdff dff_A_eZkA2yIW6_1(.dout(w_n1408_0[1]),.din(w_dff_A_eZkA2yIW6_1),.clk(gclk));
	jdff dff_A_IjDgqFsP6_1(.dout(w_dff_A_eZkA2yIW6_1),.din(w_dff_A_IjDgqFsP6_1),.clk(gclk));
	jdff dff_A_05DUFI563_1(.dout(w_dff_A_IjDgqFsP6_1),.din(w_dff_A_05DUFI563_1),.clk(gclk));
	jdff dff_A_WPxaR21L2_1(.dout(w_dff_A_05DUFI563_1),.din(w_dff_A_WPxaR21L2_1),.clk(gclk));
	jdff dff_A_K8H2s6xj3_1(.dout(w_dff_A_WPxaR21L2_1),.din(w_dff_A_K8H2s6xj3_1),.clk(gclk));
	jdff dff_A_MWmQHqrw8_1(.dout(w_dff_A_K8H2s6xj3_1),.din(w_dff_A_MWmQHqrw8_1),.clk(gclk));
	jdff dff_A_H227V6P77_1(.dout(w_dff_A_MWmQHqrw8_1),.din(w_dff_A_H227V6P77_1),.clk(gclk));
	jdff dff_B_qwYIpRNY4_1(.din(n1403),.dout(w_dff_B_qwYIpRNY4_1),.clk(gclk));
	jdff dff_B_oUKrvhW93_1(.din(w_dff_B_qwYIpRNY4_1),.dout(w_dff_B_oUKrvhW93_1),.clk(gclk));
	jdff dff_B_yJorNVda5_1(.din(w_dff_B_oUKrvhW93_1),.dout(w_dff_B_yJorNVda5_1),.clk(gclk));
	jdff dff_B_mp19wXpG4_1(.din(w_dff_B_yJorNVda5_1),.dout(w_dff_B_mp19wXpG4_1),.clk(gclk));
	jdff dff_B_j7ri32Ll5_1(.din(w_dff_B_mp19wXpG4_1),.dout(w_dff_B_j7ri32Ll5_1),.clk(gclk));
	jdff dff_B_rqgIY5ES8_1(.din(w_dff_B_j7ri32Ll5_1),.dout(w_dff_B_rqgIY5ES8_1),.clk(gclk));
	jdff dff_B_EKprS7Q16_0(.din(n1405),.dout(w_dff_B_EKprS7Q16_0),.clk(gclk));
	jdff dff_B_bGDSMlsM5_0(.din(w_dff_B_EKprS7Q16_0),.dout(w_dff_B_bGDSMlsM5_0),.clk(gclk));
	jdff dff_B_CnVb1Lwf1_0(.din(w_dff_B_bGDSMlsM5_0),.dout(w_dff_B_CnVb1Lwf1_0),.clk(gclk));
	jdff dff_A_TabvV23X2_1(.dout(w_n1402_0[1]),.din(w_dff_A_TabvV23X2_1),.clk(gclk));
	jdff dff_A_vswOw34m7_1(.dout(w_dff_A_TabvV23X2_1),.din(w_dff_A_vswOw34m7_1),.clk(gclk));
	jdff dff_A_M1TycP0p7_1(.dout(w_dff_A_vswOw34m7_1),.din(w_dff_A_M1TycP0p7_1),.clk(gclk));
	jdff dff_A_dfIKLkOG9_1(.dout(w_dff_A_M1TycP0p7_1),.din(w_dff_A_dfIKLkOG9_1),.clk(gclk));
	jdff dff_A_DdevqCW49_1(.dout(w_dff_A_dfIKLkOG9_1),.din(w_dff_A_DdevqCW49_1),.clk(gclk));
	jdff dff_A_MLEKQuC59_1(.dout(w_dff_A_DdevqCW49_1),.din(w_dff_A_MLEKQuC59_1),.clk(gclk));
	jdff dff_A_ngUTuCte4_1(.dout(w_dff_A_MLEKQuC59_1),.din(w_dff_A_ngUTuCte4_1),.clk(gclk));
	jdff dff_A_x3DqQd8p4_1(.dout(w_dff_A_ngUTuCte4_1),.din(w_dff_A_x3DqQd8p4_1),.clk(gclk));
	jdff dff_A_Sg5V6eJQ8_1(.dout(w_dff_A_x3DqQd8p4_1),.din(w_dff_A_Sg5V6eJQ8_1),.clk(gclk));
	jdff dff_A_o9f56Jhc7_1(.dout(w_dff_A_Sg5V6eJQ8_1),.din(w_dff_A_o9f56Jhc7_1),.clk(gclk));
	jdff dff_A_39Do16BY4_1(.dout(w_dff_A_o9f56Jhc7_1),.din(w_dff_A_39Do16BY4_1),.clk(gclk));
	jdff dff_A_ahBHxoSc6_1(.dout(w_dff_A_39Do16BY4_1),.din(w_dff_A_ahBHxoSc6_1),.clk(gclk));
	jdff dff_A_n6i6XZTi2_1(.dout(w_dff_A_ahBHxoSc6_1),.din(w_dff_A_n6i6XZTi2_1),.clk(gclk));
	jdff dff_A_oWXDgH8R3_1(.dout(w_dff_A_n6i6XZTi2_1),.din(w_dff_A_oWXDgH8R3_1),.clk(gclk));
	jdff dff_A_07VbPBFq4_1(.dout(w_dff_A_oWXDgH8R3_1),.din(w_dff_A_07VbPBFq4_1),.clk(gclk));
	jdff dff_B_1eGYARXL9_0(.din(n1549),.dout(w_dff_B_1eGYARXL9_0),.clk(gclk));
	jdff dff_B_JC4Q6jwA2_0(.din(n1548),.dout(w_dff_B_JC4Q6jwA2_0),.clk(gclk));
	jdff dff_B_wwtBx1AL7_1(.din(n1311),.dout(w_dff_B_wwtBx1AL7_1),.clk(gclk));
	jdff dff_B_Zd7shYUE7_1(.din(w_dff_B_wwtBx1AL7_1),.dout(w_dff_B_Zd7shYUE7_1),.clk(gclk));
	jdff dff_B_4RDfK5419_1(.din(w_dff_B_Zd7shYUE7_1),.dout(w_dff_B_4RDfK5419_1),.clk(gclk));
	jdff dff_B_cpxQha6Z2_1(.din(w_dff_B_4RDfK5419_1),.dout(w_dff_B_cpxQha6Z2_1),.clk(gclk));
	jdff dff_B_kyDp6uk88_1(.din(w_dff_B_cpxQha6Z2_1),.dout(w_dff_B_kyDp6uk88_1),.clk(gclk));
	jdff dff_B_oJVVuy8x8_1(.din(w_dff_B_kyDp6uk88_1),.dout(w_dff_B_oJVVuy8x8_1),.clk(gclk));
	jdff dff_B_SEwrgOtF6_1(.din(w_dff_B_oJVVuy8x8_1),.dout(w_dff_B_SEwrgOtF6_1),.clk(gclk));
	jdff dff_B_NudPdGMP0_1(.din(w_dff_B_SEwrgOtF6_1),.dout(w_dff_B_NudPdGMP0_1),.clk(gclk));
	jdff dff_B_tVNopkYn6_1(.din(w_dff_B_NudPdGMP0_1),.dout(w_dff_B_tVNopkYn6_1),.clk(gclk));
	jdff dff_B_eDtWO0qj3_1(.din(w_dff_B_tVNopkYn6_1),.dout(w_dff_B_eDtWO0qj3_1),.clk(gclk));
	jdff dff_B_hMF0gLGw1_1(.din(w_dff_B_eDtWO0qj3_1),.dout(w_dff_B_hMF0gLGw1_1),.clk(gclk));
	jdff dff_B_R7AEYJd50_1(.din(w_dff_B_hMF0gLGw1_1),.dout(w_dff_B_R7AEYJd50_1),.clk(gclk));
	jdff dff_B_eZ81QOBf4_0(.din(n1545),.dout(w_dff_B_eZ81QOBf4_0),.clk(gclk));
	jdff dff_A_3BncMQJW6_1(.dout(w_n1543_0[1]),.din(w_dff_A_3BncMQJW6_1),.clk(gclk));
	jdff dff_B_4FNzd9Pc5_2(.din(n1543),.dout(w_dff_B_4FNzd9Pc5_2),.clk(gclk));
	jdff dff_B_24mtxUlb8_2(.din(w_dff_B_4FNzd9Pc5_2),.dout(w_dff_B_24mtxUlb8_2),.clk(gclk));
	jdff dff_B_kBZpwD7o1_0(.din(n1542),.dout(w_dff_B_kBZpwD7o1_0),.clk(gclk));
	jdff dff_B_hm3K74fN6_0(.din(w_dff_B_kBZpwD7o1_0),.dout(w_dff_B_hm3K74fN6_0),.clk(gclk));
	jdff dff_B_XEqBx23A8_0(.din(w_dff_B_hm3K74fN6_0),.dout(w_dff_B_XEqBx23A8_0),.clk(gclk));
	jdff dff_B_4xMheUue8_0(.din(w_dff_B_XEqBx23A8_0),.dout(w_dff_B_4xMheUue8_0),.clk(gclk));
	jdff dff_B_FkQP94Gv6_0(.din(n1541),.dout(w_dff_B_FkQP94Gv6_0),.clk(gclk));
	jdff dff_B_CO0nfNWu6_1(.din(n1538),.dout(w_dff_B_CO0nfNWu6_1),.clk(gclk));
	jdff dff_B_QDA88Cd25_1(.din(w_dff_B_CO0nfNWu6_1),.dout(w_dff_B_QDA88Cd25_1),.clk(gclk));
	jdff dff_B_EU2ykJhL3_1(.din(w_dff_B_QDA88Cd25_1),.dout(w_dff_B_EU2ykJhL3_1),.clk(gclk));
	jdff dff_A_h2VvtMUM2_0(.dout(w_n1536_0[0]),.din(w_dff_A_h2VvtMUM2_0),.clk(gclk));
	jdff dff_A_WMngvtCD5_0(.dout(w_dff_A_h2VvtMUM2_0),.din(w_dff_A_WMngvtCD5_0),.clk(gclk));
	jdff dff_A_mRLmi6Zn1_0(.dout(w_dff_A_WMngvtCD5_0),.din(w_dff_A_mRLmi6Zn1_0),.clk(gclk));
	jdff dff_A_W85UgazU7_0(.dout(w_dff_A_mRLmi6Zn1_0),.din(w_dff_A_W85UgazU7_0),.clk(gclk));
	jdff dff_A_9CJyk6me6_1(.dout(w_n1426_0[1]),.din(w_dff_A_9CJyk6me6_1),.clk(gclk));
	jdff dff_A_JfAr3Uyd2_1(.dout(w_dff_A_9CJyk6me6_1),.din(w_dff_A_JfAr3Uyd2_1),.clk(gclk));
	jdff dff_A_aTcH09wp5_1(.dout(w_dff_A_JfAr3Uyd2_1),.din(w_dff_A_aTcH09wp5_1),.clk(gclk));
	jdff dff_A_pHS2QGSq2_1(.dout(w_dff_A_aTcH09wp5_1),.din(w_dff_A_pHS2QGSq2_1),.clk(gclk));
	jdff dff_A_ipZqOBiQ8_1(.dout(w_dff_A_pHS2QGSq2_1),.din(w_dff_A_ipZqOBiQ8_1),.clk(gclk));
	jdff dff_A_oTx87bls5_1(.dout(w_dff_A_ipZqOBiQ8_1),.din(w_dff_A_oTx87bls5_1),.clk(gclk));
	jdff dff_A_iqqYYH0K0_1(.dout(w_dff_A_oTx87bls5_1),.din(w_dff_A_iqqYYH0K0_1),.clk(gclk));
	jdff dff_A_vygkvrDe7_1(.dout(w_dff_A_iqqYYH0K0_1),.din(w_dff_A_vygkvrDe7_1),.clk(gclk));
	jdff dff_A_bRsDcaSe0_1(.dout(w_dff_A_vygkvrDe7_1),.din(w_dff_A_bRsDcaSe0_1),.clk(gclk));
	jdff dff_A_TF5cqGEb7_1(.dout(w_dff_A_bRsDcaSe0_1),.din(w_dff_A_TF5cqGEb7_1),.clk(gclk));
	jdff dff_A_8IWkgJBx5_1(.dout(w_dff_A_TF5cqGEb7_1),.din(w_dff_A_8IWkgJBx5_1),.clk(gclk));
	jdff dff_A_LoRLtfpl3_1(.dout(w_dff_A_8IWkgJBx5_1),.din(w_dff_A_LoRLtfpl3_1),.clk(gclk));
	jdff dff_A_UEjyKK6E7_1(.dout(w_dff_A_LoRLtfpl3_1),.din(w_dff_A_UEjyKK6E7_1),.clk(gclk));
	jdff dff_A_TR24fotw6_1(.dout(w_dff_A_UEjyKK6E7_1),.din(w_dff_A_TR24fotw6_1),.clk(gclk));
	jdff dff_A_tVeRf5z89_1(.dout(w_dff_A_TR24fotw6_1),.din(w_dff_A_tVeRf5z89_1),.clk(gclk));
	jdff dff_A_mdctKRx36_1(.dout(w_dff_A_tVeRf5z89_1),.din(w_dff_A_mdctKRx36_1),.clk(gclk));
	jdff dff_B_uMxn8nPI8_0(.din(n1533),.dout(w_dff_B_uMxn8nPI8_0),.clk(gclk));
	jdff dff_B_0VGiGqZB7_0(.din(w_dff_B_uMxn8nPI8_0),.dout(w_dff_B_0VGiGqZB7_0),.clk(gclk));
	jdff dff_B_M3G9IcnN5_0(.din(w_dff_B_0VGiGqZB7_0),.dout(w_dff_B_M3G9IcnN5_0),.clk(gclk));
	jdff dff_B_mrMzToCv7_0(.din(w_dff_B_M3G9IcnN5_0),.dout(w_dff_B_mrMzToCv7_0),.clk(gclk));
	jdff dff_B_bLVqyfKW6_0(.din(n1532),.dout(w_dff_B_bLVqyfKW6_0),.clk(gclk));
	jdff dff_B_d6WT5pj18_0(.din(w_dff_B_bLVqyfKW6_0),.dout(w_dff_B_d6WT5pj18_0),.clk(gclk));
	jdff dff_B_qoeLEU5k2_0(.din(w_dff_B_d6WT5pj18_0),.dout(w_dff_B_qoeLEU5k2_0),.clk(gclk));
	jdff dff_A_qdiTRg3f2_1(.dout(w_n1419_0[1]),.din(w_dff_A_qdiTRg3f2_1),.clk(gclk));
	jdff dff_A_PVUmlWos8_1(.dout(w_dff_A_qdiTRg3f2_1),.din(w_dff_A_PVUmlWos8_1),.clk(gclk));
	jdff dff_A_reUXqUeJ4_1(.dout(w_dff_A_PVUmlWos8_1),.din(w_dff_A_reUXqUeJ4_1),.clk(gclk));
	jdff dff_A_5EqcL14M4_1(.dout(w_dff_A_reUXqUeJ4_1),.din(w_dff_A_5EqcL14M4_1),.clk(gclk));
	jdff dff_A_HQovdrkH7_1(.dout(w_dff_A_5EqcL14M4_1),.din(w_dff_A_HQovdrkH7_1),.clk(gclk));
	jdff dff_A_5tmnPJWJ9_1(.dout(w_dff_A_HQovdrkH7_1),.din(w_dff_A_5tmnPJWJ9_1),.clk(gclk));
	jdff dff_A_cZzw0s9p4_1(.dout(w_dff_A_5tmnPJWJ9_1),.din(w_dff_A_cZzw0s9p4_1),.clk(gclk));
	jdff dff_A_VqPGuDRg5_1(.dout(w_dff_A_cZzw0s9p4_1),.din(w_dff_A_VqPGuDRg5_1),.clk(gclk));
	jdff dff_A_mnaXM1OV5_1(.dout(w_dff_A_VqPGuDRg5_1),.din(w_dff_A_mnaXM1OV5_1),.clk(gclk));
	jdff dff_A_XV4JvTtJ0_1(.dout(w_dff_A_mnaXM1OV5_1),.din(w_dff_A_XV4JvTtJ0_1),.clk(gclk));
	jdff dff_A_WknRXqOa9_1(.dout(w_dff_A_XV4JvTtJ0_1),.din(w_dff_A_WknRXqOa9_1),.clk(gclk));
	jdff dff_A_X0XqqPhE6_1(.dout(w_dff_A_WknRXqOa9_1),.din(w_dff_A_X0XqqPhE6_1),.clk(gclk));
	jdff dff_A_EdZdUDdb8_1(.dout(w_dff_A_X0XqqPhE6_1),.din(w_dff_A_EdZdUDdb8_1),.clk(gclk));
	jdff dff_A_NXxsCLP79_1(.dout(w_dff_A_EdZdUDdb8_1),.din(w_dff_A_NXxsCLP79_1),.clk(gclk));
	jdff dff_A_Clg8QBrH5_1(.dout(w_dff_A_NXxsCLP79_1),.din(w_dff_A_Clg8QBrH5_1),.clk(gclk));
	jdff dff_A_JRCBIb8S9_1(.dout(w_dff_A_Clg8QBrH5_1),.din(w_dff_A_JRCBIb8S9_1),.clk(gclk));
	jdff dff_A_ML0wQCZb4_1(.dout(w_dff_A_JRCBIb8S9_1),.din(w_dff_A_ML0wQCZb4_1),.clk(gclk));
	jdff dff_A_9g0Gj25A9_1(.dout(w_dff_A_ML0wQCZb4_1),.din(w_dff_A_9g0Gj25A9_1),.clk(gclk));
	jdff dff_A_WmUiygcc7_1(.dout(w_dff_A_9g0Gj25A9_1),.din(w_dff_A_WmUiygcc7_1),.clk(gclk));
	jdff dff_A_NRvr2xNV3_1(.dout(w_dff_A_WmUiygcc7_1),.din(w_dff_A_NRvr2xNV3_1),.clk(gclk));
	jdff dff_B_XkcTUA521_2(.din(n1419),.dout(w_dff_B_XkcTUA521_2),.clk(gclk));
	jdff dff_A_FmgsxsHO6_2(.dout(w_n504_0[2]),.din(w_dff_A_FmgsxsHO6_2),.clk(gclk));
	jdff dff_B_Wb2jObOc6_1(.din(n502),.dout(w_dff_B_Wb2jObOc6_1),.clk(gclk));
	jdff dff_B_K91H5ioU1_0(.din(G66),.dout(w_dff_B_K91H5ioU1_0),.clk(gclk));
	jdff dff_A_pdW84Udt4_0(.dout(w_n501_0[0]),.din(w_dff_A_pdW84Udt4_0),.clk(gclk));
	jdff dff_A_KG5akhGz9_0(.dout(w_dff_A_pdW84Udt4_0),.din(w_dff_A_KG5akhGz9_0),.clk(gclk));
	jdff dff_A_CtKtQLz32_2(.dout(w_n501_0[2]),.din(w_dff_A_CtKtQLz32_2),.clk(gclk));
	jdff dff_A_qIxN32vE1_2(.dout(w_dff_A_CtKtQLz32_2),.din(w_dff_A_qIxN32vE1_2),.clk(gclk));
	jdff dff_A_9VwgKFyQ5_1(.dout(w_G4437_0[1]),.din(w_dff_A_9VwgKFyQ5_1),.clk(gclk));
	jdff dff_A_Rph632JF4_1(.dout(w_dff_A_9VwgKFyQ5_1),.din(w_dff_A_Rph632JF4_1),.clk(gclk));
	jdff dff_A_ruSKVlVn2_1(.dout(w_dff_A_Rph632JF4_1),.din(w_dff_A_ruSKVlVn2_1),.clk(gclk));
	jdff dff_A_bdb0wrOh4_1(.dout(w_dff_A_ruSKVlVn2_1),.din(w_dff_A_bdb0wrOh4_1),.clk(gclk));
	jdff dff_A_cUYEEm9U4_1(.dout(w_n1308_0[1]),.din(w_dff_A_cUYEEm9U4_1),.clk(gclk));
	jdff dff_A_Y9db0dxp5_1(.dout(w_dff_A_cUYEEm9U4_1),.din(w_dff_A_Y9db0dxp5_1),.clk(gclk));
	jdff dff_A_cAcLb03K7_1(.dout(w_dff_A_Y9db0dxp5_1),.din(w_dff_A_cAcLb03K7_1),.clk(gclk));
	jdff dff_A_VKnKUEpK1_1(.dout(w_dff_A_cAcLb03K7_1),.din(w_dff_A_VKnKUEpK1_1),.clk(gclk));
	jdff dff_A_MH9i3ecq1_1(.dout(w_dff_A_VKnKUEpK1_1),.din(w_dff_A_MH9i3ecq1_1),.clk(gclk));
	jdff dff_A_CFcnAxKv8_1(.dout(w_dff_A_MH9i3ecq1_1),.din(w_dff_A_CFcnAxKv8_1),.clk(gclk));
	jdff dff_A_3dSPtnlF5_1(.dout(w_dff_A_CFcnAxKv8_1),.din(w_dff_A_3dSPtnlF5_1),.clk(gclk));
	jdff dff_A_PlV3Rsls8_1(.dout(w_dff_A_3dSPtnlF5_1),.din(w_dff_A_PlV3Rsls8_1),.clk(gclk));
	jdff dff_A_rWD19SEB3_1(.dout(w_dff_A_PlV3Rsls8_1),.din(w_dff_A_rWD19SEB3_1),.clk(gclk));
	jdff dff_A_0q8P4K7e5_1(.dout(w_dff_A_rWD19SEB3_1),.din(w_dff_A_0q8P4K7e5_1),.clk(gclk));
	jdff dff_A_jlJRbxIg0_1(.dout(w_dff_A_0q8P4K7e5_1),.din(w_dff_A_jlJRbxIg0_1),.clk(gclk));
	jdff dff_A_VPXYOjKq6_1(.dout(w_dff_A_jlJRbxIg0_1),.din(w_dff_A_VPXYOjKq6_1),.clk(gclk));
	jdff dff_A_sLEVuBb67_1(.dout(w_dff_A_VPXYOjKq6_1),.din(w_dff_A_sLEVuBb67_1),.clk(gclk));
	jdff dff_A_PzXjsi4a4_1(.dout(w_dff_A_sLEVuBb67_1),.din(w_dff_A_PzXjsi4a4_1),.clk(gclk));
	jdff dff_A_KfWFhUva8_1(.dout(w_dff_A_PzXjsi4a4_1),.din(w_dff_A_KfWFhUva8_1),.clk(gclk));
	jdff dff_A_sEhCQmEg5_1(.dout(w_dff_A_KfWFhUva8_1),.din(w_dff_A_sEhCQmEg5_1),.clk(gclk));
	jdff dff_A_gcnzPzKn1_0(.dout(w_n526_0[0]),.din(w_dff_A_gcnzPzKn1_0),.clk(gclk));
	jdff dff_A_gxjgvuVr0_1(.dout(w_n526_0[1]),.din(w_dff_A_gxjgvuVr0_1),.clk(gclk));
	jdff dff_A_P1G8j8sL8_1(.dout(w_dff_A_gxjgvuVr0_1),.din(w_dff_A_P1G8j8sL8_1),.clk(gclk));
	jdff dff_A_OmPDAgAM1_1(.dout(w_dff_A_P1G8j8sL8_1),.din(w_dff_A_OmPDAgAM1_1),.clk(gclk));
	jdff dff_A_woM42a805_1(.dout(w_dff_A_OmPDAgAM1_1),.din(w_dff_A_woM42a805_1),.clk(gclk));
	jdff dff_A_Mz2LidRZ3_1(.dout(w_dff_A_woM42a805_1),.din(w_dff_A_Mz2LidRZ3_1),.clk(gclk));
	jdff dff_A_QtMsrQbs7_1(.dout(w_dff_A_Mz2LidRZ3_1),.din(w_dff_A_QtMsrQbs7_1),.clk(gclk));
	jdff dff_A_qGmwrrV43_1(.dout(w_dff_A_QtMsrQbs7_1),.din(w_dff_A_qGmwrrV43_1),.clk(gclk));
	jdff dff_A_u2yqOSGB8_1(.dout(w_dff_A_qGmwrrV43_1),.din(w_dff_A_u2yqOSGB8_1),.clk(gclk));
	jdff dff_A_FuSfG6mH8_1(.dout(w_dff_A_u2yqOSGB8_1),.din(w_dff_A_FuSfG6mH8_1),.clk(gclk));
	jdff dff_A_uEB1B4xG0_1(.dout(w_dff_A_FuSfG6mH8_1),.din(w_dff_A_uEB1B4xG0_1),.clk(gclk));
	jdff dff_A_qi908Ma83_1(.dout(w_dff_A_uEB1B4xG0_1),.din(w_dff_A_qi908Ma83_1),.clk(gclk));
	jdff dff_A_A9YZY4lC3_1(.dout(w_dff_A_qi908Ma83_1),.din(w_dff_A_A9YZY4lC3_1),.clk(gclk));
	jdff dff_A_vKpHolfe5_1(.dout(w_dff_A_A9YZY4lC3_1),.din(w_dff_A_vKpHolfe5_1),.clk(gclk));
	jdff dff_A_ilokYAdb2_1(.dout(w_dff_A_vKpHolfe5_1),.din(w_dff_A_ilokYAdb2_1),.clk(gclk));
	jdff dff_A_xxYf9NAS1_1(.dout(w_dff_A_ilokYAdb2_1),.din(w_dff_A_xxYf9NAS1_1),.clk(gclk));
	jdff dff_B_X5UPQFDB0_0(.din(n1528),.dout(w_dff_B_X5UPQFDB0_0),.clk(gclk));
	jdff dff_A_NbdGURKy2_0(.dout(w_n687_0[0]),.din(w_dff_A_NbdGURKy2_0),.clk(gclk));
	jdff dff_A_Sv7nSz9l8_0(.dout(w_dff_A_NbdGURKy2_0),.din(w_dff_A_Sv7nSz9l8_0),.clk(gclk));
	jdff dff_A_FFXW9yYQ2_0(.dout(w_n694_0[0]),.din(w_dff_A_FFXW9yYQ2_0),.clk(gclk));
	jdff dff_A_tFkBshhu5_0(.dout(w_dff_A_FFXW9yYQ2_0),.din(w_dff_A_tFkBshhu5_0),.clk(gclk));
	jdff dff_A_SPOO0Qee5_0(.dout(w_dff_A_tFkBshhu5_0),.din(w_dff_A_SPOO0Qee5_0),.clk(gclk));
	jdff dff_A_dLaasbX10_0(.dout(w_dff_A_SPOO0Qee5_0),.din(w_dff_A_dLaasbX10_0),.clk(gclk));
	jdff dff_A_ACfXfwOd5_0(.dout(w_dff_A_dLaasbX10_0),.din(w_dff_A_ACfXfwOd5_0),.clk(gclk));
	jdff dff_A_OKGU5iSW0_0(.dout(w_dff_A_ACfXfwOd5_0),.din(w_dff_A_OKGU5iSW0_0),.clk(gclk));
	jdff dff_A_HWnCfUvs6_0(.dout(w_dff_A_OKGU5iSW0_0),.din(w_dff_A_HWnCfUvs6_0),.clk(gclk));
	jdff dff_A_qa8Kysc94_0(.dout(w_dff_A_HWnCfUvs6_0),.din(w_dff_A_qa8Kysc94_0),.clk(gclk));
	jdff dff_A_WSlPrr977_0(.dout(w_dff_A_qa8Kysc94_0),.din(w_dff_A_WSlPrr977_0),.clk(gclk));
	jdff dff_A_AMiEeM2x1_0(.dout(w_dff_A_WSlPrr977_0),.din(w_dff_A_AMiEeM2x1_0),.clk(gclk));
	jdff dff_A_4KU2qdNu9_0(.dout(w_dff_A_AMiEeM2x1_0),.din(w_dff_A_4KU2qdNu9_0),.clk(gclk));
	jdff dff_A_cP1V2UuK0_0(.dout(w_dff_A_4KU2qdNu9_0),.din(w_dff_A_cP1V2UuK0_0),.clk(gclk));
	jdff dff_A_EgStRu3Z1_0(.dout(w_dff_A_cP1V2UuK0_0),.din(w_dff_A_EgStRu3Z1_0),.clk(gclk));
	jdff dff_A_fZaJ32m37_0(.dout(w_dff_A_EgStRu3Z1_0),.din(w_dff_A_fZaJ32m37_0),.clk(gclk));
	jdff dff_A_DoHWcUNe7_0(.dout(w_dff_A_fZaJ32m37_0),.din(w_dff_A_DoHWcUNe7_0),.clk(gclk));
	jdff dff_A_RF0FdYnX6_0(.dout(w_dff_A_DoHWcUNe7_0),.din(w_dff_A_RF0FdYnX6_0),.clk(gclk));
	jdff dff_B_0gubTSiJ7_1(.din(n691),.dout(w_dff_B_0gubTSiJ7_1),.clk(gclk));
	jdff dff_A_X3wpJNbL7_2(.dout(w_n524_1[2]),.din(w_dff_A_X3wpJNbL7_2),.clk(gclk));
	jdff dff_A_xa0iUHlC0_2(.dout(w_dff_A_X3wpJNbL7_2),.din(w_dff_A_xa0iUHlC0_2),.clk(gclk));
	jdff dff_A_F4pBuDFz7_2(.dout(w_dff_A_xa0iUHlC0_2),.din(w_dff_A_F4pBuDFz7_2),.clk(gclk));
	jdff dff_A_3WTyAe7S4_2(.dout(w_dff_A_F4pBuDFz7_2),.din(w_dff_A_3WTyAe7S4_2),.clk(gclk));
	jdff dff_A_6C1fHsB43_2(.dout(w_dff_A_3WTyAe7S4_2),.din(w_dff_A_6C1fHsB43_2),.clk(gclk));
	jdff dff_A_ndzhgdq44_2(.dout(w_dff_A_6C1fHsB43_2),.din(w_dff_A_ndzhgdq44_2),.clk(gclk));
	jdff dff_A_8oZU5jxL3_2(.dout(w_dff_A_ndzhgdq44_2),.din(w_dff_A_8oZU5jxL3_2),.clk(gclk));
	jdff dff_A_YXHTOKGL7_2(.dout(w_dff_A_8oZU5jxL3_2),.din(w_dff_A_YXHTOKGL7_2),.clk(gclk));
	jdff dff_A_nxsvG44V5_2(.dout(w_dff_A_YXHTOKGL7_2),.din(w_dff_A_nxsvG44V5_2),.clk(gclk));
	jdff dff_A_GkxlOikL3_2(.dout(w_dff_A_nxsvG44V5_2),.din(w_dff_A_GkxlOikL3_2),.clk(gclk));
	jdff dff_A_RiUiXrFZ1_2(.dout(w_dff_A_GkxlOikL3_2),.din(w_dff_A_RiUiXrFZ1_2),.clk(gclk));
	jdff dff_A_n5DF96ap2_2(.dout(w_dff_A_RiUiXrFZ1_2),.din(w_dff_A_n5DF96ap2_2),.clk(gclk));
	jdff dff_A_egbsKCSp0_2(.dout(w_dff_A_n5DF96ap2_2),.din(w_dff_A_egbsKCSp0_2),.clk(gclk));
	jdff dff_A_bGYEB6pl8_2(.dout(w_dff_A_egbsKCSp0_2),.din(w_dff_A_bGYEB6pl8_2),.clk(gclk));
	jdff dff_A_0Z6mcsHj6_2(.dout(w_dff_A_bGYEB6pl8_2),.din(w_dff_A_0Z6mcsHj6_2),.clk(gclk));
	jdff dff_A_tnuH08Or1_2(.dout(w_dff_A_0Z6mcsHj6_2),.din(w_dff_A_tnuH08Or1_2),.clk(gclk));
	jdff dff_A_rPeFpmjZ9_2(.dout(w_dff_A_tnuH08Or1_2),.din(w_dff_A_rPeFpmjZ9_2),.clk(gclk));
	jdff dff_A_WpnNlCOD7_0(.dout(w_n518_1[0]),.din(w_dff_A_WpnNlCOD7_0),.clk(gclk));
	jdff dff_A_lIoSxRE81_0(.dout(w_dff_A_WpnNlCOD7_0),.din(w_dff_A_lIoSxRE81_0),.clk(gclk));
	jdff dff_A_V1kp8t771_0(.dout(w_dff_A_lIoSxRE81_0),.din(w_dff_A_V1kp8t771_0),.clk(gclk));
	jdff dff_A_7QRC78JY0_0(.dout(w_dff_A_V1kp8t771_0),.din(w_dff_A_7QRC78JY0_0),.clk(gclk));
	jdff dff_A_Lw0NA0X93_0(.dout(w_dff_A_7QRC78JY0_0),.din(w_dff_A_Lw0NA0X93_0),.clk(gclk));
	jdff dff_A_UZoUoleR8_0(.dout(w_dff_A_Lw0NA0X93_0),.din(w_dff_A_UZoUoleR8_0),.clk(gclk));
	jdff dff_A_E761DXP95_0(.dout(w_dff_A_UZoUoleR8_0),.din(w_dff_A_E761DXP95_0),.clk(gclk));
	jdff dff_A_QaSYnA678_0(.dout(w_dff_A_E761DXP95_0),.din(w_dff_A_QaSYnA678_0),.clk(gclk));
	jdff dff_A_eUgnv7qh7_0(.dout(w_dff_A_QaSYnA678_0),.din(w_dff_A_eUgnv7qh7_0),.clk(gclk));
	jdff dff_A_m9MJl1UE7_0(.dout(w_dff_A_eUgnv7qh7_0),.din(w_dff_A_m9MJl1UE7_0),.clk(gclk));
	jdff dff_A_5U7xi0fk0_0(.dout(w_dff_A_m9MJl1UE7_0),.din(w_dff_A_5U7xi0fk0_0),.clk(gclk));
	jdff dff_A_PzPvBfxc1_0(.dout(w_dff_A_5U7xi0fk0_0),.din(w_dff_A_PzPvBfxc1_0),.clk(gclk));
	jdff dff_A_VU7ydF1Q8_0(.dout(w_dff_A_PzPvBfxc1_0),.din(w_dff_A_VU7ydF1Q8_0),.clk(gclk));
	jdff dff_A_eUTDHlIA4_0(.dout(w_dff_A_VU7ydF1Q8_0),.din(w_dff_A_eUTDHlIA4_0),.clk(gclk));
	jdff dff_A_txV26H1W3_0(.dout(w_dff_A_eUTDHlIA4_0),.din(w_dff_A_txV26H1W3_0),.clk(gclk));
	jdff dff_A_zSSjrwjo9_0(.dout(w_dff_A_txV26H1W3_0),.din(w_dff_A_zSSjrwjo9_0),.clk(gclk));
	jdff dff_A_6BYmRLtj1_0(.dout(w_dff_A_zSSjrwjo9_0),.din(w_dff_A_6BYmRLtj1_0),.clk(gclk));
	jdff dff_A_lCny2K5N7_0(.dout(w_dff_A_6BYmRLtj1_0),.din(w_dff_A_lCny2K5N7_0),.clk(gclk));
	jdff dff_B_1BBgLLMX6_1(.din(n515),.dout(w_dff_B_1BBgLLMX6_1),.clk(gclk));
	jdff dff_B_ZDKRkgen7_0(.din(G35),.dout(w_dff_B_ZDKRkgen7_0),.clk(gclk));
	jdff dff_B_DR692JWO3_2(.din(n514),.dout(w_dff_B_DR692JWO3_2),.clk(gclk));
	jdff dff_B_o50higMX4_2(.din(w_dff_B_DR692JWO3_2),.dout(w_dff_B_o50higMX4_2),.clk(gclk));
	jdff dff_A_GhDTW6uW7_0(.dout(w_G4420_1[0]),.din(w_dff_A_GhDTW6uW7_0),.clk(gclk));
	jdff dff_A_yfxtB0Mj6_0(.dout(w_dff_A_GhDTW6uW7_0),.din(w_dff_A_yfxtB0Mj6_0),.clk(gclk));
	jdff dff_A_5gr2MZxc3_0(.dout(w_dff_A_yfxtB0Mj6_0),.din(w_dff_A_5gr2MZxc3_0),.clk(gclk));
	jdff dff_A_QOT75w8e3_0(.dout(w_dff_A_5gr2MZxc3_0),.din(w_dff_A_QOT75w8e3_0),.clk(gclk));
	jdff dff_B_hfhO92eX9_1(.din(n521),.dout(w_dff_B_hfhO92eX9_1),.clk(gclk));
	jdff dff_B_Tf4sktAQ5_0(.din(G32),.dout(w_dff_B_Tf4sktAQ5_0),.clk(gclk));
	jdff dff_B_RoOexd8W5_2(.din(n520),.dout(w_dff_B_RoOexd8W5_2),.clk(gclk));
	jdff dff_B_s3BtrIMB0_2(.din(w_dff_B_RoOexd8W5_2),.dout(w_dff_B_s3BtrIMB0_2),.clk(gclk));
	jdff dff_A_9ccwibTO2_1(.dout(w_n690_0[1]),.din(w_dff_A_9ccwibTO2_1),.clk(gclk));
	jdff dff_B_xsOrJPyQ6_2(.din(n690),.dout(w_dff_B_xsOrJPyQ6_2),.clk(gclk));
	jdff dff_A_OJnxlWYq1_2(.dout(w_n513_0[2]),.din(w_dff_A_OJnxlWYq1_2),.clk(gclk));
	jdff dff_A_qSmO3sxM0_2(.dout(w_dff_A_OJnxlWYq1_2),.din(w_dff_A_qSmO3sxM0_2),.clk(gclk));
	jdff dff_A_9LQtxqQs0_2(.dout(w_dff_A_qSmO3sxM0_2),.din(w_dff_A_9LQtxqQs0_2),.clk(gclk));
	jdff dff_A_cyokqCZy9_2(.dout(w_dff_A_9LQtxqQs0_2),.din(w_dff_A_cyokqCZy9_2),.clk(gclk));
	jdff dff_A_VgXoLfYa4_2(.dout(w_dff_A_cyokqCZy9_2),.din(w_dff_A_VgXoLfYa4_2),.clk(gclk));
	jdff dff_B_S7QK8PnQ1_1(.din(n510),.dout(w_dff_B_S7QK8PnQ1_1),.clk(gclk));
	jdff dff_B_GlAauAlX5_0(.din(G50),.dout(w_dff_B_GlAauAlX5_0),.clk(gclk));
	jdff dff_A_4t9OGUoO9_1(.dout(w_n509_0[1]),.din(w_dff_A_4t9OGUoO9_1),.clk(gclk));
	jdff dff_A_ze2TbJmO2_1(.dout(w_dff_A_4t9OGUoO9_1),.din(w_dff_A_ze2TbJmO2_1),.clk(gclk));
	jdff dff_A_McacbpMI7_2(.dout(w_n509_0[2]),.din(w_dff_A_McacbpMI7_2),.clk(gclk));
	jdff dff_A_DSMLlou83_2(.dout(w_dff_A_McacbpMI7_2),.din(w_dff_A_DSMLlou83_2),.clk(gclk));
	jdff dff_A_lhwAhZoi6_1(.dout(w_G4432_0[1]),.din(w_dff_A_lhwAhZoi6_1),.clk(gclk));
	jdff dff_A_QUdhUQBY9_1(.dout(w_dff_A_lhwAhZoi6_1),.din(w_dff_A_QUdhUQBY9_1),.clk(gclk));
	jdff dff_A_AzityleY0_1(.dout(w_dff_A_QUdhUQBY9_1),.din(w_dff_A_AzityleY0_1),.clk(gclk));
	jdff dff_A_ttAswpf56_1(.dout(w_dff_A_AzityleY0_1),.din(w_dff_A_ttAswpf56_1),.clk(gclk));
	jdff dff_A_TLQRb0oS4_1(.dout(w_n1309_0[1]),.din(w_dff_A_TLQRb0oS4_1),.clk(gclk));
	jdff dff_A_fojp8nj44_1(.dout(w_dff_A_TLQRb0oS4_1),.din(w_dff_A_fojp8nj44_1),.clk(gclk));
	jdff dff_A_TiY8jbIF4_1(.dout(w_dff_A_fojp8nj44_1),.din(w_dff_A_TiY8jbIF4_1),.clk(gclk));
	jdff dff_A_Uy6kw2GG4_1(.dout(w_dff_A_TiY8jbIF4_1),.din(w_dff_A_Uy6kw2GG4_1),.clk(gclk));
	jdff dff_A_QAA4dzyl1_1(.dout(w_n572_1[1]),.din(w_dff_A_QAA4dzyl1_1),.clk(gclk));
	jdff dff_A_icwwhiNp2_1(.dout(w_dff_A_QAA4dzyl1_1),.din(w_dff_A_icwwhiNp2_1),.clk(gclk));
	jdff dff_A_BzJeaHSw9_1(.dout(w_dff_A_icwwhiNp2_1),.din(w_dff_A_BzJeaHSw9_1),.clk(gclk));
	jdff dff_A_O2xbLzO42_1(.dout(w_dff_A_BzJeaHSw9_1),.din(w_dff_A_O2xbLzO42_1),.clk(gclk));
	jdff dff_A_qmdxOz5k3_1(.dout(w_dff_A_O2xbLzO42_1),.din(w_dff_A_qmdxOz5k3_1),.clk(gclk));
	jdff dff_B_a6OhZh6Y1_1(.din(n532),.dout(w_dff_B_a6OhZh6Y1_1),.clk(gclk));
	jdff dff_B_f82gaWqz6_1(.din(w_dff_B_a6OhZh6Y1_1),.dout(w_dff_B_f82gaWqz6_1),.clk(gclk));
	jdff dff_B_tH0iE8Zk9_1(.din(w_dff_B_f82gaWqz6_1),.dout(w_dff_B_tH0iE8Zk9_1),.clk(gclk));
	jdff dff_B_1xEumEkB4_1(.din(w_dff_B_tH0iE8Zk9_1),.dout(w_dff_B_1xEumEkB4_1),.clk(gclk));
	jdff dff_B_qjwCuMP90_1(.din(w_dff_B_1xEumEkB4_1),.dout(w_dff_B_qjwCuMP90_1),.clk(gclk));
	jdff dff_B_0H8kGMJe9_1(.din(w_dff_B_qjwCuMP90_1),.dout(w_dff_B_0H8kGMJe9_1),.clk(gclk));
	jdff dff_B_0osHwrEi3_1(.din(w_dff_B_0H8kGMJe9_1),.dout(w_dff_B_0osHwrEi3_1),.clk(gclk));
	jdff dff_B_zL3CkYRw0_1(.din(w_dff_B_0osHwrEi3_1),.dout(w_dff_B_zL3CkYRw0_1),.clk(gclk));
	jdff dff_B_w5dep8MM1_1(.din(w_dff_B_zL3CkYRw0_1),.dout(w_dff_B_w5dep8MM1_1),.clk(gclk));
	jdff dff_B_14DQgkg33_1(.din(n535),.dout(w_dff_B_14DQgkg33_1),.clk(gclk));
	jdff dff_B_iS5JGtt31_1(.din(w_dff_B_14DQgkg33_1),.dout(w_dff_B_iS5JGtt31_1),.clk(gclk));
	jdff dff_B_1LTYs2VH4_1(.din(w_dff_B_iS5JGtt31_1),.dout(w_dff_B_1LTYs2VH4_1),.clk(gclk));
	jdff dff_B_CXbr2tSP6_1(.din(w_dff_B_1LTYs2VH4_1),.dout(w_dff_B_CXbr2tSP6_1),.clk(gclk));
	jdff dff_B_6gyHgv593_1(.din(w_dff_B_CXbr2tSP6_1),.dout(w_dff_B_6gyHgv593_1),.clk(gclk));
	jdff dff_B_o9pz9yqM5_1(.din(w_dff_B_6gyHgv593_1),.dout(w_dff_B_o9pz9yqM5_1),.clk(gclk));
	jdff dff_A_7qvt01Gw7_1(.dout(w_n570_1[1]),.din(w_dff_A_7qvt01Gw7_1),.clk(gclk));
	jdff dff_A_EeAwhK9t6_1(.dout(w_dff_A_7qvt01Gw7_1),.din(w_dff_A_EeAwhK9t6_1),.clk(gclk));
	jdff dff_A_jVlUQMio7_1(.dout(w_dff_A_EeAwhK9t6_1),.din(w_dff_A_jVlUQMio7_1),.clk(gclk));
	jdff dff_A_HybwZxUB0_1(.dout(w_dff_A_jVlUQMio7_1),.din(w_dff_A_HybwZxUB0_1),.clk(gclk));
	jdff dff_A_45QPxJd27_1(.dout(w_dff_A_HybwZxUB0_1),.din(w_dff_A_45QPxJd27_1),.clk(gclk));
	jdff dff_A_9zizjlgD3_1(.dout(w_dff_A_45QPxJd27_1),.din(w_dff_A_9zizjlgD3_1),.clk(gclk));
	jdff dff_A_a2DMK6Mh4_1(.dout(w_dff_A_9zizjlgD3_1),.din(w_dff_A_a2DMK6Mh4_1),.clk(gclk));
	jdff dff_B_yiMi5WIJ2_1(.din(n540),.dout(w_dff_B_yiMi5WIJ2_1),.clk(gclk));
	jdff dff_B_RPzbXaBE0_1(.din(w_dff_B_yiMi5WIJ2_1),.dout(w_dff_B_RPzbXaBE0_1),.clk(gclk));
	jdff dff_B_oicmsVBS8_1(.din(w_dff_B_RPzbXaBE0_1),.dout(w_dff_B_oicmsVBS8_1),.clk(gclk));
	jdff dff_B_EEYomzKA0_1(.din(w_dff_B_oicmsVBS8_1),.dout(w_dff_B_EEYomzKA0_1),.clk(gclk));
	jdff dff_B_Z9Yjz69g1_1(.din(w_dff_B_EEYomzKA0_1),.dout(w_dff_B_Z9Yjz69g1_1),.clk(gclk));
	jdff dff_B_nPL5O5D18_1(.din(w_dff_B_Z9Yjz69g1_1),.dout(w_dff_B_nPL5O5D18_1),.clk(gclk));
	jdff dff_B_aKKKoBAO2_1(.din(w_dff_B_nPL5O5D18_1),.dout(w_dff_B_aKKKoBAO2_1),.clk(gclk));
	jdff dff_B_Me8b3bQA0_1(.din(n543),.dout(w_dff_B_Me8b3bQA0_1),.clk(gclk));
	jdff dff_B_zoefxJOB6_1(.din(w_dff_B_Me8b3bQA0_1),.dout(w_dff_B_zoefxJOB6_1),.clk(gclk));
	jdff dff_B_oRD1y27v5_1(.din(w_dff_B_zoefxJOB6_1),.dout(w_dff_B_oRD1y27v5_1),.clk(gclk));
	jdff dff_B_Hit352gK4_1(.din(w_dff_B_oRD1y27v5_1),.dout(w_dff_B_Hit352gK4_1),.clk(gclk));
	jdff dff_B_LBb1e79w3_1(.din(n551),.dout(w_dff_B_LBb1e79w3_1),.clk(gclk));
	jdff dff_B_Md0cH27z3_1(.din(w_dff_B_LBb1e79w3_1),.dout(w_dff_B_Md0cH27z3_1),.clk(gclk));
	jdff dff_A_j7Vpwvjf1_0(.dout(w_n566_0[0]),.din(w_dff_A_j7Vpwvjf1_0),.clk(gclk));
	jdff dff_A_nMqu4bjN2_0(.dout(w_dff_A_j7Vpwvjf1_0),.din(w_dff_A_nMqu4bjN2_0),.clk(gclk));
	jdff dff_A_cU02PYpS4_0(.dout(w_dff_A_nMqu4bjN2_0),.din(w_dff_A_cU02PYpS4_0),.clk(gclk));
	jdff dff_A_RgqDsN3a3_0(.dout(w_dff_A_cU02PYpS4_0),.din(w_dff_A_RgqDsN3a3_0),.clk(gclk));
	jdff dff_A_6Lo7wcKL3_0(.dout(w_dff_A_RgqDsN3a3_0),.din(w_dff_A_6Lo7wcKL3_0),.clk(gclk));
	jdff dff_A_2ImJFL3k4_0(.dout(w_dff_A_6Lo7wcKL3_0),.din(w_dff_A_2ImJFL3k4_0),.clk(gclk));
	jdff dff_A_BrNc2Zwt0_0(.dout(w_dff_A_2ImJFL3k4_0),.din(w_dff_A_BrNc2Zwt0_0),.clk(gclk));
	jdff dff_A_ZB5F9ZHS6_0(.dout(w_dff_A_BrNc2Zwt0_0),.din(w_dff_A_ZB5F9ZHS6_0),.clk(gclk));
	jdff dff_A_wY4cOqzB6_0(.dout(w_dff_A_ZB5F9ZHS6_0),.din(w_dff_A_wY4cOqzB6_0),.clk(gclk));
	jdff dff_A_ujQXfP9L6_0(.dout(w_dff_A_wY4cOqzB6_0),.din(w_dff_A_ujQXfP9L6_0),.clk(gclk));
	jdff dff_A_TRgHmW7P3_0(.dout(w_dff_A_ujQXfP9L6_0),.din(w_dff_A_TRgHmW7P3_0),.clk(gclk));
	jdff dff_A_h6jXJq6t3_1(.dout(w_n564_0[1]),.din(w_dff_A_h6jXJq6t3_1),.clk(gclk));
	jdff dff_A_MhbFbLx72_1(.dout(w_dff_A_h6jXJq6t3_1),.din(w_dff_A_MhbFbLx72_1),.clk(gclk));
	jdff dff_A_KdPodqNV8_1(.dout(w_dff_A_MhbFbLx72_1),.din(w_dff_A_KdPodqNV8_1),.clk(gclk));
	jdff dff_A_a4AEExw83_1(.dout(w_dff_A_KdPodqNV8_1),.din(w_dff_A_a4AEExw83_1),.clk(gclk));
	jdff dff_A_fuN38Th80_1(.dout(w_dff_A_a4AEExw83_1),.din(w_dff_A_fuN38Th80_1),.clk(gclk));
	jdff dff_A_XYunfvvK4_1(.dout(w_dff_A_fuN38Th80_1),.din(w_dff_A_XYunfvvK4_1),.clk(gclk));
	jdff dff_A_CIq3GO9s4_1(.dout(w_dff_A_XYunfvvK4_1),.din(w_dff_A_CIq3GO9s4_1),.clk(gclk));
	jdff dff_A_4NkmOesI3_1(.dout(w_dff_A_CIq3GO9s4_1),.din(w_dff_A_4NkmOesI3_1),.clk(gclk));
	jdff dff_A_gxjmdQNJ1_1(.dout(w_dff_A_4NkmOesI3_1),.din(w_dff_A_gxjmdQNJ1_1),.clk(gclk));
	jdff dff_A_BfOUIvdr8_1(.dout(w_dff_A_gxjmdQNJ1_1),.din(w_dff_A_BfOUIvdr8_1),.clk(gclk));
	jdff dff_A_nbD5zfLn8_1(.dout(w_dff_A_BfOUIvdr8_1),.din(w_dff_A_nbD5zfLn8_1),.clk(gclk));
	jdff dff_A_Nx1p4Kpj3_1(.dout(w_dff_A_nbD5zfLn8_1),.din(w_dff_A_Nx1p4Kpj3_1),.clk(gclk));
	jdff dff_A_DfWVp4ef4_1(.dout(w_dff_A_Nx1p4Kpj3_1),.din(w_dff_A_DfWVp4ef4_1),.clk(gclk));
	jdff dff_A_MGkzqXCE2_1(.dout(w_dff_A_DfWVp4ef4_1),.din(w_dff_A_MGkzqXCE2_1),.clk(gclk));
	jdff dff_A_hFM6fXmV7_1(.dout(w_dff_A_MGkzqXCE2_1),.din(w_dff_A_hFM6fXmV7_1),.clk(gclk));
	jdff dff_A_kkEaQzo72_2(.dout(w_n564_0[2]),.din(w_dff_A_kkEaQzo72_2),.clk(gclk));
	jdff dff_A_md8RtMPF9_2(.dout(w_dff_A_kkEaQzo72_2),.din(w_dff_A_md8RtMPF9_2),.clk(gclk));
	jdff dff_A_9H7CSzP19_0(.dout(w_n558_0[0]),.din(w_dff_A_9H7CSzP19_0),.clk(gclk));
	jdff dff_A_oQuHNRS80_1(.dout(w_n556_0[1]),.din(w_dff_A_oQuHNRS80_1),.clk(gclk));
	jdff dff_A_R95kl5eb2_2(.dout(w_n556_0[2]),.din(w_dff_A_R95kl5eb2_2),.clk(gclk));
	jdff dff_A_gKKIKIjz5_2(.dout(w_dff_A_R95kl5eb2_2),.din(w_dff_A_gKKIKIjz5_2),.clk(gclk));
	jdff dff_A_dGv0HnBV7_2(.dout(w_dff_A_gKKIKIjz5_2),.din(w_dff_A_dGv0HnBV7_2),.clk(gclk));
	jdff dff_A_xtbKG4df1_0(.dout(w_n550_0[0]),.din(w_dff_A_xtbKG4df1_0),.clk(gclk));
	jdff dff_A_itcAS2LG7_0(.dout(w_dff_A_xtbKG4df1_0),.din(w_dff_A_itcAS2LG7_0),.clk(gclk));
	jdff dff_A_VWIuIhjw6_0(.dout(w_dff_A_itcAS2LG7_0),.din(w_dff_A_VWIuIhjw6_0),.clk(gclk));
	jdff dff_A_u9hrOZe56_0(.dout(w_dff_A_VWIuIhjw6_0),.din(w_dff_A_u9hrOZe56_0),.clk(gclk));
	jdff dff_A_HAQrLaVw1_0(.dout(w_dff_A_u9hrOZe56_0),.din(w_dff_A_HAQrLaVw1_0),.clk(gclk));
	jdff dff_A_E4QIsxER2_1(.dout(w_n548_0[1]),.din(w_dff_A_E4QIsxER2_1),.clk(gclk));
	jdff dff_A_QisLD6h50_1(.dout(w_dff_A_E4QIsxER2_1),.din(w_dff_A_QisLD6h50_1),.clk(gclk));
	jdff dff_A_GngKVSlr5_1(.dout(w_dff_A_QisLD6h50_1),.din(w_dff_A_GngKVSlr5_1),.clk(gclk));
	jdff dff_A_yLqtJmZL3_1(.dout(w_dff_A_GngKVSlr5_1),.din(w_dff_A_yLqtJmZL3_1),.clk(gclk));
	jdff dff_A_3WoZ6Qs11_1(.dout(w_dff_A_yLqtJmZL3_1),.din(w_dff_A_3WoZ6Qs11_1),.clk(gclk));
	jdff dff_A_aMyWZKbS1_1(.dout(w_n1310_0[1]),.din(w_dff_A_aMyWZKbS1_1),.clk(gclk));
	jdff dff_A_oKs18H4K4_1(.dout(w_dff_A_aMyWZKbS1_1),.din(w_dff_A_oKs18H4K4_1),.clk(gclk));
	jdff dff_B_iS4GFBys8_2(.din(n1310),.dout(w_dff_B_iS4GFBys8_2),.clk(gclk));
	jdff dff_B_OC3cbWcf6_2(.din(w_dff_B_iS4GFBys8_2),.dout(w_dff_B_OC3cbWcf6_2),.clk(gclk));
	jdff dff_B_hsmlqB6f6_2(.din(w_dff_B_OC3cbWcf6_2),.dout(w_dff_B_hsmlqB6f6_2),.clk(gclk));
	jdff dff_B_7CLyjbwD3_2(.din(w_dff_B_hsmlqB6f6_2),.dout(w_dff_B_7CLyjbwD3_2),.clk(gclk));
	jdff dff_B_6GTJuSD64_2(.din(w_dff_B_7CLyjbwD3_2),.dout(w_dff_B_6GTJuSD64_2),.clk(gclk));
	jdff dff_B_qZe0Y4ZI8_2(.din(w_dff_B_6GTJuSD64_2),.dout(w_dff_B_qZe0Y4ZI8_2),.clk(gclk));
	jdff dff_B_yU4cyUmK7_2(.din(w_dff_B_qZe0Y4ZI8_2),.dout(w_dff_B_yU4cyUmK7_2),.clk(gclk));
	jdff dff_B_jm3SBMPv0_2(.din(w_dff_B_yU4cyUmK7_2),.dout(w_dff_B_jm3SBMPv0_2),.clk(gclk));
	jdff dff_A_V9Yu8TzO9_0(.dout(w_n581_0[0]),.din(w_dff_A_V9Yu8TzO9_0),.clk(gclk));
	jdff dff_A_QQEgXUCX7_0(.dout(w_dff_A_V9Yu8TzO9_0),.din(w_dff_A_QQEgXUCX7_0),.clk(gclk));
	jdff dff_A_Ydu3eo0F2_0(.dout(w_dff_A_QQEgXUCX7_0),.din(w_dff_A_Ydu3eo0F2_0),.clk(gclk));
	jdff dff_A_nVS25w047_0(.dout(w_dff_A_Ydu3eo0F2_0),.din(w_dff_A_nVS25w047_0),.clk(gclk));
	jdff dff_A_XWCBOf1L4_0(.dout(w_dff_A_nVS25w047_0),.din(w_dff_A_XWCBOf1L4_0),.clk(gclk));
	jdff dff_A_13P1wu2X7_0(.dout(w_dff_A_XWCBOf1L4_0),.din(w_dff_A_13P1wu2X7_0),.clk(gclk));
	jdff dff_A_ljIFcQ6O6_0(.dout(w_dff_A_13P1wu2X7_0),.din(w_dff_A_ljIFcQ6O6_0),.clk(gclk));
	jdff dff_A_fcEi5dX74_2(.dout(w_n581_0[2]),.din(w_dff_A_fcEi5dX74_2),.clk(gclk));
	jdff dff_A_pFRmMylo5_2(.dout(w_dff_A_fcEi5dX74_2),.din(w_dff_A_pFRmMylo5_2),.clk(gclk));
	jdff dff_A_Y0RvLGZH2_2(.dout(w_dff_A_pFRmMylo5_2),.din(w_dff_A_Y0RvLGZH2_2),.clk(gclk));
	jdff dff_A_addw5Elf2_2(.dout(w_dff_A_Y0RvLGZH2_2),.din(w_dff_A_addw5Elf2_2),.clk(gclk));
	jdff dff_A_aOM5wPos3_2(.dout(w_dff_A_addw5Elf2_2),.din(w_dff_A_aOM5wPos3_2),.clk(gclk));
	jdff dff_A_a0xwW19R2_2(.dout(w_dff_A_aOM5wPos3_2),.din(w_dff_A_a0xwW19R2_2),.clk(gclk));
	jdff dff_A_m7BPBVeD9_2(.dout(w_dff_A_a0xwW19R2_2),.din(w_dff_A_m7BPBVeD9_2),.clk(gclk));
	jdff dff_A_pglbKG1h6_2(.dout(w_dff_A_m7BPBVeD9_2),.din(w_dff_A_pglbKG1h6_2),.clk(gclk));
	jdff dff_A_PQfki17f3_2(.dout(w_dff_A_pglbKG1h6_2),.din(w_dff_A_PQfki17f3_2),.clk(gclk));
	jdff dff_A_BbqT1xbR5_2(.dout(w_dff_A_PQfki17f3_2),.din(w_dff_A_BbqT1xbR5_2),.clk(gclk));
	jdff dff_A_2EevMicO9_2(.dout(w_dff_A_BbqT1xbR5_2),.din(w_dff_A_2EevMicO9_2),.clk(gclk));
	jdff dff_A_j45oVpwh7_0(.dout(w_n580_0[0]),.din(w_dff_A_j45oVpwh7_0),.clk(gclk));
	jdff dff_A_jiux9eNi8_0(.dout(w_dff_A_j45oVpwh7_0),.din(w_dff_A_jiux9eNi8_0),.clk(gclk));
	jdff dff_A_bplawuSj0_0(.dout(w_dff_A_jiux9eNi8_0),.din(w_dff_A_bplawuSj0_0),.clk(gclk));
	jdff dff_A_y4JmTDcA8_0(.dout(w_dff_A_bplawuSj0_0),.din(w_dff_A_y4JmTDcA8_0),.clk(gclk));
	jdff dff_A_WfVSZ6Rn1_0(.dout(w_dff_A_y4JmTDcA8_0),.din(w_dff_A_WfVSZ6Rn1_0),.clk(gclk));
	jdff dff_A_amHkDlX56_0(.dout(w_dff_A_WfVSZ6Rn1_0),.din(w_dff_A_amHkDlX56_0),.clk(gclk));
	jdff dff_A_IYP4Qtpr2_0(.dout(w_dff_A_amHkDlX56_0),.din(w_dff_A_IYP4Qtpr2_0),.clk(gclk));
	jdff dff_A_f47I2eI74_1(.dout(w_n580_0[1]),.din(w_dff_A_f47I2eI74_1),.clk(gclk));
	jdff dff_A_9iXGh8Hf9_1(.dout(w_dff_A_f47I2eI74_1),.din(w_dff_A_9iXGh8Hf9_1),.clk(gclk));
	jdff dff_A_rXPU0POp2_1(.dout(w_dff_A_9iXGh8Hf9_1),.din(w_dff_A_rXPU0POp2_1),.clk(gclk));
	jdff dff_A_YSOuSMyB4_1(.dout(w_dff_A_rXPU0POp2_1),.din(w_dff_A_YSOuSMyB4_1),.clk(gclk));
	jdff dff_A_HwNhSJvh4_1(.dout(w_dff_A_YSOuSMyB4_1),.din(w_dff_A_HwNhSJvh4_1),.clk(gclk));
	jdff dff_A_eYogqwxd6_1(.dout(w_dff_A_HwNhSJvh4_1),.din(w_dff_A_eYogqwxd6_1),.clk(gclk));
	jdff dff_A_VANahx7h4_1(.dout(w_dff_A_eYogqwxd6_1),.din(w_dff_A_VANahx7h4_1),.clk(gclk));
	jdff dff_A_q7M6kJU42_1(.dout(w_dff_A_VANahx7h4_1),.din(w_dff_A_q7M6kJU42_1),.clk(gclk));
	jdff dff_A_q4eSgDJJ1_1(.dout(w_dff_A_q7M6kJU42_1),.din(w_dff_A_q4eSgDJJ1_1),.clk(gclk));
	jdff dff_A_vULS35Ya7_1(.dout(w_dff_A_q4eSgDJJ1_1),.din(w_dff_A_vULS35Ya7_1),.clk(gclk));
	jdff dff_A_vjUkS9AR4_1(.dout(w_dff_A_vULS35Ya7_1),.din(w_dff_A_vjUkS9AR4_1),.clk(gclk));
	jdff dff_A_nSimRdzg0_1(.dout(w_dff_A_vjUkS9AR4_1),.din(w_dff_A_nSimRdzg0_1),.clk(gclk));
	jdff dff_A_m1xlhcAx1_0(.dout(w_n578_0[0]),.din(w_dff_A_m1xlhcAx1_0),.clk(gclk));
	jdff dff_A_eWSBL3Rl6_1(.dout(w_n578_0[1]),.din(w_dff_A_eWSBL3Rl6_1),.clk(gclk));
	jdff dff_A_tDpN4mup8_1(.dout(w_dff_A_eWSBL3Rl6_1),.din(w_dff_A_tDpN4mup8_1),.clk(gclk));
	jdff dff_A_IvD4zRpv4_1(.dout(w_dff_A_tDpN4mup8_1),.din(w_dff_A_IvD4zRpv4_1),.clk(gclk));
	jdff dff_A_STxpAMYJ6_1(.dout(w_dff_A_IvD4zRpv4_1),.din(w_dff_A_STxpAMYJ6_1),.clk(gclk));
	jdff dff_A_Zz1qrTBt0_1(.dout(w_dff_A_STxpAMYJ6_1),.din(w_dff_A_Zz1qrTBt0_1),.clk(gclk));
	jdff dff_A_UPRVCcTd1_1(.dout(w_dff_A_Zz1qrTBt0_1),.din(w_dff_A_UPRVCcTd1_1),.clk(gclk));
	jdff dff_A_GWv2Ifkk4_1(.dout(w_dff_A_UPRVCcTd1_1),.din(w_dff_A_GWv2Ifkk4_1),.clk(gclk));
	jdff dff_A_3n4UuHX64_1(.dout(w_dff_A_GWv2Ifkk4_1),.din(w_dff_A_3n4UuHX64_1),.clk(gclk));
	jdff dff_A_eXxIkS7S1_1(.dout(w_dff_A_3n4UuHX64_1),.din(w_dff_A_eXxIkS7S1_1),.clk(gclk));
	jdff dff_A_rVEXEA3D4_1(.dout(w_dff_A_eXxIkS7S1_1),.din(w_dff_A_rVEXEA3D4_1),.clk(gclk));
	jdff dff_A_f10blSsZ4_1(.dout(w_dff_A_rVEXEA3D4_1),.din(w_dff_A_f10blSsZ4_1),.clk(gclk));
	jdff dff_A_mqsdTUsB8_1(.dout(w_dff_A_f10blSsZ4_1),.din(w_dff_A_mqsdTUsB8_1),.clk(gclk));
	jdff dff_A_yJoL8IxM9_1(.dout(w_dff_A_mqsdTUsB8_1),.din(w_dff_A_yJoL8IxM9_1),.clk(gclk));
	jdff dff_A_pnN4e0tt2_1(.dout(w_dff_A_yJoL8IxM9_1),.din(w_dff_A_pnN4e0tt2_1),.clk(gclk));
	jdff dff_A_icuiq9cj9_1(.dout(w_dff_A_pnN4e0tt2_1),.din(w_dff_A_icuiq9cj9_1),.clk(gclk));
	jdff dff_A_Jy21ZVUD4_1(.dout(w_dff_A_icuiq9cj9_1),.din(w_dff_A_Jy21ZVUD4_1),.clk(gclk));
	jdff dff_B_lncsuzpc2_1(.din(n545),.dout(w_dff_B_lncsuzpc2_1),.clk(gclk));
	jdff dff_B_NdacBAVQ8_0(.din(G94),.dout(w_dff_B_NdacBAVQ8_0),.clk(gclk));
	jdff dff_B_MCOGhzGZ9_2(.din(n544),.dout(w_dff_B_MCOGhzGZ9_2),.clk(gclk));
	jdff dff_B_JLLYtHSi6_2(.din(w_dff_B_MCOGhzGZ9_2),.dout(w_dff_B_JLLYtHSi6_2),.clk(gclk));
	jdff dff_A_jsUAqiQy4_0(.dout(w_G4405_1[0]),.din(w_dff_A_jsUAqiQy4_0),.clk(gclk));
	jdff dff_A_Nwk7wgF06_0(.dout(w_dff_A_jsUAqiQy4_0),.din(w_dff_A_Nwk7wgF06_0),.clk(gclk));
	jdff dff_A_5POAQ0Lp3_0(.dout(w_dff_A_Nwk7wgF06_0),.din(w_dff_A_5POAQ0Lp3_0),.clk(gclk));
	jdff dff_A_KsBxcwTl2_0(.dout(w_dff_A_5POAQ0Lp3_0),.din(w_dff_A_KsBxcwTl2_0),.clk(gclk));
	jdff dff_B_eBTD6XLU8_1(.din(n537),.dout(w_dff_B_eBTD6XLU8_1),.clk(gclk));
	jdff dff_B_VTqLAKE61_0(.din(G121),.dout(w_dff_B_VTqLAKE61_0),.clk(gclk));
	jdff dff_A_fD6XjZkR4_1(.dout(w_n536_0[1]),.din(w_dff_A_fD6XjZkR4_1),.clk(gclk));
	jdff dff_A_hOgeOUPF7_1(.dout(w_dff_A_fD6XjZkR4_1),.din(w_dff_A_hOgeOUPF7_1),.clk(gclk));
	jdff dff_A_wLnxcjBH0_2(.dout(w_n536_0[2]),.din(w_dff_A_wLnxcjBH0_2),.clk(gclk));
	jdff dff_A_iC5C8OjB4_2(.dout(w_dff_A_wLnxcjBH0_2),.din(w_dff_A_iC5C8OjB4_2),.clk(gclk));
	jdff dff_A_DeYJNhYT6_1(.dout(w_G4410_0[1]),.din(w_dff_A_DeYJNhYT6_1),.clk(gclk));
	jdff dff_A_YXAAON592_1(.dout(w_dff_A_DeYJNhYT6_1),.din(w_dff_A_YXAAON592_1),.clk(gclk));
	jdff dff_A_yT4V3izG7_1(.dout(w_dff_A_YXAAON592_1),.din(w_dff_A_yT4V3izG7_1),.clk(gclk));
	jdff dff_A_RQNKq2ED1_1(.dout(w_dff_A_yT4V3izG7_1),.din(w_dff_A_RQNKq2ED1_1),.clk(gclk));
	jdff dff_A_H1TkR1ev1_0(.dout(w_n576_0[0]),.din(w_dff_A_H1TkR1ev1_0),.clk(gclk));
	jdff dff_A_w25X416A8_0(.dout(w_dff_A_H1TkR1ev1_0),.din(w_dff_A_w25X416A8_0),.clk(gclk));
	jdff dff_A_lUCU7CAt0_0(.dout(w_dff_A_w25X416A8_0),.din(w_dff_A_lUCU7CAt0_0),.clk(gclk));
	jdff dff_A_VOURb8ns2_0(.dout(w_dff_A_lUCU7CAt0_0),.din(w_dff_A_VOURb8ns2_0),.clk(gclk));
	jdff dff_A_Q1cYFrFu1_0(.dout(w_dff_A_VOURb8ns2_0),.din(w_dff_A_Q1cYFrFu1_0),.clk(gclk));
	jdff dff_A_xwFz6suw3_0(.dout(w_dff_A_Q1cYFrFu1_0),.din(w_dff_A_xwFz6suw3_0),.clk(gclk));
	jdff dff_A_e9mg32bY4_0(.dout(w_dff_A_xwFz6suw3_0),.din(w_dff_A_e9mg32bY4_0),.clk(gclk));
	jdff dff_A_kGhswp7n5_0(.dout(w_dff_A_e9mg32bY4_0),.din(w_dff_A_kGhswp7n5_0),.clk(gclk));
	jdff dff_A_XH39Dzng4_0(.dout(w_dff_A_kGhswp7n5_0),.din(w_dff_A_XH39Dzng4_0),.clk(gclk));
	jdff dff_A_UhNbnvkD5_0(.dout(w_dff_A_XH39Dzng4_0),.din(w_dff_A_UhNbnvkD5_0),.clk(gclk));
	jdff dff_A_F7SLceJQ5_0(.dout(w_dff_A_UhNbnvkD5_0),.din(w_dff_A_F7SLceJQ5_0),.clk(gclk));
	jdff dff_A_fviSfmSJ5_0(.dout(w_dff_A_F7SLceJQ5_0),.din(w_dff_A_fviSfmSJ5_0),.clk(gclk));
	jdff dff_A_LqCO2wEt1_0(.dout(w_dff_A_fviSfmSJ5_0),.din(w_dff_A_LqCO2wEt1_0),.clk(gclk));
	jdff dff_A_L8Jt8ksO4_0(.dout(w_n575_1[0]),.din(w_dff_A_L8Jt8ksO4_0),.clk(gclk));
	jdff dff_A_4y45Qwkg8_0(.dout(w_dff_A_L8Jt8ksO4_0),.din(w_dff_A_4y45Qwkg8_0),.clk(gclk));
	jdff dff_A_yAcqsvcv1_0(.dout(w_dff_A_4y45Qwkg8_0),.din(w_dff_A_yAcqsvcv1_0),.clk(gclk));
	jdff dff_A_hnsfD6Wa9_0(.dout(w_dff_A_yAcqsvcv1_0),.din(w_dff_A_hnsfD6Wa9_0),.clk(gclk));
	jdff dff_A_Ec1vrAUN4_0(.dout(w_dff_A_hnsfD6Wa9_0),.din(w_dff_A_Ec1vrAUN4_0),.clk(gclk));
	jdff dff_A_Q4gWlfxQ5_0(.dout(w_dff_A_Ec1vrAUN4_0),.din(w_dff_A_Q4gWlfxQ5_0),.clk(gclk));
	jdff dff_A_tc4wjIme4_0(.dout(w_dff_A_Q4gWlfxQ5_0),.din(w_dff_A_tc4wjIme4_0),.clk(gclk));
	jdff dff_A_WKkDVb398_0(.dout(w_dff_A_tc4wjIme4_0),.din(w_dff_A_WKkDVb398_0),.clk(gclk));
	jdff dff_A_zWBuL2iM5_0(.dout(w_dff_A_WKkDVb398_0),.din(w_dff_A_zWBuL2iM5_0),.clk(gclk));
	jdff dff_A_7nbNurT41_0(.dout(w_dff_A_zWBuL2iM5_0),.din(w_dff_A_7nbNurT41_0),.clk(gclk));
	jdff dff_A_1UPCQan38_0(.dout(w_dff_A_7nbNurT41_0),.din(w_dff_A_1UPCQan38_0),.clk(gclk));
	jdff dff_A_Db3vSDXQ2_0(.dout(w_dff_A_1UPCQan38_0),.din(w_dff_A_Db3vSDXQ2_0),.clk(gclk));
	jdff dff_A_fgRorDQ94_0(.dout(w_dff_A_Db3vSDXQ2_0),.din(w_dff_A_fgRorDQ94_0),.clk(gclk));
	jdff dff_A_834GmKxn6_0(.dout(w_dff_A_fgRorDQ94_0),.din(w_dff_A_834GmKxn6_0),.clk(gclk));
	jdff dff_A_mr411PyE1_2(.dout(w_n575_0[2]),.din(w_dff_A_mr411PyE1_2),.clk(gclk));
	jdff dff_A_diwNUycN8_2(.dout(w_dff_A_mr411PyE1_2),.din(w_dff_A_diwNUycN8_2),.clk(gclk));
	jdff dff_A_z8Of0bIP4_2(.dout(w_dff_A_diwNUycN8_2),.din(w_dff_A_z8Of0bIP4_2),.clk(gclk));
	jdff dff_A_cL81nsjY6_2(.dout(w_dff_A_z8Of0bIP4_2),.din(w_dff_A_cL81nsjY6_2),.clk(gclk));
	jdff dff_A_i3EjHGms9_2(.dout(w_dff_A_cL81nsjY6_2),.din(w_dff_A_i3EjHGms9_2),.clk(gclk));
	jdff dff_A_65K3OV268_2(.dout(w_dff_A_i3EjHGms9_2),.din(w_dff_A_65K3OV268_2),.clk(gclk));
	jdff dff_A_eq2zt1Y13_2(.dout(w_dff_A_65K3OV268_2),.din(w_dff_A_eq2zt1Y13_2),.clk(gclk));
	jdff dff_A_OtOJedEa0_2(.dout(w_dff_A_eq2zt1Y13_2),.din(w_dff_A_OtOJedEa0_2),.clk(gclk));
	jdff dff_A_TBsNULbG4_2(.dout(w_dff_A_OtOJedEa0_2),.din(w_dff_A_TBsNULbG4_2),.clk(gclk));
	jdff dff_A_7AA5fqZw8_2(.dout(w_dff_A_TBsNULbG4_2),.din(w_dff_A_7AA5fqZw8_2),.clk(gclk));
	jdff dff_A_AzHJQS0M2_2(.dout(w_dff_A_7AA5fqZw8_2),.din(w_dff_A_AzHJQS0M2_2),.clk(gclk));
	jdff dff_A_eg8aB7iI1_2(.dout(w_dff_A_AzHJQS0M2_2),.din(w_dff_A_eg8aB7iI1_2),.clk(gclk));
	jdff dff_A_rGfyodch6_2(.dout(w_dff_A_eg8aB7iI1_2),.din(w_dff_A_rGfyodch6_2),.clk(gclk));
	jdff dff_A_vgM6wKl89_2(.dout(w_dff_A_rGfyodch6_2),.din(w_dff_A_vgM6wKl89_2),.clk(gclk));
	jdff dff_B_zfeiiKV59_1(.din(n561),.dout(w_dff_B_zfeiiKV59_1),.clk(gclk));
	jdff dff_B_B9vMYkRe1_0(.din(G118),.dout(w_dff_B_B9vMYkRe1_0),.clk(gclk));
	jdff dff_B_qmQ8RXc35_2(.din(n560),.dout(w_dff_B_qmQ8RXc35_2),.clk(gclk));
	jdff dff_B_mbNgPm2M9_2(.din(w_dff_B_qmQ8RXc35_2),.dout(w_dff_B_mbNgPm2M9_2),.clk(gclk));
	jdff dff_A_fBS8ixlD8_2(.dout(w_G4394_0[2]),.din(w_dff_A_fBS8ixlD8_2),.clk(gclk));
	jdff dff_A_UaorlTs97_2(.dout(w_dff_A_fBS8ixlD8_2),.din(w_dff_A_UaorlTs97_2),.clk(gclk));
	jdff dff_A_WWwU03BM3_2(.dout(w_dff_A_UaorlTs97_2),.din(w_dff_A_WWwU03BM3_2),.clk(gclk));
	jdff dff_A_E5eUml0l6_2(.dout(w_dff_A_WWwU03BM3_2),.din(w_dff_A_E5eUml0l6_2),.clk(gclk));
	jdff dff_A_YjrnoYQ10_1(.dout(w_n574_0[1]),.din(w_dff_A_YjrnoYQ10_1),.clk(gclk));
	jdff dff_A_6V5Tyu9B5_1(.dout(w_dff_A_YjrnoYQ10_1),.din(w_dff_A_6V5Tyu9B5_1),.clk(gclk));
	jdff dff_A_IrR3M08e7_1(.dout(w_dff_A_6V5Tyu9B5_1),.din(w_dff_A_IrR3M08e7_1),.clk(gclk));
	jdff dff_A_CjzTuaok6_1(.dout(w_dff_A_IrR3M08e7_1),.din(w_dff_A_CjzTuaok6_1),.clk(gclk));
	jdff dff_A_Ai8doFeD4_1(.dout(w_dff_A_CjzTuaok6_1),.din(w_dff_A_Ai8doFeD4_1),.clk(gclk));
	jdff dff_A_B4W2SeIN8_1(.dout(w_dff_A_Ai8doFeD4_1),.din(w_dff_A_B4W2SeIN8_1),.clk(gclk));
	jdff dff_A_h7He2goE9_1(.dout(w_dff_A_B4W2SeIN8_1),.din(w_dff_A_h7He2goE9_1),.clk(gclk));
	jdff dff_A_C3wFZKjy1_1(.dout(w_dff_A_h7He2goE9_1),.din(w_dff_A_C3wFZKjy1_1),.clk(gclk));
	jdff dff_A_aoA6KkSh8_1(.dout(w_dff_A_C3wFZKjy1_1),.din(w_dff_A_aoA6KkSh8_1),.clk(gclk));
	jdff dff_A_lwRixicT2_1(.dout(w_dff_A_aoA6KkSh8_1),.din(w_dff_A_lwRixicT2_1),.clk(gclk));
	jdff dff_A_JcXsaGgX0_1(.dout(w_dff_A_lwRixicT2_1),.din(w_dff_A_JcXsaGgX0_1),.clk(gclk));
	jdff dff_A_kkzKgLQU8_1(.dout(w_dff_A_JcXsaGgX0_1),.din(w_dff_A_kkzKgLQU8_1),.clk(gclk));
	jdff dff_A_ytGAotxk2_1(.dout(w_dff_A_kkzKgLQU8_1),.din(w_dff_A_ytGAotxk2_1),.clk(gclk));
	jdff dff_A_UbRdQzBQ3_1(.dout(w_dff_A_ytGAotxk2_1),.din(w_dff_A_UbRdQzBQ3_1),.clk(gclk));
	jdff dff_A_FI0vtvFW6_1(.dout(w_dff_A_UbRdQzBQ3_1),.din(w_dff_A_FI0vtvFW6_1),.clk(gclk));
	jdff dff_A_XafuP8tA7_1(.dout(w_dff_A_FI0vtvFW6_1),.din(w_dff_A_XafuP8tA7_1),.clk(gclk));
	jdff dff_B_Ay4BhMt72_1(.din(n553),.dout(w_dff_B_Ay4BhMt72_1),.clk(gclk));
	jdff dff_B_d32fgfP58_0(.din(G97),.dout(w_dff_B_d32fgfP58_0),.clk(gclk));
	jdff dff_B_XMHt8AVL9_2(.din(n552),.dout(w_dff_B_XMHt8AVL9_2),.clk(gclk));
	jdff dff_B_o3YYZP3c6_2(.din(w_dff_B_XMHt8AVL9_2),.dout(w_dff_B_o3YYZP3c6_2),.clk(gclk));
	jdff dff_A_psUMw5Bv8_0(.dout(w_G4400_1[0]),.din(w_dff_A_psUMw5Bv8_0),.clk(gclk));
	jdff dff_A_ew2MzLwk9_0(.dout(w_dff_A_psUMw5Bv8_0),.din(w_dff_A_ew2MzLwk9_0),.clk(gclk));
	jdff dff_A_8ek1yGCB3_0(.dout(w_dff_A_ew2MzLwk9_0),.din(w_dff_A_8ek1yGCB3_0),.clk(gclk));
	jdff dff_A_pTOs2fBc6_0(.dout(w_dff_A_8ek1yGCB3_0),.din(w_dff_A_pTOs2fBc6_0),.clk(gclk));
	jdff dff_A_6MdOfsxL0_0(.dout(w_n573_1[0]),.din(w_dff_A_6MdOfsxL0_0),.clk(gclk));
	jdff dff_A_AIIYD2so7_0(.dout(w_dff_A_6MdOfsxL0_0),.din(w_dff_A_AIIYD2so7_0),.clk(gclk));
	jdff dff_A_REoYckIc9_0(.dout(w_dff_A_AIIYD2so7_0),.din(w_dff_A_REoYckIc9_0),.clk(gclk));
	jdff dff_A_KUOvir0x7_0(.dout(w_dff_A_REoYckIc9_0),.din(w_dff_A_KUOvir0x7_0),.clk(gclk));
	jdff dff_A_d40E8XcC7_0(.dout(w_dff_A_KUOvir0x7_0),.din(w_dff_A_d40E8XcC7_0),.clk(gclk));
	jdff dff_A_ynijqlNQ3_0(.dout(w_dff_A_d40E8XcC7_0),.din(w_dff_A_ynijqlNQ3_0),.clk(gclk));
	jdff dff_A_Kpdj06vu8_0(.dout(w_dff_A_ynijqlNQ3_0),.din(w_dff_A_Kpdj06vu8_0),.clk(gclk));
	jdff dff_A_7xQjhrrT7_0(.dout(w_dff_A_Kpdj06vu8_0),.din(w_dff_A_7xQjhrrT7_0),.clk(gclk));
	jdff dff_A_INjiewfE2_0(.dout(w_dff_A_7xQjhrrT7_0),.din(w_dff_A_INjiewfE2_0),.clk(gclk));
	jdff dff_A_ejd5kZHd0_0(.dout(w_dff_A_INjiewfE2_0),.din(w_dff_A_ejd5kZHd0_0),.clk(gclk));
	jdff dff_A_6p5yPW499_0(.dout(w_dff_A_ejd5kZHd0_0),.din(w_dff_A_6p5yPW499_0),.clk(gclk));
	jdff dff_A_4AXJbFjP3_0(.dout(w_dff_A_6p5yPW499_0),.din(w_dff_A_4AXJbFjP3_0),.clk(gclk));
	jdff dff_A_gvkPwK1R6_0(.dout(w_dff_A_4AXJbFjP3_0),.din(w_dff_A_gvkPwK1R6_0),.clk(gclk));
	jdff dff_A_hguD7QRp5_0(.dout(w_dff_A_gvkPwK1R6_0),.din(w_dff_A_hguD7QRp5_0),.clk(gclk));
	jdff dff_A_tYjulFFW0_1(.dout(w_n573_0[1]),.din(w_dff_A_tYjulFFW0_1),.clk(gclk));
	jdff dff_A_txsL6BBs8_1(.dout(w_dff_A_tYjulFFW0_1),.din(w_dff_A_txsL6BBs8_1),.clk(gclk));
	jdff dff_A_zkIvd3R72_1(.dout(w_dff_A_txsL6BBs8_1),.din(w_dff_A_zkIvd3R72_1),.clk(gclk));
	jdff dff_A_iDFAnv7Y7_2(.dout(w_n573_0[2]),.din(w_dff_A_iDFAnv7Y7_2),.clk(gclk));
	jdff dff_A_Pvhb6ZV98_2(.dout(w_dff_A_iDFAnv7Y7_2),.din(w_dff_A_Pvhb6ZV98_2),.clk(gclk));
	jdff dff_B_S8Z1ZWjF1_3(.din(n573),.dout(w_dff_B_S8Z1ZWjF1_3),.clk(gclk));
	jdff dff_B_w0b9mGea6_3(.din(w_dff_B_S8Z1ZWjF1_3),.dout(w_dff_B_w0b9mGea6_3),.clk(gclk));
	jdff dff_B_hpaCQnrD8_1(.din(n529),.dout(w_dff_B_hpaCQnrD8_1),.clk(gclk));
	jdff dff_B_zO4tm7vU4_0(.din(G47),.dout(w_dff_B_zO4tm7vU4_0),.clk(gclk));
	jdff dff_B_TXLOIQC71_2(.din(n528),.dout(w_dff_B_TXLOIQC71_2),.clk(gclk));
	jdff dff_B_6kXN9UvO1_2(.din(w_dff_B_TXLOIQC71_2),.dout(w_dff_B_6kXN9UvO1_2),.clk(gclk));
	jdff dff_A_a3ffRSgg9_0(.dout(w_G4415_1[0]),.din(w_dff_A_a3ffRSgg9_0),.clk(gclk));
	jdff dff_A_nM7jgZub7_0(.dout(w_dff_A_a3ffRSgg9_0),.din(w_dff_A_nM7jgZub7_0),.clk(gclk));
	jdff dff_A_I120n9PQ1_0(.dout(w_dff_A_nM7jgZub7_0),.din(w_dff_A_I120n9PQ1_0),.clk(gclk));
	jdff dff_A_9AKXfkfi4_0(.dout(w_dff_A_I120n9PQ1_0),.din(w_dff_A_9AKXfkfi4_0),.clk(gclk));
	jdff dff_B_aV689boM3_1(.din(n589),.dout(w_dff_B_aV689boM3_1),.clk(gclk));
	jdff dff_B_EMrRo1jj1_1(.din(w_dff_B_aV689boM3_1),.dout(w_dff_B_EMrRo1jj1_1),.clk(gclk));
	jdff dff_B_LFNDJRb97_1(.din(w_dff_B_EMrRo1jj1_1),.dout(w_dff_B_LFNDJRb97_1),.clk(gclk));
	jdff dff_B_PaXEQWEA3_1(.din(w_dff_B_LFNDJRb97_1),.dout(w_dff_B_PaXEQWEA3_1),.clk(gclk));
	jdff dff_B_yKZFxwnm6_1(.din(w_dff_B_PaXEQWEA3_1),.dout(w_dff_B_yKZFxwnm6_1),.clk(gclk));
	jdff dff_B_8AhLXQQP6_1(.din(w_dff_B_yKZFxwnm6_1),.dout(w_dff_B_8AhLXQQP6_1),.clk(gclk));
	jdff dff_B_MdLgWlRM9_1(.din(w_dff_B_8AhLXQQP6_1),.dout(w_dff_B_MdLgWlRM9_1),.clk(gclk));
	jdff dff_B_xiawR7N49_1(.din(w_dff_B_MdLgWlRM9_1),.dout(w_dff_B_xiawR7N49_1),.clk(gclk));
	jdff dff_B_T6NLPMsr0_1(.din(w_dff_B_xiawR7N49_1),.dout(w_dff_B_T6NLPMsr0_1),.clk(gclk));
	jdff dff_B_VXnoGf3b7_1(.din(w_dff_B_T6NLPMsr0_1),.dout(w_dff_B_VXnoGf3b7_1),.clk(gclk));
	jdff dff_B_XvmBW3hC8_1(.din(n620),.dout(w_dff_B_XvmBW3hC8_1),.clk(gclk));
	jdff dff_B_skb62kuA6_1(.din(w_dff_B_XvmBW3hC8_1),.dout(w_dff_B_skb62kuA6_1),.clk(gclk));
	jdff dff_B_P7LsQFV40_1(.din(w_dff_B_skb62kuA6_1),.dout(w_dff_B_P7LsQFV40_1),.clk(gclk));
	jdff dff_B_DN46X9li4_1(.din(w_dff_B_P7LsQFV40_1),.dout(w_dff_B_DN46X9li4_1),.clk(gclk));
	jdff dff_B_W5HpanmD0_1(.din(n621),.dout(w_dff_B_W5HpanmD0_1),.clk(gclk));
	jdff dff_B_FNWAFQOO8_1(.din(w_dff_B_W5HpanmD0_1),.dout(w_dff_B_FNWAFQOO8_1),.clk(gclk));
	jdff dff_B_xZN7lzeh2_1(.din(w_dff_B_FNWAFQOO8_1),.dout(w_dff_B_xZN7lzeh2_1),.clk(gclk));
	jdff dff_B_arJKPxfw8_1(.din(w_dff_B_xZN7lzeh2_1),.dout(w_dff_B_arJKPxfw8_1),.clk(gclk));
	jdff dff_A_2ydoM0Lz3_0(.dout(w_G4526_2[0]),.din(w_dff_A_2ydoM0Lz3_0),.clk(gclk));
	jdff dff_A_0Q5F53ju8_0(.dout(w_dff_A_2ydoM0Lz3_0),.din(w_dff_A_0Q5F53ju8_0),.clk(gclk));
	jdff dff_A_eGfvfQ5k5_0(.dout(w_dff_A_0Q5F53ju8_0),.din(w_dff_A_eGfvfQ5k5_0),.clk(gclk));
	jdff dff_A_sYy0gg4E5_1(.dout(w_G4526_2[1]),.din(w_dff_A_sYy0gg4E5_1),.clk(gclk));
	jdff dff_A_HTS5qAX63_1(.dout(w_dff_A_sYy0gg4E5_1),.din(w_dff_A_HTS5qAX63_1),.clk(gclk));
	jdff dff_A_rWmUNWKg4_1(.dout(w_dff_A_HTS5qAX63_1),.din(w_dff_A_rWmUNWKg4_1),.clk(gclk));
	jdff dff_A_1qpZwEpq4_1(.dout(w_dff_A_rWmUNWKg4_1),.din(w_dff_A_1qpZwEpq4_1),.clk(gclk));
	jdff dff_A_fj54Z1BF9_1(.dout(w_dff_A_1qpZwEpq4_1),.din(w_dff_A_fj54Z1BF9_1),.clk(gclk));
	jdff dff_A_HL8nOjL58_1(.dout(w_dff_A_fj54Z1BF9_1),.din(w_dff_A_HL8nOjL58_1),.clk(gclk));
	jdff dff_A_dzxADrtF4_1(.dout(w_dff_A_HL8nOjL58_1),.din(w_dff_A_dzxADrtF4_1),.clk(gclk));
	jdff dff_A_U4zVM82Y9_0(.dout(w_n588_0[0]),.din(w_dff_A_U4zVM82Y9_0),.clk(gclk));
	jdff dff_A_n9LvWGKt4_0(.dout(w_dff_A_U4zVM82Y9_0),.din(w_dff_A_n9LvWGKt4_0),.clk(gclk));
	jdff dff_A_M2ofONVP6_0(.dout(w_dff_A_n9LvWGKt4_0),.din(w_dff_A_M2ofONVP6_0),.clk(gclk));
	jdff dff_A_p6MopZZu3_0(.dout(w_dff_A_M2ofONVP6_0),.din(w_dff_A_p6MopZZu3_0),.clk(gclk));
	jdff dff_A_ahdM1dSZ2_0(.dout(w_dff_A_p6MopZZu3_0),.din(w_dff_A_ahdM1dSZ2_0),.clk(gclk));
	jdff dff_A_Z2ePpNmk0_0(.dout(w_dff_A_ahdM1dSZ2_0),.din(w_dff_A_Z2ePpNmk0_0),.clk(gclk));
	jdff dff_A_TutWKrlk6_0(.dout(w_dff_A_Z2ePpNmk0_0),.din(w_dff_A_TutWKrlk6_0),.clk(gclk));
	jdff dff_A_npGINIGV7_0(.dout(w_dff_A_TutWKrlk6_0),.din(w_dff_A_npGINIGV7_0),.clk(gclk));
	jdff dff_A_iIlM0pb63_0(.dout(w_dff_A_npGINIGV7_0),.din(w_dff_A_iIlM0pb63_0),.clk(gclk));
	jdff dff_A_SApXtcds4_0(.dout(w_dff_A_iIlM0pb63_0),.din(w_dff_A_SApXtcds4_0),.clk(gclk));
	jdff dff_A_I8ZCmTMw6_0(.dout(w_dff_A_SApXtcds4_0),.din(w_dff_A_I8ZCmTMw6_0),.clk(gclk));
	jdff dff_A_zL1CMt5T3_1(.dout(w_n586_0[1]),.din(w_dff_A_zL1CMt5T3_1),.clk(gclk));
	jdff dff_A_zdNmMN4z5_1(.dout(w_dff_A_zL1CMt5T3_1),.din(w_dff_A_zdNmMN4z5_1),.clk(gclk));
	jdff dff_A_Kutyw1wQ0_1(.dout(w_dff_A_zdNmMN4z5_1),.din(w_dff_A_Kutyw1wQ0_1),.clk(gclk));
	jdff dff_A_cVl90BdP7_1(.dout(w_dff_A_Kutyw1wQ0_1),.din(w_dff_A_cVl90BdP7_1),.clk(gclk));
	jdff dff_A_tWk0h5Mk6_1(.dout(w_dff_A_cVl90BdP7_1),.din(w_dff_A_tWk0h5Mk6_1),.clk(gclk));
	jdff dff_A_ONqJEs5t9_1(.dout(w_dff_A_tWk0h5Mk6_1),.din(w_dff_A_ONqJEs5t9_1),.clk(gclk));
	jdff dff_A_2RymdssX3_1(.dout(w_dff_A_ONqJEs5t9_1),.din(w_dff_A_2RymdssX3_1),.clk(gclk));
	jdff dff_A_gnpfGqTm5_1(.dout(w_dff_A_2RymdssX3_1),.din(w_dff_A_gnpfGqTm5_1),.clk(gclk));
	jdff dff_A_JJmyLzV54_1(.dout(w_dff_A_gnpfGqTm5_1),.din(w_dff_A_JJmyLzV54_1),.clk(gclk));
	jdff dff_A_7g1m9XmN6_1(.dout(w_dff_A_JJmyLzV54_1),.din(w_dff_A_7g1m9XmN6_1),.clk(gclk));
	jdff dff_A_MTC5u9nW3_1(.dout(w_dff_A_7g1m9XmN6_1),.din(w_dff_A_MTC5u9nW3_1),.clk(gclk));
	jdff dff_A_Kvr04JiN4_1(.dout(w_dff_A_MTC5u9nW3_1),.din(w_dff_A_Kvr04JiN4_1),.clk(gclk));
	jdff dff_A_UOjkKZjf8_1(.dout(w_dff_A_Kvr04JiN4_1),.din(w_dff_A_UOjkKZjf8_1),.clk(gclk));
	jdff dff_A_vf1lO32r1_2(.dout(w_n586_0[2]),.din(w_dff_A_vf1lO32r1_2),.clk(gclk));
	jdff dff_A_I6NJZyvv3_2(.dout(w_dff_A_vf1lO32r1_2),.din(w_dff_A_I6NJZyvv3_2),.clk(gclk));
	jdff dff_A_tpefdaWu0_2(.dout(w_dff_A_I6NJZyvv3_2),.din(w_dff_A_tpefdaWu0_2),.clk(gclk));
	jdff dff_A_xg2SzjY73_2(.dout(w_dff_A_tpefdaWu0_2),.din(w_dff_A_xg2SzjY73_2),.clk(gclk));
	jdff dff_A_HtcKTuk79_2(.dout(w_dff_A_xg2SzjY73_2),.din(w_dff_A_HtcKTuk79_2),.clk(gclk));
	jdff dff_A_z767cB1A0_2(.dout(w_dff_A_HtcKTuk79_2),.din(w_dff_A_z767cB1A0_2),.clk(gclk));
	jdff dff_A_LwSPtd0c8_2(.dout(w_dff_A_z767cB1A0_2),.din(w_dff_A_LwSPtd0c8_2),.clk(gclk));
	jdff dff_A_68v2XJIJ9_2(.dout(w_dff_A_LwSPtd0c8_2),.din(w_dff_A_68v2XJIJ9_2),.clk(gclk));
	jdff dff_A_uNmMGJuS4_2(.dout(w_dff_A_68v2XJIJ9_2),.din(w_dff_A_uNmMGJuS4_2),.clk(gclk));
	jdff dff_A_Sm5KmY0V8_2(.dout(w_dff_A_uNmMGJuS4_2),.din(w_dff_A_Sm5KmY0V8_2),.clk(gclk));
	jdff dff_A_zAvLW0qS0_2(.dout(w_dff_A_Sm5KmY0V8_2),.din(w_dff_A_zAvLW0qS0_2),.clk(gclk));
	jdff dff_A_3mdVLWpU8_2(.dout(w_dff_A_zAvLW0qS0_2),.din(w_dff_A_3mdVLWpU8_2),.clk(gclk));
	jdff dff_A_Jif3DlyP9_2(.dout(w_dff_A_3mdVLWpU8_2),.din(w_dff_A_Jif3DlyP9_2),.clk(gclk));
	jdff dff_B_sazdHijE6_0(.din(n1631),.dout(w_dff_B_sazdHijE6_0),.clk(gclk));
	jdff dff_B_SrJEm8ST2_0(.din(w_dff_B_sazdHijE6_0),.dout(w_dff_B_SrJEm8ST2_0),.clk(gclk));
	jdff dff_B_Q71OLlIm8_0(.din(w_dff_B_SrJEm8ST2_0),.dout(w_dff_B_Q71OLlIm8_0),.clk(gclk));
	jdff dff_B_yLAvauhF0_0(.din(w_dff_B_Q71OLlIm8_0),.dout(w_dff_B_yLAvauhF0_0),.clk(gclk));
	jdff dff_B_roJCGVcF8_0(.din(w_dff_B_yLAvauhF0_0),.dout(w_dff_B_roJCGVcF8_0),.clk(gclk));
	jdff dff_B_8LVKQobM8_0(.din(w_dff_B_roJCGVcF8_0),.dout(w_dff_B_8LVKQobM8_0),.clk(gclk));
	jdff dff_B_bzKPX9cf4_0(.din(w_dff_B_8LVKQobM8_0),.dout(w_dff_B_bzKPX9cf4_0),.clk(gclk));
	jdff dff_B_d1aAI8ly4_0(.din(w_dff_B_bzKPX9cf4_0),.dout(w_dff_B_d1aAI8ly4_0),.clk(gclk));
	jdff dff_B_Az2yaSxJ4_0(.din(w_dff_B_d1aAI8ly4_0),.dout(w_dff_B_Az2yaSxJ4_0),.clk(gclk));
	jdff dff_B_ozeg8SWK8_0(.din(w_dff_B_Az2yaSxJ4_0),.dout(w_dff_B_ozeg8SWK8_0),.clk(gclk));
	jdff dff_B_dE3sVdpW8_0(.din(w_dff_B_ozeg8SWK8_0),.dout(w_dff_B_dE3sVdpW8_0),.clk(gclk));
	jdff dff_B_N05BqhbP3_1(.din(n1621),.dout(w_dff_B_N05BqhbP3_1),.clk(gclk));
	jdff dff_B_NIqczoov3_1(.din(w_dff_B_N05BqhbP3_1),.dout(w_dff_B_NIqczoov3_1),.clk(gclk));
	jdff dff_B_qI4S16l17_1(.din(n1622),.dout(w_dff_B_qI4S16l17_1),.clk(gclk));
	jdff dff_A_3xDhesA69_0(.dout(w_n1620_0[0]),.din(w_dff_A_3xDhesA69_0),.clk(gclk));
	jdff dff_A_o1ibeUd56_0(.dout(w_dff_A_3xDhesA69_0),.din(w_dff_A_o1ibeUd56_0),.clk(gclk));
	jdff dff_B_pLSfkFdq2_0(.din(n1617),.dout(w_dff_B_pLSfkFdq2_0),.clk(gclk));
	jdff dff_B_r2mzG9rG0_0(.din(w_dff_B_pLSfkFdq2_0),.dout(w_dff_B_r2mzG9rG0_0),.clk(gclk));
	jdff dff_B_6dtNDip40_1(.din(n1611),.dout(w_dff_B_6dtNDip40_1),.clk(gclk));
	jdff dff_B_9hQjcZU16_1(.din(w_dff_B_6dtNDip40_1),.dout(w_dff_B_9hQjcZU16_1),.clk(gclk));
	jdff dff_B_pGs50NTd7_1(.din(n1608),.dout(w_dff_B_pGs50NTd7_1),.clk(gclk));
	jdff dff_B_9fCmHICZ8_0(.din(n1609),.dout(w_dff_B_9fCmHICZ8_0),.clk(gclk));
	jdff dff_B_2NxGL0PU0_0(.din(w_dff_B_9fCmHICZ8_0),.dout(w_dff_B_2NxGL0PU0_0),.clk(gclk));
	jdff dff_B_oOQZMAY02_0(.din(w_dff_B_2NxGL0PU0_0),.dout(w_dff_B_oOQZMAY02_0),.clk(gclk));
	jdff dff_B_uBDpo2xi1_0(.din(w_dff_B_oOQZMAY02_0),.dout(w_dff_B_uBDpo2xi1_0),.clk(gclk));
	jdff dff_B_fEle8DqW2_0(.din(w_dff_B_uBDpo2xi1_0),.dout(w_dff_B_fEle8DqW2_0),.clk(gclk));
	jdff dff_A_T9LZAj526_0(.dout(w_n1607_0[0]),.din(w_dff_A_T9LZAj526_0),.clk(gclk));
	jdff dff_A_OtQD0IBF3_0(.dout(w_dff_A_T9LZAj526_0),.din(w_dff_A_OtQD0IBF3_0),.clk(gclk));
	jdff dff_A_6NPsbDMG0_0(.dout(w_dff_A_OtQD0IBF3_0),.din(w_dff_A_6NPsbDMG0_0),.clk(gclk));
	jdff dff_B_5Ifwxcif7_0(.din(n1606),.dout(w_dff_B_5Ifwxcif7_0),.clk(gclk));
	jdff dff_A_UWlumCSz6_0(.dout(w_n1605_0[0]),.din(w_dff_A_UWlumCSz6_0),.clk(gclk));
	jdff dff_A_r61HzQDy6_0(.dout(w_dff_A_UWlumCSz6_0),.din(w_dff_A_r61HzQDy6_0),.clk(gclk));
	jdff dff_A_tf5p52Ec4_0(.dout(w_dff_A_r61HzQDy6_0),.din(w_dff_A_tf5p52Ec4_0),.clk(gclk));
	jdff dff_A_dPrAgsv13_0(.dout(w_dff_A_tf5p52Ec4_0),.din(w_dff_A_dPrAgsv13_0),.clk(gclk));
	jdff dff_A_dOaRQNjy6_0(.dout(w_dff_A_dPrAgsv13_0),.din(w_dff_A_dOaRQNjy6_0),.clk(gclk));
	jdff dff_B_NWmQF8Ab9_0(.din(n1603),.dout(w_dff_B_NWmQF8Ab9_0),.clk(gclk));
	jdff dff_B_YtMXNCep7_1(.din(n1588),.dout(w_dff_B_YtMXNCep7_1),.clk(gclk));
	jdff dff_A_cU7m0Lw71_1(.dout(w_n1597_0[1]),.din(w_dff_A_cU7m0Lw71_1),.clk(gclk));
	jdff dff_B_w8rOjI4n1_2(.din(n1597),.dout(w_dff_B_w8rOjI4n1_2),.clk(gclk));
	jdff dff_B_3XopZPmy5_0(.din(n1596),.dout(w_dff_B_3XopZPmy5_0),.clk(gclk));
	jdff dff_B_vR2uCBVR6_0(.din(n1595),.dout(w_dff_B_vR2uCBVR6_0),.clk(gclk));
	jdff dff_B_3KXtXQqc2_0(.din(w_dff_B_vR2uCBVR6_0),.dout(w_dff_B_3KXtXQqc2_0),.clk(gclk));
	jdff dff_B_ZmV7R1xK6_0(.din(w_dff_B_3KXtXQqc2_0),.dout(w_dff_B_ZmV7R1xK6_0),.clk(gclk));
	jdff dff_B_0XqqsElB1_0(.din(n1592),.dout(w_dff_B_0XqqsElB1_0),.clk(gclk));
	jdff dff_A_LuCcrrTp7_1(.dout(w_n1106_0[1]),.din(w_dff_A_LuCcrrTp7_1),.clk(gclk));
	jdff dff_A_YmjYPiIJ5_1(.dout(w_dff_A_LuCcrrTp7_1),.din(w_dff_A_YmjYPiIJ5_1),.clk(gclk));
	jdff dff_A_4RzCVLNv9_1(.dout(w_dff_A_YmjYPiIJ5_1),.din(w_dff_A_4RzCVLNv9_1),.clk(gclk));
	jdff dff_A_RvvrxBSi0_1(.dout(w_dff_A_4RzCVLNv9_1),.din(w_dff_A_RvvrxBSi0_1),.clk(gclk));
	jdff dff_A_C86U8i2H1_1(.dout(w_dff_A_RvvrxBSi0_1),.din(w_dff_A_C86U8i2H1_1),.clk(gclk));
	jdff dff_A_b9c2Mbgn9_1(.dout(w_dff_A_C86U8i2H1_1),.din(w_dff_A_b9c2Mbgn9_1),.clk(gclk));
	jdff dff_A_r3qnJ5C00_1(.dout(w_dff_A_b9c2Mbgn9_1),.din(w_dff_A_r3qnJ5C00_1),.clk(gclk));
	jdff dff_A_QtZCvjht7_1(.dout(w_dff_A_r3qnJ5C00_1),.din(w_dff_A_QtZCvjht7_1),.clk(gclk));
	jdff dff_A_BZUMQKgO2_1(.dout(w_dff_A_QtZCvjht7_1),.din(w_dff_A_BZUMQKgO2_1),.clk(gclk));
	jdff dff_A_Da3PXiuw3_1(.dout(w_dff_A_BZUMQKgO2_1),.din(w_dff_A_Da3PXiuw3_1),.clk(gclk));
	jdff dff_A_GpkEY0jh0_1(.dout(w_n619_0[1]),.din(w_dff_A_GpkEY0jh0_1),.clk(gclk));
	jdff dff_A_J8hwEzkF8_1(.dout(w_dff_A_GpkEY0jh0_1),.din(w_dff_A_J8hwEzkF8_1),.clk(gclk));
	jdff dff_A_xIQ7gbAj8_1(.dout(w_dff_A_J8hwEzkF8_1),.din(w_dff_A_xIQ7gbAj8_1),.clk(gclk));
	jdff dff_A_HG3c8mgp8_1(.dout(w_dff_A_xIQ7gbAj8_1),.din(w_dff_A_HG3c8mgp8_1),.clk(gclk));
	jdff dff_A_9j1YVS9y4_1(.dout(w_dff_A_HG3c8mgp8_1),.din(w_dff_A_9j1YVS9y4_1),.clk(gclk));
	jdff dff_B_9MsAzG8q7_1(.din(n607),.dout(w_dff_B_9MsAzG8q7_1),.clk(gclk));
	jdff dff_B_Q8FR69JP3_1(.din(w_dff_B_9MsAzG8q7_1),.dout(w_dff_B_Q8FR69JP3_1),.clk(gclk));
	jdff dff_A_SXs6JVZ94_0(.dout(w_n618_0[0]),.din(w_dff_A_SXs6JVZ94_0),.clk(gclk));
	jdff dff_A_Av51p9Z88_0(.dout(w_dff_A_SXs6JVZ94_0),.din(w_dff_A_Av51p9Z88_0),.clk(gclk));
	jdff dff_A_3GBMsHpT0_0(.dout(w_dff_A_Av51p9Z88_0),.din(w_dff_A_3GBMsHpT0_0),.clk(gclk));
	jdff dff_A_h8BPYLPv4_0(.dout(w_dff_A_3GBMsHpT0_0),.din(w_dff_A_h8BPYLPv4_0),.clk(gclk));
	jdff dff_A_4HO5pGpq3_0(.dout(w_dff_A_h8BPYLPv4_0),.din(w_dff_A_4HO5pGpq3_0),.clk(gclk));
	jdff dff_B_R97nAaRo7_1(.din(n611),.dout(w_dff_B_R97nAaRo7_1),.clk(gclk));
	jdff dff_B_1aY1013Z9_1(.din(w_dff_B_R97nAaRo7_1),.dout(w_dff_B_1aY1013Z9_1),.clk(gclk));
	jdff dff_A_Rq9lncRI9_0(.dout(w_n605_0[0]),.din(w_dff_A_Rq9lncRI9_0),.clk(gclk));
	jdff dff_A_tPE7GcZP7_0(.dout(w_dff_A_Rq9lncRI9_0),.din(w_dff_A_tPE7GcZP7_0),.clk(gclk));
	jdff dff_A_2CcqA3Wp5_1(.dout(w_n605_0[1]),.din(w_dff_A_2CcqA3Wp5_1),.clk(gclk));
	jdff dff_A_A4Tkes5G2_1(.dout(w_dff_A_2CcqA3Wp5_1),.din(w_dff_A_A4Tkes5G2_1),.clk(gclk));
	jdff dff_A_5mzia1uA7_1(.dout(w_dff_A_A4Tkes5G2_1),.din(w_dff_A_5mzia1uA7_1),.clk(gclk));
	jdff dff_A_TNobmL449_1(.dout(w_dff_A_5mzia1uA7_1),.din(w_dff_A_TNobmL449_1),.clk(gclk));
	jdff dff_A_AZoqO2o88_1(.dout(w_dff_A_TNobmL449_1),.din(w_dff_A_AZoqO2o88_1),.clk(gclk));
	jdff dff_A_tYXA1acM7_1(.dout(w_dff_A_AZoqO2o88_1),.din(w_dff_A_tYXA1acM7_1),.clk(gclk));
	jdff dff_A_794GiRhN5_1(.dout(w_dff_A_tYXA1acM7_1),.din(w_dff_A_794GiRhN5_1),.clk(gclk));
	jdff dff_A_gnJKtLYn9_1(.dout(w_dff_A_794GiRhN5_1),.din(w_dff_A_gnJKtLYn9_1),.clk(gclk));
	jdff dff_A_0KXMix2R7_1(.dout(w_dff_A_gnJKtLYn9_1),.din(w_dff_A_0KXMix2R7_1),.clk(gclk));
	jdff dff_A_a6MHcINx3_0(.dout(w_n604_0[0]),.din(w_dff_A_a6MHcINx3_0),.clk(gclk));
	jdff dff_A_P0ECXsiM0_0(.dout(w_dff_A_a6MHcINx3_0),.din(w_dff_A_P0ECXsiM0_0),.clk(gclk));
	jdff dff_A_K58WcmBV6_0(.dout(w_dff_A_P0ECXsiM0_0),.din(w_dff_A_K58WcmBV6_0),.clk(gclk));
	jdff dff_A_f7lECtP44_0(.dout(w_dff_A_K58WcmBV6_0),.din(w_dff_A_f7lECtP44_0),.clk(gclk));
	jdff dff_A_9nNDEB4q5_0(.dout(w_dff_A_f7lECtP44_0),.din(w_dff_A_9nNDEB4q5_0),.clk(gclk));
	jdff dff_A_tvzVDIrl0_0(.dout(w_dff_A_9nNDEB4q5_0),.din(w_dff_A_tvzVDIrl0_0),.clk(gclk));
	jdff dff_A_4odcy0QT3_0(.dout(w_dff_A_tvzVDIrl0_0),.din(w_dff_A_4odcy0QT3_0),.clk(gclk));
	jdff dff_A_emGEHPlv5_0(.dout(w_dff_A_4odcy0QT3_0),.din(w_dff_A_emGEHPlv5_0),.clk(gclk));
	jdff dff_A_FLmQyZFF2_0(.dout(w_dff_A_emGEHPlv5_0),.din(w_dff_A_FLmQyZFF2_0),.clk(gclk));
	jdff dff_A_eybIkGQx0_0(.dout(w_dff_A_FLmQyZFF2_0),.din(w_dff_A_eybIkGQx0_0),.clk(gclk));
	jdff dff_A_dDpbM4O12_1(.dout(w_n594_0[1]),.din(w_dff_A_dDpbM4O12_1),.clk(gclk));
	jdff dff_A_L6t83EmZ4_1(.dout(w_dff_A_dDpbM4O12_1),.din(w_dff_A_L6t83EmZ4_1),.clk(gclk));
	jdff dff_A_fzUHu6em2_1(.dout(w_dff_A_L6t83EmZ4_1),.din(w_dff_A_fzUHu6em2_1),.clk(gclk));
	jdff dff_A_6BKBDSwR7_1(.dout(w_dff_A_fzUHu6em2_1),.din(w_dff_A_6BKBDSwR7_1),.clk(gclk));
	jdff dff_A_S8jMWJYh0_1(.dout(w_dff_A_6BKBDSwR7_1),.din(w_dff_A_S8jMWJYh0_1),.clk(gclk));
	jdff dff_A_baKVXvgD7_1(.dout(w_dff_A_S8jMWJYh0_1),.din(w_dff_A_baKVXvgD7_1),.clk(gclk));
	jdff dff_A_LVitKlWq9_1(.dout(w_dff_A_baKVXvgD7_1),.din(w_dff_A_LVitKlWq9_1),.clk(gclk));
	jdff dff_A_HZOXCUEY6_1(.dout(w_dff_A_LVitKlWq9_1),.din(w_dff_A_HZOXCUEY6_1),.clk(gclk));
	jdff dff_A_wlaO9dSU5_1(.dout(w_dff_A_HZOXCUEY6_1),.din(w_dff_A_wlaO9dSU5_1),.clk(gclk));
	jdff dff_A_bykxBIGm9_1(.dout(w_dff_A_wlaO9dSU5_1),.din(w_dff_A_bykxBIGm9_1),.clk(gclk));
	jdff dff_A_7SqSx9tl8_1(.dout(w_dff_A_bykxBIGm9_1),.din(w_dff_A_7SqSx9tl8_1),.clk(gclk));
	jdff dff_A_kmmA1FoC8_1(.dout(w_dff_A_7SqSx9tl8_1),.din(w_dff_A_kmmA1FoC8_1),.clk(gclk));
	jdff dff_A_R7HIKgfX4_2(.dout(w_n594_0[2]),.din(w_dff_A_R7HIKgfX4_2),.clk(gclk));
	jdff dff_B_vH4nvQFC5_1(.din(n650),.dout(w_dff_B_vH4nvQFC5_1),.clk(gclk));
	jdff dff_B_AjURoX3e3_1(.din(w_dff_B_vH4nvQFC5_1),.dout(w_dff_B_AjURoX3e3_1),.clk(gclk));
	jdff dff_B_H3ACOtNF0_1(.din(w_dff_B_AjURoX3e3_1),.dout(w_dff_B_H3ACOtNF0_1),.clk(gclk));
	jdff dff_B_KOksx7kp3_1(.din(w_dff_B_H3ACOtNF0_1),.dout(w_dff_B_KOksx7kp3_1),.clk(gclk));
	jdff dff_A_Bwoqm0jQ7_0(.dout(w_n666_0[0]),.din(w_dff_A_Bwoqm0jQ7_0),.clk(gclk));
	jdff dff_A_9oJWk3Pj8_0(.dout(w_n664_0[0]),.din(w_dff_A_9oJWk3Pj8_0),.clk(gclk));
	jdff dff_A_nBMtiG5B5_0(.dout(w_dff_A_9oJWk3Pj8_0),.din(w_dff_A_nBMtiG5B5_0),.clk(gclk));
	jdff dff_B_eLWVEYyq7_2(.din(n664),.dout(w_dff_B_eLWVEYyq7_2),.clk(gclk));
	jdff dff_A_UqyDJu4D5_1(.dout(w_n662_0[1]),.din(w_dff_A_UqyDJu4D5_1),.clk(gclk));
	jdff dff_A_Icd7JuWI5_1(.dout(w_n661_0[1]),.din(w_dff_A_Icd7JuWI5_1),.clk(gclk));
	jdff dff_A_RwBj1TKk8_1(.dout(w_dff_A_Icd7JuWI5_1),.din(w_dff_A_RwBj1TKk8_1),.clk(gclk));
	jdff dff_A_kXj7iwpq7_1(.dout(w_dff_A_RwBj1TKk8_1),.din(w_dff_A_kXj7iwpq7_1),.clk(gclk));
	jdff dff_A_yUGoHWWg2_2(.dout(w_n661_0[2]),.din(w_dff_A_yUGoHWWg2_2),.clk(gclk));
	jdff dff_B_pTaV3zpz2_1(.din(n658),.dout(w_dff_B_pTaV3zpz2_1),.clk(gclk));
	jdff dff_A_kF5LMZdN8_1(.dout(w_n657_0[1]),.din(w_dff_A_kF5LMZdN8_1),.clk(gclk));
	jdff dff_A_A1OPI00p8_1(.dout(w_dff_A_kF5LMZdN8_1),.din(w_dff_A_A1OPI00p8_1),.clk(gclk));
	jdff dff_A_v4wmxwJL6_2(.dout(w_n657_0[2]),.din(w_dff_A_v4wmxwJL6_2),.clk(gclk));
	jdff dff_A_2GrllwjR3_2(.dout(w_dff_A_v4wmxwJL6_2),.din(w_dff_A_2GrllwjR3_2),.clk(gclk));
	jdff dff_A_PZOFBsFT3_0(.dout(w_n653_0[0]),.din(w_dff_A_PZOFBsFT3_0),.clk(gclk));
	jdff dff_A_kjJgJEyu9_0(.dout(w_dff_A_PZOFBsFT3_0),.din(w_dff_A_kjJgJEyu9_0),.clk(gclk));
	jdff dff_A_UjSvI0Ny8_0(.dout(w_dff_A_kjJgJEyu9_0),.din(w_dff_A_UjSvI0Ny8_0),.clk(gclk));
	jdff dff_B_5lt25F7C8_2(.din(n653),.dout(w_dff_B_5lt25F7C8_2),.clk(gclk));
	jdff dff_B_uoIN38tW4_2(.din(w_dff_B_5lt25F7C8_2),.dout(w_dff_B_uoIN38tW4_2),.clk(gclk));
	jdff dff_B_aEhxahxj8_2(.din(w_dff_B_uoIN38tW4_2),.dout(w_dff_B_aEhxahxj8_2),.clk(gclk));
	jdff dff_A_Rkv4QTmw4_0(.dout(w_n1094_0[0]),.din(w_dff_A_Rkv4QTmw4_0),.clk(gclk));
	jdff dff_A_dEMNL1jD3_1(.dout(w_n1094_0[1]),.din(w_dff_A_dEMNL1jD3_1),.clk(gclk));
	jdff dff_A_dlGEQ5aM2_1(.dout(w_dff_A_dEMNL1jD3_1),.din(w_dff_A_dlGEQ5aM2_1),.clk(gclk));
	jdff dff_B_uHsnKISb7_3(.din(n1094),.dout(w_dff_B_uHsnKISb7_3),.clk(gclk));
	jdff dff_B_HCaRfry94_3(.din(w_dff_B_uHsnKISb7_3),.dout(w_dff_B_HCaRfry94_3),.clk(gclk));
	jdff dff_B_CHuIJ1FZ5_3(.din(w_dff_B_HCaRfry94_3),.dout(w_dff_B_CHuIJ1FZ5_3),.clk(gclk));
	jdff dff_B_YKTqkjlu3_3(.din(w_dff_B_CHuIJ1FZ5_3),.dout(w_dff_B_YKTqkjlu3_3),.clk(gclk));
	jdff dff_B_GBC6tgsS0_3(.din(w_dff_B_YKTqkjlu3_3),.dout(w_dff_B_GBC6tgsS0_3),.clk(gclk));
	jdff dff_B_fNNYFwtv6_3(.din(w_dff_B_GBC6tgsS0_3),.dout(w_dff_B_fNNYFwtv6_3),.clk(gclk));
	jdff dff_B_vRBwmbzP8_3(.din(w_dff_B_fNNYFwtv6_3),.dout(w_dff_B_vRBwmbzP8_3),.clk(gclk));
	jdff dff_B_Zzbkcf9B6_3(.din(w_dff_B_vRBwmbzP8_3),.dout(w_dff_B_Zzbkcf9B6_3),.clk(gclk));
	jdff dff_B_jM3c1MzT9_3(.din(w_dff_B_Zzbkcf9B6_3),.dout(w_dff_B_jM3c1MzT9_3),.clk(gclk));
	jdff dff_B_EsOLP7h00_3(.din(w_dff_B_jM3c1MzT9_3),.dout(w_dff_B_EsOLP7h00_3),.clk(gclk));
	jdff dff_B_18wAMXjE5_3(.din(w_dff_B_EsOLP7h00_3),.dout(w_dff_B_18wAMXjE5_3),.clk(gclk));
	jdff dff_A_ZB8TSSX78_0(.dout(w_G4526_1[0]),.din(w_dff_A_ZB8TSSX78_0),.clk(gclk));
	jdff dff_A_e4bLKr3j3_0(.dout(w_dff_A_ZB8TSSX78_0),.din(w_dff_A_e4bLKr3j3_0),.clk(gclk));
	jdff dff_A_C5lxxWGP2_0(.dout(w_dff_A_e4bLKr3j3_0),.din(w_dff_A_C5lxxWGP2_0),.clk(gclk));
	jdff dff_A_SFO0hwky9_0(.dout(w_dff_A_C5lxxWGP2_0),.din(w_dff_A_SFO0hwky9_0),.clk(gclk));
	jdff dff_A_NT4AtEq80_0(.dout(w_dff_A_SFO0hwky9_0),.din(w_dff_A_NT4AtEq80_0),.clk(gclk));
	jdff dff_A_fQAJd3EL8_0(.dout(w_dff_A_NT4AtEq80_0),.din(w_dff_A_fQAJd3EL8_0),.clk(gclk));
	jdff dff_A_5yjwNBpz2_0(.dout(w_dff_A_fQAJd3EL8_0),.din(w_dff_A_5yjwNBpz2_0),.clk(gclk));
	jdff dff_A_SelS453N1_0(.dout(w_dff_A_5yjwNBpz2_0),.din(w_dff_A_SelS453N1_0),.clk(gclk));
	jdff dff_A_qrO3UpGs9_0(.dout(w_dff_A_SelS453N1_0),.din(w_dff_A_qrO3UpGs9_0),.clk(gclk));
	jdff dff_A_p2bKUdqv7_0(.dout(w_dff_A_qrO3UpGs9_0),.din(w_dff_A_p2bKUdqv7_0),.clk(gclk));
	jdff dff_A_WH1e1dBZ8_0(.dout(w_dff_A_p2bKUdqv7_0),.din(w_dff_A_WH1e1dBZ8_0),.clk(gclk));
	jdff dff_A_4Iu5KSXc9_0(.dout(w_dff_A_WH1e1dBZ8_0),.din(w_dff_A_4Iu5KSXc9_0),.clk(gclk));
	jdff dff_A_rkpjtdP25_0(.dout(w_dff_A_4Iu5KSXc9_0),.din(w_dff_A_rkpjtdP25_0),.clk(gclk));
	jdff dff_A_WgW83LfH5_0(.dout(w_dff_A_rkpjtdP25_0),.din(w_dff_A_WgW83LfH5_0),.clk(gclk));
	jdff dff_A_XxhC2lv49_2(.dout(w_G4526_1[2]),.din(w_dff_A_XxhC2lv49_2),.clk(gclk));
	jdff dff_A_KjHWuwaD6_2(.dout(w_dff_A_XxhC2lv49_2),.din(w_dff_A_KjHWuwaD6_2),.clk(gclk));
	jdff dff_A_wROp01Cy2_2(.dout(w_dff_A_KjHWuwaD6_2),.din(w_dff_A_wROp01Cy2_2),.clk(gclk));
	jdff dff_A_N2XdCU0N8_2(.dout(w_dff_A_wROp01Cy2_2),.din(w_dff_A_N2XdCU0N8_2),.clk(gclk));
	jdff dff_A_vIdPQ6qN6_2(.dout(w_dff_A_N2XdCU0N8_2),.din(w_dff_A_vIdPQ6qN6_2),.clk(gclk));
	jdff dff_A_kaQKAcE87_1(.dout(w_G4526_0[1]),.din(w_dff_A_kaQKAcE87_1),.clk(gclk));
	jdff dff_A_pQu3n5bo0_1(.dout(w_dff_A_kaQKAcE87_1),.din(w_dff_A_pQu3n5bo0_1),.clk(gclk));
	jdff dff_A_rof2vaeC3_1(.dout(w_dff_A_pQu3n5bo0_1),.din(w_dff_A_rof2vaeC3_1),.clk(gclk));
	jdff dff_A_KzlUK4uX4_1(.dout(w_dff_A_rof2vaeC3_1),.din(w_dff_A_KzlUK4uX4_1),.clk(gclk));
	jdff dff_A_AAVX09nF5_1(.dout(w_dff_A_KzlUK4uX4_1),.din(w_dff_A_AAVX09nF5_1),.clk(gclk));
	jdff dff_A_WFnPfGsW1_2(.dout(w_G4526_0[2]),.din(w_dff_A_WFnPfGsW1_2),.clk(gclk));
	jdff dff_A_9fMpdCo01_2(.dout(w_dff_A_WFnPfGsW1_2),.din(w_dff_A_9fMpdCo01_2),.clk(gclk));
	jdff dff_A_xeuuFKas7_2(.dout(w_dff_A_9fMpdCo01_2),.din(w_dff_A_xeuuFKas7_2),.clk(gclk));
	jdff dff_A_n39KGL7a6_2(.dout(w_dff_A_xeuuFKas7_2),.din(w_dff_A_n39KGL7a6_2),.clk(gclk));
	jdff dff_A_1wZzwL965_2(.dout(w_dff_A_n39KGL7a6_2),.din(w_dff_A_1wZzwL965_2),.clk(gclk));
	jdff dff_A_GbpiApuL1_2(.dout(w_dff_A_1wZzwL965_2),.din(w_dff_A_GbpiApuL1_2),.clk(gclk));
	jdff dff_A_iubDQSNR7_2(.dout(w_dff_A_GbpiApuL1_2),.din(w_dff_A_iubDQSNR7_2),.clk(gclk));
	jdff dff_A_zIkDMXcZ8_2(.dout(w_dff_A_iubDQSNR7_2),.din(w_dff_A_zIkDMXcZ8_2),.clk(gclk));
	jdff dff_A_8se1Bysi3_2(.dout(w_dff_A_zIkDMXcZ8_2),.din(w_dff_A_8se1Bysi3_2),.clk(gclk));
	jdff dff_A_dKJHBT0a7_2(.dout(w_dff_A_8se1Bysi3_2),.din(w_dff_A_dKJHBT0a7_2),.clk(gclk));
	jdff dff_A_5gsDfRXy5_2(.dout(w_dff_A_dKJHBT0a7_2),.din(w_dff_A_5gsDfRXy5_2),.clk(gclk));
	jdff dff_A_CThn5KxT9_2(.dout(w_dff_A_5gsDfRXy5_2),.din(w_dff_A_CThn5KxT9_2),.clk(gclk));
	jdff dff_A_M4E1PaT90_2(.dout(w_dff_A_CThn5KxT9_2),.din(w_dff_A_M4E1PaT90_2),.clk(gclk));
	jdff dff_B_B17T1vBb1_0(.din(n1586),.dout(w_dff_B_B17T1vBb1_0),.clk(gclk));
	jdff dff_B_ivaSIiH18_0(.din(w_dff_B_B17T1vBb1_0),.dout(w_dff_B_ivaSIiH18_0),.clk(gclk));
	jdff dff_B_x4WMh0ub5_1(.din(n1582),.dout(w_dff_B_x4WMh0ub5_1),.clk(gclk));
	jdff dff_B_mGxIXwGq5_1(.din(w_dff_B_x4WMh0ub5_1),.dout(w_dff_B_mGxIXwGq5_1),.clk(gclk));
	jdff dff_B_JV2A6PtL3_0(.din(n1584),.dout(w_dff_B_JV2A6PtL3_0),.clk(gclk));
	jdff dff_A_aUsyYBN80_0(.dout(w_n610_0[0]),.din(w_dff_A_aUsyYBN80_0),.clk(gclk));
	jdff dff_A_iag1hkad3_0(.dout(w_dff_A_aUsyYBN80_0),.din(w_dff_A_iag1hkad3_0),.clk(gclk));
	jdff dff_A_8w9F53vG1_1(.dout(w_n590_0[1]),.din(w_dff_A_8w9F53vG1_1),.clk(gclk));
	jdff dff_A_9ZEcId8N2_1(.dout(w_dff_A_8w9F53vG1_1),.din(w_dff_A_9ZEcId8N2_1),.clk(gclk));
	jdff dff_A_pQHBUbia0_2(.dout(w_n590_0[2]),.din(w_dff_A_pQHBUbia0_2),.clk(gclk));
	jdff dff_A_agWuWEKK0_2(.dout(w_dff_A_pQHBUbia0_2),.din(w_dff_A_agWuWEKK0_2),.clk(gclk));
	jdff dff_A_xCO3wEwh1_1(.dout(w_n615_0[1]),.din(w_dff_A_xCO3wEwh1_1),.clk(gclk));
	jdff dff_A_X7auKSNU3_1(.dout(w_dff_A_xCO3wEwh1_1),.din(w_dff_A_X7auKSNU3_1),.clk(gclk));
	jdff dff_A_LkTghKlY6_1(.dout(w_dff_A_X7auKSNU3_1),.din(w_dff_A_LkTghKlY6_1),.clk(gclk));
	jdff dff_A_VZOYcmTX5_1(.dout(w_dff_A_LkTghKlY6_1),.din(w_dff_A_VZOYcmTX5_1),.clk(gclk));
	jdff dff_A_TrvEIaVe4_1(.dout(w_dff_A_VZOYcmTX5_1),.din(w_dff_A_TrvEIaVe4_1),.clk(gclk));
	jdff dff_A_nwt7supn4_1(.dout(w_dff_A_TrvEIaVe4_1),.din(w_dff_A_nwt7supn4_1),.clk(gclk));
	jdff dff_A_QRLz4kkM9_1(.dout(w_dff_A_nwt7supn4_1),.din(w_dff_A_QRLz4kkM9_1),.clk(gclk));
	jdff dff_A_ge2KhoMZ4_1(.dout(w_dff_A_QRLz4kkM9_1),.din(w_dff_A_ge2KhoMZ4_1),.clk(gclk));
	jdff dff_A_6QjljWL94_1(.dout(w_dff_A_ge2KhoMZ4_1),.din(w_dff_A_6QjljWL94_1),.clk(gclk));
	jdff dff_B_bDqZolpk9_2(.din(n600),.dout(w_dff_B_bDqZolpk9_2),.clk(gclk));
	jdff dff_B_BXVAVGHI5_2(.din(w_dff_B_bDqZolpk9_2),.dout(w_dff_B_BXVAVGHI5_2),.clk(gclk));
	jdff dff_A_NJ16sLVB1_1(.dout(w_n612_0[1]),.din(w_dff_A_NJ16sLVB1_1),.clk(gclk));
	jdff dff_A_PWYghY9h1_1(.dout(w_n609_0[1]),.din(w_dff_A_PWYghY9h1_1),.clk(gclk));
	jdff dff_B_XqLl8wJC5_2(.din(n609),.dout(w_dff_B_XqLl8wJC5_2),.clk(gclk));
	jdff dff_B_tJHYdyLG7_2(.din(w_dff_B_XqLl8wJC5_2),.dout(w_dff_B_tJHYdyLG7_2),.clk(gclk));
	jdff dff_B_0Y1cWcdy6_1(.din(n591),.dout(w_dff_B_0Y1cWcdy6_1),.clk(gclk));
	jdff dff_B_Vz2Xni5H6_0(.din(G124),.dout(w_dff_B_Vz2Xni5H6_0),.clk(gclk));
	jdff dff_A_C4MMxLEe2_1(.dout(w_G3743_0[1]),.din(w_dff_A_C4MMxLEe2_1),.clk(gclk));
	jdff dff_A_pDhCs61i9_1(.dout(w_dff_A_C4MMxLEe2_1),.din(w_dff_A_pDhCs61i9_1),.clk(gclk));
	jdff dff_A_1GwjxuQt0_1(.dout(w_dff_A_pDhCs61i9_1),.din(w_dff_A_1GwjxuQt0_1),.clk(gclk));
	jdff dff_A_ggo8CN6V0_1(.dout(w_dff_A_1GwjxuQt0_1),.din(w_dff_A_ggo8CN6V0_1),.clk(gclk));
	jdff dff_A_689w9I3n8_1(.dout(w_n1084_0[1]),.din(w_dff_A_689w9I3n8_1),.clk(gclk));
	jdff dff_A_K5ZrTf5f6_2(.dout(w_n1084_0[2]),.din(w_dff_A_K5ZrTf5f6_2),.clk(gclk));
	jdff dff_A_Hn9NuiWs7_2(.dout(w_dff_A_K5ZrTf5f6_2),.din(w_dff_A_Hn9NuiWs7_2),.clk(gclk));
	jdff dff_A_oezZcvdH4_2(.dout(w_dff_A_Hn9NuiWs7_2),.din(w_dff_A_oezZcvdH4_2),.clk(gclk));
	jdff dff_A_rewglPAF1_2(.dout(w_dff_A_oezZcvdH4_2),.din(w_dff_A_rewglPAF1_2),.clk(gclk));
	jdff dff_A_kvJ3T86d4_2(.dout(w_dff_A_rewglPAF1_2),.din(w_dff_A_kvJ3T86d4_2),.clk(gclk));
	jdff dff_A_fJWjDWHI5_2(.dout(w_dff_A_kvJ3T86d4_2),.din(w_dff_A_fJWjDWHI5_2),.clk(gclk));
	jdff dff_A_QGWFhGrH0_2(.dout(w_dff_A_fJWjDWHI5_2),.din(w_dff_A_QGWFhGrH0_2),.clk(gclk));
	jdff dff_A_kWpWYWT03_2(.dout(w_dff_A_QGWFhGrH0_2),.din(w_dff_A_kWpWYWT03_2),.clk(gclk));
	jdff dff_A_fO1wqDCy3_2(.dout(w_dff_A_kWpWYWT03_2),.din(w_dff_A_fO1wqDCy3_2),.clk(gclk));
	jdff dff_A_rXWtukPu0_2(.dout(w_dff_A_fO1wqDCy3_2),.din(w_dff_A_rXWtukPu0_2),.clk(gclk));
	jdff dff_A_WRFvq4cH9_2(.dout(w_dff_A_rXWtukPu0_2),.din(w_dff_A_WRFvq4cH9_2),.clk(gclk));
	jdff dff_A_zIaVZtZh8_2(.dout(w_dff_A_WRFvq4cH9_2),.din(w_dff_A_zIaVZtZh8_2),.clk(gclk));
	jdff dff_B_izFmWNtm7_1(.din(n583),.dout(w_dff_B_izFmWNtm7_1),.clk(gclk));
	jdff dff_B_pbQHyWMd6_0(.din(G100),.dout(w_dff_B_pbQHyWMd6_0),.clk(gclk));
	jdff dff_A_10QKI3Aw8_0(.dout(w_n582_0[0]),.din(w_dff_A_10QKI3Aw8_0),.clk(gclk));
	jdff dff_A_bSEYi0OK8_0(.dout(w_dff_A_10QKI3Aw8_0),.din(w_dff_A_bSEYi0OK8_0),.clk(gclk));
	jdff dff_A_zKkWUVVK3_2(.dout(w_n582_0[2]),.din(w_dff_A_zKkWUVVK3_2),.clk(gclk));
	jdff dff_A_ouNZOQcj1_2(.dout(w_dff_A_zKkWUVVK3_2),.din(w_dff_A_ouNZOQcj1_2),.clk(gclk));
	jdff dff_A_WlxqNpyP9_1(.dout(w_G3749_0[1]),.din(w_dff_A_WlxqNpyP9_1),.clk(gclk));
	jdff dff_A_JwtNIGmY0_1(.dout(w_dff_A_WlxqNpyP9_1),.din(w_dff_A_JwtNIGmY0_1),.clk(gclk));
	jdff dff_A_ysaxURk58_1(.dout(w_dff_A_JwtNIGmY0_1),.din(w_dff_A_ysaxURk58_1),.clk(gclk));
	jdff dff_A_zBnmxytd5_1(.dout(w_dff_A_ysaxURk58_1),.din(w_dff_A_zBnmxytd5_1),.clk(gclk));
	jdff dff_A_pDtEMtL68_1(.dout(w_n1108_0[1]),.din(w_dff_A_pDtEMtL68_1),.clk(gclk));
	jdff dff_A_O7Jo6SXl6_1(.dout(w_dff_A_pDtEMtL68_1),.din(w_dff_A_O7Jo6SXl6_1),.clk(gclk));
	jdff dff_A_3wySArqs6_1(.dout(w_dff_A_O7Jo6SXl6_1),.din(w_dff_A_3wySArqs6_1),.clk(gclk));
	jdff dff_A_NYHHFhxm7_1(.dout(w_dff_A_3wySArqs6_1),.din(w_dff_A_NYHHFhxm7_1),.clk(gclk));
	jdff dff_A_KayMGbHT1_1(.dout(w_dff_A_NYHHFhxm7_1),.din(w_dff_A_KayMGbHT1_1),.clk(gclk));
	jdff dff_A_lLFT9WMi5_1(.dout(w_dff_A_KayMGbHT1_1),.din(w_dff_A_lLFT9WMi5_1),.clk(gclk));
	jdff dff_A_wKof2ftZ0_1(.dout(w_dff_A_lLFT9WMi5_1),.din(w_dff_A_wKof2ftZ0_1),.clk(gclk));
	jdff dff_A_Zpy5zA207_1(.dout(w_dff_A_wKof2ftZ0_1),.din(w_dff_A_Zpy5zA207_1),.clk(gclk));
	jdff dff_A_ym1Eibhz7_1(.dout(w_dff_A_Zpy5zA207_1),.din(w_dff_A_ym1Eibhz7_1),.clk(gclk));
	jdff dff_B_lULSSn2v6_1(.din(n601),.dout(w_dff_B_lULSSn2v6_1),.clk(gclk));
	jdff dff_B_0p2ojq8i8_0(.din(G130),.dout(w_dff_B_0p2ojq8i8_0),.clk(gclk));
	jdff dff_A_SsXq4vV18_2(.dout(w_G3729_0[2]),.din(w_dff_A_SsXq4vV18_2),.clk(gclk));
	jdff dff_A_fzEbCmmv1_2(.dout(w_dff_A_SsXq4vV18_2),.din(w_dff_A_fzEbCmmv1_2),.clk(gclk));
	jdff dff_A_Myy3nlgI8_2(.dout(w_dff_A_fzEbCmmv1_2),.din(w_dff_A_Myy3nlgI8_2),.clk(gclk));
	jdff dff_A_Uq2Gp1T96_2(.dout(w_dff_A_Myy3nlgI8_2),.din(w_dff_A_Uq2Gp1T96_2),.clk(gclk));
	jdff dff_A_IcAFC0mS5_1(.dout(w_n1105_0[1]),.din(w_dff_A_IcAFC0mS5_1),.clk(gclk));
	jdff dff_A_EZ39tuNI9_1(.dout(w_dff_A_IcAFC0mS5_1),.din(w_dff_A_EZ39tuNI9_1),.clk(gclk));
	jdff dff_A_OCosiyvZ4_1(.dout(w_dff_A_EZ39tuNI9_1),.din(w_dff_A_OCosiyvZ4_1),.clk(gclk));
	jdff dff_A_BUTLgfjH3_1(.dout(w_dff_A_OCosiyvZ4_1),.din(w_dff_A_BUTLgfjH3_1),.clk(gclk));
	jdff dff_A_AP5bIcxU3_1(.dout(w_dff_A_BUTLgfjH3_1),.din(w_dff_A_AP5bIcxU3_1),.clk(gclk));
	jdff dff_A_FtDVlJMR1_1(.dout(w_dff_A_AP5bIcxU3_1),.din(w_dff_A_FtDVlJMR1_1),.clk(gclk));
	jdff dff_A_CqddQdSg5_1(.dout(w_dff_A_FtDVlJMR1_1),.din(w_dff_A_CqddQdSg5_1),.clk(gclk));
	jdff dff_A_JN1pSXGJ2_1(.dout(w_dff_A_CqddQdSg5_1),.din(w_dff_A_JN1pSXGJ2_1),.clk(gclk));
	jdff dff_A_kCk5ZQvw1_1(.dout(w_dff_A_JN1pSXGJ2_1),.din(w_dff_A_kCk5ZQvw1_1),.clk(gclk));
	jdff dff_A_eNTiblVA7_1(.dout(w_dff_A_kCk5ZQvw1_1),.din(w_dff_A_eNTiblVA7_1),.clk(gclk));
	jdff dff_B_dqPP4jvQ7_2(.din(n1105),.dout(w_dff_B_dqPP4jvQ7_2),.clk(gclk));
	jdff dff_B_XueDhB7k7_1(.din(n596),.dout(w_dff_B_XueDhB7k7_1),.clk(gclk));
	jdff dff_B_XAFmI2px1_0(.din(G127),.dout(w_dff_B_XAFmI2px1_0),.clk(gclk));
	jdff dff_A_G4DRRie31_1(.dout(w_n595_0[1]),.din(w_dff_A_G4DRRie31_1),.clk(gclk));
	jdff dff_A_hKABPv192_1(.dout(w_dff_A_G4DRRie31_1),.din(w_dff_A_hKABPv192_1),.clk(gclk));
	jdff dff_A_SqMPRcZC1_2(.dout(w_n595_0[2]),.din(w_dff_A_SqMPRcZC1_2),.clk(gclk));
	jdff dff_A_OtRZhWkL0_2(.dout(w_dff_A_SqMPRcZC1_2),.din(w_dff_A_OtRZhWkL0_2),.clk(gclk));
	jdff dff_A_BuLXbkO42_1(.dout(w_G3737_0[1]),.din(w_dff_A_BuLXbkO42_1),.clk(gclk));
	jdff dff_A_7NPCYtjt2_1(.dout(w_dff_A_BuLXbkO42_1),.din(w_dff_A_7NPCYtjt2_1),.clk(gclk));
	jdff dff_A_cHu6eCAS9_1(.dout(w_dff_A_7NPCYtjt2_1),.din(w_dff_A_cHu6eCAS9_1),.clk(gclk));
	jdff dff_A_wq8328gB9_1(.dout(w_dff_A_cHu6eCAS9_1),.din(w_dff_A_wq8328gB9_1),.clk(gclk));
	jdff dff_B_LtWNy6fy1_1(.din(n1087),.dout(w_dff_B_LtWNy6fy1_1),.clk(gclk));
	jdff dff_B_rO78xemd1_1(.din(w_dff_B_LtWNy6fy1_1),.dout(w_dff_B_rO78xemd1_1),.clk(gclk));
	jdff dff_B_QrSECUrD8_1(.din(w_dff_B_rO78xemd1_1),.dout(w_dff_B_QrSECUrD8_1),.clk(gclk));
	jdff dff_B_t2W9AHbf2_1(.din(w_dff_B_QrSECUrD8_1),.dout(w_dff_B_t2W9AHbf2_1),.clk(gclk));
	jdff dff_B_xEOXWKi15_1(.din(w_dff_B_t2W9AHbf2_1),.dout(w_dff_B_xEOXWKi15_1),.clk(gclk));
	jdff dff_B_bqNfjuoh2_1(.din(w_dff_B_xEOXWKi15_1),.dout(w_dff_B_bqNfjuoh2_1),.clk(gclk));
	jdff dff_B_iuGSE1wl9_1(.din(n1088),.dout(w_dff_B_iuGSE1wl9_1),.clk(gclk));
	jdff dff_B_bxk3BgJ65_1(.din(w_dff_B_iuGSE1wl9_1),.dout(w_dff_B_bxk3BgJ65_1),.clk(gclk));
	jdff dff_B_45VyFlQB5_1(.din(w_dff_B_bxk3BgJ65_1),.dout(w_dff_B_45VyFlQB5_1),.clk(gclk));
	jdff dff_B_ZdHS22Za8_1(.din(n1062),.dout(w_dff_B_ZdHS22Za8_1),.clk(gclk));
	jdff dff_B_Tjb98FfF9_1(.din(w_dff_B_ZdHS22Za8_1),.dout(w_dff_B_Tjb98FfF9_1),.clk(gclk));
	jdff dff_B_8t3jpyCn9_1(.din(n1063),.dout(w_dff_B_8t3jpyCn9_1),.clk(gclk));
	jdff dff_B_q4V9eCAW1_1(.din(n1064),.dout(w_dff_B_q4V9eCAW1_1),.clk(gclk));
	jdff dff_A_cysCXh4O1_1(.dout(w_n656_0[1]),.din(w_dff_A_cysCXh4O1_1),.clk(gclk));
	jdff dff_A_bU3HxgH34_1(.dout(w_dff_A_cysCXh4O1_1),.din(w_dff_A_bU3HxgH34_1),.clk(gclk));
	jdff dff_A_FTVzuvmY1_1(.dout(w_n655_0[1]),.din(w_dff_A_FTVzuvmY1_1),.clk(gclk));
	jdff dff_A_Ynu68b1n4_1(.dout(w_dff_A_FTVzuvmY1_1),.din(w_dff_A_Ynu68b1n4_1),.clk(gclk));
	jdff dff_A_PDijplF23_1(.dout(w_dff_A_Ynu68b1n4_1),.din(w_dff_A_PDijplF23_1),.clk(gclk));
	jdff dff_A_OGbbccXe7_1(.dout(w_n654_0[1]),.din(w_dff_A_OGbbccXe7_1),.clk(gclk));
	jdff dff_A_FuBjQKpz4_1(.dout(w_dff_A_OGbbccXe7_1),.din(w_dff_A_FuBjQKpz4_1),.clk(gclk));
	jdff dff_A_reYAtjlZ6_1(.dout(w_dff_A_FuBjQKpz4_1),.din(w_dff_A_reYAtjlZ6_1),.clk(gclk));
	jdff dff_A_6P3ypGPy3_1(.dout(w_dff_A_reYAtjlZ6_1),.din(w_dff_A_6P3ypGPy3_1),.clk(gclk));
	jdff dff_A_NUufaEzV0_1(.dout(w_dff_A_6P3ypGPy3_1),.din(w_dff_A_NUufaEzV0_1),.clk(gclk));
	jdff dff_A_2vpKgsog9_1(.dout(w_dff_A_NUufaEzV0_1),.din(w_dff_A_2vpKgsog9_1),.clk(gclk));
	jdff dff_A_ce8Cg8FA8_1(.dout(w_dff_A_2vpKgsog9_1),.din(w_dff_A_ce8Cg8FA8_1),.clk(gclk));
	jdff dff_A_qPcqFAnM7_2(.dout(w_n654_0[2]),.din(w_dff_A_qPcqFAnM7_2),.clk(gclk));
	jdff dff_A_b96WBDRe8_2(.dout(w_dff_A_qPcqFAnM7_2),.din(w_dff_A_b96WBDRe8_2),.clk(gclk));
	jdff dff_A_JmNaSGB24_2(.dout(w_dff_A_b96WBDRe8_2),.din(w_dff_A_JmNaSGB24_2),.clk(gclk));
	jdff dff_A_zA6O4Agt9_2(.dout(w_dff_A_JmNaSGB24_2),.din(w_dff_A_zA6O4Agt9_2),.clk(gclk));
	jdff dff_A_XI4CKZxJ1_0(.dout(w_n652_0[0]),.din(w_dff_A_XI4CKZxJ1_0),.clk(gclk));
	jdff dff_A_kG63O8gK8_0(.dout(w_dff_A_XI4CKZxJ1_0),.din(w_dff_A_kG63O8gK8_0),.clk(gclk));
	jdff dff_A_hkHSszR17_0(.dout(w_dff_A_kG63O8gK8_0),.din(w_dff_A_hkHSszR17_0),.clk(gclk));
	jdff dff_A_nJFI4ewU7_0(.dout(w_dff_A_hkHSszR17_0),.din(w_dff_A_nJFI4ewU7_0),.clk(gclk));
	jdff dff_A_tgb0i89Y2_0(.dout(w_n649_0[0]),.din(w_dff_A_tgb0i89Y2_0),.clk(gclk));
	jdff dff_A_0e2A0Xbb2_0(.dout(w_dff_A_tgb0i89Y2_0),.din(w_dff_A_0e2A0Xbb2_0),.clk(gclk));
	jdff dff_A_vjFv8mU73_0(.dout(w_dff_A_0e2A0Xbb2_0),.din(w_dff_A_vjFv8mU73_0),.clk(gclk));
	jdff dff_A_wcqp9dnb6_0(.dout(w_dff_A_vjFv8mU73_0),.din(w_dff_A_wcqp9dnb6_0),.clk(gclk));
	jdff dff_A_9aQUFTwP0_0(.dout(w_dff_A_wcqp9dnb6_0),.din(w_dff_A_9aQUFTwP0_0),.clk(gclk));
	jdff dff_A_9fFv3bbF7_1(.dout(w_n647_0[1]),.din(w_dff_A_9fFv3bbF7_1),.clk(gclk));
	jdff dff_A_ryOVwv122_1(.dout(w_dff_A_9fFv3bbF7_1),.din(w_dff_A_ryOVwv122_1),.clk(gclk));
	jdff dff_A_uuO3hIu62_1(.dout(w_dff_A_ryOVwv122_1),.din(w_dff_A_uuO3hIu62_1),.clk(gclk));
	jdff dff_A_lAilQdBT7_1(.dout(w_dff_A_uuO3hIu62_1),.din(w_dff_A_lAilQdBT7_1),.clk(gclk));
	jdff dff_A_igMw3oUG4_1(.dout(w_dff_A_lAilQdBT7_1),.din(w_dff_A_igMw3oUG4_1),.clk(gclk));
	jdff dff_A_LWSNA2DT0_1(.dout(w_dff_A_igMw3oUG4_1),.din(w_dff_A_LWSNA2DT0_1),.clk(gclk));
	jdff dff_A_wGTAaL9u6_1(.dout(w_dff_A_LWSNA2DT0_1),.din(w_dff_A_wGTAaL9u6_1),.clk(gclk));
	jdff dff_A_5np9xzlW8_0(.dout(w_n1086_0[0]),.din(w_dff_A_5np9xzlW8_0),.clk(gclk));
	jdff dff_B_ddE4oc3f2_2(.din(n1086),.dout(w_dff_B_ddE4oc3f2_2),.clk(gclk));
	jdff dff_B_IrzrFxNw3_2(.din(w_dff_B_ddE4oc3f2_2),.dout(w_dff_B_IrzrFxNw3_2),.clk(gclk));
	jdff dff_A_I66KZtkK6_1(.dout(w_n646_0[1]),.din(w_dff_A_I66KZtkK6_1),.clk(gclk));
	jdff dff_A_vpPwzcMV9_1(.dout(w_dff_A_I66KZtkK6_1),.din(w_dff_A_vpPwzcMV9_1),.clk(gclk));
	jdff dff_A_Xub83BwO5_1(.dout(w_dff_A_vpPwzcMV9_1),.din(w_dff_A_Xub83BwO5_1),.clk(gclk));
	jdff dff_A_Q4gslOok1_1(.dout(w_n642_0[1]),.din(w_dff_A_Q4gslOok1_1),.clk(gclk));
	jdff dff_A_VjQZaMGs4_1(.dout(w_dff_A_Q4gslOok1_1),.din(w_dff_A_VjQZaMGs4_1),.clk(gclk));
	jdff dff_B_NUMZYu669_3(.din(n642),.dout(w_dff_B_NUMZYu669_3),.clk(gclk));
	jdff dff_A_tj16hwk92_0(.dout(w_G29_0[0]),.din(w_dff_A_tj16hwk92_0),.clk(gclk));
	jdff dff_A_3SL7naHL2_0(.dout(w_G3705_1[0]),.din(w_dff_A_3SL7naHL2_0),.clk(gclk));
	jdff dff_A_L4pp5dTu2_0(.dout(w_dff_A_3SL7naHL2_0),.din(w_dff_A_L4pp5dTu2_0),.clk(gclk));
	jdff dff_A_4z0juuWj9_0(.dout(w_dff_A_L4pp5dTu2_0),.din(w_dff_A_4z0juuWj9_0),.clk(gclk));
	jdff dff_A_eorgmWoP0_2(.dout(w_G3705_1[2]),.din(w_dff_A_eorgmWoP0_2),.clk(gclk));
	jdff dff_A_EIYJuf6S6_2(.dout(w_dff_A_eorgmWoP0_2),.din(w_dff_A_EIYJuf6S6_2),.clk(gclk));
	jdff dff_A_YPFFoyh43_2(.dout(w_dff_A_EIYJuf6S6_2),.din(w_dff_A_YPFFoyh43_2),.clk(gclk));
	jdff dff_A_V0MKqD0R2_2(.dout(w_G3705_0[2]),.din(w_dff_A_V0MKqD0R2_2),.clk(gclk));
	jdff dff_A_zSq0MprW8_2(.dout(w_dff_A_V0MKqD0R2_2),.din(w_dff_A_zSq0MprW8_2),.clk(gclk));
	jdff dff_A_w8ug4njh8_2(.dout(w_dff_A_zSq0MprW8_2),.din(w_dff_A_w8ug4njh8_2),.clk(gclk));
	jdff dff_A_8QWeCkZB8_0(.dout(w_n357_0[0]),.din(w_dff_A_8QWeCkZB8_0),.clk(gclk));
	jdff dff_A_qoaZTQKb9_0(.dout(w_dff_A_8QWeCkZB8_0),.din(w_dff_A_qoaZTQKb9_0),.clk(gclk));
	jdff dff_A_8u8zz0hI7_0(.dout(w_dff_A_qoaZTQKb9_0),.din(w_dff_A_8u8zz0hI7_0),.clk(gclk));
	jdff dff_B_bRLAOsI35_3(.din(n354),.dout(w_dff_B_bRLAOsI35_3),.clk(gclk));
	jdff dff_A_ox4zSsWX7_0(.dout(w_G41_0[0]),.din(w_dff_A_ox4zSsWX7_0),.clk(gclk));
	jdff dff_A_8S7dEa0i4_1(.dout(w_G3701_1[1]),.din(w_dff_A_8S7dEa0i4_1),.clk(gclk));
	jdff dff_A_Pqsjnv4v5_0(.dout(w_G3701_0[0]),.din(w_dff_A_Pqsjnv4v5_0),.clk(gclk));
	jdff dff_A_xcezbmkX0_1(.dout(w_n636_0[1]),.din(w_dff_A_xcezbmkX0_1),.clk(gclk));
	jdff dff_A_ueHqDwNa9_1(.dout(w_dff_A_xcezbmkX0_1),.din(w_dff_A_ueHqDwNa9_1),.clk(gclk));
	jdff dff_A_J7rztvn01_1(.dout(w_dff_A_ueHqDwNa9_1),.din(w_dff_A_J7rztvn01_1),.clk(gclk));
	jdff dff_A_gg61SxAS4_1(.dout(w_dff_A_J7rztvn01_1),.din(w_dff_A_gg61SxAS4_1),.clk(gclk));
	jdff dff_A_ZKNFV40b0_2(.dout(w_n636_0[2]),.din(w_dff_A_ZKNFV40b0_2),.clk(gclk));
	jdff dff_A_fEUrzPyw6_2(.dout(w_dff_A_ZKNFV40b0_2),.din(w_dff_A_fEUrzPyw6_2),.clk(gclk));
	jdff dff_B_C6xg2Z3Z4_1(.din(n633),.dout(w_dff_B_C6xg2Z3Z4_1),.clk(gclk));
	jdff dff_B_imc1wVcA6_0(.din(G26),.dout(w_dff_B_imc1wVcA6_0),.clk(gclk));
	jdff dff_A_h8yjWpDz5_1(.dout(w_G18_42[1]),.din(w_dff_A_h8yjWpDz5_1),.clk(gclk));
	jdff dff_A_xz0LDdqJ7_0(.dout(w_n632_0[0]),.din(w_dff_A_xz0LDdqJ7_0),.clk(gclk));
	jdff dff_A_oKX0JHAy5_0(.dout(w_dff_A_xz0LDdqJ7_0),.din(w_dff_A_oKX0JHAy5_0),.clk(gclk));
	jdff dff_A_CKSZqIIO0_2(.dout(w_n632_0[2]),.din(w_dff_A_CKSZqIIO0_2),.clk(gclk));
	jdff dff_A_nAx8PBdD7_2(.dout(w_dff_A_CKSZqIIO0_2),.din(w_dff_A_nAx8PBdD7_2),.clk(gclk));
	jdff dff_A_EtjwFWbC2_1(.dout(w_n631_0[1]),.din(w_dff_A_EtjwFWbC2_1),.clk(gclk));
	jdff dff_A_xJI09LtI7_1(.dout(w_dff_A_EtjwFWbC2_1),.din(w_dff_A_xJI09LtI7_1),.clk(gclk));
	jdff dff_A_DkSJbuj46_1(.dout(w_dff_A_xJI09LtI7_1),.din(w_dff_A_DkSJbuj46_1),.clk(gclk));
	jdff dff_A_J8W2vvAm2_1(.dout(w_dff_A_DkSJbuj46_1),.din(w_dff_A_J8W2vvAm2_1),.clk(gclk));
	jdff dff_A_9Y44Fhkp4_1(.dout(w_dff_A_J8W2vvAm2_1),.din(w_dff_A_9Y44Fhkp4_1),.clk(gclk));
	jdff dff_A_EXP6f9nN5_1(.dout(w_dff_A_9Y44Fhkp4_1),.din(w_dff_A_EXP6f9nN5_1),.clk(gclk));
	jdff dff_A_tikeZxdx1_1(.dout(w_dff_A_EXP6f9nN5_1),.din(w_dff_A_tikeZxdx1_1),.clk(gclk));
	jdff dff_A_WtEFTgVK8_2(.dout(w_n631_0[2]),.din(w_dff_A_WtEFTgVK8_2),.clk(gclk));
	jdff dff_A_6fV3kaxC7_2(.dout(w_dff_A_WtEFTgVK8_2),.din(w_dff_A_6fV3kaxC7_2),.clk(gclk));
	jdff dff_A_FSv2gqVb9_2(.dout(w_dff_A_6fV3kaxC7_2),.din(w_dff_A_FSv2gqVb9_2),.clk(gclk));
	jdff dff_B_eSI8rUsk5_1(.din(n628),.dout(w_dff_B_eSI8rUsk5_1),.clk(gclk));
	jdff dff_B_qWV7iYu50_0(.din(G23),.dout(w_dff_B_qWV7iYu50_0),.clk(gclk));
	jdff dff_A_9I9RuQo60_1(.dout(w_n627_0[1]),.din(w_dff_A_9I9RuQo60_1),.clk(gclk));
	jdff dff_A_imEWMNjW5_1(.dout(w_dff_A_9I9RuQo60_1),.din(w_dff_A_imEWMNjW5_1),.clk(gclk));
	jdff dff_A_lZJY7RlZ8_2(.dout(w_n627_0[2]),.din(w_dff_A_lZJY7RlZ8_2),.clk(gclk));
	jdff dff_A_woTKomL55_2(.dout(w_dff_A_lZJY7RlZ8_2),.din(w_dff_A_woTKomL55_2),.clk(gclk));
	jdff dff_A_1G0kWD285_1(.dout(w_G3717_0[1]),.din(w_dff_A_1G0kWD285_1),.clk(gclk));
	jdff dff_A_hyOa1aWo8_1(.dout(w_dff_A_1G0kWD285_1),.din(w_dff_A_hyOa1aWo8_1),.clk(gclk));
	jdff dff_A_PNL2GcxS9_1(.dout(w_dff_A_hyOa1aWo8_1),.din(w_dff_A_PNL2GcxS9_1),.clk(gclk));
	jdff dff_A_x0EMkzxd8_1(.dout(w_dff_A_PNL2GcxS9_1),.din(w_dff_A_x0EMkzxd8_1),.clk(gclk));
	jdff dff_A_jObMJrur8_0(.dout(w_n626_1[0]),.din(w_dff_A_jObMJrur8_0),.clk(gclk));
	jdff dff_A_mKzlczDt4_0(.dout(w_dff_A_jObMJrur8_0),.din(w_dff_A_mKzlczDt4_0),.clk(gclk));
	jdff dff_A_KtpsS1Dp0_0(.dout(w_dff_A_mKzlczDt4_0),.din(w_dff_A_KtpsS1Dp0_0),.clk(gclk));
	jdff dff_A_KEHmf4lu0_0(.dout(w_dff_A_KtpsS1Dp0_0),.din(w_dff_A_KEHmf4lu0_0),.clk(gclk));
	jdff dff_A_Gs5W5Cso5_0(.dout(w_dff_A_KEHmf4lu0_0),.din(w_dff_A_Gs5W5Cso5_0),.clk(gclk));
	jdff dff_A_ZBMCsjP81_0(.dout(w_n626_0[0]),.din(w_dff_A_ZBMCsjP81_0),.clk(gclk));
	jdff dff_A_DhWvulUT0_0(.dout(w_dff_A_ZBMCsjP81_0),.din(w_dff_A_DhWvulUT0_0),.clk(gclk));
	jdff dff_A_iimobAsk6_0(.dout(w_dff_A_DhWvulUT0_0),.din(w_dff_A_iimobAsk6_0),.clk(gclk));
	jdff dff_A_3kVY6l0E9_0(.dout(w_dff_A_iimobAsk6_0),.din(w_dff_A_3kVY6l0E9_0),.clk(gclk));
	jdff dff_A_XNShdIJK8_1(.dout(w_n626_0[1]),.din(w_dff_A_XNShdIJK8_1),.clk(gclk));
	jdff dff_A_haP4sgFU1_1(.dout(w_dff_A_XNShdIJK8_1),.din(w_dff_A_haP4sgFU1_1),.clk(gclk));
	jdff dff_A_Qcljl5nJ4_1(.dout(w_dff_A_haP4sgFU1_1),.din(w_dff_A_Qcljl5nJ4_1),.clk(gclk));
	jdff dff_A_wND6vBd05_1(.dout(w_dff_A_Qcljl5nJ4_1),.din(w_dff_A_wND6vBd05_1),.clk(gclk));
	jdff dff_B_A084MN4E7_1(.din(n623),.dout(w_dff_B_A084MN4E7_1),.clk(gclk));
	jdff dff_B_uNyvENmp2_0(.din(G103),.dout(w_dff_B_uNyvENmp2_0),.clk(gclk));
	jdff dff_A_sd1wNqVa8_2(.dout(w_G18_49[2]),.din(w_dff_A_sd1wNqVa8_2),.clk(gclk));
	jdff dff_A_QttmMOPF5_1(.dout(w_n622_0[1]),.din(w_dff_A_QttmMOPF5_1),.clk(gclk));
	jdff dff_A_Ovq9bdPh2_1(.dout(w_dff_A_QttmMOPF5_1),.din(w_dff_A_Ovq9bdPh2_1),.clk(gclk));
	jdff dff_A_zoLh1nev8_2(.dout(w_n622_0[2]),.din(w_dff_A_zoLh1nev8_2),.clk(gclk));
	jdff dff_A_erNsfYQU8_2(.dout(w_dff_A_zoLh1nev8_2),.din(w_dff_A_erNsfYQU8_2),.clk(gclk));
	jdff dff_A_nAynoQZb3_1(.dout(w_G3723_0[1]),.din(w_dff_A_nAynoQZb3_1),.clk(gclk));
	jdff dff_A_8rwikamZ4_1(.dout(w_dff_A_nAynoQZb3_1),.din(w_dff_A_8rwikamZ4_1),.clk(gclk));
	jdff dff_A_OQjVDZsr1_1(.dout(w_dff_A_8rwikamZ4_1),.din(w_dff_A_OQjVDZsr1_1),.clk(gclk));
	jdff dff_A_RgggCuSl6_1(.dout(w_dff_A_OQjVDZsr1_1),.din(w_dff_A_RgggCuSl6_1),.clk(gclk));
	jdff dff_A_StDwqhMe5_1(.dout(w_dff_A_SeHU1hgo8_0),.din(w_dff_A_StDwqhMe5_1),.clk(gclk));
	jdff dff_A_SeHU1hgo8_0(.dout(w_dff_A_T3vqXCwM2_0),.din(w_dff_A_SeHU1hgo8_0),.clk(gclk));
	jdff dff_A_T3vqXCwM2_0(.dout(w_dff_A_KoxgZOEF1_0),.din(w_dff_A_T3vqXCwM2_0),.clk(gclk));
	jdff dff_A_KoxgZOEF1_0(.dout(w_dff_A_bWecyCwf2_0),.din(w_dff_A_KoxgZOEF1_0),.clk(gclk));
	jdff dff_A_bWecyCwf2_0(.dout(w_dff_A_AzJeX3xC8_0),.din(w_dff_A_bWecyCwf2_0),.clk(gclk));
	jdff dff_A_AzJeX3xC8_0(.dout(w_dff_A_sL5HqlXH6_0),.din(w_dff_A_AzJeX3xC8_0),.clk(gclk));
	jdff dff_A_sL5HqlXH6_0(.dout(w_dff_A_jEGO6G9f3_0),.din(w_dff_A_sL5HqlXH6_0),.clk(gclk));
	jdff dff_A_jEGO6G9f3_0(.dout(w_dff_A_ol50RqS85_0),.din(w_dff_A_jEGO6G9f3_0),.clk(gclk));
	jdff dff_A_ol50RqS85_0(.dout(w_dff_A_V7E4IWB67_0),.din(w_dff_A_ol50RqS85_0),.clk(gclk));
	jdff dff_A_V7E4IWB67_0(.dout(w_dff_A_WAdk7IEB6_0),.din(w_dff_A_V7E4IWB67_0),.clk(gclk));
	jdff dff_A_WAdk7IEB6_0(.dout(w_dff_A_VOrFJZH17_0),.din(w_dff_A_WAdk7IEB6_0),.clk(gclk));
	jdff dff_A_VOrFJZH17_0(.dout(w_dff_A_2mO9BGRa1_0),.din(w_dff_A_VOrFJZH17_0),.clk(gclk));
	jdff dff_A_2mO9BGRa1_0(.dout(w_dff_A_7MkaPO6t1_0),.din(w_dff_A_2mO9BGRa1_0),.clk(gclk));
	jdff dff_A_7MkaPO6t1_0(.dout(w_dff_A_yGAzjzMr3_0),.din(w_dff_A_7MkaPO6t1_0),.clk(gclk));
	jdff dff_A_yGAzjzMr3_0(.dout(w_dff_A_QldLZweh7_0),.din(w_dff_A_yGAzjzMr3_0),.clk(gclk));
	jdff dff_A_QldLZweh7_0(.dout(w_dff_A_LRwXOCGr6_0),.din(w_dff_A_QldLZweh7_0),.clk(gclk));
	jdff dff_A_LRwXOCGr6_0(.dout(w_dff_A_cUxzD6Z81_0),.din(w_dff_A_LRwXOCGr6_0),.clk(gclk));
	jdff dff_A_cUxzD6Z81_0(.dout(w_dff_A_w1EMWtID4_0),.din(w_dff_A_cUxzD6Z81_0),.clk(gclk));
	jdff dff_A_w1EMWtID4_0(.dout(w_dff_A_ICd6E9qD0_0),.din(w_dff_A_w1EMWtID4_0),.clk(gclk));
	jdff dff_A_ICd6E9qD0_0(.dout(w_dff_A_Iewlz38u3_0),.din(w_dff_A_ICd6E9qD0_0),.clk(gclk));
	jdff dff_A_Iewlz38u3_0(.dout(w_dff_A_UpIfp7D50_0),.din(w_dff_A_Iewlz38u3_0),.clk(gclk));
	jdff dff_A_UpIfp7D50_0(.dout(w_dff_A_TTQnkFMr2_0),.din(w_dff_A_UpIfp7D50_0),.clk(gclk));
	jdff dff_A_TTQnkFMr2_0(.dout(w_dff_A_u2fcHUyK2_0),.din(w_dff_A_TTQnkFMr2_0),.clk(gclk));
	jdff dff_A_u2fcHUyK2_0(.dout(w_dff_A_KLwZPYX23_0),.din(w_dff_A_u2fcHUyK2_0),.clk(gclk));
	jdff dff_A_KLwZPYX23_0(.dout(w_dff_A_YP5NO6vp6_0),.din(w_dff_A_KLwZPYX23_0),.clk(gclk));
	jdff dff_A_YP5NO6vp6_0(.dout(w_dff_A_gV3La4kk8_0),.din(w_dff_A_YP5NO6vp6_0),.clk(gclk));
	jdff dff_A_gV3La4kk8_0(.dout(w_dff_A_eB55MZVj0_0),.din(w_dff_A_gV3La4kk8_0),.clk(gclk));
	jdff dff_A_eB55MZVj0_0(.dout(w_dff_A_hKEjw8si9_0),.din(w_dff_A_eB55MZVj0_0),.clk(gclk));
	jdff dff_A_hKEjw8si9_0(.dout(w_dff_A_TGt4jsAn4_0),.din(w_dff_A_hKEjw8si9_0),.clk(gclk));
	jdff dff_A_TGt4jsAn4_0(.dout(w_dff_A_fe7BH65t8_0),.din(w_dff_A_TGt4jsAn4_0),.clk(gclk));
	jdff dff_A_fe7BH65t8_0(.dout(w_dff_A_NxO8nnaY3_0),.din(w_dff_A_fe7BH65t8_0),.clk(gclk));
	jdff dff_A_NxO8nnaY3_0(.dout(w_dff_A_zwJRnC6v8_0),.din(w_dff_A_NxO8nnaY3_0),.clk(gclk));
	jdff dff_A_zwJRnC6v8_0(.dout(w_dff_A_5W9wWePd1_0),.din(w_dff_A_zwJRnC6v8_0),.clk(gclk));
	jdff dff_A_5W9wWePd1_0(.dout(w_dff_A_WjqOJxsZ7_0),.din(w_dff_A_5W9wWePd1_0),.clk(gclk));
	jdff dff_A_WjqOJxsZ7_0(.dout(w_dff_A_7qk2mgLd2_0),.din(w_dff_A_WjqOJxsZ7_0),.clk(gclk));
	jdff dff_A_7qk2mgLd2_0(.dout(w_dff_A_KhKWKH7s8_0),.din(w_dff_A_7qk2mgLd2_0),.clk(gclk));
	jdff dff_A_KhKWKH7s8_0(.dout(w_dff_A_3r7eKSVv3_0),.din(w_dff_A_KhKWKH7s8_0),.clk(gclk));
	jdff dff_A_3r7eKSVv3_0(.dout(G2),.din(w_dff_A_3r7eKSVv3_0),.clk(gclk));
	jdff dff_A_lnaQpt5X0_1(.dout(w_dff_A_akETpjd88_0),.din(w_dff_A_lnaQpt5X0_1),.clk(gclk));
	jdff dff_A_akETpjd88_0(.dout(w_dff_A_BRWlUsTg0_0),.din(w_dff_A_akETpjd88_0),.clk(gclk));
	jdff dff_A_BRWlUsTg0_0(.dout(w_dff_A_jbhnCSo23_0),.din(w_dff_A_BRWlUsTg0_0),.clk(gclk));
	jdff dff_A_jbhnCSo23_0(.dout(w_dff_A_CvAgXfbh8_0),.din(w_dff_A_jbhnCSo23_0),.clk(gclk));
	jdff dff_A_CvAgXfbh8_0(.dout(w_dff_A_JOO9heH96_0),.din(w_dff_A_CvAgXfbh8_0),.clk(gclk));
	jdff dff_A_JOO9heH96_0(.dout(w_dff_A_cb9wsTnb1_0),.din(w_dff_A_JOO9heH96_0),.clk(gclk));
	jdff dff_A_cb9wsTnb1_0(.dout(w_dff_A_H4a7cb6z9_0),.din(w_dff_A_cb9wsTnb1_0),.clk(gclk));
	jdff dff_A_H4a7cb6z9_0(.dout(w_dff_A_0h2NUQrw5_0),.din(w_dff_A_H4a7cb6z9_0),.clk(gclk));
	jdff dff_A_0h2NUQrw5_0(.dout(w_dff_A_Er9z4s6r0_0),.din(w_dff_A_0h2NUQrw5_0),.clk(gclk));
	jdff dff_A_Er9z4s6r0_0(.dout(w_dff_A_nuuhhDUB4_0),.din(w_dff_A_Er9z4s6r0_0),.clk(gclk));
	jdff dff_A_nuuhhDUB4_0(.dout(w_dff_A_Y0tSrl9Y2_0),.din(w_dff_A_nuuhhDUB4_0),.clk(gclk));
	jdff dff_A_Y0tSrl9Y2_0(.dout(w_dff_A_c3mtIW6s2_0),.din(w_dff_A_Y0tSrl9Y2_0),.clk(gclk));
	jdff dff_A_c3mtIW6s2_0(.dout(w_dff_A_ZAyTBcY43_0),.din(w_dff_A_c3mtIW6s2_0),.clk(gclk));
	jdff dff_A_ZAyTBcY43_0(.dout(w_dff_A_Jb4htPzv0_0),.din(w_dff_A_ZAyTBcY43_0),.clk(gclk));
	jdff dff_A_Jb4htPzv0_0(.dout(w_dff_A_Kno6wHgd8_0),.din(w_dff_A_Jb4htPzv0_0),.clk(gclk));
	jdff dff_A_Kno6wHgd8_0(.dout(w_dff_A_asZ4ybZH5_0),.din(w_dff_A_Kno6wHgd8_0),.clk(gclk));
	jdff dff_A_asZ4ybZH5_0(.dout(w_dff_A_JcMTuyK20_0),.din(w_dff_A_asZ4ybZH5_0),.clk(gclk));
	jdff dff_A_JcMTuyK20_0(.dout(w_dff_A_E9klAfIO8_0),.din(w_dff_A_JcMTuyK20_0),.clk(gclk));
	jdff dff_A_E9klAfIO8_0(.dout(w_dff_A_aFhFIG2k8_0),.din(w_dff_A_E9klAfIO8_0),.clk(gclk));
	jdff dff_A_aFhFIG2k8_0(.dout(w_dff_A_pC5ZSHLp6_0),.din(w_dff_A_aFhFIG2k8_0),.clk(gclk));
	jdff dff_A_pC5ZSHLp6_0(.dout(w_dff_A_dcZZo00o8_0),.din(w_dff_A_pC5ZSHLp6_0),.clk(gclk));
	jdff dff_A_dcZZo00o8_0(.dout(w_dff_A_57l2aB2k0_0),.din(w_dff_A_dcZZo00o8_0),.clk(gclk));
	jdff dff_A_57l2aB2k0_0(.dout(w_dff_A_cZa7Y2LU5_0),.din(w_dff_A_57l2aB2k0_0),.clk(gclk));
	jdff dff_A_cZa7Y2LU5_0(.dout(w_dff_A_VtBhzFD22_0),.din(w_dff_A_cZa7Y2LU5_0),.clk(gclk));
	jdff dff_A_VtBhzFD22_0(.dout(w_dff_A_ZEnx1QJh6_0),.din(w_dff_A_VtBhzFD22_0),.clk(gclk));
	jdff dff_A_ZEnx1QJh6_0(.dout(w_dff_A_4lPC5YK68_0),.din(w_dff_A_ZEnx1QJh6_0),.clk(gclk));
	jdff dff_A_4lPC5YK68_0(.dout(w_dff_A_vR5xfdH05_0),.din(w_dff_A_4lPC5YK68_0),.clk(gclk));
	jdff dff_A_vR5xfdH05_0(.dout(w_dff_A_5pce0cdr3_0),.din(w_dff_A_vR5xfdH05_0),.clk(gclk));
	jdff dff_A_5pce0cdr3_0(.dout(w_dff_A_ULxU10nX0_0),.din(w_dff_A_5pce0cdr3_0),.clk(gclk));
	jdff dff_A_ULxU10nX0_0(.dout(w_dff_A_vRm0XJat8_0),.din(w_dff_A_ULxU10nX0_0),.clk(gclk));
	jdff dff_A_vRm0XJat8_0(.dout(w_dff_A_NoNuQYZl5_0),.din(w_dff_A_vRm0XJat8_0),.clk(gclk));
	jdff dff_A_NoNuQYZl5_0(.dout(w_dff_A_kqJI1BYN8_0),.din(w_dff_A_NoNuQYZl5_0),.clk(gclk));
	jdff dff_A_kqJI1BYN8_0(.dout(w_dff_A_33yiYwlA9_0),.din(w_dff_A_kqJI1BYN8_0),.clk(gclk));
	jdff dff_A_33yiYwlA9_0(.dout(w_dff_A_FetlggL45_0),.din(w_dff_A_33yiYwlA9_0),.clk(gclk));
	jdff dff_A_FetlggL45_0(.dout(w_dff_A_qErBFBCE0_0),.din(w_dff_A_FetlggL45_0),.clk(gclk));
	jdff dff_A_qErBFBCE0_0(.dout(w_dff_A_h2R4569f1_0),.din(w_dff_A_qErBFBCE0_0),.clk(gclk));
	jdff dff_A_h2R4569f1_0(.dout(w_dff_A_Ka7CPswc2_0),.din(w_dff_A_h2R4569f1_0),.clk(gclk));
	jdff dff_A_Ka7CPswc2_0(.dout(G3),.din(w_dff_A_Ka7CPswc2_0),.clk(gclk));
	jdff dff_A_nByzfYml7_1(.dout(w_dff_A_J2dNTYMk9_0),.din(w_dff_A_nByzfYml7_1),.clk(gclk));
	jdff dff_A_J2dNTYMk9_0(.dout(w_dff_A_JlQzPGxX6_0),.din(w_dff_A_J2dNTYMk9_0),.clk(gclk));
	jdff dff_A_JlQzPGxX6_0(.dout(w_dff_A_hNT8dqZ58_0),.din(w_dff_A_JlQzPGxX6_0),.clk(gclk));
	jdff dff_A_hNT8dqZ58_0(.dout(w_dff_A_RilbSa9c8_0),.din(w_dff_A_hNT8dqZ58_0),.clk(gclk));
	jdff dff_A_RilbSa9c8_0(.dout(w_dff_A_92Y45FwU6_0),.din(w_dff_A_RilbSa9c8_0),.clk(gclk));
	jdff dff_A_92Y45FwU6_0(.dout(w_dff_A_r1OWdJB38_0),.din(w_dff_A_92Y45FwU6_0),.clk(gclk));
	jdff dff_A_r1OWdJB38_0(.dout(w_dff_A_d3Oa4mE99_0),.din(w_dff_A_r1OWdJB38_0),.clk(gclk));
	jdff dff_A_d3Oa4mE99_0(.dout(w_dff_A_m8qSEMKx5_0),.din(w_dff_A_d3Oa4mE99_0),.clk(gclk));
	jdff dff_A_m8qSEMKx5_0(.dout(w_dff_A_Kol595Eo5_0),.din(w_dff_A_m8qSEMKx5_0),.clk(gclk));
	jdff dff_A_Kol595Eo5_0(.dout(w_dff_A_JTDHGrp79_0),.din(w_dff_A_Kol595Eo5_0),.clk(gclk));
	jdff dff_A_JTDHGrp79_0(.dout(w_dff_A_uwkSKMaW8_0),.din(w_dff_A_JTDHGrp79_0),.clk(gclk));
	jdff dff_A_uwkSKMaW8_0(.dout(w_dff_A_vfBdUksM7_0),.din(w_dff_A_uwkSKMaW8_0),.clk(gclk));
	jdff dff_A_vfBdUksM7_0(.dout(w_dff_A_02ugSumQ8_0),.din(w_dff_A_vfBdUksM7_0),.clk(gclk));
	jdff dff_A_02ugSumQ8_0(.dout(w_dff_A_7VOvqwFU2_0),.din(w_dff_A_02ugSumQ8_0),.clk(gclk));
	jdff dff_A_7VOvqwFU2_0(.dout(w_dff_A_ZBMacSA12_0),.din(w_dff_A_7VOvqwFU2_0),.clk(gclk));
	jdff dff_A_ZBMacSA12_0(.dout(w_dff_A_MugumP369_0),.din(w_dff_A_ZBMacSA12_0),.clk(gclk));
	jdff dff_A_MugumP369_0(.dout(w_dff_A_1giOurUF3_0),.din(w_dff_A_MugumP369_0),.clk(gclk));
	jdff dff_A_1giOurUF3_0(.dout(w_dff_A_cor92Twd7_0),.din(w_dff_A_1giOurUF3_0),.clk(gclk));
	jdff dff_A_cor92Twd7_0(.dout(w_dff_A_3AHtEvjq0_0),.din(w_dff_A_cor92Twd7_0),.clk(gclk));
	jdff dff_A_3AHtEvjq0_0(.dout(w_dff_A_oDe15tqa7_0),.din(w_dff_A_3AHtEvjq0_0),.clk(gclk));
	jdff dff_A_oDe15tqa7_0(.dout(w_dff_A_LzM80Iw81_0),.din(w_dff_A_oDe15tqa7_0),.clk(gclk));
	jdff dff_A_LzM80Iw81_0(.dout(w_dff_A_O3R5Eqsw7_0),.din(w_dff_A_LzM80Iw81_0),.clk(gclk));
	jdff dff_A_O3R5Eqsw7_0(.dout(w_dff_A_ax8DhLVl6_0),.din(w_dff_A_O3R5Eqsw7_0),.clk(gclk));
	jdff dff_A_ax8DhLVl6_0(.dout(w_dff_A_XmvNloMl0_0),.din(w_dff_A_ax8DhLVl6_0),.clk(gclk));
	jdff dff_A_XmvNloMl0_0(.dout(w_dff_A_v7bhiMPO1_0),.din(w_dff_A_XmvNloMl0_0),.clk(gclk));
	jdff dff_A_v7bhiMPO1_0(.dout(w_dff_A_b14A3KCN9_0),.din(w_dff_A_v7bhiMPO1_0),.clk(gclk));
	jdff dff_A_b14A3KCN9_0(.dout(w_dff_A_A8Uh0u299_0),.din(w_dff_A_b14A3KCN9_0),.clk(gclk));
	jdff dff_A_A8Uh0u299_0(.dout(w_dff_A_3vw78fWU2_0),.din(w_dff_A_A8Uh0u299_0),.clk(gclk));
	jdff dff_A_3vw78fWU2_0(.dout(w_dff_A_IVFV1qeD7_0),.din(w_dff_A_3vw78fWU2_0),.clk(gclk));
	jdff dff_A_IVFV1qeD7_0(.dout(w_dff_A_cDn6Vza06_0),.din(w_dff_A_IVFV1qeD7_0),.clk(gclk));
	jdff dff_A_cDn6Vza06_0(.dout(w_dff_A_U3Ur1uFB9_0),.din(w_dff_A_cDn6Vza06_0),.clk(gclk));
	jdff dff_A_U3Ur1uFB9_0(.dout(w_dff_A_gjmkPsRA6_0),.din(w_dff_A_U3Ur1uFB9_0),.clk(gclk));
	jdff dff_A_gjmkPsRA6_0(.dout(w_dff_A_bm8orVMl7_0),.din(w_dff_A_gjmkPsRA6_0),.clk(gclk));
	jdff dff_A_bm8orVMl7_0(.dout(w_dff_A_eTtD0IZL0_0),.din(w_dff_A_bm8orVMl7_0),.clk(gclk));
	jdff dff_A_eTtD0IZL0_0(.dout(w_dff_A_v33XOql27_0),.din(w_dff_A_eTtD0IZL0_0),.clk(gclk));
	jdff dff_A_v33XOql27_0(.dout(w_dff_A_mSnL3nEr0_0),.din(w_dff_A_v33XOql27_0),.clk(gclk));
	jdff dff_A_mSnL3nEr0_0(.dout(w_dff_A_PC9rFL5d2_0),.din(w_dff_A_mSnL3nEr0_0),.clk(gclk));
	jdff dff_A_PC9rFL5d2_0(.dout(G450),.din(w_dff_A_PC9rFL5d2_0),.clk(gclk));
	jdff dff_A_X1gH7vPc7_1(.dout(w_dff_A_ydkh7xRL8_0),.din(w_dff_A_X1gH7vPc7_1),.clk(gclk));
	jdff dff_A_ydkh7xRL8_0(.dout(w_dff_A_FCvaEbTU9_0),.din(w_dff_A_ydkh7xRL8_0),.clk(gclk));
	jdff dff_A_FCvaEbTU9_0(.dout(w_dff_A_yJcuvwvd0_0),.din(w_dff_A_FCvaEbTU9_0),.clk(gclk));
	jdff dff_A_yJcuvwvd0_0(.dout(w_dff_A_CLlJzujA7_0),.din(w_dff_A_yJcuvwvd0_0),.clk(gclk));
	jdff dff_A_CLlJzujA7_0(.dout(w_dff_A_25TzLaDL2_0),.din(w_dff_A_CLlJzujA7_0),.clk(gclk));
	jdff dff_A_25TzLaDL2_0(.dout(w_dff_A_GCGFgT1b1_0),.din(w_dff_A_25TzLaDL2_0),.clk(gclk));
	jdff dff_A_GCGFgT1b1_0(.dout(w_dff_A_svYKQF5g5_0),.din(w_dff_A_GCGFgT1b1_0),.clk(gclk));
	jdff dff_A_svYKQF5g5_0(.dout(w_dff_A_7bwT5q4B2_0),.din(w_dff_A_svYKQF5g5_0),.clk(gclk));
	jdff dff_A_7bwT5q4B2_0(.dout(w_dff_A_cfzUSbMH7_0),.din(w_dff_A_7bwT5q4B2_0),.clk(gclk));
	jdff dff_A_cfzUSbMH7_0(.dout(w_dff_A_zverzQER2_0),.din(w_dff_A_cfzUSbMH7_0),.clk(gclk));
	jdff dff_A_zverzQER2_0(.dout(w_dff_A_0N9Zz3165_0),.din(w_dff_A_zverzQER2_0),.clk(gclk));
	jdff dff_A_0N9Zz3165_0(.dout(w_dff_A_q3lNx0fH3_0),.din(w_dff_A_0N9Zz3165_0),.clk(gclk));
	jdff dff_A_q3lNx0fH3_0(.dout(w_dff_A_S9xkrVUq0_0),.din(w_dff_A_q3lNx0fH3_0),.clk(gclk));
	jdff dff_A_S9xkrVUq0_0(.dout(w_dff_A_KzOr32x21_0),.din(w_dff_A_S9xkrVUq0_0),.clk(gclk));
	jdff dff_A_KzOr32x21_0(.dout(w_dff_A_cbP674Kv9_0),.din(w_dff_A_KzOr32x21_0),.clk(gclk));
	jdff dff_A_cbP674Kv9_0(.dout(w_dff_A_atdhSgYQ0_0),.din(w_dff_A_cbP674Kv9_0),.clk(gclk));
	jdff dff_A_atdhSgYQ0_0(.dout(w_dff_A_XEooD6Y84_0),.din(w_dff_A_atdhSgYQ0_0),.clk(gclk));
	jdff dff_A_XEooD6Y84_0(.dout(w_dff_A_PMEDLE3F2_0),.din(w_dff_A_XEooD6Y84_0),.clk(gclk));
	jdff dff_A_PMEDLE3F2_0(.dout(w_dff_A_unq1obuO9_0),.din(w_dff_A_PMEDLE3F2_0),.clk(gclk));
	jdff dff_A_unq1obuO9_0(.dout(w_dff_A_9pChAC9s5_0),.din(w_dff_A_unq1obuO9_0),.clk(gclk));
	jdff dff_A_9pChAC9s5_0(.dout(w_dff_A_OxLpBcm77_0),.din(w_dff_A_9pChAC9s5_0),.clk(gclk));
	jdff dff_A_OxLpBcm77_0(.dout(w_dff_A_DNwDOW2w1_0),.din(w_dff_A_OxLpBcm77_0),.clk(gclk));
	jdff dff_A_DNwDOW2w1_0(.dout(w_dff_A_MmIfOmpd2_0),.din(w_dff_A_DNwDOW2w1_0),.clk(gclk));
	jdff dff_A_MmIfOmpd2_0(.dout(w_dff_A_UhhXUQQY4_0),.din(w_dff_A_MmIfOmpd2_0),.clk(gclk));
	jdff dff_A_UhhXUQQY4_0(.dout(w_dff_A_xN8E6Ghb2_0),.din(w_dff_A_UhhXUQQY4_0),.clk(gclk));
	jdff dff_A_xN8E6Ghb2_0(.dout(w_dff_A_PXYf0dZq4_0),.din(w_dff_A_xN8E6Ghb2_0),.clk(gclk));
	jdff dff_A_PXYf0dZq4_0(.dout(w_dff_A_hfN5wi7i8_0),.din(w_dff_A_PXYf0dZq4_0),.clk(gclk));
	jdff dff_A_hfN5wi7i8_0(.dout(w_dff_A_oPajINVY9_0),.din(w_dff_A_hfN5wi7i8_0),.clk(gclk));
	jdff dff_A_oPajINVY9_0(.dout(w_dff_A_pnYtcv6T3_0),.din(w_dff_A_oPajINVY9_0),.clk(gclk));
	jdff dff_A_pnYtcv6T3_0(.dout(w_dff_A_YkqGDftS9_0),.din(w_dff_A_pnYtcv6T3_0),.clk(gclk));
	jdff dff_A_YkqGDftS9_0(.dout(w_dff_A_RtToPjVr3_0),.din(w_dff_A_YkqGDftS9_0),.clk(gclk));
	jdff dff_A_RtToPjVr3_0(.dout(w_dff_A_ilREnJUH4_0),.din(w_dff_A_RtToPjVr3_0),.clk(gclk));
	jdff dff_A_ilREnJUH4_0(.dout(w_dff_A_FeK7bATw0_0),.din(w_dff_A_ilREnJUH4_0),.clk(gclk));
	jdff dff_A_FeK7bATw0_0(.dout(w_dff_A_lKYIe5Vw6_0),.din(w_dff_A_FeK7bATw0_0),.clk(gclk));
	jdff dff_A_lKYIe5Vw6_0(.dout(w_dff_A_wWOuanCo7_0),.din(w_dff_A_lKYIe5Vw6_0),.clk(gclk));
	jdff dff_A_wWOuanCo7_0(.dout(w_dff_A_E4l51J4X3_0),.din(w_dff_A_wWOuanCo7_0),.clk(gclk));
	jdff dff_A_E4l51J4X3_0(.dout(w_dff_A_f9ECAxSt3_0),.din(w_dff_A_E4l51J4X3_0),.clk(gclk));
	jdff dff_A_f9ECAxSt3_0(.dout(G448),.din(w_dff_A_f9ECAxSt3_0),.clk(gclk));
	jdff dff_A_uLsdXGj77_1(.dout(w_dff_A_NX1FLLKx8_0),.din(w_dff_A_uLsdXGj77_1),.clk(gclk));
	jdff dff_A_NX1FLLKx8_0(.dout(w_dff_A_i1fIY9VA9_0),.din(w_dff_A_NX1FLLKx8_0),.clk(gclk));
	jdff dff_A_i1fIY9VA9_0(.dout(w_dff_A_vinnMVKQ3_0),.din(w_dff_A_i1fIY9VA9_0),.clk(gclk));
	jdff dff_A_vinnMVKQ3_0(.dout(w_dff_A_Z6MLrGcd7_0),.din(w_dff_A_vinnMVKQ3_0),.clk(gclk));
	jdff dff_A_Z6MLrGcd7_0(.dout(w_dff_A_8HtCx68v9_0),.din(w_dff_A_Z6MLrGcd7_0),.clk(gclk));
	jdff dff_A_8HtCx68v9_0(.dout(w_dff_A_gZq3zVus4_0),.din(w_dff_A_8HtCx68v9_0),.clk(gclk));
	jdff dff_A_gZq3zVus4_0(.dout(w_dff_A_l7tOmevN2_0),.din(w_dff_A_gZq3zVus4_0),.clk(gclk));
	jdff dff_A_l7tOmevN2_0(.dout(w_dff_A_OgqSDkSL2_0),.din(w_dff_A_l7tOmevN2_0),.clk(gclk));
	jdff dff_A_OgqSDkSL2_0(.dout(w_dff_A_lPJuA1QS4_0),.din(w_dff_A_OgqSDkSL2_0),.clk(gclk));
	jdff dff_A_lPJuA1QS4_0(.dout(w_dff_A_nn0FKwip9_0),.din(w_dff_A_lPJuA1QS4_0),.clk(gclk));
	jdff dff_A_nn0FKwip9_0(.dout(w_dff_A_NsBrquGu9_0),.din(w_dff_A_nn0FKwip9_0),.clk(gclk));
	jdff dff_A_NsBrquGu9_0(.dout(w_dff_A_CSnJrBrw5_0),.din(w_dff_A_NsBrquGu9_0),.clk(gclk));
	jdff dff_A_CSnJrBrw5_0(.dout(w_dff_A_gP7CTIag1_0),.din(w_dff_A_CSnJrBrw5_0),.clk(gclk));
	jdff dff_A_gP7CTIag1_0(.dout(w_dff_A_L5iHt3dr8_0),.din(w_dff_A_gP7CTIag1_0),.clk(gclk));
	jdff dff_A_L5iHt3dr8_0(.dout(w_dff_A_K6JvbFWp4_0),.din(w_dff_A_L5iHt3dr8_0),.clk(gclk));
	jdff dff_A_K6JvbFWp4_0(.dout(w_dff_A_9fcGjbCy8_0),.din(w_dff_A_K6JvbFWp4_0),.clk(gclk));
	jdff dff_A_9fcGjbCy8_0(.dout(w_dff_A_wS6cb22j4_0),.din(w_dff_A_9fcGjbCy8_0),.clk(gclk));
	jdff dff_A_wS6cb22j4_0(.dout(w_dff_A_GX3cdPUI3_0),.din(w_dff_A_wS6cb22j4_0),.clk(gclk));
	jdff dff_A_GX3cdPUI3_0(.dout(w_dff_A_Lkvpz61y5_0),.din(w_dff_A_GX3cdPUI3_0),.clk(gclk));
	jdff dff_A_Lkvpz61y5_0(.dout(w_dff_A_GQehuQGn9_0),.din(w_dff_A_Lkvpz61y5_0),.clk(gclk));
	jdff dff_A_GQehuQGn9_0(.dout(w_dff_A_BMg5TUVv2_0),.din(w_dff_A_GQehuQGn9_0),.clk(gclk));
	jdff dff_A_BMg5TUVv2_0(.dout(w_dff_A_wZ2f8pTL6_0),.din(w_dff_A_BMg5TUVv2_0),.clk(gclk));
	jdff dff_A_wZ2f8pTL6_0(.dout(w_dff_A_83ZOiplb4_0),.din(w_dff_A_wZ2f8pTL6_0),.clk(gclk));
	jdff dff_A_83ZOiplb4_0(.dout(w_dff_A_cE5GgqAB8_0),.din(w_dff_A_83ZOiplb4_0),.clk(gclk));
	jdff dff_A_cE5GgqAB8_0(.dout(w_dff_A_GgNHQkRp9_0),.din(w_dff_A_cE5GgqAB8_0),.clk(gclk));
	jdff dff_A_GgNHQkRp9_0(.dout(w_dff_A_vIWR0YOL4_0),.din(w_dff_A_GgNHQkRp9_0),.clk(gclk));
	jdff dff_A_vIWR0YOL4_0(.dout(w_dff_A_w0W6kF634_0),.din(w_dff_A_vIWR0YOL4_0),.clk(gclk));
	jdff dff_A_w0W6kF634_0(.dout(w_dff_A_8os3EzAM6_0),.din(w_dff_A_w0W6kF634_0),.clk(gclk));
	jdff dff_A_8os3EzAM6_0(.dout(w_dff_A_7nuPcMTJ8_0),.din(w_dff_A_8os3EzAM6_0),.clk(gclk));
	jdff dff_A_7nuPcMTJ8_0(.dout(w_dff_A_fXIeBo3c7_0),.din(w_dff_A_7nuPcMTJ8_0),.clk(gclk));
	jdff dff_A_fXIeBo3c7_0(.dout(w_dff_A_DTuzhzlB3_0),.din(w_dff_A_fXIeBo3c7_0),.clk(gclk));
	jdff dff_A_DTuzhzlB3_0(.dout(w_dff_A_vbAbtqJV7_0),.din(w_dff_A_DTuzhzlB3_0),.clk(gclk));
	jdff dff_A_vbAbtqJV7_0(.dout(w_dff_A_FDpsTSAO0_0),.din(w_dff_A_vbAbtqJV7_0),.clk(gclk));
	jdff dff_A_FDpsTSAO0_0(.dout(w_dff_A_3PMa9iHI6_0),.din(w_dff_A_FDpsTSAO0_0),.clk(gclk));
	jdff dff_A_3PMa9iHI6_0(.dout(w_dff_A_cPOODtLB6_0),.din(w_dff_A_3PMa9iHI6_0),.clk(gclk));
	jdff dff_A_cPOODtLB6_0(.dout(w_dff_A_cH04DPs96_0),.din(w_dff_A_cPOODtLB6_0),.clk(gclk));
	jdff dff_A_cH04DPs96_0(.dout(w_dff_A_ybJM6jXC5_0),.din(w_dff_A_cH04DPs96_0),.clk(gclk));
	jdff dff_A_ybJM6jXC5_0(.dout(G444),.din(w_dff_A_ybJM6jXC5_0),.clk(gclk));
	jdff dff_A_2l1hqVy46_1(.dout(w_dff_A_9d3UVCu13_0),.din(w_dff_A_2l1hqVy46_1),.clk(gclk));
	jdff dff_A_9d3UVCu13_0(.dout(w_dff_A_KGfjFnLn0_0),.din(w_dff_A_9d3UVCu13_0),.clk(gclk));
	jdff dff_A_KGfjFnLn0_0(.dout(w_dff_A_Z6Fss6RC9_0),.din(w_dff_A_KGfjFnLn0_0),.clk(gclk));
	jdff dff_A_Z6Fss6RC9_0(.dout(w_dff_A_tf6WkaWM4_0),.din(w_dff_A_Z6Fss6RC9_0),.clk(gclk));
	jdff dff_A_tf6WkaWM4_0(.dout(w_dff_A_Jau20yRE0_0),.din(w_dff_A_tf6WkaWM4_0),.clk(gclk));
	jdff dff_A_Jau20yRE0_0(.dout(w_dff_A_H4CrkWjr8_0),.din(w_dff_A_Jau20yRE0_0),.clk(gclk));
	jdff dff_A_H4CrkWjr8_0(.dout(w_dff_A_qMt4R6XX4_0),.din(w_dff_A_H4CrkWjr8_0),.clk(gclk));
	jdff dff_A_qMt4R6XX4_0(.dout(w_dff_A_tRWnFen94_0),.din(w_dff_A_qMt4R6XX4_0),.clk(gclk));
	jdff dff_A_tRWnFen94_0(.dout(w_dff_A_pPyLbdqA5_0),.din(w_dff_A_tRWnFen94_0),.clk(gclk));
	jdff dff_A_pPyLbdqA5_0(.dout(w_dff_A_aFPXLgXY1_0),.din(w_dff_A_pPyLbdqA5_0),.clk(gclk));
	jdff dff_A_aFPXLgXY1_0(.dout(w_dff_A_8MX3tftK2_0),.din(w_dff_A_aFPXLgXY1_0),.clk(gclk));
	jdff dff_A_8MX3tftK2_0(.dout(w_dff_A_mSxr0lMG2_0),.din(w_dff_A_8MX3tftK2_0),.clk(gclk));
	jdff dff_A_mSxr0lMG2_0(.dout(w_dff_A_CAYi5kPi8_0),.din(w_dff_A_mSxr0lMG2_0),.clk(gclk));
	jdff dff_A_CAYi5kPi8_0(.dout(w_dff_A_tk7VeiD46_0),.din(w_dff_A_CAYi5kPi8_0),.clk(gclk));
	jdff dff_A_tk7VeiD46_0(.dout(w_dff_A_2YjvvqZ29_0),.din(w_dff_A_tk7VeiD46_0),.clk(gclk));
	jdff dff_A_2YjvvqZ29_0(.dout(w_dff_A_oYZRwpwO7_0),.din(w_dff_A_2YjvvqZ29_0),.clk(gclk));
	jdff dff_A_oYZRwpwO7_0(.dout(w_dff_A_dic5qb4a4_0),.din(w_dff_A_oYZRwpwO7_0),.clk(gclk));
	jdff dff_A_dic5qb4a4_0(.dout(w_dff_A_OmWpxsGv9_0),.din(w_dff_A_dic5qb4a4_0),.clk(gclk));
	jdff dff_A_OmWpxsGv9_0(.dout(w_dff_A_bZp5g0I93_0),.din(w_dff_A_OmWpxsGv9_0),.clk(gclk));
	jdff dff_A_bZp5g0I93_0(.dout(w_dff_A_kinliT5j2_0),.din(w_dff_A_bZp5g0I93_0),.clk(gclk));
	jdff dff_A_kinliT5j2_0(.dout(w_dff_A_5Hc9Ldb98_0),.din(w_dff_A_kinliT5j2_0),.clk(gclk));
	jdff dff_A_5Hc9Ldb98_0(.dout(w_dff_A_Dwc2Xno58_0),.din(w_dff_A_5Hc9Ldb98_0),.clk(gclk));
	jdff dff_A_Dwc2Xno58_0(.dout(w_dff_A_rmc3rdFx6_0),.din(w_dff_A_Dwc2Xno58_0),.clk(gclk));
	jdff dff_A_rmc3rdFx6_0(.dout(w_dff_A_3HQ4aECa5_0),.din(w_dff_A_rmc3rdFx6_0),.clk(gclk));
	jdff dff_A_3HQ4aECa5_0(.dout(w_dff_A_6L5t83EB3_0),.din(w_dff_A_3HQ4aECa5_0),.clk(gclk));
	jdff dff_A_6L5t83EB3_0(.dout(w_dff_A_jNTqtUKP1_0),.din(w_dff_A_6L5t83EB3_0),.clk(gclk));
	jdff dff_A_jNTqtUKP1_0(.dout(w_dff_A_e5cC8NpR5_0),.din(w_dff_A_jNTqtUKP1_0),.clk(gclk));
	jdff dff_A_e5cC8NpR5_0(.dout(w_dff_A_vFOy2fyY4_0),.din(w_dff_A_e5cC8NpR5_0),.clk(gclk));
	jdff dff_A_vFOy2fyY4_0(.dout(w_dff_A_8EL24QTX0_0),.din(w_dff_A_vFOy2fyY4_0),.clk(gclk));
	jdff dff_A_8EL24QTX0_0(.dout(w_dff_A_nqbQipO56_0),.din(w_dff_A_8EL24QTX0_0),.clk(gclk));
	jdff dff_A_nqbQipO56_0(.dout(w_dff_A_5cxFsShh1_0),.din(w_dff_A_nqbQipO56_0),.clk(gclk));
	jdff dff_A_5cxFsShh1_0(.dout(w_dff_A_nowipb605_0),.din(w_dff_A_5cxFsShh1_0),.clk(gclk));
	jdff dff_A_nowipb605_0(.dout(w_dff_A_SHE8aMfO7_0),.din(w_dff_A_nowipb605_0),.clk(gclk));
	jdff dff_A_SHE8aMfO7_0(.dout(w_dff_A_5wO5d7hK3_0),.din(w_dff_A_SHE8aMfO7_0),.clk(gclk));
	jdff dff_A_5wO5d7hK3_0(.dout(w_dff_A_dfNJmO6F8_0),.din(w_dff_A_5wO5d7hK3_0),.clk(gclk));
	jdff dff_A_dfNJmO6F8_0(.dout(w_dff_A_q2Ks7Jvr8_0),.din(w_dff_A_dfNJmO6F8_0),.clk(gclk));
	jdff dff_A_q2Ks7Jvr8_0(.dout(w_dff_A_2rX7MfhW7_0),.din(w_dff_A_q2Ks7Jvr8_0),.clk(gclk));
	jdff dff_A_2rX7MfhW7_0(.dout(G442),.din(w_dff_A_2rX7MfhW7_0),.clk(gclk));
	jdff dff_A_HiWLfWKP7_1(.dout(w_dff_A_0UCvrhVi4_0),.din(w_dff_A_HiWLfWKP7_1),.clk(gclk));
	jdff dff_A_0UCvrhVi4_0(.dout(w_dff_A_n8cv8puG5_0),.din(w_dff_A_0UCvrhVi4_0),.clk(gclk));
	jdff dff_A_n8cv8puG5_0(.dout(w_dff_A_RYvqZK1l1_0),.din(w_dff_A_n8cv8puG5_0),.clk(gclk));
	jdff dff_A_RYvqZK1l1_0(.dout(w_dff_A_ENzhW5jK9_0),.din(w_dff_A_RYvqZK1l1_0),.clk(gclk));
	jdff dff_A_ENzhW5jK9_0(.dout(w_dff_A_dVMDnWrn3_0),.din(w_dff_A_ENzhW5jK9_0),.clk(gclk));
	jdff dff_A_dVMDnWrn3_0(.dout(w_dff_A_8e1c2y0W5_0),.din(w_dff_A_dVMDnWrn3_0),.clk(gclk));
	jdff dff_A_8e1c2y0W5_0(.dout(w_dff_A_xRJmrmeE0_0),.din(w_dff_A_8e1c2y0W5_0),.clk(gclk));
	jdff dff_A_xRJmrmeE0_0(.dout(w_dff_A_ATMFP5mw9_0),.din(w_dff_A_xRJmrmeE0_0),.clk(gclk));
	jdff dff_A_ATMFP5mw9_0(.dout(w_dff_A_fNIQnVzC4_0),.din(w_dff_A_ATMFP5mw9_0),.clk(gclk));
	jdff dff_A_fNIQnVzC4_0(.dout(w_dff_A_C12bCA4o3_0),.din(w_dff_A_fNIQnVzC4_0),.clk(gclk));
	jdff dff_A_C12bCA4o3_0(.dout(w_dff_A_8ZbMhV4i6_0),.din(w_dff_A_C12bCA4o3_0),.clk(gclk));
	jdff dff_A_8ZbMhV4i6_0(.dout(w_dff_A_y9pz8Om91_0),.din(w_dff_A_8ZbMhV4i6_0),.clk(gclk));
	jdff dff_A_y9pz8Om91_0(.dout(w_dff_A_9NF812NG2_0),.din(w_dff_A_y9pz8Om91_0),.clk(gclk));
	jdff dff_A_9NF812NG2_0(.dout(w_dff_A_iqBQPIcQ3_0),.din(w_dff_A_9NF812NG2_0),.clk(gclk));
	jdff dff_A_iqBQPIcQ3_0(.dout(w_dff_A_RCkWIBlx8_0),.din(w_dff_A_iqBQPIcQ3_0),.clk(gclk));
	jdff dff_A_RCkWIBlx8_0(.dout(w_dff_A_bY3ubHh02_0),.din(w_dff_A_RCkWIBlx8_0),.clk(gclk));
	jdff dff_A_bY3ubHh02_0(.dout(w_dff_A_QfxCFLnc7_0),.din(w_dff_A_bY3ubHh02_0),.clk(gclk));
	jdff dff_A_QfxCFLnc7_0(.dout(w_dff_A_xfmKH9L01_0),.din(w_dff_A_QfxCFLnc7_0),.clk(gclk));
	jdff dff_A_xfmKH9L01_0(.dout(w_dff_A_KpNIUVEs0_0),.din(w_dff_A_xfmKH9L01_0),.clk(gclk));
	jdff dff_A_KpNIUVEs0_0(.dout(w_dff_A_MIrF1B9i2_0),.din(w_dff_A_KpNIUVEs0_0),.clk(gclk));
	jdff dff_A_MIrF1B9i2_0(.dout(w_dff_A_HzGvQglx0_0),.din(w_dff_A_MIrF1B9i2_0),.clk(gclk));
	jdff dff_A_HzGvQglx0_0(.dout(w_dff_A_4twZSC3O2_0),.din(w_dff_A_HzGvQglx0_0),.clk(gclk));
	jdff dff_A_4twZSC3O2_0(.dout(w_dff_A_kSagvAEW3_0),.din(w_dff_A_4twZSC3O2_0),.clk(gclk));
	jdff dff_A_kSagvAEW3_0(.dout(w_dff_A_IolfRFdE2_0),.din(w_dff_A_kSagvAEW3_0),.clk(gclk));
	jdff dff_A_IolfRFdE2_0(.dout(w_dff_A_GriAU1Pt1_0),.din(w_dff_A_IolfRFdE2_0),.clk(gclk));
	jdff dff_A_GriAU1Pt1_0(.dout(w_dff_A_667x8J2q8_0),.din(w_dff_A_GriAU1Pt1_0),.clk(gclk));
	jdff dff_A_667x8J2q8_0(.dout(w_dff_A_vLmPdVaY4_0),.din(w_dff_A_667x8J2q8_0),.clk(gclk));
	jdff dff_A_vLmPdVaY4_0(.dout(w_dff_A_9cXdnejb2_0),.din(w_dff_A_vLmPdVaY4_0),.clk(gclk));
	jdff dff_A_9cXdnejb2_0(.dout(w_dff_A_c9vUUgNJ6_0),.din(w_dff_A_9cXdnejb2_0),.clk(gclk));
	jdff dff_A_c9vUUgNJ6_0(.dout(w_dff_A_dSk0q1FY6_0),.din(w_dff_A_c9vUUgNJ6_0),.clk(gclk));
	jdff dff_A_dSk0q1FY6_0(.dout(w_dff_A_p8LBrKaF4_0),.din(w_dff_A_dSk0q1FY6_0),.clk(gclk));
	jdff dff_A_p8LBrKaF4_0(.dout(w_dff_A_LmEwFyAl4_0),.din(w_dff_A_p8LBrKaF4_0),.clk(gclk));
	jdff dff_A_LmEwFyAl4_0(.dout(w_dff_A_ipSodC7T5_0),.din(w_dff_A_LmEwFyAl4_0),.clk(gclk));
	jdff dff_A_ipSodC7T5_0(.dout(w_dff_A_frVC1RHd9_0),.din(w_dff_A_ipSodC7T5_0),.clk(gclk));
	jdff dff_A_frVC1RHd9_0(.dout(w_dff_A_9SQwtwIr4_0),.din(w_dff_A_frVC1RHd9_0),.clk(gclk));
	jdff dff_A_9SQwtwIr4_0(.dout(w_dff_A_pYiQIiIQ6_0),.din(w_dff_A_9SQwtwIr4_0),.clk(gclk));
	jdff dff_A_pYiQIiIQ6_0(.dout(w_dff_A_S2TA1OUr4_0),.din(w_dff_A_pYiQIiIQ6_0),.clk(gclk));
	jdff dff_A_S2TA1OUr4_0(.dout(G440),.din(w_dff_A_S2TA1OUr4_0),.clk(gclk));
	jdff dff_A_kvGxlUzO4_1(.dout(w_dff_A_HQiO5ttM3_0),.din(w_dff_A_kvGxlUzO4_1),.clk(gclk));
	jdff dff_A_HQiO5ttM3_0(.dout(w_dff_A_wDMwpEe39_0),.din(w_dff_A_HQiO5ttM3_0),.clk(gclk));
	jdff dff_A_wDMwpEe39_0(.dout(w_dff_A_D25LVPdq9_0),.din(w_dff_A_wDMwpEe39_0),.clk(gclk));
	jdff dff_A_D25LVPdq9_0(.dout(w_dff_A_LdqQ8GS96_0),.din(w_dff_A_D25LVPdq9_0),.clk(gclk));
	jdff dff_A_LdqQ8GS96_0(.dout(w_dff_A_g5SNYsFV2_0),.din(w_dff_A_LdqQ8GS96_0),.clk(gclk));
	jdff dff_A_g5SNYsFV2_0(.dout(w_dff_A_7VIbVF2i0_0),.din(w_dff_A_g5SNYsFV2_0),.clk(gclk));
	jdff dff_A_7VIbVF2i0_0(.dout(w_dff_A_u5gsozjE8_0),.din(w_dff_A_7VIbVF2i0_0),.clk(gclk));
	jdff dff_A_u5gsozjE8_0(.dout(w_dff_A_bYkPkdv60_0),.din(w_dff_A_u5gsozjE8_0),.clk(gclk));
	jdff dff_A_bYkPkdv60_0(.dout(w_dff_A_h6GV5PaT1_0),.din(w_dff_A_bYkPkdv60_0),.clk(gclk));
	jdff dff_A_h6GV5PaT1_0(.dout(w_dff_A_5GOGn6aE4_0),.din(w_dff_A_h6GV5PaT1_0),.clk(gclk));
	jdff dff_A_5GOGn6aE4_0(.dout(w_dff_A_4RwAOoPy3_0),.din(w_dff_A_5GOGn6aE4_0),.clk(gclk));
	jdff dff_A_4RwAOoPy3_0(.dout(w_dff_A_PO8kIc2X7_0),.din(w_dff_A_4RwAOoPy3_0),.clk(gclk));
	jdff dff_A_PO8kIc2X7_0(.dout(w_dff_A_G0oO1yNn5_0),.din(w_dff_A_PO8kIc2X7_0),.clk(gclk));
	jdff dff_A_G0oO1yNn5_0(.dout(w_dff_A_wcG2Op2J1_0),.din(w_dff_A_G0oO1yNn5_0),.clk(gclk));
	jdff dff_A_wcG2Op2J1_0(.dout(w_dff_A_GH70SxUr8_0),.din(w_dff_A_wcG2Op2J1_0),.clk(gclk));
	jdff dff_A_GH70SxUr8_0(.dout(w_dff_A_CcWFvBEL0_0),.din(w_dff_A_GH70SxUr8_0),.clk(gclk));
	jdff dff_A_CcWFvBEL0_0(.dout(w_dff_A_sf5jpRQu8_0),.din(w_dff_A_CcWFvBEL0_0),.clk(gclk));
	jdff dff_A_sf5jpRQu8_0(.dout(w_dff_A_0WgsX7tT0_0),.din(w_dff_A_sf5jpRQu8_0),.clk(gclk));
	jdff dff_A_0WgsX7tT0_0(.dout(w_dff_A_nnPg39Tz2_0),.din(w_dff_A_0WgsX7tT0_0),.clk(gclk));
	jdff dff_A_nnPg39Tz2_0(.dout(w_dff_A_SHnaC6LD5_0),.din(w_dff_A_nnPg39Tz2_0),.clk(gclk));
	jdff dff_A_SHnaC6LD5_0(.dout(w_dff_A_WaTtFhQm2_0),.din(w_dff_A_SHnaC6LD5_0),.clk(gclk));
	jdff dff_A_WaTtFhQm2_0(.dout(w_dff_A_hD38IotZ8_0),.din(w_dff_A_WaTtFhQm2_0),.clk(gclk));
	jdff dff_A_hD38IotZ8_0(.dout(w_dff_A_rGzf70ts7_0),.din(w_dff_A_hD38IotZ8_0),.clk(gclk));
	jdff dff_A_rGzf70ts7_0(.dout(w_dff_A_xRDBuaYF9_0),.din(w_dff_A_rGzf70ts7_0),.clk(gclk));
	jdff dff_A_xRDBuaYF9_0(.dout(w_dff_A_xcQvfbi58_0),.din(w_dff_A_xRDBuaYF9_0),.clk(gclk));
	jdff dff_A_xcQvfbi58_0(.dout(w_dff_A_SQGo8CdU4_0),.din(w_dff_A_xcQvfbi58_0),.clk(gclk));
	jdff dff_A_SQGo8CdU4_0(.dout(w_dff_A_LWbBRtU55_0),.din(w_dff_A_SQGo8CdU4_0),.clk(gclk));
	jdff dff_A_LWbBRtU55_0(.dout(w_dff_A_SvM85YHX4_0),.din(w_dff_A_LWbBRtU55_0),.clk(gclk));
	jdff dff_A_SvM85YHX4_0(.dout(w_dff_A_c7snQ1q51_0),.din(w_dff_A_SvM85YHX4_0),.clk(gclk));
	jdff dff_A_c7snQ1q51_0(.dout(w_dff_A_14omzql55_0),.din(w_dff_A_c7snQ1q51_0),.clk(gclk));
	jdff dff_A_14omzql55_0(.dout(w_dff_A_uIKWQI7U1_0),.din(w_dff_A_14omzql55_0),.clk(gclk));
	jdff dff_A_uIKWQI7U1_0(.dout(w_dff_A_GTQTm0DE4_0),.din(w_dff_A_uIKWQI7U1_0),.clk(gclk));
	jdff dff_A_GTQTm0DE4_0(.dout(w_dff_A_wYryfeQU2_0),.din(w_dff_A_GTQTm0DE4_0),.clk(gclk));
	jdff dff_A_wYryfeQU2_0(.dout(w_dff_A_R2ME4zqR4_0),.din(w_dff_A_wYryfeQU2_0),.clk(gclk));
	jdff dff_A_R2ME4zqR4_0(.dout(w_dff_A_V5LgGH9N4_0),.din(w_dff_A_R2ME4zqR4_0),.clk(gclk));
	jdff dff_A_V5LgGH9N4_0(.dout(w_dff_A_wCgTN6nU2_0),.din(w_dff_A_V5LgGH9N4_0),.clk(gclk));
	jdff dff_A_wCgTN6nU2_0(.dout(w_dff_A_pp9IsZJP3_0),.din(w_dff_A_wCgTN6nU2_0),.clk(gclk));
	jdff dff_A_pp9IsZJP3_0(.dout(G438),.din(w_dff_A_pp9IsZJP3_0),.clk(gclk));
	jdff dff_A_fKxVyEvG8_1(.dout(w_dff_A_F92hdeRJ0_0),.din(w_dff_A_fKxVyEvG8_1),.clk(gclk));
	jdff dff_A_F92hdeRJ0_0(.dout(w_dff_A_lh4qTxSA6_0),.din(w_dff_A_F92hdeRJ0_0),.clk(gclk));
	jdff dff_A_lh4qTxSA6_0(.dout(w_dff_A_Lj4aZEHl3_0),.din(w_dff_A_lh4qTxSA6_0),.clk(gclk));
	jdff dff_A_Lj4aZEHl3_0(.dout(w_dff_A_Ch9i7imW9_0),.din(w_dff_A_Lj4aZEHl3_0),.clk(gclk));
	jdff dff_A_Ch9i7imW9_0(.dout(w_dff_A_kCkxOE5N3_0),.din(w_dff_A_Ch9i7imW9_0),.clk(gclk));
	jdff dff_A_kCkxOE5N3_0(.dout(w_dff_A_dnWzRb6X7_0),.din(w_dff_A_kCkxOE5N3_0),.clk(gclk));
	jdff dff_A_dnWzRb6X7_0(.dout(w_dff_A_2SrkhawT5_0),.din(w_dff_A_dnWzRb6X7_0),.clk(gclk));
	jdff dff_A_2SrkhawT5_0(.dout(w_dff_A_J4ggTXvG5_0),.din(w_dff_A_2SrkhawT5_0),.clk(gclk));
	jdff dff_A_J4ggTXvG5_0(.dout(w_dff_A_laU8SMs35_0),.din(w_dff_A_J4ggTXvG5_0),.clk(gclk));
	jdff dff_A_laU8SMs35_0(.dout(w_dff_A_z1f7J1W22_0),.din(w_dff_A_laU8SMs35_0),.clk(gclk));
	jdff dff_A_z1f7J1W22_0(.dout(w_dff_A_FsoH9K6T3_0),.din(w_dff_A_z1f7J1W22_0),.clk(gclk));
	jdff dff_A_FsoH9K6T3_0(.dout(w_dff_A_IoUyw4J14_0),.din(w_dff_A_FsoH9K6T3_0),.clk(gclk));
	jdff dff_A_IoUyw4J14_0(.dout(w_dff_A_QURQmPgQ3_0),.din(w_dff_A_IoUyw4J14_0),.clk(gclk));
	jdff dff_A_QURQmPgQ3_0(.dout(w_dff_A_aLGroFPl3_0),.din(w_dff_A_QURQmPgQ3_0),.clk(gclk));
	jdff dff_A_aLGroFPl3_0(.dout(w_dff_A_LfcpGE3l3_0),.din(w_dff_A_aLGroFPl3_0),.clk(gclk));
	jdff dff_A_LfcpGE3l3_0(.dout(w_dff_A_EqJmcoBQ9_0),.din(w_dff_A_LfcpGE3l3_0),.clk(gclk));
	jdff dff_A_EqJmcoBQ9_0(.dout(w_dff_A_LUMKoF214_0),.din(w_dff_A_EqJmcoBQ9_0),.clk(gclk));
	jdff dff_A_LUMKoF214_0(.dout(w_dff_A_3yUQLkN69_0),.din(w_dff_A_LUMKoF214_0),.clk(gclk));
	jdff dff_A_3yUQLkN69_0(.dout(w_dff_A_bqDVKuKK3_0),.din(w_dff_A_3yUQLkN69_0),.clk(gclk));
	jdff dff_A_bqDVKuKK3_0(.dout(w_dff_A_SAUFHYGW9_0),.din(w_dff_A_bqDVKuKK3_0),.clk(gclk));
	jdff dff_A_SAUFHYGW9_0(.dout(w_dff_A_TAfyRZJC0_0),.din(w_dff_A_SAUFHYGW9_0),.clk(gclk));
	jdff dff_A_TAfyRZJC0_0(.dout(w_dff_A_LBPJll499_0),.din(w_dff_A_TAfyRZJC0_0),.clk(gclk));
	jdff dff_A_LBPJll499_0(.dout(w_dff_A_c2nudf8R7_0),.din(w_dff_A_LBPJll499_0),.clk(gclk));
	jdff dff_A_c2nudf8R7_0(.dout(w_dff_A_KcmDLKqn1_0),.din(w_dff_A_c2nudf8R7_0),.clk(gclk));
	jdff dff_A_KcmDLKqn1_0(.dout(w_dff_A_s16URw4I2_0),.din(w_dff_A_KcmDLKqn1_0),.clk(gclk));
	jdff dff_A_s16URw4I2_0(.dout(w_dff_A_5JPYUQsM5_0),.din(w_dff_A_s16URw4I2_0),.clk(gclk));
	jdff dff_A_5JPYUQsM5_0(.dout(w_dff_A_Idu8qWNB6_0),.din(w_dff_A_5JPYUQsM5_0),.clk(gclk));
	jdff dff_A_Idu8qWNB6_0(.dout(w_dff_A_1WWExI6x8_0),.din(w_dff_A_Idu8qWNB6_0),.clk(gclk));
	jdff dff_A_1WWExI6x8_0(.dout(w_dff_A_0mnoZRSQ5_0),.din(w_dff_A_1WWExI6x8_0),.clk(gclk));
	jdff dff_A_0mnoZRSQ5_0(.dout(w_dff_A_CF2GSWek0_0),.din(w_dff_A_0mnoZRSQ5_0),.clk(gclk));
	jdff dff_A_CF2GSWek0_0(.dout(w_dff_A_VQpVfuAR4_0),.din(w_dff_A_CF2GSWek0_0),.clk(gclk));
	jdff dff_A_VQpVfuAR4_0(.dout(w_dff_A_e170Ure11_0),.din(w_dff_A_VQpVfuAR4_0),.clk(gclk));
	jdff dff_A_e170Ure11_0(.dout(w_dff_A_3VILppcH7_0),.din(w_dff_A_e170Ure11_0),.clk(gclk));
	jdff dff_A_3VILppcH7_0(.dout(w_dff_A_l4NAm9en6_0),.din(w_dff_A_3VILppcH7_0),.clk(gclk));
	jdff dff_A_l4NAm9en6_0(.dout(w_dff_A_fDmTOJTi1_0),.din(w_dff_A_l4NAm9en6_0),.clk(gclk));
	jdff dff_A_fDmTOJTi1_0(.dout(w_dff_A_hph6m4e00_0),.din(w_dff_A_fDmTOJTi1_0),.clk(gclk));
	jdff dff_A_hph6m4e00_0(.dout(w_dff_A_PSZgYxFA9_0),.din(w_dff_A_hph6m4e00_0),.clk(gclk));
	jdff dff_A_PSZgYxFA9_0(.dout(G496),.din(w_dff_A_PSZgYxFA9_0),.clk(gclk));
	jdff dff_A_AcwEvtBl8_1(.dout(w_dff_A_6OWjTLXC6_0),.din(w_dff_A_AcwEvtBl8_1),.clk(gclk));
	jdff dff_A_6OWjTLXC6_0(.dout(w_dff_A_rpdzzsy26_0),.din(w_dff_A_6OWjTLXC6_0),.clk(gclk));
	jdff dff_A_rpdzzsy26_0(.dout(w_dff_A_RRnxiAJm6_0),.din(w_dff_A_rpdzzsy26_0),.clk(gclk));
	jdff dff_A_RRnxiAJm6_0(.dout(w_dff_A_Prlg8BjP1_0),.din(w_dff_A_RRnxiAJm6_0),.clk(gclk));
	jdff dff_A_Prlg8BjP1_0(.dout(w_dff_A_3bCnMy7x4_0),.din(w_dff_A_Prlg8BjP1_0),.clk(gclk));
	jdff dff_A_3bCnMy7x4_0(.dout(w_dff_A_LGjH8Pn65_0),.din(w_dff_A_3bCnMy7x4_0),.clk(gclk));
	jdff dff_A_LGjH8Pn65_0(.dout(w_dff_A_VYde3mL26_0),.din(w_dff_A_LGjH8Pn65_0),.clk(gclk));
	jdff dff_A_VYde3mL26_0(.dout(w_dff_A_aBaFFw074_0),.din(w_dff_A_VYde3mL26_0),.clk(gclk));
	jdff dff_A_aBaFFw074_0(.dout(w_dff_A_YqWJ6E5b9_0),.din(w_dff_A_aBaFFw074_0),.clk(gclk));
	jdff dff_A_YqWJ6E5b9_0(.dout(w_dff_A_ZRs2QVpA7_0),.din(w_dff_A_YqWJ6E5b9_0),.clk(gclk));
	jdff dff_A_ZRs2QVpA7_0(.dout(w_dff_A_9oebRl9I6_0),.din(w_dff_A_ZRs2QVpA7_0),.clk(gclk));
	jdff dff_A_9oebRl9I6_0(.dout(w_dff_A_hpjYXzxN6_0),.din(w_dff_A_9oebRl9I6_0),.clk(gclk));
	jdff dff_A_hpjYXzxN6_0(.dout(w_dff_A_OBgwRlmI9_0),.din(w_dff_A_hpjYXzxN6_0),.clk(gclk));
	jdff dff_A_OBgwRlmI9_0(.dout(w_dff_A_EnWHsSSQ6_0),.din(w_dff_A_OBgwRlmI9_0),.clk(gclk));
	jdff dff_A_EnWHsSSQ6_0(.dout(w_dff_A_ZqKAs4xj1_0),.din(w_dff_A_EnWHsSSQ6_0),.clk(gclk));
	jdff dff_A_ZqKAs4xj1_0(.dout(w_dff_A_mcCDbzoh3_0),.din(w_dff_A_ZqKAs4xj1_0),.clk(gclk));
	jdff dff_A_mcCDbzoh3_0(.dout(w_dff_A_4APlkpIW4_0),.din(w_dff_A_mcCDbzoh3_0),.clk(gclk));
	jdff dff_A_4APlkpIW4_0(.dout(w_dff_A_yGrE6SZE2_0),.din(w_dff_A_4APlkpIW4_0),.clk(gclk));
	jdff dff_A_yGrE6SZE2_0(.dout(w_dff_A_ch7R156V2_0),.din(w_dff_A_yGrE6SZE2_0),.clk(gclk));
	jdff dff_A_ch7R156V2_0(.dout(w_dff_A_bbSEe4Wi5_0),.din(w_dff_A_ch7R156V2_0),.clk(gclk));
	jdff dff_A_bbSEe4Wi5_0(.dout(w_dff_A_ebmEU7UJ1_0),.din(w_dff_A_bbSEe4Wi5_0),.clk(gclk));
	jdff dff_A_ebmEU7UJ1_0(.dout(w_dff_A_ww67YbTu2_0),.din(w_dff_A_ebmEU7UJ1_0),.clk(gclk));
	jdff dff_A_ww67YbTu2_0(.dout(w_dff_A_HNskSIVu3_0),.din(w_dff_A_ww67YbTu2_0),.clk(gclk));
	jdff dff_A_HNskSIVu3_0(.dout(w_dff_A_VKUvB8OA4_0),.din(w_dff_A_HNskSIVu3_0),.clk(gclk));
	jdff dff_A_VKUvB8OA4_0(.dout(w_dff_A_XE5PC3Zx2_0),.din(w_dff_A_VKUvB8OA4_0),.clk(gclk));
	jdff dff_A_XE5PC3Zx2_0(.dout(w_dff_A_iRRtSOHo3_0),.din(w_dff_A_XE5PC3Zx2_0),.clk(gclk));
	jdff dff_A_iRRtSOHo3_0(.dout(w_dff_A_UhSxZrF77_0),.din(w_dff_A_iRRtSOHo3_0),.clk(gclk));
	jdff dff_A_UhSxZrF77_0(.dout(w_dff_A_kTeJyuOT2_0),.din(w_dff_A_UhSxZrF77_0),.clk(gclk));
	jdff dff_A_kTeJyuOT2_0(.dout(w_dff_A_vWv3fmiR5_0),.din(w_dff_A_kTeJyuOT2_0),.clk(gclk));
	jdff dff_A_vWv3fmiR5_0(.dout(w_dff_A_w1lbupO53_0),.din(w_dff_A_vWv3fmiR5_0),.clk(gclk));
	jdff dff_A_w1lbupO53_0(.dout(w_dff_A_nBVCXKhB1_0),.din(w_dff_A_w1lbupO53_0),.clk(gclk));
	jdff dff_A_nBVCXKhB1_0(.dout(w_dff_A_QbV8s2JN4_0),.din(w_dff_A_nBVCXKhB1_0),.clk(gclk));
	jdff dff_A_QbV8s2JN4_0(.dout(w_dff_A_0d02QCDj3_0),.din(w_dff_A_QbV8s2JN4_0),.clk(gclk));
	jdff dff_A_0d02QCDj3_0(.dout(w_dff_A_Cy6LBfrM8_0),.din(w_dff_A_0d02QCDj3_0),.clk(gclk));
	jdff dff_A_Cy6LBfrM8_0(.dout(w_dff_A_K8hUt43B8_0),.din(w_dff_A_Cy6LBfrM8_0),.clk(gclk));
	jdff dff_A_K8hUt43B8_0(.dout(w_dff_A_JecLXnvU4_0),.din(w_dff_A_K8hUt43B8_0),.clk(gclk));
	jdff dff_A_JecLXnvU4_0(.dout(w_dff_A_NGD2okon1_0),.din(w_dff_A_JecLXnvU4_0),.clk(gclk));
	jdff dff_A_NGD2okon1_0(.dout(G494),.din(w_dff_A_NGD2okon1_0),.clk(gclk));
	jdff dff_A_z4lHrBEn5_1(.dout(w_dff_A_wMXkQfNZ7_0),.din(w_dff_A_z4lHrBEn5_1),.clk(gclk));
	jdff dff_A_wMXkQfNZ7_0(.dout(w_dff_A_PIHhjbMF1_0),.din(w_dff_A_wMXkQfNZ7_0),.clk(gclk));
	jdff dff_A_PIHhjbMF1_0(.dout(w_dff_A_7XwEtK6h9_0),.din(w_dff_A_PIHhjbMF1_0),.clk(gclk));
	jdff dff_A_7XwEtK6h9_0(.dout(w_dff_A_VeQmwW8d0_0),.din(w_dff_A_7XwEtK6h9_0),.clk(gclk));
	jdff dff_A_VeQmwW8d0_0(.dout(w_dff_A_1IcuaTuF8_0),.din(w_dff_A_VeQmwW8d0_0),.clk(gclk));
	jdff dff_A_1IcuaTuF8_0(.dout(w_dff_A_Q0bxyaBG9_0),.din(w_dff_A_1IcuaTuF8_0),.clk(gclk));
	jdff dff_A_Q0bxyaBG9_0(.dout(w_dff_A_AC23EK8I0_0),.din(w_dff_A_Q0bxyaBG9_0),.clk(gclk));
	jdff dff_A_AC23EK8I0_0(.dout(w_dff_A_1YFYwp1q0_0),.din(w_dff_A_AC23EK8I0_0),.clk(gclk));
	jdff dff_A_1YFYwp1q0_0(.dout(w_dff_A_0uSb1EZf5_0),.din(w_dff_A_1YFYwp1q0_0),.clk(gclk));
	jdff dff_A_0uSb1EZf5_0(.dout(w_dff_A_fba7M4lh6_0),.din(w_dff_A_0uSb1EZf5_0),.clk(gclk));
	jdff dff_A_fba7M4lh6_0(.dout(w_dff_A_1V4bVSun7_0),.din(w_dff_A_fba7M4lh6_0),.clk(gclk));
	jdff dff_A_1V4bVSun7_0(.dout(w_dff_A_GWUFa7EB2_0),.din(w_dff_A_1V4bVSun7_0),.clk(gclk));
	jdff dff_A_GWUFa7EB2_0(.dout(w_dff_A_ydN3znsn0_0),.din(w_dff_A_GWUFa7EB2_0),.clk(gclk));
	jdff dff_A_ydN3znsn0_0(.dout(w_dff_A_Wwalok0z5_0),.din(w_dff_A_ydN3znsn0_0),.clk(gclk));
	jdff dff_A_Wwalok0z5_0(.dout(w_dff_A_hVfJakKe3_0),.din(w_dff_A_Wwalok0z5_0),.clk(gclk));
	jdff dff_A_hVfJakKe3_0(.dout(w_dff_A_c6vz4bpA5_0),.din(w_dff_A_hVfJakKe3_0),.clk(gclk));
	jdff dff_A_c6vz4bpA5_0(.dout(w_dff_A_eAhWjZ4y4_0),.din(w_dff_A_c6vz4bpA5_0),.clk(gclk));
	jdff dff_A_eAhWjZ4y4_0(.dout(w_dff_A_5QBs58y93_0),.din(w_dff_A_eAhWjZ4y4_0),.clk(gclk));
	jdff dff_A_5QBs58y93_0(.dout(w_dff_A_QME7xHGK3_0),.din(w_dff_A_5QBs58y93_0),.clk(gclk));
	jdff dff_A_QME7xHGK3_0(.dout(w_dff_A_KUCDi4qU8_0),.din(w_dff_A_QME7xHGK3_0),.clk(gclk));
	jdff dff_A_KUCDi4qU8_0(.dout(w_dff_A_bKhBPAJF1_0),.din(w_dff_A_KUCDi4qU8_0),.clk(gclk));
	jdff dff_A_bKhBPAJF1_0(.dout(w_dff_A_M1Vyk1d97_0),.din(w_dff_A_bKhBPAJF1_0),.clk(gclk));
	jdff dff_A_M1Vyk1d97_0(.dout(w_dff_A_n9aHY8JG4_0),.din(w_dff_A_M1Vyk1d97_0),.clk(gclk));
	jdff dff_A_n9aHY8JG4_0(.dout(w_dff_A_jnuSaW5o8_0),.din(w_dff_A_n9aHY8JG4_0),.clk(gclk));
	jdff dff_A_jnuSaW5o8_0(.dout(w_dff_A_WUqwmtjw0_0),.din(w_dff_A_jnuSaW5o8_0),.clk(gclk));
	jdff dff_A_WUqwmtjw0_0(.dout(w_dff_A_KQt9Ye494_0),.din(w_dff_A_WUqwmtjw0_0),.clk(gclk));
	jdff dff_A_KQt9Ye494_0(.dout(w_dff_A_mNYPkUIT3_0),.din(w_dff_A_KQt9Ye494_0),.clk(gclk));
	jdff dff_A_mNYPkUIT3_0(.dout(w_dff_A_WPAyqyhM6_0),.din(w_dff_A_mNYPkUIT3_0),.clk(gclk));
	jdff dff_A_WPAyqyhM6_0(.dout(w_dff_A_sDJbfh4v8_0),.din(w_dff_A_WPAyqyhM6_0),.clk(gclk));
	jdff dff_A_sDJbfh4v8_0(.dout(w_dff_A_eF4yq6ZG2_0),.din(w_dff_A_sDJbfh4v8_0),.clk(gclk));
	jdff dff_A_eF4yq6ZG2_0(.dout(w_dff_A_rRUU0rwy4_0),.din(w_dff_A_eF4yq6ZG2_0),.clk(gclk));
	jdff dff_A_rRUU0rwy4_0(.dout(w_dff_A_SRz56pQD2_0),.din(w_dff_A_rRUU0rwy4_0),.clk(gclk));
	jdff dff_A_SRz56pQD2_0(.dout(w_dff_A_U23LyN9s0_0),.din(w_dff_A_SRz56pQD2_0),.clk(gclk));
	jdff dff_A_U23LyN9s0_0(.dout(w_dff_A_houm0qa04_0),.din(w_dff_A_U23LyN9s0_0),.clk(gclk));
	jdff dff_A_houm0qa04_0(.dout(w_dff_A_EWxXOe9A8_0),.din(w_dff_A_houm0qa04_0),.clk(gclk));
	jdff dff_A_EWxXOe9A8_0(.dout(w_dff_A_RA96IEze4_0),.din(w_dff_A_EWxXOe9A8_0),.clk(gclk));
	jdff dff_A_RA96IEze4_0(.dout(w_dff_A_8oeq2vBk5_0),.din(w_dff_A_RA96IEze4_0),.clk(gclk));
	jdff dff_A_8oeq2vBk5_0(.dout(G492),.din(w_dff_A_8oeq2vBk5_0),.clk(gclk));
	jdff dff_A_36IIFIIA7_1(.dout(w_dff_A_FkmA8tq38_0),.din(w_dff_A_36IIFIIA7_1),.clk(gclk));
	jdff dff_A_FkmA8tq38_0(.dout(w_dff_A_9aGlH3DO0_0),.din(w_dff_A_FkmA8tq38_0),.clk(gclk));
	jdff dff_A_9aGlH3DO0_0(.dout(w_dff_A_lMSm5W6U6_0),.din(w_dff_A_9aGlH3DO0_0),.clk(gclk));
	jdff dff_A_lMSm5W6U6_0(.dout(w_dff_A_prz6a1sx7_0),.din(w_dff_A_lMSm5W6U6_0),.clk(gclk));
	jdff dff_A_prz6a1sx7_0(.dout(w_dff_A_3cQzEwjl6_0),.din(w_dff_A_prz6a1sx7_0),.clk(gclk));
	jdff dff_A_3cQzEwjl6_0(.dout(w_dff_A_A3wrVfxj6_0),.din(w_dff_A_3cQzEwjl6_0),.clk(gclk));
	jdff dff_A_A3wrVfxj6_0(.dout(w_dff_A_ngJ6Fizn9_0),.din(w_dff_A_A3wrVfxj6_0),.clk(gclk));
	jdff dff_A_ngJ6Fizn9_0(.dout(w_dff_A_ePkytt8P6_0),.din(w_dff_A_ngJ6Fizn9_0),.clk(gclk));
	jdff dff_A_ePkytt8P6_0(.dout(w_dff_A_nKeN6kf55_0),.din(w_dff_A_ePkytt8P6_0),.clk(gclk));
	jdff dff_A_nKeN6kf55_0(.dout(w_dff_A_ukFQpkC67_0),.din(w_dff_A_nKeN6kf55_0),.clk(gclk));
	jdff dff_A_ukFQpkC67_0(.dout(w_dff_A_9wB1IUS94_0),.din(w_dff_A_ukFQpkC67_0),.clk(gclk));
	jdff dff_A_9wB1IUS94_0(.dout(w_dff_A_0sQPsP7I3_0),.din(w_dff_A_9wB1IUS94_0),.clk(gclk));
	jdff dff_A_0sQPsP7I3_0(.dout(w_dff_A_IYpIvJiJ2_0),.din(w_dff_A_0sQPsP7I3_0),.clk(gclk));
	jdff dff_A_IYpIvJiJ2_0(.dout(w_dff_A_OvqoPMTn3_0),.din(w_dff_A_IYpIvJiJ2_0),.clk(gclk));
	jdff dff_A_OvqoPMTn3_0(.dout(w_dff_A_9QwibUCc8_0),.din(w_dff_A_OvqoPMTn3_0),.clk(gclk));
	jdff dff_A_9QwibUCc8_0(.dout(w_dff_A_R1ICejDp3_0),.din(w_dff_A_9QwibUCc8_0),.clk(gclk));
	jdff dff_A_R1ICejDp3_0(.dout(w_dff_A_oN2D5d8m5_0),.din(w_dff_A_R1ICejDp3_0),.clk(gclk));
	jdff dff_A_oN2D5d8m5_0(.dout(w_dff_A_YuYOUTou0_0),.din(w_dff_A_oN2D5d8m5_0),.clk(gclk));
	jdff dff_A_YuYOUTou0_0(.dout(w_dff_A_U6BGYJb88_0),.din(w_dff_A_YuYOUTou0_0),.clk(gclk));
	jdff dff_A_U6BGYJb88_0(.dout(w_dff_A_47TVOq246_0),.din(w_dff_A_U6BGYJb88_0),.clk(gclk));
	jdff dff_A_47TVOq246_0(.dout(w_dff_A_PbVCMIuH5_0),.din(w_dff_A_47TVOq246_0),.clk(gclk));
	jdff dff_A_PbVCMIuH5_0(.dout(w_dff_A_ufFMvqlb0_0),.din(w_dff_A_PbVCMIuH5_0),.clk(gclk));
	jdff dff_A_ufFMvqlb0_0(.dout(w_dff_A_1M54oIVD0_0),.din(w_dff_A_ufFMvqlb0_0),.clk(gclk));
	jdff dff_A_1M54oIVD0_0(.dout(w_dff_A_BrK1dTY31_0),.din(w_dff_A_1M54oIVD0_0),.clk(gclk));
	jdff dff_A_BrK1dTY31_0(.dout(w_dff_A_YaIfHXcC6_0),.din(w_dff_A_BrK1dTY31_0),.clk(gclk));
	jdff dff_A_YaIfHXcC6_0(.dout(w_dff_A_gcwgr0Rl8_0),.din(w_dff_A_YaIfHXcC6_0),.clk(gclk));
	jdff dff_A_gcwgr0Rl8_0(.dout(w_dff_A_ybpOetFU3_0),.din(w_dff_A_gcwgr0Rl8_0),.clk(gclk));
	jdff dff_A_ybpOetFU3_0(.dout(w_dff_A_6hEOK7Eq8_0),.din(w_dff_A_ybpOetFU3_0),.clk(gclk));
	jdff dff_A_6hEOK7Eq8_0(.dout(w_dff_A_4Yhz2anG0_0),.din(w_dff_A_6hEOK7Eq8_0),.clk(gclk));
	jdff dff_A_4Yhz2anG0_0(.dout(w_dff_A_zRVHWq2I9_0),.din(w_dff_A_4Yhz2anG0_0),.clk(gclk));
	jdff dff_A_zRVHWq2I9_0(.dout(w_dff_A_32HSNbuY5_0),.din(w_dff_A_zRVHWq2I9_0),.clk(gclk));
	jdff dff_A_32HSNbuY5_0(.dout(w_dff_A_xA2Dcb131_0),.din(w_dff_A_32HSNbuY5_0),.clk(gclk));
	jdff dff_A_xA2Dcb131_0(.dout(w_dff_A_cd7WkMJc1_0),.din(w_dff_A_xA2Dcb131_0),.clk(gclk));
	jdff dff_A_cd7WkMJc1_0(.dout(w_dff_A_P6yfV3Ci3_0),.din(w_dff_A_cd7WkMJc1_0),.clk(gclk));
	jdff dff_A_P6yfV3Ci3_0(.dout(w_dff_A_DKS9rln26_0),.din(w_dff_A_P6yfV3Ci3_0),.clk(gclk));
	jdff dff_A_DKS9rln26_0(.dout(w_dff_A_gKtsmjWV7_0),.din(w_dff_A_DKS9rln26_0),.clk(gclk));
	jdff dff_A_gKtsmjWV7_0(.dout(w_dff_A_Kcmhynvt0_0),.din(w_dff_A_gKtsmjWV7_0),.clk(gclk));
	jdff dff_A_Kcmhynvt0_0(.dout(G490),.din(w_dff_A_Kcmhynvt0_0),.clk(gclk));
	jdff dff_A_DXzas7OV3_1(.dout(w_dff_A_DitevIQt4_0),.din(w_dff_A_DXzas7OV3_1),.clk(gclk));
	jdff dff_A_DitevIQt4_0(.dout(w_dff_A_gXqQdEKN7_0),.din(w_dff_A_DitevIQt4_0),.clk(gclk));
	jdff dff_A_gXqQdEKN7_0(.dout(w_dff_A_cqb7lCs85_0),.din(w_dff_A_gXqQdEKN7_0),.clk(gclk));
	jdff dff_A_cqb7lCs85_0(.dout(w_dff_A_KZ6waLow6_0),.din(w_dff_A_cqb7lCs85_0),.clk(gclk));
	jdff dff_A_KZ6waLow6_0(.dout(w_dff_A_KeltLhp16_0),.din(w_dff_A_KZ6waLow6_0),.clk(gclk));
	jdff dff_A_KeltLhp16_0(.dout(w_dff_A_Wt7Ebn225_0),.din(w_dff_A_KeltLhp16_0),.clk(gclk));
	jdff dff_A_Wt7Ebn225_0(.dout(w_dff_A_mlvYLxPi1_0),.din(w_dff_A_Wt7Ebn225_0),.clk(gclk));
	jdff dff_A_mlvYLxPi1_0(.dout(w_dff_A_M0xobwCI7_0),.din(w_dff_A_mlvYLxPi1_0),.clk(gclk));
	jdff dff_A_M0xobwCI7_0(.dout(w_dff_A_D25uNUG66_0),.din(w_dff_A_M0xobwCI7_0),.clk(gclk));
	jdff dff_A_D25uNUG66_0(.dout(w_dff_A_Cn9l1ycb3_0),.din(w_dff_A_D25uNUG66_0),.clk(gclk));
	jdff dff_A_Cn9l1ycb3_0(.dout(w_dff_A_nYnI3YW30_0),.din(w_dff_A_Cn9l1ycb3_0),.clk(gclk));
	jdff dff_A_nYnI3YW30_0(.dout(w_dff_A_XlR2KVD69_0),.din(w_dff_A_nYnI3YW30_0),.clk(gclk));
	jdff dff_A_XlR2KVD69_0(.dout(w_dff_A_lFNeG9137_0),.din(w_dff_A_XlR2KVD69_0),.clk(gclk));
	jdff dff_A_lFNeG9137_0(.dout(w_dff_A_7s3CsHRd6_0),.din(w_dff_A_lFNeG9137_0),.clk(gclk));
	jdff dff_A_7s3CsHRd6_0(.dout(w_dff_A_szt6NtZ92_0),.din(w_dff_A_7s3CsHRd6_0),.clk(gclk));
	jdff dff_A_szt6NtZ92_0(.dout(w_dff_A_AQOP14g49_0),.din(w_dff_A_szt6NtZ92_0),.clk(gclk));
	jdff dff_A_AQOP14g49_0(.dout(w_dff_A_aC1yb7r84_0),.din(w_dff_A_AQOP14g49_0),.clk(gclk));
	jdff dff_A_aC1yb7r84_0(.dout(w_dff_A_0AJZRDpq0_0),.din(w_dff_A_aC1yb7r84_0),.clk(gclk));
	jdff dff_A_0AJZRDpq0_0(.dout(w_dff_A_IOWH5kqj7_0),.din(w_dff_A_0AJZRDpq0_0),.clk(gclk));
	jdff dff_A_IOWH5kqj7_0(.dout(w_dff_A_CuRnAuZp7_0),.din(w_dff_A_IOWH5kqj7_0),.clk(gclk));
	jdff dff_A_CuRnAuZp7_0(.dout(w_dff_A_O6yepDJU3_0),.din(w_dff_A_CuRnAuZp7_0),.clk(gclk));
	jdff dff_A_O6yepDJU3_0(.dout(w_dff_A_lkxaeDzS6_0),.din(w_dff_A_O6yepDJU3_0),.clk(gclk));
	jdff dff_A_lkxaeDzS6_0(.dout(w_dff_A_oPkwPXyi7_0),.din(w_dff_A_lkxaeDzS6_0),.clk(gclk));
	jdff dff_A_oPkwPXyi7_0(.dout(w_dff_A_M3HGtLT02_0),.din(w_dff_A_oPkwPXyi7_0),.clk(gclk));
	jdff dff_A_M3HGtLT02_0(.dout(w_dff_A_F3Ojr0sb4_0),.din(w_dff_A_M3HGtLT02_0),.clk(gclk));
	jdff dff_A_F3Ojr0sb4_0(.dout(w_dff_A_7Xl7WXQP8_0),.din(w_dff_A_F3Ojr0sb4_0),.clk(gclk));
	jdff dff_A_7Xl7WXQP8_0(.dout(w_dff_A_KsFnX82u9_0),.din(w_dff_A_7Xl7WXQP8_0),.clk(gclk));
	jdff dff_A_KsFnX82u9_0(.dout(w_dff_A_5KInHmCx2_0),.din(w_dff_A_KsFnX82u9_0),.clk(gclk));
	jdff dff_A_5KInHmCx2_0(.dout(w_dff_A_MSMhMbcC5_0),.din(w_dff_A_5KInHmCx2_0),.clk(gclk));
	jdff dff_A_MSMhMbcC5_0(.dout(w_dff_A_lEu24tQd8_0),.din(w_dff_A_MSMhMbcC5_0),.clk(gclk));
	jdff dff_A_lEu24tQd8_0(.dout(w_dff_A_6FfYaLH39_0),.din(w_dff_A_lEu24tQd8_0),.clk(gclk));
	jdff dff_A_6FfYaLH39_0(.dout(w_dff_A_NT84FmHo9_0),.din(w_dff_A_6FfYaLH39_0),.clk(gclk));
	jdff dff_A_NT84FmHo9_0(.dout(w_dff_A_2fnemDXS9_0),.din(w_dff_A_NT84FmHo9_0),.clk(gclk));
	jdff dff_A_2fnemDXS9_0(.dout(w_dff_A_hADZS1ol7_0),.din(w_dff_A_2fnemDXS9_0),.clk(gclk));
	jdff dff_A_hADZS1ol7_0(.dout(w_dff_A_HFGnETG61_0),.din(w_dff_A_hADZS1ol7_0),.clk(gclk));
	jdff dff_A_HFGnETG61_0(.dout(w_dff_A_J3VE4y9D9_0),.din(w_dff_A_HFGnETG61_0),.clk(gclk));
	jdff dff_A_J3VE4y9D9_0(.dout(w_dff_A_oSWjikhs8_0),.din(w_dff_A_J3VE4y9D9_0),.clk(gclk));
	jdff dff_A_oSWjikhs8_0(.dout(G488),.din(w_dff_A_oSWjikhs8_0),.clk(gclk));
	jdff dff_A_8wLrcBEf7_1(.dout(w_dff_A_MBtpf6nG4_0),.din(w_dff_A_8wLrcBEf7_1),.clk(gclk));
	jdff dff_A_MBtpf6nG4_0(.dout(w_dff_A_zTds5Dbw1_0),.din(w_dff_A_MBtpf6nG4_0),.clk(gclk));
	jdff dff_A_zTds5Dbw1_0(.dout(w_dff_A_dLAi06If4_0),.din(w_dff_A_zTds5Dbw1_0),.clk(gclk));
	jdff dff_A_dLAi06If4_0(.dout(w_dff_A_i9I3egDZ9_0),.din(w_dff_A_dLAi06If4_0),.clk(gclk));
	jdff dff_A_i9I3egDZ9_0(.dout(w_dff_A_5gnGIPUa4_0),.din(w_dff_A_i9I3egDZ9_0),.clk(gclk));
	jdff dff_A_5gnGIPUa4_0(.dout(w_dff_A_7Nvh6Vgj4_0),.din(w_dff_A_5gnGIPUa4_0),.clk(gclk));
	jdff dff_A_7Nvh6Vgj4_0(.dout(w_dff_A_erCiyXWt7_0),.din(w_dff_A_7Nvh6Vgj4_0),.clk(gclk));
	jdff dff_A_erCiyXWt7_0(.dout(w_dff_A_TYHneHoA3_0),.din(w_dff_A_erCiyXWt7_0),.clk(gclk));
	jdff dff_A_TYHneHoA3_0(.dout(w_dff_A_FWqguuIS8_0),.din(w_dff_A_TYHneHoA3_0),.clk(gclk));
	jdff dff_A_FWqguuIS8_0(.dout(w_dff_A_Kz9cUupp4_0),.din(w_dff_A_FWqguuIS8_0),.clk(gclk));
	jdff dff_A_Kz9cUupp4_0(.dout(w_dff_A_LhcF0VFA1_0),.din(w_dff_A_Kz9cUupp4_0),.clk(gclk));
	jdff dff_A_LhcF0VFA1_0(.dout(w_dff_A_TWLJK79o0_0),.din(w_dff_A_LhcF0VFA1_0),.clk(gclk));
	jdff dff_A_TWLJK79o0_0(.dout(w_dff_A_AhAOzCav7_0),.din(w_dff_A_TWLJK79o0_0),.clk(gclk));
	jdff dff_A_AhAOzCav7_0(.dout(w_dff_A_pJDYz61E3_0),.din(w_dff_A_AhAOzCav7_0),.clk(gclk));
	jdff dff_A_pJDYz61E3_0(.dout(w_dff_A_MgswgbaL1_0),.din(w_dff_A_pJDYz61E3_0),.clk(gclk));
	jdff dff_A_MgswgbaL1_0(.dout(w_dff_A_mBbmJr9x4_0),.din(w_dff_A_MgswgbaL1_0),.clk(gclk));
	jdff dff_A_mBbmJr9x4_0(.dout(w_dff_A_mwi9elKe0_0),.din(w_dff_A_mBbmJr9x4_0),.clk(gclk));
	jdff dff_A_mwi9elKe0_0(.dout(w_dff_A_8h8XM6yw7_0),.din(w_dff_A_mwi9elKe0_0),.clk(gclk));
	jdff dff_A_8h8XM6yw7_0(.dout(w_dff_A_0Fb1Z5739_0),.din(w_dff_A_8h8XM6yw7_0),.clk(gclk));
	jdff dff_A_0Fb1Z5739_0(.dout(w_dff_A_QdUUU36t8_0),.din(w_dff_A_0Fb1Z5739_0),.clk(gclk));
	jdff dff_A_QdUUU36t8_0(.dout(w_dff_A_UZ1PALCw1_0),.din(w_dff_A_QdUUU36t8_0),.clk(gclk));
	jdff dff_A_UZ1PALCw1_0(.dout(w_dff_A_K0ll3kxt0_0),.din(w_dff_A_UZ1PALCw1_0),.clk(gclk));
	jdff dff_A_K0ll3kxt0_0(.dout(w_dff_A_tdS0yNrO9_0),.din(w_dff_A_K0ll3kxt0_0),.clk(gclk));
	jdff dff_A_tdS0yNrO9_0(.dout(w_dff_A_fUBM5kay7_0),.din(w_dff_A_tdS0yNrO9_0),.clk(gclk));
	jdff dff_A_fUBM5kay7_0(.dout(w_dff_A_1LCeM0fm7_0),.din(w_dff_A_fUBM5kay7_0),.clk(gclk));
	jdff dff_A_1LCeM0fm7_0(.dout(w_dff_A_a6FGzUCU1_0),.din(w_dff_A_1LCeM0fm7_0),.clk(gclk));
	jdff dff_A_a6FGzUCU1_0(.dout(w_dff_A_cDyH5COV3_0),.din(w_dff_A_a6FGzUCU1_0),.clk(gclk));
	jdff dff_A_cDyH5COV3_0(.dout(w_dff_A_anFDywGS0_0),.din(w_dff_A_cDyH5COV3_0),.clk(gclk));
	jdff dff_A_anFDywGS0_0(.dout(w_dff_A_PqpMyNmQ3_0),.din(w_dff_A_anFDywGS0_0),.clk(gclk));
	jdff dff_A_PqpMyNmQ3_0(.dout(w_dff_A_NJDgWsIe4_0),.din(w_dff_A_PqpMyNmQ3_0),.clk(gclk));
	jdff dff_A_NJDgWsIe4_0(.dout(w_dff_A_A4NiK8Pt5_0),.din(w_dff_A_NJDgWsIe4_0),.clk(gclk));
	jdff dff_A_A4NiK8Pt5_0(.dout(w_dff_A_JZ2xUKIN3_0),.din(w_dff_A_A4NiK8Pt5_0),.clk(gclk));
	jdff dff_A_JZ2xUKIN3_0(.dout(w_dff_A_wjYWRq041_0),.din(w_dff_A_JZ2xUKIN3_0),.clk(gclk));
	jdff dff_A_wjYWRq041_0(.dout(w_dff_A_RCutgdgV5_0),.din(w_dff_A_wjYWRq041_0),.clk(gclk));
	jdff dff_A_RCutgdgV5_0(.dout(w_dff_A_RuGhyXir1_0),.din(w_dff_A_RCutgdgV5_0),.clk(gclk));
	jdff dff_A_RuGhyXir1_0(.dout(w_dff_A_MySFxhTV8_0),.din(w_dff_A_RuGhyXir1_0),.clk(gclk));
	jdff dff_A_MySFxhTV8_0(.dout(w_dff_A_es4GlcNn2_0),.din(w_dff_A_MySFxhTV8_0),.clk(gclk));
	jdff dff_A_es4GlcNn2_0(.dout(G486),.din(w_dff_A_es4GlcNn2_0),.clk(gclk));
	jdff dff_A_0XQfGMjy7_1(.dout(w_dff_A_GmWmMbMS4_0),.din(w_dff_A_0XQfGMjy7_1),.clk(gclk));
	jdff dff_A_GmWmMbMS4_0(.dout(w_dff_A_xfon8w0f5_0),.din(w_dff_A_GmWmMbMS4_0),.clk(gclk));
	jdff dff_A_xfon8w0f5_0(.dout(w_dff_A_dpXPvg7D6_0),.din(w_dff_A_xfon8w0f5_0),.clk(gclk));
	jdff dff_A_dpXPvg7D6_0(.dout(w_dff_A_CVj0Pjvs7_0),.din(w_dff_A_dpXPvg7D6_0),.clk(gclk));
	jdff dff_A_CVj0Pjvs7_0(.dout(w_dff_A_qAfRDUAY1_0),.din(w_dff_A_CVj0Pjvs7_0),.clk(gclk));
	jdff dff_A_qAfRDUAY1_0(.dout(w_dff_A_QfNvzWUm6_0),.din(w_dff_A_qAfRDUAY1_0),.clk(gclk));
	jdff dff_A_QfNvzWUm6_0(.dout(w_dff_A_eNVXP6yO2_0),.din(w_dff_A_QfNvzWUm6_0),.clk(gclk));
	jdff dff_A_eNVXP6yO2_0(.dout(w_dff_A_OLvJPhHz4_0),.din(w_dff_A_eNVXP6yO2_0),.clk(gclk));
	jdff dff_A_OLvJPhHz4_0(.dout(w_dff_A_hcvwTh5I5_0),.din(w_dff_A_OLvJPhHz4_0),.clk(gclk));
	jdff dff_A_hcvwTh5I5_0(.dout(w_dff_A_bCeKO90o8_0),.din(w_dff_A_hcvwTh5I5_0),.clk(gclk));
	jdff dff_A_bCeKO90o8_0(.dout(w_dff_A_s8ITB5Uc1_0),.din(w_dff_A_bCeKO90o8_0),.clk(gclk));
	jdff dff_A_s8ITB5Uc1_0(.dout(w_dff_A_RjgeXgxr9_0),.din(w_dff_A_s8ITB5Uc1_0),.clk(gclk));
	jdff dff_A_RjgeXgxr9_0(.dout(w_dff_A_u3rMyb6D9_0),.din(w_dff_A_RjgeXgxr9_0),.clk(gclk));
	jdff dff_A_u3rMyb6D9_0(.dout(w_dff_A_Tn0hMPUG9_0),.din(w_dff_A_u3rMyb6D9_0),.clk(gclk));
	jdff dff_A_Tn0hMPUG9_0(.dout(w_dff_A_SWymwAb43_0),.din(w_dff_A_Tn0hMPUG9_0),.clk(gclk));
	jdff dff_A_SWymwAb43_0(.dout(w_dff_A_bzW8e2QY6_0),.din(w_dff_A_SWymwAb43_0),.clk(gclk));
	jdff dff_A_bzW8e2QY6_0(.dout(w_dff_A_siXEcYW97_0),.din(w_dff_A_bzW8e2QY6_0),.clk(gclk));
	jdff dff_A_siXEcYW97_0(.dout(w_dff_A_Ecx6SjWU4_0),.din(w_dff_A_siXEcYW97_0),.clk(gclk));
	jdff dff_A_Ecx6SjWU4_0(.dout(w_dff_A_VwCWuPYR3_0),.din(w_dff_A_Ecx6SjWU4_0),.clk(gclk));
	jdff dff_A_VwCWuPYR3_0(.dout(w_dff_A_eZclCqGA6_0),.din(w_dff_A_VwCWuPYR3_0),.clk(gclk));
	jdff dff_A_eZclCqGA6_0(.dout(w_dff_A_jL2jo5bH9_0),.din(w_dff_A_eZclCqGA6_0),.clk(gclk));
	jdff dff_A_jL2jo5bH9_0(.dout(w_dff_A_AOQ49JsI8_0),.din(w_dff_A_jL2jo5bH9_0),.clk(gclk));
	jdff dff_A_AOQ49JsI8_0(.dout(w_dff_A_iZMLTyxH9_0),.din(w_dff_A_AOQ49JsI8_0),.clk(gclk));
	jdff dff_A_iZMLTyxH9_0(.dout(w_dff_A_oKnyiuwN2_0),.din(w_dff_A_iZMLTyxH9_0),.clk(gclk));
	jdff dff_A_oKnyiuwN2_0(.dout(w_dff_A_9fE7aXkZ7_0),.din(w_dff_A_oKnyiuwN2_0),.clk(gclk));
	jdff dff_A_9fE7aXkZ7_0(.dout(w_dff_A_H9OV5D8P3_0),.din(w_dff_A_9fE7aXkZ7_0),.clk(gclk));
	jdff dff_A_H9OV5D8P3_0(.dout(w_dff_A_tS1YKY697_0),.din(w_dff_A_H9OV5D8P3_0),.clk(gclk));
	jdff dff_A_tS1YKY697_0(.dout(w_dff_A_CDkfbcBc1_0),.din(w_dff_A_tS1YKY697_0),.clk(gclk));
	jdff dff_A_CDkfbcBc1_0(.dout(w_dff_A_b8Mrjkzo9_0),.din(w_dff_A_CDkfbcBc1_0),.clk(gclk));
	jdff dff_A_b8Mrjkzo9_0(.dout(w_dff_A_efP6I1qo1_0),.din(w_dff_A_b8Mrjkzo9_0),.clk(gclk));
	jdff dff_A_efP6I1qo1_0(.dout(w_dff_A_Ty0eUYJ12_0),.din(w_dff_A_efP6I1qo1_0),.clk(gclk));
	jdff dff_A_Ty0eUYJ12_0(.dout(w_dff_A_xDMHUktA4_0),.din(w_dff_A_Ty0eUYJ12_0),.clk(gclk));
	jdff dff_A_xDMHUktA4_0(.dout(w_dff_A_mDxoQrm45_0),.din(w_dff_A_xDMHUktA4_0),.clk(gclk));
	jdff dff_A_mDxoQrm45_0(.dout(w_dff_A_uCFJA9Sx9_0),.din(w_dff_A_mDxoQrm45_0),.clk(gclk));
	jdff dff_A_uCFJA9Sx9_0(.dout(w_dff_A_xQXYupyA1_0),.din(w_dff_A_uCFJA9Sx9_0),.clk(gclk));
	jdff dff_A_xQXYupyA1_0(.dout(w_dff_A_vNexCwex3_0),.din(w_dff_A_xQXYupyA1_0),.clk(gclk));
	jdff dff_A_vNexCwex3_0(.dout(w_dff_A_gZjphLfx4_0),.din(w_dff_A_vNexCwex3_0),.clk(gclk));
	jdff dff_A_gZjphLfx4_0(.dout(G484),.din(w_dff_A_gZjphLfx4_0),.clk(gclk));
	jdff dff_A_azIhLlon4_1(.dout(w_dff_A_aX7lGb0V6_0),.din(w_dff_A_azIhLlon4_1),.clk(gclk));
	jdff dff_A_aX7lGb0V6_0(.dout(w_dff_A_BVr18Mkg6_0),.din(w_dff_A_aX7lGb0V6_0),.clk(gclk));
	jdff dff_A_BVr18Mkg6_0(.dout(w_dff_A_7IjS7lU89_0),.din(w_dff_A_BVr18Mkg6_0),.clk(gclk));
	jdff dff_A_7IjS7lU89_0(.dout(w_dff_A_f0wHBvQ86_0),.din(w_dff_A_7IjS7lU89_0),.clk(gclk));
	jdff dff_A_f0wHBvQ86_0(.dout(w_dff_A_5gzUUM279_0),.din(w_dff_A_f0wHBvQ86_0),.clk(gclk));
	jdff dff_A_5gzUUM279_0(.dout(w_dff_A_nTOv59km5_0),.din(w_dff_A_5gzUUM279_0),.clk(gclk));
	jdff dff_A_nTOv59km5_0(.dout(w_dff_A_O0HAABJw1_0),.din(w_dff_A_nTOv59km5_0),.clk(gclk));
	jdff dff_A_O0HAABJw1_0(.dout(w_dff_A_aOl1XXUs2_0),.din(w_dff_A_O0HAABJw1_0),.clk(gclk));
	jdff dff_A_aOl1XXUs2_0(.dout(w_dff_A_fhLYO8NA7_0),.din(w_dff_A_aOl1XXUs2_0),.clk(gclk));
	jdff dff_A_fhLYO8NA7_0(.dout(w_dff_A_xaMWc1gD3_0),.din(w_dff_A_fhLYO8NA7_0),.clk(gclk));
	jdff dff_A_xaMWc1gD3_0(.dout(w_dff_A_SyVGQfqx2_0),.din(w_dff_A_xaMWc1gD3_0),.clk(gclk));
	jdff dff_A_SyVGQfqx2_0(.dout(w_dff_A_19Y0Xrxv7_0),.din(w_dff_A_SyVGQfqx2_0),.clk(gclk));
	jdff dff_A_19Y0Xrxv7_0(.dout(w_dff_A_QXfnmOgn3_0),.din(w_dff_A_19Y0Xrxv7_0),.clk(gclk));
	jdff dff_A_QXfnmOgn3_0(.dout(w_dff_A_MDxKriLN4_0),.din(w_dff_A_QXfnmOgn3_0),.clk(gclk));
	jdff dff_A_MDxKriLN4_0(.dout(w_dff_A_KwSkPwEL1_0),.din(w_dff_A_MDxKriLN4_0),.clk(gclk));
	jdff dff_A_KwSkPwEL1_0(.dout(w_dff_A_fGAuh8jG0_0),.din(w_dff_A_KwSkPwEL1_0),.clk(gclk));
	jdff dff_A_fGAuh8jG0_0(.dout(w_dff_A_Vl3eqJhC7_0),.din(w_dff_A_fGAuh8jG0_0),.clk(gclk));
	jdff dff_A_Vl3eqJhC7_0(.dout(w_dff_A_9JF6gBlC6_0),.din(w_dff_A_Vl3eqJhC7_0),.clk(gclk));
	jdff dff_A_9JF6gBlC6_0(.dout(w_dff_A_3wCsGf8m6_0),.din(w_dff_A_9JF6gBlC6_0),.clk(gclk));
	jdff dff_A_3wCsGf8m6_0(.dout(w_dff_A_E5FGXIej3_0),.din(w_dff_A_3wCsGf8m6_0),.clk(gclk));
	jdff dff_A_E5FGXIej3_0(.dout(w_dff_A_vuSVhI3f8_0),.din(w_dff_A_E5FGXIej3_0),.clk(gclk));
	jdff dff_A_vuSVhI3f8_0(.dout(w_dff_A_sgL9W5m90_0),.din(w_dff_A_vuSVhI3f8_0),.clk(gclk));
	jdff dff_A_sgL9W5m90_0(.dout(w_dff_A_lgmrrzQR3_0),.din(w_dff_A_sgL9W5m90_0),.clk(gclk));
	jdff dff_A_lgmrrzQR3_0(.dout(w_dff_A_jvqZIyvX9_0),.din(w_dff_A_lgmrrzQR3_0),.clk(gclk));
	jdff dff_A_jvqZIyvX9_0(.dout(w_dff_A_92QMTkZo8_0),.din(w_dff_A_jvqZIyvX9_0),.clk(gclk));
	jdff dff_A_92QMTkZo8_0(.dout(w_dff_A_DhptXEy64_0),.din(w_dff_A_92QMTkZo8_0),.clk(gclk));
	jdff dff_A_DhptXEy64_0(.dout(w_dff_A_kbsjlWvv7_0),.din(w_dff_A_DhptXEy64_0),.clk(gclk));
	jdff dff_A_kbsjlWvv7_0(.dout(w_dff_A_xMmYfnOj8_0),.din(w_dff_A_kbsjlWvv7_0),.clk(gclk));
	jdff dff_A_xMmYfnOj8_0(.dout(w_dff_A_GRJr3iAi0_0),.din(w_dff_A_xMmYfnOj8_0),.clk(gclk));
	jdff dff_A_GRJr3iAi0_0(.dout(w_dff_A_ZWEhvrVo6_0),.din(w_dff_A_GRJr3iAi0_0),.clk(gclk));
	jdff dff_A_ZWEhvrVo6_0(.dout(w_dff_A_UP7ljwom8_0),.din(w_dff_A_ZWEhvrVo6_0),.clk(gclk));
	jdff dff_A_UP7ljwom8_0(.dout(w_dff_A_uvrF2HIT8_0),.din(w_dff_A_UP7ljwom8_0),.clk(gclk));
	jdff dff_A_uvrF2HIT8_0(.dout(w_dff_A_lWV9yiZL0_0),.din(w_dff_A_uvrF2HIT8_0),.clk(gclk));
	jdff dff_A_lWV9yiZL0_0(.dout(w_dff_A_I2oZQKlL1_0),.din(w_dff_A_lWV9yiZL0_0),.clk(gclk));
	jdff dff_A_I2oZQKlL1_0(.dout(w_dff_A_Z2UxhWsj7_0),.din(w_dff_A_I2oZQKlL1_0),.clk(gclk));
	jdff dff_A_Z2UxhWsj7_0(.dout(w_dff_A_IjTnKPUP4_0),.din(w_dff_A_Z2UxhWsj7_0),.clk(gclk));
	jdff dff_A_IjTnKPUP4_0(.dout(w_dff_A_0bdAFRdb1_0),.din(w_dff_A_IjTnKPUP4_0),.clk(gclk));
	jdff dff_A_0bdAFRdb1_0(.dout(G482),.din(w_dff_A_0bdAFRdb1_0),.clk(gclk));
	jdff dff_A_OfRm1bFs5_1(.dout(w_dff_A_6KmIy3PK6_0),.din(w_dff_A_OfRm1bFs5_1),.clk(gclk));
	jdff dff_A_6KmIy3PK6_0(.dout(w_dff_A_aYfHaKv06_0),.din(w_dff_A_6KmIy3PK6_0),.clk(gclk));
	jdff dff_A_aYfHaKv06_0(.dout(w_dff_A_ZejgaIp97_0),.din(w_dff_A_aYfHaKv06_0),.clk(gclk));
	jdff dff_A_ZejgaIp97_0(.dout(w_dff_A_yzGc5Yw31_0),.din(w_dff_A_ZejgaIp97_0),.clk(gclk));
	jdff dff_A_yzGc5Yw31_0(.dout(w_dff_A_xqMcAvkU1_0),.din(w_dff_A_yzGc5Yw31_0),.clk(gclk));
	jdff dff_A_xqMcAvkU1_0(.dout(w_dff_A_R59MYq8p2_0),.din(w_dff_A_xqMcAvkU1_0),.clk(gclk));
	jdff dff_A_R59MYq8p2_0(.dout(w_dff_A_tiPOHG574_0),.din(w_dff_A_R59MYq8p2_0),.clk(gclk));
	jdff dff_A_tiPOHG574_0(.dout(w_dff_A_zkTwiCE67_0),.din(w_dff_A_tiPOHG574_0),.clk(gclk));
	jdff dff_A_zkTwiCE67_0(.dout(w_dff_A_2Z5sOrnG3_0),.din(w_dff_A_zkTwiCE67_0),.clk(gclk));
	jdff dff_A_2Z5sOrnG3_0(.dout(w_dff_A_0g1jZ2Ei2_0),.din(w_dff_A_2Z5sOrnG3_0),.clk(gclk));
	jdff dff_A_0g1jZ2Ei2_0(.dout(w_dff_A_sxPu2aiE8_0),.din(w_dff_A_0g1jZ2Ei2_0),.clk(gclk));
	jdff dff_A_sxPu2aiE8_0(.dout(w_dff_A_qXHISY2e5_0),.din(w_dff_A_sxPu2aiE8_0),.clk(gclk));
	jdff dff_A_qXHISY2e5_0(.dout(w_dff_A_5V6AmOpN0_0),.din(w_dff_A_qXHISY2e5_0),.clk(gclk));
	jdff dff_A_5V6AmOpN0_0(.dout(w_dff_A_IeZXgIph9_0),.din(w_dff_A_5V6AmOpN0_0),.clk(gclk));
	jdff dff_A_IeZXgIph9_0(.dout(w_dff_A_6HeGVw1M1_0),.din(w_dff_A_IeZXgIph9_0),.clk(gclk));
	jdff dff_A_6HeGVw1M1_0(.dout(w_dff_A_bxVfAVKx8_0),.din(w_dff_A_6HeGVw1M1_0),.clk(gclk));
	jdff dff_A_bxVfAVKx8_0(.dout(w_dff_A_UF25iH2F4_0),.din(w_dff_A_bxVfAVKx8_0),.clk(gclk));
	jdff dff_A_UF25iH2F4_0(.dout(w_dff_A_7lydPKM67_0),.din(w_dff_A_UF25iH2F4_0),.clk(gclk));
	jdff dff_A_7lydPKM67_0(.dout(w_dff_A_12i31rrE7_0),.din(w_dff_A_7lydPKM67_0),.clk(gclk));
	jdff dff_A_12i31rrE7_0(.dout(w_dff_A_aZccxvds0_0),.din(w_dff_A_12i31rrE7_0),.clk(gclk));
	jdff dff_A_aZccxvds0_0(.dout(w_dff_A_Jg6GTRmk2_0),.din(w_dff_A_aZccxvds0_0),.clk(gclk));
	jdff dff_A_Jg6GTRmk2_0(.dout(w_dff_A_uO8ThcsR6_0),.din(w_dff_A_Jg6GTRmk2_0),.clk(gclk));
	jdff dff_A_uO8ThcsR6_0(.dout(w_dff_A_ryiJoZyX0_0),.din(w_dff_A_uO8ThcsR6_0),.clk(gclk));
	jdff dff_A_ryiJoZyX0_0(.dout(w_dff_A_x43oecP31_0),.din(w_dff_A_ryiJoZyX0_0),.clk(gclk));
	jdff dff_A_x43oecP31_0(.dout(w_dff_A_LcnKBECF8_0),.din(w_dff_A_x43oecP31_0),.clk(gclk));
	jdff dff_A_LcnKBECF8_0(.dout(w_dff_A_askDIDOz1_0),.din(w_dff_A_LcnKBECF8_0),.clk(gclk));
	jdff dff_A_askDIDOz1_0(.dout(w_dff_A_yp5eiI6D2_0),.din(w_dff_A_askDIDOz1_0),.clk(gclk));
	jdff dff_A_yp5eiI6D2_0(.dout(w_dff_A_0pgN7H7a9_0),.din(w_dff_A_yp5eiI6D2_0),.clk(gclk));
	jdff dff_A_0pgN7H7a9_0(.dout(w_dff_A_J0Cl8Llt1_0),.din(w_dff_A_0pgN7H7a9_0),.clk(gclk));
	jdff dff_A_J0Cl8Llt1_0(.dout(w_dff_A_MsnsuOBh0_0),.din(w_dff_A_J0Cl8Llt1_0),.clk(gclk));
	jdff dff_A_MsnsuOBh0_0(.dout(w_dff_A_JlaKHGbb1_0),.din(w_dff_A_MsnsuOBh0_0),.clk(gclk));
	jdff dff_A_JlaKHGbb1_0(.dout(w_dff_A_7H0JS3R56_0),.din(w_dff_A_JlaKHGbb1_0),.clk(gclk));
	jdff dff_A_7H0JS3R56_0(.dout(w_dff_A_S70F4loh0_0),.din(w_dff_A_7H0JS3R56_0),.clk(gclk));
	jdff dff_A_S70F4loh0_0(.dout(w_dff_A_L0KI4wXP4_0),.din(w_dff_A_S70F4loh0_0),.clk(gclk));
	jdff dff_A_L0KI4wXP4_0(.dout(w_dff_A_NrQNIThS3_0),.din(w_dff_A_L0KI4wXP4_0),.clk(gclk));
	jdff dff_A_NrQNIThS3_0(.dout(w_dff_A_B7IuYAhl5_0),.din(w_dff_A_NrQNIThS3_0),.clk(gclk));
	jdff dff_A_B7IuYAhl5_0(.dout(w_dff_A_M8AkHDF90_0),.din(w_dff_A_B7IuYAhl5_0),.clk(gclk));
	jdff dff_A_M8AkHDF90_0(.dout(G480),.din(w_dff_A_M8AkHDF90_0),.clk(gclk));
	jdff dff_A_4CAs5RJf1_1(.dout(w_dff_A_QMx2GvSa2_0),.din(w_dff_A_4CAs5RJf1_1),.clk(gclk));
	jdff dff_A_QMx2GvSa2_0(.dout(w_dff_A_pSrOzuj04_0),.din(w_dff_A_QMx2GvSa2_0),.clk(gclk));
	jdff dff_A_pSrOzuj04_0(.dout(w_dff_A_w6mjS1H76_0),.din(w_dff_A_pSrOzuj04_0),.clk(gclk));
	jdff dff_A_w6mjS1H76_0(.dout(w_dff_A_KIIoL9qz8_0),.din(w_dff_A_w6mjS1H76_0),.clk(gclk));
	jdff dff_A_KIIoL9qz8_0(.dout(w_dff_A_geGPXntj4_0),.din(w_dff_A_KIIoL9qz8_0),.clk(gclk));
	jdff dff_A_geGPXntj4_0(.dout(w_dff_A_8ZxDRM5e6_0),.din(w_dff_A_geGPXntj4_0),.clk(gclk));
	jdff dff_A_8ZxDRM5e6_0(.dout(w_dff_A_Jn6DX5Do3_0),.din(w_dff_A_8ZxDRM5e6_0),.clk(gclk));
	jdff dff_A_Jn6DX5Do3_0(.dout(w_dff_A_Q8F5g7S29_0),.din(w_dff_A_Jn6DX5Do3_0),.clk(gclk));
	jdff dff_A_Q8F5g7S29_0(.dout(w_dff_A_UxBbbfbk4_0),.din(w_dff_A_Q8F5g7S29_0),.clk(gclk));
	jdff dff_A_UxBbbfbk4_0(.dout(w_dff_A_AjFpM39c8_0),.din(w_dff_A_UxBbbfbk4_0),.clk(gclk));
	jdff dff_A_AjFpM39c8_0(.dout(w_dff_A_1m3PDwZa2_0),.din(w_dff_A_AjFpM39c8_0),.clk(gclk));
	jdff dff_A_1m3PDwZa2_0(.dout(w_dff_A_vmH4HACf8_0),.din(w_dff_A_1m3PDwZa2_0),.clk(gclk));
	jdff dff_A_vmH4HACf8_0(.dout(w_dff_A_xwXVKDmV3_0),.din(w_dff_A_vmH4HACf8_0),.clk(gclk));
	jdff dff_A_xwXVKDmV3_0(.dout(w_dff_A_eAEiSS7W8_0),.din(w_dff_A_xwXVKDmV3_0),.clk(gclk));
	jdff dff_A_eAEiSS7W8_0(.dout(w_dff_A_YO3aOyis2_0),.din(w_dff_A_eAEiSS7W8_0),.clk(gclk));
	jdff dff_A_YO3aOyis2_0(.dout(w_dff_A_8tlymgnb3_0),.din(w_dff_A_YO3aOyis2_0),.clk(gclk));
	jdff dff_A_8tlymgnb3_0(.dout(w_dff_A_kZWwcbLK3_0),.din(w_dff_A_8tlymgnb3_0),.clk(gclk));
	jdff dff_A_kZWwcbLK3_0(.dout(w_dff_A_QN2zhAZ00_0),.din(w_dff_A_kZWwcbLK3_0),.clk(gclk));
	jdff dff_A_QN2zhAZ00_0(.dout(w_dff_A_Iw8tVeJe3_0),.din(w_dff_A_QN2zhAZ00_0),.clk(gclk));
	jdff dff_A_Iw8tVeJe3_0(.dout(w_dff_A_A3NyS7Sa5_0),.din(w_dff_A_Iw8tVeJe3_0),.clk(gclk));
	jdff dff_A_A3NyS7Sa5_0(.dout(w_dff_A_4b5jcwNx0_0),.din(w_dff_A_A3NyS7Sa5_0),.clk(gclk));
	jdff dff_A_4b5jcwNx0_0(.dout(w_dff_A_sch38MpP0_0),.din(w_dff_A_4b5jcwNx0_0),.clk(gclk));
	jdff dff_A_sch38MpP0_0(.dout(w_dff_A_oTwkmGe08_0),.din(w_dff_A_sch38MpP0_0),.clk(gclk));
	jdff dff_A_oTwkmGe08_0(.dout(w_dff_A_zgtpWmSx4_0),.din(w_dff_A_oTwkmGe08_0),.clk(gclk));
	jdff dff_A_zgtpWmSx4_0(.dout(w_dff_A_4x3UBLSF8_0),.din(w_dff_A_zgtpWmSx4_0),.clk(gclk));
	jdff dff_A_4x3UBLSF8_0(.dout(w_dff_A_yxhFuPQj5_0),.din(w_dff_A_4x3UBLSF8_0),.clk(gclk));
	jdff dff_A_yxhFuPQj5_0(.dout(w_dff_A_OLMT80EA4_0),.din(w_dff_A_yxhFuPQj5_0),.clk(gclk));
	jdff dff_A_OLMT80EA4_0(.dout(w_dff_A_8owFwn9k2_0),.din(w_dff_A_OLMT80EA4_0),.clk(gclk));
	jdff dff_A_8owFwn9k2_0(.dout(w_dff_A_XP7bJKId0_0),.din(w_dff_A_8owFwn9k2_0),.clk(gclk));
	jdff dff_A_XP7bJKId0_0(.dout(w_dff_A_5aZy4HNv7_0),.din(w_dff_A_XP7bJKId0_0),.clk(gclk));
	jdff dff_A_5aZy4HNv7_0(.dout(w_dff_A_s5UK2fwQ1_0),.din(w_dff_A_5aZy4HNv7_0),.clk(gclk));
	jdff dff_A_s5UK2fwQ1_0(.dout(w_dff_A_dIiYmdtN4_0),.din(w_dff_A_s5UK2fwQ1_0),.clk(gclk));
	jdff dff_A_dIiYmdtN4_0(.dout(w_dff_A_OZgHfJat0_0),.din(w_dff_A_dIiYmdtN4_0),.clk(gclk));
	jdff dff_A_OZgHfJat0_0(.dout(w_dff_A_4XJbp7bv6_0),.din(w_dff_A_OZgHfJat0_0),.clk(gclk));
	jdff dff_A_4XJbp7bv6_0(.dout(w_dff_A_gPxA2HPg8_0),.din(w_dff_A_4XJbp7bv6_0),.clk(gclk));
	jdff dff_A_gPxA2HPg8_0(.dout(w_dff_A_pGa0lBVM3_0),.din(w_dff_A_gPxA2HPg8_0),.clk(gclk));
	jdff dff_A_pGa0lBVM3_0(.dout(w_dff_A_L3bN9oRH5_0),.din(w_dff_A_pGa0lBVM3_0),.clk(gclk));
	jdff dff_A_L3bN9oRH5_0(.dout(G560),.din(w_dff_A_L3bN9oRH5_0),.clk(gclk));
	jdff dff_A_C0h2PJSo2_1(.dout(w_dff_A_3ZlSs3ql0_0),.din(w_dff_A_C0h2PJSo2_1),.clk(gclk));
	jdff dff_A_3ZlSs3ql0_0(.dout(w_dff_A_u4y4jl7v3_0),.din(w_dff_A_3ZlSs3ql0_0),.clk(gclk));
	jdff dff_A_u4y4jl7v3_0(.dout(w_dff_A_s6AQ10ey3_0),.din(w_dff_A_u4y4jl7v3_0),.clk(gclk));
	jdff dff_A_s6AQ10ey3_0(.dout(w_dff_A_nxrKI0JN5_0),.din(w_dff_A_s6AQ10ey3_0),.clk(gclk));
	jdff dff_A_nxrKI0JN5_0(.dout(w_dff_A_4ln3jjCC8_0),.din(w_dff_A_nxrKI0JN5_0),.clk(gclk));
	jdff dff_A_4ln3jjCC8_0(.dout(w_dff_A_5Yh2akrM3_0),.din(w_dff_A_4ln3jjCC8_0),.clk(gclk));
	jdff dff_A_5Yh2akrM3_0(.dout(w_dff_A_yFRi18p44_0),.din(w_dff_A_5Yh2akrM3_0),.clk(gclk));
	jdff dff_A_yFRi18p44_0(.dout(w_dff_A_oYyNcA7M6_0),.din(w_dff_A_yFRi18p44_0),.clk(gclk));
	jdff dff_A_oYyNcA7M6_0(.dout(w_dff_A_oNu8gdjv7_0),.din(w_dff_A_oYyNcA7M6_0),.clk(gclk));
	jdff dff_A_oNu8gdjv7_0(.dout(w_dff_A_RTGOMqj45_0),.din(w_dff_A_oNu8gdjv7_0),.clk(gclk));
	jdff dff_A_RTGOMqj45_0(.dout(w_dff_A_9SOpOpus0_0),.din(w_dff_A_RTGOMqj45_0),.clk(gclk));
	jdff dff_A_9SOpOpus0_0(.dout(w_dff_A_ABGEGEJA6_0),.din(w_dff_A_9SOpOpus0_0),.clk(gclk));
	jdff dff_A_ABGEGEJA6_0(.dout(w_dff_A_SIe8LqtX6_0),.din(w_dff_A_ABGEGEJA6_0),.clk(gclk));
	jdff dff_A_SIe8LqtX6_0(.dout(w_dff_A_iVpJPaOb8_0),.din(w_dff_A_SIe8LqtX6_0),.clk(gclk));
	jdff dff_A_iVpJPaOb8_0(.dout(w_dff_A_6BmYJTgU8_0),.din(w_dff_A_iVpJPaOb8_0),.clk(gclk));
	jdff dff_A_6BmYJTgU8_0(.dout(w_dff_A_GrpZCmGt9_0),.din(w_dff_A_6BmYJTgU8_0),.clk(gclk));
	jdff dff_A_GrpZCmGt9_0(.dout(w_dff_A_Ij9f2J918_0),.din(w_dff_A_GrpZCmGt9_0),.clk(gclk));
	jdff dff_A_Ij9f2J918_0(.dout(w_dff_A_RLU4wszg0_0),.din(w_dff_A_Ij9f2J918_0),.clk(gclk));
	jdff dff_A_RLU4wszg0_0(.dout(w_dff_A_LgTtKnGd6_0),.din(w_dff_A_RLU4wszg0_0),.clk(gclk));
	jdff dff_A_LgTtKnGd6_0(.dout(w_dff_A_6anem5Lo0_0),.din(w_dff_A_LgTtKnGd6_0),.clk(gclk));
	jdff dff_A_6anem5Lo0_0(.dout(w_dff_A_we5WbZM39_0),.din(w_dff_A_6anem5Lo0_0),.clk(gclk));
	jdff dff_A_we5WbZM39_0(.dout(w_dff_A_2CQsupRd5_0),.din(w_dff_A_we5WbZM39_0),.clk(gclk));
	jdff dff_A_2CQsupRd5_0(.dout(w_dff_A_ps2xr9Xj4_0),.din(w_dff_A_2CQsupRd5_0),.clk(gclk));
	jdff dff_A_ps2xr9Xj4_0(.dout(w_dff_A_O9lqSmp91_0),.din(w_dff_A_ps2xr9Xj4_0),.clk(gclk));
	jdff dff_A_O9lqSmp91_0(.dout(w_dff_A_WVvNACZO4_0),.din(w_dff_A_O9lqSmp91_0),.clk(gclk));
	jdff dff_A_WVvNACZO4_0(.dout(w_dff_A_Vk368qoA7_0),.din(w_dff_A_WVvNACZO4_0),.clk(gclk));
	jdff dff_A_Vk368qoA7_0(.dout(w_dff_A_7zsfv1wu5_0),.din(w_dff_A_Vk368qoA7_0),.clk(gclk));
	jdff dff_A_7zsfv1wu5_0(.dout(w_dff_A_bLGWfnQL5_0),.din(w_dff_A_7zsfv1wu5_0),.clk(gclk));
	jdff dff_A_bLGWfnQL5_0(.dout(w_dff_A_dAcC6USf3_0),.din(w_dff_A_bLGWfnQL5_0),.clk(gclk));
	jdff dff_A_dAcC6USf3_0(.dout(w_dff_A_JIUqB4bi5_0),.din(w_dff_A_dAcC6USf3_0),.clk(gclk));
	jdff dff_A_JIUqB4bi5_0(.dout(w_dff_A_vEfoIVrU5_0),.din(w_dff_A_JIUqB4bi5_0),.clk(gclk));
	jdff dff_A_vEfoIVrU5_0(.dout(w_dff_A_4ED88eQB2_0),.din(w_dff_A_vEfoIVrU5_0),.clk(gclk));
	jdff dff_A_4ED88eQB2_0(.dout(w_dff_A_fptj2er38_0),.din(w_dff_A_4ED88eQB2_0),.clk(gclk));
	jdff dff_A_fptj2er38_0(.dout(w_dff_A_hPEzMaVO1_0),.din(w_dff_A_fptj2er38_0),.clk(gclk));
	jdff dff_A_hPEzMaVO1_0(.dout(w_dff_A_TttMYAGY1_0),.din(w_dff_A_hPEzMaVO1_0),.clk(gclk));
	jdff dff_A_TttMYAGY1_0(.dout(w_dff_A_0ZNHaH8t7_0),.din(w_dff_A_TttMYAGY1_0),.clk(gclk));
	jdff dff_A_0ZNHaH8t7_0(.dout(w_dff_A_1kvOQdXn9_0),.din(w_dff_A_0ZNHaH8t7_0),.clk(gclk));
	jdff dff_A_1kvOQdXn9_0(.dout(G542),.din(w_dff_A_1kvOQdXn9_0),.clk(gclk));
	jdff dff_A_pxhHMs847_1(.dout(w_dff_A_VsW5jftS6_0),.din(w_dff_A_pxhHMs847_1),.clk(gclk));
	jdff dff_A_VsW5jftS6_0(.dout(w_dff_A_JgySY6F13_0),.din(w_dff_A_VsW5jftS6_0),.clk(gclk));
	jdff dff_A_JgySY6F13_0(.dout(w_dff_A_9sVR3Bsm9_0),.din(w_dff_A_JgySY6F13_0),.clk(gclk));
	jdff dff_A_9sVR3Bsm9_0(.dout(w_dff_A_4IHpVARz4_0),.din(w_dff_A_9sVR3Bsm9_0),.clk(gclk));
	jdff dff_A_4IHpVARz4_0(.dout(w_dff_A_jeD6TjU52_0),.din(w_dff_A_4IHpVARz4_0),.clk(gclk));
	jdff dff_A_jeD6TjU52_0(.dout(w_dff_A_udeU1dBJ2_0),.din(w_dff_A_jeD6TjU52_0),.clk(gclk));
	jdff dff_A_udeU1dBJ2_0(.dout(w_dff_A_WadM1TZy1_0),.din(w_dff_A_udeU1dBJ2_0),.clk(gclk));
	jdff dff_A_WadM1TZy1_0(.dout(w_dff_A_iG0Oa1QY8_0),.din(w_dff_A_WadM1TZy1_0),.clk(gclk));
	jdff dff_A_iG0Oa1QY8_0(.dout(w_dff_A_yqICLXAO0_0),.din(w_dff_A_iG0Oa1QY8_0),.clk(gclk));
	jdff dff_A_yqICLXAO0_0(.dout(w_dff_A_XR9DT6Ab2_0),.din(w_dff_A_yqICLXAO0_0),.clk(gclk));
	jdff dff_A_XR9DT6Ab2_0(.dout(w_dff_A_W7zwRZey1_0),.din(w_dff_A_XR9DT6Ab2_0),.clk(gclk));
	jdff dff_A_W7zwRZey1_0(.dout(w_dff_A_5CeLt9wu6_0),.din(w_dff_A_W7zwRZey1_0),.clk(gclk));
	jdff dff_A_5CeLt9wu6_0(.dout(w_dff_A_zCdns82z9_0),.din(w_dff_A_5CeLt9wu6_0),.clk(gclk));
	jdff dff_A_zCdns82z9_0(.dout(w_dff_A_o19kE1385_0),.din(w_dff_A_zCdns82z9_0),.clk(gclk));
	jdff dff_A_o19kE1385_0(.dout(w_dff_A_CRP9tPGI1_0),.din(w_dff_A_o19kE1385_0),.clk(gclk));
	jdff dff_A_CRP9tPGI1_0(.dout(w_dff_A_BYt7de0p9_0),.din(w_dff_A_CRP9tPGI1_0),.clk(gclk));
	jdff dff_A_BYt7de0p9_0(.dout(w_dff_A_uR1WvLjb3_0),.din(w_dff_A_BYt7de0p9_0),.clk(gclk));
	jdff dff_A_uR1WvLjb3_0(.dout(w_dff_A_3dSBGSdb4_0),.din(w_dff_A_uR1WvLjb3_0),.clk(gclk));
	jdff dff_A_3dSBGSdb4_0(.dout(w_dff_A_PYstLBrc4_0),.din(w_dff_A_3dSBGSdb4_0),.clk(gclk));
	jdff dff_A_PYstLBrc4_0(.dout(w_dff_A_qS2eEVGC4_0),.din(w_dff_A_PYstLBrc4_0),.clk(gclk));
	jdff dff_A_qS2eEVGC4_0(.dout(w_dff_A_rO4RnK5C1_0),.din(w_dff_A_qS2eEVGC4_0),.clk(gclk));
	jdff dff_A_rO4RnK5C1_0(.dout(w_dff_A_iTjdMU746_0),.din(w_dff_A_rO4RnK5C1_0),.clk(gclk));
	jdff dff_A_iTjdMU746_0(.dout(w_dff_A_iBVr8gmg1_0),.din(w_dff_A_iTjdMU746_0),.clk(gclk));
	jdff dff_A_iBVr8gmg1_0(.dout(w_dff_A_TNdRy4995_0),.din(w_dff_A_iBVr8gmg1_0),.clk(gclk));
	jdff dff_A_TNdRy4995_0(.dout(w_dff_A_bdntXmWL8_0),.din(w_dff_A_TNdRy4995_0),.clk(gclk));
	jdff dff_A_bdntXmWL8_0(.dout(w_dff_A_C6YvucMg7_0),.din(w_dff_A_bdntXmWL8_0),.clk(gclk));
	jdff dff_A_C6YvucMg7_0(.dout(w_dff_A_5jVqDDGp3_0),.din(w_dff_A_C6YvucMg7_0),.clk(gclk));
	jdff dff_A_5jVqDDGp3_0(.dout(w_dff_A_Ofw10gvI4_0),.din(w_dff_A_5jVqDDGp3_0),.clk(gclk));
	jdff dff_A_Ofw10gvI4_0(.dout(w_dff_A_lYmDq50Z4_0),.din(w_dff_A_Ofw10gvI4_0),.clk(gclk));
	jdff dff_A_lYmDq50Z4_0(.dout(w_dff_A_hsfvckSQ1_0),.din(w_dff_A_lYmDq50Z4_0),.clk(gclk));
	jdff dff_A_hsfvckSQ1_0(.dout(w_dff_A_LBYiaKUj8_0),.din(w_dff_A_hsfvckSQ1_0),.clk(gclk));
	jdff dff_A_LBYiaKUj8_0(.dout(w_dff_A_ecvZcZ1M3_0),.din(w_dff_A_LBYiaKUj8_0),.clk(gclk));
	jdff dff_A_ecvZcZ1M3_0(.dout(w_dff_A_cK3SquUy9_0),.din(w_dff_A_ecvZcZ1M3_0),.clk(gclk));
	jdff dff_A_cK3SquUy9_0(.dout(w_dff_A_AO3odD4Z5_0),.din(w_dff_A_cK3SquUy9_0),.clk(gclk));
	jdff dff_A_AO3odD4Z5_0(.dout(w_dff_A_pDZLOiEj7_0),.din(w_dff_A_AO3odD4Z5_0),.clk(gclk));
	jdff dff_A_pDZLOiEj7_0(.dout(w_dff_A_GjZBSWIH4_0),.din(w_dff_A_pDZLOiEj7_0),.clk(gclk));
	jdff dff_A_GjZBSWIH4_0(.dout(w_dff_A_Im9h7vRQ0_0),.din(w_dff_A_GjZBSWIH4_0),.clk(gclk));
	jdff dff_A_Im9h7vRQ0_0(.dout(G558),.din(w_dff_A_Im9h7vRQ0_0),.clk(gclk));
	jdff dff_A_PaiAskYr6_1(.dout(w_dff_A_PEa039RS9_0),.din(w_dff_A_PaiAskYr6_1),.clk(gclk));
	jdff dff_A_PEa039RS9_0(.dout(w_dff_A_HjVD2Ytw1_0),.din(w_dff_A_PEa039RS9_0),.clk(gclk));
	jdff dff_A_HjVD2Ytw1_0(.dout(w_dff_A_yT9STdds6_0),.din(w_dff_A_HjVD2Ytw1_0),.clk(gclk));
	jdff dff_A_yT9STdds6_0(.dout(w_dff_A_RFgEf2nd3_0),.din(w_dff_A_yT9STdds6_0),.clk(gclk));
	jdff dff_A_RFgEf2nd3_0(.dout(w_dff_A_NzQEx5ya8_0),.din(w_dff_A_RFgEf2nd3_0),.clk(gclk));
	jdff dff_A_NzQEx5ya8_0(.dout(w_dff_A_kikej6Xq9_0),.din(w_dff_A_NzQEx5ya8_0),.clk(gclk));
	jdff dff_A_kikej6Xq9_0(.dout(w_dff_A_h2d6Zx2W3_0),.din(w_dff_A_kikej6Xq9_0),.clk(gclk));
	jdff dff_A_h2d6Zx2W3_0(.dout(w_dff_A_LCDAcrbe1_0),.din(w_dff_A_h2d6Zx2W3_0),.clk(gclk));
	jdff dff_A_LCDAcrbe1_0(.dout(w_dff_A_fMLPRsZ55_0),.din(w_dff_A_LCDAcrbe1_0),.clk(gclk));
	jdff dff_A_fMLPRsZ55_0(.dout(w_dff_A_7aDMI00h7_0),.din(w_dff_A_fMLPRsZ55_0),.clk(gclk));
	jdff dff_A_7aDMI00h7_0(.dout(w_dff_A_SFh5HPZa5_0),.din(w_dff_A_7aDMI00h7_0),.clk(gclk));
	jdff dff_A_SFh5HPZa5_0(.dout(w_dff_A_Mm7RvVhS7_0),.din(w_dff_A_SFh5HPZa5_0),.clk(gclk));
	jdff dff_A_Mm7RvVhS7_0(.dout(w_dff_A_Jpov4B8I8_0),.din(w_dff_A_Mm7RvVhS7_0),.clk(gclk));
	jdff dff_A_Jpov4B8I8_0(.dout(w_dff_A_cjL4xQIG5_0),.din(w_dff_A_Jpov4B8I8_0),.clk(gclk));
	jdff dff_A_cjL4xQIG5_0(.dout(w_dff_A_PSSwYHHx5_0),.din(w_dff_A_cjL4xQIG5_0),.clk(gclk));
	jdff dff_A_PSSwYHHx5_0(.dout(w_dff_A_2oZDLeZX0_0),.din(w_dff_A_PSSwYHHx5_0),.clk(gclk));
	jdff dff_A_2oZDLeZX0_0(.dout(w_dff_A_4KsZuqwr2_0),.din(w_dff_A_2oZDLeZX0_0),.clk(gclk));
	jdff dff_A_4KsZuqwr2_0(.dout(w_dff_A_iwURB6rR4_0),.din(w_dff_A_4KsZuqwr2_0),.clk(gclk));
	jdff dff_A_iwURB6rR4_0(.dout(w_dff_A_h5hsiT301_0),.din(w_dff_A_iwURB6rR4_0),.clk(gclk));
	jdff dff_A_h5hsiT301_0(.dout(w_dff_A_EAP9Fzxq8_0),.din(w_dff_A_h5hsiT301_0),.clk(gclk));
	jdff dff_A_EAP9Fzxq8_0(.dout(w_dff_A_MTzjLy4Z3_0),.din(w_dff_A_EAP9Fzxq8_0),.clk(gclk));
	jdff dff_A_MTzjLy4Z3_0(.dout(w_dff_A_QyV2OEZm1_0),.din(w_dff_A_MTzjLy4Z3_0),.clk(gclk));
	jdff dff_A_QyV2OEZm1_0(.dout(w_dff_A_LzccGiWz1_0),.din(w_dff_A_QyV2OEZm1_0),.clk(gclk));
	jdff dff_A_LzccGiWz1_0(.dout(w_dff_A_4z79Vr0M3_0),.din(w_dff_A_LzccGiWz1_0),.clk(gclk));
	jdff dff_A_4z79Vr0M3_0(.dout(w_dff_A_Mq503fkA3_0),.din(w_dff_A_4z79Vr0M3_0),.clk(gclk));
	jdff dff_A_Mq503fkA3_0(.dout(w_dff_A_jZeqrxm32_0),.din(w_dff_A_Mq503fkA3_0),.clk(gclk));
	jdff dff_A_jZeqrxm32_0(.dout(w_dff_A_czPnHY5l5_0),.din(w_dff_A_jZeqrxm32_0),.clk(gclk));
	jdff dff_A_czPnHY5l5_0(.dout(w_dff_A_6O0aTqTv1_0),.din(w_dff_A_czPnHY5l5_0),.clk(gclk));
	jdff dff_A_6O0aTqTv1_0(.dout(w_dff_A_pjbuSGrh8_0),.din(w_dff_A_6O0aTqTv1_0),.clk(gclk));
	jdff dff_A_pjbuSGrh8_0(.dout(w_dff_A_hCIu31mj5_0),.din(w_dff_A_pjbuSGrh8_0),.clk(gclk));
	jdff dff_A_hCIu31mj5_0(.dout(w_dff_A_L8q86LG33_0),.din(w_dff_A_hCIu31mj5_0),.clk(gclk));
	jdff dff_A_L8q86LG33_0(.dout(w_dff_A_lBlhLQ2q3_0),.din(w_dff_A_L8q86LG33_0),.clk(gclk));
	jdff dff_A_lBlhLQ2q3_0(.dout(w_dff_A_7udL8dx51_0),.din(w_dff_A_lBlhLQ2q3_0),.clk(gclk));
	jdff dff_A_7udL8dx51_0(.dout(w_dff_A_UKvZ8OJJ2_0),.din(w_dff_A_7udL8dx51_0),.clk(gclk));
	jdff dff_A_UKvZ8OJJ2_0(.dout(w_dff_A_XrhJPh4c1_0),.din(w_dff_A_UKvZ8OJJ2_0),.clk(gclk));
	jdff dff_A_XrhJPh4c1_0(.dout(w_dff_A_SPebHgFh5_0),.din(w_dff_A_XrhJPh4c1_0),.clk(gclk));
	jdff dff_A_SPebHgFh5_0(.dout(w_dff_A_FWlxy7J35_0),.din(w_dff_A_SPebHgFh5_0),.clk(gclk));
	jdff dff_A_FWlxy7J35_0(.dout(G556),.din(w_dff_A_FWlxy7J35_0),.clk(gclk));
	jdff dff_A_Nu4uyITW4_1(.dout(w_dff_A_KYGZMWuo6_0),.din(w_dff_A_Nu4uyITW4_1),.clk(gclk));
	jdff dff_A_KYGZMWuo6_0(.dout(w_dff_A_V4M1shWF4_0),.din(w_dff_A_KYGZMWuo6_0),.clk(gclk));
	jdff dff_A_V4M1shWF4_0(.dout(w_dff_A_mYA8b5aI6_0),.din(w_dff_A_V4M1shWF4_0),.clk(gclk));
	jdff dff_A_mYA8b5aI6_0(.dout(w_dff_A_rOxpbbnc1_0),.din(w_dff_A_mYA8b5aI6_0),.clk(gclk));
	jdff dff_A_rOxpbbnc1_0(.dout(w_dff_A_uIPU12619_0),.din(w_dff_A_rOxpbbnc1_0),.clk(gclk));
	jdff dff_A_uIPU12619_0(.dout(w_dff_A_4uOo96oq0_0),.din(w_dff_A_uIPU12619_0),.clk(gclk));
	jdff dff_A_4uOo96oq0_0(.dout(w_dff_A_oUpgZ5rd5_0),.din(w_dff_A_4uOo96oq0_0),.clk(gclk));
	jdff dff_A_oUpgZ5rd5_0(.dout(w_dff_A_yN3MoL568_0),.din(w_dff_A_oUpgZ5rd5_0),.clk(gclk));
	jdff dff_A_yN3MoL568_0(.dout(w_dff_A_Szwxe2ap6_0),.din(w_dff_A_yN3MoL568_0),.clk(gclk));
	jdff dff_A_Szwxe2ap6_0(.dout(w_dff_A_pMU5co2v7_0),.din(w_dff_A_Szwxe2ap6_0),.clk(gclk));
	jdff dff_A_pMU5co2v7_0(.dout(w_dff_A_XbsXp4Hc6_0),.din(w_dff_A_pMU5co2v7_0),.clk(gclk));
	jdff dff_A_XbsXp4Hc6_0(.dout(w_dff_A_6zhj1UlZ9_0),.din(w_dff_A_XbsXp4Hc6_0),.clk(gclk));
	jdff dff_A_6zhj1UlZ9_0(.dout(w_dff_A_PYzorhCM0_0),.din(w_dff_A_6zhj1UlZ9_0),.clk(gclk));
	jdff dff_A_PYzorhCM0_0(.dout(w_dff_A_IpYh18977_0),.din(w_dff_A_PYzorhCM0_0),.clk(gclk));
	jdff dff_A_IpYh18977_0(.dout(w_dff_A_WJTv4oxh6_0),.din(w_dff_A_IpYh18977_0),.clk(gclk));
	jdff dff_A_WJTv4oxh6_0(.dout(w_dff_A_7zD783ES2_0),.din(w_dff_A_WJTv4oxh6_0),.clk(gclk));
	jdff dff_A_7zD783ES2_0(.dout(w_dff_A_THVfvlSd4_0),.din(w_dff_A_7zD783ES2_0),.clk(gclk));
	jdff dff_A_THVfvlSd4_0(.dout(w_dff_A_8k2dkvxx0_0),.din(w_dff_A_THVfvlSd4_0),.clk(gclk));
	jdff dff_A_8k2dkvxx0_0(.dout(w_dff_A_pVcpbkyG8_0),.din(w_dff_A_8k2dkvxx0_0),.clk(gclk));
	jdff dff_A_pVcpbkyG8_0(.dout(w_dff_A_jcA1LeCl9_0),.din(w_dff_A_pVcpbkyG8_0),.clk(gclk));
	jdff dff_A_jcA1LeCl9_0(.dout(w_dff_A_ER5x3I9I6_0),.din(w_dff_A_jcA1LeCl9_0),.clk(gclk));
	jdff dff_A_ER5x3I9I6_0(.dout(w_dff_A_cDRioxeM9_0),.din(w_dff_A_ER5x3I9I6_0),.clk(gclk));
	jdff dff_A_cDRioxeM9_0(.dout(w_dff_A_ABZ6XXaD7_0),.din(w_dff_A_cDRioxeM9_0),.clk(gclk));
	jdff dff_A_ABZ6XXaD7_0(.dout(w_dff_A_gZZUu6lb2_0),.din(w_dff_A_ABZ6XXaD7_0),.clk(gclk));
	jdff dff_A_gZZUu6lb2_0(.dout(w_dff_A_sLQNeUj59_0),.din(w_dff_A_gZZUu6lb2_0),.clk(gclk));
	jdff dff_A_sLQNeUj59_0(.dout(w_dff_A_ceg1PngX7_0),.din(w_dff_A_sLQNeUj59_0),.clk(gclk));
	jdff dff_A_ceg1PngX7_0(.dout(w_dff_A_w16ZXeoN1_0),.din(w_dff_A_ceg1PngX7_0),.clk(gclk));
	jdff dff_A_w16ZXeoN1_0(.dout(w_dff_A_oagw8f2y1_0),.din(w_dff_A_w16ZXeoN1_0),.clk(gclk));
	jdff dff_A_oagw8f2y1_0(.dout(w_dff_A_CqzgH1EY3_0),.din(w_dff_A_oagw8f2y1_0),.clk(gclk));
	jdff dff_A_CqzgH1EY3_0(.dout(w_dff_A_wrhauYB39_0),.din(w_dff_A_CqzgH1EY3_0),.clk(gclk));
	jdff dff_A_wrhauYB39_0(.dout(w_dff_A_tQKxpYIC2_0),.din(w_dff_A_wrhauYB39_0),.clk(gclk));
	jdff dff_A_tQKxpYIC2_0(.dout(w_dff_A_RzdnuyV65_0),.din(w_dff_A_tQKxpYIC2_0),.clk(gclk));
	jdff dff_A_RzdnuyV65_0(.dout(w_dff_A_aH1I6zrz7_0),.din(w_dff_A_RzdnuyV65_0),.clk(gclk));
	jdff dff_A_aH1I6zrz7_0(.dout(w_dff_A_TRsc783g3_0),.din(w_dff_A_aH1I6zrz7_0),.clk(gclk));
	jdff dff_A_TRsc783g3_0(.dout(w_dff_A_im4eF1Z26_0),.din(w_dff_A_TRsc783g3_0),.clk(gclk));
	jdff dff_A_im4eF1Z26_0(.dout(w_dff_A_jd4bV5Tj0_0),.din(w_dff_A_im4eF1Z26_0),.clk(gclk));
	jdff dff_A_jd4bV5Tj0_0(.dout(w_dff_A_JKCsMSY77_0),.din(w_dff_A_jd4bV5Tj0_0),.clk(gclk));
	jdff dff_A_JKCsMSY77_0(.dout(G554),.din(w_dff_A_JKCsMSY77_0),.clk(gclk));
	jdff dff_A_Ol3YBVCw1_1(.dout(w_dff_A_3xSYrUPJ1_0),.din(w_dff_A_Ol3YBVCw1_1),.clk(gclk));
	jdff dff_A_3xSYrUPJ1_0(.dout(w_dff_A_SUusDXpc7_0),.din(w_dff_A_3xSYrUPJ1_0),.clk(gclk));
	jdff dff_A_SUusDXpc7_0(.dout(w_dff_A_UOfqOoHs5_0),.din(w_dff_A_SUusDXpc7_0),.clk(gclk));
	jdff dff_A_UOfqOoHs5_0(.dout(w_dff_A_qsE9DeKb3_0),.din(w_dff_A_UOfqOoHs5_0),.clk(gclk));
	jdff dff_A_qsE9DeKb3_0(.dout(w_dff_A_HuUsKLXL9_0),.din(w_dff_A_qsE9DeKb3_0),.clk(gclk));
	jdff dff_A_HuUsKLXL9_0(.dout(w_dff_A_g31GadDR8_0),.din(w_dff_A_HuUsKLXL9_0),.clk(gclk));
	jdff dff_A_g31GadDR8_0(.dout(w_dff_A_FdiocZBN3_0),.din(w_dff_A_g31GadDR8_0),.clk(gclk));
	jdff dff_A_FdiocZBN3_0(.dout(w_dff_A_FMYTCX8M9_0),.din(w_dff_A_FdiocZBN3_0),.clk(gclk));
	jdff dff_A_FMYTCX8M9_0(.dout(w_dff_A_nF5Gf2cQ6_0),.din(w_dff_A_FMYTCX8M9_0),.clk(gclk));
	jdff dff_A_nF5Gf2cQ6_0(.dout(w_dff_A_55I86xLm8_0),.din(w_dff_A_nF5Gf2cQ6_0),.clk(gclk));
	jdff dff_A_55I86xLm8_0(.dout(w_dff_A_mACA9E8N1_0),.din(w_dff_A_55I86xLm8_0),.clk(gclk));
	jdff dff_A_mACA9E8N1_0(.dout(w_dff_A_V49O5pIP8_0),.din(w_dff_A_mACA9E8N1_0),.clk(gclk));
	jdff dff_A_V49O5pIP8_0(.dout(w_dff_A_9SMjUDta9_0),.din(w_dff_A_V49O5pIP8_0),.clk(gclk));
	jdff dff_A_9SMjUDta9_0(.dout(w_dff_A_a9xdFmh85_0),.din(w_dff_A_9SMjUDta9_0),.clk(gclk));
	jdff dff_A_a9xdFmh85_0(.dout(w_dff_A_9lYXErQp7_0),.din(w_dff_A_a9xdFmh85_0),.clk(gclk));
	jdff dff_A_9lYXErQp7_0(.dout(w_dff_A_C5MZFXZ75_0),.din(w_dff_A_9lYXErQp7_0),.clk(gclk));
	jdff dff_A_C5MZFXZ75_0(.dout(w_dff_A_bpCqdoll5_0),.din(w_dff_A_C5MZFXZ75_0),.clk(gclk));
	jdff dff_A_bpCqdoll5_0(.dout(w_dff_A_L4yJ4DLO0_0),.din(w_dff_A_bpCqdoll5_0),.clk(gclk));
	jdff dff_A_L4yJ4DLO0_0(.dout(w_dff_A_QPFjJrQi9_0),.din(w_dff_A_L4yJ4DLO0_0),.clk(gclk));
	jdff dff_A_QPFjJrQi9_0(.dout(w_dff_A_fEJvXimn8_0),.din(w_dff_A_QPFjJrQi9_0),.clk(gclk));
	jdff dff_A_fEJvXimn8_0(.dout(w_dff_A_5IUykv0K0_0),.din(w_dff_A_fEJvXimn8_0),.clk(gclk));
	jdff dff_A_5IUykv0K0_0(.dout(w_dff_A_VsHqff184_0),.din(w_dff_A_5IUykv0K0_0),.clk(gclk));
	jdff dff_A_VsHqff184_0(.dout(w_dff_A_0UGzpnuI2_0),.din(w_dff_A_VsHqff184_0),.clk(gclk));
	jdff dff_A_0UGzpnuI2_0(.dout(w_dff_A_zjP89fBS5_0),.din(w_dff_A_0UGzpnuI2_0),.clk(gclk));
	jdff dff_A_zjP89fBS5_0(.dout(w_dff_A_6QF1TzX20_0),.din(w_dff_A_zjP89fBS5_0),.clk(gclk));
	jdff dff_A_6QF1TzX20_0(.dout(w_dff_A_jZB9fzoP3_0),.din(w_dff_A_6QF1TzX20_0),.clk(gclk));
	jdff dff_A_jZB9fzoP3_0(.dout(w_dff_A_57zNAon70_0),.din(w_dff_A_jZB9fzoP3_0),.clk(gclk));
	jdff dff_A_57zNAon70_0(.dout(w_dff_A_bwdy6hBL9_0),.din(w_dff_A_57zNAon70_0),.clk(gclk));
	jdff dff_A_bwdy6hBL9_0(.dout(w_dff_A_MAliRglB3_0),.din(w_dff_A_bwdy6hBL9_0),.clk(gclk));
	jdff dff_A_MAliRglB3_0(.dout(w_dff_A_qiO91mHu9_0),.din(w_dff_A_MAliRglB3_0),.clk(gclk));
	jdff dff_A_qiO91mHu9_0(.dout(w_dff_A_GFjYQP9P8_0),.din(w_dff_A_qiO91mHu9_0),.clk(gclk));
	jdff dff_A_GFjYQP9P8_0(.dout(w_dff_A_8oHigkgq9_0),.din(w_dff_A_GFjYQP9P8_0),.clk(gclk));
	jdff dff_A_8oHigkgq9_0(.dout(w_dff_A_B7zQoqDe2_0),.din(w_dff_A_8oHigkgq9_0),.clk(gclk));
	jdff dff_A_B7zQoqDe2_0(.dout(w_dff_A_wk72eYIK2_0),.din(w_dff_A_B7zQoqDe2_0),.clk(gclk));
	jdff dff_A_wk72eYIK2_0(.dout(w_dff_A_C0aK5UtC3_0),.din(w_dff_A_wk72eYIK2_0),.clk(gclk));
	jdff dff_A_C0aK5UtC3_0(.dout(w_dff_A_3Ntfvrp73_0),.din(w_dff_A_C0aK5UtC3_0),.clk(gclk));
	jdff dff_A_3Ntfvrp73_0(.dout(w_dff_A_9BShlmBg5_0),.din(w_dff_A_3Ntfvrp73_0),.clk(gclk));
	jdff dff_A_9BShlmBg5_0(.dout(G552),.din(w_dff_A_9BShlmBg5_0),.clk(gclk));
	jdff dff_A_vskJrkeb7_1(.dout(w_dff_A_UXRGTtyt8_0),.din(w_dff_A_vskJrkeb7_1),.clk(gclk));
	jdff dff_A_UXRGTtyt8_0(.dout(w_dff_A_IkSHepBD2_0),.din(w_dff_A_UXRGTtyt8_0),.clk(gclk));
	jdff dff_A_IkSHepBD2_0(.dout(w_dff_A_zFEDy7cc2_0),.din(w_dff_A_IkSHepBD2_0),.clk(gclk));
	jdff dff_A_zFEDy7cc2_0(.dout(w_dff_A_rA0VUDm33_0),.din(w_dff_A_zFEDy7cc2_0),.clk(gclk));
	jdff dff_A_rA0VUDm33_0(.dout(w_dff_A_xiplURXD8_0),.din(w_dff_A_rA0VUDm33_0),.clk(gclk));
	jdff dff_A_xiplURXD8_0(.dout(w_dff_A_8mkM6KpS5_0),.din(w_dff_A_xiplURXD8_0),.clk(gclk));
	jdff dff_A_8mkM6KpS5_0(.dout(w_dff_A_PR9l0QZ11_0),.din(w_dff_A_8mkM6KpS5_0),.clk(gclk));
	jdff dff_A_PR9l0QZ11_0(.dout(w_dff_A_SEXLDF4N1_0),.din(w_dff_A_PR9l0QZ11_0),.clk(gclk));
	jdff dff_A_SEXLDF4N1_0(.dout(w_dff_A_KBiiob3w8_0),.din(w_dff_A_SEXLDF4N1_0),.clk(gclk));
	jdff dff_A_KBiiob3w8_0(.dout(w_dff_A_9WPEtNDk8_0),.din(w_dff_A_KBiiob3w8_0),.clk(gclk));
	jdff dff_A_9WPEtNDk8_0(.dout(w_dff_A_KJ3QnQ0p9_0),.din(w_dff_A_9WPEtNDk8_0),.clk(gclk));
	jdff dff_A_KJ3QnQ0p9_0(.dout(w_dff_A_lktW1RCq9_0),.din(w_dff_A_KJ3QnQ0p9_0),.clk(gclk));
	jdff dff_A_lktW1RCq9_0(.dout(w_dff_A_vqgQ8fcO2_0),.din(w_dff_A_lktW1RCq9_0),.clk(gclk));
	jdff dff_A_vqgQ8fcO2_0(.dout(w_dff_A_3gaC2I0l1_0),.din(w_dff_A_vqgQ8fcO2_0),.clk(gclk));
	jdff dff_A_3gaC2I0l1_0(.dout(w_dff_A_u4c3Jyrf9_0),.din(w_dff_A_3gaC2I0l1_0),.clk(gclk));
	jdff dff_A_u4c3Jyrf9_0(.dout(w_dff_A_e5XpNalE0_0),.din(w_dff_A_u4c3Jyrf9_0),.clk(gclk));
	jdff dff_A_e5XpNalE0_0(.dout(w_dff_A_haPEPRUE0_0),.din(w_dff_A_e5XpNalE0_0),.clk(gclk));
	jdff dff_A_haPEPRUE0_0(.dout(w_dff_A_5836id9O3_0),.din(w_dff_A_haPEPRUE0_0),.clk(gclk));
	jdff dff_A_5836id9O3_0(.dout(w_dff_A_DiVwlFmt9_0),.din(w_dff_A_5836id9O3_0),.clk(gclk));
	jdff dff_A_DiVwlFmt9_0(.dout(w_dff_A_vTIAIXSj4_0),.din(w_dff_A_DiVwlFmt9_0),.clk(gclk));
	jdff dff_A_vTIAIXSj4_0(.dout(w_dff_A_VPgE7vpf6_0),.din(w_dff_A_vTIAIXSj4_0),.clk(gclk));
	jdff dff_A_VPgE7vpf6_0(.dout(w_dff_A_AXCSkW7H8_0),.din(w_dff_A_VPgE7vpf6_0),.clk(gclk));
	jdff dff_A_AXCSkW7H8_0(.dout(w_dff_A_GQlxiqb36_0),.din(w_dff_A_AXCSkW7H8_0),.clk(gclk));
	jdff dff_A_GQlxiqb36_0(.dout(w_dff_A_fvYAw2d11_0),.din(w_dff_A_GQlxiqb36_0),.clk(gclk));
	jdff dff_A_fvYAw2d11_0(.dout(w_dff_A_fzBALfbb9_0),.din(w_dff_A_fvYAw2d11_0),.clk(gclk));
	jdff dff_A_fzBALfbb9_0(.dout(w_dff_A_z5Ba6lRk8_0),.din(w_dff_A_fzBALfbb9_0),.clk(gclk));
	jdff dff_A_z5Ba6lRk8_0(.dout(w_dff_A_RwwqTgD14_0),.din(w_dff_A_z5Ba6lRk8_0),.clk(gclk));
	jdff dff_A_RwwqTgD14_0(.dout(w_dff_A_JSUOVrrD5_0),.din(w_dff_A_RwwqTgD14_0),.clk(gclk));
	jdff dff_A_JSUOVrrD5_0(.dout(w_dff_A_P6epez6C6_0),.din(w_dff_A_JSUOVrrD5_0),.clk(gclk));
	jdff dff_A_P6epez6C6_0(.dout(w_dff_A_wp7nBcW56_0),.din(w_dff_A_P6epez6C6_0),.clk(gclk));
	jdff dff_A_wp7nBcW56_0(.dout(w_dff_A_wKKZ6bcq6_0),.din(w_dff_A_wp7nBcW56_0),.clk(gclk));
	jdff dff_A_wKKZ6bcq6_0(.dout(w_dff_A_orWLLVAh9_0),.din(w_dff_A_wKKZ6bcq6_0),.clk(gclk));
	jdff dff_A_orWLLVAh9_0(.dout(w_dff_A_oPsjac513_0),.din(w_dff_A_orWLLVAh9_0),.clk(gclk));
	jdff dff_A_oPsjac513_0(.dout(w_dff_A_onglniyU2_0),.din(w_dff_A_oPsjac513_0),.clk(gclk));
	jdff dff_A_onglniyU2_0(.dout(w_dff_A_eZ0JpgUC2_0),.din(w_dff_A_onglniyU2_0),.clk(gclk));
	jdff dff_A_eZ0JpgUC2_0(.dout(w_dff_A_ZIEpFpLb1_0),.din(w_dff_A_eZ0JpgUC2_0),.clk(gclk));
	jdff dff_A_ZIEpFpLb1_0(.dout(w_dff_A_JpkdzXt20_0),.din(w_dff_A_ZIEpFpLb1_0),.clk(gclk));
	jdff dff_A_JpkdzXt20_0(.dout(G550),.din(w_dff_A_JpkdzXt20_0),.clk(gclk));
	jdff dff_A_RaK8syet9_1(.dout(w_dff_A_Pb0FOVEH6_0),.din(w_dff_A_RaK8syet9_1),.clk(gclk));
	jdff dff_A_Pb0FOVEH6_0(.dout(w_dff_A_cNh3RjrQ9_0),.din(w_dff_A_Pb0FOVEH6_0),.clk(gclk));
	jdff dff_A_cNh3RjrQ9_0(.dout(w_dff_A_ubaG4VGD3_0),.din(w_dff_A_cNh3RjrQ9_0),.clk(gclk));
	jdff dff_A_ubaG4VGD3_0(.dout(w_dff_A_L3uNG30D4_0),.din(w_dff_A_ubaG4VGD3_0),.clk(gclk));
	jdff dff_A_L3uNG30D4_0(.dout(w_dff_A_IBFinrlo6_0),.din(w_dff_A_L3uNG30D4_0),.clk(gclk));
	jdff dff_A_IBFinrlo6_0(.dout(w_dff_A_CXm6vD924_0),.din(w_dff_A_IBFinrlo6_0),.clk(gclk));
	jdff dff_A_CXm6vD924_0(.dout(w_dff_A_Ko6wFLrb9_0),.din(w_dff_A_CXm6vD924_0),.clk(gclk));
	jdff dff_A_Ko6wFLrb9_0(.dout(w_dff_A_O95VmH619_0),.din(w_dff_A_Ko6wFLrb9_0),.clk(gclk));
	jdff dff_A_O95VmH619_0(.dout(w_dff_A_FuicjDch4_0),.din(w_dff_A_O95VmH619_0),.clk(gclk));
	jdff dff_A_FuicjDch4_0(.dout(w_dff_A_9zh2Pvub1_0),.din(w_dff_A_FuicjDch4_0),.clk(gclk));
	jdff dff_A_9zh2Pvub1_0(.dout(w_dff_A_5B7ZAKeH5_0),.din(w_dff_A_9zh2Pvub1_0),.clk(gclk));
	jdff dff_A_5B7ZAKeH5_0(.dout(w_dff_A_kyiH4Rgi2_0),.din(w_dff_A_5B7ZAKeH5_0),.clk(gclk));
	jdff dff_A_kyiH4Rgi2_0(.dout(w_dff_A_R6e2XuF09_0),.din(w_dff_A_kyiH4Rgi2_0),.clk(gclk));
	jdff dff_A_R6e2XuF09_0(.dout(w_dff_A_BaCSXDmo4_0),.din(w_dff_A_R6e2XuF09_0),.clk(gclk));
	jdff dff_A_BaCSXDmo4_0(.dout(w_dff_A_xk4RxYvX4_0),.din(w_dff_A_BaCSXDmo4_0),.clk(gclk));
	jdff dff_A_xk4RxYvX4_0(.dout(w_dff_A_LcaHG0SP1_0),.din(w_dff_A_xk4RxYvX4_0),.clk(gclk));
	jdff dff_A_LcaHG0SP1_0(.dout(w_dff_A_E7OIItkO5_0),.din(w_dff_A_LcaHG0SP1_0),.clk(gclk));
	jdff dff_A_E7OIItkO5_0(.dout(w_dff_A_TMCGoWJI1_0),.din(w_dff_A_E7OIItkO5_0),.clk(gclk));
	jdff dff_A_TMCGoWJI1_0(.dout(w_dff_A_cRBGF4Ah5_0),.din(w_dff_A_TMCGoWJI1_0),.clk(gclk));
	jdff dff_A_cRBGF4Ah5_0(.dout(w_dff_A_wAmiWsAq9_0),.din(w_dff_A_cRBGF4Ah5_0),.clk(gclk));
	jdff dff_A_wAmiWsAq9_0(.dout(w_dff_A_OPHZwJFJ1_0),.din(w_dff_A_wAmiWsAq9_0),.clk(gclk));
	jdff dff_A_OPHZwJFJ1_0(.dout(w_dff_A_2HsX3HrD8_0),.din(w_dff_A_OPHZwJFJ1_0),.clk(gclk));
	jdff dff_A_2HsX3HrD8_0(.dout(w_dff_A_y8o5wT4a7_0),.din(w_dff_A_2HsX3HrD8_0),.clk(gclk));
	jdff dff_A_y8o5wT4a7_0(.dout(w_dff_A_ocYDhLiT6_0),.din(w_dff_A_y8o5wT4a7_0),.clk(gclk));
	jdff dff_A_ocYDhLiT6_0(.dout(w_dff_A_qdlBs3d92_0),.din(w_dff_A_ocYDhLiT6_0),.clk(gclk));
	jdff dff_A_qdlBs3d92_0(.dout(w_dff_A_egPTUtCl0_0),.din(w_dff_A_qdlBs3d92_0),.clk(gclk));
	jdff dff_A_egPTUtCl0_0(.dout(w_dff_A_2qERvLwG6_0),.din(w_dff_A_egPTUtCl0_0),.clk(gclk));
	jdff dff_A_2qERvLwG6_0(.dout(w_dff_A_Rfq5qPW86_0),.din(w_dff_A_2qERvLwG6_0),.clk(gclk));
	jdff dff_A_Rfq5qPW86_0(.dout(w_dff_A_PbSay1IH1_0),.din(w_dff_A_Rfq5qPW86_0),.clk(gclk));
	jdff dff_A_PbSay1IH1_0(.dout(w_dff_A_YJjrWvDO5_0),.din(w_dff_A_PbSay1IH1_0),.clk(gclk));
	jdff dff_A_YJjrWvDO5_0(.dout(w_dff_A_ICQVzuXr5_0),.din(w_dff_A_YJjrWvDO5_0),.clk(gclk));
	jdff dff_A_ICQVzuXr5_0(.dout(w_dff_A_PjGBXlrt5_0),.din(w_dff_A_ICQVzuXr5_0),.clk(gclk));
	jdff dff_A_PjGBXlrt5_0(.dout(w_dff_A_KEQio50c4_0),.din(w_dff_A_PjGBXlrt5_0),.clk(gclk));
	jdff dff_A_KEQio50c4_0(.dout(w_dff_A_cw6n8IGT6_0),.din(w_dff_A_KEQio50c4_0),.clk(gclk));
	jdff dff_A_cw6n8IGT6_0(.dout(w_dff_A_SOWjsBFD4_0),.din(w_dff_A_cw6n8IGT6_0),.clk(gclk));
	jdff dff_A_SOWjsBFD4_0(.dout(w_dff_A_e5wWdgSw4_0),.din(w_dff_A_SOWjsBFD4_0),.clk(gclk));
	jdff dff_A_e5wWdgSw4_0(.dout(w_dff_A_kzLLaeop0_0),.din(w_dff_A_e5wWdgSw4_0),.clk(gclk));
	jdff dff_A_kzLLaeop0_0(.dout(G548),.din(w_dff_A_kzLLaeop0_0),.clk(gclk));
	jdff dff_A_rcmF46MD0_1(.dout(w_dff_A_TIKAjhuU9_0),.din(w_dff_A_rcmF46MD0_1),.clk(gclk));
	jdff dff_A_TIKAjhuU9_0(.dout(w_dff_A_ZRN1dQRs5_0),.din(w_dff_A_TIKAjhuU9_0),.clk(gclk));
	jdff dff_A_ZRN1dQRs5_0(.dout(w_dff_A_myDFnknc2_0),.din(w_dff_A_ZRN1dQRs5_0),.clk(gclk));
	jdff dff_A_myDFnknc2_0(.dout(w_dff_A_Pr60PBI84_0),.din(w_dff_A_myDFnknc2_0),.clk(gclk));
	jdff dff_A_Pr60PBI84_0(.dout(w_dff_A_v9xMhqA74_0),.din(w_dff_A_Pr60PBI84_0),.clk(gclk));
	jdff dff_A_v9xMhqA74_0(.dout(w_dff_A_sTaudX3u8_0),.din(w_dff_A_v9xMhqA74_0),.clk(gclk));
	jdff dff_A_sTaudX3u8_0(.dout(w_dff_A_WkRKEYxj7_0),.din(w_dff_A_sTaudX3u8_0),.clk(gclk));
	jdff dff_A_WkRKEYxj7_0(.dout(w_dff_A_8p3Y9tIm7_0),.din(w_dff_A_WkRKEYxj7_0),.clk(gclk));
	jdff dff_A_8p3Y9tIm7_0(.dout(w_dff_A_63qalUZc9_0),.din(w_dff_A_8p3Y9tIm7_0),.clk(gclk));
	jdff dff_A_63qalUZc9_0(.dout(w_dff_A_Y0gpKUP46_0),.din(w_dff_A_63qalUZc9_0),.clk(gclk));
	jdff dff_A_Y0gpKUP46_0(.dout(w_dff_A_Nl6H9Dbz0_0),.din(w_dff_A_Y0gpKUP46_0),.clk(gclk));
	jdff dff_A_Nl6H9Dbz0_0(.dout(w_dff_A_VBNYUmul2_0),.din(w_dff_A_Nl6H9Dbz0_0),.clk(gclk));
	jdff dff_A_VBNYUmul2_0(.dout(w_dff_A_OZfGCYwu9_0),.din(w_dff_A_VBNYUmul2_0),.clk(gclk));
	jdff dff_A_OZfGCYwu9_0(.dout(w_dff_A_cJtEl5kD8_0),.din(w_dff_A_OZfGCYwu9_0),.clk(gclk));
	jdff dff_A_cJtEl5kD8_0(.dout(w_dff_A_iEHPrY3h4_0),.din(w_dff_A_cJtEl5kD8_0),.clk(gclk));
	jdff dff_A_iEHPrY3h4_0(.dout(w_dff_A_hmaNOJpJ2_0),.din(w_dff_A_iEHPrY3h4_0),.clk(gclk));
	jdff dff_A_hmaNOJpJ2_0(.dout(w_dff_A_UPoEbzff2_0),.din(w_dff_A_hmaNOJpJ2_0),.clk(gclk));
	jdff dff_A_UPoEbzff2_0(.dout(w_dff_A_JGzFKfVt4_0),.din(w_dff_A_UPoEbzff2_0),.clk(gclk));
	jdff dff_A_JGzFKfVt4_0(.dout(w_dff_A_RAiL0qDq9_0),.din(w_dff_A_JGzFKfVt4_0),.clk(gclk));
	jdff dff_A_RAiL0qDq9_0(.dout(w_dff_A_xq0VoqIJ2_0),.din(w_dff_A_RAiL0qDq9_0),.clk(gclk));
	jdff dff_A_xq0VoqIJ2_0(.dout(w_dff_A_OyMd5xR60_0),.din(w_dff_A_xq0VoqIJ2_0),.clk(gclk));
	jdff dff_A_OyMd5xR60_0(.dout(w_dff_A_JmEGPCpi9_0),.din(w_dff_A_OyMd5xR60_0),.clk(gclk));
	jdff dff_A_JmEGPCpi9_0(.dout(w_dff_A_gJSuG6s35_0),.din(w_dff_A_JmEGPCpi9_0),.clk(gclk));
	jdff dff_A_gJSuG6s35_0(.dout(w_dff_A_ARddEvWE7_0),.din(w_dff_A_gJSuG6s35_0),.clk(gclk));
	jdff dff_A_ARddEvWE7_0(.dout(w_dff_A_DbDzDBwI0_0),.din(w_dff_A_ARddEvWE7_0),.clk(gclk));
	jdff dff_A_DbDzDBwI0_0(.dout(w_dff_A_Lupy8mqA7_0),.din(w_dff_A_DbDzDBwI0_0),.clk(gclk));
	jdff dff_A_Lupy8mqA7_0(.dout(w_dff_A_0VTU5TVu6_0),.din(w_dff_A_Lupy8mqA7_0),.clk(gclk));
	jdff dff_A_0VTU5TVu6_0(.dout(w_dff_A_SDITtrK46_0),.din(w_dff_A_0VTU5TVu6_0),.clk(gclk));
	jdff dff_A_SDITtrK46_0(.dout(w_dff_A_FVF7AGru3_0),.din(w_dff_A_SDITtrK46_0),.clk(gclk));
	jdff dff_A_FVF7AGru3_0(.dout(w_dff_A_ICynjAzX7_0),.din(w_dff_A_FVF7AGru3_0),.clk(gclk));
	jdff dff_A_ICynjAzX7_0(.dout(w_dff_A_66klPyMA8_0),.din(w_dff_A_ICynjAzX7_0),.clk(gclk));
	jdff dff_A_66klPyMA8_0(.dout(w_dff_A_V3PxxPoI9_0),.din(w_dff_A_66klPyMA8_0),.clk(gclk));
	jdff dff_A_V3PxxPoI9_0(.dout(w_dff_A_1cnWBF4V9_0),.din(w_dff_A_V3PxxPoI9_0),.clk(gclk));
	jdff dff_A_1cnWBF4V9_0(.dout(w_dff_A_ycaRZFlL9_0),.din(w_dff_A_1cnWBF4V9_0),.clk(gclk));
	jdff dff_A_ycaRZFlL9_0(.dout(w_dff_A_pbDOYEnG0_0),.din(w_dff_A_ycaRZFlL9_0),.clk(gclk));
	jdff dff_A_pbDOYEnG0_0(.dout(w_dff_A_bX0Ptm3l1_0),.din(w_dff_A_pbDOYEnG0_0),.clk(gclk));
	jdff dff_A_bX0Ptm3l1_0(.dout(w_dff_A_ObZeEgSA1_0),.din(w_dff_A_bX0Ptm3l1_0),.clk(gclk));
	jdff dff_A_ObZeEgSA1_0(.dout(G546),.din(w_dff_A_ObZeEgSA1_0),.clk(gclk));
	jdff dff_A_dxxPtiY89_1(.dout(w_dff_A_G97i5TXp7_0),.din(w_dff_A_dxxPtiY89_1),.clk(gclk));
	jdff dff_A_G97i5TXp7_0(.dout(w_dff_A_VHRF8OEO2_0),.din(w_dff_A_G97i5TXp7_0),.clk(gclk));
	jdff dff_A_VHRF8OEO2_0(.dout(w_dff_A_I3eEu5BT4_0),.din(w_dff_A_VHRF8OEO2_0),.clk(gclk));
	jdff dff_A_I3eEu5BT4_0(.dout(w_dff_A_0ANP60F64_0),.din(w_dff_A_I3eEu5BT4_0),.clk(gclk));
	jdff dff_A_0ANP60F64_0(.dout(w_dff_A_PmBYg4Oq2_0),.din(w_dff_A_0ANP60F64_0),.clk(gclk));
	jdff dff_A_PmBYg4Oq2_0(.dout(w_dff_A_XfqgMaMf9_0),.din(w_dff_A_PmBYg4Oq2_0),.clk(gclk));
	jdff dff_A_XfqgMaMf9_0(.dout(w_dff_A_QdgbZmrm1_0),.din(w_dff_A_XfqgMaMf9_0),.clk(gclk));
	jdff dff_A_QdgbZmrm1_0(.dout(w_dff_A_b1Dk2QaW7_0),.din(w_dff_A_QdgbZmrm1_0),.clk(gclk));
	jdff dff_A_b1Dk2QaW7_0(.dout(w_dff_A_yuhXJrgn8_0),.din(w_dff_A_b1Dk2QaW7_0),.clk(gclk));
	jdff dff_A_yuhXJrgn8_0(.dout(w_dff_A_wxgERnc01_0),.din(w_dff_A_yuhXJrgn8_0),.clk(gclk));
	jdff dff_A_wxgERnc01_0(.dout(w_dff_A_T692Kb5M9_0),.din(w_dff_A_wxgERnc01_0),.clk(gclk));
	jdff dff_A_T692Kb5M9_0(.dout(w_dff_A_E21QNLKS4_0),.din(w_dff_A_T692Kb5M9_0),.clk(gclk));
	jdff dff_A_E21QNLKS4_0(.dout(w_dff_A_W4iO5Nsn4_0),.din(w_dff_A_E21QNLKS4_0),.clk(gclk));
	jdff dff_A_W4iO5Nsn4_0(.dout(w_dff_A_eGycNfi15_0),.din(w_dff_A_W4iO5Nsn4_0),.clk(gclk));
	jdff dff_A_eGycNfi15_0(.dout(w_dff_A_nW0dzScY3_0),.din(w_dff_A_eGycNfi15_0),.clk(gclk));
	jdff dff_A_nW0dzScY3_0(.dout(w_dff_A_Outscrxx1_0),.din(w_dff_A_nW0dzScY3_0),.clk(gclk));
	jdff dff_A_Outscrxx1_0(.dout(w_dff_A_VMIh675L0_0),.din(w_dff_A_Outscrxx1_0),.clk(gclk));
	jdff dff_A_VMIh675L0_0(.dout(w_dff_A_ORckzife0_0),.din(w_dff_A_VMIh675L0_0),.clk(gclk));
	jdff dff_A_ORckzife0_0(.dout(w_dff_A_uxMBtKj98_0),.din(w_dff_A_ORckzife0_0),.clk(gclk));
	jdff dff_A_uxMBtKj98_0(.dout(w_dff_A_EvTsR43w5_0),.din(w_dff_A_uxMBtKj98_0),.clk(gclk));
	jdff dff_A_EvTsR43w5_0(.dout(w_dff_A_POHudtj46_0),.din(w_dff_A_EvTsR43w5_0),.clk(gclk));
	jdff dff_A_POHudtj46_0(.dout(w_dff_A_Cn5eg88Q0_0),.din(w_dff_A_POHudtj46_0),.clk(gclk));
	jdff dff_A_Cn5eg88Q0_0(.dout(w_dff_A_kCv8v0yV1_0),.din(w_dff_A_Cn5eg88Q0_0),.clk(gclk));
	jdff dff_A_kCv8v0yV1_0(.dout(w_dff_A_BkYbtoU89_0),.din(w_dff_A_kCv8v0yV1_0),.clk(gclk));
	jdff dff_A_BkYbtoU89_0(.dout(w_dff_A_2s01hytV1_0),.din(w_dff_A_BkYbtoU89_0),.clk(gclk));
	jdff dff_A_2s01hytV1_0(.dout(w_dff_A_x0MQOnZ92_0),.din(w_dff_A_2s01hytV1_0),.clk(gclk));
	jdff dff_A_x0MQOnZ92_0(.dout(w_dff_A_YFmCDhea8_0),.din(w_dff_A_x0MQOnZ92_0),.clk(gclk));
	jdff dff_A_YFmCDhea8_0(.dout(w_dff_A_JE7Bxocw3_0),.din(w_dff_A_YFmCDhea8_0),.clk(gclk));
	jdff dff_A_JE7Bxocw3_0(.dout(w_dff_A_MSq3OtVs5_0),.din(w_dff_A_JE7Bxocw3_0),.clk(gclk));
	jdff dff_A_MSq3OtVs5_0(.dout(w_dff_A_LVicT9iL1_0),.din(w_dff_A_MSq3OtVs5_0),.clk(gclk));
	jdff dff_A_LVicT9iL1_0(.dout(w_dff_A_yykhCNPr0_0),.din(w_dff_A_LVicT9iL1_0),.clk(gclk));
	jdff dff_A_yykhCNPr0_0(.dout(w_dff_A_kbhJRXdQ6_0),.din(w_dff_A_yykhCNPr0_0),.clk(gclk));
	jdff dff_A_kbhJRXdQ6_0(.dout(w_dff_A_2tqiUYdu1_0),.din(w_dff_A_kbhJRXdQ6_0),.clk(gclk));
	jdff dff_A_2tqiUYdu1_0(.dout(w_dff_A_DKAYhMC89_0),.din(w_dff_A_2tqiUYdu1_0),.clk(gclk));
	jdff dff_A_DKAYhMC89_0(.dout(w_dff_A_bjHWOuXD7_0),.din(w_dff_A_DKAYhMC89_0),.clk(gclk));
	jdff dff_A_bjHWOuXD7_0(.dout(w_dff_A_RDsF7P6a8_0),.din(w_dff_A_bjHWOuXD7_0),.clk(gclk));
	jdff dff_A_RDsF7P6a8_0(.dout(w_dff_A_QYJkjfVl0_0),.din(w_dff_A_RDsF7P6a8_0),.clk(gclk));
	jdff dff_A_QYJkjfVl0_0(.dout(G544),.din(w_dff_A_QYJkjfVl0_0),.clk(gclk));
	jdff dff_A_k9lEreo95_1(.dout(w_dff_A_0nwAKcp88_0),.din(w_dff_A_k9lEreo95_1),.clk(gclk));
	jdff dff_A_0nwAKcp88_0(.dout(w_dff_A_jGNhNoDc3_0),.din(w_dff_A_0nwAKcp88_0),.clk(gclk));
	jdff dff_A_jGNhNoDc3_0(.dout(w_dff_A_ejCxPrz08_0),.din(w_dff_A_jGNhNoDc3_0),.clk(gclk));
	jdff dff_A_ejCxPrz08_0(.dout(w_dff_A_w4MTPZZ84_0),.din(w_dff_A_ejCxPrz08_0),.clk(gclk));
	jdff dff_A_w4MTPZZ84_0(.dout(w_dff_A_Sgf2csNq0_0),.din(w_dff_A_w4MTPZZ84_0),.clk(gclk));
	jdff dff_A_Sgf2csNq0_0(.dout(w_dff_A_8cjCODhm6_0),.din(w_dff_A_Sgf2csNq0_0),.clk(gclk));
	jdff dff_A_8cjCODhm6_0(.dout(w_dff_A_DreVlXB93_0),.din(w_dff_A_8cjCODhm6_0),.clk(gclk));
	jdff dff_A_DreVlXB93_0(.dout(w_dff_A_QvaNNxVW7_0),.din(w_dff_A_DreVlXB93_0),.clk(gclk));
	jdff dff_A_QvaNNxVW7_0(.dout(w_dff_A_Eae8EmhX1_0),.din(w_dff_A_QvaNNxVW7_0),.clk(gclk));
	jdff dff_A_Eae8EmhX1_0(.dout(w_dff_A_KDUKBNT96_0),.din(w_dff_A_Eae8EmhX1_0),.clk(gclk));
	jdff dff_A_KDUKBNT96_0(.dout(w_dff_A_CJS2jRgH4_0),.din(w_dff_A_KDUKBNT96_0),.clk(gclk));
	jdff dff_A_CJS2jRgH4_0(.dout(w_dff_A_0pg6gr2N2_0),.din(w_dff_A_CJS2jRgH4_0),.clk(gclk));
	jdff dff_A_0pg6gr2N2_0(.dout(w_dff_A_rUgAKxQk2_0),.din(w_dff_A_0pg6gr2N2_0),.clk(gclk));
	jdff dff_A_rUgAKxQk2_0(.dout(w_dff_A_F62ckR6d5_0),.din(w_dff_A_rUgAKxQk2_0),.clk(gclk));
	jdff dff_A_F62ckR6d5_0(.dout(w_dff_A_hqze5srK4_0),.din(w_dff_A_F62ckR6d5_0),.clk(gclk));
	jdff dff_A_hqze5srK4_0(.dout(w_dff_A_DYinpXFB0_0),.din(w_dff_A_hqze5srK4_0),.clk(gclk));
	jdff dff_A_DYinpXFB0_0(.dout(w_dff_A_USTYARax8_0),.din(w_dff_A_DYinpXFB0_0),.clk(gclk));
	jdff dff_A_USTYARax8_0(.dout(w_dff_A_weaCHrdm0_0),.din(w_dff_A_USTYARax8_0),.clk(gclk));
	jdff dff_A_weaCHrdm0_0(.dout(w_dff_A_lIvf3hr91_0),.din(w_dff_A_weaCHrdm0_0),.clk(gclk));
	jdff dff_A_lIvf3hr91_0(.dout(w_dff_A_uy2MvhMz9_0),.din(w_dff_A_lIvf3hr91_0),.clk(gclk));
	jdff dff_A_uy2MvhMz9_0(.dout(w_dff_A_4Non3de70_0),.din(w_dff_A_uy2MvhMz9_0),.clk(gclk));
	jdff dff_A_4Non3de70_0(.dout(w_dff_A_MPeLjYBn4_0),.din(w_dff_A_4Non3de70_0),.clk(gclk));
	jdff dff_A_MPeLjYBn4_0(.dout(w_dff_A_VpYkl1ja7_0),.din(w_dff_A_MPeLjYBn4_0),.clk(gclk));
	jdff dff_A_VpYkl1ja7_0(.dout(w_dff_A_uRS1m2v22_0),.din(w_dff_A_VpYkl1ja7_0),.clk(gclk));
	jdff dff_A_uRS1m2v22_0(.dout(w_dff_A_dcCxrZNW1_0),.din(w_dff_A_uRS1m2v22_0),.clk(gclk));
	jdff dff_A_dcCxrZNW1_0(.dout(w_dff_A_Zx2B5KrL4_0),.din(w_dff_A_dcCxrZNW1_0),.clk(gclk));
	jdff dff_A_Zx2B5KrL4_0(.dout(w_dff_A_qJJSCMbZ0_0),.din(w_dff_A_Zx2B5KrL4_0),.clk(gclk));
	jdff dff_A_qJJSCMbZ0_0(.dout(w_dff_A_XFyMPW0X9_0),.din(w_dff_A_qJJSCMbZ0_0),.clk(gclk));
	jdff dff_A_XFyMPW0X9_0(.dout(w_dff_A_B7epnpWG3_0),.din(w_dff_A_XFyMPW0X9_0),.clk(gclk));
	jdff dff_A_B7epnpWG3_0(.dout(w_dff_A_JUZHmBjy2_0),.din(w_dff_A_B7epnpWG3_0),.clk(gclk));
	jdff dff_A_JUZHmBjy2_0(.dout(w_dff_A_VXZs3TAF0_0),.din(w_dff_A_JUZHmBjy2_0),.clk(gclk));
	jdff dff_A_VXZs3TAF0_0(.dout(w_dff_A_MAqTSXBt9_0),.din(w_dff_A_VXZs3TAF0_0),.clk(gclk));
	jdff dff_A_MAqTSXBt9_0(.dout(w_dff_A_QOjK9iD20_0),.din(w_dff_A_MAqTSXBt9_0),.clk(gclk));
	jdff dff_A_QOjK9iD20_0(.dout(w_dff_A_U2EDWbT94_0),.din(w_dff_A_QOjK9iD20_0),.clk(gclk));
	jdff dff_A_U2EDWbT94_0(.dout(w_dff_A_KkTw2BSX2_0),.din(w_dff_A_U2EDWbT94_0),.clk(gclk));
	jdff dff_A_KkTw2BSX2_0(.dout(w_dff_A_CP1kEolh0_0),.din(w_dff_A_KkTw2BSX2_0),.clk(gclk));
	jdff dff_A_CP1kEolh0_0(.dout(w_dff_A_19ElGh7A7_0),.din(w_dff_A_CP1kEolh0_0),.clk(gclk));
	jdff dff_A_19ElGh7A7_0(.dout(G540),.din(w_dff_A_19ElGh7A7_0),.clk(gclk));
	jdff dff_A_OvoAegEm6_1(.dout(w_dff_A_ydkyoe2X6_0),.din(w_dff_A_OvoAegEm6_1),.clk(gclk));
	jdff dff_A_ydkyoe2X6_0(.dout(w_dff_A_wh0eUoIo5_0),.din(w_dff_A_ydkyoe2X6_0),.clk(gclk));
	jdff dff_A_wh0eUoIo5_0(.dout(w_dff_A_7d98hpyX4_0),.din(w_dff_A_wh0eUoIo5_0),.clk(gclk));
	jdff dff_A_7d98hpyX4_0(.dout(w_dff_A_rgZN6Zkb7_0),.din(w_dff_A_7d98hpyX4_0),.clk(gclk));
	jdff dff_A_rgZN6Zkb7_0(.dout(w_dff_A_xVug889p9_0),.din(w_dff_A_rgZN6Zkb7_0),.clk(gclk));
	jdff dff_A_xVug889p9_0(.dout(w_dff_A_ZZBzL6wA1_0),.din(w_dff_A_xVug889p9_0),.clk(gclk));
	jdff dff_A_ZZBzL6wA1_0(.dout(w_dff_A_GpDI3p6U6_0),.din(w_dff_A_ZZBzL6wA1_0),.clk(gclk));
	jdff dff_A_GpDI3p6U6_0(.dout(w_dff_A_aVuUX56V4_0),.din(w_dff_A_GpDI3p6U6_0),.clk(gclk));
	jdff dff_A_aVuUX56V4_0(.dout(w_dff_A_qwj7MtCH2_0),.din(w_dff_A_aVuUX56V4_0),.clk(gclk));
	jdff dff_A_qwj7MtCH2_0(.dout(w_dff_A_X6n74ntP7_0),.din(w_dff_A_qwj7MtCH2_0),.clk(gclk));
	jdff dff_A_X6n74ntP7_0(.dout(w_dff_A_M2xpWZOp0_0),.din(w_dff_A_X6n74ntP7_0),.clk(gclk));
	jdff dff_A_M2xpWZOp0_0(.dout(w_dff_A_KrfvbOPY0_0),.din(w_dff_A_M2xpWZOp0_0),.clk(gclk));
	jdff dff_A_KrfvbOPY0_0(.dout(w_dff_A_mZ4nhya30_0),.din(w_dff_A_KrfvbOPY0_0),.clk(gclk));
	jdff dff_A_mZ4nhya30_0(.dout(w_dff_A_KhIoE2iT8_0),.din(w_dff_A_mZ4nhya30_0),.clk(gclk));
	jdff dff_A_KhIoE2iT8_0(.dout(w_dff_A_Ujr24iPF8_0),.din(w_dff_A_KhIoE2iT8_0),.clk(gclk));
	jdff dff_A_Ujr24iPF8_0(.dout(w_dff_A_B8fAShn17_0),.din(w_dff_A_Ujr24iPF8_0),.clk(gclk));
	jdff dff_A_B8fAShn17_0(.dout(w_dff_A_Ih6dd4rl0_0),.din(w_dff_A_B8fAShn17_0),.clk(gclk));
	jdff dff_A_Ih6dd4rl0_0(.dout(w_dff_A_raRKZkES9_0),.din(w_dff_A_Ih6dd4rl0_0),.clk(gclk));
	jdff dff_A_raRKZkES9_0(.dout(w_dff_A_yIUv6Glp2_0),.din(w_dff_A_raRKZkES9_0),.clk(gclk));
	jdff dff_A_yIUv6Glp2_0(.dout(w_dff_A_NWV0efjI5_0),.din(w_dff_A_yIUv6Glp2_0),.clk(gclk));
	jdff dff_A_NWV0efjI5_0(.dout(w_dff_A_5vsPEcrY6_0),.din(w_dff_A_NWV0efjI5_0),.clk(gclk));
	jdff dff_A_5vsPEcrY6_0(.dout(w_dff_A_yuhaGSUP4_0),.din(w_dff_A_5vsPEcrY6_0),.clk(gclk));
	jdff dff_A_yuhaGSUP4_0(.dout(w_dff_A_WbIpVahl1_0),.din(w_dff_A_yuhaGSUP4_0),.clk(gclk));
	jdff dff_A_WbIpVahl1_0(.dout(w_dff_A_5nQjm3KJ8_0),.din(w_dff_A_WbIpVahl1_0),.clk(gclk));
	jdff dff_A_5nQjm3KJ8_0(.dout(w_dff_A_mbRarS1g5_0),.din(w_dff_A_5nQjm3KJ8_0),.clk(gclk));
	jdff dff_A_mbRarS1g5_0(.dout(w_dff_A_N5QgfnDu5_0),.din(w_dff_A_mbRarS1g5_0),.clk(gclk));
	jdff dff_A_N5QgfnDu5_0(.dout(w_dff_A_Pb2yFNHE9_0),.din(w_dff_A_N5QgfnDu5_0),.clk(gclk));
	jdff dff_A_Pb2yFNHE9_0(.dout(w_dff_A_Czc2e6Vp5_0),.din(w_dff_A_Pb2yFNHE9_0),.clk(gclk));
	jdff dff_A_Czc2e6Vp5_0(.dout(w_dff_A_hKmT7x8c4_0),.din(w_dff_A_Czc2e6Vp5_0),.clk(gclk));
	jdff dff_A_hKmT7x8c4_0(.dout(w_dff_A_DDidJ2n95_0),.din(w_dff_A_hKmT7x8c4_0),.clk(gclk));
	jdff dff_A_DDidJ2n95_0(.dout(w_dff_A_I59aTpTO1_0),.din(w_dff_A_DDidJ2n95_0),.clk(gclk));
	jdff dff_A_I59aTpTO1_0(.dout(w_dff_A_18OEmnbb0_0),.din(w_dff_A_I59aTpTO1_0),.clk(gclk));
	jdff dff_A_18OEmnbb0_0(.dout(w_dff_A_L3RXcbDh0_0),.din(w_dff_A_18OEmnbb0_0),.clk(gclk));
	jdff dff_A_L3RXcbDh0_0(.dout(w_dff_A_4I5IVXMF3_0),.din(w_dff_A_L3RXcbDh0_0),.clk(gclk));
	jdff dff_A_4I5IVXMF3_0(.dout(w_dff_A_EWOwMrOK0_0),.din(w_dff_A_4I5IVXMF3_0),.clk(gclk));
	jdff dff_A_EWOwMrOK0_0(.dout(w_dff_A_0VpkrRIy8_0),.din(w_dff_A_EWOwMrOK0_0),.clk(gclk));
	jdff dff_A_0VpkrRIy8_0(.dout(w_dff_A_y10T6j0N4_0),.din(w_dff_A_0VpkrRIy8_0),.clk(gclk));
	jdff dff_A_y10T6j0N4_0(.dout(G538),.din(w_dff_A_y10T6j0N4_0),.clk(gclk));
	jdff dff_A_tWFx69fK7_1(.dout(w_dff_A_rBXTNuUt5_0),.din(w_dff_A_tWFx69fK7_1),.clk(gclk));
	jdff dff_A_rBXTNuUt5_0(.dout(w_dff_A_o1iutIEO7_0),.din(w_dff_A_rBXTNuUt5_0),.clk(gclk));
	jdff dff_A_o1iutIEO7_0(.dout(w_dff_A_gOWLBNeg9_0),.din(w_dff_A_o1iutIEO7_0),.clk(gclk));
	jdff dff_A_gOWLBNeg9_0(.dout(w_dff_A_UGtPa2xC2_0),.din(w_dff_A_gOWLBNeg9_0),.clk(gclk));
	jdff dff_A_UGtPa2xC2_0(.dout(w_dff_A_nNwuuTzu5_0),.din(w_dff_A_UGtPa2xC2_0),.clk(gclk));
	jdff dff_A_nNwuuTzu5_0(.dout(w_dff_A_cqqhmPMK6_0),.din(w_dff_A_nNwuuTzu5_0),.clk(gclk));
	jdff dff_A_cqqhmPMK6_0(.dout(w_dff_A_ikMW08vh6_0),.din(w_dff_A_cqqhmPMK6_0),.clk(gclk));
	jdff dff_A_ikMW08vh6_0(.dout(w_dff_A_RU6Ktixm8_0),.din(w_dff_A_ikMW08vh6_0),.clk(gclk));
	jdff dff_A_RU6Ktixm8_0(.dout(w_dff_A_RlfKC6hj9_0),.din(w_dff_A_RU6Ktixm8_0),.clk(gclk));
	jdff dff_A_RlfKC6hj9_0(.dout(w_dff_A_fNk6dXlS5_0),.din(w_dff_A_RlfKC6hj9_0),.clk(gclk));
	jdff dff_A_fNk6dXlS5_0(.dout(w_dff_A_EYhkACvk6_0),.din(w_dff_A_fNk6dXlS5_0),.clk(gclk));
	jdff dff_A_EYhkACvk6_0(.dout(w_dff_A_KdJX0QZ25_0),.din(w_dff_A_EYhkACvk6_0),.clk(gclk));
	jdff dff_A_KdJX0QZ25_0(.dout(w_dff_A_TV58zjAa9_0),.din(w_dff_A_KdJX0QZ25_0),.clk(gclk));
	jdff dff_A_TV58zjAa9_0(.dout(w_dff_A_zBTMu70L5_0),.din(w_dff_A_TV58zjAa9_0),.clk(gclk));
	jdff dff_A_zBTMu70L5_0(.dout(w_dff_A_EsETY64J9_0),.din(w_dff_A_zBTMu70L5_0),.clk(gclk));
	jdff dff_A_EsETY64J9_0(.dout(w_dff_A_xvGjPyfh0_0),.din(w_dff_A_EsETY64J9_0),.clk(gclk));
	jdff dff_A_xvGjPyfh0_0(.dout(w_dff_A_65jCh6314_0),.din(w_dff_A_xvGjPyfh0_0),.clk(gclk));
	jdff dff_A_65jCh6314_0(.dout(w_dff_A_yY971RDm1_0),.din(w_dff_A_65jCh6314_0),.clk(gclk));
	jdff dff_A_yY971RDm1_0(.dout(w_dff_A_wcM56EJB3_0),.din(w_dff_A_yY971RDm1_0),.clk(gclk));
	jdff dff_A_wcM56EJB3_0(.dout(w_dff_A_tFAjRxPB6_0),.din(w_dff_A_wcM56EJB3_0),.clk(gclk));
	jdff dff_A_tFAjRxPB6_0(.dout(w_dff_A_QHXXRhc95_0),.din(w_dff_A_tFAjRxPB6_0),.clk(gclk));
	jdff dff_A_QHXXRhc95_0(.dout(w_dff_A_FzEdkxbu0_0),.din(w_dff_A_QHXXRhc95_0),.clk(gclk));
	jdff dff_A_FzEdkxbu0_0(.dout(w_dff_A_dmwX4KAX6_0),.din(w_dff_A_FzEdkxbu0_0),.clk(gclk));
	jdff dff_A_dmwX4KAX6_0(.dout(w_dff_A_LZUxxINK8_0),.din(w_dff_A_dmwX4KAX6_0),.clk(gclk));
	jdff dff_A_LZUxxINK8_0(.dout(w_dff_A_XqCnE4RS6_0),.din(w_dff_A_LZUxxINK8_0),.clk(gclk));
	jdff dff_A_XqCnE4RS6_0(.dout(w_dff_A_234JKLKH4_0),.din(w_dff_A_XqCnE4RS6_0),.clk(gclk));
	jdff dff_A_234JKLKH4_0(.dout(w_dff_A_g1iWwlxg0_0),.din(w_dff_A_234JKLKH4_0),.clk(gclk));
	jdff dff_A_g1iWwlxg0_0(.dout(w_dff_A_OyIrr8827_0),.din(w_dff_A_g1iWwlxg0_0),.clk(gclk));
	jdff dff_A_OyIrr8827_0(.dout(w_dff_A_6vm2bBBs2_0),.din(w_dff_A_OyIrr8827_0),.clk(gclk));
	jdff dff_A_6vm2bBBs2_0(.dout(w_dff_A_W5AHB6tU7_0),.din(w_dff_A_6vm2bBBs2_0),.clk(gclk));
	jdff dff_A_W5AHB6tU7_0(.dout(w_dff_A_dQ0E8VZA2_0),.din(w_dff_A_W5AHB6tU7_0),.clk(gclk));
	jdff dff_A_dQ0E8VZA2_0(.dout(w_dff_A_OTO4CLrO6_0),.din(w_dff_A_dQ0E8VZA2_0),.clk(gclk));
	jdff dff_A_OTO4CLrO6_0(.dout(w_dff_A_hBNXpWWr1_0),.din(w_dff_A_OTO4CLrO6_0),.clk(gclk));
	jdff dff_A_hBNXpWWr1_0(.dout(w_dff_A_k2jTy2Qw9_0),.din(w_dff_A_hBNXpWWr1_0),.clk(gclk));
	jdff dff_A_k2jTy2Qw9_0(.dout(w_dff_A_JtbBrwXu8_0),.din(w_dff_A_k2jTy2Qw9_0),.clk(gclk));
	jdff dff_A_JtbBrwXu8_0(.dout(w_dff_A_PxN5ufQQ4_0),.din(w_dff_A_JtbBrwXu8_0),.clk(gclk));
	jdff dff_A_PxN5ufQQ4_0(.dout(w_dff_A_IRFD80KQ9_0),.din(w_dff_A_PxN5ufQQ4_0),.clk(gclk));
	jdff dff_A_IRFD80KQ9_0(.dout(G536),.din(w_dff_A_IRFD80KQ9_0),.clk(gclk));
	jdff dff_A_WpSOD8rp3_1(.dout(w_dff_A_CdT4sQSo2_0),.din(w_dff_A_WpSOD8rp3_1),.clk(gclk));
	jdff dff_A_CdT4sQSo2_0(.dout(w_dff_A_HMHE3DiA7_0),.din(w_dff_A_CdT4sQSo2_0),.clk(gclk));
	jdff dff_A_HMHE3DiA7_0(.dout(w_dff_A_x67nYRTP7_0),.din(w_dff_A_HMHE3DiA7_0),.clk(gclk));
	jdff dff_A_x67nYRTP7_0(.dout(w_dff_A_mcfY7cTk4_0),.din(w_dff_A_x67nYRTP7_0),.clk(gclk));
	jdff dff_A_mcfY7cTk4_0(.dout(w_dff_A_fSiYOQJI0_0),.din(w_dff_A_mcfY7cTk4_0),.clk(gclk));
	jdff dff_A_fSiYOQJI0_0(.dout(w_dff_A_38EpSSyU5_0),.din(w_dff_A_fSiYOQJI0_0),.clk(gclk));
	jdff dff_A_38EpSSyU5_0(.dout(w_dff_A_g6CO0Dzi9_0),.din(w_dff_A_38EpSSyU5_0),.clk(gclk));
	jdff dff_A_g6CO0Dzi9_0(.dout(w_dff_A_00OqCLVW3_0),.din(w_dff_A_g6CO0Dzi9_0),.clk(gclk));
	jdff dff_A_00OqCLVW3_0(.dout(w_dff_A_TsAWrXEj4_0),.din(w_dff_A_00OqCLVW3_0),.clk(gclk));
	jdff dff_A_TsAWrXEj4_0(.dout(w_dff_A_IlTOizfN3_0),.din(w_dff_A_TsAWrXEj4_0),.clk(gclk));
	jdff dff_A_IlTOizfN3_0(.dout(w_dff_A_RISActYd1_0),.din(w_dff_A_IlTOizfN3_0),.clk(gclk));
	jdff dff_A_RISActYd1_0(.dout(w_dff_A_H5j4OuP52_0),.din(w_dff_A_RISActYd1_0),.clk(gclk));
	jdff dff_A_H5j4OuP52_0(.dout(w_dff_A_adGiQ2RC5_0),.din(w_dff_A_H5j4OuP52_0),.clk(gclk));
	jdff dff_A_adGiQ2RC5_0(.dout(w_dff_A_FiyPuiCJ2_0),.din(w_dff_A_adGiQ2RC5_0),.clk(gclk));
	jdff dff_A_FiyPuiCJ2_0(.dout(w_dff_A_XFCBeme97_0),.din(w_dff_A_FiyPuiCJ2_0),.clk(gclk));
	jdff dff_A_XFCBeme97_0(.dout(w_dff_A_CkcwRHEs5_0),.din(w_dff_A_XFCBeme97_0),.clk(gclk));
	jdff dff_A_CkcwRHEs5_0(.dout(w_dff_A_Tv2cXZev3_0),.din(w_dff_A_CkcwRHEs5_0),.clk(gclk));
	jdff dff_A_Tv2cXZev3_0(.dout(w_dff_A_J507qUcA2_0),.din(w_dff_A_Tv2cXZev3_0),.clk(gclk));
	jdff dff_A_J507qUcA2_0(.dout(w_dff_A_MEHbksYP3_0),.din(w_dff_A_J507qUcA2_0),.clk(gclk));
	jdff dff_A_MEHbksYP3_0(.dout(w_dff_A_GjJV2pwR2_0),.din(w_dff_A_MEHbksYP3_0),.clk(gclk));
	jdff dff_A_GjJV2pwR2_0(.dout(w_dff_A_a93uWquw8_0),.din(w_dff_A_GjJV2pwR2_0),.clk(gclk));
	jdff dff_A_a93uWquw8_0(.dout(w_dff_A_eYCmwouk4_0),.din(w_dff_A_a93uWquw8_0),.clk(gclk));
	jdff dff_A_eYCmwouk4_0(.dout(w_dff_A_AFiznRLh2_0),.din(w_dff_A_eYCmwouk4_0),.clk(gclk));
	jdff dff_A_AFiznRLh2_0(.dout(w_dff_A_h5VXymDw1_0),.din(w_dff_A_AFiznRLh2_0),.clk(gclk));
	jdff dff_A_h5VXymDw1_0(.dout(w_dff_A_TZ63m7H05_0),.din(w_dff_A_h5VXymDw1_0),.clk(gclk));
	jdff dff_A_TZ63m7H05_0(.dout(w_dff_A_hrfWgdWW8_0),.din(w_dff_A_TZ63m7H05_0),.clk(gclk));
	jdff dff_A_hrfWgdWW8_0(.dout(w_dff_A_UgHRdBhH4_0),.din(w_dff_A_hrfWgdWW8_0),.clk(gclk));
	jdff dff_A_UgHRdBhH4_0(.dout(w_dff_A_B6M3UwiU8_0),.din(w_dff_A_UgHRdBhH4_0),.clk(gclk));
	jdff dff_A_B6M3UwiU8_0(.dout(w_dff_A_FR305U978_0),.din(w_dff_A_B6M3UwiU8_0),.clk(gclk));
	jdff dff_A_FR305U978_0(.dout(w_dff_A_GWB1OvPB0_0),.din(w_dff_A_FR305U978_0),.clk(gclk));
	jdff dff_A_GWB1OvPB0_0(.dout(w_dff_A_1KLeYKf19_0),.din(w_dff_A_GWB1OvPB0_0),.clk(gclk));
	jdff dff_A_1KLeYKf19_0(.dout(w_dff_A_pA7G6NbE5_0),.din(w_dff_A_1KLeYKf19_0),.clk(gclk));
	jdff dff_A_pA7G6NbE5_0(.dout(w_dff_A_FOwIA3GO4_0),.din(w_dff_A_pA7G6NbE5_0),.clk(gclk));
	jdff dff_A_FOwIA3GO4_0(.dout(w_dff_A_3Lcnqqwp8_0),.din(w_dff_A_FOwIA3GO4_0),.clk(gclk));
	jdff dff_A_3Lcnqqwp8_0(.dout(w_dff_A_qi1yUlle9_0),.din(w_dff_A_3Lcnqqwp8_0),.clk(gclk));
	jdff dff_A_qi1yUlle9_0(.dout(w_dff_A_g93qrmQt4_0),.din(w_dff_A_qi1yUlle9_0),.clk(gclk));
	jdff dff_A_g93qrmQt4_0(.dout(w_dff_A_lMOuGJNH0_0),.din(w_dff_A_g93qrmQt4_0),.clk(gclk));
	jdff dff_A_lMOuGJNH0_0(.dout(G534),.din(w_dff_A_lMOuGJNH0_0),.clk(gclk));
	jdff dff_A_0Bt12MFX2_1(.dout(w_dff_A_rz54Zfzl8_0),.din(w_dff_A_0Bt12MFX2_1),.clk(gclk));
	jdff dff_A_rz54Zfzl8_0(.dout(w_dff_A_QOlJGFcz9_0),.din(w_dff_A_rz54Zfzl8_0),.clk(gclk));
	jdff dff_A_QOlJGFcz9_0(.dout(w_dff_A_mMDuSWno3_0),.din(w_dff_A_QOlJGFcz9_0),.clk(gclk));
	jdff dff_A_mMDuSWno3_0(.dout(w_dff_A_HKdk1ZV48_0),.din(w_dff_A_mMDuSWno3_0),.clk(gclk));
	jdff dff_A_HKdk1ZV48_0(.dout(w_dff_A_u2bfEMbj0_0),.din(w_dff_A_HKdk1ZV48_0),.clk(gclk));
	jdff dff_A_u2bfEMbj0_0(.dout(w_dff_A_wn1z2M069_0),.din(w_dff_A_u2bfEMbj0_0),.clk(gclk));
	jdff dff_A_wn1z2M069_0(.dout(w_dff_A_BQyIudlE2_0),.din(w_dff_A_wn1z2M069_0),.clk(gclk));
	jdff dff_A_BQyIudlE2_0(.dout(w_dff_A_UuF8KJMG0_0),.din(w_dff_A_BQyIudlE2_0),.clk(gclk));
	jdff dff_A_UuF8KJMG0_0(.dout(w_dff_A_vrQXckRA3_0),.din(w_dff_A_UuF8KJMG0_0),.clk(gclk));
	jdff dff_A_vrQXckRA3_0(.dout(w_dff_A_htRr66EF8_0),.din(w_dff_A_vrQXckRA3_0),.clk(gclk));
	jdff dff_A_htRr66EF8_0(.dout(w_dff_A_tPtjB26c0_0),.din(w_dff_A_htRr66EF8_0),.clk(gclk));
	jdff dff_A_tPtjB26c0_0(.dout(w_dff_A_A0nrnv027_0),.din(w_dff_A_tPtjB26c0_0),.clk(gclk));
	jdff dff_A_A0nrnv027_0(.dout(w_dff_A_cBlnpneQ5_0),.din(w_dff_A_A0nrnv027_0),.clk(gclk));
	jdff dff_A_cBlnpneQ5_0(.dout(w_dff_A_sGINlGaG2_0),.din(w_dff_A_cBlnpneQ5_0),.clk(gclk));
	jdff dff_A_sGINlGaG2_0(.dout(w_dff_A_9ejt6TRu9_0),.din(w_dff_A_sGINlGaG2_0),.clk(gclk));
	jdff dff_A_9ejt6TRu9_0(.dout(w_dff_A_FTc2yuNf2_0),.din(w_dff_A_9ejt6TRu9_0),.clk(gclk));
	jdff dff_A_FTc2yuNf2_0(.dout(w_dff_A_Qo0qyAeu0_0),.din(w_dff_A_FTc2yuNf2_0),.clk(gclk));
	jdff dff_A_Qo0qyAeu0_0(.dout(w_dff_A_GYg1aoAD3_0),.din(w_dff_A_Qo0qyAeu0_0),.clk(gclk));
	jdff dff_A_GYg1aoAD3_0(.dout(w_dff_A_oUYbyAmX5_0),.din(w_dff_A_GYg1aoAD3_0),.clk(gclk));
	jdff dff_A_oUYbyAmX5_0(.dout(w_dff_A_v2oLe0R57_0),.din(w_dff_A_oUYbyAmX5_0),.clk(gclk));
	jdff dff_A_v2oLe0R57_0(.dout(w_dff_A_wfmD05pD2_0),.din(w_dff_A_v2oLe0R57_0),.clk(gclk));
	jdff dff_A_wfmD05pD2_0(.dout(w_dff_A_Q70oevZG8_0),.din(w_dff_A_wfmD05pD2_0),.clk(gclk));
	jdff dff_A_Q70oevZG8_0(.dout(w_dff_A_j9sDj5rm9_0),.din(w_dff_A_Q70oevZG8_0),.clk(gclk));
	jdff dff_A_j9sDj5rm9_0(.dout(w_dff_A_W7AnjYws3_0),.din(w_dff_A_j9sDj5rm9_0),.clk(gclk));
	jdff dff_A_W7AnjYws3_0(.dout(w_dff_A_Y0mNZce09_0),.din(w_dff_A_W7AnjYws3_0),.clk(gclk));
	jdff dff_A_Y0mNZce09_0(.dout(w_dff_A_hQAGEpKD2_0),.din(w_dff_A_Y0mNZce09_0),.clk(gclk));
	jdff dff_A_hQAGEpKD2_0(.dout(w_dff_A_vQBBfBVH8_0),.din(w_dff_A_hQAGEpKD2_0),.clk(gclk));
	jdff dff_A_vQBBfBVH8_0(.dout(w_dff_A_LpnxXwLD7_0),.din(w_dff_A_vQBBfBVH8_0),.clk(gclk));
	jdff dff_A_LpnxXwLD7_0(.dout(w_dff_A_MWFhbBBb3_0),.din(w_dff_A_LpnxXwLD7_0),.clk(gclk));
	jdff dff_A_MWFhbBBb3_0(.dout(w_dff_A_Ns6dSFxd8_0),.din(w_dff_A_MWFhbBBb3_0),.clk(gclk));
	jdff dff_A_Ns6dSFxd8_0(.dout(w_dff_A_A3DMHh212_0),.din(w_dff_A_Ns6dSFxd8_0),.clk(gclk));
	jdff dff_A_A3DMHh212_0(.dout(w_dff_A_Gorq8wbJ5_0),.din(w_dff_A_A3DMHh212_0),.clk(gclk));
	jdff dff_A_Gorq8wbJ5_0(.dout(w_dff_A_WotqE8j32_0),.din(w_dff_A_Gorq8wbJ5_0),.clk(gclk));
	jdff dff_A_WotqE8j32_0(.dout(w_dff_A_wD6MLlh62_0),.din(w_dff_A_WotqE8j32_0),.clk(gclk));
	jdff dff_A_wD6MLlh62_0(.dout(w_dff_A_IHPxW33Q6_0),.din(w_dff_A_wD6MLlh62_0),.clk(gclk));
	jdff dff_A_IHPxW33Q6_0(.dout(w_dff_A_thYjKvrw5_0),.din(w_dff_A_IHPxW33Q6_0),.clk(gclk));
	jdff dff_A_thYjKvrw5_0(.dout(w_dff_A_SfYhXbFh8_0),.din(w_dff_A_thYjKvrw5_0),.clk(gclk));
	jdff dff_A_SfYhXbFh8_0(.dout(G532),.din(w_dff_A_SfYhXbFh8_0),.clk(gclk));
	jdff dff_A_Btoykzj63_1(.dout(w_dff_A_DBPTFWA46_0),.din(w_dff_A_Btoykzj63_1),.clk(gclk));
	jdff dff_A_DBPTFWA46_0(.dout(w_dff_A_1iZsiXTt0_0),.din(w_dff_A_DBPTFWA46_0),.clk(gclk));
	jdff dff_A_1iZsiXTt0_0(.dout(w_dff_A_10uOhHhX1_0),.din(w_dff_A_1iZsiXTt0_0),.clk(gclk));
	jdff dff_A_10uOhHhX1_0(.dout(w_dff_A_BKq4JrHR1_0),.din(w_dff_A_10uOhHhX1_0),.clk(gclk));
	jdff dff_A_BKq4JrHR1_0(.dout(w_dff_A_Ptj17vIZ4_0),.din(w_dff_A_BKq4JrHR1_0),.clk(gclk));
	jdff dff_A_Ptj17vIZ4_0(.dout(w_dff_A_7lme9fO97_0),.din(w_dff_A_Ptj17vIZ4_0),.clk(gclk));
	jdff dff_A_7lme9fO97_0(.dout(w_dff_A_6QkS7RX48_0),.din(w_dff_A_7lme9fO97_0),.clk(gclk));
	jdff dff_A_6QkS7RX48_0(.dout(w_dff_A_GO9a7j7J8_0),.din(w_dff_A_6QkS7RX48_0),.clk(gclk));
	jdff dff_A_GO9a7j7J8_0(.dout(w_dff_A_93u88cEs6_0),.din(w_dff_A_GO9a7j7J8_0),.clk(gclk));
	jdff dff_A_93u88cEs6_0(.dout(w_dff_A_05SoZ6GH4_0),.din(w_dff_A_93u88cEs6_0),.clk(gclk));
	jdff dff_A_05SoZ6GH4_0(.dout(w_dff_A_MS2eqpsR2_0),.din(w_dff_A_05SoZ6GH4_0),.clk(gclk));
	jdff dff_A_MS2eqpsR2_0(.dout(w_dff_A_PXDy0tFB9_0),.din(w_dff_A_MS2eqpsR2_0),.clk(gclk));
	jdff dff_A_PXDy0tFB9_0(.dout(w_dff_A_GvDIfDeg8_0),.din(w_dff_A_PXDy0tFB9_0),.clk(gclk));
	jdff dff_A_GvDIfDeg8_0(.dout(w_dff_A_BvgvXHtP6_0),.din(w_dff_A_GvDIfDeg8_0),.clk(gclk));
	jdff dff_A_BvgvXHtP6_0(.dout(w_dff_A_tDA1uXjO3_0),.din(w_dff_A_BvgvXHtP6_0),.clk(gclk));
	jdff dff_A_tDA1uXjO3_0(.dout(w_dff_A_uJD1uhaZ6_0),.din(w_dff_A_tDA1uXjO3_0),.clk(gclk));
	jdff dff_A_uJD1uhaZ6_0(.dout(w_dff_A_l6BGa1Kh6_0),.din(w_dff_A_uJD1uhaZ6_0),.clk(gclk));
	jdff dff_A_l6BGa1Kh6_0(.dout(w_dff_A_1h69Ug5y4_0),.din(w_dff_A_l6BGa1Kh6_0),.clk(gclk));
	jdff dff_A_1h69Ug5y4_0(.dout(w_dff_A_lGcKFsVI7_0),.din(w_dff_A_1h69Ug5y4_0),.clk(gclk));
	jdff dff_A_lGcKFsVI7_0(.dout(w_dff_A_gP1jGYPA2_0),.din(w_dff_A_lGcKFsVI7_0),.clk(gclk));
	jdff dff_A_gP1jGYPA2_0(.dout(w_dff_A_9pX1HmKe5_0),.din(w_dff_A_gP1jGYPA2_0),.clk(gclk));
	jdff dff_A_9pX1HmKe5_0(.dout(w_dff_A_OgPKySg30_0),.din(w_dff_A_9pX1HmKe5_0),.clk(gclk));
	jdff dff_A_OgPKySg30_0(.dout(w_dff_A_WW5Y83WK3_0),.din(w_dff_A_OgPKySg30_0),.clk(gclk));
	jdff dff_A_WW5Y83WK3_0(.dout(w_dff_A_fb7eTxiX1_0),.din(w_dff_A_WW5Y83WK3_0),.clk(gclk));
	jdff dff_A_fb7eTxiX1_0(.dout(w_dff_A_tuH7XCB63_0),.din(w_dff_A_fb7eTxiX1_0),.clk(gclk));
	jdff dff_A_tuH7XCB63_0(.dout(w_dff_A_eJFWAKch7_0),.din(w_dff_A_tuH7XCB63_0),.clk(gclk));
	jdff dff_A_eJFWAKch7_0(.dout(w_dff_A_2cYrZ14W2_0),.din(w_dff_A_eJFWAKch7_0),.clk(gclk));
	jdff dff_A_2cYrZ14W2_0(.dout(w_dff_A_Gzc1oqwx2_0),.din(w_dff_A_2cYrZ14W2_0),.clk(gclk));
	jdff dff_A_Gzc1oqwx2_0(.dout(w_dff_A_sJdCtwPd5_0),.din(w_dff_A_Gzc1oqwx2_0),.clk(gclk));
	jdff dff_A_sJdCtwPd5_0(.dout(w_dff_A_UkTyILvP7_0),.din(w_dff_A_sJdCtwPd5_0),.clk(gclk));
	jdff dff_A_UkTyILvP7_0(.dout(w_dff_A_1WsKbfvO8_0),.din(w_dff_A_UkTyILvP7_0),.clk(gclk));
	jdff dff_A_1WsKbfvO8_0(.dout(w_dff_A_cSIiDGfg7_0),.din(w_dff_A_1WsKbfvO8_0),.clk(gclk));
	jdff dff_A_cSIiDGfg7_0(.dout(w_dff_A_uTekU42l4_0),.din(w_dff_A_cSIiDGfg7_0),.clk(gclk));
	jdff dff_A_uTekU42l4_0(.dout(w_dff_A_lxZTtf413_0),.din(w_dff_A_uTekU42l4_0),.clk(gclk));
	jdff dff_A_lxZTtf413_0(.dout(w_dff_A_86D7dpH85_0),.din(w_dff_A_lxZTtf413_0),.clk(gclk));
	jdff dff_A_86D7dpH85_0(.dout(w_dff_A_phxFdKTc5_0),.din(w_dff_A_86D7dpH85_0),.clk(gclk));
	jdff dff_A_phxFdKTc5_0(.dout(w_dff_A_wiS1sg8g9_0),.din(w_dff_A_phxFdKTc5_0),.clk(gclk));
	jdff dff_A_wiS1sg8g9_0(.dout(G530),.din(w_dff_A_wiS1sg8g9_0),.clk(gclk));
	jdff dff_A_Mp0c0e9T0_1(.dout(w_dff_A_QAN1kA3n9_0),.din(w_dff_A_Mp0c0e9T0_1),.clk(gclk));
	jdff dff_A_QAN1kA3n9_0(.dout(w_dff_A_ZLWJaSWH5_0),.din(w_dff_A_QAN1kA3n9_0),.clk(gclk));
	jdff dff_A_ZLWJaSWH5_0(.dout(w_dff_A_9iINOz5i0_0),.din(w_dff_A_ZLWJaSWH5_0),.clk(gclk));
	jdff dff_A_9iINOz5i0_0(.dout(w_dff_A_UHSRuxXA0_0),.din(w_dff_A_9iINOz5i0_0),.clk(gclk));
	jdff dff_A_UHSRuxXA0_0(.dout(w_dff_A_bobjiQpk6_0),.din(w_dff_A_UHSRuxXA0_0),.clk(gclk));
	jdff dff_A_bobjiQpk6_0(.dout(w_dff_A_06zGBEtv9_0),.din(w_dff_A_bobjiQpk6_0),.clk(gclk));
	jdff dff_A_06zGBEtv9_0(.dout(w_dff_A_zawuMBcn0_0),.din(w_dff_A_06zGBEtv9_0),.clk(gclk));
	jdff dff_A_zawuMBcn0_0(.dout(w_dff_A_LHrGMtDa1_0),.din(w_dff_A_zawuMBcn0_0),.clk(gclk));
	jdff dff_A_LHrGMtDa1_0(.dout(w_dff_A_YmhHv6QF0_0),.din(w_dff_A_LHrGMtDa1_0),.clk(gclk));
	jdff dff_A_YmhHv6QF0_0(.dout(w_dff_A_vZ6Yf7Ir1_0),.din(w_dff_A_YmhHv6QF0_0),.clk(gclk));
	jdff dff_A_vZ6Yf7Ir1_0(.dout(w_dff_A_UW4jf6w40_0),.din(w_dff_A_vZ6Yf7Ir1_0),.clk(gclk));
	jdff dff_A_UW4jf6w40_0(.dout(w_dff_A_1vubCZQV2_0),.din(w_dff_A_UW4jf6w40_0),.clk(gclk));
	jdff dff_A_1vubCZQV2_0(.dout(w_dff_A_jrvG67F59_0),.din(w_dff_A_1vubCZQV2_0),.clk(gclk));
	jdff dff_A_jrvG67F59_0(.dout(w_dff_A_gK1eM2kv2_0),.din(w_dff_A_jrvG67F59_0),.clk(gclk));
	jdff dff_A_gK1eM2kv2_0(.dout(w_dff_A_IIAWXZjE5_0),.din(w_dff_A_gK1eM2kv2_0),.clk(gclk));
	jdff dff_A_IIAWXZjE5_0(.dout(w_dff_A_Cwa9wFxL1_0),.din(w_dff_A_IIAWXZjE5_0),.clk(gclk));
	jdff dff_A_Cwa9wFxL1_0(.dout(w_dff_A_nA96BF973_0),.din(w_dff_A_Cwa9wFxL1_0),.clk(gclk));
	jdff dff_A_nA96BF973_0(.dout(w_dff_A_V3UQUgxY9_0),.din(w_dff_A_nA96BF973_0),.clk(gclk));
	jdff dff_A_V3UQUgxY9_0(.dout(w_dff_A_E4GdjO9Q8_0),.din(w_dff_A_V3UQUgxY9_0),.clk(gclk));
	jdff dff_A_E4GdjO9Q8_0(.dout(w_dff_A_tAHhD5eq9_0),.din(w_dff_A_E4GdjO9Q8_0),.clk(gclk));
	jdff dff_A_tAHhD5eq9_0(.dout(w_dff_A_bHB88nvE1_0),.din(w_dff_A_tAHhD5eq9_0),.clk(gclk));
	jdff dff_A_bHB88nvE1_0(.dout(w_dff_A_9XwpDm3b1_0),.din(w_dff_A_bHB88nvE1_0),.clk(gclk));
	jdff dff_A_9XwpDm3b1_0(.dout(w_dff_A_kCFIHhXa8_0),.din(w_dff_A_9XwpDm3b1_0),.clk(gclk));
	jdff dff_A_kCFIHhXa8_0(.dout(w_dff_A_tOIP03Re8_0),.din(w_dff_A_kCFIHhXa8_0),.clk(gclk));
	jdff dff_A_tOIP03Re8_0(.dout(w_dff_A_dyv9nxPW5_0),.din(w_dff_A_tOIP03Re8_0),.clk(gclk));
	jdff dff_A_dyv9nxPW5_0(.dout(w_dff_A_xKrQk2kV3_0),.din(w_dff_A_dyv9nxPW5_0),.clk(gclk));
	jdff dff_A_xKrQk2kV3_0(.dout(w_dff_A_aa9KrGIT1_0),.din(w_dff_A_xKrQk2kV3_0),.clk(gclk));
	jdff dff_A_aa9KrGIT1_0(.dout(w_dff_A_kbFOTB0W7_0),.din(w_dff_A_aa9KrGIT1_0),.clk(gclk));
	jdff dff_A_kbFOTB0W7_0(.dout(w_dff_A_69HdGNk67_0),.din(w_dff_A_kbFOTB0W7_0),.clk(gclk));
	jdff dff_A_69HdGNk67_0(.dout(w_dff_A_1YYDhmyB3_0),.din(w_dff_A_69HdGNk67_0),.clk(gclk));
	jdff dff_A_1YYDhmyB3_0(.dout(w_dff_A_lOghKWBG3_0),.din(w_dff_A_1YYDhmyB3_0),.clk(gclk));
	jdff dff_A_lOghKWBG3_0(.dout(w_dff_A_CcIk14aE8_0),.din(w_dff_A_lOghKWBG3_0),.clk(gclk));
	jdff dff_A_CcIk14aE8_0(.dout(w_dff_A_qh42paZS2_0),.din(w_dff_A_CcIk14aE8_0),.clk(gclk));
	jdff dff_A_qh42paZS2_0(.dout(w_dff_A_9kBu6i9W7_0),.din(w_dff_A_qh42paZS2_0),.clk(gclk));
	jdff dff_A_9kBu6i9W7_0(.dout(w_dff_A_RkerbP610_0),.din(w_dff_A_9kBu6i9W7_0),.clk(gclk));
	jdff dff_A_RkerbP610_0(.dout(w_dff_A_Pzq9DuDH9_0),.din(w_dff_A_RkerbP610_0),.clk(gclk));
	jdff dff_A_Pzq9DuDH9_0(.dout(w_dff_A_qWJuqif76_0),.din(w_dff_A_Pzq9DuDH9_0),.clk(gclk));
	jdff dff_A_qWJuqif76_0(.dout(G528),.din(w_dff_A_qWJuqif76_0),.clk(gclk));
	jdff dff_A_ReeCzHam0_1(.dout(w_dff_A_VAtd6ojO6_0),.din(w_dff_A_ReeCzHam0_1),.clk(gclk));
	jdff dff_A_VAtd6ojO6_0(.dout(w_dff_A_fgLIz7579_0),.din(w_dff_A_VAtd6ojO6_0),.clk(gclk));
	jdff dff_A_fgLIz7579_0(.dout(w_dff_A_e6psGgm19_0),.din(w_dff_A_fgLIz7579_0),.clk(gclk));
	jdff dff_A_e6psGgm19_0(.dout(w_dff_A_HU1Er5R40_0),.din(w_dff_A_e6psGgm19_0),.clk(gclk));
	jdff dff_A_HU1Er5R40_0(.dout(w_dff_A_p0ejQOe19_0),.din(w_dff_A_HU1Er5R40_0),.clk(gclk));
	jdff dff_A_p0ejQOe19_0(.dout(w_dff_A_OakH9ahz8_0),.din(w_dff_A_p0ejQOe19_0),.clk(gclk));
	jdff dff_A_OakH9ahz8_0(.dout(w_dff_A_namE0PEt9_0),.din(w_dff_A_OakH9ahz8_0),.clk(gclk));
	jdff dff_A_namE0PEt9_0(.dout(w_dff_A_bKBHiHXY7_0),.din(w_dff_A_namE0PEt9_0),.clk(gclk));
	jdff dff_A_bKBHiHXY7_0(.dout(w_dff_A_5JS1xSX60_0),.din(w_dff_A_bKBHiHXY7_0),.clk(gclk));
	jdff dff_A_5JS1xSX60_0(.dout(w_dff_A_BdGG74w49_0),.din(w_dff_A_5JS1xSX60_0),.clk(gclk));
	jdff dff_A_BdGG74w49_0(.dout(w_dff_A_LxevbDgk3_0),.din(w_dff_A_BdGG74w49_0),.clk(gclk));
	jdff dff_A_LxevbDgk3_0(.dout(w_dff_A_dyX5QeVm6_0),.din(w_dff_A_LxevbDgk3_0),.clk(gclk));
	jdff dff_A_dyX5QeVm6_0(.dout(w_dff_A_7wrVGsvS6_0),.din(w_dff_A_dyX5QeVm6_0),.clk(gclk));
	jdff dff_A_7wrVGsvS6_0(.dout(w_dff_A_mdvTV2M94_0),.din(w_dff_A_7wrVGsvS6_0),.clk(gclk));
	jdff dff_A_mdvTV2M94_0(.dout(w_dff_A_ZOXB797B5_0),.din(w_dff_A_mdvTV2M94_0),.clk(gclk));
	jdff dff_A_ZOXB797B5_0(.dout(w_dff_A_XqDhwwTU2_0),.din(w_dff_A_ZOXB797B5_0),.clk(gclk));
	jdff dff_A_XqDhwwTU2_0(.dout(w_dff_A_FN2meJcS4_0),.din(w_dff_A_XqDhwwTU2_0),.clk(gclk));
	jdff dff_A_FN2meJcS4_0(.dout(w_dff_A_UWDI1rcn2_0),.din(w_dff_A_FN2meJcS4_0),.clk(gclk));
	jdff dff_A_UWDI1rcn2_0(.dout(w_dff_A_nQ5FjT9j2_0),.din(w_dff_A_UWDI1rcn2_0),.clk(gclk));
	jdff dff_A_nQ5FjT9j2_0(.dout(w_dff_A_VMdq6R6P3_0),.din(w_dff_A_nQ5FjT9j2_0),.clk(gclk));
	jdff dff_A_VMdq6R6P3_0(.dout(w_dff_A_UcPK5xLx8_0),.din(w_dff_A_VMdq6R6P3_0),.clk(gclk));
	jdff dff_A_UcPK5xLx8_0(.dout(w_dff_A_VaMgQ7rf1_0),.din(w_dff_A_UcPK5xLx8_0),.clk(gclk));
	jdff dff_A_VaMgQ7rf1_0(.dout(w_dff_A_3KRlIzmx2_0),.din(w_dff_A_VaMgQ7rf1_0),.clk(gclk));
	jdff dff_A_3KRlIzmx2_0(.dout(w_dff_A_1iZOStDw8_0),.din(w_dff_A_3KRlIzmx2_0),.clk(gclk));
	jdff dff_A_1iZOStDw8_0(.dout(w_dff_A_WlBN6Pna2_0),.din(w_dff_A_1iZOStDw8_0),.clk(gclk));
	jdff dff_A_WlBN6Pna2_0(.dout(w_dff_A_wYWfktBK4_0),.din(w_dff_A_WlBN6Pna2_0),.clk(gclk));
	jdff dff_A_wYWfktBK4_0(.dout(w_dff_A_c278mtd82_0),.din(w_dff_A_wYWfktBK4_0),.clk(gclk));
	jdff dff_A_c278mtd82_0(.dout(w_dff_A_6Kt4kC7J3_0),.din(w_dff_A_c278mtd82_0),.clk(gclk));
	jdff dff_A_6Kt4kC7J3_0(.dout(w_dff_A_JxCayiBq8_0),.din(w_dff_A_6Kt4kC7J3_0),.clk(gclk));
	jdff dff_A_JxCayiBq8_0(.dout(w_dff_A_2EzZnyBp1_0),.din(w_dff_A_JxCayiBq8_0),.clk(gclk));
	jdff dff_A_2EzZnyBp1_0(.dout(w_dff_A_tJsHhYII5_0),.din(w_dff_A_2EzZnyBp1_0),.clk(gclk));
	jdff dff_A_tJsHhYII5_0(.dout(w_dff_A_BDPAqsf18_0),.din(w_dff_A_tJsHhYII5_0),.clk(gclk));
	jdff dff_A_BDPAqsf18_0(.dout(w_dff_A_LDtMW9hx8_0),.din(w_dff_A_BDPAqsf18_0),.clk(gclk));
	jdff dff_A_LDtMW9hx8_0(.dout(w_dff_A_9K7Cq7G98_0),.din(w_dff_A_LDtMW9hx8_0),.clk(gclk));
	jdff dff_A_9K7Cq7G98_0(.dout(w_dff_A_vSWIXsnq3_0),.din(w_dff_A_9K7Cq7G98_0),.clk(gclk));
	jdff dff_A_vSWIXsnq3_0(.dout(w_dff_A_JsxhfXln5_0),.din(w_dff_A_vSWIXsnq3_0),.clk(gclk));
	jdff dff_A_JsxhfXln5_0(.dout(w_dff_A_R8bl4UCH7_0),.din(w_dff_A_JsxhfXln5_0),.clk(gclk));
	jdff dff_A_R8bl4UCH7_0(.dout(G526),.din(w_dff_A_R8bl4UCH7_0),.clk(gclk));
	jdff dff_A_wNDkqV9X6_1(.dout(w_dff_A_r0WQzJi04_0),.din(w_dff_A_wNDkqV9X6_1),.clk(gclk));
	jdff dff_A_r0WQzJi04_0(.dout(w_dff_A_L7TZ5b2t1_0),.din(w_dff_A_r0WQzJi04_0),.clk(gclk));
	jdff dff_A_L7TZ5b2t1_0(.dout(w_dff_A_S8GueEaO6_0),.din(w_dff_A_L7TZ5b2t1_0),.clk(gclk));
	jdff dff_A_S8GueEaO6_0(.dout(w_dff_A_d2iAScxU8_0),.din(w_dff_A_S8GueEaO6_0),.clk(gclk));
	jdff dff_A_d2iAScxU8_0(.dout(w_dff_A_PeyvzLzQ4_0),.din(w_dff_A_d2iAScxU8_0),.clk(gclk));
	jdff dff_A_PeyvzLzQ4_0(.dout(w_dff_A_ajzfxveW1_0),.din(w_dff_A_PeyvzLzQ4_0),.clk(gclk));
	jdff dff_A_ajzfxveW1_0(.dout(w_dff_A_Iy9YAmz36_0),.din(w_dff_A_ajzfxveW1_0),.clk(gclk));
	jdff dff_A_Iy9YAmz36_0(.dout(w_dff_A_W35tNQns1_0),.din(w_dff_A_Iy9YAmz36_0),.clk(gclk));
	jdff dff_A_W35tNQns1_0(.dout(w_dff_A_lWT33Ufv7_0),.din(w_dff_A_W35tNQns1_0),.clk(gclk));
	jdff dff_A_lWT33Ufv7_0(.dout(w_dff_A_ScI156pN7_0),.din(w_dff_A_lWT33Ufv7_0),.clk(gclk));
	jdff dff_A_ScI156pN7_0(.dout(w_dff_A_FAqIWjmC6_0),.din(w_dff_A_ScI156pN7_0),.clk(gclk));
	jdff dff_A_FAqIWjmC6_0(.dout(w_dff_A_fyOoPG2X5_0),.din(w_dff_A_FAqIWjmC6_0),.clk(gclk));
	jdff dff_A_fyOoPG2X5_0(.dout(w_dff_A_3OgmrwKD1_0),.din(w_dff_A_fyOoPG2X5_0),.clk(gclk));
	jdff dff_A_3OgmrwKD1_0(.dout(w_dff_A_Fs0ju9HF8_0),.din(w_dff_A_3OgmrwKD1_0),.clk(gclk));
	jdff dff_A_Fs0ju9HF8_0(.dout(w_dff_A_uCWLPIYQ2_0),.din(w_dff_A_Fs0ju9HF8_0),.clk(gclk));
	jdff dff_A_uCWLPIYQ2_0(.dout(w_dff_A_LW9T8MCW7_0),.din(w_dff_A_uCWLPIYQ2_0),.clk(gclk));
	jdff dff_A_LW9T8MCW7_0(.dout(w_dff_A_IYKKslCv1_0),.din(w_dff_A_LW9T8MCW7_0),.clk(gclk));
	jdff dff_A_IYKKslCv1_0(.dout(w_dff_A_4nNAy4ns5_0),.din(w_dff_A_IYKKslCv1_0),.clk(gclk));
	jdff dff_A_4nNAy4ns5_0(.dout(w_dff_A_oCRZZGWp7_0),.din(w_dff_A_4nNAy4ns5_0),.clk(gclk));
	jdff dff_A_oCRZZGWp7_0(.dout(w_dff_A_XsdgfgUC7_0),.din(w_dff_A_oCRZZGWp7_0),.clk(gclk));
	jdff dff_A_XsdgfgUC7_0(.dout(w_dff_A_xABX73f49_0),.din(w_dff_A_XsdgfgUC7_0),.clk(gclk));
	jdff dff_A_xABX73f49_0(.dout(w_dff_A_zyGl4EHl4_0),.din(w_dff_A_xABX73f49_0),.clk(gclk));
	jdff dff_A_zyGl4EHl4_0(.dout(w_dff_A_e3Ydfltt6_0),.din(w_dff_A_zyGl4EHl4_0),.clk(gclk));
	jdff dff_A_e3Ydfltt6_0(.dout(w_dff_A_Y83BffQe9_0),.din(w_dff_A_e3Ydfltt6_0),.clk(gclk));
	jdff dff_A_Y83BffQe9_0(.dout(w_dff_A_sKtdNFkT7_0),.din(w_dff_A_Y83BffQe9_0),.clk(gclk));
	jdff dff_A_sKtdNFkT7_0(.dout(w_dff_A_tJtXXvJM5_0),.din(w_dff_A_sKtdNFkT7_0),.clk(gclk));
	jdff dff_A_tJtXXvJM5_0(.dout(w_dff_A_stbY7ACb3_0),.din(w_dff_A_tJtXXvJM5_0),.clk(gclk));
	jdff dff_A_stbY7ACb3_0(.dout(w_dff_A_mHiYY7PV6_0),.din(w_dff_A_stbY7ACb3_0),.clk(gclk));
	jdff dff_A_mHiYY7PV6_0(.dout(w_dff_A_pxrAQ3mi1_0),.din(w_dff_A_mHiYY7PV6_0),.clk(gclk));
	jdff dff_A_pxrAQ3mi1_0(.dout(w_dff_A_vDJsEelS6_0),.din(w_dff_A_pxrAQ3mi1_0),.clk(gclk));
	jdff dff_A_vDJsEelS6_0(.dout(w_dff_A_nMMYk4NR7_0),.din(w_dff_A_vDJsEelS6_0),.clk(gclk));
	jdff dff_A_nMMYk4NR7_0(.dout(w_dff_A_f6L6XOUy6_0),.din(w_dff_A_nMMYk4NR7_0),.clk(gclk));
	jdff dff_A_f6L6XOUy6_0(.dout(w_dff_A_7l4D5zCO0_0),.din(w_dff_A_f6L6XOUy6_0),.clk(gclk));
	jdff dff_A_7l4D5zCO0_0(.dout(w_dff_A_TooqVmUK2_0),.din(w_dff_A_7l4D5zCO0_0),.clk(gclk));
	jdff dff_A_TooqVmUK2_0(.dout(w_dff_A_fTxHXQjX8_0),.din(w_dff_A_TooqVmUK2_0),.clk(gclk));
	jdff dff_A_fTxHXQjX8_0(.dout(w_dff_A_HTCSvGZZ3_0),.din(w_dff_A_fTxHXQjX8_0),.clk(gclk));
	jdff dff_A_HTCSvGZZ3_0(.dout(w_dff_A_4hC2oC508_0),.din(w_dff_A_HTCSvGZZ3_0),.clk(gclk));
	jdff dff_A_4hC2oC508_0(.dout(G524),.din(w_dff_A_4hC2oC508_0),.clk(gclk));
	jdff dff_A_TnC3fYtR3_1(.dout(w_dff_A_OusjvvD54_0),.din(w_dff_A_TnC3fYtR3_1),.clk(gclk));
	jdff dff_A_OusjvvD54_0(.dout(w_dff_A_X91AlhYc5_0),.din(w_dff_A_OusjvvD54_0),.clk(gclk));
	jdff dff_A_X91AlhYc5_0(.dout(w_dff_A_MyYDfWOG7_0),.din(w_dff_A_X91AlhYc5_0),.clk(gclk));
	jdff dff_A_MyYDfWOG7_0(.dout(w_dff_A_Ugd1jy1D7_0),.din(w_dff_A_MyYDfWOG7_0),.clk(gclk));
	jdff dff_A_Ugd1jy1D7_0(.dout(w_dff_A_DkDYaxly0_0),.din(w_dff_A_Ugd1jy1D7_0),.clk(gclk));
	jdff dff_A_DkDYaxly0_0(.dout(w_dff_A_CUQTXiKE8_0),.din(w_dff_A_DkDYaxly0_0),.clk(gclk));
	jdff dff_A_CUQTXiKE8_0(.dout(w_dff_A_7NUqq3zw5_0),.din(w_dff_A_CUQTXiKE8_0),.clk(gclk));
	jdff dff_A_7NUqq3zw5_0(.dout(w_dff_A_vLtl5ggm3_0),.din(w_dff_A_7NUqq3zw5_0),.clk(gclk));
	jdff dff_A_vLtl5ggm3_0(.dout(w_dff_A_njdB9fOO3_0),.din(w_dff_A_vLtl5ggm3_0),.clk(gclk));
	jdff dff_A_njdB9fOO3_0(.dout(w_dff_A_fCkscxnd0_0),.din(w_dff_A_njdB9fOO3_0),.clk(gclk));
	jdff dff_A_fCkscxnd0_0(.dout(w_dff_A_IqkPXJAb0_0),.din(w_dff_A_fCkscxnd0_0),.clk(gclk));
	jdff dff_A_IqkPXJAb0_0(.dout(w_dff_A_er7grrb98_0),.din(w_dff_A_IqkPXJAb0_0),.clk(gclk));
	jdff dff_A_er7grrb98_0(.dout(w_dff_A_OKNEDAyD6_0),.din(w_dff_A_er7grrb98_0),.clk(gclk));
	jdff dff_A_OKNEDAyD6_0(.dout(w_dff_A_aaO32Qjc1_0),.din(w_dff_A_OKNEDAyD6_0),.clk(gclk));
	jdff dff_A_aaO32Qjc1_0(.dout(w_dff_A_j6ckGRFj5_0),.din(w_dff_A_aaO32Qjc1_0),.clk(gclk));
	jdff dff_A_j6ckGRFj5_0(.dout(w_dff_A_j9CNGlJS8_0),.din(w_dff_A_j6ckGRFj5_0),.clk(gclk));
	jdff dff_A_j9CNGlJS8_0(.dout(w_dff_A_qJBXjZCB1_0),.din(w_dff_A_j9CNGlJS8_0),.clk(gclk));
	jdff dff_A_qJBXjZCB1_0(.dout(w_dff_A_K2dViIzc0_0),.din(w_dff_A_qJBXjZCB1_0),.clk(gclk));
	jdff dff_A_K2dViIzc0_0(.dout(w_dff_A_RxcO7qo52_0),.din(w_dff_A_K2dViIzc0_0),.clk(gclk));
	jdff dff_A_RxcO7qo52_0(.dout(w_dff_A_RUL3SLqx6_0),.din(w_dff_A_RxcO7qo52_0),.clk(gclk));
	jdff dff_A_RUL3SLqx6_0(.dout(w_dff_A_DlqLsbAj3_0),.din(w_dff_A_RUL3SLqx6_0),.clk(gclk));
	jdff dff_A_DlqLsbAj3_0(.dout(w_dff_A_VAF0i8ZA2_0),.din(w_dff_A_DlqLsbAj3_0),.clk(gclk));
	jdff dff_A_VAF0i8ZA2_0(.dout(w_dff_A_aWDQUBIU0_0),.din(w_dff_A_VAF0i8ZA2_0),.clk(gclk));
	jdff dff_A_aWDQUBIU0_0(.dout(w_dff_A_ojutfHwt4_0),.din(w_dff_A_aWDQUBIU0_0),.clk(gclk));
	jdff dff_A_ojutfHwt4_0(.dout(w_dff_A_mPYCv19x1_0),.din(w_dff_A_ojutfHwt4_0),.clk(gclk));
	jdff dff_A_mPYCv19x1_0(.dout(w_dff_A_8hb3iYw81_0),.din(w_dff_A_mPYCv19x1_0),.clk(gclk));
	jdff dff_A_8hb3iYw81_0(.dout(w_dff_A_3zIjocPC5_0),.din(w_dff_A_8hb3iYw81_0),.clk(gclk));
	jdff dff_A_3zIjocPC5_0(.dout(w_dff_A_PypNKC9r3_0),.din(w_dff_A_3zIjocPC5_0),.clk(gclk));
	jdff dff_A_PypNKC9r3_0(.dout(w_dff_A_xW0JxjF53_0),.din(w_dff_A_PypNKC9r3_0),.clk(gclk));
	jdff dff_A_xW0JxjF53_0(.dout(w_dff_A_4VMtYlsa4_0),.din(w_dff_A_xW0JxjF53_0),.clk(gclk));
	jdff dff_A_4VMtYlsa4_0(.dout(w_dff_A_ivYYIrsJ4_0),.din(w_dff_A_4VMtYlsa4_0),.clk(gclk));
	jdff dff_A_ivYYIrsJ4_0(.dout(w_dff_A_ftxL8Nqp4_0),.din(w_dff_A_ivYYIrsJ4_0),.clk(gclk));
	jdff dff_A_ftxL8Nqp4_0(.dout(w_dff_A_q3D0uZNR4_0),.din(w_dff_A_ftxL8Nqp4_0),.clk(gclk));
	jdff dff_A_q3D0uZNR4_0(.dout(w_dff_A_wB1HIsRx4_0),.din(w_dff_A_q3D0uZNR4_0),.clk(gclk));
	jdff dff_A_wB1HIsRx4_0(.dout(w_dff_A_TqJ2Mjfy5_0),.din(w_dff_A_wB1HIsRx4_0),.clk(gclk));
	jdff dff_A_TqJ2Mjfy5_0(.dout(w_dff_A_Uj2ECwpB9_0),.din(w_dff_A_TqJ2Mjfy5_0),.clk(gclk));
	jdff dff_A_Uj2ECwpB9_0(.dout(w_dff_A_Xetz9aSM4_0),.din(w_dff_A_Uj2ECwpB9_0),.clk(gclk));
	jdff dff_A_Xetz9aSM4_0(.dout(G279),.din(w_dff_A_Xetz9aSM4_0),.clk(gclk));
	jdff dff_A_3rxkWg5S9_1(.dout(w_dff_A_LE2rjmPW1_0),.din(w_dff_A_3rxkWg5S9_1),.clk(gclk));
	jdff dff_A_LE2rjmPW1_0(.dout(w_dff_A_QytUHVI58_0),.din(w_dff_A_LE2rjmPW1_0),.clk(gclk));
	jdff dff_A_QytUHVI58_0(.dout(w_dff_A_KorsMJiw9_0),.din(w_dff_A_QytUHVI58_0),.clk(gclk));
	jdff dff_A_KorsMJiw9_0(.dout(w_dff_A_pgbKMHN99_0),.din(w_dff_A_KorsMJiw9_0),.clk(gclk));
	jdff dff_A_pgbKMHN99_0(.dout(w_dff_A_BXE8Vq7z6_0),.din(w_dff_A_pgbKMHN99_0),.clk(gclk));
	jdff dff_A_BXE8Vq7z6_0(.dout(w_dff_A_04mTBibP3_0),.din(w_dff_A_BXE8Vq7z6_0),.clk(gclk));
	jdff dff_A_04mTBibP3_0(.dout(w_dff_A_KaB9jzjV7_0),.din(w_dff_A_04mTBibP3_0),.clk(gclk));
	jdff dff_A_KaB9jzjV7_0(.dout(w_dff_A_9pC5nFss3_0),.din(w_dff_A_KaB9jzjV7_0),.clk(gclk));
	jdff dff_A_9pC5nFss3_0(.dout(w_dff_A_CwEBZBp51_0),.din(w_dff_A_9pC5nFss3_0),.clk(gclk));
	jdff dff_A_CwEBZBp51_0(.dout(w_dff_A_l9Vh7Do05_0),.din(w_dff_A_CwEBZBp51_0),.clk(gclk));
	jdff dff_A_l9Vh7Do05_0(.dout(w_dff_A_vOvfAFlI4_0),.din(w_dff_A_l9Vh7Do05_0),.clk(gclk));
	jdff dff_A_vOvfAFlI4_0(.dout(w_dff_A_YIdbzm4r7_0),.din(w_dff_A_vOvfAFlI4_0),.clk(gclk));
	jdff dff_A_YIdbzm4r7_0(.dout(w_dff_A_mZUaz71h5_0),.din(w_dff_A_YIdbzm4r7_0),.clk(gclk));
	jdff dff_A_mZUaz71h5_0(.dout(w_dff_A_HPPW8HyZ8_0),.din(w_dff_A_mZUaz71h5_0),.clk(gclk));
	jdff dff_A_HPPW8HyZ8_0(.dout(w_dff_A_wR0eZlHq0_0),.din(w_dff_A_HPPW8HyZ8_0),.clk(gclk));
	jdff dff_A_wR0eZlHq0_0(.dout(w_dff_A_rimFFKaY6_0),.din(w_dff_A_wR0eZlHq0_0),.clk(gclk));
	jdff dff_A_rimFFKaY6_0(.dout(w_dff_A_RkKW1rvY3_0),.din(w_dff_A_rimFFKaY6_0),.clk(gclk));
	jdff dff_A_RkKW1rvY3_0(.dout(w_dff_A_QhWst42O8_0),.din(w_dff_A_RkKW1rvY3_0),.clk(gclk));
	jdff dff_A_QhWst42O8_0(.dout(w_dff_A_PKO1MUXk5_0),.din(w_dff_A_QhWst42O8_0),.clk(gclk));
	jdff dff_A_PKO1MUXk5_0(.dout(w_dff_A_OwNzPaYB5_0),.din(w_dff_A_PKO1MUXk5_0),.clk(gclk));
	jdff dff_A_OwNzPaYB5_0(.dout(w_dff_A_7UITA4t27_0),.din(w_dff_A_OwNzPaYB5_0),.clk(gclk));
	jdff dff_A_7UITA4t27_0(.dout(w_dff_A_CXJqxKHW3_0),.din(w_dff_A_7UITA4t27_0),.clk(gclk));
	jdff dff_A_CXJqxKHW3_0(.dout(w_dff_A_I73LU5FT4_0),.din(w_dff_A_CXJqxKHW3_0),.clk(gclk));
	jdff dff_A_I73LU5FT4_0(.dout(w_dff_A_4ltZu5ML1_0),.din(w_dff_A_I73LU5FT4_0),.clk(gclk));
	jdff dff_A_4ltZu5ML1_0(.dout(w_dff_A_9Tkyn4VC7_0),.din(w_dff_A_4ltZu5ML1_0),.clk(gclk));
	jdff dff_A_9Tkyn4VC7_0(.dout(w_dff_A_Lg4ALZlf9_0),.din(w_dff_A_9Tkyn4VC7_0),.clk(gclk));
	jdff dff_A_Lg4ALZlf9_0(.dout(w_dff_A_hKpMjOIw7_0),.din(w_dff_A_Lg4ALZlf9_0),.clk(gclk));
	jdff dff_A_hKpMjOIw7_0(.dout(w_dff_A_nLo2os3J5_0),.din(w_dff_A_hKpMjOIw7_0),.clk(gclk));
	jdff dff_A_nLo2os3J5_0(.dout(w_dff_A_KA2T3DwW2_0),.din(w_dff_A_nLo2os3J5_0),.clk(gclk));
	jdff dff_A_KA2T3DwW2_0(.dout(w_dff_A_f4BbQmFp5_0),.din(w_dff_A_KA2T3DwW2_0),.clk(gclk));
	jdff dff_A_f4BbQmFp5_0(.dout(w_dff_A_K06CakgD0_0),.din(w_dff_A_f4BbQmFp5_0),.clk(gclk));
	jdff dff_A_K06CakgD0_0(.dout(w_dff_A_eKKYvRWU5_0),.din(w_dff_A_K06CakgD0_0),.clk(gclk));
	jdff dff_A_eKKYvRWU5_0(.dout(w_dff_A_YHgJ9OAa6_0),.din(w_dff_A_eKKYvRWU5_0),.clk(gclk));
	jdff dff_A_YHgJ9OAa6_0(.dout(w_dff_A_qtR2F5Pr4_0),.din(w_dff_A_YHgJ9OAa6_0),.clk(gclk));
	jdff dff_A_qtR2F5Pr4_0(.dout(w_dff_A_zKxJyPZ97_0),.din(w_dff_A_qtR2F5Pr4_0),.clk(gclk));
	jdff dff_A_zKxJyPZ97_0(.dout(w_dff_A_xK5nuJMO5_0),.din(w_dff_A_zKxJyPZ97_0),.clk(gclk));
	jdff dff_A_xK5nuJMO5_0(.dout(w_dff_A_NIFIvBQ92_0),.din(w_dff_A_xK5nuJMO5_0),.clk(gclk));
	jdff dff_A_NIFIvBQ92_0(.dout(G436),.din(w_dff_A_NIFIvBQ92_0),.clk(gclk));
	jdff dff_A_VGhsnYzH9_1(.dout(w_dff_A_k0kxFyxg5_0),.din(w_dff_A_VGhsnYzH9_1),.clk(gclk));
	jdff dff_A_k0kxFyxg5_0(.dout(w_dff_A_0Kub6lVs4_0),.din(w_dff_A_k0kxFyxg5_0),.clk(gclk));
	jdff dff_A_0Kub6lVs4_0(.dout(w_dff_A_vpkqxgEZ9_0),.din(w_dff_A_0Kub6lVs4_0),.clk(gclk));
	jdff dff_A_vpkqxgEZ9_0(.dout(w_dff_A_3D01UMmf6_0),.din(w_dff_A_vpkqxgEZ9_0),.clk(gclk));
	jdff dff_A_3D01UMmf6_0(.dout(w_dff_A_EHtETE1Z0_0),.din(w_dff_A_3D01UMmf6_0),.clk(gclk));
	jdff dff_A_EHtETE1Z0_0(.dout(w_dff_A_Pv3fbyyt1_0),.din(w_dff_A_EHtETE1Z0_0),.clk(gclk));
	jdff dff_A_Pv3fbyyt1_0(.dout(w_dff_A_4E9fniZY7_0),.din(w_dff_A_Pv3fbyyt1_0),.clk(gclk));
	jdff dff_A_4E9fniZY7_0(.dout(w_dff_A_MYc4JEl05_0),.din(w_dff_A_4E9fniZY7_0),.clk(gclk));
	jdff dff_A_MYc4JEl05_0(.dout(w_dff_A_oe8rHOUi9_0),.din(w_dff_A_MYc4JEl05_0),.clk(gclk));
	jdff dff_A_oe8rHOUi9_0(.dout(w_dff_A_OWaAt6vZ5_0),.din(w_dff_A_oe8rHOUi9_0),.clk(gclk));
	jdff dff_A_OWaAt6vZ5_0(.dout(w_dff_A_jkL1XRRL0_0),.din(w_dff_A_OWaAt6vZ5_0),.clk(gclk));
	jdff dff_A_jkL1XRRL0_0(.dout(w_dff_A_pOnNXAhg8_0),.din(w_dff_A_jkL1XRRL0_0),.clk(gclk));
	jdff dff_A_pOnNXAhg8_0(.dout(w_dff_A_MNOt3Rpk5_0),.din(w_dff_A_pOnNXAhg8_0),.clk(gclk));
	jdff dff_A_MNOt3Rpk5_0(.dout(w_dff_A_8bnmCgFn2_0),.din(w_dff_A_MNOt3Rpk5_0),.clk(gclk));
	jdff dff_A_8bnmCgFn2_0(.dout(w_dff_A_GFqcIxkx0_0),.din(w_dff_A_8bnmCgFn2_0),.clk(gclk));
	jdff dff_A_GFqcIxkx0_0(.dout(w_dff_A_hK3okQKZ0_0),.din(w_dff_A_GFqcIxkx0_0),.clk(gclk));
	jdff dff_A_hK3okQKZ0_0(.dout(w_dff_A_6zYNJLny9_0),.din(w_dff_A_hK3okQKZ0_0),.clk(gclk));
	jdff dff_A_6zYNJLny9_0(.dout(w_dff_A_MEoDZomE2_0),.din(w_dff_A_6zYNJLny9_0),.clk(gclk));
	jdff dff_A_MEoDZomE2_0(.dout(w_dff_A_JnNj51JT8_0),.din(w_dff_A_MEoDZomE2_0),.clk(gclk));
	jdff dff_A_JnNj51JT8_0(.dout(w_dff_A_JprOozQS7_0),.din(w_dff_A_JnNj51JT8_0),.clk(gclk));
	jdff dff_A_JprOozQS7_0(.dout(w_dff_A_Ip0iVPii6_0),.din(w_dff_A_JprOozQS7_0),.clk(gclk));
	jdff dff_A_Ip0iVPii6_0(.dout(w_dff_A_R0sbkSL78_0),.din(w_dff_A_Ip0iVPii6_0),.clk(gclk));
	jdff dff_A_R0sbkSL78_0(.dout(w_dff_A_tllcEnYY0_0),.din(w_dff_A_R0sbkSL78_0),.clk(gclk));
	jdff dff_A_tllcEnYY0_0(.dout(w_dff_A_0tEM0fhe1_0),.din(w_dff_A_tllcEnYY0_0),.clk(gclk));
	jdff dff_A_0tEM0fhe1_0(.dout(w_dff_A_SMqhLXjc6_0),.din(w_dff_A_0tEM0fhe1_0),.clk(gclk));
	jdff dff_A_SMqhLXjc6_0(.dout(w_dff_A_qgBiWEHo1_0),.din(w_dff_A_SMqhLXjc6_0),.clk(gclk));
	jdff dff_A_qgBiWEHo1_0(.dout(w_dff_A_Fp9Uf06n7_0),.din(w_dff_A_qgBiWEHo1_0),.clk(gclk));
	jdff dff_A_Fp9Uf06n7_0(.dout(w_dff_A_nSo6I93q6_0),.din(w_dff_A_Fp9Uf06n7_0),.clk(gclk));
	jdff dff_A_nSo6I93q6_0(.dout(w_dff_A_acXF0J0C6_0),.din(w_dff_A_nSo6I93q6_0),.clk(gclk));
	jdff dff_A_acXF0J0C6_0(.dout(w_dff_A_VCkrEa8s3_0),.din(w_dff_A_acXF0J0C6_0),.clk(gclk));
	jdff dff_A_VCkrEa8s3_0(.dout(w_dff_A_dJHNVGkm4_0),.din(w_dff_A_VCkrEa8s3_0),.clk(gclk));
	jdff dff_A_dJHNVGkm4_0(.dout(w_dff_A_cgUuihUD0_0),.din(w_dff_A_dJHNVGkm4_0),.clk(gclk));
	jdff dff_A_cgUuihUD0_0(.dout(w_dff_A_ntG72hgR0_0),.din(w_dff_A_cgUuihUD0_0),.clk(gclk));
	jdff dff_A_ntG72hgR0_0(.dout(w_dff_A_uYXQn4582_0),.din(w_dff_A_ntG72hgR0_0),.clk(gclk));
	jdff dff_A_uYXQn4582_0(.dout(w_dff_A_28I0bMga3_0),.din(w_dff_A_uYXQn4582_0),.clk(gclk));
	jdff dff_A_28I0bMga3_0(.dout(w_dff_A_FIyxzINt4_0),.din(w_dff_A_28I0bMga3_0),.clk(gclk));
	jdff dff_A_FIyxzINt4_0(.dout(w_dff_A_dMSxsxpb2_0),.din(w_dff_A_FIyxzINt4_0),.clk(gclk));
	jdff dff_A_dMSxsxpb2_0(.dout(G478),.din(w_dff_A_dMSxsxpb2_0),.clk(gclk));
	jdff dff_A_JFXSKKkp5_1(.dout(w_dff_A_KmRG8YSZ8_0),.din(w_dff_A_JFXSKKkp5_1),.clk(gclk));
	jdff dff_A_KmRG8YSZ8_0(.dout(w_dff_A_Hmd9HzlN3_0),.din(w_dff_A_KmRG8YSZ8_0),.clk(gclk));
	jdff dff_A_Hmd9HzlN3_0(.dout(w_dff_A_cjGxqako2_0),.din(w_dff_A_Hmd9HzlN3_0),.clk(gclk));
	jdff dff_A_cjGxqako2_0(.dout(w_dff_A_tyW7NXjR8_0),.din(w_dff_A_cjGxqako2_0),.clk(gclk));
	jdff dff_A_tyW7NXjR8_0(.dout(w_dff_A_aWyQiUHD4_0),.din(w_dff_A_tyW7NXjR8_0),.clk(gclk));
	jdff dff_A_aWyQiUHD4_0(.dout(w_dff_A_CBYYRz818_0),.din(w_dff_A_aWyQiUHD4_0),.clk(gclk));
	jdff dff_A_CBYYRz818_0(.dout(w_dff_A_Rf3WrN775_0),.din(w_dff_A_CBYYRz818_0),.clk(gclk));
	jdff dff_A_Rf3WrN775_0(.dout(w_dff_A_tgxb4eBv7_0),.din(w_dff_A_Rf3WrN775_0),.clk(gclk));
	jdff dff_A_tgxb4eBv7_0(.dout(w_dff_A_astaUZVK0_0),.din(w_dff_A_tgxb4eBv7_0),.clk(gclk));
	jdff dff_A_astaUZVK0_0(.dout(w_dff_A_EbzHxp4j0_0),.din(w_dff_A_astaUZVK0_0),.clk(gclk));
	jdff dff_A_EbzHxp4j0_0(.dout(w_dff_A_TbGuQqq25_0),.din(w_dff_A_EbzHxp4j0_0),.clk(gclk));
	jdff dff_A_TbGuQqq25_0(.dout(w_dff_A_dns6CZ698_0),.din(w_dff_A_TbGuQqq25_0),.clk(gclk));
	jdff dff_A_dns6CZ698_0(.dout(w_dff_A_5nmK8d0p2_0),.din(w_dff_A_dns6CZ698_0),.clk(gclk));
	jdff dff_A_5nmK8d0p2_0(.dout(w_dff_A_OQJ8q4XR8_0),.din(w_dff_A_5nmK8d0p2_0),.clk(gclk));
	jdff dff_A_OQJ8q4XR8_0(.dout(w_dff_A_AWSAZYem2_0),.din(w_dff_A_OQJ8q4XR8_0),.clk(gclk));
	jdff dff_A_AWSAZYem2_0(.dout(w_dff_A_k3YahAFL4_0),.din(w_dff_A_AWSAZYem2_0),.clk(gclk));
	jdff dff_A_k3YahAFL4_0(.dout(w_dff_A_56F7Au5a4_0),.din(w_dff_A_k3YahAFL4_0),.clk(gclk));
	jdff dff_A_56F7Au5a4_0(.dout(w_dff_A_zlQKHLze9_0),.din(w_dff_A_56F7Au5a4_0),.clk(gclk));
	jdff dff_A_zlQKHLze9_0(.dout(w_dff_A_kxFPVAmC5_0),.din(w_dff_A_zlQKHLze9_0),.clk(gclk));
	jdff dff_A_kxFPVAmC5_0(.dout(w_dff_A_cUiNiaLE9_0),.din(w_dff_A_kxFPVAmC5_0),.clk(gclk));
	jdff dff_A_cUiNiaLE9_0(.dout(w_dff_A_LqlnNlhh8_0),.din(w_dff_A_cUiNiaLE9_0),.clk(gclk));
	jdff dff_A_LqlnNlhh8_0(.dout(w_dff_A_EoJ7s8AD2_0),.din(w_dff_A_LqlnNlhh8_0),.clk(gclk));
	jdff dff_A_EoJ7s8AD2_0(.dout(w_dff_A_XVGMf8mF1_0),.din(w_dff_A_EoJ7s8AD2_0),.clk(gclk));
	jdff dff_A_XVGMf8mF1_0(.dout(w_dff_A_xhiXXSCI6_0),.din(w_dff_A_XVGMf8mF1_0),.clk(gclk));
	jdff dff_A_xhiXXSCI6_0(.dout(w_dff_A_RsnUzjIM7_0),.din(w_dff_A_xhiXXSCI6_0),.clk(gclk));
	jdff dff_A_RsnUzjIM7_0(.dout(w_dff_A_nubtNemo2_0),.din(w_dff_A_RsnUzjIM7_0),.clk(gclk));
	jdff dff_A_nubtNemo2_0(.dout(w_dff_A_nEZtyRX62_0),.din(w_dff_A_nubtNemo2_0),.clk(gclk));
	jdff dff_A_nEZtyRX62_0(.dout(w_dff_A_ME7rmiYF4_0),.din(w_dff_A_nEZtyRX62_0),.clk(gclk));
	jdff dff_A_ME7rmiYF4_0(.dout(w_dff_A_Z058oID48_0),.din(w_dff_A_ME7rmiYF4_0),.clk(gclk));
	jdff dff_A_Z058oID48_0(.dout(w_dff_A_wOc3JKWb7_0),.din(w_dff_A_Z058oID48_0),.clk(gclk));
	jdff dff_A_wOc3JKWb7_0(.dout(w_dff_A_oIxqCI0V0_0),.din(w_dff_A_wOc3JKWb7_0),.clk(gclk));
	jdff dff_A_oIxqCI0V0_0(.dout(w_dff_A_i0LZDUdt2_0),.din(w_dff_A_oIxqCI0V0_0),.clk(gclk));
	jdff dff_A_i0LZDUdt2_0(.dout(w_dff_A_WHKvjddF5_0),.din(w_dff_A_i0LZDUdt2_0),.clk(gclk));
	jdff dff_A_WHKvjddF5_0(.dout(w_dff_A_m07byV5r5_0),.din(w_dff_A_WHKvjddF5_0),.clk(gclk));
	jdff dff_A_m07byV5r5_0(.dout(w_dff_A_0Lf6114F7_0),.din(w_dff_A_m07byV5r5_0),.clk(gclk));
	jdff dff_A_0Lf6114F7_0(.dout(w_dff_A_MEU3uGmb7_0),.din(w_dff_A_0Lf6114F7_0),.clk(gclk));
	jdff dff_A_MEU3uGmb7_0(.dout(w_dff_A_Vj3nW6U86_0),.din(w_dff_A_MEU3uGmb7_0),.clk(gclk));
	jdff dff_A_Vj3nW6U86_0(.dout(G522),.din(w_dff_A_Vj3nW6U86_0),.clk(gclk));
	jdff dff_A_158BVJfx5_2(.dout(w_dff_A_CLL2gg4d5_0),.din(w_dff_A_158BVJfx5_2),.clk(gclk));
	jdff dff_A_CLL2gg4d5_0(.dout(w_dff_A_9oE5xXgH8_0),.din(w_dff_A_CLL2gg4d5_0),.clk(gclk));
	jdff dff_A_9oE5xXgH8_0(.dout(w_dff_A_5Dm0OX310_0),.din(w_dff_A_9oE5xXgH8_0),.clk(gclk));
	jdff dff_A_5Dm0OX310_0(.dout(w_dff_A_xacIzu1s5_0),.din(w_dff_A_5Dm0OX310_0),.clk(gclk));
	jdff dff_A_xacIzu1s5_0(.dout(w_dff_A_pemjsvk11_0),.din(w_dff_A_xacIzu1s5_0),.clk(gclk));
	jdff dff_A_pemjsvk11_0(.dout(w_dff_A_VZZHPRUb7_0),.din(w_dff_A_pemjsvk11_0),.clk(gclk));
	jdff dff_A_VZZHPRUb7_0(.dout(w_dff_A_CFT6vBDo3_0),.din(w_dff_A_VZZHPRUb7_0),.clk(gclk));
	jdff dff_A_CFT6vBDo3_0(.dout(w_dff_A_b8zK4la92_0),.din(w_dff_A_CFT6vBDo3_0),.clk(gclk));
	jdff dff_A_b8zK4la92_0(.dout(w_dff_A_3Xb9YTFB0_0),.din(w_dff_A_b8zK4la92_0),.clk(gclk));
	jdff dff_A_3Xb9YTFB0_0(.dout(w_dff_A_3sKgfhgL1_0),.din(w_dff_A_3Xb9YTFB0_0),.clk(gclk));
	jdff dff_A_3sKgfhgL1_0(.dout(w_dff_A_miJLNjiY1_0),.din(w_dff_A_3sKgfhgL1_0),.clk(gclk));
	jdff dff_A_miJLNjiY1_0(.dout(w_dff_A_Ih7lLUxj2_0),.din(w_dff_A_miJLNjiY1_0),.clk(gclk));
	jdff dff_A_Ih7lLUxj2_0(.dout(w_dff_A_wZ1HvS8d8_0),.din(w_dff_A_Ih7lLUxj2_0),.clk(gclk));
	jdff dff_A_wZ1HvS8d8_0(.dout(w_dff_A_8D0Z7R2P1_0),.din(w_dff_A_wZ1HvS8d8_0),.clk(gclk));
	jdff dff_A_8D0Z7R2P1_0(.dout(w_dff_A_ku5aXqcm2_0),.din(w_dff_A_8D0Z7R2P1_0),.clk(gclk));
	jdff dff_A_ku5aXqcm2_0(.dout(w_dff_A_j4LrhcMD0_0),.din(w_dff_A_ku5aXqcm2_0),.clk(gclk));
	jdff dff_A_j4LrhcMD0_0(.dout(w_dff_A_RCMzzZ511_0),.din(w_dff_A_j4LrhcMD0_0),.clk(gclk));
	jdff dff_A_RCMzzZ511_0(.dout(w_dff_A_ZmeHSxo71_0),.din(w_dff_A_RCMzzZ511_0),.clk(gclk));
	jdff dff_A_ZmeHSxo71_0(.dout(w_dff_A_MNGIbMlA0_0),.din(w_dff_A_ZmeHSxo71_0),.clk(gclk));
	jdff dff_A_MNGIbMlA0_0(.dout(w_dff_A_EySmUv1b4_0),.din(w_dff_A_MNGIbMlA0_0),.clk(gclk));
	jdff dff_A_EySmUv1b4_0(.dout(w_dff_A_fkQkFkf26_0),.din(w_dff_A_EySmUv1b4_0),.clk(gclk));
	jdff dff_A_fkQkFkf26_0(.dout(w_dff_A_QC3yvEuU0_0),.din(w_dff_A_fkQkFkf26_0),.clk(gclk));
	jdff dff_A_QC3yvEuU0_0(.dout(w_dff_A_mOYl6UFY1_0),.din(w_dff_A_QC3yvEuU0_0),.clk(gclk));
	jdff dff_A_mOYl6UFY1_0(.dout(w_dff_A_nh36QvYs6_0),.din(w_dff_A_mOYl6UFY1_0),.clk(gclk));
	jdff dff_A_nh36QvYs6_0(.dout(w_dff_A_etqlJ6TU7_0),.din(w_dff_A_nh36QvYs6_0),.clk(gclk));
	jdff dff_A_etqlJ6TU7_0(.dout(w_dff_A_NjIgqH7Q1_0),.din(w_dff_A_etqlJ6TU7_0),.clk(gclk));
	jdff dff_A_NjIgqH7Q1_0(.dout(w_dff_A_TGmHPZnS2_0),.din(w_dff_A_NjIgqH7Q1_0),.clk(gclk));
	jdff dff_A_TGmHPZnS2_0(.dout(w_dff_A_EEN8P03i3_0),.din(w_dff_A_TGmHPZnS2_0),.clk(gclk));
	jdff dff_A_EEN8P03i3_0(.dout(w_dff_A_rl3A3UPi4_0),.din(w_dff_A_EEN8P03i3_0),.clk(gclk));
	jdff dff_A_rl3A3UPi4_0(.dout(w_dff_A_bYRWAxlR4_0),.din(w_dff_A_rl3A3UPi4_0),.clk(gclk));
	jdff dff_A_bYRWAxlR4_0(.dout(w_dff_A_o4VX0bgv8_0),.din(w_dff_A_bYRWAxlR4_0),.clk(gclk));
	jdff dff_A_o4VX0bgv8_0(.dout(w_dff_A_iRGSMRKl2_0),.din(w_dff_A_o4VX0bgv8_0),.clk(gclk));
	jdff dff_A_iRGSMRKl2_0(.dout(w_dff_A_Md8CSjuT2_0),.din(w_dff_A_iRGSMRKl2_0),.clk(gclk));
	jdff dff_A_Md8CSjuT2_0(.dout(w_dff_A_sYVzjdXt8_0),.din(w_dff_A_Md8CSjuT2_0),.clk(gclk));
	jdff dff_A_sYVzjdXt8_0(.dout(w_dff_A_J7k3LctK6_0),.din(w_dff_A_sYVzjdXt8_0),.clk(gclk));
	jdff dff_A_J7k3LctK6_0(.dout(w_dff_A_FVVC0TFo0_0),.din(w_dff_A_J7k3LctK6_0),.clk(gclk));
	jdff dff_A_FVVC0TFo0_0(.dout(w_dff_A_kWgYBNDK3_0),.din(w_dff_A_FVVC0TFo0_0),.clk(gclk));
	jdff dff_A_kWgYBNDK3_0(.dout(G402),.din(w_dff_A_kWgYBNDK3_0),.clk(gclk));
	jdff dff_A_GynMmCSi4_1(.dout(w_dff_A_vj1i6Q4W4_0),.din(w_dff_A_GynMmCSi4_1),.clk(gclk));
	jdff dff_A_vj1i6Q4W4_0(.dout(w_dff_A_9iyTVvLU4_0),.din(w_dff_A_vj1i6Q4W4_0),.clk(gclk));
	jdff dff_A_9iyTVvLU4_0(.dout(w_dff_A_BIS7cSYb4_0),.din(w_dff_A_9iyTVvLU4_0),.clk(gclk));
	jdff dff_A_BIS7cSYb4_0(.dout(w_dff_A_DSrrF1LD0_0),.din(w_dff_A_BIS7cSYb4_0),.clk(gclk));
	jdff dff_A_DSrrF1LD0_0(.dout(w_dff_A_VIcrETCE7_0),.din(w_dff_A_DSrrF1LD0_0),.clk(gclk));
	jdff dff_A_VIcrETCE7_0(.dout(w_dff_A_ZWUV3q6f1_0),.din(w_dff_A_VIcrETCE7_0),.clk(gclk));
	jdff dff_A_ZWUV3q6f1_0(.dout(w_dff_A_TJ3rlJPR7_0),.din(w_dff_A_ZWUV3q6f1_0),.clk(gclk));
	jdff dff_A_TJ3rlJPR7_0(.dout(w_dff_A_88fEcWo73_0),.din(w_dff_A_TJ3rlJPR7_0),.clk(gclk));
	jdff dff_A_88fEcWo73_0(.dout(w_dff_A_e4qr6Kim1_0),.din(w_dff_A_88fEcWo73_0),.clk(gclk));
	jdff dff_A_e4qr6Kim1_0(.dout(w_dff_A_DIRzeKGR5_0),.din(w_dff_A_e4qr6Kim1_0),.clk(gclk));
	jdff dff_A_DIRzeKGR5_0(.dout(w_dff_A_qqwVFXsz4_0),.din(w_dff_A_DIRzeKGR5_0),.clk(gclk));
	jdff dff_A_qqwVFXsz4_0(.dout(w_dff_A_xqHEpXaw2_0),.din(w_dff_A_qqwVFXsz4_0),.clk(gclk));
	jdff dff_A_xqHEpXaw2_0(.dout(w_dff_A_WY0X2efS1_0),.din(w_dff_A_xqHEpXaw2_0),.clk(gclk));
	jdff dff_A_WY0X2efS1_0(.dout(w_dff_A_hJ3ZGWct2_0),.din(w_dff_A_WY0X2efS1_0),.clk(gclk));
	jdff dff_A_hJ3ZGWct2_0(.dout(w_dff_A_nawroWYY6_0),.din(w_dff_A_hJ3ZGWct2_0),.clk(gclk));
	jdff dff_A_nawroWYY6_0(.dout(w_dff_A_aTs9Zv9f3_0),.din(w_dff_A_nawroWYY6_0),.clk(gclk));
	jdff dff_A_aTs9Zv9f3_0(.dout(w_dff_A_q8GdOi1s4_0),.din(w_dff_A_aTs9Zv9f3_0),.clk(gclk));
	jdff dff_A_q8GdOi1s4_0(.dout(w_dff_A_VvfLsch44_0),.din(w_dff_A_q8GdOi1s4_0),.clk(gclk));
	jdff dff_A_VvfLsch44_0(.dout(w_dff_A_XimVxw858_0),.din(w_dff_A_VvfLsch44_0),.clk(gclk));
	jdff dff_A_XimVxw858_0(.dout(w_dff_A_667T2w5h1_0),.din(w_dff_A_XimVxw858_0),.clk(gclk));
	jdff dff_A_667T2w5h1_0(.dout(w_dff_A_HR4KjMBJ0_0),.din(w_dff_A_667T2w5h1_0),.clk(gclk));
	jdff dff_A_HR4KjMBJ0_0(.dout(w_dff_A_0RwHo2li2_0),.din(w_dff_A_HR4KjMBJ0_0),.clk(gclk));
	jdff dff_A_0RwHo2li2_0(.dout(w_dff_A_JcJogVNy6_0),.din(w_dff_A_0RwHo2li2_0),.clk(gclk));
	jdff dff_A_JcJogVNy6_0(.dout(w_dff_A_YAUbcyV69_0),.din(w_dff_A_JcJogVNy6_0),.clk(gclk));
	jdff dff_A_YAUbcyV69_0(.dout(w_dff_A_Gs4iSEBu7_0),.din(w_dff_A_YAUbcyV69_0),.clk(gclk));
	jdff dff_A_Gs4iSEBu7_0(.dout(w_dff_A_Pkj2Y5nd5_0),.din(w_dff_A_Gs4iSEBu7_0),.clk(gclk));
	jdff dff_A_Pkj2Y5nd5_0(.dout(w_dff_A_WFMLinim1_0),.din(w_dff_A_Pkj2Y5nd5_0),.clk(gclk));
	jdff dff_A_WFMLinim1_0(.dout(w_dff_A_RcIwekHA4_0),.din(w_dff_A_WFMLinim1_0),.clk(gclk));
	jdff dff_A_RcIwekHA4_0(.dout(w_dff_A_0xaU0Cuh0_0),.din(w_dff_A_RcIwekHA4_0),.clk(gclk));
	jdff dff_A_0xaU0Cuh0_0(.dout(w_dff_A_HTAEPPW28_0),.din(w_dff_A_0xaU0Cuh0_0),.clk(gclk));
	jdff dff_A_HTAEPPW28_0(.dout(w_dff_A_Rdlf2Vif7_0),.din(w_dff_A_HTAEPPW28_0),.clk(gclk));
	jdff dff_A_Rdlf2Vif7_0(.dout(w_dff_A_PXw3ExlL2_0),.din(w_dff_A_Rdlf2Vif7_0),.clk(gclk));
	jdff dff_A_PXw3ExlL2_0(.dout(w_dff_A_aCpWcBb56_0),.din(w_dff_A_PXw3ExlL2_0),.clk(gclk));
	jdff dff_A_aCpWcBb56_0(.dout(w_dff_A_CpcPe3Hn7_0),.din(w_dff_A_aCpWcBb56_0),.clk(gclk));
	jdff dff_A_CpcPe3Hn7_0(.dout(w_dff_A_ao8jql5i9_0),.din(w_dff_A_CpcPe3Hn7_0),.clk(gclk));
	jdff dff_A_ao8jql5i9_0(.dout(G404),.din(w_dff_A_ao8jql5i9_0),.clk(gclk));
	jdff dff_A_QtSapZun2_1(.dout(w_dff_A_Ni8tMVZk0_0),.din(w_dff_A_QtSapZun2_1),.clk(gclk));
	jdff dff_A_Ni8tMVZk0_0(.dout(w_dff_A_Yr13wJqq8_0),.din(w_dff_A_Ni8tMVZk0_0),.clk(gclk));
	jdff dff_A_Yr13wJqq8_0(.dout(w_dff_A_5HzB6MDS0_0),.din(w_dff_A_Yr13wJqq8_0),.clk(gclk));
	jdff dff_A_5HzB6MDS0_0(.dout(w_dff_A_Mmh4FKkW1_0),.din(w_dff_A_5HzB6MDS0_0),.clk(gclk));
	jdff dff_A_Mmh4FKkW1_0(.dout(w_dff_A_NUUm0Deu7_0),.din(w_dff_A_Mmh4FKkW1_0),.clk(gclk));
	jdff dff_A_NUUm0Deu7_0(.dout(w_dff_A_Eg47cOYr6_0),.din(w_dff_A_NUUm0Deu7_0),.clk(gclk));
	jdff dff_A_Eg47cOYr6_0(.dout(w_dff_A_DHI7KS9M8_0),.din(w_dff_A_Eg47cOYr6_0),.clk(gclk));
	jdff dff_A_DHI7KS9M8_0(.dout(w_dff_A_vF4yevS25_0),.din(w_dff_A_DHI7KS9M8_0),.clk(gclk));
	jdff dff_A_vF4yevS25_0(.dout(w_dff_A_a2Re9Td98_0),.din(w_dff_A_vF4yevS25_0),.clk(gclk));
	jdff dff_A_a2Re9Td98_0(.dout(w_dff_A_rtUhi4762_0),.din(w_dff_A_a2Re9Td98_0),.clk(gclk));
	jdff dff_A_rtUhi4762_0(.dout(w_dff_A_9rU4JBHW4_0),.din(w_dff_A_rtUhi4762_0),.clk(gclk));
	jdff dff_A_9rU4JBHW4_0(.dout(w_dff_A_EbPVg9GJ5_0),.din(w_dff_A_9rU4JBHW4_0),.clk(gclk));
	jdff dff_A_EbPVg9GJ5_0(.dout(w_dff_A_tXaxjFRS5_0),.din(w_dff_A_EbPVg9GJ5_0),.clk(gclk));
	jdff dff_A_tXaxjFRS5_0(.dout(w_dff_A_1etpoojM9_0),.din(w_dff_A_tXaxjFRS5_0),.clk(gclk));
	jdff dff_A_1etpoojM9_0(.dout(w_dff_A_ffGf5HGF1_0),.din(w_dff_A_1etpoojM9_0),.clk(gclk));
	jdff dff_A_ffGf5HGF1_0(.dout(w_dff_A_mdA6x57w6_0),.din(w_dff_A_ffGf5HGF1_0),.clk(gclk));
	jdff dff_A_mdA6x57w6_0(.dout(w_dff_A_pM1xlMzH9_0),.din(w_dff_A_mdA6x57w6_0),.clk(gclk));
	jdff dff_A_pM1xlMzH9_0(.dout(w_dff_A_BQVMZrRw0_0),.din(w_dff_A_pM1xlMzH9_0),.clk(gclk));
	jdff dff_A_BQVMZrRw0_0(.dout(w_dff_A_qB8ix4dM5_0),.din(w_dff_A_BQVMZrRw0_0),.clk(gclk));
	jdff dff_A_qB8ix4dM5_0(.dout(w_dff_A_UckGQ84b8_0),.din(w_dff_A_qB8ix4dM5_0),.clk(gclk));
	jdff dff_A_UckGQ84b8_0(.dout(w_dff_A_3DyiCViY7_0),.din(w_dff_A_UckGQ84b8_0),.clk(gclk));
	jdff dff_A_3DyiCViY7_0(.dout(w_dff_A_lI64x69H9_0),.din(w_dff_A_3DyiCViY7_0),.clk(gclk));
	jdff dff_A_lI64x69H9_0(.dout(w_dff_A_xABE00sC0_0),.din(w_dff_A_lI64x69H9_0),.clk(gclk));
	jdff dff_A_xABE00sC0_0(.dout(w_dff_A_9ifPF6r31_0),.din(w_dff_A_xABE00sC0_0),.clk(gclk));
	jdff dff_A_9ifPF6r31_0(.dout(w_dff_A_aUxtXqlF6_0),.din(w_dff_A_9ifPF6r31_0),.clk(gclk));
	jdff dff_A_aUxtXqlF6_0(.dout(w_dff_A_rsRX30xy1_0),.din(w_dff_A_aUxtXqlF6_0),.clk(gclk));
	jdff dff_A_rsRX30xy1_0(.dout(w_dff_A_FHMB4Ax24_0),.din(w_dff_A_rsRX30xy1_0),.clk(gclk));
	jdff dff_A_FHMB4Ax24_0(.dout(w_dff_A_4XAdbL8E9_0),.din(w_dff_A_FHMB4Ax24_0),.clk(gclk));
	jdff dff_A_4XAdbL8E9_0(.dout(w_dff_A_61Kaltr52_0),.din(w_dff_A_4XAdbL8E9_0),.clk(gclk));
	jdff dff_A_61Kaltr52_0(.dout(w_dff_A_xLSKHv535_0),.din(w_dff_A_61Kaltr52_0),.clk(gclk));
	jdff dff_A_xLSKHv535_0(.dout(w_dff_A_QUvfsMu10_0),.din(w_dff_A_xLSKHv535_0),.clk(gclk));
	jdff dff_A_QUvfsMu10_0(.dout(w_dff_A_k9lcU8oD2_0),.din(w_dff_A_QUvfsMu10_0),.clk(gclk));
	jdff dff_A_k9lcU8oD2_0(.dout(w_dff_A_SeTd8ZPF5_0),.din(w_dff_A_k9lcU8oD2_0),.clk(gclk));
	jdff dff_A_SeTd8ZPF5_0(.dout(w_dff_A_G0pdch835_0),.din(w_dff_A_SeTd8ZPF5_0),.clk(gclk));
	jdff dff_A_G0pdch835_0(.dout(w_dff_A_1efeAtYx5_0),.din(w_dff_A_G0pdch835_0),.clk(gclk));
	jdff dff_A_1efeAtYx5_0(.dout(G406),.din(w_dff_A_1efeAtYx5_0),.clk(gclk));
	jdff dff_A_iYRibRUl1_1(.dout(w_dff_A_DtfApZ644_0),.din(w_dff_A_iYRibRUl1_1),.clk(gclk));
	jdff dff_A_DtfApZ644_0(.dout(w_dff_A_spBeFz7Q1_0),.din(w_dff_A_DtfApZ644_0),.clk(gclk));
	jdff dff_A_spBeFz7Q1_0(.dout(w_dff_A_zggI7YUb0_0),.din(w_dff_A_spBeFz7Q1_0),.clk(gclk));
	jdff dff_A_zggI7YUb0_0(.dout(w_dff_A_uqnBezBm3_0),.din(w_dff_A_zggI7YUb0_0),.clk(gclk));
	jdff dff_A_uqnBezBm3_0(.dout(w_dff_A_4M7CeSQk3_0),.din(w_dff_A_uqnBezBm3_0),.clk(gclk));
	jdff dff_A_4M7CeSQk3_0(.dout(w_dff_A_DJ6AhKP72_0),.din(w_dff_A_4M7CeSQk3_0),.clk(gclk));
	jdff dff_A_DJ6AhKP72_0(.dout(w_dff_A_BFztI4Bh1_0),.din(w_dff_A_DJ6AhKP72_0),.clk(gclk));
	jdff dff_A_BFztI4Bh1_0(.dout(w_dff_A_cqJA7KfR5_0),.din(w_dff_A_BFztI4Bh1_0),.clk(gclk));
	jdff dff_A_cqJA7KfR5_0(.dout(w_dff_A_zsGQi5M20_0),.din(w_dff_A_cqJA7KfR5_0),.clk(gclk));
	jdff dff_A_zsGQi5M20_0(.dout(w_dff_A_UlVdO9237_0),.din(w_dff_A_zsGQi5M20_0),.clk(gclk));
	jdff dff_A_UlVdO9237_0(.dout(w_dff_A_wUk8zebQ7_0),.din(w_dff_A_UlVdO9237_0),.clk(gclk));
	jdff dff_A_wUk8zebQ7_0(.dout(w_dff_A_pmgoKI551_0),.din(w_dff_A_wUk8zebQ7_0),.clk(gclk));
	jdff dff_A_pmgoKI551_0(.dout(w_dff_A_rM84gTKC2_0),.din(w_dff_A_pmgoKI551_0),.clk(gclk));
	jdff dff_A_rM84gTKC2_0(.dout(w_dff_A_HrFf6mQx3_0),.din(w_dff_A_rM84gTKC2_0),.clk(gclk));
	jdff dff_A_HrFf6mQx3_0(.dout(w_dff_A_YfYXewFo9_0),.din(w_dff_A_HrFf6mQx3_0),.clk(gclk));
	jdff dff_A_YfYXewFo9_0(.dout(w_dff_A_r2MSjyaJ9_0),.din(w_dff_A_YfYXewFo9_0),.clk(gclk));
	jdff dff_A_r2MSjyaJ9_0(.dout(w_dff_A_jcBqriGy5_0),.din(w_dff_A_r2MSjyaJ9_0),.clk(gclk));
	jdff dff_A_jcBqriGy5_0(.dout(w_dff_A_jwfMJWPO3_0),.din(w_dff_A_jcBqriGy5_0),.clk(gclk));
	jdff dff_A_jwfMJWPO3_0(.dout(w_dff_A_l0XUuEHd6_0),.din(w_dff_A_jwfMJWPO3_0),.clk(gclk));
	jdff dff_A_l0XUuEHd6_0(.dout(w_dff_A_TLmp5ND70_0),.din(w_dff_A_l0XUuEHd6_0),.clk(gclk));
	jdff dff_A_TLmp5ND70_0(.dout(w_dff_A_CQbFnLfr6_0),.din(w_dff_A_TLmp5ND70_0),.clk(gclk));
	jdff dff_A_CQbFnLfr6_0(.dout(w_dff_A_SKbKcetk1_0),.din(w_dff_A_CQbFnLfr6_0),.clk(gclk));
	jdff dff_A_SKbKcetk1_0(.dout(w_dff_A_L6IqURT07_0),.din(w_dff_A_SKbKcetk1_0),.clk(gclk));
	jdff dff_A_L6IqURT07_0(.dout(w_dff_A_1RlyPywy1_0),.din(w_dff_A_L6IqURT07_0),.clk(gclk));
	jdff dff_A_1RlyPywy1_0(.dout(w_dff_A_YM7WnGRF9_0),.din(w_dff_A_1RlyPywy1_0),.clk(gclk));
	jdff dff_A_YM7WnGRF9_0(.dout(w_dff_A_EIe6eaZE5_0),.din(w_dff_A_YM7WnGRF9_0),.clk(gclk));
	jdff dff_A_EIe6eaZE5_0(.dout(w_dff_A_lslajPSF1_0),.din(w_dff_A_EIe6eaZE5_0),.clk(gclk));
	jdff dff_A_lslajPSF1_0(.dout(w_dff_A_e8ZfvcSP1_0),.din(w_dff_A_lslajPSF1_0),.clk(gclk));
	jdff dff_A_e8ZfvcSP1_0(.dout(w_dff_A_9SlHEK3L8_0),.din(w_dff_A_e8ZfvcSP1_0),.clk(gclk));
	jdff dff_A_9SlHEK3L8_0(.dout(w_dff_A_CIp6Cpqx5_0),.din(w_dff_A_9SlHEK3L8_0),.clk(gclk));
	jdff dff_A_CIp6Cpqx5_0(.dout(w_dff_A_c906w5Tr0_0),.din(w_dff_A_CIp6Cpqx5_0),.clk(gclk));
	jdff dff_A_c906w5Tr0_0(.dout(w_dff_A_KzHKDdGE1_0),.din(w_dff_A_c906w5Tr0_0),.clk(gclk));
	jdff dff_A_KzHKDdGE1_0(.dout(w_dff_A_UBBuUfUc6_0),.din(w_dff_A_KzHKDdGE1_0),.clk(gclk));
	jdff dff_A_UBBuUfUc6_0(.dout(w_dff_A_6wW9gcSs6_0),.din(w_dff_A_UBBuUfUc6_0),.clk(gclk));
	jdff dff_A_6wW9gcSs6_0(.dout(w_dff_A_kJxTHZ8z4_0),.din(w_dff_A_6wW9gcSs6_0),.clk(gclk));
	jdff dff_A_kJxTHZ8z4_0(.dout(G408),.din(w_dff_A_kJxTHZ8z4_0),.clk(gclk));
	jdff dff_A_tsINoMcR6_1(.dout(w_dff_A_XIOyU0On8_0),.din(w_dff_A_tsINoMcR6_1),.clk(gclk));
	jdff dff_A_XIOyU0On8_0(.dout(w_dff_A_DKq3e43b4_0),.din(w_dff_A_XIOyU0On8_0),.clk(gclk));
	jdff dff_A_DKq3e43b4_0(.dout(w_dff_A_czLKlFlI1_0),.din(w_dff_A_DKq3e43b4_0),.clk(gclk));
	jdff dff_A_czLKlFlI1_0(.dout(w_dff_A_kneUDeSo9_0),.din(w_dff_A_czLKlFlI1_0),.clk(gclk));
	jdff dff_A_kneUDeSo9_0(.dout(w_dff_A_asRLFjFv8_0),.din(w_dff_A_kneUDeSo9_0),.clk(gclk));
	jdff dff_A_asRLFjFv8_0(.dout(w_dff_A_dmSL62r85_0),.din(w_dff_A_asRLFjFv8_0),.clk(gclk));
	jdff dff_A_dmSL62r85_0(.dout(w_dff_A_WGYuRayh3_0),.din(w_dff_A_dmSL62r85_0),.clk(gclk));
	jdff dff_A_WGYuRayh3_0(.dout(w_dff_A_t6Yo5nF36_0),.din(w_dff_A_WGYuRayh3_0),.clk(gclk));
	jdff dff_A_t6Yo5nF36_0(.dout(w_dff_A_ff0bDvq20_0),.din(w_dff_A_t6Yo5nF36_0),.clk(gclk));
	jdff dff_A_ff0bDvq20_0(.dout(w_dff_A_YprfJ5oT0_0),.din(w_dff_A_ff0bDvq20_0),.clk(gclk));
	jdff dff_A_YprfJ5oT0_0(.dout(w_dff_A_joTFkHDa9_0),.din(w_dff_A_YprfJ5oT0_0),.clk(gclk));
	jdff dff_A_joTFkHDa9_0(.dout(w_dff_A_e3zsG0NN4_0),.din(w_dff_A_joTFkHDa9_0),.clk(gclk));
	jdff dff_A_e3zsG0NN4_0(.dout(w_dff_A_GiAcPx413_0),.din(w_dff_A_e3zsG0NN4_0),.clk(gclk));
	jdff dff_A_GiAcPx413_0(.dout(w_dff_A_dK4zzXzr1_0),.din(w_dff_A_GiAcPx413_0),.clk(gclk));
	jdff dff_A_dK4zzXzr1_0(.dout(w_dff_A_Ht2WsStZ1_0),.din(w_dff_A_dK4zzXzr1_0),.clk(gclk));
	jdff dff_A_Ht2WsStZ1_0(.dout(w_dff_A_cQMboIm72_0),.din(w_dff_A_Ht2WsStZ1_0),.clk(gclk));
	jdff dff_A_cQMboIm72_0(.dout(w_dff_A_8ON1Eriq9_0),.din(w_dff_A_cQMboIm72_0),.clk(gclk));
	jdff dff_A_8ON1Eriq9_0(.dout(w_dff_A_v8lLApdP1_0),.din(w_dff_A_8ON1Eriq9_0),.clk(gclk));
	jdff dff_A_v8lLApdP1_0(.dout(w_dff_A_zuxOMWEg1_0),.din(w_dff_A_v8lLApdP1_0),.clk(gclk));
	jdff dff_A_zuxOMWEg1_0(.dout(w_dff_A_XM4UcsAw0_0),.din(w_dff_A_zuxOMWEg1_0),.clk(gclk));
	jdff dff_A_XM4UcsAw0_0(.dout(w_dff_A_2hzFlrvq5_0),.din(w_dff_A_XM4UcsAw0_0),.clk(gclk));
	jdff dff_A_2hzFlrvq5_0(.dout(w_dff_A_MfntoeHo8_0),.din(w_dff_A_2hzFlrvq5_0),.clk(gclk));
	jdff dff_A_MfntoeHo8_0(.dout(w_dff_A_sNo8GWjO7_0),.din(w_dff_A_MfntoeHo8_0),.clk(gclk));
	jdff dff_A_sNo8GWjO7_0(.dout(w_dff_A_gQqToHrd4_0),.din(w_dff_A_sNo8GWjO7_0),.clk(gclk));
	jdff dff_A_gQqToHrd4_0(.dout(w_dff_A_dmv0xlOx5_0),.din(w_dff_A_gQqToHrd4_0),.clk(gclk));
	jdff dff_A_dmv0xlOx5_0(.dout(w_dff_A_Axk2z5rC2_0),.din(w_dff_A_dmv0xlOx5_0),.clk(gclk));
	jdff dff_A_Axk2z5rC2_0(.dout(w_dff_A_YnNXsQSi6_0),.din(w_dff_A_Axk2z5rC2_0),.clk(gclk));
	jdff dff_A_YnNXsQSi6_0(.dout(w_dff_A_HYgM8sFp3_0),.din(w_dff_A_YnNXsQSi6_0),.clk(gclk));
	jdff dff_A_HYgM8sFp3_0(.dout(w_dff_A_4jlBtAG66_0),.din(w_dff_A_HYgM8sFp3_0),.clk(gclk));
	jdff dff_A_4jlBtAG66_0(.dout(w_dff_A_qu88kCpS4_0),.din(w_dff_A_4jlBtAG66_0),.clk(gclk));
	jdff dff_A_qu88kCpS4_0(.dout(w_dff_A_vZjIRnTp8_0),.din(w_dff_A_qu88kCpS4_0),.clk(gclk));
	jdff dff_A_vZjIRnTp8_0(.dout(w_dff_A_YBpAlVzF8_0),.din(w_dff_A_vZjIRnTp8_0),.clk(gclk));
	jdff dff_A_YBpAlVzF8_0(.dout(w_dff_A_wUcfwBcW0_0),.din(w_dff_A_YBpAlVzF8_0),.clk(gclk));
	jdff dff_A_wUcfwBcW0_0(.dout(w_dff_A_97LBmKt26_0),.din(w_dff_A_wUcfwBcW0_0),.clk(gclk));
	jdff dff_A_97LBmKt26_0(.dout(w_dff_A_E8Kfagdu4_0),.din(w_dff_A_97LBmKt26_0),.clk(gclk));
	jdff dff_A_E8Kfagdu4_0(.dout(G410),.din(w_dff_A_E8Kfagdu4_0),.clk(gclk));
	jdff dff_A_qBosUjhi3_1(.dout(w_dff_A_XmgoDoCt4_0),.din(w_dff_A_qBosUjhi3_1),.clk(gclk));
	jdff dff_A_XmgoDoCt4_0(.dout(w_dff_A_itObX5ox0_0),.din(w_dff_A_XmgoDoCt4_0),.clk(gclk));
	jdff dff_A_itObX5ox0_0(.dout(w_dff_A_Rpp4e2bC3_0),.din(w_dff_A_itObX5ox0_0),.clk(gclk));
	jdff dff_A_Rpp4e2bC3_0(.dout(w_dff_A_lTkrdVcb8_0),.din(w_dff_A_Rpp4e2bC3_0),.clk(gclk));
	jdff dff_A_lTkrdVcb8_0(.dout(w_dff_A_D5p6PecJ3_0),.din(w_dff_A_lTkrdVcb8_0),.clk(gclk));
	jdff dff_A_D5p6PecJ3_0(.dout(w_dff_A_JXSZ5SvE0_0),.din(w_dff_A_D5p6PecJ3_0),.clk(gclk));
	jdff dff_A_JXSZ5SvE0_0(.dout(w_dff_A_3Z2f4XkW7_0),.din(w_dff_A_JXSZ5SvE0_0),.clk(gclk));
	jdff dff_A_3Z2f4XkW7_0(.dout(w_dff_A_A9OrukCD7_0),.din(w_dff_A_3Z2f4XkW7_0),.clk(gclk));
	jdff dff_A_A9OrukCD7_0(.dout(w_dff_A_NAYmCd8j7_0),.din(w_dff_A_A9OrukCD7_0),.clk(gclk));
	jdff dff_A_NAYmCd8j7_0(.dout(w_dff_A_xupyWn3O3_0),.din(w_dff_A_NAYmCd8j7_0),.clk(gclk));
	jdff dff_A_xupyWn3O3_0(.dout(w_dff_A_H4RuCvSp8_0),.din(w_dff_A_xupyWn3O3_0),.clk(gclk));
	jdff dff_A_H4RuCvSp8_0(.dout(w_dff_A_zZ1EwvVA0_0),.din(w_dff_A_H4RuCvSp8_0),.clk(gclk));
	jdff dff_A_zZ1EwvVA0_0(.dout(w_dff_A_czCWPgKP9_0),.din(w_dff_A_zZ1EwvVA0_0),.clk(gclk));
	jdff dff_A_czCWPgKP9_0(.dout(w_dff_A_xNdcvHzM6_0),.din(w_dff_A_czCWPgKP9_0),.clk(gclk));
	jdff dff_A_xNdcvHzM6_0(.dout(w_dff_A_j87HSMIm3_0),.din(w_dff_A_xNdcvHzM6_0),.clk(gclk));
	jdff dff_A_j87HSMIm3_0(.dout(w_dff_A_GmbMW3xD9_0),.din(w_dff_A_j87HSMIm3_0),.clk(gclk));
	jdff dff_A_GmbMW3xD9_0(.dout(w_dff_A_C18XUQQa7_0),.din(w_dff_A_GmbMW3xD9_0),.clk(gclk));
	jdff dff_A_C18XUQQa7_0(.dout(w_dff_A_naa32m2T6_0),.din(w_dff_A_C18XUQQa7_0),.clk(gclk));
	jdff dff_A_naa32m2T6_0(.dout(w_dff_A_cOfx9NFv1_0),.din(w_dff_A_naa32m2T6_0),.clk(gclk));
	jdff dff_A_cOfx9NFv1_0(.dout(w_dff_A_4hpYc9fY4_0),.din(w_dff_A_cOfx9NFv1_0),.clk(gclk));
	jdff dff_A_4hpYc9fY4_0(.dout(w_dff_A_XsJpSv5p8_0),.din(w_dff_A_4hpYc9fY4_0),.clk(gclk));
	jdff dff_A_XsJpSv5p8_0(.dout(w_dff_A_fqUaLZyf4_0),.din(w_dff_A_XsJpSv5p8_0),.clk(gclk));
	jdff dff_A_fqUaLZyf4_0(.dout(w_dff_A_8RZ7vtGk9_0),.din(w_dff_A_fqUaLZyf4_0),.clk(gclk));
	jdff dff_A_8RZ7vtGk9_0(.dout(w_dff_A_ODlXNWHL3_0),.din(w_dff_A_8RZ7vtGk9_0),.clk(gclk));
	jdff dff_A_ODlXNWHL3_0(.dout(w_dff_A_4swP6WIa2_0),.din(w_dff_A_ODlXNWHL3_0),.clk(gclk));
	jdff dff_A_4swP6WIa2_0(.dout(w_dff_A_d6Mo7nOM4_0),.din(w_dff_A_4swP6WIa2_0),.clk(gclk));
	jdff dff_A_d6Mo7nOM4_0(.dout(w_dff_A_KTfYlTgG4_0),.din(w_dff_A_d6Mo7nOM4_0),.clk(gclk));
	jdff dff_A_KTfYlTgG4_0(.dout(w_dff_A_Zyw4Hh4c6_0),.din(w_dff_A_KTfYlTgG4_0),.clk(gclk));
	jdff dff_A_Zyw4Hh4c6_0(.dout(w_dff_A_n2kFEPZK1_0),.din(w_dff_A_Zyw4Hh4c6_0),.clk(gclk));
	jdff dff_A_n2kFEPZK1_0(.dout(w_dff_A_aJ1zcPEv6_0),.din(w_dff_A_n2kFEPZK1_0),.clk(gclk));
	jdff dff_A_aJ1zcPEv6_0(.dout(w_dff_A_6irygS6R2_0),.din(w_dff_A_aJ1zcPEv6_0),.clk(gclk));
	jdff dff_A_6irygS6R2_0(.dout(w_dff_A_bolcnoIS3_0),.din(w_dff_A_6irygS6R2_0),.clk(gclk));
	jdff dff_A_bolcnoIS3_0(.dout(w_dff_A_uSEjDQWZ8_0),.din(w_dff_A_bolcnoIS3_0),.clk(gclk));
	jdff dff_A_uSEjDQWZ8_0(.dout(w_dff_A_KL8TYi5m6_0),.din(w_dff_A_uSEjDQWZ8_0),.clk(gclk));
	jdff dff_A_KL8TYi5m6_0(.dout(w_dff_A_kQwDryEX1_0),.din(w_dff_A_KL8TYi5m6_0),.clk(gclk));
	jdff dff_A_kQwDryEX1_0(.dout(w_dff_A_xbTcNRte5_0),.din(w_dff_A_kQwDryEX1_0),.clk(gclk));
	jdff dff_A_xbTcNRte5_0(.dout(w_dff_A_lAwUlNW61_0),.din(w_dff_A_xbTcNRte5_0),.clk(gclk));
	jdff dff_A_lAwUlNW61_0(.dout(G432),.din(w_dff_A_lAwUlNW61_0),.clk(gclk));
	jdff dff_A_7CPkUKba1_1(.dout(w_dff_A_hFHRnq6W9_0),.din(w_dff_A_7CPkUKba1_1),.clk(gclk));
	jdff dff_A_hFHRnq6W9_0(.dout(w_dff_A_cRkVY68A8_0),.din(w_dff_A_hFHRnq6W9_0),.clk(gclk));
	jdff dff_A_cRkVY68A8_0(.dout(w_dff_A_IwjzF4j26_0),.din(w_dff_A_cRkVY68A8_0),.clk(gclk));
	jdff dff_A_IwjzF4j26_0(.dout(w_dff_A_JdS5G9fi0_0),.din(w_dff_A_IwjzF4j26_0),.clk(gclk));
	jdff dff_A_JdS5G9fi0_0(.dout(w_dff_A_fOQ4OWmk6_0),.din(w_dff_A_JdS5G9fi0_0),.clk(gclk));
	jdff dff_A_fOQ4OWmk6_0(.dout(w_dff_A_mLoOTjCq3_0),.din(w_dff_A_fOQ4OWmk6_0),.clk(gclk));
	jdff dff_A_mLoOTjCq3_0(.dout(w_dff_A_HsuMZptG0_0),.din(w_dff_A_mLoOTjCq3_0),.clk(gclk));
	jdff dff_A_HsuMZptG0_0(.dout(w_dff_A_ND3CZ08G8_0),.din(w_dff_A_HsuMZptG0_0),.clk(gclk));
	jdff dff_A_ND3CZ08G8_0(.dout(w_dff_A_9BvbREtT2_0),.din(w_dff_A_ND3CZ08G8_0),.clk(gclk));
	jdff dff_A_9BvbREtT2_0(.dout(w_dff_A_a4PKNzHV1_0),.din(w_dff_A_9BvbREtT2_0),.clk(gclk));
	jdff dff_A_a4PKNzHV1_0(.dout(w_dff_A_5NBegsxh8_0),.din(w_dff_A_a4PKNzHV1_0),.clk(gclk));
	jdff dff_A_5NBegsxh8_0(.dout(w_dff_A_dF4jaW3N3_0),.din(w_dff_A_5NBegsxh8_0),.clk(gclk));
	jdff dff_A_dF4jaW3N3_0(.dout(w_dff_A_99JjSqbQ1_0),.din(w_dff_A_dF4jaW3N3_0),.clk(gclk));
	jdff dff_A_99JjSqbQ1_0(.dout(w_dff_A_p2BmPM2V6_0),.din(w_dff_A_99JjSqbQ1_0),.clk(gclk));
	jdff dff_A_p2BmPM2V6_0(.dout(w_dff_A_4ZozXwag7_0),.din(w_dff_A_p2BmPM2V6_0),.clk(gclk));
	jdff dff_A_4ZozXwag7_0(.dout(w_dff_A_htkz3Bcv2_0),.din(w_dff_A_4ZozXwag7_0),.clk(gclk));
	jdff dff_A_htkz3Bcv2_0(.dout(w_dff_A_btiXgu8q3_0),.din(w_dff_A_htkz3Bcv2_0),.clk(gclk));
	jdff dff_A_btiXgu8q3_0(.dout(w_dff_A_FnFL6dh00_0),.din(w_dff_A_btiXgu8q3_0),.clk(gclk));
	jdff dff_A_FnFL6dh00_0(.dout(w_dff_A_afGZXWsr7_0),.din(w_dff_A_FnFL6dh00_0),.clk(gclk));
	jdff dff_A_afGZXWsr7_0(.dout(w_dff_A_v2n8Ng6n3_0),.din(w_dff_A_afGZXWsr7_0),.clk(gclk));
	jdff dff_A_v2n8Ng6n3_0(.dout(w_dff_A_d2BlWLgO1_0),.din(w_dff_A_v2n8Ng6n3_0),.clk(gclk));
	jdff dff_A_d2BlWLgO1_0(.dout(w_dff_A_0Q0zobza8_0),.din(w_dff_A_d2BlWLgO1_0),.clk(gclk));
	jdff dff_A_0Q0zobza8_0(.dout(w_dff_A_bgYQnZzi9_0),.din(w_dff_A_0Q0zobza8_0),.clk(gclk));
	jdff dff_A_bgYQnZzi9_0(.dout(w_dff_A_5H3xuNUW5_0),.din(w_dff_A_bgYQnZzi9_0),.clk(gclk));
	jdff dff_A_5H3xuNUW5_0(.dout(w_dff_A_S7AHO3mo4_0),.din(w_dff_A_5H3xuNUW5_0),.clk(gclk));
	jdff dff_A_S7AHO3mo4_0(.dout(w_dff_A_jtWoDO2h5_0),.din(w_dff_A_S7AHO3mo4_0),.clk(gclk));
	jdff dff_A_jtWoDO2h5_0(.dout(w_dff_A_gBOFoBxy4_0),.din(w_dff_A_jtWoDO2h5_0),.clk(gclk));
	jdff dff_A_gBOFoBxy4_0(.dout(w_dff_A_RhFHycWi4_0),.din(w_dff_A_gBOFoBxy4_0),.clk(gclk));
	jdff dff_A_RhFHycWi4_0(.dout(w_dff_A_DT78MEPQ2_0),.din(w_dff_A_RhFHycWi4_0),.clk(gclk));
	jdff dff_A_DT78MEPQ2_0(.dout(w_dff_A_Oc6JN0xg0_0),.din(w_dff_A_DT78MEPQ2_0),.clk(gclk));
	jdff dff_A_Oc6JN0xg0_0(.dout(w_dff_A_HdxBD7nt4_0),.din(w_dff_A_Oc6JN0xg0_0),.clk(gclk));
	jdff dff_A_HdxBD7nt4_0(.dout(w_dff_A_bInwR5Tk5_0),.din(w_dff_A_HdxBD7nt4_0),.clk(gclk));
	jdff dff_A_bInwR5Tk5_0(.dout(w_dff_A_JFFF6dnL9_0),.din(w_dff_A_bInwR5Tk5_0),.clk(gclk));
	jdff dff_A_JFFF6dnL9_0(.dout(w_dff_A_xooZ55Ga8_0),.din(w_dff_A_JFFF6dnL9_0),.clk(gclk));
	jdff dff_A_xooZ55Ga8_0(.dout(w_dff_A_A4jbgDlv0_0),.din(w_dff_A_xooZ55Ga8_0),.clk(gclk));
	jdff dff_A_A4jbgDlv0_0(.dout(w_dff_A_GgnUw7223_0),.din(w_dff_A_A4jbgDlv0_0),.clk(gclk));
	jdff dff_A_GgnUw7223_0(.dout(w_dff_A_DK5nqAm15_0),.din(w_dff_A_GgnUw7223_0),.clk(gclk));
	jdff dff_A_DK5nqAm15_0(.dout(G446),.din(w_dff_A_DK5nqAm15_0),.clk(gclk));
	jdff dff_A_ssThCr5Y4_2(.dout(w_dff_A_M4P5kbJ74_0),.din(w_dff_A_ssThCr5Y4_2),.clk(gclk));
	jdff dff_A_M4P5kbJ74_0(.dout(w_dff_A_jl8WAa2z7_0),.din(w_dff_A_M4P5kbJ74_0),.clk(gclk));
	jdff dff_A_jl8WAa2z7_0(.dout(w_dff_A_5NHkHYdl1_0),.din(w_dff_A_jl8WAa2z7_0),.clk(gclk));
	jdff dff_A_5NHkHYdl1_0(.dout(w_dff_A_p1QNopHh9_0),.din(w_dff_A_5NHkHYdl1_0),.clk(gclk));
	jdff dff_A_p1QNopHh9_0(.dout(w_dff_A_CKsYa0bN9_0),.din(w_dff_A_p1QNopHh9_0),.clk(gclk));
	jdff dff_A_CKsYa0bN9_0(.dout(w_dff_A_fUcmldH32_0),.din(w_dff_A_CKsYa0bN9_0),.clk(gclk));
	jdff dff_A_fUcmldH32_0(.dout(w_dff_A_YXJAhgpv8_0),.din(w_dff_A_fUcmldH32_0),.clk(gclk));
	jdff dff_A_YXJAhgpv8_0(.dout(w_dff_A_bw2fKbEw5_0),.din(w_dff_A_YXJAhgpv8_0),.clk(gclk));
	jdff dff_A_bw2fKbEw5_0(.dout(w_dff_A_FJJLuoSa8_0),.din(w_dff_A_bw2fKbEw5_0),.clk(gclk));
	jdff dff_A_FJJLuoSa8_0(.dout(w_dff_A_o7Hz3tdQ5_0),.din(w_dff_A_FJJLuoSa8_0),.clk(gclk));
	jdff dff_A_o7Hz3tdQ5_0(.dout(w_dff_A_kzHlWNOg3_0),.din(w_dff_A_o7Hz3tdQ5_0),.clk(gclk));
	jdff dff_A_kzHlWNOg3_0(.dout(w_dff_A_PUqeC5lp1_0),.din(w_dff_A_kzHlWNOg3_0),.clk(gclk));
	jdff dff_A_PUqeC5lp1_0(.dout(w_dff_A_P07lZhrt0_0),.din(w_dff_A_PUqeC5lp1_0),.clk(gclk));
	jdff dff_A_P07lZhrt0_0(.dout(w_dff_A_totwC3zQ5_0),.din(w_dff_A_P07lZhrt0_0),.clk(gclk));
	jdff dff_A_totwC3zQ5_0(.dout(w_dff_A_cMqDTa7Z0_0),.din(w_dff_A_totwC3zQ5_0),.clk(gclk));
	jdff dff_A_cMqDTa7Z0_0(.dout(w_dff_A_iBdouH5S5_0),.din(w_dff_A_cMqDTa7Z0_0),.clk(gclk));
	jdff dff_A_iBdouH5S5_0(.dout(w_dff_A_3VKFQcpz6_0),.din(w_dff_A_iBdouH5S5_0),.clk(gclk));
	jdff dff_A_3VKFQcpz6_0(.dout(w_dff_A_T9P5G9uA4_0),.din(w_dff_A_3VKFQcpz6_0),.clk(gclk));
	jdff dff_A_T9P5G9uA4_0(.dout(w_dff_A_5rr3c4HZ8_0),.din(w_dff_A_T9P5G9uA4_0),.clk(gclk));
	jdff dff_A_5rr3c4HZ8_0(.dout(w_dff_A_d8ncZiCq3_0),.din(w_dff_A_5rr3c4HZ8_0),.clk(gclk));
	jdff dff_A_d8ncZiCq3_0(.dout(w_dff_A_KYIgKngs5_0),.din(w_dff_A_d8ncZiCq3_0),.clk(gclk));
	jdff dff_A_KYIgKngs5_0(.dout(w_dff_A_qTx1po8g7_0),.din(w_dff_A_KYIgKngs5_0),.clk(gclk));
	jdff dff_A_qTx1po8g7_0(.dout(w_dff_A_0tW622NM2_0),.din(w_dff_A_qTx1po8g7_0),.clk(gclk));
	jdff dff_A_0tW622NM2_0(.dout(w_dff_A_sdiKqK4P3_0),.din(w_dff_A_0tW622NM2_0),.clk(gclk));
	jdff dff_A_sdiKqK4P3_0(.dout(w_dff_A_gzziJXjC0_0),.din(w_dff_A_sdiKqK4P3_0),.clk(gclk));
	jdff dff_A_gzziJXjC0_0(.dout(w_dff_A_USJhQbOg3_0),.din(w_dff_A_gzziJXjC0_0),.clk(gclk));
	jdff dff_A_USJhQbOg3_0(.dout(w_dff_A_LBF6doIT2_0),.din(w_dff_A_USJhQbOg3_0),.clk(gclk));
	jdff dff_A_LBF6doIT2_0(.dout(w_dff_A_fBpDS66K8_0),.din(w_dff_A_LBF6doIT2_0),.clk(gclk));
	jdff dff_A_fBpDS66K8_0(.dout(w_dff_A_icL07ajY8_0),.din(w_dff_A_fBpDS66K8_0),.clk(gclk));
	jdff dff_A_icL07ajY8_0(.dout(w_dff_A_SS5zIw232_0),.din(w_dff_A_icL07ajY8_0),.clk(gclk));
	jdff dff_A_SS5zIw232_0(.dout(w_dff_A_qCEiOyxe6_0),.din(w_dff_A_SS5zIw232_0),.clk(gclk));
	jdff dff_A_qCEiOyxe6_0(.dout(w_dff_A_S4fqUD1W6_0),.din(w_dff_A_qCEiOyxe6_0),.clk(gclk));
	jdff dff_A_S4fqUD1W6_0(.dout(w_dff_A_VMd4BWbO7_0),.din(w_dff_A_S4fqUD1W6_0),.clk(gclk));
	jdff dff_A_VMd4BWbO7_0(.dout(w_dff_A_72TtIEga5_0),.din(w_dff_A_VMd4BWbO7_0),.clk(gclk));
	jdff dff_A_72TtIEga5_0(.dout(w_dff_A_GRCmtOQz2_0),.din(w_dff_A_72TtIEga5_0),.clk(gclk));
	jdff dff_A_GRCmtOQz2_0(.dout(w_dff_A_bM2a9uym8_0),.din(w_dff_A_GRCmtOQz2_0),.clk(gclk));
	jdff dff_A_bM2a9uym8_0(.dout(G284),.din(w_dff_A_bM2a9uym8_0),.clk(gclk));
	jdff dff_A_2CM4RefF3_1(.dout(w_dff_A_n5yoZDCf8_0),.din(w_dff_A_2CM4RefF3_1),.clk(gclk));
	jdff dff_A_n5yoZDCf8_0(.dout(w_dff_A_bKF5IE3v5_0),.din(w_dff_A_n5yoZDCf8_0),.clk(gclk));
	jdff dff_A_bKF5IE3v5_0(.dout(w_dff_A_4zRKyYlP0_0),.din(w_dff_A_bKF5IE3v5_0),.clk(gclk));
	jdff dff_A_4zRKyYlP0_0(.dout(w_dff_A_VWD6FnwO0_0),.din(w_dff_A_4zRKyYlP0_0),.clk(gclk));
	jdff dff_A_VWD6FnwO0_0(.dout(w_dff_A_c7AkPyDO7_0),.din(w_dff_A_VWD6FnwO0_0),.clk(gclk));
	jdff dff_A_c7AkPyDO7_0(.dout(w_dff_A_NU8Yegop7_0),.din(w_dff_A_c7AkPyDO7_0),.clk(gclk));
	jdff dff_A_NU8Yegop7_0(.dout(w_dff_A_FjyWPSxX2_0),.din(w_dff_A_NU8Yegop7_0),.clk(gclk));
	jdff dff_A_FjyWPSxX2_0(.dout(w_dff_A_qX7D6fDA9_0),.din(w_dff_A_FjyWPSxX2_0),.clk(gclk));
	jdff dff_A_qX7D6fDA9_0(.dout(w_dff_A_jiIR7V6H0_0),.din(w_dff_A_qX7D6fDA9_0),.clk(gclk));
	jdff dff_A_jiIR7V6H0_0(.dout(w_dff_A_u69AqvrK0_0),.din(w_dff_A_jiIR7V6H0_0),.clk(gclk));
	jdff dff_A_u69AqvrK0_0(.dout(w_dff_A_TSC8EBos4_0),.din(w_dff_A_u69AqvrK0_0),.clk(gclk));
	jdff dff_A_TSC8EBos4_0(.dout(w_dff_A_TMTyYm9x4_0),.din(w_dff_A_TSC8EBos4_0),.clk(gclk));
	jdff dff_A_TMTyYm9x4_0(.dout(w_dff_A_iVmQubmu0_0),.din(w_dff_A_TMTyYm9x4_0),.clk(gclk));
	jdff dff_A_iVmQubmu0_0(.dout(w_dff_A_4kYU3pSG2_0),.din(w_dff_A_iVmQubmu0_0),.clk(gclk));
	jdff dff_A_4kYU3pSG2_0(.dout(w_dff_A_TOO6hyuv1_0),.din(w_dff_A_4kYU3pSG2_0),.clk(gclk));
	jdff dff_A_TOO6hyuv1_0(.dout(w_dff_A_pqZdBcaF9_0),.din(w_dff_A_TOO6hyuv1_0),.clk(gclk));
	jdff dff_A_pqZdBcaF9_0(.dout(w_dff_A_Fbjf0KqF1_0),.din(w_dff_A_pqZdBcaF9_0),.clk(gclk));
	jdff dff_A_Fbjf0KqF1_0(.dout(w_dff_A_dB48OhgZ7_0),.din(w_dff_A_Fbjf0KqF1_0),.clk(gclk));
	jdff dff_A_dB48OhgZ7_0(.dout(w_dff_A_zCkggYEu9_0),.din(w_dff_A_dB48OhgZ7_0),.clk(gclk));
	jdff dff_A_zCkggYEu9_0(.dout(w_dff_A_XrWLbXV64_0),.din(w_dff_A_zCkggYEu9_0),.clk(gclk));
	jdff dff_A_XrWLbXV64_0(.dout(w_dff_A_nDeGW0gs1_0),.din(w_dff_A_XrWLbXV64_0),.clk(gclk));
	jdff dff_A_nDeGW0gs1_0(.dout(w_dff_A_AWxxHpcb5_0),.din(w_dff_A_nDeGW0gs1_0),.clk(gclk));
	jdff dff_A_AWxxHpcb5_0(.dout(w_dff_A_KMlUbPeh0_0),.din(w_dff_A_AWxxHpcb5_0),.clk(gclk));
	jdff dff_A_KMlUbPeh0_0(.dout(w_dff_A_uLqjC8R84_0),.din(w_dff_A_KMlUbPeh0_0),.clk(gclk));
	jdff dff_A_uLqjC8R84_0(.dout(w_dff_A_Wiwszthh8_0),.din(w_dff_A_uLqjC8R84_0),.clk(gclk));
	jdff dff_A_Wiwszthh8_0(.dout(w_dff_A_GQtNPTjH2_0),.din(w_dff_A_Wiwszthh8_0),.clk(gclk));
	jdff dff_A_GQtNPTjH2_0(.dout(w_dff_A_ul6SvONu8_0),.din(w_dff_A_GQtNPTjH2_0),.clk(gclk));
	jdff dff_A_ul6SvONu8_0(.dout(w_dff_A_3C3pdOhQ0_0),.din(w_dff_A_ul6SvONu8_0),.clk(gclk));
	jdff dff_A_3C3pdOhQ0_0(.dout(w_dff_A_gwXh8D4n5_0),.din(w_dff_A_3C3pdOhQ0_0),.clk(gclk));
	jdff dff_A_gwXh8D4n5_0(.dout(w_dff_A_CwSzkxRm1_0),.din(w_dff_A_gwXh8D4n5_0),.clk(gclk));
	jdff dff_A_CwSzkxRm1_0(.dout(w_dff_A_N1pluRYG2_0),.din(w_dff_A_CwSzkxRm1_0),.clk(gclk));
	jdff dff_A_N1pluRYG2_0(.dout(w_dff_A_Xa6DPwYr3_0),.din(w_dff_A_N1pluRYG2_0),.clk(gclk));
	jdff dff_A_Xa6DPwYr3_0(.dout(w_dff_A_GU7r6nvd5_0),.din(w_dff_A_Xa6DPwYr3_0),.clk(gclk));
	jdff dff_A_GU7r6nvd5_0(.dout(w_dff_A_mrVNT3gD6_0),.din(w_dff_A_GU7r6nvd5_0),.clk(gclk));
	jdff dff_A_mrVNT3gD6_0(.dout(w_dff_A_coFlINwc6_0),.din(w_dff_A_mrVNT3gD6_0),.clk(gclk));
	jdff dff_A_coFlINwc6_0(.dout(w_dff_A_2i4GnoHT7_0),.din(w_dff_A_coFlINwc6_0),.clk(gclk));
	jdff dff_A_2i4GnoHT7_0(.dout(w_dff_A_GEUJn6gc6_0),.din(w_dff_A_2i4GnoHT7_0),.clk(gclk));
	jdff dff_A_GEUJn6gc6_0(.dout(G286),.din(w_dff_A_GEUJn6gc6_0),.clk(gclk));
	jdff dff_A_ZwTqURVo7_2(.dout(w_dff_A_plbNHkHT8_0),.din(w_dff_A_ZwTqURVo7_2),.clk(gclk));
	jdff dff_A_plbNHkHT8_0(.dout(w_dff_A_62v67yL61_0),.din(w_dff_A_plbNHkHT8_0),.clk(gclk));
	jdff dff_A_62v67yL61_0(.dout(w_dff_A_lzLj9gwB7_0),.din(w_dff_A_62v67yL61_0),.clk(gclk));
	jdff dff_A_lzLj9gwB7_0(.dout(w_dff_A_AMqU5Q7T1_0),.din(w_dff_A_lzLj9gwB7_0),.clk(gclk));
	jdff dff_A_AMqU5Q7T1_0(.dout(w_dff_A_rKxjZvUk8_0),.din(w_dff_A_AMqU5Q7T1_0),.clk(gclk));
	jdff dff_A_rKxjZvUk8_0(.dout(w_dff_A_IokWATAQ4_0),.din(w_dff_A_rKxjZvUk8_0),.clk(gclk));
	jdff dff_A_IokWATAQ4_0(.dout(w_dff_A_BgZ99lLa4_0),.din(w_dff_A_IokWATAQ4_0),.clk(gclk));
	jdff dff_A_BgZ99lLa4_0(.dout(w_dff_A_pJnvJxP37_0),.din(w_dff_A_BgZ99lLa4_0),.clk(gclk));
	jdff dff_A_pJnvJxP37_0(.dout(w_dff_A_yxQp2DIN4_0),.din(w_dff_A_pJnvJxP37_0),.clk(gclk));
	jdff dff_A_yxQp2DIN4_0(.dout(w_dff_A_ocwSjP7n9_0),.din(w_dff_A_yxQp2DIN4_0),.clk(gclk));
	jdff dff_A_ocwSjP7n9_0(.dout(w_dff_A_tgOR6fJn0_0),.din(w_dff_A_ocwSjP7n9_0),.clk(gclk));
	jdff dff_A_tgOR6fJn0_0(.dout(w_dff_A_h4ApIzZf9_0),.din(w_dff_A_tgOR6fJn0_0),.clk(gclk));
	jdff dff_A_h4ApIzZf9_0(.dout(w_dff_A_EKQhDHtQ6_0),.din(w_dff_A_h4ApIzZf9_0),.clk(gclk));
	jdff dff_A_EKQhDHtQ6_0(.dout(w_dff_A_rTmEYGpL2_0),.din(w_dff_A_EKQhDHtQ6_0),.clk(gclk));
	jdff dff_A_rTmEYGpL2_0(.dout(w_dff_A_Oh1EcsKi0_0),.din(w_dff_A_rTmEYGpL2_0),.clk(gclk));
	jdff dff_A_Oh1EcsKi0_0(.dout(w_dff_A_QbVMJAyt6_0),.din(w_dff_A_Oh1EcsKi0_0),.clk(gclk));
	jdff dff_A_QbVMJAyt6_0(.dout(w_dff_A_x38VK13U7_0),.din(w_dff_A_QbVMJAyt6_0),.clk(gclk));
	jdff dff_A_x38VK13U7_0(.dout(w_dff_A_Lf3y1ZlA5_0),.din(w_dff_A_x38VK13U7_0),.clk(gclk));
	jdff dff_A_Lf3y1ZlA5_0(.dout(w_dff_A_pkU8CXXw0_0),.din(w_dff_A_Lf3y1ZlA5_0),.clk(gclk));
	jdff dff_A_pkU8CXXw0_0(.dout(w_dff_A_yUQyUETs8_0),.din(w_dff_A_pkU8CXXw0_0),.clk(gclk));
	jdff dff_A_yUQyUETs8_0(.dout(w_dff_A_kq3u3yqe7_0),.din(w_dff_A_yUQyUETs8_0),.clk(gclk));
	jdff dff_A_kq3u3yqe7_0(.dout(w_dff_A_v9ZiQGw37_0),.din(w_dff_A_kq3u3yqe7_0),.clk(gclk));
	jdff dff_A_v9ZiQGw37_0(.dout(w_dff_A_4ryWWJ1Q2_0),.din(w_dff_A_v9ZiQGw37_0),.clk(gclk));
	jdff dff_A_4ryWWJ1Q2_0(.dout(w_dff_A_wzbqZFOy7_0),.din(w_dff_A_4ryWWJ1Q2_0),.clk(gclk));
	jdff dff_A_wzbqZFOy7_0(.dout(w_dff_A_j1ezqyNl7_0),.din(w_dff_A_wzbqZFOy7_0),.clk(gclk));
	jdff dff_A_j1ezqyNl7_0(.dout(w_dff_A_blHQsdka1_0),.din(w_dff_A_j1ezqyNl7_0),.clk(gclk));
	jdff dff_A_blHQsdka1_0(.dout(w_dff_A_5eU4ibM80_0),.din(w_dff_A_blHQsdka1_0),.clk(gclk));
	jdff dff_A_5eU4ibM80_0(.dout(w_dff_A_AHgRfG8G2_0),.din(w_dff_A_5eU4ibM80_0),.clk(gclk));
	jdff dff_A_AHgRfG8G2_0(.dout(w_dff_A_frXSsZH08_0),.din(w_dff_A_AHgRfG8G2_0),.clk(gclk));
	jdff dff_A_frXSsZH08_0(.dout(w_dff_A_0vJJS7Pc9_0),.din(w_dff_A_frXSsZH08_0),.clk(gclk));
	jdff dff_A_0vJJS7Pc9_0(.dout(w_dff_A_EqH1qAAp1_0),.din(w_dff_A_0vJJS7Pc9_0),.clk(gclk));
	jdff dff_A_EqH1qAAp1_0(.dout(w_dff_A_uUWmgIk26_0),.din(w_dff_A_EqH1qAAp1_0),.clk(gclk));
	jdff dff_A_uUWmgIk26_0(.dout(w_dff_A_Xwr63UvT2_0),.din(w_dff_A_uUWmgIk26_0),.clk(gclk));
	jdff dff_A_Xwr63UvT2_0(.dout(w_dff_A_aNtfbfzQ8_0),.din(w_dff_A_Xwr63UvT2_0),.clk(gclk));
	jdff dff_A_aNtfbfzQ8_0(.dout(w_dff_A_n5p0vNWm1_0),.din(w_dff_A_aNtfbfzQ8_0),.clk(gclk));
	jdff dff_A_n5p0vNWm1_0(.dout(w_dff_A_16veWjrJ2_0),.din(w_dff_A_n5p0vNWm1_0),.clk(gclk));
	jdff dff_A_16veWjrJ2_0(.dout(G289),.din(w_dff_A_16veWjrJ2_0),.clk(gclk));
	jdff dff_A_x6bwFvue0_2(.dout(w_dff_A_vJTDuolT8_0),.din(w_dff_A_x6bwFvue0_2),.clk(gclk));
	jdff dff_A_vJTDuolT8_0(.dout(w_dff_A_mVRE5PBb3_0),.din(w_dff_A_vJTDuolT8_0),.clk(gclk));
	jdff dff_A_mVRE5PBb3_0(.dout(w_dff_A_j4HHhwUy1_0),.din(w_dff_A_mVRE5PBb3_0),.clk(gclk));
	jdff dff_A_j4HHhwUy1_0(.dout(w_dff_A_8ymnaPga4_0),.din(w_dff_A_j4HHhwUy1_0),.clk(gclk));
	jdff dff_A_8ymnaPga4_0(.dout(w_dff_A_gMawEEuw6_0),.din(w_dff_A_8ymnaPga4_0),.clk(gclk));
	jdff dff_A_gMawEEuw6_0(.dout(w_dff_A_kkOSS41X7_0),.din(w_dff_A_gMawEEuw6_0),.clk(gclk));
	jdff dff_A_kkOSS41X7_0(.dout(w_dff_A_FokBI5dd4_0),.din(w_dff_A_kkOSS41X7_0),.clk(gclk));
	jdff dff_A_FokBI5dd4_0(.dout(w_dff_A_eKfA5OVK9_0),.din(w_dff_A_FokBI5dd4_0),.clk(gclk));
	jdff dff_A_eKfA5OVK9_0(.dout(w_dff_A_oLhL8F5V8_0),.din(w_dff_A_eKfA5OVK9_0),.clk(gclk));
	jdff dff_A_oLhL8F5V8_0(.dout(w_dff_A_xm5UzF4w4_0),.din(w_dff_A_oLhL8F5V8_0),.clk(gclk));
	jdff dff_A_xm5UzF4w4_0(.dout(w_dff_A_xirkfDEl9_0),.din(w_dff_A_xm5UzF4w4_0),.clk(gclk));
	jdff dff_A_xirkfDEl9_0(.dout(w_dff_A_VSyMBy6L9_0),.din(w_dff_A_xirkfDEl9_0),.clk(gclk));
	jdff dff_A_VSyMBy6L9_0(.dout(w_dff_A_hwPy5vzu4_0),.din(w_dff_A_VSyMBy6L9_0),.clk(gclk));
	jdff dff_A_hwPy5vzu4_0(.dout(w_dff_A_bVZYnrVS2_0),.din(w_dff_A_hwPy5vzu4_0),.clk(gclk));
	jdff dff_A_bVZYnrVS2_0(.dout(w_dff_A_qKLwvFUP1_0),.din(w_dff_A_bVZYnrVS2_0),.clk(gclk));
	jdff dff_A_qKLwvFUP1_0(.dout(w_dff_A_PWdW3zAt4_0),.din(w_dff_A_qKLwvFUP1_0),.clk(gclk));
	jdff dff_A_PWdW3zAt4_0(.dout(w_dff_A_xPZrV0SC3_0),.din(w_dff_A_PWdW3zAt4_0),.clk(gclk));
	jdff dff_A_xPZrV0SC3_0(.dout(w_dff_A_fJaFXqRS8_0),.din(w_dff_A_xPZrV0SC3_0),.clk(gclk));
	jdff dff_A_fJaFXqRS8_0(.dout(w_dff_A_TPgnHYr46_0),.din(w_dff_A_fJaFXqRS8_0),.clk(gclk));
	jdff dff_A_TPgnHYr46_0(.dout(w_dff_A_xAKLmj6O5_0),.din(w_dff_A_TPgnHYr46_0),.clk(gclk));
	jdff dff_A_xAKLmj6O5_0(.dout(w_dff_A_QWWWZ0AH4_0),.din(w_dff_A_xAKLmj6O5_0),.clk(gclk));
	jdff dff_A_QWWWZ0AH4_0(.dout(w_dff_A_s6o5VFmK0_0),.din(w_dff_A_QWWWZ0AH4_0),.clk(gclk));
	jdff dff_A_s6o5VFmK0_0(.dout(w_dff_A_gXKFYeAi4_0),.din(w_dff_A_s6o5VFmK0_0),.clk(gclk));
	jdff dff_A_gXKFYeAi4_0(.dout(w_dff_A_KfUohfH77_0),.din(w_dff_A_gXKFYeAi4_0),.clk(gclk));
	jdff dff_A_KfUohfH77_0(.dout(w_dff_A_IxFXTg752_0),.din(w_dff_A_KfUohfH77_0),.clk(gclk));
	jdff dff_A_IxFXTg752_0(.dout(w_dff_A_fjgkxzkq0_0),.din(w_dff_A_IxFXTg752_0),.clk(gclk));
	jdff dff_A_fjgkxzkq0_0(.dout(w_dff_A_cR61TyC04_0),.din(w_dff_A_fjgkxzkq0_0),.clk(gclk));
	jdff dff_A_cR61TyC04_0(.dout(w_dff_A_lJS3UL8m0_0),.din(w_dff_A_cR61TyC04_0),.clk(gclk));
	jdff dff_A_lJS3UL8m0_0(.dout(w_dff_A_jzmgkfkQ5_0),.din(w_dff_A_lJS3UL8m0_0),.clk(gclk));
	jdff dff_A_jzmgkfkQ5_0(.dout(w_dff_A_T7UAfG1r1_0),.din(w_dff_A_jzmgkfkQ5_0),.clk(gclk));
	jdff dff_A_T7UAfG1r1_0(.dout(w_dff_A_PVcoIPhT0_0),.din(w_dff_A_T7UAfG1r1_0),.clk(gclk));
	jdff dff_A_PVcoIPhT0_0(.dout(w_dff_A_of390Vzo3_0),.din(w_dff_A_PVcoIPhT0_0),.clk(gclk));
	jdff dff_A_of390Vzo3_0(.dout(w_dff_A_GDUSIUm76_0),.din(w_dff_A_of390Vzo3_0),.clk(gclk));
	jdff dff_A_GDUSIUm76_0(.dout(w_dff_A_hYnJaZzd3_0),.din(w_dff_A_GDUSIUm76_0),.clk(gclk));
	jdff dff_A_hYnJaZzd3_0(.dout(w_dff_A_3SV0BPMb8_0),.din(w_dff_A_hYnJaZzd3_0),.clk(gclk));
	jdff dff_A_3SV0BPMb8_0(.dout(G292),.din(w_dff_A_3SV0BPMb8_0),.clk(gclk));
	jdff dff_A_0w6Csyvn8_1(.dout(w_dff_A_aJRzz02e8_0),.din(w_dff_A_0w6Csyvn8_1),.clk(gclk));
	jdff dff_A_aJRzz02e8_0(.dout(w_dff_A_ySSvZSMX1_0),.din(w_dff_A_aJRzz02e8_0),.clk(gclk));
	jdff dff_A_ySSvZSMX1_0(.dout(w_dff_A_817qS1Yx7_0),.din(w_dff_A_ySSvZSMX1_0),.clk(gclk));
	jdff dff_A_817qS1Yx7_0(.dout(w_dff_A_vwTRdGvn7_0),.din(w_dff_A_817qS1Yx7_0),.clk(gclk));
	jdff dff_A_vwTRdGvn7_0(.dout(w_dff_A_NmgrfalF8_0),.din(w_dff_A_vwTRdGvn7_0),.clk(gclk));
	jdff dff_A_NmgrfalF8_0(.dout(w_dff_A_DMZsHzAL7_0),.din(w_dff_A_NmgrfalF8_0),.clk(gclk));
	jdff dff_A_DMZsHzAL7_0(.dout(w_dff_A_wcMw7NWP6_0),.din(w_dff_A_DMZsHzAL7_0),.clk(gclk));
	jdff dff_A_wcMw7NWP6_0(.dout(w_dff_A_3gaDqzmV2_0),.din(w_dff_A_wcMw7NWP6_0),.clk(gclk));
	jdff dff_A_3gaDqzmV2_0(.dout(w_dff_A_WOxNUutk7_0),.din(w_dff_A_3gaDqzmV2_0),.clk(gclk));
	jdff dff_A_WOxNUutk7_0(.dout(w_dff_A_Tpyuw7Lb4_0),.din(w_dff_A_WOxNUutk7_0),.clk(gclk));
	jdff dff_A_Tpyuw7Lb4_0(.dout(w_dff_A_vGyNWZlW9_0),.din(w_dff_A_Tpyuw7Lb4_0),.clk(gclk));
	jdff dff_A_vGyNWZlW9_0(.dout(w_dff_A_vY89ozsT9_0),.din(w_dff_A_vGyNWZlW9_0),.clk(gclk));
	jdff dff_A_vY89ozsT9_0(.dout(w_dff_A_W92VnVZr5_0),.din(w_dff_A_vY89ozsT9_0),.clk(gclk));
	jdff dff_A_W92VnVZr5_0(.dout(w_dff_A_1S4h1ec35_0),.din(w_dff_A_W92VnVZr5_0),.clk(gclk));
	jdff dff_A_1S4h1ec35_0(.dout(w_dff_A_nQYf6h6r3_0),.din(w_dff_A_1S4h1ec35_0),.clk(gclk));
	jdff dff_A_nQYf6h6r3_0(.dout(w_dff_A_XFgQYpmq3_0),.din(w_dff_A_nQYf6h6r3_0),.clk(gclk));
	jdff dff_A_XFgQYpmq3_0(.dout(w_dff_A_dTAP4cXN1_0),.din(w_dff_A_XFgQYpmq3_0),.clk(gclk));
	jdff dff_A_dTAP4cXN1_0(.dout(w_dff_A_vCjQO0hF3_0),.din(w_dff_A_dTAP4cXN1_0),.clk(gclk));
	jdff dff_A_vCjQO0hF3_0(.dout(w_dff_A_32bftMGQ8_0),.din(w_dff_A_vCjQO0hF3_0),.clk(gclk));
	jdff dff_A_32bftMGQ8_0(.dout(w_dff_A_T4hKSIS77_0),.din(w_dff_A_32bftMGQ8_0),.clk(gclk));
	jdff dff_A_T4hKSIS77_0(.dout(w_dff_A_REX2j62H4_0),.din(w_dff_A_T4hKSIS77_0),.clk(gclk));
	jdff dff_A_REX2j62H4_0(.dout(w_dff_A_Gq3lznHz2_0),.din(w_dff_A_REX2j62H4_0),.clk(gclk));
	jdff dff_A_Gq3lznHz2_0(.dout(w_dff_A_QhEIEVDd9_0),.din(w_dff_A_Gq3lznHz2_0),.clk(gclk));
	jdff dff_A_QhEIEVDd9_0(.dout(w_dff_A_bHzDProK3_0),.din(w_dff_A_QhEIEVDd9_0),.clk(gclk));
	jdff dff_A_bHzDProK3_0(.dout(w_dff_A_ykyFEO5f6_0),.din(w_dff_A_bHzDProK3_0),.clk(gclk));
	jdff dff_A_ykyFEO5f6_0(.dout(w_dff_A_lNTfgc6s7_0),.din(w_dff_A_ykyFEO5f6_0),.clk(gclk));
	jdff dff_A_lNTfgc6s7_0(.dout(w_dff_A_oOdCMo2h3_0),.din(w_dff_A_lNTfgc6s7_0),.clk(gclk));
	jdff dff_A_oOdCMo2h3_0(.dout(w_dff_A_ZESI0Ss79_0),.din(w_dff_A_oOdCMo2h3_0),.clk(gclk));
	jdff dff_A_ZESI0Ss79_0(.dout(w_dff_A_EWfjLcQY6_0),.din(w_dff_A_ZESI0Ss79_0),.clk(gclk));
	jdff dff_A_EWfjLcQY6_0(.dout(w_dff_A_qmZVpdSi9_0),.din(w_dff_A_EWfjLcQY6_0),.clk(gclk));
	jdff dff_A_qmZVpdSi9_0(.dout(w_dff_A_2vQLWaaH3_0),.din(w_dff_A_qmZVpdSi9_0),.clk(gclk));
	jdff dff_A_2vQLWaaH3_0(.dout(w_dff_A_03PM1Ut50_0),.din(w_dff_A_2vQLWaaH3_0),.clk(gclk));
	jdff dff_A_03PM1Ut50_0(.dout(w_dff_A_UhMHdjPL6_0),.din(w_dff_A_03PM1Ut50_0),.clk(gclk));
	jdff dff_A_UhMHdjPL6_0(.dout(w_dff_A_uz1hkg592_0),.din(w_dff_A_UhMHdjPL6_0),.clk(gclk));
	jdff dff_A_uz1hkg592_0(.dout(w_dff_A_cCEHWIOR6_0),.din(w_dff_A_uz1hkg592_0),.clk(gclk));
	jdff dff_A_cCEHWIOR6_0(.dout(w_dff_A_9Pj9fEaC9_0),.din(w_dff_A_cCEHWIOR6_0),.clk(gclk));
	jdff dff_A_9Pj9fEaC9_0(.dout(w_dff_A_vT7Mf1cx5_0),.din(w_dff_A_9Pj9fEaC9_0),.clk(gclk));
	jdff dff_A_vT7Mf1cx5_0(.dout(G341),.din(w_dff_A_vT7Mf1cx5_0),.clk(gclk));
	jdff dff_A_UKxWtnJd8_2(.dout(w_dff_A_RuP9411f3_0),.din(w_dff_A_UKxWtnJd8_2),.clk(gclk));
	jdff dff_A_RuP9411f3_0(.dout(w_dff_A_ALhJE6hN7_0),.din(w_dff_A_RuP9411f3_0),.clk(gclk));
	jdff dff_A_ALhJE6hN7_0(.dout(w_dff_A_GbNS7SoF3_0),.din(w_dff_A_ALhJE6hN7_0),.clk(gclk));
	jdff dff_A_GbNS7SoF3_0(.dout(w_dff_A_cn5ShnvJ9_0),.din(w_dff_A_GbNS7SoF3_0),.clk(gclk));
	jdff dff_A_cn5ShnvJ9_0(.dout(w_dff_A_qwTw1RaX2_0),.din(w_dff_A_cn5ShnvJ9_0),.clk(gclk));
	jdff dff_A_qwTw1RaX2_0(.dout(w_dff_A_PNs8KCUb1_0),.din(w_dff_A_qwTw1RaX2_0),.clk(gclk));
	jdff dff_A_PNs8KCUb1_0(.dout(w_dff_A_93QzkCA82_0),.din(w_dff_A_PNs8KCUb1_0),.clk(gclk));
	jdff dff_A_93QzkCA82_0(.dout(w_dff_A_xglkL6wa8_0),.din(w_dff_A_93QzkCA82_0),.clk(gclk));
	jdff dff_A_xglkL6wa8_0(.dout(w_dff_A_LXbpOo1Z0_0),.din(w_dff_A_xglkL6wa8_0),.clk(gclk));
	jdff dff_A_LXbpOo1Z0_0(.dout(w_dff_A_Xvh2uMQd3_0),.din(w_dff_A_LXbpOo1Z0_0),.clk(gclk));
	jdff dff_A_Xvh2uMQd3_0(.dout(w_dff_A_LRBna6GA3_0),.din(w_dff_A_Xvh2uMQd3_0),.clk(gclk));
	jdff dff_A_LRBna6GA3_0(.dout(w_dff_A_AESoj9m69_0),.din(w_dff_A_LRBna6GA3_0),.clk(gclk));
	jdff dff_A_AESoj9m69_0(.dout(w_dff_A_SXECSwnZ7_0),.din(w_dff_A_AESoj9m69_0),.clk(gclk));
	jdff dff_A_SXECSwnZ7_0(.dout(w_dff_A_DKCrPw4f9_0),.din(w_dff_A_SXECSwnZ7_0),.clk(gclk));
	jdff dff_A_DKCrPw4f9_0(.dout(w_dff_A_eXmqM5jx6_0),.din(w_dff_A_DKCrPw4f9_0),.clk(gclk));
	jdff dff_A_eXmqM5jx6_0(.dout(w_dff_A_w4oSo3Yn8_0),.din(w_dff_A_eXmqM5jx6_0),.clk(gclk));
	jdff dff_A_w4oSo3Yn8_0(.dout(w_dff_A_91V8v4Y38_0),.din(w_dff_A_w4oSo3Yn8_0),.clk(gclk));
	jdff dff_A_91V8v4Y38_0(.dout(w_dff_A_nULIvwbz1_0),.din(w_dff_A_91V8v4Y38_0),.clk(gclk));
	jdff dff_A_nULIvwbz1_0(.dout(w_dff_A_2c8d4vxf3_0),.din(w_dff_A_nULIvwbz1_0),.clk(gclk));
	jdff dff_A_2c8d4vxf3_0(.dout(w_dff_A_rND2kL1W5_0),.din(w_dff_A_2c8d4vxf3_0),.clk(gclk));
	jdff dff_A_rND2kL1W5_0(.dout(w_dff_A_vZpAs4mw8_0),.din(w_dff_A_rND2kL1W5_0),.clk(gclk));
	jdff dff_A_vZpAs4mw8_0(.dout(w_dff_A_BZ0hxsoU0_0),.din(w_dff_A_vZpAs4mw8_0),.clk(gclk));
	jdff dff_A_BZ0hxsoU0_0(.dout(w_dff_A_BDOGNpk46_0),.din(w_dff_A_BZ0hxsoU0_0),.clk(gclk));
	jdff dff_A_BDOGNpk46_0(.dout(w_dff_A_TZznJtTl5_0),.din(w_dff_A_BDOGNpk46_0),.clk(gclk));
	jdff dff_A_TZznJtTl5_0(.dout(w_dff_A_ZYFuPgoN6_0),.din(w_dff_A_TZznJtTl5_0),.clk(gclk));
	jdff dff_A_ZYFuPgoN6_0(.dout(w_dff_A_c1vNB3sB2_0),.din(w_dff_A_ZYFuPgoN6_0),.clk(gclk));
	jdff dff_A_c1vNB3sB2_0(.dout(w_dff_A_tmxk6DYN5_0),.din(w_dff_A_c1vNB3sB2_0),.clk(gclk));
	jdff dff_A_tmxk6DYN5_0(.dout(w_dff_A_Flz6wzH57_0),.din(w_dff_A_tmxk6DYN5_0),.clk(gclk));
	jdff dff_A_Flz6wzH57_0(.dout(w_dff_A_WzZOrcEQ3_0),.din(w_dff_A_Flz6wzH57_0),.clk(gclk));
	jdff dff_A_WzZOrcEQ3_0(.dout(w_dff_A_Pd7S7EJy4_0),.din(w_dff_A_WzZOrcEQ3_0),.clk(gclk));
	jdff dff_A_Pd7S7EJy4_0(.dout(w_dff_A_fVJNAEaJ9_0),.din(w_dff_A_Pd7S7EJy4_0),.clk(gclk));
	jdff dff_A_fVJNAEaJ9_0(.dout(w_dff_A_j7TRNiBv1_0),.din(w_dff_A_fVJNAEaJ9_0),.clk(gclk));
	jdff dff_A_j7TRNiBv1_0(.dout(w_dff_A_jWybCdhP2_0),.din(w_dff_A_j7TRNiBv1_0),.clk(gclk));
	jdff dff_A_jWybCdhP2_0(.dout(w_dff_A_RWyN0RFi0_0),.din(w_dff_A_jWybCdhP2_0),.clk(gclk));
	jdff dff_A_RWyN0RFi0_0(.dout(w_dff_A_jQgGwhbs3_0),.din(w_dff_A_RWyN0RFi0_0),.clk(gclk));
	jdff dff_A_jQgGwhbs3_0(.dout(G281),.din(w_dff_A_jQgGwhbs3_0),.clk(gclk));
	jdff dff_A_M0HT7wKV8_1(.dout(w_dff_A_XEH1iaR35_0),.din(w_dff_A_M0HT7wKV8_1),.clk(gclk));
	jdff dff_A_XEH1iaR35_0(.dout(w_dff_A_CqiTVAVZ2_0),.din(w_dff_A_XEH1iaR35_0),.clk(gclk));
	jdff dff_A_CqiTVAVZ2_0(.dout(w_dff_A_bsfuE8Sl1_0),.din(w_dff_A_CqiTVAVZ2_0),.clk(gclk));
	jdff dff_A_bsfuE8Sl1_0(.dout(w_dff_A_zWxyzn3l5_0),.din(w_dff_A_bsfuE8Sl1_0),.clk(gclk));
	jdff dff_A_zWxyzn3l5_0(.dout(w_dff_A_WzuUtemE3_0),.din(w_dff_A_zWxyzn3l5_0),.clk(gclk));
	jdff dff_A_WzuUtemE3_0(.dout(w_dff_A_paBSIU5t2_0),.din(w_dff_A_WzuUtemE3_0),.clk(gclk));
	jdff dff_A_paBSIU5t2_0(.dout(w_dff_A_nu7sBOC97_0),.din(w_dff_A_paBSIU5t2_0),.clk(gclk));
	jdff dff_A_nu7sBOC97_0(.dout(w_dff_A_HzvtWlB31_0),.din(w_dff_A_nu7sBOC97_0),.clk(gclk));
	jdff dff_A_HzvtWlB31_0(.dout(w_dff_A_kuGB9u1T4_0),.din(w_dff_A_HzvtWlB31_0),.clk(gclk));
	jdff dff_A_kuGB9u1T4_0(.dout(w_dff_A_q0C6jZsZ7_0),.din(w_dff_A_kuGB9u1T4_0),.clk(gclk));
	jdff dff_A_q0C6jZsZ7_0(.dout(w_dff_A_ATNOlEmw6_0),.din(w_dff_A_q0C6jZsZ7_0),.clk(gclk));
	jdff dff_A_ATNOlEmw6_0(.dout(w_dff_A_l78yR6Lg3_0),.din(w_dff_A_ATNOlEmw6_0),.clk(gclk));
	jdff dff_A_l78yR6Lg3_0(.dout(w_dff_A_WeboNXlf9_0),.din(w_dff_A_l78yR6Lg3_0),.clk(gclk));
	jdff dff_A_WeboNXlf9_0(.dout(w_dff_A_6Xgt1Nuk4_0),.din(w_dff_A_WeboNXlf9_0),.clk(gclk));
	jdff dff_A_6Xgt1Nuk4_0(.dout(w_dff_A_BxZix9QQ3_0),.din(w_dff_A_6Xgt1Nuk4_0),.clk(gclk));
	jdff dff_A_BxZix9QQ3_0(.dout(w_dff_A_FwZWJJCL2_0),.din(w_dff_A_BxZix9QQ3_0),.clk(gclk));
	jdff dff_A_FwZWJJCL2_0(.dout(w_dff_A_lID18ov26_0),.din(w_dff_A_FwZWJJCL2_0),.clk(gclk));
	jdff dff_A_lID18ov26_0(.dout(w_dff_A_AjzjY1pl6_0),.din(w_dff_A_lID18ov26_0),.clk(gclk));
	jdff dff_A_AjzjY1pl6_0(.dout(w_dff_A_oNu8Qi0D7_0),.din(w_dff_A_AjzjY1pl6_0),.clk(gclk));
	jdff dff_A_oNu8Qi0D7_0(.dout(w_dff_A_aZE4mLlt9_0),.din(w_dff_A_oNu8Qi0D7_0),.clk(gclk));
	jdff dff_A_aZE4mLlt9_0(.dout(w_dff_A_bZMU7YKQ7_0),.din(w_dff_A_aZE4mLlt9_0),.clk(gclk));
	jdff dff_A_bZMU7YKQ7_0(.dout(w_dff_A_RR9XyXBC3_0),.din(w_dff_A_bZMU7YKQ7_0),.clk(gclk));
	jdff dff_A_RR9XyXBC3_0(.dout(w_dff_A_wrF4K1iO4_0),.din(w_dff_A_RR9XyXBC3_0),.clk(gclk));
	jdff dff_A_wrF4K1iO4_0(.dout(w_dff_A_x9NQhUqe8_0),.din(w_dff_A_wrF4K1iO4_0),.clk(gclk));
	jdff dff_A_x9NQhUqe8_0(.dout(w_dff_A_gOZDgZ043_0),.din(w_dff_A_x9NQhUqe8_0),.clk(gclk));
	jdff dff_A_gOZDgZ043_0(.dout(w_dff_A_ZjsyHjk21_0),.din(w_dff_A_gOZDgZ043_0),.clk(gclk));
	jdff dff_A_ZjsyHjk21_0(.dout(w_dff_A_S0Qy6RCn4_0),.din(w_dff_A_ZjsyHjk21_0),.clk(gclk));
	jdff dff_A_S0Qy6RCn4_0(.dout(w_dff_A_d9rpGd3U9_0),.din(w_dff_A_S0Qy6RCn4_0),.clk(gclk));
	jdff dff_A_d9rpGd3U9_0(.dout(w_dff_A_BUfKz0sK4_0),.din(w_dff_A_d9rpGd3U9_0),.clk(gclk));
	jdff dff_A_BUfKz0sK4_0(.dout(w_dff_A_xK4mRano6_0),.din(w_dff_A_BUfKz0sK4_0),.clk(gclk));
	jdff dff_A_xK4mRano6_0(.dout(w_dff_A_2RJVWX3P4_0),.din(w_dff_A_xK4mRano6_0),.clk(gclk));
	jdff dff_A_2RJVWX3P4_0(.dout(w_dff_A_KniBZR9T5_0),.din(w_dff_A_2RJVWX3P4_0),.clk(gclk));
	jdff dff_A_KniBZR9T5_0(.dout(w_dff_A_sAHh03771_0),.din(w_dff_A_KniBZR9T5_0),.clk(gclk));
	jdff dff_A_sAHh03771_0(.dout(w_dff_A_iQckNP664_0),.din(w_dff_A_sAHh03771_0),.clk(gclk));
	jdff dff_A_iQckNP664_0(.dout(w_dff_A_v3a1Duhj4_0),.din(w_dff_A_iQckNP664_0),.clk(gclk));
	jdff dff_A_v3a1Duhj4_0(.dout(w_dff_A_KWBqBybj2_0),.din(w_dff_A_v3a1Duhj4_0),.clk(gclk));
	jdff dff_A_KWBqBybj2_0(.dout(w_dff_A_vcCgEMvk3_0),.din(w_dff_A_KWBqBybj2_0),.clk(gclk));
	jdff dff_A_vcCgEMvk3_0(.dout(G453),.din(w_dff_A_vcCgEMvk3_0),.clk(gclk));
	jdff dff_A_EbglPHaX6_2(.dout(w_dff_A_swV84blL3_0),.din(w_dff_A_EbglPHaX6_2),.clk(gclk));
	jdff dff_A_swV84blL3_0(.dout(w_dff_A_MoTpyETq4_0),.din(w_dff_A_swV84blL3_0),.clk(gclk));
	jdff dff_A_MoTpyETq4_0(.dout(w_dff_A_befxaSdt5_0),.din(w_dff_A_MoTpyETq4_0),.clk(gclk));
	jdff dff_A_befxaSdt5_0(.dout(w_dff_A_nj1S3wB41_0),.din(w_dff_A_befxaSdt5_0),.clk(gclk));
	jdff dff_A_nj1S3wB41_0(.dout(w_dff_A_7C4MqCvJ4_0),.din(w_dff_A_nj1S3wB41_0),.clk(gclk));
	jdff dff_A_7C4MqCvJ4_0(.dout(w_dff_A_NJpT3PZq6_0),.din(w_dff_A_7C4MqCvJ4_0),.clk(gclk));
	jdff dff_A_NJpT3PZq6_0(.dout(w_dff_A_rUUp3FX02_0),.din(w_dff_A_NJpT3PZq6_0),.clk(gclk));
	jdff dff_A_rUUp3FX02_0(.dout(w_dff_A_fSutrgXe6_0),.din(w_dff_A_rUUp3FX02_0),.clk(gclk));
	jdff dff_A_fSutrgXe6_0(.dout(w_dff_A_VgcIlFzG8_0),.din(w_dff_A_fSutrgXe6_0),.clk(gclk));
	jdff dff_A_VgcIlFzG8_0(.dout(w_dff_A_69izWaog9_0),.din(w_dff_A_VgcIlFzG8_0),.clk(gclk));
	jdff dff_A_69izWaog9_0(.dout(w_dff_A_Cdzp4wZp7_0),.din(w_dff_A_69izWaog9_0),.clk(gclk));
	jdff dff_A_Cdzp4wZp7_0(.dout(w_dff_A_virqKLAN5_0),.din(w_dff_A_Cdzp4wZp7_0),.clk(gclk));
	jdff dff_A_virqKLAN5_0(.dout(w_dff_A_5ENM3xos9_0),.din(w_dff_A_virqKLAN5_0),.clk(gclk));
	jdff dff_A_5ENM3xos9_0(.dout(w_dff_A_V2tqs1vF0_0),.din(w_dff_A_5ENM3xos9_0),.clk(gclk));
	jdff dff_A_V2tqs1vF0_0(.dout(w_dff_A_wk30Ygv81_0),.din(w_dff_A_V2tqs1vF0_0),.clk(gclk));
	jdff dff_A_wk30Ygv81_0(.dout(w_dff_A_110pMlfj1_0),.din(w_dff_A_wk30Ygv81_0),.clk(gclk));
	jdff dff_A_110pMlfj1_0(.dout(w_dff_A_hWdkipOI8_0),.din(w_dff_A_110pMlfj1_0),.clk(gclk));
	jdff dff_A_hWdkipOI8_0(.dout(w_dff_A_GQm3qUCT1_0),.din(w_dff_A_hWdkipOI8_0),.clk(gclk));
	jdff dff_A_GQm3qUCT1_0(.dout(w_dff_A_iIUXtAtb7_0),.din(w_dff_A_GQm3qUCT1_0),.clk(gclk));
	jdff dff_A_iIUXtAtb7_0(.dout(w_dff_A_ZsJAKTfe5_0),.din(w_dff_A_iIUXtAtb7_0),.clk(gclk));
	jdff dff_A_ZsJAKTfe5_0(.dout(w_dff_A_qXeYCbkh8_0),.din(w_dff_A_ZsJAKTfe5_0),.clk(gclk));
	jdff dff_A_qXeYCbkh8_0(.dout(w_dff_A_RFNpAnF93_0),.din(w_dff_A_qXeYCbkh8_0),.clk(gclk));
	jdff dff_A_RFNpAnF93_0(.dout(w_dff_A_EjXHQbSF4_0),.din(w_dff_A_RFNpAnF93_0),.clk(gclk));
	jdff dff_A_EjXHQbSF4_0(.dout(w_dff_A_40eeJVPZ1_0),.din(w_dff_A_EjXHQbSF4_0),.clk(gclk));
	jdff dff_A_40eeJVPZ1_0(.dout(w_dff_A_5QtKENZk9_0),.din(w_dff_A_40eeJVPZ1_0),.clk(gclk));
	jdff dff_A_5QtKENZk9_0(.dout(w_dff_A_wkcGo9BV7_0),.din(w_dff_A_5QtKENZk9_0),.clk(gclk));
	jdff dff_A_wkcGo9BV7_0(.dout(w_dff_A_Oit6hlsp3_0),.din(w_dff_A_wkcGo9BV7_0),.clk(gclk));
	jdff dff_A_Oit6hlsp3_0(.dout(w_dff_A_RmnDTltQ2_0),.din(w_dff_A_Oit6hlsp3_0),.clk(gclk));
	jdff dff_A_RmnDTltQ2_0(.dout(w_dff_A_EtNNyMz02_0),.din(w_dff_A_RmnDTltQ2_0),.clk(gclk));
	jdff dff_A_EtNNyMz02_0(.dout(w_dff_A_rIrObztX0_0),.din(w_dff_A_EtNNyMz02_0),.clk(gclk));
	jdff dff_A_rIrObztX0_0(.dout(w_dff_A_9dE3pU650_0),.din(w_dff_A_rIrObztX0_0),.clk(gclk));
	jdff dff_A_9dE3pU650_0(.dout(w_dff_A_6L9Z9La10_0),.din(w_dff_A_9dE3pU650_0),.clk(gclk));
	jdff dff_A_6L9Z9La10_0(.dout(w_dff_A_rfwuTdbL8_0),.din(w_dff_A_6L9Z9La10_0),.clk(gclk));
	jdff dff_A_rfwuTdbL8_0(.dout(w_dff_A_XcD2rOzf0_0),.din(w_dff_A_rfwuTdbL8_0),.clk(gclk));
	jdff dff_A_XcD2rOzf0_0(.dout(w_dff_A_siWTAYaz3_0),.din(w_dff_A_XcD2rOzf0_0),.clk(gclk));
	jdff dff_A_siWTAYaz3_0(.dout(w_dff_A_POP02OC74_0),.din(w_dff_A_siWTAYaz3_0),.clk(gclk));
	jdff dff_A_POP02OC74_0(.dout(w_dff_A_rz4eBgoh6_0),.din(w_dff_A_POP02OC74_0),.clk(gclk));
	jdff dff_A_rz4eBgoh6_0(.dout(G278),.din(w_dff_A_rz4eBgoh6_0),.clk(gclk));
	jdff dff_A_S8QuRzkE0_2(.dout(w_dff_A_dseyb2v74_0),.din(w_dff_A_S8QuRzkE0_2),.clk(gclk));
	jdff dff_A_dseyb2v74_0(.dout(w_dff_A_OUFirTFu9_0),.din(w_dff_A_dseyb2v74_0),.clk(gclk));
	jdff dff_A_OUFirTFu9_0(.dout(w_dff_A_0TFd1sSJ4_0),.din(w_dff_A_OUFirTFu9_0),.clk(gclk));
	jdff dff_A_0TFd1sSJ4_0(.dout(w_dff_A_kXRCpNYU6_0),.din(w_dff_A_0TFd1sSJ4_0),.clk(gclk));
	jdff dff_A_kXRCpNYU6_0(.dout(w_dff_A_YUdKZbFq6_0),.din(w_dff_A_kXRCpNYU6_0),.clk(gclk));
	jdff dff_A_YUdKZbFq6_0(.dout(w_dff_A_W5OsBaa58_0),.din(w_dff_A_YUdKZbFq6_0),.clk(gclk));
	jdff dff_A_W5OsBaa58_0(.dout(w_dff_A_uu9vKEwQ8_0),.din(w_dff_A_W5OsBaa58_0),.clk(gclk));
	jdff dff_A_uu9vKEwQ8_0(.dout(w_dff_A_FMlwMk116_0),.din(w_dff_A_uu9vKEwQ8_0),.clk(gclk));
	jdff dff_A_FMlwMk116_0(.dout(w_dff_A_XAK0UxfS4_0),.din(w_dff_A_FMlwMk116_0),.clk(gclk));
	jdff dff_A_XAK0UxfS4_0(.dout(w_dff_A_fvgllW6Q1_0),.din(w_dff_A_XAK0UxfS4_0),.clk(gclk));
	jdff dff_A_fvgllW6Q1_0(.dout(w_dff_A_XCi5mrWq6_0),.din(w_dff_A_fvgllW6Q1_0),.clk(gclk));
	jdff dff_A_XCi5mrWq6_0(.dout(w_dff_A_vMeoGz8n2_0),.din(w_dff_A_XCi5mrWq6_0),.clk(gclk));
	jdff dff_A_vMeoGz8n2_0(.dout(w_dff_A_0Bdpm1em9_0),.din(w_dff_A_vMeoGz8n2_0),.clk(gclk));
	jdff dff_A_0Bdpm1em9_0(.dout(w_dff_A_3nVUNd1z4_0),.din(w_dff_A_0Bdpm1em9_0),.clk(gclk));
	jdff dff_A_3nVUNd1z4_0(.dout(w_dff_A_q6yS1vd01_0),.din(w_dff_A_3nVUNd1z4_0),.clk(gclk));
	jdff dff_A_q6yS1vd01_0(.dout(w_dff_A_VeUuPMa17_0),.din(w_dff_A_q6yS1vd01_0),.clk(gclk));
	jdff dff_A_VeUuPMa17_0(.dout(w_dff_A_XNT9SGAd2_0),.din(w_dff_A_VeUuPMa17_0),.clk(gclk));
	jdff dff_A_XNT9SGAd2_0(.dout(w_dff_A_x7xCGkqj3_0),.din(w_dff_A_XNT9SGAd2_0),.clk(gclk));
	jdff dff_A_x7xCGkqj3_0(.dout(w_dff_A_T0wCi8o12_0),.din(w_dff_A_x7xCGkqj3_0),.clk(gclk));
	jdff dff_A_T0wCi8o12_0(.dout(w_dff_A_Cely64dP6_0),.din(w_dff_A_T0wCi8o12_0),.clk(gclk));
	jdff dff_A_Cely64dP6_0(.dout(w_dff_A_nrExZfeL0_0),.din(w_dff_A_Cely64dP6_0),.clk(gclk));
	jdff dff_A_nrExZfeL0_0(.dout(w_dff_A_rQYLfaUN2_0),.din(w_dff_A_nrExZfeL0_0),.clk(gclk));
	jdff dff_A_rQYLfaUN2_0(.dout(w_dff_A_12TaG0F05_0),.din(w_dff_A_rQYLfaUN2_0),.clk(gclk));
	jdff dff_A_12TaG0F05_0(.dout(w_dff_A_5a9NCTDT6_0),.din(w_dff_A_12TaG0F05_0),.clk(gclk));
	jdff dff_A_5a9NCTDT6_0(.dout(w_dff_A_aFXjbadQ2_0),.din(w_dff_A_5a9NCTDT6_0),.clk(gclk));
	jdff dff_A_aFXjbadQ2_0(.dout(w_dff_A_BBfr5o794_0),.din(w_dff_A_aFXjbadQ2_0),.clk(gclk));
	jdff dff_A_BBfr5o794_0(.dout(w_dff_A_B5YKQYA75_0),.din(w_dff_A_BBfr5o794_0),.clk(gclk));
	jdff dff_A_B5YKQYA75_0(.dout(w_dff_A_tHYkYDFq7_0),.din(w_dff_A_B5YKQYA75_0),.clk(gclk));
	jdff dff_A_tHYkYDFq7_0(.dout(w_dff_A_OxPfMyx55_0),.din(w_dff_A_tHYkYDFq7_0),.clk(gclk));
	jdff dff_A_OxPfMyx55_0(.dout(w_dff_A_MvRVSvZU6_0),.din(w_dff_A_OxPfMyx55_0),.clk(gclk));
	jdff dff_A_MvRVSvZU6_0(.dout(w_dff_A_T99Xbd8v0_0),.din(w_dff_A_MvRVSvZU6_0),.clk(gclk));
	jdff dff_A_T99Xbd8v0_0(.dout(w_dff_A_0ioXxkSG6_0),.din(w_dff_A_T99Xbd8v0_0),.clk(gclk));
	jdff dff_A_0ioXxkSG6_0(.dout(G373),.din(w_dff_A_0ioXxkSG6_0),.clk(gclk));
	jdff dff_A_C7Y9DVay5_2(.dout(w_dff_A_nzl4gXeX9_0),.din(w_dff_A_C7Y9DVay5_2),.clk(gclk));
	jdff dff_A_nzl4gXeX9_0(.dout(w_dff_A_H3VhH1vY2_0),.din(w_dff_A_nzl4gXeX9_0),.clk(gclk));
	jdff dff_A_H3VhH1vY2_0(.dout(w_dff_A_JZLqlW553_0),.din(w_dff_A_H3VhH1vY2_0),.clk(gclk));
	jdff dff_A_JZLqlW553_0(.dout(w_dff_A_kfVPIFvh6_0),.din(w_dff_A_JZLqlW553_0),.clk(gclk));
	jdff dff_A_kfVPIFvh6_0(.dout(w_dff_A_xZOhCyG66_0),.din(w_dff_A_kfVPIFvh6_0),.clk(gclk));
	jdff dff_A_xZOhCyG66_0(.dout(w_dff_A_enRZMrRj2_0),.din(w_dff_A_xZOhCyG66_0),.clk(gclk));
	jdff dff_A_enRZMrRj2_0(.dout(w_dff_A_5ULdjhRT0_0),.din(w_dff_A_enRZMrRj2_0),.clk(gclk));
	jdff dff_A_5ULdjhRT0_0(.dout(w_dff_A_ViaN4srH4_0),.din(w_dff_A_5ULdjhRT0_0),.clk(gclk));
	jdff dff_A_ViaN4srH4_0(.dout(w_dff_A_9D32lsUc0_0),.din(w_dff_A_ViaN4srH4_0),.clk(gclk));
	jdff dff_A_9D32lsUc0_0(.dout(w_dff_A_xeF3ArdW7_0),.din(w_dff_A_9D32lsUc0_0),.clk(gclk));
	jdff dff_A_xeF3ArdW7_0(.dout(G258),.din(w_dff_A_xeF3ArdW7_0),.clk(gclk));
	jdff dff_A_6veNz4KY3_2(.dout(w_dff_A_9HZvrbM50_0),.din(w_dff_A_6veNz4KY3_2),.clk(gclk));
	jdff dff_A_9HZvrbM50_0(.dout(w_dff_A_Iofqhzvn3_0),.din(w_dff_A_9HZvrbM50_0),.clk(gclk));
	jdff dff_A_Iofqhzvn3_0(.dout(w_dff_A_Rpdsh7GX8_0),.din(w_dff_A_Iofqhzvn3_0),.clk(gclk));
	jdff dff_A_Rpdsh7GX8_0(.dout(w_dff_A_ShHN4Y151_0),.din(w_dff_A_Rpdsh7GX8_0),.clk(gclk));
	jdff dff_A_ShHN4Y151_0(.dout(w_dff_A_KT01SSCm0_0),.din(w_dff_A_ShHN4Y151_0),.clk(gclk));
	jdff dff_A_KT01SSCm0_0(.dout(w_dff_A_jUpYjNDe8_0),.din(w_dff_A_KT01SSCm0_0),.clk(gclk));
	jdff dff_A_jUpYjNDe8_0(.dout(w_dff_A_koFrxztT6_0),.din(w_dff_A_jUpYjNDe8_0),.clk(gclk));
	jdff dff_A_koFrxztT6_0(.dout(w_dff_A_Q3yJPoNu6_0),.din(w_dff_A_koFrxztT6_0),.clk(gclk));
	jdff dff_A_Q3yJPoNu6_0(.dout(w_dff_A_jfYRn6PI6_0),.din(w_dff_A_Q3yJPoNu6_0),.clk(gclk));
	jdff dff_A_jfYRn6PI6_0(.dout(w_dff_A_pJJ0Ihlt6_0),.din(w_dff_A_jfYRn6PI6_0),.clk(gclk));
	jdff dff_A_pJJ0Ihlt6_0(.dout(G264),.din(w_dff_A_pJJ0Ihlt6_0),.clk(gclk));
	jdff dff_A_oa0XxNvS3_2(.dout(w_dff_A_bB4avgpf0_0),.din(w_dff_A_oa0XxNvS3_2),.clk(gclk));
	jdff dff_A_bB4avgpf0_0(.dout(w_dff_A_Nt3WlxA69_0),.din(w_dff_A_bB4avgpf0_0),.clk(gclk));
	jdff dff_A_Nt3WlxA69_0(.dout(w_dff_A_IzCSaNRG4_0),.din(w_dff_A_Nt3WlxA69_0),.clk(gclk));
	jdff dff_A_IzCSaNRG4_0(.dout(w_dff_A_VqUfarth3_0),.din(w_dff_A_IzCSaNRG4_0),.clk(gclk));
	jdff dff_A_VqUfarth3_0(.dout(w_dff_A_CP0LNn3C8_0),.din(w_dff_A_VqUfarth3_0),.clk(gclk));
	jdff dff_A_CP0LNn3C8_0(.dout(w_dff_A_wBzVYZfD6_0),.din(w_dff_A_CP0LNn3C8_0),.clk(gclk));
	jdff dff_A_wBzVYZfD6_0(.dout(w_dff_A_Wko3XSpy7_0),.din(w_dff_A_wBzVYZfD6_0),.clk(gclk));
	jdff dff_A_Wko3XSpy7_0(.dout(w_dff_A_M0lcvcBX0_0),.din(w_dff_A_Wko3XSpy7_0),.clk(gclk));
	jdff dff_A_M0lcvcBX0_0(.dout(w_dff_A_yFOsYNUg9_0),.din(w_dff_A_M0lcvcBX0_0),.clk(gclk));
	jdff dff_A_yFOsYNUg9_0(.dout(w_dff_A_NED2kRvc1_0),.din(w_dff_A_yFOsYNUg9_0),.clk(gclk));
	jdff dff_A_NED2kRvc1_0(.dout(w_dff_A_Y3lDAcRw4_0),.din(w_dff_A_NED2kRvc1_0),.clk(gclk));
	jdff dff_A_Y3lDAcRw4_0(.dout(w_dff_A_jOZt3TJ25_0),.din(w_dff_A_Y3lDAcRw4_0),.clk(gclk));
	jdff dff_A_jOZt3TJ25_0(.dout(w_dff_A_JERUK1X57_0),.din(w_dff_A_jOZt3TJ25_0),.clk(gclk));
	jdff dff_A_JERUK1X57_0(.dout(w_dff_A_Ngvebk253_0),.din(w_dff_A_JERUK1X57_0),.clk(gclk));
	jdff dff_A_Ngvebk253_0(.dout(w_dff_A_w1ntX4QK4_0),.din(w_dff_A_Ngvebk253_0),.clk(gclk));
	jdff dff_A_w1ntX4QK4_0(.dout(w_dff_A_AYdDzrQq9_0),.din(w_dff_A_w1ntX4QK4_0),.clk(gclk));
	jdff dff_A_AYdDzrQq9_0(.dout(w_dff_A_hToYVN4Y9_0),.din(w_dff_A_AYdDzrQq9_0),.clk(gclk));
	jdff dff_A_hToYVN4Y9_0(.dout(w_dff_A_mcyC9mh01_0),.din(w_dff_A_hToYVN4Y9_0),.clk(gclk));
	jdff dff_A_mcyC9mh01_0(.dout(w_dff_A_KuuqqpVz0_0),.din(w_dff_A_mcyC9mh01_0),.clk(gclk));
	jdff dff_A_KuuqqpVz0_0(.dout(w_dff_A_cBOkQEx37_0),.din(w_dff_A_KuuqqpVz0_0),.clk(gclk));
	jdff dff_A_cBOkQEx37_0(.dout(w_dff_A_NXSWMPmp2_0),.din(w_dff_A_cBOkQEx37_0),.clk(gclk));
	jdff dff_A_NXSWMPmp2_0(.dout(w_dff_A_ftUV2bVH7_0),.din(w_dff_A_NXSWMPmp2_0),.clk(gclk));
	jdff dff_A_ftUV2bVH7_0(.dout(w_dff_A_sdKYZNvW4_0),.din(w_dff_A_ftUV2bVH7_0),.clk(gclk));
	jdff dff_A_sdKYZNvW4_0(.dout(w_dff_A_Ij8AChXO0_0),.din(w_dff_A_sdKYZNvW4_0),.clk(gclk));
	jdff dff_A_Ij8AChXO0_0(.dout(G388),.din(w_dff_A_Ij8AChXO0_0),.clk(gclk));
	jdff dff_A_NyvscHrC9_2(.dout(w_dff_A_x8uJ3uU14_0),.din(w_dff_A_NyvscHrC9_2),.clk(gclk));
	jdff dff_A_x8uJ3uU14_0(.dout(w_dff_A_uWUq719U4_0),.din(w_dff_A_x8uJ3uU14_0),.clk(gclk));
	jdff dff_A_uWUq719U4_0(.dout(w_dff_A_Ra96J6TQ9_0),.din(w_dff_A_uWUq719U4_0),.clk(gclk));
	jdff dff_A_Ra96J6TQ9_0(.dout(w_dff_A_oYmIiRKo1_0),.din(w_dff_A_Ra96J6TQ9_0),.clk(gclk));
	jdff dff_A_oYmIiRKo1_0(.dout(w_dff_A_Ag0jBzgQ0_0),.din(w_dff_A_oYmIiRKo1_0),.clk(gclk));
	jdff dff_A_Ag0jBzgQ0_0(.dout(w_dff_A_6y2qeYlc9_0),.din(w_dff_A_Ag0jBzgQ0_0),.clk(gclk));
	jdff dff_A_6y2qeYlc9_0(.dout(w_dff_A_63ytucfX7_0),.din(w_dff_A_6y2qeYlc9_0),.clk(gclk));
	jdff dff_A_63ytucfX7_0(.dout(w_dff_A_DV8plbpk4_0),.din(w_dff_A_63ytucfX7_0),.clk(gclk));
	jdff dff_A_DV8plbpk4_0(.dout(w_dff_A_D56M6mj31_0),.din(w_dff_A_DV8plbpk4_0),.clk(gclk));
	jdff dff_A_D56M6mj31_0(.dout(w_dff_A_7vvA95Gx0_0),.din(w_dff_A_D56M6mj31_0),.clk(gclk));
	jdff dff_A_7vvA95Gx0_0(.dout(w_dff_A_7Pro7rEs1_0),.din(w_dff_A_7vvA95Gx0_0),.clk(gclk));
	jdff dff_A_7Pro7rEs1_0(.dout(w_dff_A_I7WGF6fh4_0),.din(w_dff_A_7Pro7rEs1_0),.clk(gclk));
	jdff dff_A_I7WGF6fh4_0(.dout(w_dff_A_QpadcRY80_0),.din(w_dff_A_I7WGF6fh4_0),.clk(gclk));
	jdff dff_A_QpadcRY80_0(.dout(w_dff_A_l7Pn9xLV6_0),.din(w_dff_A_QpadcRY80_0),.clk(gclk));
	jdff dff_A_l7Pn9xLV6_0(.dout(w_dff_A_sdWqi4Go1_0),.din(w_dff_A_l7Pn9xLV6_0),.clk(gclk));
	jdff dff_A_sdWqi4Go1_0(.dout(w_dff_A_oz2mxFWJ6_0),.din(w_dff_A_sdWqi4Go1_0),.clk(gclk));
	jdff dff_A_oz2mxFWJ6_0(.dout(w_dff_A_UDnVxWWn3_0),.din(w_dff_A_oz2mxFWJ6_0),.clk(gclk));
	jdff dff_A_UDnVxWWn3_0(.dout(w_dff_A_AldomAwp8_0),.din(w_dff_A_UDnVxWWn3_0),.clk(gclk));
	jdff dff_A_AldomAwp8_0(.dout(w_dff_A_8gjEDqU79_0),.din(w_dff_A_AldomAwp8_0),.clk(gclk));
	jdff dff_A_8gjEDqU79_0(.dout(w_dff_A_F6GX7V5k7_0),.din(w_dff_A_8gjEDqU79_0),.clk(gclk));
	jdff dff_A_F6GX7V5k7_0(.dout(w_dff_A_ylmtbOf76_0),.din(w_dff_A_F6GX7V5k7_0),.clk(gclk));
	jdff dff_A_ylmtbOf76_0(.dout(w_dff_A_rXriJFTA6_0),.din(w_dff_A_ylmtbOf76_0),.clk(gclk));
	jdff dff_A_rXriJFTA6_0(.dout(w_dff_A_I33HmPdM2_0),.din(w_dff_A_rXriJFTA6_0),.clk(gclk));
	jdff dff_A_I33HmPdM2_0(.dout(w_dff_A_fjmmPZfX7_0),.din(w_dff_A_I33HmPdM2_0),.clk(gclk));
	jdff dff_A_fjmmPZfX7_0(.dout(w_dff_A_rPh0qnnX6_0),.din(w_dff_A_fjmmPZfX7_0),.clk(gclk));
	jdff dff_A_rPh0qnnX6_0(.dout(w_dff_A_MLSieQRb5_0),.din(w_dff_A_rPh0qnnX6_0),.clk(gclk));
	jdff dff_A_MLSieQRb5_0(.dout(G391),.din(w_dff_A_MLSieQRb5_0),.clk(gclk));
	jdff dff_A_lPzfP2la9_2(.dout(w_dff_A_VEC37Kb97_0),.din(w_dff_A_lPzfP2la9_2),.clk(gclk));
	jdff dff_A_VEC37Kb97_0(.dout(w_dff_A_yKwTG61T1_0),.din(w_dff_A_VEC37Kb97_0),.clk(gclk));
	jdff dff_A_yKwTG61T1_0(.dout(w_dff_A_U29S5hfu4_0),.din(w_dff_A_yKwTG61T1_0),.clk(gclk));
	jdff dff_A_U29S5hfu4_0(.dout(w_dff_A_v6cvdGue5_0),.din(w_dff_A_U29S5hfu4_0),.clk(gclk));
	jdff dff_A_v6cvdGue5_0(.dout(w_dff_A_PgLsNzlD8_0),.din(w_dff_A_v6cvdGue5_0),.clk(gclk));
	jdff dff_A_PgLsNzlD8_0(.dout(w_dff_A_IwHeJo6u7_0),.din(w_dff_A_PgLsNzlD8_0),.clk(gclk));
	jdff dff_A_IwHeJo6u7_0(.dout(w_dff_A_eepxyCLY5_0),.din(w_dff_A_IwHeJo6u7_0),.clk(gclk));
	jdff dff_A_eepxyCLY5_0(.dout(w_dff_A_KoOHLsFp7_0),.din(w_dff_A_eepxyCLY5_0),.clk(gclk));
	jdff dff_A_KoOHLsFp7_0(.dout(w_dff_A_GeuJQvZH1_0),.din(w_dff_A_KoOHLsFp7_0),.clk(gclk));
	jdff dff_A_GeuJQvZH1_0(.dout(w_dff_A_w9WqPI5b7_0),.din(w_dff_A_GeuJQvZH1_0),.clk(gclk));
	jdff dff_A_w9WqPI5b7_0(.dout(w_dff_A_h6KY3otM4_0),.din(w_dff_A_w9WqPI5b7_0),.clk(gclk));
	jdff dff_A_h6KY3otM4_0(.dout(w_dff_A_pQXfIaEc7_0),.din(w_dff_A_h6KY3otM4_0),.clk(gclk));
	jdff dff_A_pQXfIaEc7_0(.dout(w_dff_A_OGfNbo279_0),.din(w_dff_A_pQXfIaEc7_0),.clk(gclk));
	jdff dff_A_OGfNbo279_0(.dout(w_dff_A_OPysQK8j9_0),.din(w_dff_A_OGfNbo279_0),.clk(gclk));
	jdff dff_A_OPysQK8j9_0(.dout(w_dff_A_YKfG7xbx4_0),.din(w_dff_A_OPysQK8j9_0),.clk(gclk));
	jdff dff_A_YKfG7xbx4_0(.dout(w_dff_A_046HKjwD5_0),.din(w_dff_A_YKfG7xbx4_0),.clk(gclk));
	jdff dff_A_046HKjwD5_0(.dout(w_dff_A_nyu2S2zC0_0),.din(w_dff_A_046HKjwD5_0),.clk(gclk));
	jdff dff_A_nyu2S2zC0_0(.dout(w_dff_A_8ePTkFr49_0),.din(w_dff_A_nyu2S2zC0_0),.clk(gclk));
	jdff dff_A_8ePTkFr49_0(.dout(w_dff_A_Efgp4oSm6_0),.din(w_dff_A_8ePTkFr49_0),.clk(gclk));
	jdff dff_A_Efgp4oSm6_0(.dout(w_dff_A_6fJC1h071_0),.din(w_dff_A_Efgp4oSm6_0),.clk(gclk));
	jdff dff_A_6fJC1h071_0(.dout(w_dff_A_948eRYST5_0),.din(w_dff_A_6fJC1h071_0),.clk(gclk));
	jdff dff_A_948eRYST5_0(.dout(w_dff_A_0Ee2ZB4q3_0),.din(w_dff_A_948eRYST5_0),.clk(gclk));
	jdff dff_A_0Ee2ZB4q3_0(.dout(w_dff_A_s3R6TkFj3_0),.din(w_dff_A_0Ee2ZB4q3_0),.clk(gclk));
	jdff dff_A_s3R6TkFj3_0(.dout(w_dff_A_zKOEIkDr2_0),.din(w_dff_A_s3R6TkFj3_0),.clk(gclk));
	jdff dff_A_zKOEIkDr2_0(.dout(w_dff_A_2z1wE9Tr7_0),.din(w_dff_A_zKOEIkDr2_0),.clk(gclk));
	jdff dff_A_2z1wE9Tr7_0(.dout(w_dff_A_CreCEGnX4_0),.din(w_dff_A_2z1wE9Tr7_0),.clk(gclk));
	jdff dff_A_CreCEGnX4_0(.dout(w_dff_A_ZVuNEt8t7_0),.din(w_dff_A_CreCEGnX4_0),.clk(gclk));
	jdff dff_A_ZVuNEt8t7_0(.dout(w_dff_A_IQkVbZHN5_0),.din(w_dff_A_ZVuNEt8t7_0),.clk(gclk));
	jdff dff_A_IQkVbZHN5_0(.dout(w_dff_A_tL4B5Qt22_0),.din(w_dff_A_IQkVbZHN5_0),.clk(gclk));
	jdff dff_A_tL4B5Qt22_0(.dout(G394),.din(w_dff_A_tL4B5Qt22_0),.clk(gclk));
	jdff dff_A_JmJfu1Jx3_2(.dout(w_dff_A_prcnguFT9_0),.din(w_dff_A_JmJfu1Jx3_2),.clk(gclk));
	jdff dff_A_prcnguFT9_0(.dout(w_dff_A_XKV3xiQI6_0),.din(w_dff_A_prcnguFT9_0),.clk(gclk));
	jdff dff_A_XKV3xiQI6_0(.dout(w_dff_A_sfGrFQKw2_0),.din(w_dff_A_XKV3xiQI6_0),.clk(gclk));
	jdff dff_A_sfGrFQKw2_0(.dout(w_dff_A_1TmbwBDk6_0),.din(w_dff_A_sfGrFQKw2_0),.clk(gclk));
	jdff dff_A_1TmbwBDk6_0(.dout(w_dff_A_GlJUvyaM9_0),.din(w_dff_A_1TmbwBDk6_0),.clk(gclk));
	jdff dff_A_GlJUvyaM9_0(.dout(w_dff_A_4vpgJdKb8_0),.din(w_dff_A_GlJUvyaM9_0),.clk(gclk));
	jdff dff_A_4vpgJdKb8_0(.dout(w_dff_A_E6RaSHGq9_0),.din(w_dff_A_4vpgJdKb8_0),.clk(gclk));
	jdff dff_A_E6RaSHGq9_0(.dout(w_dff_A_Z5vwzN8A5_0),.din(w_dff_A_E6RaSHGq9_0),.clk(gclk));
	jdff dff_A_Z5vwzN8A5_0(.dout(w_dff_A_HaUUTyqT3_0),.din(w_dff_A_Z5vwzN8A5_0),.clk(gclk));
	jdff dff_A_HaUUTyqT3_0(.dout(w_dff_A_Oqd4VR4j8_0),.din(w_dff_A_HaUUTyqT3_0),.clk(gclk));
	jdff dff_A_Oqd4VR4j8_0(.dout(w_dff_A_XrCT66DO4_0),.din(w_dff_A_Oqd4VR4j8_0),.clk(gclk));
	jdff dff_A_XrCT66DO4_0(.dout(w_dff_A_fD6h7s5w5_0),.din(w_dff_A_XrCT66DO4_0),.clk(gclk));
	jdff dff_A_fD6h7s5w5_0(.dout(w_dff_A_sBgo36vb4_0),.din(w_dff_A_fD6h7s5w5_0),.clk(gclk));
	jdff dff_A_sBgo36vb4_0(.dout(w_dff_A_P6AVwomB9_0),.din(w_dff_A_sBgo36vb4_0),.clk(gclk));
	jdff dff_A_P6AVwomB9_0(.dout(w_dff_A_LGhfym0w3_0),.din(w_dff_A_P6AVwomB9_0),.clk(gclk));
	jdff dff_A_LGhfym0w3_0(.dout(w_dff_A_ismxpB1d4_0),.din(w_dff_A_LGhfym0w3_0),.clk(gclk));
	jdff dff_A_ismxpB1d4_0(.dout(w_dff_A_Qa4lUHWV6_0),.din(w_dff_A_ismxpB1d4_0),.clk(gclk));
	jdff dff_A_Qa4lUHWV6_0(.dout(w_dff_A_P5bnf5xA4_0),.din(w_dff_A_Qa4lUHWV6_0),.clk(gclk));
	jdff dff_A_P5bnf5xA4_0(.dout(w_dff_A_TLWD8j7q8_0),.din(w_dff_A_P5bnf5xA4_0),.clk(gclk));
	jdff dff_A_TLWD8j7q8_0(.dout(w_dff_A_PmPFXRkm5_0),.din(w_dff_A_TLWD8j7q8_0),.clk(gclk));
	jdff dff_A_PmPFXRkm5_0(.dout(w_dff_A_1DEqSVSh8_0),.din(w_dff_A_PmPFXRkm5_0),.clk(gclk));
	jdff dff_A_1DEqSVSh8_0(.dout(w_dff_A_hvLRLS7Y4_0),.din(w_dff_A_1DEqSVSh8_0),.clk(gclk));
	jdff dff_A_hvLRLS7Y4_0(.dout(w_dff_A_hBdyxDej5_0),.din(w_dff_A_hvLRLS7Y4_0),.clk(gclk));
	jdff dff_A_hBdyxDej5_0(.dout(w_dff_A_uVOIUjPU9_0),.din(w_dff_A_hBdyxDej5_0),.clk(gclk));
	jdff dff_A_uVOIUjPU9_0(.dout(w_dff_A_LcmR00Rp7_0),.din(w_dff_A_uVOIUjPU9_0),.clk(gclk));
	jdff dff_A_LcmR00Rp7_0(.dout(w_dff_A_RLqxLHBO8_0),.din(w_dff_A_LcmR00Rp7_0),.clk(gclk));
	jdff dff_A_RLqxLHBO8_0(.dout(w_dff_A_nTjrgZKe8_0),.din(w_dff_A_RLqxLHBO8_0),.clk(gclk));
	jdff dff_A_nTjrgZKe8_0(.dout(w_dff_A_FFcBnvFW4_0),.din(w_dff_A_nTjrgZKe8_0),.clk(gclk));
	jdff dff_A_FFcBnvFW4_0(.dout(w_dff_A_TQEAN2BS3_0),.din(w_dff_A_FFcBnvFW4_0),.clk(gclk));
	jdff dff_A_TQEAN2BS3_0(.dout(w_dff_A_yAlJLw6x9_0),.din(w_dff_A_TQEAN2BS3_0),.clk(gclk));
	jdff dff_A_yAlJLw6x9_0(.dout(G397),.din(w_dff_A_yAlJLw6x9_0),.clk(gclk));
	jdff dff_A_SGZG573Y4_2(.dout(w_dff_A_9mPUOZh00_0),.din(w_dff_A_SGZG573Y4_2),.clk(gclk));
	jdff dff_A_9mPUOZh00_0(.dout(w_dff_A_Jnwu2Yhf4_0),.din(w_dff_A_9mPUOZh00_0),.clk(gclk));
	jdff dff_A_Jnwu2Yhf4_0(.dout(w_dff_A_joi2S2HD0_0),.din(w_dff_A_Jnwu2Yhf4_0),.clk(gclk));
	jdff dff_A_joi2S2HD0_0(.dout(w_dff_A_Jr2FxMJX9_0),.din(w_dff_A_joi2S2HD0_0),.clk(gclk));
	jdff dff_A_Jr2FxMJX9_0(.dout(w_dff_A_qzv6Kkxg3_0),.din(w_dff_A_Jr2FxMJX9_0),.clk(gclk));
	jdff dff_A_qzv6Kkxg3_0(.dout(w_dff_A_rov2lSPR2_0),.din(w_dff_A_qzv6Kkxg3_0),.clk(gclk));
	jdff dff_A_rov2lSPR2_0(.dout(w_dff_A_QmAp1mWZ8_0),.din(w_dff_A_rov2lSPR2_0),.clk(gclk));
	jdff dff_A_QmAp1mWZ8_0(.dout(w_dff_A_QZwkynxl6_0),.din(w_dff_A_QmAp1mWZ8_0),.clk(gclk));
	jdff dff_A_QZwkynxl6_0(.dout(w_dff_A_Iu7M7jYm4_0),.din(w_dff_A_QZwkynxl6_0),.clk(gclk));
	jdff dff_A_Iu7M7jYm4_0(.dout(w_dff_A_pOGcSKCK9_0),.din(w_dff_A_Iu7M7jYm4_0),.clk(gclk));
	jdff dff_A_pOGcSKCK9_0(.dout(w_dff_A_mYyUNWY12_0),.din(w_dff_A_pOGcSKCK9_0),.clk(gclk));
	jdff dff_A_mYyUNWY12_0(.dout(w_dff_A_dSTkFMBC4_0),.din(w_dff_A_mYyUNWY12_0),.clk(gclk));
	jdff dff_A_dSTkFMBC4_0(.dout(w_dff_A_fJTZhBr26_0),.din(w_dff_A_dSTkFMBC4_0),.clk(gclk));
	jdff dff_A_fJTZhBr26_0(.dout(w_dff_A_5JsqUKxw8_0),.din(w_dff_A_fJTZhBr26_0),.clk(gclk));
	jdff dff_A_5JsqUKxw8_0(.dout(w_dff_A_3Rh7J9tu3_0),.din(w_dff_A_5JsqUKxw8_0),.clk(gclk));
	jdff dff_A_3Rh7J9tu3_0(.dout(w_dff_A_bnz3u5M11_0),.din(w_dff_A_3Rh7J9tu3_0),.clk(gclk));
	jdff dff_A_bnz3u5M11_0(.dout(w_dff_A_xMdH4bvC6_0),.din(w_dff_A_bnz3u5M11_0),.clk(gclk));
	jdff dff_A_xMdH4bvC6_0(.dout(w_dff_A_w14rmFCR8_0),.din(w_dff_A_xMdH4bvC6_0),.clk(gclk));
	jdff dff_A_w14rmFCR8_0(.dout(w_dff_A_YIe0BZdp2_0),.din(w_dff_A_w14rmFCR8_0),.clk(gclk));
	jdff dff_A_YIe0BZdp2_0(.dout(G376),.din(w_dff_A_YIe0BZdp2_0),.clk(gclk));
	jdff dff_A_1iQksQaM0_2(.dout(w_dff_A_hJfgijJH7_0),.din(w_dff_A_1iQksQaM0_2),.clk(gclk));
	jdff dff_A_hJfgijJH7_0(.dout(w_dff_A_ENMl7Ul43_0),.din(w_dff_A_hJfgijJH7_0),.clk(gclk));
	jdff dff_A_ENMl7Ul43_0(.dout(w_dff_A_DExDC5NA7_0),.din(w_dff_A_ENMl7Ul43_0),.clk(gclk));
	jdff dff_A_DExDC5NA7_0(.dout(w_dff_A_lvtQbmGm9_0),.din(w_dff_A_DExDC5NA7_0),.clk(gclk));
	jdff dff_A_lvtQbmGm9_0(.dout(w_dff_A_Dn1W2jZo5_0),.din(w_dff_A_lvtQbmGm9_0),.clk(gclk));
	jdff dff_A_Dn1W2jZo5_0(.dout(w_dff_A_oRVU4bwl0_0),.din(w_dff_A_Dn1W2jZo5_0),.clk(gclk));
	jdff dff_A_oRVU4bwl0_0(.dout(w_dff_A_3EwZXQr04_0),.din(w_dff_A_oRVU4bwl0_0),.clk(gclk));
	jdff dff_A_3EwZXQr04_0(.dout(w_dff_A_AdfZZQkV9_0),.din(w_dff_A_3EwZXQr04_0),.clk(gclk));
	jdff dff_A_AdfZZQkV9_0(.dout(w_dff_A_cPHzPg2Q5_0),.din(w_dff_A_AdfZZQkV9_0),.clk(gclk));
	jdff dff_A_cPHzPg2Q5_0(.dout(w_dff_A_Utf0xcYh7_0),.din(w_dff_A_cPHzPg2Q5_0),.clk(gclk));
	jdff dff_A_Utf0xcYh7_0(.dout(w_dff_A_g5xImQhC7_0),.din(w_dff_A_Utf0xcYh7_0),.clk(gclk));
	jdff dff_A_g5xImQhC7_0(.dout(w_dff_A_ASQRqqgS8_0),.din(w_dff_A_g5xImQhC7_0),.clk(gclk));
	jdff dff_A_ASQRqqgS8_0(.dout(w_dff_A_npwC4EFi4_0),.din(w_dff_A_ASQRqqgS8_0),.clk(gclk));
	jdff dff_A_npwC4EFi4_0(.dout(w_dff_A_TttgXi3p2_0),.din(w_dff_A_npwC4EFi4_0),.clk(gclk));
	jdff dff_A_TttgXi3p2_0(.dout(w_dff_A_xz1zoii98_0),.din(w_dff_A_TttgXi3p2_0),.clk(gclk));
	jdff dff_A_xz1zoii98_0(.dout(w_dff_A_QZu0Vnbb5_0),.din(w_dff_A_xz1zoii98_0),.clk(gclk));
	jdff dff_A_QZu0Vnbb5_0(.dout(w_dff_A_cuTUdWVQ7_0),.din(w_dff_A_QZu0Vnbb5_0),.clk(gclk));
	jdff dff_A_cuTUdWVQ7_0(.dout(w_dff_A_DmhPxgal5_0),.din(w_dff_A_cuTUdWVQ7_0),.clk(gclk));
	jdff dff_A_DmhPxgal5_0(.dout(w_dff_A_TU3bReNd5_0),.din(w_dff_A_DmhPxgal5_0),.clk(gclk));
	jdff dff_A_TU3bReNd5_0(.dout(w_dff_A_CtZh37QI7_0),.din(w_dff_A_TU3bReNd5_0),.clk(gclk));
	jdff dff_A_CtZh37QI7_0(.dout(w_dff_A_Pvsn6F9o5_0),.din(w_dff_A_CtZh37QI7_0),.clk(gclk));
	jdff dff_A_Pvsn6F9o5_0(.dout(G379),.din(w_dff_A_Pvsn6F9o5_0),.clk(gclk));
	jdff dff_A_8hS9m2Y73_2(.dout(w_dff_A_81labtvY2_0),.din(w_dff_A_8hS9m2Y73_2),.clk(gclk));
	jdff dff_A_81labtvY2_0(.dout(w_dff_A_akV4xtHz7_0),.din(w_dff_A_81labtvY2_0),.clk(gclk));
	jdff dff_A_akV4xtHz7_0(.dout(w_dff_A_nIGbZKFp1_0),.din(w_dff_A_akV4xtHz7_0),.clk(gclk));
	jdff dff_A_nIGbZKFp1_0(.dout(w_dff_A_lUNlwOxw3_0),.din(w_dff_A_nIGbZKFp1_0),.clk(gclk));
	jdff dff_A_lUNlwOxw3_0(.dout(w_dff_A_gSSZ0jMX7_0),.din(w_dff_A_lUNlwOxw3_0),.clk(gclk));
	jdff dff_A_gSSZ0jMX7_0(.dout(w_dff_A_rcRwI3k86_0),.din(w_dff_A_gSSZ0jMX7_0),.clk(gclk));
	jdff dff_A_rcRwI3k86_0(.dout(w_dff_A_4noCiurx9_0),.din(w_dff_A_rcRwI3k86_0),.clk(gclk));
	jdff dff_A_4noCiurx9_0(.dout(w_dff_A_k94ta9Te0_0),.din(w_dff_A_4noCiurx9_0),.clk(gclk));
	jdff dff_A_k94ta9Te0_0(.dout(w_dff_A_9ipDSy589_0),.din(w_dff_A_k94ta9Te0_0),.clk(gclk));
	jdff dff_A_9ipDSy589_0(.dout(w_dff_A_uEyHgZvI9_0),.din(w_dff_A_9ipDSy589_0),.clk(gclk));
	jdff dff_A_uEyHgZvI9_0(.dout(w_dff_A_PSRTnObD1_0),.din(w_dff_A_uEyHgZvI9_0),.clk(gclk));
	jdff dff_A_PSRTnObD1_0(.dout(w_dff_A_mvSPDdfY6_0),.din(w_dff_A_PSRTnObD1_0),.clk(gclk));
	jdff dff_A_mvSPDdfY6_0(.dout(w_dff_A_QN6sim7e1_0),.din(w_dff_A_mvSPDdfY6_0),.clk(gclk));
	jdff dff_A_QN6sim7e1_0(.dout(w_dff_A_JP63ReqE8_0),.din(w_dff_A_QN6sim7e1_0),.clk(gclk));
	jdff dff_A_JP63ReqE8_0(.dout(w_dff_A_y2sS8QCS1_0),.din(w_dff_A_JP63ReqE8_0),.clk(gclk));
	jdff dff_A_y2sS8QCS1_0(.dout(w_dff_A_a5EPy4Eo6_0),.din(w_dff_A_y2sS8QCS1_0),.clk(gclk));
	jdff dff_A_a5EPy4Eo6_0(.dout(w_dff_A_5o1x4bdg3_0),.din(w_dff_A_a5EPy4Eo6_0),.clk(gclk));
	jdff dff_A_5o1x4bdg3_0(.dout(w_dff_A_3ICkKOD14_0),.din(w_dff_A_5o1x4bdg3_0),.clk(gclk));
	jdff dff_A_3ICkKOD14_0(.dout(w_dff_A_C1hkKMUJ3_0),.din(w_dff_A_3ICkKOD14_0),.clk(gclk));
	jdff dff_A_C1hkKMUJ3_0(.dout(w_dff_A_JZvHAGLw5_0),.din(w_dff_A_C1hkKMUJ3_0),.clk(gclk));
	jdff dff_A_JZvHAGLw5_0(.dout(w_dff_A_fyaugnMa2_0),.din(w_dff_A_JZvHAGLw5_0),.clk(gclk));
	jdff dff_A_fyaugnMa2_0(.dout(G382),.din(w_dff_A_fyaugnMa2_0),.clk(gclk));
	jdff dff_A_QdpmjzBx0_2(.dout(w_dff_A_iZEIChW01_0),.din(w_dff_A_QdpmjzBx0_2),.clk(gclk));
	jdff dff_A_iZEIChW01_0(.dout(w_dff_A_mn0c5MFP5_0),.din(w_dff_A_iZEIChW01_0),.clk(gclk));
	jdff dff_A_mn0c5MFP5_0(.dout(w_dff_A_Dj3tBW0L8_0),.din(w_dff_A_mn0c5MFP5_0),.clk(gclk));
	jdff dff_A_Dj3tBW0L8_0(.dout(w_dff_A_7kaOGsd84_0),.din(w_dff_A_Dj3tBW0L8_0),.clk(gclk));
	jdff dff_A_7kaOGsd84_0(.dout(w_dff_A_0cWbSjBm6_0),.din(w_dff_A_7kaOGsd84_0),.clk(gclk));
	jdff dff_A_0cWbSjBm6_0(.dout(w_dff_A_MIY5zbxi1_0),.din(w_dff_A_0cWbSjBm6_0),.clk(gclk));
	jdff dff_A_MIY5zbxi1_0(.dout(w_dff_A_wTQvmoWW0_0),.din(w_dff_A_MIY5zbxi1_0),.clk(gclk));
	jdff dff_A_wTQvmoWW0_0(.dout(w_dff_A_GAteg4uW2_0),.din(w_dff_A_wTQvmoWW0_0),.clk(gclk));
	jdff dff_A_GAteg4uW2_0(.dout(w_dff_A_xVQkVIfh8_0),.din(w_dff_A_GAteg4uW2_0),.clk(gclk));
	jdff dff_A_xVQkVIfh8_0(.dout(w_dff_A_HGnJh86x2_0),.din(w_dff_A_xVQkVIfh8_0),.clk(gclk));
	jdff dff_A_HGnJh86x2_0(.dout(w_dff_A_OJvHaqSg2_0),.din(w_dff_A_HGnJh86x2_0),.clk(gclk));
	jdff dff_A_OJvHaqSg2_0(.dout(w_dff_A_vxK1JuXe5_0),.din(w_dff_A_OJvHaqSg2_0),.clk(gclk));
	jdff dff_A_vxK1JuXe5_0(.dout(w_dff_A_lI7zYVwi0_0),.din(w_dff_A_vxK1JuXe5_0),.clk(gclk));
	jdff dff_A_lI7zYVwi0_0(.dout(w_dff_A_qgijVHmm8_0),.din(w_dff_A_lI7zYVwi0_0),.clk(gclk));
	jdff dff_A_qgijVHmm8_0(.dout(w_dff_A_bQjDTPrO9_0),.din(w_dff_A_qgijVHmm8_0),.clk(gclk));
	jdff dff_A_bQjDTPrO9_0(.dout(w_dff_A_vHHhn0rE8_0),.din(w_dff_A_bQjDTPrO9_0),.clk(gclk));
	jdff dff_A_vHHhn0rE8_0(.dout(w_dff_A_moKsCxe35_0),.din(w_dff_A_vHHhn0rE8_0),.clk(gclk));
	jdff dff_A_moKsCxe35_0(.dout(w_dff_A_fbVCFjhV8_0),.din(w_dff_A_moKsCxe35_0),.clk(gclk));
	jdff dff_A_fbVCFjhV8_0(.dout(w_dff_A_yxYhDQmB1_0),.din(w_dff_A_fbVCFjhV8_0),.clk(gclk));
	jdff dff_A_yxYhDQmB1_0(.dout(w_dff_A_VEG1LvX42_0),.din(w_dff_A_yxYhDQmB1_0),.clk(gclk));
	jdff dff_A_VEG1LvX42_0(.dout(w_dff_A_DH8muabI7_0),.din(w_dff_A_VEG1LvX42_0),.clk(gclk));
	jdff dff_A_DH8muabI7_0(.dout(w_dff_A_lvIBfCit0_0),.din(w_dff_A_DH8muabI7_0),.clk(gclk));
	jdff dff_A_lvIBfCit0_0(.dout(w_dff_A_i6ELr4Gm8_0),.din(w_dff_A_lvIBfCit0_0),.clk(gclk));
	jdff dff_A_i6ELr4Gm8_0(.dout(G385),.din(w_dff_A_i6ELr4Gm8_0),.clk(gclk));
	jdff dff_A_bjP8Gnko9_1(.dout(w_dff_A_JygE6xV54_0),.din(w_dff_A_bjP8Gnko9_1),.clk(gclk));
	jdff dff_A_JygE6xV54_0(.dout(w_dff_A_H4LIQZcz0_0),.din(w_dff_A_JygE6xV54_0),.clk(gclk));
	jdff dff_A_H4LIQZcz0_0(.dout(w_dff_A_9BdYvwWZ5_0),.din(w_dff_A_H4LIQZcz0_0),.clk(gclk));
	jdff dff_A_9BdYvwWZ5_0(.dout(w_dff_A_xjFsUMIC1_0),.din(w_dff_A_9BdYvwWZ5_0),.clk(gclk));
	jdff dff_A_xjFsUMIC1_0(.dout(w_dff_A_nBEVTmQl0_0),.din(w_dff_A_xjFsUMIC1_0),.clk(gclk));
	jdff dff_A_nBEVTmQl0_0(.dout(w_dff_A_ZTRW8m1r2_0),.din(w_dff_A_nBEVTmQl0_0),.clk(gclk));
	jdff dff_A_ZTRW8m1r2_0(.dout(w_dff_A_vY0xZFyl9_0),.din(w_dff_A_ZTRW8m1r2_0),.clk(gclk));
	jdff dff_A_vY0xZFyl9_0(.dout(w_dff_A_Mt9v6H714_0),.din(w_dff_A_vY0xZFyl9_0),.clk(gclk));
	jdff dff_A_Mt9v6H714_0(.dout(w_dff_A_0YXCL5Ik2_0),.din(w_dff_A_Mt9v6H714_0),.clk(gclk));
	jdff dff_A_0YXCL5Ik2_0(.dout(w_dff_A_CBiBBm4n5_0),.din(w_dff_A_0YXCL5Ik2_0),.clk(gclk));
	jdff dff_A_CBiBBm4n5_0(.dout(w_dff_A_iBsDKZqG6_0),.din(w_dff_A_CBiBBm4n5_0),.clk(gclk));
	jdff dff_A_iBsDKZqG6_0(.dout(w_dff_A_7WFgkYER7_0),.din(w_dff_A_iBsDKZqG6_0),.clk(gclk));
	jdff dff_A_7WFgkYER7_0(.dout(w_dff_A_FsukPbtM5_0),.din(w_dff_A_7WFgkYER7_0),.clk(gclk));
	jdff dff_A_FsukPbtM5_0(.dout(w_dff_A_GugBEpix2_0),.din(w_dff_A_FsukPbtM5_0),.clk(gclk));
	jdff dff_A_GugBEpix2_0(.dout(w_dff_A_V0skxr0F7_0),.din(w_dff_A_GugBEpix2_0),.clk(gclk));
	jdff dff_A_V0skxr0F7_0(.dout(w_dff_A_XfMIXKrl8_0),.din(w_dff_A_V0skxr0F7_0),.clk(gclk));
	jdff dff_A_XfMIXKrl8_0(.dout(w_dff_A_Ll27CUwy3_0),.din(w_dff_A_XfMIXKrl8_0),.clk(gclk));
	jdff dff_A_Ll27CUwy3_0(.dout(w_dff_A_NzGWomL06_0),.din(w_dff_A_Ll27CUwy3_0),.clk(gclk));
	jdff dff_A_NzGWomL06_0(.dout(w_dff_A_UUfhRLOj5_0),.din(w_dff_A_NzGWomL06_0),.clk(gclk));
	jdff dff_A_UUfhRLOj5_0(.dout(w_dff_A_o6KxQzLL7_0),.din(w_dff_A_UUfhRLOj5_0),.clk(gclk));
	jdff dff_A_o6KxQzLL7_0(.dout(w_dff_A_GfGoUerw9_0),.din(w_dff_A_o6KxQzLL7_0),.clk(gclk));
	jdff dff_A_GfGoUerw9_0(.dout(w_dff_A_r2wZF0K61_0),.din(w_dff_A_GfGoUerw9_0),.clk(gclk));
	jdff dff_A_r2wZF0K61_0(.dout(w_dff_A_H9WEcLuX7_0),.din(w_dff_A_r2wZF0K61_0),.clk(gclk));
	jdff dff_A_H9WEcLuX7_0(.dout(w_dff_A_cplgJl6L5_0),.din(w_dff_A_H9WEcLuX7_0),.clk(gclk));
	jdff dff_A_cplgJl6L5_0(.dout(w_dff_A_kgzbzXtT2_0),.din(w_dff_A_cplgJl6L5_0),.clk(gclk));
	jdff dff_A_kgzbzXtT2_0(.dout(w_dff_A_KY6aIAwW6_0),.din(w_dff_A_kgzbzXtT2_0),.clk(gclk));
	jdff dff_A_KY6aIAwW6_0(.dout(w_dff_A_vfpGiafr1_0),.din(w_dff_A_KY6aIAwW6_0),.clk(gclk));
	jdff dff_A_vfpGiafr1_0(.dout(G412),.din(w_dff_A_vfpGiafr1_0),.clk(gclk));
	jdff dff_A_I8w0B8AP8_1(.dout(w_dff_A_lvMnoDQb4_0),.din(w_dff_A_I8w0B8AP8_1),.clk(gclk));
	jdff dff_A_lvMnoDQb4_0(.dout(w_dff_A_quCktKZK7_0),.din(w_dff_A_lvMnoDQb4_0),.clk(gclk));
	jdff dff_A_quCktKZK7_0(.dout(w_dff_A_X2cIBIdp3_0),.din(w_dff_A_quCktKZK7_0),.clk(gclk));
	jdff dff_A_X2cIBIdp3_0(.dout(w_dff_A_t4blgWWg3_0),.din(w_dff_A_X2cIBIdp3_0),.clk(gclk));
	jdff dff_A_t4blgWWg3_0(.dout(w_dff_A_Of6vaUcI3_0),.din(w_dff_A_t4blgWWg3_0),.clk(gclk));
	jdff dff_A_Of6vaUcI3_0(.dout(w_dff_A_WCLfFFzk4_0),.din(w_dff_A_Of6vaUcI3_0),.clk(gclk));
	jdff dff_A_WCLfFFzk4_0(.dout(w_dff_A_hEk6ocyy6_0),.din(w_dff_A_WCLfFFzk4_0),.clk(gclk));
	jdff dff_A_hEk6ocyy6_0(.dout(w_dff_A_WBawVD2a9_0),.din(w_dff_A_hEk6ocyy6_0),.clk(gclk));
	jdff dff_A_WBawVD2a9_0(.dout(w_dff_A_VycTajte5_0),.din(w_dff_A_WBawVD2a9_0),.clk(gclk));
	jdff dff_A_VycTajte5_0(.dout(w_dff_A_YhKGf7wL9_0),.din(w_dff_A_VycTajte5_0),.clk(gclk));
	jdff dff_A_YhKGf7wL9_0(.dout(w_dff_A_Kz6Ru4PS6_0),.din(w_dff_A_YhKGf7wL9_0),.clk(gclk));
	jdff dff_A_Kz6Ru4PS6_0(.dout(w_dff_A_L0UlO98V6_0),.din(w_dff_A_Kz6Ru4PS6_0),.clk(gclk));
	jdff dff_A_L0UlO98V6_0(.dout(w_dff_A_gR1jdJvZ9_0),.din(w_dff_A_L0UlO98V6_0),.clk(gclk));
	jdff dff_A_gR1jdJvZ9_0(.dout(w_dff_A_nExZUtR06_0),.din(w_dff_A_gR1jdJvZ9_0),.clk(gclk));
	jdff dff_A_nExZUtR06_0(.dout(w_dff_A_5BU2K0yv5_0),.din(w_dff_A_nExZUtR06_0),.clk(gclk));
	jdff dff_A_5BU2K0yv5_0(.dout(w_dff_A_hT4K5FmC9_0),.din(w_dff_A_5BU2K0yv5_0),.clk(gclk));
	jdff dff_A_hT4K5FmC9_0(.dout(w_dff_A_5LoUhNRd9_0),.din(w_dff_A_hT4K5FmC9_0),.clk(gclk));
	jdff dff_A_5LoUhNRd9_0(.dout(w_dff_A_h0ewkhsh3_0),.din(w_dff_A_5LoUhNRd9_0),.clk(gclk));
	jdff dff_A_h0ewkhsh3_0(.dout(w_dff_A_btY6XhyT9_0),.din(w_dff_A_h0ewkhsh3_0),.clk(gclk));
	jdff dff_A_btY6XhyT9_0(.dout(w_dff_A_A5zHOWMX2_0),.din(w_dff_A_btY6XhyT9_0),.clk(gclk));
	jdff dff_A_A5zHOWMX2_0(.dout(w_dff_A_E7nqzzLD2_0),.din(w_dff_A_A5zHOWMX2_0),.clk(gclk));
	jdff dff_A_E7nqzzLD2_0(.dout(w_dff_A_aYNRGjsY9_0),.din(w_dff_A_E7nqzzLD2_0),.clk(gclk));
	jdff dff_A_aYNRGjsY9_0(.dout(w_dff_A_2uwE9oa72_0),.din(w_dff_A_aYNRGjsY9_0),.clk(gclk));
	jdff dff_A_2uwE9oa72_0(.dout(w_dff_A_52KrNaZP3_0),.din(w_dff_A_2uwE9oa72_0),.clk(gclk));
	jdff dff_A_52KrNaZP3_0(.dout(w_dff_A_Udi0OLKP8_0),.din(w_dff_A_52KrNaZP3_0),.clk(gclk));
	jdff dff_A_Udi0OLKP8_0(.dout(w_dff_A_pC563uJb1_0),.din(w_dff_A_Udi0OLKP8_0),.clk(gclk));
	jdff dff_A_pC563uJb1_0(.dout(w_dff_A_3jAjF1Gz6_0),.din(w_dff_A_pC563uJb1_0),.clk(gclk));
	jdff dff_A_3jAjF1Gz6_0(.dout(w_dff_A_wwd0LvTI7_0),.din(w_dff_A_3jAjF1Gz6_0),.clk(gclk));
	jdff dff_A_wwd0LvTI7_0(.dout(w_dff_A_fl9wfYSL3_0),.din(w_dff_A_wwd0LvTI7_0),.clk(gclk));
	jdff dff_A_fl9wfYSL3_0(.dout(G414),.din(w_dff_A_fl9wfYSL3_0),.clk(gclk));
	jdff dff_A_qkkR41lL2_1(.dout(w_dff_A_7ljZlT9V9_0),.din(w_dff_A_qkkR41lL2_1),.clk(gclk));
	jdff dff_A_7ljZlT9V9_0(.dout(w_dff_A_shnOCCR11_0),.din(w_dff_A_7ljZlT9V9_0),.clk(gclk));
	jdff dff_A_shnOCCR11_0(.dout(w_dff_A_czG8FT767_0),.din(w_dff_A_shnOCCR11_0),.clk(gclk));
	jdff dff_A_czG8FT767_0(.dout(w_dff_A_al6xBKIX6_0),.din(w_dff_A_czG8FT767_0),.clk(gclk));
	jdff dff_A_al6xBKIX6_0(.dout(w_dff_A_R7QPpjgf2_0),.din(w_dff_A_al6xBKIX6_0),.clk(gclk));
	jdff dff_A_R7QPpjgf2_0(.dout(w_dff_A_pPRppIca7_0),.din(w_dff_A_R7QPpjgf2_0),.clk(gclk));
	jdff dff_A_pPRppIca7_0(.dout(w_dff_A_zO4s8VNy2_0),.din(w_dff_A_pPRppIca7_0),.clk(gclk));
	jdff dff_A_zO4s8VNy2_0(.dout(w_dff_A_NTX6bz143_0),.din(w_dff_A_zO4s8VNy2_0),.clk(gclk));
	jdff dff_A_NTX6bz143_0(.dout(w_dff_A_GhGmbBTX1_0),.din(w_dff_A_NTX6bz143_0),.clk(gclk));
	jdff dff_A_GhGmbBTX1_0(.dout(w_dff_A_uhyNS0uH7_0),.din(w_dff_A_GhGmbBTX1_0),.clk(gclk));
	jdff dff_A_uhyNS0uH7_0(.dout(w_dff_A_MKOz98611_0),.din(w_dff_A_uhyNS0uH7_0),.clk(gclk));
	jdff dff_A_MKOz98611_0(.dout(w_dff_A_2LBlAj0V3_0),.din(w_dff_A_MKOz98611_0),.clk(gclk));
	jdff dff_A_2LBlAj0V3_0(.dout(w_dff_A_S74WIrSZ4_0),.din(w_dff_A_2LBlAj0V3_0),.clk(gclk));
	jdff dff_A_S74WIrSZ4_0(.dout(w_dff_A_qBBnIvzr8_0),.din(w_dff_A_S74WIrSZ4_0),.clk(gclk));
	jdff dff_A_qBBnIvzr8_0(.dout(w_dff_A_6AmY8qAZ4_0),.din(w_dff_A_qBBnIvzr8_0),.clk(gclk));
	jdff dff_A_6AmY8qAZ4_0(.dout(w_dff_A_Sr5tra2P7_0),.din(w_dff_A_6AmY8qAZ4_0),.clk(gclk));
	jdff dff_A_Sr5tra2P7_0(.dout(w_dff_A_slxDaHWE6_0),.din(w_dff_A_Sr5tra2P7_0),.clk(gclk));
	jdff dff_A_slxDaHWE6_0(.dout(w_dff_A_386anNwP6_0),.din(w_dff_A_slxDaHWE6_0),.clk(gclk));
	jdff dff_A_386anNwP6_0(.dout(w_dff_A_u4bbuj2R2_0),.din(w_dff_A_386anNwP6_0),.clk(gclk));
	jdff dff_A_u4bbuj2R2_0(.dout(w_dff_A_BG3MG6e71_0),.din(w_dff_A_u4bbuj2R2_0),.clk(gclk));
	jdff dff_A_BG3MG6e71_0(.dout(w_dff_A_XtDUCDlA7_0),.din(w_dff_A_BG3MG6e71_0),.clk(gclk));
	jdff dff_A_XtDUCDlA7_0(.dout(w_dff_A_1P1c9G1b8_0),.din(w_dff_A_XtDUCDlA7_0),.clk(gclk));
	jdff dff_A_1P1c9G1b8_0(.dout(w_dff_A_M23WeA3w0_0),.din(w_dff_A_1P1c9G1b8_0),.clk(gclk));
	jdff dff_A_M23WeA3w0_0(.dout(w_dff_A_y5ZnVpJd4_0),.din(w_dff_A_M23WeA3w0_0),.clk(gclk));
	jdff dff_A_y5ZnVpJd4_0(.dout(w_dff_A_kBitKUpS4_0),.din(w_dff_A_y5ZnVpJd4_0),.clk(gclk));
	jdff dff_A_kBitKUpS4_0(.dout(w_dff_A_mG0QgLiw8_0),.din(w_dff_A_kBitKUpS4_0),.clk(gclk));
	jdff dff_A_mG0QgLiw8_0(.dout(w_dff_A_IMH9stej5_0),.din(w_dff_A_mG0QgLiw8_0),.clk(gclk));
	jdff dff_A_IMH9stej5_0(.dout(w_dff_A_ku4bgICf8_0),.din(w_dff_A_IMH9stej5_0),.clk(gclk));
	jdff dff_A_ku4bgICf8_0(.dout(G416),.din(w_dff_A_ku4bgICf8_0),.clk(gclk));
	jdff dff_A_ILSvZBEJ4_2(.dout(w_dff_A_OVLSzOC91_0),.din(w_dff_A_ILSvZBEJ4_2),.clk(gclk));
	jdff dff_A_OVLSzOC91_0(.dout(w_dff_A_ZyDKHbNT6_0),.din(w_dff_A_OVLSzOC91_0),.clk(gclk));
	jdff dff_A_ZyDKHbNT6_0(.dout(w_dff_A_01A7bkPs6_0),.din(w_dff_A_ZyDKHbNT6_0),.clk(gclk));
	jdff dff_A_01A7bkPs6_0(.dout(w_dff_A_SdsYbdir9_0),.din(w_dff_A_01A7bkPs6_0),.clk(gclk));
	jdff dff_A_SdsYbdir9_0(.dout(w_dff_A_yUIXDO435_0),.din(w_dff_A_SdsYbdir9_0),.clk(gclk));
	jdff dff_A_yUIXDO435_0(.dout(w_dff_A_SFTo6Cfo7_0),.din(w_dff_A_yUIXDO435_0),.clk(gclk));
	jdff dff_A_SFTo6Cfo7_0(.dout(w_dff_A_QK4jZoz99_0),.din(w_dff_A_SFTo6Cfo7_0),.clk(gclk));
	jdff dff_A_QK4jZoz99_0(.dout(w_dff_A_2krjyInS3_0),.din(w_dff_A_QK4jZoz99_0),.clk(gclk));
	jdff dff_A_2krjyInS3_0(.dout(w_dff_A_P125zpNw4_0),.din(w_dff_A_2krjyInS3_0),.clk(gclk));
	jdff dff_A_P125zpNw4_0(.dout(w_dff_A_ediNWG1J7_0),.din(w_dff_A_P125zpNw4_0),.clk(gclk));
	jdff dff_A_ediNWG1J7_0(.dout(G249),.din(w_dff_A_ediNWG1J7_0),.clk(gclk));
	jdff dff_A_xfiKRwPP3_2(.dout(w_dff_A_aK0GLROY2_0),.din(w_dff_A_xfiKRwPP3_2),.clk(gclk));
	jdff dff_A_aK0GLROY2_0(.dout(w_dff_A_36wbyAAn1_0),.din(w_dff_A_aK0GLROY2_0),.clk(gclk));
	jdff dff_A_36wbyAAn1_0(.dout(w_dff_A_i6rV34jg1_0),.din(w_dff_A_36wbyAAn1_0),.clk(gclk));
	jdff dff_A_i6rV34jg1_0(.dout(w_dff_A_vfccntIk7_0),.din(w_dff_A_i6rV34jg1_0),.clk(gclk));
	jdff dff_A_vfccntIk7_0(.dout(w_dff_A_NZNHqxuW7_0),.din(w_dff_A_vfccntIk7_0),.clk(gclk));
	jdff dff_A_NZNHqxuW7_0(.dout(w_dff_A_fycggT6y2_0),.din(w_dff_A_NZNHqxuW7_0),.clk(gclk));
	jdff dff_A_fycggT6y2_0(.dout(w_dff_A_4o1FDuoc5_0),.din(w_dff_A_fycggT6y2_0),.clk(gclk));
	jdff dff_A_4o1FDuoc5_0(.dout(w_dff_A_FjvKrP1L7_0),.din(w_dff_A_4o1FDuoc5_0),.clk(gclk));
	jdff dff_A_FjvKrP1L7_0(.dout(w_dff_A_led1xBmg1_0),.din(w_dff_A_FjvKrP1L7_0),.clk(gclk));
	jdff dff_A_led1xBmg1_0(.dout(w_dff_A_X39QseWh6_0),.din(w_dff_A_led1xBmg1_0),.clk(gclk));
	jdff dff_A_X39QseWh6_0(.dout(G295),.din(w_dff_A_X39QseWh6_0),.clk(gclk));
	jdff dff_A_zrcXL1rl7_2(.dout(w_dff_A_V6rEcdFt9_0),.din(w_dff_A_zrcXL1rl7_2),.clk(gclk));
	jdff dff_A_V6rEcdFt9_0(.dout(w_dff_A_YVfZ5NnC0_0),.din(w_dff_A_V6rEcdFt9_0),.clk(gclk));
	jdff dff_A_YVfZ5NnC0_0(.dout(w_dff_A_742KAgvO1_0),.din(w_dff_A_YVfZ5NnC0_0),.clk(gclk));
	jdff dff_A_742KAgvO1_0(.dout(G324),.din(w_dff_A_742KAgvO1_0),.clk(gclk));
	jdff dff_A_qDtSjULd9_1(.dout(w_dff_A_ugdaHuIq3_0),.din(w_dff_A_qDtSjULd9_1),.clk(gclk));
	jdff dff_A_ugdaHuIq3_0(.dout(w_dff_A_KsYWvMPz2_0),.din(w_dff_A_ugdaHuIq3_0),.clk(gclk));
	jdff dff_A_KsYWvMPz2_0(.dout(w_dff_A_pzKquxwd5_0),.din(w_dff_A_KsYWvMPz2_0),.clk(gclk));
	jdff dff_A_pzKquxwd5_0(.dout(w_dff_A_xPDRx4bs8_0),.din(w_dff_A_pzKquxwd5_0),.clk(gclk));
	jdff dff_A_xPDRx4bs8_0(.dout(w_dff_A_1XTG5deb9_0),.din(w_dff_A_xPDRx4bs8_0),.clk(gclk));
	jdff dff_A_1XTG5deb9_0(.dout(w_dff_A_uDtlWOCu5_0),.din(w_dff_A_1XTG5deb9_0),.clk(gclk));
	jdff dff_A_uDtlWOCu5_0(.dout(w_dff_A_VLrYmf5Z1_0),.din(w_dff_A_uDtlWOCu5_0),.clk(gclk));
	jdff dff_A_VLrYmf5Z1_0(.dout(w_dff_A_spldhYxi7_0),.din(w_dff_A_VLrYmf5Z1_0),.clk(gclk));
	jdff dff_A_spldhYxi7_0(.dout(w_dff_A_KhQG3VGM0_0),.din(w_dff_A_spldhYxi7_0),.clk(gclk));
	jdff dff_A_KhQG3VGM0_0(.dout(w_dff_A_n5Qvx2W22_0),.din(w_dff_A_KhQG3VGM0_0),.clk(gclk));
	jdff dff_A_n5Qvx2W22_0(.dout(w_dff_A_8S4rUr0x5_0),.din(w_dff_A_n5Qvx2W22_0),.clk(gclk));
	jdff dff_A_8S4rUr0x5_0(.dout(w_dff_A_PYLW6zl73_0),.din(w_dff_A_8S4rUr0x5_0),.clk(gclk));
	jdff dff_A_PYLW6zl73_0(.dout(w_dff_A_mGLUpW3V3_0),.din(w_dff_A_PYLW6zl73_0),.clk(gclk));
	jdff dff_A_mGLUpW3V3_0(.dout(w_dff_A_FIEAXlDu9_0),.din(w_dff_A_mGLUpW3V3_0),.clk(gclk));
	jdff dff_A_FIEAXlDu9_0(.dout(w_dff_A_1tJXCDZH5_0),.din(w_dff_A_FIEAXlDu9_0),.clk(gclk));
	jdff dff_A_1tJXCDZH5_0(.dout(w_dff_A_l5gMOBei4_0),.din(w_dff_A_1tJXCDZH5_0),.clk(gclk));
	jdff dff_A_l5gMOBei4_0(.dout(w_dff_A_8qXkLzQl9_0),.din(w_dff_A_l5gMOBei4_0),.clk(gclk));
	jdff dff_A_8qXkLzQl9_0(.dout(w_dff_A_5sNSkv1N1_0),.din(w_dff_A_8qXkLzQl9_0),.clk(gclk));
	jdff dff_A_5sNSkv1N1_0(.dout(w_dff_A_ASJ4J5SQ2_0),.din(w_dff_A_5sNSkv1N1_0),.clk(gclk));
	jdff dff_A_ASJ4J5SQ2_0(.dout(w_dff_A_w4VHtvYt5_0),.din(w_dff_A_ASJ4J5SQ2_0),.clk(gclk));
	jdff dff_A_w4VHtvYt5_0(.dout(G252),.din(w_dff_A_w4VHtvYt5_0),.clk(gclk));
	jdff dff_A_gwDlvvGS8_2(.dout(w_dff_A_pyMSuIju5_0),.din(w_dff_A_gwDlvvGS8_2),.clk(gclk));
	jdff dff_A_pyMSuIju5_0(.dout(w_dff_A_HvPMqq5t9_0),.din(w_dff_A_pyMSuIju5_0),.clk(gclk));
	jdff dff_A_HvPMqq5t9_0(.dout(w_dff_A_UGyAlJ6Y0_0),.din(w_dff_A_HvPMqq5t9_0),.clk(gclk));
	jdff dff_A_UGyAlJ6Y0_0(.dout(w_dff_A_XSrtizU08_0),.din(w_dff_A_UGyAlJ6Y0_0),.clk(gclk));
	jdff dff_A_XSrtizU08_0(.dout(w_dff_A_8lN7DabA1_0),.din(w_dff_A_XSrtizU08_0),.clk(gclk));
	jdff dff_A_8lN7DabA1_0(.dout(G310),.din(w_dff_A_8lN7DabA1_0),.clk(gclk));
	jdff dff_A_HM3MKpQL8_2(.dout(w_dff_A_R6jWaAUu3_0),.din(w_dff_A_HM3MKpQL8_2),.clk(gclk));
	jdff dff_A_R6jWaAUu3_0(.dout(w_dff_A_MBiSDkNg6_0),.din(w_dff_A_R6jWaAUu3_0),.clk(gclk));
	jdff dff_A_MBiSDkNg6_0(.dout(w_dff_A_TiLs4IDp0_0),.din(w_dff_A_MBiSDkNg6_0),.clk(gclk));
	jdff dff_A_TiLs4IDp0_0(.dout(w_dff_A_f2y4bC435_0),.din(w_dff_A_TiLs4IDp0_0),.clk(gclk));
	jdff dff_A_f2y4bC435_0(.dout(G313),.din(w_dff_A_f2y4bC435_0),.clk(gclk));
	jdff dff_A_90iJhh3S3_2(.dout(w_dff_A_wMVTovFG7_0),.din(w_dff_A_90iJhh3S3_2),.clk(gclk));
	jdff dff_A_wMVTovFG7_0(.dout(w_dff_A_sNDuGX0S8_0),.din(w_dff_A_wMVTovFG7_0),.clk(gclk));
	jdff dff_A_sNDuGX0S8_0(.dout(w_dff_A_cNEKW8gF0_0),.din(w_dff_A_sNDuGX0S8_0),.clk(gclk));
	jdff dff_A_cNEKW8gF0_0(.dout(w_dff_A_uimQMgSQ5_0),.din(w_dff_A_cNEKW8gF0_0),.clk(gclk));
	jdff dff_A_uimQMgSQ5_0(.dout(w_dff_A_QhnLDcRO1_0),.din(w_dff_A_uimQMgSQ5_0),.clk(gclk));
	jdff dff_A_QhnLDcRO1_0(.dout(w_dff_A_QndRye4D9_0),.din(w_dff_A_QhnLDcRO1_0),.clk(gclk));
	jdff dff_A_QndRye4D9_0(.dout(w_dff_A_Qp3H3yc01_0),.din(w_dff_A_QndRye4D9_0),.clk(gclk));
	jdff dff_A_Qp3H3yc01_0(.dout(w_dff_A_eTQMF5Qy7_0),.din(w_dff_A_Qp3H3yc01_0),.clk(gclk));
	jdff dff_A_eTQMF5Qy7_0(.dout(G316),.din(w_dff_A_eTQMF5Qy7_0),.clk(gclk));
	jdff dff_A_3fDqDu737_2(.dout(w_dff_A_7KFerPuq5_0),.din(w_dff_A_3fDqDu737_2),.clk(gclk));
	jdff dff_A_7KFerPuq5_0(.dout(w_dff_A_5Zm3OgNo7_0),.din(w_dff_A_7KFerPuq5_0),.clk(gclk));
	jdff dff_A_5Zm3OgNo7_0(.dout(w_dff_A_1rPRtXIg7_0),.din(w_dff_A_5Zm3OgNo7_0),.clk(gclk));
	jdff dff_A_1rPRtXIg7_0(.dout(w_dff_A_LUjSBSBl2_0),.din(w_dff_A_1rPRtXIg7_0),.clk(gclk));
	jdff dff_A_LUjSBSBl2_0(.dout(w_dff_A_xgQlfr3r4_0),.din(w_dff_A_LUjSBSBl2_0),.clk(gclk));
	jdff dff_A_xgQlfr3r4_0(.dout(w_dff_A_CdS7RY2u4_0),.din(w_dff_A_xgQlfr3r4_0),.clk(gclk));
	jdff dff_A_CdS7RY2u4_0(.dout(w_dff_A_q2DaGNrb1_0),.din(w_dff_A_CdS7RY2u4_0),.clk(gclk));
	jdff dff_A_q2DaGNrb1_0(.dout(w_dff_A_eOEDl1WL5_0),.din(w_dff_A_q2DaGNrb1_0),.clk(gclk));
	jdff dff_A_eOEDl1WL5_0(.dout(G319),.din(w_dff_A_eOEDl1WL5_0),.clk(gclk));
	jdff dff_A_F5JBNVEW3_2(.dout(w_dff_A_Phw1tJnA6_0),.din(w_dff_A_F5JBNVEW3_2),.clk(gclk));
	jdff dff_A_Phw1tJnA6_0(.dout(G327),.din(w_dff_A_Phw1tJnA6_0),.clk(gclk));
	jdff dff_A_4qm3SZjK2_2(.dout(w_dff_A_WDRkfbAT3_0),.din(w_dff_A_4qm3SZjK2_2),.clk(gclk));
	jdff dff_A_WDRkfbAT3_0(.dout(G330),.din(w_dff_A_WDRkfbAT3_0),.clk(gclk));
	jdff dff_A_LuZMZecF1_2(.dout(w_dff_A_8FT8dgJl5_0),.din(w_dff_A_LuZMZecF1_2),.clk(gclk));
	jdff dff_A_8FT8dgJl5_0(.dout(G336),.din(w_dff_A_8FT8dgJl5_0),.clk(gclk));
	jdff dff_A_DpK9MJgg0_2(.dout(w_dff_A_XmzPJ8Z65_0),.din(w_dff_A_DpK9MJgg0_2),.clk(gclk));
	jdff dff_A_XmzPJ8Z65_0(.dout(w_dff_A_e8tpRDF93_0),.din(w_dff_A_XmzPJ8Z65_0),.clk(gclk));
	jdff dff_A_e8tpRDF93_0(.dout(w_dff_A_4bsi1gVk1_0),.din(w_dff_A_e8tpRDF93_0),.clk(gclk));
	jdff dff_A_4bsi1gVk1_0(.dout(w_dff_A_RwTLNT8w2_0),.din(w_dff_A_4bsi1gVk1_0),.clk(gclk));
	jdff dff_A_RwTLNT8w2_0(.dout(w_dff_A_WfdH0IHe9_0),.din(w_dff_A_RwTLNT8w2_0),.clk(gclk));
	jdff dff_A_WfdH0IHe9_0(.dout(w_dff_A_0MxlA2ET8_0),.din(w_dff_A_WfdH0IHe9_0),.clk(gclk));
	jdff dff_A_0MxlA2ET8_0(.dout(w_dff_A_fkKoHX4M6_0),.din(w_dff_A_0MxlA2ET8_0),.clk(gclk));
	jdff dff_A_fkKoHX4M6_0(.dout(w_dff_A_tVu4vRE77_0),.din(w_dff_A_fkKoHX4M6_0),.clk(gclk));
	jdff dff_A_tVu4vRE77_0(.dout(w_dff_A_sPJrOy6n7_0),.din(w_dff_A_tVu4vRE77_0),.clk(gclk));
	jdff dff_A_sPJrOy6n7_0(.dout(w_dff_A_MSlCcuJr7_0),.din(w_dff_A_sPJrOy6n7_0),.clk(gclk));
	jdff dff_A_MSlCcuJr7_0(.dout(w_dff_A_5Faf9DTs9_0),.din(w_dff_A_MSlCcuJr7_0),.clk(gclk));
	jdff dff_A_5Faf9DTs9_0(.dout(w_dff_A_ZD0wqzCR0_0),.din(w_dff_A_5Faf9DTs9_0),.clk(gclk));
	jdff dff_A_ZD0wqzCR0_0(.dout(w_dff_A_uN8TCNXs0_0),.din(w_dff_A_ZD0wqzCR0_0),.clk(gclk));
	jdff dff_A_uN8TCNXs0_0(.dout(w_dff_A_OJOU4HGP3_0),.din(w_dff_A_uN8TCNXs0_0),.clk(gclk));
	jdff dff_A_OJOU4HGP3_0(.dout(w_dff_A_vrTN3nrh9_0),.din(w_dff_A_OJOU4HGP3_0),.clk(gclk));
	jdff dff_A_vrTN3nrh9_0(.dout(w_dff_A_Yu8avxCL4_0),.din(w_dff_A_vrTN3nrh9_0),.clk(gclk));
	jdff dff_A_Yu8avxCL4_0(.dout(w_dff_A_2dEyfsHJ7_0),.din(w_dff_A_Yu8avxCL4_0),.clk(gclk));
	jdff dff_A_2dEyfsHJ7_0(.dout(w_dff_A_Ztvpptee8_0),.din(w_dff_A_2dEyfsHJ7_0),.clk(gclk));
	jdff dff_A_Ztvpptee8_0(.dout(w_dff_A_MexYlLuv6_0),.din(w_dff_A_Ztvpptee8_0),.clk(gclk));
	jdff dff_A_MexYlLuv6_0(.dout(w_dff_A_skz1TVNd4_0),.din(w_dff_A_MexYlLuv6_0),.clk(gclk));
	jdff dff_A_skz1TVNd4_0(.dout(w_dff_A_ja4VovS83_0),.din(w_dff_A_skz1TVNd4_0),.clk(gclk));
	jdff dff_A_ja4VovS83_0(.dout(w_dff_A_cO5F2zJo7_0),.din(w_dff_A_ja4VovS83_0),.clk(gclk));
	jdff dff_A_cO5F2zJo7_0(.dout(w_dff_A_EvNvKbhg4_0),.din(w_dff_A_cO5F2zJo7_0),.clk(gclk));
	jdff dff_A_EvNvKbhg4_0(.dout(w_dff_A_7S3hWtba7_0),.din(w_dff_A_EvNvKbhg4_0),.clk(gclk));
	jdff dff_A_7S3hWtba7_0(.dout(G418),.din(w_dff_A_7S3hWtba7_0),.clk(gclk));
	jdff dff_A_66Kxv2s37_2(.dout(w_dff_A_5FuhfzB66_0),.din(w_dff_A_66Kxv2s37_2),.clk(gclk));
	jdff dff_A_5FuhfzB66_0(.dout(w_dff_A_9k1mbw330_0),.din(w_dff_A_5FuhfzB66_0),.clk(gclk));
	jdff dff_A_9k1mbw330_0(.dout(w_dff_A_0o1hTSuY3_0),.din(w_dff_A_9k1mbw330_0),.clk(gclk));
	jdff dff_A_0o1hTSuY3_0(.dout(w_dff_A_u2QOunfA3_0),.din(w_dff_A_0o1hTSuY3_0),.clk(gclk));
	jdff dff_A_u2QOunfA3_0(.dout(w_dff_A_5HB4DTtw9_0),.din(w_dff_A_u2QOunfA3_0),.clk(gclk));
	jdff dff_A_5HB4DTtw9_0(.dout(G298),.din(w_dff_A_5HB4DTtw9_0),.clk(gclk));
	jdff dff_A_Zf5g3S756_2(.dout(w_dff_A_WL258vLB9_0),.din(w_dff_A_Zf5g3S756_2),.clk(gclk));
	jdff dff_A_WL258vLB9_0(.dout(w_dff_A_nyc2roSQ8_0),.din(w_dff_A_WL258vLB9_0),.clk(gclk));
	jdff dff_A_nyc2roSQ8_0(.dout(w_dff_A_wgWE2OIF4_0),.din(w_dff_A_nyc2roSQ8_0),.clk(gclk));
	jdff dff_A_wgWE2OIF4_0(.dout(w_dff_A_EQdiu7Rs7_0),.din(w_dff_A_wgWE2OIF4_0),.clk(gclk));
	jdff dff_A_EQdiu7Rs7_0(.dout(w_dff_A_7s1UEE4E9_0),.din(w_dff_A_EQdiu7Rs7_0),.clk(gclk));
	jdff dff_A_7s1UEE4E9_0(.dout(G301),.din(w_dff_A_7s1UEE4E9_0),.clk(gclk));
	jdff dff_A_5ZJ7pWXu5_2(.dout(w_dff_A_B9hm0S602_0),.din(w_dff_A_5ZJ7pWXu5_2),.clk(gclk));
	jdff dff_A_B9hm0S602_0(.dout(w_dff_A_62ACiwer7_0),.din(w_dff_A_B9hm0S602_0),.clk(gclk));
	jdff dff_A_62ACiwer7_0(.dout(w_dff_A_33B314zn1_0),.din(w_dff_A_62ACiwer7_0),.clk(gclk));
	jdff dff_A_33B314zn1_0(.dout(w_dff_A_1ORmC1Rr9_0),.din(w_dff_A_33B314zn1_0),.clk(gclk));
	jdff dff_A_1ORmC1Rr9_0(.dout(w_dff_A_UD0mHw0Y8_0),.din(w_dff_A_1ORmC1Rr9_0),.clk(gclk));
	jdff dff_A_UD0mHw0Y8_0(.dout(G304),.din(w_dff_A_UD0mHw0Y8_0),.clk(gclk));
	jdff dff_A_xlZ8L1W07_2(.dout(w_dff_A_8RsmyaiI5_0),.din(w_dff_A_xlZ8L1W07_2),.clk(gclk));
	jdff dff_A_8RsmyaiI5_0(.dout(w_dff_A_t1a9Lv1z5_0),.din(w_dff_A_8RsmyaiI5_0),.clk(gclk));
	jdff dff_A_t1a9Lv1z5_0(.dout(w_dff_A_1mvlSIxx1_0),.din(w_dff_A_t1a9Lv1z5_0),.clk(gclk));
	jdff dff_A_1mvlSIxx1_0(.dout(w_dff_A_OPuVijkx7_0),.din(w_dff_A_1mvlSIxx1_0),.clk(gclk));
	jdff dff_A_OPuVijkx7_0(.dout(w_dff_A_pN6rLBLl2_0),.din(w_dff_A_OPuVijkx7_0),.clk(gclk));
	jdff dff_A_pN6rLBLl2_0(.dout(w_dff_A_Enrz0vw03_0),.din(w_dff_A_pN6rLBLl2_0),.clk(gclk));
	jdff dff_A_Enrz0vw03_0(.dout(w_dff_A_ZNa2zk2F9_0),.din(w_dff_A_Enrz0vw03_0),.clk(gclk));
	jdff dff_A_ZNa2zk2F9_0(.dout(G307),.din(w_dff_A_ZNa2zk2F9_0),.clk(gclk));
	jdff dff_A_NpO6pto17_2(.dout(w_dff_A_yGWClJHQ3_0),.din(w_dff_A_NpO6pto17_2),.clk(gclk));
	jdff dff_A_yGWClJHQ3_0(.dout(w_dff_A_KVuEHkkb2_0),.din(w_dff_A_yGWClJHQ3_0),.clk(gclk));
	jdff dff_A_KVuEHkkb2_0(.dout(w_dff_A_Tx2EeQEC5_0),.din(w_dff_A_KVuEHkkb2_0),.clk(gclk));
	jdff dff_A_Tx2EeQEC5_0(.dout(w_dff_A_TRwoNDg73_0),.din(w_dff_A_Tx2EeQEC5_0),.clk(gclk));
	jdff dff_A_TRwoNDg73_0(.dout(w_dff_A_hikfPZ1u3_0),.din(w_dff_A_TRwoNDg73_0),.clk(gclk));
	jdff dff_A_hikfPZ1u3_0(.dout(w_dff_A_7TrXXuFg1_0),.din(w_dff_A_hikfPZ1u3_0),.clk(gclk));
	jdff dff_A_7TrXXuFg1_0(.dout(w_dff_A_xNhO77ex5_0),.din(w_dff_A_7TrXXuFg1_0),.clk(gclk));
	jdff dff_A_xNhO77ex5_0(.dout(w_dff_A_LNfNVx5v9_0),.din(w_dff_A_xNhO77ex5_0),.clk(gclk));
	jdff dff_A_LNfNVx5v9_0(.dout(w_dff_A_lNXZEEmI6_0),.din(w_dff_A_LNfNVx5v9_0),.clk(gclk));
	jdff dff_A_lNXZEEmI6_0(.dout(w_dff_A_sxzLpbNr9_0),.din(w_dff_A_lNXZEEmI6_0),.clk(gclk));
	jdff dff_A_sxzLpbNr9_0(.dout(w_dff_A_QgfBEcCl0_0),.din(w_dff_A_sxzLpbNr9_0),.clk(gclk));
	jdff dff_A_QgfBEcCl0_0(.dout(w_dff_A_H4nuQuD29_0),.din(w_dff_A_QgfBEcCl0_0),.clk(gclk));
	jdff dff_A_H4nuQuD29_0(.dout(w_dff_A_RmMNSInv4_0),.din(w_dff_A_H4nuQuD29_0),.clk(gclk));
	jdff dff_A_RmMNSInv4_0(.dout(w_dff_A_Cn0gG3nw8_0),.din(w_dff_A_RmMNSInv4_0),.clk(gclk));
	jdff dff_A_Cn0gG3nw8_0(.dout(w_dff_A_oEcxtlaH3_0),.din(w_dff_A_Cn0gG3nw8_0),.clk(gclk));
	jdff dff_A_oEcxtlaH3_0(.dout(w_dff_A_kBA3nHEg5_0),.din(w_dff_A_oEcxtlaH3_0),.clk(gclk));
	jdff dff_A_kBA3nHEg5_0(.dout(w_dff_A_z4pndscK5_0),.din(w_dff_A_kBA3nHEg5_0),.clk(gclk));
	jdff dff_A_z4pndscK5_0(.dout(w_dff_A_zg3xNFJl1_0),.din(w_dff_A_z4pndscK5_0),.clk(gclk));
	jdff dff_A_zg3xNFJl1_0(.dout(w_dff_A_Izr64Mtx0_0),.din(w_dff_A_zg3xNFJl1_0),.clk(gclk));
	jdff dff_A_Izr64Mtx0_0(.dout(G344),.din(w_dff_A_Izr64Mtx0_0),.clk(gclk));
	jdff dff_A_5xWKymr18_2(.dout(w_dff_A_HlcRKYcW8_0),.din(w_dff_A_5xWKymr18_2),.clk(gclk));
	jdff dff_A_HlcRKYcW8_0(.dout(G419),.din(w_dff_A_HlcRKYcW8_0),.clk(gclk));
	jdff dff_A_TNQyhMuw3_2(.dout(w_dff_A_kyRgxR5R7_0),.din(w_dff_A_TNQyhMuw3_2),.clk(gclk));
	jdff dff_A_kyRgxR5R7_0(.dout(G471),.din(w_dff_A_kyRgxR5R7_0),.clk(gclk));
	jdff dff_A_gjRLzgIm3_2(.dout(w_dff_A_JXazmYKP2_0),.din(w_dff_A_gjRLzgIm3_2),.clk(gclk));
	jdff dff_A_JXazmYKP2_0(.dout(w_dff_A_bEIjtywn2_0),.din(w_dff_A_JXazmYKP2_0),.clk(gclk));
	jdff dff_A_bEIjtywn2_0(.dout(w_dff_A_tPHdV3u70_0),.din(w_dff_A_bEIjtywn2_0),.clk(gclk));
	jdff dff_A_tPHdV3u70_0(.dout(w_dff_A_Lca0kmFz9_0),.din(w_dff_A_tPHdV3u70_0),.clk(gclk));
	jdff dff_A_Lca0kmFz9_0(.dout(w_dff_A_X3BxciBC4_0),.din(w_dff_A_Lca0kmFz9_0),.clk(gclk));
	jdff dff_A_X3BxciBC4_0(.dout(w_dff_A_VfdZ5erP6_0),.din(w_dff_A_X3BxciBC4_0),.clk(gclk));
	jdff dff_A_VfdZ5erP6_0(.dout(w_dff_A_nvN9YVzL6_0),.din(w_dff_A_VfdZ5erP6_0),.clk(gclk));
	jdff dff_A_nvN9YVzL6_0(.dout(w_dff_A_Ng5PWTK74_0),.din(w_dff_A_nvN9YVzL6_0),.clk(gclk));
	jdff dff_A_Ng5PWTK74_0(.dout(w_dff_A_SRISsozN2_0),.din(w_dff_A_Ng5PWTK74_0),.clk(gclk));
	jdff dff_A_SRISsozN2_0(.dout(w_dff_A_zK39wwoO4_0),.din(w_dff_A_SRISsozN2_0),.clk(gclk));
	jdff dff_A_zK39wwoO4_0(.dout(w_dff_A_n9IPYTyO1_0),.din(w_dff_A_zK39wwoO4_0),.clk(gclk));
	jdff dff_A_n9IPYTyO1_0(.dout(w_dff_A_4k3rMu2f9_0),.din(w_dff_A_n9IPYTyO1_0),.clk(gclk));
	jdff dff_A_4k3rMu2f9_0(.dout(w_dff_A_MAHEbFBd1_0),.din(w_dff_A_4k3rMu2f9_0),.clk(gclk));
	jdff dff_A_MAHEbFBd1_0(.dout(w_dff_A_Bmfi1Pd85_0),.din(w_dff_A_MAHEbFBd1_0),.clk(gclk));
	jdff dff_A_Bmfi1Pd85_0(.dout(w_dff_A_JWsvIb9c8_0),.din(w_dff_A_Bmfi1Pd85_0),.clk(gclk));
	jdff dff_A_JWsvIb9c8_0(.dout(w_dff_A_fy6XihzP7_0),.din(w_dff_A_JWsvIb9c8_0),.clk(gclk));
	jdff dff_A_fy6XihzP7_0(.dout(w_dff_A_6wJk8jyM6_0),.din(w_dff_A_fy6XihzP7_0),.clk(gclk));
	jdff dff_A_6wJk8jyM6_0(.dout(G359),.din(w_dff_A_6wJk8jyM6_0),.clk(gclk));
	jdff dff_A_A4XOy4fh6_2(.dout(w_dff_A_gTN6iNlU9_0),.din(w_dff_A_A4XOy4fh6_2),.clk(gclk));
	jdff dff_A_gTN6iNlU9_0(.dout(w_dff_A_GCu76aiM2_0),.din(w_dff_A_gTN6iNlU9_0),.clk(gclk));
	jdff dff_A_GCu76aiM2_0(.dout(w_dff_A_Vc4je3797_0),.din(w_dff_A_GCu76aiM2_0),.clk(gclk));
	jdff dff_A_Vc4je3797_0(.dout(w_dff_A_LcOUrM4m3_0),.din(w_dff_A_Vc4je3797_0),.clk(gclk));
	jdff dff_A_LcOUrM4m3_0(.dout(w_dff_A_Wp5C6Slw5_0),.din(w_dff_A_LcOUrM4m3_0),.clk(gclk));
	jdff dff_A_Wp5C6Slw5_0(.dout(w_dff_A_j7MCRLo46_0),.din(w_dff_A_Wp5C6Slw5_0),.clk(gclk));
	jdff dff_A_j7MCRLo46_0(.dout(w_dff_A_DBJGPkYD5_0),.din(w_dff_A_j7MCRLo46_0),.clk(gclk));
	jdff dff_A_DBJGPkYD5_0(.dout(w_dff_A_13cYZlMt2_0),.din(w_dff_A_DBJGPkYD5_0),.clk(gclk));
	jdff dff_A_13cYZlMt2_0(.dout(w_dff_A_zTHqLjhk6_0),.din(w_dff_A_13cYZlMt2_0),.clk(gclk));
	jdff dff_A_zTHqLjhk6_0(.dout(w_dff_A_6L7oKnnq6_0),.din(w_dff_A_zTHqLjhk6_0),.clk(gclk));
	jdff dff_A_6L7oKnnq6_0(.dout(w_dff_A_XyI0mOA96_0),.din(w_dff_A_6L7oKnnq6_0),.clk(gclk));
	jdff dff_A_XyI0mOA96_0(.dout(w_dff_A_CpHfLnY25_0),.din(w_dff_A_XyI0mOA96_0),.clk(gclk));
	jdff dff_A_CpHfLnY25_0(.dout(w_dff_A_ZqUBEiYz9_0),.din(w_dff_A_CpHfLnY25_0),.clk(gclk));
	jdff dff_A_ZqUBEiYz9_0(.dout(w_dff_A_8yoyiDDb7_0),.din(w_dff_A_ZqUBEiYz9_0),.clk(gclk));
	jdff dff_A_8yoyiDDb7_0(.dout(w_dff_A_0RTInmma9_0),.din(w_dff_A_8yoyiDDb7_0),.clk(gclk));
	jdff dff_A_0RTInmma9_0(.dout(w_dff_A_OhYKUvWI1_0),.din(w_dff_A_0RTInmma9_0),.clk(gclk));
	jdff dff_A_OhYKUvWI1_0(.dout(w_dff_A_UPZ5k5Xb9_0),.din(w_dff_A_OhYKUvWI1_0),.clk(gclk));
	jdff dff_A_UPZ5k5Xb9_0(.dout(G362),.din(w_dff_A_UPZ5k5Xb9_0),.clk(gclk));
	jdff dff_A_aqO8jZ6A6_2(.dout(w_dff_A_AZzDua9b3_0),.din(w_dff_A_aqO8jZ6A6_2),.clk(gclk));
	jdff dff_A_AZzDua9b3_0(.dout(w_dff_A_6YO4tzXl6_0),.din(w_dff_A_AZzDua9b3_0),.clk(gclk));
	jdff dff_A_6YO4tzXl6_0(.dout(w_dff_A_o0UazIW82_0),.din(w_dff_A_6YO4tzXl6_0),.clk(gclk));
	jdff dff_A_o0UazIW82_0(.dout(w_dff_A_YOBdtfMA2_0),.din(w_dff_A_o0UazIW82_0),.clk(gclk));
	jdff dff_A_YOBdtfMA2_0(.dout(w_dff_A_uCogFCmT3_0),.din(w_dff_A_YOBdtfMA2_0),.clk(gclk));
	jdff dff_A_uCogFCmT3_0(.dout(w_dff_A_xWT3jQs29_0),.din(w_dff_A_uCogFCmT3_0),.clk(gclk));
	jdff dff_A_xWT3jQs29_0(.dout(w_dff_A_72h9EVtj2_0),.din(w_dff_A_xWT3jQs29_0),.clk(gclk));
	jdff dff_A_72h9EVtj2_0(.dout(w_dff_A_YzK76lN63_0),.din(w_dff_A_72h9EVtj2_0),.clk(gclk));
	jdff dff_A_YzK76lN63_0(.dout(w_dff_A_TCxdCZHY1_0),.din(w_dff_A_YzK76lN63_0),.clk(gclk));
	jdff dff_A_TCxdCZHY1_0(.dout(w_dff_A_2UzDimiZ9_0),.din(w_dff_A_TCxdCZHY1_0),.clk(gclk));
	jdff dff_A_2UzDimiZ9_0(.dout(w_dff_A_7PP1sbCB6_0),.din(w_dff_A_2UzDimiZ9_0),.clk(gclk));
	jdff dff_A_7PP1sbCB6_0(.dout(w_dff_A_fQgQo2ye7_0),.din(w_dff_A_7PP1sbCB6_0),.clk(gclk));
	jdff dff_A_fQgQo2ye7_0(.dout(w_dff_A_5VkYQ8El0_0),.din(w_dff_A_fQgQo2ye7_0),.clk(gclk));
	jdff dff_A_5VkYQ8El0_0(.dout(w_dff_A_YGpfq2Jd9_0),.din(w_dff_A_5VkYQ8El0_0),.clk(gclk));
	jdff dff_A_YGpfq2Jd9_0(.dout(w_dff_A_aOSDakV86_0),.din(w_dff_A_YGpfq2Jd9_0),.clk(gclk));
	jdff dff_A_aOSDakV86_0(.dout(w_dff_A_Li7dGMDe5_0),.din(w_dff_A_aOSDakV86_0),.clk(gclk));
	jdff dff_A_Li7dGMDe5_0(.dout(w_dff_A_6NQCOJIc2_0),.din(w_dff_A_Li7dGMDe5_0),.clk(gclk));
	jdff dff_A_6NQCOJIc2_0(.dout(G365),.din(w_dff_A_6NQCOJIc2_0),.clk(gclk));
	jdff dff_A_7pKYbPVy4_2(.dout(w_dff_A_WBGl0WpB8_0),.din(w_dff_A_7pKYbPVy4_2),.clk(gclk));
	jdff dff_A_WBGl0WpB8_0(.dout(w_dff_A_WhsXkAvs8_0),.din(w_dff_A_WBGl0WpB8_0),.clk(gclk));
	jdff dff_A_WhsXkAvs8_0(.dout(w_dff_A_CDe5Np1a1_0),.din(w_dff_A_WhsXkAvs8_0),.clk(gclk));
	jdff dff_A_CDe5Np1a1_0(.dout(w_dff_A_akKupNvi7_0),.din(w_dff_A_CDe5Np1a1_0),.clk(gclk));
	jdff dff_A_akKupNvi7_0(.dout(w_dff_A_iWlaiOJf0_0),.din(w_dff_A_akKupNvi7_0),.clk(gclk));
	jdff dff_A_iWlaiOJf0_0(.dout(w_dff_A_eQUQsWTy3_0),.din(w_dff_A_iWlaiOJf0_0),.clk(gclk));
	jdff dff_A_eQUQsWTy3_0(.dout(w_dff_A_adO26Uvs3_0),.din(w_dff_A_eQUQsWTy3_0),.clk(gclk));
	jdff dff_A_adO26Uvs3_0(.dout(w_dff_A_LgSqa9uP7_0),.din(w_dff_A_adO26Uvs3_0),.clk(gclk));
	jdff dff_A_LgSqa9uP7_0(.dout(w_dff_A_eHYOdJuD0_0),.din(w_dff_A_LgSqa9uP7_0),.clk(gclk));
	jdff dff_A_eHYOdJuD0_0(.dout(w_dff_A_06QDEm150_0),.din(w_dff_A_eHYOdJuD0_0),.clk(gclk));
	jdff dff_A_06QDEm150_0(.dout(w_dff_A_Uk1kWr2b3_0),.din(w_dff_A_06QDEm150_0),.clk(gclk));
	jdff dff_A_Uk1kWr2b3_0(.dout(w_dff_A_jphJM6sA5_0),.din(w_dff_A_Uk1kWr2b3_0),.clk(gclk));
	jdff dff_A_jphJM6sA5_0(.dout(w_dff_A_KZnSz4oG9_0),.din(w_dff_A_jphJM6sA5_0),.clk(gclk));
	jdff dff_A_KZnSz4oG9_0(.dout(w_dff_A_FsiRgk9F2_0),.din(w_dff_A_KZnSz4oG9_0),.clk(gclk));
	jdff dff_A_FsiRgk9F2_0(.dout(w_dff_A_npPxXng34_0),.din(w_dff_A_FsiRgk9F2_0),.clk(gclk));
	jdff dff_A_npPxXng34_0(.dout(w_dff_A_tggbj35D0_0),.din(w_dff_A_npPxXng34_0),.clk(gclk));
	jdff dff_A_tggbj35D0_0(.dout(w_dff_A_f6zmQDRH2_0),.din(w_dff_A_tggbj35D0_0),.clk(gclk));
	jdff dff_A_f6zmQDRH2_0(.dout(G368),.din(w_dff_A_f6zmQDRH2_0),.clk(gclk));
	jdff dff_A_QExPo0Wj9_2(.dout(w_dff_A_zjSrlHje7_0),.din(w_dff_A_QExPo0Wj9_2),.clk(gclk));
	jdff dff_A_zjSrlHje7_0(.dout(w_dff_A_64PeerYV0_0),.din(w_dff_A_zjSrlHje7_0),.clk(gclk));
	jdff dff_A_64PeerYV0_0(.dout(w_dff_A_joX9QhWi4_0),.din(w_dff_A_64PeerYV0_0),.clk(gclk));
	jdff dff_A_joX9QhWi4_0(.dout(w_dff_A_F4x6EZGn9_0),.din(w_dff_A_joX9QhWi4_0),.clk(gclk));
	jdff dff_A_F4x6EZGn9_0(.dout(w_dff_A_I58el1FW9_0),.din(w_dff_A_F4x6EZGn9_0),.clk(gclk));
	jdff dff_A_I58el1FW9_0(.dout(w_dff_A_n7JEDQ8V9_0),.din(w_dff_A_I58el1FW9_0),.clk(gclk));
	jdff dff_A_n7JEDQ8V9_0(.dout(w_dff_A_Muat5UCv8_0),.din(w_dff_A_n7JEDQ8V9_0),.clk(gclk));
	jdff dff_A_Muat5UCv8_0(.dout(w_dff_A_npOvNuPR5_0),.din(w_dff_A_Muat5UCv8_0),.clk(gclk));
	jdff dff_A_npOvNuPR5_0(.dout(w_dff_A_cigL26PG5_0),.din(w_dff_A_npOvNuPR5_0),.clk(gclk));
	jdff dff_A_cigL26PG5_0(.dout(w_dff_A_v1AWzzSo9_0),.din(w_dff_A_cigL26PG5_0),.clk(gclk));
	jdff dff_A_v1AWzzSo9_0(.dout(w_dff_A_6D9PtInS1_0),.din(w_dff_A_v1AWzzSo9_0),.clk(gclk));
	jdff dff_A_6D9PtInS1_0(.dout(w_dff_A_77ssRZCb2_0),.din(w_dff_A_6D9PtInS1_0),.clk(gclk));
	jdff dff_A_77ssRZCb2_0(.dout(G347),.din(w_dff_A_77ssRZCb2_0),.clk(gclk));
	jdff dff_A_RRVhlcbP2_2(.dout(w_dff_A_Y3duYJiR3_0),.din(w_dff_A_RRVhlcbP2_2),.clk(gclk));
	jdff dff_A_Y3duYJiR3_0(.dout(w_dff_A_XZea749D9_0),.din(w_dff_A_Y3duYJiR3_0),.clk(gclk));
	jdff dff_A_XZea749D9_0(.dout(w_dff_A_cd9govl93_0),.din(w_dff_A_XZea749D9_0),.clk(gclk));
	jdff dff_A_cd9govl93_0(.dout(w_dff_A_BiAC9qPC4_0),.din(w_dff_A_cd9govl93_0),.clk(gclk));
	jdff dff_A_BiAC9qPC4_0(.dout(w_dff_A_SdAU7V2Q1_0),.din(w_dff_A_BiAC9qPC4_0),.clk(gclk));
	jdff dff_A_SdAU7V2Q1_0(.dout(w_dff_A_tVFX3nj97_0),.din(w_dff_A_SdAU7V2Q1_0),.clk(gclk));
	jdff dff_A_tVFX3nj97_0(.dout(w_dff_A_Xy2JumR71_0),.din(w_dff_A_tVFX3nj97_0),.clk(gclk));
	jdff dff_A_Xy2JumR71_0(.dout(w_dff_A_eZlrCZqr9_0),.din(w_dff_A_Xy2JumR71_0),.clk(gclk));
	jdff dff_A_eZlrCZqr9_0(.dout(w_dff_A_hvHvB2zE9_0),.din(w_dff_A_eZlrCZqr9_0),.clk(gclk));
	jdff dff_A_hvHvB2zE9_0(.dout(w_dff_A_fYKJRhen9_0),.din(w_dff_A_hvHvB2zE9_0),.clk(gclk));
	jdff dff_A_fYKJRhen9_0(.dout(w_dff_A_lCZJMyYO7_0),.din(w_dff_A_fYKJRhen9_0),.clk(gclk));
	jdff dff_A_lCZJMyYO7_0(.dout(w_dff_A_ko2P7GjQ4_0),.din(w_dff_A_lCZJMyYO7_0),.clk(gclk));
	jdff dff_A_ko2P7GjQ4_0(.dout(w_dff_A_Dtcr2t8E9_0),.din(w_dff_A_ko2P7GjQ4_0),.clk(gclk));
	jdff dff_A_Dtcr2t8E9_0(.dout(G350),.din(w_dff_A_Dtcr2t8E9_0),.clk(gclk));
	jdff dff_A_lnookEJx5_2(.dout(w_dff_A_hFSAKiyw3_0),.din(w_dff_A_lnookEJx5_2),.clk(gclk));
	jdff dff_A_hFSAKiyw3_0(.dout(w_dff_A_JEcEXyYJ5_0),.din(w_dff_A_hFSAKiyw3_0),.clk(gclk));
	jdff dff_A_JEcEXyYJ5_0(.dout(w_dff_A_xGtgUL8o3_0),.din(w_dff_A_JEcEXyYJ5_0),.clk(gclk));
	jdff dff_A_xGtgUL8o3_0(.dout(w_dff_A_nB9rpTsv6_0),.din(w_dff_A_xGtgUL8o3_0),.clk(gclk));
	jdff dff_A_nB9rpTsv6_0(.dout(w_dff_A_WQGQdT9K8_0),.din(w_dff_A_nB9rpTsv6_0),.clk(gclk));
	jdff dff_A_WQGQdT9K8_0(.dout(w_dff_A_pl2xJzib4_0),.din(w_dff_A_WQGQdT9K8_0),.clk(gclk));
	jdff dff_A_pl2xJzib4_0(.dout(w_dff_A_wnqCkNDS2_0),.din(w_dff_A_pl2xJzib4_0),.clk(gclk));
	jdff dff_A_wnqCkNDS2_0(.dout(w_dff_A_HwJX9iCr2_0),.din(w_dff_A_wnqCkNDS2_0),.clk(gclk));
	jdff dff_A_HwJX9iCr2_0(.dout(w_dff_A_z4uEjMGn0_0),.din(w_dff_A_HwJX9iCr2_0),.clk(gclk));
	jdff dff_A_z4uEjMGn0_0(.dout(w_dff_A_3WBHduyB5_0),.din(w_dff_A_z4uEjMGn0_0),.clk(gclk));
	jdff dff_A_3WBHduyB5_0(.dout(w_dff_A_klBuYOAh1_0),.din(w_dff_A_3WBHduyB5_0),.clk(gclk));
	jdff dff_A_klBuYOAh1_0(.dout(w_dff_A_8Wg1UBbA2_0),.din(w_dff_A_klBuYOAh1_0),.clk(gclk));
	jdff dff_A_8Wg1UBbA2_0(.dout(w_dff_A_o2PvDGlQ1_0),.din(w_dff_A_8Wg1UBbA2_0),.clk(gclk));
	jdff dff_A_o2PvDGlQ1_0(.dout(w_dff_A_RrFeEEwF1_0),.din(w_dff_A_o2PvDGlQ1_0),.clk(gclk));
	jdff dff_A_RrFeEEwF1_0(.dout(w_dff_A_wX30sGNI9_0),.din(w_dff_A_RrFeEEwF1_0),.clk(gclk));
	jdff dff_A_wX30sGNI9_0(.dout(G353),.din(w_dff_A_wX30sGNI9_0),.clk(gclk));
	jdff dff_A_fSEwKRmD3_2(.dout(w_dff_A_tdsQ6rES9_0),.din(w_dff_A_fSEwKRmD3_2),.clk(gclk));
	jdff dff_A_tdsQ6rES9_0(.dout(w_dff_A_hLvOlyGW9_0),.din(w_dff_A_tdsQ6rES9_0),.clk(gclk));
	jdff dff_A_hLvOlyGW9_0(.dout(w_dff_A_Hwn6ljTY8_0),.din(w_dff_A_hLvOlyGW9_0),.clk(gclk));
	jdff dff_A_Hwn6ljTY8_0(.dout(w_dff_A_6oZDhHqT0_0),.din(w_dff_A_Hwn6ljTY8_0),.clk(gclk));
	jdff dff_A_6oZDhHqT0_0(.dout(w_dff_A_LAsdIJpO2_0),.din(w_dff_A_6oZDhHqT0_0),.clk(gclk));
	jdff dff_A_LAsdIJpO2_0(.dout(w_dff_A_ZTTy8cRz9_0),.din(w_dff_A_LAsdIJpO2_0),.clk(gclk));
	jdff dff_A_ZTTy8cRz9_0(.dout(w_dff_A_oaqnHzPb4_0),.din(w_dff_A_ZTTy8cRz9_0),.clk(gclk));
	jdff dff_A_oaqnHzPb4_0(.dout(w_dff_A_asSJdhsN3_0),.din(w_dff_A_oaqnHzPb4_0),.clk(gclk));
	jdff dff_A_asSJdhsN3_0(.dout(w_dff_A_icCUAyOh3_0),.din(w_dff_A_asSJdhsN3_0),.clk(gclk));
	jdff dff_A_icCUAyOh3_0(.dout(w_dff_A_zGpUNtdD2_0),.din(w_dff_A_icCUAyOh3_0),.clk(gclk));
	jdff dff_A_zGpUNtdD2_0(.dout(w_dff_A_UpoGRkq93_0),.din(w_dff_A_zGpUNtdD2_0),.clk(gclk));
	jdff dff_A_UpoGRkq93_0(.dout(w_dff_A_bK9inClz4_0),.din(w_dff_A_UpoGRkq93_0),.clk(gclk));
	jdff dff_A_bK9inClz4_0(.dout(w_dff_A_557gcgzR0_0),.din(w_dff_A_bK9inClz4_0),.clk(gclk));
	jdff dff_A_557gcgzR0_0(.dout(w_dff_A_iFGbiI5M0_0),.din(w_dff_A_557gcgzR0_0),.clk(gclk));
	jdff dff_A_iFGbiI5M0_0(.dout(w_dff_A_CMGYIz2W0_0),.din(w_dff_A_iFGbiI5M0_0),.clk(gclk));
	jdff dff_A_CMGYIz2W0_0(.dout(w_dff_A_G4LGUiy17_0),.din(w_dff_A_CMGYIz2W0_0),.clk(gclk));
	jdff dff_A_G4LGUiy17_0(.dout(w_dff_A_C2zreAzv5_0),.din(w_dff_A_G4LGUiy17_0),.clk(gclk));
	jdff dff_A_C2zreAzv5_0(.dout(G356),.din(w_dff_A_C2zreAzv5_0),.clk(gclk));
	jdff dff_A_kjGGFBjr5_2(.dout(w_dff_A_mIhX1E8q9_0),.din(w_dff_A_kjGGFBjr5_2),.clk(gclk));
	jdff dff_A_mIhX1E8q9_0(.dout(w_dff_A_63iv9Lgt4_0),.din(w_dff_A_mIhX1E8q9_0),.clk(gclk));
	jdff dff_A_63iv9Lgt4_0(.dout(w_dff_A_syg62Qgg5_0),.din(w_dff_A_63iv9Lgt4_0),.clk(gclk));
	jdff dff_A_syg62Qgg5_0(.dout(w_dff_A_XbNGlsgT6_0),.din(w_dff_A_syg62Qgg5_0),.clk(gclk));
	jdff dff_A_XbNGlsgT6_0(.dout(w_dff_A_ocJ5WiQt8_0),.din(w_dff_A_XbNGlsgT6_0),.clk(gclk));
	jdff dff_A_ocJ5WiQt8_0(.dout(G321),.din(w_dff_A_ocJ5WiQt8_0),.clk(gclk));
	jdff dff_A_3AVLPWfs6_2(.dout(G338),.din(w_dff_A_3AVLPWfs6_2),.clk(gclk));
	jdff dff_A_oM4MwWtI5_2(.dout(w_dff_A_o8QafsO16_0),.din(w_dff_A_oM4MwWtI5_2),.clk(gclk));
	jdff dff_A_o8QafsO16_0(.dout(w_dff_A_Jqd4xWpb1_0),.din(w_dff_A_o8QafsO16_0),.clk(gclk));
	jdff dff_A_Jqd4xWpb1_0(.dout(w_dff_A_Yo2qFoKU9_0),.din(w_dff_A_Jqd4xWpb1_0),.clk(gclk));
	jdff dff_A_Yo2qFoKU9_0(.dout(w_dff_A_pom0h5kE6_0),.din(w_dff_A_Yo2qFoKU9_0),.clk(gclk));
	jdff dff_A_pom0h5kE6_0(.dout(w_dff_A_OozD2UhM1_0),.din(w_dff_A_pom0h5kE6_0),.clk(gclk));
	jdff dff_A_OozD2UhM1_0(.dout(w_dff_A_BgCpmlhe9_0),.din(w_dff_A_OozD2UhM1_0),.clk(gclk));
	jdff dff_A_BgCpmlhe9_0(.dout(w_dff_A_QBrIUpQs0_0),.din(w_dff_A_BgCpmlhe9_0),.clk(gclk));
	jdff dff_A_QBrIUpQs0_0(.dout(w_dff_A_NpIy8QxP0_0),.din(w_dff_A_QBrIUpQs0_0),.clk(gclk));
	jdff dff_A_NpIy8QxP0_0(.dout(w_dff_A_eRzlU6yE5_0),.din(w_dff_A_NpIy8QxP0_0),.clk(gclk));
	jdff dff_A_eRzlU6yE5_0(.dout(w_dff_A_bi5YO1QB7_0),.din(w_dff_A_eRzlU6yE5_0),.clk(gclk));
	jdff dff_A_bi5YO1QB7_0(.dout(w_dff_A_patlHC8c3_0),.din(w_dff_A_bi5YO1QB7_0),.clk(gclk));
	jdff dff_A_patlHC8c3_0(.dout(w_dff_A_HCOqsXlx4_0),.din(w_dff_A_patlHC8c3_0),.clk(gclk));
	jdff dff_A_HCOqsXlx4_0(.dout(w_dff_A_caS97pzf2_0),.din(w_dff_A_HCOqsXlx4_0),.clk(gclk));
	jdff dff_A_caS97pzf2_0(.dout(w_dff_A_5HZDyfup5_0),.din(w_dff_A_caS97pzf2_0),.clk(gclk));
	jdff dff_A_5HZDyfup5_0(.dout(w_dff_A_04DFZzRO4_0),.din(w_dff_A_5HZDyfup5_0),.clk(gclk));
	jdff dff_A_04DFZzRO4_0(.dout(w_dff_A_iBbCuLEp4_0),.din(w_dff_A_04DFZzRO4_0),.clk(gclk));
	jdff dff_A_iBbCuLEp4_0(.dout(G370),.din(w_dff_A_iBbCuLEp4_0),.clk(gclk));
	jdff dff_A_SZHKifOh5_2(.dout(w_dff_A_xrM9NinU7_0),.din(w_dff_A_SZHKifOh5_2),.clk(gclk));
	jdff dff_A_xrM9NinU7_0(.dout(w_dff_A_faxxTd5s3_0),.din(w_dff_A_xrM9NinU7_0),.clk(gclk));
	jdff dff_A_faxxTd5s3_0(.dout(w_dff_A_4ctQpcnd2_0),.din(w_dff_A_faxxTd5s3_0),.clk(gclk));
	jdff dff_A_4ctQpcnd2_0(.dout(w_dff_A_iDNk4g734_0),.din(w_dff_A_4ctQpcnd2_0),.clk(gclk));
	jdff dff_A_iDNk4g734_0(.dout(w_dff_A_PSY8VEdo3_0),.din(w_dff_A_iDNk4g734_0),.clk(gclk));
	jdff dff_A_PSY8VEdo3_0(.dout(w_dff_A_eOFAMxXJ6_0),.din(w_dff_A_PSY8VEdo3_0),.clk(gclk));
	jdff dff_A_eOFAMxXJ6_0(.dout(w_dff_A_QS29gxdM5_0),.din(w_dff_A_eOFAMxXJ6_0),.clk(gclk));
	jdff dff_A_QS29gxdM5_0(.dout(w_dff_A_UqQwMQpd0_0),.din(w_dff_A_QS29gxdM5_0),.clk(gclk));
	jdff dff_A_UqQwMQpd0_0(.dout(w_dff_A_sNl1j9sY2_0),.din(w_dff_A_UqQwMQpd0_0),.clk(gclk));
	jdff dff_A_sNl1j9sY2_0(.dout(w_dff_A_eVXWxF4r8_0),.din(w_dff_A_sNl1j9sY2_0),.clk(gclk));
	jdff dff_A_eVXWxF4r8_0(.dout(w_dff_A_LVLxvjpj1_0),.din(w_dff_A_eVXWxF4r8_0),.clk(gclk));
	jdff dff_A_LVLxvjpj1_0(.dout(w_dff_A_utWrhI8o3_0),.din(w_dff_A_LVLxvjpj1_0),.clk(gclk));
	jdff dff_A_utWrhI8o3_0(.dout(w_dff_A_j3c1f5To7_0),.din(w_dff_A_utWrhI8o3_0),.clk(gclk));
	jdff dff_A_j3c1f5To7_0(.dout(w_dff_A_EnSTdf7g6_0),.din(w_dff_A_j3c1f5To7_0),.clk(gclk));
	jdff dff_A_EnSTdf7g6_0(.dout(w_dff_A_1vJFTEEo4_0),.din(w_dff_A_EnSTdf7g6_0),.clk(gclk));
	jdff dff_A_1vJFTEEo4_0(.dout(w_dff_A_Jt6aMDQ94_0),.din(w_dff_A_1vJFTEEo4_0),.clk(gclk));
	jdff dff_A_Jt6aMDQ94_0(.dout(w_dff_A_9ZIm3fD33_0),.din(w_dff_A_Jt6aMDQ94_0),.clk(gclk));
	jdff dff_A_9ZIm3fD33_0(.dout(w_dff_A_2MSuZMVk5_0),.din(w_dff_A_9ZIm3fD33_0),.clk(gclk));
	jdff dff_A_2MSuZMVk5_0(.dout(w_dff_A_Tm1UH8M69_0),.din(w_dff_A_2MSuZMVk5_0),.clk(gclk));
	jdff dff_A_Tm1UH8M69_0(.dout(w_dff_A_qp69ew1k3_0),.din(w_dff_A_Tm1UH8M69_0),.clk(gclk));
	jdff dff_A_qp69ew1k3_0(.dout(G399),.din(w_dff_A_qp69ew1k3_0),.clk(gclk));
endmodule

