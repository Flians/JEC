/*

c432:
	jxor: 1
	jspl: 84
	jspl3: 48
	jnot: 47
	jdff: 1154
	jand: 104
	jor: 104

Summary:
	jxor: 1
	jspl: 84
	jspl3: 48
	jnot: 47
	jdff: 1154
	jand: 104
	jor: 104
*/

module c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n43;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G4gat_0;
	wire [2:0] w_G8gat_0;
	wire [2:0] w_G11gat_0;
	wire [2:0] w_G14gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G21gat_0;
	wire [2:0] w_G24gat_0;
	wire [1:0] w_G27gat_0;
	wire [2:0] w_G30gat_0;
	wire [2:0] w_G34gat_0;
	wire [1:0] w_G40gat_0;
	wire [1:0] w_G43gat_0;
	wire [2:0] w_G47gat_0;
	wire [1:0] w_G50gat_0;
	wire [1:0] w_G53gat_0;
	wire [2:0] w_G56gat_0;
	wire [1:0] w_G56gat_1;
	wire [1:0] w_G60gat_0;
	wire [2:0] w_G63gat_0;
	wire [2:0] w_G66gat_0;
	wire [2:0] w_G69gat_0;
	wire [2:0] w_G73gat_0;
	wire [2:0] w_G76gat_0;
	wire [1:0] w_G79gat_0;
	wire [2:0] w_G82gat_0;
	wire [2:0] w_G86gat_0;
	wire [2:0] w_G89gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G95gat_0;
	wire [2:0] w_G99gat_0;
	wire [1:0] w_G102gat_0;
	wire [1:0] w_G105gat_0;
	wire [2:0] w_G108gat_0;
	wire [2:0] w_G112gat_0;
	wire [1:0] w_G115gat_0;
	wire [2:0] w_G223gat_0;
	wire [2:0] w_G223gat_1;
	wire [2:0] w_G223gat_2;
	wire [2:0] w_G223gat_3;
	wire w_G223gat_4;
	wire G223gat_fa_;
	wire [2:0] w_G329gat_0;
	wire [2:0] w_G329gat_1;
	wire [2:0] w_G329gat_2;
	wire [2:0] w_G329gat_3;
	wire w_G329gat_4;
	wire G329gat_fa_;
	wire [2:0] w_G370gat_0;
	wire [1:0] w_G370gat_1;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire [1:0] w_n43_0;
	wire [1:0] w_n44_0;
	wire [1:0] w_n45_0;
	wire [2:0] w_n46_0;
	wire [1:0] w_n47_0;
	wire [1:0] w_n49_0;
	wire [1:0] w_n51_0;
	wire [1:0] w_n54_0;
	wire [1:0] w_n57_0;
	wire [1:0] w_n60_0;
	wire [1:0] w_n62_0;
	wire [1:0] w_n64_0;
	wire [1:0] w_n70_0;
	wire [1:0] w_n73_0;
	wire [1:0] w_n75_0;
	wire [1:0] w_n78_0;
	wire [1:0] w_n80_0;
	wire [1:0] w_n81_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n86_0;
	wire [1:0] w_n88_0;
	wire [2:0] w_n93_0;
	wire [2:0] w_n93_1;
	wire [2:0] w_n93_2;
	wire [2:0] w_n93_3;
	wire [1:0] w_n95_0;
	wire [1:0] w_n102_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n106_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n111_0;
	wire [1:0] w_n113_0;
	wire [1:0] w_n117_0;
	wire [2:0] w_n119_0;
	wire [1:0] w_n120_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n123_0;
	wire [1:0] w_n125_0;
	wire [1:0] w_n127_0;
	wire [2:0] w_n131_0;
	wire [1:0] w_n138_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n141_0;
	wire [1:0] w_n144_0;
	wire [1:0] w_n145_0;
	wire [1:0] w_n147_0;
	wire [1:0] w_n149_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n156_0;
	wire [1:0] w_n159_0;
	wire [1:0] w_n164_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n173_0;
	wire [2:0] w_n181_0;
	wire [2:0] w_n181_1;
	wire [2:0] w_n181_2;
	wire [1:0] w_n183_0;
	wire [1:0] w_n185_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n202_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n206_0;
	wire [1:0] w_n209_0;
	wire [1:0] w_n211_0;
	wire [1:0] w_n222_0;
	wire [1:0] w_n227_0;
	wire [1:0] w_n230_0;
	wire [2:0] w_n246_0;
	wire [2:0] w_n246_1;
	wire [2:0] w_n246_2;
	wire [1:0] w_n248_0;
	wire [1:0] w_n250_0;
	wire [1:0] w_n251_0;
	wire [1:0] w_n253_0;
	wire [1:0] w_n254_0;
	wire [1:0] w_n257_0;
	wire [1:0] w_n264_0;
	wire [1:0] w_n265_0;
	wire [1:0] w_n269_0;
	wire [1:0] w_n271_0;
	wire [1:0] w_n281_0;
	wire [1:0] w_n288_0;
	wire [1:0] w_n290_0;
	wire w_dff_B_nNqmRsp24_0;
	wire w_dff_B_DPvU5Quz3_0;
	wire w_dff_B_y6Q9Vrdi5_0;
	wire w_dff_B_LEU6kzmi3_0;
	wire w_dff_B_MbNAgu3c0_0;
	wire w_dff_B_iPSNwcO46_0;
	wire w_dff_B_hlDujAZe1_0;
	wire w_dff_B_S8fN2eSL6_0;
	wire w_dff_B_fn3dAsWe4_0;
	wire w_dff_B_gm120Oud6_2;
	wire w_dff_A_CGsl3pof0_0;
	wire w_dff_B_26IILePm0_2;
	wire w_dff_A_q7Tu8nTb4_1;
	wire w_dff_B_NKNZqV8m2_1;
	wire w_dff_B_JcokKGtz9_1;
	wire w_dff_B_GlRJCYin5_1;
	wire w_dff_B_1wOjlkoT3_1;
	wire w_dff_B_QU1k9qCM4_1;
	wire w_dff_B_HXxjs9fd1_1;
	wire w_dff_B_0UYRfxd18_1;
	wire w_dff_B_MQvrzUcL1_1;
	wire w_dff_B_gYK1ymEv1_1;
	wire w_dff_B_iDH25Nws7_1;
	wire w_dff_B_M4gRjj490_1;
	wire w_dff_B_Pd4PdKN34_1;
	wire w_dff_B_11ePEZrX5_1;
	wire w_dff_B_PmLR5C9Z9_1;
	wire w_dff_B_HzFvrYs33_1;
	wire w_dff_B_rNUSAL3o8_1;
	wire w_dff_B_ek5lLYeP0_1;
	wire w_dff_B_u2pTCMcv7_1;
	wire w_dff_B_Jo5vL0Ub8_1;
	wire w_dff_B_vHqkHYop4_1;
	wire w_dff_B_3e5MOXWc9_1;
	wire w_dff_B_3vLTyasL5_1;
	wire w_dff_B_RuN9JMrB1_1;
	wire w_dff_B_m2yO53ZN7_1;
	wire w_dff_B_SFkrwljf0_2;
	wire w_dff_A_JFZSl3S94_0;
	wire w_dff_A_StAWxQvm3_0;
	wire w_dff_A_IoJGLttf4_0;
	wire w_dff_B_MTftNmki7_1;
	wire w_dff_A_M7m9KzrF2_0;
	wire w_dff_A_eeWmzvKG2_0;
	wire w_dff_A_tSs5Q0CR8_0;
	wire w_dff_A_gitFoMzA3_0;
	wire w_dff_A_KGuYjPc29_0;
	wire w_dff_A_XTA5sNUR6_0;
	wire w_dff_B_hTfrpH2X9_1;
	wire w_dff_B_Hni7MjoT2_1;
	wire w_dff_B_s6XJgI8S8_1;
	wire w_dff_B_OgWkF7Jl6_1;
	wire w_dff_B_zEtFVFdN7_1;
	wire w_dff_B_XL0xSoKd8_1;
	wire w_dff_B_JAMoUcrp2_1;
	wire w_dff_B_52tih4US5_0;
	wire w_dff_B_a3R5Amyo4_0;
	wire w_dff_B_DS6bcRlE0_0;
	wire w_dff_B_yMwr3pGu7_0;
	wire w_dff_A_cnSOicKp4_1;
	wire w_dff_A_3iMvnEdv2_1;
	wire w_dff_A_PP6xv8B28_1;
	wire w_dff_A_G1zTjTjC7_1;
	wire w_dff_A_USMqUlZT0_1;
	wire w_dff_B_9IqYxDq65_1;
	wire w_dff_B_rbsEoq272_0;
	wire w_dff_A_6w3XrPb50_0;
	wire w_dff_A_P6xyLfQo8_0;
	wire w_dff_A_TbntlUCQ0_0;
	wire w_dff_A_niiZHyDf9_0;
	wire w_dff_A_eNncHZYl5_0;
	wire w_dff_A_iNsHqmcB9_0;
	wire w_dff_A_75bDSFoY0_0;
	wire w_dff_A_NHcGcBLA5_0;
	wire w_dff_A_RILjHrJd7_0;
	wire w_dff_A_X4OhDqV63_0;
	wire w_dff_A_6I3Xz4tf1_0;
	wire w_dff_B_cdYsUHPR7_2;
	wire w_dff_B_PigP3P9I7_2;
	wire w_dff_B_t3QDEiRX2_2;
	wire w_dff_B_lyURepkx2_2;
	wire w_dff_B_3B9PK8623_2;
	wire w_dff_B_klbztqoW1_2;
	wire w_dff_B_Ay7FmcZt3_2;
	wire w_dff_B_a4PjgekG0_2;
	wire w_dff_B_0sLZaZ0C9_2;
	wire w_dff_B_Dwxc4tOo5_2;
	wire w_dff_B_53WsXVy56_2;
	wire w_dff_B_ZKIIDDwF9_2;
	wire w_dff_B_VLULyZFX3_2;
	wire w_dff_B_meL2PgNV6_2;
	wire w_dff_A_pna7zWFq8_0;
	wire w_dff_A_6SuufCPf4_0;
	wire w_dff_A_foeaykq62_0;
	wire w_dff_A_4znjuRdk8_0;
	wire w_dff_A_OwzA9siF2_0;
	wire w_dff_A_QICiSLGL9_0;
	wire w_dff_A_XkXZ0vP80_0;
	wire w_dff_A_oOu6h61c0_0;
	wire w_dff_A_iDlsSKQD2_0;
	wire w_dff_A_6CgZkNlh1_0;
	wire w_dff_A_zs8YKF2e3_0;
	wire w_dff_B_d8WufGIU6_2;
	wire w_dff_B_HS906qcc6_2;
	wire w_dff_B_emxqyXlt3_2;
	wire w_dff_B_GShhl6df7_2;
	wire w_dff_B_IzvDEbq43_2;
	wire w_dff_B_Qfzo6o843_2;
	wire w_dff_B_xAKdQLAb0_2;
	wire w_dff_B_IOM21WA49_2;
	wire w_dff_B_hPfCIXVH7_2;
	wire w_dff_B_NdxVDHo48_2;
	wire w_dff_B_2ZOsculb0_2;
	wire w_dff_B_PkP4nR5V3_2;
	wire w_dff_B_gN3uTzN49_2;
	wire w_dff_B_i1S2LK491_2;
	wire w_dff_B_hSN3jX8C9_1;
	wire w_dff_B_UN0gIONJ9_1;
	wire w_dff_B_quwS2UZ37_1;
	wire w_dff_B_eMfrHHK78_1;
	wire w_dff_B_bQEPOnxS9_1;
	wire w_dff_B_GUzvpdtD6_1;
	wire w_dff_B_jhOqW2AQ2_1;
	wire w_dff_B_H7cAMaLf2_1;
	wire w_dff_B_KzVFbklm1_1;
	wire w_dff_B_bvFIEeEr2_1;
	wire w_dff_B_IpfMBLA47_1;
	wire w_dff_B_8nLJvSQB1_1;
	wire w_dff_B_OtfSRp3W8_1;
	wire w_dff_B_CSHAgvXc6_1;
	wire w_dff_B_ahpQh7Hq2_1;
	wire w_dff_B_H9eeFopC3_1;
	wire w_dff_B_3ybyy3hW3_1;
	wire w_dff_B_ZERgL2zy9_1;
	wire w_dff_B_0FtBJo2C0_1;
	wire w_dff_B_eMTLxAtr9_1;
	wire w_dff_B_X8pu3I4w2_1;
	wire w_dff_B_FppoivKJ5_1;
	wire w_dff_B_JqgPeDQ92_1;
	wire w_dff_B_Pm1mYZYb5_1;
	wire w_dff_B_9eoe5DiQ4_1;
	wire w_dff_B_y119Gm4e1_1;
	wire w_dff_B_PPTVKxs89_1;
	wire w_dff_B_6hCX4gzq3_1;
	wire w_dff_A_hbIzBRil4_0;
	wire w_dff_A_xWkEArkY2_0;
	wire w_dff_A_VzSf0tvp2_0;
	wire w_dff_A_MOnorS0Q2_0;
	wire w_dff_A_LoqwA0X89_0;
	wire w_dff_B_o1HFGAr20_2;
	wire w_dff_B_kwWDYk5C7_2;
	wire w_dff_B_TAQ6QRbC4_2;
	wire w_dff_B_D2DJvxiQ0_2;
	wire w_dff_B_8tIFyV6u7_2;
	wire w_dff_B_ShlRA1jJ9_2;
	wire w_dff_B_MFHLqJBc9_2;
	wire w_dff_B_Tbepjkxg3_2;
	wire w_dff_B_WkuYxLfV3_2;
	wire w_dff_B_xXizeWOv0_2;
	wire w_dff_B_yogZZlHe7_2;
	wire w_dff_B_aggZKSxg1_2;
	wire w_dff_B_waK8gA0f1_2;
	wire w_dff_B_Sj0dESrj1_2;
	wire w_dff_B_j2A0JnKG7_2;
	wire w_dff_A_z3SpAsBY9_0;
	wire w_dff_A_h4vlfbh53_0;
	wire w_dff_A_iOmNIkL74_0;
	wire w_dff_A_kvCzikRY8_0;
	wire w_dff_A_JHX29h7K1_0;
	wire w_dff_B_TXVJFZdx9_2;
	wire w_dff_B_CdOhYngW4_2;
	wire w_dff_B_srtBb4KE9_2;
	wire w_dff_B_E5b1TohV2_2;
	wire w_dff_B_lBgeFI7Q9_2;
	wire w_dff_B_BpaOmRlf2_2;
	wire w_dff_B_RD9Kn9XY6_2;
	wire w_dff_B_TQK1Qdis4_2;
	wire w_dff_B_e1Jzoar65_2;
	wire w_dff_B_OvTt47YR2_2;
	wire w_dff_B_vxLDuHaH6_2;
	wire w_dff_B_8OCXqUup1_2;
	wire w_dff_B_tmfxmr9z1_2;
	wire w_dff_B_y9kN6HzJ7_2;
	wire w_dff_A_KrIZNGa98_0;
	wire w_dff_A_6YdQI9NW3_0;
	wire w_dff_A_FyMZjLpX9_0;
	wire w_dff_A_JzvDndrG6_0;
	wire w_dff_A_EYG2HVQB7_0;
	wire w_dff_A_zLTzD8dK1_0;
	wire w_dff_A_L5OcRHyo7_0;
	wire w_dff_A_UvEyALCO5_0;
	wire w_dff_A_p31a5J3T1_0;
	wire w_dff_B_wE7cgOgy0_1;
	wire w_dff_B_dcHqjuw37_0;
	wire w_dff_A_ouB13RQR3_0;
	wire w_dff_A_Xwi1K41p4_0;
	wire w_dff_A_sZGuDTaw4_0;
	wire w_dff_A_g0aJYL8b2_0;
	wire w_dff_A_FD32KFaa3_0;
	wire w_dff_A_SDE9snpP9_0;
	wire w_dff_A_eoze8ZM17_0;
	wire w_dff_A_7Hj6DsUx8_0;
	wire w_dff_A_0ywwW8Rq8_0;
	wire w_dff_A_rCoCTJoI5_0;
	wire w_dff_A_lzKY9Q687_0;
	wire w_dff_A_U7hcyydb5_0;
	wire w_dff_A_KhqhNqe23_0;
	wire w_dff_A_gBUzPPL46_0;
	wire w_dff_A_7gL6YP9d9_0;
	wire w_dff_A_eV8Lx7100_0;
	wire w_dff_A_wGbATrVY0_0;
	wire w_dff_A_vuYSf4N41_0;
	wire w_dff_A_YmlLkxql5_0;
	wire w_dff_A_R8I8AAsQ5_0;
	wire w_dff_A_gs1alE2z3_0;
	wire w_dff_A_r1CjFEzp9_0;
	wire w_dff_A_i36nh8WP6_0;
	wire w_dff_A_5OMAwbl14_0;
	wire w_dff_A_uE08Gi2I7_0;
	wire w_dff_A_LTfavr4G4_0;
	wire w_dff_A_5HCok42Z6_0;
	wire w_dff_A_h6tCBzkt0_0;
	wire w_dff_A_bojiUxdi7_0;
	wire w_dff_A_XBgUQi9j7_0;
	wire w_dff_A_k09LsJHf9_0;
	wire w_dff_A_cCbtaSj38_0;
	wire w_dff_A_SSwdXTSp0_0;
	wire w_dff_A_eg0q4qZl8_0;
	wire w_dff_A_jDkb1jpo9_0;
	wire w_dff_A_bL9BbCqS1_0;
	wire w_dff_A_C8SQykNj3_0;
	wire w_dff_A_leS70mqm1_0;
	wire w_dff_A_vVYN5yWg5_0;
	wire w_dff_A_S0Kla4y45_0;
	wire w_dff_A_pRex8mM39_0;
	wire w_dff_A_5xBYIMNA9_0;
	wire w_dff_A_4EjLBTNK1_0;
	wire w_dff_A_6ytp8to95_0;
	wire w_dff_A_cpPAdx7b7_0;
	wire w_dff_A_7VkWFbcc8_0;
	wire w_dff_A_Gnv9MqAk3_0;
	wire w_dff_A_KNZphkKF2_0;
	wire w_dff_A_NeCADXen4_0;
	wire w_dff_A_EdgOFw2R9_0;
	wire w_dff_A_uJTzLuYp8_0;
	wire w_dff_A_7jw3osed7_0;
	wire w_dff_A_0Wzhe35b9_0;
	wire w_dff_A_BqV46oBm3_0;
	wire w_dff_A_00MwMpVh8_0;
	wire w_dff_A_7LgXY2hr6_0;
	wire w_dff_A_bSa6l7RW6_1;
	wire w_dff_A_1Z6Vvesv4_1;
	wire w_dff_A_WeZ7fiuu0_1;
	wire w_dff_A_t0VpaKQb1_1;
	wire w_dff_A_DbMQ5Kkp5_1;
	wire w_dff_A_ZYuRGBwP4_1;
	wire w_dff_A_Z8JZutAt6_1;
	wire w_dff_A_YD7r77AC1_1;
	wire w_dff_A_R7E24HdF0_1;
	wire w_dff_A_bK8Fm5t88_1;
	wire w_dff_A_R4i0rjYk5_1;
	wire w_dff_A_VdhXtesf8_1;
	wire w_dff_A_tZOwrxrb9_1;
	wire w_dff_A_JrmgusHO7_1;
	wire w_dff_A_GGlQsEAT7_1;
	wire w_dff_A_BUrvsHja4_0;
	wire w_dff_A_OcWXa17Y1_0;
	wire w_dff_A_BG0cQmZT7_0;
	wire w_dff_A_aahn85jA5_0;
	wire w_dff_A_FEBuYrZW5_0;
	wire w_dff_A_FJ3P9wKY4_0;
	wire w_dff_A_JPLY7oM47_0;
	wire w_dff_A_R3oU3nPo4_0;
	wire w_dff_A_YYq9HJgt7_0;
	wire w_dff_A_1RlXYkc87_0;
	wire w_dff_A_QY9Ipw8V4_0;
	wire w_dff_A_dCJ7UnOL5_0;
	wire w_dff_A_75P5qZAy0_0;
	wire w_dff_A_WOxpT6gn6_0;
	wire w_dff_A_T2b1KUU77_0;
	wire w_dff_A_JCh726ST6_0;
	wire w_dff_A_UX51u8a68_0;
	wire w_dff_A_RfRUVYcJ2_0;
	wire w_dff_A_hOAqRrwN1_0;
	wire w_dff_A_kdlP9fvG4_0;
	wire w_dff_A_qhVJUMCa5_0;
	wire w_dff_A_lObfZyCr0_0;
	wire w_dff_A_yoQXhp4u4_0;
	wire w_dff_A_FfMTUyTq9_0;
	wire w_dff_A_F7lAHMbZ5_0;
	wire w_dff_A_KIT2oVfE1_0;
	wire w_dff_A_JKE684fO2_1;
	wire w_dff_A_rSt4TXBy7_1;
	wire w_dff_A_J6Hzp2vL6_1;
	wire w_dff_A_FeEW38KQ2_1;
	wire w_dff_A_n5vkYsBO7_1;
	wire w_dff_A_BS9zWpGs5_1;
	wire w_dff_A_pEoz1OBv7_1;
	wire w_dff_A_Fu2Vs6AE0_1;
	wire w_dff_A_bDYQFhP55_1;
	wire w_dff_A_2VPGrUa42_1;
	wire w_dff_A_suCVm50r3_1;
	wire w_dff_A_NIBZlJdj7_1;
	wire w_dff_A_3eQYcUjq8_1;
	wire w_dff_A_TYCpRd5N7_1;
	wire w_dff_A_WU7QAd689_1;
	wire w_dff_B_WK9KEog83_1;
	wire w_dff_B_grZPPI3n8_1;
	wire w_dff_B_02OmAt9I1_1;
	wire w_dff_B_2gCBTnE53_1;
	wire w_dff_B_a1GBCKnw2_1;
	wire w_dff_A_yhAsLHUh1_0;
	wire w_dff_A_j2SRVSWZ7_0;
	wire w_dff_A_oqPGa1lA9_0;
	wire w_dff_A_lcDkJHCH7_0;
	wire w_dff_A_fVVl20bv9_0;
	wire w_dff_A_SuT3eh386_0;
	wire w_dff_A_1nE3g42z8_0;
	wire w_dff_A_Eu7zaKVF5_0;
	wire w_dff_A_TcFdt9j46_0;
	wire w_dff_A_SdzTQ94W1_0;
	wire w_dff_A_hvrce2D24_0;
	wire w_dff_A_LfaykFyx0_0;
	wire w_dff_A_qVdxKEMW5_0;
	wire w_dff_A_SILs09bL3_0;
	wire w_dff_A_VkoZPS2k8_0;
	wire w_dff_A_SOsuPz846_0;
	wire w_dff_A_pHj5P0KO3_0;
	wire w_dff_A_Jodl1kHr9_0;
	wire w_dff_A_xv87rs4a3_0;
	wire w_dff_A_uKZwDS0q6_0;
	wire w_dff_A_jMIz7C8h3_1;
	wire w_dff_A_1IdMa42O0_1;
	wire w_dff_A_d0ncg8xV9_1;
	wire w_dff_A_LuDJ4YAm5_1;
	wire w_dff_A_hVDIqeOx4_1;
	wire w_dff_A_O21Mcrh82_1;
	wire w_dff_A_htWH4NPe7_1;
	wire w_dff_A_gMJmElbO0_1;
	wire w_dff_A_FXJaqxkI0_1;
	wire w_dff_A_xL0Lr6kL9_1;
	wire w_dff_A_hW2S2Ij85_1;
	wire w_dff_A_hb7DXibW9_1;
	wire w_dff_A_3T6DmOyr0_1;
	wire w_dff_A_X4d6cjKk8_1;
	wire w_dff_A_UYPDyGoW5_1;
	wire w_dff_A_qCQw9XKY0_0;
	wire w_dff_A_JtjTntn92_0;
	wire w_dff_A_YyI3E8jL9_0;
	wire w_dff_A_3vPeYXJb3_0;
	wire w_dff_A_7hDGEycb2_0;
	wire w_dff_A_YFNNmnBs3_0;
	wire w_dff_A_owZ2ONHU0_0;
	wire w_dff_A_rAyouTn90_0;
	wire w_dff_A_iRmxoRdw8_0;
	wire w_dff_A_DOevHaDy3_0;
	wire w_dff_A_nwdt9Yh96_0;
	wire w_dff_A_xQXq5qmb4_0;
	wire w_dff_A_dkjsXZhx2_0;
	wire w_dff_A_snA76Se24_0;
	wire w_dff_A_keiPrwBc3_0;
	wire w_dff_A_sqAm8OBq6_1;
	wire w_dff_B_cKZQaniF9_0;
	wire w_dff_B_k9o0KQBQ9_0;
	wire w_dff_B_DBInkPzr8_0;
	wire w_dff_B_h1tH2DaY1_0;
	wire w_dff_B_5iIZ9mmT2_0;
	wire w_dff_B_nDQgQQTX0_0;
	wire w_dff_A_rFP2X7Ot3_0;
	wire w_dff_A_PmNy3l3S7_0;
	wire w_dff_A_OGUA7Yfg2_0;
	wire w_dff_A_l1MvIUxs8_0;
	wire w_dff_A_uN1BM3qe9_0;
	wire w_dff_A_h2gruX1q6_0;
	wire w_dff_A_ZiyjYaVi2_0;
	wire w_dff_A_Qp59nlcQ9_0;
	wire w_dff_A_lMmH3DMV3_0;
	wire w_dff_A_vyzQ50Oe2_0;
	wire w_dff_A_Fdwi0p8x5_0;
	wire w_dff_A_z7sg22NV4_0;
	wire w_dff_B_ySC9SCAy7_2;
	wire w_dff_B_YAXGXf4H5_2;
	wire w_dff_B_gufyE0UY3_2;
	wire w_dff_B_0PpXGkgc6_2;
	wire w_dff_B_NNMPcNyT2_2;
	wire w_dff_B_VXg5wxDF6_2;
	wire w_dff_B_jxoo1BoU7_2;
	wire w_dff_A_iEsle1um8_0;
	wire w_dff_A_xtvhbAgz7_0;
	wire w_dff_A_gVfjfpbx0_0;
	wire w_dff_A_6tRiK9bI8_0;
	wire w_dff_A_utqPZN1V2_0;
	wire w_dff_A_KWQOLJYA8_0;
	wire w_dff_A_akBvbjZh2_0;
	wire w_dff_A_S4qFHhA64_0;
	wire w_dff_A_uSayjKQ25_0;
	wire w_dff_A_awbMIBy38_0;
	wire w_dff_A_Rm7ITCFT2_0;
	wire w_dff_A_n6exB7d33_0;
	wire w_dff_A_LVZ3uWFS9_0;
	wire w_dff_A_sJFh9Q6L0_0;
	wire w_dff_A_J5W4BsEu8_0;
	wire w_dff_A_EBA9LwQz5_0;
	wire w_dff_A_oBwHkyDm1_0;
	wire w_dff_A_95gPHotj2_0;
	wire w_dff_A_Am5UDLDt8_0;
	wire w_dff_A_Znhp1xeO2_0;
	wire w_dff_A_ib5ffShs1_0;
	wire w_dff_B_4DXugcxX7_1;
	wire w_dff_B_8kMUfIEC2_1;
	wire w_dff_B_GKh9iShf2_1;
	wire w_dff_B_8JOGPEdp3_1;
	wire w_dff_B_oOLbckUF0_1;
	wire w_dff_B_GWdQCYAe2_1;
	wire w_dff_B_aYB5X7vv5_1;
	wire w_dff_B_FGBvw4r15_1;
	wire w_dff_A_MDjoAOsQ5_0;
	wire w_dff_A_UMWgwLFp8_0;
	wire w_dff_A_pJjipAp56_0;
	wire w_dff_A_l28gomvj3_0;
	wire w_dff_A_MxVc0yor4_0;
	wire w_dff_A_0mAW1mXN5_0;
	wire w_dff_A_FXI92NMi3_0;
	wire w_dff_A_VjGIC8EB9_0;
	wire w_dff_A_OT3PLfim4_0;
	wire w_dff_A_tJ0B2s2A0_0;
	wire w_dff_A_pSc3zSWP5_0;
	wire w_dff_A_uBhXGZHN2_0;
	wire w_dff_A_pbXfR2hO7_0;
	wire w_dff_A_IPgss1P70_0;
	wire w_dff_A_G0aVskIx5_0;
	wire w_dff_A_WBxZLyLk5_0;
	wire w_dff_A_oZeyjCbM9_0;
	wire w_dff_A_om0J4qJz5_0;
	wire w_dff_B_pxpFaRoM0_2;
	wire w_dff_B_6LQsEQ8l5_2;
	wire w_dff_B_ArjxqDzQ1_2;
	wire w_dff_B_J165GFxe3_2;
	wire w_dff_B_oCTUljJ76_2;
	wire w_dff_B_J3FBaEnX3_2;
	wire w_dff_B_gy8RwmTF8_2;
	wire w_dff_A_Q2aHZ2AR8_0;
	wire w_dff_A_VQSOghpU7_0;
	wire w_dff_A_g50Uylmq0_0;
	wire w_dff_A_xkWLDgEz5_0;
	wire w_dff_A_aBGkLZjJ0_0;
	wire w_dff_A_q0TIis069_0;
	wire w_dff_A_W4ZZ7MPk2_0;
	wire w_dff_A_SgDemcaX1_0;
	wire w_dff_A_WbnqLGQM2_0;
	wire w_dff_A_lViaLDAp8_0;
	wire w_dff_A_Gz1Wo5EE2_0;
	wire w_dff_B_zVvm2PVc8_2;
	wire w_dff_B_VkmgccGa7_2;
	wire w_dff_B_SB6gz8lS6_2;
	wire w_dff_B_qa13KKWe8_2;
	wire w_dff_B_DPQ5NdHZ5_2;
	wire w_dff_B_02drxMj56_2;
	wire w_dff_B_MMpWv6I94_2;
	wire w_dff_B_MK2UGFni2_1;
	wire w_dff_B_zMVnDgUe7_0;
	wire w_dff_A_6xLzEwn20_0;
	wire w_dff_A_M1ji5M4c3_0;
	wire w_dff_A_zFp14LDU7_0;
	wire w_dff_A_B811KskL6_0;
	wire w_dff_A_xl9l1zNu8_0;
	wire w_dff_A_7P26Z4cx2_0;
	wire w_dff_A_MlnUQfpg3_0;
	wire w_dff_A_bZQqt8Il9_0;
	wire w_dff_A_Lqj3nDNG1_0;
	wire w_dff_A_B9Sli7pD7_0;
	wire w_dff_A_8SBupB3J0_0;
	wire w_dff_B_WGfXzdsH6_2;
	wire w_dff_B_sKb7Wm967_2;
	wire w_dff_B_CfkeuXU98_2;
	wire w_dff_B_bbl0mFmM6_2;
	wire w_dff_B_adIJcoHX8_2;
	wire w_dff_B_Yr9IKhTo4_2;
	wire w_dff_B_OfkeaqDE0_2;
	wire w_dff_A_PC08HT9Y0_0;
	wire w_dff_A_oo98AnT41_0;
	wire w_dff_A_anNQlfgt9_0;
	wire w_dff_A_WbEqaL9H4_0;
	wire w_dff_A_0PmFYCQ70_0;
	wire w_dff_A_I1ALeByX7_0;
	wire w_dff_A_05yPVrX25_0;
	wire w_dff_A_UOb6IWM88_0;
	wire w_dff_A_u7b3FYz57_0;
	wire w_dff_A_nCEn706y7_0;
	wire w_dff_A_HaGm7f1e2_0;
	wire w_dff_B_KANx3TDy8_2;
	wire w_dff_B_M3GEBIT96_2;
	wire w_dff_B_jVrQqdLO8_2;
	wire w_dff_B_zNnCM56m1_2;
	wire w_dff_B_VQbypCJw3_2;
	wire w_dff_B_GtN1Zagn7_2;
	wire w_dff_B_mr0pUf0l2_2;
	wire w_dff_B_HzekDwx63_1;
	wire w_dff_B_TVhoArzx1_1;
	wire w_dff_B_sWJOKgQ53_1;
	wire w_dff_B_tsOyWqJd5_1;
	wire w_dff_B_FgBqOXf90_1;
	wire w_dff_B_vbGj5EFR3_1;
	wire w_dff_B_XXQEqsMp7_1;
	wire w_dff_A_y0KjvieU4_0;
	wire w_dff_A_VCGhisw99_0;
	wire w_dff_A_aDHjhZMm0_0;
	wire w_dff_A_6b0YLsRo1_0;
	wire w_dff_A_nNo8Umco1_0;
	wire w_dff_A_zc5jePtT9_0;
	wire w_dff_A_7tOG5CNC9_0;
	wire w_dff_A_fmpfwvpc6_0;
	wire w_dff_A_6tR1FPKT0_0;
	wire w_dff_A_oFE9Iqmq0_0;
	wire w_dff_A_ACXJhbV32_0;
	wire w_dff_B_EXmU3giR8_2;
	wire w_dff_B_TmpCBnNW7_2;
	wire w_dff_B_Lf1dolqs8_2;
	wire w_dff_B_uZwg1S0t8_2;
	wire w_dff_B_XNUlyNiK9_2;
	wire w_dff_B_0QiJThQf3_2;
	wire w_dff_B_Ubacgs9I4_2;
	wire w_dff_A_cLZeErEF5_1;
	wire w_dff_A_YJwq2Zvq8_1;
	wire w_dff_A_p8rYGSep5_1;
	wire w_dff_A_qn3GcS4x5_1;
	wire w_dff_A_OE8rw2Yl7_1;
	wire w_dff_A_cQrg6etf2_1;
	wire w_dff_A_y3CrpwWQ9_1;
	wire w_dff_A_EPYoHhSd8_1;
	wire w_dff_A_zp8dRXpZ3_1;
	wire w_dff_A_c3n6djoO9_1;
	wire w_dff_A_jNKQiOuQ6_1;
	wire w_dff_A_W90tvkBv7_1;
	wire w_dff_A_4LIxEHvP0_1;
	wire w_dff_A_W4yJQrOz5_1;
	wire w_dff_A_3J53RKR44_1;
	wire w_dff_A_UVCWxBSj6_0;
	wire w_dff_A_uCLvcsCq4_0;
	wire w_dff_A_cAK5wk6x4_0;
	wire w_dff_A_jsGd9WQB7_0;
	wire w_dff_A_Vo0RVpcN6_0;
	wire w_dff_B_Gzw5Bwni2_2;
	wire w_dff_B_SCuL5UL08_2;
	wire w_dff_B_JEb5hJMN2_2;
	wire w_dff_B_7DjrZRPu5_2;
	wire w_dff_B_5tfaG7j98_2;
	wire w_dff_B_CXhyXXLJ0_2;
	wire w_dff_B_xvGXlgaU1_2;
	wire w_dff_B_7eXvcIPj8_2;
	wire w_dff_B_Z0lqTgGg8_2;
	wire w_dff_B_WK8PQyOj0_2;
	wire w_dff_B_bWlwbmt07_2;
	wire w_dff_B_HXvx0jsb8_2;
	wire w_dff_B_xnxbckoe6_2;
	wire w_dff_B_0peKtRbm5_2;
	wire w_dff_A_spVL2x6z2_0;
	wire w_dff_A_Ec7nvYtZ2_0;
	wire w_dff_A_ppdqxHB96_0;
	wire w_dff_A_eDkZ3wto8_0;
	wire w_dff_A_e1lXdjTl6_0;
	wire w_dff_A_q2quDH244_0;
	wire w_dff_A_L8wjvI4q6_0;
	wire w_dff_A_GA8xiqQi5_0;
	wire w_dff_A_rTaC778S1_0;
	wire w_dff_A_Sn06y3j33_0;
	wire w_dff_A_QPh8TyZT5_0;
	wire w_dff_A_mtt4fRf73_0;
	wire w_dff_A_9gw6BSS25_0;
	wire w_dff_A_ekmdJ2sK3_0;
	wire w_dff_A_YkuPxYKQ6_0;
	wire w_dff_A_bjcClbaR1_0;
	wire w_dff_A_traNO1Cg9_0;
	wire w_dff_A_k1h1GkCY5_0;
	wire w_dff_A_J94BjYdu6_0;
	wire w_dff_A_TsK5Cy9C6_0;
	wire w_dff_A_YwWieT7T5_0;
	wire w_dff_B_5CHZjteE6_1;
	wire w_dff_B_N5FF0fRm0_1;
	wire w_dff_A_sSdwTqtN8_0;
	wire w_dff_A_NC9vZe4y4_0;
	wire w_dff_A_dsRlYXKa0_0;
	wire w_dff_A_A0nPH3QQ1_0;
	wire w_dff_A_mMGUuize7_0;
	wire w_dff_A_hhjqW6sl3_0;
	wire w_dff_A_Apq31EEP4_0;
	wire w_dff_A_oV3Xayi37_0;
	wire w_dff_A_gfoqQjDK5_1;
	wire w_dff_A_CAMTCoCg0_1;
	wire w_dff_A_eMgtIPQW1_1;
	wire w_dff_A_K2l6bWI91_1;
	wire w_dff_A_N0irNl0C0_1;
	wire w_dff_A_tIbzckN32_1;
	wire w_dff_A_Wn8GzLHn2_1;
	wire w_dff_A_Zrqt1NQW4_1;
	wire w_dff_A_7xjnVOMN3_1;
	wire w_dff_A_9q5YkO6C6_1;
	wire w_dff_A_ZLJNJwzp0_1;
	wire w_dff_A_3ZHAhX0v1_1;
	wire w_dff_A_PMjxuwGC4_1;
	wire w_dff_A_AD4xuczk8_0;
	wire w_dff_A_UKfqoEhy9_0;
	wire w_dff_A_4oeBmz9q3_0;
	wire w_dff_A_hZXzDmHd0_0;
	wire w_dff_A_PyJBH4GW3_0;
	wire w_dff_A_8ZaN7ty78_0;
	wire w_dff_A_un6aqxhM5_0;
	wire w_dff_A_w1JLPekb1_0;
	wire w_dff_A_zkcMRtOO9_0;
	wire w_dff_A_xa1Nrk0b1_0;
	wire w_dff_A_hyZBNk011_0;
	wire w_dff_A_sCBP5Tky8_0;
	wire w_dff_A_7GdUoFLc2_0;
	wire w_dff_A_ZXVf5Nzp2_0;
	wire w_dff_A_mhJoslKp5_0;
	wire w_dff_A_F7oiPhA36_0;
	wire w_dff_A_5di2L4su3_0;
	wire w_dff_A_0Dd4OR8I1_0;
	wire w_dff_A_XzwxnOKp0_0;
	wire w_dff_A_FHuc58tC3_1;
	wire w_dff_A_vihw9c6K3_1;
	wire w_dff_A_0LU4okXJ3_1;
	wire w_dff_A_tslWGU1S1_1;
	wire w_dff_A_s4Ani3Gk5_1;
	wire w_dff_A_qZV14EGE8_1;
	wire w_dff_A_VfnyHQxD8_1;
	wire w_dff_A_kD7MLEVY8_1;
	wire w_dff_A_QDLByZa57_0;
	wire w_dff_A_BSgXFtMW4_0;
	wire w_dff_A_7CAeB6Wl0_0;
	wire w_dff_A_6gHQvYU45_0;
	wire w_dff_A_gi9H9yxK9_0;
	wire w_dff_A_SkawIwLd5_0;
	wire w_dff_A_R2gKMqU40_0;
	wire w_dff_A_JG3Heh8G4_0;
	wire w_dff_A_Y6eOtt9B1_0;
	wire w_dff_A_eF8DZN3L3_0;
	wire w_dff_A_6YCfdz0H4_0;
	wire w_dff_A_Yv0B43UV0_0;
	wire w_dff_A_KLS6JTbl0_0;
	wire w_dff_A_NH9UMk1G5_0;
	wire w_dff_A_hBBQgif57_0;
	wire w_dff_A_lmmQJEJx9_0;
	wire w_dff_A_p1brhldv6_0;
	wire w_dff_A_rNRGTngr3_0;
	wire w_dff_A_KrUqlXWO1_0;
	wire w_dff_A_lG4fbDm27_1;
	wire w_dff_A_AaH5f4xM2_1;
	wire w_dff_A_c59gx8zd7_1;
	wire w_dff_A_PnsqMdEa7_1;
	wire w_dff_A_8F9UQrgo7_1;
	wire w_dff_A_FHIs6XF06_1;
	wire w_dff_A_vsBdrI9I9_1;
	wire w_dff_A_L69zbemZ6_1;
	wire w_dff_A_yKJPnWMB9_1;
	wire w_dff_A_3ADpAWyi0_1;
	wire w_dff_A_oNCdNQzd2_1;
	wire w_dff_A_oZE6wGQp2_1;
	wire w_dff_A_L0rw6R8r0_1;
	wire w_dff_A_K1wdPRtT1_1;
	wire w_dff_A_JkqTa2vl0_1;
	wire w_dff_A_IiKOOlhv4_1;
	wire w_dff_A_QZk5PW4p2_0;
	wire w_dff_A_EO0z2ifm0_0;
	wire w_dff_A_uMldxBtI8_0;
	wire w_dff_A_arf4bEHa4_0;
	wire w_dff_A_JvWzoQW80_0;
	wire w_dff_B_F0JguZzJ5_2;
	wire w_dff_B_m3dJybvj1_2;
	wire w_dff_B_e7g7yZtB6_2;
	wire w_dff_B_asvh0jIs2_2;
	wire w_dff_B_vspyw1L60_2;
	wire w_dff_B_ulGm0nvv1_2;
	wire w_dff_B_WmSvZ7f01_2;
	wire w_dff_A_mzHtWNOf6_0;
	wire w_dff_A_nvkOzMxY0_0;
	wire w_dff_A_6KASFCUD7_0;
	wire w_dff_A_IYPetPUa0_0;
	wire w_dff_A_AM18Ao5n8_0;
	wire w_dff_A_hpFyGLSH4_0;
	wire w_dff_A_ntwLmnvx3_0;
	wire w_dff_A_tQwx1AAg8_0;
	wire w_dff_A_SN515lfE4_0;
	wire w_dff_A_qfXVdmSh4_0;
	wire w_dff_A_m4TbpFLn5_0;
	wire w_dff_A_ZY1y03VH3_0;
	wire w_dff_A_NKLuK1yq9_0;
	wire w_dff_B_je38FjIa0_1;
	wire w_dff_B_322Gjxrg7_0;
	wire w_dff_A_t04fUksS7_0;
	wire w_dff_A_o2uHKknx3_0;
	wire w_dff_A_qQTO3HbX5_0;
	wire w_dff_A_x4HZyByn8_0;
	wire w_dff_A_NczRzFiI9_0;
	wire w_dff_A_KIgzyAMf8_0;
	wire w_dff_B_dDO3Yzt54_1;
	wire w_dff_B_hw3qssex4_1;
	wire w_dff_B_NMbbV1YO5_1;
	wire w_dff_B_1lcgFhYH1_1;
	wire w_dff_B_ppddoFWA0_1;
	wire w_dff_B_bG9ClS3E6_1;
	wire w_dff_A_A5pOeaCf2_0;
	wire w_dff_A_pQNcgboV1_0;
	wire w_dff_A_ZOHyfuig1_0;
	wire w_dff_A_CNUZ71yK0_0;
	wire w_dff_A_rYrtoSBl9_0;
	wire w_dff_A_NNo3Tlci1_0;
	wire w_dff_A_h2Y9ZJzD2_0;
	wire w_dff_A_o85ay8Vw5_0;
	wire w_dff_A_wefd0r991_0;
	wire w_dff_A_Pts60yJD2_0;
	wire w_dff_A_mAKc8hN59_0;
	wire w_dff_A_fP25fRNS7_0;
	wire w_dff_A_l6NYPA6D1_0;
	wire w_dff_A_GfC7Bp2N2_1;
	wire w_dff_A_YVj5YIYD5_1;
	wire w_dff_A_NeWIEbjl9_1;
	wire w_dff_A_FgzBJMXg7_1;
	wire w_dff_A_yKc3S2P46_1;
	wire w_dff_A_0ckAmdGe6_1;
	wire w_dff_A_NU9uRoma3_1;
	wire w_dff_A_tqBIb0nN5_1;
	wire w_dff_A_dJOGWLWu1_0;
	wire w_dff_A_eeH93Aek3_0;
	wire w_dff_A_7vuqptF97_0;
	wire w_dff_A_6EfTsEgy0_0;
	wire w_dff_A_4Io0qKV22_0;
	wire w_dff_A_Hpp4eHyo1_0;
	wire w_dff_A_2MCyHMoD3_0;
	wire w_dff_A_zGokofoE6_0;
	wire w_dff_A_cj9R3qHv7_0;
	wire w_dff_A_bK50tSnb9_0;
	wire w_dff_A_bQ0gpzmo7_0;
	wire w_dff_A_tmxd6p482_0;
	wire w_dff_A_14R76Bzs5_0;
	wire w_dff_A_dUG3WhLy4_0;
	wire w_dff_A_kR7ACrt62_0;
	wire w_dff_A_yYWLwLlL7_0;
	wire w_dff_A_qXerH0iI8_0;
	wire w_dff_A_MoqWAgef6_0;
	wire w_dff_A_WxwdJJR06_0;
	wire w_dff_A_zwgpQTjc8_1;
	wire w_dff_A_pJ75RshI2_1;
	wire w_dff_A_EWEHM0VO0_1;
	wire w_dff_A_GHSz4eE30_1;
	wire w_dff_A_I7mCkaqp6_1;
	wire w_dff_A_UFtWY4da2_1;
	wire w_dff_A_gOOdI2ru9_1;
	wire w_dff_A_KVLsXlA68_1;
	wire w_dff_A_tSNHuSQF0_0;
	wire w_dff_A_73BhENhZ9_0;
	wire w_dff_A_evqLtQAD5_0;
	wire w_dff_A_e44ds8NR4_0;
	wire w_dff_A_sHaAYpWX2_0;
	wire w_dff_A_IB1VLXnM4_0;
	wire w_dff_A_Zwvh3ak07_1;
	wire w_dff_A_OVs73K2D2_1;
	wire w_dff_A_X67GF4lf1_1;
	wire w_dff_A_6sKgfne63_1;
	wire w_dff_A_fmbGG5rq0_1;
	wire w_dff_A_0h4uRpNu1_1;
	wire w_dff_A_xVbnUlJz2_0;
	wire w_dff_A_ZEWq0X020_0;
	wire w_dff_A_lrmNfJTA2_0;
	wire w_dff_A_6bJhwbl34_0;
	wire w_dff_A_HnTWAOgu1_0;
	wire w_dff_A_pEGBuJJz2_0;
	wire w_dff_A_rx6gk8z21_0;
	wire w_dff_A_lQ3WEhM69_0;
	wire w_dff_A_qGFULiEO4_1;
	wire w_dff_A_TAST8Uue5_1;
	wire w_dff_A_v2sdafcS2_1;
	wire w_dff_A_TNGkTsMo6_1;
	wire w_dff_A_ugHHWuQG4_1;
	wire w_dff_A_nlXoKio41_1;
	wire w_dff_A_s4aL91iV2_1;
	wire w_dff_A_t7842EW06_1;
	wire w_dff_A_vACIrymr1_1;
	wire w_dff_A_GI8wvvPZ6_1;
	wire w_dff_A_jynH119r0_1;
	wire w_dff_A_Na2a7yxM4_1;
	wire w_dff_A_SJ41GHkM6_1;
	wire w_dff_A_GZjtroyw6_0;
	wire w_dff_A_gBvb6wRA4_0;
	wire w_dff_A_UtLjcSU38_0;
	wire w_dff_A_SmABoodp9_0;
	wire w_dff_A_ZxKtvrd09_0;
	wire w_dff_A_LzcbsiGM9_0;
	wire w_dff_B_oFHjK9Vy2_1;
	wire w_dff_B_uy7Ipox02_1;
	wire w_dff_A_8vpAUUyx1_0;
	wire w_dff_A_rVlhmgEL9_0;
	wire w_dff_A_3ZJcno1i2_0;
	wire w_dff_A_blzEouPS7_0;
	wire w_dff_A_LdfUle2X1_0;
	wire w_dff_A_wktOnP1n7_0;
	wire w_dff_A_23rckZjR5_0;
	wire w_dff_A_DGM5D3ml6_0;
	wire w_dff_A_7tjp1Vyz8_0;
	wire w_dff_A_8L0BALgF9_0;
	wire w_dff_A_v1P0GAct8_0;
	wire w_dff_A_EQDqglJl5_0;
	wire w_dff_A_9dS6k8xR5_0;
	wire w_dff_A_4Ne3XgsQ3_0;
	wire w_dff_A_dfHDav1S5_0;
	wire w_dff_A_qsYE7pvN0_0;
	wire w_dff_A_k0qdTbHE4_0;
	wire w_dff_A_8wKpf4oa0_0;
	wire w_dff_A_lHlGuDJ27_0;
	wire w_dff_A_QnNiPzO00_0;
	wire w_dff_A_mDmrsqG29_0;
	wire w_dff_A_7Wkvu69p4_0;
	wire w_dff_A_wbAVqUWU0_0;
	wire w_dff_A_1RKxfJyf4_0;
	wire w_dff_A_nEZUbuOp2_0;
	wire w_dff_A_4azKf7PR2_0;
	wire w_dff_A_2z0aG76x2_0;
	wire w_dff_A_u22NVl2Z9_0;
	wire w_dff_A_OD6Iv26o4_0;
	wire w_dff_A_IToyDlht6_0;
	wire w_dff_A_Z8kEapOt6_0;
	wire w_dff_A_kp91eHvW8_0;
	wire w_dff_A_RvKDN4TZ1_0;
	wire w_dff_A_kkFSYdNl7_0;
	wire w_dff_A_Jq7fBqOF2_0;
	wire w_dff_A_s5VjoMFf9_0;
	wire w_dff_A_2EOcIFN52_0;
	wire w_dff_A_e2SsFd7f5_0;
	wire w_dff_A_jTcb8ZOl1_0;
	wire w_dff_A_YBtA6iDe4_0;
	wire w_dff_A_Xyt4i8y75_0;
	wire w_dff_A_fqhsjAks2_0;
	wire w_dff_A_KVWmTdjA8_0;
	wire w_dff_A_kpwza5SJ1_0;
	wire w_dff_A_ZOOuc7Ci6_0;
	wire w_dff_A_d1rrIRyd8_1;
	wire w_dff_A_yjLcObeY9_1;
	wire w_dff_A_hZcBfOUz8_1;
	wire w_dff_A_u8lwkm4s9_1;
	wire w_dff_A_hNl5FUOt7_1;
	wire w_dff_A_uAHsQf6v4_1;
	wire w_dff_A_SaVx8Hky1_1;
	wire w_dff_A_QBYLUvGz0_1;
	wire w_dff_A_LJPjatJ13_0;
	wire w_dff_A_eNBbkTo37_0;
	wire w_dff_A_JG7WXW0r9_0;
	wire w_dff_A_0TYQFC2b0_0;
	wire w_dff_A_wG5NK1E20_0;
	wire w_dff_B_ZMbGXRTG6_2;
	wire w_dff_B_iUlywCdM6_2;
	wire w_dff_B_7WNg8MN43_2;
	wire w_dff_B_WoxK1Frj3_2;
	wire w_dff_B_YN3ImGOS9_2;
	wire w_dff_B_hcPfypnS0_2;
	wire w_dff_B_44Sdazhr1_2;
	wire w_dff_A_2j5m2UZt0_0;
	wire w_dff_A_cS4Ucj8e9_0;
	wire w_dff_A_wKpgph9G5_0;
	wire w_dff_A_crOzn7BM3_0;
	wire w_dff_A_slbOCpSC2_0;
	wire w_dff_A_vpWnXkot6_0;
	wire w_dff_A_60jqn3kM3_0;
	wire w_dff_A_kYfuFxKh5_0;
	wire w_dff_A_xukxow173_0;
	wire w_dff_A_BiqpwgVM3_0;
	wire w_dff_A_onrBnMrm3_0;
	wire w_dff_A_yJgxfflI4_0;
	wire w_dff_A_PMAB5Jus3_0;
	wire w_dff_A_hj99hYJI9_1;
	wire w_dff_A_nZ1NBaOT1_1;
	wire w_dff_A_08BxUcFA2_1;
	wire w_dff_A_bAh2j8pu0_1;
	wire w_dff_A_OemU1Rgk7_1;
	wire w_dff_A_7w73e4kj4_1;
	wire w_dff_A_pvqPqSX98_1;
	wire w_dff_A_vx0g4e2i9_1;
	wire w_dff_A_V9ZXIcU37_0;
	wire w_dff_A_ZZpuQu4K5_0;
	wire w_dff_A_rEmuxZFv2_0;
	wire w_dff_A_ku63wcS59_0;
	wire w_dff_A_kS8OMkNR1_0;
	wire w_dff_A_4YgwA3ay8_0;
	wire w_dff_B_YfLa0vRk4_1;
	wire w_dff_B_PLZnYOXY2_1;
	wire w_dff_A_Bn9j67c56_0;
	wire w_dff_A_URLQiw6p2_0;
	wire w_dff_A_ZpXDOWGU0_0;
	wire w_dff_A_u0vo2dOR2_0;
	wire w_dff_A_cCb31esJ6_0;
	wire w_dff_A_cP0Dv3z61_0;
	wire w_dff_A_dB0buItk9_0;
	wire w_dff_A_6fK1W0AF1_0;
	wire w_dff_A_9QbkHJCp9_0;
	wire w_dff_A_AP9W7KQp1_0;
	wire w_dff_A_cqasrydz0_0;
	wire w_dff_A_bTT3B0U15_0;
	wire w_dff_A_RFTucnJE8_0;
	wire w_dff_A_hxkmzegh6_2;
	wire w_dff_A_60zA4AUF4_0;
	wire w_dff_A_UC10F9uH3_0;
	wire w_dff_A_vHH5HqRt0_0;
	wire w_dff_A_w6jy9CZx0_0;
	wire w_dff_A_vZIGNYMV3_0;
	wire w_dff_A_ywEvo4Ck3_0;
	wire w_dff_A_9NmUiCia9_1;
	wire w_dff_A_IQ8Cochu7_0;
	wire w_dff_A_NK2fXNy09_0;
	wire w_dff_A_7So5Ycq72_0;
	wire w_dff_A_njPNXPUC9_0;
	wire w_dff_A_sSX6e2yF5_0;
	wire w_dff_A_kHTV6ebl3_0;
	wire w_dff_A_UpOzULii4_0;
	wire w_dff_A_jw7dUq1X5_0;
	wire w_dff_A_YTJkIzR18_0;
	wire w_dff_A_VogTLJuw5_0;
	wire w_dff_A_CJvyBEDg6_0;
	wire w_dff_A_d3OR2Mk21_0;
	wire w_dff_A_k1PxBuxu6_0;
	wire w_dff_A_TsWW9uRX3_2;
	wire w_dff_A_xj5ZsRTa2_0;
	wire w_dff_A_lOImutZS3_0;
	wire w_dff_A_DUQ7apof3_0;
	wire w_dff_A_0xnoinQb8_0;
	wire w_dff_A_THf5n9Jx2_0;
	wire w_dff_A_EdeihZfi9_0;
	wire w_dff_A_TxQgQLVW1_1;
	wire w_dff_A_eMg2oYDa2_0;
	wire w_dff_A_yQOA5XwW1_0;
	wire w_dff_A_kfhgffsh9_0;
	wire w_dff_A_Wcuqr8lv2_0;
	wire w_dff_A_vlbRyPbg6_0;
	wire w_dff_A_ZT6PXlUK2_0;
	wire w_dff_A_SZMwVZMi4_0;
	wire w_dff_A_Eck8mjQ39_0;
	wire w_dff_A_9FKcUddG1_0;
	wire w_dff_A_UwJK3hhG1_0;
	wire w_dff_A_WFYITHG53_0;
	wire w_dff_A_bmvNrT030_0;
	wire w_dff_A_7PR6cJPe7_0;
	wire w_dff_A_CvptQvyC1_2;
	wire w_dff_A_xAE2yBz56_0;
	wire w_dff_A_AY3xOjbm3_0;
	wire w_dff_A_p90pGOqB0_0;
	wire w_dff_A_4WhCyM904_0;
	wire w_dff_A_TeTrPhwU8_0;
	wire w_dff_A_EWXebSuV4_0;
	wire w_dff_A_7wzDnKAk5_1;
	wire w_dff_A_NpKpEWfM1_0;
	wire w_dff_A_QA7CqL0h7_0;
	wire w_dff_A_dq4eVbYY9_0;
	wire w_dff_A_n9TvJP6c8_0;
	wire w_dff_A_MXoh95nB9_0;
	wire w_dff_A_exi9foQy0_0;
	wire w_dff_A_Vz87ur456_0;
	wire w_dff_A_RZyyhAbN0_0;
	wire w_dff_A_rsUOLE0u5_0;
	wire w_dff_A_5yNGVIWc8_0;
	wire w_dff_A_v3c8etSx2_0;
	wire w_dff_A_rQXTpGPf5_0;
	wire w_dff_A_SpSs8p8F2_0;
	wire w_dff_A_xnFEGC1b9_0;
	wire w_dff_A_DdSMJzfb4_0;
	wire w_dff_A_kUH8qIxF8_0;
	wire w_dff_A_fUx3ADay4_0;
	wire w_dff_A_bihIuxL99_0;
	wire w_dff_A_QkEetc6U8_0;
	wire w_dff_A_rRV5Ak2s0_0;
	wire w_dff_A_hwWOZ2qg2_0;
	wire w_dff_A_Su3yF4Rz7_0;
	wire w_dff_A_IvWgaa469_0;
	wire w_dff_A_fGlpwA8o1_0;
	wire w_dff_A_iuKWqCDK1_0;
	wire w_dff_A_KLo7KpIM1_1;
	wire w_dff_A_8wcGsKQx9_1;
	wire w_dff_A_dLuEru8m7_1;
	wire w_dff_A_LU6UkSEE9_1;
	wire w_dff_A_YTewSvrr7_1;
	wire w_dff_A_ebOJZH0D9_1;
	wire w_dff_A_VabbyFyh1_1;
	wire w_dff_A_tyvo7vN59_1;
	wire w_dff_A_tHuw6Rx03_1;
	wire w_dff_A_d4TMXWAz4_1;
	wire w_dff_A_7oq7v2Oe7_1;
	wire w_dff_A_Fdx6kx4w0_1;
	wire w_dff_A_k5GyKWBM9_1;
	wire w_dff_A_5M1BU1WW1_1;
	wire w_dff_A_wO1R5bKD2_1;
	wire w_dff_A_macC6PVE0_1;
	wire w_dff_A_nxnwmZGd1_1;
	wire w_dff_A_gqGFj5658_1;
	wire w_dff_A_c2IuFEPq5_1;
	wire w_dff_A_sgoJJj325_1;
	wire w_dff_A_MNKC2Dk62_1;
	wire w_dff_A_z0lqQNYb6_1;
	wire w_dff_A_3HySTJXS6_1;
	wire w_dff_A_BzjL9RWB2_2;
	wire w_dff_A_sc7G6lZl4_2;
	wire w_dff_A_uXNkjymG2_2;
	wire w_dff_A_vW0lIcPc0_2;
	wire w_dff_A_AdlW5dGu1_2;
	wire w_dff_A_zmE76EGO9_2;
	wire w_dff_A_67DigGNO6_2;
	wire w_dff_A_38dReck29_0;
	wire w_dff_A_IBe76F2N6_0;
	wire w_dff_A_LBJHi2yA5_0;
	wire w_dff_A_cSrLcZQX1_0;
	wire w_dff_A_k2PzWjou7_0;
	wire w_dff_A_wiqJSjdl0_0;
	wire w_dff_A_LPwi6se02_0;
	wire w_dff_A_SlVvIL6N8_0;
	wire w_dff_A_tr8YxxJk1_0;
	wire w_dff_A_7B3ZcoPL1_0;
	wire w_dff_A_ZosyvRvQ5_0;
	wire w_dff_A_2nEkXE7m1_0;
	wire w_dff_A_c3bypZTb4_0;
	wire w_dff_A_WQrXtqZC6_0;
	wire w_dff_A_eiXD1ttD4_2;
	wire w_dff_A_asXunjx04_0;
	wire w_dff_A_w17O8rej4_0;
	wire w_dff_A_HEQ2d7nX4_0;
	wire w_dff_A_QtG5Up7k5_0;
	wire w_dff_A_120NDMG06_0;
	wire w_dff_A_S3XhaID98_0;
	wire w_dff_A_PvHrowcr3_1;
	wire w_dff_A_MabweP9I7_0;
	wire w_dff_A_AyaUzMts8_0;
	wire w_dff_A_JoXecjJZ5_0;
	wire w_dff_A_YyEC9TrN8_0;
	wire w_dff_A_lbWiKf2i3_0;
	wire w_dff_A_zabAMT5S6_0;
	wire w_dff_A_rk0Ef1XQ4_0;
	wire w_dff_A_0btwrpQX6_0;
	wire w_dff_A_2cq9wl740_0;
	wire w_dff_A_gOSXiN7N7_0;
	wire w_dff_A_eqpzt1Md9_0;
	wire w_dff_A_vcgU7BgU1_0;
	wire w_dff_A_DdvFNv9v8_0;
	wire w_dff_A_algeuzM07_2;
	wire w_dff_A_eM82LuXd5_0;
	wire w_dff_A_TEopAfeD2_0;
	wire w_dff_A_xP0569zs8_0;
	wire w_dff_A_BeR21p7D0_0;
	wire w_dff_A_R35Guu1I3_0;
	wire w_dff_A_F4ECU3Yl1_0;
	wire w_dff_A_eBSbcp988_1;
	wire w_dff_A_Cnq4Y3gi7_0;
	wire w_dff_A_XgR4sJ4e5_0;
	wire w_dff_A_xdOwZ12M2_0;
	wire w_dff_A_coqpr0cX2_0;
	wire w_dff_A_PgZmOUSo7_0;
	wire w_dff_A_EnKYUt7C8_0;
	wire w_dff_A_wM6M0nWR5_0;
	wire w_dff_A_rGilqM3G7_0;
	wire w_dff_A_xTJRYaT95_0;
	wire w_dff_A_05zSM0OU7_0;
	wire w_dff_A_741alT7e3_0;
	wire w_dff_A_2Y9OrBWF5_0;
	wire w_dff_A_o1hoiLYi4_0;
	wire w_dff_A_RrmSmg7E5_2;
	wire w_dff_A_d9v12Sb57_0;
	wire w_dff_A_pljv0OjR5_0;
	wire w_dff_A_AEXiYSKt0_0;
	wire w_dff_A_kRJdjUmV6_0;
	wire w_dff_A_CBjgYnE14_1;
	wire w_dff_B_G0rNMgmM4_1;
	wire w_dff_A_oDpvd1uY3_0;
	wire w_dff_A_DkMJvmm33_0;
	wire w_dff_A_Eb2Yup1z2_0;
	wire w_dff_A_OhgP6H9w5_0;
	wire w_dff_A_pM4Ofpgb7_0;
	wire w_dff_A_05Ai5toY8_0;
	wire w_dff_A_vfRa9laY8_0;
	wire w_dff_A_8Cs8PhPB6_0;
	wire w_dff_A_hhT4Jx8v0_0;
	wire w_dff_A_c6qjtPui5_0;
	wire w_dff_A_22k1zkSY4_0;
	wire w_dff_A_eUT9tNhY0_0;
	wire w_dff_A_oft2wnYa5_0;
	wire w_dff_A_HoANK5OL6_1;
	wire w_dff_A_RxVzK2DL7_1;
	wire w_dff_A_4r98Dtqy5_1;
	wire w_dff_A_MnNDID1c5_1;
	wire w_dff_A_LkRv3Zqz5_1;
	wire w_dff_A_MBsFD3iu8_1;
	wire w_dff_A_nfpFi98I8_1;
	wire w_dff_A_eimXMdMg7_1;
	wire w_dff_A_OmXIee1c6_2;
	wire w_dff_A_zVidtoy64_0;
	wire w_dff_A_nU0cGZB42_0;
	wire w_dff_A_UDmQ15sN3_0;
	wire w_dff_A_Klm7WHf28_0;
	wire w_dff_A_hsvJpFM39_0;
	wire w_dff_A_UUJHy9aY1_0;
	wire w_dff_A_MD3643T96_0;
	wire w_dff_A_lGW3MMVj8_0;
	wire w_dff_A_erP4FJQC0_0;
	wire w_dff_A_5USV3o975_0;
	wire w_dff_A_8Lhq2fEL2_0;
	wire w_dff_A_qfLvVxkS1_0;
	wire w_dff_A_s0FqWuix1_0;
	wire w_dff_A_a6GzlPaf0_0;
	wire w_dff_A_JweVlmwy5_0;
	wire w_dff_A_bZLERgLv8_0;
	wire w_dff_A_FNl4fuHc6_0;
	wire w_dff_A_NkcHCvcA7_0;
	wire w_dff_A_G3IE0QgD5_0;
	wire w_dff_A_5YwW0yUb5_0;
	wire w_dff_A_3sOePMWg6_0;
	wire w_dff_A_F8UourEb8_0;
	wire w_dff_A_hnHpacdE9_1;
	wire w_dff_A_vQF300D38_1;
	wire w_dff_A_ejRr1Wao7_0;
	wire w_dff_A_aNUq5zKg5_0;
	wire w_dff_A_JqVg5MQE1_0;
	wire w_dff_A_XnQmRbMn9_0;
	wire w_dff_A_NgOxlcCU6_0;
	wire w_dff_A_GDlDXedd5_0;
	wire w_dff_A_VUpbDg4h6_0;
	wire w_dff_A_jI60A05b1_0;
	wire w_dff_A_KkAXZY2U1_0;
	wire w_dff_A_IPn330I22_0;
	wire w_dff_A_34aUbV7e2_0;
	wire w_dff_A_5F54Zuqg9_0;
	wire w_dff_A_LnLCDlFK8_0;
	wire w_dff_A_cVlkYZFJ1_0;
	wire w_dff_A_9xuIsWKI1_0;
	wire w_dff_A_oMk0Sfed2_0;
	wire w_dff_A_i8ye4iiK7_0;
	wire w_dff_A_eNw8VwPP9_0;
	wire w_dff_A_vttDMYKt0_0;
	wire w_dff_A_baacOaEL2_0;
	wire w_dff_A_qQJGeCWt3_1;
	wire w_dff_A_KlqEYryB7_0;
	wire w_dff_A_xdCspEKk1_0;
	wire w_dff_A_gLfy1ggQ9_0;
	wire w_dff_A_Ofb9KTck9_0;
	wire w_dff_A_fzonw2D54_0;
	wire w_dff_A_GRjqZ6qO6_0;
	wire w_dff_A_y8LDHsvB4_0;
	wire w_dff_A_rC33axc43_0;
	wire w_dff_A_gBKVROkF6_0;
	wire w_dff_A_BmxIRDOu0_0;
	wire w_dff_A_XVm4blHM1_0;
	wire w_dff_A_n5Eu2lKB6_0;
	wire w_dff_A_FJBVPdWa6_0;
	wire w_dff_A_VpmklDhU3_2;
	wire w_dff_A_FigXqfKP0_0;
	wire w_dff_A_lATlPhVO1_0;
	wire w_dff_A_7hPv0BTi1_0;
	wire w_dff_A_a949ANRM9_0;
	wire w_dff_A_ndvlgC9D9_0;
	wire w_dff_A_WuH62Us75_0;
	wire w_dff_A_EIdOR7m34_1;
	wire w_dff_A_7aVGoP6A3_0;
	jnot g000(.din(w_G102gat_0[1]),.dout(n43),.clk(gclk));
	jand g001(.dina(w_G108gat_0[2]),.dinb(w_n43_0[1]),.dout(n44),.clk(gclk));
	jnot g002(.din(w_G43gat_0[1]),.dout(n45),.clk(gclk));
	jor g003(.dina(w_n45_0[1]),.dinb(w_dff_B_G0rNMgmM4_1),.dout(n46),.clk(gclk));
	jnot g004(.din(w_n46_0[2]),.dout(n47),.clk(gclk));
	jor g005(.dina(w_n47_0[1]),.dinb(w_n44_0[1]),.dout(n48),.clk(gclk));
	jnot g006(.din(w_G63gat_0[2]),.dout(n49),.clk(gclk));
	jand g007(.dina(w_G69gat_0[2]),.dinb(w_n49_0[1]),.dout(n50),.clk(gclk));
	jnot g008(.din(w_G11gat_0[2]),.dout(n51),.clk(gclk));
	jand g009(.dina(w_G17gat_0[2]),.dinb(w_n51_0[1]),.dout(n52),.clk(gclk));
	jor g010(.dina(n52),.dinb(n50),.dout(n53),.clk(gclk));
	jnot g011(.din(w_G24gat_0[2]),.dout(n54),.clk(gclk));
	jand g012(.dina(w_G30gat_0[2]),.dinb(w_n54_0[1]),.dout(n55),.clk(gclk));
	jnot g013(.din(w_G50gat_0[1]),.dout(n56),.clk(gclk));
	jand g014(.dina(w_G56gat_1[1]),.dinb(n56),.dout(n57),.clk(gclk));
	jor g015(.dina(w_n57_0[1]),.dinb(n55),.dout(n58),.clk(gclk));
	jor g016(.dina(n58),.dinb(n53),.dout(n59),.clk(gclk));
	jnot g017(.din(w_G1gat_0[2]),.dout(n60),.clk(gclk));
	jand g018(.dina(w_G4gat_0[2]),.dinb(w_n60_0[1]),.dout(n61),.clk(gclk));
	jnot g019(.din(w_G89gat_0[2]),.dout(n62),.clk(gclk));
	jand g020(.dina(w_G95gat_0[2]),.dinb(w_n62_0[1]),.dout(n63),.clk(gclk));
	jnot g021(.din(w_G76gat_0[2]),.dout(n64),.clk(gclk));
	jand g022(.dina(w_G82gat_0[2]),.dinb(w_n64_0[1]),.dout(n65),.clk(gclk));
	jor g023(.dina(n65),.dinb(n63),.dout(n66),.clk(gclk));
	jor g024(.dina(n66),.dinb(w_dff_B_uy7Ipox02_1),.dout(n67),.clk(gclk));
	jor g025(.dina(n67),.dinb(n59),.dout(n68),.clk(gclk));
	jor g026(.dina(n68),.dinb(w_dff_B_oFHjK9Vy2_1),.dout(G223gat_fa_),.clk(gclk));
	jnot g027(.din(w_G21gat_0[2]),.dout(n70),.clk(gclk));
	jnot g028(.din(w_n44_0[0]),.dout(n71),.clk(gclk));
	jand g029(.dina(w_n46_0[1]),.dinb(n71),.dout(n72),.clk(gclk));
	jnot g030(.din(w_G69gat_0[1]),.dout(n73),.clk(gclk));
	jor g031(.dina(w_n73_0[1]),.dinb(w_G63gat_0[1]),.dout(n74),.clk(gclk));
	jnot g032(.din(w_G17gat_0[1]),.dout(n75),.clk(gclk));
	jor g033(.dina(w_n75_0[1]),.dinb(w_G11gat_0[1]),.dout(n76),.clk(gclk));
	jand g034(.dina(n76),.dinb(n74),.dout(n77),.clk(gclk));
	jnot g035(.din(w_G30gat_0[1]),.dout(n78),.clk(gclk));
	jor g036(.dina(w_n78_0[1]),.dinb(w_G24gat_0[1]),.dout(n79),.clk(gclk));
	jnot g037(.din(w_G56gat_1[0]),.dout(n80),.clk(gclk));
	jor g038(.dina(w_n80_0[1]),.dinb(w_G50gat_0[0]),.dout(n81),.clk(gclk));
	jand g039(.dina(w_n81_0[1]),.dinb(n79),.dout(n82),.clk(gclk));
	jand g040(.dina(n82),.dinb(n77),.dout(n83),.clk(gclk));
	jnot g041(.din(w_G4gat_0[1]),.dout(n84),.clk(gclk));
	jor g042(.dina(w_n84_0[1]),.dinb(w_G1gat_0[1]),.dout(n85),.clk(gclk));
	jnot g043(.din(w_G95gat_0[1]),.dout(n86),.clk(gclk));
	jor g044(.dina(w_n86_0[1]),.dinb(w_G89gat_0[1]),.dout(n87),.clk(gclk));
	jnot g045(.din(w_G82gat_0[1]),.dout(n88),.clk(gclk));
	jor g046(.dina(w_n88_0[1]),.dinb(w_G76gat_0[1]),.dout(n89),.clk(gclk));
	jand g047(.dina(n89),.dinb(n87),.dout(n90),.clk(gclk));
	jand g048(.dina(n90),.dinb(w_dff_B_PLZnYOXY2_1),.dout(n91),.clk(gclk));
	jand g049(.dina(n91),.dinb(n83),.dout(n92),.clk(gclk));
	jand g050(.dina(n92),.dinb(w_dff_B_YfLa0vRk4_1),.dout(n93),.clk(gclk));
	jor g051(.dina(w_n93_3[2]),.dinb(w_n51_0[0]),.dout(n94),.clk(gclk));
	jand g052(.dina(n94),.dinb(w_G17gat_0[0]),.dout(n95),.clk(gclk));
	jand g053(.dina(w_n95_0[1]),.dinb(w_n70_0[1]),.dout(n96),.clk(gclk));
	jnot g054(.din(w_G99gat_0[2]),.dout(n97),.clk(gclk));
	jor g055(.dina(w_n93_3[1]),.dinb(w_n62_0[0]),.dout(n98),.clk(gclk));
	jand g056(.dina(n98),.dinb(w_G95gat_0[0]),.dout(n99),.clk(gclk));
	jand g057(.dina(n99),.dinb(w_dff_B_XXQEqsMp7_1),.dout(n100),.clk(gclk));
	jor g058(.dina(n100),.dinb(n96),.dout(n101),.clk(gclk));
	jnot g059(.din(w_G73gat_0[2]),.dout(n102),.clk(gclk));
	jor g060(.dina(w_n93_3[0]),.dinb(w_n49_0[0]),.dout(n103),.clk(gclk));
	jand g061(.dina(n103),.dinb(w_G69gat_0[0]),.dout(n104),.clk(gclk));
	jand g062(.dina(w_n104_0[1]),.dinb(w_n102_0[1]),.dout(n105),.clk(gclk));
	jnot g063(.din(w_G34gat_0[2]),.dout(n106),.clk(gclk));
	jor g064(.dina(w_n93_2[2]),.dinb(w_n54_0[0]),.dout(n107),.clk(gclk));
	jand g065(.dina(n107),.dinb(w_G30gat_0[0]),.dout(n108),.clk(gclk));
	jand g066(.dina(w_n108_0[1]),.dinb(w_n106_0[1]),.dout(n109),.clk(gclk));
	jor g067(.dina(n109),.dinb(n105),.dout(n110),.clk(gclk));
	jnot g068(.din(w_G112gat_0[2]),.dout(n111),.clk(gclk));
	jor g069(.dina(w_n93_2[1]),.dinb(w_n43_0[0]),.dout(n112),.clk(gclk));
	jand g070(.dina(n112),.dinb(w_G108gat_0[1]),.dout(n113),.clk(gclk));
	jand g071(.dina(w_n113_0[1]),.dinb(w_n111_0[1]),.dout(n114),.clk(gclk));
	jor g072(.dina(w_dff_B_zMVnDgUe7_0),.dinb(n110),.dout(n115),.clk(gclk));
	jor g073(.dina(n115),.dinb(w_dff_B_MK2UGFni2_1),.dout(n116),.clk(gclk));
	jnot g074(.din(w_G60gat_0[1]),.dout(n117),.clk(gclk));
	jxor g075(.dina(w_n93_2[0]),.dinb(w_n57_0[0]),.dout(n118),.clk(gclk));
	jand g076(.dina(n118),.dinb(w_G56gat_0[2]),.dout(n119),.clk(gclk));
	jand g077(.dina(w_n119_0[2]),.dinb(w_n117_0[1]),.dout(n120),.clk(gclk));
	jnot g078(.din(w_G86gat_0[2]),.dout(n121),.clk(gclk));
	jor g079(.dina(w_n93_1[2]),.dinb(w_n64_0[0]),.dout(n122),.clk(gclk));
	jand g080(.dina(n122),.dinb(w_G82gat_0[0]),.dout(n123),.clk(gclk));
	jand g081(.dina(w_n123_0[1]),.dinb(w_n121_0[1]),.dout(n124),.clk(gclk));
	jnot g082(.din(w_G8gat_0[2]),.dout(n125),.clk(gclk));
	jor g083(.dina(w_n93_1[1]),.dinb(w_n60_0[0]),.dout(n126),.clk(gclk));
	jand g084(.dina(n126),.dinb(w_G4gat_0[0]),.dout(n127),.clk(gclk));
	jand g085(.dina(w_n127_0[1]),.dinb(w_n125_0[1]),.dout(n128),.clk(gclk));
	jnot g086(.din(w_G47gat_0[2]),.dout(n129),.clk(gclk));
	jor g087(.dina(w_n93_1[0]),.dinb(w_n47_0[0]),.dout(n130),.clk(gclk));
	jand g088(.dina(n130),.dinb(w_G43gat_0[0]),.dout(n131),.clk(gclk));
	jand g089(.dina(w_n131_0[2]),.dinb(w_dff_B_FGBvw4r15_1),.dout(n132),.clk(gclk));
	jor g090(.dina(n132),.dinb(n128),.dout(n133),.clk(gclk));
	jor g091(.dina(n133),.dinb(w_dff_B_4DXugcxX7_1),.dout(n134),.clk(gclk));
	jor g092(.dina(n134),.dinb(w_n120_0[1]),.dout(n135),.clk(gclk));
	jor g093(.dina(n135),.dinb(n116),.dout(G329gat_fa_),.clk(gclk));
	jand g094(.dina(w_G223gat_4),.dinb(w_G89gat_0[0]),.dout(n137),.clk(gclk));
	jor g095(.dina(n137),.dinb(w_n86_0[0]),.dout(n138),.clk(gclk));
	jand g096(.dina(w_G329gat_4),.dinb(w_G99gat_0[1]),.dout(n139),.clk(gclk));
	jor g097(.dina(n139),.dinb(w_n138_0[1]),.dout(n140),.clk(gclk));
	jor g098(.dina(w_n140_0[1]),.dinb(w_G105gat_0[1]),.dout(n141),.clk(gclk));
	jnot g099(.din(w_n141_0[1]),.dout(n142),.clk(gclk));
	jand g100(.dina(w_G329gat_3[2]),.dinb(w_G47gat_0[1]),.dout(n143),.clk(gclk));
	jnot g101(.din(n143),.dout(n144),.clk(gclk));
	jnot g102(.din(w_G53gat_0[1]),.dout(n145),.clk(gclk));
	jand g103(.dina(w_n131_0[1]),.dinb(w_n145_0[1]),.dout(n146),.clk(gclk));
	jand g104(.dina(w_dff_B_nDQgQQTX0_0),.dinb(w_n144_0[1]),.dout(n147),.clk(gclk));
	jor g105(.dina(w_n147_0[1]),.dinb(n142),.dout(n148),.clk(gclk));
	jnot g106(.din(w_G40gat_0[1]),.dout(n149),.clk(gclk));
	jand g107(.dina(w_G223gat_3[2]),.dinb(w_G11gat_0[0]),.dout(n150),.clk(gclk));
	jor g108(.dina(n150),.dinb(w_n75_0[0]),.dout(n151),.clk(gclk));
	jor g109(.dina(w_n151_0[1]),.dinb(w_G21gat_0[1]),.dout(n152),.clk(gclk));
	jor g110(.dina(w_n138_0[0]),.dinb(w_G99gat_0[0]),.dout(n153),.clk(gclk));
	jand g111(.dina(n153),.dinb(n152),.dout(n154),.clk(gclk));
	jand g112(.dina(w_G223gat_3[1]),.dinb(w_G63gat_0[0]),.dout(n155),.clk(gclk));
	jor g113(.dina(n155),.dinb(w_n73_0[0]),.dout(n156),.clk(gclk));
	jor g114(.dina(w_n156_0[1]),.dinb(w_G73gat_0[1]),.dout(n157),.clk(gclk));
	jand g115(.dina(w_G223gat_3[0]),.dinb(w_G24gat_0[0]),.dout(n158),.clk(gclk));
	jor g116(.dina(n158),.dinb(w_n78_0[0]),.dout(n159),.clk(gclk));
	jor g117(.dina(w_n159_0[1]),.dinb(w_G34gat_0[1]),.dout(n160),.clk(gclk));
	jand g118(.dina(n160),.dinb(n157),.dout(n161),.clk(gclk));
	jnot g119(.din(w_G108gat_0[0]),.dout(n162),.clk(gclk));
	jand g120(.dina(w_G223gat_2[2]),.dinb(w_G102gat_0[0]),.dout(n163),.clk(gclk));
	jor g121(.dina(n163),.dinb(w_dff_B_bG9ClS3E6_1),.dout(n164),.clk(gclk));
	jor g122(.dina(w_n164_0[1]),.dinb(w_G112gat_0[1]),.dout(n165),.clk(gclk));
	jand g123(.dina(w_dff_B_322Gjxrg7_0),.dinb(n161),.dout(n166),.clk(gclk));
	jand g124(.dina(n166),.dinb(w_dff_B_je38FjIa0_1),.dout(n167),.clk(gclk));
	jnot g125(.din(w_n120_0[0]),.dout(n168),.clk(gclk));
	jand g126(.dina(w_G223gat_2[1]),.dinb(w_G76gat_0[0]),.dout(n169),.clk(gclk));
	jor g127(.dina(n169),.dinb(w_n88_0[0]),.dout(n170),.clk(gclk));
	jor g128(.dina(w_n170_0[1]),.dinb(w_G86gat_0[1]),.dout(n171),.clk(gclk));
	jand g129(.dina(w_G223gat_2[0]),.dinb(w_G1gat_0[0]),.dout(n172),.clk(gclk));
	jor g130(.dina(n172),.dinb(w_n84_0[0]),.dout(n173),.clk(gclk));
	jor g131(.dina(w_n173_0[1]),.dinb(w_G8gat_0[1]),.dout(n174),.clk(gclk));
	jand g132(.dina(w_G223gat_1[2]),.dinb(w_n46_0[0]),.dout(n175),.clk(gclk));
	jor g133(.dina(n175),.dinb(w_n45_0[0]),.dout(n176),.clk(gclk));
	jor g134(.dina(n176),.dinb(w_G47gat_0[0]),.dout(n177),.clk(gclk));
	jand g135(.dina(n177),.dinb(n174),.dout(n178),.clk(gclk));
	jand g136(.dina(n178),.dinb(w_dff_B_N5FF0fRm0_1),.dout(n179),.clk(gclk));
	jand g137(.dina(n179),.dinb(w_dff_B_5CHZjteE6_1),.dout(n180),.clk(gclk));
	jand g138(.dina(n180),.dinb(n167),.dout(n181),.clk(gclk));
	jor g139(.dina(w_n181_2[2]),.dinb(w_n106_0[0]),.dout(n182),.clk(gclk));
	jand g140(.dina(n182),.dinb(w_n108_0[0]),.dout(n183),.clk(gclk));
	jand g141(.dina(w_n183_0[1]),.dinb(w_n149_0[1]),.dout(n184),.clk(gclk));
	jnot g142(.din(w_G66gat_0[2]),.dout(n185),.clk(gclk));
	jor g143(.dina(w_n181_2[1]),.dinb(w_n117_0[0]),.dout(n186),.clk(gclk));
	jand g144(.dina(n186),.dinb(w_n119_0[1]),.dout(n187),.clk(gclk));
	jand g145(.dina(n187),.dinb(w_n185_0[1]),.dout(n188),.clk(gclk));
	jor g146(.dina(n188),.dinb(n184),.dout(n189),.clk(gclk));
	jnot g147(.din(w_G14gat_0[2]),.dout(n190),.clk(gclk));
	jor g148(.dina(w_n181_2[0]),.dinb(w_n125_0[0]),.dout(n191),.clk(gclk));
	jand g149(.dina(n191),.dinb(w_n127_0[0]),.dout(n192),.clk(gclk));
	jand g150(.dina(n192),.dinb(w_dff_B_6hCX4gzq3_1),.dout(n193),.clk(gclk));
	jnot g151(.din(w_G92gat_0[2]),.dout(n194),.clk(gclk));
	jor g152(.dina(w_n181_1[2]),.dinb(w_n121_0[0]),.dout(n195),.clk(gclk));
	jand g153(.dina(n195),.dinb(w_n123_0[0]),.dout(n196),.clk(gclk));
	jand g154(.dina(n196),.dinb(w_dff_B_CSHAgvXc6_1),.dout(n197),.clk(gclk));
	jor g155(.dina(n197),.dinb(n193),.dout(n198),.clk(gclk));
	jor g156(.dina(n198),.dinb(n189),.dout(n199),.clk(gclk));
	jnot g157(.din(w_G79gat_0[1]),.dout(n200),.clk(gclk));
	jor g158(.dina(w_n181_1[1]),.dinb(w_n102_0[0]),.dout(n201),.clk(gclk));
	jand g159(.dina(n201),.dinb(w_n104_0[0]),.dout(n202),.clk(gclk));
	jand g160(.dina(w_n202_0[1]),.dinb(w_n200_0[1]),.dout(n203),.clk(gclk));
	jnot g161(.din(w_G115gat_0[1]),.dout(n204),.clk(gclk));
	jor g162(.dina(w_n181_1[0]),.dinb(w_n111_0[0]),.dout(n205),.clk(gclk));
	jand g163(.dina(n205),.dinb(w_n113_0[0]),.dout(n206),.clk(gclk));
	jand g164(.dina(w_n206_0[1]),.dinb(w_n204_0[1]),.dout(n207),.clk(gclk));
	jor g165(.dina(n207),.dinb(n203),.dout(n208),.clk(gclk));
	jnot g166(.din(w_G27gat_0[1]),.dout(n209),.clk(gclk));
	jor g167(.dina(w_n181_0[2]),.dinb(w_n70_0[0]),.dout(n210),.clk(gclk));
	jand g168(.dina(n210),.dinb(w_n95_0[0]),.dout(n211),.clk(gclk));
	jand g169(.dina(w_n211_0[1]),.dinb(w_n209_0[1]),.dout(n212),.clk(gclk));
	jor g170(.dina(w_dff_B_rbsEoq272_0),.dinb(n208),.dout(n213),.clk(gclk));
	jor g171(.dina(n213),.dinb(n199),.dout(n214),.clk(gclk));
	jor g172(.dina(n214),.dinb(w_dff_B_9IqYxDq65_1),.dout(G370gat_fa_),.clk(gclk));
	jnot g173(.din(w_n147_0[0]),.dout(n216),.clk(gclk));
	jand g174(.dina(n216),.dinb(w_n141_0[0]),.dout(n217),.clk(gclk));
	jand g175(.dina(w_G329gat_3[1]),.dinb(w_G34gat_0[0]),.dout(n218),.clk(gclk));
	jor g176(.dina(n218),.dinb(w_n159_0[0]),.dout(n219),.clk(gclk));
	jor g177(.dina(n219),.dinb(w_G40gat_0[0]),.dout(n220),.clk(gclk));
	jnot g178(.din(w_n119_0[0]),.dout(n221),.clk(gclk));
	jand g179(.dina(w_G329gat_3[0]),.dinb(w_G60gat_0[0]),.dout(n222),.clk(gclk));
	jor g180(.dina(w_n222_0[1]),.dinb(w_dff_B_a1GBCKnw2_1),.dout(n223),.clk(gclk));
	jor g181(.dina(n223),.dinb(w_G66gat_0[1]),.dout(n224),.clk(gclk));
	jand g182(.dina(n224),.dinb(n220),.dout(n225),.clk(gclk));
	jand g183(.dina(w_G329gat_2[2]),.dinb(w_G8gat_0[0]),.dout(n226),.clk(gclk));
	jor g184(.dina(n226),.dinb(w_n173_0[0]),.dout(n227),.clk(gclk));
	jor g185(.dina(w_n227_0[1]),.dinb(w_G14gat_0[1]),.dout(n228),.clk(gclk));
	jand g186(.dina(w_G329gat_2[1]),.dinb(w_G86gat_0[0]),.dout(n229),.clk(gclk));
	jor g187(.dina(n229),.dinb(w_n170_0[0]),.dout(n230),.clk(gclk));
	jor g188(.dina(w_n230_0[1]),.dinb(w_G92gat_0[1]),.dout(n231),.clk(gclk));
	jand g189(.dina(n231),.dinb(n228),.dout(n232),.clk(gclk));
	jand g190(.dina(n232),.dinb(n225),.dout(n233),.clk(gclk));
	jand g191(.dina(w_G329gat_2[0]),.dinb(w_G73gat_0[0]),.dout(n234),.clk(gclk));
	jor g192(.dina(n234),.dinb(w_n156_0[0]),.dout(n235),.clk(gclk));
	jor g193(.dina(n235),.dinb(w_G79gat_0[0]),.dout(n236),.clk(gclk));
	jand g194(.dina(w_G329gat_1[2]),.dinb(w_G112gat_0[0]),.dout(n237),.clk(gclk));
	jor g195(.dina(n237),.dinb(w_n164_0[0]),.dout(n238),.clk(gclk));
	jor g196(.dina(n238),.dinb(w_G115gat_0[0]),.dout(n239),.clk(gclk));
	jand g197(.dina(n239),.dinb(n236),.dout(n240),.clk(gclk));
	jand g198(.dina(w_G329gat_1[1]),.dinb(w_G21gat_0[0]),.dout(n241),.clk(gclk));
	jor g199(.dina(n241),.dinb(w_n151_0[0]),.dout(n242),.clk(gclk));
	jor g200(.dina(n242),.dinb(w_G27gat_0[0]),.dout(n243),.clk(gclk));
	jand g201(.dina(w_dff_B_dcHqjuw37_0),.dinb(n240),.dout(n244),.clk(gclk));
	jand g202(.dina(n244),.dinb(n233),.dout(n245),.clk(gclk));
	jand g203(.dina(n245),.dinb(w_dff_B_wE7cgOgy0_1),.dout(n246),.clk(gclk));
	jor g204(.dina(w_n246_2[2]),.dinb(w_n209_0[0]),.dout(n247),.clk(gclk));
	jand g205(.dina(n247),.dinb(w_n211_0[0]),.dout(n248),.clk(gclk));
	jor g206(.dina(w_n246_2[1]),.dinb(w_n149_0[0]),.dout(n249),.clk(gclk));
	jand g207(.dina(n249),.dinb(w_n183_0[0]),.dout(n250),.clk(gclk));
	jor g208(.dina(w_n250_0[1]),.dinb(w_n248_0[1]),.dout(n251),.clk(gclk));
	jor g209(.dina(w_n246_2[0]),.dinb(w_n145_0[0]),.dout(n252),.clk(gclk));
	jand g210(.dina(w_n144_0[0]),.dinb(w_n131_0[0]),.dout(n253),.clk(gclk));
	jand g211(.dina(w_n253_0[1]),.dinb(n252),.dout(n254),.clk(gclk));
	jor g212(.dina(w_n246_1[2]),.dinb(w_n185_0[0]),.dout(n255),.clk(gclk));
	jand g213(.dina(w_G223gat_1[1]),.dinb(w_n81_0[0]),.dout(n256),.clk(gclk));
	jor g214(.dina(w_n222_0[0]),.dinb(w_dff_B_JAMoUcrp2_1),.dout(n257),.clk(gclk));
	jnot g215(.din(w_n257_0[1]),.dout(n258),.clk(gclk));
	jand g216(.dina(w_dff_B_fn3dAsWe4_0),.dinb(n255),.dout(n259),.clk(gclk));
	jand g217(.dina(n259),.dinb(w_G56gat_0[1]),.dout(n260),.clk(gclk));
	jor g218(.dina(n260),.dinb(w_n254_0[1]),.dout(n261),.clk(gclk));
	jor g219(.dina(n261),.dinb(w_n251_0[1]),.dout(G430gat_fa_),.clk(gclk));
	jand g220(.dina(w_G370gat_1[1]),.dinb(w_G92gat_0[0]),.dout(n263),.clk(gclk));
	jor g221(.dina(n263),.dinb(w_n230_0[0]),.dout(n264),.clk(gclk));
	jnot g222(.din(w_n264_0[1]),.dout(n265),.clk(gclk));
	jnot g223(.din(w_n140_0[0]),.dout(n266),.clk(gclk));
	jnot g224(.din(w_G105gat_0[0]),.dout(n267),.clk(gclk));
	jor g225(.dina(w_n246_1[1]),.dinb(w_dff_B_m2yO53ZN7_1),.dout(n268),.clk(gclk));
	jand g226(.dina(n268),.dinb(w_dff_B_QU1k9qCM4_1),.dout(n269),.clk(gclk));
	jor g227(.dina(w_n246_1[0]),.dinb(w_n200_0[0]),.dout(n270),.clk(gclk));
	jand g228(.dina(n270),.dinb(w_n202_0[0]),.dout(n271),.clk(gclk));
	jor g229(.dina(w_n246_0[2]),.dinb(w_n204_0[0]),.dout(n272),.clk(gclk));
	jand g230(.dina(n272),.dinb(w_n206_0[0]),.dout(n273),.clk(gclk));
	jor g231(.dina(n273),.dinb(w_n271_0[1]),.dout(n274),.clk(gclk));
	jor g232(.dina(n274),.dinb(w_n269_0[1]),.dout(n275),.clk(gclk));
	jor g233(.dina(n275),.dinb(w_n265_0[1]),.dout(n276),.clk(gclk));
	jor g234(.dina(n276),.dinb(w_G430gat_0),.dout(n277),.clk(gclk));
	jand g235(.dina(w_G370gat_1[0]),.dinb(w_G14gat_0[0]),.dout(n278),.clk(gclk));
	jor g236(.dina(n278),.dinb(w_n227_0[0]),.dout(n279),.clk(gclk));
	jand g237(.dina(w_dff_B_LEU6kzmi3_0),.dinb(n277),.dout(G421gat),.clk(gclk));
	jnot g238(.din(w_n250_0[0]),.dout(n281),.clk(gclk));
	jand g239(.dina(w_G370gat_0[2]),.dinb(w_G53gat_0[0]),.dout(n282),.clk(gclk));
	jnot g240(.din(w_n253_0[0]),.dout(n283),.clk(gclk));
	jor g241(.dina(w_dff_B_yMwr3pGu7_0),.dinb(n282),.dout(n284),.clk(gclk));
	jand g242(.dina(w_G370gat_0[1]),.dinb(w_G66gat_0[0]),.dout(n285),.clk(gclk));
	jor g243(.dina(w_n257_0[0]),.dinb(n285),.dout(n286),.clk(gclk));
	jor g244(.dina(n286),.dinb(w_n80_0[0]),.dout(n287),.clk(gclk));
	jand g245(.dina(n287),.dinb(w_dff_B_MTftNmki7_1),.dout(n288),.clk(gclk));
	jand g246(.dina(w_n288_0[1]),.dinb(w_n281_0[1]),.dout(n289),.clk(gclk));
	jand g247(.dina(n289),.dinb(w_n271_0[0]),.dout(n290),.clk(gclk));
	jand g248(.dina(w_n265_0[0]),.dinb(w_n288_0[0]),.dout(n291),.clk(gclk));
	jor g249(.dina(n291),.dinb(w_n251_0[0]),.dout(n292),.clk(gclk));
	jor g250(.dina(n292),.dinb(w_n290_0[1]),.dout(G431gat),.clk(gclk));
	jand g251(.dina(w_n269_0[0]),.dinb(w_n264_0[0]),.dout(n294),.clk(gclk));
	jor g252(.dina(n294),.dinb(w_n254_0[0]),.dout(n295),.clk(gclk));
	jand g253(.dina(n295),.dinb(w_n281_0[0]),.dout(n296),.clk(gclk));
	jor g254(.dina(n296),.dinb(w_n248_0[0]),.dout(n297),.clk(gclk));
	jor g255(.dina(n297),.dinb(w_n290_0[0]),.dout(G432gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_EWXebSuV4_0),.doutb(w_dff_A_7wzDnKAk5_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_dff_A_7PR6cJPe7_0),.doutb(w_G4gat_0[1]),.doutc(w_dff_A_CvptQvyC1_2),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_XzwxnOKp0_0),.doutb(w_dff_A_kD7MLEVY8_1),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G11gat_0(.douta(w_dff_A_F4ECU3Yl1_0),.doutb(w_dff_A_eBSbcp988_1),.doutc(w_G11gat_0[2]),.din(G11gat));
	jspl3 jspl3_w_G14gat_0(.douta(w_dff_A_KIT2oVfE1_0),.doutb(w_dff_A_WU7QAd689_1),.doutc(w_G14gat_0[2]),.din(G14gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_dff_A_DdvFNv9v8_0),.doutb(w_G17gat_0[1]),.doutc(w_dff_A_algeuzM07_2),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_dff_A_ZOOuc7Ci6_0),.doutb(w_dff_A_QBYLUvGz0_1),.doutc(w_G21gat_0[2]),.din(G21gat));
	jspl3 jspl3_w_G24gat_0(.douta(w_dff_A_S3XhaID98_0),.doutb(w_dff_A_PvHrowcr3_1),.doutc(w_G24gat_0[2]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_dff_A_7gL6YP9d9_0),.doutb(w_G27gat_0[1]),.din(G27gat));
	jspl3 jspl3_w_G30gat_0(.douta(w_dff_A_WQrXtqZC6_0),.doutb(w_G30gat_0[1]),.doutc(w_dff_A_eiXD1ttD4_2),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_dff_A_WxwdJJR06_0),.doutb(w_dff_A_KVLsXlA68_1),.doutc(w_G34gat_0[2]),.din(G34gat));
	jspl jspl_w_G40gat_0(.douta(w_dff_A_keiPrwBc3_0),.doutb(w_G40gat_0[1]),.din(G40gat));
	jspl jspl_w_G43gat_0(.douta(w_dff_A_oft2wnYa5_0),.doutb(w_G43gat_0[1]),.din(G43gat));
	jspl3 jspl3_w_G47gat_0(.douta(w_dff_A_oV3Xayi37_0),.doutb(w_dff_A_PMjxuwGC4_1),.doutc(w_G47gat_0[2]),.din(G47gat));
	jspl jspl_w_G50gat_0(.douta(w_dff_A_38dReck29_0),.doutb(w_G50gat_0[1]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_dff_A_Znhp1xeO2_0),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_G56gat_0[0]),.doutb(w_dff_A_3HySTJXS6_1),.doutc(w_dff_A_67DigGNO6_2),.din(G56gat));
	jspl jspl_w_G56gat_1(.douta(w_G56gat_1[0]),.doutb(w_dff_A_KLo7KpIM1_1),.din(w_G56gat_0[0]));
	jspl jspl_w_G60gat_0(.douta(w_dff_A_NKLuK1yq9_0),.doutb(w_G60gat_0[1]),.din(G60gat));
	jspl3 jspl3_w_G63gat_0(.douta(w_dff_A_F8UourEb8_0),.doutb(w_dff_A_hnHpacdE9_1),.doutc(w_G63gat_0[2]),.din(G63gat));
	jspl3 jspl3_w_G66gat_0(.douta(w_dff_A_uKZwDS0q6_0),.doutb(w_dff_A_UYPDyGoW5_1),.doutc(w_G66gat_0[2]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_dff_A_o1hoiLYi4_0),.doutb(w_G69gat_0[1]),.doutc(w_dff_A_RrmSmg7E5_2),.din(G69gat));
	jspl3 jspl3_w_G73gat_0(.douta(w_dff_A_PMAB5Jus3_0),.doutb(w_dff_A_vx0g4e2i9_1),.doutc(w_G73gat_0[2]),.din(G73gat));
	jspl3 jspl3_w_G76gat_0(.douta(w_dff_A_ywEvo4Ck3_0),.doutb(w_dff_A_9NmUiCia9_1),.doutc(w_G76gat_0[2]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_dff_A_YkuPxYKQ6_0),.doutb(w_G79gat_0[1]),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_dff_A_RFTucnJE8_0),.doutb(w_G82gat_0[1]),.doutc(w_dff_A_hxkmzegh6_2),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_dff_A_KrUqlXWO1_0),.doutb(w_dff_A_L69zbemZ6_1),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G89gat_0(.douta(w_dff_A_EdeihZfi9_0),.doutb(w_dff_A_TxQgQLVW1_1),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_7LgXY2hr6_0),.doutb(w_dff_A_GGlQsEAT7_1),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_dff_A_k1PxBuxu6_0),.doutb(w_G95gat_0[1]),.doutc(w_dff_A_TsWW9uRX3_2),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_lQ3WEhM69_0),.doutb(w_dff_A_SJ41GHkM6_1),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl jspl_w_G102gat_0(.douta(w_dff_A_8Lhq2fEL2_0),.doutb(w_G102gat_0[1]),.din(G102gat));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_dff_A_3J53RKR44_1),.din(G105gat));
	jspl3 jspl3_w_G108gat_0(.douta(w_G108gat_0[0]),.doutb(w_dff_A_eimXMdMg7_1),.doutc(w_dff_A_OmXIee1c6_2),.din(G108gat));
	jspl3 jspl3_w_G112gat_0(.douta(w_dff_A_l6NYPA6D1_0),.doutb(w_dff_A_tqBIb0nN5_1),.doutc(w_G112gat_0[2]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_dff_A_XBgUQi9j7_0),.doutb(w_G115gat_0[1]),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(w_G223gat_3[2]),.din(w_G223gat_0[2]));
	jspl jspl_w_G223gat_4(.douta(w_G223gat_4),.doutb(w_dff_A_vQF300D38_1),.din(w_G223gat_1[0]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl jspl_w_G329gat_4(.douta(w_G329gat_4),.doutb(w_dff_A_qQJGeCWt3_1),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_dff_A_VpmklDhU3_2),.din(w_G370gat_0[0]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(w_dff_A_EIdOR7m34_1),.din(G430gat_fa_));
	jspl jspl_w_n43_0(.douta(w_dff_A_hsvJpFM39_0),.doutb(w_n43_0[1]),.din(n43));
	jspl jspl_w_n44_0(.douta(w_n44_0[0]),.doutb(w_dff_A_HoANK5OL6_1),.din(n44));
	jspl jspl_w_n45_0(.douta(w_dff_A_05Ai5toY8_0),.doutb(w_n45_0[1]),.din(n45));
	jspl3 jspl3_w_n46_0(.douta(w_dff_A_kRJdjUmV6_0),.doutb(w_dff_A_CBjgYnE14_1),.doutc(w_n46_0[2]),.din(n46));
	jspl jspl_w_n47_0(.douta(w_dff_A_kp91eHvW8_0),.doutb(w_n47_0[1]),.din(n47));
	jspl jspl_w_n49_0(.douta(w_dff_A_bZLERgLv8_0),.doutb(w_n49_0[1]),.din(n49));
	jspl jspl_w_n51_0(.douta(w_dff_A_OD6Iv26o4_0),.doutb(w_n51_0[1]),.din(n51));
	jspl jspl_w_n54_0(.douta(w_dff_A_1RKxfJyf4_0),.doutb(w_n54_0[1]),.din(n54));
	jspl jspl_w_n57_0(.douta(w_dff_A_lHlGuDJ27_0),.doutb(w_n57_0[1]),.din(n57));
	jspl jspl_w_n60_0(.douta(w_dff_A_dfHDav1S5_0),.doutb(w_n60_0[1]),.din(n60));
	jspl jspl_w_n62_0(.douta(w_dff_A_8L0BALgF9_0),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n64_0(.douta(w_dff_A_LdfUle2X1_0),.doutb(w_n64_0[1]),.din(n64));
	jspl jspl_w_n70_0(.douta(w_dff_A_ACXJhbV32_0),.doutb(w_n70_0[1]),.din(w_dff_B_Ubacgs9I4_2));
	jspl jspl_w_n73_0(.douta(w_dff_A_EnKYUt7C8_0),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n75_0(.douta(w_dff_A_zabAMT5S6_0),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n78_0(.douta(w_dff_A_LPwi6se02_0),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n80_0(.douta(w_dff_A_iuKWqCDK1_0),.doutb(w_n80_0[1]),.din(n80));
	jspl jspl_w_n81_0(.douta(w_dff_A_n9TvJP6c8_0),.doutb(w_n81_0[1]),.din(n81));
	jspl jspl_w_n84_0(.douta(w_dff_A_ZT6PXlUK2_0),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_dff_A_kHTV6ebl3_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_dff_A_cP0Dv3z61_0),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl3 jspl3_w_n93_1(.douta(w_n93_1[0]),.doutb(w_n93_1[1]),.doutc(w_n93_1[2]),.din(w_n93_0[0]));
	jspl3 jspl3_w_n93_2(.douta(w_n93_2[0]),.doutb(w_n93_2[1]),.doutc(w_n93_2[2]),.din(w_n93_0[1]));
	jspl3 jspl3_w_n93_3(.douta(w_n93_3[0]),.doutb(w_n93_3[1]),.doutc(w_n93_3[2]),.din(w_n93_0[2]));
	jspl jspl_w_n95_0(.douta(w_dff_A_zc5jePtT9_0),.doutb(w_n95_0[1]),.din(n95));
	jspl jspl_w_n102_0(.douta(w_dff_A_wG5NK1E20_0),.doutb(w_n102_0[1]),.din(w_dff_B_44Sdazhr1_2));
	jspl jspl_w_n104_0(.douta(w_dff_A_4YgwA3ay8_0),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n106_0(.douta(w_dff_A_HaGm7f1e2_0),.doutb(w_n106_0[1]),.din(w_dff_B_mr0pUf0l2_2));
	jspl jspl_w_n108_0(.douta(w_dff_A_I1ALeByX7_0),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n111_0(.douta(w_dff_A_8SBupB3J0_0),.doutb(w_n111_0[1]),.din(w_dff_B_OfkeaqDE0_2));
	jspl jspl_w_n113_0(.douta(w_dff_A_7P26Z4cx2_0),.doutb(w_n113_0[1]),.din(n113));
	jspl jspl_w_n117_0(.douta(w_dff_A_JvWzoQW80_0),.doutb(w_n117_0[1]),.din(w_dff_B_WmSvZ7f01_2));
	jspl3 jspl3_w_n119_0(.douta(w_n119_0[0]),.doutb(w_dff_A_IiKOOlhv4_1),.doutc(w_n119_0[2]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_dff_A_3ADpAWyi0_1),.din(n120));
	jspl jspl_w_n121_0(.douta(w_dff_A_Gz1Wo5EE2_0),.doutb(w_n121_0[1]),.din(w_dff_B_MMpWv6I94_2));
	jspl jspl_w_n123_0(.douta(w_dff_A_q0TIis069_0),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n125_0(.douta(w_dff_A_om0J4qJz5_0),.doutb(w_n125_0[1]),.din(w_dff_B_gy8RwmTF8_2));
	jspl jspl_w_n127_0(.douta(w_dff_A_pbXfR2hO7_0),.doutb(w_n127_0[1]),.din(n127));
	jspl3 jspl3_w_n131_0(.douta(w_dff_A_FXI92NMi3_0),.doutb(w_n131_0[1]),.doutc(w_n131_0[2]),.din(n131));
	jspl jspl_w_n138_0(.douta(w_n138_0[0]),.doutb(w_dff_A_0h4uRpNu1_1),.din(n138));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n141_0(.douta(w_dff_A_ib5ffShs1_0),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(n144));
	jspl jspl_w_n145_0(.douta(w_dff_A_z7sg22NV4_0),.doutb(w_n145_0[1]),.din(w_dff_B_jxoo1BoU7_2));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_dff_A_sqAm8OBq6_1),.din(n147));
	jspl jspl_w_n149_0(.douta(w_dff_A_JHX29h7K1_0),.doutb(w_n149_0[1]),.din(w_dff_B_y9kN6HzJ7_2));
	jspl jspl_w_n151_0(.douta(w_dff_A_LzcbsiGM9_0),.doutb(w_n151_0[1]),.din(n151));
	jspl jspl_w_n156_0(.douta(w_dff_A_IB1VLXnM4_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n159_0(.douta(w_dff_A_Hpp4eHyo1_0),.doutb(w_n159_0[1]),.din(n159));
	jspl jspl_w_n164_0(.douta(w_dff_A_KIgzyAMf8_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n170_0(.douta(w_dff_A_SkawIwLd5_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n173_0(.douta(w_dff_A_8ZaN7ty78_0),.doutb(w_n173_0[1]),.din(n173));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n181_2(.douta(w_n181_2[0]),.doutb(w_n181_2[1]),.doutc(w_n181_2[2]),.din(w_n181_0[1]));
	jspl jspl_w_n183_0(.douta(w_dff_A_zLTzD8dK1_0),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n185_0(.douta(w_dff_A_LoqwA0X89_0),.doutb(w_n185_0[1]),.din(w_dff_B_Sj0dESrj1_2));
	jspl jspl_w_n200_0(.douta(w_dff_A_Vo0RVpcN6_0),.doutb(w_n200_0[1]),.din(w_dff_B_0peKtRbm5_2));
	jspl jspl_w_n202_0(.douta(w_dff_A_YwWieT7T5_0),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n204_0(.douta(w_dff_A_zs8YKF2e3_0),.doutb(w_n204_0[1]),.din(w_dff_B_i1S2LK491_2));
	jspl jspl_w_n206_0(.douta(w_dff_A_QICiSLGL9_0),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n209_0(.douta(w_dff_A_6I3Xz4tf1_0),.doutb(w_n209_0[1]),.din(w_dff_B_meL2PgNV6_2));
	jspl jspl_w_n211_0(.douta(w_dff_A_iNsHqmcB9_0),.doutb(w_n211_0[1]),.din(n211));
	jspl jspl_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n227_0(.douta(w_dff_A_FJ3P9wKY4_0),.doutb(w_n227_0[1]),.din(n227));
	jspl jspl_w_n230_0(.douta(w_dff_A_bL9BbCqS1_0),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl3 jspl3_w_n246_1(.douta(w_n246_1[0]),.doutb(w_n246_1[1]),.doutc(w_n246_1[2]),.din(w_n246_0[0]));
	jspl3 jspl3_w_n246_2(.douta(w_n246_2[0]),.doutb(w_n246_2[1]),.doutc(w_n246_2[2]),.din(w_n246_0[1]));
	jspl jspl_w_n248_0(.douta(w_dff_A_IoJGLttf4_0),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_dff_A_CGsl3pof0_0),.doutb(w_n251_0[1]),.din(w_dff_B_26IILePm0_2));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_dff_A_USMqUlZT0_1),.din(n253));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(w_dff_B_SFkrwljf0_2));
	jspl jspl_w_n257_0(.douta(w_dff_A_XTA5sNUR6_0),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(w_dff_B_gm120Oud6_2));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_dff_A_q7Tu8nTb4_1),.din(n269));
	jspl jspl_w_n271_0(.douta(w_dff_A_p31a5J3T1_0),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.din(w_dff_B_j2A0JnKG7_2));
	jspl jspl_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.din(n288));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(n290));
	jdff dff_B_nNqmRsp24_0(.din(n279),.dout(w_dff_B_nNqmRsp24_0),.clk(gclk));
	jdff dff_B_DPvU5Quz3_0(.din(w_dff_B_nNqmRsp24_0),.dout(w_dff_B_DPvU5Quz3_0),.clk(gclk));
	jdff dff_B_y6Q9Vrdi5_0(.din(w_dff_B_DPvU5Quz3_0),.dout(w_dff_B_y6Q9Vrdi5_0),.clk(gclk));
	jdff dff_B_LEU6kzmi3_0(.din(w_dff_B_y6Q9Vrdi5_0),.dout(w_dff_B_LEU6kzmi3_0),.clk(gclk));
	jdff dff_B_MbNAgu3c0_0(.din(n258),.dout(w_dff_B_MbNAgu3c0_0),.clk(gclk));
	jdff dff_B_iPSNwcO46_0(.din(w_dff_B_MbNAgu3c0_0),.dout(w_dff_B_iPSNwcO46_0),.clk(gclk));
	jdff dff_B_hlDujAZe1_0(.din(w_dff_B_iPSNwcO46_0),.dout(w_dff_B_hlDujAZe1_0),.clk(gclk));
	jdff dff_B_S8fN2eSL6_0(.din(w_dff_B_hlDujAZe1_0),.dout(w_dff_B_S8fN2eSL6_0),.clk(gclk));
	jdff dff_B_fn3dAsWe4_0(.din(w_dff_B_S8fN2eSL6_0),.dout(w_dff_B_fn3dAsWe4_0),.clk(gclk));
	jdff dff_B_gm120Oud6_2(.din(n265),.dout(w_dff_B_gm120Oud6_2),.clk(gclk));
	jdff dff_A_CGsl3pof0_0(.dout(w_n251_0[0]),.din(w_dff_A_CGsl3pof0_0),.clk(gclk));
	jdff dff_B_26IILePm0_2(.din(n251),.dout(w_dff_B_26IILePm0_2),.clk(gclk));
	jdff dff_A_q7Tu8nTb4_1(.dout(w_n269_0[1]),.din(w_dff_A_q7Tu8nTb4_1),.clk(gclk));
	jdff dff_B_NKNZqV8m2_1(.din(n266),.dout(w_dff_B_NKNZqV8m2_1),.clk(gclk));
	jdff dff_B_JcokKGtz9_1(.din(w_dff_B_NKNZqV8m2_1),.dout(w_dff_B_JcokKGtz9_1),.clk(gclk));
	jdff dff_B_GlRJCYin5_1(.din(w_dff_B_JcokKGtz9_1),.dout(w_dff_B_GlRJCYin5_1),.clk(gclk));
	jdff dff_B_1wOjlkoT3_1(.din(w_dff_B_GlRJCYin5_1),.dout(w_dff_B_1wOjlkoT3_1),.clk(gclk));
	jdff dff_B_QU1k9qCM4_1(.din(w_dff_B_1wOjlkoT3_1),.dout(w_dff_B_QU1k9qCM4_1),.clk(gclk));
	jdff dff_B_HXxjs9fd1_1(.din(n267),.dout(w_dff_B_HXxjs9fd1_1),.clk(gclk));
	jdff dff_B_0UYRfxd18_1(.din(w_dff_B_HXxjs9fd1_1),.dout(w_dff_B_0UYRfxd18_1),.clk(gclk));
	jdff dff_B_MQvrzUcL1_1(.din(w_dff_B_0UYRfxd18_1),.dout(w_dff_B_MQvrzUcL1_1),.clk(gclk));
	jdff dff_B_gYK1ymEv1_1(.din(w_dff_B_MQvrzUcL1_1),.dout(w_dff_B_gYK1ymEv1_1),.clk(gclk));
	jdff dff_B_iDH25Nws7_1(.din(w_dff_B_gYK1ymEv1_1),.dout(w_dff_B_iDH25Nws7_1),.clk(gclk));
	jdff dff_B_M4gRjj490_1(.din(w_dff_B_iDH25Nws7_1),.dout(w_dff_B_M4gRjj490_1),.clk(gclk));
	jdff dff_B_Pd4PdKN34_1(.din(w_dff_B_M4gRjj490_1),.dout(w_dff_B_Pd4PdKN34_1),.clk(gclk));
	jdff dff_B_11ePEZrX5_1(.din(w_dff_B_Pd4PdKN34_1),.dout(w_dff_B_11ePEZrX5_1),.clk(gclk));
	jdff dff_B_PmLR5C9Z9_1(.din(w_dff_B_11ePEZrX5_1),.dout(w_dff_B_PmLR5C9Z9_1),.clk(gclk));
	jdff dff_B_HzFvrYs33_1(.din(w_dff_B_PmLR5C9Z9_1),.dout(w_dff_B_HzFvrYs33_1),.clk(gclk));
	jdff dff_B_rNUSAL3o8_1(.din(w_dff_B_HzFvrYs33_1),.dout(w_dff_B_rNUSAL3o8_1),.clk(gclk));
	jdff dff_B_ek5lLYeP0_1(.din(w_dff_B_rNUSAL3o8_1),.dout(w_dff_B_ek5lLYeP0_1),.clk(gclk));
	jdff dff_B_u2pTCMcv7_1(.din(w_dff_B_ek5lLYeP0_1),.dout(w_dff_B_u2pTCMcv7_1),.clk(gclk));
	jdff dff_B_Jo5vL0Ub8_1(.din(w_dff_B_u2pTCMcv7_1),.dout(w_dff_B_Jo5vL0Ub8_1),.clk(gclk));
	jdff dff_B_vHqkHYop4_1(.din(w_dff_B_Jo5vL0Ub8_1),.dout(w_dff_B_vHqkHYop4_1),.clk(gclk));
	jdff dff_B_3e5MOXWc9_1(.din(w_dff_B_vHqkHYop4_1),.dout(w_dff_B_3e5MOXWc9_1),.clk(gclk));
	jdff dff_B_3vLTyasL5_1(.din(w_dff_B_3e5MOXWc9_1),.dout(w_dff_B_3vLTyasL5_1),.clk(gclk));
	jdff dff_B_RuN9JMrB1_1(.din(w_dff_B_3vLTyasL5_1),.dout(w_dff_B_RuN9JMrB1_1),.clk(gclk));
	jdff dff_B_m2yO53ZN7_1(.din(w_dff_B_RuN9JMrB1_1),.dout(w_dff_B_m2yO53ZN7_1),.clk(gclk));
	jdff dff_B_SFkrwljf0_2(.din(n254),.dout(w_dff_B_SFkrwljf0_2),.clk(gclk));
	jdff dff_A_JFZSl3S94_0(.dout(w_n248_0[0]),.din(w_dff_A_JFZSl3S94_0),.clk(gclk));
	jdff dff_A_StAWxQvm3_0(.dout(w_dff_A_JFZSl3S94_0),.din(w_dff_A_StAWxQvm3_0),.clk(gclk));
	jdff dff_A_IoJGLttf4_0(.dout(w_dff_A_StAWxQvm3_0),.din(w_dff_A_IoJGLttf4_0),.clk(gclk));
	jdff dff_B_MTftNmki7_1(.din(n284),.dout(w_dff_B_MTftNmki7_1),.clk(gclk));
	jdff dff_A_M7m9KzrF2_0(.dout(w_n257_0[0]),.din(w_dff_A_M7m9KzrF2_0),.clk(gclk));
	jdff dff_A_eeWmzvKG2_0(.dout(w_dff_A_M7m9KzrF2_0),.din(w_dff_A_eeWmzvKG2_0),.clk(gclk));
	jdff dff_A_tSs5Q0CR8_0(.dout(w_dff_A_eeWmzvKG2_0),.din(w_dff_A_tSs5Q0CR8_0),.clk(gclk));
	jdff dff_A_gitFoMzA3_0(.dout(w_dff_A_tSs5Q0CR8_0),.din(w_dff_A_gitFoMzA3_0),.clk(gclk));
	jdff dff_A_KGuYjPc29_0(.dout(w_dff_A_gitFoMzA3_0),.din(w_dff_A_KGuYjPc29_0),.clk(gclk));
	jdff dff_A_XTA5sNUR6_0(.dout(w_dff_A_KGuYjPc29_0),.din(w_dff_A_XTA5sNUR6_0),.clk(gclk));
	jdff dff_B_hTfrpH2X9_1(.din(n256),.dout(w_dff_B_hTfrpH2X9_1),.clk(gclk));
	jdff dff_B_Hni7MjoT2_1(.din(w_dff_B_hTfrpH2X9_1),.dout(w_dff_B_Hni7MjoT2_1),.clk(gclk));
	jdff dff_B_s6XJgI8S8_1(.din(w_dff_B_Hni7MjoT2_1),.dout(w_dff_B_s6XJgI8S8_1),.clk(gclk));
	jdff dff_B_OgWkF7Jl6_1(.din(w_dff_B_s6XJgI8S8_1),.dout(w_dff_B_OgWkF7Jl6_1),.clk(gclk));
	jdff dff_B_zEtFVFdN7_1(.din(w_dff_B_OgWkF7Jl6_1),.dout(w_dff_B_zEtFVFdN7_1),.clk(gclk));
	jdff dff_B_XL0xSoKd8_1(.din(w_dff_B_zEtFVFdN7_1),.dout(w_dff_B_XL0xSoKd8_1),.clk(gclk));
	jdff dff_B_JAMoUcrp2_1(.din(w_dff_B_XL0xSoKd8_1),.dout(w_dff_B_JAMoUcrp2_1),.clk(gclk));
	jdff dff_B_52tih4US5_0(.din(n283),.dout(w_dff_B_52tih4US5_0),.clk(gclk));
	jdff dff_B_a3R5Amyo4_0(.din(w_dff_B_52tih4US5_0),.dout(w_dff_B_a3R5Amyo4_0),.clk(gclk));
	jdff dff_B_DS6bcRlE0_0(.din(w_dff_B_a3R5Amyo4_0),.dout(w_dff_B_DS6bcRlE0_0),.clk(gclk));
	jdff dff_B_yMwr3pGu7_0(.din(w_dff_B_DS6bcRlE0_0),.dout(w_dff_B_yMwr3pGu7_0),.clk(gclk));
	jdff dff_A_cnSOicKp4_1(.dout(w_n253_0[1]),.din(w_dff_A_cnSOicKp4_1),.clk(gclk));
	jdff dff_A_3iMvnEdv2_1(.dout(w_dff_A_cnSOicKp4_1),.din(w_dff_A_3iMvnEdv2_1),.clk(gclk));
	jdff dff_A_PP6xv8B28_1(.dout(w_dff_A_3iMvnEdv2_1),.din(w_dff_A_PP6xv8B28_1),.clk(gclk));
	jdff dff_A_G1zTjTjC7_1(.dout(w_dff_A_PP6xv8B28_1),.din(w_dff_A_G1zTjTjC7_1),.clk(gclk));
	jdff dff_A_USMqUlZT0_1(.dout(w_dff_A_G1zTjTjC7_1),.din(w_dff_A_USMqUlZT0_1),.clk(gclk));
	jdff dff_B_9IqYxDq65_1(.din(n148),.dout(w_dff_B_9IqYxDq65_1),.clk(gclk));
	jdff dff_B_rbsEoq272_0(.din(n212),.dout(w_dff_B_rbsEoq272_0),.clk(gclk));
	jdff dff_A_6w3XrPb50_0(.dout(w_n211_0[0]),.din(w_dff_A_6w3XrPb50_0),.clk(gclk));
	jdff dff_A_P6xyLfQo8_0(.dout(w_dff_A_6w3XrPb50_0),.din(w_dff_A_P6xyLfQo8_0),.clk(gclk));
	jdff dff_A_TbntlUCQ0_0(.dout(w_dff_A_P6xyLfQo8_0),.din(w_dff_A_TbntlUCQ0_0),.clk(gclk));
	jdff dff_A_niiZHyDf9_0(.dout(w_dff_A_TbntlUCQ0_0),.din(w_dff_A_niiZHyDf9_0),.clk(gclk));
	jdff dff_A_eNncHZYl5_0(.dout(w_dff_A_niiZHyDf9_0),.din(w_dff_A_eNncHZYl5_0),.clk(gclk));
	jdff dff_A_iNsHqmcB9_0(.dout(w_dff_A_eNncHZYl5_0),.din(w_dff_A_iNsHqmcB9_0),.clk(gclk));
	jdff dff_A_75bDSFoY0_0(.dout(w_n209_0[0]),.din(w_dff_A_75bDSFoY0_0),.clk(gclk));
	jdff dff_A_NHcGcBLA5_0(.dout(w_dff_A_75bDSFoY0_0),.din(w_dff_A_NHcGcBLA5_0),.clk(gclk));
	jdff dff_A_RILjHrJd7_0(.dout(w_dff_A_NHcGcBLA5_0),.din(w_dff_A_RILjHrJd7_0),.clk(gclk));
	jdff dff_A_X4OhDqV63_0(.dout(w_dff_A_RILjHrJd7_0),.din(w_dff_A_X4OhDqV63_0),.clk(gclk));
	jdff dff_A_6I3Xz4tf1_0(.dout(w_dff_A_X4OhDqV63_0),.din(w_dff_A_6I3Xz4tf1_0),.clk(gclk));
	jdff dff_B_cdYsUHPR7_2(.din(n209),.dout(w_dff_B_cdYsUHPR7_2),.clk(gclk));
	jdff dff_B_PigP3P9I7_2(.din(w_dff_B_cdYsUHPR7_2),.dout(w_dff_B_PigP3P9I7_2),.clk(gclk));
	jdff dff_B_t3QDEiRX2_2(.din(w_dff_B_PigP3P9I7_2),.dout(w_dff_B_t3QDEiRX2_2),.clk(gclk));
	jdff dff_B_lyURepkx2_2(.din(w_dff_B_t3QDEiRX2_2),.dout(w_dff_B_lyURepkx2_2),.clk(gclk));
	jdff dff_B_3B9PK8623_2(.din(w_dff_B_lyURepkx2_2),.dout(w_dff_B_3B9PK8623_2),.clk(gclk));
	jdff dff_B_klbztqoW1_2(.din(w_dff_B_3B9PK8623_2),.dout(w_dff_B_klbztqoW1_2),.clk(gclk));
	jdff dff_B_Ay7FmcZt3_2(.din(w_dff_B_klbztqoW1_2),.dout(w_dff_B_Ay7FmcZt3_2),.clk(gclk));
	jdff dff_B_a4PjgekG0_2(.din(w_dff_B_Ay7FmcZt3_2),.dout(w_dff_B_a4PjgekG0_2),.clk(gclk));
	jdff dff_B_0sLZaZ0C9_2(.din(w_dff_B_a4PjgekG0_2),.dout(w_dff_B_0sLZaZ0C9_2),.clk(gclk));
	jdff dff_B_Dwxc4tOo5_2(.din(w_dff_B_0sLZaZ0C9_2),.dout(w_dff_B_Dwxc4tOo5_2),.clk(gclk));
	jdff dff_B_53WsXVy56_2(.din(w_dff_B_Dwxc4tOo5_2),.dout(w_dff_B_53WsXVy56_2),.clk(gclk));
	jdff dff_B_ZKIIDDwF9_2(.din(w_dff_B_53WsXVy56_2),.dout(w_dff_B_ZKIIDDwF9_2),.clk(gclk));
	jdff dff_B_VLULyZFX3_2(.din(w_dff_B_ZKIIDDwF9_2),.dout(w_dff_B_VLULyZFX3_2),.clk(gclk));
	jdff dff_B_meL2PgNV6_2(.din(w_dff_B_VLULyZFX3_2),.dout(w_dff_B_meL2PgNV6_2),.clk(gclk));
	jdff dff_A_pna7zWFq8_0(.dout(w_n206_0[0]),.din(w_dff_A_pna7zWFq8_0),.clk(gclk));
	jdff dff_A_6SuufCPf4_0(.dout(w_dff_A_pna7zWFq8_0),.din(w_dff_A_6SuufCPf4_0),.clk(gclk));
	jdff dff_A_foeaykq62_0(.dout(w_dff_A_6SuufCPf4_0),.din(w_dff_A_foeaykq62_0),.clk(gclk));
	jdff dff_A_4znjuRdk8_0(.dout(w_dff_A_foeaykq62_0),.din(w_dff_A_4znjuRdk8_0),.clk(gclk));
	jdff dff_A_OwzA9siF2_0(.dout(w_dff_A_4znjuRdk8_0),.din(w_dff_A_OwzA9siF2_0),.clk(gclk));
	jdff dff_A_QICiSLGL9_0(.dout(w_dff_A_OwzA9siF2_0),.din(w_dff_A_QICiSLGL9_0),.clk(gclk));
	jdff dff_A_XkXZ0vP80_0(.dout(w_n204_0[0]),.din(w_dff_A_XkXZ0vP80_0),.clk(gclk));
	jdff dff_A_oOu6h61c0_0(.dout(w_dff_A_XkXZ0vP80_0),.din(w_dff_A_oOu6h61c0_0),.clk(gclk));
	jdff dff_A_iDlsSKQD2_0(.dout(w_dff_A_oOu6h61c0_0),.din(w_dff_A_iDlsSKQD2_0),.clk(gclk));
	jdff dff_A_6CgZkNlh1_0(.dout(w_dff_A_iDlsSKQD2_0),.din(w_dff_A_6CgZkNlh1_0),.clk(gclk));
	jdff dff_A_zs8YKF2e3_0(.dout(w_dff_A_6CgZkNlh1_0),.din(w_dff_A_zs8YKF2e3_0),.clk(gclk));
	jdff dff_B_d8WufGIU6_2(.din(n204),.dout(w_dff_B_d8WufGIU6_2),.clk(gclk));
	jdff dff_B_HS906qcc6_2(.din(w_dff_B_d8WufGIU6_2),.dout(w_dff_B_HS906qcc6_2),.clk(gclk));
	jdff dff_B_emxqyXlt3_2(.din(w_dff_B_HS906qcc6_2),.dout(w_dff_B_emxqyXlt3_2),.clk(gclk));
	jdff dff_B_GShhl6df7_2(.din(w_dff_B_emxqyXlt3_2),.dout(w_dff_B_GShhl6df7_2),.clk(gclk));
	jdff dff_B_IzvDEbq43_2(.din(w_dff_B_GShhl6df7_2),.dout(w_dff_B_IzvDEbq43_2),.clk(gclk));
	jdff dff_B_Qfzo6o843_2(.din(w_dff_B_IzvDEbq43_2),.dout(w_dff_B_Qfzo6o843_2),.clk(gclk));
	jdff dff_B_xAKdQLAb0_2(.din(w_dff_B_Qfzo6o843_2),.dout(w_dff_B_xAKdQLAb0_2),.clk(gclk));
	jdff dff_B_IOM21WA49_2(.din(w_dff_B_xAKdQLAb0_2),.dout(w_dff_B_IOM21WA49_2),.clk(gclk));
	jdff dff_B_hPfCIXVH7_2(.din(w_dff_B_IOM21WA49_2),.dout(w_dff_B_hPfCIXVH7_2),.clk(gclk));
	jdff dff_B_NdxVDHo48_2(.din(w_dff_B_hPfCIXVH7_2),.dout(w_dff_B_NdxVDHo48_2),.clk(gclk));
	jdff dff_B_2ZOsculb0_2(.din(w_dff_B_NdxVDHo48_2),.dout(w_dff_B_2ZOsculb0_2),.clk(gclk));
	jdff dff_B_PkP4nR5V3_2(.din(w_dff_B_2ZOsculb0_2),.dout(w_dff_B_PkP4nR5V3_2),.clk(gclk));
	jdff dff_B_gN3uTzN49_2(.din(w_dff_B_PkP4nR5V3_2),.dout(w_dff_B_gN3uTzN49_2),.clk(gclk));
	jdff dff_B_i1S2LK491_2(.din(w_dff_B_gN3uTzN49_2),.dout(w_dff_B_i1S2LK491_2),.clk(gclk));
	jdff dff_B_hSN3jX8C9_1(.din(n194),.dout(w_dff_B_hSN3jX8C9_1),.clk(gclk));
	jdff dff_B_UN0gIONJ9_1(.din(w_dff_B_hSN3jX8C9_1),.dout(w_dff_B_UN0gIONJ9_1),.clk(gclk));
	jdff dff_B_quwS2UZ37_1(.din(w_dff_B_UN0gIONJ9_1),.dout(w_dff_B_quwS2UZ37_1),.clk(gclk));
	jdff dff_B_eMfrHHK78_1(.din(w_dff_B_quwS2UZ37_1),.dout(w_dff_B_eMfrHHK78_1),.clk(gclk));
	jdff dff_B_bQEPOnxS9_1(.din(w_dff_B_eMfrHHK78_1),.dout(w_dff_B_bQEPOnxS9_1),.clk(gclk));
	jdff dff_B_GUzvpdtD6_1(.din(w_dff_B_bQEPOnxS9_1),.dout(w_dff_B_GUzvpdtD6_1),.clk(gclk));
	jdff dff_B_jhOqW2AQ2_1(.din(w_dff_B_GUzvpdtD6_1),.dout(w_dff_B_jhOqW2AQ2_1),.clk(gclk));
	jdff dff_B_H7cAMaLf2_1(.din(w_dff_B_jhOqW2AQ2_1),.dout(w_dff_B_H7cAMaLf2_1),.clk(gclk));
	jdff dff_B_KzVFbklm1_1(.din(w_dff_B_H7cAMaLf2_1),.dout(w_dff_B_KzVFbklm1_1),.clk(gclk));
	jdff dff_B_bvFIEeEr2_1(.din(w_dff_B_KzVFbklm1_1),.dout(w_dff_B_bvFIEeEr2_1),.clk(gclk));
	jdff dff_B_IpfMBLA47_1(.din(w_dff_B_bvFIEeEr2_1),.dout(w_dff_B_IpfMBLA47_1),.clk(gclk));
	jdff dff_B_8nLJvSQB1_1(.din(w_dff_B_IpfMBLA47_1),.dout(w_dff_B_8nLJvSQB1_1),.clk(gclk));
	jdff dff_B_OtfSRp3W8_1(.din(w_dff_B_8nLJvSQB1_1),.dout(w_dff_B_OtfSRp3W8_1),.clk(gclk));
	jdff dff_B_CSHAgvXc6_1(.din(w_dff_B_OtfSRp3W8_1),.dout(w_dff_B_CSHAgvXc6_1),.clk(gclk));
	jdff dff_B_ahpQh7Hq2_1(.din(n190),.dout(w_dff_B_ahpQh7Hq2_1),.clk(gclk));
	jdff dff_B_H9eeFopC3_1(.din(w_dff_B_ahpQh7Hq2_1),.dout(w_dff_B_H9eeFopC3_1),.clk(gclk));
	jdff dff_B_3ybyy3hW3_1(.din(w_dff_B_H9eeFopC3_1),.dout(w_dff_B_3ybyy3hW3_1),.clk(gclk));
	jdff dff_B_ZERgL2zy9_1(.din(w_dff_B_3ybyy3hW3_1),.dout(w_dff_B_ZERgL2zy9_1),.clk(gclk));
	jdff dff_B_0FtBJo2C0_1(.din(w_dff_B_ZERgL2zy9_1),.dout(w_dff_B_0FtBJo2C0_1),.clk(gclk));
	jdff dff_B_eMTLxAtr9_1(.din(w_dff_B_0FtBJo2C0_1),.dout(w_dff_B_eMTLxAtr9_1),.clk(gclk));
	jdff dff_B_X8pu3I4w2_1(.din(w_dff_B_eMTLxAtr9_1),.dout(w_dff_B_X8pu3I4w2_1),.clk(gclk));
	jdff dff_B_FppoivKJ5_1(.din(w_dff_B_X8pu3I4w2_1),.dout(w_dff_B_FppoivKJ5_1),.clk(gclk));
	jdff dff_B_JqgPeDQ92_1(.din(w_dff_B_FppoivKJ5_1),.dout(w_dff_B_JqgPeDQ92_1),.clk(gclk));
	jdff dff_B_Pm1mYZYb5_1(.din(w_dff_B_JqgPeDQ92_1),.dout(w_dff_B_Pm1mYZYb5_1),.clk(gclk));
	jdff dff_B_9eoe5DiQ4_1(.din(w_dff_B_Pm1mYZYb5_1),.dout(w_dff_B_9eoe5DiQ4_1),.clk(gclk));
	jdff dff_B_y119Gm4e1_1(.din(w_dff_B_9eoe5DiQ4_1),.dout(w_dff_B_y119Gm4e1_1),.clk(gclk));
	jdff dff_B_PPTVKxs89_1(.din(w_dff_B_y119Gm4e1_1),.dout(w_dff_B_PPTVKxs89_1),.clk(gclk));
	jdff dff_B_6hCX4gzq3_1(.din(w_dff_B_PPTVKxs89_1),.dout(w_dff_B_6hCX4gzq3_1),.clk(gclk));
	jdff dff_A_hbIzBRil4_0(.dout(w_n185_0[0]),.din(w_dff_A_hbIzBRil4_0),.clk(gclk));
	jdff dff_A_xWkEArkY2_0(.dout(w_dff_A_hbIzBRil4_0),.din(w_dff_A_xWkEArkY2_0),.clk(gclk));
	jdff dff_A_VzSf0tvp2_0(.dout(w_dff_A_xWkEArkY2_0),.din(w_dff_A_VzSf0tvp2_0),.clk(gclk));
	jdff dff_A_MOnorS0Q2_0(.dout(w_dff_A_VzSf0tvp2_0),.din(w_dff_A_MOnorS0Q2_0),.clk(gclk));
	jdff dff_A_LoqwA0X89_0(.dout(w_dff_A_MOnorS0Q2_0),.din(w_dff_A_LoqwA0X89_0),.clk(gclk));
	jdff dff_B_o1HFGAr20_2(.din(n185),.dout(w_dff_B_o1HFGAr20_2),.clk(gclk));
	jdff dff_B_kwWDYk5C7_2(.din(w_dff_B_o1HFGAr20_2),.dout(w_dff_B_kwWDYk5C7_2),.clk(gclk));
	jdff dff_B_TAQ6QRbC4_2(.din(w_dff_B_kwWDYk5C7_2),.dout(w_dff_B_TAQ6QRbC4_2),.clk(gclk));
	jdff dff_B_D2DJvxiQ0_2(.din(w_dff_B_TAQ6QRbC4_2),.dout(w_dff_B_D2DJvxiQ0_2),.clk(gclk));
	jdff dff_B_8tIFyV6u7_2(.din(w_dff_B_D2DJvxiQ0_2),.dout(w_dff_B_8tIFyV6u7_2),.clk(gclk));
	jdff dff_B_ShlRA1jJ9_2(.din(w_dff_B_8tIFyV6u7_2),.dout(w_dff_B_ShlRA1jJ9_2),.clk(gclk));
	jdff dff_B_MFHLqJBc9_2(.din(w_dff_B_ShlRA1jJ9_2),.dout(w_dff_B_MFHLqJBc9_2),.clk(gclk));
	jdff dff_B_Tbepjkxg3_2(.din(w_dff_B_MFHLqJBc9_2),.dout(w_dff_B_Tbepjkxg3_2),.clk(gclk));
	jdff dff_B_WkuYxLfV3_2(.din(w_dff_B_Tbepjkxg3_2),.dout(w_dff_B_WkuYxLfV3_2),.clk(gclk));
	jdff dff_B_xXizeWOv0_2(.din(w_dff_B_WkuYxLfV3_2),.dout(w_dff_B_xXizeWOv0_2),.clk(gclk));
	jdff dff_B_yogZZlHe7_2(.din(w_dff_B_xXizeWOv0_2),.dout(w_dff_B_yogZZlHe7_2),.clk(gclk));
	jdff dff_B_aggZKSxg1_2(.din(w_dff_B_yogZZlHe7_2),.dout(w_dff_B_aggZKSxg1_2),.clk(gclk));
	jdff dff_B_waK8gA0f1_2(.din(w_dff_B_aggZKSxg1_2),.dout(w_dff_B_waK8gA0f1_2),.clk(gclk));
	jdff dff_B_Sj0dESrj1_2(.din(w_dff_B_waK8gA0f1_2),.dout(w_dff_B_Sj0dESrj1_2),.clk(gclk));
	jdff dff_B_j2A0JnKG7_2(.din(n281),.dout(w_dff_B_j2A0JnKG7_2),.clk(gclk));
	jdff dff_A_z3SpAsBY9_0(.dout(w_n149_0[0]),.din(w_dff_A_z3SpAsBY9_0),.clk(gclk));
	jdff dff_A_h4vlfbh53_0(.dout(w_dff_A_z3SpAsBY9_0),.din(w_dff_A_h4vlfbh53_0),.clk(gclk));
	jdff dff_A_iOmNIkL74_0(.dout(w_dff_A_h4vlfbh53_0),.din(w_dff_A_iOmNIkL74_0),.clk(gclk));
	jdff dff_A_kvCzikRY8_0(.dout(w_dff_A_iOmNIkL74_0),.din(w_dff_A_kvCzikRY8_0),.clk(gclk));
	jdff dff_A_JHX29h7K1_0(.dout(w_dff_A_kvCzikRY8_0),.din(w_dff_A_JHX29h7K1_0),.clk(gclk));
	jdff dff_B_TXVJFZdx9_2(.din(n149),.dout(w_dff_B_TXVJFZdx9_2),.clk(gclk));
	jdff dff_B_CdOhYngW4_2(.din(w_dff_B_TXVJFZdx9_2),.dout(w_dff_B_CdOhYngW4_2),.clk(gclk));
	jdff dff_B_srtBb4KE9_2(.din(w_dff_B_CdOhYngW4_2),.dout(w_dff_B_srtBb4KE9_2),.clk(gclk));
	jdff dff_B_E5b1TohV2_2(.din(w_dff_B_srtBb4KE9_2),.dout(w_dff_B_E5b1TohV2_2),.clk(gclk));
	jdff dff_B_lBgeFI7Q9_2(.din(w_dff_B_E5b1TohV2_2),.dout(w_dff_B_lBgeFI7Q9_2),.clk(gclk));
	jdff dff_B_BpaOmRlf2_2(.din(w_dff_B_lBgeFI7Q9_2),.dout(w_dff_B_BpaOmRlf2_2),.clk(gclk));
	jdff dff_B_RD9Kn9XY6_2(.din(w_dff_B_BpaOmRlf2_2),.dout(w_dff_B_RD9Kn9XY6_2),.clk(gclk));
	jdff dff_B_TQK1Qdis4_2(.din(w_dff_B_RD9Kn9XY6_2),.dout(w_dff_B_TQK1Qdis4_2),.clk(gclk));
	jdff dff_B_e1Jzoar65_2(.din(w_dff_B_TQK1Qdis4_2),.dout(w_dff_B_e1Jzoar65_2),.clk(gclk));
	jdff dff_B_OvTt47YR2_2(.din(w_dff_B_e1Jzoar65_2),.dout(w_dff_B_OvTt47YR2_2),.clk(gclk));
	jdff dff_B_vxLDuHaH6_2(.din(w_dff_B_OvTt47YR2_2),.dout(w_dff_B_vxLDuHaH6_2),.clk(gclk));
	jdff dff_B_8OCXqUup1_2(.din(w_dff_B_vxLDuHaH6_2),.dout(w_dff_B_8OCXqUup1_2),.clk(gclk));
	jdff dff_B_tmfxmr9z1_2(.din(w_dff_B_8OCXqUup1_2),.dout(w_dff_B_tmfxmr9z1_2),.clk(gclk));
	jdff dff_B_y9kN6HzJ7_2(.din(w_dff_B_tmfxmr9z1_2),.dout(w_dff_B_y9kN6HzJ7_2),.clk(gclk));
	jdff dff_A_KrIZNGa98_0(.dout(w_n183_0[0]),.din(w_dff_A_KrIZNGa98_0),.clk(gclk));
	jdff dff_A_6YdQI9NW3_0(.dout(w_dff_A_KrIZNGa98_0),.din(w_dff_A_6YdQI9NW3_0),.clk(gclk));
	jdff dff_A_FyMZjLpX9_0(.dout(w_dff_A_6YdQI9NW3_0),.din(w_dff_A_FyMZjLpX9_0),.clk(gclk));
	jdff dff_A_JzvDndrG6_0(.dout(w_dff_A_FyMZjLpX9_0),.din(w_dff_A_JzvDndrG6_0),.clk(gclk));
	jdff dff_A_EYG2HVQB7_0(.dout(w_dff_A_JzvDndrG6_0),.din(w_dff_A_EYG2HVQB7_0),.clk(gclk));
	jdff dff_A_zLTzD8dK1_0(.dout(w_dff_A_EYG2HVQB7_0),.din(w_dff_A_zLTzD8dK1_0),.clk(gclk));
	jdff dff_A_L5OcRHyo7_0(.dout(w_n271_0[0]),.din(w_dff_A_L5OcRHyo7_0),.clk(gclk));
	jdff dff_A_UvEyALCO5_0(.dout(w_dff_A_L5OcRHyo7_0),.din(w_dff_A_UvEyALCO5_0),.clk(gclk));
	jdff dff_A_p31a5J3T1_0(.dout(w_dff_A_UvEyALCO5_0),.din(w_dff_A_p31a5J3T1_0),.clk(gclk));
	jdff dff_B_wE7cgOgy0_1(.din(n217),.dout(w_dff_B_wE7cgOgy0_1),.clk(gclk));
	jdff dff_B_dcHqjuw37_0(.din(n243),.dout(w_dff_B_dcHqjuw37_0),.clk(gclk));
	jdff dff_A_ouB13RQR3_0(.dout(w_G27gat_0[0]),.din(w_dff_A_ouB13RQR3_0),.clk(gclk));
	jdff dff_A_Xwi1K41p4_0(.dout(w_dff_A_ouB13RQR3_0),.din(w_dff_A_Xwi1K41p4_0),.clk(gclk));
	jdff dff_A_sZGuDTaw4_0(.dout(w_dff_A_Xwi1K41p4_0),.din(w_dff_A_sZGuDTaw4_0),.clk(gclk));
	jdff dff_A_g0aJYL8b2_0(.dout(w_dff_A_sZGuDTaw4_0),.din(w_dff_A_g0aJYL8b2_0),.clk(gclk));
	jdff dff_A_FD32KFaa3_0(.dout(w_dff_A_g0aJYL8b2_0),.din(w_dff_A_FD32KFaa3_0),.clk(gclk));
	jdff dff_A_SDE9snpP9_0(.dout(w_dff_A_FD32KFaa3_0),.din(w_dff_A_SDE9snpP9_0),.clk(gclk));
	jdff dff_A_eoze8ZM17_0(.dout(w_dff_A_SDE9snpP9_0),.din(w_dff_A_eoze8ZM17_0),.clk(gclk));
	jdff dff_A_7Hj6DsUx8_0(.dout(w_dff_A_eoze8ZM17_0),.din(w_dff_A_7Hj6DsUx8_0),.clk(gclk));
	jdff dff_A_0ywwW8Rq8_0(.dout(w_dff_A_7Hj6DsUx8_0),.din(w_dff_A_0ywwW8Rq8_0),.clk(gclk));
	jdff dff_A_rCoCTJoI5_0(.dout(w_dff_A_0ywwW8Rq8_0),.din(w_dff_A_rCoCTJoI5_0),.clk(gclk));
	jdff dff_A_lzKY9Q687_0(.dout(w_dff_A_rCoCTJoI5_0),.din(w_dff_A_lzKY9Q687_0),.clk(gclk));
	jdff dff_A_U7hcyydb5_0(.dout(w_dff_A_lzKY9Q687_0),.din(w_dff_A_U7hcyydb5_0),.clk(gclk));
	jdff dff_A_KhqhNqe23_0(.dout(w_dff_A_U7hcyydb5_0),.din(w_dff_A_KhqhNqe23_0),.clk(gclk));
	jdff dff_A_gBUzPPL46_0(.dout(w_dff_A_KhqhNqe23_0),.din(w_dff_A_gBUzPPL46_0),.clk(gclk));
	jdff dff_A_7gL6YP9d9_0(.dout(w_dff_A_gBUzPPL46_0),.din(w_dff_A_7gL6YP9d9_0),.clk(gclk));
	jdff dff_A_eV8Lx7100_0(.dout(w_G115gat_0[0]),.din(w_dff_A_eV8Lx7100_0),.clk(gclk));
	jdff dff_A_wGbATrVY0_0(.dout(w_dff_A_eV8Lx7100_0),.din(w_dff_A_wGbATrVY0_0),.clk(gclk));
	jdff dff_A_vuYSf4N41_0(.dout(w_dff_A_wGbATrVY0_0),.din(w_dff_A_vuYSf4N41_0),.clk(gclk));
	jdff dff_A_YmlLkxql5_0(.dout(w_dff_A_vuYSf4N41_0),.din(w_dff_A_YmlLkxql5_0),.clk(gclk));
	jdff dff_A_R8I8AAsQ5_0(.dout(w_dff_A_YmlLkxql5_0),.din(w_dff_A_R8I8AAsQ5_0),.clk(gclk));
	jdff dff_A_gs1alE2z3_0(.dout(w_dff_A_R8I8AAsQ5_0),.din(w_dff_A_gs1alE2z3_0),.clk(gclk));
	jdff dff_A_r1CjFEzp9_0(.dout(w_dff_A_gs1alE2z3_0),.din(w_dff_A_r1CjFEzp9_0),.clk(gclk));
	jdff dff_A_i36nh8WP6_0(.dout(w_dff_A_r1CjFEzp9_0),.din(w_dff_A_i36nh8WP6_0),.clk(gclk));
	jdff dff_A_5OMAwbl14_0(.dout(w_dff_A_i36nh8WP6_0),.din(w_dff_A_5OMAwbl14_0),.clk(gclk));
	jdff dff_A_uE08Gi2I7_0(.dout(w_dff_A_5OMAwbl14_0),.din(w_dff_A_uE08Gi2I7_0),.clk(gclk));
	jdff dff_A_LTfavr4G4_0(.dout(w_dff_A_uE08Gi2I7_0),.din(w_dff_A_LTfavr4G4_0),.clk(gclk));
	jdff dff_A_5HCok42Z6_0(.dout(w_dff_A_LTfavr4G4_0),.din(w_dff_A_5HCok42Z6_0),.clk(gclk));
	jdff dff_A_h6tCBzkt0_0(.dout(w_dff_A_5HCok42Z6_0),.din(w_dff_A_h6tCBzkt0_0),.clk(gclk));
	jdff dff_A_bojiUxdi7_0(.dout(w_dff_A_h6tCBzkt0_0),.din(w_dff_A_bojiUxdi7_0),.clk(gclk));
	jdff dff_A_XBgUQi9j7_0(.dout(w_dff_A_bojiUxdi7_0),.din(w_dff_A_XBgUQi9j7_0),.clk(gclk));
	jdff dff_A_k09LsJHf9_0(.dout(w_n230_0[0]),.din(w_dff_A_k09LsJHf9_0),.clk(gclk));
	jdff dff_A_cCbtaSj38_0(.dout(w_dff_A_k09LsJHf9_0),.din(w_dff_A_cCbtaSj38_0),.clk(gclk));
	jdff dff_A_SSwdXTSp0_0(.dout(w_dff_A_cCbtaSj38_0),.din(w_dff_A_SSwdXTSp0_0),.clk(gclk));
	jdff dff_A_eg0q4qZl8_0(.dout(w_dff_A_SSwdXTSp0_0),.din(w_dff_A_eg0q4qZl8_0),.clk(gclk));
	jdff dff_A_jDkb1jpo9_0(.dout(w_dff_A_eg0q4qZl8_0),.din(w_dff_A_jDkb1jpo9_0),.clk(gclk));
	jdff dff_A_bL9BbCqS1_0(.dout(w_dff_A_jDkb1jpo9_0),.din(w_dff_A_bL9BbCqS1_0),.clk(gclk));
	jdff dff_A_C8SQykNj3_0(.dout(w_G92gat_0[0]),.din(w_dff_A_C8SQykNj3_0),.clk(gclk));
	jdff dff_A_leS70mqm1_0(.dout(w_dff_A_C8SQykNj3_0),.din(w_dff_A_leS70mqm1_0),.clk(gclk));
	jdff dff_A_vVYN5yWg5_0(.dout(w_dff_A_leS70mqm1_0),.din(w_dff_A_vVYN5yWg5_0),.clk(gclk));
	jdff dff_A_S0Kla4y45_0(.dout(w_dff_A_vVYN5yWg5_0),.din(w_dff_A_S0Kla4y45_0),.clk(gclk));
	jdff dff_A_pRex8mM39_0(.dout(w_dff_A_S0Kla4y45_0),.din(w_dff_A_pRex8mM39_0),.clk(gclk));
	jdff dff_A_5xBYIMNA9_0(.dout(w_dff_A_pRex8mM39_0),.din(w_dff_A_5xBYIMNA9_0),.clk(gclk));
	jdff dff_A_4EjLBTNK1_0(.dout(w_dff_A_5xBYIMNA9_0),.din(w_dff_A_4EjLBTNK1_0),.clk(gclk));
	jdff dff_A_6ytp8to95_0(.dout(w_dff_A_4EjLBTNK1_0),.din(w_dff_A_6ytp8to95_0),.clk(gclk));
	jdff dff_A_cpPAdx7b7_0(.dout(w_dff_A_6ytp8to95_0),.din(w_dff_A_cpPAdx7b7_0),.clk(gclk));
	jdff dff_A_7VkWFbcc8_0(.dout(w_dff_A_cpPAdx7b7_0),.din(w_dff_A_7VkWFbcc8_0),.clk(gclk));
	jdff dff_A_Gnv9MqAk3_0(.dout(w_dff_A_7VkWFbcc8_0),.din(w_dff_A_Gnv9MqAk3_0),.clk(gclk));
	jdff dff_A_KNZphkKF2_0(.dout(w_dff_A_Gnv9MqAk3_0),.din(w_dff_A_KNZphkKF2_0),.clk(gclk));
	jdff dff_A_NeCADXen4_0(.dout(w_dff_A_KNZphkKF2_0),.din(w_dff_A_NeCADXen4_0),.clk(gclk));
	jdff dff_A_EdgOFw2R9_0(.dout(w_dff_A_NeCADXen4_0),.din(w_dff_A_EdgOFw2R9_0),.clk(gclk));
	jdff dff_A_uJTzLuYp8_0(.dout(w_dff_A_EdgOFw2R9_0),.din(w_dff_A_uJTzLuYp8_0),.clk(gclk));
	jdff dff_A_7jw3osed7_0(.dout(w_dff_A_uJTzLuYp8_0),.din(w_dff_A_7jw3osed7_0),.clk(gclk));
	jdff dff_A_0Wzhe35b9_0(.dout(w_dff_A_7jw3osed7_0),.din(w_dff_A_0Wzhe35b9_0),.clk(gclk));
	jdff dff_A_BqV46oBm3_0(.dout(w_dff_A_0Wzhe35b9_0),.din(w_dff_A_BqV46oBm3_0),.clk(gclk));
	jdff dff_A_00MwMpVh8_0(.dout(w_dff_A_BqV46oBm3_0),.din(w_dff_A_00MwMpVh8_0),.clk(gclk));
	jdff dff_A_7LgXY2hr6_0(.dout(w_dff_A_00MwMpVh8_0),.din(w_dff_A_7LgXY2hr6_0),.clk(gclk));
	jdff dff_A_bSa6l7RW6_1(.dout(w_G92gat_0[1]),.din(w_dff_A_bSa6l7RW6_1),.clk(gclk));
	jdff dff_A_1Z6Vvesv4_1(.dout(w_dff_A_bSa6l7RW6_1),.din(w_dff_A_1Z6Vvesv4_1),.clk(gclk));
	jdff dff_A_WeZ7fiuu0_1(.dout(w_dff_A_1Z6Vvesv4_1),.din(w_dff_A_WeZ7fiuu0_1),.clk(gclk));
	jdff dff_A_t0VpaKQb1_1(.dout(w_dff_A_WeZ7fiuu0_1),.din(w_dff_A_t0VpaKQb1_1),.clk(gclk));
	jdff dff_A_DbMQ5Kkp5_1(.dout(w_dff_A_t0VpaKQb1_1),.din(w_dff_A_DbMQ5Kkp5_1),.clk(gclk));
	jdff dff_A_ZYuRGBwP4_1(.dout(w_dff_A_DbMQ5Kkp5_1),.din(w_dff_A_ZYuRGBwP4_1),.clk(gclk));
	jdff dff_A_Z8JZutAt6_1(.dout(w_dff_A_ZYuRGBwP4_1),.din(w_dff_A_Z8JZutAt6_1),.clk(gclk));
	jdff dff_A_YD7r77AC1_1(.dout(w_dff_A_Z8JZutAt6_1),.din(w_dff_A_YD7r77AC1_1),.clk(gclk));
	jdff dff_A_R7E24HdF0_1(.dout(w_dff_A_YD7r77AC1_1),.din(w_dff_A_R7E24HdF0_1),.clk(gclk));
	jdff dff_A_bK8Fm5t88_1(.dout(w_dff_A_R7E24HdF0_1),.din(w_dff_A_bK8Fm5t88_1),.clk(gclk));
	jdff dff_A_R4i0rjYk5_1(.dout(w_dff_A_bK8Fm5t88_1),.din(w_dff_A_R4i0rjYk5_1),.clk(gclk));
	jdff dff_A_VdhXtesf8_1(.dout(w_dff_A_R4i0rjYk5_1),.din(w_dff_A_VdhXtesf8_1),.clk(gclk));
	jdff dff_A_tZOwrxrb9_1(.dout(w_dff_A_VdhXtesf8_1),.din(w_dff_A_tZOwrxrb9_1),.clk(gclk));
	jdff dff_A_JrmgusHO7_1(.dout(w_dff_A_tZOwrxrb9_1),.din(w_dff_A_JrmgusHO7_1),.clk(gclk));
	jdff dff_A_GGlQsEAT7_1(.dout(w_dff_A_JrmgusHO7_1),.din(w_dff_A_GGlQsEAT7_1),.clk(gclk));
	jdff dff_A_BUrvsHja4_0(.dout(w_n227_0[0]),.din(w_dff_A_BUrvsHja4_0),.clk(gclk));
	jdff dff_A_OcWXa17Y1_0(.dout(w_dff_A_BUrvsHja4_0),.din(w_dff_A_OcWXa17Y1_0),.clk(gclk));
	jdff dff_A_BG0cQmZT7_0(.dout(w_dff_A_OcWXa17Y1_0),.din(w_dff_A_BG0cQmZT7_0),.clk(gclk));
	jdff dff_A_aahn85jA5_0(.dout(w_dff_A_BG0cQmZT7_0),.din(w_dff_A_aahn85jA5_0),.clk(gclk));
	jdff dff_A_FEBuYrZW5_0(.dout(w_dff_A_aahn85jA5_0),.din(w_dff_A_FEBuYrZW5_0),.clk(gclk));
	jdff dff_A_FJ3P9wKY4_0(.dout(w_dff_A_FEBuYrZW5_0),.din(w_dff_A_FJ3P9wKY4_0),.clk(gclk));
	jdff dff_A_JPLY7oM47_0(.dout(w_G14gat_0[0]),.din(w_dff_A_JPLY7oM47_0),.clk(gclk));
	jdff dff_A_R3oU3nPo4_0(.dout(w_dff_A_JPLY7oM47_0),.din(w_dff_A_R3oU3nPo4_0),.clk(gclk));
	jdff dff_A_YYq9HJgt7_0(.dout(w_dff_A_R3oU3nPo4_0),.din(w_dff_A_YYq9HJgt7_0),.clk(gclk));
	jdff dff_A_1RlXYkc87_0(.dout(w_dff_A_YYq9HJgt7_0),.din(w_dff_A_1RlXYkc87_0),.clk(gclk));
	jdff dff_A_QY9Ipw8V4_0(.dout(w_dff_A_1RlXYkc87_0),.din(w_dff_A_QY9Ipw8V4_0),.clk(gclk));
	jdff dff_A_dCJ7UnOL5_0(.dout(w_dff_A_QY9Ipw8V4_0),.din(w_dff_A_dCJ7UnOL5_0),.clk(gclk));
	jdff dff_A_75P5qZAy0_0(.dout(w_dff_A_dCJ7UnOL5_0),.din(w_dff_A_75P5qZAy0_0),.clk(gclk));
	jdff dff_A_WOxpT6gn6_0(.dout(w_dff_A_75P5qZAy0_0),.din(w_dff_A_WOxpT6gn6_0),.clk(gclk));
	jdff dff_A_T2b1KUU77_0(.dout(w_dff_A_WOxpT6gn6_0),.din(w_dff_A_T2b1KUU77_0),.clk(gclk));
	jdff dff_A_JCh726ST6_0(.dout(w_dff_A_T2b1KUU77_0),.din(w_dff_A_JCh726ST6_0),.clk(gclk));
	jdff dff_A_UX51u8a68_0(.dout(w_dff_A_JCh726ST6_0),.din(w_dff_A_UX51u8a68_0),.clk(gclk));
	jdff dff_A_RfRUVYcJ2_0(.dout(w_dff_A_UX51u8a68_0),.din(w_dff_A_RfRUVYcJ2_0),.clk(gclk));
	jdff dff_A_hOAqRrwN1_0(.dout(w_dff_A_RfRUVYcJ2_0),.din(w_dff_A_hOAqRrwN1_0),.clk(gclk));
	jdff dff_A_kdlP9fvG4_0(.dout(w_dff_A_hOAqRrwN1_0),.din(w_dff_A_kdlP9fvG4_0),.clk(gclk));
	jdff dff_A_qhVJUMCa5_0(.dout(w_dff_A_kdlP9fvG4_0),.din(w_dff_A_qhVJUMCa5_0),.clk(gclk));
	jdff dff_A_lObfZyCr0_0(.dout(w_dff_A_qhVJUMCa5_0),.din(w_dff_A_lObfZyCr0_0),.clk(gclk));
	jdff dff_A_yoQXhp4u4_0(.dout(w_dff_A_lObfZyCr0_0),.din(w_dff_A_yoQXhp4u4_0),.clk(gclk));
	jdff dff_A_FfMTUyTq9_0(.dout(w_dff_A_yoQXhp4u4_0),.din(w_dff_A_FfMTUyTq9_0),.clk(gclk));
	jdff dff_A_F7lAHMbZ5_0(.dout(w_dff_A_FfMTUyTq9_0),.din(w_dff_A_F7lAHMbZ5_0),.clk(gclk));
	jdff dff_A_KIT2oVfE1_0(.dout(w_dff_A_F7lAHMbZ5_0),.din(w_dff_A_KIT2oVfE1_0),.clk(gclk));
	jdff dff_A_JKE684fO2_1(.dout(w_G14gat_0[1]),.din(w_dff_A_JKE684fO2_1),.clk(gclk));
	jdff dff_A_rSt4TXBy7_1(.dout(w_dff_A_JKE684fO2_1),.din(w_dff_A_rSt4TXBy7_1),.clk(gclk));
	jdff dff_A_J6Hzp2vL6_1(.dout(w_dff_A_rSt4TXBy7_1),.din(w_dff_A_J6Hzp2vL6_1),.clk(gclk));
	jdff dff_A_FeEW38KQ2_1(.dout(w_dff_A_J6Hzp2vL6_1),.din(w_dff_A_FeEW38KQ2_1),.clk(gclk));
	jdff dff_A_n5vkYsBO7_1(.dout(w_dff_A_FeEW38KQ2_1),.din(w_dff_A_n5vkYsBO7_1),.clk(gclk));
	jdff dff_A_BS9zWpGs5_1(.dout(w_dff_A_n5vkYsBO7_1),.din(w_dff_A_BS9zWpGs5_1),.clk(gclk));
	jdff dff_A_pEoz1OBv7_1(.dout(w_dff_A_BS9zWpGs5_1),.din(w_dff_A_pEoz1OBv7_1),.clk(gclk));
	jdff dff_A_Fu2Vs6AE0_1(.dout(w_dff_A_pEoz1OBv7_1),.din(w_dff_A_Fu2Vs6AE0_1),.clk(gclk));
	jdff dff_A_bDYQFhP55_1(.dout(w_dff_A_Fu2Vs6AE0_1),.din(w_dff_A_bDYQFhP55_1),.clk(gclk));
	jdff dff_A_2VPGrUa42_1(.dout(w_dff_A_bDYQFhP55_1),.din(w_dff_A_2VPGrUa42_1),.clk(gclk));
	jdff dff_A_suCVm50r3_1(.dout(w_dff_A_2VPGrUa42_1),.din(w_dff_A_suCVm50r3_1),.clk(gclk));
	jdff dff_A_NIBZlJdj7_1(.dout(w_dff_A_suCVm50r3_1),.din(w_dff_A_NIBZlJdj7_1),.clk(gclk));
	jdff dff_A_3eQYcUjq8_1(.dout(w_dff_A_NIBZlJdj7_1),.din(w_dff_A_3eQYcUjq8_1),.clk(gclk));
	jdff dff_A_TYCpRd5N7_1(.dout(w_dff_A_3eQYcUjq8_1),.din(w_dff_A_TYCpRd5N7_1),.clk(gclk));
	jdff dff_A_WU7QAd689_1(.dout(w_dff_A_TYCpRd5N7_1),.din(w_dff_A_WU7QAd689_1),.clk(gclk));
	jdff dff_B_WK9KEog83_1(.din(n221),.dout(w_dff_B_WK9KEog83_1),.clk(gclk));
	jdff dff_B_grZPPI3n8_1(.din(w_dff_B_WK9KEog83_1),.dout(w_dff_B_grZPPI3n8_1),.clk(gclk));
	jdff dff_B_02OmAt9I1_1(.din(w_dff_B_grZPPI3n8_1),.dout(w_dff_B_02OmAt9I1_1),.clk(gclk));
	jdff dff_B_2gCBTnE53_1(.din(w_dff_B_02OmAt9I1_1),.dout(w_dff_B_2gCBTnE53_1),.clk(gclk));
	jdff dff_B_a1GBCKnw2_1(.din(w_dff_B_2gCBTnE53_1),.dout(w_dff_B_a1GBCKnw2_1),.clk(gclk));
	jdff dff_A_yhAsLHUh1_0(.dout(w_G66gat_0[0]),.din(w_dff_A_yhAsLHUh1_0),.clk(gclk));
	jdff dff_A_j2SRVSWZ7_0(.dout(w_dff_A_yhAsLHUh1_0),.din(w_dff_A_j2SRVSWZ7_0),.clk(gclk));
	jdff dff_A_oqPGa1lA9_0(.dout(w_dff_A_j2SRVSWZ7_0),.din(w_dff_A_oqPGa1lA9_0),.clk(gclk));
	jdff dff_A_lcDkJHCH7_0(.dout(w_dff_A_oqPGa1lA9_0),.din(w_dff_A_lcDkJHCH7_0),.clk(gclk));
	jdff dff_A_fVVl20bv9_0(.dout(w_dff_A_lcDkJHCH7_0),.din(w_dff_A_fVVl20bv9_0),.clk(gclk));
	jdff dff_A_SuT3eh386_0(.dout(w_dff_A_fVVl20bv9_0),.din(w_dff_A_SuT3eh386_0),.clk(gclk));
	jdff dff_A_1nE3g42z8_0(.dout(w_dff_A_SuT3eh386_0),.din(w_dff_A_1nE3g42z8_0),.clk(gclk));
	jdff dff_A_Eu7zaKVF5_0(.dout(w_dff_A_1nE3g42z8_0),.din(w_dff_A_Eu7zaKVF5_0),.clk(gclk));
	jdff dff_A_TcFdt9j46_0(.dout(w_dff_A_Eu7zaKVF5_0),.din(w_dff_A_TcFdt9j46_0),.clk(gclk));
	jdff dff_A_SdzTQ94W1_0(.dout(w_dff_A_TcFdt9j46_0),.din(w_dff_A_SdzTQ94W1_0),.clk(gclk));
	jdff dff_A_hvrce2D24_0(.dout(w_dff_A_SdzTQ94W1_0),.din(w_dff_A_hvrce2D24_0),.clk(gclk));
	jdff dff_A_LfaykFyx0_0(.dout(w_dff_A_hvrce2D24_0),.din(w_dff_A_LfaykFyx0_0),.clk(gclk));
	jdff dff_A_qVdxKEMW5_0(.dout(w_dff_A_LfaykFyx0_0),.din(w_dff_A_qVdxKEMW5_0),.clk(gclk));
	jdff dff_A_SILs09bL3_0(.dout(w_dff_A_qVdxKEMW5_0),.din(w_dff_A_SILs09bL3_0),.clk(gclk));
	jdff dff_A_VkoZPS2k8_0(.dout(w_dff_A_SILs09bL3_0),.din(w_dff_A_VkoZPS2k8_0),.clk(gclk));
	jdff dff_A_SOsuPz846_0(.dout(w_dff_A_VkoZPS2k8_0),.din(w_dff_A_SOsuPz846_0),.clk(gclk));
	jdff dff_A_pHj5P0KO3_0(.dout(w_dff_A_SOsuPz846_0),.din(w_dff_A_pHj5P0KO3_0),.clk(gclk));
	jdff dff_A_Jodl1kHr9_0(.dout(w_dff_A_pHj5P0KO3_0),.din(w_dff_A_Jodl1kHr9_0),.clk(gclk));
	jdff dff_A_xv87rs4a3_0(.dout(w_dff_A_Jodl1kHr9_0),.din(w_dff_A_xv87rs4a3_0),.clk(gclk));
	jdff dff_A_uKZwDS0q6_0(.dout(w_dff_A_xv87rs4a3_0),.din(w_dff_A_uKZwDS0q6_0),.clk(gclk));
	jdff dff_A_jMIz7C8h3_1(.dout(w_G66gat_0[1]),.din(w_dff_A_jMIz7C8h3_1),.clk(gclk));
	jdff dff_A_1IdMa42O0_1(.dout(w_dff_A_jMIz7C8h3_1),.din(w_dff_A_1IdMa42O0_1),.clk(gclk));
	jdff dff_A_d0ncg8xV9_1(.dout(w_dff_A_1IdMa42O0_1),.din(w_dff_A_d0ncg8xV9_1),.clk(gclk));
	jdff dff_A_LuDJ4YAm5_1(.dout(w_dff_A_d0ncg8xV9_1),.din(w_dff_A_LuDJ4YAm5_1),.clk(gclk));
	jdff dff_A_hVDIqeOx4_1(.dout(w_dff_A_LuDJ4YAm5_1),.din(w_dff_A_hVDIqeOx4_1),.clk(gclk));
	jdff dff_A_O21Mcrh82_1(.dout(w_dff_A_hVDIqeOx4_1),.din(w_dff_A_O21Mcrh82_1),.clk(gclk));
	jdff dff_A_htWH4NPe7_1(.dout(w_dff_A_O21Mcrh82_1),.din(w_dff_A_htWH4NPe7_1),.clk(gclk));
	jdff dff_A_gMJmElbO0_1(.dout(w_dff_A_htWH4NPe7_1),.din(w_dff_A_gMJmElbO0_1),.clk(gclk));
	jdff dff_A_FXJaqxkI0_1(.dout(w_dff_A_gMJmElbO0_1),.din(w_dff_A_FXJaqxkI0_1),.clk(gclk));
	jdff dff_A_xL0Lr6kL9_1(.dout(w_dff_A_FXJaqxkI0_1),.din(w_dff_A_xL0Lr6kL9_1),.clk(gclk));
	jdff dff_A_hW2S2Ij85_1(.dout(w_dff_A_xL0Lr6kL9_1),.din(w_dff_A_hW2S2Ij85_1),.clk(gclk));
	jdff dff_A_hb7DXibW9_1(.dout(w_dff_A_hW2S2Ij85_1),.din(w_dff_A_hb7DXibW9_1),.clk(gclk));
	jdff dff_A_3T6DmOyr0_1(.dout(w_dff_A_hb7DXibW9_1),.din(w_dff_A_3T6DmOyr0_1),.clk(gclk));
	jdff dff_A_X4d6cjKk8_1(.dout(w_dff_A_3T6DmOyr0_1),.din(w_dff_A_X4d6cjKk8_1),.clk(gclk));
	jdff dff_A_UYPDyGoW5_1(.dout(w_dff_A_X4d6cjKk8_1),.din(w_dff_A_UYPDyGoW5_1),.clk(gclk));
	jdff dff_A_qCQw9XKY0_0(.dout(w_G40gat_0[0]),.din(w_dff_A_qCQw9XKY0_0),.clk(gclk));
	jdff dff_A_JtjTntn92_0(.dout(w_dff_A_qCQw9XKY0_0),.din(w_dff_A_JtjTntn92_0),.clk(gclk));
	jdff dff_A_YyI3E8jL9_0(.dout(w_dff_A_JtjTntn92_0),.din(w_dff_A_YyI3E8jL9_0),.clk(gclk));
	jdff dff_A_3vPeYXJb3_0(.dout(w_dff_A_YyI3E8jL9_0),.din(w_dff_A_3vPeYXJb3_0),.clk(gclk));
	jdff dff_A_7hDGEycb2_0(.dout(w_dff_A_3vPeYXJb3_0),.din(w_dff_A_7hDGEycb2_0),.clk(gclk));
	jdff dff_A_YFNNmnBs3_0(.dout(w_dff_A_7hDGEycb2_0),.din(w_dff_A_YFNNmnBs3_0),.clk(gclk));
	jdff dff_A_owZ2ONHU0_0(.dout(w_dff_A_YFNNmnBs3_0),.din(w_dff_A_owZ2ONHU0_0),.clk(gclk));
	jdff dff_A_rAyouTn90_0(.dout(w_dff_A_owZ2ONHU0_0),.din(w_dff_A_rAyouTn90_0),.clk(gclk));
	jdff dff_A_iRmxoRdw8_0(.dout(w_dff_A_rAyouTn90_0),.din(w_dff_A_iRmxoRdw8_0),.clk(gclk));
	jdff dff_A_DOevHaDy3_0(.dout(w_dff_A_iRmxoRdw8_0),.din(w_dff_A_DOevHaDy3_0),.clk(gclk));
	jdff dff_A_nwdt9Yh96_0(.dout(w_dff_A_DOevHaDy3_0),.din(w_dff_A_nwdt9Yh96_0),.clk(gclk));
	jdff dff_A_xQXq5qmb4_0(.dout(w_dff_A_nwdt9Yh96_0),.din(w_dff_A_xQXq5qmb4_0),.clk(gclk));
	jdff dff_A_dkjsXZhx2_0(.dout(w_dff_A_xQXq5qmb4_0),.din(w_dff_A_dkjsXZhx2_0),.clk(gclk));
	jdff dff_A_snA76Se24_0(.dout(w_dff_A_dkjsXZhx2_0),.din(w_dff_A_snA76Se24_0),.clk(gclk));
	jdff dff_A_keiPrwBc3_0(.dout(w_dff_A_snA76Se24_0),.din(w_dff_A_keiPrwBc3_0),.clk(gclk));
	jdff dff_A_sqAm8OBq6_1(.dout(w_n147_0[1]),.din(w_dff_A_sqAm8OBq6_1),.clk(gclk));
	jdff dff_B_cKZQaniF9_0(.din(n146),.dout(w_dff_B_cKZQaniF9_0),.clk(gclk));
	jdff dff_B_k9o0KQBQ9_0(.din(w_dff_B_cKZQaniF9_0),.dout(w_dff_B_k9o0KQBQ9_0),.clk(gclk));
	jdff dff_B_DBInkPzr8_0(.din(w_dff_B_k9o0KQBQ9_0),.dout(w_dff_B_DBInkPzr8_0),.clk(gclk));
	jdff dff_B_h1tH2DaY1_0(.din(w_dff_B_DBInkPzr8_0),.dout(w_dff_B_h1tH2DaY1_0),.clk(gclk));
	jdff dff_B_5iIZ9mmT2_0(.din(w_dff_B_h1tH2DaY1_0),.dout(w_dff_B_5iIZ9mmT2_0),.clk(gclk));
	jdff dff_B_nDQgQQTX0_0(.din(w_dff_B_5iIZ9mmT2_0),.dout(w_dff_B_nDQgQQTX0_0),.clk(gclk));
	jdff dff_A_rFP2X7Ot3_0(.dout(w_n145_0[0]),.din(w_dff_A_rFP2X7Ot3_0),.clk(gclk));
	jdff dff_A_PmNy3l3S7_0(.dout(w_dff_A_rFP2X7Ot3_0),.din(w_dff_A_PmNy3l3S7_0),.clk(gclk));
	jdff dff_A_OGUA7Yfg2_0(.dout(w_dff_A_PmNy3l3S7_0),.din(w_dff_A_OGUA7Yfg2_0),.clk(gclk));
	jdff dff_A_l1MvIUxs8_0(.dout(w_dff_A_OGUA7Yfg2_0),.din(w_dff_A_l1MvIUxs8_0),.clk(gclk));
	jdff dff_A_uN1BM3qe9_0(.dout(w_dff_A_l1MvIUxs8_0),.din(w_dff_A_uN1BM3qe9_0),.clk(gclk));
	jdff dff_A_h2gruX1q6_0(.dout(w_dff_A_uN1BM3qe9_0),.din(w_dff_A_h2gruX1q6_0),.clk(gclk));
	jdff dff_A_ZiyjYaVi2_0(.dout(w_dff_A_h2gruX1q6_0),.din(w_dff_A_ZiyjYaVi2_0),.clk(gclk));
	jdff dff_A_Qp59nlcQ9_0(.dout(w_dff_A_ZiyjYaVi2_0),.din(w_dff_A_Qp59nlcQ9_0),.clk(gclk));
	jdff dff_A_lMmH3DMV3_0(.dout(w_dff_A_Qp59nlcQ9_0),.din(w_dff_A_lMmH3DMV3_0),.clk(gclk));
	jdff dff_A_vyzQ50Oe2_0(.dout(w_dff_A_lMmH3DMV3_0),.din(w_dff_A_vyzQ50Oe2_0),.clk(gclk));
	jdff dff_A_Fdwi0p8x5_0(.dout(w_dff_A_vyzQ50Oe2_0),.din(w_dff_A_Fdwi0p8x5_0),.clk(gclk));
	jdff dff_A_z7sg22NV4_0(.dout(w_dff_A_Fdwi0p8x5_0),.din(w_dff_A_z7sg22NV4_0),.clk(gclk));
	jdff dff_B_ySC9SCAy7_2(.din(n145),.dout(w_dff_B_ySC9SCAy7_2),.clk(gclk));
	jdff dff_B_YAXGXf4H5_2(.din(w_dff_B_ySC9SCAy7_2),.dout(w_dff_B_YAXGXf4H5_2),.clk(gclk));
	jdff dff_B_gufyE0UY3_2(.din(w_dff_B_YAXGXf4H5_2),.dout(w_dff_B_gufyE0UY3_2),.clk(gclk));
	jdff dff_B_0PpXGkgc6_2(.din(w_dff_B_gufyE0UY3_2),.dout(w_dff_B_0PpXGkgc6_2),.clk(gclk));
	jdff dff_B_NNMPcNyT2_2(.din(w_dff_B_0PpXGkgc6_2),.dout(w_dff_B_NNMPcNyT2_2),.clk(gclk));
	jdff dff_B_VXg5wxDF6_2(.din(w_dff_B_NNMPcNyT2_2),.dout(w_dff_B_VXg5wxDF6_2),.clk(gclk));
	jdff dff_B_jxoo1BoU7_2(.din(w_dff_B_VXg5wxDF6_2),.dout(w_dff_B_jxoo1BoU7_2),.clk(gclk));
	jdff dff_A_iEsle1um8_0(.dout(w_G53gat_0[0]),.din(w_dff_A_iEsle1um8_0),.clk(gclk));
	jdff dff_A_xtvhbAgz7_0(.dout(w_dff_A_iEsle1um8_0),.din(w_dff_A_xtvhbAgz7_0),.clk(gclk));
	jdff dff_A_gVfjfpbx0_0(.dout(w_dff_A_xtvhbAgz7_0),.din(w_dff_A_gVfjfpbx0_0),.clk(gclk));
	jdff dff_A_6tRiK9bI8_0(.dout(w_dff_A_gVfjfpbx0_0),.din(w_dff_A_6tRiK9bI8_0),.clk(gclk));
	jdff dff_A_utqPZN1V2_0(.dout(w_dff_A_6tRiK9bI8_0),.din(w_dff_A_utqPZN1V2_0),.clk(gclk));
	jdff dff_A_KWQOLJYA8_0(.dout(w_dff_A_utqPZN1V2_0),.din(w_dff_A_KWQOLJYA8_0),.clk(gclk));
	jdff dff_A_akBvbjZh2_0(.dout(w_dff_A_KWQOLJYA8_0),.din(w_dff_A_akBvbjZh2_0),.clk(gclk));
	jdff dff_A_S4qFHhA64_0(.dout(w_dff_A_akBvbjZh2_0),.din(w_dff_A_S4qFHhA64_0),.clk(gclk));
	jdff dff_A_uSayjKQ25_0(.dout(w_dff_A_S4qFHhA64_0),.din(w_dff_A_uSayjKQ25_0),.clk(gclk));
	jdff dff_A_awbMIBy38_0(.dout(w_dff_A_uSayjKQ25_0),.din(w_dff_A_awbMIBy38_0),.clk(gclk));
	jdff dff_A_Rm7ITCFT2_0(.dout(w_dff_A_awbMIBy38_0),.din(w_dff_A_Rm7ITCFT2_0),.clk(gclk));
	jdff dff_A_n6exB7d33_0(.dout(w_dff_A_Rm7ITCFT2_0),.din(w_dff_A_n6exB7d33_0),.clk(gclk));
	jdff dff_A_LVZ3uWFS9_0(.dout(w_dff_A_n6exB7d33_0),.din(w_dff_A_LVZ3uWFS9_0),.clk(gclk));
	jdff dff_A_sJFh9Q6L0_0(.dout(w_dff_A_LVZ3uWFS9_0),.din(w_dff_A_sJFh9Q6L0_0),.clk(gclk));
	jdff dff_A_J5W4BsEu8_0(.dout(w_dff_A_sJFh9Q6L0_0),.din(w_dff_A_J5W4BsEu8_0),.clk(gclk));
	jdff dff_A_EBA9LwQz5_0(.dout(w_dff_A_J5W4BsEu8_0),.din(w_dff_A_EBA9LwQz5_0),.clk(gclk));
	jdff dff_A_oBwHkyDm1_0(.dout(w_dff_A_EBA9LwQz5_0),.din(w_dff_A_oBwHkyDm1_0),.clk(gclk));
	jdff dff_A_95gPHotj2_0(.dout(w_dff_A_oBwHkyDm1_0),.din(w_dff_A_95gPHotj2_0),.clk(gclk));
	jdff dff_A_Am5UDLDt8_0(.dout(w_dff_A_95gPHotj2_0),.din(w_dff_A_Am5UDLDt8_0),.clk(gclk));
	jdff dff_A_Znhp1xeO2_0(.dout(w_dff_A_Am5UDLDt8_0),.din(w_dff_A_Znhp1xeO2_0),.clk(gclk));
	jdff dff_A_ib5ffShs1_0(.dout(w_n141_0[0]),.din(w_dff_A_ib5ffShs1_0),.clk(gclk));
	jdff dff_B_4DXugcxX7_1(.din(n124),.dout(w_dff_B_4DXugcxX7_1),.clk(gclk));
	jdff dff_B_8kMUfIEC2_1(.din(n129),.dout(w_dff_B_8kMUfIEC2_1),.clk(gclk));
	jdff dff_B_GKh9iShf2_1(.din(w_dff_B_8kMUfIEC2_1),.dout(w_dff_B_GKh9iShf2_1),.clk(gclk));
	jdff dff_B_8JOGPEdp3_1(.din(w_dff_B_GKh9iShf2_1),.dout(w_dff_B_8JOGPEdp3_1),.clk(gclk));
	jdff dff_B_oOLbckUF0_1(.din(w_dff_B_8JOGPEdp3_1),.dout(w_dff_B_oOLbckUF0_1),.clk(gclk));
	jdff dff_B_GWdQCYAe2_1(.din(w_dff_B_oOLbckUF0_1),.dout(w_dff_B_GWdQCYAe2_1),.clk(gclk));
	jdff dff_B_aYB5X7vv5_1(.din(w_dff_B_GWdQCYAe2_1),.dout(w_dff_B_aYB5X7vv5_1),.clk(gclk));
	jdff dff_B_FGBvw4r15_1(.din(w_dff_B_aYB5X7vv5_1),.dout(w_dff_B_FGBvw4r15_1),.clk(gclk));
	jdff dff_A_MDjoAOsQ5_0(.dout(w_n131_0[0]),.din(w_dff_A_MDjoAOsQ5_0),.clk(gclk));
	jdff dff_A_UMWgwLFp8_0(.dout(w_dff_A_MDjoAOsQ5_0),.din(w_dff_A_UMWgwLFp8_0),.clk(gclk));
	jdff dff_A_pJjipAp56_0(.dout(w_dff_A_UMWgwLFp8_0),.din(w_dff_A_pJjipAp56_0),.clk(gclk));
	jdff dff_A_l28gomvj3_0(.dout(w_dff_A_pJjipAp56_0),.din(w_dff_A_l28gomvj3_0),.clk(gclk));
	jdff dff_A_MxVc0yor4_0(.dout(w_dff_A_l28gomvj3_0),.din(w_dff_A_MxVc0yor4_0),.clk(gclk));
	jdff dff_A_0mAW1mXN5_0(.dout(w_dff_A_MxVc0yor4_0),.din(w_dff_A_0mAW1mXN5_0),.clk(gclk));
	jdff dff_A_FXI92NMi3_0(.dout(w_dff_A_0mAW1mXN5_0),.din(w_dff_A_FXI92NMi3_0),.clk(gclk));
	jdff dff_A_VjGIC8EB9_0(.dout(w_n127_0[0]),.din(w_dff_A_VjGIC8EB9_0),.clk(gclk));
	jdff dff_A_OT3PLfim4_0(.dout(w_dff_A_VjGIC8EB9_0),.din(w_dff_A_OT3PLfim4_0),.clk(gclk));
	jdff dff_A_tJ0B2s2A0_0(.dout(w_dff_A_OT3PLfim4_0),.din(w_dff_A_tJ0B2s2A0_0),.clk(gclk));
	jdff dff_A_pSc3zSWP5_0(.dout(w_dff_A_tJ0B2s2A0_0),.din(w_dff_A_pSc3zSWP5_0),.clk(gclk));
	jdff dff_A_uBhXGZHN2_0(.dout(w_dff_A_pSc3zSWP5_0),.din(w_dff_A_uBhXGZHN2_0),.clk(gclk));
	jdff dff_A_pbXfR2hO7_0(.dout(w_dff_A_uBhXGZHN2_0),.din(w_dff_A_pbXfR2hO7_0),.clk(gclk));
	jdff dff_A_IPgss1P70_0(.dout(w_n125_0[0]),.din(w_dff_A_IPgss1P70_0),.clk(gclk));
	jdff dff_A_G0aVskIx5_0(.dout(w_dff_A_IPgss1P70_0),.din(w_dff_A_G0aVskIx5_0),.clk(gclk));
	jdff dff_A_WBxZLyLk5_0(.dout(w_dff_A_G0aVskIx5_0),.din(w_dff_A_WBxZLyLk5_0),.clk(gclk));
	jdff dff_A_oZeyjCbM9_0(.dout(w_dff_A_WBxZLyLk5_0),.din(w_dff_A_oZeyjCbM9_0),.clk(gclk));
	jdff dff_A_om0J4qJz5_0(.dout(w_dff_A_oZeyjCbM9_0),.din(w_dff_A_om0J4qJz5_0),.clk(gclk));
	jdff dff_B_pxpFaRoM0_2(.din(n125),.dout(w_dff_B_pxpFaRoM0_2),.clk(gclk));
	jdff dff_B_6LQsEQ8l5_2(.din(w_dff_B_pxpFaRoM0_2),.dout(w_dff_B_6LQsEQ8l5_2),.clk(gclk));
	jdff dff_B_ArjxqDzQ1_2(.din(w_dff_B_6LQsEQ8l5_2),.dout(w_dff_B_ArjxqDzQ1_2),.clk(gclk));
	jdff dff_B_J165GFxe3_2(.din(w_dff_B_ArjxqDzQ1_2),.dout(w_dff_B_J165GFxe3_2),.clk(gclk));
	jdff dff_B_oCTUljJ76_2(.din(w_dff_B_J165GFxe3_2),.dout(w_dff_B_oCTUljJ76_2),.clk(gclk));
	jdff dff_B_J3FBaEnX3_2(.din(w_dff_B_oCTUljJ76_2),.dout(w_dff_B_J3FBaEnX3_2),.clk(gclk));
	jdff dff_B_gy8RwmTF8_2(.din(w_dff_B_J3FBaEnX3_2),.dout(w_dff_B_gy8RwmTF8_2),.clk(gclk));
	jdff dff_A_Q2aHZ2AR8_0(.dout(w_n123_0[0]),.din(w_dff_A_Q2aHZ2AR8_0),.clk(gclk));
	jdff dff_A_VQSOghpU7_0(.dout(w_dff_A_Q2aHZ2AR8_0),.din(w_dff_A_VQSOghpU7_0),.clk(gclk));
	jdff dff_A_g50Uylmq0_0(.dout(w_dff_A_VQSOghpU7_0),.din(w_dff_A_g50Uylmq0_0),.clk(gclk));
	jdff dff_A_xkWLDgEz5_0(.dout(w_dff_A_g50Uylmq0_0),.din(w_dff_A_xkWLDgEz5_0),.clk(gclk));
	jdff dff_A_aBGkLZjJ0_0(.dout(w_dff_A_xkWLDgEz5_0),.din(w_dff_A_aBGkLZjJ0_0),.clk(gclk));
	jdff dff_A_q0TIis069_0(.dout(w_dff_A_aBGkLZjJ0_0),.din(w_dff_A_q0TIis069_0),.clk(gclk));
	jdff dff_A_W4ZZ7MPk2_0(.dout(w_n121_0[0]),.din(w_dff_A_W4ZZ7MPk2_0),.clk(gclk));
	jdff dff_A_SgDemcaX1_0(.dout(w_dff_A_W4ZZ7MPk2_0),.din(w_dff_A_SgDemcaX1_0),.clk(gclk));
	jdff dff_A_WbnqLGQM2_0(.dout(w_dff_A_SgDemcaX1_0),.din(w_dff_A_WbnqLGQM2_0),.clk(gclk));
	jdff dff_A_lViaLDAp8_0(.dout(w_dff_A_WbnqLGQM2_0),.din(w_dff_A_lViaLDAp8_0),.clk(gclk));
	jdff dff_A_Gz1Wo5EE2_0(.dout(w_dff_A_lViaLDAp8_0),.din(w_dff_A_Gz1Wo5EE2_0),.clk(gclk));
	jdff dff_B_zVvm2PVc8_2(.din(n121),.dout(w_dff_B_zVvm2PVc8_2),.clk(gclk));
	jdff dff_B_VkmgccGa7_2(.din(w_dff_B_zVvm2PVc8_2),.dout(w_dff_B_VkmgccGa7_2),.clk(gclk));
	jdff dff_B_SB6gz8lS6_2(.din(w_dff_B_VkmgccGa7_2),.dout(w_dff_B_SB6gz8lS6_2),.clk(gclk));
	jdff dff_B_qa13KKWe8_2(.din(w_dff_B_SB6gz8lS6_2),.dout(w_dff_B_qa13KKWe8_2),.clk(gclk));
	jdff dff_B_DPQ5NdHZ5_2(.din(w_dff_B_qa13KKWe8_2),.dout(w_dff_B_DPQ5NdHZ5_2),.clk(gclk));
	jdff dff_B_02drxMj56_2(.din(w_dff_B_DPQ5NdHZ5_2),.dout(w_dff_B_02drxMj56_2),.clk(gclk));
	jdff dff_B_MMpWv6I94_2(.din(w_dff_B_02drxMj56_2),.dout(w_dff_B_MMpWv6I94_2),.clk(gclk));
	jdff dff_B_MK2UGFni2_1(.din(n101),.dout(w_dff_B_MK2UGFni2_1),.clk(gclk));
	jdff dff_B_zMVnDgUe7_0(.din(n114),.dout(w_dff_B_zMVnDgUe7_0),.clk(gclk));
	jdff dff_A_6xLzEwn20_0(.dout(w_n113_0[0]),.din(w_dff_A_6xLzEwn20_0),.clk(gclk));
	jdff dff_A_M1ji5M4c3_0(.dout(w_dff_A_6xLzEwn20_0),.din(w_dff_A_M1ji5M4c3_0),.clk(gclk));
	jdff dff_A_zFp14LDU7_0(.dout(w_dff_A_M1ji5M4c3_0),.din(w_dff_A_zFp14LDU7_0),.clk(gclk));
	jdff dff_A_B811KskL6_0(.dout(w_dff_A_zFp14LDU7_0),.din(w_dff_A_B811KskL6_0),.clk(gclk));
	jdff dff_A_xl9l1zNu8_0(.dout(w_dff_A_B811KskL6_0),.din(w_dff_A_xl9l1zNu8_0),.clk(gclk));
	jdff dff_A_7P26Z4cx2_0(.dout(w_dff_A_xl9l1zNu8_0),.din(w_dff_A_7P26Z4cx2_0),.clk(gclk));
	jdff dff_A_MlnUQfpg3_0(.dout(w_n111_0[0]),.din(w_dff_A_MlnUQfpg3_0),.clk(gclk));
	jdff dff_A_bZQqt8Il9_0(.dout(w_dff_A_MlnUQfpg3_0),.din(w_dff_A_bZQqt8Il9_0),.clk(gclk));
	jdff dff_A_Lqj3nDNG1_0(.dout(w_dff_A_bZQqt8Il9_0),.din(w_dff_A_Lqj3nDNG1_0),.clk(gclk));
	jdff dff_A_B9Sli7pD7_0(.dout(w_dff_A_Lqj3nDNG1_0),.din(w_dff_A_B9Sli7pD7_0),.clk(gclk));
	jdff dff_A_8SBupB3J0_0(.dout(w_dff_A_B9Sli7pD7_0),.din(w_dff_A_8SBupB3J0_0),.clk(gclk));
	jdff dff_B_WGfXzdsH6_2(.din(n111),.dout(w_dff_B_WGfXzdsH6_2),.clk(gclk));
	jdff dff_B_sKb7Wm967_2(.din(w_dff_B_WGfXzdsH6_2),.dout(w_dff_B_sKb7Wm967_2),.clk(gclk));
	jdff dff_B_CfkeuXU98_2(.din(w_dff_B_sKb7Wm967_2),.dout(w_dff_B_CfkeuXU98_2),.clk(gclk));
	jdff dff_B_bbl0mFmM6_2(.din(w_dff_B_CfkeuXU98_2),.dout(w_dff_B_bbl0mFmM6_2),.clk(gclk));
	jdff dff_B_adIJcoHX8_2(.din(w_dff_B_bbl0mFmM6_2),.dout(w_dff_B_adIJcoHX8_2),.clk(gclk));
	jdff dff_B_Yr9IKhTo4_2(.din(w_dff_B_adIJcoHX8_2),.dout(w_dff_B_Yr9IKhTo4_2),.clk(gclk));
	jdff dff_B_OfkeaqDE0_2(.din(w_dff_B_Yr9IKhTo4_2),.dout(w_dff_B_OfkeaqDE0_2),.clk(gclk));
	jdff dff_A_PC08HT9Y0_0(.dout(w_n108_0[0]),.din(w_dff_A_PC08HT9Y0_0),.clk(gclk));
	jdff dff_A_oo98AnT41_0(.dout(w_dff_A_PC08HT9Y0_0),.din(w_dff_A_oo98AnT41_0),.clk(gclk));
	jdff dff_A_anNQlfgt9_0(.dout(w_dff_A_oo98AnT41_0),.din(w_dff_A_anNQlfgt9_0),.clk(gclk));
	jdff dff_A_WbEqaL9H4_0(.dout(w_dff_A_anNQlfgt9_0),.din(w_dff_A_WbEqaL9H4_0),.clk(gclk));
	jdff dff_A_0PmFYCQ70_0(.dout(w_dff_A_WbEqaL9H4_0),.din(w_dff_A_0PmFYCQ70_0),.clk(gclk));
	jdff dff_A_I1ALeByX7_0(.dout(w_dff_A_0PmFYCQ70_0),.din(w_dff_A_I1ALeByX7_0),.clk(gclk));
	jdff dff_A_05yPVrX25_0(.dout(w_n106_0[0]),.din(w_dff_A_05yPVrX25_0),.clk(gclk));
	jdff dff_A_UOb6IWM88_0(.dout(w_dff_A_05yPVrX25_0),.din(w_dff_A_UOb6IWM88_0),.clk(gclk));
	jdff dff_A_u7b3FYz57_0(.dout(w_dff_A_UOb6IWM88_0),.din(w_dff_A_u7b3FYz57_0),.clk(gclk));
	jdff dff_A_nCEn706y7_0(.dout(w_dff_A_u7b3FYz57_0),.din(w_dff_A_nCEn706y7_0),.clk(gclk));
	jdff dff_A_HaGm7f1e2_0(.dout(w_dff_A_nCEn706y7_0),.din(w_dff_A_HaGm7f1e2_0),.clk(gclk));
	jdff dff_B_KANx3TDy8_2(.din(n106),.dout(w_dff_B_KANx3TDy8_2),.clk(gclk));
	jdff dff_B_M3GEBIT96_2(.din(w_dff_B_KANx3TDy8_2),.dout(w_dff_B_M3GEBIT96_2),.clk(gclk));
	jdff dff_B_jVrQqdLO8_2(.din(w_dff_B_M3GEBIT96_2),.dout(w_dff_B_jVrQqdLO8_2),.clk(gclk));
	jdff dff_B_zNnCM56m1_2(.din(w_dff_B_jVrQqdLO8_2),.dout(w_dff_B_zNnCM56m1_2),.clk(gclk));
	jdff dff_B_VQbypCJw3_2(.din(w_dff_B_zNnCM56m1_2),.dout(w_dff_B_VQbypCJw3_2),.clk(gclk));
	jdff dff_B_GtN1Zagn7_2(.din(w_dff_B_VQbypCJw3_2),.dout(w_dff_B_GtN1Zagn7_2),.clk(gclk));
	jdff dff_B_mr0pUf0l2_2(.din(w_dff_B_GtN1Zagn7_2),.dout(w_dff_B_mr0pUf0l2_2),.clk(gclk));
	jdff dff_B_HzekDwx63_1(.din(n97),.dout(w_dff_B_HzekDwx63_1),.clk(gclk));
	jdff dff_B_TVhoArzx1_1(.din(w_dff_B_HzekDwx63_1),.dout(w_dff_B_TVhoArzx1_1),.clk(gclk));
	jdff dff_B_sWJOKgQ53_1(.din(w_dff_B_TVhoArzx1_1),.dout(w_dff_B_sWJOKgQ53_1),.clk(gclk));
	jdff dff_B_tsOyWqJd5_1(.din(w_dff_B_sWJOKgQ53_1),.dout(w_dff_B_tsOyWqJd5_1),.clk(gclk));
	jdff dff_B_FgBqOXf90_1(.din(w_dff_B_tsOyWqJd5_1),.dout(w_dff_B_FgBqOXf90_1),.clk(gclk));
	jdff dff_B_vbGj5EFR3_1(.din(w_dff_B_FgBqOXf90_1),.dout(w_dff_B_vbGj5EFR3_1),.clk(gclk));
	jdff dff_B_XXQEqsMp7_1(.din(w_dff_B_vbGj5EFR3_1),.dout(w_dff_B_XXQEqsMp7_1),.clk(gclk));
	jdff dff_A_y0KjvieU4_0(.dout(w_n95_0[0]),.din(w_dff_A_y0KjvieU4_0),.clk(gclk));
	jdff dff_A_VCGhisw99_0(.dout(w_dff_A_y0KjvieU4_0),.din(w_dff_A_VCGhisw99_0),.clk(gclk));
	jdff dff_A_aDHjhZMm0_0(.dout(w_dff_A_VCGhisw99_0),.din(w_dff_A_aDHjhZMm0_0),.clk(gclk));
	jdff dff_A_6b0YLsRo1_0(.dout(w_dff_A_aDHjhZMm0_0),.din(w_dff_A_6b0YLsRo1_0),.clk(gclk));
	jdff dff_A_nNo8Umco1_0(.dout(w_dff_A_6b0YLsRo1_0),.din(w_dff_A_nNo8Umco1_0),.clk(gclk));
	jdff dff_A_zc5jePtT9_0(.dout(w_dff_A_nNo8Umco1_0),.din(w_dff_A_zc5jePtT9_0),.clk(gclk));
	jdff dff_A_7tOG5CNC9_0(.dout(w_n70_0[0]),.din(w_dff_A_7tOG5CNC9_0),.clk(gclk));
	jdff dff_A_fmpfwvpc6_0(.dout(w_dff_A_7tOG5CNC9_0),.din(w_dff_A_fmpfwvpc6_0),.clk(gclk));
	jdff dff_A_6tR1FPKT0_0(.dout(w_dff_A_fmpfwvpc6_0),.din(w_dff_A_6tR1FPKT0_0),.clk(gclk));
	jdff dff_A_oFE9Iqmq0_0(.dout(w_dff_A_6tR1FPKT0_0),.din(w_dff_A_oFE9Iqmq0_0),.clk(gclk));
	jdff dff_A_ACXJhbV32_0(.dout(w_dff_A_oFE9Iqmq0_0),.din(w_dff_A_ACXJhbV32_0),.clk(gclk));
	jdff dff_B_EXmU3giR8_2(.din(n70),.dout(w_dff_B_EXmU3giR8_2),.clk(gclk));
	jdff dff_B_TmpCBnNW7_2(.din(w_dff_B_EXmU3giR8_2),.dout(w_dff_B_TmpCBnNW7_2),.clk(gclk));
	jdff dff_B_Lf1dolqs8_2(.din(w_dff_B_TmpCBnNW7_2),.dout(w_dff_B_Lf1dolqs8_2),.clk(gclk));
	jdff dff_B_uZwg1S0t8_2(.din(w_dff_B_Lf1dolqs8_2),.dout(w_dff_B_uZwg1S0t8_2),.clk(gclk));
	jdff dff_B_XNUlyNiK9_2(.din(w_dff_B_uZwg1S0t8_2),.dout(w_dff_B_XNUlyNiK9_2),.clk(gclk));
	jdff dff_B_0QiJThQf3_2(.din(w_dff_B_XNUlyNiK9_2),.dout(w_dff_B_0QiJThQf3_2),.clk(gclk));
	jdff dff_B_Ubacgs9I4_2(.din(w_dff_B_0QiJThQf3_2),.dout(w_dff_B_Ubacgs9I4_2),.clk(gclk));
	jdff dff_A_cLZeErEF5_1(.dout(w_G105gat_0[1]),.din(w_dff_A_cLZeErEF5_1),.clk(gclk));
	jdff dff_A_YJwq2Zvq8_1(.dout(w_dff_A_cLZeErEF5_1),.din(w_dff_A_YJwq2Zvq8_1),.clk(gclk));
	jdff dff_A_p8rYGSep5_1(.dout(w_dff_A_YJwq2Zvq8_1),.din(w_dff_A_p8rYGSep5_1),.clk(gclk));
	jdff dff_A_qn3GcS4x5_1(.dout(w_dff_A_p8rYGSep5_1),.din(w_dff_A_qn3GcS4x5_1),.clk(gclk));
	jdff dff_A_OE8rw2Yl7_1(.dout(w_dff_A_qn3GcS4x5_1),.din(w_dff_A_OE8rw2Yl7_1),.clk(gclk));
	jdff dff_A_cQrg6etf2_1(.dout(w_dff_A_OE8rw2Yl7_1),.din(w_dff_A_cQrg6etf2_1),.clk(gclk));
	jdff dff_A_y3CrpwWQ9_1(.dout(w_dff_A_cQrg6etf2_1),.din(w_dff_A_y3CrpwWQ9_1),.clk(gclk));
	jdff dff_A_EPYoHhSd8_1(.dout(w_dff_A_y3CrpwWQ9_1),.din(w_dff_A_EPYoHhSd8_1),.clk(gclk));
	jdff dff_A_zp8dRXpZ3_1(.dout(w_dff_A_EPYoHhSd8_1),.din(w_dff_A_zp8dRXpZ3_1),.clk(gclk));
	jdff dff_A_c3n6djoO9_1(.dout(w_dff_A_zp8dRXpZ3_1),.din(w_dff_A_c3n6djoO9_1),.clk(gclk));
	jdff dff_A_jNKQiOuQ6_1(.dout(w_dff_A_c3n6djoO9_1),.din(w_dff_A_jNKQiOuQ6_1),.clk(gclk));
	jdff dff_A_W90tvkBv7_1(.dout(w_dff_A_jNKQiOuQ6_1),.din(w_dff_A_W90tvkBv7_1),.clk(gclk));
	jdff dff_A_4LIxEHvP0_1(.dout(w_dff_A_W90tvkBv7_1),.din(w_dff_A_4LIxEHvP0_1),.clk(gclk));
	jdff dff_A_W4yJQrOz5_1(.dout(w_dff_A_4LIxEHvP0_1),.din(w_dff_A_W4yJQrOz5_1),.clk(gclk));
	jdff dff_A_3J53RKR44_1(.dout(w_dff_A_W4yJQrOz5_1),.din(w_dff_A_3J53RKR44_1),.clk(gclk));
	jdff dff_A_UVCWxBSj6_0(.dout(w_n200_0[0]),.din(w_dff_A_UVCWxBSj6_0),.clk(gclk));
	jdff dff_A_uCLvcsCq4_0(.dout(w_dff_A_UVCWxBSj6_0),.din(w_dff_A_uCLvcsCq4_0),.clk(gclk));
	jdff dff_A_cAK5wk6x4_0(.dout(w_dff_A_uCLvcsCq4_0),.din(w_dff_A_cAK5wk6x4_0),.clk(gclk));
	jdff dff_A_jsGd9WQB7_0(.dout(w_dff_A_cAK5wk6x4_0),.din(w_dff_A_jsGd9WQB7_0),.clk(gclk));
	jdff dff_A_Vo0RVpcN6_0(.dout(w_dff_A_jsGd9WQB7_0),.din(w_dff_A_Vo0RVpcN6_0),.clk(gclk));
	jdff dff_B_Gzw5Bwni2_2(.din(n200),.dout(w_dff_B_Gzw5Bwni2_2),.clk(gclk));
	jdff dff_B_SCuL5UL08_2(.din(w_dff_B_Gzw5Bwni2_2),.dout(w_dff_B_SCuL5UL08_2),.clk(gclk));
	jdff dff_B_JEb5hJMN2_2(.din(w_dff_B_SCuL5UL08_2),.dout(w_dff_B_JEb5hJMN2_2),.clk(gclk));
	jdff dff_B_7DjrZRPu5_2(.din(w_dff_B_JEb5hJMN2_2),.dout(w_dff_B_7DjrZRPu5_2),.clk(gclk));
	jdff dff_B_5tfaG7j98_2(.din(w_dff_B_7DjrZRPu5_2),.dout(w_dff_B_5tfaG7j98_2),.clk(gclk));
	jdff dff_B_CXhyXXLJ0_2(.din(w_dff_B_5tfaG7j98_2),.dout(w_dff_B_CXhyXXLJ0_2),.clk(gclk));
	jdff dff_B_xvGXlgaU1_2(.din(w_dff_B_CXhyXXLJ0_2),.dout(w_dff_B_xvGXlgaU1_2),.clk(gclk));
	jdff dff_B_7eXvcIPj8_2(.din(w_dff_B_xvGXlgaU1_2),.dout(w_dff_B_7eXvcIPj8_2),.clk(gclk));
	jdff dff_B_Z0lqTgGg8_2(.din(w_dff_B_7eXvcIPj8_2),.dout(w_dff_B_Z0lqTgGg8_2),.clk(gclk));
	jdff dff_B_WK8PQyOj0_2(.din(w_dff_B_Z0lqTgGg8_2),.dout(w_dff_B_WK8PQyOj0_2),.clk(gclk));
	jdff dff_B_bWlwbmt07_2(.din(w_dff_B_WK8PQyOj0_2),.dout(w_dff_B_bWlwbmt07_2),.clk(gclk));
	jdff dff_B_HXvx0jsb8_2(.din(w_dff_B_bWlwbmt07_2),.dout(w_dff_B_HXvx0jsb8_2),.clk(gclk));
	jdff dff_B_xnxbckoe6_2(.din(w_dff_B_HXvx0jsb8_2),.dout(w_dff_B_xnxbckoe6_2),.clk(gclk));
	jdff dff_B_0peKtRbm5_2(.din(w_dff_B_xnxbckoe6_2),.dout(w_dff_B_0peKtRbm5_2),.clk(gclk));
	jdff dff_A_spVL2x6z2_0(.dout(w_G79gat_0[0]),.din(w_dff_A_spVL2x6z2_0),.clk(gclk));
	jdff dff_A_Ec7nvYtZ2_0(.dout(w_dff_A_spVL2x6z2_0),.din(w_dff_A_Ec7nvYtZ2_0),.clk(gclk));
	jdff dff_A_ppdqxHB96_0(.dout(w_dff_A_Ec7nvYtZ2_0),.din(w_dff_A_ppdqxHB96_0),.clk(gclk));
	jdff dff_A_eDkZ3wto8_0(.dout(w_dff_A_ppdqxHB96_0),.din(w_dff_A_eDkZ3wto8_0),.clk(gclk));
	jdff dff_A_e1lXdjTl6_0(.dout(w_dff_A_eDkZ3wto8_0),.din(w_dff_A_e1lXdjTl6_0),.clk(gclk));
	jdff dff_A_q2quDH244_0(.dout(w_dff_A_e1lXdjTl6_0),.din(w_dff_A_q2quDH244_0),.clk(gclk));
	jdff dff_A_L8wjvI4q6_0(.dout(w_dff_A_q2quDH244_0),.din(w_dff_A_L8wjvI4q6_0),.clk(gclk));
	jdff dff_A_GA8xiqQi5_0(.dout(w_dff_A_L8wjvI4q6_0),.din(w_dff_A_GA8xiqQi5_0),.clk(gclk));
	jdff dff_A_rTaC778S1_0(.dout(w_dff_A_GA8xiqQi5_0),.din(w_dff_A_rTaC778S1_0),.clk(gclk));
	jdff dff_A_Sn06y3j33_0(.dout(w_dff_A_rTaC778S1_0),.din(w_dff_A_Sn06y3j33_0),.clk(gclk));
	jdff dff_A_QPh8TyZT5_0(.dout(w_dff_A_Sn06y3j33_0),.din(w_dff_A_QPh8TyZT5_0),.clk(gclk));
	jdff dff_A_mtt4fRf73_0(.dout(w_dff_A_QPh8TyZT5_0),.din(w_dff_A_mtt4fRf73_0),.clk(gclk));
	jdff dff_A_9gw6BSS25_0(.dout(w_dff_A_mtt4fRf73_0),.din(w_dff_A_9gw6BSS25_0),.clk(gclk));
	jdff dff_A_ekmdJ2sK3_0(.dout(w_dff_A_9gw6BSS25_0),.din(w_dff_A_ekmdJ2sK3_0),.clk(gclk));
	jdff dff_A_YkuPxYKQ6_0(.dout(w_dff_A_ekmdJ2sK3_0),.din(w_dff_A_YkuPxYKQ6_0),.clk(gclk));
	jdff dff_A_bjcClbaR1_0(.dout(w_n202_0[0]),.din(w_dff_A_bjcClbaR1_0),.clk(gclk));
	jdff dff_A_traNO1Cg9_0(.dout(w_dff_A_bjcClbaR1_0),.din(w_dff_A_traNO1Cg9_0),.clk(gclk));
	jdff dff_A_k1h1GkCY5_0(.dout(w_dff_A_traNO1Cg9_0),.din(w_dff_A_k1h1GkCY5_0),.clk(gclk));
	jdff dff_A_J94BjYdu6_0(.dout(w_dff_A_k1h1GkCY5_0),.din(w_dff_A_J94BjYdu6_0),.clk(gclk));
	jdff dff_A_TsK5Cy9C6_0(.dout(w_dff_A_J94BjYdu6_0),.din(w_dff_A_TsK5Cy9C6_0),.clk(gclk));
	jdff dff_A_YwWieT7T5_0(.dout(w_dff_A_TsK5Cy9C6_0),.din(w_dff_A_YwWieT7T5_0),.clk(gclk));
	jdff dff_B_5CHZjteE6_1(.din(n168),.dout(w_dff_B_5CHZjteE6_1),.clk(gclk));
	jdff dff_B_N5FF0fRm0_1(.din(n171),.dout(w_dff_B_N5FF0fRm0_1),.clk(gclk));
	jdff dff_A_sSdwTqtN8_0(.dout(w_G47gat_0[0]),.din(w_dff_A_sSdwTqtN8_0),.clk(gclk));
	jdff dff_A_NC9vZe4y4_0(.dout(w_dff_A_sSdwTqtN8_0),.din(w_dff_A_NC9vZe4y4_0),.clk(gclk));
	jdff dff_A_dsRlYXKa0_0(.dout(w_dff_A_NC9vZe4y4_0),.din(w_dff_A_dsRlYXKa0_0),.clk(gclk));
	jdff dff_A_A0nPH3QQ1_0(.dout(w_dff_A_dsRlYXKa0_0),.din(w_dff_A_A0nPH3QQ1_0),.clk(gclk));
	jdff dff_A_mMGUuize7_0(.dout(w_dff_A_A0nPH3QQ1_0),.din(w_dff_A_mMGUuize7_0),.clk(gclk));
	jdff dff_A_hhjqW6sl3_0(.dout(w_dff_A_mMGUuize7_0),.din(w_dff_A_hhjqW6sl3_0),.clk(gclk));
	jdff dff_A_Apq31EEP4_0(.dout(w_dff_A_hhjqW6sl3_0),.din(w_dff_A_Apq31EEP4_0),.clk(gclk));
	jdff dff_A_oV3Xayi37_0(.dout(w_dff_A_Apq31EEP4_0),.din(w_dff_A_oV3Xayi37_0),.clk(gclk));
	jdff dff_A_gfoqQjDK5_1(.dout(w_G47gat_0[1]),.din(w_dff_A_gfoqQjDK5_1),.clk(gclk));
	jdff dff_A_CAMTCoCg0_1(.dout(w_dff_A_gfoqQjDK5_1),.din(w_dff_A_CAMTCoCg0_1),.clk(gclk));
	jdff dff_A_eMgtIPQW1_1(.dout(w_dff_A_CAMTCoCg0_1),.din(w_dff_A_eMgtIPQW1_1),.clk(gclk));
	jdff dff_A_K2l6bWI91_1(.dout(w_dff_A_eMgtIPQW1_1),.din(w_dff_A_K2l6bWI91_1),.clk(gclk));
	jdff dff_A_N0irNl0C0_1(.dout(w_dff_A_K2l6bWI91_1),.din(w_dff_A_N0irNl0C0_1),.clk(gclk));
	jdff dff_A_tIbzckN32_1(.dout(w_dff_A_N0irNl0C0_1),.din(w_dff_A_tIbzckN32_1),.clk(gclk));
	jdff dff_A_Wn8GzLHn2_1(.dout(w_dff_A_tIbzckN32_1),.din(w_dff_A_Wn8GzLHn2_1),.clk(gclk));
	jdff dff_A_Zrqt1NQW4_1(.dout(w_dff_A_Wn8GzLHn2_1),.din(w_dff_A_Zrqt1NQW4_1),.clk(gclk));
	jdff dff_A_7xjnVOMN3_1(.dout(w_dff_A_Zrqt1NQW4_1),.din(w_dff_A_7xjnVOMN3_1),.clk(gclk));
	jdff dff_A_9q5YkO6C6_1(.dout(w_dff_A_7xjnVOMN3_1),.din(w_dff_A_9q5YkO6C6_1),.clk(gclk));
	jdff dff_A_ZLJNJwzp0_1(.dout(w_dff_A_9q5YkO6C6_1),.din(w_dff_A_ZLJNJwzp0_1),.clk(gclk));
	jdff dff_A_3ZHAhX0v1_1(.dout(w_dff_A_ZLJNJwzp0_1),.din(w_dff_A_3ZHAhX0v1_1),.clk(gclk));
	jdff dff_A_PMjxuwGC4_1(.dout(w_dff_A_3ZHAhX0v1_1),.din(w_dff_A_PMjxuwGC4_1),.clk(gclk));
	jdff dff_A_AD4xuczk8_0(.dout(w_n173_0[0]),.din(w_dff_A_AD4xuczk8_0),.clk(gclk));
	jdff dff_A_UKfqoEhy9_0(.dout(w_dff_A_AD4xuczk8_0),.din(w_dff_A_UKfqoEhy9_0),.clk(gclk));
	jdff dff_A_4oeBmz9q3_0(.dout(w_dff_A_UKfqoEhy9_0),.din(w_dff_A_4oeBmz9q3_0),.clk(gclk));
	jdff dff_A_hZXzDmHd0_0(.dout(w_dff_A_4oeBmz9q3_0),.din(w_dff_A_hZXzDmHd0_0),.clk(gclk));
	jdff dff_A_PyJBH4GW3_0(.dout(w_dff_A_hZXzDmHd0_0),.din(w_dff_A_PyJBH4GW3_0),.clk(gclk));
	jdff dff_A_8ZaN7ty78_0(.dout(w_dff_A_PyJBH4GW3_0),.din(w_dff_A_8ZaN7ty78_0),.clk(gclk));
	jdff dff_A_un6aqxhM5_0(.dout(w_G8gat_0[0]),.din(w_dff_A_un6aqxhM5_0),.clk(gclk));
	jdff dff_A_w1JLPekb1_0(.dout(w_dff_A_un6aqxhM5_0),.din(w_dff_A_w1JLPekb1_0),.clk(gclk));
	jdff dff_A_zkcMRtOO9_0(.dout(w_dff_A_w1JLPekb1_0),.din(w_dff_A_zkcMRtOO9_0),.clk(gclk));
	jdff dff_A_xa1Nrk0b1_0(.dout(w_dff_A_zkcMRtOO9_0),.din(w_dff_A_xa1Nrk0b1_0),.clk(gclk));
	jdff dff_A_hyZBNk011_0(.dout(w_dff_A_xa1Nrk0b1_0),.din(w_dff_A_hyZBNk011_0),.clk(gclk));
	jdff dff_A_sCBP5Tky8_0(.dout(w_dff_A_hyZBNk011_0),.din(w_dff_A_sCBP5Tky8_0),.clk(gclk));
	jdff dff_A_7GdUoFLc2_0(.dout(w_dff_A_sCBP5Tky8_0),.din(w_dff_A_7GdUoFLc2_0),.clk(gclk));
	jdff dff_A_ZXVf5Nzp2_0(.dout(w_dff_A_7GdUoFLc2_0),.din(w_dff_A_ZXVf5Nzp2_0),.clk(gclk));
	jdff dff_A_mhJoslKp5_0(.dout(w_dff_A_ZXVf5Nzp2_0),.din(w_dff_A_mhJoslKp5_0),.clk(gclk));
	jdff dff_A_F7oiPhA36_0(.dout(w_dff_A_mhJoslKp5_0),.din(w_dff_A_F7oiPhA36_0),.clk(gclk));
	jdff dff_A_5di2L4su3_0(.dout(w_dff_A_F7oiPhA36_0),.din(w_dff_A_5di2L4su3_0),.clk(gclk));
	jdff dff_A_0Dd4OR8I1_0(.dout(w_dff_A_5di2L4su3_0),.din(w_dff_A_0Dd4OR8I1_0),.clk(gclk));
	jdff dff_A_XzwxnOKp0_0(.dout(w_dff_A_0Dd4OR8I1_0),.din(w_dff_A_XzwxnOKp0_0),.clk(gclk));
	jdff dff_A_FHuc58tC3_1(.dout(w_G8gat_0[1]),.din(w_dff_A_FHuc58tC3_1),.clk(gclk));
	jdff dff_A_vihw9c6K3_1(.dout(w_dff_A_FHuc58tC3_1),.din(w_dff_A_vihw9c6K3_1),.clk(gclk));
	jdff dff_A_0LU4okXJ3_1(.dout(w_dff_A_vihw9c6K3_1),.din(w_dff_A_0LU4okXJ3_1),.clk(gclk));
	jdff dff_A_tslWGU1S1_1(.dout(w_dff_A_0LU4okXJ3_1),.din(w_dff_A_tslWGU1S1_1),.clk(gclk));
	jdff dff_A_s4Ani3Gk5_1(.dout(w_dff_A_tslWGU1S1_1),.din(w_dff_A_s4Ani3Gk5_1),.clk(gclk));
	jdff dff_A_qZV14EGE8_1(.dout(w_dff_A_s4Ani3Gk5_1),.din(w_dff_A_qZV14EGE8_1),.clk(gclk));
	jdff dff_A_VfnyHQxD8_1(.dout(w_dff_A_qZV14EGE8_1),.din(w_dff_A_VfnyHQxD8_1),.clk(gclk));
	jdff dff_A_kD7MLEVY8_1(.dout(w_dff_A_VfnyHQxD8_1),.din(w_dff_A_kD7MLEVY8_1),.clk(gclk));
	jdff dff_A_QDLByZa57_0(.dout(w_n170_0[0]),.din(w_dff_A_QDLByZa57_0),.clk(gclk));
	jdff dff_A_BSgXFtMW4_0(.dout(w_dff_A_QDLByZa57_0),.din(w_dff_A_BSgXFtMW4_0),.clk(gclk));
	jdff dff_A_7CAeB6Wl0_0(.dout(w_dff_A_BSgXFtMW4_0),.din(w_dff_A_7CAeB6Wl0_0),.clk(gclk));
	jdff dff_A_6gHQvYU45_0(.dout(w_dff_A_7CAeB6Wl0_0),.din(w_dff_A_6gHQvYU45_0),.clk(gclk));
	jdff dff_A_gi9H9yxK9_0(.dout(w_dff_A_6gHQvYU45_0),.din(w_dff_A_gi9H9yxK9_0),.clk(gclk));
	jdff dff_A_SkawIwLd5_0(.dout(w_dff_A_gi9H9yxK9_0),.din(w_dff_A_SkawIwLd5_0),.clk(gclk));
	jdff dff_A_R2gKMqU40_0(.dout(w_G86gat_0[0]),.din(w_dff_A_R2gKMqU40_0),.clk(gclk));
	jdff dff_A_JG3Heh8G4_0(.dout(w_dff_A_R2gKMqU40_0),.din(w_dff_A_JG3Heh8G4_0),.clk(gclk));
	jdff dff_A_Y6eOtt9B1_0(.dout(w_dff_A_JG3Heh8G4_0),.din(w_dff_A_Y6eOtt9B1_0),.clk(gclk));
	jdff dff_A_eF8DZN3L3_0(.dout(w_dff_A_Y6eOtt9B1_0),.din(w_dff_A_eF8DZN3L3_0),.clk(gclk));
	jdff dff_A_6YCfdz0H4_0(.dout(w_dff_A_eF8DZN3L3_0),.din(w_dff_A_6YCfdz0H4_0),.clk(gclk));
	jdff dff_A_Yv0B43UV0_0(.dout(w_dff_A_6YCfdz0H4_0),.din(w_dff_A_Yv0B43UV0_0),.clk(gclk));
	jdff dff_A_KLS6JTbl0_0(.dout(w_dff_A_Yv0B43UV0_0),.din(w_dff_A_KLS6JTbl0_0),.clk(gclk));
	jdff dff_A_NH9UMk1G5_0(.dout(w_dff_A_KLS6JTbl0_0),.din(w_dff_A_NH9UMk1G5_0),.clk(gclk));
	jdff dff_A_hBBQgif57_0(.dout(w_dff_A_NH9UMk1G5_0),.din(w_dff_A_hBBQgif57_0),.clk(gclk));
	jdff dff_A_lmmQJEJx9_0(.dout(w_dff_A_hBBQgif57_0),.din(w_dff_A_lmmQJEJx9_0),.clk(gclk));
	jdff dff_A_p1brhldv6_0(.dout(w_dff_A_lmmQJEJx9_0),.din(w_dff_A_p1brhldv6_0),.clk(gclk));
	jdff dff_A_rNRGTngr3_0(.dout(w_dff_A_p1brhldv6_0),.din(w_dff_A_rNRGTngr3_0),.clk(gclk));
	jdff dff_A_KrUqlXWO1_0(.dout(w_dff_A_rNRGTngr3_0),.din(w_dff_A_KrUqlXWO1_0),.clk(gclk));
	jdff dff_A_lG4fbDm27_1(.dout(w_G86gat_0[1]),.din(w_dff_A_lG4fbDm27_1),.clk(gclk));
	jdff dff_A_AaH5f4xM2_1(.dout(w_dff_A_lG4fbDm27_1),.din(w_dff_A_AaH5f4xM2_1),.clk(gclk));
	jdff dff_A_c59gx8zd7_1(.dout(w_dff_A_AaH5f4xM2_1),.din(w_dff_A_c59gx8zd7_1),.clk(gclk));
	jdff dff_A_PnsqMdEa7_1(.dout(w_dff_A_c59gx8zd7_1),.din(w_dff_A_PnsqMdEa7_1),.clk(gclk));
	jdff dff_A_8F9UQrgo7_1(.dout(w_dff_A_PnsqMdEa7_1),.din(w_dff_A_8F9UQrgo7_1),.clk(gclk));
	jdff dff_A_FHIs6XF06_1(.dout(w_dff_A_8F9UQrgo7_1),.din(w_dff_A_FHIs6XF06_1),.clk(gclk));
	jdff dff_A_vsBdrI9I9_1(.dout(w_dff_A_FHIs6XF06_1),.din(w_dff_A_vsBdrI9I9_1),.clk(gclk));
	jdff dff_A_L69zbemZ6_1(.dout(w_dff_A_vsBdrI9I9_1),.din(w_dff_A_L69zbemZ6_1),.clk(gclk));
	jdff dff_A_yKJPnWMB9_1(.dout(w_n120_0[1]),.din(w_dff_A_yKJPnWMB9_1),.clk(gclk));
	jdff dff_A_3ADpAWyi0_1(.dout(w_dff_A_yKJPnWMB9_1),.din(w_dff_A_3ADpAWyi0_1),.clk(gclk));
	jdff dff_A_oNCdNQzd2_1(.dout(w_n119_0[1]),.din(w_dff_A_oNCdNQzd2_1),.clk(gclk));
	jdff dff_A_oZE6wGQp2_1(.dout(w_dff_A_oNCdNQzd2_1),.din(w_dff_A_oZE6wGQp2_1),.clk(gclk));
	jdff dff_A_L0rw6R8r0_1(.dout(w_dff_A_oZE6wGQp2_1),.din(w_dff_A_L0rw6R8r0_1),.clk(gclk));
	jdff dff_A_K1wdPRtT1_1(.dout(w_dff_A_L0rw6R8r0_1),.din(w_dff_A_K1wdPRtT1_1),.clk(gclk));
	jdff dff_A_JkqTa2vl0_1(.dout(w_dff_A_K1wdPRtT1_1),.din(w_dff_A_JkqTa2vl0_1),.clk(gclk));
	jdff dff_A_IiKOOlhv4_1(.dout(w_dff_A_JkqTa2vl0_1),.din(w_dff_A_IiKOOlhv4_1),.clk(gclk));
	jdff dff_A_QZk5PW4p2_0(.dout(w_n117_0[0]),.din(w_dff_A_QZk5PW4p2_0),.clk(gclk));
	jdff dff_A_EO0z2ifm0_0(.dout(w_dff_A_QZk5PW4p2_0),.din(w_dff_A_EO0z2ifm0_0),.clk(gclk));
	jdff dff_A_uMldxBtI8_0(.dout(w_dff_A_EO0z2ifm0_0),.din(w_dff_A_uMldxBtI8_0),.clk(gclk));
	jdff dff_A_arf4bEHa4_0(.dout(w_dff_A_uMldxBtI8_0),.din(w_dff_A_arf4bEHa4_0),.clk(gclk));
	jdff dff_A_JvWzoQW80_0(.dout(w_dff_A_arf4bEHa4_0),.din(w_dff_A_JvWzoQW80_0),.clk(gclk));
	jdff dff_B_F0JguZzJ5_2(.din(n117),.dout(w_dff_B_F0JguZzJ5_2),.clk(gclk));
	jdff dff_B_m3dJybvj1_2(.din(w_dff_B_F0JguZzJ5_2),.dout(w_dff_B_m3dJybvj1_2),.clk(gclk));
	jdff dff_B_e7g7yZtB6_2(.din(w_dff_B_m3dJybvj1_2),.dout(w_dff_B_e7g7yZtB6_2),.clk(gclk));
	jdff dff_B_asvh0jIs2_2(.din(w_dff_B_e7g7yZtB6_2),.dout(w_dff_B_asvh0jIs2_2),.clk(gclk));
	jdff dff_B_vspyw1L60_2(.din(w_dff_B_asvh0jIs2_2),.dout(w_dff_B_vspyw1L60_2),.clk(gclk));
	jdff dff_B_ulGm0nvv1_2(.din(w_dff_B_vspyw1L60_2),.dout(w_dff_B_ulGm0nvv1_2),.clk(gclk));
	jdff dff_B_WmSvZ7f01_2(.din(w_dff_B_ulGm0nvv1_2),.dout(w_dff_B_WmSvZ7f01_2),.clk(gclk));
	jdff dff_A_mzHtWNOf6_0(.dout(w_G60gat_0[0]),.din(w_dff_A_mzHtWNOf6_0),.clk(gclk));
	jdff dff_A_nvkOzMxY0_0(.dout(w_dff_A_mzHtWNOf6_0),.din(w_dff_A_nvkOzMxY0_0),.clk(gclk));
	jdff dff_A_6KASFCUD7_0(.dout(w_dff_A_nvkOzMxY0_0),.din(w_dff_A_6KASFCUD7_0),.clk(gclk));
	jdff dff_A_IYPetPUa0_0(.dout(w_dff_A_6KASFCUD7_0),.din(w_dff_A_IYPetPUa0_0),.clk(gclk));
	jdff dff_A_AM18Ao5n8_0(.dout(w_dff_A_IYPetPUa0_0),.din(w_dff_A_AM18Ao5n8_0),.clk(gclk));
	jdff dff_A_hpFyGLSH4_0(.dout(w_dff_A_AM18Ao5n8_0),.din(w_dff_A_hpFyGLSH4_0),.clk(gclk));
	jdff dff_A_ntwLmnvx3_0(.dout(w_dff_A_hpFyGLSH4_0),.din(w_dff_A_ntwLmnvx3_0),.clk(gclk));
	jdff dff_A_tQwx1AAg8_0(.dout(w_dff_A_ntwLmnvx3_0),.din(w_dff_A_tQwx1AAg8_0),.clk(gclk));
	jdff dff_A_SN515lfE4_0(.dout(w_dff_A_tQwx1AAg8_0),.din(w_dff_A_SN515lfE4_0),.clk(gclk));
	jdff dff_A_qfXVdmSh4_0(.dout(w_dff_A_SN515lfE4_0),.din(w_dff_A_qfXVdmSh4_0),.clk(gclk));
	jdff dff_A_m4TbpFLn5_0(.dout(w_dff_A_qfXVdmSh4_0),.din(w_dff_A_m4TbpFLn5_0),.clk(gclk));
	jdff dff_A_ZY1y03VH3_0(.dout(w_dff_A_m4TbpFLn5_0),.din(w_dff_A_ZY1y03VH3_0),.clk(gclk));
	jdff dff_A_NKLuK1yq9_0(.dout(w_dff_A_ZY1y03VH3_0),.din(w_dff_A_NKLuK1yq9_0),.clk(gclk));
	jdff dff_B_je38FjIa0_1(.din(n154),.dout(w_dff_B_je38FjIa0_1),.clk(gclk));
	jdff dff_B_322Gjxrg7_0(.din(n165),.dout(w_dff_B_322Gjxrg7_0),.clk(gclk));
	jdff dff_A_t04fUksS7_0(.dout(w_n164_0[0]),.din(w_dff_A_t04fUksS7_0),.clk(gclk));
	jdff dff_A_o2uHKknx3_0(.dout(w_dff_A_t04fUksS7_0),.din(w_dff_A_o2uHKknx3_0),.clk(gclk));
	jdff dff_A_qQTO3HbX5_0(.dout(w_dff_A_o2uHKknx3_0),.din(w_dff_A_qQTO3HbX5_0),.clk(gclk));
	jdff dff_A_x4HZyByn8_0(.dout(w_dff_A_qQTO3HbX5_0),.din(w_dff_A_x4HZyByn8_0),.clk(gclk));
	jdff dff_A_NczRzFiI9_0(.dout(w_dff_A_x4HZyByn8_0),.din(w_dff_A_NczRzFiI9_0),.clk(gclk));
	jdff dff_A_KIgzyAMf8_0(.dout(w_dff_A_NczRzFiI9_0),.din(w_dff_A_KIgzyAMf8_0),.clk(gclk));
	jdff dff_B_dDO3Yzt54_1(.din(n162),.dout(w_dff_B_dDO3Yzt54_1),.clk(gclk));
	jdff dff_B_hw3qssex4_1(.din(w_dff_B_dDO3Yzt54_1),.dout(w_dff_B_hw3qssex4_1),.clk(gclk));
	jdff dff_B_NMbbV1YO5_1(.din(w_dff_B_hw3qssex4_1),.dout(w_dff_B_NMbbV1YO5_1),.clk(gclk));
	jdff dff_B_1lcgFhYH1_1(.din(w_dff_B_NMbbV1YO5_1),.dout(w_dff_B_1lcgFhYH1_1),.clk(gclk));
	jdff dff_B_ppddoFWA0_1(.din(w_dff_B_1lcgFhYH1_1),.dout(w_dff_B_ppddoFWA0_1),.clk(gclk));
	jdff dff_B_bG9ClS3E6_1(.din(w_dff_B_ppddoFWA0_1),.dout(w_dff_B_bG9ClS3E6_1),.clk(gclk));
	jdff dff_A_A5pOeaCf2_0(.dout(w_G112gat_0[0]),.din(w_dff_A_A5pOeaCf2_0),.clk(gclk));
	jdff dff_A_pQNcgboV1_0(.dout(w_dff_A_A5pOeaCf2_0),.din(w_dff_A_pQNcgboV1_0),.clk(gclk));
	jdff dff_A_ZOHyfuig1_0(.dout(w_dff_A_pQNcgboV1_0),.din(w_dff_A_ZOHyfuig1_0),.clk(gclk));
	jdff dff_A_CNUZ71yK0_0(.dout(w_dff_A_ZOHyfuig1_0),.din(w_dff_A_CNUZ71yK0_0),.clk(gclk));
	jdff dff_A_rYrtoSBl9_0(.dout(w_dff_A_CNUZ71yK0_0),.din(w_dff_A_rYrtoSBl9_0),.clk(gclk));
	jdff dff_A_NNo3Tlci1_0(.dout(w_dff_A_rYrtoSBl9_0),.din(w_dff_A_NNo3Tlci1_0),.clk(gclk));
	jdff dff_A_h2Y9ZJzD2_0(.dout(w_dff_A_NNo3Tlci1_0),.din(w_dff_A_h2Y9ZJzD2_0),.clk(gclk));
	jdff dff_A_o85ay8Vw5_0(.dout(w_dff_A_h2Y9ZJzD2_0),.din(w_dff_A_o85ay8Vw5_0),.clk(gclk));
	jdff dff_A_wefd0r991_0(.dout(w_dff_A_o85ay8Vw5_0),.din(w_dff_A_wefd0r991_0),.clk(gclk));
	jdff dff_A_Pts60yJD2_0(.dout(w_dff_A_wefd0r991_0),.din(w_dff_A_Pts60yJD2_0),.clk(gclk));
	jdff dff_A_mAKc8hN59_0(.dout(w_dff_A_Pts60yJD2_0),.din(w_dff_A_mAKc8hN59_0),.clk(gclk));
	jdff dff_A_fP25fRNS7_0(.dout(w_dff_A_mAKc8hN59_0),.din(w_dff_A_fP25fRNS7_0),.clk(gclk));
	jdff dff_A_l6NYPA6D1_0(.dout(w_dff_A_fP25fRNS7_0),.din(w_dff_A_l6NYPA6D1_0),.clk(gclk));
	jdff dff_A_GfC7Bp2N2_1(.dout(w_G112gat_0[1]),.din(w_dff_A_GfC7Bp2N2_1),.clk(gclk));
	jdff dff_A_YVj5YIYD5_1(.dout(w_dff_A_GfC7Bp2N2_1),.din(w_dff_A_YVj5YIYD5_1),.clk(gclk));
	jdff dff_A_NeWIEbjl9_1(.dout(w_dff_A_YVj5YIYD5_1),.din(w_dff_A_NeWIEbjl9_1),.clk(gclk));
	jdff dff_A_FgzBJMXg7_1(.dout(w_dff_A_NeWIEbjl9_1),.din(w_dff_A_FgzBJMXg7_1),.clk(gclk));
	jdff dff_A_yKc3S2P46_1(.dout(w_dff_A_FgzBJMXg7_1),.din(w_dff_A_yKc3S2P46_1),.clk(gclk));
	jdff dff_A_0ckAmdGe6_1(.dout(w_dff_A_yKc3S2P46_1),.din(w_dff_A_0ckAmdGe6_1),.clk(gclk));
	jdff dff_A_NU9uRoma3_1(.dout(w_dff_A_0ckAmdGe6_1),.din(w_dff_A_NU9uRoma3_1),.clk(gclk));
	jdff dff_A_tqBIb0nN5_1(.dout(w_dff_A_NU9uRoma3_1),.din(w_dff_A_tqBIb0nN5_1),.clk(gclk));
	jdff dff_A_dJOGWLWu1_0(.dout(w_n159_0[0]),.din(w_dff_A_dJOGWLWu1_0),.clk(gclk));
	jdff dff_A_eeH93Aek3_0(.dout(w_dff_A_dJOGWLWu1_0),.din(w_dff_A_eeH93Aek3_0),.clk(gclk));
	jdff dff_A_7vuqptF97_0(.dout(w_dff_A_eeH93Aek3_0),.din(w_dff_A_7vuqptF97_0),.clk(gclk));
	jdff dff_A_6EfTsEgy0_0(.dout(w_dff_A_7vuqptF97_0),.din(w_dff_A_6EfTsEgy0_0),.clk(gclk));
	jdff dff_A_4Io0qKV22_0(.dout(w_dff_A_6EfTsEgy0_0),.din(w_dff_A_4Io0qKV22_0),.clk(gclk));
	jdff dff_A_Hpp4eHyo1_0(.dout(w_dff_A_4Io0qKV22_0),.din(w_dff_A_Hpp4eHyo1_0),.clk(gclk));
	jdff dff_A_2MCyHMoD3_0(.dout(w_G34gat_0[0]),.din(w_dff_A_2MCyHMoD3_0),.clk(gclk));
	jdff dff_A_zGokofoE6_0(.dout(w_dff_A_2MCyHMoD3_0),.din(w_dff_A_zGokofoE6_0),.clk(gclk));
	jdff dff_A_cj9R3qHv7_0(.dout(w_dff_A_zGokofoE6_0),.din(w_dff_A_cj9R3qHv7_0),.clk(gclk));
	jdff dff_A_bK50tSnb9_0(.dout(w_dff_A_cj9R3qHv7_0),.din(w_dff_A_bK50tSnb9_0),.clk(gclk));
	jdff dff_A_bQ0gpzmo7_0(.dout(w_dff_A_bK50tSnb9_0),.din(w_dff_A_bQ0gpzmo7_0),.clk(gclk));
	jdff dff_A_tmxd6p482_0(.dout(w_dff_A_bQ0gpzmo7_0),.din(w_dff_A_tmxd6p482_0),.clk(gclk));
	jdff dff_A_14R76Bzs5_0(.dout(w_dff_A_tmxd6p482_0),.din(w_dff_A_14R76Bzs5_0),.clk(gclk));
	jdff dff_A_dUG3WhLy4_0(.dout(w_dff_A_14R76Bzs5_0),.din(w_dff_A_dUG3WhLy4_0),.clk(gclk));
	jdff dff_A_kR7ACrt62_0(.dout(w_dff_A_dUG3WhLy4_0),.din(w_dff_A_kR7ACrt62_0),.clk(gclk));
	jdff dff_A_yYWLwLlL7_0(.dout(w_dff_A_kR7ACrt62_0),.din(w_dff_A_yYWLwLlL7_0),.clk(gclk));
	jdff dff_A_qXerH0iI8_0(.dout(w_dff_A_yYWLwLlL7_0),.din(w_dff_A_qXerH0iI8_0),.clk(gclk));
	jdff dff_A_MoqWAgef6_0(.dout(w_dff_A_qXerH0iI8_0),.din(w_dff_A_MoqWAgef6_0),.clk(gclk));
	jdff dff_A_WxwdJJR06_0(.dout(w_dff_A_MoqWAgef6_0),.din(w_dff_A_WxwdJJR06_0),.clk(gclk));
	jdff dff_A_zwgpQTjc8_1(.dout(w_G34gat_0[1]),.din(w_dff_A_zwgpQTjc8_1),.clk(gclk));
	jdff dff_A_pJ75RshI2_1(.dout(w_dff_A_zwgpQTjc8_1),.din(w_dff_A_pJ75RshI2_1),.clk(gclk));
	jdff dff_A_EWEHM0VO0_1(.dout(w_dff_A_pJ75RshI2_1),.din(w_dff_A_EWEHM0VO0_1),.clk(gclk));
	jdff dff_A_GHSz4eE30_1(.dout(w_dff_A_EWEHM0VO0_1),.din(w_dff_A_GHSz4eE30_1),.clk(gclk));
	jdff dff_A_I7mCkaqp6_1(.dout(w_dff_A_GHSz4eE30_1),.din(w_dff_A_I7mCkaqp6_1),.clk(gclk));
	jdff dff_A_UFtWY4da2_1(.dout(w_dff_A_I7mCkaqp6_1),.din(w_dff_A_UFtWY4da2_1),.clk(gclk));
	jdff dff_A_gOOdI2ru9_1(.dout(w_dff_A_UFtWY4da2_1),.din(w_dff_A_gOOdI2ru9_1),.clk(gclk));
	jdff dff_A_KVLsXlA68_1(.dout(w_dff_A_gOOdI2ru9_1),.din(w_dff_A_KVLsXlA68_1),.clk(gclk));
	jdff dff_A_tSNHuSQF0_0(.dout(w_n156_0[0]),.din(w_dff_A_tSNHuSQF0_0),.clk(gclk));
	jdff dff_A_73BhENhZ9_0(.dout(w_dff_A_tSNHuSQF0_0),.din(w_dff_A_73BhENhZ9_0),.clk(gclk));
	jdff dff_A_evqLtQAD5_0(.dout(w_dff_A_73BhENhZ9_0),.din(w_dff_A_evqLtQAD5_0),.clk(gclk));
	jdff dff_A_e44ds8NR4_0(.dout(w_dff_A_evqLtQAD5_0),.din(w_dff_A_e44ds8NR4_0),.clk(gclk));
	jdff dff_A_sHaAYpWX2_0(.dout(w_dff_A_e44ds8NR4_0),.din(w_dff_A_sHaAYpWX2_0),.clk(gclk));
	jdff dff_A_IB1VLXnM4_0(.dout(w_dff_A_sHaAYpWX2_0),.din(w_dff_A_IB1VLXnM4_0),.clk(gclk));
	jdff dff_A_Zwvh3ak07_1(.dout(w_n138_0[1]),.din(w_dff_A_Zwvh3ak07_1),.clk(gclk));
	jdff dff_A_OVs73K2D2_1(.dout(w_dff_A_Zwvh3ak07_1),.din(w_dff_A_OVs73K2D2_1),.clk(gclk));
	jdff dff_A_X67GF4lf1_1(.dout(w_dff_A_OVs73K2D2_1),.din(w_dff_A_X67GF4lf1_1),.clk(gclk));
	jdff dff_A_6sKgfne63_1(.dout(w_dff_A_X67GF4lf1_1),.din(w_dff_A_6sKgfne63_1),.clk(gclk));
	jdff dff_A_fmbGG5rq0_1(.dout(w_dff_A_6sKgfne63_1),.din(w_dff_A_fmbGG5rq0_1),.clk(gclk));
	jdff dff_A_0h4uRpNu1_1(.dout(w_dff_A_fmbGG5rq0_1),.din(w_dff_A_0h4uRpNu1_1),.clk(gclk));
	jdff dff_A_xVbnUlJz2_0(.dout(w_G99gat_0[0]),.din(w_dff_A_xVbnUlJz2_0),.clk(gclk));
	jdff dff_A_ZEWq0X020_0(.dout(w_dff_A_xVbnUlJz2_0),.din(w_dff_A_ZEWq0X020_0),.clk(gclk));
	jdff dff_A_lrmNfJTA2_0(.dout(w_dff_A_ZEWq0X020_0),.din(w_dff_A_lrmNfJTA2_0),.clk(gclk));
	jdff dff_A_6bJhwbl34_0(.dout(w_dff_A_lrmNfJTA2_0),.din(w_dff_A_6bJhwbl34_0),.clk(gclk));
	jdff dff_A_HnTWAOgu1_0(.dout(w_dff_A_6bJhwbl34_0),.din(w_dff_A_HnTWAOgu1_0),.clk(gclk));
	jdff dff_A_pEGBuJJz2_0(.dout(w_dff_A_HnTWAOgu1_0),.din(w_dff_A_pEGBuJJz2_0),.clk(gclk));
	jdff dff_A_rx6gk8z21_0(.dout(w_dff_A_pEGBuJJz2_0),.din(w_dff_A_rx6gk8z21_0),.clk(gclk));
	jdff dff_A_lQ3WEhM69_0(.dout(w_dff_A_rx6gk8z21_0),.din(w_dff_A_lQ3WEhM69_0),.clk(gclk));
	jdff dff_A_qGFULiEO4_1(.dout(w_G99gat_0[1]),.din(w_dff_A_qGFULiEO4_1),.clk(gclk));
	jdff dff_A_TAST8Uue5_1(.dout(w_dff_A_qGFULiEO4_1),.din(w_dff_A_TAST8Uue5_1),.clk(gclk));
	jdff dff_A_v2sdafcS2_1(.dout(w_dff_A_TAST8Uue5_1),.din(w_dff_A_v2sdafcS2_1),.clk(gclk));
	jdff dff_A_TNGkTsMo6_1(.dout(w_dff_A_v2sdafcS2_1),.din(w_dff_A_TNGkTsMo6_1),.clk(gclk));
	jdff dff_A_ugHHWuQG4_1(.dout(w_dff_A_TNGkTsMo6_1),.din(w_dff_A_ugHHWuQG4_1),.clk(gclk));
	jdff dff_A_nlXoKio41_1(.dout(w_dff_A_ugHHWuQG4_1),.din(w_dff_A_nlXoKio41_1),.clk(gclk));
	jdff dff_A_s4aL91iV2_1(.dout(w_dff_A_nlXoKio41_1),.din(w_dff_A_s4aL91iV2_1),.clk(gclk));
	jdff dff_A_t7842EW06_1(.dout(w_dff_A_s4aL91iV2_1),.din(w_dff_A_t7842EW06_1),.clk(gclk));
	jdff dff_A_vACIrymr1_1(.dout(w_dff_A_t7842EW06_1),.din(w_dff_A_vACIrymr1_1),.clk(gclk));
	jdff dff_A_GI8wvvPZ6_1(.dout(w_dff_A_vACIrymr1_1),.din(w_dff_A_GI8wvvPZ6_1),.clk(gclk));
	jdff dff_A_jynH119r0_1(.dout(w_dff_A_GI8wvvPZ6_1),.din(w_dff_A_jynH119r0_1),.clk(gclk));
	jdff dff_A_Na2a7yxM4_1(.dout(w_dff_A_jynH119r0_1),.din(w_dff_A_Na2a7yxM4_1),.clk(gclk));
	jdff dff_A_SJ41GHkM6_1(.dout(w_dff_A_Na2a7yxM4_1),.din(w_dff_A_SJ41GHkM6_1),.clk(gclk));
	jdff dff_A_GZjtroyw6_0(.dout(w_n151_0[0]),.din(w_dff_A_GZjtroyw6_0),.clk(gclk));
	jdff dff_A_gBvb6wRA4_0(.dout(w_dff_A_GZjtroyw6_0),.din(w_dff_A_gBvb6wRA4_0),.clk(gclk));
	jdff dff_A_UtLjcSU38_0(.dout(w_dff_A_gBvb6wRA4_0),.din(w_dff_A_UtLjcSU38_0),.clk(gclk));
	jdff dff_A_SmABoodp9_0(.dout(w_dff_A_UtLjcSU38_0),.din(w_dff_A_SmABoodp9_0),.clk(gclk));
	jdff dff_A_ZxKtvrd09_0(.dout(w_dff_A_SmABoodp9_0),.din(w_dff_A_ZxKtvrd09_0),.clk(gclk));
	jdff dff_A_LzcbsiGM9_0(.dout(w_dff_A_ZxKtvrd09_0),.din(w_dff_A_LzcbsiGM9_0),.clk(gclk));
	jdff dff_B_oFHjK9Vy2_1(.din(n48),.dout(w_dff_B_oFHjK9Vy2_1),.clk(gclk));
	jdff dff_B_uy7Ipox02_1(.din(n61),.dout(w_dff_B_uy7Ipox02_1),.clk(gclk));
	jdff dff_A_8vpAUUyx1_0(.dout(w_n64_0[0]),.din(w_dff_A_8vpAUUyx1_0),.clk(gclk));
	jdff dff_A_rVlhmgEL9_0(.dout(w_dff_A_8vpAUUyx1_0),.din(w_dff_A_rVlhmgEL9_0),.clk(gclk));
	jdff dff_A_3ZJcno1i2_0(.dout(w_dff_A_rVlhmgEL9_0),.din(w_dff_A_3ZJcno1i2_0),.clk(gclk));
	jdff dff_A_blzEouPS7_0(.dout(w_dff_A_3ZJcno1i2_0),.din(w_dff_A_blzEouPS7_0),.clk(gclk));
	jdff dff_A_LdfUle2X1_0(.dout(w_dff_A_blzEouPS7_0),.din(w_dff_A_LdfUle2X1_0),.clk(gclk));
	jdff dff_A_wktOnP1n7_0(.dout(w_n62_0[0]),.din(w_dff_A_wktOnP1n7_0),.clk(gclk));
	jdff dff_A_23rckZjR5_0(.dout(w_dff_A_wktOnP1n7_0),.din(w_dff_A_23rckZjR5_0),.clk(gclk));
	jdff dff_A_DGM5D3ml6_0(.dout(w_dff_A_23rckZjR5_0),.din(w_dff_A_DGM5D3ml6_0),.clk(gclk));
	jdff dff_A_7tjp1Vyz8_0(.dout(w_dff_A_DGM5D3ml6_0),.din(w_dff_A_7tjp1Vyz8_0),.clk(gclk));
	jdff dff_A_8L0BALgF9_0(.dout(w_dff_A_7tjp1Vyz8_0),.din(w_dff_A_8L0BALgF9_0),.clk(gclk));
	jdff dff_A_v1P0GAct8_0(.dout(w_n60_0[0]),.din(w_dff_A_v1P0GAct8_0),.clk(gclk));
	jdff dff_A_EQDqglJl5_0(.dout(w_dff_A_v1P0GAct8_0),.din(w_dff_A_EQDqglJl5_0),.clk(gclk));
	jdff dff_A_9dS6k8xR5_0(.dout(w_dff_A_EQDqglJl5_0),.din(w_dff_A_9dS6k8xR5_0),.clk(gclk));
	jdff dff_A_4Ne3XgsQ3_0(.dout(w_dff_A_9dS6k8xR5_0),.din(w_dff_A_4Ne3XgsQ3_0),.clk(gclk));
	jdff dff_A_dfHDav1S5_0(.dout(w_dff_A_4Ne3XgsQ3_0),.din(w_dff_A_dfHDav1S5_0),.clk(gclk));
	jdff dff_A_qsYE7pvN0_0(.dout(w_n57_0[0]),.din(w_dff_A_qsYE7pvN0_0),.clk(gclk));
	jdff dff_A_k0qdTbHE4_0(.dout(w_dff_A_qsYE7pvN0_0),.din(w_dff_A_k0qdTbHE4_0),.clk(gclk));
	jdff dff_A_8wKpf4oa0_0(.dout(w_dff_A_k0qdTbHE4_0),.din(w_dff_A_8wKpf4oa0_0),.clk(gclk));
	jdff dff_A_lHlGuDJ27_0(.dout(w_dff_A_8wKpf4oa0_0),.din(w_dff_A_lHlGuDJ27_0),.clk(gclk));
	jdff dff_A_QnNiPzO00_0(.dout(w_n54_0[0]),.din(w_dff_A_QnNiPzO00_0),.clk(gclk));
	jdff dff_A_mDmrsqG29_0(.dout(w_dff_A_QnNiPzO00_0),.din(w_dff_A_mDmrsqG29_0),.clk(gclk));
	jdff dff_A_7Wkvu69p4_0(.dout(w_dff_A_mDmrsqG29_0),.din(w_dff_A_7Wkvu69p4_0),.clk(gclk));
	jdff dff_A_wbAVqUWU0_0(.dout(w_dff_A_7Wkvu69p4_0),.din(w_dff_A_wbAVqUWU0_0),.clk(gclk));
	jdff dff_A_1RKxfJyf4_0(.dout(w_dff_A_wbAVqUWU0_0),.din(w_dff_A_1RKxfJyf4_0),.clk(gclk));
	jdff dff_A_nEZUbuOp2_0(.dout(w_n51_0[0]),.din(w_dff_A_nEZUbuOp2_0),.clk(gclk));
	jdff dff_A_4azKf7PR2_0(.dout(w_dff_A_nEZUbuOp2_0),.din(w_dff_A_4azKf7PR2_0),.clk(gclk));
	jdff dff_A_2z0aG76x2_0(.dout(w_dff_A_4azKf7PR2_0),.din(w_dff_A_2z0aG76x2_0),.clk(gclk));
	jdff dff_A_u22NVl2Z9_0(.dout(w_dff_A_2z0aG76x2_0),.din(w_dff_A_u22NVl2Z9_0),.clk(gclk));
	jdff dff_A_OD6Iv26o4_0(.dout(w_dff_A_u22NVl2Z9_0),.din(w_dff_A_OD6Iv26o4_0),.clk(gclk));
	jdff dff_A_IToyDlht6_0(.dout(w_n47_0[0]),.din(w_dff_A_IToyDlht6_0),.clk(gclk));
	jdff dff_A_Z8kEapOt6_0(.dout(w_dff_A_IToyDlht6_0),.din(w_dff_A_Z8kEapOt6_0),.clk(gclk));
	jdff dff_A_kp91eHvW8_0(.dout(w_dff_A_Z8kEapOt6_0),.din(w_dff_A_kp91eHvW8_0),.clk(gclk));
	jdff dff_A_RvKDN4TZ1_0(.dout(w_G21gat_0[0]),.din(w_dff_A_RvKDN4TZ1_0),.clk(gclk));
	jdff dff_A_kkFSYdNl7_0(.dout(w_dff_A_RvKDN4TZ1_0),.din(w_dff_A_kkFSYdNl7_0),.clk(gclk));
	jdff dff_A_Jq7fBqOF2_0(.dout(w_dff_A_kkFSYdNl7_0),.din(w_dff_A_Jq7fBqOF2_0),.clk(gclk));
	jdff dff_A_s5VjoMFf9_0(.dout(w_dff_A_Jq7fBqOF2_0),.din(w_dff_A_s5VjoMFf9_0),.clk(gclk));
	jdff dff_A_2EOcIFN52_0(.dout(w_dff_A_s5VjoMFf9_0),.din(w_dff_A_2EOcIFN52_0),.clk(gclk));
	jdff dff_A_e2SsFd7f5_0(.dout(w_dff_A_2EOcIFN52_0),.din(w_dff_A_e2SsFd7f5_0),.clk(gclk));
	jdff dff_A_jTcb8ZOl1_0(.dout(w_dff_A_e2SsFd7f5_0),.din(w_dff_A_jTcb8ZOl1_0),.clk(gclk));
	jdff dff_A_YBtA6iDe4_0(.dout(w_dff_A_jTcb8ZOl1_0),.din(w_dff_A_YBtA6iDe4_0),.clk(gclk));
	jdff dff_A_Xyt4i8y75_0(.dout(w_dff_A_YBtA6iDe4_0),.din(w_dff_A_Xyt4i8y75_0),.clk(gclk));
	jdff dff_A_fqhsjAks2_0(.dout(w_dff_A_Xyt4i8y75_0),.din(w_dff_A_fqhsjAks2_0),.clk(gclk));
	jdff dff_A_KVWmTdjA8_0(.dout(w_dff_A_fqhsjAks2_0),.din(w_dff_A_KVWmTdjA8_0),.clk(gclk));
	jdff dff_A_kpwza5SJ1_0(.dout(w_dff_A_KVWmTdjA8_0),.din(w_dff_A_kpwza5SJ1_0),.clk(gclk));
	jdff dff_A_ZOOuc7Ci6_0(.dout(w_dff_A_kpwza5SJ1_0),.din(w_dff_A_ZOOuc7Ci6_0),.clk(gclk));
	jdff dff_A_d1rrIRyd8_1(.dout(w_G21gat_0[1]),.din(w_dff_A_d1rrIRyd8_1),.clk(gclk));
	jdff dff_A_yjLcObeY9_1(.dout(w_dff_A_d1rrIRyd8_1),.din(w_dff_A_yjLcObeY9_1),.clk(gclk));
	jdff dff_A_hZcBfOUz8_1(.dout(w_dff_A_yjLcObeY9_1),.din(w_dff_A_hZcBfOUz8_1),.clk(gclk));
	jdff dff_A_u8lwkm4s9_1(.dout(w_dff_A_hZcBfOUz8_1),.din(w_dff_A_u8lwkm4s9_1),.clk(gclk));
	jdff dff_A_hNl5FUOt7_1(.dout(w_dff_A_u8lwkm4s9_1),.din(w_dff_A_hNl5FUOt7_1),.clk(gclk));
	jdff dff_A_uAHsQf6v4_1(.dout(w_dff_A_hNl5FUOt7_1),.din(w_dff_A_uAHsQf6v4_1),.clk(gclk));
	jdff dff_A_SaVx8Hky1_1(.dout(w_dff_A_uAHsQf6v4_1),.din(w_dff_A_SaVx8Hky1_1),.clk(gclk));
	jdff dff_A_QBYLUvGz0_1(.dout(w_dff_A_SaVx8Hky1_1),.din(w_dff_A_QBYLUvGz0_1),.clk(gclk));
	jdff dff_A_LJPjatJ13_0(.dout(w_n102_0[0]),.din(w_dff_A_LJPjatJ13_0),.clk(gclk));
	jdff dff_A_eNBbkTo37_0(.dout(w_dff_A_LJPjatJ13_0),.din(w_dff_A_eNBbkTo37_0),.clk(gclk));
	jdff dff_A_JG7WXW0r9_0(.dout(w_dff_A_eNBbkTo37_0),.din(w_dff_A_JG7WXW0r9_0),.clk(gclk));
	jdff dff_A_0TYQFC2b0_0(.dout(w_dff_A_JG7WXW0r9_0),.din(w_dff_A_0TYQFC2b0_0),.clk(gclk));
	jdff dff_A_wG5NK1E20_0(.dout(w_dff_A_0TYQFC2b0_0),.din(w_dff_A_wG5NK1E20_0),.clk(gclk));
	jdff dff_B_ZMbGXRTG6_2(.din(n102),.dout(w_dff_B_ZMbGXRTG6_2),.clk(gclk));
	jdff dff_B_iUlywCdM6_2(.din(w_dff_B_ZMbGXRTG6_2),.dout(w_dff_B_iUlywCdM6_2),.clk(gclk));
	jdff dff_B_7WNg8MN43_2(.din(w_dff_B_iUlywCdM6_2),.dout(w_dff_B_7WNg8MN43_2),.clk(gclk));
	jdff dff_B_WoxK1Frj3_2(.din(w_dff_B_7WNg8MN43_2),.dout(w_dff_B_WoxK1Frj3_2),.clk(gclk));
	jdff dff_B_YN3ImGOS9_2(.din(w_dff_B_WoxK1Frj3_2),.dout(w_dff_B_YN3ImGOS9_2),.clk(gclk));
	jdff dff_B_hcPfypnS0_2(.din(w_dff_B_YN3ImGOS9_2),.dout(w_dff_B_hcPfypnS0_2),.clk(gclk));
	jdff dff_B_44Sdazhr1_2(.din(w_dff_B_hcPfypnS0_2),.dout(w_dff_B_44Sdazhr1_2),.clk(gclk));
	jdff dff_A_2j5m2UZt0_0(.dout(w_G73gat_0[0]),.din(w_dff_A_2j5m2UZt0_0),.clk(gclk));
	jdff dff_A_cS4Ucj8e9_0(.dout(w_dff_A_2j5m2UZt0_0),.din(w_dff_A_cS4Ucj8e9_0),.clk(gclk));
	jdff dff_A_wKpgph9G5_0(.dout(w_dff_A_cS4Ucj8e9_0),.din(w_dff_A_wKpgph9G5_0),.clk(gclk));
	jdff dff_A_crOzn7BM3_0(.dout(w_dff_A_wKpgph9G5_0),.din(w_dff_A_crOzn7BM3_0),.clk(gclk));
	jdff dff_A_slbOCpSC2_0(.dout(w_dff_A_crOzn7BM3_0),.din(w_dff_A_slbOCpSC2_0),.clk(gclk));
	jdff dff_A_vpWnXkot6_0(.dout(w_dff_A_slbOCpSC2_0),.din(w_dff_A_vpWnXkot6_0),.clk(gclk));
	jdff dff_A_60jqn3kM3_0(.dout(w_dff_A_vpWnXkot6_0),.din(w_dff_A_60jqn3kM3_0),.clk(gclk));
	jdff dff_A_kYfuFxKh5_0(.dout(w_dff_A_60jqn3kM3_0),.din(w_dff_A_kYfuFxKh5_0),.clk(gclk));
	jdff dff_A_xukxow173_0(.dout(w_dff_A_kYfuFxKh5_0),.din(w_dff_A_xukxow173_0),.clk(gclk));
	jdff dff_A_BiqpwgVM3_0(.dout(w_dff_A_xukxow173_0),.din(w_dff_A_BiqpwgVM3_0),.clk(gclk));
	jdff dff_A_onrBnMrm3_0(.dout(w_dff_A_BiqpwgVM3_0),.din(w_dff_A_onrBnMrm3_0),.clk(gclk));
	jdff dff_A_yJgxfflI4_0(.dout(w_dff_A_onrBnMrm3_0),.din(w_dff_A_yJgxfflI4_0),.clk(gclk));
	jdff dff_A_PMAB5Jus3_0(.dout(w_dff_A_yJgxfflI4_0),.din(w_dff_A_PMAB5Jus3_0),.clk(gclk));
	jdff dff_A_hj99hYJI9_1(.dout(w_G73gat_0[1]),.din(w_dff_A_hj99hYJI9_1),.clk(gclk));
	jdff dff_A_nZ1NBaOT1_1(.dout(w_dff_A_hj99hYJI9_1),.din(w_dff_A_nZ1NBaOT1_1),.clk(gclk));
	jdff dff_A_08BxUcFA2_1(.dout(w_dff_A_nZ1NBaOT1_1),.din(w_dff_A_08BxUcFA2_1),.clk(gclk));
	jdff dff_A_bAh2j8pu0_1(.dout(w_dff_A_08BxUcFA2_1),.din(w_dff_A_bAh2j8pu0_1),.clk(gclk));
	jdff dff_A_OemU1Rgk7_1(.dout(w_dff_A_bAh2j8pu0_1),.din(w_dff_A_OemU1Rgk7_1),.clk(gclk));
	jdff dff_A_7w73e4kj4_1(.dout(w_dff_A_OemU1Rgk7_1),.din(w_dff_A_7w73e4kj4_1),.clk(gclk));
	jdff dff_A_pvqPqSX98_1(.dout(w_dff_A_7w73e4kj4_1),.din(w_dff_A_pvqPqSX98_1),.clk(gclk));
	jdff dff_A_vx0g4e2i9_1(.dout(w_dff_A_pvqPqSX98_1),.din(w_dff_A_vx0g4e2i9_1),.clk(gclk));
	jdff dff_A_V9ZXIcU37_0(.dout(w_n104_0[0]),.din(w_dff_A_V9ZXIcU37_0),.clk(gclk));
	jdff dff_A_ZZpuQu4K5_0(.dout(w_dff_A_V9ZXIcU37_0),.din(w_dff_A_ZZpuQu4K5_0),.clk(gclk));
	jdff dff_A_rEmuxZFv2_0(.dout(w_dff_A_ZZpuQu4K5_0),.din(w_dff_A_rEmuxZFv2_0),.clk(gclk));
	jdff dff_A_ku63wcS59_0(.dout(w_dff_A_rEmuxZFv2_0),.din(w_dff_A_ku63wcS59_0),.clk(gclk));
	jdff dff_A_kS8OMkNR1_0(.dout(w_dff_A_ku63wcS59_0),.din(w_dff_A_kS8OMkNR1_0),.clk(gclk));
	jdff dff_A_4YgwA3ay8_0(.dout(w_dff_A_kS8OMkNR1_0),.din(w_dff_A_4YgwA3ay8_0),.clk(gclk));
	jdff dff_B_YfLa0vRk4_1(.din(n72),.dout(w_dff_B_YfLa0vRk4_1),.clk(gclk));
	jdff dff_B_PLZnYOXY2_1(.din(n85),.dout(w_dff_B_PLZnYOXY2_1),.clk(gclk));
	jdff dff_A_Bn9j67c56_0(.dout(w_n88_0[0]),.din(w_dff_A_Bn9j67c56_0),.clk(gclk));
	jdff dff_A_URLQiw6p2_0(.dout(w_dff_A_Bn9j67c56_0),.din(w_dff_A_URLQiw6p2_0),.clk(gclk));
	jdff dff_A_ZpXDOWGU0_0(.dout(w_dff_A_URLQiw6p2_0),.din(w_dff_A_ZpXDOWGU0_0),.clk(gclk));
	jdff dff_A_u0vo2dOR2_0(.dout(w_dff_A_ZpXDOWGU0_0),.din(w_dff_A_u0vo2dOR2_0),.clk(gclk));
	jdff dff_A_cCb31esJ6_0(.dout(w_dff_A_u0vo2dOR2_0),.din(w_dff_A_cCb31esJ6_0),.clk(gclk));
	jdff dff_A_cP0Dv3z61_0(.dout(w_dff_A_cCb31esJ6_0),.din(w_dff_A_cP0Dv3z61_0),.clk(gclk));
	jdff dff_A_dB0buItk9_0(.dout(w_G82gat_0[0]),.din(w_dff_A_dB0buItk9_0),.clk(gclk));
	jdff dff_A_6fK1W0AF1_0(.dout(w_dff_A_dB0buItk9_0),.din(w_dff_A_6fK1W0AF1_0),.clk(gclk));
	jdff dff_A_9QbkHJCp9_0(.dout(w_dff_A_6fK1W0AF1_0),.din(w_dff_A_9QbkHJCp9_0),.clk(gclk));
	jdff dff_A_AP9W7KQp1_0(.dout(w_dff_A_9QbkHJCp9_0),.din(w_dff_A_AP9W7KQp1_0),.clk(gclk));
	jdff dff_A_cqasrydz0_0(.dout(w_dff_A_AP9W7KQp1_0),.din(w_dff_A_cqasrydz0_0),.clk(gclk));
	jdff dff_A_bTT3B0U15_0(.dout(w_dff_A_cqasrydz0_0),.din(w_dff_A_bTT3B0U15_0),.clk(gclk));
	jdff dff_A_RFTucnJE8_0(.dout(w_dff_A_bTT3B0U15_0),.din(w_dff_A_RFTucnJE8_0),.clk(gclk));
	jdff dff_A_hxkmzegh6_2(.dout(w_G82gat_0[2]),.din(w_dff_A_hxkmzegh6_2),.clk(gclk));
	jdff dff_A_60zA4AUF4_0(.dout(w_G76gat_0[0]),.din(w_dff_A_60zA4AUF4_0),.clk(gclk));
	jdff dff_A_UC10F9uH3_0(.dout(w_dff_A_60zA4AUF4_0),.din(w_dff_A_UC10F9uH3_0),.clk(gclk));
	jdff dff_A_vHH5HqRt0_0(.dout(w_dff_A_UC10F9uH3_0),.din(w_dff_A_vHH5HqRt0_0),.clk(gclk));
	jdff dff_A_w6jy9CZx0_0(.dout(w_dff_A_vHH5HqRt0_0),.din(w_dff_A_w6jy9CZx0_0),.clk(gclk));
	jdff dff_A_vZIGNYMV3_0(.dout(w_dff_A_w6jy9CZx0_0),.din(w_dff_A_vZIGNYMV3_0),.clk(gclk));
	jdff dff_A_ywEvo4Ck3_0(.dout(w_dff_A_vZIGNYMV3_0),.din(w_dff_A_ywEvo4Ck3_0),.clk(gclk));
	jdff dff_A_9NmUiCia9_1(.dout(w_G76gat_0[1]),.din(w_dff_A_9NmUiCia9_1),.clk(gclk));
	jdff dff_A_IQ8Cochu7_0(.dout(w_n86_0[0]),.din(w_dff_A_IQ8Cochu7_0),.clk(gclk));
	jdff dff_A_NK2fXNy09_0(.dout(w_dff_A_IQ8Cochu7_0),.din(w_dff_A_NK2fXNy09_0),.clk(gclk));
	jdff dff_A_7So5Ycq72_0(.dout(w_dff_A_NK2fXNy09_0),.din(w_dff_A_7So5Ycq72_0),.clk(gclk));
	jdff dff_A_njPNXPUC9_0(.dout(w_dff_A_7So5Ycq72_0),.din(w_dff_A_njPNXPUC9_0),.clk(gclk));
	jdff dff_A_sSX6e2yF5_0(.dout(w_dff_A_njPNXPUC9_0),.din(w_dff_A_sSX6e2yF5_0),.clk(gclk));
	jdff dff_A_kHTV6ebl3_0(.dout(w_dff_A_sSX6e2yF5_0),.din(w_dff_A_kHTV6ebl3_0),.clk(gclk));
	jdff dff_A_UpOzULii4_0(.dout(w_G95gat_0[0]),.din(w_dff_A_UpOzULii4_0),.clk(gclk));
	jdff dff_A_jw7dUq1X5_0(.dout(w_dff_A_UpOzULii4_0),.din(w_dff_A_jw7dUq1X5_0),.clk(gclk));
	jdff dff_A_YTJkIzR18_0(.dout(w_dff_A_jw7dUq1X5_0),.din(w_dff_A_YTJkIzR18_0),.clk(gclk));
	jdff dff_A_VogTLJuw5_0(.dout(w_dff_A_YTJkIzR18_0),.din(w_dff_A_VogTLJuw5_0),.clk(gclk));
	jdff dff_A_CJvyBEDg6_0(.dout(w_dff_A_VogTLJuw5_0),.din(w_dff_A_CJvyBEDg6_0),.clk(gclk));
	jdff dff_A_d3OR2Mk21_0(.dout(w_dff_A_CJvyBEDg6_0),.din(w_dff_A_d3OR2Mk21_0),.clk(gclk));
	jdff dff_A_k1PxBuxu6_0(.dout(w_dff_A_d3OR2Mk21_0),.din(w_dff_A_k1PxBuxu6_0),.clk(gclk));
	jdff dff_A_TsWW9uRX3_2(.dout(w_G95gat_0[2]),.din(w_dff_A_TsWW9uRX3_2),.clk(gclk));
	jdff dff_A_xj5ZsRTa2_0(.dout(w_G89gat_0[0]),.din(w_dff_A_xj5ZsRTa2_0),.clk(gclk));
	jdff dff_A_lOImutZS3_0(.dout(w_dff_A_xj5ZsRTa2_0),.din(w_dff_A_lOImutZS3_0),.clk(gclk));
	jdff dff_A_DUQ7apof3_0(.dout(w_dff_A_lOImutZS3_0),.din(w_dff_A_DUQ7apof3_0),.clk(gclk));
	jdff dff_A_0xnoinQb8_0(.dout(w_dff_A_DUQ7apof3_0),.din(w_dff_A_0xnoinQb8_0),.clk(gclk));
	jdff dff_A_THf5n9Jx2_0(.dout(w_dff_A_0xnoinQb8_0),.din(w_dff_A_THf5n9Jx2_0),.clk(gclk));
	jdff dff_A_EdeihZfi9_0(.dout(w_dff_A_THf5n9Jx2_0),.din(w_dff_A_EdeihZfi9_0),.clk(gclk));
	jdff dff_A_TxQgQLVW1_1(.dout(w_G89gat_0[1]),.din(w_dff_A_TxQgQLVW1_1),.clk(gclk));
	jdff dff_A_eMg2oYDa2_0(.dout(w_n84_0[0]),.din(w_dff_A_eMg2oYDa2_0),.clk(gclk));
	jdff dff_A_yQOA5XwW1_0(.dout(w_dff_A_eMg2oYDa2_0),.din(w_dff_A_yQOA5XwW1_0),.clk(gclk));
	jdff dff_A_kfhgffsh9_0(.dout(w_dff_A_yQOA5XwW1_0),.din(w_dff_A_kfhgffsh9_0),.clk(gclk));
	jdff dff_A_Wcuqr8lv2_0(.dout(w_dff_A_kfhgffsh9_0),.din(w_dff_A_Wcuqr8lv2_0),.clk(gclk));
	jdff dff_A_vlbRyPbg6_0(.dout(w_dff_A_Wcuqr8lv2_0),.din(w_dff_A_vlbRyPbg6_0),.clk(gclk));
	jdff dff_A_ZT6PXlUK2_0(.dout(w_dff_A_vlbRyPbg6_0),.din(w_dff_A_ZT6PXlUK2_0),.clk(gclk));
	jdff dff_A_SZMwVZMi4_0(.dout(w_G4gat_0[0]),.din(w_dff_A_SZMwVZMi4_0),.clk(gclk));
	jdff dff_A_Eck8mjQ39_0(.dout(w_dff_A_SZMwVZMi4_0),.din(w_dff_A_Eck8mjQ39_0),.clk(gclk));
	jdff dff_A_9FKcUddG1_0(.dout(w_dff_A_Eck8mjQ39_0),.din(w_dff_A_9FKcUddG1_0),.clk(gclk));
	jdff dff_A_UwJK3hhG1_0(.dout(w_dff_A_9FKcUddG1_0),.din(w_dff_A_UwJK3hhG1_0),.clk(gclk));
	jdff dff_A_WFYITHG53_0(.dout(w_dff_A_UwJK3hhG1_0),.din(w_dff_A_WFYITHG53_0),.clk(gclk));
	jdff dff_A_bmvNrT030_0(.dout(w_dff_A_WFYITHG53_0),.din(w_dff_A_bmvNrT030_0),.clk(gclk));
	jdff dff_A_7PR6cJPe7_0(.dout(w_dff_A_bmvNrT030_0),.din(w_dff_A_7PR6cJPe7_0),.clk(gclk));
	jdff dff_A_CvptQvyC1_2(.dout(w_G4gat_0[2]),.din(w_dff_A_CvptQvyC1_2),.clk(gclk));
	jdff dff_A_xAE2yBz56_0(.dout(w_G1gat_0[0]),.din(w_dff_A_xAE2yBz56_0),.clk(gclk));
	jdff dff_A_AY3xOjbm3_0(.dout(w_dff_A_xAE2yBz56_0),.din(w_dff_A_AY3xOjbm3_0),.clk(gclk));
	jdff dff_A_p90pGOqB0_0(.dout(w_dff_A_AY3xOjbm3_0),.din(w_dff_A_p90pGOqB0_0),.clk(gclk));
	jdff dff_A_4WhCyM904_0(.dout(w_dff_A_p90pGOqB0_0),.din(w_dff_A_4WhCyM904_0),.clk(gclk));
	jdff dff_A_TeTrPhwU8_0(.dout(w_dff_A_4WhCyM904_0),.din(w_dff_A_TeTrPhwU8_0),.clk(gclk));
	jdff dff_A_EWXebSuV4_0(.dout(w_dff_A_TeTrPhwU8_0),.din(w_dff_A_EWXebSuV4_0),.clk(gclk));
	jdff dff_A_7wzDnKAk5_1(.dout(w_G1gat_0[1]),.din(w_dff_A_7wzDnKAk5_1),.clk(gclk));
	jdff dff_A_NpKpEWfM1_0(.dout(w_n81_0[0]),.din(w_dff_A_NpKpEWfM1_0),.clk(gclk));
	jdff dff_A_QA7CqL0h7_0(.dout(w_dff_A_NpKpEWfM1_0),.din(w_dff_A_QA7CqL0h7_0),.clk(gclk));
	jdff dff_A_dq4eVbYY9_0(.dout(w_dff_A_QA7CqL0h7_0),.din(w_dff_A_dq4eVbYY9_0),.clk(gclk));
	jdff dff_A_n9TvJP6c8_0(.dout(w_dff_A_dq4eVbYY9_0),.din(w_dff_A_n9TvJP6c8_0),.clk(gclk));
	jdff dff_A_MXoh95nB9_0(.dout(w_n80_0[0]),.din(w_dff_A_MXoh95nB9_0),.clk(gclk));
	jdff dff_A_exi9foQy0_0(.dout(w_dff_A_MXoh95nB9_0),.din(w_dff_A_exi9foQy0_0),.clk(gclk));
	jdff dff_A_Vz87ur456_0(.dout(w_dff_A_exi9foQy0_0),.din(w_dff_A_Vz87ur456_0),.clk(gclk));
	jdff dff_A_RZyyhAbN0_0(.dout(w_dff_A_Vz87ur456_0),.din(w_dff_A_RZyyhAbN0_0),.clk(gclk));
	jdff dff_A_rsUOLE0u5_0(.dout(w_dff_A_RZyyhAbN0_0),.din(w_dff_A_rsUOLE0u5_0),.clk(gclk));
	jdff dff_A_5yNGVIWc8_0(.dout(w_dff_A_rsUOLE0u5_0),.din(w_dff_A_5yNGVIWc8_0),.clk(gclk));
	jdff dff_A_v3c8etSx2_0(.dout(w_dff_A_5yNGVIWc8_0),.din(w_dff_A_v3c8etSx2_0),.clk(gclk));
	jdff dff_A_rQXTpGPf5_0(.dout(w_dff_A_v3c8etSx2_0),.din(w_dff_A_rQXTpGPf5_0),.clk(gclk));
	jdff dff_A_SpSs8p8F2_0(.dout(w_dff_A_rQXTpGPf5_0),.din(w_dff_A_SpSs8p8F2_0),.clk(gclk));
	jdff dff_A_xnFEGC1b9_0(.dout(w_dff_A_SpSs8p8F2_0),.din(w_dff_A_xnFEGC1b9_0),.clk(gclk));
	jdff dff_A_DdSMJzfb4_0(.dout(w_dff_A_xnFEGC1b9_0),.din(w_dff_A_DdSMJzfb4_0),.clk(gclk));
	jdff dff_A_kUH8qIxF8_0(.dout(w_dff_A_DdSMJzfb4_0),.din(w_dff_A_kUH8qIxF8_0),.clk(gclk));
	jdff dff_A_fUx3ADay4_0(.dout(w_dff_A_kUH8qIxF8_0),.din(w_dff_A_fUx3ADay4_0),.clk(gclk));
	jdff dff_A_bihIuxL99_0(.dout(w_dff_A_fUx3ADay4_0),.din(w_dff_A_bihIuxL99_0),.clk(gclk));
	jdff dff_A_QkEetc6U8_0(.dout(w_dff_A_bihIuxL99_0),.din(w_dff_A_QkEetc6U8_0),.clk(gclk));
	jdff dff_A_rRV5Ak2s0_0(.dout(w_dff_A_QkEetc6U8_0),.din(w_dff_A_rRV5Ak2s0_0),.clk(gclk));
	jdff dff_A_hwWOZ2qg2_0(.dout(w_dff_A_rRV5Ak2s0_0),.din(w_dff_A_hwWOZ2qg2_0),.clk(gclk));
	jdff dff_A_Su3yF4Rz7_0(.dout(w_dff_A_hwWOZ2qg2_0),.din(w_dff_A_Su3yF4Rz7_0),.clk(gclk));
	jdff dff_A_IvWgaa469_0(.dout(w_dff_A_Su3yF4Rz7_0),.din(w_dff_A_IvWgaa469_0),.clk(gclk));
	jdff dff_A_fGlpwA8o1_0(.dout(w_dff_A_IvWgaa469_0),.din(w_dff_A_fGlpwA8o1_0),.clk(gclk));
	jdff dff_A_iuKWqCDK1_0(.dout(w_dff_A_fGlpwA8o1_0),.din(w_dff_A_iuKWqCDK1_0),.clk(gclk));
	jdff dff_A_KLo7KpIM1_1(.dout(w_G56gat_1[1]),.din(w_dff_A_KLo7KpIM1_1),.clk(gclk));
	jdff dff_A_8wcGsKQx9_1(.dout(w_G56gat_0[1]),.din(w_dff_A_8wcGsKQx9_1),.clk(gclk));
	jdff dff_A_dLuEru8m7_1(.dout(w_dff_A_8wcGsKQx9_1),.din(w_dff_A_dLuEru8m7_1),.clk(gclk));
	jdff dff_A_LU6UkSEE9_1(.dout(w_dff_A_dLuEru8m7_1),.din(w_dff_A_LU6UkSEE9_1),.clk(gclk));
	jdff dff_A_YTewSvrr7_1(.dout(w_dff_A_LU6UkSEE9_1),.din(w_dff_A_YTewSvrr7_1),.clk(gclk));
	jdff dff_A_ebOJZH0D9_1(.dout(w_dff_A_YTewSvrr7_1),.din(w_dff_A_ebOJZH0D9_1),.clk(gclk));
	jdff dff_A_VabbyFyh1_1(.dout(w_dff_A_ebOJZH0D9_1),.din(w_dff_A_VabbyFyh1_1),.clk(gclk));
	jdff dff_A_tyvo7vN59_1(.dout(w_dff_A_VabbyFyh1_1),.din(w_dff_A_tyvo7vN59_1),.clk(gclk));
	jdff dff_A_tHuw6Rx03_1(.dout(w_dff_A_tyvo7vN59_1),.din(w_dff_A_tHuw6Rx03_1),.clk(gclk));
	jdff dff_A_d4TMXWAz4_1(.dout(w_dff_A_tHuw6Rx03_1),.din(w_dff_A_d4TMXWAz4_1),.clk(gclk));
	jdff dff_A_7oq7v2Oe7_1(.dout(w_dff_A_d4TMXWAz4_1),.din(w_dff_A_7oq7v2Oe7_1),.clk(gclk));
	jdff dff_A_Fdx6kx4w0_1(.dout(w_dff_A_7oq7v2Oe7_1),.din(w_dff_A_Fdx6kx4w0_1),.clk(gclk));
	jdff dff_A_k5GyKWBM9_1(.dout(w_dff_A_Fdx6kx4w0_1),.din(w_dff_A_k5GyKWBM9_1),.clk(gclk));
	jdff dff_A_5M1BU1WW1_1(.dout(w_dff_A_k5GyKWBM9_1),.din(w_dff_A_5M1BU1WW1_1),.clk(gclk));
	jdff dff_A_wO1R5bKD2_1(.dout(w_dff_A_5M1BU1WW1_1),.din(w_dff_A_wO1R5bKD2_1),.clk(gclk));
	jdff dff_A_macC6PVE0_1(.dout(w_dff_A_wO1R5bKD2_1),.din(w_dff_A_macC6PVE0_1),.clk(gclk));
	jdff dff_A_nxnwmZGd1_1(.dout(w_dff_A_macC6PVE0_1),.din(w_dff_A_nxnwmZGd1_1),.clk(gclk));
	jdff dff_A_gqGFj5658_1(.dout(w_dff_A_nxnwmZGd1_1),.din(w_dff_A_gqGFj5658_1),.clk(gclk));
	jdff dff_A_c2IuFEPq5_1(.dout(w_dff_A_gqGFj5658_1),.din(w_dff_A_c2IuFEPq5_1),.clk(gclk));
	jdff dff_A_sgoJJj325_1(.dout(w_dff_A_c2IuFEPq5_1),.din(w_dff_A_sgoJJj325_1),.clk(gclk));
	jdff dff_A_MNKC2Dk62_1(.dout(w_dff_A_sgoJJj325_1),.din(w_dff_A_MNKC2Dk62_1),.clk(gclk));
	jdff dff_A_z0lqQNYb6_1(.dout(w_dff_A_MNKC2Dk62_1),.din(w_dff_A_z0lqQNYb6_1),.clk(gclk));
	jdff dff_A_3HySTJXS6_1(.dout(w_dff_A_z0lqQNYb6_1),.din(w_dff_A_3HySTJXS6_1),.clk(gclk));
	jdff dff_A_BzjL9RWB2_2(.dout(w_G56gat_0[2]),.din(w_dff_A_BzjL9RWB2_2),.clk(gclk));
	jdff dff_A_sc7G6lZl4_2(.dout(w_dff_A_BzjL9RWB2_2),.din(w_dff_A_sc7G6lZl4_2),.clk(gclk));
	jdff dff_A_uXNkjymG2_2(.dout(w_dff_A_sc7G6lZl4_2),.din(w_dff_A_uXNkjymG2_2),.clk(gclk));
	jdff dff_A_vW0lIcPc0_2(.dout(w_dff_A_uXNkjymG2_2),.din(w_dff_A_vW0lIcPc0_2),.clk(gclk));
	jdff dff_A_AdlW5dGu1_2(.dout(w_dff_A_vW0lIcPc0_2),.din(w_dff_A_AdlW5dGu1_2),.clk(gclk));
	jdff dff_A_zmE76EGO9_2(.dout(w_dff_A_AdlW5dGu1_2),.din(w_dff_A_zmE76EGO9_2),.clk(gclk));
	jdff dff_A_67DigGNO6_2(.dout(w_dff_A_zmE76EGO9_2),.din(w_dff_A_67DigGNO6_2),.clk(gclk));
	jdff dff_A_38dReck29_0(.dout(w_G50gat_0[0]),.din(w_dff_A_38dReck29_0),.clk(gclk));
	jdff dff_A_IBe76F2N6_0(.dout(w_n78_0[0]),.din(w_dff_A_IBe76F2N6_0),.clk(gclk));
	jdff dff_A_LBJHi2yA5_0(.dout(w_dff_A_IBe76F2N6_0),.din(w_dff_A_LBJHi2yA5_0),.clk(gclk));
	jdff dff_A_cSrLcZQX1_0(.dout(w_dff_A_LBJHi2yA5_0),.din(w_dff_A_cSrLcZQX1_0),.clk(gclk));
	jdff dff_A_k2PzWjou7_0(.dout(w_dff_A_cSrLcZQX1_0),.din(w_dff_A_k2PzWjou7_0),.clk(gclk));
	jdff dff_A_wiqJSjdl0_0(.dout(w_dff_A_k2PzWjou7_0),.din(w_dff_A_wiqJSjdl0_0),.clk(gclk));
	jdff dff_A_LPwi6se02_0(.dout(w_dff_A_wiqJSjdl0_0),.din(w_dff_A_LPwi6se02_0),.clk(gclk));
	jdff dff_A_SlVvIL6N8_0(.dout(w_G30gat_0[0]),.din(w_dff_A_SlVvIL6N8_0),.clk(gclk));
	jdff dff_A_tr8YxxJk1_0(.dout(w_dff_A_SlVvIL6N8_0),.din(w_dff_A_tr8YxxJk1_0),.clk(gclk));
	jdff dff_A_7B3ZcoPL1_0(.dout(w_dff_A_tr8YxxJk1_0),.din(w_dff_A_7B3ZcoPL1_0),.clk(gclk));
	jdff dff_A_ZosyvRvQ5_0(.dout(w_dff_A_7B3ZcoPL1_0),.din(w_dff_A_ZosyvRvQ5_0),.clk(gclk));
	jdff dff_A_2nEkXE7m1_0(.dout(w_dff_A_ZosyvRvQ5_0),.din(w_dff_A_2nEkXE7m1_0),.clk(gclk));
	jdff dff_A_c3bypZTb4_0(.dout(w_dff_A_2nEkXE7m1_0),.din(w_dff_A_c3bypZTb4_0),.clk(gclk));
	jdff dff_A_WQrXtqZC6_0(.dout(w_dff_A_c3bypZTb4_0),.din(w_dff_A_WQrXtqZC6_0),.clk(gclk));
	jdff dff_A_eiXD1ttD4_2(.dout(w_G30gat_0[2]),.din(w_dff_A_eiXD1ttD4_2),.clk(gclk));
	jdff dff_A_asXunjx04_0(.dout(w_G24gat_0[0]),.din(w_dff_A_asXunjx04_0),.clk(gclk));
	jdff dff_A_w17O8rej4_0(.dout(w_dff_A_asXunjx04_0),.din(w_dff_A_w17O8rej4_0),.clk(gclk));
	jdff dff_A_HEQ2d7nX4_0(.dout(w_dff_A_w17O8rej4_0),.din(w_dff_A_HEQ2d7nX4_0),.clk(gclk));
	jdff dff_A_QtG5Up7k5_0(.dout(w_dff_A_HEQ2d7nX4_0),.din(w_dff_A_QtG5Up7k5_0),.clk(gclk));
	jdff dff_A_120NDMG06_0(.dout(w_dff_A_QtG5Up7k5_0),.din(w_dff_A_120NDMG06_0),.clk(gclk));
	jdff dff_A_S3XhaID98_0(.dout(w_dff_A_120NDMG06_0),.din(w_dff_A_S3XhaID98_0),.clk(gclk));
	jdff dff_A_PvHrowcr3_1(.dout(w_G24gat_0[1]),.din(w_dff_A_PvHrowcr3_1),.clk(gclk));
	jdff dff_A_MabweP9I7_0(.dout(w_n75_0[0]),.din(w_dff_A_MabweP9I7_0),.clk(gclk));
	jdff dff_A_AyaUzMts8_0(.dout(w_dff_A_MabweP9I7_0),.din(w_dff_A_AyaUzMts8_0),.clk(gclk));
	jdff dff_A_JoXecjJZ5_0(.dout(w_dff_A_AyaUzMts8_0),.din(w_dff_A_JoXecjJZ5_0),.clk(gclk));
	jdff dff_A_YyEC9TrN8_0(.dout(w_dff_A_JoXecjJZ5_0),.din(w_dff_A_YyEC9TrN8_0),.clk(gclk));
	jdff dff_A_lbWiKf2i3_0(.dout(w_dff_A_YyEC9TrN8_0),.din(w_dff_A_lbWiKf2i3_0),.clk(gclk));
	jdff dff_A_zabAMT5S6_0(.dout(w_dff_A_lbWiKf2i3_0),.din(w_dff_A_zabAMT5S6_0),.clk(gclk));
	jdff dff_A_rk0Ef1XQ4_0(.dout(w_G17gat_0[0]),.din(w_dff_A_rk0Ef1XQ4_0),.clk(gclk));
	jdff dff_A_0btwrpQX6_0(.dout(w_dff_A_rk0Ef1XQ4_0),.din(w_dff_A_0btwrpQX6_0),.clk(gclk));
	jdff dff_A_2cq9wl740_0(.dout(w_dff_A_0btwrpQX6_0),.din(w_dff_A_2cq9wl740_0),.clk(gclk));
	jdff dff_A_gOSXiN7N7_0(.dout(w_dff_A_2cq9wl740_0),.din(w_dff_A_gOSXiN7N7_0),.clk(gclk));
	jdff dff_A_eqpzt1Md9_0(.dout(w_dff_A_gOSXiN7N7_0),.din(w_dff_A_eqpzt1Md9_0),.clk(gclk));
	jdff dff_A_vcgU7BgU1_0(.dout(w_dff_A_eqpzt1Md9_0),.din(w_dff_A_vcgU7BgU1_0),.clk(gclk));
	jdff dff_A_DdvFNv9v8_0(.dout(w_dff_A_vcgU7BgU1_0),.din(w_dff_A_DdvFNv9v8_0),.clk(gclk));
	jdff dff_A_algeuzM07_2(.dout(w_G17gat_0[2]),.din(w_dff_A_algeuzM07_2),.clk(gclk));
	jdff dff_A_eM82LuXd5_0(.dout(w_G11gat_0[0]),.din(w_dff_A_eM82LuXd5_0),.clk(gclk));
	jdff dff_A_TEopAfeD2_0(.dout(w_dff_A_eM82LuXd5_0),.din(w_dff_A_TEopAfeD2_0),.clk(gclk));
	jdff dff_A_xP0569zs8_0(.dout(w_dff_A_TEopAfeD2_0),.din(w_dff_A_xP0569zs8_0),.clk(gclk));
	jdff dff_A_BeR21p7D0_0(.dout(w_dff_A_xP0569zs8_0),.din(w_dff_A_BeR21p7D0_0),.clk(gclk));
	jdff dff_A_R35Guu1I3_0(.dout(w_dff_A_BeR21p7D0_0),.din(w_dff_A_R35Guu1I3_0),.clk(gclk));
	jdff dff_A_F4ECU3Yl1_0(.dout(w_dff_A_R35Guu1I3_0),.din(w_dff_A_F4ECU3Yl1_0),.clk(gclk));
	jdff dff_A_eBSbcp988_1(.dout(w_G11gat_0[1]),.din(w_dff_A_eBSbcp988_1),.clk(gclk));
	jdff dff_A_Cnq4Y3gi7_0(.dout(w_n73_0[0]),.din(w_dff_A_Cnq4Y3gi7_0),.clk(gclk));
	jdff dff_A_XgR4sJ4e5_0(.dout(w_dff_A_Cnq4Y3gi7_0),.din(w_dff_A_XgR4sJ4e5_0),.clk(gclk));
	jdff dff_A_xdOwZ12M2_0(.dout(w_dff_A_XgR4sJ4e5_0),.din(w_dff_A_xdOwZ12M2_0),.clk(gclk));
	jdff dff_A_coqpr0cX2_0(.dout(w_dff_A_xdOwZ12M2_0),.din(w_dff_A_coqpr0cX2_0),.clk(gclk));
	jdff dff_A_PgZmOUSo7_0(.dout(w_dff_A_coqpr0cX2_0),.din(w_dff_A_PgZmOUSo7_0),.clk(gclk));
	jdff dff_A_EnKYUt7C8_0(.dout(w_dff_A_PgZmOUSo7_0),.din(w_dff_A_EnKYUt7C8_0),.clk(gclk));
	jdff dff_A_wM6M0nWR5_0(.dout(w_G69gat_0[0]),.din(w_dff_A_wM6M0nWR5_0),.clk(gclk));
	jdff dff_A_rGilqM3G7_0(.dout(w_dff_A_wM6M0nWR5_0),.din(w_dff_A_rGilqM3G7_0),.clk(gclk));
	jdff dff_A_xTJRYaT95_0(.dout(w_dff_A_rGilqM3G7_0),.din(w_dff_A_xTJRYaT95_0),.clk(gclk));
	jdff dff_A_05zSM0OU7_0(.dout(w_dff_A_xTJRYaT95_0),.din(w_dff_A_05zSM0OU7_0),.clk(gclk));
	jdff dff_A_741alT7e3_0(.dout(w_dff_A_05zSM0OU7_0),.din(w_dff_A_741alT7e3_0),.clk(gclk));
	jdff dff_A_2Y9OrBWF5_0(.dout(w_dff_A_741alT7e3_0),.din(w_dff_A_2Y9OrBWF5_0),.clk(gclk));
	jdff dff_A_o1hoiLYi4_0(.dout(w_dff_A_2Y9OrBWF5_0),.din(w_dff_A_o1hoiLYi4_0),.clk(gclk));
	jdff dff_A_RrmSmg7E5_2(.dout(w_G69gat_0[2]),.din(w_dff_A_RrmSmg7E5_2),.clk(gclk));
	jdff dff_A_d9v12Sb57_0(.dout(w_n46_0[0]),.din(w_dff_A_d9v12Sb57_0),.clk(gclk));
	jdff dff_A_pljv0OjR5_0(.dout(w_dff_A_d9v12Sb57_0),.din(w_dff_A_pljv0OjR5_0),.clk(gclk));
	jdff dff_A_AEXiYSKt0_0(.dout(w_dff_A_pljv0OjR5_0),.din(w_dff_A_AEXiYSKt0_0),.clk(gclk));
	jdff dff_A_kRJdjUmV6_0(.dout(w_dff_A_AEXiYSKt0_0),.din(w_dff_A_kRJdjUmV6_0),.clk(gclk));
	jdff dff_A_CBjgYnE14_1(.dout(w_n46_0[1]),.din(w_dff_A_CBjgYnE14_1),.clk(gclk));
	jdff dff_B_G0rNMgmM4_1(.din(G37gat),.dout(w_dff_B_G0rNMgmM4_1),.clk(gclk));
	jdff dff_A_oDpvd1uY3_0(.dout(w_n45_0[0]),.din(w_dff_A_oDpvd1uY3_0),.clk(gclk));
	jdff dff_A_DkMJvmm33_0(.dout(w_dff_A_oDpvd1uY3_0),.din(w_dff_A_DkMJvmm33_0),.clk(gclk));
	jdff dff_A_Eb2Yup1z2_0(.dout(w_dff_A_DkMJvmm33_0),.din(w_dff_A_Eb2Yup1z2_0),.clk(gclk));
	jdff dff_A_OhgP6H9w5_0(.dout(w_dff_A_Eb2Yup1z2_0),.din(w_dff_A_OhgP6H9w5_0),.clk(gclk));
	jdff dff_A_pM4Ofpgb7_0(.dout(w_dff_A_OhgP6H9w5_0),.din(w_dff_A_pM4Ofpgb7_0),.clk(gclk));
	jdff dff_A_05Ai5toY8_0(.dout(w_dff_A_pM4Ofpgb7_0),.din(w_dff_A_05Ai5toY8_0),.clk(gclk));
	jdff dff_A_vfRa9laY8_0(.dout(w_G43gat_0[0]),.din(w_dff_A_vfRa9laY8_0),.clk(gclk));
	jdff dff_A_8Cs8PhPB6_0(.dout(w_dff_A_vfRa9laY8_0),.din(w_dff_A_8Cs8PhPB6_0),.clk(gclk));
	jdff dff_A_hhT4Jx8v0_0(.dout(w_dff_A_8Cs8PhPB6_0),.din(w_dff_A_hhT4Jx8v0_0),.clk(gclk));
	jdff dff_A_c6qjtPui5_0(.dout(w_dff_A_hhT4Jx8v0_0),.din(w_dff_A_c6qjtPui5_0),.clk(gclk));
	jdff dff_A_22k1zkSY4_0(.dout(w_dff_A_c6qjtPui5_0),.din(w_dff_A_22k1zkSY4_0),.clk(gclk));
	jdff dff_A_eUT9tNhY0_0(.dout(w_dff_A_22k1zkSY4_0),.din(w_dff_A_eUT9tNhY0_0),.clk(gclk));
	jdff dff_A_oft2wnYa5_0(.dout(w_dff_A_eUT9tNhY0_0),.din(w_dff_A_oft2wnYa5_0),.clk(gclk));
	jdff dff_A_HoANK5OL6_1(.dout(w_n44_0[1]),.din(w_dff_A_HoANK5OL6_1),.clk(gclk));
	jdff dff_A_RxVzK2DL7_1(.dout(w_G108gat_0[1]),.din(w_dff_A_RxVzK2DL7_1),.clk(gclk));
	jdff dff_A_4r98Dtqy5_1(.dout(w_dff_A_RxVzK2DL7_1),.din(w_dff_A_4r98Dtqy5_1),.clk(gclk));
	jdff dff_A_MnNDID1c5_1(.dout(w_dff_A_4r98Dtqy5_1),.din(w_dff_A_MnNDID1c5_1),.clk(gclk));
	jdff dff_A_LkRv3Zqz5_1(.dout(w_dff_A_MnNDID1c5_1),.din(w_dff_A_LkRv3Zqz5_1),.clk(gclk));
	jdff dff_A_MBsFD3iu8_1(.dout(w_dff_A_LkRv3Zqz5_1),.din(w_dff_A_MBsFD3iu8_1),.clk(gclk));
	jdff dff_A_nfpFi98I8_1(.dout(w_dff_A_MBsFD3iu8_1),.din(w_dff_A_nfpFi98I8_1),.clk(gclk));
	jdff dff_A_eimXMdMg7_1(.dout(w_dff_A_nfpFi98I8_1),.din(w_dff_A_eimXMdMg7_1),.clk(gclk));
	jdff dff_A_OmXIee1c6_2(.dout(w_G108gat_0[2]),.din(w_dff_A_OmXIee1c6_2),.clk(gclk));
	jdff dff_A_zVidtoy64_0(.dout(w_n43_0[0]),.din(w_dff_A_zVidtoy64_0),.clk(gclk));
	jdff dff_A_nU0cGZB42_0(.dout(w_dff_A_zVidtoy64_0),.din(w_dff_A_nU0cGZB42_0),.clk(gclk));
	jdff dff_A_UDmQ15sN3_0(.dout(w_dff_A_nU0cGZB42_0),.din(w_dff_A_UDmQ15sN3_0),.clk(gclk));
	jdff dff_A_Klm7WHf28_0(.dout(w_dff_A_UDmQ15sN3_0),.din(w_dff_A_Klm7WHf28_0),.clk(gclk));
	jdff dff_A_hsvJpFM39_0(.dout(w_dff_A_Klm7WHf28_0),.din(w_dff_A_hsvJpFM39_0),.clk(gclk));
	jdff dff_A_UUJHy9aY1_0(.dout(w_G102gat_0[0]),.din(w_dff_A_UUJHy9aY1_0),.clk(gclk));
	jdff dff_A_MD3643T96_0(.dout(w_dff_A_UUJHy9aY1_0),.din(w_dff_A_MD3643T96_0),.clk(gclk));
	jdff dff_A_lGW3MMVj8_0(.dout(w_dff_A_MD3643T96_0),.din(w_dff_A_lGW3MMVj8_0),.clk(gclk));
	jdff dff_A_erP4FJQC0_0(.dout(w_dff_A_lGW3MMVj8_0),.din(w_dff_A_erP4FJQC0_0),.clk(gclk));
	jdff dff_A_5USV3o975_0(.dout(w_dff_A_erP4FJQC0_0),.din(w_dff_A_5USV3o975_0),.clk(gclk));
	jdff dff_A_8Lhq2fEL2_0(.dout(w_dff_A_5USV3o975_0),.din(w_dff_A_8Lhq2fEL2_0),.clk(gclk));
	jdff dff_A_qfLvVxkS1_0(.dout(w_n49_0[0]),.din(w_dff_A_qfLvVxkS1_0),.clk(gclk));
	jdff dff_A_s0FqWuix1_0(.dout(w_dff_A_qfLvVxkS1_0),.din(w_dff_A_s0FqWuix1_0),.clk(gclk));
	jdff dff_A_a6GzlPaf0_0(.dout(w_dff_A_s0FqWuix1_0),.din(w_dff_A_a6GzlPaf0_0),.clk(gclk));
	jdff dff_A_JweVlmwy5_0(.dout(w_dff_A_a6GzlPaf0_0),.din(w_dff_A_JweVlmwy5_0),.clk(gclk));
	jdff dff_A_bZLERgLv8_0(.dout(w_dff_A_JweVlmwy5_0),.din(w_dff_A_bZLERgLv8_0),.clk(gclk));
	jdff dff_A_FNl4fuHc6_0(.dout(w_G63gat_0[0]),.din(w_dff_A_FNl4fuHc6_0),.clk(gclk));
	jdff dff_A_NkcHCvcA7_0(.dout(w_dff_A_FNl4fuHc6_0),.din(w_dff_A_NkcHCvcA7_0),.clk(gclk));
	jdff dff_A_G3IE0QgD5_0(.dout(w_dff_A_NkcHCvcA7_0),.din(w_dff_A_G3IE0QgD5_0),.clk(gclk));
	jdff dff_A_5YwW0yUb5_0(.dout(w_dff_A_G3IE0QgD5_0),.din(w_dff_A_5YwW0yUb5_0),.clk(gclk));
	jdff dff_A_3sOePMWg6_0(.dout(w_dff_A_5YwW0yUb5_0),.din(w_dff_A_3sOePMWg6_0),.clk(gclk));
	jdff dff_A_F8UourEb8_0(.dout(w_dff_A_3sOePMWg6_0),.din(w_dff_A_F8UourEb8_0),.clk(gclk));
	jdff dff_A_hnHpacdE9_1(.dout(w_G63gat_0[1]),.din(w_dff_A_hnHpacdE9_1),.clk(gclk));
	jdff dff_A_vQF300D38_1(.dout(w_dff_A_ejRr1Wao7_0),.din(w_dff_A_vQF300D38_1),.clk(gclk));
	jdff dff_A_ejRr1Wao7_0(.dout(w_dff_A_aNUq5zKg5_0),.din(w_dff_A_ejRr1Wao7_0),.clk(gclk));
	jdff dff_A_aNUq5zKg5_0(.dout(w_dff_A_JqVg5MQE1_0),.din(w_dff_A_aNUq5zKg5_0),.clk(gclk));
	jdff dff_A_JqVg5MQE1_0(.dout(w_dff_A_XnQmRbMn9_0),.din(w_dff_A_JqVg5MQE1_0),.clk(gclk));
	jdff dff_A_XnQmRbMn9_0(.dout(w_dff_A_NgOxlcCU6_0),.din(w_dff_A_XnQmRbMn9_0),.clk(gclk));
	jdff dff_A_NgOxlcCU6_0(.dout(w_dff_A_GDlDXedd5_0),.din(w_dff_A_NgOxlcCU6_0),.clk(gclk));
	jdff dff_A_GDlDXedd5_0(.dout(w_dff_A_VUpbDg4h6_0),.din(w_dff_A_GDlDXedd5_0),.clk(gclk));
	jdff dff_A_VUpbDg4h6_0(.dout(w_dff_A_jI60A05b1_0),.din(w_dff_A_VUpbDg4h6_0),.clk(gclk));
	jdff dff_A_jI60A05b1_0(.dout(w_dff_A_KkAXZY2U1_0),.din(w_dff_A_jI60A05b1_0),.clk(gclk));
	jdff dff_A_KkAXZY2U1_0(.dout(w_dff_A_IPn330I22_0),.din(w_dff_A_KkAXZY2U1_0),.clk(gclk));
	jdff dff_A_IPn330I22_0(.dout(w_dff_A_34aUbV7e2_0),.din(w_dff_A_IPn330I22_0),.clk(gclk));
	jdff dff_A_34aUbV7e2_0(.dout(w_dff_A_5F54Zuqg9_0),.din(w_dff_A_34aUbV7e2_0),.clk(gclk));
	jdff dff_A_5F54Zuqg9_0(.dout(w_dff_A_LnLCDlFK8_0),.din(w_dff_A_5F54Zuqg9_0),.clk(gclk));
	jdff dff_A_LnLCDlFK8_0(.dout(w_dff_A_cVlkYZFJ1_0),.din(w_dff_A_LnLCDlFK8_0),.clk(gclk));
	jdff dff_A_cVlkYZFJ1_0(.dout(w_dff_A_9xuIsWKI1_0),.din(w_dff_A_cVlkYZFJ1_0),.clk(gclk));
	jdff dff_A_9xuIsWKI1_0(.dout(w_dff_A_oMk0Sfed2_0),.din(w_dff_A_9xuIsWKI1_0),.clk(gclk));
	jdff dff_A_oMk0Sfed2_0(.dout(w_dff_A_i8ye4iiK7_0),.din(w_dff_A_oMk0Sfed2_0),.clk(gclk));
	jdff dff_A_i8ye4iiK7_0(.dout(w_dff_A_eNw8VwPP9_0),.din(w_dff_A_i8ye4iiK7_0),.clk(gclk));
	jdff dff_A_eNw8VwPP9_0(.dout(w_dff_A_vttDMYKt0_0),.din(w_dff_A_eNw8VwPP9_0),.clk(gclk));
	jdff dff_A_vttDMYKt0_0(.dout(w_dff_A_baacOaEL2_0),.din(w_dff_A_vttDMYKt0_0),.clk(gclk));
	jdff dff_A_baacOaEL2_0(.dout(G223gat),.din(w_dff_A_baacOaEL2_0),.clk(gclk));
	jdff dff_A_qQJGeCWt3_1(.dout(w_dff_A_KlqEYryB7_0),.din(w_dff_A_qQJGeCWt3_1),.clk(gclk));
	jdff dff_A_KlqEYryB7_0(.dout(w_dff_A_xdCspEKk1_0),.din(w_dff_A_KlqEYryB7_0),.clk(gclk));
	jdff dff_A_xdCspEKk1_0(.dout(w_dff_A_gLfy1ggQ9_0),.din(w_dff_A_xdCspEKk1_0),.clk(gclk));
	jdff dff_A_gLfy1ggQ9_0(.dout(w_dff_A_Ofb9KTck9_0),.din(w_dff_A_gLfy1ggQ9_0),.clk(gclk));
	jdff dff_A_Ofb9KTck9_0(.dout(w_dff_A_fzonw2D54_0),.din(w_dff_A_Ofb9KTck9_0),.clk(gclk));
	jdff dff_A_fzonw2D54_0(.dout(w_dff_A_GRjqZ6qO6_0),.din(w_dff_A_fzonw2D54_0),.clk(gclk));
	jdff dff_A_GRjqZ6qO6_0(.dout(w_dff_A_y8LDHsvB4_0),.din(w_dff_A_GRjqZ6qO6_0),.clk(gclk));
	jdff dff_A_y8LDHsvB4_0(.dout(w_dff_A_rC33axc43_0),.din(w_dff_A_y8LDHsvB4_0),.clk(gclk));
	jdff dff_A_rC33axc43_0(.dout(w_dff_A_gBKVROkF6_0),.din(w_dff_A_rC33axc43_0),.clk(gclk));
	jdff dff_A_gBKVROkF6_0(.dout(w_dff_A_BmxIRDOu0_0),.din(w_dff_A_gBKVROkF6_0),.clk(gclk));
	jdff dff_A_BmxIRDOu0_0(.dout(w_dff_A_XVm4blHM1_0),.din(w_dff_A_BmxIRDOu0_0),.clk(gclk));
	jdff dff_A_XVm4blHM1_0(.dout(w_dff_A_n5Eu2lKB6_0),.din(w_dff_A_XVm4blHM1_0),.clk(gclk));
	jdff dff_A_n5Eu2lKB6_0(.dout(w_dff_A_FJBVPdWa6_0),.din(w_dff_A_n5Eu2lKB6_0),.clk(gclk));
	jdff dff_A_FJBVPdWa6_0(.dout(G329gat),.din(w_dff_A_FJBVPdWa6_0),.clk(gclk));
	jdff dff_A_VpmklDhU3_2(.dout(w_dff_A_FigXqfKP0_0),.din(w_dff_A_VpmklDhU3_2),.clk(gclk));
	jdff dff_A_FigXqfKP0_0(.dout(w_dff_A_lATlPhVO1_0),.din(w_dff_A_FigXqfKP0_0),.clk(gclk));
	jdff dff_A_lATlPhVO1_0(.dout(w_dff_A_7hPv0BTi1_0),.din(w_dff_A_lATlPhVO1_0),.clk(gclk));
	jdff dff_A_7hPv0BTi1_0(.dout(w_dff_A_a949ANRM9_0),.din(w_dff_A_7hPv0BTi1_0),.clk(gclk));
	jdff dff_A_a949ANRM9_0(.dout(w_dff_A_ndvlgC9D9_0),.din(w_dff_A_a949ANRM9_0),.clk(gclk));
	jdff dff_A_ndvlgC9D9_0(.dout(w_dff_A_WuH62Us75_0),.din(w_dff_A_ndvlgC9D9_0),.clk(gclk));
	jdff dff_A_WuH62Us75_0(.dout(G370gat),.din(w_dff_A_WuH62Us75_0),.clk(gclk));
	jdff dff_A_EIdOR7m34_1(.dout(w_dff_A_7aVGoP6A3_0),.din(w_dff_A_EIdOR7m34_1),.clk(gclk));
	jdff dff_A_7aVGoP6A3_0(.dout(G430gat),.din(w_dff_A_7aVGoP6A3_0),.clk(gclk));
endmodule

