/*

c1908:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jdff: 153
	jand: 128
	jor: 102

Summary:
	jxor: 74
	jspl: 106
	jspl3: 95
	jnot: 41
	jdff: 153
	jand: 128
	jor: 102

The maximum logic level gap of any gate:
	c1908: 17
*/

module rf_c1908(gclk, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57);
	input gclk;
	input G101;
	input G104;
	input G107;
	input G110;
	input G113;
	input G116;
	input G119;
	input G122;
	input G125;
	input G128;
	input G131;
	input G134;
	input G137;
	input G140;
	input G143;
	input G146;
	input G210;
	input G214;
	input G217;
	input G221;
	input G224;
	input G227;
	input G234;
	input G237;
	input G469;
	input G472;
	input G475;
	input G478;
	input G898;
	input G900;
	input G902;
	input G952;
	input G953;
	output G3;
	output G6;
	output G9;
	output G12;
	output G30;
	output G45;
	output G48;
	output G15;
	output G18;
	output G21;
	output G24;
	output G27;
	output G33;
	output G36;
	output G39;
	output G42;
	output G75;
	output G51;
	output G54;
	output G60;
	output G63;
	output G66;
	output G69;
	output G72;
	output G57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n188;
	wire n189;
	wire n190;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n202;
	wire n204;
	wire n205;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n222;
	wire n224;
	wire n225;
	wire n226;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire[2:0] w_G101_0;
	wire[2:0] w_G104_0;
	wire[2:0] w_G107_0;
	wire[2:0] w_G110_0;
	wire[1:0] w_G110_1;
	wire[1:0] w_G113_0;
	wire[2:0] w_G116_0;
	wire[2:0] w_G119_0;
	wire[2:0] w_G122_0;
	wire[1:0] w_G122_1;
	wire[2:0] w_G125_0;
	wire[2:0] w_G128_0;
	wire[1:0] w_G128_1;
	wire[1:0] w_G131_0;
	wire[2:0] w_G134_0;
	wire[2:0] w_G137_0;
	wire[2:0] w_G140_0;
	wire[2:0] w_G143_0;
	wire[1:0] w_G143_1;
	wire[2:0] w_G146_0;
	wire[2:0] w_G210_0;
	wire[1:0] w_G214_0;
	wire[2:0] w_G217_0;
	wire[1:0] w_G221_0;
	wire[1:0] w_G224_0;
	wire[1:0] w_G227_0;
	wire[2:0] w_G234_0;
	wire[2:0] w_G237_0;
	wire[2:0] w_G469_0;
	wire[1:0] w_G472_0;
	wire[2:0] w_G475_0;
	wire[2:0] w_G478_0;
	wire[2:0] w_G902_0;
	wire[2:0] w_G902_1;
	wire[2:0] w_G902_2;
	wire[2:0] w_G902_3;
	wire[2:0] w_G952_0;
	wire[2:0] w_G953_0;
	wire[2:0] w_G953_1;
	wire[1:0] w_n59_0;
	wire[2:0] w_n60_0;
	wire[2:0] w_n61_0;
	wire[2:0] w_n61_1;
	wire[2:0] w_n61_2;
	wire[2:0] w_n61_3;
	wire[1:0] w_n62_0;
	wire[1:0] w_n67_0;
	wire[1:0] w_n68_0;
	wire[2:0] w_n70_0;
	wire[2:0] w_n70_1;
	wire[2:0] w_n70_2;
	wire[1:0] w_n70_3;
	wire[1:0] w_n71_0;
	wire[1:0] w_n73_0;
	wire[2:0] w_n74_0;
	wire[1:0] w_n74_1;
	wire[1:0] w_n77_0;
	wire[1:0] w_n79_0;
	wire[2:0] w_n81_0;
	wire[1:0] w_n82_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[2:0] w_n90_0;
	wire[2:0] w_n92_0;
	wire[2:0] w_n92_1;
	wire[2:0] w_n93_0;
	wire[1:0] w_n94_0;
	wire[2:0] w_n95_0;
	wire[2:0] w_n96_0;
	wire[1:0] w_n97_0;
	wire[1:0] w_n101_0;
	wire[1:0] w_n103_0;
	wire[2:0] w_n107_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n109_0;
	wire[2:0] w_n110_0;
	wire[2:0] w_n112_0;
	wire[1:0] w_n112_1;
	wire[2:0] w_n117_0;
	wire[1:0] w_n118_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[2:0] w_n121_0;
	wire[1:0] w_n121_1;
	wire[1:0] w_n122_0;
	wire[2:0] w_n130_0;
	wire[1:0] w_n131_0;
	wire[2:0] w_n132_0;
	wire[2:0] w_n141_0;
	wire[1:0] w_n142_0;
	wire[2:0] w_n143_0;
	wire[1:0] w_n143_1;
	wire[2:0] w_n144_0;
	wire[2:0] w_n144_1;
	wire[1:0] w_n145_0;
	wire[1:0] w_n146_0;
	wire[1:0] w_n147_0;
	wire[2:0] w_n151_0;
	wire[1:0] w_n152_0;
	wire[2:0] w_n153_0;
	wire[2:0] w_n154_0;
	wire[1:0] w_n154_1;
	wire[2:0] w_n155_0;
	wire[1:0] w_n156_0;
	wire[2:0] w_n158_0;
	wire[1:0] w_n158_1;
	wire[2:0] w_n159_0;
	wire[1:0] w_n159_1;
	wire[1:0] w_n160_0;
	wire[2:0] w_n161_0;
	wire[1:0] w_n162_0;
	wire[2:0] w_n163_0;
	wire[1:0] w_n164_0;
	wire[2:0] w_n166_0;
	wire[1:0] w_n166_1;
	wire[1:0] w_n167_0;
	wire[2:0] w_n168_0;
	wire[1:0] w_n169_0;
	wire[1:0] w_n172_0;
	wire[2:0] w_n174_0;
	wire[1:0] w_n174_1;
	wire[1:0] w_n175_0;
	wire[1:0] w_n177_0;
	wire[2:0] w_n179_0;
	wire[1:0] w_n180_0;
	wire[2:0] w_n181_0;
	wire[2:0] w_n183_0;
	wire[2:0] w_n184_0;
	wire[1:0] w_n184_1;
	wire[2:0] w_n185_0;
	wire[1:0] w_n186_0;
	wire[2:0] w_n188_0;
	wire[1:0] w_n189_0;
	wire[1:0] w_n190_0;
	wire[2:0] w_n192_0;
	wire[1:0] w_n193_0;
	wire[2:0] w_n196_0;
	wire[2:0] w_n197_0;
	wire[1:0] w_n197_1;
	wire[2:0] w_n198_0;
	wire[1:0] w_n198_1;
	wire[1:0] w_n199_0;
	wire[1:0] w_n200_0;
	wire[1:0] w_n202_0;
	wire[1:0] w_n205_0;
	wire[1:0] w_n207_0;
	wire[1:0] w_n210_0;
	wire[1:0] w_n212_0;
	wire[1:0] w_n213_0;
	wire[2:0] w_n216_0;
	wire[2:0] w_n217_0;
	wire[2:0] w_n218_0;
	wire[1:0] w_n218_1;
	wire[1:0] w_n219_0;
	wire[1:0] w_n220_0;
	wire[1:0] w_n222_0;
	wire[1:0] w_n226_0;
	wire[1:0] w_n228_0;
	wire[2:0] w_n244_0;
	wire[2:0] w_n244_1;
	wire[2:0] w_n244_2;
	wire[1:0] w_n252_0;
	wire[2:0] w_n253_0;
	wire[2:0] w_n254_0;
	wire[1:0] w_n254_1;
	wire[2:0] w_n273_0;
	wire[1:0] w_n274_0;
	wire[1:0] w_n275_0;
	wire[2:0] w_n276_0;
	wire[1:0] w_n276_1;
	wire[1:0] w_n277_0;
	wire[1:0] w_n278_0;
	wire[1:0] w_n280_0;
	wire[2:0] w_n281_0;
	wire[1:0] w_n282_0;
	wire[1:0] w_n286_0;
	wire[2:0] w_n288_0;
	wire[1:0] w_n289_0;
	wire[2:0] w_n290_0;
	wire[1:0] w_n291_0;
	wire[1:0] w_n295_0;
	wire[1:0] w_n308_0;
	wire[1:0] w_n309_0;
	wire[2:0] w_n311_0;
	wire[2:0] w_n314_0;
	wire[1:0] w_n315_0;
	wire[1:0] w_n318_0;
	wire[1:0] w_n325_0;
	wire[1:0] w_n334_0;
	wire[2:0] w_n335_0;
	wire[2:0] w_n335_1;
	wire[1:0] w_n335_2;
	wire[1:0] w_n336_0;
	wire[2:0] w_n340_0;
	wire[2:0] w_n340_1;
	wire[1:0] w_n340_2;
	wire[1:0] w_n346_0;
	wire[1:0] w_n355_0;
	wire[1:0] w_n364_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n395_0;
	wire w_dff_B_ZVKO1Mo51_0;
	wire w_dff_B_Bnhasfkr6_0;
	wire w_dff_B_P396Rp8F4_0;
	wire w_dff_B_GO4wAQ8u2_0;
	wire w_dff_B_hos9PQp09_0;
	wire w_dff_B_2orChbYK1_1;
	wire w_dff_B_kjsma4km9_1;
	wire w_dff_B_CqM0mfmv2_1;
	wire w_dff_B_kssSIq840_1;
	wire w_dff_B_29RFV7IF1_1;
	wire w_dff_B_dzWAwNCf7_1;
	wire w_dff_B_BZfl0Bnq5_1;
	wire w_dff_B_6RKKJuU99_1;
	wire w_dff_B_b0kIoAb76_1;
	wire w_dff_B_Le1XJwK91_1;
	wire w_dff_B_wfNoYcMm6_1;
	wire w_dff_B_fI246dkN2_1;
	wire w_dff_B_WWxgCCjf9_1;
	wire w_dff_B_42RkquX53_1;
	wire w_dff_B_VMt0Omiv0_1;
	wire w_dff_B_mzcgcshM3_1;
	wire w_dff_B_QiucouSo8_1;
	wire w_dff_B_WpLdC2yf9_1;
	wire w_dff_B_sOwajJPg5_1;
	wire w_dff_B_LumDwg734_1;
	wire w_dff_B_Kw5aBqFC1_0;
	wire w_dff_B_DheBu80T7_0;
	wire w_dff_B_8F8oQlE15_0;
	wire w_dff_B_4zXuBon64_0;
	wire w_dff_B_5Bc3Cq8z0_0;
	wire w_dff_B_xU9fo7k41_0;
	wire w_dff_B_hW7WgSM70_0;
	wire w_dff_B_EtTbpHWJ2_0;
	wire w_dff_B_3EXQ8fe84_0;
	wire w_dff_B_zJp7DNCj6_0;
	wire w_dff_B_dlWi642E9_0;
	wire w_dff_B_9rmQ04lU6_1;
	wire w_dff_A_fuse14T61_2;
	wire w_dff_A_9MUfrTW15_0;
	wire w_dff_A_dKF5pgqF8_0;
	wire w_dff_A_GbxA3kj26_0;
	wire w_dff_A_BHlsa0a93_0;
	wire w_dff_A_U0ssrYvD0_0;
	wire w_dff_A_kzR5NI6S3_0;
	wire w_dff_A_2gaEHoHJ9_2;
	wire w_dff_A_hVjHpR7I4_0;
	wire w_dff_A_UvkMzsCG6_0;
	wire w_dff_A_DZ5w9hss0_0;
	wire w_dff_A_YbYzecui7_0;
	wire w_dff_A_aC57sAI99_0;
	wire w_dff_A_dYt9jr318_0;
	wire w_dff_A_P8R2qX6l0_2;
	wire w_dff_A_sBFpdlpI2_0;
	wire w_dff_A_wZeA5PC48_0;
	wire w_dff_A_LUesZXVF2_0;
	wire w_dff_A_EvlSyBMq0_0;
	wire w_dff_A_QM9OZKLr8_0;
	wire w_dff_A_F7gG8OG23_0;
	wire w_dff_A_Iv1cyd7k5_2;
	wire w_dff_A_VlePD7MI0_0;
	wire w_dff_A_HYZxUNkd7_0;
	wire w_dff_A_iLKjr7Zx3_0;
	wire w_dff_A_y4IhiKIr6_0;
	wire w_dff_A_blTbcDJf5_0;
	wire w_dff_A_0lztIxwK2_0;
	wire w_dff_A_8PLLfsFp3_2;
	wire w_dff_A_KbdHPIkd9_0;
	wire w_dff_A_YAy6vcNW3_0;
	wire w_dff_A_MfXzEgtD1_0;
	wire w_dff_A_7enoBNa54_0;
	wire w_dff_A_9mzdA1ar1_0;
	wire w_dff_A_Yhxa399s3_0;
	wire w_dff_A_uKogXNzU7_2;
	wire w_dff_A_GmLMgmTL9_0;
	wire w_dff_A_LgLqwJ3d3_0;
	wire w_dff_A_19AiRCiG9_0;
	wire w_dff_A_x3Y4IHRn3_0;
	wire w_dff_A_nN8uEuiz3_0;
	wire w_dff_A_iijZsxpL1_0;
	wire w_dff_A_b9MQohhs2_2;
	wire w_dff_A_hzsudhFQ2_0;
	wire w_dff_A_44GvxLGf9_0;
	wire w_dff_A_lK6scgeg4_0;
	wire w_dff_A_7U93AYXO2_0;
	wire w_dff_A_1SbbXg5O1_0;
	wire w_dff_A_TTlaiYnO7_0;
	wire w_dff_A_30rl8IDl4_2;
	wire w_dff_A_dN4c5WwJ6_0;
	wire w_dff_A_2LSmskpI0_0;
	wire w_dff_A_TtEBxQGL1_0;
	wire w_dff_A_Z6NaGQ060_0;
	wire w_dff_A_NxsNfYrg8_0;
	wire w_dff_A_AspwU5ia6_0;
	wire w_dff_A_cPpb56RY3_2;
	wire w_dff_A_K82LTB7q9_0;
	wire w_dff_A_rCdHRB3a0_0;
	wire w_dff_A_iem2k9aV8_0;
	wire w_dff_A_nNwrKDRC4_0;
	wire w_dff_A_cFG1oKhb9_0;
	wire w_dff_A_MTLeesBI4_0;
	wire w_dff_A_vWFS0OZ25_2;
	wire w_dff_A_LodlJLby4_0;
	wire w_dff_A_2EtwuHP34_0;
	wire w_dff_A_EVhoD0Uo5_0;
	wire w_dff_A_JebwlGQM1_0;
	wire w_dff_A_lhgDSYtn2_0;
	wire w_dff_A_mhT7ScXv4_0;
	wire w_dff_A_fXWr2Uu04_2;
	wire w_dff_A_Cf4oJ98q5_0;
	wire w_dff_A_6q7OG8m15_0;
	wire w_dff_A_xH1dtE183_0;
	wire w_dff_A_C0HrwjsY5_0;
	wire w_dff_A_KZMoV3PV7_0;
	wire w_dff_A_H4dd3DQS0_0;
	wire w_dff_A_E9NAXxXK0_2;
	wire w_dff_A_03NK2lHB4_0;
	wire w_dff_A_k7YLEW7A6_0;
	wire w_dff_A_Zy92Q7jn2_0;
	wire w_dff_A_Q7HRDvYK1_0;
	wire w_dff_A_qel2dIz33_0;
	wire w_dff_A_ITyeNT9e2_0;
	wire w_dff_A_jF9YHq5j2_2;
	wire w_dff_A_iwZpseBI0_0;
	wire w_dff_A_RNmSBhdL7_0;
	wire w_dff_A_J57e2zIl8_0;
	wire w_dff_A_dPAcUBw47_0;
	wire w_dff_A_mE8iwXT05_0;
	wire w_dff_A_Bhg3h0bn3_0;
	wire w_dff_A_CObwD37Y6_2;
	wire w_dff_A_NkBrZtAD0_0;
	wire w_dff_A_ccYvgVl96_0;
	wire w_dff_A_ZmxJS0DB0_0;
	wire w_dff_A_uGB2f2br7_0;
	wire w_dff_A_gQJYD8Bv5_0;
	wire w_dff_A_q3v43UeU5_0;
	wire w_dff_A_9pyUhmRS8_2;
	wire w_dff_A_bEYpzb9h4_0;
	wire w_dff_A_ZP19CT7t9_0;
	wire w_dff_A_ihkGyJKt2_0;
	wire w_dff_A_yBM0Ovkd0_0;
	wire w_dff_A_kwbLCVc64_0;
	wire w_dff_A_m0SgaP3O1_0;
	wire w_dff_A_bMjqVEuP0_2;
	wire w_dff_A_eBQQkB3P1_0;
	wire w_dff_A_E0SZC2Xx1_0;
	wire w_dff_A_LEo8QUvu2_0;
	wire w_dff_A_pKqBkQWa2_0;
	wire w_dff_A_XygrURur2_0;
	wire w_dff_A_9BAqzG8j3_0;
	wire w_dff_A_T9z38KbT5_2;
	wire w_dff_A_wZn0xXb02_2;
	wire w_dff_A_EFbnONC66_2;
	wire w_dff_A_q1bJJ9db2_0;
	jnot g000(.din(w_G146_0[2]),.dout(n58),.clk(gclk));
	jxor g001(.dina(w_G140_0[2]),.dinb(w_G125_0[2]),.dout(n59),.clk(gclk));
	jxor g002(.dina(w_n59_0[1]),.dinb(n58),.dout(n60),.clk(gclk));
	jnot g003(.din(w_G953_1[2]),.dout(n61),.clk(gclk));
	jand g004(.dina(w_n61_3[2]),.dinb(w_G234_0[2]),.dout(n62),.clk(gclk));
	jand g005(.dina(w_n62_0[1]),.dinb(w_G221_0[1]),.dout(n63),.clk(gclk));
	jxor g006(.dina(n63),.dinb(w_G137_0[2]),.dout(n64),.clk(gclk));
	jxor g007(.dina(w_G128_1[1]),.dinb(w_G119_0[2]),.dout(n65),.clk(gclk));
	jxor g008(.dina(n65),.dinb(n64),.dout(n66),.clk(gclk));
	jxor g009(.dina(n66),.dinb(w_G110_1[1]),.dout(n67),.clk(gclk));
	jxor g010(.dina(w_n67_0[1]),.dinb(w_n60_0[2]),.dout(n68),.clk(gclk));
	jor g011(.dina(w_n68_0[1]),.dinb(w_G902_3[2]),.dout(n69),.clk(gclk));
	jnot g012(.din(w_G902_3[1]),.dout(n70),.clk(gclk));
	jand g013(.dina(w_n70_3[1]),.dinb(w_G234_0[1]),.dout(n71),.clk(gclk));
	jnot g014(.din(w_n71_0[1]),.dout(n72),.clk(gclk));
	jand g015(.dina(n72),.dinb(w_G217_0[2]),.dout(n73),.clk(gclk));
	jxor g016(.dina(w_n73_0[1]),.dinb(n69),.dout(n74),.clk(gclk));
	jnot g017(.din(w_G134_0[2]),.dout(n75),.clk(gclk));
	jxor g018(.dina(w_G137_0[1]),.dinb(n75),.dout(n76),.clk(gclk));
	jnot g019(.din(w_G131_0[1]),.dout(n77),.clk(gclk));
	jxor g020(.dina(w_G146_0[1]),.dinb(w_G143_1[1]),.dout(n78),.clk(gclk));
	jxor g021(.dina(n78),.dinb(w_G128_1[0]),.dout(n79),.clk(gclk));
	jxor g022(.dina(w_n79_0[1]),.dinb(w_n77_0[1]),.dout(n80),.clk(gclk));
	jxor g023(.dina(n80),.dinb(n76),.dout(n81),.clk(gclk));
	jnot g024(.din(w_G113_0[1]),.dout(n82),.clk(gclk));
	jxor g025(.dina(w_G119_0[1]),.dinb(w_G116_0[2]),.dout(n83),.clk(gclk));
	jxor g026(.dina(n83),.dinb(w_n82_0[1]),.dout(n84),.clk(gclk));
	jnot g027(.din(w_G210_0[2]),.dout(n85),.clk(gclk));
	jor g028(.dina(w_G953_1[1]),.dinb(w_G237_0[2]),.dout(n86),.clk(gclk));
	jor g029(.dina(w_n86_0[1]),.dinb(n85),.dout(n87),.clk(gclk));
	jxor g030(.dina(n87),.dinb(w_G101_0[2]),.dout(n88),.clk(gclk));
	jxor g031(.dina(n88),.dinb(w_n84_0[1]),.dout(n89),.clk(gclk));
	jxor g032(.dina(n89),.dinb(w_n81_0[2]),.dout(n90),.clk(gclk));
	jand g033(.dina(w_n90_0[2]),.dinb(w_n70_3[0]),.dout(n91),.clk(gclk));
	jxor g034(.dina(n91),.dinb(w_G472_0[1]),.dout(n92),.clk(gclk));
	jand g035(.dina(w_n92_1[2]),.dinb(w_n74_1[1]),.dout(n93),.clk(gclk));
	jor g036(.dina(w_G902_3[0]),.dinb(w_G237_0[1]),.dout(n94),.clk(gclk));
	jand g037(.dina(w_n94_0[1]),.dinb(w_G214_0[1]),.dout(n95),.clk(gclk));
	jnot g038(.din(w_n95_0[2]),.dout(n96),.clk(gclk));
	jand g039(.dina(w_n94_0[0]),.dinb(w_G210_0[1]),.dout(n97),.clk(gclk));
	jnot g040(.din(w_G110_1[0]),.dout(n98),.clk(gclk));
	jxor g041(.dina(w_G122_1[1]),.dinb(n98),.dout(n99),.clk(gclk));
	jxor g042(.dina(w_G107_0[2]),.dinb(w_G104_0[2]),.dout(n100),.clk(gclk));
	jxor g043(.dina(n100),.dinb(w_G101_0[1]),.dout(n101),.clk(gclk));
	jxor g044(.dina(w_n101_0[1]),.dinb(w_n84_0[0]),.dout(n102),.clk(gclk));
	jxor g045(.dina(n102),.dinb(n99),.dout(n103),.clk(gclk));
	jand g046(.dina(w_n61_3[1]),.dinb(w_G224_0[1]),.dout(n104),.clk(gclk));
	jxor g047(.dina(w_n79_0[0]),.dinb(w_G125_0[1]),.dout(n105),.clk(gclk));
	jxor g048(.dina(n105),.dinb(n104),.dout(n106),.clk(gclk));
	jxor g049(.dina(n106),.dinb(w_n103_0[1]),.dout(n107),.clk(gclk));
	jand g050(.dina(w_n107_0[2]),.dinb(w_n70_2[2]),.dout(n108),.clk(gclk));
	jxor g051(.dina(w_n108_0[1]),.dinb(w_n97_0[1]),.dout(n109),.clk(gclk));
	jand g052(.dina(w_n109_0[1]),.dinb(w_n96_0[2]),.dout(n110),.clk(gclk));
	jnot g053(.din(w_G221_0[0]),.dout(n111),.clk(gclk));
	jor g054(.dina(w_n71_0[0]),.dinb(n111),.dout(n112),.clk(gclk));
	jxor g055(.dina(w_G140_0[1]),.dinb(w_G110_0[2]),.dout(n113),.clk(gclk));
	jand g056(.dina(w_n61_3[0]),.dinb(w_G227_0[1]),.dout(n114),.clk(gclk));
	jxor g057(.dina(n114),.dinb(w_n101_0[0]),.dout(n115),.clk(gclk));
	jxor g058(.dina(n115),.dinb(n113),.dout(n116),.clk(gclk));
	jxor g059(.dina(n116),.dinb(w_n81_0[1]),.dout(n117),.clk(gclk));
	jand g060(.dina(w_n117_0[2]),.dinb(w_n70_2[1]),.dout(n118),.clk(gclk));
	jxor g061(.dina(w_n118_0[1]),.dinb(w_G469_0[2]),.dout(n119),.clk(gclk));
	jand g062(.dina(w_n119_0[1]),.dinb(w_n112_1[1]),.dout(n120),.clk(gclk));
	jand g063(.dina(w_n120_0[1]),.dinb(w_n110_0[2]),.dout(n121),.clk(gclk));
	jand g064(.dina(w_n121_1[1]),.dinb(w_n93_0[2]),.dout(n122),.clk(gclk));
	jnot g065(.din(w_G478_0[2]),.dout(n123),.clk(gclk));
	jxor g066(.dina(w_G143_1[0]),.dinb(w_G128_0[2]),.dout(n124),.clk(gclk));
	jand g067(.dina(w_n62_0[0]),.dinb(w_G217_0[1]),.dout(n125),.clk(gclk));
	jxor g068(.dina(w_G122_1[0]),.dinb(w_G116_0[1]),.dout(n126),.clk(gclk));
	jxor g069(.dina(w_G134_0[1]),.dinb(w_G107_0[1]),.dout(n127),.clk(gclk));
	jxor g070(.dina(n127),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g071(.dina(n128),.dinb(n125),.dout(n129),.clk(gclk));
	jxor g072(.dina(n129),.dinb(n124),.dout(n130),.clk(gclk));
	jand g073(.dina(w_n130_0[2]),.dinb(w_n70_2[0]),.dout(n131),.clk(gclk));
	jxor g074(.dina(w_n131_0[1]),.dinb(n123),.dout(n132),.clk(gclk));
	jnot g075(.din(w_G475_0[2]),.dout(n133),.clk(gclk));
	jxor g076(.dina(w_G143_0[2]),.dinb(w_n77_0[0]),.dout(n134),.clk(gclk));
	jxor g077(.dina(w_G122_0[2]),.dinb(w_n82_0[0]),.dout(n135),.clk(gclk));
	jxor g078(.dina(n135),.dinb(w_G104_0[1]),.dout(n136),.clk(gclk));
	jnot g079(.din(w_G214_0[0]),.dout(n137),.clk(gclk));
	jor g080(.dina(w_n86_0[0]),.dinb(n137),.dout(n138),.clk(gclk));
	jxor g081(.dina(n138),.dinb(w_n60_0[1]),.dout(n139),.clk(gclk));
	jxor g082(.dina(n139),.dinb(n136),.dout(n140),.clk(gclk));
	jxor g083(.dina(n140),.dinb(n134),.dout(n141),.clk(gclk));
	jand g084(.dina(w_n141_0[2]),.dinb(w_n70_1[2]),.dout(n142),.clk(gclk));
	jxor g085(.dina(w_n142_0[1]),.dinb(n133),.dout(n143),.clk(gclk));
	jand g086(.dina(w_n143_1[1]),.dinb(w_n132_0[2]),.dout(n144),.clk(gclk));
	jor g087(.dina(w_n61_2[2]),.dinb(G898),.dout(n145),.clk(gclk));
	jand g088(.dina(w_G237_0[0]),.dinb(w_G234_0[0]),.dout(n146),.clk(gclk));
	jor g089(.dina(w_n146_0[1]),.dinb(w_n70_1[1]),.dout(n147),.clk(gclk));
	jor g090(.dina(w_n147_0[1]),.dinb(w_n145_0[1]),.dout(n148),.clk(gclk));
	jnot g091(.din(w_n146_0[0]),.dout(n149),.clk(gclk));
	jand g092(.dina(w_n61_2[1]),.dinb(w_G952_0[2]),.dout(n150),.clk(gclk));
	jand g093(.dina(n150),.dinb(n149),.dout(n151),.clk(gclk));
	jnot g094(.din(w_n151_0[2]),.dout(n152),.clk(gclk));
	jand g095(.dina(w_n152_0[1]),.dinb(n148),.dout(n153),.clk(gclk));
	jnot g096(.din(w_n153_0[2]),.dout(n154),.clk(gclk));
	jand g097(.dina(w_n154_1[1]),.dinb(w_n144_1[2]),.dout(n155),.clk(gclk));
	jand g098(.dina(w_n155_0[2]),.dinb(w_n122_0[1]),.dout(n156),.clk(gclk));
	jxor g099(.dina(w_n156_0[1]),.dinb(w_G101_0[0]),.dout(w_dff_A_fuse14T61_2),.clk(gclk));
	jnot g100(.din(w_n92_1[1]),.dout(n158),.clk(gclk));
	jand g101(.dina(w_n158_1[1]),.dinb(w_n74_1[0]),.dout(n159),.clk(gclk));
	jand g102(.dina(w_n159_1[1]),.dinb(w_n121_1[0]),.dout(n160),.clk(gclk));
	jxor g103(.dina(w_n142_0[0]),.dinb(w_G475_0[1]),.dout(n161),.clk(gclk));
	jand g104(.dina(w_n161_0[2]),.dinb(w_n132_0[1]),.dout(n162),.clk(gclk));
	jand g105(.dina(w_n162_0[1]),.dinb(w_n154_1[0]),.dout(n163),.clk(gclk));
	jand g106(.dina(w_n163_0[2]),.dinb(w_n160_0[1]),.dout(n164),.clk(gclk));
	jxor g107(.dina(w_n164_0[1]),.dinb(w_G104_0[0]),.dout(w_dff_A_2gaEHoHJ9_2),.clk(gclk));
	jxor g108(.dina(w_n131_0[0]),.dinb(w_G478_0[1]),.dout(n166),.clk(gclk));
	jand g109(.dina(w_n143_1[0]),.dinb(w_n166_1[1]),.dout(n167),.clk(gclk));
	jand g110(.dina(w_n167_0[1]),.dinb(w_n154_0[2]),.dout(n168),.clk(gclk));
	jand g111(.dina(w_n168_0[2]),.dinb(w_n160_0[0]),.dout(n169),.clk(gclk));
	jxor g112(.dina(w_n169_0[1]),.dinb(w_G107_0[0]),.dout(w_dff_A_P8R2qX6l0_2),.clk(gclk));
	jnot g113(.din(w_n60_0[0]),.dout(n171),.clk(gclk));
	jxor g114(.dina(w_n67_0[0]),.dinb(n171),.dout(n172),.clk(gclk));
	jand g115(.dina(w_n172_0[1]),.dinb(w_n70_1[0]),.dout(n173),.clk(gclk));
	jxor g116(.dina(w_n73_0[0]),.dinb(n173),.dout(n174),.clk(gclk));
	jand g117(.dina(w_n158_1[0]),.dinb(w_n174_1[1]),.dout(n175),.clk(gclk));
	jand g118(.dina(w_n175_0[1]),.dinb(w_n155_0[1]),.dout(n176),.clk(gclk));
	jand g119(.dina(n176),.dinb(w_n121_0[2]),.dout(n177),.clk(gclk));
	jxor g120(.dina(w_n177_0[1]),.dinb(w_G110_0[1]),.dout(w_dff_A_Iv1cyd7k5_2),.clk(gclk));
	jand g121(.dina(w_n92_1[0]),.dinb(w_n174_1[0]),.dout(n179),.clk(gclk));
	jand g122(.dina(w_n179_0[2]),.dinb(w_n121_0[1]),.dout(n180),.clk(gclk));
	jor g123(.dina(w_n61_2[0]),.dinb(G900),.dout(n181),.clk(gclk));
	jor g124(.dina(w_n181_0[2]),.dinb(w_n147_0[0]),.dout(n182),.clk(gclk));
	jand g125(.dina(n182),.dinb(w_n152_0[0]),.dout(n183),.clk(gclk));
	jnot g126(.din(w_n183_0[2]),.dout(n184),.clk(gclk));
	jand g127(.dina(w_n184_1[1]),.dinb(w_n167_0[0]),.dout(n185),.clk(gclk));
	jand g128(.dina(w_n185_0[2]),.dinb(w_n180_0[1]),.dout(n186),.clk(gclk));
	jxor g129(.dina(w_n186_0[1]),.dinb(w_G128_0[1]),.dout(w_dff_A_8PLLfsFp3_2),.clk(gclk));
	jand g130(.dina(w_n161_0[1]),.dinb(w_n166_1[0]),.dout(n188),.clk(gclk));
	jand g131(.dina(w_n188_0[2]),.dinb(w_n184_1[0]),.dout(n189),.clk(gclk));
	jand g132(.dina(w_n189_0[1]),.dinb(w_n122_0[0]),.dout(n190),.clk(gclk));
	jxor g133(.dina(w_n190_0[1]),.dinb(w_G143_0[1]),.dout(w_dff_A_uKogXNzU7_2),.clk(gclk));
	jand g134(.dina(w_n184_0[2]),.dinb(w_n162_0[0]),.dout(n192),.clk(gclk));
	jand g135(.dina(w_n192_0[2]),.dinb(w_n180_0[0]),.dout(n193),.clk(gclk));
	jxor g136(.dina(w_n193_0[1]),.dinb(w_G146_0[0]),.dout(w_dff_A_b9MQohhs2_2),.clk(gclk));
	jnot g137(.din(w_G469_0[1]),.dout(n195),.clk(gclk));
	jxor g138(.dina(w_n118_0[0]),.dinb(n195),.dout(n196),.clk(gclk));
	jand g139(.dina(w_n196_0[2]),.dinb(w_n112_1[0]),.dout(n197),.clk(gclk));
	jand g140(.dina(w_n197_1[1]),.dinb(w_n110_0[1]),.dout(n198),.clk(gclk));
	jand g141(.dina(w_n198_1[1]),.dinb(w_n93_0[1]),.dout(n199),.clk(gclk));
	jand g142(.dina(w_n199_0[1]),.dinb(w_n163_0[1]),.dout(n200),.clk(gclk));
	jxor g143(.dina(w_n200_0[1]),.dinb(w_G113_0[0]),.dout(w_dff_A_30rl8IDl4_2),.clk(gclk));
	jand g144(.dina(w_n199_0[0]),.dinb(w_n168_0[1]),.dout(n202),.clk(gclk));
	jxor g145(.dina(w_n202_0[1]),.dinb(w_G116_0[0]),.dout(w_dff_A_cPpb56RY3_2),.clk(gclk));
	jand g146(.dina(w_n198_1[0]),.dinb(w_n179_0[1]),.dout(n204),.clk(gclk));
	jand g147(.dina(n204),.dinb(w_n155_0[0]),.dout(n205),.clk(gclk));
	jxor g148(.dina(w_n205_0[1]),.dinb(w_G119_0[0]),.dout(w_dff_A_vWFS0OZ25_2),.clk(gclk));
	jand g149(.dina(w_n197_1[0]),.dinb(w_n159_1[0]),.dout(n207),.clk(gclk));
	jand g150(.dina(w_n154_0[1]),.dinb(w_n110_0[0]),.dout(n208),.clk(gclk));
	jand g151(.dina(n208),.dinb(w_n188_0[1]),.dout(n209),.clk(gclk));
	jand g152(.dina(n209),.dinb(w_n207_0[1]),.dout(n210),.clk(gclk));
	jxor g153(.dina(w_n210_0[1]),.dinb(w_G122_0[1]),.dout(w_dff_A_fXWr2Uu04_2),.clk(gclk));
	jand g154(.dina(w_n192_0[1]),.dinb(w_n175_0[0]),.dout(n212),.clk(gclk));
	jand g155(.dina(w_n212_0[1]),.dinb(w_n198_0[2]),.dout(n213),.clk(gclk));
	jxor g156(.dina(w_n213_0[1]),.dinb(w_G125_0[0]),.dout(w_dff_A_E9NAXxXK0_2),.clk(gclk));
	jnot g157(.din(w_n97_0[0]),.dout(n215),.clk(gclk));
	jxor g158(.dina(w_n108_0[0]),.dinb(n215),.dout(n216),.clk(gclk));
	jand g159(.dina(w_n216_0[2]),.dinb(w_n96_0[1]),.dout(n217),.clk(gclk));
	jand g160(.dina(w_n217_0[2]),.dinb(w_n120_0[0]),.dout(n218),.clk(gclk));
	jand g161(.dina(w_n218_1[1]),.dinb(w_n93_0[0]),.dout(n219),.clk(gclk));
	jand g162(.dina(w_n219_0[1]),.dinb(w_n192_0[0]),.dout(n220),.clk(gclk));
	jxor g163(.dina(w_n220_0[1]),.dinb(w_G131_0[0]),.dout(w_dff_A_jF9YHq5j2_2),.clk(gclk));
	jand g164(.dina(w_n219_0[0]),.dinb(w_n185_0[1]),.dout(n222),.clk(gclk));
	jxor g165(.dina(w_n222_0[1]),.dinb(w_G134_0[0]),.dout(w_dff_A_CObwD37Y6_2),.clk(gclk));
	jand g166(.dina(w_n184_0[1]),.dinb(w_n144_1[1]),.dout(n224),.clk(gclk));
	jand g167(.dina(n224),.dinb(w_n179_0[0]),.dout(n225),.clk(gclk));
	jand g168(.dina(n225),.dinb(w_n218_1[0]),.dout(n226),.clk(gclk));
	jxor g169(.dina(w_n226_0[1]),.dinb(w_G137_0[0]),.dout(w_dff_A_9pyUhmRS8_2),.clk(gclk));
	jand g170(.dina(w_n218_0[2]),.dinb(w_n212_0[0]),.dout(n228),.clk(gclk));
	jxor g171(.dina(w_n228_0[1]),.dinb(w_G140_0[0]),.dout(w_dff_A_bMjqVEuP0_2),.clk(gclk));
	jor g172(.dina(w_n177_0[0]),.dinb(w_n169_0[0]),.dout(n230),.clk(gclk));
	jor g173(.dina(w_n202_0[0]),.dinb(w_n164_0[0]),.dout(n231),.clk(gclk));
	jor g174(.dina(n231),.dinb(n230),.dout(n232),.clk(gclk));
	jor g175(.dina(w_n205_0[0]),.dinb(w_n156_0[0]),.dout(n233),.clk(gclk));
	jor g176(.dina(w_n210_0[0]),.dinb(w_n200_0[0]),.dout(n234),.clk(gclk));
	jor g177(.dina(n234),.dinb(n233),.dout(n235),.clk(gclk));
	jor g178(.dina(n235),.dinb(n232),.dout(n236),.clk(gclk));
	jor g179(.dina(w_n220_0[0]),.dinb(w_n193_0[0]),.dout(n237),.clk(gclk));
	jor g180(.dina(w_n222_0[0]),.dinb(w_n186_0[0]),.dout(n238),.clk(gclk));
	jor g181(.dina(n238),.dinb(n237),.dout(n239),.clk(gclk));
	jor g182(.dina(w_n228_0[0]),.dinb(w_n190_0[0]),.dout(n240),.clk(gclk));
	jor g183(.dina(w_n226_0[0]),.dinb(w_n213_0[0]),.dout(n241),.clk(gclk));
	jor g184(.dina(n241),.dinb(n240),.dout(n242),.clk(gclk));
	jor g185(.dina(n242),.dinb(n239),.dout(n243),.clk(gclk));
	jor g186(.dina(n243),.dinb(n236),.dout(n244),.clk(gclk));
	jor g187(.dina(w_n218_0[1]),.dinb(w_n198_0[1]),.dout(n245),.clk(gclk));
	jand g188(.dina(n245),.dinb(w_n144_1[0]),.dout(n246),.clk(gclk));
	jand g189(.dina(w_n217_0[1]),.dinb(w_n197_0[2]),.dout(n247),.clk(gclk));
	jxor g190(.dina(w_n143_0[2]),.dinb(w_n132_0[0]),.dout(n248),.clk(gclk));
	jand g191(.dina(n248),.dinb(n247),.dout(n249),.clk(gclk));
	jor g192(.dina(n249),.dinb(n246),.dout(n250),.clk(gclk));
	jand g193(.dina(n250),.dinb(w_n159_0[2]),.dout(n251),.clk(gclk));
	jand g194(.dina(w_n217_0[0]),.dinb(w_n144_0[2]),.dout(n252),.clk(gclk));
	jor g195(.dina(w_n92_0[2]),.dinb(w_n174_0[2]),.dout(n253),.clk(gclk));
	jor g196(.dina(w_n158_0[2]),.dinb(w_n74_0[2]),.dout(n254),.clk(gclk));
	jand g197(.dina(w_n197_0[1]),.dinb(w_n254_1[1]),.dout(n255),.clk(gclk));
	jand g198(.dina(n255),.dinb(w_n253_0[2]),.dout(n256),.clk(gclk));
	jand g199(.dina(n256),.dinb(w_n252_0[1]),.dout(n257),.clk(gclk));
	jor g200(.dina(n257),.dinb(n251),.dout(n258),.clk(gclk));
	jand g201(.dina(n258),.dinb(w_n151_0[1]),.dout(n259),.clk(gclk));
	jxor g202(.dina(w_n112_0[2]),.dinb(w_n96_0[0]),.dout(n260),.clk(gclk));
	jand g203(.dina(n260),.dinb(w_n151_0[0]),.dout(n261),.clk(gclk));
	jand g204(.dina(n261),.dinb(w_n196_0[1]),.dout(n262),.clk(gclk));
	jand g205(.dina(n262),.dinb(w_n216_0[1]),.dout(n263),.clk(gclk));
	jand g206(.dina(w_n159_0[1]),.dinb(w_n144_0[1]),.dout(n264),.clk(gclk));
	jand g207(.dina(n264),.dinb(n263),.dout(n265),.clk(gclk));
	jor g208(.dina(n265),.dinb(n259),.dout(n266),.clk(gclk));
	jor g209(.dina(n266),.dinb(w_n244_2[2]),.dout(n267),.clk(gclk));
	jand g210(.dina(n267),.dinb(w_G952_0[1]),.dout(n268),.clk(gclk));
	jand g211(.dina(w_n252_0[0]),.dinb(w_n207_0[0]),.dout(n269),.clk(gclk));
	jor g212(.dina(n269),.dinb(w_G953_1[0]),.dout(n270),.clk(gclk));
	jor g213(.dina(w_dff_B_hos9PQp09_0),.dinb(n268),.dout(w_dff_A_T9z38KbT5_2),.clk(gclk));
	jnot g214(.din(w_n107_0[1]),.dout(n272),.clk(gclk));
	jor g215(.dina(w_n216_0[0]),.dinb(w_n95_0[1]),.dout(n273),.clk(gclk));
	jnot g216(.din(w_n112_0[1]),.dout(n274),.clk(gclk));
	jor g217(.dina(w_n196_0[0]),.dinb(w_n274_0[1]),.dout(n275),.clk(gclk));
	jor g218(.dina(w_n275_0[1]),.dinb(w_n273_0[2]),.dout(n276),.clk(gclk));
	jor g219(.dina(w_n253_0[1]),.dinb(w_n276_1[1]),.dout(n277),.clk(gclk));
	jnot g220(.din(w_n168_0[0]),.dout(n278),.clk(gclk));
	jor g221(.dina(w_n278_0[1]),.dinb(w_n277_0[1]),.dout(n279),.clk(gclk));
	jor g222(.dina(w_n161_0[0]),.dinb(w_n166_0[2]),.dout(n280),.clk(gclk));
	jor g223(.dina(w_n153_0[1]),.dinb(w_n280_0[1]),.dout(n281),.clk(gclk));
	jor g224(.dina(w_n92_0[1]),.dinb(w_n74_0[1]),.dout(n282),.clk(gclk));
	jor g225(.dina(w_n282_0[1]),.dinb(w_n281_0[2]),.dout(n283),.clk(gclk));
	jor g226(.dina(n283),.dinb(w_n276_1[0]),.dout(n284),.clk(gclk));
	jand g227(.dina(n284),.dinb(n279),.dout(n285),.clk(gclk));
	jnot g228(.din(w_n163_0[0]),.dout(n286),.clk(gclk));
	jor g229(.dina(w_n286_0[1]),.dinb(w_n277_0[0]),.dout(n287),.clk(gclk));
	jor g230(.dina(w_n158_0[1]),.dinb(w_n174_0[1]),.dout(n288),.clk(gclk));
	jor g231(.dina(w_n119_0[0]),.dinb(w_n274_0[0]),.dout(n289),.clk(gclk));
	jor g232(.dina(w_n289_0[1]),.dinb(w_n273_0[1]),.dout(n290),.clk(gclk));
	jor g233(.dina(w_n290_0[2]),.dinb(w_n288_0[2]),.dout(n291),.clk(gclk));
	jor g234(.dina(w_n291_0[1]),.dinb(w_n278_0[0]),.dout(n292),.clk(gclk));
	jand g235(.dina(n292),.dinb(n287),.dout(n293),.clk(gclk));
	jand g236(.dina(n293),.dinb(n285),.dout(n294),.clk(gclk));
	jor g237(.dina(w_n276_0[2]),.dinb(w_n288_0[1]),.dout(n295),.clk(gclk));
	jor g238(.dina(w_n281_0[1]),.dinb(w_n295_0[1]),.dout(n296),.clk(gclk));
	jor g239(.dina(w_n290_0[1]),.dinb(w_n254_1[0]),.dout(n297),.clk(gclk));
	jor g240(.dina(n297),.dinb(w_n281_0[0]),.dout(n298),.clk(gclk));
	jand g241(.dina(n298),.dinb(n296),.dout(n299),.clk(gclk));
	jor g242(.dina(w_n291_0[0]),.dinb(w_n286_0[0]),.dout(n300),.clk(gclk));
	jor g243(.dina(w_n289_0[0]),.dinb(w_n253_0[0]),.dout(n301),.clk(gclk));
	jnot g244(.din(w_n188_0[0]),.dout(n302),.clk(gclk));
	jor g245(.dina(w_n153_0[0]),.dinb(w_n273_0[0]),.dout(n303),.clk(gclk));
	jor g246(.dina(n303),.dinb(n302),.dout(n304),.clk(gclk));
	jor g247(.dina(n304),.dinb(n301),.dout(n305),.clk(gclk));
	jand g248(.dina(n305),.dinb(n300),.dout(n306),.clk(gclk));
	jand g249(.dina(n306),.dinb(n299),.dout(n307),.clk(gclk));
	jand g250(.dina(n307),.dinb(n294),.dout(n308),.clk(gclk));
	jor g251(.dina(w_n254_0[2]),.dinb(w_n276_0[1]),.dout(n309),.clk(gclk));
	jor g252(.dina(w_n143_0[1]),.dinb(w_n166_0[1]),.dout(n310),.clk(gclk));
	jor g253(.dina(w_n183_0[1]),.dinb(n310),.dout(n311),.clk(gclk));
	jor g254(.dina(w_n311_0[2]),.dinb(w_n309_0[1]),.dout(n312),.clk(gclk));
	jor g255(.dina(w_n109_0[0]),.dinb(w_n95_0[0]),.dout(n313),.clk(gclk));
	jor g256(.dina(n313),.dinb(w_n275_0[0]),.dout(n314),.clk(gclk));
	jor g257(.dina(w_n314_0[2]),.dinb(w_n288_0[0]),.dout(n315),.clk(gclk));
	jor g258(.dina(w_n315_0[1]),.dinb(w_n311_0[1]),.dout(n316),.clk(gclk));
	jand g259(.dina(n316),.dinb(n312),.dout(n317),.clk(gclk));
	jnot g260(.din(w_n185_0[0]),.dout(n318),.clk(gclk));
	jor g261(.dina(w_n318_0[1]),.dinb(w_n309_0[0]),.dout(n319),.clk(gclk));
	jor g262(.dina(w_n315_0[0]),.dinb(w_n318_0[0]),.dout(n320),.clk(gclk));
	jand g263(.dina(n320),.dinb(n319),.dout(n321),.clk(gclk));
	jand g264(.dina(n321),.dinb(n317),.dout(n322),.clk(gclk));
	jnot g265(.din(w_n189_0[0]),.dout(n323),.clk(gclk));
	jor g266(.dina(n323),.dinb(w_n295_0[0]),.dout(n324),.clk(gclk));
	jor g267(.dina(w_n311_0[0]),.dinb(w_n282_0[0]),.dout(n325),.clk(gclk));
	jor g268(.dina(w_n314_0[1]),.dinb(w_n325_0[1]),.dout(n326),.clk(gclk));
	jand g269(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jor g270(.dina(w_n325_0[0]),.dinb(w_n290_0[0]),.dout(n328),.clk(gclk));
	jor g271(.dina(w_n183_0[0]),.dinb(w_n280_0[0]),.dout(n329),.clk(gclk));
	jor g272(.dina(n329),.dinb(w_n254_0[1]),.dout(n330),.clk(gclk));
	jor g273(.dina(n330),.dinb(w_n314_0[0]),.dout(n331),.clk(gclk));
	jand g274(.dina(n331),.dinb(n328),.dout(n332),.clk(gclk));
	jand g275(.dina(n332),.dinb(n327),.dout(n333),.clk(gclk));
	jand g276(.dina(n333),.dinb(n322),.dout(n334),.clk(gclk));
	jand g277(.dina(w_n334_0[1]),.dinb(w_n308_0[1]),.dout(n335),.clk(gclk));
	jand g278(.dina(w_G902_2[2]),.dinb(w_G210_0[0]),.dout(n336),.clk(gclk));
	jnot g279(.din(w_n336_0[1]),.dout(n337),.clk(gclk));
	jor g280(.dina(n337),.dinb(w_n335_2[1]),.dout(n338),.clk(gclk));
	jor g281(.dina(n338),.dinb(n272),.dout(n339),.clk(gclk));
	jor g282(.dina(w_n61_1[2]),.dinb(w_G952_0[0]),.dout(n340),.clk(gclk));
	jand g283(.dina(w_n336_0[0]),.dinb(w_n244_2[1]),.dout(n341),.clk(gclk));
	jor g284(.dina(n341),.dinb(w_n107_0[0]),.dout(n342),.clk(gclk));
	jand g285(.dina(n342),.dinb(w_n340_2[1]),.dout(n343),.clk(gclk));
	jand g286(.dina(n343),.dinb(w_dff_B_2orChbYK1_1),.dout(G51),.clk(gclk));
	jnot g287(.din(w_n117_0[1]),.dout(n345),.clk(gclk));
	jand g288(.dina(w_G902_2[1]),.dinb(w_G469_0[0]),.dout(n346),.clk(gclk));
	jnot g289(.din(w_n346_0[1]),.dout(n347),.clk(gclk));
	jor g290(.dina(n347),.dinb(w_n335_2[0]),.dout(n348),.clk(gclk));
	jor g291(.dina(n348),.dinb(n345),.dout(n349),.clk(gclk));
	jand g292(.dina(w_n346_0[0]),.dinb(w_n244_2[0]),.dout(n350),.clk(gclk));
	jor g293(.dina(n350),.dinb(w_n117_0[0]),.dout(n351),.clk(gclk));
	jand g294(.dina(n351),.dinb(w_n340_2[0]),.dout(n352),.clk(gclk));
	jand g295(.dina(n352),.dinb(w_dff_B_kjsma4km9_1),.dout(G54),.clk(gclk));
	jnot g296(.din(w_n141_0[1]),.dout(n354),.clk(gclk));
	jand g297(.dina(w_G902_2[0]),.dinb(w_G475_0[0]),.dout(n355),.clk(gclk));
	jnot g298(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jor g299(.dina(n356),.dinb(w_n335_1[2]),.dout(n357),.clk(gclk));
	jor g300(.dina(n357),.dinb(n354),.dout(n358),.clk(gclk));
	jand g301(.dina(w_n355_0[0]),.dinb(w_n244_1[2]),.dout(n359),.clk(gclk));
	jor g302(.dina(n359),.dinb(w_n141_0[0]),.dout(n360),.clk(gclk));
	jand g303(.dina(n360),.dinb(w_n340_1[2]),.dout(n361),.clk(gclk));
	jand g304(.dina(n361),.dinb(w_dff_B_CqM0mfmv2_1),.dout(G60),.clk(gclk));
	jnot g305(.din(w_n130_0[1]),.dout(n363),.clk(gclk));
	jand g306(.dina(w_G902_1[2]),.dinb(w_G478_0[0]),.dout(n364),.clk(gclk));
	jnot g307(.din(w_n364_0[1]),.dout(n365),.clk(gclk));
	jor g308(.dina(n365),.dinb(w_n335_1[1]),.dout(n366),.clk(gclk));
	jor g309(.dina(n366),.dinb(n363),.dout(n367),.clk(gclk));
	jand g310(.dina(w_n364_0[0]),.dinb(w_n244_1[1]),.dout(n368),.clk(gclk));
	jor g311(.dina(n368),.dinb(w_n130_0[0]),.dout(n369),.clk(gclk));
	jand g312(.dina(n369),.dinb(w_n340_1[1]),.dout(n370),.clk(gclk));
	jand g313(.dina(n370),.dinb(w_dff_B_kssSIq840_1),.dout(G63),.clk(gclk));
	jand g314(.dina(w_G902_1[1]),.dinb(w_G217_0[0]),.dout(n372),.clk(gclk));
	jand g315(.dina(w_n372_0[1]),.dinb(w_n244_1[0]),.dout(n373),.clk(gclk));
	jor g316(.dina(n373),.dinb(w_n172_0[0]),.dout(n374),.clk(gclk));
	jnot g317(.din(w_n372_0[0]),.dout(n375),.clk(gclk));
	jor g318(.dina(n375),.dinb(w_n335_1[0]),.dout(n376),.clk(gclk));
	jor g319(.dina(n376),.dinb(w_n68_0[0]),.dout(n377),.clk(gclk));
	jand g320(.dina(n377),.dinb(w_n340_1[0]),.dout(n378),.clk(gclk));
	jand g321(.dina(n378),.dinb(w_dff_B_29RFV7IF1_1),.dout(G66),.clk(gclk));
	jnot g322(.din(w_n145_0[0]),.dout(n380),.clk(gclk));
	jor g323(.dina(w_n308_0[0]),.dinb(w_G953_0[2]),.dout(n381),.clk(gclk));
	jor g324(.dina(w_n61_1[1]),.dinb(w_G224_0[0]),.dout(n382),.clk(gclk));
	jand g325(.dina(n382),.dinb(n381),.dout(n383),.clk(gclk));
	jxor g326(.dina(n383),.dinb(w_n103_0[0]),.dout(n384),.clk(gclk));
	jor g327(.dina(n384),.dinb(w_dff_B_LumDwg734_1),.dout(w_dff_A_wZn0xXb02_2),.clk(gclk));
	jor g328(.dina(w_n334_0[0]),.dinb(w_G953_0[1]),.dout(n386),.clk(gclk));
	jor g329(.dina(w_n61_1[0]),.dinb(w_G227_0[0]),.dout(n387),.clk(gclk));
	jand g330(.dina(n387),.dinb(w_n181_0[1]),.dout(n388),.clk(gclk));
	jand g331(.dina(n388),.dinb(n386),.dout(n389),.clk(gclk));
	jnot g332(.din(w_n181_0[0]),.dout(n390),.clk(gclk));
	jxor g333(.dina(w_n81_0[0]),.dinb(w_n59_0[0]),.dout(n391),.clk(gclk));
	jor g334(.dina(n391),.dinb(n390),.dout(n392),.clk(gclk));
	jxor g335(.dina(w_dff_B_dlWi642E9_0),.dinb(n389),.dout(w_dff_A_EFbnONC66_2),.clk(gclk));
	jnot g336(.din(w_n90_0[1]),.dout(n394),.clk(gclk));
	jand g337(.dina(w_G902_1[0]),.dinb(w_G472_0[0]),.dout(n395),.clk(gclk));
	jnot g338(.din(w_n395_0[1]),.dout(n396),.clk(gclk));
	jor g339(.dina(n396),.dinb(w_n335_0[2]),.dout(n397),.clk(gclk));
	jor g340(.dina(n397),.dinb(n394),.dout(n398),.clk(gclk));
	jand g341(.dina(w_n395_0[0]),.dinb(w_n244_0[2]),.dout(n399),.clk(gclk));
	jor g342(.dina(n399),.dinb(w_n90_0[0]),.dout(n400),.clk(gclk));
	jand g343(.dina(n400),.dinb(w_n340_0[2]),.dout(n401),.clk(gclk));
	jand g344(.dina(n401),.dinb(w_dff_B_9rmQ04lU6_1),.dout(G57),.clk(gclk));
	jspl3 jspl3_w_G101_0(.douta(w_G101_0[0]),.doutb(w_G101_0[1]),.doutc(w_G101_0[2]),.din(G101));
	jspl3 jspl3_w_G104_0(.douta(w_G104_0[0]),.doutb(w_G104_0[1]),.doutc(w_G104_0[2]),.din(G104));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_G107_0[1]),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G110_0(.douta(w_G110_0[0]),.doutb(w_G110_0[1]),.doutc(w_G110_0[2]),.din(G110));
	jspl jspl_w_G110_1(.douta(w_G110_1[0]),.doutb(w_G110_1[1]),.din(w_G110_0[0]));
	jspl jspl_w_G113_0(.douta(w_G113_0[0]),.doutb(w_G113_0[1]),.din(G113));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_G116_0[1]),.doutc(w_G116_0[2]),.din(G116));
	jspl3 jspl3_w_G119_0(.douta(w_G119_0[0]),.doutb(w_G119_0[1]),.doutc(w_G119_0[2]),.din(G119));
	jspl3 jspl3_w_G122_0(.douta(w_G122_0[0]),.doutb(w_G122_0[1]),.doutc(w_G122_0[2]),.din(G122));
	jspl jspl_w_G122_1(.douta(w_G122_1[0]),.doutb(w_G122_1[1]),.din(w_G122_0[0]));
	jspl3 jspl3_w_G125_0(.douta(w_G125_0[0]),.doutb(w_G125_0[1]),.doutc(w_G125_0[2]),.din(G125));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(G128));
	jspl jspl_w_G128_1(.douta(w_G128_1[0]),.doutb(w_G128_1[1]),.din(w_G128_0[0]));
	jspl jspl_w_G131_0(.douta(w_G131_0[0]),.doutb(w_G131_0[1]),.din(G131));
	jspl3 jspl3_w_G134_0(.douta(w_G134_0[0]),.doutb(w_G134_0[1]),.doutc(w_G134_0[2]),.din(G134));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G140_0(.douta(w_G140_0[0]),.doutb(w_G140_0[1]),.doutc(w_G140_0[2]),.din(G140));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(G143));
	jspl jspl_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.din(w_G143_0[0]));
	jspl3 jspl3_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.doutc(w_G146_0[2]),.din(G146));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_G210_0[2]),.din(G210));
	jspl jspl_w_G214_0(.douta(w_G214_0[0]),.doutb(w_G214_0[1]),.din(G214));
	jspl3 jspl3_w_G217_0(.douta(w_G217_0[0]),.doutb(w_G217_0[1]),.doutc(w_G217_0[2]),.din(G217));
	jspl jspl_w_G221_0(.douta(w_G221_0[0]),.doutb(w_G221_0[1]),.din(G221));
	jspl jspl_w_G224_0(.douta(w_G224_0[0]),.doutb(w_G224_0[1]),.din(G224));
	jspl jspl_w_G227_0(.douta(w_G227_0[0]),.doutb(w_G227_0[1]),.din(G227));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_G234_0[2]),.din(G234));
	jspl3 jspl3_w_G237_0(.douta(w_G237_0[0]),.doutb(w_G237_0[1]),.doutc(w_G237_0[2]),.din(G237));
	jspl3 jspl3_w_G469_0(.douta(w_G469_0[0]),.doutb(w_G469_0[1]),.doutc(w_G469_0[2]),.din(G469));
	jspl jspl_w_G472_0(.douta(w_G472_0[0]),.doutb(w_G472_0[1]),.din(G472));
	jspl3 jspl3_w_G475_0(.douta(w_G475_0[0]),.doutb(w_G475_0[1]),.doutc(w_G475_0[2]),.din(G475));
	jspl3 jspl3_w_G478_0(.douta(w_G478_0[0]),.doutb(w_G478_0[1]),.doutc(w_G478_0[2]),.din(G478));
	jspl3 jspl3_w_G902_0(.douta(w_G902_0[0]),.doutb(w_G902_0[1]),.doutc(w_G902_0[2]),.din(G902));
	jspl3 jspl3_w_G902_1(.douta(w_G902_1[0]),.doutb(w_G902_1[1]),.doutc(w_G902_1[2]),.din(w_G902_0[0]));
	jspl3 jspl3_w_G902_2(.douta(w_G902_2[0]),.doutb(w_G902_2[1]),.doutc(w_G902_2[2]),.din(w_G902_0[1]));
	jspl3 jspl3_w_G902_3(.douta(w_G902_3[0]),.doutb(w_G902_3[1]),.doutc(w_G902_3[2]),.din(w_G902_0[2]));
	jspl3 jspl3_w_G952_0(.douta(w_G952_0[0]),.doutb(w_G952_0[1]),.doutc(w_G952_0[2]),.din(G952));
	jspl3 jspl3_w_G953_0(.douta(w_G953_0[0]),.doutb(w_G953_0[1]),.doutc(w_G953_0[2]),.din(G953));
	jspl3 jspl3_w_G953_1(.douta(w_G953_1[0]),.doutb(w_G953_1[1]),.doutc(w_G953_1[2]),.din(w_G953_0[0]));
	jspl jspl_w_n59_0(.douta(w_n59_0[0]),.doutb(w_n59_0[1]),.din(n59));
	jspl3 jspl3_w_n60_0(.douta(w_n60_0[0]),.doutb(w_n60_0[1]),.doutc(w_n60_0[2]),.din(n60));
	jspl3 jspl3_w_n61_0(.douta(w_n61_0[0]),.doutb(w_n61_0[1]),.doutc(w_n61_0[2]),.din(n61));
	jspl3 jspl3_w_n61_1(.douta(w_n61_1[0]),.doutb(w_n61_1[1]),.doutc(w_n61_1[2]),.din(w_n61_0[0]));
	jspl3 jspl3_w_n61_2(.douta(w_n61_2[0]),.doutb(w_n61_2[1]),.doutc(w_n61_2[2]),.din(w_n61_0[1]));
	jspl3 jspl3_w_n61_3(.douta(w_n61_3[0]),.doutb(w_n61_3[1]),.doutc(w_n61_3[2]),.din(w_n61_0[2]));
	jspl jspl_w_n62_0(.douta(w_n62_0[0]),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n68_0(.douta(w_n68_0[0]),.doutb(w_n68_0[1]),.din(n68));
	jspl3 jspl3_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.doutc(w_n70_0[2]),.din(n70));
	jspl3 jspl3_w_n70_1(.douta(w_n70_1[0]),.doutb(w_n70_1[1]),.doutc(w_n70_1[2]),.din(w_n70_0[0]));
	jspl3 jspl3_w_n70_2(.douta(w_n70_2[0]),.doutb(w_n70_2[1]),.doutc(w_n70_2[2]),.din(w_n70_0[1]));
	jspl jspl_w_n70_3(.douta(w_n70_3[0]),.doutb(w_n70_3[1]),.din(w_n70_0[2]));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(n73));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n79_0(.douta(w_n79_0[0]),.doutb(w_n79_0[1]),.din(n79));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl jspl_w_n82_0(.douta(w_n82_0[0]),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl3 jspl3_w_n92_1(.douta(w_n92_1[0]),.doutb(w_n92_1[1]),.doutc(w_n92_1[2]),.din(w_n92_0[0]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl3 jspl3_w_n95_0(.douta(w_n95_0[0]),.doutb(w_n95_0[1]),.doutc(w_n95_0[2]),.din(n95));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.doutc(w_n96_0[2]),.din(n96));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.din(n103));
	jspl3 jspl3_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.doutc(w_n107_0[2]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.doutc(w_n110_0[2]),.din(n110));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl jspl_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.din(n118));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl jspl_w_n121_1(.douta(w_n121_1[0]),.doutb(w_n121_1[1]),.din(w_n121_0[0]));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.din(n122));
	jspl3 jspl3_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.doutc(w_n130_0[2]),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl3 jspl3_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.doutc(w_n143_0[2]),.din(n143));
	jspl jspl_w_n143_1(.douta(w_n143_1[0]),.doutb(w_n143_1[1]),.din(w_n143_0[0]));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n144_1(.douta(w_n144_1[0]),.doutb(w_n144_1[1]),.doutc(w_n144_1[2]),.din(w_n144_0[0]));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.doutc(w_n151_0[2]),.din(n151));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_n154_0[2]),.din(n154));
	jspl jspl_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.din(w_n154_0[0]));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.doutc(w_n158_0[2]),.din(n158));
	jspl jspl_w_n158_1(.douta(w_n158_1[0]),.doutb(w_n158_1[1]),.din(w_n158_0[0]));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_n163_0[2]),.din(n163));
	jspl jspl_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.din(n164));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl jspl_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.din(w_n166_0[0]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl3 jspl3_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.doutc(w_n174_0[2]),.din(n174));
	jspl jspl_w_n174_1(.douta(w_n174_1[0]),.doutb(w_n174_1[1]),.din(w_n174_0[0]));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_n179_0[1]),.doutc(w_n179_0[2]),.din(n179));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n183_0(.douta(w_n183_0[0]),.doutb(w_n183_0[1]),.doutc(w_n183_0[2]),.din(n183));
	jspl3 jspl3_w_n184_0(.douta(w_n184_0[0]),.doutb(w_n184_0[1]),.doutc(w_n184_0[2]),.din(n184));
	jspl jspl_w_n184_1(.douta(w_n184_1[0]),.doutb(w_n184_1[1]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.doutc(w_n185_0[2]),.din(n185));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl3 jspl3_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.doutc(w_n188_0[2]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.doutc(w_n192_0[2]),.din(n192));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.din(n193));
	jspl3 jspl3_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.doutc(w_n196_0[2]),.din(n196));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_n197_1[0]),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_n198_0[2]),.din(n198));
	jspl jspl_w_n198_1(.douta(w_n198_1[0]),.doutb(w_n198_1[1]),.din(w_n198_0[0]));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(n202));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.doutc(w_n216_0[2]),.din(n216));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_n218_0[2]),.din(n218));
	jspl jspl_w_n218_1(.douta(w_n218_1[0]),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.din(n222));
	jspl jspl_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl3 jspl3_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.doutc(w_n244_0[2]),.din(n244));
	jspl3 jspl3_w_n244_1(.douta(w_n244_1[0]),.doutb(w_n244_1[1]),.doutc(w_n244_1[2]),.din(w_n244_0[0]));
	jspl3 jspl3_w_n244_2(.douta(w_n244_2[0]),.doutb(w_n244_2[1]),.doutc(w_n244_2[2]),.din(w_n244_0[1]));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl3 jspl3_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.doutc(w_n253_0[2]),.din(n253));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl jspl_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.doutc(w_n273_0[2]),.din(n273));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl3 jspl3_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.doutc(w_n276_0[2]),.din(n276));
	jspl jspl_w_n276_1(.douta(w_n276_1[0]),.doutb(w_n276_1[1]),.din(w_n276_0[0]));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.din(n278));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.doutc(w_n281_0[2]),.din(n281));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.din(n286));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.din(n289));
	jspl3 jspl3_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.doutc(w_n290_0[2]),.din(n290));
	jspl jspl_w_n291_0(.douta(w_n291_0[0]),.doutb(w_n291_0[1]),.din(n291));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(n295));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(n309));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.doutc(w_n311_0[2]),.din(n311));
	jspl3 jspl3_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.doutc(w_n314_0[2]),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.doutc(w_n335_1[2]),.din(w_n335_0[0]));
	jspl jspl_w_n335_2(.douta(w_n335_2[0]),.doutb(w_n335_2[1]),.din(w_n335_0[1]));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl3 jspl3_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.doutc(w_n340_0[2]),.din(n340));
	jspl3 jspl3_w_n340_1(.douta(w_n340_1[0]),.doutb(w_n340_1[1]),.doutc(w_n340_1[2]),.din(w_n340_0[0]));
	jspl jspl_w_n340_2(.douta(w_n340_2[0]),.doutb(w_n340_2[1]),.din(w_n340_0[1]));
	jspl jspl_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n395_0(.douta(w_n395_0[0]),.doutb(w_n395_0[1]),.din(n395));
	jdff dff_B_ZVKO1Mo51_0(.din(n270),.dout(w_dff_B_ZVKO1Mo51_0),.clk(gclk));
	jdff dff_B_Bnhasfkr6_0(.din(w_dff_B_ZVKO1Mo51_0),.dout(w_dff_B_Bnhasfkr6_0),.clk(gclk));
	jdff dff_B_P396Rp8F4_0(.din(w_dff_B_Bnhasfkr6_0),.dout(w_dff_B_P396Rp8F4_0),.clk(gclk));
	jdff dff_B_GO4wAQ8u2_0(.din(w_dff_B_P396Rp8F4_0),.dout(w_dff_B_GO4wAQ8u2_0),.clk(gclk));
	jdff dff_B_hos9PQp09_0(.din(w_dff_B_GO4wAQ8u2_0),.dout(w_dff_B_hos9PQp09_0),.clk(gclk));
	jdff dff_B_2orChbYK1_1(.din(n339),.dout(w_dff_B_2orChbYK1_1),.clk(gclk));
	jdff dff_B_kjsma4km9_1(.din(n349),.dout(w_dff_B_kjsma4km9_1),.clk(gclk));
	jdff dff_B_CqM0mfmv2_1(.din(n358),.dout(w_dff_B_CqM0mfmv2_1),.clk(gclk));
	jdff dff_B_kssSIq840_1(.din(n367),.dout(w_dff_B_kssSIq840_1),.clk(gclk));
	jdff dff_B_29RFV7IF1_1(.din(n374),.dout(w_dff_B_29RFV7IF1_1),.clk(gclk));
	jdff dff_B_dzWAwNCf7_1(.din(n380),.dout(w_dff_B_dzWAwNCf7_1),.clk(gclk));
	jdff dff_B_BZfl0Bnq5_1(.din(w_dff_B_dzWAwNCf7_1),.dout(w_dff_B_BZfl0Bnq5_1),.clk(gclk));
	jdff dff_B_6RKKJuU99_1(.din(w_dff_B_BZfl0Bnq5_1),.dout(w_dff_B_6RKKJuU99_1),.clk(gclk));
	jdff dff_B_b0kIoAb76_1(.din(w_dff_B_6RKKJuU99_1),.dout(w_dff_B_b0kIoAb76_1),.clk(gclk));
	jdff dff_B_Le1XJwK91_1(.din(w_dff_B_b0kIoAb76_1),.dout(w_dff_B_Le1XJwK91_1),.clk(gclk));
	jdff dff_B_wfNoYcMm6_1(.din(w_dff_B_Le1XJwK91_1),.dout(w_dff_B_wfNoYcMm6_1),.clk(gclk));
	jdff dff_B_fI246dkN2_1(.din(w_dff_B_wfNoYcMm6_1),.dout(w_dff_B_fI246dkN2_1),.clk(gclk));
	jdff dff_B_WWxgCCjf9_1(.din(w_dff_B_fI246dkN2_1),.dout(w_dff_B_WWxgCCjf9_1),.clk(gclk));
	jdff dff_B_42RkquX53_1(.din(w_dff_B_WWxgCCjf9_1),.dout(w_dff_B_42RkquX53_1),.clk(gclk));
	jdff dff_B_VMt0Omiv0_1(.din(w_dff_B_42RkquX53_1),.dout(w_dff_B_VMt0Omiv0_1),.clk(gclk));
	jdff dff_B_mzcgcshM3_1(.din(w_dff_B_VMt0Omiv0_1),.dout(w_dff_B_mzcgcshM3_1),.clk(gclk));
	jdff dff_B_QiucouSo8_1(.din(w_dff_B_mzcgcshM3_1),.dout(w_dff_B_QiucouSo8_1),.clk(gclk));
	jdff dff_B_WpLdC2yf9_1(.din(w_dff_B_QiucouSo8_1),.dout(w_dff_B_WpLdC2yf9_1),.clk(gclk));
	jdff dff_B_sOwajJPg5_1(.din(w_dff_B_WpLdC2yf9_1),.dout(w_dff_B_sOwajJPg5_1),.clk(gclk));
	jdff dff_B_LumDwg734_1(.din(w_dff_B_sOwajJPg5_1),.dout(w_dff_B_LumDwg734_1),.clk(gclk));
	jdff dff_B_Kw5aBqFC1_0(.din(n392),.dout(w_dff_B_Kw5aBqFC1_0),.clk(gclk));
	jdff dff_B_DheBu80T7_0(.din(w_dff_B_Kw5aBqFC1_0),.dout(w_dff_B_DheBu80T7_0),.clk(gclk));
	jdff dff_B_8F8oQlE15_0(.din(w_dff_B_DheBu80T7_0),.dout(w_dff_B_8F8oQlE15_0),.clk(gclk));
	jdff dff_B_4zXuBon64_0(.din(w_dff_B_8F8oQlE15_0),.dout(w_dff_B_4zXuBon64_0),.clk(gclk));
	jdff dff_B_5Bc3Cq8z0_0(.din(w_dff_B_4zXuBon64_0),.dout(w_dff_B_5Bc3Cq8z0_0),.clk(gclk));
	jdff dff_B_xU9fo7k41_0(.din(w_dff_B_5Bc3Cq8z0_0),.dout(w_dff_B_xU9fo7k41_0),.clk(gclk));
	jdff dff_B_hW7WgSM70_0(.din(w_dff_B_xU9fo7k41_0),.dout(w_dff_B_hW7WgSM70_0),.clk(gclk));
	jdff dff_B_EtTbpHWJ2_0(.din(w_dff_B_hW7WgSM70_0),.dout(w_dff_B_EtTbpHWJ2_0),.clk(gclk));
	jdff dff_B_3EXQ8fe84_0(.din(w_dff_B_EtTbpHWJ2_0),.dout(w_dff_B_3EXQ8fe84_0),.clk(gclk));
	jdff dff_B_zJp7DNCj6_0(.din(w_dff_B_3EXQ8fe84_0),.dout(w_dff_B_zJp7DNCj6_0),.clk(gclk));
	jdff dff_B_dlWi642E9_0(.din(w_dff_B_zJp7DNCj6_0),.dout(w_dff_B_dlWi642E9_0),.clk(gclk));
	jdff dff_B_9rmQ04lU6_1(.din(n398),.dout(w_dff_B_9rmQ04lU6_1),.clk(gclk));
	jdff dff_A_fuse14T61_2(.dout(w_dff_A_9MUfrTW15_0),.din(w_dff_A_fuse14T61_2),.clk(gclk));
	jdff dff_A_9MUfrTW15_0(.dout(w_dff_A_dKF5pgqF8_0),.din(w_dff_A_9MUfrTW15_0),.clk(gclk));
	jdff dff_A_dKF5pgqF8_0(.dout(w_dff_A_GbxA3kj26_0),.din(w_dff_A_dKF5pgqF8_0),.clk(gclk));
	jdff dff_A_GbxA3kj26_0(.dout(w_dff_A_BHlsa0a93_0),.din(w_dff_A_GbxA3kj26_0),.clk(gclk));
	jdff dff_A_BHlsa0a93_0(.dout(w_dff_A_U0ssrYvD0_0),.din(w_dff_A_BHlsa0a93_0),.clk(gclk));
	jdff dff_A_U0ssrYvD0_0(.dout(w_dff_A_kzR5NI6S3_0),.din(w_dff_A_U0ssrYvD0_0),.clk(gclk));
	jdff dff_A_kzR5NI6S3_0(.dout(G3),.din(w_dff_A_kzR5NI6S3_0),.clk(gclk));
	jdff dff_A_2gaEHoHJ9_2(.dout(w_dff_A_hVjHpR7I4_0),.din(w_dff_A_2gaEHoHJ9_2),.clk(gclk));
	jdff dff_A_hVjHpR7I4_0(.dout(w_dff_A_UvkMzsCG6_0),.din(w_dff_A_hVjHpR7I4_0),.clk(gclk));
	jdff dff_A_UvkMzsCG6_0(.dout(w_dff_A_DZ5w9hss0_0),.din(w_dff_A_UvkMzsCG6_0),.clk(gclk));
	jdff dff_A_DZ5w9hss0_0(.dout(w_dff_A_YbYzecui7_0),.din(w_dff_A_DZ5w9hss0_0),.clk(gclk));
	jdff dff_A_YbYzecui7_0(.dout(w_dff_A_aC57sAI99_0),.din(w_dff_A_YbYzecui7_0),.clk(gclk));
	jdff dff_A_aC57sAI99_0(.dout(w_dff_A_dYt9jr318_0),.din(w_dff_A_aC57sAI99_0),.clk(gclk));
	jdff dff_A_dYt9jr318_0(.dout(G6),.din(w_dff_A_dYt9jr318_0),.clk(gclk));
	jdff dff_A_P8R2qX6l0_2(.dout(w_dff_A_sBFpdlpI2_0),.din(w_dff_A_P8R2qX6l0_2),.clk(gclk));
	jdff dff_A_sBFpdlpI2_0(.dout(w_dff_A_wZeA5PC48_0),.din(w_dff_A_sBFpdlpI2_0),.clk(gclk));
	jdff dff_A_wZeA5PC48_0(.dout(w_dff_A_LUesZXVF2_0),.din(w_dff_A_wZeA5PC48_0),.clk(gclk));
	jdff dff_A_LUesZXVF2_0(.dout(w_dff_A_EvlSyBMq0_0),.din(w_dff_A_LUesZXVF2_0),.clk(gclk));
	jdff dff_A_EvlSyBMq0_0(.dout(w_dff_A_QM9OZKLr8_0),.din(w_dff_A_EvlSyBMq0_0),.clk(gclk));
	jdff dff_A_QM9OZKLr8_0(.dout(w_dff_A_F7gG8OG23_0),.din(w_dff_A_QM9OZKLr8_0),.clk(gclk));
	jdff dff_A_F7gG8OG23_0(.dout(G9),.din(w_dff_A_F7gG8OG23_0),.clk(gclk));
	jdff dff_A_Iv1cyd7k5_2(.dout(w_dff_A_VlePD7MI0_0),.din(w_dff_A_Iv1cyd7k5_2),.clk(gclk));
	jdff dff_A_VlePD7MI0_0(.dout(w_dff_A_HYZxUNkd7_0),.din(w_dff_A_VlePD7MI0_0),.clk(gclk));
	jdff dff_A_HYZxUNkd7_0(.dout(w_dff_A_iLKjr7Zx3_0),.din(w_dff_A_HYZxUNkd7_0),.clk(gclk));
	jdff dff_A_iLKjr7Zx3_0(.dout(w_dff_A_y4IhiKIr6_0),.din(w_dff_A_iLKjr7Zx3_0),.clk(gclk));
	jdff dff_A_y4IhiKIr6_0(.dout(w_dff_A_blTbcDJf5_0),.din(w_dff_A_y4IhiKIr6_0),.clk(gclk));
	jdff dff_A_blTbcDJf5_0(.dout(w_dff_A_0lztIxwK2_0),.din(w_dff_A_blTbcDJf5_0),.clk(gclk));
	jdff dff_A_0lztIxwK2_0(.dout(G12),.din(w_dff_A_0lztIxwK2_0),.clk(gclk));
	jdff dff_A_8PLLfsFp3_2(.dout(w_dff_A_KbdHPIkd9_0),.din(w_dff_A_8PLLfsFp3_2),.clk(gclk));
	jdff dff_A_KbdHPIkd9_0(.dout(w_dff_A_YAy6vcNW3_0),.din(w_dff_A_KbdHPIkd9_0),.clk(gclk));
	jdff dff_A_YAy6vcNW3_0(.dout(w_dff_A_MfXzEgtD1_0),.din(w_dff_A_YAy6vcNW3_0),.clk(gclk));
	jdff dff_A_MfXzEgtD1_0(.dout(w_dff_A_7enoBNa54_0),.din(w_dff_A_MfXzEgtD1_0),.clk(gclk));
	jdff dff_A_7enoBNa54_0(.dout(w_dff_A_9mzdA1ar1_0),.din(w_dff_A_7enoBNa54_0),.clk(gclk));
	jdff dff_A_9mzdA1ar1_0(.dout(w_dff_A_Yhxa399s3_0),.din(w_dff_A_9mzdA1ar1_0),.clk(gclk));
	jdff dff_A_Yhxa399s3_0(.dout(G30),.din(w_dff_A_Yhxa399s3_0),.clk(gclk));
	jdff dff_A_uKogXNzU7_2(.dout(w_dff_A_GmLMgmTL9_0),.din(w_dff_A_uKogXNzU7_2),.clk(gclk));
	jdff dff_A_GmLMgmTL9_0(.dout(w_dff_A_LgLqwJ3d3_0),.din(w_dff_A_GmLMgmTL9_0),.clk(gclk));
	jdff dff_A_LgLqwJ3d3_0(.dout(w_dff_A_19AiRCiG9_0),.din(w_dff_A_LgLqwJ3d3_0),.clk(gclk));
	jdff dff_A_19AiRCiG9_0(.dout(w_dff_A_x3Y4IHRn3_0),.din(w_dff_A_19AiRCiG9_0),.clk(gclk));
	jdff dff_A_x3Y4IHRn3_0(.dout(w_dff_A_nN8uEuiz3_0),.din(w_dff_A_x3Y4IHRn3_0),.clk(gclk));
	jdff dff_A_nN8uEuiz3_0(.dout(w_dff_A_iijZsxpL1_0),.din(w_dff_A_nN8uEuiz3_0),.clk(gclk));
	jdff dff_A_iijZsxpL1_0(.dout(G45),.din(w_dff_A_iijZsxpL1_0),.clk(gclk));
	jdff dff_A_b9MQohhs2_2(.dout(w_dff_A_hzsudhFQ2_0),.din(w_dff_A_b9MQohhs2_2),.clk(gclk));
	jdff dff_A_hzsudhFQ2_0(.dout(w_dff_A_44GvxLGf9_0),.din(w_dff_A_hzsudhFQ2_0),.clk(gclk));
	jdff dff_A_44GvxLGf9_0(.dout(w_dff_A_lK6scgeg4_0),.din(w_dff_A_44GvxLGf9_0),.clk(gclk));
	jdff dff_A_lK6scgeg4_0(.dout(w_dff_A_7U93AYXO2_0),.din(w_dff_A_lK6scgeg4_0),.clk(gclk));
	jdff dff_A_7U93AYXO2_0(.dout(w_dff_A_1SbbXg5O1_0),.din(w_dff_A_7U93AYXO2_0),.clk(gclk));
	jdff dff_A_1SbbXg5O1_0(.dout(w_dff_A_TTlaiYnO7_0),.din(w_dff_A_1SbbXg5O1_0),.clk(gclk));
	jdff dff_A_TTlaiYnO7_0(.dout(G48),.din(w_dff_A_TTlaiYnO7_0),.clk(gclk));
	jdff dff_A_30rl8IDl4_2(.dout(w_dff_A_dN4c5WwJ6_0),.din(w_dff_A_30rl8IDl4_2),.clk(gclk));
	jdff dff_A_dN4c5WwJ6_0(.dout(w_dff_A_2LSmskpI0_0),.din(w_dff_A_dN4c5WwJ6_0),.clk(gclk));
	jdff dff_A_2LSmskpI0_0(.dout(w_dff_A_TtEBxQGL1_0),.din(w_dff_A_2LSmskpI0_0),.clk(gclk));
	jdff dff_A_TtEBxQGL1_0(.dout(w_dff_A_Z6NaGQ060_0),.din(w_dff_A_TtEBxQGL1_0),.clk(gclk));
	jdff dff_A_Z6NaGQ060_0(.dout(w_dff_A_NxsNfYrg8_0),.din(w_dff_A_Z6NaGQ060_0),.clk(gclk));
	jdff dff_A_NxsNfYrg8_0(.dout(w_dff_A_AspwU5ia6_0),.din(w_dff_A_NxsNfYrg8_0),.clk(gclk));
	jdff dff_A_AspwU5ia6_0(.dout(G15),.din(w_dff_A_AspwU5ia6_0),.clk(gclk));
	jdff dff_A_cPpb56RY3_2(.dout(w_dff_A_K82LTB7q9_0),.din(w_dff_A_cPpb56RY3_2),.clk(gclk));
	jdff dff_A_K82LTB7q9_0(.dout(w_dff_A_rCdHRB3a0_0),.din(w_dff_A_K82LTB7q9_0),.clk(gclk));
	jdff dff_A_rCdHRB3a0_0(.dout(w_dff_A_iem2k9aV8_0),.din(w_dff_A_rCdHRB3a0_0),.clk(gclk));
	jdff dff_A_iem2k9aV8_0(.dout(w_dff_A_nNwrKDRC4_0),.din(w_dff_A_iem2k9aV8_0),.clk(gclk));
	jdff dff_A_nNwrKDRC4_0(.dout(w_dff_A_cFG1oKhb9_0),.din(w_dff_A_nNwrKDRC4_0),.clk(gclk));
	jdff dff_A_cFG1oKhb9_0(.dout(w_dff_A_MTLeesBI4_0),.din(w_dff_A_cFG1oKhb9_0),.clk(gclk));
	jdff dff_A_MTLeesBI4_0(.dout(G18),.din(w_dff_A_MTLeesBI4_0),.clk(gclk));
	jdff dff_A_vWFS0OZ25_2(.dout(w_dff_A_LodlJLby4_0),.din(w_dff_A_vWFS0OZ25_2),.clk(gclk));
	jdff dff_A_LodlJLby4_0(.dout(w_dff_A_2EtwuHP34_0),.din(w_dff_A_LodlJLby4_0),.clk(gclk));
	jdff dff_A_2EtwuHP34_0(.dout(w_dff_A_EVhoD0Uo5_0),.din(w_dff_A_2EtwuHP34_0),.clk(gclk));
	jdff dff_A_EVhoD0Uo5_0(.dout(w_dff_A_JebwlGQM1_0),.din(w_dff_A_EVhoD0Uo5_0),.clk(gclk));
	jdff dff_A_JebwlGQM1_0(.dout(w_dff_A_lhgDSYtn2_0),.din(w_dff_A_JebwlGQM1_0),.clk(gclk));
	jdff dff_A_lhgDSYtn2_0(.dout(w_dff_A_mhT7ScXv4_0),.din(w_dff_A_lhgDSYtn2_0),.clk(gclk));
	jdff dff_A_mhT7ScXv4_0(.dout(G21),.din(w_dff_A_mhT7ScXv4_0),.clk(gclk));
	jdff dff_A_fXWr2Uu04_2(.dout(w_dff_A_Cf4oJ98q5_0),.din(w_dff_A_fXWr2Uu04_2),.clk(gclk));
	jdff dff_A_Cf4oJ98q5_0(.dout(w_dff_A_6q7OG8m15_0),.din(w_dff_A_Cf4oJ98q5_0),.clk(gclk));
	jdff dff_A_6q7OG8m15_0(.dout(w_dff_A_xH1dtE183_0),.din(w_dff_A_6q7OG8m15_0),.clk(gclk));
	jdff dff_A_xH1dtE183_0(.dout(w_dff_A_C0HrwjsY5_0),.din(w_dff_A_xH1dtE183_0),.clk(gclk));
	jdff dff_A_C0HrwjsY5_0(.dout(w_dff_A_KZMoV3PV7_0),.din(w_dff_A_C0HrwjsY5_0),.clk(gclk));
	jdff dff_A_KZMoV3PV7_0(.dout(w_dff_A_H4dd3DQS0_0),.din(w_dff_A_KZMoV3PV7_0),.clk(gclk));
	jdff dff_A_H4dd3DQS0_0(.dout(G24),.din(w_dff_A_H4dd3DQS0_0),.clk(gclk));
	jdff dff_A_E9NAXxXK0_2(.dout(w_dff_A_03NK2lHB4_0),.din(w_dff_A_E9NAXxXK0_2),.clk(gclk));
	jdff dff_A_03NK2lHB4_0(.dout(w_dff_A_k7YLEW7A6_0),.din(w_dff_A_03NK2lHB4_0),.clk(gclk));
	jdff dff_A_k7YLEW7A6_0(.dout(w_dff_A_Zy92Q7jn2_0),.din(w_dff_A_k7YLEW7A6_0),.clk(gclk));
	jdff dff_A_Zy92Q7jn2_0(.dout(w_dff_A_Q7HRDvYK1_0),.din(w_dff_A_Zy92Q7jn2_0),.clk(gclk));
	jdff dff_A_Q7HRDvYK1_0(.dout(w_dff_A_qel2dIz33_0),.din(w_dff_A_Q7HRDvYK1_0),.clk(gclk));
	jdff dff_A_qel2dIz33_0(.dout(w_dff_A_ITyeNT9e2_0),.din(w_dff_A_qel2dIz33_0),.clk(gclk));
	jdff dff_A_ITyeNT9e2_0(.dout(G27),.din(w_dff_A_ITyeNT9e2_0),.clk(gclk));
	jdff dff_A_jF9YHq5j2_2(.dout(w_dff_A_iwZpseBI0_0),.din(w_dff_A_jF9YHq5j2_2),.clk(gclk));
	jdff dff_A_iwZpseBI0_0(.dout(w_dff_A_RNmSBhdL7_0),.din(w_dff_A_iwZpseBI0_0),.clk(gclk));
	jdff dff_A_RNmSBhdL7_0(.dout(w_dff_A_J57e2zIl8_0),.din(w_dff_A_RNmSBhdL7_0),.clk(gclk));
	jdff dff_A_J57e2zIl8_0(.dout(w_dff_A_dPAcUBw47_0),.din(w_dff_A_J57e2zIl8_0),.clk(gclk));
	jdff dff_A_dPAcUBw47_0(.dout(w_dff_A_mE8iwXT05_0),.din(w_dff_A_dPAcUBw47_0),.clk(gclk));
	jdff dff_A_mE8iwXT05_0(.dout(w_dff_A_Bhg3h0bn3_0),.din(w_dff_A_mE8iwXT05_0),.clk(gclk));
	jdff dff_A_Bhg3h0bn3_0(.dout(G33),.din(w_dff_A_Bhg3h0bn3_0),.clk(gclk));
	jdff dff_A_CObwD37Y6_2(.dout(w_dff_A_NkBrZtAD0_0),.din(w_dff_A_CObwD37Y6_2),.clk(gclk));
	jdff dff_A_NkBrZtAD0_0(.dout(w_dff_A_ccYvgVl96_0),.din(w_dff_A_NkBrZtAD0_0),.clk(gclk));
	jdff dff_A_ccYvgVl96_0(.dout(w_dff_A_ZmxJS0DB0_0),.din(w_dff_A_ccYvgVl96_0),.clk(gclk));
	jdff dff_A_ZmxJS0DB0_0(.dout(w_dff_A_uGB2f2br7_0),.din(w_dff_A_ZmxJS0DB0_0),.clk(gclk));
	jdff dff_A_uGB2f2br7_0(.dout(w_dff_A_gQJYD8Bv5_0),.din(w_dff_A_uGB2f2br7_0),.clk(gclk));
	jdff dff_A_gQJYD8Bv5_0(.dout(w_dff_A_q3v43UeU5_0),.din(w_dff_A_gQJYD8Bv5_0),.clk(gclk));
	jdff dff_A_q3v43UeU5_0(.dout(G36),.din(w_dff_A_q3v43UeU5_0),.clk(gclk));
	jdff dff_A_9pyUhmRS8_2(.dout(w_dff_A_bEYpzb9h4_0),.din(w_dff_A_9pyUhmRS8_2),.clk(gclk));
	jdff dff_A_bEYpzb9h4_0(.dout(w_dff_A_ZP19CT7t9_0),.din(w_dff_A_bEYpzb9h4_0),.clk(gclk));
	jdff dff_A_ZP19CT7t9_0(.dout(w_dff_A_ihkGyJKt2_0),.din(w_dff_A_ZP19CT7t9_0),.clk(gclk));
	jdff dff_A_ihkGyJKt2_0(.dout(w_dff_A_yBM0Ovkd0_0),.din(w_dff_A_ihkGyJKt2_0),.clk(gclk));
	jdff dff_A_yBM0Ovkd0_0(.dout(w_dff_A_kwbLCVc64_0),.din(w_dff_A_yBM0Ovkd0_0),.clk(gclk));
	jdff dff_A_kwbLCVc64_0(.dout(w_dff_A_m0SgaP3O1_0),.din(w_dff_A_kwbLCVc64_0),.clk(gclk));
	jdff dff_A_m0SgaP3O1_0(.dout(G39),.din(w_dff_A_m0SgaP3O1_0),.clk(gclk));
	jdff dff_A_bMjqVEuP0_2(.dout(w_dff_A_eBQQkB3P1_0),.din(w_dff_A_bMjqVEuP0_2),.clk(gclk));
	jdff dff_A_eBQQkB3P1_0(.dout(w_dff_A_E0SZC2Xx1_0),.din(w_dff_A_eBQQkB3P1_0),.clk(gclk));
	jdff dff_A_E0SZC2Xx1_0(.dout(w_dff_A_LEo8QUvu2_0),.din(w_dff_A_E0SZC2Xx1_0),.clk(gclk));
	jdff dff_A_LEo8QUvu2_0(.dout(w_dff_A_pKqBkQWa2_0),.din(w_dff_A_LEo8QUvu2_0),.clk(gclk));
	jdff dff_A_pKqBkQWa2_0(.dout(w_dff_A_XygrURur2_0),.din(w_dff_A_pKqBkQWa2_0),.clk(gclk));
	jdff dff_A_XygrURur2_0(.dout(w_dff_A_9BAqzG8j3_0),.din(w_dff_A_XygrURur2_0),.clk(gclk));
	jdff dff_A_9BAqzG8j3_0(.dout(G42),.din(w_dff_A_9BAqzG8j3_0),.clk(gclk));
	jdff dff_A_T9z38KbT5_2(.dout(G75),.din(w_dff_A_T9z38KbT5_2),.clk(gclk));
	jdff dff_A_wZn0xXb02_2(.dout(G69),.din(w_dff_A_wZn0xXb02_2),.clk(gclk));
	jdff dff_A_EFbnONC66_2(.dout(w_dff_A_q1bJJ9db2_0),.din(w_dff_A_EFbnONC66_2),.clk(gclk));
	jdff dff_A_q1bJJ9db2_0(.dout(G72),.din(w_dff_A_q1bJJ9db2_0),.clk(gclk));
endmodule

