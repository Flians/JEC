/*

c5315:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jdff: 6080
	jand: 606
	jor: 486

Summary:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jdff: 6080
	jand: 606
	jor: 486
*/

module c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[1:0] w_G1_2;
	wire[2:0] w_G4_0;
	wire[1:0] w_G11_0;
	wire[1:0] w_G14_0;
	wire[1:0] w_G17_0;
	wire[1:0] w_G20_0;
	wire[1:0] w_G37_0;
	wire[1:0] w_G40_0;
	wire[1:0] w_G43_0;
	wire[1:0] w_G46_0;
	wire[1:0] w_G49_0;
	wire[2:0] w_G54_0;
	wire[1:0] w_G61_0;
	wire[1:0] w_G64_0;
	wire[1:0] w_G67_0;
	wire[1:0] w_G70_0;
	wire[1:0] w_G73_0;
	wire[1:0] w_G76_0;
	wire[1:0] w_G91_0;
	wire[1:0] w_G100_0;
	wire[1:0] w_G103_0;
	wire[1:0] w_G106_0;
	wire[1:0] w_G109_0;
	wire[1:0] w_G123_0;
	wire[2:0] w_G137_0;
	wire[2:0] w_G137_1;
	wire[2:0] w_G137_2;
	wire[2:0] w_G137_3;
	wire[2:0] w_G137_4;
	wire[2:0] w_G137_5;
	wire[2:0] w_G137_6;
	wire[2:0] w_G137_7;
	wire[2:0] w_G137_8;
	wire[1:0] w_G137_9;
	wire[2:0] w_G141_0;
	wire[2:0] w_G141_1;
	wire[2:0] w_G141_2;
	wire[1:0] w_G146_0;
	wire[1:0] w_G149_0;
	wire[1:0] w_G152_0;
	wire[1:0] w_G155_0;
	wire[1:0] w_G158_0;
	wire[1:0] w_G161_0;
	wire[1:0] w_G164_0;
	wire[1:0] w_G167_0;
	wire[1:0] w_G170_0;
	wire[1:0] w_G173_0;
	wire[1:0] w_G182_0;
	wire[1:0] w_G185_0;
	wire[1:0] w_G188_0;
	wire[1:0] w_G191_0;
	wire[1:0] w_G194_0;
	wire[1:0] w_G197_0;
	wire[1:0] w_G200_0;
	wire[1:0] w_G203_0;
	wire[2:0] w_G206_0;
	wire[2:0] w_G206_1;
	wire[2:0] w_G210_0;
	wire[2:0] w_G210_1;
	wire[1:0] w_G210_2;
	wire[2:0] w_G218_0;
	wire[2:0] w_G218_1;
	wire[1:0] w_G218_2;
	wire[2:0] w_G226_0;
	wire[2:0] w_G226_1;
	wire[1:0] w_G226_2;
	wire[2:0] w_G234_0;
	wire[2:0] w_G234_1;
	wire[1:0] w_G234_2;
	wire[2:0] w_G242_0;
	wire[1:0] w_G242_1;
	wire[1:0] w_G245_0;
	wire[2:0] w_G248_0;
	wire[2:0] w_G248_1;
	wire[2:0] w_G248_2;
	wire[2:0] w_G248_3;
	wire[2:0] w_G248_4;
	wire[2:0] w_G248_5;
	wire[2:0] w_G251_0;
	wire[2:0] w_G251_1;
	wire[2:0] w_G251_2;
	wire[2:0] w_G251_3;
	wire[2:0] w_G251_4;
	wire[1:0] w_G251_5;
	wire[2:0] w_G254_0;
	wire[1:0] w_G254_1;
	wire[2:0] w_G257_0;
	wire[2:0] w_G257_1;
	wire[1:0] w_G257_2;
	wire[2:0] w_G265_0;
	wire[2:0] w_G265_1;
	wire[2:0] w_G273_0;
	wire[2:0] w_G273_1;
	wire[1:0] w_G273_2;
	wire[2:0] w_G281_0;
	wire[2:0] w_G281_1;
	wire[1:0] w_G281_2;
	wire[1:0] w_G289_0;
	wire[2:0] w_G293_0;
	wire[2:0] w_G299_0;
	wire[2:0] w_G302_0;
	wire[2:0] w_G308_0;
	wire[2:0] w_G308_1;
	wire[2:0] w_G316_0;
	wire[1:0] w_G316_1;
	wire[2:0] w_G324_0;
	wire[2:0] w_G324_1;
	wire[1:0] w_G331_0;
	wire[2:0] w_G332_0;
	wire[2:0] w_G332_1;
	wire[2:0] w_G332_2;
	wire[2:0] w_G332_3;
	wire[2:0] w_G335_0;
	wire[1:0] w_G338_0;
	wire[2:0] w_G341_0;
	wire[2:0] w_G341_1;
	wire[2:0] w_G341_2;
	wire[1:0] w_G348_0;
	wire[2:0] w_G351_0;
	wire[2:0] w_G351_1;
	wire[2:0] w_G351_2;
	wire[1:0] w_G358_0;
	wire[2:0] w_G361_0;
	wire[1:0] w_G361_1;
	wire[1:0] w_G366_0;
	wire[1:0] w_G369_0;
	wire[2:0] w_G374_0;
	wire[2:0] w_G374_1;
	wire[2:0] w_G389_0;
	wire[2:0] w_G389_1;
	wire[2:0] w_G400_0;
	wire[2:0] w_G400_1;
	wire[2:0] w_G411_0;
	wire[2:0] w_G411_1;
	wire[1:0] w_G411_2;
	wire[2:0] w_G422_0;
	wire[1:0] w_G422_1;
	wire[2:0] w_G435_0;
	wire[2:0] w_G435_1;
	wire[2:0] w_G446_0;
	wire[2:0] w_G446_1;
	wire[2:0] w_G457_0;
	wire[2:0] w_G457_1;
	wire[2:0] w_G468_0;
	wire[2:0] w_G468_1;
	wire[2:0] w_G479_0;
	wire[2:0] w_G490_0;
	wire[1:0] w_G490_1;
	wire[2:0] w_G503_0;
	wire[2:0] w_G503_1;
	wire[1:0] w_G503_2;
	wire[2:0] w_G514_0;
	wire[2:0] w_G514_1;
	wire[1:0] w_G514_2;
	wire[2:0] w_G523_0;
	wire[2:0] w_G523_1;
	wire[2:0] w_G534_0;
	wire[2:0] w_G534_1;
	wire[1:0] w_G534_2;
	wire[2:0] w_G545_0;
	wire[2:0] w_G549_0;
	wire[1:0] w_G552_0;
	wire[1:0] w_G559_0;
	wire[1:0] w_G562_0;
	wire[2:0] w_G1497_0;
	wire[2:0] w_G1689_0;
	wire[2:0] w_G1689_1;
	wire[2:0] w_G1689_2;
	wire[2:0] w_G1689_3;
	wire[2:0] w_G1689_4;
	wire[1:0] w_G1689_5;
	wire[2:0] w_G1690_0;
	wire[1:0] w_G1690_1;
	wire[2:0] w_G1691_0;
	wire[2:0] w_G1691_1;
	wire[2:0] w_G1691_2;
	wire[2:0] w_G1691_3;
	wire[2:0] w_G1691_4;
	wire[1:0] w_G1691_5;
	wire[2:0] w_G1694_0;
	wire[1:0] w_G1694_1;
	wire[2:0] w_G2174_0;
	wire[2:0] w_G2358_0;
	wire[2:0] w_G2358_1;
	wire[2:0] w_G2358_2;
	wire[1:0] w_G3173_0;
	wire[2:0] w_G3546_0;
	wire[2:0] w_G3546_1;
	wire[2:0] w_G3546_2;
	wire[2:0] w_G3546_3;
	wire[2:0] w_G3546_4;
	wire[1:0] w_G3546_5;
	wire[2:0] w_G3548_0;
	wire[2:0] w_G3548_1;
	wire[2:0] w_G3548_2;
	wire[2:0] w_G3548_3;
	wire[2:0] w_G3548_4;
	wire[1:0] w_G3552_0;
	wire[1:0] w_G3717_0;
	wire[2:0] w_G3724_0;
	wire[2:0] w_G4087_0;
	wire[2:0] w_G4087_1;
	wire[2:0] w_G4087_2;
	wire[2:0] w_G4087_3;
	wire[2:0] w_G4087_4;
	wire[2:0] w_G4088_0;
	wire[2:0] w_G4088_1;
	wire[2:0] w_G4088_2;
	wire[2:0] w_G4088_3;
	wire[2:0] w_G4088_4;
	wire[2:0] w_G4088_5;
	wire[2:0] w_G4088_6;
	wire[2:0] w_G4088_7;
	wire[2:0] w_G4088_8;
	wire[2:0] w_G4088_9;
	wire[2:0] w_G4089_0;
	wire[2:0] w_G4089_1;
	wire[2:0] w_G4089_2;
	wire[2:0] w_G4089_3;
	wire[2:0] w_G4089_4;
	wire[2:0] w_G4089_5;
	wire[2:0] w_G4089_6;
	wire[2:0] w_G4089_7;
	wire[2:0] w_G4089_8;
	wire[2:0] w_G4089_9;
	wire[2:0] w_G4090_0;
	wire[2:0] w_G4090_1;
	wire[2:0] w_G4090_2;
	wire[2:0] w_G4090_3;
	wire[2:0] w_G4090_4;
	wire[2:0] w_G4091_0;
	wire[2:0] w_G4091_1;
	wire[2:0] w_G4091_2;
	wire[2:0] w_G4091_3;
	wire[2:0] w_G4091_4;
	wire[2:0] w_G4091_5;
	wire[1:0] w_G4091_6;
	wire[2:0] w_G4092_0;
	wire[2:0] w_G4092_1;
	wire[2:0] w_G4092_2;
	wire[2:0] w_G4092_3;
	wire[2:0] w_G4092_4;
	wire[2:0] w_G4092_5;
	wire[2:0] w_G4092_6;
	wire[2:0] w_G4092_7;
	wire[2:0] w_G4092_8;
	wire[2:0] w_G4092_9;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire[2:0] w_G809_0;
	wire[2:0] w_G809_1;
	wire[2:0] w_G809_2;
	wire[1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G623_0;
	wire G623_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G998_0;
	wire G998_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G865_0;
	wire G865_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire[1:0] w_n316_0;
	wire[1:0] w_n318_0;
	wire[2:0] w_n326_0;
	wire[2:0] w_n326_1;
	wire[1:0] w_n326_2;
	wire[1:0] w_n333_0;
	wire[1:0] w_n336_0;
	wire[1:0] w_n361_0;
	wire[1:0] w_n365_0;
	wire[2:0] w_n366_0;
	wire[2:0] w_n366_1;
	wire[2:0] w_n369_0;
	wire[2:0] w_n369_1;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[2:0] w_n374_0;
	wire[1:0] w_n374_1;
	wire[2:0] w_n375_0;
	wire[2:0] w_n375_1;
	wire[2:0] w_n375_2;
	wire[2:0] w_n375_3;
	wire[2:0] w_n375_4;
	wire[2:0] w_n377_0;
	wire[1:0] w_n377_1;
	wire[2:0] w_n378_0;
	wire[2:0] w_n378_1;
	wire[2:0] w_n378_2;
	wire[2:0] w_n378_3;
	wire[2:0] w_n378_4;
	wire[1:0] w_n386_0;
	wire[2:0] w_n387_0;
	wire[1:0] w_n387_1;
	wire[2:0] w_n389_0;
	wire[1:0] w_n389_1;
	wire[1:0] w_n397_0;
	wire[1:0] w_n401_0;
	wire[2:0] w_n402_0;
	wire[2:0] w_n406_0;
	wire[2:0] w_n406_1;
	wire[2:0] w_n406_2;
	wire[2:0] w_n406_3;
	wire[2:0] w_n406_4;
	wire[1:0] w_n406_5;
	wire[2:0] w_n408_0;
	wire[2:0] w_n408_1;
	wire[2:0] w_n408_2;
	wire[2:0] w_n408_3;
	wire[2:0] w_n408_4;
	wire[2:0] w_n408_5;
	wire[2:0] w_n412_0;
	wire[1:0] w_n414_0;
	wire[1:0] w_n415_0;
	wire[2:0] w_n423_0;
	wire[2:0] w_n425_0;
	wire[2:0] w_n428_0;
	wire[1:0] w_n428_1;
	wire[1:0] w_n429_0;
	wire[2:0] w_n433_0;
	wire[2:0] w_n435_0;
	wire[2:0] w_n435_1;
	wire[1:0] w_n435_2;
	wire[1:0] w_n437_0;
	wire[1:0] w_n445_0;
	wire[2:0] w_n449_0;
	wire[2:0] w_n449_1;
	wire[2:0] w_n451_0;
	wire[1:0] w_n459_0;
	wire[2:0] w_n460_0;
	wire[2:0] w_n460_1;
	wire[2:0] w_n462_0;
	wire[1:0] w_n470_0;
	wire[2:0] w_n471_0;
	wire[2:0] w_n471_1;
	wire[2:0] w_n473_0;
	wire[1:0] w_n473_1;
	wire[1:0] w_n481_0;
	wire[2:0] w_n483_0;
	wire[2:0] w_n483_1;
	wire[1:0] w_n483_2;
	wire[2:0] w_n485_0;
	wire[1:0] w_n485_1;
	wire[1:0] w_n493_0;
	wire[2:0] w_n494_0;
	wire[2:0] w_n494_1;
	wire[2:0] w_n496_0;
	wire[1:0] w_n496_1;
	wire[1:0] w_n504_0;
	wire[2:0] w_n507_0;
	wire[2:0] w_n507_1;
	wire[2:0] w_n509_0;
	wire[1:0] w_n517_0;
	wire[2:0] w_n518_0;
	wire[2:0] w_n518_1;
	wire[2:0] w_n520_0;
	wire[1:0] w_n528_0;
	wire[2:0] w_n530_0;
	wire[2:0] w_n530_1;
	wire[2:0] w_n532_0;
	wire[1:0] w_n532_1;
	wire[1:0] w_n540_0;
	wire[1:0] w_n543_0;
	wire[2:0] w_n551_0;
	wire[2:0] w_n556_0;
	wire[2:0] w_n556_1;
	wire[2:0] w_n556_2;
	wire[2:0] w_n556_3;
	wire[2:0] w_n556_4;
	wire[2:0] w_n556_5;
	wire[2:0] w_n556_6;
	wire[2:0] w_n556_7;
	wire[1:0] w_n556_8;
	wire[1:0] w_n557_0;
	wire[1:0] w_n559_0;
	wire[2:0] w_n560_0;
	wire[2:0] w_n561_0;
	wire[1:0] w_n561_1;
	wire[1:0] w_n562_0;
	wire[1:0] w_n564_0;
	wire[2:0] w_n565_0;
	wire[2:0] w_n566_0;
	wire[2:0] w_n567_0;
	wire[1:0] w_n569_0;
	wire[1:0] w_n571_0;
	wire[2:0] w_n572_0;
	wire[2:0] w_n573_0;
	wire[2:0] w_n574_0;
	wire[2:0] w_n578_0;
	wire[1:0] w_n578_1;
	wire[2:0] w_n579_0;
	wire[1:0] w_n579_1;
	wire[1:0] w_n581_0;
	wire[2:0] w_n586_0;
	wire[1:0] w_n586_1;
	wire[1:0] w_n587_0;
	wire[2:0] w_n588_0;
	wire[1:0] w_n588_1;
	wire[2:0] w_n591_0;
	wire[1:0] w_n591_1;
	wire[2:0] w_n592_0;
	wire[2:0] w_n596_0;
	wire[1:0] w_n596_1;
	wire[2:0] w_n597_0;
	wire[2:0] w_n601_0;
	wire[1:0] w_n601_1;
	wire[2:0] w_n602_0;
	wire[1:0] w_n603_0;
	wire[2:0] w_n607_0;
	wire[1:0] w_n607_1;
	wire[2:0] w_n608_0;
	wire[2:0] w_n609_0;
	wire[2:0] w_n611_0;
	wire[2:0] w_n613_0;
	wire[2:0] w_n613_1;
	wire[2:0] w_n613_2;
	wire[2:0] w_n613_3;
	wire[2:0] w_n613_4;
	wire[2:0] w_n613_5;
	wire[2:0] w_n617_0;
	wire[1:0] w_n617_1;
	wire[2:0] w_n618_0;
	wire[2:0] w_n619_0;
	wire[2:0] w_n619_1;
	wire[2:0] w_n620_0;
	wire[1:0] w_n620_1;
	wire[1:0] w_n621_0;
	wire[1:0] w_n623_0;
	wire[2:0] w_n624_0;
	wire[1:0] w_n625_0;
	wire[2:0] w_n627_0;
	wire[1:0] w_n627_1;
	wire[2:0] w_n628_0;
	wire[1:0] w_n631_0;
	wire[1:0] w_n632_0;
	wire[2:0] w_n635_0;
	wire[1:0] w_n635_1;
	wire[2:0] w_n636_0;
	wire[2:0] w_n637_0;
	wire[1:0] w_n638_0;
	wire[2:0] w_n639_0;
	wire[1:0] w_n640_0;
	wire[2:0] w_n641_0;
	wire[2:0] w_n641_1;
	wire[2:0] w_n644_0;
	wire[2:0] w_n648_0;
	wire[1:0] w_n648_1;
	wire[1:0] w_n649_0;
	wire[1:0] w_n650_0;
	wire[2:0] w_n653_0;
	wire[2:0] w_n654_0;
	wire[2:0] w_n654_1;
	wire[2:0] w_n654_2;
	wire[2:0] w_n658_0;
	wire[1:0] w_n658_1;
	wire[1:0] w_n659_0;
	wire[2:0] w_n660_0;
	wire[1:0] w_n660_1;
	wire[1:0] w_n661_0;
	wire[1:0] w_n670_0;
	wire[1:0] w_n680_0;
	wire[2:0] w_n682_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n685_0;
	wire[1:0] w_n686_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n692_0;
	wire[2:0] w_n694_0;
	wire[2:0] w_n695_0;
	wire[2:0] w_n699_0;
	wire[1:0] w_n701_0;
	wire[2:0] w_n703_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n709_0;
	wire[1:0] w_n710_0;
	wire[1:0] w_n711_0;
	wire[2:0] w_n713_0;
	wire[2:0] w_n715_0;
	wire[1:0] w_n717_0;
	wire[1:0] w_n719_0;
	wire[1:0] w_n720_0;
	wire[1:0] w_n721_0;
	wire[1:0] w_n722_0;
	wire[2:0] w_n725_0;
	wire[1:0] w_n726_0;
	wire[1:0] w_n728_0;
	wire[2:0] w_n733_0;
	wire[2:0] w_n735_0;
	wire[2:0] w_n737_0;
	wire[1:0] w_n737_1;
	wire[1:0] w_n738_0;
	wire[2:0] w_n742_0;
	wire[1:0] w_n745_0;
	wire[2:0] w_n746_0;
	wire[1:0] w_n747_0;
	wire[2:0] w_n749_0;
	wire[2:0] w_n749_1;
	wire[2:0] w_n749_2;
	wire[2:0] w_n749_3;
	wire[2:0] w_n749_4;
	wire[2:0] w_n749_5;
	wire[2:0] w_n749_6;
	wire[2:0] w_n749_7;
	wire[2:0] w_n749_8;
	wire[2:0] w_n749_9;
	wire[2:0] w_n749_10;
	wire[2:0] w_n749_11;
	wire[2:0] w_n749_12;
	wire[1:0] w_n749_13;
	wire[2:0] w_n750_0;
	wire[2:0] w_n750_1;
	wire[2:0] w_n750_2;
	wire[2:0] w_n750_3;
	wire[2:0] w_n750_4;
	wire[2:0] w_n750_5;
	wire[2:0] w_n750_6;
	wire[2:0] w_n750_7;
	wire[2:0] w_n750_8;
	wire[2:0] w_n753_0;
	wire[1:0] w_n753_1;
	wire[1:0] w_n755_0;
	wire[2:0] w_n763_0;
	wire[1:0] w_n767_0;
	wire[1:0] w_n779_0;
	wire[2:0] w_n786_0;
	wire[2:0] w_n788_0;
	wire[2:0] w_n790_0;
	wire[2:0] w_n792_0;
	wire[2:0] w_n795_0;
	wire[1:0] w_n795_1;
	wire[2:0] w_n797_0;
	wire[2:0] w_n797_1;
	wire[2:0] w_n797_2;
	wire[2:0] w_n797_3;
	wire[2:0] w_n797_4;
	wire[2:0] w_n797_5;
	wire[2:0] w_n797_6;
	wire[2:0] w_n797_7;
	wire[2:0] w_n797_8;
	wire[1:0] w_n797_9;
	wire[2:0] w_n798_0;
	wire[1:0] w_n798_1;
	wire[2:0] w_n800_0;
	wire[2:0] w_n800_1;
	wire[2:0] w_n800_2;
	wire[2:0] w_n800_3;
	wire[1:0] w_n800_4;
	wire[2:0] w_n801_0;
	wire[1:0] w_n801_1;
	wire[2:0] w_n814_0;
	wire[2:0] w_n819_0;
	wire[1:0] w_n821_0;
	wire[1:0] w_n824_0;
	wire[1:0] w_n827_0;
	wire[1:0] w_n836_0;
	wire[1:0] w_n847_0;
	wire[2:0] w_n852_0;
	wire[2:0] w_n852_1;
	wire[2:0] w_n852_2;
	wire[2:0] w_n852_3;
	wire[2:0] w_n852_4;
	wire[2:0] w_n852_5;
	wire[2:0] w_n852_6;
	wire[2:0] w_n852_7;
	wire[2:0] w_n852_8;
	wire[1:0] w_n852_9;
	wire[2:0] w_n854_0;
	wire[2:0] w_n854_1;
	wire[2:0] w_n854_2;
	wire[2:0] w_n854_3;
	wire[1:0] w_n854_4;
	wire[2:0] w_n865_0;
	wire[1:0] w_n867_0;
	wire[1:0] w_n868_0;
	wire[1:0] w_n870_0;
	wire[1:0] w_n871_0;
	wire[1:0] w_n880_0;
	wire[1:0] w_n890_0;
	wire[1:0] w_n901_0;
	wire[2:0] w_n923_0;
	wire[1:0] w_n935_0;
	wire[2:0] w_n938_0;
	wire[2:0] w_n940_0;
	wire[1:0] w_n940_1;
	wire[1:0] w_n944_0;
	wire[1:0] w_n949_0;
	wire[1:0] w_n953_0;
	wire[2:0] w_n954_0;
	wire[1:0] w_n957_0;
	wire[1:0] w_n962_0;
	wire[1:0] w_n964_0;
	wire[1:0] w_n969_0;
	wire[2:0] w_n977_0;
	wire[1:0] w_n981_0;
	wire[1:0] w_n986_0;
	wire[1:0] w_n989_0;
	wire[2:0] w_n993_0;
	wire[2:0] w_n993_1;
	wire[2:0] w_n993_2;
	wire[2:0] w_n993_3;
	wire[2:0] w_n993_4;
	wire[2:0] w_n994_0;
	wire[2:0] w_n994_1;
	wire[2:0] w_n994_2;
	wire[2:0] w_n994_3;
	wire[1:0] w_n994_4;
	wire[2:0] w_n996_0;
	wire[2:0] w_n996_1;
	wire[2:0] w_n996_2;
	wire[2:0] w_n996_3;
	wire[1:0] w_n996_4;
	wire[2:0] w_n999_0;
	wire[2:0] w_n999_1;
	wire[2:0] w_n999_2;
	wire[2:0] w_n999_3;
	wire[2:0] w_n1007_0;
	wire[2:0] w_n1007_1;
	wire[2:0] w_n1007_2;
	wire[2:0] w_n1007_3;
	wire[2:0] w_n1008_0;
	wire[2:0] w_n1008_1;
	wire[2:0] w_n1008_2;
	wire[2:0] w_n1008_3;
	wire[2:0] w_n1008_4;
	wire[2:0] w_n1012_0;
	wire[2:0] w_n1012_1;
	wire[2:0] w_n1012_2;
	wire[2:0] w_n1012_3;
	wire[1:0] w_n1012_4;
	wire[2:0] w_n1014_0;
	wire[2:0] w_n1014_1;
	wire[2:0] w_n1014_2;
	wire[2:0] w_n1014_3;
	wire[1:0] w_n1014_4;
	wire[2:0] w_n1019_0;
	wire[1:0] w_n1019_1;
	wire[2:0] w_n1021_0;
	wire[1:0] w_n1021_1;
	wire[2:0] w_n1030_0;
	wire[1:0] w_n1030_1;
	wire[2:0] w_n1032_0;
	wire[1:0] w_n1032_1;
	wire[2:0] w_n1041_0;
	wire[1:0] w_n1041_1;
	wire[2:0] w_n1043_0;
	wire[1:0] w_n1043_1;
	wire[2:0] w_n1052_0;
	wire[1:0] w_n1052_1;
	wire[2:0] w_n1054_0;
	wire[1:0] w_n1054_1;
	wire[1:0] w_n1177_0;
	wire[1:0] w_n1179_0;
	wire[2:0] w_n1196_0;
	wire[2:0] w_n1196_1;
	wire[2:0] w_n1201_0;
	wire[2:0] w_n1205_0;
	wire[2:0] w_n1205_1;
	wire[2:0] w_n1213_0;
	wire[2:0] w_n1213_1;
	wire[2:0] w_n1236_0;
	wire[2:0] w_n1236_1;
	wire[2:0] w_n1251_0;
	wire[2:0] w_n1251_1;
	wire[2:0] w_n1279_0;
	wire[1:0] w_n1279_1;
	wire[2:0] w_n1297_0;
	wire[1:0] w_n1297_1;
	wire[2:0] w_n1299_0;
	wire[1:0] w_n1299_1;
	wire[2:0] w_n1410_0;
	wire[2:0] w_n1412_0;
	wire[1:0] w_n1416_0;
	wire[1:0] w_n1422_0;
	wire[1:0] w_n1425_0;
	wire[1:0] w_n1428_0;
	wire[1:0] w_n1429_0;
	wire[1:0] w_n1451_0;
	wire[1:0] w_n1503_0;
	wire[1:0] w_n1504_0;
	wire[1:0] w_n1592_0;
	wire[1:0] w_n1593_0;
	wire[1:0] w_n1596_0;
	wire[1:0] w_n1599_0;
	wire[1:0] w_n1603_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1609_0;
	wire[2:0] w_n1611_0;
	wire[1:0] w_n1613_0;
	wire[1:0] w_n1615_0;
	wire[1:0] w_n1618_0;
	wire[1:0] w_n1633_0;
	wire[1:0] w_n1637_0;
	wire[1:0] w_n1643_0;
	wire[1:0] w_n1652_0;
	wire[1:0] w_n1665_0;
	wire[2:0] w_n1674_0;
	wire[1:0] w_n1675_0;
	wire[2:0] w_n1679_0;
	wire[1:0] w_n1680_0;
	wire[1:0] w_n1694_0;
	wire[1:0] w_n1695_0;
	wire[1:0] w_n1698_0;
	wire w_dff_B_5pseY3ze5_1;
	wire w_dff_B_5d0LIbSn2_0;
	wire w_dff_B_gZLfCesE0_1;
	wire w_dff_B_XXGaiOMy4_1;
	wire w_dff_B_uZZ3q6Nx0_2;
	wire w_dff_B_3l13xEUy4_1;
	wire w_dff_B_uWMWTVN67_1;
	wire w_dff_B_0UaRHFHX3_0;
	wire w_dff_B_1gs4QHJx1_1;
	wire w_dff_B_rtRIxOw27_1;
	wire w_dff_B_fcKXeWTj0_0;
	wire w_dff_B_U8XNJdiR0_1;
	wire w_dff_A_QQ8poydE2_0;
	wire w_dff_A_Vom0CuN06_0;
	wire w_dff_A_nxHYnxi72_0;
	wire w_dff_A_QsBAZN6D1_0;
	wire w_dff_A_p77QdkLy9_1;
	wire w_dff_A_XtZe12Jn2_1;
	wire w_dff_A_nZjOPtI04_1;
	wire w_dff_A_4zSc1LyP2_1;
	wire w_dff_B_49CQMAWp8_1;
	wire w_dff_B_mV6sOTPV5_0;
	wire w_dff_B_dxVJs3kJ3_1;
	wire w_dff_B_JNlV6HdC8_1;
	wire w_dff_B_24q7TdUc7_1;
	wire w_dff_B_TonoSrvx8_1;
	wire w_dff_A_sfF8rck74_0;
	wire w_dff_A_LxfFmvmr5_1;
	wire w_dff_A_RnnwGZJ82_1;
	wire w_dff_A_wf2fsBPP2_1;
	wire w_dff_A_x0BvDMD32_1;
	wire w_dff_A_4zGRtotu7_1;
	wire w_dff_A_LO9HR7Du4_2;
	wire w_dff_A_9sIB7H2L7_2;
	wire w_dff_A_LAtJFuWb8_2;
	wire w_dff_A_TccOO6vn9_2;
	wire w_dff_B_JiQHGNmO2_1;
	wire w_dff_B_hKIdI6aE7_2;
	wire w_dff_B_fOGWVeyJ0_2;
	wire w_dff_B_Apk4W4Cq7_2;
	wire w_dff_B_HaW6KD374_2;
	wire w_dff_B_5scfG8PG4_1;
	wire w_dff_B_C0HkSu132_1;
	wire w_dff_B_OtJkf61N6_1;
	wire w_dff_B_lNqwqNLr0_1;
	wire w_dff_B_t2G5m4Xl0_1;
	wire w_dff_B_9A2iSTBK3_1;
	wire w_dff_B_gcvUXHpN5_1;
	wire w_dff_B_dM0hsl3E7_1;
	wire w_dff_B_kovXpwa96_1;
	wire w_dff_B_v9eAHOge7_1;
	wire w_dff_B_cb2UIZEQ3_1;
	wire w_dff_A_TBJLgtFH8_1;
	wire w_dff_A_wK0ga2Vk4_1;
	wire w_dff_B_Y78scTpD4_3;
	wire w_dff_B_7f7BGebr2_2;
	wire w_dff_B_59QTf0HI5_2;
	wire w_dff_B_ip4JU1t60_1;
	wire w_dff_B_lgf4lBax9_1;
	wire w_dff_A_h1J2x2Ra4_0;
	wire w_dff_A_75yJteUV9_0;
	wire w_dff_A_1nYH5uZI8_0;
	wire w_dff_A_szz1ylTx7_0;
	wire w_dff_A_q7uSuu5a5_0;
	wire w_dff_B_OW6jf2Sd3_0;
	wire w_dff_B_WgOLK0H23_0;
	wire w_dff_B_cEH97czM1_0;
	wire w_dff_B_dJCb12AO3_0;
	wire w_dff_B_r7lcnJvL4_0;
	wire w_dff_B_7vEWjXbf7_0;
	wire w_dff_B_pjcJhtvT5_0;
	wire w_dff_B_9Z1qVH0j7_0;
	wire w_dff_B_aCMTOUZe0_0;
	wire w_dff_B_YQx7uU1H6_0;
	wire w_dff_B_6UaTBp6x0_0;
	wire w_dff_A_yvkTFnJ01_1;
	wire w_dff_A_QbrgWKe19_1;
	wire w_dff_A_cRhSMklw6_1;
	wire w_dff_A_Hmk375zk1_1;
	wire w_dff_A_XS65W3Tb0_1;
	wire w_dff_A_XLu2d7qV7_1;
	wire w_dff_A_ffpR4mWY8_1;
	wire w_dff_A_hfbZ9uG27_1;
	wire w_dff_A_NKHrKRDb4_1;
	wire w_dff_A_jwufuSU28_1;
	wire w_dff_B_dxadoulk7_0;
	wire w_dff_B_nflMTdIG9_0;
	wire w_dff_B_xvDPDxmy0_0;
	wire w_dff_B_o0ptTId29_0;
	wire w_dff_B_qOKjY7rs7_0;
	wire w_dff_B_yVBOucxr8_0;
	wire w_dff_B_AYQD91Uo5_0;
	wire w_dff_B_uhReZfBD9_0;
	wire w_dff_B_adVclcQ96_0;
	wire w_dff_B_9jj3DoR38_0;
	wire w_dff_B_D334u1qO2_2;
	wire w_dff_B_0IFzQppa9_0;
	wire w_dff_A_BM69SWUv2_1;
	wire w_dff_A_M8Q9Df9q4_1;
	wire w_dff_A_ASZC6nE61_1;
	wire w_dff_A_NASzT5FX1_1;
	wire w_dff_A_ATEQW8G72_1;
	wire w_dff_A_1GaqXvWj0_1;
	wire w_dff_A_IvliJj7m2_1;
	wire w_dff_A_1jJHwIJK8_1;
	wire w_dff_A_4MVfoLgo8_1;
	wire w_dff_A_nQHq9kuD5_1;
	wire w_dff_B_QIMtgdLF5_0;
	wire w_dff_B_MCoew3nT4_1;
	wire w_dff_B_KbbBnvZI2_1;
	wire w_dff_B_RH5sCLMh0_1;
	wire w_dff_B_LNKh3xgB8_0;
	wire w_dff_B_MsSxupwE8_1;
	wire w_dff_B_gwZZCsGf6_1;
	wire w_dff_B_xUjzgfDb8_1;
	wire w_dff_B_AG9aNpSz3_1;
	wire w_dff_B_cA5UtwHA5_1;
	wire w_dff_B_hTywLHFX4_1;
	wire w_dff_B_AUY7s4db5_1;
	wire w_dff_B_Qya5qyKF1_1;
	wire w_dff_B_EN9kUsYt2_1;
	wire w_dff_B_LGtJH1MA6_1;
	wire w_dff_B_rLse5twH7_1;
	wire w_dff_B_dyr2GmnC0_1;
	wire w_dff_B_QOBSfU5f1_1;
	wire w_dff_B_WGGjwLHl1_1;
	wire w_dff_B_oNDzFxhm3_1;
	wire w_dff_B_1dDUVuTi6_1;
	wire w_dff_B_Ynynngap4_1;
	wire w_dff_B_96gCK1kk3_1;
	wire w_dff_B_Bj8SxTbY3_1;
	wire w_dff_B_OHythTkV1_1;
	wire w_dff_B_E5dUUKBX6_1;
	wire w_dff_B_SGWjoghx5_1;
	wire w_dff_B_8CAnK0on1_1;
	wire w_dff_B_atnPbo0f4_1;
	wire w_dff_B_L1Ma3WVe6_1;
	wire w_dff_B_j6UYEdby3_1;
	wire w_dff_B_2ozp6x2H3_1;
	wire w_dff_B_zHVZMFQC0_1;
	wire w_dff_B_wixnft3X6_1;
	wire w_dff_B_LB8GxHHJ9_0;
	wire w_dff_B_umFULM2S3_0;
	wire w_dff_B_xcyEfhkz8_0;
	wire w_dff_B_IHGACzIj0_0;
	wire w_dff_B_kshCvsy17_0;
	wire w_dff_B_2T2lo8qZ5_0;
	wire w_dff_B_iakkHnI28_0;
	wire w_dff_B_pGe9HiPR0_0;
	wire w_dff_B_wnqpi1zG9_0;
	wire w_dff_B_dzUXXO4t5_0;
	wire w_dff_B_jYwc0CJA9_0;
	wire w_dff_B_Er9MKswT7_1;
	wire w_dff_B_QwwoiTRd0_2;
	wire w_dff_B_4NfCGkbl4_2;
	wire w_dff_B_eZ8BiIdW9_2;
	wire w_dff_B_hG0UErfk8_1;
	wire w_dff_B_SaMigYhO5_1;
	wire w_dff_B_sObn9bEK3_1;
	wire w_dff_B_zUVC3qY25_1;
	wire w_dff_B_tcmkMNDz8_1;
	wire w_dff_B_n1ABL9mY3_1;
	wire w_dff_B_dyaOGlLv3_1;
	wire w_dff_B_8ZKG8dxr1_1;
	wire w_dff_B_zK5ZTSk17_0;
	wire w_dff_B_QgSZRQ2D7_1;
	wire w_dff_B_vfk6ABnv7_1;
	wire w_dff_A_rnixLMeT4_0;
	wire w_dff_A_QmtQyr2u7_0;
	wire w_dff_B_fSWHe2016_1;
	wire w_dff_B_6cjba8ES8_1;
	wire w_dff_B_412dZbzB8_1;
	wire w_dff_B_Evl6tKCs9_1;
	wire w_dff_B_9CjPmnQA1_1;
	wire w_dff_A_7iOJvDjX4_0;
	wire w_dff_A_vRVddJJz5_0;
	wire w_dff_A_CxBDqyPT0_0;
	wire w_dff_A_jdCE27XT0_0;
	wire w_dff_A_u4v0WMYu4_0;
	wire w_dff_A_ZXn6SsW18_0;
	wire w_dff_A_HOGXNGNK0_0;
	wire w_dff_A_jeVpKP5m4_0;
	wire w_dff_A_AVD6DKrQ3_0;
	wire w_dff_A_XotcTJEI5_0;
	wire w_dff_A_YzDgD4NE9_0;
	wire w_dff_B_tNxFShYp2_1;
	wire w_dff_B_QCr6Roxr9_1;
	wire w_dff_B_hem3m85J9_0;
	wire w_dff_B_jB9kaDXI6_0;
	wire w_dff_B_imStMAos3_0;
	wire w_dff_B_qpRosqnp9_0;
	wire w_dff_B_lPeYGUcP2_0;
	wire w_dff_B_xLM2x2TL0_0;
	wire w_dff_B_afLguixQ7_0;
	wire w_dff_B_J8SFRSD43_0;
	wire w_dff_B_TWNIPGHf4_0;
	wire w_dff_B_G0CDObb12_0;
	wire w_dff_B_6GrgtVyM6_0;
	wire w_dff_B_Lb0MexbC2_0;
	wire w_dff_B_Yw796fOH8_0;
	wire w_dff_B_DUIetwC06_0;
	wire w_dff_B_sfwCod1Y0_0;
	wire w_dff_B_XbfJ5Bvn5_0;
	wire w_dff_B_0j02iMEa7_1;
	wire w_dff_A_vdnHW2mK9_0;
	wire w_dff_A_CNfTMicX7_0;
	wire w_dff_A_DiHdsEXo0_0;
	wire w_dff_A_eCkujpTU6_0;
	wire w_dff_A_KOlomuab5_0;
	wire w_dff_A_HjnkrWBB2_0;
	wire w_dff_A_7SbTxlr39_0;
	wire w_dff_B_aZnhjJwS1_0;
	wire w_dff_B_HGXdE1JU2_0;
	wire w_dff_B_wbHK1kru7_0;
	wire w_dff_B_1ORWIEv39_0;
	wire w_dff_B_whN8cBP94_0;
	wire w_dff_B_JmR7KTY56_0;
	wire w_dff_B_Xzul8GGG7_0;
	wire w_dff_B_ezuhTk814_0;
	wire w_dff_B_dnpunXcO3_0;
	wire w_dff_B_xCa9bdv23_0;
	wire w_dff_B_kQjoGtDh7_0;
	wire w_dff_B_EO0LESZg7_0;
	wire w_dff_B_8LpmW8yO4_0;
	wire w_dff_B_CE7e9NrA5_0;
	wire w_dff_B_MzogfC1j1_0;
	wire w_dff_B_ewZDUYYX1_1;
	wire w_dff_B_Hp4BtsS16_1;
	wire w_dff_A_1SidvPKG3_0;
	wire w_dff_A_gQlOEQWk7_0;
	wire w_dff_A_FoGlKVWx7_0;
	wire w_dff_A_VSuBAylf6_0;
	wire w_dff_A_9Pp4vPt31_0;
	wire w_dff_A_fweZvjD31_0;
	wire w_dff_A_qZRtGKRU3_0;
	wire w_dff_A_MuP6YyT31_0;
	wire w_dff_A_pP6kBUgi0_0;
	wire w_dff_A_EEv23slt9_0;
	wire w_dff_A_ok7JKiik8_0;
	wire w_dff_A_Jftb7nTX1_0;
	wire w_dff_A_m5XKEMfx7_0;
	wire w_dff_A_JjJ0bDPt0_0;
	wire w_dff_A_neKuS7Eu8_0;
	wire w_dff_A_9iDDQStT0_2;
	wire w_dff_A_aaEC14nC7_2;
	wire w_dff_A_zWgHIMGW7_2;
	wire w_dff_A_LPEzXf2q2_2;
	wire w_dff_A_jAa0sGrV2_2;
	wire w_dff_A_KdxEX8AO0_2;
	wire w_dff_A_XHQqgWwY6_2;
	wire w_dff_A_fpgmwc9O5_2;
	wire w_dff_A_xEIdpfM55_2;
	wire w_dff_A_rjsII0Je5_2;
	wire w_dff_A_MOpea18H8_2;
	wire w_dff_A_oe67f4Qu4_2;
	wire w_dff_A_01MzUA0w5_2;
	wire w_dff_A_jNCimEpT6_2;
	wire w_dff_A_3ssK2ygp8_2;
	wire w_dff_A_zDaWfg2a1_2;
	wire w_dff_A_ZAGSIkLI4_0;
	wire w_dff_A_v4x7lXO91_0;
	wire w_dff_A_FdnfLvON5_0;
	wire w_dff_A_CpOhPon59_0;
	wire w_dff_A_Qfb5vhqN4_0;
	wire w_dff_A_gEPDidKX5_0;
	wire w_dff_A_Ppaf1Vnl2_0;
	wire w_dff_A_jeZCQKRq0_0;
	wire w_dff_A_6QQgHyQG6_0;
	wire w_dff_A_ZqnhYi1e2_0;
	wire w_dff_A_mwdqPnKb4_0;
	wire w_dff_A_bKBLcDTV3_0;
	wire w_dff_A_WkEANbXK0_0;
	wire w_dff_A_ou2QQ6fy9_2;
	wire w_dff_A_c5Dp73J89_2;
	wire w_dff_A_Hix2Sr1j7_2;
	wire w_dff_A_RlbRqm319_2;
	wire w_dff_A_SIXkhWH32_2;
	wire w_dff_A_kOVtR4pq6_2;
	wire w_dff_A_REWzpq9E4_2;
	wire w_dff_A_UlP05Wkw8_2;
	wire w_dff_A_RGWDA76O5_2;
	wire w_dff_A_HrUtZ42O6_2;
	wire w_dff_A_7vAGRxiF9_2;
	wire w_dff_A_PThipe6u7_2;
	wire w_dff_A_ydXySLI27_2;
	wire w_dff_A_dpNgruTi0_2;
	wire w_dff_A_DhSM3jhv1_2;
	wire w_dff_B_PpPZ4mCF7_0;
	wire w_dff_B_buytFbIi2_0;
	wire w_dff_B_SUfuZQEe8_0;
	wire w_dff_B_d4GLyjtf2_0;
	wire w_dff_B_crnmLoxB9_0;
	wire w_dff_B_Zv9QWa687_0;
	wire w_dff_B_SnANx2NB0_0;
	wire w_dff_B_mhTozrtV2_0;
	wire w_dff_B_dsIZujJ90_0;
	wire w_dff_B_xhMl4xgP7_0;
	wire w_dff_B_mkGZjtUB5_0;
	wire w_dff_B_3nORkulA1_0;
	wire w_dff_B_Yerqif9U3_0;
	wire w_dff_B_GSF4OTTx6_1;
	wire w_dff_A_n29bVcSe6_1;
	wire w_dff_A_bJHrf9zj4_1;
	wire w_dff_A_bXIbCL2N4_1;
	wire w_dff_A_PnZuGu2T4_1;
	wire w_dff_A_puB3p0UK8_1;
	wire w_dff_A_g03S2BFt7_1;
	wire w_dff_A_m6QhEtQX8_1;
	wire w_dff_A_zmH8t6tw7_1;
	wire w_dff_A_B5ruK8Uz3_1;
	wire w_dff_A_fxnPmKbg2_1;
	wire w_dff_A_VFQbVcPE5_1;
	wire w_dff_A_ktRA898b1_1;
	wire w_dff_A_axkdoY4Q0_1;
	wire w_dff_A_7M0IHwGm2_1;
	wire w_dff_A_bxoWGViU6_1;
	wire w_dff_A_01JYIkab4_1;
	wire w_dff_A_UUIxNnyx7_1;
	wire w_dff_A_gvF91yLG1_1;
	wire w_dff_A_veiMbtOw5_1;
	wire w_dff_A_wBADW5Wd7_1;
	wire w_dff_A_n1dyIVjz4_1;
	wire w_dff_A_25f27IqB4_1;
	wire w_dff_A_c8QfGWm31_1;
	wire w_dff_A_9sSALoD26_1;
	wire w_dff_A_SGXCpmyO5_1;
	wire w_dff_B_dYn8RS1x1_0;
	wire w_dff_B_lH2NefW04_0;
	wire w_dff_B_eQRB0NKi3_0;
	wire w_dff_B_wsr3lvtj0_0;
	wire w_dff_B_rTMxEox44_0;
	wire w_dff_B_rAXi5MGZ2_0;
	wire w_dff_B_f3Ordk8G1_0;
	wire w_dff_B_4cf75ATx5_0;
	wire w_dff_B_qtS4LE9L9_0;
	wire w_dff_B_6e6VC4629_0;
	wire w_dff_B_1bNeTI3B4_0;
	wire w_dff_B_cmGXKS7h8_0;
	wire w_dff_B_2ufFjAIS4_0;
	wire w_dff_B_NXlOkNV54_0;
	wire w_dff_B_Vs09V1U34_1;
	wire w_dff_B_OVdatxwx6_1;
	wire w_dff_B_XPkTXUtv3_1;
	wire w_dff_A_nbDlv0sp1_0;
	wire w_dff_A_UWVHTOkT5_2;
	wire w_dff_A_LYsHmIKq1_2;
	wire w_dff_B_Vok9Jdl50_1;
	wire w_dff_B_pbBmfKE70_1;
	wire w_dff_B_cm38cG3f5_1;
	wire w_dff_B_VnpyObGo1_1;
	wire w_dff_B_PCmAm8xV7_1;
	wire w_dff_B_RPERlSfS4_1;
	wire w_dff_B_wlMOJKNq7_1;
	wire w_dff_B_GSrExPpn2_1;
	wire w_dff_B_fmHxdKZr7_1;
	wire w_dff_B_TpOQrr2C8_1;
	wire w_dff_B_XXZ18Gv14_1;
	wire w_dff_B_WXInNCAx2_1;
	wire w_dff_B_shGYiVLn1_1;
	wire w_dff_B_WBzlmFzL0_1;
	wire w_dff_B_IZm3Gvzd0_1;
	wire w_dff_A_VW3jl7Ex2_0;
	wire w_dff_A_79Oez01Q9_0;
	wire w_dff_A_D2NTLLU55_0;
	wire w_dff_A_eYo1lnmW7_0;
	wire w_dff_A_6JZNvong7_0;
	wire w_dff_A_CiWSb2bP5_0;
	wire w_dff_A_1AhnXBIo2_0;
	wire w_dff_A_Y9uM1MYt2_0;
	wire w_dff_B_7alQrAGz6_1;
	wire w_dff_B_JwnPyo986_1;
	wire w_dff_B_lHCNbdw67_2;
	wire w_dff_B_Or7ieCL40_1;
	wire w_dff_B_jyW51YLO6_1;
	wire w_dff_B_Ti1HaDSO1_1;
	wire w_dff_B_VK6F6Gs06_1;
	wire w_dff_B_LqmTnlO72_1;
	wire w_dff_B_6kmkD8AC8_1;
	wire w_dff_B_n506kiGD5_1;
	wire w_dff_B_xL2ZF1gM3_1;
	wire w_dff_B_ZH1SJDAf2_1;
	wire w_dff_B_dpwT5ush0_1;
	wire w_dff_B_uu52JJP23_1;
	wire w_dff_B_ke0txx4M7_1;
	wire w_dff_B_BaNWfyXH9_1;
	wire w_dff_B_3PqhCcif5_1;
	wire w_dff_B_OTTsIfBA1_0;
	wire w_dff_B_O6sgrkC04_1;
	wire w_dff_B_z2wmbyYC3_1;
	wire w_dff_A_6ugtbfPB3_1;
	wire w_dff_A_oh1lAM2o7_1;
	wire w_dff_A_u3l2NVtL2_1;
	wire w_dff_A_s6fVlPWS9_1;
	wire w_dff_A_qweThpfB5_1;
	wire w_dff_A_OU2kOwBn0_1;
	wire w_dff_A_zPAMdFSs7_1;
	wire w_dff_A_yCh42Enh1_1;
	wire w_dff_A_gdzIDZF52_1;
	wire w_dff_A_mTP01M8b7_1;
	wire w_dff_A_hwpktazI0_1;
	wire w_dff_A_bEnidND31_1;
	wire w_dff_A_wMdmBG4W9_1;
	wire w_dff_A_PgdRUJlY1_1;
	wire w_dff_A_fbZ2eGkt8_1;
	wire w_dff_B_2S5587Jz0_2;
	wire w_dff_A_z3IMOOoq7_1;
	wire w_dff_A_a4w9YAAH5_1;
	wire w_dff_A_tzjLVKs71_1;
	wire w_dff_A_IaYJB8XB0_1;
	wire w_dff_A_yWUBgGhE0_1;
	wire w_dff_A_U3azGVav7_1;
	wire w_dff_A_34zAk1gL3_1;
	wire w_dff_A_aQsWuZ0H7_1;
	wire w_dff_A_oK0W2Tqd0_1;
	wire w_dff_A_8Y5jKg274_1;
	wire w_dff_A_r9bJ7dDD4_1;
	wire w_dff_A_xNCVyGLH7_1;
	wire w_dff_A_lIpPLIlz4_1;
	wire w_dff_A_PJktRTXK0_1;
	wire w_dff_A_wbLq5Ln62_1;
	wire w_dff_A_WeY6qbfv3_1;
	wire w_dff_B_XLnPo97s6_1;
	wire w_dff_B_9Hi7TPf16_1;
	wire w_dff_B_nx7no1rL6_1;
	wire w_dff_B_B6MzBm4y3_1;
	wire w_dff_B_2Oqfe33G1_1;
	wire w_dff_B_9lMLVFMa8_1;
	wire w_dff_B_2GOZwkDz6_1;
	wire w_dff_B_CvbipimJ4_1;
	wire w_dff_B_1UWSti0X0_1;
	wire w_dff_B_TzLFqooJ8_1;
	wire w_dff_B_iadIqWnp5_1;
	wire w_dff_B_CMFnyfac9_1;
	wire w_dff_B_1pUSJGLJ6_1;
	wire w_dff_B_f9HXrqET1_1;
	wire w_dff_A_QIGa4Vxw0_0;
	wire w_dff_A_jR5m4kYB0_0;
	wire w_dff_A_YBwAHMoQ3_0;
	wire w_dff_A_VUc2TGVB7_0;
	wire w_dff_A_M4JBrh589_0;
	wire w_dff_A_XTX7mUEQ6_0;
	wire w_dff_A_JkH3f71n7_0;
	wire w_dff_A_0xeiQsgV3_0;
	wire w_dff_A_zgYvJxwK8_0;
	wire w_dff_A_8Y89BlU08_0;
	wire w_dff_A_TPAe0JcF3_0;
	wire w_dff_A_VSekOTg48_0;
	wire w_dff_A_jcig5Us53_2;
	wire w_dff_A_D6EBUCPr5_2;
	wire w_dff_A_KeX40C7E4_2;
	wire w_dff_A_Nx206cUP8_2;
	wire w_dff_A_2iImcXw27_2;
	wire w_dff_A_T0lbkzxz2_2;
	wire w_dff_A_XFKTu5Ma0_2;
	wire w_dff_A_wWADclJz7_2;
	wire w_dff_A_r2F5r87r9_2;
	wire w_dff_A_0nm2xijW1_2;
	wire w_dff_A_x0KPSQ9a9_2;
	wire w_dff_A_pqzAX0Kb3_2;
	wire w_dff_A_gQ0ePflD6_2;
	wire w_dff_B_kXvSSlQq3_2;
	wire w_dff_A_EVSU5lyt1_0;
	wire w_dff_A_9dcVJLK39_0;
	wire w_dff_A_ScFoQiCK6_0;
	wire w_dff_A_UaGggClO3_0;
	wire w_dff_A_ODBnUjcP9_0;
	wire w_dff_A_aq99JOlU2_0;
	wire w_dff_A_WdATVlpF8_0;
	wire w_dff_A_U8WVisHU5_0;
	wire w_dff_A_6ZccGNd50_0;
	wire w_dff_A_uCiFszMf5_0;
	wire w_dff_A_vsvynI6l4_0;
	wire w_dff_A_Cq8pswRj8_0;
	wire w_dff_A_ttTEApFA6_0;
	wire w_dff_A_ljERb6es5_2;
	wire w_dff_A_pDi6sdYw2_2;
	wire w_dff_A_4GRQRVfW1_2;
	wire w_dff_A_Zf8PCDGj7_2;
	wire w_dff_A_dcOF4l9u1_2;
	wire w_dff_A_blIdSm9Z9_2;
	wire w_dff_A_njF9yI397_2;
	wire w_dff_A_hKxsYyVD2_2;
	wire w_dff_A_Dd0CuaQU7_2;
	wire w_dff_A_MfHzTLBw5_2;
	wire w_dff_A_bUuxeHB43_2;
	wire w_dff_A_X0pE9JoL7_2;
	wire w_dff_A_pdByMsJz9_2;
	wire w_dff_A_D48t4b391_2;
	wire w_dff_A_AtGQZzA59_2;
	wire w_dff_B_jTMkOXTe0_0;
	wire w_dff_B_AnWszdc59_0;
	wire w_dff_B_nDCKo3bF5_0;
	wire w_dff_B_rFulOtJ36_0;
	wire w_dff_B_0rAR0gjE5_0;
	wire w_dff_B_jBCxrajO0_0;
	wire w_dff_B_PZTJQhVQ7_0;
	wire w_dff_B_smqajFHb2_0;
	wire w_dff_B_BANfFmOR9_0;
	wire w_dff_B_8MOYsacq3_0;
	wire w_dff_B_15W2sopy9_0;
	wire w_dff_B_3yet1Eid8_0;
	wire w_dff_B_bccQQaUr7_0;
	wire w_dff_B_LKSFC2wQ7_0;
	wire w_dff_A_klxH40F92_1;
	wire w_dff_A_7JjJKAlK5_2;
	wire w_dff_B_OdJBfi1i5_2;
	wire w_dff_B_VgSWLDu21_1;
	wire w_dff_B_X2FQN6vl5_1;
	wire w_dff_B_e1PvzZF09_1;
	wire w_dff_A_PJpeYuDT6_2;
	wire w_dff_A_tfvNvX5W5_2;
	wire w_dff_B_ASjmq8333_0;
	wire w_dff_B_Hj3oGY198_0;
	wire w_dff_B_rDbHduqH3_0;
	wire w_dff_B_nBDadRNt4_0;
	wire w_dff_B_jggZGPEQ4_0;
	wire w_dff_B_HsfYJFYe5_0;
	wire w_dff_B_Lk9noBZP0_0;
	wire w_dff_B_EIfO8b2u0_0;
	wire w_dff_B_xPAqGxKl7_0;
	wire w_dff_B_JOPDo2TI9_0;
	wire w_dff_B_ipUpO3rW9_0;
	wire w_dff_B_aDUJAUWH2_0;
	wire w_dff_B_Fjx6FOmC5_0;
	wire w_dff_B_mH6hBIym7_0;
	wire w_dff_B_URYxDwxI2_0;
	wire w_dff_B_BcTWHefg0_0;
	wire w_dff_B_JeJ532NP3_1;
	wire w_dff_B_KfFW1Fkk3_0;
	wire w_dff_B_ywbCWTgM4_0;
	wire w_dff_B_prB4rSPH2_0;
	wire w_dff_B_4TUwwte84_0;
	wire w_dff_B_GIcoci6S0_0;
	wire w_dff_B_PYiQKGSz9_0;
	wire w_dff_B_Pr2RB04Y5_0;
	wire w_dff_B_5TMt0c0u6_0;
	wire w_dff_B_S8q2Y4OC4_0;
	wire w_dff_B_HnqMlbLq3_0;
	wire w_dff_B_G7x6S2a65_0;
	wire w_dff_B_VxYJZoC49_0;
	wire w_dff_B_ZTwiHh5O9_0;
	wire w_dff_B_YAFkuvKh2_0;
	wire w_dff_A_Ni8pVGn12_0;
	wire w_dff_A_EFk0UZYV1_0;
	wire w_dff_A_iItlQ5sG3_0;
	wire w_dff_A_sZ7qQDgD8_1;
	wire w_dff_A_O9LgnZvy7_1;
	wire w_dff_A_jLVWflxl8_1;
	wire w_dff_A_2d3zzqSu0_1;
	wire w_dff_A_o7fd8FI87_1;
	wire w_dff_A_WjqiIhQa3_1;
	wire w_dff_A_CZiGEFGF6_1;
	wire w_dff_A_zBqjoj2v6_0;
	wire w_dff_A_O75CPJQW1_0;
	wire w_dff_A_PDtPIIxj8_0;
	wire w_dff_A_sPNwTG3r6_0;
	wire w_dff_A_QuEJt7JU6_0;
	wire w_dff_A_m4anppy54_1;
	wire w_dff_A_mWAL1dEc8_1;
	wire w_dff_A_pe7FpfbB5_1;
	wire w_dff_A_UK5h9lDg4_1;
	wire w_dff_A_umvdPpb11_1;
	wire w_dff_A_9ya0V2IF3_1;
	wire w_dff_A_90mI8wQY7_1;
	wire w_dff_B_WgLtXsRa3_0;
	wire w_dff_B_dpcbcZS22_0;
	wire w_dff_B_FXWbEvUQ8_0;
	wire w_dff_B_IwjpEjEa5_0;
	wire w_dff_B_yvqEcoX00_0;
	wire w_dff_B_hi1waNrn4_0;
	wire w_dff_B_UvOcAHl45_0;
	wire w_dff_B_PzumL7cK2_0;
	wire w_dff_B_uvcy7Fap1_0;
	wire w_dff_B_qhTRHxet7_0;
	wire w_dff_B_823xxaS29_0;
	wire w_dff_B_93Pkxbgz0_0;
	wire w_dff_B_qeCi42wT9_0;
	wire w_dff_B_3QEbJYIQ0_1;
	wire w_dff_A_GqhGK6Ko6_2;
	wire w_dff_A_iozQxqyE8_2;
	wire w_dff_A_RkhToDx10_2;
	wire w_dff_B_kqndtGmv5_0;
	wire w_dff_B_becFu0ta7_0;
	wire w_dff_B_WoZs7mQy0_0;
	wire w_dff_B_rCpMffo45_0;
	wire w_dff_B_l0rf3xqv1_0;
	wire w_dff_B_GkCLHMos6_0;
	wire w_dff_B_jJdAtBfJ7_0;
	wire w_dff_B_H8GxjWtT6_0;
	wire w_dff_B_Z2I8Q26F6_0;
	wire w_dff_B_qb0oIRn35_0;
	wire w_dff_B_llJ7JzUh5_0;
	wire w_dff_B_EcZf0wcu0_0;
	wire w_dff_B_Zp7KqYat4_0;
	wire w_dff_B_P8C265hN7_0;
	wire w_dff_A_TGCFqqnx8_0;
	wire w_dff_A_IhOTjENe3_0;
	wire w_dff_A_qCkbwAAw0_1;
	wire w_dff_B_Mg9EJ5kz0_1;
	wire w_dff_B_LLmtF0zo3_1;
	wire w_dff_B_qJu1NlfA0_1;
	wire w_dff_B_rvQOjbCt1_1;
	wire w_dff_B_Svymtap50_1;
	wire w_dff_B_4tNpsCiz0_1;
	wire w_dff_B_Zk5OPS667_1;
	wire w_dff_B_EKj1OGyS0_1;
	wire w_dff_B_JPxczKMH0_1;
	wire w_dff_B_lihhcyfF2_1;
	wire w_dff_B_nTKZW1Cr2_1;
	wire w_dff_B_0Qevwsqk0_1;
	wire w_dff_B_v8txGR5D8_1;
	wire w_dff_B_OGJYKypv5_1;
	wire w_dff_B_Jum9HHgx3_1;
	wire w_dff_B_34ILIyfT2_1;
	wire w_dff_B_YPte2gEs3_1;
	wire w_dff_B_EA3HTJ9z4_1;
	wire w_dff_B_vx3EQJt79_1;
	wire w_dff_B_3sRK3wxY0_1;
	wire w_dff_B_YlHWyepJ5_1;
	wire w_dff_B_5iW68SO90_1;
	wire w_dff_B_gXd6knBH9_1;
	wire w_dff_B_ZTf8MQTh6_1;
	wire w_dff_B_EEeSmgZ44_1;
	wire w_dff_B_FfwXozkg9_1;
	wire w_dff_B_kSkScJmV4_1;
	wire w_dff_B_UQrUsxZJ0_1;
	wire w_dff_B_APgQFSPT5_1;
	wire w_dff_B_Ddu4rOUr7_1;
	wire w_dff_B_UWwOies06_1;
	wire w_dff_B_FamlHe4h4_1;
	wire w_dff_B_M5ccVy9N4_1;
	wire w_dff_B_b0B1pIhC7_1;
	wire w_dff_B_ZFXfjuh32_1;
	wire w_dff_B_auqaRaO50_1;
	wire w_dff_B_8hmBxek14_1;
	wire w_dff_B_N33P6Y9g5_1;
	wire w_dff_B_7EHHcQ7p9_1;
	wire w_dff_B_RUU5PmNh1_1;
	wire w_dff_B_60Q6r02i0_1;
	wire w_dff_B_VBLEOHd63_1;
	wire w_dff_B_dDaX9vin5_1;
	wire w_dff_B_bvhI34cd3_1;
	wire w_dff_B_L8i3cC3X1_0;
	wire w_dff_B_VhaICDBA5_0;
	wire w_dff_B_Vj2hRPJ01_0;
	wire w_dff_B_Xsa2AxOe3_0;
	wire w_dff_B_9QOCPZyK3_0;
	wire w_dff_B_qH1jI7nu0_0;
	wire w_dff_B_HCIzJQ130_1;
	wire w_dff_B_6jRaOUUu8_1;
	wire w_dff_B_ha0atSkg5_1;
	wire w_dff_B_l2sgmT7n1_1;
	wire w_dff_B_9llXinuz3_1;
	wire w_dff_B_w1vflgpN3_1;
	wire w_dff_B_DbDIyK689_1;
	wire w_dff_B_7lpTNgCX8_1;
	wire w_dff_B_PiyvcPOW4_1;
	wire w_dff_B_JgNojHL90_1;
	wire w_dff_B_YBylxNfk1_1;
	wire w_dff_B_AO4fSm5S0_1;
	wire w_dff_B_iQuXzvXk5_1;
	wire w_dff_B_3Z7GaG621_1;
	wire w_dff_B_wyxXsqek5_1;
	wire w_dff_B_Zoh1sYfm8_1;
	wire w_dff_B_qcUKq5av0_1;
	wire w_dff_B_DowEpmwH5_1;
	wire w_dff_B_WwJ0NSWx1_1;
	wire w_dff_B_JfwrxIuU8_0;
	wire w_dff_B_RXLcMShc3_0;
	wire w_dff_B_ZNulepyy7_0;
	wire w_dff_B_9p04cYS64_0;
	wire w_dff_B_9wyuRh0q9_0;
	wire w_dff_B_mXSWqqI47_0;
	wire w_dff_B_iLPynGW98_1;
	wire w_dff_B_Xl5HX38I0_1;
	wire w_dff_B_1sVHQLs98_1;
	wire w_dff_B_qakfyPmS7_1;
	wire w_dff_B_33vZx0Wk4_2;
	wire w_dff_B_nOEfcpdq6_2;
	wire w_dff_B_Z7RccH1E0_2;
	wire w_dff_B_2uabgvoB1_0;
	wire w_dff_B_6yuWUfCZ6_0;
	wire w_dff_B_GoDZdDgy7_0;
	wire w_dff_B_YLSk5S105_0;
	wire w_dff_B_x8W7rtEd7_0;
	wire w_dff_B_caJdmGw79_0;
	wire w_dff_B_Mpn6ZRof5_0;
	wire w_dff_B_fssDAQDr5_0;
	wire w_dff_B_I09pJjqL9_0;
	wire w_dff_B_K7L63pMg9_0;
	wire w_dff_B_9pBGq7fL8_0;
	wire w_dff_B_0mHdEneZ3_0;
	wire w_dff_B_KoFZQHj32_0;
	wire w_dff_B_focYSCPh7_2;
	wire w_dff_B_y55UpSa60_2;
	wire w_dff_B_bLSBvltT6_2;
	wire w_dff_B_WevrzoMI7_0;
	wire w_dff_B_fCcYb1HK3_1;
	wire w_dff_B_u3X9cDNy1_1;
	wire w_dff_B_K1lhKfP65_1;
	wire w_dff_B_170aO85v8_1;
	wire w_dff_B_cpKPO1eC0_1;
	wire w_dff_B_4xRmqUBc3_1;
	wire w_dff_B_Zo5UtX9N0_0;
	wire w_dff_B_PgKBBWqC0_0;
	wire w_dff_B_3XH3aMG67_1;
	wire w_dff_B_aQUqQRTG7_1;
	wire w_dff_A_Fpaig06N3_0;
	wire w_dff_A_S3xNVy6Y3_0;
	wire w_dff_B_Bm6FwsJ27_1;
	wire w_dff_B_et0bOagX2_1;
	wire w_dff_B_yaRqtMlG8_1;
	wire w_dff_A_jx8wBfJg7_0;
	wire w_dff_A_GPrWgRHY4_1;
	wire w_dff_A_W3h0h3592_1;
	wire w_dff_A_b6OH5gk64_1;
	wire w_dff_A_3lodQBnn5_1;
	wire w_dff_A_IIYIDKfM5_1;
	wire w_dff_A_0UNvS99k5_1;
	wire w_dff_B_HH3jiI268_1;
	wire w_dff_B_uEG2tnnx6_1;
	wire w_dff_B_gT9CoaJA8_1;
	wire w_dff_B_PVwQTJdm6_1;
	wire w_dff_B_e3NDGQlq6_1;
	wire w_dff_B_Cy1N3WdK5_1;
	wire w_dff_B_IwJouphq5_1;
	wire w_dff_B_W86gbJTr4_1;
	wire w_dff_B_OhH9u7m70_0;
	wire w_dff_B_eMz8smkY6_0;
	wire w_dff_B_zszzuhX94_0;
	wire w_dff_B_5OSjEKub0_0;
	wire w_dff_B_ndtQ8J8A2_1;
	wire w_dff_B_1zB6cnra8_1;
	wire w_dff_B_6ggxj0f47_0;
	wire w_dff_B_bXxiS1Vt8_0;
	wire w_dff_B_gIJJEWgu0_0;
	wire w_dff_B_xI1S3T0I1_0;
	wire w_dff_A_A1X0X5sl5_0;
	wire w_dff_A_r1D25C2M4_0;
	wire w_dff_A_gUq2Ekrx3_0;
	wire w_dff_A_dCKwEEz49_0;
	wire w_dff_A_OFptFf4R2_0;
	wire w_dff_A_rRRegyjH1_0;
	wire w_dff_A_LHqCxxok4_0;
	wire w_dff_A_ggZuIP4t4_0;
	wire w_dff_A_aEzecLA27_0;
	wire w_dff_A_FZrxiTix6_0;
	wire w_dff_A_jxpmN3le4_2;
	wire w_dff_A_2ievJ18M9_2;
	wire w_dff_A_awc91F4R1_2;
	wire w_dff_B_ueIeBsUt2_1;
	wire w_dff_B_3PWJPcsw6_1;
	wire w_dff_A_bW5mP7gb9_1;
	wire w_dff_A_2FQneTPi2_1;
	wire w_dff_A_HsfrBfd07_1;
	wire w_dff_A_rpRPwpt80_1;
	wire w_dff_A_kkjYvLWy1_2;
	wire w_dff_A_BkSHWRxp6_0;
	wire w_dff_A_D5l59Qyj7_0;
	wire w_dff_A_a8XZ43Js4_1;
	wire w_dff_A_5YLdQIJG0_1;
	wire w_dff_B_WkgTgB8s2_0;
	wire w_dff_B_jj7QTbvu5_0;
	wire w_dff_B_G8YWFHHL2_0;
	wire w_dff_B_X7tN8g4a7_0;
	wire w_dff_B_Q3toTGed4_0;
	wire w_dff_B_RTKBsLD81_0;
	wire w_dff_B_OTbKmBll2_0;
	wire w_dff_B_0strUoqp1_0;
	wire w_dff_B_gHsL6Q9M2_0;
	wire w_dff_B_hAveu1Gn1_0;
	wire w_dff_B_4O5FlavO8_0;
	wire w_dff_B_2iqz4Qca6_0;
	wire w_dff_B_hrPZbIHP1_0;
	wire w_dff_B_1lHDzU4e3_2;
	wire w_dff_B_iSPI2NTX6_2;
	wire w_dff_B_D4nHgDTr3_2;
	wire w_dff_B_SMMNfKzr1_1;
	wire w_dff_B_fqoEoEid8_1;
	wire w_dff_B_u34MmkyJ4_1;
	wire w_dff_B_n9ADeJyW6_1;
	wire w_dff_B_loUnZsCX4_1;
	wire w_dff_B_LGSufPLq9_1;
	wire w_dff_B_aDsq1VDI1_1;
	wire w_dff_B_zJDkO5pI3_1;
	wire w_dff_B_G7gUarwH4_0;
	wire w_dff_B_mBbYEeAf7_0;
	wire w_dff_B_tjkDXg8y1_0;
	wire w_dff_B_ebyXWjon0_1;
	wire w_dff_B_u09SE55u4_1;
	wire w_dff_B_L7NYPyV12_1;
	wire w_dff_B_x4PZrSTy0_1;
	wire w_dff_B_shPkzRl94_1;
	wire w_dff_B_whuvM3Q51_1;
	wire w_dff_B_Q531J5yL6_1;
	wire w_dff_B_oUFeRytN2_1;
	wire w_dff_B_w8b7rGUl0_1;
	wire w_dff_B_EOjIbgGb2_1;
	wire w_dff_B_vS45smQj3_1;
	wire w_dff_B_2qKPxEwx7_1;
	wire w_dff_B_KthAG3j72_1;
	wire w_dff_B_UygP64ca7_1;
	wire w_dff_B_vO0YA87X3_1;
	wire w_dff_A_BkmynQCa8_0;
	wire w_dff_A_L7OWDQXr2_0;
	wire w_dff_A_8dO28ARF5_0;
	wire w_dff_A_6yGPh6Yv3_0;
	wire w_dff_A_QodupDsy5_0;
	wire w_dff_B_6pT1L4yy1_1;
	wire w_dff_B_6bDH561l7_1;
	wire w_dff_B_kbMravUl7_1;
	wire w_dff_B_gzn3ppYX3_1;
	wire w_dff_B_L5gyn8Za0_0;
	wire w_dff_B_ofQbNUbt5_0;
	wire w_dff_B_XBsHMG8d2_0;
	wire w_dff_B_qHGkKn6b1_0;
	wire w_dff_B_NPBVLA1n1_0;
	wire w_dff_B_r5x4ks831_0;
	wire w_dff_B_n4OzFfxW7_0;
	wire w_dff_B_RXu676aU5_0;
	wire w_dff_B_ykUVoXwi4_0;
	wire w_dff_B_AmiUrmva0_0;
	wire w_dff_B_l9L4pKaY8_0;
	wire w_dff_B_JJ9BEM7M2_0;
	wire w_dff_B_yHemKvBF0_0;
	wire w_dff_B_zBKxwZd23_0;
	wire w_dff_B_TqW49frs3_2;
	wire w_dff_B_jiFN7tWL0_2;
	wire w_dff_B_dil3UexK9_2;
	wire w_dff_B_enXgUU5g4_1;
	wire w_dff_B_sF91ZaHz1_1;
	wire w_dff_B_KuakVzVa2_1;
	wire w_dff_B_Kp0eYmnF7_1;
	wire w_dff_B_AbMsTt9T4_1;
	wire w_dff_B_feve4orU4_1;
	wire w_dff_B_vzEfQoki3_1;
	wire w_dff_B_EMjRTHoL2_1;
	wire w_dff_B_5HsUXeEf0_0;
	wire w_dff_B_yefxkvvk1_0;
	wire w_dff_B_u4BizK8s4_0;
	wire w_dff_B_fte8Gnki9_0;
	wire w_dff_B_4tWlY9bq3_1;
	wire w_dff_B_Icuqqmhk5_1;
	wire w_dff_A_ToPV5wHw3_2;
	wire w_dff_A_2Ag8oVJY1_2;
	wire w_dff_A_sXs48mAJ2_2;
	wire w_dff_A_pkrpol0q8_0;
	wire w_dff_A_Rc4alZ5s4_0;
	wire w_dff_A_nZHAwGjk1_0;
	wire w_dff_A_1awNcfCx8_0;
	wire w_dff_A_UqfCelNO3_0;
	wire w_dff_A_hjTmyCYm9_1;
	wire w_dff_A_Q826vMP53_2;
	wire w_dff_A_1d6GvdyF2_2;
	wire w_dff_B_JKC03qpZ6_1;
	wire w_dff_B_I2URrG8P0_1;
	wire w_dff_A_Xf4DBYUo9_0;
	wire w_dff_A_KBPGaox53_0;
	wire w_dff_A_7kP6WV9w4_1;
	wire w_dff_B_fDChoKtb0_1;
	wire w_dff_B_x5qi5khF1_1;
	wire w_dff_B_GJS68R1O6_1;
	wire w_dff_B_iKAp5iwP1_1;
	wire w_dff_B_ltgUwjIp9_1;
	wire w_dff_B_rbnADBru1_1;
	wire w_dff_B_ATgaZu0P8_1;
	wire w_dff_B_o9FCPZlq3_1;
	wire w_dff_B_lXbCqQiA8_1;
	wire w_dff_B_3xas6Zzu6_0;
	wire w_dff_B_qP4G1cQn3_0;
	wire w_dff_B_hqjbsfWB2_0;
	wire w_dff_B_XFTdOrUM3_0;
	wire w_dff_B_h26Tk7ao5_0;
	wire w_dff_B_YwyUonoH8_0;
	wire w_dff_B_xP1DKWMQ0_1;
	wire w_dff_A_YBRV6JoW0_0;
	wire w_dff_A_wmEkHaAt4_1;
	wire w_dff_A_sGjd8nTr1_0;
	wire w_dff_A_K6riXqK07_2;
	wire w_dff_A_aIHJe3SX5_1;
	wire w_dff_A_fsG94DFF4_2;
	wire w_dff_A_Q8gasQY60_0;
	wire w_dff_A_oo1MVGZV9_0;
	wire w_dff_A_n4GJO1j45_0;
	wire w_dff_A_Vg2LN1cI2_0;
	wire w_dff_A_4YVVfOtG6_0;
	wire w_dff_A_d0YTLvCK5_0;
	wire w_dff_A_hFWOoDh04_0;
	wire w_dff_A_dG2T47mw8_1;
	wire w_dff_A_butyZvEC9_1;
	wire w_dff_A_NhU4K2DY7_2;
	wire w_dff_A_rAsnwgLK2_2;
	wire w_dff_A_wmGJVR450_2;
	wire w_dff_A_edRtoikW4_2;
	wire w_dff_A_wBk3dmqZ4_2;
	wire w_dff_B_6WPuEnl14_3;
	wire w_dff_B_CabbYQKU6_3;
	wire w_dff_A_3t32s8AQ0_0;
	wire w_dff_A_2vAXRqdl8_0;
	wire w_dff_A_KdetSORu4_0;
	wire w_dff_A_wEzJNpno8_0;
	wire w_dff_A_Bi8XuIGL9_2;
	wire w_dff_A_NzwxeOLa6_2;
	wire w_dff_A_ZzP2sz4o8_2;
	wire w_dff_B_UQ6NEMru6_1;
	wire w_dff_B_0QuqJQqF4_1;
	wire w_dff_B_q6jkLf9D4_1;
	wire w_dff_B_gvWWt8179_1;
	wire w_dff_B_HCVvmeyx9_1;
	wire w_dff_B_Towb3JhV2_1;
	wire w_dff_B_DvYmC1dl7_1;
	wire w_dff_B_X4A99RoH5_1;
	wire w_dff_B_JmXHJZjB7_1;
	wire w_dff_B_iZKQKn2k8_1;
	wire w_dff_B_dlWD6ODR7_1;
	wire w_dff_B_mPyDFJ913_1;
	wire w_dff_B_p2ZINNA54_1;
	wire w_dff_B_G3tm66WX3_1;
	wire w_dff_B_hH16Nipb3_1;
	wire w_dff_B_qmmAf7A57_1;
	wire w_dff_B_DjZx3B481_1;
	wire w_dff_B_JpgqzGnk3_1;
	wire w_dff_B_xmQ7M9xF6_1;
	wire w_dff_B_Ivd7VMH57_1;
	wire w_dff_B_XhjxZbDM4_1;
	wire w_dff_B_6mQgSj0s0_1;
	wire w_dff_B_Jc6CjSTS4_1;
	wire w_dff_B_ZqqnOma20_1;
	wire w_dff_B_YH5U34AS3_1;
	wire w_dff_B_QU4SmOqC5_1;
	wire w_dff_B_8DMwpq5A1_1;
	wire w_dff_B_AS9Mmiq39_1;
	wire w_dff_B_WW3sFcDx4_1;
	wire w_dff_B_Pzz3Wyd36_1;
	wire w_dff_B_dIuZ8OO31_0;
	wire w_dff_B_KFEIgUKM1_0;
	wire w_dff_B_fj5SL7Wz5_0;
	wire w_dff_B_Noki1fYK8_0;
	wire w_dff_B_snpjvWNa3_0;
	wire w_dff_B_p2Syoab75_0;
	wire w_dff_B_82ZWVWhY8_0;
	wire w_dff_B_f4vuB5h31_0;
	wire w_dff_B_yqVOazlv2_0;
	wire w_dff_B_32nEx41T3_0;
	wire w_dff_B_aCFUkeCV3_0;
	wire w_dff_B_Dm3ZAoIg6_0;
	wire w_dff_B_IdJBzlcj5_0;
	wire w_dff_B_yVH7W18P1_0;
	wire w_dff_B_VC63psti9_0;
	wire w_dff_B_2fXFua545_0;
	wire w_dff_B_YBD5ZGiK7_1;
	wire w_dff_B_ueT7NGUG0_1;
	wire w_dff_B_twTMpFZ06_1;
	wire w_dff_B_n8RVwXTT6_1;
	wire w_dff_B_d8bkvUs89_1;
	wire w_dff_B_q9dJCnUC4_1;
	wire w_dff_B_AsmfxMTM7_1;
	wire w_dff_B_MPqOTiqy8_1;
	wire w_dff_B_oO0itrCv6_1;
	wire w_dff_A_frpBbFp05_0;
	wire w_dff_A_aitynTe77_0;
	wire w_dff_A_LVeLffIQ7_0;
	wire w_dff_A_aaGYHJJX7_0;
	wire w_dff_A_sXkJnJh31_0;
	wire w_dff_A_W9KmvIw12_0;
	wire w_dff_A_Ed2tEucy6_0;
	wire w_dff_A_IYpiv8BJ8_0;
	wire w_dff_A_JJOQs7Wi4_0;
	wire w_dff_A_RqAIpejz8_0;
	wire w_dff_A_64TXrpuB7_0;
	wire w_dff_B_OOPdKPrC6_2;
	wire w_dff_B_Y02DkMOs8_2;
	wire w_dff_B_BP0FHnd11_2;
	wire w_dff_B_QLVd4Pmh4_2;
	wire w_dff_B_504jPPon2_2;
	wire w_dff_A_5vksmMD30_0;
	wire w_dff_A_KNKfWtxB6_1;
	wire w_dff_A_tCh7tCAi7_2;
	wire w_dff_A_dKM9fRZC2_2;
	wire w_dff_A_w6FAsZmD5_2;
	wire w_dff_A_HSDjMAYL4_2;
	wire w_dff_A_KHTTcMNu5_0;
	wire w_dff_A_oPjllWo38_0;
	wire w_dff_A_EcjYyVXo1_0;
	wire w_dff_A_fTJeBMfM6_0;
	wire w_dff_A_1kcaw7ez7_0;
	wire w_dff_A_DnJ5DBzF1_0;
	wire w_dff_A_faTBR8PZ7_0;
	wire w_dff_A_aqGYU6qh7_0;
	wire w_dff_A_hF4QMVNa8_0;
	wire w_dff_A_EMneLXFc6_0;
	wire w_dff_A_5GDr8oCN8_0;
	wire w_dff_B_3ZtdagPq9_1;
	wire w_dff_B_u0WOS3Pc4_1;
	wire w_dff_B_V53cg0X02_1;
	wire w_dff_B_K8TahF035_1;
	wire w_dff_B_btmOODy13_1;
	wire w_dff_B_qEQQpsKk5_0;
	wire w_dff_B_r9MmtNCY7_0;
	wire w_dff_B_MS3xUnKy5_0;
	wire w_dff_B_xC81aw5z5_0;
	wire w_dff_B_eh53O0zL0_0;
	wire w_dff_A_PcpneghQ7_0;
	wire w_dff_A_2cTOs3ML8_0;
	wire w_dff_B_T9BYHnEv1_0;
	wire w_dff_B_6lPqW0NK3_1;
	wire w_dff_B_TJmzSrc90_1;
	wire w_dff_B_odN55ZPf6_1;
	wire w_dff_B_z8WZTYfZ4_0;
	wire w_dff_B_qe1eSGki3_1;
	wire w_dff_B_lJIOTZQH6_0;
	wire w_dff_B_4gwmfbNS1_1;
	wire w_dff_B_uu6sxKaR8_1;
	wire w_dff_B_7wKi2Shd7_1;
	wire w_dff_B_RV9gjbcG5_0;
	wire w_dff_B_FcX5Hktv6_0;
	wire w_dff_B_2ri51vPv3_0;
	wire w_dff_B_GktndBhK1_0;
	wire w_dff_B_fJLKRzUl4_1;
	wire w_dff_A_lNYH5L6n4_0;
	wire w_dff_A_mwcxET8O5_0;
	wire w_dff_A_yPcGyAXE4_0;
	wire w_dff_A_h3X8GGaS8_0;
	wire w_dff_B_L0gb3Hkz2_1;
	wire w_dff_B_yyP4thTY9_1;
	wire w_dff_B_S0xTrdX29_1;
	wire w_dff_B_da3s2Xhl4_1;
	wire w_dff_B_LYANNG6m0_1;
	wire w_dff_B_cS5Q11L10_1;
	wire w_dff_B_eeGo6B2W3_1;
	wire w_dff_B_GjL4teN95_1;
	wire w_dff_B_zTLMdmw39_1;
	wire w_dff_B_9ra4wDRl9_1;
	wire w_dff_B_Fh2gQ6be0_1;
	wire w_dff_B_Juy0Tt2p6_1;
	wire w_dff_B_PWnJhhAO2_1;
	wire w_dff_B_vRy6dq1h5_1;
	wire w_dff_B_vSFtWIEC2_1;
	wire w_dff_B_1g47Foue8_1;
	wire w_dff_B_kAndRELX8_1;
	wire w_dff_B_6EBdFV0W8_1;
	wire w_dff_B_ziHDoDNs1_1;
	wire w_dff_B_xPNZux7h1_1;
	wire w_dff_B_X36jGgTQ2_1;
	wire w_dff_B_QrhlCgfN8_1;
	wire w_dff_B_eBNDRAH97_1;
	wire w_dff_B_Oa4FPMrk7_1;
	wire w_dff_B_yXaaSN0r9_1;
	wire w_dff_B_EllftlNr1_1;
	wire w_dff_A_E29owVpO8_2;
	wire w_dff_A_fLvleYC64_2;
	wire w_dff_A_4caMF2zU4_2;
	wire w_dff_A_vf3Gj3wd1_2;
	wire w_dff_A_jkbpH5wQ5_2;
	wire w_dff_A_KDIgANww9_2;
	wire w_dff_A_RyklNXlN7_2;
	wire w_dff_A_oOfK8kwV9_2;
	wire w_dff_A_9shosCWL7_2;
	wire w_dff_A_s4vdH9qE5_2;
	wire w_dff_A_KgpDjXJt6_2;
	wire w_dff_A_dlwQqz3t3_2;
	wire w_dff_A_eJ7z3tGy4_2;
	wire w_dff_A_VsuE2nZs8_2;
	wire w_dff_A_C4BKBJs97_2;
	wire w_dff_A_AlozjURd2_2;
	wire w_dff_A_r60OqSVx4_2;
	wire w_dff_A_VMaU69V91_2;
	wire w_dff_A_aPSaX0Ac6_2;
	wire w_dff_A_4OA7GnSW0_2;
	wire w_dff_A_s9qkZEY39_2;
	wire w_dff_A_N0O1RP3f7_2;
	wire w_dff_A_6l7D93C82_2;
	wire w_dff_A_VDxF2ZcP8_2;
	wire w_dff_A_Uy0iffnN3_2;
	wire w_dff_B_ZRoBCCT49_0;
	wire w_dff_B_fmSecLm54_0;
	wire w_dff_B_zgNCQm5D1_0;
	wire w_dff_B_FHmxkujZ1_0;
	wire w_dff_B_amlKhovH2_0;
	wire w_dff_B_ccDsk3zu6_0;
	wire w_dff_B_hn76hPMW8_0;
	wire w_dff_B_0HX4qyA17_0;
	wire w_dff_B_wbCmYHaw6_0;
	wire w_dff_B_BObX65gH8_0;
	wire w_dff_B_Rv7rYFht8_0;
	wire w_dff_B_4eeXoA0X8_0;
	wire w_dff_B_OA0MvQRM5_0;
	wire w_dff_B_qvNlr5RR8_0;
	wire w_dff_B_CGoMiKOQ9_0;
	wire w_dff_B_YEdl7OfL6_0;
	wire w_dff_B_yp8qlzjU5_0;
	wire w_dff_B_YQtkHUAk7_0;
	wire w_dff_B_Z9IXGwA60_0;
	wire w_dff_B_ipqgx8Tu0_0;
	wire w_dff_B_Oc5FpvzU5_0;
	wire w_dff_B_613TrTLX7_2;
	wire w_dff_B_fVB9cpGC4_1;
	wire w_dff_B_5kW2X1Jt1_1;
	wire w_dff_A_vmu3grkC7_0;
	wire w_dff_A_P0qOsKlY4_0;
	wire w_dff_A_DXKRFzAL8_0;
	wire w_dff_A_CyFPFsgZ5_0;
	wire w_dff_A_Ak71Hu3n0_0;
	wire w_dff_A_1cpvF5ce9_0;
	wire w_dff_A_mWPLGSTW8_0;
	wire w_dff_A_LYZ5Ozx56_0;
	wire w_dff_A_N8kS113w0_0;
	wire w_dff_A_Tz8aNJD11_0;
	wire w_dff_A_msNELFM06_0;
	wire w_dff_A_gYhWE2PL5_0;
	wire w_dff_A_ZOR8hdyJ7_0;
	wire w_dff_A_swTQvqRQ1_0;
	wire w_dff_A_UMTYZDQ84_0;
	wire w_dff_A_8dg1W2673_0;
	wire w_dff_A_3nVv4tEd8_0;
	wire w_dff_A_eiblXQ9W4_0;
	wire w_dff_A_Klmtffqm4_0;
	wire w_dff_A_e2azE1u77_0;
	wire w_dff_A_ilKoLCXX7_2;
	wire w_dff_A_j9wGIjuJ3_2;
	wire w_dff_A_iv4jWVui0_2;
	wire w_dff_A_slBwO6yM4_2;
	wire w_dff_A_m865teEJ0_2;
	wire w_dff_A_cCAvu9o55_2;
	wire w_dff_A_vz4vnveJ1_2;
	wire w_dff_A_ndDbO4cl5_2;
	wire w_dff_A_hPePvWMc1_2;
	wire w_dff_A_PBISrbJt7_2;
	wire w_dff_A_yraG014I1_2;
	wire w_dff_A_VTL4K4AN2_0;
	wire w_dff_A_cZycAh8e0_0;
	wire w_dff_A_L2OUdAyE3_0;
	wire w_dff_A_FHyPy2w78_0;
	wire w_dff_A_H9OFNDI03_0;
	wire w_dff_A_6p5mLKqQ5_0;
	wire w_dff_A_XMqXqIrL6_0;
	wire w_dff_A_hIqNW8aG6_0;
	wire w_dff_A_OH0nMXVi0_0;
	wire w_dff_A_YKE7TXah8_0;
	wire w_dff_A_mRTnXCtn3_0;
	wire w_dff_A_NUax58OZ8_0;
	wire w_dff_A_IXgFBrHy9_0;
	wire w_dff_A_ykhlCQX31_0;
	wire w_dff_A_5aeUg1Co1_0;
	wire w_dff_A_Yd56h4Yw5_0;
	wire w_dff_A_A0EatiEj7_0;
	wire w_dff_A_2gT5xT5g5_0;
	wire w_dff_A_rqTnFF352_0;
	wire w_dff_A_DnGrOMJs5_0;
	wire w_dff_A_mZPRQKzC3_2;
	wire w_dff_A_uDSmtvhE7_2;
	wire w_dff_A_0rz0RcBA5_2;
	wire w_dff_A_WwdrCMyo0_2;
	wire w_dff_A_P5KRAUwM4_2;
	wire w_dff_A_AV0x3rVB6_2;
	wire w_dff_A_uQ4ODTvv1_2;
	wire w_dff_A_zep5KxRb6_2;
	wire w_dff_A_ldWFV7vf9_2;
	wire w_dff_A_NZMNoHdR2_2;
	wire w_dff_A_m3suCFgq3_2;
	wire w_dff_A_n8vnFEGM9_2;
	wire w_dff_A_5gIW36ZP4_2;
	wire w_dff_A_wDrieCip9_2;
	wire w_dff_B_26vXIsBq6_0;
	wire w_dff_B_237LmwaP1_0;
	wire w_dff_B_HYqnMS4b3_0;
	wire w_dff_B_KIlfmhqN7_0;
	wire w_dff_B_b0aBPuSw9_0;
	wire w_dff_B_Q9E1as2H0_0;
	wire w_dff_B_melxdjnz5_0;
	wire w_dff_B_NvLChvnn6_0;
	wire w_dff_B_X4ZlOaTY1_0;
	wire w_dff_B_tybX5DEv3_0;
	wire w_dff_B_DqusuIoh6_0;
	wire w_dff_B_by69jzI17_0;
	wire w_dff_B_nvGFCjNw2_0;
	wire w_dff_B_OVYSqZTJ5_0;
	wire w_dff_B_JVYlG0v43_0;
	wire w_dff_B_4vBj07Vh5_0;
	wire w_dff_B_2YsL8ecb2_0;
	wire w_dff_B_XRI0FZX86_0;
	wire w_dff_B_0mBTJR4Q8_0;
	wire w_dff_B_ucBX0RAq0_0;
	wire w_dff_B_Kldu5qHO6_1;
	wire w_dff_B_gocFImUT3_1;
	wire w_dff_A_fW0wnGPG7_1;
	wire w_dff_A_c2JOarfZ8_1;
	wire w_dff_A_f4wIRi5n4_1;
	wire w_dff_A_G7U2y4mg0_1;
	wire w_dff_A_eb5TBan76_1;
	wire w_dff_A_NaHnANhF3_1;
	wire w_dff_A_AEMtDXUi3_1;
	wire w_dff_A_CfQ9ro8Z8_1;
	wire w_dff_A_Kdko3opX3_1;
	wire w_dff_A_JaJAejEe3_1;
	wire w_dff_A_OHDH7wRu3_1;
	wire w_dff_A_Kx6c7k823_1;
	wire w_dff_A_Epcwrcqr2_1;
	wire w_dff_A_gnIEyZ3w4_1;
	wire w_dff_A_FQO6eSNF1_1;
	wire w_dff_A_4eWSPZKd2_1;
	wire w_dff_A_H6tcGR0p0_1;
	wire w_dff_A_Bc2Y3kNT6_1;
	wire w_dff_A_bxqxQOu92_1;
	wire w_dff_A_qr1zaZfW9_1;
	wire w_dff_A_ouVm1GKL6_1;
	wire w_dff_A_Ddie4o278_1;
	wire w_dff_A_WnITRA3p3_1;
	wire w_dff_A_96QPoJ9O4_1;
	wire w_dff_A_6HbkPmG85_1;
	wire w_dff_A_zhxWjCru4_1;
	wire w_dff_A_y4arpHE37_1;
	wire w_dff_A_QlFPTUxj5_1;
	wire w_dff_A_WIEMXsFY3_1;
	wire w_dff_A_pDA50E2E5_1;
	wire w_dff_A_8AnJhNNe4_1;
	wire w_dff_A_ReZifjbl4_1;
	wire w_dff_A_d5Cz99bG2_1;
	wire w_dff_A_9ZZjS1ph8_1;
	wire w_dff_A_lH7F1bdL0_1;
	wire w_dff_A_oOFGgjiW7_1;
	wire w_dff_A_nrZt1lOM6_1;
	wire w_dff_A_cNzuEArp5_1;
	wire w_dff_B_7UjudSZW9_0;
	wire w_dff_B_DcadDWTU5_0;
	wire w_dff_B_gX3TpLfj4_0;
	wire w_dff_B_Vo5jpYLr7_0;
	wire w_dff_B_tOna3Ym00_0;
	wire w_dff_B_tgNBYLqh4_0;
	wire w_dff_B_7yaZaOhd8_0;
	wire w_dff_B_4vDqfosu3_0;
	wire w_dff_B_mOLvacjo2_0;
	wire w_dff_B_2PpFbc1B8_0;
	wire w_dff_B_WE21cq7c4_0;
	wire w_dff_B_VflmCJ1O8_0;
	wire w_dff_B_t6KdXIAc2_0;
	wire w_dff_B_Ea27ydjA8_0;
	wire w_dff_B_8mtSHyKK6_0;
	wire w_dff_B_VT34JV8y1_0;
	wire w_dff_B_oZPXF36v3_0;
	wire w_dff_B_8pkK5WnP2_0;
	wire w_dff_B_4ZDBi9CO4_0;
	wire w_dff_B_ckn15Wxm8_0;
	wire w_dff_B_0D6r4phK0_1;
	wire w_dff_A_F6kEEoLb0_2;
	wire w_dff_B_vp73fETp6_0;
	wire w_dff_B_tLVzxb7o8_0;
	wire w_dff_B_LnGzdbko1_0;
	wire w_dff_B_OJeBpcXP6_0;
	wire w_dff_B_ndmMawgf5_0;
	wire w_dff_B_5LIcaxSZ6_0;
	wire w_dff_B_vjChEcSU9_0;
	wire w_dff_B_9LRB2zkL8_0;
	wire w_dff_B_pGcqzuNM2_0;
	wire w_dff_B_CPZiW7jH9_0;
	wire w_dff_B_lcrO5USL6_0;
	wire w_dff_B_drPAWo4y3_0;
	wire w_dff_B_uZW28TeO5_0;
	wire w_dff_B_L9wP2SIE6_0;
	wire w_dff_B_6B1BSFVf9_0;
	wire w_dff_B_8LweTrcT8_0;
	wire w_dff_B_zpWxDfUm7_0;
	wire w_dff_B_ovcS07R84_0;
	wire w_dff_B_ZPD2HFVt2_0;
	wire w_dff_B_gnu0io0Y0_1;
	wire w_dff_B_Mguj03XS6_1;
	wire w_dff_B_Y0iBS1MF6_1;
	wire w_dff_A_c8Kmh86T8_0;
	wire w_dff_A_mcKseCPZ0_0;
	wire w_dff_A_gzFjyGFk8_0;
	wire w_dff_A_aTbMuSXF5_0;
	wire w_dff_A_dkModUv92_0;
	wire w_dff_A_mmi0TJ2l1_0;
	wire w_dff_A_ZzFSyu8U7_0;
	wire w_dff_A_xJs2sFMc6_0;
	wire w_dff_A_6TiupRoT3_0;
	wire w_dff_A_hP8Luy1H1_0;
	wire w_dff_A_WTS0IMSz4_0;
	wire w_dff_A_t9DcpFOp2_0;
	wire w_dff_A_4fcaJOul6_0;
	wire w_dff_A_yxrj8M9C6_0;
	wire w_dff_A_JQAb2F3x3_0;
	wire w_dff_A_OE3fPINj8_0;
	wire w_dff_A_D21QqSyu6_0;
	wire w_dff_A_0PAbTmFU7_0;
	wire w_dff_A_l5VQZLGs8_2;
	wire w_dff_A_Wi8FS5Qf4_2;
	wire w_dff_A_MgFTMBNo6_2;
	wire w_dff_A_Zw79KdCA2_2;
	wire w_dff_A_gMiMV8FR9_2;
	wire w_dff_A_ix6r8cx42_2;
	wire w_dff_A_8RyrBXgn9_2;
	wire w_dff_A_4KYwUy5x1_2;
	wire w_dff_A_Dmet1Hgc7_2;
	wire w_dff_A_MAyHAZ0z1_2;
	wire w_dff_A_b185gkc21_2;
	wire w_dff_A_aTCTlvJy2_2;
	wire w_dff_A_2RMoAcWF9_2;
	wire w_dff_A_PiGyPitN2_2;
	wire w_dff_A_MHh1cXZs6_2;
	wire w_dff_A_l4R2yFE22_2;
	wire w_dff_A_PJVQDKlL0_2;
	wire w_dff_A_C4ifFUPk4_2;
	wire w_dff_A_qOvYg6Ov9_2;
	wire w_dff_A_qESsbqie3_0;
	wire w_dff_A_YJTwBiIT3_0;
	wire w_dff_A_a3otgkqM4_0;
	wire w_dff_A_fL0tGpx44_0;
	wire w_dff_A_Q93y5Iik5_0;
	wire w_dff_A_45hqZKf57_0;
	wire w_dff_A_dQRPsQqf2_0;
	wire w_dff_A_OEbN8EXk5_0;
	wire w_dff_A_DRJflWKr9_0;
	wire w_dff_A_gSLcyW3V2_0;
	wire w_dff_A_Z3HRJwEi0_0;
	wire w_dff_A_M5wqTL3w1_0;
	wire w_dff_A_HyEHA1b12_0;
	wire w_dff_A_z966KQDq9_0;
	wire w_dff_A_Fa0uN8os5_0;
	wire w_dff_A_vH4D8Mmr4_0;
	wire w_dff_A_n56Cg8U79_0;
	wire w_dff_A_g60qJbka0_2;
	wire w_dff_A_Z7AbxlRT4_2;
	wire w_dff_A_sLlhvxc51_2;
	wire w_dff_A_nTKTtuIH6_2;
	wire w_dff_A_1LACJbbj5_2;
	wire w_dff_A_tGuooKm99_2;
	wire w_dff_A_HMeDhRlP1_2;
	wire w_dff_A_Z9An5mDf6_2;
	wire w_dff_A_nwo6rMuK4_2;
	wire w_dff_A_GIRc0fds5_2;
	wire w_dff_A_WNH877zU8_2;
	wire w_dff_A_LkUCL5xp3_2;
	wire w_dff_A_CotZHC4G3_2;
	wire w_dff_A_ubrXqq9h7_2;
	wire w_dff_A_h6ODVTHe3_2;
	wire w_dff_A_Rkj2NQzS1_2;
	wire w_dff_A_y4MCU1Or5_2;
	wire w_dff_A_OGv8jIoD3_2;
	wire w_dff_A_GLLu1T570_2;
	wire w_dff_A_3MTawk6p2_2;
	wire w_dff_B_sLQnThb07_0;
	wire w_dff_B_FpPR17FD1_0;
	wire w_dff_B_fDzXJuTr2_0;
	wire w_dff_B_clEgHPOm1_0;
	wire w_dff_B_huIMoZ791_0;
	wire w_dff_B_4T6hSof15_0;
	wire w_dff_B_mP2gaJKY6_0;
	wire w_dff_B_ZFDINmTe2_0;
	wire w_dff_B_2f4Odfvv7_0;
	wire w_dff_B_1MX9Kp512_0;
	wire w_dff_B_DzZl1J0C9_0;
	wire w_dff_B_uLmsER0w4_0;
	wire w_dff_B_HB9Uenv55_0;
	wire w_dff_B_0GPm6Bc90_0;
	wire w_dff_B_99IbGpKN5_0;
	wire w_dff_B_5cShaHcV2_0;
	wire w_dff_B_679P78Q55_0;
	wire w_dff_B_5zcaT43A4_0;
	wire w_dff_B_k5gzeLve0_0;
	wire w_dff_B_sS6HhTvr8_0;
	wire w_dff_B_BpkAsc1y6_2;
	wire w_dff_B_tnKmZ8XB9_1;
	wire w_dff_B_Xq6EIfTl7_1;
	wire w_dff_A_YwCVStrG5_1;
	wire w_dff_A_iqM4HQ2X9_1;
	wire w_dff_A_3sqNHz3t1_1;
	wire w_dff_A_CbzZsDXQ2_1;
	wire w_dff_A_eaVJy22C3_1;
	wire w_dff_A_iQS3qMlv3_1;
	wire w_dff_A_W1kud2fI7_1;
	wire w_dff_A_F0ZOs3nt1_1;
	wire w_dff_A_8V78MCKm0_1;
	wire w_dff_A_R51gQHhk2_1;
	wire w_dff_A_UIZHmYXx2_1;
	wire w_dff_A_QISS2oXA3_1;
	wire w_dff_A_tBzkUQdT8_1;
	wire w_dff_A_UBf3TArc6_1;
	wire w_dff_A_5h51zdDZ3_1;
	wire w_dff_A_6Lp0Fj9l6_1;
	wire w_dff_A_dzJ10lsn6_1;
	wire w_dff_A_DPVYKORw1_1;
	wire w_dff_A_bn9BiymC4_1;
	wire w_dff_A_d0PDyUJm9_2;
	wire w_dff_A_y2a2Dp8J0_2;
	wire w_dff_A_LAJorAAD2_2;
	wire w_dff_A_vew6i1Ws8_2;
	wire w_dff_A_nsPb19gP9_2;
	wire w_dff_A_DvmywXrd9_2;
	wire w_dff_A_qoXdwmNy8_2;
	wire w_dff_A_CISUJWI08_2;
	wire w_dff_A_LUfgd2Hd7_2;
	wire w_dff_A_dEneHv9m8_2;
	wire w_dff_A_i0Yk1vAb5_2;
	wire w_dff_A_1rX1K71I0_2;
	wire w_dff_A_LrGycIDG9_2;
	wire w_dff_A_Snd94FQK2_2;
	wire w_dff_A_om8VqVgx9_2;
	wire w_dff_A_Az5eyil72_2;
	wire w_dff_A_Js4HmcVz2_2;
	wire w_dff_A_Q2nWyxKH7_2;
	wire w_dff_A_3Je4OfGt1_2;
	wire w_dff_A_l7yjVuJE0_2;
	wire w_dff_A_YoMJhFeU5_1;
	wire w_dff_A_udvKaqGj0_1;
	wire w_dff_A_gD303vOn0_1;
	wire w_dff_A_wB0nvP2l9_1;
	wire w_dff_A_qDASnoKV9_1;
	wire w_dff_A_qvhKjY1a3_1;
	wire w_dff_A_xvay0Dri8_1;
	wire w_dff_A_Gzin9HnS2_1;
	wire w_dff_A_BzPsx90L0_1;
	wire w_dff_A_jFyLk3b71_1;
	wire w_dff_A_7aNaPJP95_1;
	wire w_dff_A_SnlfO4Ny4_1;
	wire w_dff_A_Wxc2EWao9_1;
	wire w_dff_A_vl56YY354_1;
	wire w_dff_A_yFPcyPHm1_1;
	wire w_dff_A_E9Ao7VvB8_1;
	wire w_dff_A_gocVw8n22_1;
	wire w_dff_A_epruyMLi0_1;
	wire w_dff_A_AZUk2N372_1;
	wire w_dff_A_sSo3SwRo0_2;
	wire w_dff_A_9qiF0ob89_2;
	wire w_dff_A_G5sR4Sco4_2;
	wire w_dff_A_Oedmlh5m1_2;
	wire w_dff_A_7kD2yT968_2;
	wire w_dff_A_hbjkuKhH9_2;
	wire w_dff_A_1avGh9X24_2;
	wire w_dff_A_q9DS2HfD8_2;
	wire w_dff_A_KSBaIyKx3_2;
	wire w_dff_A_00t9mj1C0_2;
	wire w_dff_A_nr47YXuu8_2;
	wire w_dff_A_IRWHGHsC2_2;
	wire w_dff_A_2HsNTUVT5_2;
	wire w_dff_A_hZw2nYKR1_2;
	wire w_dff_A_ePxzCj0Z4_2;
	wire w_dff_A_0Z7jcUqa5_2;
	wire w_dff_A_SwmEI5h61_2;
	wire w_dff_A_EzcBz4r93_2;
	wire w_dff_A_hoBTjbXv9_2;
	wire w_dff_A_4PPCRYOm0_2;
	wire w_dff_B_YIHEzFLr0_0;
	wire w_dff_B_jdUK9P8A4_0;
	wire w_dff_B_8VbUnEOV0_0;
	wire w_dff_B_g9gjqgJv5_0;
	wire w_dff_B_iI5WRS1v9_0;
	wire w_dff_B_6JDFyqZo5_0;
	wire w_dff_B_GlVtUsFp6_0;
	wire w_dff_B_8ahMyhzz3_0;
	wire w_dff_B_mksuzE8m9_0;
	wire w_dff_B_nqkE2MRd7_0;
	wire w_dff_B_1xVD6u4R2_0;
	wire w_dff_B_MjtRJtDF1_0;
	wire w_dff_B_ryiqz1h99_0;
	wire w_dff_B_HP1w4vLn7_0;
	wire w_dff_B_sO7Fx42m4_0;
	wire w_dff_B_M9Muah9E5_0;
	wire w_dff_B_af4HBjBw3_0;
	wire w_dff_B_28uQhLBD8_0;
	wire w_dff_B_O2kpaOd25_0;
	wire w_dff_B_KRwNmUJd6_0;
	wire w_dff_A_uRkmLDwz7_2;
	wire w_dff_B_BGVVzNqh7_2;
	wire w_dff_B_VwyDH8wE1_1;
	wire w_dff_B_XOjiSMhh1_0;
	wire w_dff_B_Z8tTqNO08_0;
	wire w_dff_B_EPscGlBm4_0;
	wire w_dff_B_ZSuExcoD5_0;
	wire w_dff_B_Z9FwUdeg9_0;
	wire w_dff_B_rxgoapfK8_0;
	wire w_dff_B_cg5CIlMC6_0;
	wire w_dff_B_9CDAg0i09_0;
	wire w_dff_B_ko5wrpcG1_0;
	wire w_dff_B_eL2xxCXb3_0;
	wire w_dff_B_TdetwKw54_0;
	wire w_dff_B_it33mLoO2_0;
	wire w_dff_B_CgJk59Z23_0;
	wire w_dff_B_DiUfPGgd6_0;
	wire w_dff_B_zJalZ0Rc6_0;
	wire w_dff_B_2Qzm5fIQ3_0;
	wire w_dff_B_SZYu7Suh5_0;
	wire w_dff_B_P9BQJHRS3_0;
	wire w_dff_B_ZMLXcoSU6_0;
	wire w_dff_B_t85foF892_2;
	wire w_dff_B_SitaWkjy3_1;
	wire w_dff_B_hOIKizSm7_1;
	wire w_dff_B_ZdDAzTRd3_1;
	wire w_dff_A_by2ZWpO37_0;
	wire w_dff_A_ie0b4jAk4_0;
	wire w_dff_A_esGKByTC7_0;
	wire w_dff_A_hZs1WtX98_0;
	wire w_dff_A_K1Rw60c30_0;
	wire w_dff_A_VF7lNyY25_0;
	wire w_dff_A_ILcIecHr3_0;
	wire w_dff_A_mQIQYFXF7_0;
	wire w_dff_A_ahNcR6lG6_0;
	wire w_dff_A_2ayUgYl83_0;
	wire w_dff_A_8yTjE47g1_0;
	wire w_dff_A_a3TyolLG8_0;
	wire w_dff_A_c4RUVjH83_0;
	wire w_dff_A_TaHuFmQ14_0;
	wire w_dff_A_T8Pmqg4G4_0;
	wire w_dff_A_KvoQN0Ve8_0;
	wire w_dff_A_LGZ0akvm4_0;
	wire w_dff_A_fxyaCb5N2_0;
	wire w_dff_A_XbjMvyRI0_2;
	wire w_dff_A_T2bA6jRM9_2;
	wire w_dff_A_AKOBf5E62_2;
	wire w_dff_A_y8fZEZoG9_2;
	wire w_dff_A_8l70AWw09_2;
	wire w_dff_A_8yeNDHZb9_2;
	wire w_dff_A_pTbMdTeW4_2;
	wire w_dff_A_DTl5ZaCh6_2;
	wire w_dff_A_niERBPN88_2;
	wire w_dff_A_sHfpWgE41_2;
	wire w_dff_A_U0dCrpGY6_2;
	wire w_dff_A_y4Ho3ifi1_2;
	wire w_dff_A_olHhnR640_2;
	wire w_dff_A_wq7z9bw63_2;
	wire w_dff_A_jYAnm2Ef5_2;
	wire w_dff_A_idF6996p9_2;
	wire w_dff_A_TN4Wuusu5_2;
	wire w_dff_A_uvaYWoK85_2;
	wire w_dff_A_HFOfGJ697_2;
	wire w_dff_A_PbS1Dyty5_0;
	wire w_dff_A_qJUwRZle8_0;
	wire w_dff_A_RXQT9YT18_0;
	wire w_dff_A_OtAELsg52_0;
	wire w_dff_A_asBKpU700_0;
	wire w_dff_A_7imHS2CW0_0;
	wire w_dff_A_z4Qm6UW55_0;
	wire w_dff_A_Eg5EPzsk6_0;
	wire w_dff_A_KIvcsf1l0_0;
	wire w_dff_A_3hLwwdsr3_0;
	wire w_dff_A_rkMHbOso7_0;
	wire w_dff_A_7jqmFCAY6_0;
	wire w_dff_A_GIN3W9H24_0;
	wire w_dff_A_QumNV0cR9_0;
	wire w_dff_A_2XITXUSG1_0;
	wire w_dff_A_D1Nz5B0M1_0;
	wire w_dff_A_KR9zwP2a9_0;
	wire w_dff_A_ofsxSK8w5_2;
	wire w_dff_A_2eh89Xiw1_2;
	wire w_dff_A_FxuohrWp6_2;
	wire w_dff_A_iCoN45B83_2;
	wire w_dff_A_LTHvzbjP6_2;
	wire w_dff_A_6CLnFoqv8_2;
	wire w_dff_A_i9sVupR50_2;
	wire w_dff_A_klecAp9m1_2;
	wire w_dff_A_iUvccvH48_2;
	wire w_dff_A_3adhuu0b5_2;
	wire w_dff_A_i3ApvijZ2_2;
	wire w_dff_A_nU4ZQWXR0_2;
	wire w_dff_A_p3UwHcrX3_2;
	wire w_dff_A_OkLzUhR09_2;
	wire w_dff_A_AWvzkvRJ0_2;
	wire w_dff_A_S61aay9x6_2;
	wire w_dff_A_TttGYNRt5_2;
	wire w_dff_A_lkiDT9Ip1_2;
	wire w_dff_A_QVJf2g3j8_2;
	wire w_dff_A_u9j9nshs9_2;
	wire w_dff_B_mshRwsy15_0;
	wire w_dff_B_5OUtjts12_0;
	wire w_dff_B_VYbzqxtc2_0;
	wire w_dff_B_IU7kvnLJ1_0;
	wire w_dff_B_YgT2FB157_0;
	wire w_dff_B_3K9M6PQ34_0;
	wire w_dff_B_B6TgXyfQ6_0;
	wire w_dff_B_HaxRkJZa8_0;
	wire w_dff_B_w7AOvR1R4_0;
	wire w_dff_B_OF7SeKIn9_0;
	wire w_dff_B_MCjGfvfv8_0;
	wire w_dff_B_3nJ1XFp51_0;
	wire w_dff_B_bjWvK6MY7_0;
	wire w_dff_B_hfGImiBG3_0;
	wire w_dff_B_3jmRfZ6H2_0;
	wire w_dff_B_oSGRjATN5_0;
	wire w_dff_B_Ds0udzs05_0;
	wire w_dff_B_eVq55WOs0_0;
	wire w_dff_B_ZwbUsRCP6_0;
	wire w_dff_B_G4jUsiup6_1;
	wire w_dff_B_4t4hdD2x4_1;
	wire w_dff_B_iodepxmR8_1;
	wire w_dff_A_GSyRofOQ7_0;
	wire w_dff_A_hgh9N07M2_0;
	wire w_dff_A_u9sRUKwF3_0;
	wire w_dff_A_Tyr7VT9b3_0;
	wire w_dff_A_Q1yahVas4_0;
	wire w_dff_A_ofsuAHg40_0;
	wire w_dff_A_BCdCY5Bq5_1;
	wire w_dff_A_ECxU1y2h3_0;
	wire w_dff_A_4CVT1Hot5_0;
	wire w_dff_A_ctnCsLVJ4_0;
	wire w_dff_A_wZh9lAPx0_0;
	wire w_dff_A_8mUEnxPQ0_1;
	wire w_dff_A_logOGiod7_1;
	wire w_dff_A_ifnZ00NC1_0;
	wire w_dff_A_D1Ua89gJ3_0;
	wire w_dff_A_k64mAtH56_0;
	wire w_dff_A_SLZgQgE55_0;
	wire w_dff_A_BwyTTUWD1_0;
	wire w_dff_A_f5mbHDtI7_0;
	wire w_dff_A_9zUtyW7p6_1;
	wire w_dff_B_XjaC9nKG1_0;
	wire w_dff_B_ZEDC7mwH7_0;
	wire w_dff_B_EkORrSbH4_0;
	wire w_dff_B_NvgGy6PA7_0;
	wire w_dff_B_8tzfis8M8_0;
	wire w_dff_B_0PaRI3PM5_0;
	wire w_dff_B_JTsamusx0_0;
	wire w_dff_B_HjvntQIJ4_0;
	wire w_dff_B_wrYh4IKt1_0;
	wire w_dff_B_GOTQGqsC4_0;
	wire w_dff_B_5sRSuzAU3_0;
	wire w_dff_B_bB6CWHQR7_0;
	wire w_dff_B_f1w60ZHt1_0;
	wire w_dff_B_1f3yI4xk6_0;
	wire w_dff_B_FOvcNYLR7_0;
	wire w_dff_B_PKY53IIb3_0;
	wire w_dff_B_TCGNstJk9_0;
	wire w_dff_B_RiYAOghw7_0;
	wire w_dff_B_MSnu5F2k2_0;
	wire w_dff_B_A9RfTUUr4_0;
	wire w_dff_B_pXPjkzqj2_1;
	wire w_dff_B_rVKnJ34T9_1;
	wire w_dff_B_Hkk4bdr51_1;
	wire w_dff_B_5SSN6Lbr9_1;
	wire w_dff_B_B44k5oz26_1;
	wire w_dff_B_Sl64ll7i0_1;
	wire w_dff_B_q7pKPDPL3_1;
	wire w_dff_B_HiWYwMmy0_1;
	wire w_dff_B_VptNvT6w3_1;
	wire w_dff_B_O5t6VBUW4_1;
	wire w_dff_B_R1GJTSVh0_1;
	wire w_dff_B_AeROLd9g8_1;
	wire w_dff_B_OtN8yW254_1;
	wire w_dff_B_xMoW2Dhx7_1;
	wire w_dff_B_nc1BxIhm3_1;
	wire w_dff_B_9OE8mQuF3_1;
	wire w_dff_B_2fhg3qiy4_1;
	wire w_dff_B_HvNa44bQ7_1;
	wire w_dff_B_62WZ5jra6_1;
	wire w_dff_B_KUFA6Oyb8_1;
	wire w_dff_B_dzStsXEr1_1;
	wire w_dff_A_UJV9MCdP1_0;
	wire w_dff_A_LZMJYExx1_1;
	wire w_dff_B_CWFOGWVM9_0;
	wire w_dff_B_wh8zH6Xi6_1;
	wire w_dff_B_72Kzoy8E7_1;
	wire w_dff_B_Q6iNnIcH9_1;
	wire w_dff_B_ksA3Qrcc9_1;
	wire w_dff_B_wevj9OWe1_1;
	wire w_dff_B_Hyvlp0Q17_1;
	wire w_dff_B_VO9tCWRW9_1;
	wire w_dff_B_6qWfUCn13_1;
	wire w_dff_B_rF5XBp3F5_1;
	wire w_dff_B_q2oX5MxI5_1;
	wire w_dff_B_Zf2qB9y65_1;
	wire w_dff_B_opxgwODg5_1;
	wire w_dff_B_2Qs9TehO5_1;
	wire w_dff_B_mkKF3TOm3_1;
	wire w_dff_B_CF0ODAgd0_1;
	wire w_dff_B_ITanyA184_1;
	wire w_dff_B_TnTWAq0f1_1;
	wire w_dff_B_avgwYtql8_1;
	wire w_dff_B_iOkN3Tgq2_1;
	wire w_dff_B_uDgQeQAK7_1;
	wire w_dff_B_7pe10V1S7_1;
	wire w_dff_A_6wDgPfXN7_0;
	wire w_dff_A_aNM8e70a3_2;
	wire w_dff_A_qISB8Hi53_0;
	wire w_dff_A_lDSczqec3_0;
	wire w_dff_A_50ph0ZCE3_1;
	wire w_dff_A_WwQXQ3I17_0;
	wire w_dff_A_eVmXohnV6_0;
	wire w_dff_A_DbZeV6nr6_0;
	wire w_dff_A_1etL4rPz1_0;
	wire w_dff_A_bfifcuy50_0;
	wire w_dff_A_VdkDATmk3_0;
	wire w_dff_A_2kyhzeyN1_0;
	wire w_dff_A_gPS5eRIT7_0;
	wire w_dff_A_SKtBkKNz4_0;
	wire w_dff_A_YWrBOHVH9_0;
	wire w_dff_A_icU0pCwP7_0;
	wire w_dff_A_8I1dSzGc2_1;
	wire w_dff_A_cTZ304fU9_1;
	wire w_dff_A_vvxP8EPU3_1;
	wire w_dff_A_aU4vB9mg4_1;
	wire w_dff_B_MiQC4BOV2_3;
	wire w_dff_B_j9vnrFtC6_3;
	wire w_dff_B_CHG1cYSZ7_3;
	wire w_dff_B_43syjiHN9_3;
	wire w_dff_B_qScJs4je2_3;
	wire w_dff_B_k72mfSlZ3_3;
	wire w_dff_B_GMYqfW2v4_3;
	wire w_dff_B_oSYOYOBo4_3;
	wire w_dff_B_p5mSOc3W6_3;
	wire w_dff_B_1G6woDmf7_0;
	wire w_dff_A_yx0qjRcw3_0;
	wire w_dff_B_V96hvkE21_0;
	wire w_dff_B_0ebIHGfR9_0;
	wire w_dff_B_JrInJpB18_0;
	wire w_dff_B_tJhIb1Y94_0;
	wire w_dff_B_iZd4IPhy2_0;
	wire w_dff_B_C8WdSPPp4_0;
	wire w_dff_B_2x7Nb5SJ0_0;
	wire w_dff_B_uxahMi3I1_0;
	wire w_dff_B_MOWosIV59_0;
	wire w_dff_B_RRjpjFhs7_0;
	wire w_dff_B_4yVWTyJK9_0;
	wire w_dff_B_EWZchb1d4_0;
	wire w_dff_B_XQUCCKxY1_0;
	wire w_dff_B_qhLkxiM24_0;
	wire w_dff_B_Peuvko154_0;
	wire w_dff_B_2IsVHzDB9_0;
	wire w_dff_B_v5HfP5tI9_0;
	wire w_dff_B_hE9dgaei3_0;
	wire w_dff_B_uQVjHuL17_0;
	wire w_dff_B_YqnsoghZ2_2;
	wire w_dff_B_L9QBeQMZ4_2;
	wire w_dff_B_nk58Ujfl0_2;
	wire w_dff_B_9dwlTRPK6_1;
	wire w_dff_B_PT7K2flI5_1;
	wire w_dff_B_loIilNij4_1;
	wire w_dff_B_rjIiuDHl2_1;
	wire w_dff_B_7TDxlIQa1_1;
	wire w_dff_B_5ihw5G2E1_1;
	wire w_dff_B_wviYuKru8_1;
	wire w_dff_B_zbm6UKsS6_1;
	wire w_dff_B_K3n1nNSV3_1;
	wire w_dff_B_ZcR4iINm1_1;
	wire w_dff_B_gMj0zf4J9_1;
	wire w_dff_B_zWezU6xw5_1;
	wire w_dff_B_gWEPWpSj1_1;
	wire w_dff_B_87kswRpq0_1;
	wire w_dff_B_Nemvtexz4_1;
	wire w_dff_B_WgBFhtdP5_1;
	wire w_dff_B_cZwe1DK44_0;
	wire w_dff_B_o9C2OPcf2_0;
	wire w_dff_B_wLPm1KOO0_0;
	wire w_dff_B_nDHwnwGW7_0;
	wire w_dff_B_EYSEgImC0_0;
	wire w_dff_B_bAtU5uxE1_0;
	wire w_dff_B_w91Uzqrj3_0;
	wire w_dff_B_GLBNoV7e9_0;
	wire w_dff_B_hcrYth2O5_0;
	wire w_dff_B_0aVBOMGB7_1;
	wire w_dff_B_NJkMpDqu5_1;
	wire w_dff_B_a8do0Dqr7_1;
	wire w_dff_B_Z0yc7H8z2_1;
	wire w_dff_A_drOFPCxq5_0;
	wire w_dff_A_8rLOe6ph0_0;
	wire w_dff_A_2058o5338_0;
	wire w_dff_A_tWvOCbwQ7_0;
	wire w_dff_A_hJmoriM15_0;
	wire w_dff_A_aQU1CCTB6_0;
	wire w_dff_A_VvUbhN3i4_1;
	wire w_dff_B_0cT48kfH1_1;
	wire w_dff_B_YqWTLaJc9_1;
	wire w_dff_B_2wtltuUq8_1;
	wire w_dff_B_EiUttOfP5_1;
	wire w_dff_B_mzEKJfeg8_1;
	wire w_dff_B_qfssFEbD9_1;
	wire w_dff_B_crIQj7qM0_1;
	wire w_dff_B_o6X1Biji3_1;
	wire w_dff_B_plA96Sp41_1;
	wire w_dff_B_wYcNF72E0_1;
	wire w_dff_B_AJAIRTUo0_1;
	wire w_dff_B_Yz38cpht3_0;
	wire w_dff_B_16grj9909_0;
	wire w_dff_B_jMmVjyZ13_0;
	wire w_dff_B_kYUGtDk47_0;
	wire w_dff_B_bRt2jkGY6_0;
	wire w_dff_B_1D18vVm55_0;
	wire w_dff_B_gq1cU9fC3_0;
	wire w_dff_A_XuHGCyMi4_1;
	wire w_dff_A_3UiLo4Hm1_1;
	wire w_dff_A_j4GCz1dc7_1;
	wire w_dff_A_Dd14Iau00_1;
	wire w_dff_A_NWcfJXEZ4_1;
	wire w_dff_B_FXQfZfv44_1;
	wire w_dff_B_ZkhZLG0U8_1;
	wire w_dff_B_6zUhAI5o8_1;
	wire w_dff_B_NHWHS9m69_1;
	wire w_dff_B_Yf1OiBcp7_1;
	wire w_dff_B_sfEVgNFW5_1;
	wire w_dff_B_cI72lTST0_1;
	wire w_dff_B_a73Lzl8l8_1;
	wire w_dff_A_YUy9gswz0_0;
	wire w_dff_A_wJ0rPfhU5_0;
	wire w_dff_A_IyJKfD3T3_0;
	wire w_dff_A_Txew2Vfp7_0;
	wire w_dff_A_vQklMjXr9_1;
	wire w_dff_A_dUMO3B2W6_1;
	wire w_dff_B_oiWrOPgC5_1;
	wire w_dff_B_uPoQbdIH4_1;
	wire w_dff_B_OBS3g2MD6_1;
	wire w_dff_B_vRpJerCc7_1;
	wire w_dff_B_eEOFLAnR3_1;
	wire w_dff_B_iG0hA9XB8_1;
	wire w_dff_B_bLBowyVr4_1;
	wire w_dff_B_Vw1PNlQ50_1;
	wire w_dff_B_B1Drztfj2_1;
	wire w_dff_B_s33XO3VT3_1;
	wire w_dff_B_Hvj9p1CS1_1;
	wire w_dff_B_Z0FtxrQn2_1;
	wire w_dff_B_HzCBsusF0_1;
	wire w_dff_B_n8thrS4o6_1;
	wire w_dff_B_y3wcn8El9_1;
	wire w_dff_B_FLllfVbz0_1;
	wire w_dff_B_FhaLKTVj6_1;
	wire w_dff_B_v0WGhzjX8_1;
	wire w_dff_B_bzeMK1fT3_1;
	wire w_dff_B_5IvycdOU8_1;
	wire w_dff_B_vUtVT9m51_1;
	wire w_dff_B_ihfIsuao4_1;
	wire w_dff_B_VWcK5Uf26_1;
	wire w_dff_B_YyvVml4o9_1;
	wire w_dff_B_Ox1teccs8_1;
	wire w_dff_B_IL0nLb354_1;
	wire w_dff_B_xBqMGKt79_1;
	wire w_dff_B_TyuQO03d8_1;
	wire w_dff_B_PmO4LLJt6_1;
	wire w_dff_B_OH7RfCxk1_1;
	wire w_dff_B_TY5Sj4AG7_1;
	wire w_dff_B_orCNM4oi7_1;
	wire w_dff_B_YQPpm5Ql9_1;
	wire w_dff_B_LDa2sPMR3_1;
	wire w_dff_B_3gr4XNVP0_1;
	wire w_dff_B_1UIdvnZ30_1;
	wire w_dff_B_0dAciVI05_1;
	wire w_dff_B_wL4MJtRq5_1;
	wire w_dff_B_CnZd14OF3_1;
	wire w_dff_B_1GFeygu12_1;
	wire w_dff_B_VbEgjxJI3_1;
	wire w_dff_B_iWrNKJ1q4_1;
	wire w_dff_B_EoFMXOvM4_1;
	wire w_dff_B_mecnd2lm6_1;
	wire w_dff_B_pWooJQ6N1_1;
	wire w_dff_B_SpJwA4xT9_1;
	wire w_dff_B_4aUXaKp82_1;
	wire w_dff_B_NSWFAZke9_1;
	wire w_dff_B_9FWr1jvA3_1;
	wire w_dff_B_LkMPGFUk7_1;
	wire w_dff_B_09uUXe1F4_1;
	wire w_dff_B_6miQpeoH1_1;
	wire w_dff_B_SUQali7o2_1;
	wire w_dff_B_TX8TZ7nS5_1;
	wire w_dff_B_ml053Y7a4_1;
	wire w_dff_B_zM4vQe9H9_1;
	wire w_dff_B_NqMwqEwj1_1;
	wire w_dff_B_uDIAkuJh8_1;
	wire w_dff_B_4Ds4lwDP6_1;
	wire w_dff_B_rugrNiAY1_1;
	wire w_dff_B_2GLPIZQU0_1;
	wire w_dff_B_wmJzhUul9_1;
	wire w_dff_B_6iZu3XYm1_1;
	wire w_dff_B_36cErOhx8_1;
	wire w_dff_B_hdVA9NAc7_1;
	wire w_dff_B_YXFtEMAb1_1;
	wire w_dff_B_Mdvbhfnk6_1;
	wire w_dff_B_BbWxzuR80_1;
	wire w_dff_B_Vn79ltD42_1;
	wire w_dff_B_6ozC2TyU9_1;
	wire w_dff_B_4rAGShJn3_1;
	wire w_dff_B_vlAIQwl63_1;
	wire w_dff_B_wMyLAZ3k7_1;
	wire w_dff_B_Q27boKAz4_1;
	wire w_dff_B_35MiG9rW5_1;
	wire w_dff_B_ir4hScXx5_0;
	wire w_dff_B_obby5ZU81_0;
	wire w_dff_B_m85n1ZBn4_0;
	wire w_dff_B_b8kt6Wkf8_0;
	wire w_dff_B_AKBW287S2_0;
	wire w_dff_B_D5xZkAnS0_0;
	wire w_dff_B_7EN0PYJH2_0;
	wire w_dff_B_x5B54nql4_0;
	wire w_dff_B_a6DELSnI0_0;
	wire w_dff_B_UTvvvdCC3_0;
	wire w_dff_B_OAYKGmcQ1_1;
	wire w_dff_B_CLR5woc61_1;
	wire w_dff_B_XX0ct9dH3_1;
	wire w_dff_B_Y7CtRPxk3_1;
	wire w_dff_B_KRGjoyy10_1;
	wire w_dff_B_0E93b3yT7_1;
	wire w_dff_B_LYFCAq8x0_1;
	wire w_dff_B_x1Br0cAA6_1;
	wire w_dff_B_moZESCAc2_1;
	wire w_dff_B_u6qAhvxI0_1;
	wire w_dff_B_CqzsS1yo9_1;
	wire w_dff_B_LkPlro0g7_1;
	wire w_dff_B_yOBdlYSZ5_1;
	wire w_dff_B_1V7xgzM43_1;
	wire w_dff_B_34l2otit6_1;
	wire w_dff_B_H0lVh1nh9_1;
	wire w_dff_B_QvouAMqL3_1;
	wire w_dff_B_8OPEYJCD1_0;
	wire w_dff_B_neZGfiL07_2;
	wire w_dff_B_ZnjI2Mea3_2;
	wire w_dff_B_F37cIesD2_2;
	wire w_dff_B_NJKycKug6_0;
	wire w_dff_B_XaZ9PEMo0_0;
	wire w_dff_B_XVgbybfh2_0;
	wire w_dff_B_GY20Zzwl9_0;
	wire w_dff_B_12NrCWhL7_0;
	wire w_dff_B_LIThVoW39_0;
	wire w_dff_B_yV6ugsuj1_0;
	wire w_dff_B_xmSoYhIA3_0;
	wire w_dff_B_xIb444Sp1_0;
	wire w_dff_B_w8M16BaX6_0;
	wire w_dff_B_ZP7sJByb6_0;
	wire w_dff_B_mxeqjROu1_0;
	wire w_dff_B_dR9Cj0wd5_0;
	wire w_dff_B_8R29XEmq1_0;
	wire w_dff_B_3t0ytUIN2_0;
	wire w_dff_B_VdFA3uXc8_0;
	wire w_dff_B_zBOwiPRE2_0;
	wire w_dff_B_R9I2p3F84_0;
	wire w_dff_B_c0egVQFZ4_0;
	wire w_dff_B_fv6coIyT0_0;
	wire w_dff_B_ZtJzWLSh7_2;
	wire w_dff_B_yNKzXfDQ4_2;
	wire w_dff_B_TFS1KFt26_2;
	wire w_dff_B_5R8yb2h83_1;
	wire w_dff_B_MuWztHRc9_1;
	wire w_dff_B_47rOcSoE7_1;
	wire w_dff_B_2mtnGLZK5_1;
	wire w_dff_B_BzZH3Vxg6_1;
	wire w_dff_B_HIwuIvE63_1;
	wire w_dff_B_aTWj3rFY0_1;
	wire w_dff_B_tU45p0v45_1;
	wire w_dff_B_thUqQi0U2_1;
	wire w_dff_B_G6K8jEA21_1;
	wire w_dff_B_BFwHCQF72_1;
	wire w_dff_B_KcQfyADH8_1;
	wire w_dff_B_4WokPKmk0_1;
	wire w_dff_B_BUurbvki8_1;
	wire w_dff_B_U2AdnZx40_1;
	wire w_dff_B_6vS3LmRH4_1;
	wire w_dff_B_4K2baa6I4_0;
	wire w_dff_B_EP8hHyTu6_0;
	wire w_dff_B_9rBKJiMz1_0;
	wire w_dff_B_bKCYm0Lj0_0;
	wire w_dff_B_ygQFlegl9_0;
	wire w_dff_B_qGnB5wcK3_0;
	wire w_dff_B_FIvrXbRt6_0;
	wire w_dff_B_PWAiMeGW4_0;
	wire w_dff_B_GwYmBqHV9_0;
	wire w_dff_B_QRj5i3yC5_0;
	wire w_dff_A_jnYcwbEQ9_1;
	wire w_dff_A_EUTT2E089_1;
	wire w_dff_A_WtRAsExu8_1;
	wire w_dff_B_zSbUmewt1_1;
	wire w_dff_B_whIVPNaU5_3;
	wire w_dff_B_19v3Jvts2_1;
	wire w_dff_A_nlNa4cWH9_0;
	wire w_dff_A_KMteQsiu9_0;
	wire w_dff_A_okgQU3dp8_0;
	wire w_dff_A_qxrxUja80_0;
	wire w_dff_A_kfHq47ow2_0;
	wire w_dff_A_FNeIz5LM0_0;
	wire w_dff_A_r2kxfEzD2_0;
	wire w_dff_A_k7px8ZIV7_0;
	wire w_dff_A_LtgjpQ8i8_0;
	wire w_dff_A_U321d9H42_0;
	wire w_dff_A_9QojdME74_0;
	wire w_dff_A_nZtcsZiB6_1;
	wire w_dff_A_DN6DoIr47_1;
	wire w_dff_B_LI1JA4KH8_1;
	wire w_dff_B_2FIk3Z3e5_1;
	wire w_dff_B_DTvxGPpS9_1;
	wire w_dff_B_i6u3ojuc0_1;
	wire w_dff_B_mtLjG21W7_1;
	wire w_dff_B_myCJoxAL4_1;
	wire w_dff_A_81UxL76d2_0;
	wire w_dff_A_Biw7FZMg8_0;
	wire w_dff_A_wZafjZe65_1;
	wire w_dff_A_PYSskl8b8_1;
	wire w_dff_A_mOsICq916_1;
	wire w_dff_B_QHGv122k0_1;
	wire w_dff_B_vTfpB1Oo6_1;
	wire w_dff_A_gg4BFt0t4_0;
	wire w_dff_A_4itjFJvj8_1;
	wire w_dff_B_qUj5qikX1_1;
	wire w_dff_B_soXvq5cY5_1;
	wire w_dff_B_FA1bullw2_1;
	wire w_dff_B_GB4S7wDx5_1;
	wire w_dff_B_yztnDgi42_1;
	wire w_dff_B_okmNacrg6_1;
	wire w_dff_B_BcDB7RYW2_1;
	wire w_dff_B_I5N7PxVN3_1;
	wire w_dff_B_YFyVXOaN4_1;
	wire w_dff_B_Ks4m6jrm6_1;
	wire w_dff_B_YzEV7fZk4_1;
	wire w_dff_B_6ciOveFz7_1;
	wire w_dff_B_YGLLw1ly6_1;
	wire w_dff_B_knVKXUQD9_1;
	wire w_dff_B_JnMTqY8m2_1;
	wire w_dff_B_hq34FAy57_1;
	wire w_dff_B_s074vNxE3_1;
	wire w_dff_B_hrsDR4cm0_1;
	wire w_dff_B_TqwmG5rH1_1;
	wire w_dff_B_grEZ1lrA2_1;
	wire w_dff_B_xPtK0Ird3_1;
	wire w_dff_B_BbqvFFVD4_1;
	wire w_dff_B_PrYZA3Vf6_1;
	wire w_dff_B_AGpDPeXA6_1;
	wire w_dff_B_viVeim727_1;
	wire w_dff_B_n8YfteQh9_1;
	wire w_dff_A_48Lg9FeE2_0;
	wire w_dff_A_PmrJgT1l0_0;
	wire w_dff_A_OvYhlNeR9_0;
	wire w_dff_A_Ht6mC1u15_0;
	wire w_dff_A_CPPaZf2j7_0;
	wire w_dff_A_kD5OqBHZ5_0;
	wire w_dff_A_HuO9a9D43_0;
	wire w_dff_A_VhgcBHLo4_0;
	wire w_dff_A_RofdZU6q4_0;
	wire w_dff_A_Z2uzUbwh6_1;
	wire w_dff_A_u4BSjaXN8_1;
	wire w_dff_A_amWxjfOZ8_1;
	wire w_dff_A_JHdr3CR71_1;
	wire w_dff_A_VlXlr4Zx1_1;
	wire w_dff_A_EKaufpOh9_1;
	wire w_dff_A_bz1X9iPL0_1;
	wire w_dff_A_slPUXqXl0_1;
	wire w_dff_A_p4crpk3Y4_1;
	wire w_dff_A_2Aco52Z85_1;
	wire w_dff_A_rCM9b6PR0_1;
	wire w_dff_A_dIDY0ASi7_1;
	wire w_dff_A_QEtZXnjq8_2;
	wire w_dff_A_nD2zMoYV7_2;
	wire w_dff_A_n9UM1KJa2_2;
	wire w_dff_A_XC1Ky63H8_2;
	wire w_dff_A_ahjHc97C7_2;
	wire w_dff_A_eu1v8Eyz1_2;
	wire w_dff_A_AOUMzYVg1_2;
	wire w_dff_A_bLirk2oD2_2;
	wire w_dff_A_EJRghaxr4_2;
	wire w_dff_A_tTXFHE0C8_2;
	wire w_dff_B_RxFp7TsG0_1;
	wire w_dff_B_znfhQR8X5_1;
	wire w_dff_A_7MpZfYVu0_0;
	wire w_dff_A_twaGs9Zc4_1;
	wire w_dff_A_2ZJ92eYq8_0;
	wire w_dff_A_NEQHZNTm8_0;
	wire w_dff_A_48O7lkU96_0;
	wire w_dff_A_7bQf64Kj1_0;
	wire w_dff_A_6P2fUvRx9_0;
	wire w_dff_A_tDErR2Fk5_0;
	wire w_dff_A_LdXCM8TE3_1;
	wire w_dff_A_5pjFRJaM5_1;
	wire w_dff_A_LFNYy1Rz5_1;
	wire w_dff_A_J5bUeEfp8_1;
	wire w_dff_A_x9SmHMpY2_1;
	wire w_dff_A_E2TeOGMc6_1;
	wire w_dff_A_BlHPAdPJ1_1;
	wire w_dff_B_cxjMtlJw8_0;
	wire w_dff_B_bZ5cU1fT1_0;
	wire w_dff_B_tsEXBXId4_0;
	wire w_dff_B_ffqNDHdl9_0;
	wire w_dff_B_ckBadHMd5_0;
	wire w_dff_B_hib07Wuo9_0;
	wire w_dff_B_lFNrILTE4_0;
	wire w_dff_B_rl3MElyJ5_0;
	wire w_dff_B_6dzn9GO70_0;
	wire w_dff_B_bZRkqF2K7_0;
	wire w_dff_B_GR5fnkDR0_0;
	wire w_dff_B_Tz2X3wya2_0;
	wire w_dff_B_33A2G5uo7_0;
	wire w_dff_B_XoFoH3AL8_0;
	wire w_dff_B_ZS5T9I4M9_0;
	wire w_dff_B_TO8jWDqr6_0;
	wire w_dff_B_wvWJ9g7h6_0;
	wire w_dff_B_m3ss79Mj7_0;
	wire w_dff_B_pD1sRVPu5_0;
	wire w_dff_B_Q00mXVOW6_0;
	wire w_dff_B_Gd68TiCk6_2;
	wire w_dff_B_O0W6fqH48_2;
	wire w_dff_B_tFRk1qYy6_2;
	wire w_dff_B_qYaEM9A89_1;
	wire w_dff_B_HcIJJcHd9_1;
	wire w_dff_B_O0DIQGRk2_1;
	wire w_dff_B_yld60UzA6_1;
	wire w_dff_B_3IgSQrui5_1;
	wire w_dff_B_qiOAYz3y8_1;
	wire w_dff_B_WlieLL8S0_1;
	wire w_dff_B_NpWqOmwQ7_1;
	wire w_dff_B_ASSwQiPh3_1;
	wire w_dff_B_38TLV40j6_1;
	wire w_dff_B_lzFDADZH4_1;
	wire w_dff_B_PDh3NrwN4_1;
	wire w_dff_B_4G2NvpMz1_1;
	wire w_dff_B_u6HFsEeJ0_1;
	wire w_dff_B_HwXft9pr8_1;
	wire w_dff_B_AMKwCWI48_1;
	wire w_dff_B_sN7HnCoS3_0;
	wire w_dff_B_dztaGO7m3_0;
	wire w_dff_B_vRp4HNDj0_0;
	wire w_dff_B_sAM8TalL7_0;
	wire w_dff_B_EorSIbqx9_0;
	wire w_dff_B_5XM3uvJJ3_0;
	wire w_dff_B_zOyDH3mQ8_0;
	wire w_dff_B_mldHocTn9_0;
	wire w_dff_B_pHvw4bJ66_0;
	wire w_dff_B_QqSS2F190_0;
	wire w_dff_B_qLenSkaw9_0;
	wire w_dff_B_0MzYLJRa4_0;
	wire w_dff_A_SG3G3CBN4_1;
	wire w_dff_A_1qyT3Zbc1_1;
	wire w_dff_A_HFuQmKcx2_2;
	wire w_dff_A_bqRP7G405_2;
	wire w_dff_B_teBg1fcI7_0;
	wire w_dff_B_JsXWV9FB2_0;
	wire w_dff_A_h5ADyBn98_0;
	wire w_dff_A_bourfFbx5_0;
	wire w_dff_A_sCcRFz7k0_0;
	wire w_dff_A_sJYbWsjZ4_0;
	wire w_dff_A_SBP5Ix5F2_0;
	wire w_dff_A_BCdrsiL09_0;
	wire w_dff_A_mTjCCKB56_0;
	wire w_dff_A_yP8gDsbq5_0;
	wire w_dff_A_TB7xn0HS8_0;
	wire w_dff_A_IaFBTQD19_1;
	wire w_dff_A_4JUUZQCO5_1;
	wire w_dff_A_04xqFnmw4_1;
	wire w_dff_A_Q3jqABZ76_1;
	wire w_dff_A_Xjp4Fyrw4_0;
	wire w_dff_A_Ia90jEnu5_2;
	wire w_dff_A_rM0uCabR7_2;
	wire w_dff_A_1CM9AJNo4_2;
	wire w_dff_A_UBpo4WQX6_2;
	wire w_dff_A_hh5e29xM8_2;
	wire w_dff_A_M33o1OnK1_2;
	wire w_dff_A_psOYotzO8_2;
	wire w_dff_A_TL9SRI464_2;
	wire w_dff_A_GUynjsb18_2;
	wire w_dff_A_DBT6MTiZ9_2;
	wire w_dff_A_M4lVm0cV4_2;
	wire w_dff_A_dOIPu4iG2_2;
	wire w_dff_A_TKAGjbmO2_2;
	wire w_dff_A_4cKtydrZ2_2;
	wire w_dff_A_rIPRvKlC4_0;
	wire w_dff_A_tVjet4u93_0;
	wire w_dff_A_OnstN0Yx8_0;
	wire w_dff_A_T3jpC6XO6_2;
	wire w_dff_A_DhcTfbY66_2;
	wire w_dff_A_yRoGyYAK2_0;
	wire w_dff_A_sXry6PBj4_0;
	wire w_dff_A_46GWPNeP7_0;
	wire w_dff_A_hKkU8OVO1_0;
	wire w_dff_A_wf6cAqmr3_0;
	wire w_dff_A_8EA8ujsr5_0;
	wire w_dff_A_Tsv6D9am1_0;
	wire w_dff_A_klfcE5ZW5_0;
	wire w_dff_A_UbutgT4e4_0;
	wire w_dff_A_XT0ifyt51_1;
	wire w_dff_A_xDJ80oeC7_1;
	wire w_dff_B_IyTF2DcU4_3;
	wire w_dff_B_WHkje4zU7_3;
	wire w_dff_B_vyq0mpfB3_3;
	wire w_dff_B_N1nOxGne4_3;
	wire w_dff_B_c1AparXY2_3;
	wire w_dff_B_0dlJOkYq9_3;
	wire w_dff_B_rtLfTblU3_3;
	wire w_dff_B_FJNAxe5d6_3;
	wire w_dff_B_V0fEmAEL9_3;
	wire w_dff_B_eebWSicJ6_3;
	wire w_dff_B_Oqq6t7dM4_3;
	wire w_dff_B_x6DPUGDY8_1;
	wire w_dff_B_DZn4P6eY6_1;
	wire w_dff_B_JqBHtfFn8_1;
	wire w_dff_B_Y8deJoUJ1_1;
	wire w_dff_B_T1WueL0q9_1;
	wire w_dff_B_fhEtG3S93_1;
	wire w_dff_B_sPtZDwYz6_1;
	wire w_dff_B_vTuHdIBO3_1;
	wire w_dff_B_Y7hqqX3B0_1;
	wire w_dff_B_nZyru5xd0_1;
	wire w_dff_B_uY9k2vfD6_1;
	wire w_dff_B_mdCuGgsK5_1;
	wire w_dff_B_dGYrlCKi3_1;
	wire w_dff_B_6Wyove6d3_1;
	wire w_dff_B_HiWT2w0S7_1;
	wire w_dff_B_KjJlP0Ik6_1;
	wire w_dff_B_xBbinTII5_1;
	wire w_dff_B_U1VjBKb27_1;
	wire w_dff_B_WcuDG3Rh0_1;
	wire w_dff_B_MZHgArMs4_1;
	wire w_dff_B_PQVlnszt2_1;
	wire w_dff_B_RkINFyKm2_1;
	wire w_dff_B_QJgowWFx3_1;
	wire w_dff_B_pW2uDacm8_1;
	wire w_dff_B_aanXl7Ko2_1;
	wire w_dff_B_AbRIiNki4_1;
	wire w_dff_B_2xpmdX743_1;
	wire w_dff_B_ME5vetwx8_1;
	wire w_dff_B_GtU33t4T5_1;
	wire w_dff_B_xrdT1GMN5_1;
	wire w_dff_B_zXT6ynzD3_1;
	wire w_dff_B_0HBF12dA9_1;
	wire w_dff_B_M8VSGcPA7_1;
	wire w_dff_B_Xfnlr1HJ1_1;
	wire w_dff_B_3WgbZ8Dl5_1;
	wire w_dff_B_m9iJzj4t6_1;
	wire w_dff_B_WIqywlki5_1;
	wire w_dff_B_VxkkGQO10_1;
	wire w_dff_B_PvmQsIGm0_1;
	wire w_dff_B_Gyu7mPT03_1;
	wire w_dff_B_zzQxdAZy6_0;
	wire w_dff_B_IKO5kJGV8_1;
	wire w_dff_B_Hm0NnoUi5_1;
	wire w_dff_A_Mo9sV4jz4_1;
	wire w_dff_B_naccYboo1_3;
	wire w_dff_B_8MPEj8T95_3;
	wire w_dff_B_LILldglh2_3;
	wire w_dff_B_aOff08097_3;
	wire w_dff_B_UYB3ZrXN6_3;
	wire w_dff_A_9yjaLKeD7_0;
	wire w_dff_A_IBBWSIUp1_1;
	wire w_dff_A_t9wquEM91_1;
	wire w_dff_B_PqvOZdZ71_3;
	wire w_dff_B_efUeAKq74_3;
	wire w_dff_B_kFqFvyp07_3;
	wire w_dff_B_se4LDacT7_3;
	wire w_dff_B_zzah0dQD8_3;
	wire w_dff_B_B5S7AWBv8_3;
	wire w_dff_B_gpdwNBUO6_3;
	wire w_dff_B_JjLzSQoQ5_3;
	wire w_dff_B_dCJ9NGDw9_3;
	wire w_dff_B_kIrk9FHa7_3;
	wire w_dff_B_xpHjaMtT7_3;
	wire w_dff_B_LeEQJQeX5_3;
	wire w_dff_B_o7daRyHo8_3;
	wire w_dff_B_20QxDwqu1_3;
	wire w_dff_B_6JI8y1nQ3_3;
	wire w_dff_A_0LASztWG5_0;
	wire w_dff_A_Mli2ce8Q1_0;
	wire w_dff_A_VRkDdy4a7_0;
	wire w_dff_A_ZM5H8oma0_0;
	wire w_dff_A_TNMG6spc9_0;
	wire w_dff_A_AOhrr9dn7_0;
	wire w_dff_A_5zR3yP6r9_1;
	wire w_dff_A_9HxEik9S3_1;
	wire w_dff_A_uRsiHsta8_1;
	wire w_dff_A_OJRTFFqW7_1;
	wire w_dff_A_2CQVESU27_1;
	wire w_dff_A_lB8jkucz9_1;
	wire w_dff_A_CclZyRgt7_0;
	wire w_dff_A_sHnMweYL9_0;
	wire w_dff_A_RzxkQFGd9_0;
	wire w_dff_A_VuzFRFpJ3_0;
	wire w_dff_A_oHcayFwH2_0;
	wire w_dff_A_wbv0D6hL1_0;
	wire w_dff_A_jqeDkZhf1_0;
	wire w_dff_A_VeGW5vE50_0;
	wire w_dff_A_WzB4BH967_0;
	wire w_dff_A_HOVFvIwm8_0;
	wire w_dff_A_JO9RWGma1_0;
	wire w_dff_A_7x2yeONB8_0;
	wire w_dff_A_Etcec46M3_0;
	wire w_dff_A_fScvVv0S0_0;
	wire w_dff_A_poGi5q4w6_1;
	wire w_dff_A_NtPI2eCN5_1;
	wire w_dff_B_6wMq7sdz6_1;
	wire w_dff_B_OUybV2HC1_1;
	wire w_dff_B_Dpc3eSHg5_0;
	wire w_dff_B_33XXtlKC0_0;
	wire w_dff_B_xPQrDetT7_0;
	wire w_dff_B_VjUnHcXl1_0;
	wire w_dff_B_NyYosQTj0_0;
	wire w_dff_B_6GiQMakZ3_0;
	wire w_dff_B_xDIgkjsQ7_0;
	wire w_dff_B_Vn6DWYu36_0;
	wire w_dff_B_Xy6Pan1d4_0;
	wire w_dff_B_E3XKDFEP0_0;
	wire w_dff_B_RGuPtAUl9_0;
	wire w_dff_B_HsBGya5a5_0;
	wire w_dff_B_FFNl50ZA3_0;
	wire w_dff_B_LfUUAna41_0;
	wire w_dff_B_9jbclwIf6_0;
	wire w_dff_B_54sFbtbX3_0;
	wire w_dff_B_bBgJxmY12_0;
	wire w_dff_B_LssX4v2H2_1;
	wire w_dff_B_aybXx0cm8_1;
	wire w_dff_B_yIyzP5Yo3_1;
	wire w_dff_B_AQMrhbqO2_0;
	wire w_dff_B_639ljYov0_0;
	wire w_dff_B_HlDp2aqp3_0;
	wire w_dff_B_6RcG2bXo2_0;
	wire w_dff_B_i48s8PXH0_0;
	wire w_dff_B_nx1Xqc5Y0_0;
	wire w_dff_B_SDKdmsel8_0;
	wire w_dff_B_QWJZBtDZ5_0;
	wire w_dff_B_RX0gvrzg4_0;
	wire w_dff_B_YPJ1XIzA3_0;
	wire w_dff_B_e0xHLQmV3_0;
	wire w_dff_B_4lCDyEm47_0;
	wire w_dff_B_3JJNPPks3_0;
	wire w_dff_B_SNRbhPRA2_0;
	wire w_dff_B_56tIiNrx0_0;
	wire w_dff_B_UF81N8mv8_0;
	wire w_dff_B_ivEnXF2Z0_0;
	wire w_dff_B_R8WvSjL46_1;
	wire w_dff_B_0jJGfgzu4_1;
	wire w_dff_B_kALI9UUy4_1;
	wire w_dff_A_s6k4vIgb7_0;
	wire w_dff_A_TGt0vwSs9_0;
	wire w_dff_A_X5Ahz7o40_0;
	wire w_dff_A_tot8P65E9_0;
	wire w_dff_A_OQJ74M3V3_0;
	wire w_dff_A_4XETqUAy6_1;
	wire w_dff_A_t69nBHlN1_1;
	wire w_dff_A_de7GXQsn2_1;
	wire w_dff_A_Nuq3dACF0_1;
	wire w_dff_A_diLxcyc94_0;
	wire w_dff_A_FdR8LCEy3_0;
	wire w_dff_A_Y34mV9nf4_0;
	wire w_dff_A_IzyPLtpV7_0;
	wire w_dff_A_UQCIH12x2_0;
	wire w_dff_A_4nQMsEJZ0_1;
	wire w_dff_A_sEYg9hlu1_1;
	wire w_dff_A_mSesgIDu5_1;
	wire w_dff_A_tnyGzhZ58_1;
	wire w_dff_A_qyUmYJxd1_0;
	wire w_dff_A_e5nWRFdM4_0;
	wire w_dff_A_xnnPnaiM2_0;
	wire w_dff_B_KpTvdyl23_1;
	wire w_dff_B_afC9Rhzc5_1;
	wire w_dff_B_1ovAACwt8_1;
	wire w_dff_B_956HnWuz3_1;
	wire w_dff_B_xc1ZUklw0_1;
	wire w_dff_B_kpz4Wosn0_1;
	wire w_dff_B_8nsS6u1d7_1;
	wire w_dff_B_5uEH2ZZq8_1;
	wire w_dff_B_S2ZwWOyy1_1;
	wire w_dff_B_dH5pHsAD8_1;
	wire w_dff_B_1D23wk9X7_1;
	wire w_dff_B_2qVySc086_1;
	wire w_dff_B_FN6Y1TDz0_1;
	wire w_dff_B_9Z9xNBnA7_1;
	wire w_dff_B_JYRFyvTf1_1;
	wire w_dff_B_2u7nNcwk6_1;
	wire w_dff_B_Hdw1ig2D4_1;
	wire w_dff_B_k6vZVOWm4_1;
	wire w_dff_B_EzSnGYyx7_1;
	wire w_dff_B_Y3yrwssN7_1;
	wire w_dff_B_df65VDdF6_1;
	wire w_dff_B_Dzxeri387_1;
	wire w_dff_B_z0n0vzl45_1;
	wire w_dff_A_BIiek8Bj7_1;
	wire w_dff_A_RptDZlU53_1;
	wire w_dff_A_NcSppiiC5_1;
	wire w_dff_A_uOwvCTMW1_1;
	wire w_dff_A_ILyyk1Ts0_1;
	wire w_dff_A_8sxACelC8_1;
	wire w_dff_A_rII7vRHv4_1;
	wire w_dff_A_6TnomH5k7_1;
	wire w_dff_A_iF88Yg0d9_1;
	wire w_dff_A_bKu8rEoc6_1;
	wire w_dff_A_K30UDXMw2_1;
	wire w_dff_A_QPyYg0kv1_1;
	wire w_dff_A_v386zVsG1_1;
	wire w_dff_A_twRL69CU3_1;
	wire w_dff_A_8NNw33gg1_2;
	wire w_dff_A_0sGD3zE15_2;
	wire w_dff_A_cLpzrqEb4_2;
	wire w_dff_A_mpZKO8EQ1_2;
	wire w_dff_A_CAhSMrq20_2;
	wire w_dff_A_DI3kWwgr6_2;
	wire w_dff_A_uxVazMlK0_2;
	wire w_dff_A_L7vU8Fzk1_2;
	wire w_dff_A_pdF860xr3_2;
	wire w_dff_A_llbMoU9z6_2;
	wire w_dff_A_V54IQlgl9_1;
	wire w_dff_A_9fu9BnWB3_1;
	wire w_dff_A_u89riaRk0_1;
	wire w_dff_A_QZvFthX22_1;
	wire w_dff_A_GJWRm6WC3_1;
	wire w_dff_A_HRt0K5jK9_1;
	wire w_dff_A_mAJinRlJ0_1;
	wire w_dff_A_AVlTkWD56_1;
	wire w_dff_A_Q0LnOjhy7_1;
	wire w_dff_A_h6pbmVRJ9_1;
	wire w_dff_A_a9eq3c733_1;
	wire w_dff_A_lIbZN6lz7_2;
	wire w_dff_A_9QX48GXi0_2;
	wire w_dff_A_Zdz5MnjK3_2;
	wire w_dff_A_aolLGTMm4_2;
	wire w_dff_B_d9uxW4Ca2_3;
	wire w_dff_B_aYP5Hrdf1_3;
	wire w_dff_B_ie2B6lhi7_3;
	wire w_dff_B_7oGvw9J40_3;
	wire w_dff_B_TRdCt46c9_3;
	wire w_dff_B_867Gc1Oh4_3;
	wire w_dff_B_GptRj8EL6_3;
	wire w_dff_B_YkdDG63U7_3;
	wire w_dff_B_x66oaevu3_3;
	wire w_dff_A_QYL6DxgV9_0;
	wire w_dff_A_OfrUFjPQ7_1;
	wire w_dff_B_A8hND6lq2_1;
	wire w_dff_B_hkA2TYSN3_1;
	wire w_dff_A_ouJpcfxc9_0;
	wire w_dff_A_12LU00iM3_0;
	wire w_dff_A_hSL1wZhs8_0;
	wire w_dff_A_HJpLEwt92_0;
	wire w_dff_A_sdQo5WV29_0;
	wire w_dff_A_RJoqGr2d3_0;
	wire w_dff_A_9ty7zU8L3_0;
	wire w_dff_A_7szxLVo21_0;
	wire w_dff_A_EnKdrWTh2_0;
	wire w_dff_A_ADFmU96c5_0;
	wire w_dff_A_BizjAxo16_0;
	wire w_dff_A_NFeBwL6s4_0;
	wire w_dff_A_iFHkitDq1_0;
	wire w_dff_A_elFdEM5y3_0;
	wire w_dff_A_zfcyOCwO3_0;
	wire w_dff_A_sNyB5mEX0_0;
	wire w_dff_A_bOSgJ2gc0_0;
	wire w_dff_A_hJMWeikJ5_0;
	wire w_dff_A_bNfrraTM5_0;
	wire w_dff_A_Suo2QwC29_0;
	wire w_dff_A_7JHi7eg18_0;
	wire w_dff_A_wZ31z6lw8_0;
	wire w_dff_A_F9pE1UfG6_1;
	wire w_dff_A_KghyqK1q7_1;
	wire w_dff_A_Hm9r92oa5_1;
	wire w_dff_A_WZAZvzlb7_1;
	wire w_dff_A_gvhV625k2_1;
	wire w_dff_A_sOYq1amW1_1;
	wire w_dff_A_N7iJ4y353_1;
	wire w_dff_A_sZcA6URo5_1;
	wire w_dff_A_8wb7EXNr3_1;
	wire w_dff_A_xmdQFswB1_1;
	wire w_dff_A_Qd0zoQ9U3_1;
	wire w_dff_A_huOUs4Y20_2;
	wire w_dff_A_q6Ybc1Cz7_1;
	wire w_dff_A_xUOYB4Xr8_2;
	wire w_dff_A_brdJO78o5_0;
	wire w_dff_A_y2a0ACGn3_0;
	wire w_dff_A_DSonxTwS0_0;
	wire w_dff_A_5jmEpHNJ9_0;
	wire w_dff_A_n5eK6xO55_0;
	wire w_dff_A_AMhzHlyw1_0;
	wire w_dff_A_LM9O3iq19_0;
	wire w_dff_A_yGc5cONx6_0;
	wire w_dff_A_nWVBq4qJ2_0;
	wire w_dff_A_w73qp5rs8_0;
	wire w_dff_A_tL4Et7y13_0;
	wire w_dff_A_4CjAXStS3_0;
	wire w_dff_A_MIxjJF3f0_0;
	wire w_dff_A_4VSsuf7r8_0;
	wire w_dff_A_Jg3el3Hr4_0;
	wire w_dff_A_oBrtqtPF7_0;
	wire w_dff_A_bV8ocIrG5_0;
	wire w_dff_A_4vUaiIPe2_0;
	wire w_dff_A_FdsMZ58L2_0;
	wire w_dff_A_gYL0V17u2_0;
	wire w_dff_A_v39QAdSF2_0;
	wire w_dff_A_SrMSNxNn8_0;
	wire w_dff_A_kH3PP8cX2_0;
	wire w_dff_B_wWgEURmU6_1;
	wire w_dff_B_6RbDTDSY8_1;
	wire w_dff_B_sjHsPvrq4_1;
	wire w_dff_B_TylWqUZJ8_1;
	wire w_dff_B_WMB2ssSy3_1;
	wire w_dff_B_deotQdSc1_1;
	wire w_dff_B_prHKaGzT1_1;
	wire w_dff_B_cmoVJNVd4_1;
	wire w_dff_B_ECow2kHo5_1;
	wire w_dff_B_UrhRL9iy3_1;
	wire w_dff_B_Drpq8IWm2_1;
	wire w_dff_B_VbuI1Wgc4_1;
	wire w_dff_B_u7BCC4MM6_1;
	wire w_dff_B_ggCWKT6J9_1;
	wire w_dff_B_K72oyMdX8_1;
	wire w_dff_B_nBpREnqN9_1;
	wire w_dff_B_HTK439Wq1_1;
	wire w_dff_B_mQkpyUbh2_1;
	wire w_dff_B_nakUJG386_1;
	wire w_dff_B_6UeAQqf66_1;
	wire w_dff_B_xEScLYl45_1;
	wire w_dff_B_KXlTl6Of8_1;
	wire w_dff_B_mpBfkQmG0_1;
	wire w_dff_A_8CO2i2n78_1;
	wire w_dff_A_m0qmgwmF4_1;
	wire w_dff_A_GABnNBn65_1;
	wire w_dff_A_dMeydbTF0_1;
	wire w_dff_A_XCxnLEyM4_1;
	wire w_dff_A_o0KZ2Ry60_1;
	wire w_dff_A_5iQzyDiR2_1;
	wire w_dff_A_nv6Uky7c9_1;
	wire w_dff_A_OhRSnYM09_1;
	wire w_dff_A_eHUfQdXt0_1;
	wire w_dff_A_1EjJS5qT2_1;
	wire w_dff_A_SBtYyH3t3_1;
	wire w_dff_A_o5DxYfoU2_1;
	wire w_dff_A_VXwxUIU01_1;
	wire w_dff_A_IqYpwzBl4_2;
	wire w_dff_A_owqyUvqg6_2;
	wire w_dff_A_FxL2PiIP3_2;
	wire w_dff_A_oPiS4LRt9_2;
	wire w_dff_A_diyjyDMc6_2;
	wire w_dff_A_BGpPLwCp0_2;
	wire w_dff_A_2oeB6MbB8_2;
	wire w_dff_A_8p5hOO8r7_2;
	wire w_dff_A_UHVhXrBV7_2;
	wire w_dff_A_nkBS7BN47_2;
	wire w_dff_A_DaTcnhiw0_1;
	wire w_dff_A_KOZClzYI2_1;
	wire w_dff_A_43adTSv83_1;
	wire w_dff_A_Tk4bY1Up4_1;
	wire w_dff_A_r54mcXYe8_1;
	wire w_dff_A_trPqvmZV0_1;
	wire w_dff_A_OJ9QNloY1_1;
	wire w_dff_A_KibaWw0P6_1;
	wire w_dff_A_Wrm4RB169_1;
	wire w_dff_A_QXVvkGMr7_1;
	wire w_dff_A_M28Bwhdm8_1;
	wire w_dff_A_rl4KCP451_2;
	wire w_dff_A_6D0AXka91_2;
	wire w_dff_A_tvVAPV5y0_2;
	wire w_dff_A_ot9sPm6n9_2;
	wire w_dff_A_sm2eBv348_2;
	wire w_dff_B_0qH55en87_3;
	wire w_dff_B_fIOicQFV5_3;
	wire w_dff_B_CTQbOwnL9_3;
	wire w_dff_B_yXMAhMSb3_3;
	wire w_dff_B_vHJR4ZOj0_3;
	wire w_dff_B_yHu6d2yL6_3;
	wire w_dff_B_38IArHka8_3;
	wire w_dff_B_6H7KQBPs7_3;
	wire w_dff_B_x6sYVZQl0_3;
	wire w_dff_A_Ha3cWrG17_0;
	wire w_dff_A_8kpK9Msz0_0;
	wire w_dff_A_26cKSgzW0_1;
	wire w_dff_B_XPvaKtdg5_1;
	wire w_dff_B_BTPIfn9Y7_1;
	wire w_dff_A_1kJQdAkM7_0;
	wire w_dff_A_xtTjGC7B2_0;
	wire w_dff_A_tumRi2mC0_0;
	wire w_dff_A_5d8H4D965_0;
	wire w_dff_A_t4LOqunI9_0;
	wire w_dff_A_lvXE7poB5_0;
	wire w_dff_A_JrSzFae68_0;
	wire w_dff_A_wl3A6yNu6_0;
	wire w_dff_A_e2NVKZAD3_0;
	wire w_dff_A_30FZuT7V4_0;
	wire w_dff_A_VFU3y2Mj3_0;
	wire w_dff_A_yYh1NV9p7_0;
	wire w_dff_A_fUWMkXjP4_0;
	wire w_dff_A_50TLP7jU3_0;
	wire w_dff_A_EZxFsrWR7_0;
	wire w_dff_A_zCOHU7d92_0;
	wire w_dff_A_ZEJQY0ik1_0;
	wire w_dff_A_mfdDrOci0_0;
	wire w_dff_A_knC7x9lC2_0;
	wire w_dff_A_VHtaA9oV7_0;
	wire w_dff_A_mL9wRMd47_0;
	wire w_dff_A_9DvEUrSW2_0;
	wire w_dff_A_hbAMZKfq7_1;
	wire w_dff_A_vmjKJRSN1_1;
	wire w_dff_A_Tiajxx3A1_1;
	wire w_dff_A_oWsllihA0_1;
	wire w_dff_A_5YVu1MZ45_1;
	wire w_dff_A_g70oY7j37_1;
	wire w_dff_A_du8J4sTC8_1;
	wire w_dff_A_p6eEK0KJ2_1;
	wire w_dff_A_I5dEYBgk2_1;
	wire w_dff_B_elWrQJ4U4_2;
	wire w_dff_A_J7W1hXpk2_1;
	wire w_dff_A_ksc0atqM3_1;
	wire w_dff_A_sRvNW2HZ1_2;
	wire w_dff_A_BYXvFlgx9_1;
	wire w_dff_A_f0KPsERX4_2;
	wire w_dff_A_5bHnMgvO1_0;
	wire w_dff_A_NcOI8saR6_0;
	wire w_dff_A_AAY4v8W08_0;
	wire w_dff_A_Y2CJTJSH4_0;
	wire w_dff_A_WXvvYtay2_0;
	wire w_dff_A_sRvXD0DF0_0;
	wire w_dff_A_rYlRiy2b1_0;
	wire w_dff_A_gDuGQ8eQ2_0;
	wire w_dff_A_x3ZlMNPZ7_0;
	wire w_dff_A_xZ2iOT8N9_0;
	wire w_dff_A_YuXCB6yR0_0;
	wire w_dff_A_5SncczX37_0;
	wire w_dff_A_xctXUhwh6_0;
	wire w_dff_A_OiIq1dkr0_0;
	wire w_dff_A_07BlpJUB8_0;
	wire w_dff_A_WcGox2sJ8_0;
	wire w_dff_A_ra6KoJbO5_0;
	wire w_dff_A_7Qshy0Zq4_0;
	wire w_dff_A_NtQSdMAy2_0;
	wire w_dff_A_lm9sZBkW6_0;
	wire w_dff_A_r609rUzY5_0;
	wire w_dff_A_r2wKOvRB6_0;
	wire w_dff_A_EoOpLKUe9_0;
	wire w_dff_B_11fBWxV75_1;
	wire w_dff_B_FXIPiwZP5_1;
	wire w_dff_B_S06WoP7R8_1;
	wire w_dff_B_btFqaB1x0_1;
	wire w_dff_B_OrAOC1Ty0_1;
	wire w_dff_B_CJRag0Yy6_1;
	wire w_dff_B_oyELLvTh7_1;
	wire w_dff_B_SYYQl30m5_1;
	wire w_dff_B_3FIhqHQg4_1;
	wire w_dff_B_TxWDfSME5_1;
	wire w_dff_B_c0yzu0w89_1;
	wire w_dff_B_XdpeJQ4V3_1;
	wire w_dff_B_AcwP5iZV3_1;
	wire w_dff_B_VHsBF9nZ9_1;
	wire w_dff_B_qesynLFK6_1;
	wire w_dff_B_A5gozeRD2_1;
	wire w_dff_B_7V00o5xe1_1;
	wire w_dff_B_otCXgSgC8_1;
	wire w_dff_B_0hJ2ADGE9_1;
	wire w_dff_B_QRkYaDOT7_1;
	wire w_dff_B_8i9nuOTJ5_1;
	wire w_dff_B_7IEUh2D10_1;
	wire w_dff_B_e9Ghi6we9_1;
	wire w_dff_B_qvliIxqM3_1;
	wire w_dff_B_9Zn9xc292_1;
	wire w_dff_B_KjZ2BQb95_1;
	wire w_dff_B_4KVRDxTW8_1;
	wire w_dff_B_ZWqa6y3m1_1;
	wire w_dff_B_lJcCMNJ15_1;
	wire w_dff_B_C4rCKfyl7_1;
	wire w_dff_B_E5hECoeZ3_1;
	wire w_dff_B_gXlz2jwY6_1;
	wire w_dff_B_6VLSEagO9_1;
	wire w_dff_B_cym21weM8_1;
	wire w_dff_B_paNP8PIy2_1;
	wire w_dff_B_GaLW9uUh6_1;
	wire w_dff_B_QZiAHxv07_1;
	wire w_dff_B_uP6EeV9O2_1;
	wire w_dff_B_7HbNEO788_1;
	wire w_dff_B_1OTuK1qe0_1;
	wire w_dff_B_TPuzgZuV2_1;
	wire w_dff_B_cvKNrSBj8_1;
	wire w_dff_B_btY59Hp39_1;
	wire w_dff_B_67NfPwbU8_1;
	wire w_dff_B_yJssm8oz1_1;
	wire w_dff_A_TRNTqb8g7_0;
	wire w_dff_A_X5YbrzOk1_0;
	wire w_dff_A_IDWv58Lr6_0;
	wire w_dff_A_ZfHDAFS63_0;
	wire w_dff_A_iQJ7qmd52_0;
	wire w_dff_A_Y3WZuILJ2_0;
	wire w_dff_A_XpehRAJP9_0;
	wire w_dff_A_zjPyLzpi2_0;
	wire w_dff_A_3NQp8nO86_0;
	wire w_dff_A_LwYGzmdy1_0;
	wire w_dff_A_S5FsDPRN0_0;
	wire w_dff_A_5uSh1v011_0;
	wire w_dff_A_yAi5FUeR2_0;
	wire w_dff_A_Ti2KgWbf0_0;
	wire w_dff_A_RiCzsvby6_0;
	wire w_dff_A_Q4yZm4bD6_1;
	wire w_dff_A_g2SDyqyM2_1;
	wire w_dff_A_oMrIZnTf2_1;
	wire w_dff_A_RPm7PPa61_1;
	wire w_dff_A_5QFWDxTx5_1;
	wire w_dff_A_wKAjSvf32_1;
	wire w_dff_A_Ndw55JCg7_1;
	wire w_dff_A_wZ1L0jbV0_1;
	wire w_dff_A_eoxyatnW6_1;
	wire w_dff_A_svDBm8Jc3_1;
	wire w_dff_A_8LsS5AGs9_1;
	wire w_dff_A_Hzv45t1J9_1;
	wire w_dff_A_l0mfcFzJ7_1;
	wire w_dff_A_mpCLWfXX3_1;
	wire w_dff_A_k114UFWy1_1;
	wire w_dff_A_isexrxmM3_1;
	wire w_dff_A_GUbHTYic0_1;
	wire w_dff_A_YxFsmCUO9_1;
	wire w_dff_A_7WzjAGkN5_1;
	wire w_dff_A_Cfa3sRpq4_1;
	wire w_dff_A_pJUeIIJh9_1;
	wire w_dff_A_g3NAHuLU2_1;
	wire w_dff_A_L9QpcrDr6_1;
	wire w_dff_A_X4UDypwM9_1;
	wire w_dff_A_BBPxCpfw1_1;
	wire w_dff_A_fyusDvm38_1;
	wire w_dff_A_r8gYdgL39_1;
	wire w_dff_A_0uuR7mHC8_1;
	wire w_dff_A_pHuy2eHG2_1;
	wire w_dff_A_79esEI9F5_1;
	wire w_dff_A_4fDZu6Ro7_1;
	wire w_dff_A_bhHgnIga9_2;
	wire w_dff_A_2ZpLNvk60_2;
	wire w_dff_A_w41nB2O55_2;
	wire w_dff_A_TbQbsKlG1_2;
	wire w_dff_A_dTJhylH06_2;
	wire w_dff_A_36FRNv1h1_2;
	wire w_dff_A_T3dr5okc6_2;
	wire w_dff_A_xxeHe6pM4_2;
	wire w_dff_A_2IVIVj9N2_2;
	wire w_dff_A_BxGFoL9k0_2;
	wire w_dff_A_jtMf4PbW9_2;
	wire w_dff_A_S2GKDEcz2_2;
	wire w_dff_A_WDIrb1ft6_2;
	wire w_dff_A_mJwO8NvT9_2;
	wire w_dff_A_RkUI6C059_2;
	wire w_dff_A_vHeYE6ai7_2;
	wire w_dff_A_4k2iyqIT3_2;
	wire w_dff_A_aCnRQ2sd0_2;
	wire w_dff_A_EHXd7r9L3_2;
	wire w_dff_A_0ShZnwgW3_2;
	wire w_dff_A_Ts5ejSxw1_1;
	wire w_dff_A_CDe73UGK4_1;
	wire w_dff_A_bByk705m9_1;
	wire w_dff_A_GfZmk5934_1;
	wire w_dff_A_3DGBthFm8_1;
	wire w_dff_A_7nPDNg0F7_1;
	wire w_dff_A_kzEOtdX72_1;
	wire w_dff_A_CfeLAbC85_1;
	wire w_dff_A_AbLKmgaf6_1;
	wire w_dff_A_juyqQyl61_1;
	wire w_dff_A_lPnI40po1_1;
	wire w_dff_A_a38Z7zQv2_1;
	wire w_dff_A_PVQH0J5H3_1;
	wire w_dff_A_vDD9AvLr0_1;
	wire w_dff_A_fxnYGVro0_1;
	wire w_dff_A_55eL2Zly2_1;
	wire w_dff_A_2bvKdXBt2_1;
	wire w_dff_A_yLxDTtHx7_1;
	wire w_dff_A_QDnuycIy2_2;
	wire w_dff_A_nVY3kyfG2_2;
	wire w_dff_A_4uFGPOqR0_2;
	wire w_dff_A_qV0CoZK13_2;
	wire w_dff_A_7ZCWIkBK5_2;
	wire w_dff_A_dXpnKGlN6_2;
	wire w_dff_A_O3hIAkMv6_2;
	wire w_dff_A_XPplqGCX4_2;
	wire w_dff_A_h47oQwxH6_2;
	wire w_dff_A_9MANMymo8_2;
	wire w_dff_A_7HUVL1Pp0_2;
	wire w_dff_A_7MZiC1pn7_1;
	wire w_dff_A_CozOhow45_1;
	wire w_dff_A_KNoEf7Di6_1;
	wire w_dff_A_iDD1DUjj3_1;
	wire w_dff_A_fJZFzTZc2_1;
	wire w_dff_A_svg15Zt01_1;
	wire w_dff_A_1IzpDqem3_1;
	wire w_dff_A_OBV2Z7rV0_1;
	wire w_dff_A_LvLFPvna1_1;
	wire w_dff_A_XlGW3R8C5_1;
	wire w_dff_A_Hr0t9hil2_1;
	wire w_dff_A_ycKLrXAJ5_1;
	wire w_dff_A_4Xxacixz3_1;
	wire w_dff_A_PIjAaaZW0_1;
	wire w_dff_A_57glIP3i7_1;
	wire w_dff_A_YxmSF84j0_1;
	wire w_dff_A_jhMcZnbt2_1;
	wire w_dff_A_DnaIkzaT3_1;
	wire w_dff_A_imHxDDda9_1;
	wire w_dff_A_6hVWXkjQ6_1;
	wire w_dff_A_xTtnHCis9_1;
	wire w_dff_A_DKnsmow48_1;
	wire w_dff_A_vfyF6Ycp1_1;
	wire w_dff_A_WFpyXQE98_1;
	wire w_dff_A_aMDjTctL1_0;
	wire w_dff_A_BwJs6p1G3_0;
	wire w_dff_A_zbC3LCll8_0;
	wire w_dff_A_ejgauGLC4_0;
	wire w_dff_A_Kw3svK8O4_0;
	wire w_dff_A_mEdP1J3l8_0;
	wire w_dff_A_IfJ6Ji1l7_0;
	wire w_dff_A_0FwZ7po26_0;
	wire w_dff_A_SXzeJC4S4_0;
	wire w_dff_A_mDWta6TW9_2;
	wire w_dff_A_hHzCmzeS4_2;
	wire w_dff_A_TtGEkeY89_2;
	wire w_dff_A_K1x60O0N4_2;
	wire w_dff_A_Uarh9PFV1_2;
	wire w_dff_A_gj7lFmNP8_2;
	wire w_dff_A_RwD8JSBg5_2;
	wire w_dff_A_wT8289un0_2;
	wire w_dff_A_Xr0Kvv8Y5_2;
	wire w_dff_A_OP52JwfC9_2;
	wire w_dff_A_Y6gUf3oU0_2;
	wire w_dff_A_9AAW29E89_2;
	wire w_dff_A_6P32KFym1_2;
	wire w_dff_A_3TKcNZZK1_2;
	wire w_dff_A_D8gzYsni2_2;
	wire w_dff_A_8ITYveoI6_2;
	wire w_dff_A_2D84yOlR5_2;
	wire w_dff_A_wc0xcGdp5_2;
	wire w_dff_A_MJEHKelT9_2;
	wire w_dff_A_TpLGOVxJ3_2;
	wire w_dff_A_Sn4d4rc53_2;
	wire w_dff_A_KG0OdvOF6_2;
	wire w_dff_A_kxet5FjL6_1;
	wire w_dff_A_o5CGr2Xd1_1;
	wire w_dff_A_3Pv0tZvA9_1;
	wire w_dff_A_Luggkojh2_1;
	wire w_dff_A_bNAwkg675_1;
	wire w_dff_A_EU1Dvvx85_1;
	wire w_dff_A_VNq02SJX2_1;
	wire w_dff_A_0403zIP21_1;
	wire w_dff_A_7vdJej4w7_1;
	wire w_dff_A_ILyRnmIo6_1;
	wire w_dff_A_1FParwAR7_1;
	wire w_dff_A_MxY3InuG6_1;
	wire w_dff_A_MjDO53oV9_1;
	wire w_dff_A_TzqSrlq20_1;
	wire w_dff_A_6gXZQCVX2_1;
	wire w_dff_A_8kdbvXo36_1;
	wire w_dff_A_rBj5yH7m2_1;
	wire w_dff_A_c2wt0MIR8_1;
	wire w_dff_A_71Hv8wWq6_1;
	wire w_dff_A_PgFreHKh6_2;
	wire w_dff_A_xafjBsPZ9_2;
	wire w_dff_A_CQU9iPEY5_2;
	wire w_dff_A_DbsFcYV09_2;
	wire w_dff_A_qiPvhrsf0_2;
	wire w_dff_A_LUvOHpZi3_2;
	wire w_dff_A_OlIIpLag3_2;
	wire w_dff_A_EHiiTA7u0_2;
	wire w_dff_A_hgA0ILHc4_2;
	wire w_dff_A_y04p6kf26_2;
	wire w_dff_A_2D4206v07_2;
	wire w_dff_A_Pfca8OpW5_2;
	wire w_dff_A_MHwIKS9y3_2;
	wire w_dff_B_GcMdmMVM2_1;
	wire w_dff_B_zMZMUDlf5_1;
	wire w_dff_B_RhyuXJLF6_1;
	wire w_dff_B_WGARJiUp5_1;
	wire w_dff_B_BvxJ2Mm64_1;
	wire w_dff_B_pLeBhFNz9_1;
	wire w_dff_B_nqh3MVxB1_1;
	wire w_dff_B_dV5BTFhk1_1;
	wire w_dff_B_P2lTB8rS3_1;
	wire w_dff_B_s9tCs7Ub1_1;
	wire w_dff_B_3Y0mdJ9U4_1;
	wire w_dff_B_0eWqvDC76_1;
	wire w_dff_B_0vl2vCaa8_1;
	wire w_dff_B_lPlH5lt62_1;
	wire w_dff_B_unJ015bL8_1;
	wire w_dff_B_O2eDBG042_1;
	wire w_dff_B_BCbxBWk33_1;
	wire w_dff_B_nUzOZrMs5_1;
	wire w_dff_B_nPxXPHIc5_1;
	wire w_dff_B_YTIhUTTB4_1;
	wire w_dff_B_NOp2b5xe5_1;
	wire w_dff_B_OMqhVrpM7_1;
	wire w_dff_B_xIkb5FXp4_1;
	wire w_dff_B_B6rP9bDy7_1;
	wire w_dff_B_JVohYFZe8_1;
	wire w_dff_B_XL1w188B3_1;
	wire w_dff_B_T7AklfjQ6_1;
	wire w_dff_B_N8Qk7xNi3_1;
	wire w_dff_B_0EcG2cvJ4_1;
	wire w_dff_B_ng0t5frc6_1;
	wire w_dff_B_FXUugAvv8_1;
	wire w_dff_B_Bt6acUxp3_1;
	wire w_dff_B_Iv9TBwiM1_1;
	wire w_dff_B_R82TuCAp8_1;
	wire w_dff_B_jFKLyiBR8_1;
	wire w_dff_B_r52Jz6kg4_1;
	wire w_dff_B_6CDC7SuT2_1;
	wire w_dff_B_GNiAnel13_1;
	wire w_dff_B_bH3FXHlC6_1;
	wire w_dff_B_FOs56RDq4_1;
	wire w_dff_B_W4xFd2Mv8_1;
	wire w_dff_B_DWwOLS1p7_1;
	wire w_dff_B_tB2tv4WR3_1;
	wire w_dff_B_ccUhAJav5_1;
	wire w_dff_B_MI2lEjEz8_1;
	wire w_dff_B_CpST3Fer2_0;
	wire w_dff_B_LxWmpUSM6_0;
	wire w_dff_B_pZcb0Kqh3_0;
	wire w_dff_B_q5nww98O8_0;
	wire w_dff_B_vqc6fzrr5_0;
	wire w_dff_B_OeVZYOW70_0;
	wire w_dff_B_SdjibiUX6_0;
	wire w_dff_B_iqEsNM4v1_0;
	wire w_dff_B_MTRkLikJ2_0;
	wire w_dff_B_ofABOZhb3_0;
	wire w_dff_B_fvXc74ma0_0;
	wire w_dff_B_AQRQ9Uxa9_0;
	wire w_dff_B_HGhr1ADv1_0;
	wire w_dff_B_MGkbql5G1_0;
	wire w_dff_B_mN4fDTrq4_0;
	wire w_dff_B_Azu6K8Sc3_0;
	wire w_dff_B_7pOQs7l51_0;
	wire w_dff_B_GpEUyCfx2_0;
	wire w_dff_B_g7SLLSYW6_0;
	wire w_dff_B_eSIga0pe3_0;
	wire w_dff_B_IrUnlNG80_0;
	wire w_dff_B_gMDbBuhw1_0;
	wire w_dff_B_eDYGrcpj3_0;
	wire w_dff_B_ryH6SxkN9_0;
	wire w_dff_B_r5rBMJ1U1_0;
	wire w_dff_B_oL51l6mP4_0;
	wire w_dff_B_wySAC3OF1_0;
	wire w_dff_B_Z6XkuS7b3_0;
	wire w_dff_B_zU9xVylp3_1;
	wire w_dff_B_3bQpT2b02_1;
	wire w_dff_B_h6IJkdMG1_1;
	wire w_dff_A_cCAn80oG9_0;
	wire w_dff_B_wFu7iZoY4_1;
	wire w_dff_B_fbBXViZA9_1;
	wire w_dff_A_H8tCWae42_1;
	wire w_dff_B_JZ7huyEY5_0;
	wire w_dff_A_iuRPSOYI0_0;
	wire w_dff_B_29o6Iq4y3_1;
	wire w_dff_A_Unoy0Uw58_0;
	wire w_dff_B_FbiuPYQL1_2;
	wire w_dff_A_N3JHm29S7_0;
	wire w_dff_A_GPJO0iP97_0;
	wire w_dff_A_c0cF66of2_0;
	wire w_dff_B_KuVIetra4_1;
	wire w_dff_B_OkaoFZ6D5_1;
	wire w_dff_B_qItMzJlr6_1;
	wire w_dff_A_XoUV0c5b2_1;
	wire w_dff_B_U9CtPUDe4_1;
	wire w_dff_B_eFO82afY2_1;
	wire w_dff_A_3iL9ABnu6_1;
	wire w_dff_B_nmS8vhuX1_1;
	wire w_dff_A_pcFGW0Pn6_0;
	wire w_dff_A_Laqa2d835_0;
	wire w_dff_A_2mXuuQ4Y2_0;
	wire w_dff_A_2g984dOy4_1;
	wire w_dff_A_ufLtg2qa8_1;
	wire w_dff_A_9GU07UWk6_1;
	wire w_dff_A_vrKrY8cu5_1;
	wire w_dff_A_i6YE0F3L3_1;
	wire w_dff_A_G2mtEQOr2_1;
	wire w_dff_A_U2mXfd1S2_1;
	wire w_dff_A_8fGymNBb2_1;
	wire w_dff_A_ECjd5M5B9_1;
	wire w_dff_A_Q38jjBbW6_1;
	wire w_dff_A_8i6JpYol0_1;
	wire w_dff_A_0Z3Tn8FY6_1;
	wire w_dff_B_oJvbEFDl0_0;
	wire w_dff_A_JPKQlNbV4_0;
	wire w_dff_A_ABbQpe6u2_0;
	wire w_dff_B_6FG4Q1yi3_0;
	wire w_dff_B_6rVycu836_0;
	wire w_dff_B_YUJFSNRH8_0;
	wire w_dff_B_IsU0fbo28_1;
	wire w_dff_B_jVmOc66Q0_1;
	wire w_dff_B_rQR8s6aN8_1;
	wire w_dff_A_N6FBxErh3_0;
	wire w_dff_A_khXuzogl9_0;
	wire w_dff_A_c21A9dki1_0;
	wire w_dff_A_5Foc6wzG5_0;
	wire w_dff_A_srcgfnHl6_0;
	wire w_dff_A_cpKxORtp9_0;
	wire w_dff_A_9PnZh8QN7_0;
	wire w_dff_A_pxtAKnMq3_0;
	wire w_dff_B_Pwwn9wzk7_1;
	wire w_dff_B_GQA8Bv4Z2_1;
	wire w_dff_B_68DvjMJx9_0;
	wire w_dff_B_94lpjmqD7_0;
	wire w_dff_A_4tImIQIC6_0;
	wire w_dff_B_ZdQHdSHF7_1;
	wire w_dff_A_rJLsUqjl8_2;
	wire w_dff_A_ZBOaviyN3_2;
	wire w_dff_A_ZlM4TwFe9_0;
	wire w_dff_A_9qjiZtE58_0;
	wire w_dff_A_0UXFHcve6_0;
	wire w_dff_A_UsjWnzyx7_0;
	wire w_dff_A_Zmwi3UTf3_1;
	wire w_dff_B_YcEiYVfb1_3;
	wire w_dff_B_4iQ1YXwM3_3;
	wire w_dff_A_CMqfPapT7_1;
	wire w_dff_A_9olhZSYh5_1;
	wire w_dff_A_fr8kjHLB5_1;
	wire w_dff_A_QSN4LlY07_1;
	wire w_dff_A_UsqvMGoB4_1;
	wire w_dff_A_NKahmuzI0_1;
	wire w_dff_A_qWlyI1sH6_2;
	wire w_dff_A_mGAL2BkJ7_2;
	wire w_dff_A_A9HHPL6c9_2;
	wire w_dff_A_9ogfngCa2_2;
	wire w_dff_A_XVAy8ZRa0_2;
	wire w_dff_A_FRIHcNj08_2;
	wire w_dff_A_igeem2lH7_2;
	wire w_dff_A_3JeCS0Rb0_1;
	wire w_dff_A_tGz2ldo26_1;
	wire w_dff_A_Aj2wo3kE8_1;
	wire w_dff_A_uNBldFdh9_1;
	wire w_dff_A_jWl5fsZ09_1;
	wire w_dff_A_4U3jWDXQ1_1;
	wire w_dff_A_sFUW312X0_2;
	wire w_dff_A_fdxC9CnN2_2;
	wire w_dff_A_qMHXqdRa3_2;
	wire w_dff_A_w7MUFPIP6_0;
	wire w_dff_B_rGgM8vH17_1;
	wire w_dff_A_pph0MgxZ3_0;
	wire w_dff_B_aMolQQ517_1;
	wire w_dff_B_HoeLbVlP7_1;
	wire w_dff_B_gjHkMSii5_1;
	wire w_dff_B_WS7nlbgh7_1;
	wire w_dff_B_EPT7mUVs7_1;
	wire w_dff_A_IotwBgAe4_2;
	wire w_dff_A_fIBMuMh99_2;
	wire w_dff_A_FbaP9dS96_2;
	wire w_dff_A_j6HjCMk69_2;
	wire w_dff_A_tSJb9xXv4_2;
	wire w_dff_A_lpXRusux6_2;
	wire w_dff_A_Z1cv1RsF6_2;
	wire w_dff_A_VJ4feSW02_2;
	wire w_dff_A_oZ9B3eiY8_2;
	wire w_dff_A_amKvZqLm9_2;
	wire w_dff_A_fb2ZOYWl2_2;
	wire w_dff_A_TOnJGDtJ1_2;
	wire w_dff_A_Fi3ptPpt7_2;
	wire w_dff_A_fh4gxAWV4_2;
	wire w_dff_A_H7atk1yL6_2;
	wire w_dff_A_p6IIo7T53_1;
	wire w_dff_A_ZuXyQCnJ5_1;
	wire w_dff_A_eKvoSu1N5_1;
	wire w_dff_A_KKEvQSj34_1;
	wire w_dff_A_D4pdAtop8_1;
	wire w_dff_A_FJSxXbdl7_1;
	wire w_dff_A_xpvPGOKX5_1;
	wire w_dff_A_D3jclvVg1_1;
	wire w_dff_A_HyqSYiZF9_1;
	wire w_dff_A_VwbmPG1e6_1;
	wire w_dff_B_9fuAt7GB5_1;
	wire w_dff_B_lUK1UlOm6_1;
	wire w_dff_B_WPPJIrq28_1;
	wire w_dff_B_qr4C19tO9_1;
	wire w_dff_B_GRuNwgC55_1;
	wire w_dff_B_NrtkYxHm3_1;
	wire w_dff_B_2IxeBqju2_1;
	wire w_dff_A_iSB1yla53_1;
	wire w_dff_B_SRgyzuye7_1;
	wire w_dff_B_B3B9hQjx5_1;
	wire w_dff_B_6y5gUE284_1;
	wire w_dff_B_hrLyDgLw7_1;
	wire w_dff_B_IFUxW3UB8_1;
	wire w_dff_B_NeZtH99f4_1;
	wire w_dff_B_PzqaW83H4_1;
	wire w_dff_A_9EaeI22C0_1;
	wire w_dff_A_hZ5D2cD50_1;
	wire w_dff_A_NcYLiKqL2_0;
	wire w_dff_A_ANjvwgwf4_0;
	wire w_dff_A_mxHttHXo8_0;
	wire w_dff_A_ci6v7xUY3_0;
	wire w_dff_A_yEJUWmDc9_1;
	wire w_dff_A_qUeNlPd81_1;
	wire w_dff_A_ITtg9bl70_2;
	wire w_dff_B_XnDd9siy9_3;
	wire w_dff_A_vnwryK2G1_0;
	wire w_dff_A_hAlFR93x7_0;
	wire w_dff_A_jEfd3TcK5_0;
	wire w_dff_A_YX2znO8M5_1;
	wire w_dff_A_gOqqgfa46_1;
	wire w_dff_A_DisGo5P51_2;
	wire w_dff_B_8Q3FfvoL7_3;
	wire w_dff_B_pbMff5Cz1_3;
	wire w_dff_B_POX1SfP90_3;
	wire w_dff_B_VnSme4hm7_3;
	wire w_dff_B_80wDeluw5_3;
	wire w_dff_B_BoJPt3mV0_3;
	wire w_dff_B_zcciXxZc3_3;
	wire w_dff_B_4vv7aUqS2_3;
	wire w_dff_B_bPFowCxE0_3;
	wire w_dff_B_X9d1K3tK5_3;
	wire w_dff_A_eJBzFm3K3_0;
	wire w_dff_A_1fyaFBeA8_0;
	wire w_dff_A_5UZS9S6D2_0;
	wire w_dff_A_n2wbnxKo6_0;
	wire w_dff_A_1dsQ5K8h8_0;
	wire w_dff_A_riFO6sSa8_0;
	wire w_dff_A_N3lgVb1j0_0;
	wire w_dff_A_fWXMmo2N7_0;
	wire w_dff_A_DaPhHxza4_0;
	wire w_dff_A_13B4Nrks8_0;
	wire w_dff_A_gZ5FYZpZ7_0;
	wire w_dff_A_YPSpdvYW5_0;
	wire w_dff_A_iO8l3Xcp1_0;
	wire w_dff_A_2wygWxmI5_1;
	wire w_dff_A_eY4OjLz98_1;
	wire w_dff_A_tr02KA827_1;
	wire w_dff_A_hXEBdvMU1_1;
	wire w_dff_A_XdB1QHq36_1;
	wire w_dff_A_kTLuUohm9_1;
	wire w_dff_A_ntI7QtOM7_1;
	wire w_dff_A_DtcriHOY9_1;
	wire w_dff_A_eAAHlm9e9_1;
	wire w_dff_A_inQvp69a0_1;
	wire w_dff_A_FPsJvK3N9_0;
	wire w_dff_B_sagk3Rbh6_0;
	wire w_dff_B_JPQ5n1MR2_0;
	wire w_dff_A_VjKBCpmZ8_0;
	wire w_dff_A_1mMfmRST8_0;
	wire w_dff_A_Mpz7Wox11_0;
	wire w_dff_B_4XfIYN468_2;
	wire w_dff_A_lLMQcsDI1_0;
	wire w_dff_A_mYnJAxXX6_0;
	wire w_dff_A_Knhhl1uN2_0;
	wire w_dff_A_HEhayoAF5_1;
	wire w_dff_A_Mm1K6Wtr8_1;
	wire w_dff_A_9nVqtLlm0_1;
	wire w_dff_A_HIQsbQFI5_1;
	wire w_dff_A_5s9HAUx73_1;
	wire w_dff_A_aWOUgwhr9_1;
	wire w_dff_A_TLALxBQU3_1;
	wire w_dff_A_b3hINvNF7_1;
	wire w_dff_A_q5eO7kLE9_0;
	wire w_dff_A_nnT4j9Jv7_0;
	wire w_dff_A_AL058DZw2_0;
	wire w_dff_A_908jh8XE2_0;
	wire w_dff_A_IIOM7Qkz1_2;
	wire w_dff_A_zyvbQmbi4_2;
	wire w_dff_A_G0NBzf615_1;
	wire w_dff_A_suv6ryfC7_1;
	wire w_dff_A_YnTQFQCz7_1;
	wire w_dff_A_KJtXCf6k5_1;
	wire w_dff_A_AGM8M7Sv0_1;
	wire w_dff_B_jb0y8H540_1;
	wire w_dff_B_w5V504Yr2_1;
	wire w_dff_A_plH1km8d8_1;
	wire w_dff_A_RWh6EijB0_1;
	wire w_dff_A_KxjkrfVe2_1;
	wire w_dff_A_wBrxynoD4_1;
	wire w_dff_A_sWBYShcs2_1;
	wire w_dff_A_sztsfTGm4_1;
	wire w_dff_A_h2ENW0g59_1;
	wire w_dff_B_yFdrxyFS0_0;
	wire w_dff_B_jWYeyIKN8_1;
	wire w_dff_A_6KzOBrkF1_2;
	wire w_dff_A_UgdAQFHI9_1;
	wire w_dff_A_nWJxO2Ho7_1;
	wire w_dff_A_mbyb7jcW9_1;
	wire w_dff_A_zutWcC9k7_1;
	wire w_dff_A_rKzJjZLt6_2;
	wire w_dff_A_aD3rUtgm9_2;
	wire w_dff_A_fIw77XNS0_2;
	wire w_dff_A_ZvPz6YQa3_2;
	wire w_dff_A_dQzCsD9g8_0;
	wire w_dff_A_v3GcPNiR7_0;
	wire w_dff_B_vw3vRAA64_3;
	wire w_dff_A_HWxL4K037_0;
	wire w_dff_B_4pBthudu4_1;
	wire w_dff_B_TkDvYJKb3_1;
	wire w_dff_A_CRbXyWah2_0;
	wire w_dff_A_VNOLxWZW2_0;
	wire w_dff_B_ONHJmS7E4_2;
	wire w_dff_A_FXZqEKHe9_0;
	wire w_dff_A_GmEHFD3f9_0;
	wire w_dff_A_HdGKWoCy4_0;
	wire w_dff_A_77MecEph4_1;
	wire w_dff_A_W8er2Mim7_1;
	wire w_dff_A_DMdqylml7_1;
	wire w_dff_A_aYMbA9d67_1;
	wire w_dff_A_xJZG6co13_1;
	wire w_dff_A_ltIQVsce8_1;
	wire w_dff_A_Pdohg5pg3_1;
	wire w_dff_A_K3cruJ2w0_2;
	wire w_dff_A_DI0ckUu57_2;
	wire w_dff_A_qpfmLGMv9_2;
	wire w_dff_A_Azp1elas1_2;
	wire w_dff_A_z5GEAU9j4_2;
	wire w_dff_B_LqUkf7YI2_0;
	wire w_dff_B_TZ9GQanc9_1;
	wire w_dff_A_AHXN0R4U7_0;
	wire w_dff_A_mio5KJpD3_1;
	wire w_dff_B_sQM3zmHS5_1;
	wire w_dff_A_GtdLA4qw5_0;
	wire w_dff_A_ShosyFsw9_1;
	wire w_dff_A_vKyo0vsz3_1;
	wire w_dff_B_D4YMhMGO0_1;
	wire w_dff_A_zCn3yGKH3_0;
	wire w_dff_A_X7X2iXnx4_0;
	wire w_dff_A_z476YpM93_2;
	wire w_dff_A_Dy7yROMc0_0;
	wire w_dff_A_IJzczlmd7_0;
	wire w_dff_A_uudzYH4a6_0;
	wire w_dff_A_DIDKx7dg3_2;
	wire w_dff_A_4Jm7U9iH9_0;
	wire w_dff_A_2JWxP9z98_1;
	wire w_dff_A_mPKOD2o62_2;
	wire w_dff_A_RsPkIsbe4_0;
	wire w_dff_A_LADkelDj8_0;
	wire w_dff_A_zizoQuCR7_0;
	wire w_dff_A_DMbad3hU7_2;
	wire w_dff_A_JGbEjWLn7_2;
	wire w_dff_A_OxQjbA5L0_2;
	wire w_dff_A_BDpeNNmD2_0;
	wire w_dff_A_X7ZMSWaE8_0;
	wire w_dff_A_FIfD5XyQ4_0;
	wire w_dff_A_MtyJ4roH9_1;
	wire w_dff_A_ckaHTcbS1_1;
	wire w_dff_A_E8mdAG5M9_2;
	wire w_dff_A_DrDwCHlH4_0;
	wire w_dff_A_xx4rnksF6_2;
	wire w_dff_B_5144iDOd1_3;
	wire w_dff_A_0RiWWR2i3_0;
	wire w_dff_A_nwJKUgmw2_0;
	wire w_dff_A_a1pkJkDq3_0;
	wire w_dff_A_cCHYyOHs7_1;
	wire w_dff_A_VpVhB3k29_1;
	wire w_dff_A_5Ds71fVU2_1;
	wire w_dff_A_hrEhE4iP4_1;
	wire w_dff_A_zh3jNfwi9_1;
	wire w_dff_A_06pQuPHL0_1;
	wire w_dff_A_6DzUmaNR4_2;
	wire w_dff_A_X3m6gHGT3_2;
	wire w_dff_A_vVYz0nIU7_2;
	wire w_dff_A_j7HvhEyZ8_1;
	wire w_dff_A_ezuIGCO32_1;
	wire w_dff_A_62MADGjn5_1;
	wire w_dff_A_dMeO5M2X8_1;
	wire w_dff_A_mqI9zWK44_1;
	wire w_dff_A_77yJpoSn1_1;
	wire w_dff_A_Hcj920qD0_1;
	wire w_dff_A_qZvNo7G69_1;
	wire w_dff_A_ysBaB5zn3_1;
	wire w_dff_A_Su4vCRfa8_1;
	wire w_dff_A_Q12d3uM86_1;
	wire w_dff_A_IPcIksHL9_0;
	wire w_dff_A_ffhFOXib9_0;
	wire w_dff_A_4vW2gdeH9_0;
	wire w_dff_A_QJgWHiKz1_2;
	wire w_dff_A_rAA9UwGv7_1;
	wire w_dff_A_SXdVppZN2_1;
	wire w_dff_A_RkwJ56zm0_1;
	wire w_dff_A_qoh4vhNv1_1;
	wire w_dff_A_nh51Fih91_1;
	wire w_dff_A_y7muOgyZ4_1;
	wire w_dff_A_3DNjikiI9_1;
	wire w_dff_A_QZDGlfHh3_1;
	wire w_dff_A_UnSMDFQx4_1;
	wire w_dff_B_XT6WQqUp7_0;
	wire w_dff_A_1BDoj2j67_1;
	wire w_dff_A_UNfn2Mjz9_1;
	wire w_dff_A_ws0VB4db8_2;
	wire w_dff_A_804CLJld9_0;
	wire w_dff_A_qAHGF4p58_0;
	wire w_dff_A_Zje9Avjg1_0;
	wire w_dff_A_zj7BXK0S0_0;
	wire w_dff_A_yshMyeTV6_2;
	wire w_dff_A_tnwJ9HxF4_2;
	wire w_dff_A_zPkn3j5y7_0;
	wire w_dff_A_fpMLpCsI5_0;
	wire w_dff_A_eybolzBm1_0;
	wire w_dff_A_9yck677m1_0;
	wire w_dff_A_ipuRDokf7_0;
	wire w_dff_A_h0ySRBKO7_0;
	wire w_dff_A_snFo9xDQ4_0;
	wire w_dff_A_8BKRwdoV7_0;
	wire w_dff_A_gBj7XBNV9_0;
	wire w_dff_A_La1cuWoT6_0;
	wire w_dff_A_hhz5Finv0_0;
	wire w_dff_A_um0Y8Tlh3_0;
	wire w_dff_A_dXCQTO4B1_0;
	wire w_dff_A_8XkyozXV8_0;
	wire w_dff_A_5AjmUA0r5_0;
	wire w_dff_A_8cAvl1RM6_0;
	wire w_dff_A_6FZFw8Wn2_0;
	wire w_dff_A_UMb2lxUr7_0;
	wire w_dff_A_UThKjtyT3_0;
	wire w_dff_A_B5jVEXVJ8_0;
	wire w_dff_A_IyFtmgwg1_2;
	wire w_dff_A_93sZyrYH7_2;
	wire w_dff_A_vwpPry2y5_2;
	wire w_dff_A_MqQyiEH24_2;
	wire w_dff_B_BkxlJdZ46_0;
	wire w_dff_B_O0ZUx5wi3_0;
	wire w_dff_B_WxdPq4aF7_0;
	wire w_dff_B_NHCck5hr7_0;
	wire w_dff_B_C8rDAqsc1_0;
	wire w_dff_B_0ap6VvY94_0;
	wire w_dff_B_YK1nnchb2_0;
	wire w_dff_B_vX0LSfgT8_0;
	wire w_dff_B_6kJ1aIoB0_0;
	wire w_dff_B_WPfkaipq5_0;
	wire w_dff_B_gGWEjK925_0;
	wire w_dff_B_KOiFVQEN6_0;
	wire w_dff_B_0wk7J7iX9_0;
	wire w_dff_B_sZlIW0VD8_0;
	wire w_dff_B_j3rZniwi8_0;
	wire w_dff_B_uq0MPfYp7_0;
	wire w_dff_B_vDw7soEk5_0;
	wire w_dff_B_vZOAtpMZ1_0;
	wire w_dff_B_d5vIGQs41_0;
	wire w_dff_B_ZqXl24ZW1_1;
	wire w_dff_B_uC3bIeM93_1;
	wire w_dff_B_MWJj8SXT8_1;
	wire w_dff_B_XZAIPmcT9_1;
	wire w_dff_B_xleXgPAa7_1;
	wire w_dff_B_lMMR4Cfn6_1;
	wire w_dff_B_CFUSpfow9_1;
	wire w_dff_B_tiupQjuw9_1;
	wire w_dff_B_bScsnL8T1_1;
	wire w_dff_B_ibd6MUij4_1;
	wire w_dff_A_5n6wNkML4_2;
	wire w_dff_A_7ToaC0wk1_2;
	wire w_dff_A_P4SEEAWN6_1;
	wire w_dff_B_CIh7LDlr1_0;
	wire w_dff_B_FsANhX6v6_1;
	wire w_dff_B_K0LZ4egM2_1;
	wire w_dff_B_DnPGAQ225_1;
	wire w_dff_B_QfmQDYsv4_1;
	wire w_dff_B_HtBxJ4xT0_1;
	wire w_dff_B_mlib1XFp3_1;
	wire w_dff_B_cWMUahs32_1;
	wire w_dff_B_LNpshacK4_0;
	wire w_dff_B_d5zF6k0X1_0;
	wire w_dff_A_psAXok7z0_1;
	wire w_dff_A_GAH6Qt1h4_1;
	wire w_dff_A_F8gxj0VY4_1;
	wire w_dff_A_WSsWGxBs5_1;
	wire w_dff_A_hEztNyTD8_1;
	wire w_dff_A_CXmnyfZQ8_1;
	wire w_dff_A_Jx6W1WJ93_1;
	wire w_dff_A_zLeIUgkS0_1;
	wire w_dff_A_NN3yA7u52_1;
	wire w_dff_A_eDMU0LZO7_1;
	wire w_dff_A_xBIqZVoy4_1;
	wire w_dff_A_HOxDukn92_1;
	wire w_dff_A_m7ftWT6w2_1;
	wire w_dff_B_85atRmAC4_2;
	wire w_dff_A_wMsnKMJ88_2;
	wire w_dff_A_uoeP3skZ5_2;
	wire w_dff_A_yNVUy8E48_2;
	wire w_dff_A_WbG1ljAS0_2;
	wire w_dff_A_BN6ZpJxo8_2;
	wire w_dff_B_Geu16LN10_1;
	wire w_dff_B_A6Ci5U740_1;
	wire w_dff_B_18LzI1ED4_1;
	wire w_dff_B_ZWyfy5xQ9_1;
	wire w_dff_B_6oCEeYCx3_1;
	wire w_dff_A_gGvEFFCe5_1;
	wire w_dff_A_i3QuapY35_1;
	wire w_dff_A_rfj2WLJI8_1;
	wire w_dff_A_ROlElPWS5_1;
	wire w_dff_A_RQf5Tvz91_1;
	wire w_dff_A_kLRNieab5_1;
	wire w_dff_A_fNtva72h0_1;
	wire w_dff_A_aglSFw1X4_0;
	wire w_dff_A_tCBNZm7E8_0;
	wire w_dff_A_HHfVC22M3_0;
	wire w_dff_A_066BfeTR1_0;
	wire w_dff_A_Z1WB7ngR6_0;
	wire w_dff_A_RyoELTp12_0;
	wire w_dff_A_ZML9gGz17_0;
	wire w_dff_A_UVhmSwRi2_0;
	wire w_dff_A_zw6mIUv48_0;
	wire w_dff_A_4TkgQVI47_0;
	wire w_dff_A_W8pUR8FL8_0;
	wire w_dff_A_AcJYINxx4_0;
	wire w_dff_A_ExtVVazX9_0;
	wire w_dff_A_GFxP12ni9_0;
	wire w_dff_A_07Q4LIuX7_0;
	wire w_dff_A_1LHGQENa9_0;
	wire w_dff_A_ufo0E6sZ2_0;
	wire w_dff_B_FpG3zss28_2;
	wire w_dff_B_Y8KYvAO46_2;
	wire w_dff_A_bZFrhxba1_1;
	wire w_dff_A_ieECgFmf2_1;
	wire w_dff_A_aiAFb0Bb7_1;
	wire w_dff_A_WU2MSFyF2_1;
	wire w_dff_A_OCMk77wF2_1;
	wire w_dff_A_DpDS1xpR7_1;
	wire w_dff_A_tMLLDGjh3_1;
	wire w_dff_A_DcebTOye1_1;
	wire w_dff_A_LtRWGmHs8_1;
	wire w_dff_A_RpA6Tcj95_1;
	wire w_dff_A_T3e2k0WO5_2;
	wire w_dff_B_D4fOFHL32_0;
	wire w_dff_B_WRS1WKld4_1;
	wire w_dff_A_hBJz7Zz76_0;
	wire w_dff_A_eLuM00936_2;
	wire w_dff_A_SvbF4Bdf8_2;
	wire w_dff_A_1NICf9Y90_2;
	wire w_dff_A_aRbml7jY4_2;
	wire w_dff_B_KjkXO6uF3_1;
	wire w_dff_B_2HPg2p4d3_1;
	wire w_dff_A_soHz0zdW4_0;
	wire w_dff_A_BuuBg4Y98_0;
	wire w_dff_A_vvtsNuvE8_0;
	wire w_dff_A_tHGNU3MT1_2;
	wire w_dff_A_aGjrNP4F6_2;
	wire w_dff_A_MmMhsMmR4_2;
	wire w_dff_A_1zbcjddR5_2;
	wire w_dff_A_aMve6OvM1_2;
	wire w_dff_A_ZZpAA2XQ4_2;
	wire w_dff_A_ccdkAcaE8_2;
	wire w_dff_B_bA6fv7q99_2;
	wire w_dff_A_Hkcjyptd3_1;
	wire w_dff_B_4gpgBaTR1_0;
	wire w_dff_B_RwubvhTj3_1;
	wire w_dff_B_vL2FhdQC8_0;
	wire w_dff_B_cgsVAW2z9_1;
	wire w_dff_A_Bq7f18HZ2_1;
	wire w_dff_A_mHZ70Jib2_0;
	wire w_dff_A_m5S8r6zo1_0;
	wire w_dff_B_DMsN892w7_2;
	wire w_dff_B_xHtQRvQv8_2;
	wire w_dff_B_FTkfTvPN9_2;
	wire w_dff_A_kz7MEoVC4_0;
	wire w_dff_A_nvuB8LKZ9_0;
	wire w_dff_A_0oBK8ZAp0_0;
	wire w_dff_A_N5RCJTb54_0;
	wire w_dff_A_URK2xtwG4_1;
	wire w_dff_A_rEhQI14U6_1;
	wire w_dff_A_LxSrrlcH4_1;
	wire w_dff_A_KeuITP3b5_1;
	wire w_dff_A_qF7txXay8_1;
	wire w_dff_A_5USy8GVJ0_1;
	wire w_dff_A_lJZaxkb85_2;
	wire w_dff_A_xW9fUiXb0_2;
	wire w_dff_A_QPI551Ni1_2;
	wire w_dff_A_rfz3GYIR9_2;
	wire w_dff_A_olY8EaMS8_2;
	wire w_dff_A_5VPYhO5W0_2;
	wire w_dff_B_nyBQTdjM8_0;
	wire w_dff_B_6PRfqFmm3_0;
	wire w_dff_B_E2p7tr5q6_0;
	wire w_dff_B_nbXMw3Mw3_0;
	wire w_dff_B_2cukDi5m9_0;
	wire w_dff_B_9tz4d4xd9_0;
	wire w_dff_B_tBGgbLg64_0;
	wire w_dff_B_SOO4Pp8b8_0;
	wire w_dff_B_Kf66Vzf82_0;
	wire w_dff_B_2psLhj9J6_0;
	wire w_dff_B_saGac2ra0_0;
	wire w_dff_B_UNIAtMf36_1;
	wire w_dff_B_9OsZINS98_1;
	wire w_dff_B_7lVXvREL6_1;
	wire w_dff_A_iKgtqary5_0;
	wire w_dff_A_pDMn4PWS6_0;
	wire w_dff_B_TGZRu1Wg8_2;
	wire w_dff_B_9t6qxJNc1_2;
	wire w_dff_B_rrJ8SN4V1_2;
	wire w_dff_B_GDBc4ZsU0_2;
	wire w_dff_B_X4yL09Gx8_2;
	wire w_dff_B_uYtmjByw1_2;
	wire w_dff_B_nXFOZ9vY9_2;
	wire w_dff_B_MLAzN9QG9_2;
	wire w_dff_B_Z8maTnec1_2;
	wire w_dff_B_eMhbkInQ9_2;
	wire w_dff_B_4180wa9x2_2;
	wire w_dff_B_r7JxUxaj9_2;
	wire w_dff_A_4uMTWYY66_0;
	wire w_dff_A_teNYVAXO2_0;
	wire w_dff_A_85z2pYkP1_0;
	wire w_dff_A_Zur9GXe36_0;
	wire w_dff_A_skKNapTl4_0;
	wire w_dff_A_UBVNAlgo3_0;
	wire w_dff_A_N8BJuBMI5_0;
	wire w_dff_A_Yrw8BFI23_0;
	wire w_dff_A_gqBH0egq3_0;
	wire w_dff_A_83IIzFRi1_0;
	wire w_dff_A_mfaNR6rt2_0;
	wire w_dff_A_TEOkXkTo7_0;
	wire w_dff_A_h9CeMrqq8_0;
	wire w_dff_A_0lGGwlJU3_0;
	wire w_dff_A_ezjoubcI2_0;
	wire w_dff_A_cPARA59N3_1;
	wire w_dff_A_R1FXdyIR7_1;
	wire w_dff_A_1njxCRKP6_1;
	wire w_dff_A_p9fMp0Yu5_1;
	wire w_dff_A_98tYvckP5_1;
	wire w_dff_A_rkkqxecX0_1;
	wire w_dff_A_wEkh6VZ99_1;
	wire w_dff_A_pv1zHmMR5_1;
	wire w_dff_A_qmZQARQv9_1;
	wire w_dff_A_kOZ4e30O9_1;
	wire w_dff_A_HGOM2LJm0_1;
	wire w_dff_A_EP0AG1Mv3_1;
	wire w_dff_B_1UoxQOPg5_1;
	wire w_dff_B_gjBGjyHe4_1;
	wire w_dff_B_3qSVlTZF9_0;
	wire w_dff_B_H6WJMbzw8_0;
	wire w_dff_B_1WSuVNJs3_0;
	wire w_dff_B_s5FvmlJb1_0;
	wire w_dff_A_jRI9t6sW0_0;
	wire w_dff_A_FcJRNiM37_0;
	wire w_dff_A_pY7wjSMf9_0;
	wire w_dff_A_xpLZ6p1m0_0;
	wire w_dff_A_NENDBLe24_0;
	wire w_dff_A_PPDwXgPR8_0;
	wire w_dff_A_hfb1qTpJ0_2;
	wire w_dff_A_yIo3iudj5_2;
	wire w_dff_A_VkK6Io6I5_2;
	wire w_dff_A_WL1htVC61_2;
	wire w_dff_A_oJqkeyL69_2;
	wire w_dff_A_SdP4WpJM4_1;
	wire w_dff_A_0XO0nWKt9_1;
	wire w_dff_A_2M7lTDwp8_1;
	wire w_dff_A_LMNkz2cr9_1;
	wire w_dff_B_fmvCkGY62_0;
	wire w_dff_B_X5fR3mvU3_1;
	wire w_dff_B_GBYNEvny9_1;
	wire w_dff_B_fTIeKDWs3_1;
	wire w_dff_B_SkzEZ1708_1;
	wire w_dff_B_W85vc1fY2_1;
	wire w_dff_B_bYjTbIzm8_1;
	wire w_dff_A_xnNU7dEY7_1;
	wire w_dff_A_dSuVNv8h2_1;
	wire w_dff_A_64xSURsP6_1;
	wire w_dff_A_TvANIoqV8_1;
	wire w_dff_A_yyqZ9IIT8_1;
	wire w_dff_A_wgGvhUbi2_1;
	wire w_dff_A_1VkHJzJt5_1;
	wire w_dff_A_O9Os1Fyr6_0;
	wire w_dff_A_wABGtHPL5_0;
	wire w_dff_A_E7y64BeT8_1;
	wire w_dff_A_rxH08Yi38_1;
	wire w_dff_A_jnfhIwPP8_2;
	wire w_dff_A_KwXpfViK5_2;
	wire w_dff_A_kTB2hiAI9_2;
	wire w_dff_A_1OUAiVoj1_2;
	wire w_dff_B_U3UaKWHr1_0;
	wire w_dff_B_7BuA7NsW1_1;
	wire w_dff_A_2vTjOU3w6_1;
	wire w_dff_A_iC3wlEyD1_1;
	wire w_dff_A_RRDptfXs3_0;
	wire w_dff_A_8aoAnBKr2_0;
	wire w_dff_B_90XiUeBv2_0;
	wire w_dff_B_7FjASU305_0;
	wire w_dff_B_xFYDrjga7_0;
	wire w_dff_A_3SbmSsG54_0;
	wire w_dff_A_iThb78dO1_1;
	wire w_dff_A_0hLVK2JU2_1;
	wire w_dff_B_ZNUr6u3F5_1;
	wire w_dff_A_OMQ6DNjv3_0;
	wire w_dff_A_YkubTpUK1_1;
	wire w_dff_A_jlXW2jXy4_1;
	wire w_dff_B_2qOmZ1NT3_1;
	wire w_dff_A_ASeZkNt49_0;
	wire w_dff_A_FyyMCPEK9_0;
	wire w_dff_A_TQ7VFzdl0_1;
	wire w_dff_B_npbHaFo88_1;
	wire w_dff_A_IWEv4cNs6_0;
	wire w_dff_A_U0oiwZ160_0;
	wire w_dff_A_VXalCOdH3_0;
	wire w_dff_A_ehmpgBWb6_1;
	wire w_dff_B_5xHzJPFB5_1;
	wire w_dff_A_UsLowW160_0;
	wire w_dff_A_7TY8sx288_0;
	wire w_dff_A_PEoHeZnd2_0;
	wire w_dff_B_9vqikBI63_0;
	wire w_dff_B_qcI4xhpd3_1;
	wire w_dff_B_1M5Qhs089_1;
	wire w_dff_A_YTqdcaIL5_0;
	wire w_dff_A_pNIdrQYI2_1;
	wire w_dff_A_N1aipDxO8_1;
	wire w_dff_B_MEJV5t838_3;
	wire w_dff_A_akd0nIm96_0;
	wire w_dff_A_D4p2fYwl0_0;
	wire w_dff_A_HIrzIPQQ3_0;
	wire w_dff_A_5NXR3OFP8_0;
	wire w_dff_A_TT2Fd5ad6_1;
	wire w_dff_A_05JR57BF6_1;
	wire w_dff_A_U8qclugG4_1;
	wire w_dff_A_92iJuFfX5_1;
	wire w_dff_A_dUzOfJsY5_1;
	wire w_dff_A_oskN5ta20_1;
	wire w_dff_A_IGdw9cT14_2;
	wire w_dff_A_ie5uQqXi4_2;
	wire w_dff_A_atSMxOPA5_2;
	wire w_dff_A_2y2w50oe2_2;
	wire w_dff_A_kvwfYG590_2;
	wire w_dff_B_9Ce1NkLg6_1;
	wire w_dff_A_6Kekg5Mn7_0;
	wire w_dff_A_ZABLnUU79_1;
	wire w_dff_A_T9ZByXAe4_1;
	wire w_dff_B_tNG1fmo45_3;
	wire w_dff_A_vk3DHFRB9_0;
	wire w_dff_A_KrTo8HK52_0;
	wire w_dff_A_3EyJadJB5_0;
	wire w_dff_A_YYWsJkFt2_0;
	wire w_dff_A_CAtbH0kG3_1;
	wire w_dff_A_UDKg6Xpi4_1;
	wire w_dff_A_7boYskag2_1;
	wire w_dff_B_Uu9M7lfg3_1;
	wire w_dff_A_5T6fR9mq7_0;
	wire w_dff_A_V2kTa9Hc7_1;
	wire w_dff_A_CBiKKZIS9_1;
	wire w_dff_A_m63lOlLZ0_2;
	wire w_dff_A_RCuN0zd90_2;
	wire w_dff_A_ceAiW7Ji5_2;
	wire w_dff_A_iNfwLSLT6_2;
	wire w_dff_A_9Ucm2QPV0_0;
	wire w_dff_B_ylgvBcdh8_1;
	wire w_dff_B_StMgBiOW8_1;
	wire w_dff_A_Jv4JdZ5u5_0;
	wire w_dff_A_bObf0x0p0_2;
	wire w_dff_A_QUtchzXp5_2;
	wire w_dff_A_cKTpejlu2_2;
	wire w_dff_B_sAWPCcwN2_3;
	wire w_dff_A_LiPYbX3r1_0;
	wire w_dff_A_h8wzHYHy1_0;
	wire w_dff_A_Y8ywuaNP0_0;
	wire w_dff_A_n7tyjkY01_1;
	wire w_dff_A_t0O7mI4e6_1;
	wire w_dff_A_V3QMQZlU8_1;
	wire w_dff_A_Aw4CuAdT5_2;
	wire w_dff_A_fy8QgxEM9_2;
	wire w_dff_A_TqHrAkxw9_2;
	wire w_dff_A_6SJLGo5A5_2;
	wire w_dff_A_L2otT6Jw9_2;
	wire w_dff_B_PlhzTukc7_1;
	wire w_dff_B_z34FMFxU3_1;
	wire w_dff_B_urOdmBcw5_1;
	wire w_dff_A_zDVZzJHB6_0;
	wire w_dff_A_h0CDLY6r9_0;
	wire w_dff_A_VNw9zwzH9_0;
	wire w_dff_A_8WUE9jgd9_1;
	wire w_dff_A_xzteHJPG2_1;
	wire w_dff_A_Bt3PYd0s2_1;
	wire w_dff_A_lHGUgZ8b5_1;
	wire w_dff_A_soqt4kU63_1;
	wire w_dff_A_J674rONt9_1;
	wire w_dff_A_5IPRpY9Y5_2;
	wire w_dff_A_hO3uPZj88_2;
	wire w_dff_A_f02csFex8_2;
	wire w_dff_A_qKmwbaOo2_0;
	wire w_dff_B_kI5zuntE0_1;
	wire w_dff_B_nIieNhIp4_1;
	wire w_dff_B_sAsxMiBZ5_1;
	wire w_dff_B_LRLQwiRy6_1;
	wire w_dff_A_6W7MCHnj4_0;
	wire w_dff_A_Dsae1irt7_1;
	wire w_dff_A_d1Rk1TxE4_1;
	wire w_dff_A_JEmkZMiG7_1;
	wire w_dff_B_MdGS8fv19_3;
	wire w_dff_A_M6dwSquL8_0;
	wire w_dff_A_6mWxIoI89_0;
	wire w_dff_A_eW6SjnNt7_0;
	wire w_dff_A_hBJWfctI0_0;
	wire w_dff_A_oei47RLu4_1;
	wire w_dff_A_DcZGlTqU3_1;
	wire w_dff_A_Lb2WQcSu6_1;
	wire w_dff_A_yApM7iip3_1;
	wire w_dff_A_chyFBETF2_1;
	wire w_dff_A_Ien8KOZI6_1;
	wire w_dff_A_neKV7vsi6_2;
	wire w_dff_A_zOuC35UD9_2;
	wire w_dff_A_nAihT9iC1_2;
	wire w_dff_A_fMLuO8Bl6_2;
	wire w_dff_A_2Fs1iHVf5_2;
	wire w_dff_B_9PHn1ibD1_1;
	wire w_dff_B_4dGYIH7l0_1;
	wire w_dff_A_m2EfBMWh9_0;
	wire w_dff_A_lyM7So0B9_1;
	wire w_dff_A_1JaE5bQI8_1;
	wire w_dff_B_rPXNYChq5_3;
	wire w_dff_A_AkSqn7jB1_0;
	wire w_dff_A_7evdrxR06_0;
	wire w_dff_A_wHxj0fRF9_0;
	wire w_dff_A_Lc2dYLdb9_0;
	wire w_dff_A_R3XFGVbj1_1;
	wire w_dff_A_sbI6OpWy7_1;
	wire w_dff_A_21gc5b9b6_1;
	wire w_dff_A_ESqOpbAI9_1;
	wire w_dff_A_WiOLTzjr3_1;
	wire w_dff_A_GQKc1rbV2_1;
	wire w_dff_A_IgQAQ7Lt9_2;
	wire w_dff_A_KfzvHsFa9_2;
	wire w_dff_A_c3nhZ7hv3_2;
	wire w_dff_A_Mr0oGODM8_2;
	wire w_dff_A_I6WA4MZP3_2;
	wire w_dff_B_XtCAGJFa0_1;
	wire w_dff_A_ZS8Xkajg5_1;
	wire w_dff_A_iRVMvfNT1_1;
	wire w_dff_A_DxScrfm78_2;
	wire w_dff_B_Kg99jZtm0_3;
	wire w_dff_A_WG9HIbrZ6_0;
	wire w_dff_A_6smh6VMm0_0;
	wire w_dff_A_tiMkaR712_0;
	wire w_dff_A_PqVa93ns6_0;
	wire w_dff_A_TlxaThbe6_1;
	wire w_dff_A_Hh6tT1RF8_1;
	wire w_dff_A_sAN6ISD43_1;
	wire w_dff_B_qOYXn8xu5_1;
	wire w_dff_A_T83XRwcv4_0;
	wire w_dff_A_EgLqHu1D1_0;
	wire w_dff_A_fN7vApHP4_2;
	wire w_dff_A_JpespLa43_1;
	wire w_dff_A_8feY9c7F4_1;
	wire w_dff_A_8Lh2rrkD9_2;
	wire w_dff_A_1vRxJY3l1_2;
	wire w_dff_A_43WpCtLJ3_2;
	wire w_dff_A_TNgrttFd5_2;
	wire w_dff_A_HdWVF1nR3_1;
	wire w_dff_A_GWO37M1N8_2;
	wire w_dff_B_6xNAJWZH8_1;
	wire w_dff_B_w3oQLA3K1_1;
	wire w_dff_A_4sti3Suj9_0;
	wire w_dff_A_eXonkdlb7_1;
	wire w_dff_A_7c7731Fg5_1;
	wire w_dff_A_pdvO5LkK8_2;
	wire w_dff_A_toLIV1WJ6_2;
	wire w_dff_B_AdYaPkP42_3;
	wire w_dff_A_VSZtUZ2U3_0;
	wire w_dff_A_8iuV7Q6Y6_0;
	wire w_dff_A_aRqKwDbl9_0;
	wire w_dff_A_n93wh5bo2_0;
	wire w_dff_A_Qh7Wzjfr2_1;
	wire w_dff_A_Ix1uHo1p1_1;
	wire w_dff_A_Gn4kNrmx8_1;
	wire w_dff_A_BO4uaQtK5_1;
	wire w_dff_A_zeXCtxqQ1_1;
	wire w_dff_A_Dw0DhlT63_1;
	wire w_dff_A_9wZqrTU88_2;
	wire w_dff_A_TK5xeshE4_2;
	wire w_dff_A_bvrIgDs56_2;
	wire w_dff_A_k06UHQ5A1_2;
	wire w_dff_A_iLESAI844_2;
	wire w_dff_A_ZPs6zkcb8_0;
	wire w_dff_A_l8cnWHa37_1;
	wire w_dff_A_USw4L3wP5_2;
	wire w_dff_B_Ql6raKPb3_1;
	wire w_dff_B_6uWvkJM58_1;
	wire w_dff_A_q5DKJWwU8_0;
	wire w_dff_A_kUArhjPR1_1;
	wire w_dff_A_1XgLJ2H39_2;
	wire w_dff_A_zHIQzKii4_1;
	wire w_dff_A_AAJrBaP18_1;
	wire w_dff_A_Q9KvcXOf2_2;
	wire w_dff_A_4IPrpr5s0_2;
	wire w_dff_B_7icCghZd5_3;
	wire w_dff_A_VCgnQjQ24_0;
	wire w_dff_A_1bSRuFLQ6_0;
	wire w_dff_A_TnqCR82Q3_0;
	wire w_dff_A_brC3Vu6C4_0;
	wire w_dff_A_8ZqrcTiy8_0;
	wire w_dff_A_ltWXsAXG3_0;
	wire w_dff_A_ug8P8f0F0_0;
	wire w_dff_A_BJ7UxRqH7_2;
	wire w_dff_A_UccuB1zX9_2;
	wire w_dff_A_ai55PT6o1_2;
	wire w_dff_A_2Rh94nuT9_1;
	wire w_dff_A_wwkj1LBC5_2;
	wire w_dff_A_clY56xZi9_2;
	wire w_dff_A_4BjCnYsa4_1;
	wire w_dff_A_njzoyN1m1_1;
	wire w_dff_A_TXctprQw6_1;
	wire w_dff_A_TZQPaEs70_1;
	wire w_dff_A_wzyPVgss4_1;
	wire w_dff_A_Q2uzrKly3_1;
	wire w_dff_A_jtu5VeW96_1;
	wire w_dff_A_c7aqkdPO9_1;
	wire w_dff_A_gjXtJhIe4_1;
	wire w_dff_A_uNcQqXEt9_1;
	wire w_dff_A_lzXJE4H84_1;
	wire w_dff_A_OYGfwP1Z3_1;
	wire w_dff_A_Vng23Yzf7_1;
	wire w_dff_A_KmbM6YnM1_1;
	wire w_dff_A_7jCuN2SO5_1;
	wire w_dff_A_B0JxwjqZ0_1;
	wire w_dff_A_BR90ggWF7_1;
	wire w_dff_A_TwZAxml05_2;
	wire w_dff_A_CAfVWKOV4_2;
	wire w_dff_A_IO2PFiQm1_2;
	wire w_dff_A_d7PL8Z2r4_2;
	wire w_dff_A_0HITXgMS0_2;
	wire w_dff_A_Roh18i988_2;
	wire w_dff_A_jfhLXF6C8_2;
	wire w_dff_A_l3hale7f1_2;
	wire w_dff_A_3vhr76GN0_1;
	wire w_dff_A_WtPchuSZ3_1;
	wire w_dff_A_AP2UQUWH2_1;
	wire w_dff_A_XjrQOuP52_1;
	wire w_dff_A_R3CgJ9rL2_2;
	wire w_dff_A_s3CCG6I42_2;
	wire w_dff_A_j0w5OR4N7_2;
	wire w_dff_A_Dq9oZTdE6_2;
	wire w_dff_A_z1Hfe0YB5_1;
	wire w_dff_A_wjIhlaw92_1;
	wire w_dff_A_HcshvQVC3_2;
	wire w_dff_A_g0hCcZSf8_2;
	wire w_dff_A_UxkExz4G1_2;
	wire w_dff_A_IOgCYga15_0;
	wire w_dff_A_86Kd2LNp4_0;
	wire w_dff_A_GN6xquat4_0;
	wire w_dff_A_14eD1Mxq5_0;
	wire w_dff_A_7ltQG4E96_0;
	wire w_dff_A_gLWajmgg3_0;
	wire w_dff_A_n6tz4ecN4_0;
	wire w_dff_A_sHtRfTck5_0;
	wire w_dff_A_wS8O3pQt5_0;
	wire w_dff_A_K1oLFTwL1_0;
	wire w_dff_A_lQ52r2gm2_0;
	wire w_dff_A_8eESOUSb4_0;
	wire w_dff_A_hln36Jja8_0;
	wire w_dff_A_yr91NgLu6_1;
	wire w_dff_A_mR1OWuD16_1;
	wire w_dff_A_4J4jjHV49_1;
	wire w_dff_A_PDU8dyMk8_1;
	wire w_dff_A_7GFOFje68_1;
	wire w_dff_A_OVOQANxh2_1;
	wire w_dff_A_0NTHthet9_1;
	wire w_dff_A_zonUQtxB9_1;
	wire w_dff_A_GLtjp44R2_1;
	wire w_dff_A_LTlLwcGZ3_1;
	wire w_dff_A_pVlcDcYX3_1;
	wire w_dff_A_0cskcqzx9_1;
	wire w_dff_A_0YbbMCGp7_1;
	wire w_dff_A_VZTMw77M2_1;
	wire w_dff_A_fGYA6cGq5_1;
	wire w_dff_A_rkY8ZJQK5_1;
	wire w_dff_A_WSYn5Wlw5_1;
	wire w_dff_A_JKDn27689_1;
	wire w_dff_A_yCTbubjL7_1;
	wire w_dff_A_TYG55EF44_1;
	wire w_dff_A_LyDSgra93_2;
	wire w_dff_A_ngEZdzKZ3_2;
	wire w_dff_A_JhkqXMBe3_2;
	wire w_dff_A_ERXfpw1o9_2;
	wire w_dff_A_GYFs6pbO1_2;
	wire w_dff_A_LCeujrmB4_2;
	wire w_dff_A_fcMhHoWx4_2;
	wire w_dff_A_4Hx3joJk7_2;
	wire w_dff_A_8YGmmi2j1_2;
	wire w_dff_A_iGCt53WG4_2;
	wire w_dff_A_C3JoLAx09_2;
	wire w_dff_A_3XBG0hhS1_2;
	wire w_dff_A_fwdwVIQH1_2;
	wire w_dff_A_zvli0YFL3_2;
	wire w_dff_A_ZT65vYE69_2;
	wire w_dff_A_HTHRu8sE3_2;
	wire w_dff_A_SlmKESRw3_2;
	wire w_dff_A_y64vHxzW0_2;
	wire w_dff_A_bIjzEVme5_2;
	wire w_dff_A_b2zXDVxs2_2;
	wire w_dff_A_4QIAdU0v9_2;
	wire w_dff_A_w1dqKSWk9_2;
	wire w_dff_A_CW0nffzh6_2;
	wire w_dff_A_NqbDsvmf2_2;
	wire w_dff_A_QjbnviA39_2;
	wire w_dff_A_LP9E1LB19_2;
	wire w_dff_A_5YG3Ifyi2_2;
	wire w_dff_A_MOuVyOFp9_2;
	wire w_dff_A_TPiTsZpu7_1;
	wire w_dff_A_hwZAhzoJ4_0;
	wire w_dff_A_8hWr8K4g5_0;
	wire w_dff_A_IW0G3zbl3_0;
	wire w_dff_A_SFV9tUrV6_0;
	wire w_dff_A_V2XmpVEJ7_0;
	wire w_dff_A_tYF0k17L9_0;
	wire w_dff_A_4Kl91n3z9_0;
	wire w_dff_A_D4IbTBJh3_0;
	wire w_dff_A_idSQuNNg4_0;
	wire w_dff_A_u0Q7WlNR5_0;
	wire w_dff_A_wh87OkOv4_0;
	wire w_dff_A_6IdwTX7I1_0;
	wire w_dff_A_0eu9l9GI7_0;
	wire w_dff_A_Fr2NndvB0_0;
	wire w_dff_A_9DaxWcVe5_0;
	wire w_dff_A_sEoFq9KD7_2;
	wire w_dff_A_fdHghczS2_2;
	wire w_dff_A_qQcbAbSF7_2;
	wire w_dff_A_YoyrKpu44_2;
	wire w_dff_A_BKE3x8si3_2;
	wire w_dff_A_I1FDdZFv7_2;
	wire w_dff_A_Ck1vgoxk8_2;
	wire w_dff_A_DBsxoXEE2_2;
	wire w_dff_A_vtwLbDZy9_2;
	wire w_dff_A_wdof90BC0_2;
	wire w_dff_A_4EUYFJ4L3_1;
	wire w_dff_A_ouFZAQwf3_1;
	wire w_dff_A_I6UTQ0tw0_1;
	wire w_dff_A_3o6uXX6Y4_1;
	wire w_dff_A_eQ2Nzjiz0_1;
	wire w_dff_A_wEBWTMQW0_1;
	wire w_dff_A_JOMmBiyi7_1;
	wire w_dff_A_ypNZPoWa5_1;
	wire w_dff_A_Q05xcyJb8_1;
	wire w_dff_A_GQQrUn1Z3_1;
	wire w_dff_A_DIcUxRg03_1;
	wire w_dff_A_sS5DdR5W9_1;
	wire w_dff_A_RcDW4DBp8_1;
	wire w_dff_A_Q5T4PhPy6_1;
	wire w_dff_A_wZLdBuM37_1;
	wire w_dff_A_DTuIgggF4_1;
	wire w_dff_A_4s07I5ZL8_1;
	wire w_dff_A_XXMmGeEz2_1;
	wire w_dff_A_LAjly4nG4_1;
	wire w_dff_A_asQoPrAi2_1;
	wire w_dff_A_nvVPJzbg4_1;
	wire w_dff_A_L6992mk66_2;
	wire w_dff_A_s5BfF6w16_2;
	wire w_dff_A_n6dlcIh69_2;
	wire w_dff_A_BGSjREbP3_2;
	wire w_dff_A_t0rquWFF1_2;
	wire w_dff_A_y5xFEzsz2_2;
	wire w_dff_A_2ZlucQDn5_2;
	wire w_dff_A_KXEVUhWT2_2;
	wire w_dff_A_HlvbUxnE9_2;
	wire w_dff_A_SKyEw6Pd4_2;
	wire w_dff_A_ByH6PFG89_2;
	wire w_dff_A_Z28xNWPq5_2;
	wire w_dff_A_OZOfdAdC6_2;
	wire w_dff_A_Lxo8zdzp5_2;
	wire w_dff_A_MCd0vN6K2_2;
	wire w_dff_A_23t6YQOa0_2;
	wire w_dff_A_pmVLIJvz9_2;
	wire w_dff_A_PisEcUlx9_2;
	wire w_dff_A_bxTVlKjW6_2;
	wire w_dff_A_zLTOu8JK5_2;
	wire w_dff_A_mpLRE0Je6_1;
	wire w_dff_A_am7yIxmf3_1;
	wire w_dff_A_rzsCQKzX1_1;
	wire w_dff_A_egFPZ24v2_1;
	wire w_dff_A_vzNTSyJY8_1;
	wire w_dff_A_1pgYDBut5_1;
	wire w_dff_A_FBWrHvsX9_1;
	wire w_dff_A_8cEyKX9r7_1;
	wire w_dff_A_u2oM8zTL1_1;
	wire w_dff_A_kPBZg1MM1_1;
	wire w_dff_A_xr7TWG8s3_1;
	wire w_dff_A_MypX9fp29_1;
	wire w_dff_A_ePr8cnFI4_1;
	wire w_dff_A_WpdWctLV6_1;
	wire w_dff_A_ZQuJxd5R4_1;
	wire w_dff_A_yuy19z7y0_1;
	wire w_dff_A_bOMjcM938_1;
	wire w_dff_A_pkIOg8DR5_1;
	wire w_dff_A_VxFFKIej9_2;
	wire w_dff_A_HqDQvGCU4_2;
	wire w_dff_A_55ETpfEB6_2;
	wire w_dff_A_9nnvYlqY6_2;
	wire w_dff_A_BFUe0ssz2_2;
	wire w_dff_A_ez6mDYfh9_2;
	wire w_dff_A_XzE95zm61_2;
	wire w_dff_A_XhWeXWgj3_2;
	wire w_dff_A_uV4raij88_2;
	wire w_dff_A_8EB01zUN2_2;
	wire w_dff_A_d18Xh9zG0_2;
	wire w_dff_A_4E7c0JBK7_1;
	wire w_dff_A_WLJRdjkR5_1;
	wire w_dff_A_JQwaCszr1_1;
	wire w_dff_A_GbYZZhVE4_1;
	wire w_dff_A_OkmxD4018_1;
	wire w_dff_A_gdG4XFfr2_1;
	wire w_dff_A_WnK7dBLg2_1;
	wire w_dff_A_kORXSVfs4_1;
	wire w_dff_A_RC3RjUy58_1;
	wire w_dff_B_vYP787lz7_2;
	wire w_dff_B_dv0Sk1rx6_2;
	wire w_dff_A_JyTimGTZ8_1;
	wire w_dff_A_tgSDKJZS0_1;
	wire w_dff_A_2FMNP6gm3_1;
	wire w_dff_A_SlXD9Zaz1_1;
	wire w_dff_A_4YxIrAtO3_1;
	wire w_dff_A_DR8HT2Cz2_1;
	wire w_dff_A_UqXC2gA67_1;
	wire w_dff_A_7Aw2yds87_1;
	wire w_dff_A_BSpXy12l8_1;
	wire w_dff_A_bxIaF5Z25_1;
	wire w_dff_A_ol4IIpzV2_1;
	wire w_dff_A_K6JfdkhC0_1;
	wire w_dff_A_9A60RQXf2_1;
	wire w_dff_A_OMbpm80E8_1;
	wire w_dff_A_i55synqN9_1;
	wire w_dff_A_QmNlyXPh1_1;
	wire w_dff_A_PIsCQWs12_1;
	wire w_dff_A_9iITZDPc3_1;
	wire w_dff_A_aaRdwr1T9_1;
	wire w_dff_A_5zpX7mQT5_1;
	wire w_dff_A_MCoDUxPh8_1;
	wire w_dff_A_4JolZxLh1_1;
	wire w_dff_A_MVuEkKuY4_1;
	wire w_dff_A_VuDmMeGV7_2;
	wire w_dff_A_Jk7SZmKU1_0;
	wire w_dff_A_FKs06vOf6_0;
	wire w_dff_A_m97GAm8A1_0;
	wire w_dff_A_jc7UkP114_0;
	wire w_dff_A_caH9ZvRL1_0;
	wire w_dff_A_kElsjG2o5_0;
	wire w_dff_A_ryM8UOrg9_0;
	wire w_dff_A_DU3H0pKq2_0;
	wire w_dff_A_Zw2VpOzO0_0;
	wire w_dff_A_ZSJKYVm82_0;
	wire w_dff_A_hjgvEmeW6_0;
	wire w_dff_A_azay8LDz1_0;
	wire w_dff_A_AK73ZF6E9_0;
	wire w_dff_A_9EMamk5B2_0;
	wire w_dff_A_7P1JnGap3_1;
	wire w_dff_A_VA0e6dU49_1;
	wire w_dff_A_3gBVCCOo6_1;
	wire w_dff_A_En2PdWcd5_1;
	wire w_dff_A_cDENqyZV9_1;
	wire w_dff_A_QmRFrdBT0_1;
	wire w_dff_A_zukXn5n45_1;
	wire w_dff_A_THYbqjPJ2_1;
	wire w_dff_A_6kFmL9K90_1;
	wire w_dff_A_MDqysnyc5_1;
	wire w_dff_A_jJf4eWaU4_1;
	wire w_dff_A_eKR2wk7F9_1;
	wire w_dff_A_4PRyniVS0_1;
	wire w_dff_A_oc9mtfTm5_1;
	wire w_dff_A_SRXyEb8c0_1;
	wire w_dff_A_gA8plgWv0_1;
	wire w_dff_A_nAlCE6Zu1_2;
	wire w_dff_A_tONs35pE1_2;
	wire w_dff_A_H0ENVOgR9_2;
	wire w_dff_A_OYPEqwMm4_2;
	wire w_dff_A_8z4UllSI9_2;
	wire w_dff_A_ttefBYj68_2;
	wire w_dff_A_XtqX9Khd7_2;
	wire w_dff_A_Qy9KWbIF1_2;
	wire w_dff_A_nKzJime58_2;
	wire w_dff_A_s8CsorvS4_2;
	wire w_dff_A_0DJTXydb5_2;
	wire w_dff_A_HxUoWY1V0_2;
	wire w_dff_A_r4M3zkXA1_2;
	wire w_dff_A_TMOLMh414_2;
	wire w_dff_A_YaTrhLx00_2;
	wire w_dff_A_Cw34PnhY4_2;
	wire w_dff_A_jtW2qP6v7_2;
	wire w_dff_A_bQxer46m5_2;
	wire w_dff_A_3n4sw47y0_2;
	wire w_dff_A_2udhEhhk6_2;
	wire w_dff_A_ZGOI0Qfx5_2;
	wire w_dff_A_qR4PjBAd9_2;
	wire w_dff_A_PSVaiqWh9_1;
	wire w_dff_A_Q0BsbUps8_1;
	wire w_dff_A_bHyQFTVD8_1;
	wire w_dff_A_tSy389Iw5_1;
	wire w_dff_A_ZdkB8XYl8_1;
	wire w_dff_A_a2PHSSgC0_1;
	wire w_dff_A_4y1WoQs30_1;
	wire w_dff_A_u1wMxsoM7_1;
	wire w_dff_A_RnSWeJMG5_1;
	wire w_dff_A_ZFfkZLAp9_1;
	wire w_dff_A_CINpUQmP2_1;
	wire w_dff_A_wfKobEfZ0_1;
	wire w_dff_A_xOC9gKt38_1;
	wire w_dff_A_QzWa2Z5n5_1;
	wire w_dff_A_ZjwBPAsB1_1;
	wire w_dff_A_9Fnp6qaA7_1;
	wire w_dff_A_CGO9D06C0_1;
	wire w_dff_A_S1zFmDVS4_1;
	wire w_dff_A_1UZ6pyuM0_1;
	wire w_dff_A_OZQKo4iO6_2;
	wire w_dff_A_c1b1bM6v6_2;
	wire w_dff_A_N5q6kPc40_2;
	wire w_dff_A_UxubReMS9_2;
	wire w_dff_A_pgvIfkwn4_2;
	wire w_dff_A_8tNVIIbT6_2;
	wire w_dff_A_uuwaA6sV0_2;
	wire w_dff_A_ZQsuTpCw2_2;
	wire w_dff_A_A5cFD2H06_2;
	wire w_dff_A_HXPeOfLY2_2;
	wire w_dff_A_REPLKCAk0_2;
	wire w_dff_A_s6N5LyGp7_2;
	wire w_dff_A_vIIwWw7D2_2;
	wire w_dff_B_poQPHa3h8_2;
	wire w_dff_B_9f5pCFcU7_2;
	wire w_dff_B_YVCPnw5W1_2;
	wire w_dff_B_03d0JNAd2_2;
	wire w_dff_B_wxCaaXBG2_2;
	wire w_dff_B_cTF7mqUj3_2;
	wire w_dff_B_3Z9z2qyF9_2;
	wire w_dff_B_WO8yaWsY6_2;
	wire w_dff_B_G7S84XVG2_2;
	wire w_dff_B_F4ejeGlL8_2;
	wire w_dff_B_gAbkvH4z9_2;
	wire w_dff_B_lzassceA1_2;
	wire w_dff_B_prZSGH047_2;
	wire w_dff_B_YpQaawxc3_2;
	wire w_dff_B_touOMwKo6_2;
	wire w_dff_B_I22Xh09X7_2;
	wire w_dff_B_UnqBlSJv9_2;
	wire w_dff_B_UUV3vhOh6_2;
	wire w_dff_B_ocsGrU6Y3_2;
	wire w_dff_B_T64IbHBO2_2;
	wire w_dff_B_N35Ki1o12_2;
	wire w_dff_B_eI2nSmHx0_2;
	wire w_dff_B_oJDt5xgE5_2;
	wire w_dff_B_ieX59DMA8_2;
	wire w_dff_B_LB8SAABg1_2;
	wire w_dff_B_I3xFUquT7_2;
	wire w_dff_B_njf0WG6e3_2;
	wire w_dff_A_5643B7op6_2;
	wire w_dff_A_1Mm6hNVS3_2;
	wire w_dff_A_QFt1YS2g4_2;
	wire w_dff_A_qLNO8SMa7_2;
	wire w_dff_A_6wQ9wlX69_2;
	wire w_dff_A_rh9CCW4X3_2;
	wire w_dff_A_HY8txvO21_2;
	wire w_dff_A_azKJV0qw6_2;
	wire w_dff_A_OyQiFhFZ3_2;
	wire w_dff_A_J24N0Do60_2;
	wire w_dff_A_5KMFeiJ76_2;
	wire w_dff_A_WuSZRG9k6_2;
	wire w_dff_A_7FYlEURy4_2;
	wire w_dff_A_5pDfpnE62_2;
	wire w_dff_A_scV9Pi6d3_2;
	wire w_dff_A_4JKI4OUM2_2;
	wire w_dff_A_aG4fRHmC3_2;
	wire w_dff_A_Ddc85VlV1_2;
	wire w_dff_A_ZnZQwgwF9_2;
	wire w_dff_A_Md0HSSz69_2;
	wire w_dff_A_POH6v1gU4_2;
	wire w_dff_A_nMEdVV4X7_2;
	wire w_dff_A_6fVhreec5_2;
	wire w_dff_A_ggIDazgF3_2;
	wire w_dff_A_MDteAlzh1_0;
	wire w_dff_A_OjM5MU2Y3_0;
	wire w_dff_A_r64M6Z4L3_0;
	wire w_dff_A_b6XHtIlt2_0;
	wire w_dff_A_vWktkhc98_0;
	wire w_dff_A_jzLh2cW58_0;
	wire w_dff_A_crX2azFC6_0;
	wire w_dff_A_yOE54uKE6_0;
	wire w_dff_A_Rv8TeEZj6_0;
	wire w_dff_A_sw2wXDE82_0;
	wire w_dff_A_9V0ji26O5_0;
	wire w_dff_A_lMp6oV2H2_0;
	wire w_dff_A_mI4bnq797_0;
	wire w_dff_A_8PRL8ZI45_0;
	wire w_dff_A_JlWSIpyw7_0;
	wire w_dff_A_5bAthwJX1_0;
	wire w_dff_A_x4dZmg6f6_0;
	wire w_dff_A_nQdMsAbm8_1;
	wire w_dff_A_XX5yG7cJ0_1;
	wire w_dff_A_zuaPrjdN7_1;
	wire w_dff_A_QHhwW1gN1_1;
	wire w_dff_A_SJG7vEhs8_1;
	wire w_dff_A_gKQP4ugM2_1;
	wire w_dff_A_9JUSLCV17_1;
	wire w_dff_A_wkBd0UsZ7_1;
	wire w_dff_A_cibIhkzl2_1;
	wire w_dff_A_khUFWdNW0_1;
	wire w_dff_A_HLjqzoFC3_1;
	wire w_dff_A_j4YTQQb54_1;
	wire w_dff_A_c02mr9Nj5_1;
	wire w_dff_A_BpFCaTCQ1_1;
	wire w_dff_A_tQnXJQLk8_1;
	wire w_dff_A_KBaZDOHP1_1;
	wire w_dff_A_O55q3XcK7_0;
	wire w_dff_A_w1WlN4AI1_0;
	wire w_dff_A_d39dEwf79_0;
	wire w_dff_A_iRFpg1AX9_0;
	wire w_dff_A_gE5dWq0S1_0;
	wire w_dff_A_ZsBMiGr98_0;
	wire w_dff_A_nwvxDHjX7_0;
	wire w_dff_A_aO9mcUsK9_0;
	wire w_dff_A_n17gOZIr2_0;
	wire w_dff_A_YFNalbol9_0;
	wire w_dff_A_YG0sqLTW2_0;
	wire w_dff_A_YpF1Lz788_0;
	wire w_dff_A_JAwS5IiX2_0;
	wire w_dff_A_CXTW5kwL9_0;
	wire w_dff_A_BH73yURA2_0;
	wire w_dff_A_vk5O05BE9_0;
	wire w_dff_A_Sdq6fSR90_0;
	wire w_dff_A_uBjr6PJN0_0;
	wire w_dff_A_oSINyjGd2_0;
	wire w_dff_A_scs8vgnV1_0;
	wire w_dff_A_DVBqqvXa1_0;
	wire w_dff_A_ZhkqUzOK5_0;
	wire w_dff_A_fiDNaUrJ2_0;
	wire w_dff_A_wAivC2bE7_0;
	wire w_dff_A_9d6KjivI6_0;
	wire w_dff_A_qDCk6K6o9_0;
	wire w_dff_A_sQ8TdCZo1_0;
	wire w_dff_A_4s92yFbR3_1;
	wire w_dff_A_iaNi7GL72_0;
	wire w_dff_A_jeeHocm09_0;
	wire w_dff_A_iEpSj3AB0_0;
	wire w_dff_A_wQ5QBoUP2_0;
	wire w_dff_A_ACyjzPfS1_0;
	wire w_dff_A_Du8rORXL4_0;
	wire w_dff_A_HCIvCoYX1_0;
	wire w_dff_A_Fs8KLIcd3_0;
	wire w_dff_A_Evrcr3Cn2_0;
	wire w_dff_A_SYf1JhFY3_0;
	wire w_dff_A_4dNXf1YS2_0;
	wire w_dff_A_l9JSuQe12_0;
	wire w_dff_A_V4cbptXz5_0;
	wire w_dff_A_heYE8yQO8_0;
	wire w_dff_A_owQF4Orj7_0;
	wire w_dff_A_gmbncTAf6_0;
	wire w_dff_A_p0EEFjqn4_0;
	wire w_dff_A_c79ofdHL9_0;
	wire w_dff_A_BsmwsAGq7_0;
	wire w_dff_A_81mxqh3e1_0;
	wire w_dff_A_f28vrxeI8_0;
	wire w_dff_A_FMJuHK8E2_0;
	wire w_dff_A_aSCv58Ye4_0;
	wire w_dff_A_Vfi4Qppj4_0;
	wire w_dff_A_t1JBGe2o0_0;
	wire w_dff_A_QtudEZHd5_0;
	wire w_dff_A_1lI57vtL8_0;
	wire w_dff_A_nC4ucAtV8_1;
	wire w_dff_A_yj1mftS23_0;
	wire w_dff_A_C808ufh08_0;
	wire w_dff_A_Sk05vxiE6_0;
	wire w_dff_A_tT5h57D99_0;
	wire w_dff_A_Ut2HIQPJ1_0;
	wire w_dff_A_kBa65aPK7_0;
	wire w_dff_A_Lda4FzC81_0;
	wire w_dff_A_0KLFGTHZ8_0;
	wire w_dff_A_BD20nFcH8_0;
	wire w_dff_A_TixNXhdh6_0;
	wire w_dff_A_9C3qfpFN7_0;
	wire w_dff_A_QLk8oJKB1_0;
	wire w_dff_A_OBdxKKiw8_0;
	wire w_dff_A_xBXelP438_0;
	wire w_dff_A_glkSImVQ6_0;
	wire w_dff_A_qFRBqL0F8_0;
	wire w_dff_A_kDerP2dF3_0;
	wire w_dff_A_7vWTjxYE3_0;
	wire w_dff_A_NF90MJWc2_0;
	wire w_dff_A_wLf5JT0f0_0;
	wire w_dff_A_czaFwE1w0_0;
	wire w_dff_A_VAl9tb9u1_0;
	wire w_dff_A_45WW4B4c5_0;
	wire w_dff_A_fwYGUm3D2_0;
	wire w_dff_A_iiHRlj2M3_0;
	wire w_dff_A_w7a0VZHC3_0;
	wire w_dff_A_5mOEKxsL9_0;
	wire w_dff_A_ep1FTgkM5_1;
	wire w_dff_A_sG5fiiKG3_0;
	wire w_dff_A_8mLk11gH5_0;
	wire w_dff_A_gEGTZFFE5_0;
	wire w_dff_A_Ex4zNjTg9_0;
	wire w_dff_A_50WgwozR5_0;
	wire w_dff_A_v9fQoIi61_0;
	wire w_dff_A_jMuvNS7h7_0;
	wire w_dff_A_8RCay6Fk4_0;
	wire w_dff_A_pudPBWr98_0;
	wire w_dff_A_8jl9caJj3_0;
	wire w_dff_A_KDPIP7dV9_0;
	wire w_dff_A_8I1KSjuQ0_0;
	wire w_dff_A_tW4BgmE30_0;
	wire w_dff_A_CEMWlLdu1_0;
	wire w_dff_A_A1QkQi018_0;
	wire w_dff_A_FqUWZ8wB4_0;
	wire w_dff_A_wmIzeUMo4_0;
	wire w_dff_A_Ai5N5ciN2_0;
	wire w_dff_A_xqazbTIo7_0;
	wire w_dff_A_nswAEyaX7_0;
	wire w_dff_A_zlEdpTdk9_0;
	wire w_dff_A_M3qfnjbV0_0;
	wire w_dff_A_wzzMYBWz1_0;
	wire w_dff_A_Ig5Xr1RJ6_0;
	wire w_dff_A_JbWVN4om8_0;
	wire w_dff_A_shGbW1mx5_0;
	wire w_dff_A_vVTXHN0Y8_1;
	wire w_dff_A_T7qej8Wr6_0;
	wire w_dff_A_00lGSYGk9_0;
	wire w_dff_A_o3xTl1vp0_0;
	wire w_dff_A_61azdeHC7_0;
	wire w_dff_A_7lUkVmbZ0_0;
	wire w_dff_A_NqiOp5g87_0;
	wire w_dff_A_PFBfGFmI6_0;
	wire w_dff_A_tgKKQzvn0_0;
	wire w_dff_A_HsB2ReTN3_0;
	wire w_dff_A_amEKxW6y8_0;
	wire w_dff_A_cbTfVXzF2_0;
	wire w_dff_A_AFQXmTym4_0;
	wire w_dff_A_Y2LEw09O5_0;
	wire w_dff_A_qXAZ85gj6_0;
	wire w_dff_A_jHVNiXGu0_0;
	wire w_dff_A_Ah5OEZOB8_0;
	wire w_dff_A_Gr2rXtPe2_0;
	wire w_dff_A_2ZorcICg0_0;
	wire w_dff_A_Ec6mxR3J3_0;
	wire w_dff_A_NfA4Wpet6_0;
	wire w_dff_A_2WIERxJT2_0;
	wire w_dff_A_prNjylbA6_0;
	wire w_dff_A_gszMv0ZJ1_0;
	wire w_dff_A_c2GUCEwU2_0;
	wire w_dff_A_QPI9oVNu0_0;
	wire w_dff_A_ayQKAA0n6_0;
	wire w_dff_A_3AcVMzYK5_1;
	wire w_dff_A_0j5bfoEz0_0;
	wire w_dff_A_5msFLLaZ2_0;
	wire w_dff_A_HQ7EyUs90_0;
	wire w_dff_A_tVzeAobB4_0;
	wire w_dff_A_46BXZkeF5_0;
	wire w_dff_A_pKa5FU5T1_0;
	wire w_dff_A_ktA3ajId1_0;
	wire w_dff_A_sVJ62UAT1_0;
	wire w_dff_A_6dTh5qJ81_0;
	wire w_dff_A_tPGzkkzL1_0;
	wire w_dff_A_IA5TMtTJ8_0;
	wire w_dff_A_pOyCgSsE2_0;
	wire w_dff_A_4hUIvpAP3_0;
	wire w_dff_A_0O0QB71m9_0;
	wire w_dff_A_vn66pJ4c5_0;
	wire w_dff_A_xHGnSItg4_0;
	wire w_dff_A_IqmN4zcM3_0;
	wire w_dff_A_pUTUQbj52_0;
	wire w_dff_A_WeKdg6F09_0;
	wire w_dff_A_EI9YwJ1u6_0;
	wire w_dff_A_bo3gmzBx1_0;
	wire w_dff_A_u698IDfd9_0;
	wire w_dff_A_KZA8eMev8_0;
	wire w_dff_A_Q0hFrD3t4_0;
	wire w_dff_A_DBz8CL4e2_0;
	wire w_dff_A_ey8ymUK49_0;
	wire w_dff_A_vJT8vmhz2_1;
	wire w_dff_A_npcMJPQN3_0;
	wire w_dff_A_M1pwvoLi1_0;
	wire w_dff_A_kkReI27O4_0;
	wire w_dff_A_Nv32qHlP3_0;
	wire w_dff_A_Q3zV6DgZ0_0;
	wire w_dff_A_PS7bCVib4_0;
	wire w_dff_A_pHzQrpJB6_0;
	wire w_dff_A_BIzqZff30_0;
	wire w_dff_A_xTc5dEBV1_0;
	wire w_dff_A_fdQWXOgn6_0;
	wire w_dff_A_ZuCcz3uN6_0;
	wire w_dff_A_CacUs3Gb8_0;
	wire w_dff_A_uvgeC17M7_0;
	wire w_dff_A_XhEB0sUY4_0;
	wire w_dff_A_ZLfHUCVs8_0;
	wire w_dff_A_H4CR3XYo6_0;
	wire w_dff_A_1LnKWEV83_0;
	wire w_dff_A_PzdUgxQs7_0;
	wire w_dff_A_UsPgI78c7_0;
	wire w_dff_A_Dj1o5tiA7_0;
	wire w_dff_A_dWu8hV7i1_0;
	wire w_dff_A_A3g2c3Ur5_0;
	wire w_dff_A_hHr3EZtt5_0;
	wire w_dff_A_k9SaaSDn3_0;
	wire w_dff_A_qMPiwV2W2_0;
	wire w_dff_A_DW3x1vES3_0;
	wire w_dff_A_izx8mPSq2_1;
	wire w_dff_A_LX1UfqQN8_0;
	wire w_dff_A_nDs8iTmV8_0;
	wire w_dff_A_Xdeug0Jp0_0;
	wire w_dff_A_BtBvgrzV4_0;
	wire w_dff_A_QMA8XHCb9_0;
	wire w_dff_A_iWmqhsGu4_0;
	wire w_dff_A_GaADXKXM5_0;
	wire w_dff_A_aiYxBukP0_0;
	wire w_dff_A_cvbiK8eE6_0;
	wire w_dff_A_7QoaRM451_0;
	wire w_dff_A_WVOGs99W8_0;
	wire w_dff_A_Ar65qGqw4_0;
	wire w_dff_A_C6Wsa84o6_0;
	wire w_dff_A_7FZ4qnfn4_0;
	wire w_dff_A_WomVql2A1_0;
	wire w_dff_A_XWfPtfUX1_0;
	wire w_dff_A_wNg1G72Z6_0;
	wire w_dff_A_zBoW7lHC5_0;
	wire w_dff_A_El2akflr1_0;
	wire w_dff_A_PYo80HcF8_0;
	wire w_dff_A_pF6sYABj2_0;
	wire w_dff_A_LO29noL97_0;
	wire w_dff_A_6vS7HMc92_0;
	wire w_dff_A_ZncOYlGO8_0;
	wire w_dff_A_cYqjTFUI8_0;
	wire w_dff_A_SpSsRYeB7_0;
	wire w_dff_A_RRZ9uML84_1;
	wire w_dff_A_6EptrX162_0;
	wire w_dff_A_G1Od5GP96_0;
	wire w_dff_A_ww2wX3W68_0;
	wire w_dff_A_eUpFYx1Q4_0;
	wire w_dff_A_9jyRWsz84_0;
	wire w_dff_A_cEOuKijU0_0;
	wire w_dff_A_U1dLwSpL4_0;
	wire w_dff_A_qJrjx8857_0;
	wire w_dff_A_6YM9uwZO4_0;
	wire w_dff_A_bMHsJKsV9_0;
	wire w_dff_A_l7qQ59Ii4_0;
	wire w_dff_A_85XxBP1b8_0;
	wire w_dff_A_SMiNRLFk5_0;
	wire w_dff_A_0aw2phkN3_0;
	wire w_dff_A_4MAuS9uP6_0;
	wire w_dff_A_eqCk8I1c9_0;
	wire w_dff_A_zQJHRcpS0_0;
	wire w_dff_A_F4v23b1g8_0;
	wire w_dff_A_ONfuArJk5_0;
	wire w_dff_A_B31WohRv9_0;
	wire w_dff_A_56J56wQp5_0;
	wire w_dff_A_M4bXR5LO2_0;
	wire w_dff_A_cSeaWL8f3_0;
	wire w_dff_A_tXdSZS8I1_0;
	wire w_dff_A_ZTusLnzd9_0;
	wire w_dff_A_niCrNmJs9_0;
	wire w_dff_A_xFbNgCE53_1;
	wire w_dff_A_5893aecq4_0;
	wire w_dff_A_GIAAGkXz9_0;
	wire w_dff_A_UwzRAMYG4_0;
	wire w_dff_A_SDc5B45W1_0;
	wire w_dff_A_r0iswRXw1_0;
	wire w_dff_A_yVCieAOq5_0;
	wire w_dff_A_3WVmII6p7_0;
	wire w_dff_A_uUYAF0u26_0;
	wire w_dff_A_14UI74mt7_0;
	wire w_dff_A_99ogk7Wt1_0;
	wire w_dff_A_QlvLiMzP3_0;
	wire w_dff_A_6jDRWn8f6_0;
	wire w_dff_A_iDhn2Ez91_0;
	wire w_dff_A_2L4os6hZ9_0;
	wire w_dff_A_bJeOn2mx4_0;
	wire w_dff_A_5RDOpVQg8_0;
	wire w_dff_A_Nw4UiyEO0_0;
	wire w_dff_A_TiAHNh6O2_0;
	wire w_dff_A_1SWJcjHW5_0;
	wire w_dff_A_8GAHJglx9_0;
	wire w_dff_A_AETZv4DY2_0;
	wire w_dff_A_5dYYkKEV6_0;
	wire w_dff_A_12FzcyT90_0;
	wire w_dff_A_ub9PuNV94_0;
	wire w_dff_A_1VprEJfk0_0;
	wire w_dff_A_Rx9e6H5w5_0;
	wire w_dff_A_myx6F0wm9_1;
	wire w_dff_A_UPbPSexA2_0;
	wire w_dff_A_SKSuOZ973_0;
	wire w_dff_A_bC6iMBGw3_0;
	wire w_dff_A_QORnzm0y5_0;
	wire w_dff_A_OWgtybLQ2_0;
	wire w_dff_A_shekAVmn9_0;
	wire w_dff_A_BlVWxxaJ9_0;
	wire w_dff_A_ttLcXXNe3_0;
	wire w_dff_A_2zaXesmB2_0;
	wire w_dff_A_17yAvfwv3_0;
	wire w_dff_A_7zb7YPEd1_0;
	wire w_dff_A_JnvVGCU53_0;
	wire w_dff_A_MR65cec07_0;
	wire w_dff_A_GUMvMTUg2_0;
	wire w_dff_A_q1ryTd3G0_0;
	wire w_dff_A_r1NabILy2_0;
	wire w_dff_A_yNOMKLxZ6_0;
	wire w_dff_A_iZ4HgfDc1_0;
	wire w_dff_A_nV6Otl9y6_0;
	wire w_dff_A_Ow890cCz1_0;
	wire w_dff_A_S2SnoV9C1_0;
	wire w_dff_A_UFtKd3I17_0;
	wire w_dff_A_RtH6a8AC7_0;
	wire w_dff_A_xkoRBOk70_0;
	wire w_dff_A_Ip0SWz022_0;
	wire w_dff_A_F2VHMPQ78_0;
	wire w_dff_A_ICrsPWT71_1;
	wire w_dff_A_PwUBf2Dt3_0;
	wire w_dff_A_ejEYJ2y29_0;
	wire w_dff_A_zUDYgoom1_0;
	wire w_dff_A_mmYMCBTp6_0;
	wire w_dff_A_hKYDvdL87_0;
	wire w_dff_A_iJoOZddR5_0;
	wire w_dff_A_mMv9XXRP0_0;
	wire w_dff_A_1lJy1rlA8_0;
	wire w_dff_A_Ek8V9XCu6_0;
	wire w_dff_A_za8WoKtK7_0;
	wire w_dff_A_jgz879Xc9_0;
	wire w_dff_A_3YbwhwE11_0;
	wire w_dff_A_ags6rIIn5_0;
	wire w_dff_A_kFUpKGHf1_0;
	wire w_dff_A_pDtrcHpW6_0;
	wire w_dff_A_MnISrHh18_0;
	wire w_dff_A_QRIQjPyF8_0;
	wire w_dff_A_sWlWgiQ21_0;
	wire w_dff_A_Tbd5q3mP1_0;
	wire w_dff_A_Af1WBMLx1_0;
	wire w_dff_A_lqXiPWlu4_0;
	wire w_dff_A_pmC392pt7_0;
	wire w_dff_A_D3CK5Nub1_0;
	wire w_dff_A_HiEfJDVg9_0;
	wire w_dff_A_WzXcBO7K7_0;
	wire w_dff_A_Js0F6f5W7_0;
	wire w_dff_A_7QTZeYzo7_2;
	wire w_dff_A_GKPCB9Sa5_0;
	wire w_dff_A_hPEAL11N7_0;
	wire w_dff_A_l86Jl5LI4_0;
	wire w_dff_A_iJg4hL9o0_0;
	wire w_dff_A_3NxsMPhs9_0;
	wire w_dff_A_LTz9gH5m4_0;
	wire w_dff_A_iIf1YJl75_0;
	wire w_dff_A_2wgJWx869_0;
	wire w_dff_A_i1KxliVk9_0;
	wire w_dff_A_qbU5CQJt0_0;
	wire w_dff_A_qAV053ju7_0;
	wire w_dff_A_tN3hkU5U5_0;
	wire w_dff_A_0IpKMhuG4_0;
	wire w_dff_A_H8Soonyh7_0;
	wire w_dff_A_I9015LC60_0;
	wire w_dff_A_Pdyd3hMk8_0;
	wire w_dff_A_JSPV5HPF4_0;
	wire w_dff_A_kGL9ChU40_0;
	wire w_dff_A_UGxOMLY81_0;
	wire w_dff_A_ZN6s2Yu81_0;
	wire w_dff_A_uDXdqO9o8_0;
	wire w_dff_A_0I6ypgUF7_0;
	wire w_dff_A_7avwLBt46_0;
	wire w_dff_A_YrTK3Fc87_0;
	wire w_dff_A_1hjW2mnA6_0;
	wire w_dff_A_C6jLwmaC6_0;
	wire w_dff_A_aACQTVri0_1;
	wire w_dff_A_LwA9mG537_0;
	wire w_dff_A_jGHiufHt5_0;
	wire w_dff_A_dQu7MDDI8_0;
	wire w_dff_A_pxAoMv8v9_0;
	wire w_dff_A_fwb8saOd2_0;
	wire w_dff_A_K7AggtN31_0;
	wire w_dff_A_cbt7OtFF1_0;
	wire w_dff_A_LFJ0a3Ok5_0;
	wire w_dff_A_JgF2gRN58_0;
	wire w_dff_A_pmc21HvS8_0;
	wire w_dff_A_GdlUhXSt2_0;
	wire w_dff_A_ruJevEXR0_0;
	wire w_dff_A_McHwuMQ00_0;
	wire w_dff_A_Akw6YEm68_0;
	wire w_dff_A_3X7OKRyH5_0;
	wire w_dff_A_PO5r0l5i0_0;
	wire w_dff_A_sgOvqIYj5_0;
	wire w_dff_A_Sb7svTrN6_0;
	wire w_dff_A_MRVGfrX30_0;
	wire w_dff_A_SMApoT755_0;
	wire w_dff_A_yFe9BGHJ4_0;
	wire w_dff_A_1SmvKHDK6_0;
	wire w_dff_A_XYOhwMu25_0;
	wire w_dff_A_IjEbgNNA6_0;
	wire w_dff_A_9bt5RQ0b4_0;
	wire w_dff_A_j8wplm9r5_0;
	wire w_dff_A_GGl98Dw74_1;
	wire w_dff_A_7fjAglrO2_0;
	wire w_dff_A_XThLXVq02_0;
	wire w_dff_A_guqdJuRK9_0;
	wire w_dff_A_1SwR83JX8_0;
	wire w_dff_A_A19UkKn51_0;
	wire w_dff_A_YQL2e9g54_0;
	wire w_dff_A_GcbbKzAH6_0;
	wire w_dff_A_wgZzcywv2_0;
	wire w_dff_A_PldWPQ5A2_0;
	wire w_dff_A_Y92iBXCG4_0;
	wire w_dff_A_XMUZeDWV4_0;
	wire w_dff_A_u3W0J0Um6_0;
	wire w_dff_A_dlgQr5Jj5_0;
	wire w_dff_A_iZUt9QcP7_0;
	wire w_dff_A_ddDbZ63u6_0;
	wire w_dff_A_kBNOjV2F0_0;
	wire w_dff_A_hXM72C1y1_0;
	wire w_dff_A_runAglZL5_0;
	wire w_dff_A_PeYKnPUy0_0;
	wire w_dff_A_kLpdds3F5_0;
	wire w_dff_A_F2BeMjGk0_0;
	wire w_dff_A_fu3FUC8D8_0;
	wire w_dff_A_NKnQs0Ww5_0;
	wire w_dff_A_rJjBTX8p7_0;
	wire w_dff_A_I6nzBz4j0_0;
	wire w_dff_A_BPa1Y1LR5_0;
	wire w_dff_A_SSAqx4n50_1;
	wire w_dff_A_cr9RgTlP6_0;
	wire w_dff_A_FB44OejC9_0;
	wire w_dff_A_SnEljJZ02_0;
	wire w_dff_A_TMteaZIn9_0;
	wire w_dff_A_qevtscPe9_0;
	wire w_dff_A_8ZexlqBd3_0;
	wire w_dff_A_NWHFzZc57_0;
	wire w_dff_A_TIoK4kMv6_0;
	wire w_dff_A_Yi6o9clo9_0;
	wire w_dff_A_dbWxIeWy7_0;
	wire w_dff_A_w29kXXER8_0;
	wire w_dff_A_tfZsEWzc3_0;
	wire w_dff_A_C2vpX75T4_0;
	wire w_dff_A_GwFpnkWH7_0;
	wire w_dff_A_wUciIsyg1_0;
	wire w_dff_A_GFDUZido9_0;
	wire w_dff_A_iuXFaMRO5_0;
	wire w_dff_A_050FeFT91_0;
	wire w_dff_A_wqbvMCEV7_0;
	wire w_dff_A_aKzwPIWl6_0;
	wire w_dff_A_YoYnhh8B7_0;
	wire w_dff_A_Djp167xu6_0;
	wire w_dff_A_O62PEz0Z7_0;
	wire w_dff_A_jipahLvn4_0;
	wire w_dff_A_gNCqqYGt2_0;
	wire w_dff_A_H6SLc7GP5_0;
	wire w_dff_A_DYNjfypZ7_1;
	wire w_dff_A_SXllwUeB1_0;
	wire w_dff_A_k5Ibsu3p7_0;
	wire w_dff_A_biIsWMuc3_0;
	wire w_dff_A_Kr1aarx15_0;
	wire w_dff_A_DkJhcVR97_0;
	wire w_dff_A_jTgN8fta8_0;
	wire w_dff_A_iML8XhOG3_0;
	wire w_dff_A_8Aet4vXu4_0;
	wire w_dff_A_Js5oazjZ3_0;
	wire w_dff_A_BOCHaZHH5_0;
	wire w_dff_A_6wdpodPw6_0;
	wire w_dff_A_zDEwES4z6_0;
	wire w_dff_A_yEzLuGhL0_0;
	wire w_dff_A_Qq2DYUyR9_0;
	wire w_dff_A_T7ZlTZ0P5_0;
	wire w_dff_A_vgb0VQIe9_0;
	wire w_dff_A_LjnDNZyK1_0;
	wire w_dff_A_OQarA5w44_0;
	wire w_dff_A_GBG7CNlC0_0;
	wire w_dff_A_KTNGYh7P9_0;
	wire w_dff_A_aUv6D9Ez0_0;
	wire w_dff_A_4Uh8XPLD4_0;
	wire w_dff_A_8oc1e8s20_0;
	wire w_dff_A_WjdJYfX37_0;
	wire w_dff_A_bLIr58ez0_0;
	wire w_dff_A_wej7VxvF9_0;
	wire w_dff_A_z8qnRYpc3_2;
	wire w_dff_A_KSXl4TP58_0;
	wire w_dff_A_4kRIGyic3_0;
	wire w_dff_A_6Mk5wrQW2_0;
	wire w_dff_A_2ri2mYmV2_0;
	wire w_dff_A_PbMBeDGo4_0;
	wire w_dff_A_id4IJGMU3_0;
	wire w_dff_A_ZDbmA7uH5_0;
	wire w_dff_A_nPJVA8tO1_0;
	wire w_dff_A_7DhbAVRD6_0;
	wire w_dff_A_Hx3PPjQL0_0;
	wire w_dff_A_AhdqAkx50_0;
	wire w_dff_A_9fliU4jh0_0;
	wire w_dff_A_pgZXVOqW9_0;
	wire w_dff_A_pBgHZpUf1_0;
	wire w_dff_A_YenyigRT8_0;
	wire w_dff_A_EU6A3Fsr0_0;
	wire w_dff_A_BZr8u2Y53_0;
	wire w_dff_A_r6Jbh0ju9_0;
	wire w_dff_A_080Svrp25_0;
	wire w_dff_A_zelzBhZh2_0;
	wire w_dff_A_tePGh3O03_0;
	wire w_dff_A_WpEobw7u0_0;
	wire w_dff_A_Hc1wxwZ89_0;
	wire w_dff_A_SXGBn3E45_0;
	wire w_dff_A_Pb3eeLyY6_0;
	wire w_dff_A_jzOhX75Q6_0;
	wire w_dff_A_OH6Zh5AK0_2;
	wire w_dff_A_N2KEKsvI8_0;
	wire w_dff_A_MIMUbMn05_0;
	wire w_dff_A_kxJNJilI8_0;
	wire w_dff_A_quTJmNWY2_0;
	wire w_dff_A_5hsWFbi39_0;
	wire w_dff_A_IfMazg3J2_0;
	wire w_dff_A_4ElZgcsd8_0;
	wire w_dff_A_TEvPyqf50_0;
	wire w_dff_A_pTX8Lrj61_0;
	wire w_dff_A_0RrTwjxH4_0;
	wire w_dff_A_H0GP8xz22_0;
	wire w_dff_A_ePVgpfCd9_0;
	wire w_dff_A_eiHZuPqO9_0;
	wire w_dff_A_fnOeO3MS8_0;
	wire w_dff_A_L9fLYnFc6_0;
	wire w_dff_A_I2pDEBjq2_0;
	wire w_dff_A_yKFCD9rK7_0;
	wire w_dff_A_iUXtmZsD8_0;
	wire w_dff_A_z8lBlD5z9_0;
	wire w_dff_A_sfhm1jSA3_0;
	wire w_dff_A_tGGJOsZT3_0;
	wire w_dff_A_9DxYxE720_0;
	wire w_dff_A_T5KojIuZ8_0;
	wire w_dff_A_qK0KQUEf0_0;
	wire w_dff_A_C9JJiO8j7_0;
	wire w_dff_A_VhL8a7Hi2_2;
	wire w_dff_A_lmDI3Xpy0_0;
	wire w_dff_A_xmJYH3i71_0;
	wire w_dff_A_X4bah6s66_0;
	wire w_dff_A_GG8xJHLR0_0;
	wire w_dff_A_Am0rr8ia6_0;
	wire w_dff_A_ziniP1yg0_0;
	wire w_dff_A_0QqbKVWN2_0;
	wire w_dff_A_qNiaCk008_0;
	wire w_dff_A_B8eWEI7M4_0;
	wire w_dff_A_Tmn3B10n1_0;
	wire w_dff_A_AdqvXExo8_0;
	wire w_dff_A_IZIvzXdC9_0;
	wire w_dff_A_I6cozvEI7_0;
	wire w_dff_A_aVQFqvYm5_0;
	wire w_dff_A_42X3hUSL4_0;
	wire w_dff_A_mnsE0i5h7_0;
	wire w_dff_A_08ZjJ4CS0_0;
	wire w_dff_A_ddxzzvO39_0;
	wire w_dff_A_w7YCfT897_0;
	wire w_dff_A_JZ6UktA11_0;
	wire w_dff_A_2J2pDMNO7_0;
	wire w_dff_A_pQCXdcjM9_0;
	wire w_dff_A_os0MY85t2_0;
	wire w_dff_A_FxIb3VD82_0;
	wire w_dff_A_DBAqT5CM5_0;
	wire w_dff_A_bVnKpyJe2_1;
	wire w_dff_A_sNMes2xq3_0;
	wire w_dff_A_gcwI9eLp5_0;
	wire w_dff_A_DhLlgaSN6_0;
	wire w_dff_A_j0Lu4hRI0_0;
	wire w_dff_A_xbCIpbPw8_0;
	wire w_dff_A_VVOeO6qV9_0;
	wire w_dff_A_AMPNKxgC4_0;
	wire w_dff_A_5vUqcwrY2_0;
	wire w_dff_A_X2FJdbXX2_0;
	wire w_dff_A_J4CyiKpG1_0;
	wire w_dff_A_0GBY2gXW5_0;
	wire w_dff_A_LZiyji1t2_0;
	wire w_dff_A_WG8yMshn7_0;
	wire w_dff_A_kpnAInKq8_0;
	wire w_dff_A_fb6p92pT0_0;
	wire w_dff_A_9CbOgmPp7_0;
	wire w_dff_A_H7bL1R8s8_0;
	wire w_dff_A_FS1QuHnS5_0;
	wire w_dff_A_wYxCKXSC5_0;
	wire w_dff_A_ByRSjIIX1_0;
	wire w_dff_A_mdZ8LgLo8_0;
	wire w_dff_A_1o1MSxgE0_0;
	wire w_dff_A_xgltJCvw2_0;
	wire w_dff_A_rcFxavpJ4_0;
	wire w_dff_A_pbKwJ33I5_0;
	wire w_dff_A_89syVh4x7_1;
	wire w_dff_A_1uvbwhDw4_0;
	wire w_dff_A_38iV7vhd5_0;
	wire w_dff_A_NLaJEFPh8_0;
	wire w_dff_A_0pXMRSfR2_0;
	wire w_dff_A_s5o6lvEh9_0;
	wire w_dff_A_NATKnATn3_0;
	wire w_dff_A_MHlUP8Er2_0;
	wire w_dff_A_kS1BFII74_0;
	wire w_dff_A_J3185Slh8_0;
	wire w_dff_A_K0N75OsA6_0;
	wire w_dff_A_EYyHNL9i5_0;
	wire w_dff_A_i1k7lZIg6_0;
	wire w_dff_A_EPBu9JjM2_0;
	wire w_dff_A_bakxyuKq1_0;
	wire w_dff_A_xJfYTcoW5_0;
	wire w_dff_A_Ti61som40_0;
	wire w_dff_A_OrvTgNDg2_0;
	wire w_dff_A_W8zT1ZWT0_0;
	wire w_dff_A_r0tORCi30_0;
	wire w_dff_A_5ieYbjB38_0;
	wire w_dff_A_yjf03Y5Q5_0;
	wire w_dff_A_7AIEKMpy6_0;
	wire w_dff_A_kl2cAbLN1_0;
	wire w_dff_A_cIFvpTN56_0;
	wire w_dff_A_RB8vrvXz7_0;
	wire w_dff_A_TrrcuXLq7_0;
	wire w_dff_A_gx8JxHGs8_0;
	wire w_dff_A_Djl8qfsF2_1;
	wire w_dff_A_uHwNA8uP4_0;
	wire w_dff_A_DdyKhmnY6_0;
	wire w_dff_A_o8HuD9hM3_0;
	wire w_dff_A_FTFAQXl47_0;
	wire w_dff_A_cbB2SOQa6_0;
	wire w_dff_A_ptTRaTXg6_0;
	wire w_dff_A_f3TOpIVJ4_0;
	wire w_dff_A_NDvHUJmN6_0;
	wire w_dff_A_ydJy0zww6_0;
	wire w_dff_A_OrkTTjHp0_0;
	wire w_dff_A_pbXFo8wI0_0;
	wire w_dff_A_FAcIb2ZA9_0;
	wire w_dff_A_DuVQZ8Zp5_0;
	wire w_dff_A_qCYSapFb8_0;
	wire w_dff_A_Ce3eQfKm3_0;
	wire w_dff_A_5yqLeVTs9_0;
	wire w_dff_A_X4Dd6mIJ0_0;
	wire w_dff_A_Xsg4b4qM0_0;
	wire w_dff_A_y0Q2HcCC9_0;
	wire w_dff_A_vswiE9ur9_0;
	wire w_dff_A_mkWQvSHp5_0;
	wire w_dff_A_1ysOx7qy7_0;
	wire w_dff_A_iYMq4zli7_0;
	wire w_dff_A_V9FvTsy90_0;
	wire w_dff_A_78Xgc0hA2_0;
	wire w_dff_A_bK7AZ3K36_0;
	wire w_dff_A_EDnwvmV64_0;
	wire w_dff_A_yjWZdSrI8_1;
	wire w_dff_A_ms8Ogwvj0_0;
	wire w_dff_A_83jEZO4Q4_0;
	wire w_dff_A_simhCqkU3_0;
	wire w_dff_A_z7IpTcvV0_0;
	wire w_dff_A_YLrRpXNn3_0;
	wire w_dff_A_9MUSjGPC7_0;
	wire w_dff_A_2V62cTiC1_0;
	wire w_dff_A_P2XWxGm99_0;
	wire w_dff_A_fCJR7X7t6_0;
	wire w_dff_A_OrE62XP96_0;
	wire w_dff_A_YbgL1t2N4_0;
	wire w_dff_A_IKaVbsgN3_0;
	wire w_dff_A_XaXi0i4v6_0;
	wire w_dff_A_dPhcw7DX7_0;
	wire w_dff_A_5SrttqCL2_0;
	wire w_dff_A_Dmy6ELkT9_0;
	wire w_dff_A_fO7YP6j59_0;
	wire w_dff_A_zbgsl6pe4_0;
	wire w_dff_A_KAM6vUaN3_0;
	wire w_dff_A_2DWTLcxA1_0;
	wire w_dff_A_Rg5ZErBR2_0;
	wire w_dff_A_CvJIUbm24_0;
	wire w_dff_A_ay0qS0rU1_0;
	wire w_dff_A_NS0MKecF1_0;
	wire w_dff_A_Y3YPvJS25_0;
	wire w_dff_A_6vBVRovC8_0;
	wire w_dff_A_IY6SMMSa5_0;
	wire w_dff_A_qN7P6uT37_1;
	wire w_dff_A_TGX3X0lo1_0;
	wire w_dff_A_aTTNi7kC6_0;
	wire w_dff_A_yoUPXft99_0;
	wire w_dff_A_k5TYflGb8_0;
	wire w_dff_A_GGgCHdBl1_0;
	wire w_dff_A_p9ZBD0Ij4_0;
	wire w_dff_A_qWaDCNBU8_0;
	wire w_dff_A_LAUJW3rj5_0;
	wire w_dff_A_spjQNx6D8_0;
	wire w_dff_A_newntnSS8_0;
	wire w_dff_A_R6nLkOSR2_0;
	wire w_dff_A_350XQWaM0_0;
	wire w_dff_A_LFiiiwHC7_0;
	wire w_dff_A_kqEd3cFC5_0;
	wire w_dff_A_VAHWTEKF6_0;
	wire w_dff_A_CCjeenWr3_0;
	wire w_dff_A_yPlqqW1x7_0;
	wire w_dff_A_vEnxif705_0;
	wire w_dff_A_jMyqDxfU2_0;
	wire w_dff_A_nq7ZcTK26_0;
	wire w_dff_A_oSAov2VM7_0;
	wire w_dff_A_FLyvadE44_0;
	wire w_dff_A_g1VTKuQY6_0;
	wire w_dff_A_7Xl50UlW7_0;
	wire w_dff_A_NPqMWFeW8_0;
	wire w_dff_A_xPevfiNR4_0;
	wire w_dff_A_QSkIBtqJ1_0;
	wire w_dff_A_PSsXJ15W0_1;
	wire w_dff_A_Ug2BgSzk9_0;
	wire w_dff_A_BBu9EIOM9_0;
	wire w_dff_A_ZMFkfpbE7_0;
	wire w_dff_A_qI1Ph0Ky6_0;
	wire w_dff_A_qDukArh07_0;
	wire w_dff_A_9U8MbDxN4_0;
	wire w_dff_A_895ieqmJ4_0;
	wire w_dff_A_uryfAE3j1_0;
	wire w_dff_A_NpFoXssA1_0;
	wire w_dff_A_HJGLyjP44_0;
	wire w_dff_A_OzFBeN273_0;
	wire w_dff_A_MC5kieKL0_0;
	wire w_dff_A_Q58p9H0s4_0;
	wire w_dff_A_agzX51c82_0;
	wire w_dff_A_RLXXXLze6_0;
	wire w_dff_A_5EE25wH68_0;
	wire w_dff_A_ylk7N2wh6_0;
	wire w_dff_A_pTINlDbJ7_0;
	wire w_dff_A_tAIuwWch8_0;
	wire w_dff_A_Y2dLup4P3_0;
	wire w_dff_A_C8dXU2ed3_0;
	wire w_dff_A_aZdJrW847_0;
	wire w_dff_A_EHyLl6oL0_0;
	wire w_dff_A_wdukhdF37_0;
	wire w_dff_A_jR4NHXAp0_0;
	wire w_dff_A_6466RNsy0_0;
	wire w_dff_A_05582kQs1_0;
	wire w_dff_A_qEhQ7mZt4_1;
	wire w_dff_A_VYiq91BK4_0;
	wire w_dff_A_Id3VjDEr4_0;
	wire w_dff_A_r7VL3lMI1_0;
	wire w_dff_A_oQmAHtLq9_0;
	wire w_dff_A_6nHge9MI2_0;
	wire w_dff_A_4tdLart07_0;
	wire w_dff_A_bMz4h6uN1_0;
	wire w_dff_A_sb8KNqAg8_0;
	wire w_dff_A_cyFhwre65_0;
	wire w_dff_A_yVQM5J398_0;
	wire w_dff_A_COp3oKn32_0;
	wire w_dff_A_CXY1px9e1_0;
	wire w_dff_A_PegklGeu8_0;
	wire w_dff_A_kXDuMQTE0_0;
	wire w_dff_A_w6Oqor3X4_0;
	wire w_dff_A_ualuFDsY8_0;
	wire w_dff_A_ObytXB1X9_0;
	wire w_dff_A_ACsoLH0A7_0;
	wire w_dff_A_tAq5Jsva7_0;
	wire w_dff_A_bysvXtS30_0;
	wire w_dff_A_9JVwg8Y61_0;
	wire w_dff_A_M5BuBABE1_0;
	wire w_dff_A_tjDV1YYa0_0;
	wire w_dff_A_iolEBKst5_0;
	wire w_dff_A_pJdVrf4L0_0;
	wire w_dff_A_du2bENbP6_0;
	wire w_dff_A_oqcc29e21_2;
	wire w_dff_A_Yqimw46x8_0;
	wire w_dff_A_t5B54jkc1_0;
	wire w_dff_A_u9HB3Ruf2_0;
	wire w_dff_A_v32F4mKa2_0;
	wire w_dff_A_QVtkJ8h12_0;
	wire w_dff_A_mas9Mo8i8_0;
	wire w_dff_A_1QJItDNs2_0;
	wire w_dff_A_U6lWPRgU2_0;
	wire w_dff_A_5PelUQCX2_0;
	wire w_dff_A_0AEkfg3q1_0;
	wire w_dff_A_xTN3EjxV8_0;
	wire w_dff_A_ZOHblKiH6_0;
	wire w_dff_A_0kqwJ3S26_0;
	wire w_dff_A_Q3AYVYiL7_0;
	wire w_dff_A_XOSBnFRT1_0;
	wire w_dff_A_c9tAdXBx3_0;
	wire w_dff_A_WnqdlrYJ9_0;
	wire w_dff_A_fdPuh2TP5_0;
	wire w_dff_A_O0VEYkna8_0;
	wire w_dff_A_4Zq9FWId0_0;
	wire w_dff_A_juj8VRgE0_0;
	wire w_dff_A_MvIbOGo68_0;
	wire w_dff_A_WDNapyno5_0;
	wire w_dff_A_XJ2fTZCO6_0;
	wire w_dff_A_CwjD3V1R2_2;
	wire w_dff_A_DS5EGWgg1_0;
	wire w_dff_A_GFwzC6XV8_0;
	wire w_dff_A_aPHB6ZpI6_0;
	wire w_dff_A_rF5evuqK8_0;
	wire w_dff_A_NdI6BpDJ8_0;
	wire w_dff_A_MDggdN5e4_0;
	wire w_dff_A_TPIh1QrY3_0;
	wire w_dff_A_Gkcfn5RK4_0;
	wire w_dff_A_D9V4I86y1_0;
	wire w_dff_A_BJIcDcHs5_0;
	wire w_dff_A_ttLtsfud7_0;
	wire w_dff_A_0UDfAeTo2_0;
	wire w_dff_A_XbXavE0S9_0;
	wire w_dff_A_TSVMNdIC4_0;
	wire w_dff_A_CI6NKT2n6_0;
	wire w_dff_A_0kPwUYkb7_0;
	wire w_dff_A_Ww5aTARl9_0;
	wire w_dff_A_ye4Yh7GD0_0;
	wire w_dff_A_5w0oXtj81_0;
	wire w_dff_A_WHCClyld9_0;
	wire w_dff_A_7VwZvmNA6_0;
	wire w_dff_A_Ka95FIKu8_0;
	wire w_dff_A_5GR9xbYu7_0;
	wire w_dff_A_jqBiUilE3_0;
	wire w_dff_A_y50DGCjn9_0;
	wire w_dff_A_Jr8Poux14_1;
	wire w_dff_A_F8bSBTaH3_0;
	wire w_dff_A_o3dv0q6f5_0;
	wire w_dff_A_cx2ZOHkk1_0;
	wire w_dff_A_qZhtsyp25_0;
	wire w_dff_A_oAEqgSbh1_0;
	wire w_dff_A_dKSe6A4v2_0;
	wire w_dff_A_AfOoE4qC9_0;
	wire w_dff_A_S5GWcIcB5_0;
	wire w_dff_A_h9cYaEAZ0_0;
	wire w_dff_A_4Zxeq7Up4_0;
	wire w_dff_A_eH7dVURb0_0;
	wire w_dff_A_8HFsyjQs2_0;
	wire w_dff_A_RIZedcK41_0;
	wire w_dff_A_1anNgPut1_0;
	wire w_dff_A_tpO0IO2S8_0;
	wire w_dff_A_GHavWRYA0_0;
	wire w_dff_A_b16INpQS9_0;
	wire w_dff_A_pcgwPvLI0_0;
	wire w_dff_A_5UoSz9aN1_0;
	wire w_dff_A_1teGdIhy7_0;
	wire w_dff_A_8z1PV1PL9_0;
	wire w_dff_A_E7ikNyBW4_0;
	wire w_dff_A_Hd6RFwKU0_0;
	wire w_dff_A_GZxFGRy99_0;
	wire w_dff_A_XYlrOvK51_0;
	wire w_dff_A_7l2rTrJ02_0;
	wire w_dff_A_0pxxqC283_0;
	wire w_dff_A_5qB1Wwgm5_1;
	wire w_dff_A_QiFcPK1d2_0;
	wire w_dff_A_KcNW2Nji3_0;
	wire w_dff_A_mY0YDJSm5_0;
	wire w_dff_A_Pai1qV8N2_0;
	wire w_dff_A_YECSUc3l7_0;
	wire w_dff_A_NiFIqM7g0_0;
	wire w_dff_A_aTPMHJjz4_0;
	wire w_dff_A_vZP94e7T5_0;
	wire w_dff_A_c5hovwXG6_0;
	wire w_dff_A_LTrnyG2e6_0;
	wire w_dff_A_pJ4DMt4b8_0;
	wire w_dff_A_my9kqod26_0;
	wire w_dff_A_z4148bWO6_0;
	wire w_dff_A_oebE02oE6_0;
	wire w_dff_A_sidP7CfN8_0;
	wire w_dff_A_5QARFbBz1_0;
	wire w_dff_A_qM7MkbBq3_0;
	wire w_dff_A_9hJpMHN12_0;
	wire w_dff_A_PHmR1R8v3_0;
	wire w_dff_A_xE7gTKhy9_0;
	wire w_dff_A_MdGHM0hg4_0;
	wire w_dff_A_BW4Rz7Wx0_0;
	wire w_dff_A_iPTIjNHM8_0;
	wire w_dff_A_gaaf1wZa8_0;
	wire w_dff_A_77sej2RW2_0;
	wire w_dff_A_Wjmm5db44_0;
	wire w_dff_A_Dyi2xxG79_0;
	wire w_dff_A_6PibwFQP0_1;
	wire w_dff_A_NAr0nbiS0_0;
	wire w_dff_A_7vcpugSA5_0;
	wire w_dff_A_PMuoWas64_0;
	wire w_dff_A_9mjG3KIa4_0;
	wire w_dff_A_WGFi5evy5_0;
	wire w_dff_A_raik2fwo0_0;
	wire w_dff_A_G1ZFgysv0_0;
	wire w_dff_A_yk23dkXe0_0;
	wire w_dff_A_oxQ6hHQa2_0;
	wire w_dff_A_NM7hZlOk6_0;
	wire w_dff_A_RURjXBRE1_0;
	wire w_dff_A_NEPMgGSQ6_0;
	wire w_dff_A_D3rzod2Y8_0;
	wire w_dff_A_CHiL6nAq2_0;
	wire w_dff_A_fVNyg9GQ7_0;
	wire w_dff_A_HV1qglns7_0;
	wire w_dff_A_gQdVYz3g4_0;
	wire w_dff_A_GGZ1bkbJ2_0;
	wire w_dff_A_48b1dG4j4_0;
	wire w_dff_A_NX0Mbq458_0;
	wire w_dff_A_lBLOVfDg7_0;
	wire w_dff_A_LqqgSHtT6_0;
	wire w_dff_A_qjoztbQ95_0;
	wire w_dff_A_x7PphQwi2_0;
	wire w_dff_A_jpb0fABL6_0;
	wire w_dff_A_5gaDKYYD1_0;
	wire w_dff_A_KRlEvn7Q5_0;
	wire w_dff_A_qMdRBAAX3_1;
	wire w_dff_A_PbAy1E7j9_0;
	wire w_dff_A_VP7Yuk048_0;
	wire w_dff_A_9JWn5wmt9_0;
	wire w_dff_A_OytqGTUF2_0;
	wire w_dff_A_iYOkjqJI0_0;
	wire w_dff_A_ngq5qNrN9_0;
	wire w_dff_A_mdTBWsOS5_0;
	wire w_dff_A_hNF3nORq8_0;
	wire w_dff_A_c9pQJQ6f5_0;
	wire w_dff_A_CxOK3SWi6_0;
	wire w_dff_A_V1rAConY6_0;
	wire w_dff_A_Rb6VoArY3_0;
	wire w_dff_A_TyodUl2B5_0;
	wire w_dff_A_kwjCYwuU4_0;
	wire w_dff_A_Gxen4T7b6_0;
	wire w_dff_A_QkFChoAe0_0;
	wire w_dff_A_PrRUgtQT1_0;
	wire w_dff_A_jflovsba6_0;
	wire w_dff_A_TOa7h5G44_0;
	wire w_dff_A_oG70jydl1_0;
	wire w_dff_A_SECA2VR75_0;
	wire w_dff_A_bQp0DKEC5_0;
	wire w_dff_A_HPPl2pon6_0;
	wire w_dff_A_4c3i4UQN2_0;
	wire w_dff_A_KWNXN5WD7_0;
	wire w_dff_A_WeWgc0Ks3_0;
	wire w_dff_A_cBoqA3M19_0;
	wire w_dff_A_Zz1Li1Zx3_1;
	wire w_dff_A_cCR9KJWS9_0;
	wire w_dff_A_IqOjfl9g1_0;
	wire w_dff_A_pK0WH2ev0_0;
	wire w_dff_A_DUvRX0o68_0;
	wire w_dff_A_0ADnCMfh8_0;
	wire w_dff_A_3RaMxQkp4_0;
	wire w_dff_A_ArgoCyNb1_0;
	wire w_dff_A_HDwlHXnf4_0;
	wire w_dff_A_Z6I7FigU6_0;
	wire w_dff_A_pWvkJEzi8_0;
	wire w_dff_A_BdFtLRAU6_0;
	wire w_dff_A_eNYZQxEt5_0;
	wire w_dff_A_IZnJYaqC9_0;
	wire w_dff_A_ICqH0h6V2_0;
	wire w_dff_A_FwWfb5WH2_0;
	wire w_dff_A_8yEdFNwL8_0;
	wire w_dff_A_Z4A7ykqo3_0;
	wire w_dff_A_KEw0JQQO1_0;
	wire w_dff_A_vyWxBQaY6_0;
	wire w_dff_A_6FoVjSK19_0;
	wire w_dff_A_dSgNEWpI3_0;
	wire w_dff_A_66KyrKr42_0;
	wire w_dff_A_tz0oaOhV2_0;
	wire w_dff_A_UZ1tRybF8_0;
	wire w_dff_A_0bfURztX9_0;
	wire w_dff_A_WsJHWIyI8_0;
	wire w_dff_A_sVE4msgX6_0;
	wire w_dff_A_AujOhDyB6_1;
	wire w_dff_A_TaYAKsDG3_0;
	wire w_dff_A_CvY2WmNa8_0;
	wire w_dff_A_IWtdi0Qj8_0;
	wire w_dff_A_NELiMDpj0_0;
	wire w_dff_A_ZPHDB9T20_0;
	wire w_dff_A_4DPSxF180_0;
	wire w_dff_A_1gPRKQvg4_0;
	wire w_dff_A_w3qxbbPi0_0;
	wire w_dff_A_RDwaEHnY7_0;
	wire w_dff_A_6eApylkC4_0;
	wire w_dff_A_J2IOZki74_0;
	wire w_dff_A_V4V9GpGs7_0;
	wire w_dff_A_8OiKwdFj1_0;
	wire w_dff_A_LPupaLFz1_0;
	wire w_dff_A_TikIZPQr3_0;
	wire w_dff_A_HCWY5qnu1_0;
	wire w_dff_A_8ixV8VVE1_0;
	wire w_dff_A_jBRbCC2h8_0;
	wire w_dff_A_iB7WVXaT5_0;
	wire w_dff_A_f0K8BVYe9_0;
	wire w_dff_A_SKy5dBIu3_0;
	wire w_dff_A_wcQfNUWc9_0;
	wire w_dff_A_xv2Ejnxx7_0;
	wire w_dff_A_qbXzBuoM0_0;
	wire w_dff_A_HiDj1bum9_0;
	wire w_dff_A_IQzfYfcm2_0;
	wire w_dff_A_pWrd5YD36_2;
	wire w_dff_A_jOtAdkIz7_0;
	wire w_dff_A_PfJ98FuH0_0;
	wire w_dff_A_mgKKCepW8_0;
	wire w_dff_A_Jzpmppu41_0;
	wire w_dff_A_ph7FrcEQ1_0;
	wire w_dff_A_k9shR9gN6_0;
	wire w_dff_A_PBJVTjTi4_0;
	wire w_dff_A_KKnSm9h82_0;
	wire w_dff_A_FtoURUJU1_0;
	wire w_dff_A_ZYYQSpt12_0;
	wire w_dff_A_CyfyQaoC9_0;
	wire w_dff_A_N3WZ1PBY1_0;
	wire w_dff_A_SW35YDbg5_0;
	wire w_dff_A_HI8RGUM81_0;
	wire w_dff_A_J9v79Wsf9_0;
	wire w_dff_A_HzN4Au3a0_0;
	wire w_dff_A_lnQSdueK3_0;
	wire w_dff_A_v5lUbtTR4_0;
	wire w_dff_A_siiUskm97_0;
	wire w_dff_A_ucsfF0rl3_0;
	wire w_dff_A_vpalG9se3_0;
	wire w_dff_A_kjjs7I8w5_0;
	wire w_dff_A_B9rike742_0;
	wire w_dff_A_N46YAxsg6_2;
	wire w_dff_A_8TcrshsE6_0;
	wire w_dff_A_3374SqzC3_0;
	wire w_dff_A_rfb9R1XU1_0;
	wire w_dff_A_25gbLvOf5_0;
	wire w_dff_A_7w2yytWT2_0;
	wire w_dff_A_JJuSxVmI3_0;
	wire w_dff_A_mMtFRIlC6_0;
	wire w_dff_A_81ut6cuy9_0;
	wire w_dff_A_TcAigBwB3_0;
	wire w_dff_A_cxziEPDK9_0;
	wire w_dff_A_P3xiG4970_0;
	wire w_dff_A_Ok59sxxA5_0;
	wire w_dff_A_qkfIa3ib4_0;
	wire w_dff_A_vQnTcW883_0;
	wire w_dff_A_GNqKwT5m5_0;
	wire w_dff_A_MpB9vjwZ8_0;
	wire w_dff_A_Ib0P5ISv5_0;
	wire w_dff_A_J5G9ejAb0_0;
	wire w_dff_A_VV0ccLqg3_0;
	wire w_dff_A_fhZ0wCzH2_0;
	wire w_dff_A_rUEVe7jm1_0;
	wire w_dff_A_n9aOoSr31_0;
	wire w_dff_A_OisW3IkR8_0;
	wire w_dff_A_2DKLk9un4_2;
	wire w_dff_A_JgRWRyUM9_0;
	wire w_dff_A_sRsUIoki6_0;
	wire w_dff_A_cLNbfYRR9_0;
	wire w_dff_A_CzXinyke2_0;
	wire w_dff_A_jlDt2KvY0_0;
	wire w_dff_A_lHKAmdl23_0;
	wire w_dff_A_meSPHwYE2_0;
	wire w_dff_A_5qWV42Zh4_0;
	wire w_dff_A_qbs43c601_0;
	wire w_dff_A_M8ughsjL8_0;
	wire w_dff_A_1zvoTGZW5_0;
	wire w_dff_A_EEj56grY2_0;
	wire w_dff_A_JEWybB8X1_0;
	wire w_dff_A_ZifTnYWB5_0;
	wire w_dff_A_zYfBxUM84_0;
	wire w_dff_A_LieJn0700_0;
	wire w_dff_A_gmSlfClF6_0;
	wire w_dff_A_o8esnD4y7_0;
	wire w_dff_A_6MMOqSuP1_0;
	wire w_dff_A_IIoEG4Ic0_0;
	wire w_dff_A_j7QSh7pg8_0;
	wire w_dff_A_DZvvssdZ8_0;
	wire w_dff_A_605ik9r09_0;
	wire w_dff_A_u4ojv5bs3_2;
	wire w_dff_A_16KvtlDM5_0;
	wire w_dff_A_AE1V1d4u8_0;
	wire w_dff_A_5JZE5UhL5_0;
	wire w_dff_A_BFqDstg08_0;
	wire w_dff_A_Baqx0k3F7_0;
	wire w_dff_A_wvgErWK60_0;
	wire w_dff_A_SWFk9gmT3_0;
	wire w_dff_A_CQR9DwNd3_0;
	wire w_dff_A_D41rGFeQ3_0;
	wire w_dff_A_ntIYE8CX3_0;
	wire w_dff_A_HLx8Hkqy9_0;
	wire w_dff_A_wq140oL94_0;
	wire w_dff_A_kBVz0q0L4_0;
	wire w_dff_A_vPg3e92w8_0;
	wire w_dff_A_2pZdvSAW8_0;
	wire w_dff_A_BfJvqf762_0;
	wire w_dff_A_b5crP4Yu0_0;
	wire w_dff_A_MgVB2XwL9_0;
	wire w_dff_A_4iW5KogW8_0;
	wire w_dff_A_DJNjM5wY4_0;
	wire w_dff_A_r4NeWXKY5_0;
	wire w_dff_A_l70H96972_0;
	wire w_dff_A_i06YsaSI0_0;
	wire w_dff_A_epPjhTZb9_0;
	wire w_dff_A_bFJAJXPe1_2;
	wire w_dff_A_HRxkIp9o4_0;
	wire w_dff_A_brxhaajo8_0;
	wire w_dff_A_rqEgMzgx2_0;
	wire w_dff_A_xtmTGpx37_0;
	wire w_dff_A_j9YDmjJY6_0;
	wire w_dff_A_qFNuSUng6_0;
	wire w_dff_A_jDpHhVf28_0;
	wire w_dff_A_SXcJ6NHi3_0;
	wire w_dff_A_iv66C4Kf9_0;
	wire w_dff_A_mXKibCkS0_0;
	wire w_dff_A_0Z5jUYvR1_0;
	wire w_dff_A_lNvV7wTx0_0;
	wire w_dff_A_nuiuHEdQ2_0;
	wire w_dff_A_LSOREHcD1_0;
	wire w_dff_A_0zWs6Ish4_0;
	wire w_dff_A_AchSd57e2_0;
	wire w_dff_A_isLWvKQ74_0;
	wire w_dff_A_2YAx5rET6_0;
	wire w_dff_A_XD4Wiv597_0;
	wire w_dff_A_93AyXj409_0;
	wire w_dff_A_Y0BA1O5Y9_0;
	wire w_dff_A_BForkMmX6_0;
	wire w_dff_A_toTyowSq4_2;
	wire w_dff_A_huRvzYvG5_0;
	wire w_dff_A_mrisWpg32_0;
	wire w_dff_A_bneBZArb2_0;
	wire w_dff_A_bHtGCzG00_0;
	wire w_dff_A_smvkZ8QC9_0;
	wire w_dff_A_FIShRQMh4_0;
	wire w_dff_A_ZHW6TmRm9_0;
	wire w_dff_A_Qx4k9JMK7_0;
	wire w_dff_A_4LjNqzSN8_0;
	wire w_dff_A_87ywqVwj9_0;
	wire w_dff_A_IgpJrgJ06_0;
	wire w_dff_A_J0E4AVTD5_0;
	wire w_dff_A_5Ltba8tL6_0;
	wire w_dff_A_R86nVaq74_0;
	wire w_dff_A_eXhXKr1I6_0;
	wire w_dff_A_2t9xbKcH2_0;
	wire w_dff_A_tJcF31Fj1_0;
	wire w_dff_A_nl8SbuXr2_0;
	wire w_dff_A_waSge6q12_0;
	wire w_dff_A_OJPwxRea2_0;
	wire w_dff_A_yxwC9F1D4_0;
	wire w_dff_A_xDV7McIN4_0;
	wire w_dff_A_OVjaSAb91_2;
	wire w_dff_A_Y9m4OCJQ8_0;
	wire w_dff_A_d3en3JWA3_0;
	wire w_dff_A_8tjISI2k2_0;
	wire w_dff_A_Jk1Oclct9_0;
	wire w_dff_A_f8fnUCoo8_0;
	wire w_dff_A_S0CLXpMb0_0;
	wire w_dff_A_IGTgyIzK7_0;
	wire w_dff_A_aicJM0Jc2_0;
	wire w_dff_A_ognLfPum9_0;
	wire w_dff_A_lzdKMGrs7_0;
	wire w_dff_A_sx8U9IIE6_0;
	wire w_dff_A_JDAyKZwk6_0;
	wire w_dff_A_kjLfUmyf6_0;
	wire w_dff_A_w7y70Prj3_0;
	wire w_dff_A_Y7Tzjf2d9_0;
	wire w_dff_A_ObMxRUlg5_0;
	wire w_dff_A_iaQv0iVY3_0;
	wire w_dff_A_FR42bIRy8_0;
	wire w_dff_A_Z3XH0dUe1_0;
	wire w_dff_A_zjRU8IB00_0;
	wire w_dff_A_NzFuA0gO8_0;
	wire w_dff_A_1wTxoZSx7_0;
	wire w_dff_A_YdWlFp8S9_2;
	wire w_dff_A_KCdz1AxZ4_0;
	wire w_dff_A_9bUfZwSh9_0;
	wire w_dff_A_DbnKsDVZ5_0;
	wire w_dff_A_JLStcglA9_0;
	wire w_dff_A_IHmy4y6X4_0;
	wire w_dff_A_z405AW0f4_0;
	wire w_dff_A_5D34Nn9Z9_0;
	wire w_dff_A_7wpAMKDJ5_0;
	wire w_dff_A_7sdL923o5_0;
	wire w_dff_A_hZszDikc8_0;
	wire w_dff_A_XHtnOvIV4_0;
	wire w_dff_A_l2TqMT775_0;
	wire w_dff_A_WtjTUU7V3_0;
	wire w_dff_A_bGyd42oc7_0;
	wire w_dff_A_boebuFR06_0;
	wire w_dff_A_ilrHZdo72_0;
	wire w_dff_A_xps0psrB4_0;
	wire w_dff_A_ADz86t9A8_0;
	wire w_dff_A_JassX8VE4_0;
	wire w_dff_A_clyvudyc4_0;
	wire w_dff_A_PiTLjypD1_0;
	wire w_dff_A_PRaWv27G2_0;
	wire w_dff_A_Cd9m9dFW8_2;
	wire w_dff_A_x1CFo4sI0_0;
	wire w_dff_A_ZO2M8zcj7_0;
	wire w_dff_A_TApE9Qia4_0;
	wire w_dff_A_cvEC4Gjj9_0;
	wire w_dff_A_69kCW8C87_0;
	wire w_dff_A_GGNGD3Ei0_0;
	wire w_dff_A_itbBHohL7_0;
	wire w_dff_A_P0SKdzAc4_0;
	wire w_dff_A_0xQlZc8H7_0;
	wire w_dff_A_r6cAHvdX3_0;
	wire w_dff_A_W8Qf7Pa14_0;
	wire w_dff_A_bn5LFuq27_0;
	wire w_dff_A_Ni8FRK3D5_0;
	wire w_dff_A_4GroKpjZ2_0;
	wire w_dff_A_HZFcZRWK7_0;
	wire w_dff_A_3hiyNlRf6_0;
	wire w_dff_A_dvsqEEWl7_0;
	wire w_dff_A_jD9Sw1kX4_0;
	wire w_dff_A_r4sKjRsk2_0;
	wire w_dff_A_ZvM57l6Z2_2;
	wire w_dff_A_WdJboYY90_0;
	wire w_dff_A_6kOSiZz19_0;
	wire w_dff_A_RG1W8S5X7_0;
	wire w_dff_A_RMyvq1En7_0;
	wire w_dff_A_qCi5ix938_0;
	wire w_dff_A_eeraTqlt9_0;
	wire w_dff_A_IPY8snXA5_0;
	wire w_dff_A_NIAZ5XQd5_0;
	wire w_dff_A_QGNLrBLj6_0;
	wire w_dff_A_2LWrXZGn6_0;
	wire w_dff_A_5tWQYmJe0_0;
	wire w_dff_A_utghDYRT6_0;
	wire w_dff_A_2p0QNLZG3_0;
	wire w_dff_A_EDWWRofg9_0;
	wire w_dff_A_n3ScF3jt9_0;
	wire w_dff_A_PiVqCAeu7_0;
	wire w_dff_A_oKIJQUEf6_0;
	wire w_dff_A_S5A92AwA3_0;
	wire w_dff_A_NVY0g9Mn7_2;
	wire w_dff_A_te31V8tb8_0;
	wire w_dff_A_7PSFedEB8_0;
	wire w_dff_A_cSiEQ6Tz3_0;
	wire w_dff_A_9wrg9FnJ0_0;
	wire w_dff_A_MtM22qNV1_0;
	wire w_dff_A_xyOHZi835_0;
	wire w_dff_A_gynlntUb3_0;
	wire w_dff_A_xFQm1ZIx9_0;
	wire w_dff_A_acEaxo339_0;
	wire w_dff_A_phwkpT6u2_0;
	wire w_dff_A_3kII0ws02_0;
	wire w_dff_A_MNbb10fD7_0;
	wire w_dff_A_9iz9nXQX7_0;
	wire w_dff_A_ILKO7dgF6_0;
	wire w_dff_A_atIJreu34_0;
	wire w_dff_A_3WiXZ4bC9_0;
	wire w_dff_A_mk7Y1tBd1_2;
	wire w_dff_A_XWkYgDBl3_0;
	wire w_dff_A_MYYB1R0X3_0;
	wire w_dff_A_EEHsWfuj6_0;
	wire w_dff_A_VrCn3CYH3_0;
	wire w_dff_A_4WCah3Wi3_0;
	wire w_dff_A_6bc9hTeH8_0;
	wire w_dff_A_AUrJXpFU8_0;
	wire w_dff_A_1Nuf7zd55_0;
	wire w_dff_A_RRrW0xeS8_0;
	wire w_dff_A_4t3pMGx94_0;
	wire w_dff_A_A1kuQrvv4_0;
	wire w_dff_A_Sg7zNRAK4_0;
	wire w_dff_A_nyCrfboS4_0;
	wire w_dff_A_GrVukXrF5_0;
	wire w_dff_A_m6xzbOsq9_0;
	wire w_dff_A_ZUlGVPQ64_0;
	wire w_dff_A_Csz3Tef33_0;
	wire w_dff_A_Bq7pFif89_2;
	wire w_dff_A_NyBMqd4Z6_0;
	wire w_dff_A_qcNk22lr4_0;
	wire w_dff_A_I8yrylqY5_0;
	wire w_dff_A_WeN5lfva2_0;
	wire w_dff_A_eeV7OZKH9_0;
	wire w_dff_A_Q1SYxoPh1_0;
	wire w_dff_A_1MwazopU0_0;
	wire w_dff_A_gcK41StV0_0;
	wire w_dff_A_ohIOO6na6_0;
	wire w_dff_A_9E7vaMOn9_0;
	wire w_dff_A_gO7jvR3r9_0;
	wire w_dff_A_3rtWMCxk3_0;
	wire w_dff_A_iOEkgF5u4_0;
	wire w_dff_A_8k6WEvqe0_0;
	wire w_dff_A_0dsAzb7T7_0;
	wire w_dff_A_fxjTDloC7_0;
	wire w_dff_A_NoDo0o8j6_0;
	wire w_dff_A_evdjIyls0_2;
	wire w_dff_A_jzBkylD54_0;
	wire w_dff_A_dOvZoZQW8_0;
	wire w_dff_A_flU1OcbQ4_0;
	wire w_dff_A_IaCaBPG70_0;
	wire w_dff_A_MNscD1Yw7_0;
	wire w_dff_A_qCZCqPYK8_0;
	wire w_dff_A_RutWYGiw4_0;
	wire w_dff_A_LINAJobM1_0;
	wire w_dff_A_Enp72iWw3_0;
	wire w_dff_A_7Xzq3iC61_0;
	wire w_dff_A_t84mrXfC6_0;
	wire w_dff_A_WQLg3pm16_0;
	wire w_dff_A_llFN5Ogb6_0;
	wire w_dff_A_IFpwLAmU4_0;
	wire w_dff_A_xc9BbSpL5_0;
	wire w_dff_A_TOOwjg3q4_0;
	wire w_dff_A_jptqbv0j0_1;
	wire w_dff_A_FtqcvtRC6_0;
	wire w_dff_A_3LSHXnf81_0;
	wire w_dff_A_gp9y5sWh5_0;
	wire w_dff_A_pYAb7dtf3_0;
	wire w_dff_A_VCTACPVm4_0;
	wire w_dff_A_DqzWFCu97_0;
	wire w_dff_A_mbaUhdEn2_0;
	wire w_dff_A_8PlfjvkJ0_0;
	wire w_dff_A_AmAi9hWm9_0;
	wire w_dff_A_Dfn5Cc469_0;
	wire w_dff_A_7Wt5ohOY3_0;
	wire w_dff_A_gE6SrsAq3_0;
	wire w_dff_A_HAroxZOP3_0;
	wire w_dff_A_tZoFuRcZ1_0;
	wire w_dff_A_GEJ6F2ho5_0;
	wire w_dff_A_i5tlMJ861_0;
	wire w_dff_A_p4bE12gd5_0;
	wire w_dff_A_4uzXs4RZ7_0;
	wire w_dff_A_7mdSQPoi2_0;
	wire w_dff_A_51ifvy761_0;
	wire w_dff_A_c0AQma3q7_0;
	wire w_dff_A_Ict1Uw3T0_0;
	wire w_dff_A_Pd8CgEzt0_1;
	wire w_dff_A_v7Pd294j0_0;
	wire w_dff_A_2S2kANZ27_0;
	wire w_dff_A_hC0YtMyi8_0;
	wire w_dff_A_YYD5lvIl2_0;
	wire w_dff_A_XLHXkMNy9_0;
	wire w_dff_A_wC4oP5EB6_0;
	wire w_dff_A_cHdSX8lB0_0;
	wire w_dff_A_OPyH4G9c4_0;
	wire w_dff_A_Nnbs9u3D5_0;
	wire w_dff_A_UHG6XuRY9_0;
	wire w_dff_A_YlzH4YUg0_0;
	wire w_dff_A_Cd08q5VN0_0;
	wire w_dff_A_PUGdYKYd2_0;
	wire w_dff_A_C5C7xX8N9_0;
	wire w_dff_A_OJ08mxmH9_0;
	wire w_dff_A_U0S7q3rb6_0;
	wire w_dff_A_4EP3LCcU4_0;
	wire w_dff_A_nqM6Xfxs1_0;
	wire w_dff_A_y6gvat6o4_0;
	wire w_dff_A_rIVKxv6q7_0;
	wire w_dff_A_2VdlY8Fw0_0;
	wire w_dff_A_RldWZnr82_0;
	wire w_dff_A_q1kryMCV0_2;
	wire w_dff_A_aRU6WpdG5_0;
	wire w_dff_A_neWwQV9V9_0;
	wire w_dff_A_ZCBEazSx6_0;
	wire w_dff_A_gZXIM8G05_0;
	wire w_dff_A_LT7T9m3H3_0;
	wire w_dff_A_3nXPjOxT4_0;
	wire w_dff_A_TVwHny2S3_0;
	wire w_dff_A_8aftCEWg1_0;
	wire w_dff_A_JKR21ULp9_0;
	wire w_dff_A_qH4se6w52_0;
	wire w_dff_A_wEQxfWDP6_0;
	wire w_dff_A_mlub69cP0_0;
	wire w_dff_A_APahAb4G9_0;
	wire w_dff_A_LaQp9IAo6_2;
	wire w_dff_A_PgdewXPo4_0;
	wire w_dff_A_0JXjAOFx6_0;
	wire w_dff_A_z9jSVDB27_0;
	wire w_dff_A_66Et3iiE7_0;
	wire w_dff_A_CjumOJ5r8_0;
	wire w_dff_A_Si0UQOSo6_0;
	wire w_dff_A_oYrTmP3u3_0;
	wire w_dff_A_8QS1SAlJ2_0;
	wire w_dff_A_65bIpZYP5_0;
	wire w_dff_A_ZhJTY5Jk0_0;
	wire w_dff_A_N8mTUgdb1_0;
	wire w_dff_A_Zrs1DhXz5_0;
	wire w_dff_A_dQPZa2Kn0_0;
	wire w_dff_A_Z1WTcebV0_0;
	wire w_dff_A_QcszTcHB2_2;
	wire w_dff_A_pIDMkYQ89_0;
	wire w_dff_A_cOkzL3up4_0;
	wire w_dff_A_u9CK4Sxx0_0;
	wire w_dff_A_PsOa3JsT8_0;
	wire w_dff_A_TsbGEXhh5_0;
	wire w_dff_A_3dlKoi9A8_0;
	wire w_dff_A_MSz5598y0_0;
	wire w_dff_A_18B72YHQ9_0;
	wire w_dff_A_r3B5LYTP4_0;
	wire w_dff_A_mvRDQt976_0;
	wire w_dff_A_nFHU9ngs0_0;
	wire w_dff_A_Y8YY6d2j0_0;
	wire w_dff_A_eHysdSF98_0;
	wire w_dff_A_wQ8OfEWM6_2;
	wire w_dff_A_aELJTW9w2_0;
	wire w_dff_A_pE0RVzCB1_0;
	wire w_dff_A_biQdVpgB5_0;
	wire w_dff_A_ZkOG7nRf2_0;
	wire w_dff_A_FAMRmQsz3_0;
	wire w_dff_A_w7XM9guO7_0;
	wire w_dff_A_pHhItWgi0_0;
	wire w_dff_A_AU7jaCK34_0;
	wire w_dff_A_0WpNeB0Z9_0;
	wire w_dff_A_PC8ItbCz1_0;
	wire w_dff_A_btSCVhcQ1_0;
	wire w_dff_A_6S4bjSJH8_0;
	wire w_dff_A_v3qbmY2d3_0;
	wire w_dff_A_Z2ObU6dd2_0;
	wire w_dff_A_JwnIrGQk0_1;
	wire w_dff_A_C4xH7tVi7_0;
	wire w_dff_A_OcGXpt8Z9_0;
	wire w_dff_A_n91V6SEJ8_0;
	wire w_dff_A_tynL68rk3_0;
	wire w_dff_A_hGwbCVo08_0;
	wire w_dff_A_8nc4jCvo7_0;
	wire w_dff_A_IKyIqu9h2_0;
	wire w_dff_A_3Ky37lAy2_0;
	wire w_dff_A_vvi2pJoo8_0;
	wire w_dff_A_2zdUVoqD6_0;
	wire w_dff_A_1CsSKF3k1_0;
	wire w_dff_A_KmtHVL3c2_0;
	wire w_dff_A_GjFEdSDm0_0;
	wire w_dff_A_QAetyHhr6_0;
	wire w_dff_A_VwPCmeLr2_0;
	wire w_dff_A_0MA9bC231_0;
	wire w_dff_A_aswn5hTa0_0;
	wire w_dff_A_8e8HGB357_0;
	wire w_dff_A_dKqdSLq24_0;
	wire w_dff_A_VFIEsrzx7_1;
	wire w_dff_A_Kk1amslp4_0;
	wire w_dff_A_ctHwxDA26_0;
	wire w_dff_A_fL1uaJKE5_0;
	wire w_dff_A_sgJBLYAJ9_0;
	wire w_dff_A_DKCyW6pd8_0;
	wire w_dff_A_8vlTKZo39_0;
	wire w_dff_A_Vb3Fqu1d0_0;
	wire w_dff_A_4mvlN60C0_0;
	wire w_dff_A_9QQMqnPi6_0;
	wire w_dff_A_XN0SEcMI0_0;
	wire w_dff_A_L97a1K454_0;
	wire w_dff_A_azqoZSDg4_0;
	wire w_dff_A_VpMHyHyO1_0;
	wire w_dff_A_LMHIKbp41_0;
	wire w_dff_A_ZyftNr317_1;
	wire w_dff_A_3untLjXb5_0;
	wire w_dff_A_SqPFw5wX7_0;
	wire w_dff_A_0IjxmDpF6_0;
	wire w_dff_A_wlmcdczE0_0;
	wire w_dff_A_v0pAfD2J4_0;
	wire w_dff_A_tAOAqvb11_0;
	wire w_dff_A_cFNv92mf3_0;
	wire w_dff_A_h0Tjdrh89_0;
	wire w_dff_A_serLEDNa0_0;
	wire w_dff_A_1IB063gI7_0;
	wire w_dff_A_WGlETsiS5_0;
	wire w_dff_A_UPp9Vnop8_0;
	wire w_dff_A_MeRrixpo5_0;
	wire w_dff_A_7vHO491q0_0;
	wire w_dff_A_1TnEsA7g0_0;
	wire w_dff_A_1grLQ4el5_0;
	wire w_dff_A_6IdK8xAF1_0;
	wire w_dff_A_mtoJbP4h4_1;
	wire w_dff_A_nvCzGaTf6_0;
	wire w_dff_A_9EtarGos9_0;
	wire w_dff_A_VEDWxJV33_0;
	wire w_dff_A_vhvYq4SF9_0;
	wire w_dff_A_SkpyfsEZ7_0;
	wire w_dff_A_7ngbVZOH2_0;
	wire w_dff_A_gQkpQBel8_0;
	wire w_dff_A_nf7oNB5I5_0;
	wire w_dff_A_Kism8BVd5_0;
	wire w_dff_A_CgLAglrU8_2;
	wire w_dff_A_LXK5wWH77_0;
	wire w_dff_A_79ufvbh97_0;
	wire w_dff_A_RZAVZjJD8_0;
	wire w_dff_A_kqVTFC2E8_0;
	wire w_dff_A_8jBoo9gs0_0;
	wire w_dff_A_kwk7g0yc3_0;
	wire w_dff_A_0jQu3geu3_0;
	wire w_dff_A_JerQidNt3_0;
	wire w_dff_A_PV84EtTp6_0;
	wire w_dff_A_dedbp4CL7_0;
	wire w_dff_A_dXcX4MYR2_0;
	wire w_dff_A_IyEev7oO5_0;
	wire w_dff_A_Pk0pOnrI0_0;
	wire w_dff_A_0TreeCMY9_1;
	wire w_dff_A_jCdOdkov6_0;
	wire w_dff_A_mu3R57fZ9_0;
	wire w_dff_A_5kOFeQuL7_0;
	wire w_dff_A_g44jRxw19_0;
	wire w_dff_A_3WNorKJD9_0;
	wire w_dff_A_HDw7VX9D5_0;
	wire w_dff_A_mK8JQec03_0;
	wire w_dff_A_T5qYpt4V1_0;
	wire w_dff_A_fOoMB7R01_0;
	wire w_dff_A_i4N3sXmR0_0;
	wire w_dff_A_tqhg0jtD8_0;
	wire w_dff_A_bJ2UM7v22_0;
	wire w_dff_A_aRP8PpQw1_1;
	wire w_dff_A_xoxA61ev1_0;
	wire w_dff_A_l8BlxnMc0_0;
	wire w_dff_A_8Wb5QN4C9_0;
	wire w_dff_A_imF7gaFM1_0;
	wire w_dff_A_sc6v5Ou48_0;
	wire w_dff_A_t9rMzcAm4_0;
	wire w_dff_A_5b7lwdYk7_0;
	wire w_dff_A_5857ocSk5_0;
	wire w_dff_A_rNpGfDUn0_0;
	wire w_dff_A_yIjaXRsn3_0;
	wire w_dff_A_5i0K9DG29_0;
	wire w_dff_A_rNxl7Uz86_0;
	wire w_dff_A_O7iZCGfN9_0;
	wire w_dff_A_cWVz6Ubw9_1;
	wire w_dff_A_gwtc3gQh9_0;
	wire w_dff_A_1Yob8p3J1_0;
	wire w_dff_A_NDy6gCHK4_0;
	wire w_dff_A_yxZRWfcC9_0;
	wire w_dff_A_b2IEnacL4_0;
	wire w_dff_A_DItqIM3H4_0;
	wire w_dff_A_fVD7jDbe1_0;
	wire w_dff_A_AdOfJN4w4_0;
	wire w_dff_A_JfhjMLSu2_0;
	wire w_dff_A_KasOH0KW7_0;
	wire w_dff_A_CcgIE2kV6_0;
	wire w_dff_A_ROHbMZeR3_0;
	wire w_dff_A_q01qvI1b7_0;
	wire w_dff_A_oAAEG4Qb2_0;
	wire w_dff_A_eB7LN01l1_0;
	wire w_dff_A_WzDV50rL1_2;
	wire w_dff_A_1WQqNT460_0;
	wire w_dff_A_SgEYbjjc6_0;
	wire w_dff_A_FZ8QYBHj0_0;
	wire w_dff_A_xl0ZOeH14_0;
	wire w_dff_A_zasEgTdG2_0;
	wire w_dff_A_n72n2s850_0;
	wire w_dff_A_rHA126FP0_0;
	wire w_dff_A_tb6ca8a54_0;
	wire w_dff_A_vwET7jYv4_0;
	wire w_dff_A_xQ3aBGyg2_0;
	wire w_dff_A_NACuYeNd7_0;
	wire w_dff_A_MPnZkezm8_0;
	wire w_dff_A_PL5MABKR8_0;
	wire w_dff_A_Xcf1pYNP1_1;
	wire w_dff_A_Xfb3PSfA2_0;
	wire w_dff_A_v0HqC36K5_0;
	wire w_dff_A_LQ0IBVtq5_0;
	wire w_dff_A_StdEhPuv8_0;
	wire w_dff_A_xxsUecIf7_0;
	wire w_dff_A_ydwbPhue5_0;
	wire w_dff_A_AsFgkaCG4_0;
	wire w_dff_A_Vq00UK2h0_0;
	wire w_dff_A_ZG74mYlJ4_0;
	wire w_dff_A_UH5QMYWn8_0;
	wire w_dff_A_TmxGSpUR0_0;
	wire w_dff_A_kFOPrfOa3_0;
	wire w_dff_A_4fYXhbSz2_1;
	wire w_dff_A_4s2xqPvZ1_0;
	wire w_dff_A_alSrChwX5_0;
	wire w_dff_A_xKfg0DK49_0;
	wire w_dff_A_CiNnPCiG6_0;
	wire w_dff_A_w1ALeF1X6_0;
	wire w_dff_A_SDXx9UyQ6_0;
	wire w_dff_A_FQLZYEwQ5_0;
	wire w_dff_A_7xFGPKkV4_0;
	wire w_dff_A_H0OqcpjM6_0;
	wire w_dff_A_kDAT9Psb4_0;
	wire w_dff_A_WkFCRsQT1_0;
	wire w_dff_A_Rq35Tq8u4_0;
	wire w_dff_A_5VGOjIgQ6_0;
	wire w_dff_A_uA1xalqg8_0;
	wire w_dff_A_cecI00zW2_1;
	wire w_dff_A_a2OhQGic0_0;
	wire w_dff_A_iiVW7oig7_0;
	wire w_dff_A_AR3vXfHt2_0;
	wire w_dff_A_tIxfdXRJ4_0;
	wire w_dff_A_QJIVTP0M3_0;
	wire w_dff_A_sqkYLEe03_0;
	wire w_dff_A_VO3EppYI0_0;
	wire w_dff_A_t097MXi33_0;
	wire w_dff_A_8tUlZekN8_0;
	wire w_dff_A_oXRdMPiV4_0;
	wire w_dff_A_r8uGsviM5_0;
	wire w_dff_A_HSH9YHwR7_0;
	wire w_dff_A_yT8r4ESN7_0;
	wire w_dff_A_hoIEO0MO1_0;
	wire w_dff_A_5JvVsRDQ2_0;
	wire w_dff_A_j4wRy3eY7_1;
	wire w_dff_A_whizhFCe3_0;
	wire w_dff_A_32kIXURn1_0;
	wire w_dff_A_hBA4Sey01_0;
	wire w_dff_A_obbFt1O36_0;
	wire w_dff_A_VCaAMLQt7_0;
	wire w_dff_A_o6UflteS0_0;
	wire w_dff_A_X5EEzZRu3_0;
	wire w_dff_A_ThuzIoiq5_0;
	wire w_dff_A_hvssTaIL6_0;
	wire w_dff_A_LGr9TRnY2_0;
	wire w_dff_A_8zm7Iq9E2_0;
	wire w_dff_A_7yQz3Z012_0;
	wire w_dff_A_vngx1fyN1_0;
	wire w_dff_A_YADLfDM62_0;
	wire w_dff_A_tFxjjqFZ0_0;
	wire w_dff_A_4uw0WhNL4_0;
	wire w_dff_A_LDVmy6xf9_1;
	wire w_dff_A_DNhCCQWP5_0;
	wire w_dff_A_hHg4PhMJ7_0;
	wire w_dff_A_Yki2C0eC2_0;
	wire w_dff_A_DF6MiZSk7_0;
	wire w_dff_A_1DpJCtoK7_0;
	wire w_dff_A_UHiBLZ2m6_0;
	wire w_dff_A_ohLDOpWV4_0;
	wire w_dff_A_O7xkq8va3_0;
	wire w_dff_A_VjHFoiEg1_0;
	wire w_dff_A_Bu9c7gBV1_0;
	wire w_dff_A_I3ofLbNy3_0;
	wire w_dff_A_Df5wHkPL5_0;
	wire w_dff_A_s3xTOZCM8_0;
	wire w_dff_A_5lTxik1F7_0;
	wire w_dff_A_0oScPgZE3_0;
	wire w_dff_A_os7iufY74_0;
	wire w_dff_A_zgFimIi60_0;
	wire w_dff_A_5Omzibjx3_0;
	wire w_dff_A_NDhWr5cn3_0;
	wire w_dff_A_XFSPDDuF1_1;
	wire w_dff_A_Gyv3mvEr2_0;
	wire w_dff_A_WPysNjOK6_0;
	wire w_dff_A_LJ2FMCiX4_0;
	wire w_dff_A_qalRgpAi5_0;
	wire w_dff_A_lRdXNXv91_0;
	wire w_dff_A_BhnySF2a4_0;
	wire w_dff_A_2KhPCSam7_0;
	wire w_dff_A_VpwJHiuj2_0;
	wire w_dff_A_JwwS0Ze11_0;
	wire w_dff_A_rWcrur6b6_0;
	wire w_dff_A_MvCoxQho3_0;
	wire w_dff_A_0lz9rzBO6_0;
	wire w_dff_A_iariGLAp4_0;
	wire w_dff_A_sNCdhDWI2_0;
	wire w_dff_A_5OZwGQr93_0;
	wire w_dff_A_90VmhJ6N4_0;
	wire w_dff_A_rwzH8ctH0_0;
	wire w_dff_A_RYcuxKUY6_0;
	wire w_dff_A_LojQ4O6a8_2;
	wire w_dff_A_fhRTsr0g6_0;
	wire w_dff_A_Qav62Bm62_0;
	wire w_dff_A_choGXKAM6_0;
	wire w_dff_A_cM2HiBzD5_0;
	wire w_dff_A_lD4PhfTP5_0;
	wire w_dff_A_aGlRU6By9_0;
	wire w_dff_A_3qAT6j0y8_0;
	wire w_dff_A_ifO26XYC5_2;
	wire w_dff_A_Ga7U7ueu8_0;
	wire w_dff_A_iADms8vr3_0;
	wire w_dff_A_FI0QRrNN2_0;
	wire w_dff_A_kJ5MLS4y0_0;
	wire w_dff_A_gP10RLMl1_0;
	wire w_dff_A_05DtLBpD9_0;
	wire w_dff_A_FG5x9kcg6_2;
	wire w_dff_A_3KjLJqhc3_0;
	wire w_dff_A_pHWukCto8_0;
	wire w_dff_A_7wbJbWma3_0;
	wire w_dff_A_tVUV7PH33_0;
	wire w_dff_A_369qkXKi3_0;
	wire w_dff_A_aPrPoqpV4_0;
	wire w_dff_A_W9Vo4v9l8_0;
	wire w_dff_A_saKgwT7n1_0;
	wire w_dff_A_WwXd2Wx76_0;
	wire w_dff_A_HS5fnaWm6_0;
	wire w_dff_A_z5rDJbAn4_0;
	wire w_dff_A_JOmnUMds0_2;
	wire w_dff_A_ThLxdI1c2_0;
	wire w_dff_A_CNOC1cE41_0;
	wire w_dff_A_0FJgxq9G5_0;
	wire w_dff_A_xdblaibq2_0;
	wire w_dff_A_o9EvYuQR7_0;
	wire w_dff_A_3SdChd5U6_0;
	wire w_dff_A_ZP9E1GS63_0;
	wire w_dff_A_6k6qiJuN0_0;
	wire w_dff_A_S8u6oNdq2_0;
	wire w_dff_A_REeoh9Ix1_0;
	wire w_dff_A_yZz67w788_0;
	wire w_dff_A_jqIyVt3z5_2;
	wire w_dff_A_a6w4mOZa7_0;
	wire w_dff_A_SU9TATiq3_0;
	wire w_dff_A_os4xKN308_0;
	wire w_dff_A_7GXsRNkE0_0;
	wire w_dff_A_6xhTyW7e6_0;
	wire w_dff_A_lWPPiM2p9_0;
	wire w_dff_A_PKe6noIS6_0;
	wire w_dff_A_BPQdP7vV4_2;
	wire w_dff_A_pV3GcW802_0;
	wire w_dff_A_aQaJ0lxD2_0;
	wire w_dff_A_HOTC0lbI8_0;
	wire w_dff_A_wC1FHTSu7_0;
	wire w_dff_A_AGE81Mej8_0;
	wire w_dff_A_fmaFpMg28_0;
	wire w_dff_A_75YbuoFO9_0;
	wire w_dff_A_JZqJ9of82_0;
	wire w_dff_A_D2cceXBm3_2;
	wire w_dff_A_aVQSBQqr3_0;
	wire w_dff_A_ekpLxEU60_0;
	wire w_dff_A_oXiNrvFE7_0;
	wire w_dff_A_gztFXmxf0_0;
	wire w_dff_A_ISA4hZLw1_0;
	wire w_dff_A_cE3UymY29_0;
	wire w_dff_A_B0TYGzQ58_0;
	wire w_dff_A_ZpEqsrB63_0;
	wire w_dff_A_RmBYI8wY6_0;
	wire w_dff_A_Y6QgWCFW9_0;
	wire w_dff_A_AEoA2Y3E4_2;
	wire w_dff_A_GDke7ttV5_0;
	wire w_dff_A_O2XduvVY3_0;
	wire w_dff_A_GWzhwAwj9_0;
	wire w_dff_A_yVCUwG0X9_0;
	wire w_dff_A_lrXr0hMv8_0;
	wire w_dff_A_GVenb3qR0_0;
	wire w_dff_A_1OVXuacQ4_0;
	wire w_dff_A_iAcPN2iP0_0;
	wire w_dff_A_5nsuGzt59_0;
	wire w_dff_A_0GA9B52D4_2;
	wire w_dff_A_7OUcHV2K3_0;
	wire w_dff_A_SoXXNMqx1_0;
	wire w_dff_A_PWbcLNIh1_0;
	wire w_dff_A_zVF2CYju0_0;
	wire w_dff_A_hIXASEkO7_0;
	wire w_dff_A_nSZhUOqs9_0;
	wire w_dff_A_8ooaBXL27_0;
	wire w_dff_A_PIbZeKxV2_2;
	wire w_dff_A_UeU8kFsv7_0;
	wire w_dff_A_ANrpXbpp0_0;
	wire w_dff_A_nmSiswmL9_0;
	wire w_dff_A_cbSy4NbF0_0;
	wire w_dff_A_JbQS280h0_0;
	wire w_dff_A_GJdXwLX77_0;
	wire w_dff_A_0p93KERt6_0;
	wire w_dff_A_im0l4GSm8_0;
	wire w_dff_A_ARx0zPuV9_2;
	wire w_dff_A_3oykOsDX5_0;
	wire w_dff_A_4aWo7xLC6_0;
	wire w_dff_A_KLBQhzhK4_0;
	wire w_dff_A_pNQ4GnV84_0;
	wire w_dff_A_VI5K4YOW2_0;
	wire w_dff_A_Tr6O11BU3_0;
	wire w_dff_A_sCvOXCik8_0;
	wire w_dff_A_xWsBFvJe6_0;
	wire w_dff_A_eyJRHqdw6_0;
	wire w_dff_A_cf8GP5E74_0;
	wire w_dff_A_ViDIITJZ5_2;
	wire w_dff_A_7BmhX4q84_0;
	wire w_dff_A_VQQhsHgK0_0;
	wire w_dff_A_xXm3HKaJ6_0;
	wire w_dff_A_G9QnRSkN4_0;
	wire w_dff_A_nu3dZDVW2_0;
	wire w_dff_A_q10fcxTz1_0;
	wire w_dff_A_TPVfqmyn0_0;
	wire w_dff_A_W7Q6ycmE1_0;
	wire w_dff_A_1RimJmaU4_0;
	wire w_dff_A_WJMGnPZm5_2;
	wire w_dff_A_jNVhEOKB2_0;
	wire w_dff_A_9twF5CGM4_0;
	wire w_dff_A_GkN6wtgT7_0;
	wire w_dff_A_aSumYti10_0;
	wire w_dff_A_KcoZXFZX4_0;
	wire w_dff_A_SSNmn5mZ1_0;
	wire w_dff_A_3gh9jhrR8_2;
	wire w_dff_A_rygam42w0_0;
	wire w_dff_A_d0Tv3I3B3_0;
	wire w_dff_A_KsLV205o3_0;
	wire w_dff_A_Ks4nR7gK1_0;
	wire w_dff_A_3roPNQ8t0_0;
	wire w_dff_A_8lQwb43X2_0;
	wire w_dff_A_1VW3DmDd3_0;
	wire w_dff_A_swGinSef6_0;
	wire w_dff_A_1uBpjeJa9_0;
	wire w_dff_A_JYKdF5A27_2;
	wire w_dff_A_criGi8qa7_0;
	wire w_dff_A_qGQ1eYVr5_0;
	wire w_dff_A_UnQd9nmp9_0;
	wire w_dff_A_2da2ZqQE7_0;
	wire w_dff_A_2c9eMvlY4_0;
	wire w_dff_A_3oWSqGQX5_0;
	wire w_dff_A_a0QAE0996_0;
	wire w_dff_A_TipkdRtq8_0;
	wire w_dff_A_F4nNpyMV2_0;
	wire w_dff_A_N23fx6Y26_2;
	wire w_dff_A_MZIpwCEs1_0;
	wire w_dff_A_4i2XggU13_0;
	wire w_dff_A_DqHzC5t82_0;
	wire w_dff_A_yKAQ5gaz3_0;
	wire w_dff_A_xjGl09qk2_0;
	wire w_dff_A_nNcdRbdL0_0;
	wire w_dff_A_KQ3abjVD8_0;
	wire w_dff_A_DbzolyGj5_0;
	wire w_dff_A_1W05j3Ma7_2;
	wire w_dff_A_HczZGVG62_0;
	wire w_dff_A_ypFB5xwd2_0;
	wire w_dff_A_VJxtsCrL3_0;
	wire w_dff_A_eEbU4kSa5_0;
	wire w_dff_A_RnW1Otv69_0;
	wire w_dff_A_vTDZFZYD2_2;
	wire w_dff_A_dzXYR51q2_0;
	wire w_dff_A_ntbpoAp36_0;
	wire w_dff_A_niYem8mS4_0;
	wire w_dff_A_V0cwFGeF1_0;
	wire w_dff_A_y6GK1rNB0_0;
	wire w_dff_A_omhyUGMP0_0;
	wire w_dff_A_DnkTZt5R7_0;
	wire w_dff_A_xzw6bPNm8_0;
	wire w_dff_A_MJBaLzfO8_0;
	wire w_dff_A_AjepxUwp4_2;
	wire w_dff_A_XCQr6ENL5_0;
	wire w_dff_A_4iUBItTP6_0;
	wire w_dff_A_5fy59RcD7_0;
	wire w_dff_A_KEY2srag6_0;
	wire w_dff_A_mjtU9AHk4_0;
	wire w_dff_A_orjcsuiy3_0;
	wire w_dff_A_pdsxLkeO1_0;
	wire w_dff_A_Jy8wTgxs7_0;
	wire w_dff_A_ljOFfVkY1_0;
	wire w_dff_A_YYfSZWDj9_2;
	wire w_dff_A_lUhqxXJL7_0;
	wire w_dff_A_YMjM2Ud85_0;
	wire w_dff_A_0UB1Df464_0;
	wire w_dff_A_9jfZYRcd1_0;
	wire w_dff_A_PdQpDT420_0;
	wire w_dff_A_E0S89ySh4_0;
	wire w_dff_A_BHXCaqFf0_0;
	wire w_dff_A_noQDTBnq8_0;
	wire w_dff_A_NtujIeyr1_2;
	wire w_dff_A_3GEXZkbc4_0;
	wire w_dff_A_5uzGkFqz9_0;
	wire w_dff_A_XYPAskFG3_0;
	wire w_dff_A_fHltWVbY3_0;
	wire w_dff_A_JuACqhWv4_0;
	wire w_dff_A_aKGtkH7S1_0;
	wire w_dff_A_bLgQBZ9M2_2;
	wire w_dff_A_Ry7IyVw57_0;
	wire w_dff_A_zKt59K149_0;
	wire w_dff_A_NSdd7evn8_0;
	wire w_dff_A_yCH3Lclx7_0;
	wire w_dff_A_yW12xv8D7_0;
	wire w_dff_A_ZmWFKoF42_0;
	wire w_dff_A_6j1meksg1_0;
	wire w_dff_A_N7k9uy9l9_0;
	wire w_dff_A_HFyqO3fr6_0;
	wire w_dff_A_IwSzkPSy1_1;
	wire w_dff_A_xmLRzduV5_0;
	wire w_dff_A_M57NM7Aw3_0;
	wire w_dff_A_SPCSwg5j3_0;
	wire w_dff_A_vGuKqxff8_0;
	wire w_dff_A_11Clv3lA0_0;
	wire w_dff_A_7dPYPCaj9_0;
	wire w_dff_A_LBerTre86_1;
	wire w_dff_A_7glTpZaY8_0;
	wire w_dff_A_sOEkLcEg6_0;
	wire w_dff_A_Dklo9zPs0_0;
	wire w_dff_A_3YWx98ka9_0;
	wire w_dff_A_3jdzWI766_0;
	wire w_dff_A_fKuXXjJx4_0;
	wire w_dff_A_rmyDQuBi2_0;
	wire w_dff_A_2FsCfOkF2_1;
	wire w_dff_A_KlbY66Mt6_0;
	wire w_dff_A_ocCd8uyj8_0;
	wire w_dff_A_fls6G7XE8_0;
	wire w_dff_A_OkihA47d8_0;
	wire w_dff_A_1fDItDbd7_0;
	wire w_dff_A_i6pwenAP1_0;
	wire w_dff_A_rvkGvTDO1_1;
	wire w_dff_A_6Cpsv1q82_0;
	wire w_dff_A_MErzE5j98_0;
	wire w_dff_A_Wqgza2RQ9_0;
	wire w_dff_A_hWOZ5pYt5_0;
	wire w_dff_A_p9EJNKVZ2_0;
	wire w_dff_A_nhz6DzGj1_0;
	wire w_dff_A_hTYwL6zP1_0;
	wire w_dff_A_06RPFrg26_0;
	wire w_dff_A_e0hzDGeR8_0;
	wire w_dff_A_hdaSVyk01_0;
	wire w_dff_A_C1ao7ope7_0;
	wire w_dff_A_GCA5ODBX8_2;
	wire w_dff_A_E1qSkLM86_0;
	wire w_dff_A_1QYWHjkS6_0;
	wire w_dff_A_Il36ld8O1_0;
	wire w_dff_A_vW0gvt8x0_0;
	wire w_dff_A_rBtOGuzq8_0;
	wire w_dff_A_nswSbyau4_0;
	wire w_dff_A_4R1SgZ0V5_0;
	wire w_dff_A_Bk3R6bQQ2_0;
	wire w_dff_A_NVyKeG0k4_0;
	wire w_dff_A_4dm6cnJD6_0;
	wire w_dff_A_krqCzVYp3_0;
	wire w_dff_A_iGMB3ghD4_0;
	wire w_dff_A_RmCZmxKB9_0;
	wire w_dff_A_6q9Z6IT89_0;
	wire w_dff_A_OqgYmzyH3_0;
	wire w_dff_A_6H9zuHzz1_0;
	wire w_dff_A_17s6VL7c5_1;
	wire w_dff_A_xJX52c8s6_0;
	wire w_dff_A_c4goXiz96_0;
	wire w_dff_A_rgA4Rmsz0_0;
	wire w_dff_A_2HcFLX1g2_0;
	wire w_dff_A_ogovuXZC5_0;
	wire w_dff_A_6AWDkRJl7_1;
	wire w_dff_A_CMvyFcM13_0;
	wire w_dff_A_KzUiaDeT1_0;
	wire w_dff_A_DzyFzZU60_0;
	wire w_dff_A_fOCbuJSH7_0;
	wire w_dff_A_xbFWoSHn1_0;
	wire w_dff_A_WDtBrpU84_0;
	wire w_dff_A_rndAmwxd1_0;
	wire w_dff_A_3FCjCRUX7_0;
	wire w_dff_A_RDGMn0975_1;
	wire w_dff_A_BO6oQZSM1_0;
	wire w_dff_A_7mTk3Ov96_0;
	wire w_dff_A_79c8EDKn7_0;
	wire w_dff_A_WASfQaS48_0;
	wire w_dff_A_q32xcWwK2_0;
	wire w_dff_A_kfyGwrzl8_0;
	wire w_dff_A_XkPdcrtq8_1;
	wire w_dff_A_gzDeM6uj5_0;
	wire w_dff_A_20ru1FE20_0;
	wire w_dff_A_L0fqvtNV9_0;
	wire w_dff_A_D6KCyxOu2_0;
	wire w_dff_A_1nW2iSBe6_0;
	wire w_dff_A_gNwfsd558_0;
	wire w_dff_A_iQi5mYeG0_0;
	wire w_dff_A_EnVzPwhT1_0;
	wire w_dff_A_dunK0EDY6_0;
	wire w_dff_A_e2RZ5Gl43_2;
	wire w_dff_A_bG2uJ3eV1_0;
	wire w_dff_A_xVvOH0tH8_0;
	wire w_dff_A_lS0zHRg66_0;
	wire w_dff_A_FqM4NOCB0_2;
	wire w_dff_A_4DvjwDJx3_0;
	wire w_dff_A_DeZOut8m1_0;
	wire w_dff_A_lz8TOsR45_2;
	wire w_dff_A_T7GgUKXY0_0;
	wire w_dff_A_PmtGzS3m3_0;
	wire w_dff_A_sgYWj5mX7_0;
	wire w_dff_A_WIFa6DUd8_2;
	wire w_dff_A_IGZem14g4_0;
	wire w_dff_A_0hmhzQZq2_0;
	wire w_dff_A_lqFU7hcd2_0;
	wire w_dff_A_qzcfvnFP9_2;
	wire w_dff_A_EaHqP5YT5_0;
	wire w_dff_A_GL5Omq3X5_0;
	wire w_dff_A_OEgS7cZX5_0;
	wire w_dff_A_YP9pzYy54_0;
	wire w_dff_A_OWe3VifZ2_2;
	wire w_dff_A_aUeO30zP0_0;
	wire w_dff_A_XIo6DZ1C0_0;
	wire w_dff_A_FRUnh6fN7_0;
	wire w_dff_A_SnzgluzA6_2;
	wire w_dff_A_HV3vwFJI0_0;
	wire w_dff_A_2k0MkZu08_0;
	wire w_dff_A_tiNEzIGs1_0;
	wire w_dff_A_xWOXwuxG9_2;
	wire w_dff_A_RMXMFMqp9_0;
	wire w_dff_A_eHIQODzU2_0;
	wire w_dff_A_qKI4RqgR6_0;
	wire w_dff_A_W9aXYAXe0_0;
	wire w_dff_A_XEra2e6U0_2;
	wire w_dff_A_zqQ1hpHe8_0;
	wire w_dff_A_gZvxIxvA7_0;
	wire w_dff_A_1gmJbbnx5_0;
	wire w_dff_A_nhdDMIc41_2;
	wire w_dff_A_c9kVy9Yk9_0;
	wire w_dff_A_iEsytF7y2_0;
	wire w_dff_A_8corv2mp0_2;
	wire w_dff_A_IQ7GLwJM3_0;
	wire w_dff_A_T1bIQLwm5_0;
	wire w_dff_A_8CLLA1Vs8_2;
	wire w_dff_A_M2kpsJKY0_0;
	wire w_dff_A_DYPsKfAw4_2;
	wire w_dff_A_EIWhP4VZ5_0;
	wire w_dff_A_KEz0mcUa8_0;
	wire w_dff_A_TC8wh8Mq3_0;
	wire w_dff_A_atPMyXnW8_2;
	wire w_dff_A_1TS8HJWG3_0;
	wire w_dff_A_BoJpPChj2_0;
	wire w_dff_A_7Un7AyR00_2;
	wire w_dff_A_e2zYwXgF4_0;
	wire w_dff_A_A9ssMPdF2_0;
	wire w_dff_A_JgJF4PTq7_2;
	wire w_dff_A_uQqnHAwU1_0;
	wire w_dff_A_PlcUNtY39_0;
	wire w_dff_A_UlPKT5TM8_2;
	wire w_dff_A_PM5GHO3P3_0;
	wire w_dff_A_qwxGPqp95_0;
	wire w_dff_A_aueYEHx92_0;
	wire w_dff_A_vETPxkNk9_0;
	wire w_dff_A_JBFDhhb70_0;
	wire w_dff_A_7huooCbl2_2;
	wire w_dff_A_A6z6T7NX4_0;
	wire w_dff_A_kKt2Q9X98_0;
	wire w_dff_A_qQ9eMm2M7_0;
	wire w_dff_A_v3AVm0XO2_0;
	wire w_dff_A_yp9N7ak12_0;
	wire w_dff_A_8I5o8ymm2_2;
	wire w_dff_A_fkiBKvyy9_2;
	jnot g0000(.din(w_G545_0[2]),.dout(w_dff_A_ep1FTgkM5_1),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(w_G366_0[1]),.dout(w_dff_A_3AcVMzYK5_1),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(w_dff_A_izx8mPSq2_1),.clk(gclk));
	jnot g0005(.din(w_G338_0[1]),.dout(w_dff_A_myx6F0wm9_1),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(w_dff_A_7QTZeYzo7_2),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(w_dff_A_aACQTVri0_1),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(w_dff_A_GGl98Dw74_1),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(w_dff_A_SSAqx4n50_1),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(w_dff_A_DYNjfypZ7_1),.clk(gclk));
	jand g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(w_dff_A_z8qnRYpc3_2),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_5pseY3ze5_1),.dout(w_dff_A_OH6Zh5AK0_2),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jor g0016(.dina(w_dff_B_5d0LIbSn2_0),.dinb(w_n316_0[1]),.dout(w_dff_A_VhL8a7Hi2_2),.clk(gclk));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(w_dff_A_bVnKpyJe2_1),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jor g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_),.clk(gclk));
	jor g0022(.dina(w_G809_3[1]),.dinb(w_dff_B_gZLfCesE0_1),.dout(w_dff_A_oqcc29e21_2),.clk(gclk));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jor g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330),.clk(gclk));
	jor g0030(.dina(n330),.dinb(w_dff_B_XXGaiOMy4_1),.dout(w_dff_A_pWrd5YD36_2),.clk(gclk));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jor g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336),.clk(gclk));
	jor g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(w_dff_A_N46YAxsg6_2),.clk(gclk));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jor g0038(.dina(w_G809_2[1]),.dinb(w_dff_B_3l13xEUy4_1),.dout(w_dff_A_u4ojv5bs3_2),.clk(gclk));
	jand g0039(.dina(w_n326_1[2]),.dinb(w_dff_B_1gs4QHJx1_1),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jor g0041(.dina(w_dff_B_0UaRHFHX3_0),.dinb(w_G809_2[0]),.dout(n342),.clk(gclk));
	jor g0042(.dina(n342),.dinb(w_dff_B_uWMWTVN67_1),.dout(n343),.clk(gclk));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(w_dff_A_bFJAJXPe1_2),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(w_dff_B_U8XNJdiR0_1),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jor g0046(.dina(w_dff_B_fcKXeWTj0_0),.dinb(w_G809_1[2]),.dout(n347),.clk(gclk));
	jor g0047(.dina(n347),.dinb(w_dff_B_rtRIxOw27_1),.dout(n348),.clk(gclk));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(w_dff_A_toTyowSq4_2),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(w_dff_B_dxVJs3kJ3_1),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jor g0051(.dina(w_dff_B_mV6sOTPV5_0),.dinb(w_G809_1[1]),.dout(n352),.clk(gclk));
	jor g0052(.dina(n352),.dinb(w_dff_B_49CQMAWp8_1),.dout(n353),.clk(gclk));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(w_dff_A_OVjaSAb91_2),.clk(gclk));
	jand g0054(.dina(w_G2358_0[2]),.dinb(G80),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_n326_0[2]),.dinb(w_dff_B_TonoSrvx8_1),.dout(n356),.clk(gclk));
	jor g0056(.dina(n356),.dinb(w_G809_1[0]),.dout(n357),.clk(gclk));
	jor g0057(.dina(n357),.dinb(w_dff_B_24q7TdUc7_1),.dout(n358),.clk(gclk));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(w_dff_A_YdWlFp8S9_2),.clk(gclk));
	jand g0059(.dina(w_G3552_0[1]),.dinb(w_G514_2[1]),.dout(n360),.clk(gclk));
	jnot g0060(.din(w_G514_2[0]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G3546_5[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(n362),.dinb(w_n361_0[1]),.dout(n363),.clk(gclk));
	jor g0063(.dina(n363),.dinb(w_dff_B_xP1DKWMQ0_1),.dout(n364),.clk(gclk));
	jnot g0064(.din(n364),.dout(n365),.clk(gclk));
	jnot g0065(.din(w_G251_5[1]),.dout(n366),.clk(gclk));
	jnot g0066(.din(w_G361_1[1]),.dout(n367),.clk(gclk));
	jand g0067(.dina(n367),.dinb(w_n366_1[2]),.dout(n368),.clk(gclk));
	jnot g0068(.din(w_G248_5[2]),.dout(n369),.clk(gclk));
	jand g0069(.dina(w_G361_1[0]),.dinb(w_n369_1[2]),.dout(n370),.clk(gclk));
	jor g0070(.dina(n370),.dinb(n368),.dout(n371),.clk(gclk));
	jnot g0071(.din(w_n371_0[1]),.dout(n372),.clk(gclk));
	jand g0072(.dina(w_n372_0[1]),.dinb(w_n365_0[1]),.dout(n373),.clk(gclk));
	jnot g0073(.din(w_G351_2[2]),.dout(n374),.clk(gclk));
	jnot g0074(.din(G3550),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_n375_4[2]),.dinb(w_n374_1[1]),.dout(n376),.clk(gclk));
	jnot g0076(.din(w_G534_2[1]),.dout(n377),.clk(gclk));
	jnot g0077(.din(w_G3552_0[0]),.dout(n378),.clk(gclk));
	jand g0078(.dina(w_n378_4[2]),.dinb(w_G351_2[1]),.dout(n379),.clk(gclk));
	jor g0079(.dina(n379),.dinb(w_n377_1[1]),.dout(n380),.clk(gclk));
	jor g0080(.dina(n380),.dinb(w_dff_B_1zB6cnra8_1),.dout(n381),.clk(gclk));
	jand g0081(.dina(w_G3546_5[0]),.dinb(w_G351_2[0]),.dout(n382),.clk(gclk));
	jand g0082(.dina(w_G3548_4[2]),.dinb(w_n374_1[0]),.dout(n383),.clk(gclk));
	jor g0083(.dina(n383),.dinb(w_dff_B_ndtQ8J8A2_1),.dout(n384),.clk(gclk));
	jor g0084(.dina(n384),.dinb(w_G534_2[0]),.dout(n385),.clk(gclk));
	jand g0085(.dina(n385),.dinb(n381),.dout(n386),.clk(gclk));
	jnot g0086(.din(w_G341_2[2]),.dout(n387),.clk(gclk));
	jand g0087(.dina(w_n375_4[1]),.dinb(w_n387_1[1]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G523_1[2]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n378_4[1]),.dinb(w_G341_2[1]),.dout(n390),.clk(gclk));
	jor g0090(.dina(n390),.dinb(w_n389_1[1]),.dout(n391),.clk(gclk));
	jor g0091(.dina(n391),.dinb(w_dff_B_6bDH561l7_1),.dout(n392),.clk(gclk));
	jand g0092(.dina(w_G3546_4[2]),.dinb(w_G341_2[0]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3548_4[1]),.dinb(w_n387_1[0]),.dout(n394),.clk(gclk));
	jor g0094(.dina(n394),.dinb(w_dff_B_6pT1L4yy1_1),.dout(n395),.clk(gclk));
	jor g0095(.dina(n395),.dinb(w_G523_1[1]),.dout(n396),.clk(gclk));
	jand g0096(.dina(n396),.dinb(n392),.dout(n397),.clk(gclk));
	jand g0097(.dina(w_n397_0[1]),.dinb(w_n386_0[1]),.dout(n398),.clk(gclk));
	jand g0098(.dina(n398),.dinb(w_dff_B_JiQHGNmO2_1),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G316_1[1]),.dinb(w_G248_5[1]),.dout(n400),.clk(gclk));
	jnot g0100(.din(w_G490_1[1]),.dout(n401),.clk(gclk));
	jnot g0101(.din(w_G316_1[0]),.dout(n402),.clk(gclk));
	jand g0102(.dina(w_n402_0[2]),.dinb(w_G251_5[0]),.dout(n403),.clk(gclk));
	jor g0103(.dina(n403),.dinb(w_n401_0[1]),.dout(n404),.clk(gclk));
	jor g0104(.dina(n404),.dinb(w_dff_B_fbBXViZA9_1),.dout(n405),.clk(gclk));
	jnot g0105(.din(w_G254_1[1]),.dout(n406),.clk(gclk));
	jand g0106(.dina(w_n402_0[1]),.dinb(w_n406_5[1]),.dout(n407),.clk(gclk));
	jnot g0107(.din(w_G242_1[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_G316_0[2]),.dinb(w_n408_5[2]),.dout(n409),.clk(gclk));
	jor g0109(.dina(n409),.dinb(n407),.dout(n410),.clk(gclk));
	jor g0110(.dina(n410),.dinb(w_G490_1[0]),.dout(n411),.clk(gclk));
	jand g0111(.dina(n411),.dinb(n405),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G308_1[2]),.dinb(w_G248_5[0]),.dout(n413),.clk(gclk));
	jnot g0113(.din(w_G479_0[2]),.dout(n414),.clk(gclk));
	jnot g0114(.din(w_G308_1[1]),.dout(n415),.clk(gclk));
	jand g0115(.dina(w_n415_0[1]),.dinb(w_G251_4[2]),.dout(n416),.clk(gclk));
	jor g0116(.dina(n416),.dinb(w_n414_0[1]),.dout(n417),.clk(gclk));
	jor g0117(.dina(n417),.dinb(w_dff_B_h6IJkdMG1_1),.dout(n418),.clk(gclk));
	jand g0118(.dina(w_n415_0[0]),.dinb(w_n406_5[0]),.dout(n419),.clk(gclk));
	jand g0119(.dina(w_G308_1[0]),.dinb(w_n408_5[1]),.dout(n420),.clk(gclk));
	jor g0120(.dina(n420),.dinb(n419),.dout(n421),.clk(gclk));
	jor g0121(.dina(n421),.dinb(w_G479_0[1]),.dout(n422),.clk(gclk));
	jand g0122(.dina(n422),.dinb(n418),.dout(n423),.clk(gclk));
	jand g0123(.dina(w_n423_0[2]),.dinb(w_n412_0[2]),.dout(n424),.clk(gclk));
	jnot g0124(.din(w_G293_0[2]),.dout(n425),.clk(gclk));
	jand g0125(.dina(w_n425_0[2]),.dinb(w_n406_4[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_G293_0[1]),.dinb(w_n408_5[0]),.dout(n427),.clk(gclk));
	jor g0127(.dina(n427),.dinb(n426),.dout(n428),.clk(gclk));
	jnot g0128(.din(w_G302_0[2]),.dout(n429),.clk(gclk));
	jand g0129(.dina(w_n429_0[1]),.dinb(w_n366_1[1]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G302_0[1]),.dinb(w_n369_1[1]),.dout(n431),.clk(gclk));
	jor g0131(.dina(n431),.dinb(n430),.dout(n432),.clk(gclk));
	jnot g0132(.din(n432),.dout(n433),.clk(gclk));
	jand g0133(.dina(w_n433_0[2]),.dinb(w_n428_1[1]),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G324_1[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n375_4[0]),.dinb(w_n435_2[1]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G503_2[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n378_4[0]),.dinb(w_G324_1[1]),.dout(n438),.clk(gclk));
	jor g0138(.dina(n438),.dinb(w_n437_0[1]),.dout(n439),.clk(gclk));
	jor g0139(.dina(n439),.dinb(w_dff_B_6jRaOUUu8_1),.dout(n440),.clk(gclk));
	jand g0140(.dina(w_G3546_4[1]),.dinb(w_G324_1[0]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3548_4[0]),.dinb(w_n435_2[0]),.dout(n442),.clk(gclk));
	jor g0142(.dina(n442),.dinb(w_dff_B_HCIzJQ130_1),.dout(n443),.clk(gclk));
	jor g0143(.dina(n443),.dinb(w_G503_2[0]),.dout(n444),.clk(gclk));
	jand g0144(.dina(n444),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(n434),.dout(n446),.clk(gclk));
	jand g0146(.dina(n446),.dinb(n424),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(n399),.dout(w_dff_A_Cd9m9dFW8_2),.clk(gclk));
	jnot g0148(.din(w_G210_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n375_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G457_1[2]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n378_3[2]),.dinb(w_G210_2[0]),.dout(n452),.clk(gclk));
	jor g0152(.dina(n452),.dinb(w_n451_0[2]),.dout(n453),.clk(gclk));
	jor g0153(.dina(n453),.dinb(w_dff_B_19v3Jvts2_1),.dout(n454),.clk(gclk));
	jand g0154(.dina(w_G3546_4[0]),.dinb(w_G210_1[2]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n456),.clk(gclk));
	jor g0156(.dina(n456),.dinb(w_dff_B_zSbUmewt1_1),.dout(n457),.clk(gclk));
	jor g0157(.dina(n457),.dinb(w_G457_1[1]),.dout(n458),.clk(gclk));
	jand g0158(.dina(n458),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n375_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n378_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jor g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464),.clk(gclk));
	jor g0164(.dina(n464),.dinb(w_dff_B_Xl5HX38I0_1),.dout(n465),.clk(gclk));
	jand g0165(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n467),.clk(gclk));
	jor g0167(.dina(n467),.dinb(w_dff_B_iLPynGW98_1),.dout(n468),.clk(gclk));
	jor g0168(.dina(n468),.dinb(w_G435_1[1]),.dout(n469),.clk(gclk));
	jand g0169(.dina(n469),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G273_2[1]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n375_3[0]),.dinb(w_n471_1[2]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G411_2[1]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n378_3[0]),.dinb(w_G273_2[0]),.dout(n474),.clk(gclk));
	jor g0174(.dina(n474),.dinb(w_n473_1[1]),.dout(n475),.clk(gclk));
	jor g0175(.dina(n475),.dinb(w_dff_B_aQUqQRTG7_1),.dout(n476),.clk(gclk));
	jand g0176(.dina(w_G3546_3[1]),.dinb(w_G273_1[2]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3548_3[0]),.dinb(w_n471_1[1]),.dout(n478),.clk(gclk));
	jor g0178(.dina(n478),.dinb(w_dff_B_3XH3aMG67_1),.dout(n479),.clk(gclk));
	jor g0179(.dina(n479),.dinb(w_G411_2[0]),.dout(n480),.clk(gclk));
	jand g0180(.dina(n480),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jnot g0182(.din(w_G265_1[2]),.dout(n483),.clk(gclk));
	jand g0183(.dina(w_n375_2[2]),.dinb(w_n483_2[1]),.dout(n484),.clk(gclk));
	jnot g0184(.din(w_G400_1[2]),.dout(n485),.clk(gclk));
	jand g0185(.dina(w_n378_2[2]),.dinb(w_G265_1[1]),.dout(n486),.clk(gclk));
	jor g0186(.dina(n486),.dinb(w_n485_1[1]),.dout(n487),.clk(gclk));
	jor g0187(.dina(n487),.dinb(w_dff_B_u09SE55u4_1),.dout(n488),.clk(gclk));
	jand g0188(.dina(w_G3546_3[0]),.dinb(w_G265_1[0]),.dout(n489),.clk(gclk));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n483_2[0]),.dout(n490),.clk(gclk));
	jor g0190(.dina(n490),.dinb(w_dff_B_ebyXWjon0_1),.dout(n491),.clk(gclk));
	jor g0191(.dina(n491),.dinb(w_G400_1[1]),.dout(n492),.clk(gclk));
	jand g0192(.dina(n492),.dinb(n488),.dout(n493),.clk(gclk));
	jnot g0193(.din(w_G226_2[1]),.dout(n494),.clk(gclk));
	jand g0194(.dina(w_n375_2[1]),.dinb(w_n494_1[2]),.dout(n495),.clk(gclk));
	jnot g0195(.din(w_G422_1[1]),.dout(n496),.clk(gclk));
	jand g0196(.dina(w_n378_2[1]),.dinb(w_G226_2[0]),.dout(n497),.clk(gclk));
	jor g0197(.dina(n497),.dinb(w_n496_1[1]),.dout(n498),.clk(gclk));
	jor g0198(.dina(n498),.dinb(w_dff_B_NJkMpDqu5_1),.dout(n499),.clk(gclk));
	jand g0199(.dina(w_G3546_2[2]),.dinb(w_G226_1[2]),.dout(n500),.clk(gclk));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n494_1[1]),.dout(n501),.clk(gclk));
	jor g0201(.dina(n501),.dinb(w_dff_B_0aVBOMGB7_1),.dout(n502),.clk(gclk));
	jor g0202(.dina(n502),.dinb(w_G422_1[0]),.dout(n503),.clk(gclk));
	jand g0203(.dina(n503),.dinb(n499),.dout(n504),.clk(gclk));
	jand g0204(.dina(w_n504_0[1]),.dinb(w_n493_0[1]),.dout(n505),.clk(gclk));
	jand g0205(.dina(n505),.dinb(n482),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[1]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n375_2[0]),.dinb(w_n507_1[2]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n378_2[0]),.dinb(w_G218_2[0]),.dout(n510),.clk(gclk));
	jor g0210(.dina(n510),.dinb(w_n509_0[2]),.dout(n511),.clk(gclk));
	jor g0211(.dina(n511),.dinb(w_dff_B_NqMwqEwj1_1),.dout(n512),.clk(gclk));
	jand g0212(.dina(w_G3546_2[1]),.dinb(w_G218_1[2]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3548_2[0]),.dinb(w_n507_1[1]),.dout(n514),.clk(gclk));
	jor g0214(.dina(n514),.dinb(w_dff_B_zM4vQe9H9_1),.dout(n515),.clk(gclk));
	jor g0215(.dina(n515),.dinb(w_G468_1[1]),.dout(n516),.clk(gclk));
	jand g0216(.dina(n516),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G257_2[1]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_n375_1[2]),.dinb(w_n518_1[2]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G389_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_n378_1[2]),.dinb(w_G257_2[0]),.dout(n521),.clk(gclk));
	jor g0221(.dina(n521),.dinb(w_n520_0[2]),.dout(n522),.clk(gclk));
	jor g0222(.dina(n522),.dinb(w_dff_B_Icuqqmhk5_1),.dout(n523),.clk(gclk));
	jand g0223(.dina(w_G3546_2[0]),.dinb(w_G257_1[2]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_G3548_1[2]),.dinb(w_n518_1[1]),.dout(n525),.clk(gclk));
	jor g0225(.dina(n525),.dinb(w_dff_B_4tWlY9bq3_1),.dout(n526),.clk(gclk));
	jor g0226(.dina(n526),.dinb(w_G389_1[1]),.dout(n527),.clk(gclk));
	jand g0227(.dina(n527),.dinb(n523),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[1]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G281_2[1]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n375_1[1]),.dinb(w_n530_1[2]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G374_1[2]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n378_1[1]),.dinb(w_G281_2[0]),.dout(n533),.clk(gclk));
	jor g0233(.dina(n533),.dinb(w_n532_1[1]),.dout(n534),.clk(gclk));
	jor g0234(.dina(n534),.dinb(w_dff_B_vfk6ABnv7_1),.dout(n535),.clk(gclk));
	jand g0235(.dina(w_G3546_1[2]),.dinb(w_G281_1[2]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3548_1[1]),.dinb(w_n530_1[1]),.dout(n537),.clk(gclk));
	jor g0237(.dina(n537),.dinb(w_dff_B_QgSZRQ2D7_1),.dout(n538),.clk(gclk));
	jor g0238(.dina(n538),.dinb(w_G374_1[1]),.dout(n539),.clk(gclk));
	jand g0239(.dina(n539),.dinb(n535),.dout(n540),.clk(gclk));
	jand g0240(.dina(w_G248_4[2]),.dinb(w_G206_1[2]),.dout(n541),.clk(gclk));
	jnot g0241(.din(w_G446_1[2]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G206_1[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_G251_4[1]),.dinb(w_n543_0[1]),.dout(n544),.clk(gclk));
	jor g0244(.dina(n544),.dinb(w_dff_B_urOdmBcw5_1),.dout(n545),.clk(gclk));
	jor g0245(.dina(n545),.dinb(w_dff_B_z34FMFxU3_1),.dout(n546),.clk(gclk));
	jand g0246(.dina(w_n406_4[1]),.dinb(w_n543_0[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_n408_4[2]),.dinb(w_G206_1[0]),.dout(n548),.clk(gclk));
	jor g0248(.dina(n548),.dinb(n547),.dout(n549),.clk(gclk));
	jor g0249(.dina(n549),.dinb(w_G446_1[1]),.dout(n550),.clk(gclk));
	jand g0250(.dina(n550),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[2]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(n506),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_n459_0[1]),.dout(w_dff_A_ZvM57l6Z2_2),.clk(gclk));
	jnot g0255(.din(w_G335_0[2]),.dout(n556),.clk(gclk));
	jand g0256(.dina(w_n556_8[1]),.dinb(w_n530_1[0]),.dout(n557),.clk(gclk));
	jnot g0257(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jor g0258(.dina(w_n556_8[0]),.dinb(w_dff_B_npbHaFo88_1),.dout(n559),.clk(gclk));
	jand g0259(.dina(w_n559_0[1]),.dinb(n558),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_0[2]),.dinb(w_G374_1[0]),.dout(n561),.clk(gclk));
	jand g0261(.dina(w_n556_7[2]),.dinb(w_n471_1[0]),.dout(n562),.clk(gclk));
	jnot g0262(.din(w_n562_0[1]),.dout(n563),.clk(gclk));
	jor g0263(.dina(w_n556_7[1]),.dinb(w_dff_B_2qOmZ1NT3_1),.dout(n564),.clk(gclk));
	jand g0264(.dina(w_n564_0[1]),.dinb(n563),.dout(n565),.clk(gclk));
	jxor g0265(.dina(w_n565_0[2]),.dinb(w_G411_1[2]),.dout(n566),.clk(gclk));
	jand g0266(.dina(w_n566_0[2]),.dinb(w_n561_1[1]),.dout(n567),.clk(gclk));
	jnot g0267(.din(w_n567_0[2]),.dout(n568),.clk(gclk));
	jand g0268(.dina(w_n556_7[0]),.dinb(w_n483_1[2]),.dout(n569),.clk(gclk));
	jnot g0269(.din(w_n569_0[1]),.dout(n570),.clk(gclk));
	jor g0270(.dina(w_n556_6[2]),.dinb(w_dff_B_5xHzJPFB5_1),.dout(n571),.clk(gclk));
	jand g0271(.dina(w_n571_0[1]),.dinb(n570),.dout(n572),.clk(gclk));
	jxor g0272(.dina(w_n572_0[2]),.dinb(w_G400_1[0]),.dout(n573),.clk(gclk));
	jnot g0273(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jand g0274(.dina(w_n556_6[1]),.dinb(w_n518_1[0]),.dout(n575),.clk(gclk));
	jnot g0275(.din(n575),.dout(n576),.clk(gclk));
	jor g0276(.dina(w_n556_6[0]),.dinb(w_dff_B_7BuA7NsW1_1),.dout(n577),.clk(gclk));
	jand g0277(.dina(w_dff_B_U3UaKWHr1_0),.dinb(n576),.dout(n578),.clk(gclk));
	jxor g0278(.dina(w_n578_1[1]),.dinb(w_n520_0[1]),.dout(n579),.clk(gclk));
	jor g0279(.dina(w_n579_1[1]),.dinb(w_n574_0[2]),.dout(n580),.clk(gclk));
	jor g0280(.dina(n580),.dinb(n568),.dout(n581),.clk(gclk));
	jnot g0281(.din(w_n581_0[1]),.dout(n582),.clk(gclk));
	jand g0282(.dina(w_n556_5[2]),.dinb(w_n460_1[0]),.dout(n583),.clk(gclk));
	jnot g0283(.din(n583),.dout(n584),.clk(gclk));
	jor g0284(.dina(w_n556_5[1]),.dinb(w_dff_B_X5fR3mvU3_1),.dout(n585),.clk(gclk));
	jand g0285(.dina(w_dff_B_fmvCkGY62_0),.dinb(n584),.dout(n586),.clk(gclk));
	jxor g0286(.dina(w_n586_1[1]),.dinb(w_G435_1[0]),.dout(n587),.clk(gclk));
	jand g0287(.dina(w_n587_0[1]),.dinb(n582),.dout(n588),.clk(gclk));
	jor g0288(.dina(w_G335_0[1]),.dinb(w_G206_0[2]),.dout(n589),.clk(gclk));
	jor g0289(.dina(w_n556_5[0]),.dinb(w_dff_B_2HPg2p4d3_1),.dout(n590),.clk(gclk));
	jand g0290(.dina(n590),.dinb(w_dff_B_KjkXO6uF3_1),.dout(n591),.clk(gclk));
	jxor g0291(.dina(w_n591_1[1]),.dinb(w_G446_1[0]),.dout(n592),.clk(gclk));
	jand g0292(.dina(w_n556_4[2]),.dinb(w_n494_1[0]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jor g0294(.dina(w_n556_4[1]),.dinb(w_dff_B_cgsVAW2z9_1),.dout(n595),.clk(gclk));
	jand g0295(.dina(w_dff_B_vL2FhdQC8_0),.dinb(n594),.dout(n596),.clk(gclk));
	jxor g0296(.dina(w_n596_1[1]),.dinb(w_n496_1[0]),.dout(n597),.clk(gclk));
	jand g0297(.dina(w_n556_4[0]),.dinb(w_n507_1[0]),.dout(n598),.clk(gclk));
	jnot g0298(.din(n598),.dout(n599),.clk(gclk));
	jor g0299(.dina(w_n556_3[2]),.dinb(w_dff_B_RwubvhTj3_1),.dout(n600),.clk(gclk));
	jand g0300(.dina(w_dff_B_4gpgBaTR1_0),.dinb(n599),.dout(n601),.clk(gclk));
	jxor g0301(.dina(w_n601_1[1]),.dinb(w_n509_0[1]),.dout(n602),.clk(gclk));
	jor g0302(.dina(w_n602_0[2]),.dinb(w_n597_0[2]),.dout(n603),.clk(gclk));
	jand g0303(.dina(w_n556_3[1]),.dinb(w_n449_1[0]),.dout(n604),.clk(gclk));
	jnot g0304(.din(n604),.dout(n605),.clk(gclk));
	jor g0305(.dina(w_n556_3[0]),.dinb(w_dff_B_WRS1WKld4_1),.dout(n606),.clk(gclk));
	jand g0306(.dina(w_dff_B_D4fOFHL32_0),.dinb(n605),.dout(n607),.clk(gclk));
	jxor g0307(.dina(w_n607_1[1]),.dinb(w_n451_0[1]),.dout(n608),.clk(gclk));
	jor g0308(.dina(w_n608_0[2]),.dinb(w_n603_0[1]),.dout(n609),.clk(gclk));
	jnot g0309(.din(w_n609_0[2]),.dout(n610),.clk(gclk));
	jand g0310(.dina(n610),.dinb(w_n592_0[2]),.dout(n611),.clk(gclk));
	jand g0311(.dina(w_n611_0[2]),.dinb(w_n588_1[1]),.dout(w_dff_A_NVY0g9Mn7_2),.clk(gclk));
	jnot g0312(.din(w_G332_3[2]),.dout(n613),.clk(gclk));
	jand g0313(.dina(w_n613_5[2]),.dinb(w_n435_1[2]),.dout(n614),.clk(gclk));
	jnot g0314(.din(n614),.dout(n615),.clk(gclk));
	jor g0315(.dina(w_n613_5[1]),.dinb(w_G331_0[1]),.dout(n616),.clk(gclk));
	jand g0316(.dina(w_dff_B_XT6WQqUp7_0),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_G503_1[2]),.dout(n618),.clk(gclk));
	jor g0318(.dina(w_G338_0[0]),.dinb(w_n613_5[0]),.dout(n619),.clk(gclk));
	jxor g0319(.dina(w_n619_1[2]),.dinb(w_G514_1[2]),.dout(n620),.clk(gclk));
	jor g0320(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n621),.clk(gclk));
	jor g0321(.dina(w_G348_0[0]),.dinb(w_n613_4[2]),.dout(n622),.clk(gclk));
	jand g0322(.dina(n622),.dinb(w_n621_0[1]),.dout(n623),.clk(gclk));
	jxor g0323(.dina(w_n623_0[1]),.dinb(w_G523_1[0]),.dout(n624),.clk(gclk));
	jor g0324(.dina(w_G351_1[2]),.dinb(w_G332_3[0]),.dout(n625),.clk(gclk));
	jor g0325(.dina(w_G358_0[0]),.dinb(w_n613_4[1]),.dout(n626),.clk(gclk));
	jand g0326(.dina(n626),.dinb(w_n625_0[1]),.dout(n627),.clk(gclk));
	jor g0327(.dina(w_n627_1[1]),.dinb(w_G534_1[2]),.dout(n628),.clk(gclk));
	jnot g0328(.din(w_n625_0[0]),.dout(n629),.clk(gclk));
	jand g0329(.dina(w_G612_0),.dinb(w_G332_2[2]),.dout(n630),.clk(gclk));
	jor g0330(.dina(n630),.dinb(n629),.dout(n631),.clk(gclk));
	jor g0331(.dina(w_n631_0[1]),.dinb(w_n377_1[0]),.dout(n632),.clk(gclk));
	jor g0332(.dina(w_G361_0[2]),.dinb(w_G332_2[1]),.dout(n633),.clk(gclk));
	jor g0333(.dina(w_G366_0[0]),.dinb(w_n613_4[0]),.dout(n634),.clk(gclk));
	jand g0334(.dina(n634),.dinb(w_dff_B_D4YMhMGO0_1),.dout(n635),.clk(gclk));
	jnot g0335(.din(w_n635_1[1]),.dout(n636),.clk(gclk));
	jand g0336(.dina(w_n636_0[2]),.dinb(w_n632_0[1]),.dout(n637),.clk(gclk));
	jand g0337(.dina(w_n637_0[2]),.dinb(w_n628_0[2]),.dout(n638),.clk(gclk));
	jand g0338(.dina(w_n638_0[1]),.dinb(w_n624_0[2]),.dout(n639),.clk(gclk));
	jand g0339(.dina(w_n639_0[2]),.dinb(w_n620_1[1]),.dout(n640),.clk(gclk));
	jand g0340(.dina(w_n640_0[1]),.dinb(w_n618_0[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n613_3[2]),.dinb(w_n425_0[1]),.dout(n642),.clk(gclk));
	jand g0342(.dina(w_G332_2[0]),.dinb(w_G593_0),.dout(n643),.clk(gclk));
	jor g0343(.dina(n643),.dinb(n642),.dout(n644),.clk(gclk));
	jand g0344(.dina(w_n613_3[1]),.dinb(w_n429_0[0]),.dout(n645),.clk(gclk));
	jnot g0345(.din(n645),.dout(n646),.clk(gclk));
	jor g0346(.dina(w_n613_3[0]),.dinb(w_dff_B_TZ9GQanc9_1),.dout(n647),.clk(gclk));
	jand g0347(.dina(w_dff_B_LqUkf7YI2_0),.dinb(n646),.dout(n648),.clk(gclk));
	jnot g0348(.din(w_n648_1[1]),.dout(n649),.clk(gclk));
	jand g0349(.dina(w_n649_0[1]),.dinb(w_n644_0[2]),.dout(n650),.clk(gclk));
	jor g0350(.dina(w_G332_1[2]),.dinb(w_G308_0[2]),.dout(n651),.clk(gclk));
	jor g0351(.dina(w_n613_2[2]),.dinb(w_dff_B_TkDvYJKb3_1),.dout(n652),.clk(gclk));
	jand g0352(.dina(n652),.dinb(w_dff_B_4pBthudu4_1),.dout(n653),.clk(gclk));
	jxor g0353(.dina(w_n653_0[2]),.dinb(w_G479_0[0]),.dout(n654),.clk(gclk));
	jand g0354(.dina(w_n613_2[1]),.dinb(w_n402_0[0]),.dout(n655),.clk(gclk));
	jnot g0355(.din(n655),.dout(n656),.clk(gclk));
	jor g0356(.dina(w_n613_2[0]),.dinb(w_dff_B_jWYeyIKN8_1),.dout(n657),.clk(gclk));
	jand g0357(.dina(w_dff_B_yFdrxyFS0_0),.dinb(n656),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_n658_1[1]),.dinb(w_G490_0[2]),.dout(n659),.clk(gclk));
	jand g0359(.dina(w_n659_0[1]),.dinb(w_n654_2[2]),.dout(n660),.clk(gclk));
	jand g0360(.dina(w_n660_1[1]),.dinb(w_n650_0[1]),.dout(n661),.clk(gclk));
	jand g0361(.dina(w_n661_0[1]),.dinb(w_n641_1[2]),.dout(w_dff_A_mk7Y1tBd1_2),.clk(gclk));
	jxor g0362(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G302_0[0]),.dinb(w_n425_0[0]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(w_dff_B_6lPqW0NK3_1),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G369_0[1]),.dinb(w_G361_0[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(n666),.dinb(w_n435_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n668),.clk(gclk));
	jxor g0368(.dina(w_dff_B_T9BYHnEv1_0),.dinb(n667),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n665),.dout(n670),.clk(gclk));
	jnot g0370(.din(w_n670_0[1]),.dout(w_dff_A_jptqbv0j0_1),.clk(gclk));
	jxor g0371(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n672),.clk(gclk));
	jxor g0372(.dina(w_G273_1[1]),.dinb(w_n483_1[1]),.dout(n673),.clk(gclk));
	jxor g0373(.dina(n673),.dinb(w_dff_B_fJLKRzUl4_1),.dout(n674),.clk(gclk));
	jxor g0374(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n675),.clk(gclk));
	jxor g0375(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n676),.clk(gclk));
	jxor g0376(.dina(n676),.dinb(n675),.dout(n677),.clk(gclk));
	jxor g0377(.dina(w_G210_1[1]),.dinb(w_G206_0[1]),.dout(n678),.clk(gclk));
	jxor g0378(.dina(w_dff_B_GktndBhK1_0),.dinb(n677),.dout(n679),.clk(gclk));
	jxor g0379(.dina(n679),.dinb(n674),.dout(n680),.clk(gclk));
	jnot g0380(.din(w_n680_0[1]),.dout(w_dff_A_Pd8CgEzt0_1),.clk(gclk));
	jand g0381(.dina(w_n586_1[0]),.dinb(w_G435_0[2]),.dout(n682),.clk(gclk));
	jnot g0382(.din(w_n586_0[2]),.dout(n683),.clk(gclk));
	jand g0383(.dina(n683),.dinb(w_n462_0[1]),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n684_0[1]),.dout(n685),.clk(gclk));
	jand g0385(.dina(w_n578_1[0]),.dinb(w_G389_1[0]),.dout(n686),.clk(gclk));
	jor g0386(.dina(w_n578_0[2]),.dinb(w_G389_0[2]),.dout(n687),.clk(gclk));
	jnot g0387(.din(w_n571_0[0]),.dout(n688),.clk(gclk));
	jor g0388(.dina(n688),.dinb(w_n569_0[0]),.dout(n689),.clk(gclk));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n485_1[0]),.dout(n690),.clk(gclk));
	jnot g0390(.din(w_n690_0[1]),.dout(n691),.clk(gclk));
	jand g0391(.dina(w_n560_0[1]),.dinb(w_G374_0[2]),.dout(n692),.clk(gclk));
	jor g0392(.dina(w_n565_0[1]),.dinb(w_G411_1[1]),.dout(n693),.clk(gclk));
	jand g0393(.dina(n693),.dinb(w_n692_0[1]),.dout(n694),.clk(gclk));
	jand g0394(.dina(w_n565_0[0]),.dinb(w_G411_1[0]),.dout(n695),.clk(gclk));
	jand g0395(.dina(w_n572_0[1]),.dinb(w_G400_0[2]),.dout(n696),.clk(gclk));
	jor g0396(.dina(n696),.dinb(w_n695_0[2]),.dout(n697),.clk(gclk));
	jor g0397(.dina(n697),.dinb(w_n694_0[2]),.dout(n698),.clk(gclk));
	jand g0398(.dina(n698),.dinb(w_dff_B_ZNUr6u3F5_1),.dout(n699),.clk(gclk));
	jand g0399(.dina(w_n699_0[2]),.dinb(w_n687_0[1]),.dout(n700),.clk(gclk));
	jor g0400(.dina(n700),.dinb(w_n686_0[1]),.dout(n701),.clk(gclk));
	jand g0401(.dina(w_n701_0[1]),.dinb(w_n685_0[1]),.dout(n702),.clk(gclk));
	jor g0402(.dina(n702),.dinb(w_n682_0[2]),.dout(n703),.clk(gclk));
	jand g0403(.dina(w_n703_0[2]),.dinb(w_n611_0[1]),.dout(n704),.clk(gclk));
	jand g0404(.dina(w_n591_1[0]),.dinb(w_G446_0[2]),.dout(n705),.clk(gclk));
	jor g0405(.dina(w_n591_0[2]),.dinb(w_G446_0[1]),.dout(n706),.clk(gclk));
	jand g0406(.dina(w_n607_1[0]),.dinb(w_G457_1[0]),.dout(n707),.clk(gclk));
	jor g0407(.dina(w_n607_0[2]),.dinb(w_G457_0[2]),.dout(n708),.clk(gclk));
	jand g0408(.dina(w_n601_1[0]),.dinb(w_G468_1[0]),.dout(n709),.clk(gclk));
	jand g0409(.dina(w_n596_1[0]),.dinb(w_G422_0[2]),.dout(n710),.clk(gclk));
	jor g0410(.dina(w_n601_0[2]),.dinb(w_G468_0[2]),.dout(n711),.clk(gclk));
	jand g0411(.dina(w_n711_0[1]),.dinb(w_n710_0[1]),.dout(n712),.clk(gclk));
	jor g0412(.dina(n712),.dinb(w_n709_0[1]),.dout(n713),.clk(gclk));
	jand g0413(.dina(w_n713_0[2]),.dinb(w_dff_B_6oCEeYCx3_1),.dout(n714),.clk(gclk));
	jor g0414(.dina(n714),.dinb(w_dff_B_18LzI1ED4_1),.dout(n715),.clk(gclk));
	jand g0415(.dina(w_n715_0[2]),.dinb(w_dff_B_cb2UIZEQ3_1),.dout(n716),.clk(gclk));
	jor g0416(.dina(n716),.dinb(w_dff_B_9A2iSTBK3_1),.dout(n717),.clk(gclk));
	jor g0417(.dina(w_n717_0[1]),.dinb(w_n704_0[1]),.dout(w_dff_A_q1kryMCV0_2),.clk(gclk));
	jand g0418(.dina(w_n617_1[0]),.dinb(w_G503_1[1]),.dout(n719),.clk(gclk));
	jor g0419(.dina(w_n617_0[2]),.dinb(w_G503_1[0]),.dout(n720),.clk(gclk));
	jor g0420(.dina(w_n619_1[1]),.dinb(w_G514_1[1]),.dout(n721),.clk(gclk));
	jand g0421(.dina(w_n619_1[0]),.dinb(w_G514_1[0]),.dout(n722),.clk(gclk));
	jnot g0422(.din(w_n621_0[0]),.dout(n723),.clk(gclk));
	jand g0423(.dina(w_G599_0),.dinb(w_G332_1[1]),.dout(n724),.clk(gclk));
	jor g0424(.dina(n724),.dinb(n723),.dout(n725),.clk(gclk));
	jand g0425(.dina(w_n725_0[2]),.dinb(w_n389_1[0]),.dout(n726),.clk(gclk));
	jnot g0426(.din(w_n726_0[1]),.dout(n727),.clk(gclk));
	jand g0427(.dina(w_n635_1[0]),.dinb(w_n628_0[1]),.dout(n728),.clk(gclk));
	jand g0428(.dina(w_n623_0[0]),.dinb(w_G523_0[2]),.dout(n729),.clk(gclk));
	jand g0429(.dina(w_n627_1[0]),.dinb(w_G534_1[1]),.dout(n730),.clk(gclk));
	jor g0430(.dina(n730),.dinb(n729),.dout(n731),.clk(gclk));
	jor g0431(.dina(n731),.dinb(w_n728_0[1]),.dout(n732),.clk(gclk));
	jand g0432(.dina(n732),.dinb(w_dff_B_sQM3zmHS5_1),.dout(n733),.clk(gclk));
	jor g0433(.dina(w_n733_0[2]),.dinb(w_n722_0[1]),.dout(n734),.clk(gclk));
	jand g0434(.dina(n734),.dinb(w_n721_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[2]),.dinb(w_n720_0[1]),.dout(n736),.clk(gclk));
	jor g0436(.dina(n736),.dinb(w_n719_0[1]),.dout(n737),.clk(gclk));
	jand g0437(.dina(w_n737_1[1]),.dinb(w_n660_1[0]),.dout(n738),.clk(gclk));
	jnot g0438(.din(w_n650_0[0]),.dout(n739),.clk(gclk));
	jnot g0439(.din(w_n653_0[1]),.dout(n740),.clk(gclk));
	jor g0440(.dina(n740),.dinb(w_n414_0[0]),.dout(n741),.clk(gclk));
	jand g0441(.dina(w_n658_1[0]),.dinb(w_G490_0[1]),.dout(n742),.clk(gclk));
	jand g0442(.dina(w_n742_0[2]),.dinb(w_n654_2[1]),.dout(n743),.clk(gclk));
	jnot g0443(.din(n743),.dout(n744),.clk(gclk));
	jand g0444(.dina(n744),.dinb(w_dff_B_w5V504Yr2_1),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_n745_0[1]),.dout(n746),.clk(gclk));
	jor g0446(.dina(w_n746_0[2]),.dinb(w_dff_B_lgf4lBax9_1),.dout(n747),.clk(gclk));
	jor g0447(.dina(w_n747_0[1]),.dinb(w_n738_0[1]),.dout(w_dff_A_LaQp9IAo6_2),.clk(gclk));
	jnot g0448(.din(w_G4091_6[1]),.dout(n749),.clk(gclk));
	jand g0449(.dina(w_G4092_9[2]),.dinb(w_n749_13[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n750_8[2]),.dinb(w_dff_B_QCr6Roxr9_1),.dout(n751),.clk(gclk));
	jnot g0451(.din(n751),.dout(n752),.clk(gclk));
	jnot g0452(.din(w_G54_0[2]),.dout(n753),.clk(gclk));
	jxor g0453(.dina(w_n635_0[2]),.dinb(w_n753_1[1]),.dout(n754),.clk(gclk));
	jnot g0454(.din(n754),.dout(n755),.clk(gclk));
	jand g0455(.dina(w_n755_0[1]),.dinb(w_G4091_6[0]),.dout(n756),.clk(gclk));
	jand g0456(.dina(w_n372_0[0]),.dinb(w_n749_13[0]),.dout(n757),.clk(gclk));
	jor g0457(.dina(n757),.dinb(w_G4092_9[1]),.dout(n758),.clk(gclk));
	jor g0458(.dina(n758),.dinb(n756),.dout(n759),.clk(gclk));
	jand g0459(.dina(n759),.dinb(w_dff_B_9CjPmnQA1_1),.dout(G822_fa_),.clk(gclk));
	jand g0460(.dina(w_n750_8[1]),.dinb(w_dff_B_3PWJPcsw6_1),.dout(n761),.clk(gclk));
	jnot g0461(.din(n761),.dout(n762),.clk(gclk));
	jxor g0462(.dina(w_n627_0[2]),.dinb(w_G534_1[0]),.dout(n763),.clk(gclk));
	jnot g0463(.din(w_n763_0[2]),.dout(n764),.clk(gclk));
	jand g0464(.dina(n764),.dinb(w_n635_0[1]),.dout(n765),.clk(gclk));
	jor g0465(.dina(n765),.dinb(w_n638_0[0]),.dout(n766),.clk(gclk));
	jnot g0466(.din(n766),.dout(n767),.clk(gclk));
	jand g0467(.dina(w_n767_0[1]),.dinb(w_n753_1[0]),.dout(n768),.clk(gclk));
	jand g0468(.dina(w_n763_0[1]),.dinb(w_G54_0[1]),.dout(n769),.clk(gclk));
	jor g0469(.dina(w_dff_B_xI1S3T0I1_0),.dinb(n768),.dout(n770),.clk(gclk));
	jand g0470(.dina(n770),.dinb(w_G4091_5[2]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n386_0[0]),.dinb(w_n749_12[2]),.dout(n772),.clk(gclk));
	jor g0472(.dina(n772),.dinb(w_G4092_9[0]),.dout(n773),.clk(gclk));
	jor g0473(.dina(w_dff_B_5OSjEKub0_0),.dinb(n771),.dout(n774),.clk(gclk));
	jand g0474(.dina(n774),.dinb(w_dff_B_W86gbJTr4_1),.dout(G838_fa_),.clk(gclk));
	jand g0475(.dina(w_n750_8[0]),.dinb(w_dff_B_6cjba8ES8_1),.dout(n776),.clk(gclk));
	jnot g0476(.din(n776),.dout(n777),.clk(gclk));
	jxor g0477(.dina(w_n561_1[0]),.dinb(w_G4_0[2]),.dout(n778),.clk(gclk));
	jnot g0478(.din(n778),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n779_0[1]),.dinb(w_G4091_5[1]),.dout(n780),.clk(gclk));
	jand g0480(.dina(w_n540_0[0]),.dinb(w_n749_12[1]),.dout(n781),.clk(gclk));
	jor g0481(.dina(n781),.dinb(w_G4092_8[2]),.dout(n782),.clk(gclk));
	jor g0482(.dina(w_dff_B_zK5ZTSk17_0),.dinb(n780),.dout(n783),.clk(gclk));
	jand g0483(.dina(n783),.dinb(w_dff_B_8ZKG8dxr1_1),.dout(G861_fa_),.clk(gclk));
	jand g0484(.dina(w_n641_1[1]),.dinb(w_G54_0[0]),.dout(n785),.clk(gclk));
	jor g0485(.dina(w_dff_B_JsXWV9FB2_0),.dinb(w_n737_1[0]),.dout(n786),.clk(gclk));
	jand g0486(.dina(w_n786_0[2]),.dinb(w_n660_0[2]),.dout(n787),.clk(gclk));
	jor g0487(.dina(n787),.dinb(w_n746_0[1]),.dout(n788),.clk(gclk));
	jnot g0488(.din(w_n788_0[2]),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n644_0[1]),.dout(n790),.clk(gclk));
	jxor g0490(.dina(w_n648_1[0]),.dinb(w_n790_0[2]),.dout(n791),.clk(gclk));
	jnot g0491(.din(n791),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_n792_0[2]),.dinb(n789),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n788_0[1]),.dinb(w_n790_0[1]),.dout(n794),.clk(gclk));
	jor g0494(.dina(w_dff_B_teBg1fcI7_0),.dinb(n793),.dout(n795),.clk(gclk));
	jnot g0495(.din(w_n795_1[1]),.dout(G623_fa_),.clk(gclk));
	jnot g0496(.din(w_G4088_9[2]),.dout(n797),.clk(gclk));
	jnot g0497(.din(w_G861_0),.dout(n798),.clk(gclk));
	jor g0498(.dina(w_n798_1[1]),.dinb(w_n797_9[1]),.dout(n799),.clk(gclk));
	jnot g0499(.din(w_G4087_4[2]),.dout(n800),.clk(gclk));
	jnot g0500(.din(w_G822_0),.dout(n801),.clk(gclk));
	jor g0501(.dina(w_n801_1[1]),.dinb(w_G4088_9[1]),.dout(n802),.clk(gclk));
	jand g0502(.dina(n802),.dinb(w_n800_4[1]),.dout(n803),.clk(gclk));
	jand g0503(.dina(w_dff_B_6UaTBp6x0_0),.dinb(n799),.dout(n804),.clk(gclk));
	jor g0504(.dina(w_n797_9[0]),.dinb(w_G61_0[1]),.dout(n805),.clk(gclk));
	jor g0505(.dina(w_G4088_9[0]),.dinb(w_G11_0[1]),.dout(n806),.clk(gclk));
	jand g0506(.dina(n806),.dinb(w_G4087_4[1]),.dout(n807),.clk(gclk));
	jand g0507(.dina(n807),.dinb(n805),.dout(n808),.clk(gclk));
	jor g0508(.dina(w_dff_B_YQx7uU1H6_0),.dinb(n804),.dout(w_dff_A_CgLAglrU8_2),.clk(gclk));
	jand g0509(.dina(w_n750_7[2]),.dinb(w_dff_B_PiyvcPOW4_1),.dout(n810),.clk(gclk));
	jnot g0510(.din(n810),.dout(n811),.clk(gclk));
	jnot g0511(.din(w_n721_0[0]),.dout(n812),.clk(gclk));
	jnot g0512(.din(w_n722_0[0]),.dout(n813),.clk(gclk));
	jand g0513(.dina(w_n631_0[0]),.dinb(w_n377_0[2]),.dout(n814),.clk(gclk));
	jor g0514(.dina(w_n636_0[1]),.dinb(w_n814_0[2]),.dout(n815),.clk(gclk));
	jor g0515(.dina(w_n725_0[1]),.dinb(w_n389_0[2]),.dout(n816),.clk(gclk));
	jand g0516(.dina(w_n632_0[0]),.dinb(n816),.dout(n817),.clk(gclk));
	jand g0517(.dina(n817),.dinb(n815),.dout(n818),.clk(gclk));
	jor g0518(.dina(n818),.dinb(w_n726_0[0]),.dout(n819),.clk(gclk));
	jand g0519(.dina(w_n819_0[2]),.dinb(w_dff_B_PzqaW83H4_1),.dout(n820),.clk(gclk));
	jor g0520(.dina(n820),.dinb(w_dff_B_hrLyDgLw7_1),.dout(n821),.clk(gclk));
	jnot g0521(.din(w_n620_1[0]),.dout(n822),.clk(gclk));
	jnot g0522(.din(w_n639_0[1]),.dout(n823),.clk(gclk));
	jor g0523(.dina(n823),.dinb(w_n753_0[2]),.dout(n824),.clk(gclk));
	jor g0524(.dina(w_n824_0[1]),.dinb(w_dff_B_DbDIyK689_1),.dout(n825),.clk(gclk));
	jand g0525(.dina(n825),.dinb(w_n821_0[1]),.dout(n826),.clk(gclk));
	jxor g0526(.dina(n826),.dinb(w_n618_0[1]),.dout(n827),.clk(gclk));
	jand g0527(.dina(w_n827_0[1]),.dinb(w_G4091_5[0]),.dout(n828),.clk(gclk));
	jand g0528(.dina(w_n445_0[0]),.dinb(w_n749_12[0]),.dout(n829),.clk(gclk));
	jor g0529(.dina(n829),.dinb(w_G4092_8[1]),.dout(n830),.clk(gclk));
	jor g0530(.dina(w_dff_B_qH1jI7nu0_0),.dinb(n828),.dout(n831),.clk(gclk));
	jand g0531(.dina(n831),.dinb(w_dff_B_bvhI34cd3_1),.dout(G832_fa_),.clk(gclk));
	jand g0532(.dina(w_n750_7[1]),.dinb(w_dff_B_0QuqJQqF4_1),.dout(n833),.clk(gclk));
	jnot g0533(.din(n833),.dout(n834),.clk(gclk));
	jand g0534(.dina(w_n824_0[0]),.dinb(w_n819_0[1]),.dout(n835),.clk(gclk));
	jxor g0535(.dina(n835),.dinb(w_n620_0[2]),.dout(n836),.clk(gclk));
	jand g0536(.dina(w_n836_0[1]),.dinb(w_G4091_4[2]),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_n365_0[0]),.dinb(w_n749_11[2]),.dout(n838),.clk(gclk));
	jor g0538(.dina(n838),.dinb(w_G4092_8[0]),.dout(n839),.clk(gclk));
	jor g0539(.dina(w_dff_B_YwyUonoH8_0),.dinb(n837),.dout(n840),.clk(gclk));
	jand g0540(.dina(n840),.dinb(w_dff_B_lXbCqQiA8_1),.dout(G834_fa_),.clk(gclk));
	jand g0541(.dina(w_n750_7[0]),.dinb(w_dff_B_gzn3ppYX3_1),.dout(n842),.clk(gclk));
	jnot g0542(.din(n842),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n397_0[0]),.dinb(w_n749_11[1]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_n637_0[1]),.dinb(w_n753_0[1]),.dout(n845),.clk(gclk));
	jor g0545(.dina(n845),.dinb(w_n814_0[1]),.dout(n846),.clk(gclk));
	jxor g0546(.dina(n846),.dinb(w_n624_0[1]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_0[1]),.dinb(w_G4091_4[1]),.dout(n848),.clk(gclk));
	jor g0548(.dina(n848),.dinb(w_G4092_7[2]),.dout(n849),.clk(gclk));
	jor g0549(.dina(n849),.dinb(w_dff_B_vO0YA87X3_1),.dout(n850),.clk(gclk));
	jand g0550(.dina(n850),.dinb(w_dff_B_vS45smQj3_1),.dout(G836_fa_),.clk(gclk));
	jnot g0551(.din(w_G4089_9[2]),.dout(n852),.clk(gclk));
	jor g0552(.dina(w_n798_1[0]),.dinb(w_n852_9[1]),.dout(n853),.clk(gclk));
	jnot g0553(.din(w_G4090_4[2]),.dout(n854),.clk(gclk));
	jor g0554(.dina(w_n801_1[0]),.dinb(w_G4089_9[1]),.dout(n855),.clk(gclk));
	jand g0555(.dina(n855),.dinb(w_n854_4[1]),.dout(n856),.clk(gclk));
	jand g0556(.dina(w_dff_B_0IFzQppa9_0),.dinb(n853),.dout(n857),.clk(gclk));
	jor g0557(.dina(w_n852_9[0]),.dinb(w_G61_0[0]),.dout(n858),.clk(gclk));
	jor g0558(.dina(w_G4089_9[0]),.dinb(w_G11_0[0]),.dout(n859),.clk(gclk));
	jand g0559(.dina(n859),.dinb(w_G4090_4[1]),.dout(n860),.clk(gclk));
	jand g0560(.dina(n860),.dinb(n858),.dout(n861),.clk(gclk));
	jor g0561(.dina(w_dff_B_9jj3DoR38_0),.dinb(n857),.dout(w_dff_A_WzDV50rL1_2),.clk(gclk));
	jand g0562(.dina(w_n750_6[2]),.dinb(w_dff_B_qakfyPmS7_1),.dout(n863),.clk(gclk));
	jnot g0563(.din(n863),.dout(n864),.clk(gclk));
	jnot g0564(.din(w_n587_0[0]),.dout(n865),.clk(gclk));
	jnot g0565(.din(w_n579_1[0]),.dout(n866),.clk(gclk));
	jand g0566(.dina(w_n567_0[1]),.dinb(w_G4_0[1]),.dout(n867),.clk(gclk));
	jand g0567(.dina(w_n867_0[1]),.dinb(w_n573_0[1]),.dout(n868),.clk(gclk));
	jand g0568(.dina(w_n868_0[1]),.dinb(w_dff_B_Hm0NnoUi5_1),.dout(n869),.clk(gclk));
	jor g0569(.dina(w_dff_B_zzQxdAZy6_0),.dinb(w_n701_0[0]),.dout(n870),.clk(gclk));
	jxor g0570(.dina(w_n870_0[1]),.dinb(w_n865_0[2]),.dout(n871),.clk(gclk));
	jand g0571(.dina(w_n871_0[1]),.dinb(w_G4091_4[0]),.dout(n872),.clk(gclk));
	jand g0572(.dina(w_n470_0[0]),.dinb(w_n749_11[0]),.dout(n873),.clk(gclk));
	jor g0573(.dina(n873),.dinb(w_G4092_7[1]),.dout(n874),.clk(gclk));
	jor g0574(.dina(w_dff_B_mXSWqqI47_0),.dinb(n872),.dout(n875),.clk(gclk));
	jand g0575(.dina(n875),.dinb(w_dff_B_WwJ0NSWx1_1),.dout(G871_fa_),.clk(gclk));
	jand g0576(.dina(w_n750_6[1]),.dinb(w_dff_B_I2URrG8P0_1),.dout(n877),.clk(gclk));
	jnot g0577(.din(n877),.dout(n878),.clk(gclk));
	jor g0578(.dina(w_n868_0[0]),.dinb(w_n699_0[1]),.dout(n879),.clk(gclk));
	jxor g0579(.dina(n879),.dinb(w_n579_0[2]),.dout(n880),.clk(gclk));
	jand g0580(.dina(w_n880_0[1]),.dinb(w_G4091_3[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n528_0[0]),.dinb(w_n749_10[2]),.dout(n882),.clk(gclk));
	jor g0582(.dina(n882),.dinb(w_G4092_7[0]),.dout(n883),.clk(gclk));
	jor g0583(.dina(w_dff_B_fte8Gnki9_0),.dinb(n881),.dout(n884),.clk(gclk));
	jand g0584(.dina(n884),.dinb(w_dff_B_EMjRTHoL2_1),.dout(G873_fa_),.clk(gclk));
	jand g0585(.dina(w_n750_6[0]),.dinb(w_dff_B_x4PZrSTy0_1),.dout(n886),.clk(gclk));
	jnot g0586(.din(n886),.dout(n887),.clk(gclk));
	jor g0587(.dina(w_n694_0[1]),.dinb(w_n695_0[1]),.dout(n888),.clk(gclk));
	jor g0588(.dina(n888),.dinb(w_n867_0[0]),.dout(n889),.clk(gclk));
	jxor g0589(.dina(n889),.dinb(w_n574_0[1]),.dout(n890),.clk(gclk));
	jand g0590(.dina(w_n890_0[1]),.dinb(w_G4091_3[1]),.dout(n891),.clk(gclk));
	jand g0591(.dina(w_n493_0[0]),.dinb(w_n749_10[1]),.dout(n892),.clk(gclk));
	jor g0592(.dina(n892),.dinb(w_G4092_6[2]),.dout(n893),.clk(gclk));
	jor g0593(.dina(w_dff_B_tjkDXg8y1_0),.dinb(n891),.dout(n894),.clk(gclk));
	jand g0594(.dina(n894),.dinb(w_dff_B_zJDkO5pI3_1),.dout(G875_fa_),.clk(gclk));
	jand g0595(.dina(w_n750_5[2]),.dinb(w_dff_B_yaRqtMlG8_1),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jnot g0597(.din(w_n566_0[1]),.dout(n898),.clk(gclk));
	jand g0598(.dina(w_n561_0[2]),.dinb(w_G4_0[0]),.dout(n899),.clk(gclk));
	jor g0599(.dina(n899),.dinb(w_n692_0[0]),.dout(n900),.clk(gclk));
	jxor g0600(.dina(n900),.dinb(w_dff_B_Bm6FwsJ27_1),.dout(n901),.clk(gclk));
	jand g0601(.dina(w_n901_0[1]),.dinb(w_G4091_3[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_n481_0[0]),.dinb(w_n749_10[0]),.dout(n903),.clk(gclk));
	jor g0603(.dina(n903),.dinb(w_G4092_6[1]),.dout(n904),.clk(gclk));
	jor g0604(.dina(w_dff_B_PgKBBWqC0_0),.dinb(n902),.dout(n905),.clk(gclk));
	jand g0605(.dina(n905),.dinb(w_dff_B_4xRmqUBc3_1),.dout(G877_fa_),.clk(gclk));
	jnot g0606(.din(w_G331_0[0]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_n619_0[2]),.dout(n908),.clk(gclk));
	jand g0608(.dina(n908),.dinb(w_dff_B_7wKi2Shd7_1),.dout(n909),.clk(gclk));
	jand g0609(.dina(w_n619_0[1]),.dinb(w_n617_0[1]),.dout(n910),.clk(gclk));
	jor g0610(.dina(n910),.dinb(w_dff_B_4gwmfbNS1_1),.dout(n911),.clk(gclk));
	jxor g0611(.dina(n911),.dinb(w_n792_0[1]),.dout(n912),.clk(gclk));
	jor g0612(.dina(w_G369_0[0]),.dinb(w_G332_1[0]),.dout(n913),.clk(gclk));
	jor g0613(.dina(w_dff_B_lJIOTZQH6_0),.dinb(w_n613_1[2]),.dout(n914),.clk(gclk));
	jand g0614(.dina(n914),.dinb(w_dff_B_qe1eSGki3_1),.dout(n915),.clk(gclk));
	jxor g0615(.dina(w_dff_B_z8WZTYfZ4_0),.dinb(w_n636_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n627_0[1]),.dinb(w_n725_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(w_n658_0[2]),.dinb(w_n653_0[0]),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_dff_B_odN55ZPf6_1),.dout(n919),.clk(gclk));
	jxor g0619(.dina(n919),.dinb(w_dff_B_TJmzSrc90_1),.dout(n920),.clk(gclk));
	jxor g0620(.dina(n920),.dinb(n912),.dout(G998_fa_),.clk(gclk));
	jnot g0621(.din(w_n564_0[0]),.dout(n922),.clk(gclk));
	jor g0622(.dina(n922),.dinb(w_n562_0[0]),.dout(n923),.clk(gclk));
	jxor g0623(.dina(w_n578_0[1]),.dinb(w_n923_0[2]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n572_0[0]),.dinb(w_n560_0[0]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jor g0626(.dina(w_G335_0[0]),.dinb(w_G289_0[0]),.dout(n927),.clk(gclk));
	jor g0627(.dina(w_n556_2[2]),.dinb(w_dff_B_LYANNG6m0_1),.dout(n928),.clk(gclk));
	jand g0628(.dina(n928),.dinb(w_dff_B_da3s2Xhl4_1),.dout(n929),.clk(gclk));
	jxor g0629(.dina(n929),.dinb(w_n591_0[1]),.dout(n930),.clk(gclk));
	jxor g0630(.dina(w_n596_0[2]),.dinb(w_n586_0[1]),.dout(n931),.clk(gclk));
	jxor g0631(.dina(w_n607_0[1]),.dinb(w_n601_0[1]),.dout(n932),.clk(gclk));
	jxor g0632(.dina(n932),.dinb(n931),.dout(n933),.clk(gclk));
	jxor g0633(.dina(n933),.dinb(w_dff_B_S0xTrdX29_1),.dout(n934),.clk(gclk));
	jxor g0634(.dina(n934),.dinb(w_dff_B_L0gb3Hkz2_1),.dout(n935),.clk(gclk));
	jnot g0635(.din(w_n935_0[1]),.dout(w_dff_A_XFSPDDuF1_1),.clk(gclk));
	jnot g0636(.din(w_n592_0[1]),.dout(n937),.clk(gclk));
	jnot g0637(.din(w_n715_0[1]),.dout(n938),.clk(gclk));
	jor g0638(.dina(w_n870_0[0]),.dinb(w_n682_0[1]),.dout(n939),.clk(gclk));
	jand g0639(.dina(n939),.dinb(w_n685_0[0]),.dout(n940),.clk(gclk));
	jnot g0640(.din(w_n940_1[1]),.dout(n941),.clk(gclk));
	jor g0641(.dina(n941),.dinb(w_n609_0[1]),.dout(n942),.clk(gclk));
	jand g0642(.dina(n942),.dinb(w_n938_0[2]),.dout(n943),.clk(gclk));
	jxor g0643(.dina(n943),.dinb(w_dff_B_Gyu7mPT03_1),.dout(n944),.clk(gclk));
	jnot g0644(.din(w_n944_0[1]),.dout(n945),.clk(gclk));
	jnot g0645(.din(w_n603_0[0]),.dout(n946),.clk(gclk));
	jand g0646(.dina(w_n940_1[0]),.dinb(w_dff_B_myCJoxAL4_1),.dout(n947),.clk(gclk));
	jor g0647(.dina(n947),.dinb(w_n713_0[1]),.dout(n948),.clk(gclk));
	jxor g0648(.dina(n948),.dinb(w_n608_0[1]),.dout(n949),.clk(gclk));
	jand g0649(.dina(w_n949_0[1]),.dinb(n945),.dout(n950),.clk(gclk));
	jnot g0650(.din(w_n602_0[1]),.dout(n951),.clk(gclk));
	jnot g0651(.din(w_n596_0[1]),.dout(n952),.clk(gclk));
	jand g0652(.dina(n952),.dinb(w_n496_0[2]),.dout(n953),.clk(gclk));
	jnot g0653(.din(w_n953_0[1]),.dout(n954),.clk(gclk));
	jor g0654(.dina(w_n940_0[2]),.dinb(w_n710_0[0]),.dout(n955),.clk(gclk));
	jand g0655(.dina(n955),.dinb(w_n954_0[2]),.dout(n956),.clk(gclk));
	jxor g0656(.dina(n956),.dinb(w_dff_B_ml053Y7a4_1),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n957_0[1]),.dout(n958),.clk(gclk));
	jand g0658(.dina(w_n890_0[0]),.dinb(w_n779_0[0]),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(w_n901_0[0]),.dout(n960),.clk(gclk));
	jand g0660(.dina(w_dff_B_LNKh3xgB8_0),.dinb(w_n871_0[0]),.dout(n961),.clk(gclk));
	jnot g0661(.din(w_n597_0[1]),.dout(n962),.clk(gclk));
	jxor g0662(.dina(w_n940_0[1]),.dinb(w_n962_0[1]),.dout(n963),.clk(gclk));
	jnot g0663(.din(n963),.dout(n964),.clk(gclk));
	jand g0664(.dina(w_n964_0[1]),.dinb(w_n880_0[0]),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(w_dff_B_RH5sCLMh0_1),.dout(n966),.clk(gclk));
	jand g0666(.dina(n966),.dinb(n958),.dout(n967),.clk(gclk));
	jand g0667(.dina(w_dff_B_QIMtgdLF5_0),.dinb(n950),.dout(w_dff_A_LojQ4O6a8_2),.clk(gclk));
	jxor g0668(.dina(w_n788_0[0]),.dinb(w_n649_0[0]),.dout(n969),.clk(gclk));
	jnot g0669(.din(w_n969_0[1]),.dout(n970),.clk(gclk));
	jand g0670(.dina(n970),.dinb(w_n755_0[0]),.dout(n971),.clk(gclk));
	jand g0671(.dina(w_n836_0[0]),.dinb(w_G623_0),.dout(n972),.clk(gclk));
	jand g0672(.dina(n972),.dinb(w_dff_B_AUY7s4db5_1),.dout(n973),.clk(gclk));
	jand g0673(.dina(w_n827_0[0]),.dinb(w_n763_0[0]),.dout(n974),.clk(gclk));
	jand g0674(.dina(n974),.dinb(w_n847_0[0]),.dout(n975),.clk(gclk));
	jnot g0675(.din(w_n658_0[1]),.dout(n976),.clk(gclk));
	jand g0676(.dina(n976),.dinb(w_n401_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(w_n977_0[2]),.dinb(w_n654_2[0]),.dout(n978),.clk(gclk));
	jor g0678(.dina(w_n977_0[1]),.dinb(w_n654_1[2]),.dout(n979),.clk(gclk));
	jnot g0679(.din(n979),.dout(n980),.clk(gclk));
	jor g0680(.dina(w_n786_0[1]),.dinb(w_n742_0[1]),.dout(n981),.clk(gclk));
	jand g0681(.dina(w_n981_0[1]),.dinb(w_dff_B_34l2otit6_1),.dout(n982),.clk(gclk));
	jnot g0682(.din(w_n981_0[0]),.dout(n983),.clk(gclk));
	jand g0683(.dina(n983),.dinb(w_n654_1[1]),.dout(n984),.clk(gclk));
	jor g0684(.dina(n984),.dinb(w_dff_B_u6qAhvxI0_1),.dout(n985),.clk(gclk));
	jor g0685(.dina(n985),.dinb(w_dff_B_moZESCAc2_1),.dout(n986),.clk(gclk));
	jnot g0686(.din(w_n986_0[1]),.dout(n987),.clk(gclk));
	jnot g0687(.din(w_n659_0[0]),.dout(n988),.clk(gclk));
	jxor g0688(.dina(w_n786_0[0]),.dinb(w_dff_B_sfEVgNFW5_1),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_n989_0[1]),.dinb(n987),.dout(n990),.clk(gclk));
	jand g0690(.dina(n990),.dinb(w_dff_B_cA5UtwHA5_1),.dout(n991),.clk(gclk));
	jand g0691(.dina(n991),.dinb(n973),.dout(w_dff_A_ifO26XYC5_2),.clk(gclk));
	jnot g0692(.din(w_G1689_5[1]),.dout(n993),.clk(gclk));
	jand g0693(.dina(w_G1690_1[1]),.dinb(w_n993_4[2]),.dout(n994),.clk(gclk));
	jand g0694(.dina(w_n994_4[1]),.dinb(w_G182_0[1]),.dout(n995),.clk(gclk));
	jand g0695(.dina(w_G1690_1[0]),.dinb(w_G1689_5[0]),.dout(n996),.clk(gclk));
	jand g0696(.dina(w_n996_4[1]),.dinb(w_G185_0[1]),.dout(n997),.clk(gclk));
	jor g0697(.dina(w_n798_0[2]),.dinb(w_n993_4[1]),.dout(n998),.clk(gclk));
	jnot g0698(.din(w_G1690_0[2]),.dout(n999),.clk(gclk));
	jor g0699(.dina(w_n801_0[2]),.dinb(w_G1689_4[2]),.dout(n1000),.clk(gclk));
	jand g0700(.dina(n1000),.dinb(w_n999_3[2]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_dff_B_LB8GxHHJ9_0),.dinb(n998),.dout(n1002),.clk(gclk));
	jor g0702(.dina(n1002),.dinb(w_dff_B_wixnft3X6_1),.dout(n1003),.clk(gclk));
	jor g0703(.dina(n1003),.dinb(w_dff_B_96gCK1kk3_1),.dout(n1004),.clk(gclk));
	jand g0704(.dina(n1004),.dinb(w_G137_9[1]),.dout(w_dff_A_FG5x9kcg6_2),.clk(gclk));
	jor g0705(.dina(w_n801_0[1]),.dinb(w_G1691_5[1]),.dout(n1006),.clk(gclk));
	jnot g0706(.din(w_G1694_1[1]),.dout(n1007),.clk(gclk));
	jnot g0707(.din(w_G1691_5[0]),.dout(n1008),.clk(gclk));
	jor g0708(.dina(w_n798_0[1]),.dinb(w_n1008_4[2]),.dout(n1009),.clk(gclk));
	jand g0709(.dina(n1009),.dinb(w_n1007_3[2]),.dout(n1010),.clk(gclk));
	jand g0710(.dina(n1010),.dinb(w_dff_B_sObn9bEK3_1),.dout(n1011),.clk(gclk));
	jand g0711(.dina(w_G1694_1[0]),.dinb(w_G1691_4[2]),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_4[1]),.dinb(w_G185_0[0]),.dout(n1013),.clk(gclk));
	jand g0713(.dina(w_G1694_0[2]),.dinb(w_n1008_4[1]),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_4[1]),.dinb(w_G182_0[0]),.dout(n1015),.clk(gclk));
	jor g0715(.dina(n1015),.dinb(w_dff_B_Er9MKswT7_1),.dout(n1016),.clk(gclk));
	jor g0716(.dina(w_dff_B_jYwc0CJA9_0),.dinb(n1011),.dout(n1017),.clk(gclk));
	jand g0717(.dina(n1017),.dinb(w_G137_9[0]),.dout(w_dff_A_JOmnUMds0_2),.clk(gclk));
	jnot g0718(.din(w_G871_0),.dout(n1019),.clk(gclk));
	jor g0719(.dina(w_n1019_1[1]),.dinb(w_n797_8[2]),.dout(n1020),.clk(gclk));
	jnot g0720(.din(w_G832_0),.dout(n1021),.clk(gclk));
	jor g0721(.dina(w_n1021_1[1]),.dinb(w_G4088_8[2]),.dout(n1022),.clk(gclk));
	jand g0722(.dina(n1022),.dinb(w_n800_4[0]),.dout(n1023),.clk(gclk));
	jand g0723(.dina(n1023),.dinb(w_dff_B_0j02iMEa7_1),.dout(n1024),.clk(gclk));
	jor g0724(.dina(w_n797_8[1]),.dinb(w_G37_0[1]),.dout(n1025),.clk(gclk));
	jor g0725(.dina(w_G4088_8[1]),.dinb(w_G43_0[1]),.dout(n1026),.clk(gclk));
	jand g0726(.dina(n1026),.dinb(w_G4087_4[0]),.dout(n1027),.clk(gclk));
	jand g0727(.dina(n1027),.dinb(n1025),.dout(n1028),.clk(gclk));
	jor g0728(.dina(w_dff_B_XbfJ5Bvn5_0),.dinb(n1024),.dout(w_dff_A_jqIyVt3z5_2),.clk(gclk));
	jnot g0729(.din(w_G873_0),.dout(n1030),.clk(gclk));
	jor g0730(.dina(w_n1030_1[1]),.dinb(w_n797_8[0]),.dout(n1031),.clk(gclk));
	jnot g0731(.din(w_G834_0),.dout(n1032),.clk(gclk));
	jor g0732(.dina(w_n1032_1[1]),.dinb(w_G4088_8[0]),.dout(n1033),.clk(gclk));
	jand g0733(.dina(n1033),.dinb(w_n800_3[2]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(n1034),.dinb(w_dff_B_Hp4BtsS16_1),.dout(n1035),.clk(gclk));
	jor g0735(.dina(w_n797_7[2]),.dinb(w_G20_0[1]),.dout(n1036),.clk(gclk));
	jor g0736(.dina(w_G4088_7[2]),.dinb(w_G76_0[1]),.dout(n1037),.clk(gclk));
	jand g0737(.dina(n1037),.dinb(w_G4087_3[2]),.dout(n1038),.clk(gclk));
	jand g0738(.dina(n1038),.dinb(n1036),.dout(n1039),.clk(gclk));
	jor g0739(.dina(w_dff_B_MzogfC1j1_0),.dinb(n1035),.dout(w_dff_A_BPQdP7vV4_2),.clk(gclk));
	jnot g0740(.din(w_G836_0),.dout(n1041),.clk(gclk));
	jor g0741(.dina(w_n1041_1[1]),.dinb(w_G4088_7[1]),.dout(n1042),.clk(gclk));
	jnot g0742(.din(w_G875_0),.dout(n1043),.clk(gclk));
	jor g0743(.dina(w_n1043_1[1]),.dinb(w_n797_7[1]),.dout(n1044),.clk(gclk));
	jand g0744(.dina(n1044),.dinb(w_n800_3[1]),.dout(n1045),.clk(gclk));
	jand g0745(.dina(n1045),.dinb(w_dff_B_GSF4OTTx6_1),.dout(n1046),.clk(gclk));
	jor g0746(.dina(w_n797_7[0]),.dinb(w_G17_0[1]),.dout(n1047),.clk(gclk));
	jor g0747(.dina(w_G4088_7[0]),.dinb(w_G73_0[1]),.dout(n1048),.clk(gclk));
	jand g0748(.dina(n1048),.dinb(w_G4087_3[1]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(n1049),.dinb(n1047),.dout(n1050),.clk(gclk));
	jor g0750(.dina(w_dff_B_Yerqif9U3_0),.dinb(n1046),.dout(w_dff_A_D2cceXBm3_2),.clk(gclk));
	jnot g0751(.din(w_G877_0),.dout(n1052),.clk(gclk));
	jor g0752(.dina(w_n1052_1[1]),.dinb(w_n797_6[2]),.dout(n1053),.clk(gclk));
	jnot g0753(.din(w_G838_0),.dout(n1054),.clk(gclk));
	jor g0754(.dina(w_n1054_1[1]),.dinb(w_G4088_6[2]),.dout(n1055),.clk(gclk));
	jand g0755(.dina(n1055),.dinb(w_n800_3[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(n1056),.dinb(w_dff_B_XPkTXUtv3_1),.dout(n1057),.clk(gclk));
	jor g0757(.dina(w_n797_6[1]),.dinb(w_G70_0[1]),.dout(n1058),.clk(gclk));
	jor g0758(.dina(w_G4088_6[1]),.dinb(w_G67_0[1]),.dout(n1059),.clk(gclk));
	jand g0759(.dina(n1059),.dinb(w_G4087_3[0]),.dout(n1060),.clk(gclk));
	jand g0760(.dina(n1060),.dinb(n1058),.dout(n1061),.clk(gclk));
	jor g0761(.dina(w_dff_B_NXlOkNV54_0),.dinb(n1057),.dout(w_dff_A_AEoA2Y3E4_2),.clk(gclk));
	jor g0762(.dina(w_G4089_8[2]),.dinb(w_G43_0[0]),.dout(n1063),.clk(gclk));
	jor g0763(.dina(w_n852_8[2]),.dinb(w_G37_0[0]),.dout(n1064),.clk(gclk));
	jand g0764(.dina(n1064),.dinb(w_G4090_4[0]),.dout(n1065),.clk(gclk));
	jand g0765(.dina(n1065),.dinb(w_dff_B_JwnPyo986_1),.dout(n1066),.clk(gclk));
	jor g0766(.dina(w_n1021_1[0]),.dinb(w_G4089_8[1]),.dout(n1067),.clk(gclk));
	jor g0767(.dina(w_n1019_1[0]),.dinb(w_n852_8[1]),.dout(n1068),.clk(gclk));
	jand g0768(.dina(n1068),.dinb(n1067),.dout(n1069),.clk(gclk));
	jand g0769(.dina(n1069),.dinb(w_n854_4[0]),.dout(n1070),.clk(gclk));
	jor g0770(.dina(n1070),.dinb(w_dff_B_IZm3Gvzd0_1),.dout(w_dff_A_0GA9B52D4_2),.clk(gclk));
	jor g0771(.dina(w_G4089_8[0]),.dinb(w_G76_0[0]),.dout(n1072),.clk(gclk));
	jor g0772(.dina(w_n852_8[0]),.dinb(w_G20_0[0]),.dout(n1073),.clk(gclk));
	jand g0773(.dina(n1073),.dinb(w_G4090_3[2]),.dout(n1074),.clk(gclk));
	jand g0774(.dina(n1074),.dinb(w_dff_B_z2wmbyYC3_1),.dout(n1075),.clk(gclk));
	jor g0775(.dina(w_n1032_1[0]),.dinb(w_G4089_7[2]),.dout(n1076),.clk(gclk));
	jor g0776(.dina(w_n1030_1[0]),.dinb(w_n852_7[2]),.dout(n1077),.clk(gclk));
	jand g0777(.dina(w_dff_B_OTTsIfBA1_0),.dinb(n1076),.dout(n1078),.clk(gclk));
	jand g0778(.dina(n1078),.dinb(w_n854_3[2]),.dout(n1079),.clk(gclk));
	jor g0779(.dina(n1079),.dinb(w_dff_B_3PqhCcif5_1),.dout(w_dff_A_PIbZeKxV2_2),.clk(gclk));
	jor g0780(.dina(w_G4089_7[1]),.dinb(w_G73_0[0]),.dout(n1081),.clk(gclk));
	jor g0781(.dina(w_n852_7[1]),.dinb(w_G17_0[0]),.dout(n1082),.clk(gclk));
	jand g0782(.dina(n1082),.dinb(w_G4090_3[1]),.dout(n1083),.clk(gclk));
	jand g0783(.dina(n1083),.dinb(w_dff_B_f9HXrqET1_1),.dout(n1084),.clk(gclk));
	jor g0784(.dina(w_n1043_1[0]),.dinb(w_n852_7[0]),.dout(n1085),.clk(gclk));
	jor g0785(.dina(w_n1041_1[0]),.dinb(w_G4089_7[0]),.dout(n1086),.clk(gclk));
	jand g0786(.dina(n1086),.dinb(n1085),.dout(n1087),.clk(gclk));
	jand g0787(.dina(n1087),.dinb(w_n854_3[1]),.dout(n1088),.clk(gclk));
	jor g0788(.dina(n1088),.dinb(w_dff_B_CMFnyfac9_1),.dout(w_dff_A_ARx0zPuV9_2),.clk(gclk));
	jor g0789(.dina(w_n1052_1[0]),.dinb(w_n852_6[2]),.dout(n1090),.clk(gclk));
	jor g0790(.dina(w_n1054_1[0]),.dinb(w_G4089_6[2]),.dout(n1091),.clk(gclk));
	jand g0791(.dina(n1091),.dinb(w_n854_3[0]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(n1092),.dinb(w_dff_B_e1PvzZF09_1),.dout(n1093),.clk(gclk));
	jor g0793(.dina(w_n852_6[1]),.dinb(w_G70_0[0]),.dout(n1094),.clk(gclk));
	jor g0794(.dina(w_G4089_6[1]),.dinb(w_G67_0[0]),.dout(n1095),.clk(gclk));
	jand g0795(.dina(n1095),.dinb(w_G4090_3[0]),.dout(n1096),.clk(gclk));
	jand g0796(.dina(n1096),.dinb(n1094),.dout(n1097),.clk(gclk));
	jor g0797(.dina(w_dff_B_LKSFC2wQ7_0),.dinb(n1093),.dout(w_dff_A_ViDIITJZ5_2),.clk(gclk));
	jor g0798(.dina(w_n1021_0[2]),.dinb(w_G1689_4[1]),.dout(n1099),.clk(gclk));
	jor g0799(.dina(w_n1019_0[2]),.dinb(w_n993_4[0]),.dout(n1100),.clk(gclk));
	jand g0800(.dina(n1100),.dinb(w_n999_3[1]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(n1101),.dinb(w_dff_B_JeJ532NP3_1),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n994_4[0]),.dinb(w_G200_0[1]),.dout(n1103),.clk(gclk));
	jand g0803(.dina(w_n996_4[0]),.dinb(w_G170_0[1]),.dout(n1104),.clk(gclk));
	jor g0804(.dina(w_dff_B_BcTWHefg0_0),.dinb(n1103),.dout(n1105),.clk(gclk));
	jor g0805(.dina(w_dff_B_URYxDwxI2_0),.dinb(n1102),.dout(n1106),.clk(gclk));
	jand g0806(.dina(n1106),.dinb(w_G137_8[2]),.dout(w_dff_A_WJMGnPZm5_2),.clk(gclk));
	jor g0807(.dina(w_n1054_0[2]),.dinb(w_G1689_4[0]),.dout(n1108),.clk(gclk));
	jor g0808(.dina(w_n1052_0[2]),.dinb(w_n993_3[2]),.dout(n1109),.clk(gclk));
	jand g0809(.dina(n1109),.dinb(w_n999_3[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(w_dff_B_YAFkuvKh2_0),.dinb(n1108),.dout(n1111),.clk(gclk));
	jand g0811(.dina(w_n994_3[2]),.dinb(w_G188_0[1]),.dout(n1112),.clk(gclk));
	jand g0812(.dina(w_n996_3[2]),.dinb(w_G158_0[1]),.dout(n1113),.clk(gclk));
	jor g0813(.dina(w_dff_B_ZTwiHh5O9_0),.dinb(n1112),.dout(n1114),.clk(gclk));
	jor g0814(.dina(w_dff_B_VxYJZoC49_0),.dinb(n1111),.dout(n1115),.clk(gclk));
	jand g0815(.dina(n1115),.dinb(w_G137_8[1]),.dout(w_dff_A_3gh9jhrR8_2),.clk(gclk));
	jor g0816(.dina(w_n1041_0[2]),.dinb(w_G1689_3[2]),.dout(n1117),.clk(gclk));
	jor g0817(.dina(w_n1043_0[2]),.dinb(w_n993_3[1]),.dout(n1118),.clk(gclk));
	jand g0818(.dina(n1118),.dinb(w_n999_2[2]),.dout(n1119),.clk(gclk));
	jand g0819(.dina(n1119),.dinb(w_dff_B_3QEbJYIQ0_1),.dout(n1120),.clk(gclk));
	jand g0820(.dina(w_n994_3[1]),.dinb(w_G155_0[1]),.dout(n1121),.clk(gclk));
	jand g0821(.dina(w_n996_3[1]),.dinb(w_G152_0[1]),.dout(n1122),.clk(gclk));
	jor g0822(.dina(w_dff_B_qeCi42wT9_0),.dinb(n1121),.dout(n1123),.clk(gclk));
	jor g0823(.dina(w_dff_B_93Pkxbgz0_0),.dinb(n1120),.dout(n1124),.clk(gclk));
	jand g0824(.dina(n1124),.dinb(w_G137_8[0]),.dout(w_dff_A_JYKdF5A27_2),.clk(gclk));
	jor g0825(.dina(w_n1032_0[2]),.dinb(w_G1689_3[1]),.dout(n1126),.clk(gclk));
	jor g0826(.dina(w_n1030_0[2]),.dinb(w_n993_3[0]),.dout(n1127),.clk(gclk));
	jand g0827(.dina(n1127),.dinb(w_n999_2[1]),.dout(n1128),.clk(gclk));
	jand g0828(.dina(n1128),.dinb(n1126),.dout(n1129),.clk(gclk));
	jand g0829(.dina(w_n994_3[0]),.dinb(w_G149_0[1]),.dout(n1130),.clk(gclk));
	jand g0830(.dina(w_n996_3[0]),.dinb(w_G146_0[1]),.dout(n1131),.clk(gclk));
	jor g0831(.dina(w_dff_B_P8C265hN7_0),.dinb(n1130),.dout(n1132),.clk(gclk));
	jor g0832(.dina(w_dff_B_Zp7KqYat4_0),.dinb(n1129),.dout(n1133),.clk(gclk));
	jand g0833(.dina(n1133),.dinb(w_G137_7[2]),.dout(w_dff_A_N23fx6Y26_2),.clk(gclk));
	jand g0834(.dina(w_n1014_4[0]),.dinb(w_G200_0[0]),.dout(n1135),.clk(gclk));
	jand g0835(.dina(w_n1012_4[0]),.dinb(w_G170_0[0]),.dout(n1136),.clk(gclk));
	jor g0836(.dina(w_n1019_0[1]),.dinb(w_n1008_4[0]),.dout(n1137),.clk(gclk));
	jor g0837(.dina(w_n1021_0[1]),.dinb(w_G1691_4[1]),.dout(n1138),.clk(gclk));
	jand g0838(.dina(n1138),.dinb(n1137),.dout(n1139),.clk(gclk));
	jand g0839(.dina(n1139),.dinb(w_n1007_3[1]),.dout(n1140),.clk(gclk));
	jor g0840(.dina(n1140),.dinb(w_dff_B_b0B1pIhC7_1),.dout(n1141),.clk(gclk));
	jor g0841(.dina(n1141),.dinb(w_dff_B_YPte2gEs3_1),.dout(n1142),.clk(gclk));
	jand g0842(.dina(n1142),.dinb(w_G137_7[1]),.dout(w_dff_A_1W05j3Ma7_2),.clk(gclk));
	jor g0843(.dina(w_n1054_0[1]),.dinb(w_G1691_4[0]),.dout(n1144),.clk(gclk));
	jor g0844(.dina(w_n1052_0[1]),.dinb(w_n1008_3[2]),.dout(n1145),.clk(gclk));
	jand g0845(.dina(n1145),.dinb(w_n1007_3[0]),.dout(n1146),.clk(gclk));
	jand g0846(.dina(w_dff_B_WevrzoMI7_0),.dinb(n1144),.dout(n1147),.clk(gclk));
	jand g0847(.dina(w_n1014_3[2]),.dinb(w_G188_0[0]),.dout(n1148),.clk(gclk));
	jand g0848(.dina(w_n1012_3[2]),.dinb(w_G158_0[0]),.dout(n1149),.clk(gclk));
	jor g0849(.dina(w_dff_B_KoFZQHj32_0),.dinb(n1148),.dout(n1150),.clk(gclk));
	jor g0850(.dina(w_dff_B_0mHdEneZ3_0),.dinb(n1147),.dout(n1151),.clk(gclk));
	jand g0851(.dina(n1151),.dinb(w_G137_7[0]),.dout(w_dff_A_vTDZFZYD2_2),.clk(gclk));
	jor g0852(.dina(w_n1041_0[1]),.dinb(w_G1691_3[2]),.dout(n1153),.clk(gclk));
	jor g0853(.dina(w_n1043_0[1]),.dinb(w_n1008_3[1]),.dout(n1154),.clk(gclk));
	jand g0854(.dina(n1154),.dinb(w_n1007_2[2]),.dout(n1155),.clk(gclk));
	jand g0855(.dina(n1155),.dinb(w_dff_B_SMMNfKzr1_1),.dout(n1156),.clk(gclk));
	jand g0856(.dina(w_n1014_3[1]),.dinb(w_G155_0[0]),.dout(n1157),.clk(gclk));
	jand g0857(.dina(w_n1012_3[1]),.dinb(w_G152_0[0]),.dout(n1158),.clk(gclk));
	jor g0858(.dina(w_dff_B_hrPZbIHP1_0),.dinb(n1157),.dout(n1159),.clk(gclk));
	jor g0859(.dina(w_dff_B_2iqz4Qca6_0),.dinb(n1156),.dout(n1160),.clk(gclk));
	jand g0860(.dina(n1160),.dinb(w_G137_6[2]),.dout(w_dff_A_AjepxUwp4_2),.clk(gclk));
	jor g0861(.dina(w_n1032_0[1]),.dinb(w_G1691_3[1]),.dout(n1162),.clk(gclk));
	jor g0862(.dina(w_n1030_0[1]),.dinb(w_n1008_3[0]),.dout(n1163),.clk(gclk));
	jand g0863(.dina(n1163),.dinb(w_n1007_2[1]),.dout(n1164),.clk(gclk));
	jand g0864(.dina(n1164),.dinb(n1162),.dout(n1165),.clk(gclk));
	jand g0865(.dina(w_n1014_3[0]),.dinb(w_G149_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n1012_3[0]),.dinb(w_G146_0[0]),.dout(n1167),.clk(gclk));
	jor g0867(.dina(w_dff_B_zBKxwZd23_0),.dinb(n1166),.dout(n1168),.clk(gclk));
	jor g0868(.dina(w_dff_B_yHemKvBF0_0),.dinb(n1165),.dout(n1169),.clk(gclk));
	jand g0869(.dina(n1169),.dinb(w_G137_6[1]),.dout(w_dff_A_YYfSZWDj9_2),.clk(gclk));
	jnot g0870(.din(G135),.dout(n1171),.clk(gclk));
	jnot g0871(.din(G4115),.dout(n1172),.clk(gclk));
	jor g0872(.dina(n1172),.dinb(n1171),.dout(n1173),.clk(gclk));
	jnot g0873(.din(w_n428_1[0]),.dout(n1174),.clk(gclk));
	jor g0874(.dina(n1174),.dinb(w_G3724_0[2]),.dout(n1175),.clk(gclk));
	jnot g0875(.din(w_G3717_0[1]),.dout(n1176),.clk(gclk));
	jnot g0876(.din(w_G3724_0[1]),.dout(n1177),.clk(gclk));
	jxor g0877(.dina(w_n790_0[0]),.dinb(w_dff_B_K8TahF035_1),.dout(n1178),.clk(gclk));
	jnot g0878(.din(n1178),.dout(n1179),.clk(gclk));
	jor g0879(.dina(w_n1179_0[1]),.dinb(w_n1177_0[1]),.dout(n1180),.clk(gclk));
	jand g0880(.dina(n1180),.dinb(w_dff_B_oO0itrCv6_1),.dout(n1181),.clk(gclk));
	jand g0881(.dina(n1181),.dinb(w_dff_B_twTMpFZ06_1),.dout(n1182),.clk(gclk));
	jor g0882(.dina(w_n795_1[0]),.dinb(w_n1177_0[0]),.dout(n1183),.clk(gclk));
	jor g0883(.dina(w_G3724_0[0]),.dinb(w_G123_0[1]),.dout(n1184),.clk(gclk));
	jand g0884(.dina(n1184),.dinb(w_G3717_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(w_dff_B_2fXFua545_0),.dinb(n1183),.dout(n1186),.clk(gclk));
	jor g0886(.dina(n1186),.dinb(w_dff_B_Pzz3Wyd36_1),.dout(n1187),.clk(gclk));
	jand g0887(.dina(n1187),.dinb(w_dff_B_Ivd7VMH57_1),.dout(w_dff_A_NtujIeyr1_2),.clk(gclk));
	jxor g0888(.dina(w_n1179_0[0]),.dinb(w_n795_0[2]),.dout(w_dff_A_bLgQBZ9M2_2),.clk(gclk));
	jand g0889(.dina(w_n750_5[1]),.dinb(w_G123_0[0]),.dout(n1190),.clk(gclk));
	jor g0890(.dina(w_n795_0[1]),.dinb(w_n749_9[2]),.dout(n1191),.clk(gclk));
	jand g0891(.dina(w_n428_0[2]),.dinb(w_n749_9[1]),.dout(n1192),.clk(gclk));
	jor g0892(.dina(n1192),.dinb(w_G4092_6[0]),.dout(n1193),.clk(gclk));
	jnot g0893(.din(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_dff_B_0MzYLJRa4_0),.dinb(n1191),.dout(n1195),.clk(gclk));
	jor g0895(.dina(n1195),.dinb(w_dff_B_AMKwCWI48_1),.dout(n1196),.clk(gclk));
	jnot g0896(.din(w_n1196_1[2]),.dout(w_dff_A_IwSzkPSy1_1),.clk(gclk));
	jand g0897(.dina(w_n750_5[0]),.dinb(w_dff_B_znfhQR8X5_1),.dout(n1198),.clk(gclk));
	jand g0898(.dina(w_n433_0[1]),.dinb(w_n749_9[0]),.dout(n1199),.clk(gclk));
	jnot g0899(.din(n1199),.dout(n1200),.clk(gclk));
	jnot g0900(.din(w_G4092_5[2]),.dout(n1201),.clk(gclk));
	jor g0901(.dina(w_n969_0[0]),.dinb(w_n749_8[2]),.dout(n1202),.clk(gclk));
	jand g0902(.dina(n1202),.dinb(w_n1201_0[2]),.dout(n1203),.clk(gclk));
	jand g0903(.dina(n1203),.dinb(w_dff_B_n8YfteQh9_1),.dout(n1204),.clk(gclk));
	jor g0904(.dina(n1204),.dinb(w_dff_B_JnMTqY8m2_1),.dout(n1205),.clk(gclk));
	jnot g0905(.din(w_n1205_1[2]),.dout(w_dff_A_LBerTre86_1),.clk(gclk));
	jand g0906(.dina(w_n750_4[2]),.dinb(w_dff_B_QvouAMqL3_1),.dout(n1207),.clk(gclk));
	jor g0907(.dina(w_n986_0[0]),.dinb(w_n749_8[1]),.dout(n1208),.clk(gclk));
	jand g0908(.dina(w_n423_0[1]),.dinb(w_n749_8[0]),.dout(n1209),.clk(gclk));
	jor g0909(.dina(n1209),.dinb(w_G4092_5[1]),.dout(n1210),.clk(gclk));
	jnot g0910(.din(n1210),.dout(n1211),.clk(gclk));
	jand g0911(.dina(w_dff_B_UTvvvdCC3_0),.dinb(n1208),.dout(n1212),.clk(gclk));
	jor g0912(.dina(n1212),.dinb(w_dff_B_35MiG9rW5_1),.dout(n1213),.clk(gclk));
	jnot g0913(.din(w_n1213_1[2]),.dout(w_dff_A_2FsCfOkF2_1),.clk(gclk));
	jand g0914(.dina(w_n750_4[1]),.dinb(w_dff_B_a73Lzl8l8_1),.dout(n1215),.clk(gclk));
	jnot g0915(.din(n1215),.dout(n1216),.clk(gclk));
	jand g0916(.dina(w_n989_0[0]),.dinb(w_G4091_2[2]),.dout(n1217),.clk(gclk));
	jand g0917(.dina(w_n412_0[1]),.dinb(w_n749_7[2]),.dout(n1218),.clk(gclk));
	jor g0918(.dina(n1218),.dinb(w_G4092_5[0]),.dout(n1219),.clk(gclk));
	jor g0919(.dina(w_dff_B_gq1cU9fC3_0),.dinb(n1217),.dout(n1220),.clk(gclk));
	jand g0920(.dina(n1220),.dinb(w_dff_B_AJAIRTUo0_1),.dout(G830_fa_),.clk(gclk));
	jand g0921(.dina(w_n680_0[0]),.dinb(w_G245_0[0]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(w_dff_B_2ri51vPv3_0),.dinb(w_n935_0[0]),.dout(n1223),.clk(gclk));
	jnot g0923(.din(w_G998_0),.dout(n1224),.clk(gclk));
	jand g0924(.dina(w_n318_0[0]),.dinb(w_G601_0),.dout(n1225),.clk(gclk));
	jand g0925(.dina(n1225),.dinb(w_G559_0[0]),.dout(n1226),.clk(gclk));
	jand g0926(.dina(w_dff_B_eh53O0zL0_0),.dinb(w_n670_0[0]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_dff_B_xC81aw5z5_0),.dinb(n1224),.dout(n1228),.clk(gclk));
	jand g0928(.dina(n1228),.dinb(w_dff_B_btmOODy13_1),.dout(w_dff_A_GCA5ODBX8_2),.clk(gclk));
	jand g0929(.dina(w_n750_4[0]),.dinb(w_dff_B_OUybV2HC1_1),.dout(n1230),.clk(gclk));
	jand g0930(.dina(w_n551_0[1]),.dinb(w_n749_7[1]),.dout(n1231),.clk(gclk));
	jnot g0931(.din(n1231),.dout(n1232),.clk(gclk));
	jor g0932(.dina(w_n944_0[0]),.dinb(w_n749_7[0]),.dout(n1233),.clk(gclk));
	jand g0933(.dina(n1233),.dinb(w_n1201_0[1]),.dout(n1234),.clk(gclk));
	jand g0934(.dina(n1234),.dinb(w_dff_B_GtU33t4T5_1),.dout(n1235),.clk(gclk));
	jor g0935(.dina(n1235),.dinb(w_dff_B_xBbinTII5_1),.dout(n1236),.clk(gclk));
	jnot g0936(.din(w_n1236_1[2]),.dout(w_dff_A_17s6VL7c5_1),.clk(gclk));
	jand g0937(.dina(w_n750_3[2]),.dinb(w_dff_B_vTfpB1Oo6_1),.dout(n1238),.clk(gclk));
	jnot g0938(.din(n1238),.dout(n1239),.clk(gclk));
	jand g0939(.dina(w_n949_0[0]),.dinb(w_G4091_2[1]),.dout(n1240),.clk(gclk));
	jand g0940(.dina(w_n459_0[0]),.dinb(w_n749_6[2]),.dout(n1241),.clk(gclk));
	jor g0941(.dina(n1241),.dinb(w_G4092_4[2]),.dout(n1242),.clk(gclk));
	jor g0942(.dina(w_dff_B_QRj5i3yC5_0),.dinb(n1240),.dout(n1243),.clk(gclk));
	jand g0943(.dina(n1243),.dinb(w_dff_B_6vS3LmRH4_1),.dout(G865_fa_),.clk(gclk));
	jand g0944(.dina(w_n750_3[1]),.dinb(w_dff_B_4Ds4lwDP6_1),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n517_0[0]),.dinb(w_n749_6[1]),.dout(n1246),.clk(gclk));
	jnot g0946(.din(n1246),.dout(n1247),.clk(gclk));
	jor g0947(.dina(w_n957_0[0]),.dinb(w_n749_6[0]),.dout(n1248),.clk(gclk));
	jand g0948(.dina(n1248),.dinb(w_n1201_0[0]),.dout(n1249),.clk(gclk));
	jand g0949(.dina(n1249),.dinb(w_dff_B_SpJwA4xT9_1),.dout(n1250),.clk(gclk));
	jor g0950(.dina(n1250),.dinb(w_dff_B_3gr4XNVP0_1),.dout(n1251),.clk(gclk));
	jnot g0951(.din(w_n1251_1[2]),.dout(w_dff_A_RDGMn0975_1),.clk(gclk));
	jand g0952(.dina(w_n750_3[0]),.dinb(w_dff_B_Z0yc7H8z2_1),.dout(n1253),.clk(gclk));
	jnot g0953(.din(n1253),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n964_0[0]),.dinb(w_G4091_2[0]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n504_0[0]),.dinb(w_n749_5[2]),.dout(n1256),.clk(gclk));
	jor g0956(.dina(n1256),.dinb(w_G4092_4[1]),.dout(n1257),.clk(gclk));
	jor g0957(.dina(w_dff_B_hcrYth2O5_0),.dinb(n1255),.dout(n1258),.clk(gclk));
	jand g0958(.dina(n1258),.dinb(w_dff_B_WgBFhtdP5_1),.dout(G869_fa_),.clk(gclk));
	jor g0959(.dina(w_G4089_6[0]),.dinb(w_G109_0[1]),.dout(n1260),.clk(gclk));
	jor g0960(.dina(w_n852_6[0]),.dinb(w_G106_0[1]),.dout(n1261),.clk(gclk));
	jand g0961(.dina(n1261),.dinb(w_G4090_2[2]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(n1262),.dinb(w_dff_B_EllftlNr1_1),.dout(n1263),.clk(gclk));
	jor g0963(.dina(w_n1236_1[1]),.dinb(w_n852_5[2]),.dout(n1264),.clk(gclk));
	jor g0964(.dina(w_n1196_1[1]),.dinb(w_G4089_5[2]),.dout(n1265),.clk(gclk));
	jand g0965(.dina(n1265),.dinb(w_n854_2[2]),.dout(n1266),.clk(gclk));
	jand g0966(.dina(n1266),.dinb(n1264),.dout(n1267),.clk(gclk));
	jor g0967(.dina(n1267),.dinb(w_dff_B_Oa4FPMrk7_1),.dout(w_dff_A_e2RZ5Gl43_2),.clk(gclk));
	jor g0968(.dina(w_n1196_1[0]),.dinb(w_G4088_6[0]),.dout(n1269),.clk(gclk));
	jor g0969(.dina(w_n1236_1[0]),.dinb(w_n797_6[0]),.dout(n1270),.clk(gclk));
	jand g0970(.dina(n1270),.dinb(w_n800_2[2]),.dout(n1271),.clk(gclk));
	jand g0971(.dina(n1271),.dinb(w_dff_B_5kW2X1Jt1_1),.dout(n1272),.clk(gclk));
	jor g0972(.dina(w_n797_5[2]),.dinb(w_G106_0[0]),.dout(n1273),.clk(gclk));
	jor g0973(.dina(w_G4088_5[2]),.dinb(w_G109_0[0]),.dout(n1274),.clk(gclk));
	jand g0974(.dina(n1274),.dinb(w_G4087_2[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(n1275),.dinb(n1273),.dout(n1276),.clk(gclk));
	jor g0976(.dina(w_dff_B_Oc5FpvzU5_0),.dinb(n1272),.dout(w_dff_A_FqM4NOCB0_2),.clk(gclk));
	jor g0977(.dina(w_n1205_1[1]),.dinb(w_G4088_5[1]),.dout(n1278),.clk(gclk));
	jnot g0978(.din(w_G865_0),.dout(n1279),.clk(gclk));
	jor g0979(.dina(w_n1279_1[1]),.dinb(w_n797_5[1]),.dout(n1280),.clk(gclk));
	jand g0980(.dina(n1280),.dinb(w_n800_2[1]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(n1281),.dinb(w_dff_B_gocFImUT3_1),.dout(n1282),.clk(gclk));
	jor g0982(.dina(w_n797_5[0]),.dinb(w_G49_0[1]),.dout(n1283),.clk(gclk));
	jor g0983(.dina(w_G4088_5[0]),.dinb(w_G46_0[1]),.dout(n1284),.clk(gclk));
	jand g0984(.dina(n1284),.dinb(w_G4087_2[1]),.dout(n1285),.clk(gclk));
	jand g0985(.dina(n1285),.dinb(n1283),.dout(n1286),.clk(gclk));
	jor g0986(.dina(w_dff_B_ucBX0RAq0_0),.dinb(n1282),.dout(w_dff_A_lz8TOsR45_2),.clk(gclk));
	jor g0987(.dina(w_n1213_1[1]),.dinb(w_G4088_4[2]),.dout(n1288),.clk(gclk));
	jor g0988(.dina(w_n1251_1[1]),.dinb(w_n797_4[2]),.dout(n1289),.clk(gclk));
	jand g0989(.dina(n1289),.dinb(w_n800_2[0]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(n1290),.dinb(w_dff_B_0D6r4phK0_1),.dout(n1291),.clk(gclk));
	jor g0991(.dina(w_n797_4[1]),.dinb(w_G103_0[1]),.dout(n1292),.clk(gclk));
	jor g0992(.dina(w_G4088_4[1]),.dinb(w_G100_0[1]),.dout(n1293),.clk(gclk));
	jand g0993(.dina(n1293),.dinb(w_G4087_2[0]),.dout(n1294),.clk(gclk));
	jand g0994(.dina(n1294),.dinb(n1292),.dout(n1295),.clk(gclk));
	jor g0995(.dina(w_dff_B_ckn15Wxm8_0),.dinb(n1291),.dout(w_dff_A_WIFa6DUd8_2),.clk(gclk));
	jnot g0996(.din(w_G830_0),.dout(n1297),.clk(gclk));
	jor g0997(.dina(w_n1297_1[1]),.dinb(w_G4088_4[0]),.dout(n1298),.clk(gclk));
	jnot g0998(.din(w_G869_0),.dout(n1299),.clk(gclk));
	jor g0999(.dina(w_n1299_1[1]),.dinb(w_n797_4[0]),.dout(n1300),.clk(gclk));
	jand g1000(.dina(n1300),.dinb(w_n800_1[2]),.dout(n1301),.clk(gclk));
	jand g1001(.dina(n1301),.dinb(w_dff_B_Y0iBS1MF6_1),.dout(n1302),.clk(gclk));
	jor g1002(.dina(w_n797_3[2]),.dinb(w_G40_0[1]),.dout(n1303),.clk(gclk));
	jor g1003(.dina(w_G4088_3[2]),.dinb(w_G91_0[1]),.dout(n1304),.clk(gclk));
	jand g1004(.dina(n1304),.dinb(w_G4087_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(n1305),.dinb(n1303),.dout(n1306),.clk(gclk));
	jor g1006(.dina(w_dff_B_ZPD2HFVt2_0),.dinb(n1302),.dout(w_dff_A_qzcfvnFP9_2),.clk(gclk));
	jor g1007(.dina(w_n1205_1[0]),.dinb(w_G4089_5[1]),.dout(n1308),.clk(gclk));
	jor g1008(.dina(w_n1279_1[0]),.dinb(w_n852_5[1]),.dout(n1309),.clk(gclk));
	jand g1009(.dina(n1309),.dinb(w_n854_2[1]),.dout(n1310),.clk(gclk));
	jand g1010(.dina(n1310),.dinb(w_dff_B_Xq6EIfTl7_1),.dout(n1311),.clk(gclk));
	jor g1011(.dina(w_n852_5[0]),.dinb(w_G49_0[0]),.dout(n1312),.clk(gclk));
	jor g1012(.dina(w_G4089_5[0]),.dinb(w_G46_0[0]),.dout(n1313),.clk(gclk));
	jand g1013(.dina(n1313),.dinb(w_G4090_2[1]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(n1314),.dinb(n1312),.dout(n1315),.clk(gclk));
	jor g1015(.dina(w_dff_B_sS6HhTvr8_0),.dinb(n1311),.dout(w_dff_A_OWe3VifZ2_2),.clk(gclk));
	jor g1016(.dina(w_n1213_1[0]),.dinb(w_G4089_4[2]),.dout(n1317),.clk(gclk));
	jor g1017(.dina(w_n1251_1[0]),.dinb(w_n852_4[2]),.dout(n1318),.clk(gclk));
	jand g1018(.dina(n1318),.dinb(w_n854_2[0]),.dout(n1319),.clk(gclk));
	jand g1019(.dina(n1319),.dinb(w_dff_B_VwyDH8wE1_1),.dout(n1320),.clk(gclk));
	jor g1020(.dina(w_n852_4[1]),.dinb(w_G103_0[0]),.dout(n1321),.clk(gclk));
	jor g1021(.dina(w_G4089_4[1]),.dinb(w_G100_0[0]),.dout(n1322),.clk(gclk));
	jand g1022(.dina(n1322),.dinb(w_G4090_2[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(n1323),.dinb(n1321),.dout(n1324),.clk(gclk));
	jor g1024(.dina(w_dff_B_KRwNmUJd6_0),.dinb(n1320),.dout(w_dff_A_SnzgluzA6_2),.clk(gclk));
	jor g1025(.dina(w_n1297_1[0]),.dinb(w_G4089_4[0]),.dout(n1326),.clk(gclk));
	jor g1026(.dina(w_n1299_1[0]),.dinb(w_n852_4[0]),.dout(n1327),.clk(gclk));
	jand g1027(.dina(n1327),.dinb(w_n854_1[2]),.dout(n1328),.clk(gclk));
	jand g1028(.dina(n1328),.dinb(w_dff_B_ZdDAzTRd3_1),.dout(n1329),.clk(gclk));
	jor g1029(.dina(w_n852_3[2]),.dinb(w_G40_0[0]),.dout(n1330),.clk(gclk));
	jor g1030(.dina(w_G4089_3[2]),.dinb(w_G91_0[0]),.dout(n1331),.clk(gclk));
	jand g1031(.dina(n1331),.dinb(w_G4090_1[2]),.dout(n1332),.clk(gclk));
	jand g1032(.dina(n1332),.dinb(n1330),.dout(n1333),.clk(gclk));
	jor g1033(.dina(w_dff_B_ZMLXcoSU6_0),.dinb(n1329),.dout(w_dff_A_xWOXwuxG9_2),.clk(gclk));
	jor g1034(.dina(w_n1297_0[2]),.dinb(w_G1689_3[0]),.dout(n1335),.clk(gclk));
	jor g1035(.dina(w_n1299_0[2]),.dinb(w_n993_2[2]),.dout(n1336),.clk(gclk));
	jand g1036(.dina(n1336),.dinb(w_n999_2[0]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(n1337),.dinb(w_dff_B_iodepxmR8_1),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n994_2[2]),.dinb(w_G203_0[1]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n996_2[2]),.dinb(w_G173_0[1]),.dout(n1340),.clk(gclk));
	jor g1040(.dina(w_dff_B_ZwbUsRCP6_0),.dinb(n1339),.dout(n1341),.clk(gclk));
	jor g1041(.dina(w_dff_B_eVq55WOs0_0),.dinb(n1338),.dout(n1342),.clk(gclk));
	jand g1042(.dina(n1342),.dinb(w_G137_6[0]),.dout(w_dff_A_XEra2e6U0_2),.clk(gclk));
	jor g1043(.dina(w_n1251_0[2]),.dinb(w_n993_2[1]),.dout(n1344),.clk(gclk));
	jor g1044(.dina(w_n1213_0[2]),.dinb(w_G1689_2[2]),.dout(n1345),.clk(gclk));
	jand g1045(.dina(n1345),.dinb(w_n999_1[2]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(n1346),.dinb(w_dff_B_pXPjkzqj2_1),.dout(n1347),.clk(gclk));
	jand g1047(.dina(w_n994_2[1]),.dinb(w_G197_0[1]),.dout(n1348),.clk(gclk));
	jand g1048(.dina(w_n996_2[1]),.dinb(w_G167_0[1]),.dout(n1349),.clk(gclk));
	jor g1049(.dina(w_dff_B_A9RfTUUr4_0),.dinb(n1348),.dout(n1350),.clk(gclk));
	jor g1050(.dina(w_dff_B_MSnu5F2k2_0),.dinb(n1347),.dout(n1351),.clk(gclk));
	jand g1051(.dina(n1351),.dinb(w_G137_5[2]),.dout(w_dff_A_nhdDMIc41_2),.clk(gclk));
	jand g1052(.dina(w_n994_2[0]),.dinb(w_G194_0[1]),.dout(n1353),.clk(gclk));
	jand g1053(.dina(w_n996_2[0]),.dinb(w_G164_0[1]),.dout(n1354),.clk(gclk));
	jor g1054(.dina(w_dff_B_CWFOGWVM9_0),.dinb(n1353),.dout(n1355),.clk(gclk));
	jor g1055(.dina(w_n1205_0[2]),.dinb(w_G1689_2[1]),.dout(n1356),.clk(gclk));
	jor g1056(.dina(w_n1279_0[2]),.dinb(w_n993_2[0]),.dout(n1357),.clk(gclk));
	jand g1057(.dina(n1357),.dinb(w_dff_B_dzStsXEr1_1),.dout(n1358),.clk(gclk));
	jand g1058(.dina(n1358),.dinb(w_n999_1[1]),.dout(n1359),.clk(gclk));
	jor g1059(.dina(n1359),.dinb(w_dff_B_KUFA6Oyb8_1),.dout(n1360),.clk(gclk));
	jand g1060(.dina(n1360),.dinb(w_G137_5[1]),.dout(w_dff_A_8corv2mp0_2),.clk(gclk));
	jand g1061(.dina(w_n994_1[2]),.dinb(w_G191_0[1]),.dout(n1362),.clk(gclk));
	jand g1062(.dina(w_n996_1[2]),.dinb(w_G161_0[1]),.dout(n1363),.clk(gclk));
	jor g1063(.dina(w_dff_B_1G6woDmf7_0),.dinb(n1362),.dout(n1364),.clk(gclk));
	jor g1064(.dina(w_n1196_0[2]),.dinb(w_G1689_2[0]),.dout(n1365),.clk(gclk));
	jor g1065(.dina(w_n1236_0[2]),.dinb(w_n993_1[2]),.dout(n1366),.clk(gclk));
	jand g1066(.dina(n1366),.dinb(w_dff_B_7pe10V1S7_1),.dout(n1367),.clk(gclk));
	jand g1067(.dina(n1367),.dinb(w_n999_1[0]),.dout(n1368),.clk(gclk));
	jor g1068(.dina(n1368),.dinb(w_dff_B_uDgQeQAK7_1),.dout(n1369),.clk(gclk));
	jand g1069(.dina(n1369),.dinb(w_G137_5[0]),.dout(w_dff_A_8CLLA1Vs8_2),.clk(gclk));
	jor g1070(.dina(w_n1297_0[1]),.dinb(w_G1691_3[0]),.dout(n1371),.clk(gclk));
	jor g1071(.dina(w_n1299_0[1]),.dinb(w_n1008_2[2]),.dout(n1372),.clk(gclk));
	jand g1072(.dina(n1372),.dinb(w_n1007_2[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(n1373),.dinb(w_dff_B_loIilNij4_1),.dout(n1374),.clk(gclk));
	jand g1074(.dina(w_n1014_2[2]),.dinb(w_G203_0[0]),.dout(n1375),.clk(gclk));
	jand g1075(.dina(w_n1012_2[2]),.dinb(w_G173_0[0]),.dout(n1376),.clk(gclk));
	jor g1076(.dina(w_dff_B_uQVjHuL17_0),.dinb(n1375),.dout(n1377),.clk(gclk));
	jor g1077(.dina(w_dff_B_hE9dgaei3_0),.dinb(n1374),.dout(n1378),.clk(gclk));
	jand g1078(.dina(n1378),.dinb(w_G137_4[2]),.dout(w_dff_A_DYPsKfAw4_2),.clk(gclk));
	jand g1079(.dina(w_n1014_2[1]),.dinb(w_G197_0[0]),.dout(n1380),.clk(gclk));
	jand g1080(.dina(w_n1012_2[1]),.dinb(w_G167_0[0]),.dout(n1381),.clk(gclk));
	jor g1081(.dina(w_dff_B_8OPEYJCD1_0),.dinb(n1380),.dout(n1382),.clk(gclk));
	jor g1082(.dina(w_n1213_0[1]),.dinb(w_G1691_2[2]),.dout(n1383),.clk(gclk));
	jor g1083(.dina(w_n1251_0[1]),.dinb(w_n1008_2[1]),.dout(n1384),.clk(gclk));
	jand g1084(.dina(n1384),.dinb(n1383),.dout(n1385),.clk(gclk));
	jand g1085(.dina(n1385),.dinb(w_n1007_1[2]),.dout(n1386),.clk(gclk));
	jor g1086(.dina(n1386),.dinb(w_dff_B_bzeMK1fT3_1),.dout(n1387),.clk(gclk));
	jand g1087(.dina(n1387),.dinb(w_G137_4[1]),.dout(w_dff_A_atPMyXnW8_2),.clk(gclk));
	jor g1088(.dina(w_n1205_0[1]),.dinb(w_G1691_2[1]),.dout(n1389),.clk(gclk));
	jor g1089(.dina(w_n1279_0[1]),.dinb(w_n1008_2[0]),.dout(n1390),.clk(gclk));
	jand g1090(.dina(n1390),.dinb(w_n1007_1[1]),.dout(n1391),.clk(gclk));
	jand g1091(.dina(n1391),.dinb(w_dff_B_MuWztHRc9_1),.dout(n1392),.clk(gclk));
	jand g1092(.dina(w_n1014_2[0]),.dinb(w_G194_0[0]),.dout(n1393),.clk(gclk));
	jand g1093(.dina(w_n1012_2[0]),.dinb(w_G164_0[0]),.dout(n1394),.clk(gclk));
	jor g1094(.dina(w_dff_B_fv6coIyT0_0),.dinb(n1393),.dout(n1395),.clk(gclk));
	jor g1095(.dina(w_dff_B_c0egVQFZ4_0),.dinb(n1392),.dout(n1396),.clk(gclk));
	jand g1096(.dina(n1396),.dinb(w_G137_4[0]),.dout(w_dff_A_7Un7AyR00_2),.clk(gclk));
	jor g1097(.dina(w_n1236_0[1]),.dinb(w_n1008_1[2]),.dout(n1398),.clk(gclk));
	jor g1098(.dina(w_n1196_0[1]),.dinb(w_G1691_2[0]),.dout(n1399),.clk(gclk));
	jand g1099(.dina(n1399),.dinb(w_n1007_1[0]),.dout(n1400),.clk(gclk));
	jand g1100(.dina(n1400),.dinb(n1398),.dout(n1401),.clk(gclk));
	jand g1101(.dina(w_n1014_1[2]),.dinb(w_G191_0[0]),.dout(n1402),.clk(gclk));
	jand g1102(.dina(w_n1012_1[2]),.dinb(w_G161_0[0]),.dout(n1403),.clk(gclk));
	jor g1103(.dina(w_dff_B_Q00mXVOW6_0),.dinb(n1402),.dout(n1404),.clk(gclk));
	jor g1104(.dina(w_dff_B_pD1sRVPu5_0),.dinb(n1401),.dout(n1405),.clk(gclk));
	jand g1105(.dina(n1405),.dinb(w_G137_3[2]),.dout(w_dff_A_JgJF4PTq7_2),.clk(gclk));
	jand g1106(.dina(w_n746_0[0]),.dinb(w_n648_0[2]),.dout(n1407),.clk(gclk));
	jxor g1107(.dina(w_n977_0[0]),.dinb(w_n654_1[0]),.dout(n1408),.clk(gclk));
	jxor g1108(.dina(n1408),.dinb(w_n644_0[0]),.dout(n1409),.clk(gclk));
	jxor g1109(.dina(w_dff_B_JPQ5n1MR2_0),.dinb(n1407),.dout(n1410),.clk(gclk));
	jor g1110(.dina(w_n1410_0[2]),.dinb(w_n737_0[2]),.dout(n1411),.clk(gclk));
	jnot g1111(.din(w_G2174_0[2]),.dout(n1412),.clk(gclk));
	jnot g1112(.din(w_n719_0[0]),.dout(n1413),.clk(gclk));
	jnot g1113(.din(w_n720_0[0]),.dout(n1414),.clk(gclk));
	jor g1114(.dina(w_n821_0[0]),.dinb(w_dff_B_2IxeBqju2_1),.dout(n1415),.clk(gclk));
	jand g1115(.dina(n1415),.dinb(w_dff_B_qr4C19tO9_1),.dout(n1416),.clk(gclk));
	jxor g1116(.dina(w_n742_0[0]),.dinb(w_n654_0[2]),.dout(n1417),.clk(gclk));
	jxor g1117(.dina(n1417),.dinb(w_n792_0[0]),.dout(n1418),.clk(gclk));
	jnot g1118(.din(w_n660_0[1]),.dout(n1419),.clk(gclk));
	jand g1119(.dina(w_n745_0[0]),.dinb(w_n648_0[1]),.dout(n1420),.clk(gclk));
	jand g1120(.dina(n1420),.dinb(w_dff_B_EPT7mUVs7_1),.dout(n1421),.clk(gclk));
	jxor g1121(.dina(n1421),.dinb(w_dff_B_gjHkMSii5_1),.dout(n1422),.clk(gclk));
	jor g1122(.dina(w_n1422_0[1]),.dinb(w_n1416_0[1]),.dout(n1423),.clk(gclk));
	jand g1123(.dina(n1423),.dinb(w_n1412_0[2]),.dout(n1424),.clk(gclk));
	jand g1124(.dina(n1424),.dinb(w_dff_B_rGgM8vH17_1),.dout(n1425),.clk(gclk));
	jnot g1125(.din(w_n1425_0[1]),.dout(n1426),.clk(gclk));
	jnot g1126(.din(w_n641_1[0]),.dout(n1427),.clk(gclk));
	jand g1127(.dina(w_n1416_0[0]),.dinb(w_dff_B_ZdQHdSHF7_1),.dout(n1428),.clk(gclk));
	jor g1128(.dina(w_n1428_0[1]),.dinb(w_n1422_0[0]),.dout(n1429),.clk(gclk));
	jnot g1129(.din(w_n1429_0[1]),.dout(n1430),.clk(gclk));
	jnot g1130(.din(w_n1410_0[1]),.dout(n1431),.clk(gclk));
	jand g1131(.dina(w_n1428_0[0]),.dinb(n1431),.dout(n1432),.clk(gclk));
	jor g1132(.dina(n1432),.dinb(w_n1412_0[1]),.dout(n1433),.clk(gclk));
	jor g1133(.dina(n1433),.dinb(n1430),.dout(n1434),.clk(gclk));
	jand g1134(.dina(n1434),.dinb(n1426),.dout(n1435),.clk(gclk));
	jor g1135(.dina(w_n728_0[0]),.dinb(w_n637_0[0]),.dout(n1436),.clk(gclk));
	jxor g1136(.dina(w_dff_B_94lpjmqD7_0),.dinb(w_n733_0[1]),.dout(n1437),.clk(gclk));
	jxor g1137(.dina(w_dff_B_68DvjMJx9_0),.dinb(w_n735_0[1]),.dout(n1438),.clk(gclk));
	jor g1138(.dina(n1438),.dinb(w_G2174_0[1]),.dout(n1439),.clk(gclk));
	jor g1139(.dina(w_n735_0[0]),.dinb(w_n640_0[0]),.dout(n1440),.clk(gclk));
	jor g1140(.dina(w_n819_0[0]),.dinb(w_n628_0[0]),.dout(n1441),.clk(gclk));
	jor g1141(.dina(w_n733_0[0]),.dinb(w_n814_0[0]),.dout(n1442),.clk(gclk));
	jor g1142(.dina(n1442),.dinb(w_n639_0[0]),.dout(n1443),.clk(gclk));
	jand g1143(.dina(n1443),.dinb(w_dff_B_GQA8Bv4Z2_1),.dout(n1444),.clk(gclk));
	jxor g1144(.dina(n1444),.dinb(n1440),.dout(n1445),.clk(gclk));
	jor g1145(.dina(n1445),.dinb(w_n1412_0[0]),.dout(n1446),.clk(gclk));
	jand g1146(.dina(n1446),.dinb(w_dff_B_Pwwn9wzk7_1),.dout(n1447),.clk(gclk));
	jxor g1147(.dina(w_n620_0[1]),.dinb(w_n618_0[0]),.dout(n1448),.clk(gclk));
	jxor g1148(.dina(w_n767_0[0]),.dinb(w_n624_0[0]),.dout(n1449),.clk(gclk));
	jxor g1149(.dina(n1449),.dinb(w_dff_B_rQR8s6aN8_1),.dout(n1450),.clk(gclk));
	jxor g1150(.dina(w_dff_B_YUJFSNRH8_0),.dinb(n1447),.dout(n1451),.clk(gclk));
	jnot g1151(.din(w_n1451_0[1]),.dout(n1452),.clk(gclk));
	jand g1152(.dina(w_dff_B_oJvbEFDl0_0),.dinb(n1435),.dout(n1453),.clk(gclk));
	jor g1153(.dina(w_n737_0[1]),.dinb(w_n641_0[2]),.dout(n1454),.clk(gclk));
	jor g1154(.dina(n1454),.dinb(w_n1410_0[0]),.dout(n1455),.clk(gclk));
	jand g1155(.dina(n1455),.dinb(w_G2174_0[0]),.dout(n1456),.clk(gclk));
	jand g1156(.dina(n1456),.dinb(w_n1429_0[0]),.dout(n1457),.clk(gclk));
	jor g1157(.dina(n1457),.dinb(w_n1425_0[0]),.dout(n1458),.clk(gclk));
	jand g1158(.dina(w_n1451_0[0]),.dinb(n1458),.dout(n1459),.clk(gclk));
	jor g1159(.dina(n1459),.dinb(w_n749_5[1]),.dout(n1460),.clk(gclk));
	jor g1160(.dina(n1460),.dinb(w_dff_B_nmS8vhuX1_1),.dout(n1461),.clk(gclk));
	jand g1161(.dina(w_G351_1[0]),.dinb(w_G248_4[1]),.dout(n1462),.clk(gclk));
	jand g1162(.dina(w_n374_0[2]),.dinb(w_G251_4[0]),.dout(n1463),.clk(gclk));
	jor g1163(.dina(n1463),.dinb(w_n377_0[1]),.dout(n1464),.clk(gclk));
	jor g1164(.dina(n1464),.dinb(w_dff_B_eFO82afY2_1),.dout(n1465),.clk(gclk));
	jand g1165(.dina(w_n374_0[1]),.dinb(w_n406_4[0]),.dout(n1466),.clk(gclk));
	jand g1166(.dina(w_G351_0[2]),.dinb(w_n408_4[1]),.dout(n1467),.clk(gclk));
	jor g1167(.dina(n1467),.dinb(n1466),.dout(n1468),.clk(gclk));
	jor g1168(.dina(n1468),.dinb(w_G534_0[2]),.dout(n1469),.clk(gclk));
	jand g1169(.dina(n1469),.dinb(n1465),.dout(n1470),.clk(gclk));
	jand g1170(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1471),.clk(gclk));
	jand g1171(.dina(w_n387_0[2]),.dinb(w_G251_3[2]),.dout(n1472),.clk(gclk));
	jor g1172(.dina(n1472),.dinb(w_n389_0[1]),.dout(n1473),.clk(gclk));
	jor g1173(.dina(n1473),.dinb(w_dff_B_qItMzJlr6_1),.dout(n1474),.clk(gclk));
	jand g1174(.dina(w_n387_0[1]),.dinb(w_n406_3[2]),.dout(n1475),.clk(gclk));
	jand g1175(.dina(w_G341_0[2]),.dinb(w_n408_4[0]),.dout(n1476),.clk(gclk));
	jor g1176(.dina(n1476),.dinb(n1475),.dout(n1477),.clk(gclk));
	jor g1177(.dina(n1477),.dinb(w_G523_0[1]),.dout(n1478),.clk(gclk));
	jand g1178(.dina(n1478),.dinb(n1474),.dout(n1479),.clk(gclk));
	jxor g1179(.dina(n1479),.dinb(n1470),.dout(n1480),.clk(gclk));
	jor g1180(.dina(w_n435_1[0]),.dinb(w_n369_1[0]),.dout(n1481),.clk(gclk));
	jor g1181(.dina(w_G324_0[2]),.dinb(w_n366_1[0]),.dout(n1482),.clk(gclk));
	jand g1182(.dina(n1482),.dinb(w_G503_0[2]),.dout(n1483),.clk(gclk));
	jand g1183(.dina(n1483),.dinb(w_dff_B_KuVIetra4_1),.dout(n1484),.clk(gclk));
	jor g1184(.dina(w_G324_0[1]),.dinb(w_G254_1[0]),.dout(n1485),.clk(gclk));
	jor g1185(.dina(w_n435_0[2]),.dinb(w_G242_1[0]),.dout(n1486),.clk(gclk));
	jand g1186(.dina(n1486),.dinb(w_dff_B_29o6Iq4y3_1),.dout(n1487),.clk(gclk));
	jand g1187(.dina(n1487),.dinb(w_n437_0[0]),.dout(n1488),.clk(gclk));
	jor g1188(.dina(n1488),.dinb(n1484),.dout(n1489),.clk(gclk));
	jor g1189(.dina(w_G514_0[2]),.dinb(w_n408_3[2]),.dout(n1490),.clk(gclk));
	jor g1190(.dina(w_n361_0[0]),.dinb(w_G248_3[2]),.dout(n1491),.clk(gclk));
	jand g1191(.dina(n1491),.dinb(n1490),.dout(n1492),.clk(gclk));
	jxor g1192(.dina(n1492),.dinb(w_n371_0[0]),.dout(n1493),.clk(gclk));
	jxor g1193(.dina(w_dff_B_JZ7huyEY5_0),.dinb(n1489),.dout(n1494),.clk(gclk));
	jxor g1194(.dina(n1494),.dinb(n1480),.dout(n1495),.clk(gclk));
	jxor g1195(.dina(w_n433_0[0]),.dinb(w_n428_0[1]),.dout(n1496),.clk(gclk));
	jxor g1196(.dina(w_n423_0[0]),.dinb(w_n412_0[0]),.dout(n1497),.clk(gclk));
	jxor g1197(.dina(n1497),.dinb(w_dff_B_zU9xVylp3_1),.dout(n1498),.clk(gclk));
	jxor g1198(.dina(n1498),.dinb(n1495),.dout(n1499),.clk(gclk));
	jand g1199(.dina(n1499),.dinb(w_n749_5[0]),.dout(n1500),.clk(gclk));
	jnot g1200(.din(n1500),.dout(n1501),.clk(gclk));
	jand g1201(.dina(w_dff_B_Z6XkuS7b3_0),.dinb(n1461),.dout(n1502),.clk(gclk));
	jor g1202(.dina(n1502),.dinb(w_G4092_4[0]),.dout(n1503),.clk(gclk));
	jnot g1203(.din(w_n750_2[2]),.dout(n1504),.clk(gclk));
	jor g1204(.dina(w_n1504_0[1]),.dinb(w_dff_B_yIyzP5Yo3_1),.dout(n1505),.clk(gclk));
	jand g1205(.dina(w_dff_B_bBgJxmY12_0),.dinb(w_n1503_0[1]),.dout(w_dff_A_UlPKT5TM8_2),.clk(gclk));
	jand g1206(.dina(w_G273_1[0]),.dinb(w_G248_3[1]),.dout(n1507),.clk(gclk));
	jand g1207(.dina(w_n471_0[2]),.dinb(w_G251_3[1]),.dout(n1508),.clk(gclk));
	jor g1208(.dina(n1508),.dinb(w_n473_1[0]),.dout(n1509),.clk(gclk));
	jor g1209(.dina(n1509),.dinb(w_dff_B_6uWvkJM58_1),.dout(n1510),.clk(gclk));
	jand g1210(.dina(w_n471_0[1]),.dinb(w_n406_3[1]),.dout(n1511),.clk(gclk));
	jand g1211(.dina(w_G273_0[2]),.dinb(w_n408_3[1]),.dout(n1512),.clk(gclk));
	jor g1212(.dina(n1512),.dinb(n1511),.dout(n1513),.clk(gclk));
	jor g1213(.dina(n1513),.dinb(w_G411_0[2]),.dout(n1514),.clk(gclk));
	jand g1214(.dina(n1514),.dinb(n1510),.dout(n1515),.clk(gclk));
	jand g1215(.dina(w_G281_1[0]),.dinb(w_G248_3[0]),.dout(n1516),.clk(gclk));
	jand g1216(.dina(w_n530_0[2]),.dinb(w_G251_3[0]),.dout(n1517),.clk(gclk));
	jor g1217(.dina(n1517),.dinb(w_n532_1[0]),.dout(n1518),.clk(gclk));
	jor g1218(.dina(n1518),.dinb(w_dff_B_w3oQLA3K1_1),.dout(n1519),.clk(gclk));
	jand g1219(.dina(w_n530_0[1]),.dinb(w_n406_3[0]),.dout(n1520),.clk(gclk));
	jand g1220(.dina(w_G281_0[2]),.dinb(w_n408_3[0]),.dout(n1521),.clk(gclk));
	jor g1221(.dina(n1521),.dinb(n1520),.dout(n1522),.clk(gclk));
	jor g1222(.dina(n1522),.dinb(w_G374_0[1]),.dout(n1523),.clk(gclk));
	jand g1223(.dina(n1523),.dinb(n1519),.dout(n1524),.clk(gclk));
	jxor g1224(.dina(n1524),.dinb(n1515),.dout(n1525),.clk(gclk));
	jor g1225(.dina(w_n483_1[0]),.dinb(w_n369_0[2]),.dout(n1526),.clk(gclk));
	jor g1226(.dina(w_G265_0[2]),.dinb(w_n366_0[2]),.dout(n1527),.clk(gclk));
	jand g1227(.dina(n1527),.dinb(w_G400_0[1]),.dout(n1528),.clk(gclk));
	jand g1228(.dina(n1528),.dinb(w_dff_B_qOYXn8xu5_1),.dout(n1529),.clk(gclk));
	jor g1229(.dina(w_G265_0[1]),.dinb(w_G254_0[2]),.dout(n1530),.clk(gclk));
	jor g1230(.dina(w_n483_0[2]),.dinb(w_G242_0[2]),.dout(n1531),.clk(gclk));
	jand g1231(.dina(n1531),.dinb(w_dff_B_XtCAGJFa0_1),.dout(n1532),.clk(gclk));
	jand g1232(.dina(n1532),.dinb(w_n485_0[2]),.dout(n1533),.clk(gclk));
	jor g1233(.dina(n1533),.dinb(n1529),.dout(n1534),.clk(gclk));
	jand g1234(.dina(w_G257_1[0]),.dinb(w_G248_2[2]),.dout(n1535),.clk(gclk));
	jand g1235(.dina(w_n518_0[2]),.dinb(w_G251_2[2]),.dout(n1536),.clk(gclk));
	jor g1236(.dina(n1536),.dinb(w_n520_0[0]),.dout(n1537),.clk(gclk));
	jor g1237(.dina(n1537),.dinb(w_dff_B_4dGYIH7l0_1),.dout(n1538),.clk(gclk));
	jand g1238(.dina(w_n518_0[1]),.dinb(w_n406_2[2]),.dout(n1539),.clk(gclk));
	jand g1239(.dina(w_G257_0[2]),.dinb(w_n408_2[2]),.dout(n1540),.clk(gclk));
	jor g1240(.dina(n1540),.dinb(n1539),.dout(n1541),.clk(gclk));
	jor g1241(.dina(n1541),.dinb(w_G389_0[1]),.dout(n1542),.clk(gclk));
	jand g1242(.dina(n1542),.dinb(n1538),.dout(n1543),.clk(gclk));
	jand g1243(.dina(w_G248_2[1]),.dinb(w_G234_1[0]),.dout(n1544),.clk(gclk));
	jand g1244(.dina(w_G251_2[1]),.dinb(w_n460_0[2]),.dout(n1545),.clk(gclk));
	jor g1245(.dina(n1545),.dinb(w_n462_0[0]),.dout(n1546),.clk(gclk));
	jor g1246(.dina(n1546),.dinb(w_dff_B_LRLQwiRy6_1),.dout(n1547),.clk(gclk));
	jand g1247(.dina(w_n406_2[1]),.dinb(w_n460_0[1]),.dout(n1548),.clk(gclk));
	jand g1248(.dina(w_n408_2[1]),.dinb(w_G234_0[2]),.dout(n1549),.clk(gclk));
	jor g1249(.dina(n1549),.dinb(n1548),.dout(n1550),.clk(gclk));
	jor g1250(.dina(n1550),.dinb(w_G435_0[1]),.dout(n1551),.clk(gclk));
	jand g1251(.dina(n1551),.dinb(n1547),.dout(n1552),.clk(gclk));
	jxor g1252(.dina(n1552),.dinb(n1543),.dout(n1553),.clk(gclk));
	jxor g1253(.dina(n1553),.dinb(w_dff_B_nIieNhIp4_1),.dout(n1554),.clk(gclk));
	jxor g1254(.dina(n1554),.dinb(w_dff_B_kI5zuntE0_1),.dout(n1555),.clk(gclk));
	jand g1255(.dina(w_G248_2[0]),.dinb(w_G226_1[0]),.dout(n1556),.clk(gclk));
	jand g1256(.dina(w_G251_2[0]),.dinb(w_n494_0[2]),.dout(n1557),.clk(gclk));
	jor g1257(.dina(n1557),.dinb(w_n496_0[1]),.dout(n1558),.clk(gclk));
	jor g1258(.dina(n1558),.dinb(w_dff_B_StMgBiOW8_1),.dout(n1559),.clk(gclk));
	jand g1259(.dina(w_n406_2[0]),.dinb(w_n494_0[1]),.dout(n1560),.clk(gclk));
	jand g1260(.dina(w_n408_2[0]),.dinb(w_G226_0[2]),.dout(n1561),.clk(gclk));
	jor g1261(.dina(n1561),.dinb(n1560),.dout(n1562),.clk(gclk));
	jor g1262(.dina(n1562),.dinb(w_G422_0[1]),.dout(n1563),.clk(gclk));
	jand g1263(.dina(n1563),.dinb(n1559),.dout(n1564),.clk(gclk));
	jxor g1264(.dina(n1564),.dinb(w_n551_0[0]),.dout(n1565),.clk(gclk));
	jor g1265(.dina(w_n369_0[1]),.dinb(w_n507_0[2]),.dout(n1566),.clk(gclk));
	jor g1266(.dina(w_n366_0[1]),.dinb(w_G218_1[0]),.dout(n1567),.clk(gclk));
	jand g1267(.dina(n1567),.dinb(w_G468_0[1]),.dout(n1568),.clk(gclk));
	jand g1268(.dina(n1568),.dinb(w_dff_B_Uu9M7lfg3_1),.dout(n1569),.clk(gclk));
	jor g1269(.dina(w_G254_0[1]),.dinb(w_G218_0[2]),.dout(n1570),.clk(gclk));
	jor g1270(.dina(w_G242_0[1]),.dinb(w_n507_0[1]),.dout(n1571),.clk(gclk));
	jand g1271(.dina(n1571),.dinb(w_dff_B_9Ce1NkLg6_1),.dout(n1572),.clk(gclk));
	jand g1272(.dina(n1572),.dinb(w_n509_0[0]),.dout(n1573),.clk(gclk));
	jor g1273(.dina(n1573),.dinb(n1569),.dout(n1574),.clk(gclk));
	jand g1274(.dina(w_G248_1[2]),.dinb(w_G210_1[0]),.dout(n1575),.clk(gclk));
	jand g1275(.dina(w_G251_1[2]),.dinb(w_n449_0[2]),.dout(n1576),.clk(gclk));
	jor g1276(.dina(n1576),.dinb(w_n451_0[0]),.dout(n1577),.clk(gclk));
	jor g1277(.dina(n1577),.dinb(w_dff_B_1M5Qhs089_1),.dout(n1578),.clk(gclk));
	jand g1278(.dina(w_n406_1[2]),.dinb(w_n449_0[1]),.dout(n1579),.clk(gclk));
	jand g1279(.dina(w_n408_1[2]),.dinb(w_G210_0[2]),.dout(n1580),.clk(gclk));
	jor g1280(.dina(n1580),.dinb(n1579),.dout(n1581),.clk(gclk));
	jor g1281(.dina(n1581),.dinb(w_G457_0[1]),.dout(n1582),.clk(gclk));
	jand g1282(.dina(n1582),.dinb(n1578),.dout(n1583),.clk(gclk));
	jxor g1283(.dina(n1583),.dinb(n1574),.dout(n1584),.clk(gclk));
	jxor g1284(.dina(n1584),.dinb(n1565),.dout(n1585),.clk(gclk));
	jxor g1285(.dina(w_dff_B_9vqikBI63_0),.dinb(n1555),.dout(n1586),.clk(gclk));
	jand g1286(.dina(n1586),.dinb(w_n749_4[2]),.dout(n1587),.clk(gclk));
	jnot g1287(.din(n1587),.dout(n1588),.clk(gclk));
	jand g1288(.dina(w_n573_0[0]),.dinb(w_n567_0[0]),.dout(n1589),.clk(gclk));
	jor g1289(.dina(w_dff_B_xFYDrjga7_0),.dinb(w_n699_0[0]),.dout(n1590),.clk(gclk));
	jnot g1290(.din(w_n559_0[0]),.dout(n1591),.clk(gclk));
	jor g1291(.dina(n1591),.dinb(w_n557_0[0]),.dout(n1592),.clk(gclk));
	jand g1292(.dina(w_n1592_0[1]),.dinb(w_n532_0[2]),.dout(n1593),.clk(gclk));
	jnot g1293(.din(w_n1593_0[1]),.dout(n1594),.clk(gclk));
	jor g1294(.dina(w_n695_0[0]),.dinb(n1594),.dout(n1595),.clk(gclk));
	jand g1295(.dina(w_n923_0[1]),.dinb(w_n473_0[2]),.dout(n1596),.clk(gclk));
	jor g1296(.dina(w_n1596_0[1]),.dinb(w_n1593_0[0]),.dout(n1597),.clk(gclk));
	jand g1297(.dina(w_dff_B_7FjASU305_0),.dinb(n1595),.dout(n1598),.clk(gclk));
	jxor g1298(.dina(w_dff_B_90XiUeBv2_0),.dinb(n1590),.dout(n1599),.clk(gclk));
	jnot g1299(.din(w_n1599_0[1]),.dout(n1600),.clk(gclk));
	jnot g1300(.din(w_n686_0[0]),.dout(n1601),.clk(gclk));
	jnot g1301(.din(w_n687_0[0]),.dout(n1602),.clk(gclk));
	jor g1302(.dina(w_n1592_0[0]),.dinb(w_n532_0[1]),.dout(n1603),.clk(gclk));
	jor g1303(.dina(w_n1596_0[0]),.dinb(w_n1603_0[1]),.dout(n1604),.clk(gclk));
	jor g1304(.dina(w_n923_0[0]),.dinb(w_n473_0[1]),.dout(n1605),.clk(gclk));
	jor g1305(.dina(w_n689_0[0]),.dinb(w_n485_0[1]),.dout(n1606),.clk(gclk));
	jand g1306(.dina(n1606),.dinb(w_n1605_0[1]),.dout(n1607),.clk(gclk));
	jand g1307(.dina(n1607),.dinb(n1604),.dout(n1608),.clk(gclk));
	jor g1308(.dina(n1608),.dinb(w_n690_0[0]),.dout(n1609),.clk(gclk));
	jor g1309(.dina(w_n1609_0[1]),.dinb(w_dff_B_bYjTbIzm8_1),.dout(n1610),.clk(gclk));
	jand g1310(.dina(n1610),.dinb(w_dff_B_SkzEZ1708_1),.dout(n1611),.clk(gclk));
	jand g1311(.dina(w_n1611_0[2]),.dinb(w_n581_0[0]),.dout(n1612),.clk(gclk));
	jxor g1312(.dina(w_n566_0[0]),.dinb(w_n561_0[1]),.dout(n1613),.clk(gclk));
	jxor g1313(.dina(w_n1613_0[1]),.dinb(w_n865_0[1]),.dout(n1614),.clk(gclk));
	jxor g1314(.dina(w_dff_B_s5FvmlJb1_0),.dinb(n1612),.dout(n1615),.clk(gclk));
	jnot g1315(.din(w_n1615_0[1]),.dout(n1616),.clk(gclk));
	jand g1316(.dina(n1616),.dinb(w_dff_B_gjBGjyHe4_1),.dout(n1617),.clk(gclk));
	jnot g1317(.din(w_G1497_0[2]),.dout(n1618),.clk(gclk));
	jand g1318(.dina(w_n1615_0[0]),.dinb(w_n1599_0[0]),.dout(n1619),.clk(gclk));
	jor g1319(.dina(n1619),.dinb(w_n1618_0[1]),.dout(n1620),.clk(gclk));
	jor g1320(.dina(n1620),.dinb(n1617),.dout(n1621),.clk(gclk));
	jand g1321(.dina(w_n1605_0[0]),.dinb(w_n1603_0[0]),.dout(n1622),.clk(gclk));
	jor g1322(.dina(n1622),.dinb(w_n694_0[0]),.dout(n1623),.clk(gclk));
	jxor g1323(.dina(w_n1613_0[0]),.dinb(w_n1609_0[0]),.dout(n1624),.clk(gclk));
	jxor g1324(.dina(n1624),.dinb(w_dff_B_7lVXvREL6_1),.dout(n1625),.clk(gclk));
	jxor g1325(.dina(w_n1611_0[1]),.dinb(w_n865_0[0]),.dout(n1626),.clk(gclk));
	jxor g1326(.dina(n1626),.dinb(w_dff_B_UNIAtMf36_1),.dout(n1627),.clk(gclk));
	jor g1327(.dina(n1627),.dinb(w_G1497_0[1]),.dout(n1628),.clk(gclk));
	jand g1328(.dina(w_dff_B_saGac2ra0_0),.dinb(n1621),.dout(n1629),.clk(gclk));
	jxor g1329(.dina(w_n579_0[1]),.dinb(w_n574_0[0]),.dout(n1630),.clk(gclk));
	jxor g1330(.dina(w_dff_B_Kf66Vzf82_0),.dinb(n1629),.dout(n1631),.clk(gclk));
	jnot g1331(.din(w_n709_0[0]),.dout(n1632),.clk(gclk));
	jand g1332(.dina(n1632),.dinb(w_n953_0[0]),.dout(n1633),.clk(gclk));
	jand g1333(.dina(w_n711_0[0]),.dinb(w_n954_0[1]),.dout(n1634),.clk(gclk));
	jor g1334(.dina(n1634),.dinb(w_n1633_0[1]),.dout(n1635),.clk(gclk));
	jxor g1335(.dina(w_n608_0[0]),.dinb(w_n592_0[0]),.dout(n1636),.clk(gclk));
	jxor g1336(.dina(n1636),.dinb(w_n602_0[0]),.dout(n1637),.clk(gclk));
	jxor g1337(.dina(w_n1637_0[1]),.dinb(n1635),.dout(n1638),.clk(gclk));
	jor g1338(.dina(w_n938_0[1]),.dinb(w_n597_0[0]),.dout(n1639),.clk(gclk));
	jand g1339(.dina(w_n609_0[0]),.dinb(w_n962_0[0]),.dout(n1640),.clk(gclk));
	jor g1340(.dina(w_dff_B_d5zF6k0X1_0),.dinb(w_n715_0[0]),.dout(n1641),.clk(gclk));
	jand g1341(.dina(w_dff_B_LNpshacK4_0),.dinb(n1639),.dout(n1642),.clk(gclk));
	jxor g1342(.dina(n1642),.dinb(w_dff_B_cWMUahs32_1),.dout(n1643),.clk(gclk));
	jand g1343(.dina(w_n1643_0[1]),.dinb(w_n703_0[1]),.dout(n1644),.clk(gclk));
	jnot g1344(.din(w_n682_0[0]),.dout(n1645),.clk(gclk));
	jor g1345(.dina(w_n1611_0[0]),.dinb(w_n684_0[0]),.dout(n1646),.clk(gclk));
	jand g1346(.dina(n1646),.dinb(w_dff_B_HtBxJ4xT0_1),.dout(n1647),.clk(gclk));
	jand g1347(.dina(w_n713_0[0]),.dinb(w_n954_0[0]),.dout(n1648),.clk(gclk));
	jor g1348(.dina(n1648),.dinb(w_n1633_0[0]),.dout(n1649),.clk(gclk));
	jxor g1349(.dina(w_dff_B_CIh7LDlr1_0),.dinb(w_n938_0[0]),.dout(n1650),.clk(gclk));
	jxor g1350(.dina(n1650),.dinb(w_n1637_0[0]),.dout(n1651),.clk(gclk));
	jand g1351(.dina(n1651),.dinb(n1647),.dout(n1652),.clk(gclk));
	jor g1352(.dina(w_n1652_0[1]),.dinb(n1644),.dout(n1653),.clk(gclk));
	jor g1353(.dina(n1653),.dinb(w_G1497_0[0]),.dout(n1654),.clk(gclk));
	jnot g1354(.din(w_n588_1[0]),.dout(n1655),.clk(gclk));
	jand g1355(.dina(w_n1652_0[0]),.dinb(w_dff_B_ibd6MUij4_1),.dout(n1656),.clk(gclk));
	jor g1356(.dina(w_n703_0[0]),.dinb(w_n588_0[2]),.dout(n1657),.clk(gclk));
	jand g1357(.dina(n1657),.dinb(w_n1643_0[0]),.dout(n1658),.clk(gclk));
	jor g1358(.dina(n1658),.dinb(n1656),.dout(n1659),.clk(gclk));
	jor g1359(.dina(n1659),.dinb(w_n1618_0[0]),.dout(n1660),.clk(gclk));
	jand g1360(.dina(n1660),.dinb(n1654),.dout(n1661),.clk(gclk));
	jxor g1361(.dina(n1661),.dinb(n1631),.dout(n1662),.clk(gclk));
	jor g1362(.dina(n1662),.dinb(w_n749_4[1]),.dout(n1663),.clk(gclk));
	jand g1363(.dina(n1663),.dinb(w_dff_B_tiupQjuw9_1),.dout(n1664),.clk(gclk));
	jor g1364(.dina(n1664),.dinb(w_G4092_3[2]),.dout(n1665),.clk(gclk));
	jor g1365(.dina(w_n1504_0[0]),.dinb(w_dff_B_kALI9UUy4_1),.dout(n1666),.clk(gclk));
	jand g1366(.dina(w_dff_B_ivEnXF2Z0_0),.dinb(w_n1665_0[1]),.dout(w_dff_A_7huooCbl2_2),.clk(gclk));
	jor g1367(.dina(w_G4088_3[1]),.dinb(w_G14_0[1]),.dout(n1668),.clk(gclk));
	jor g1368(.dina(w_n797_3[1]),.dinb(w_G64_0[1]),.dout(n1669),.clk(gclk));
	jand g1369(.dina(n1669),.dinb(w_G4087_1[1]),.dout(n1670),.clk(gclk));
	jand g1370(.dina(n1670),.dinb(w_dff_B_hkA2TYSN3_1),.dout(n1671),.clk(gclk));
	jand g1371(.dina(w_G4092_3[1]),.dinb(G97),.dout(n1672),.clk(gclk));
	jnot g1372(.din(n1672),.dout(n1673),.clk(gclk));
	jand g1373(.dina(w_dff_B_d5vIGQs41_0),.dinb(w_n1665_0[0]),.dout(n1674),.clk(gclk));
	jnot g1374(.din(w_n1674_0[2]),.dout(n1675),.clk(gclk));
	jor g1375(.dina(w_n1675_0[1]),.dinb(w_n797_3[0]),.dout(n1676),.clk(gclk));
	jand g1376(.dina(w_G4092_3[0]),.dinb(G94),.dout(n1677),.clk(gclk));
	jnot g1377(.din(n1677),.dout(n1678),.clk(gclk));
	jand g1378(.dina(w_dff_B_g7SLLSYW6_0),.dinb(w_n1503_0[0]),.dout(n1679),.clk(gclk));
	jnot g1379(.din(w_n1679_0[2]),.dout(n1680),.clk(gclk));
	jor g1380(.dina(w_n1680_0[1]),.dinb(w_G4088_3[0]),.dout(n1681),.clk(gclk));
	jand g1381(.dina(n1681),.dinb(w_n800_1[1]),.dout(n1682),.clk(gclk));
	jand g1382(.dina(n1682),.dinb(w_dff_B_z0n0vzl45_1),.dout(n1683),.clk(gclk));
	jor g1383(.dina(n1683),.dinb(w_dff_B_Dzxeri387_1),.dout(w_dff_A_8I5o8ymm2_2),.clk(gclk));
	jor g1384(.dina(w_G4089_3[1]),.dinb(w_G14_0[0]),.dout(n1685),.clk(gclk));
	jor g1385(.dina(w_n852_3[1]),.dinb(w_G64_0[0]),.dout(n1686),.clk(gclk));
	jand g1386(.dina(n1686),.dinb(w_G4090_1[1]),.dout(n1687),.clk(gclk));
	jand g1387(.dina(n1687),.dinb(w_dff_B_BTPIfn9Y7_1),.dout(n1688),.clk(gclk));
	jor g1388(.dina(w_n1675_0[0]),.dinb(w_n852_3[0]),.dout(n1689),.clk(gclk));
	jor g1389(.dina(w_n1680_0[0]),.dinb(w_G4089_3[0]),.dout(n1690),.clk(gclk));
	jand g1390(.dina(n1690),.dinb(w_n854_1[1]),.dout(n1691),.clk(gclk));
	jand g1391(.dina(n1691),.dinb(w_dff_B_mpBfkQmG0_1),.dout(n1692),.clk(gclk));
	jor g1392(.dina(n1692),.dinb(w_dff_B_KXlTl6Of8_1),.dout(w_dff_A_fkiBKvyy9_2),.clk(gclk));
	jnot g1393(.din(w_G137_3[1]),.dout(n1694),.clk(gclk));
	jnot g1394(.din(G179),.dout(n1695),.clk(gclk));
	jnot g1395(.din(w_n996_1[1]),.dout(n1696),.clk(gclk));
	jor g1396(.dina(n1696),.dinb(w_n1695_0[1]),.dout(n1697),.clk(gclk));
	jnot g1397(.din(G176),.dout(n1698),.clk(gclk));
	jnot g1398(.din(w_n994_1[1]),.dout(n1699),.clk(gclk));
	jor g1399(.dina(n1699),.dinb(w_n1698_0[1]),.dout(n1700),.clk(gclk));
	jand g1400(.dina(w_n1674_0[1]),.dinb(w_G1689_1[2]),.dout(n1701),.clk(gclk));
	jand g1401(.dina(w_n1679_0[1]),.dinb(w_n993_1[1]),.dout(n1702),.clk(gclk));
	jor g1402(.dina(n1702),.dinb(w_G1690_0[1]),.dout(n1703),.clk(gclk));
	jor g1403(.dina(n1703),.dinb(w_dff_B_yJssm8oz1_1),.dout(n1704),.clk(gclk));
	jand g1404(.dina(n1704),.dinb(w_dff_B_67NfPwbU8_1),.dout(n1705),.clk(gclk));
	jand g1405(.dina(n1705),.dinb(w_dff_B_e9Ghi6we9_1),.dout(n1706),.clk(gclk));
	jor g1406(.dina(n1706),.dinb(w_n1694_0[1]),.dout(G658),.clk(gclk));
	jnot g1407(.din(w_n1012_1[1]),.dout(n1708),.clk(gclk));
	jor g1408(.dina(n1708),.dinb(w_n1695_0[0]),.dout(n1709),.clk(gclk));
	jnot g1409(.din(w_n1014_1[1]),.dout(n1710),.clk(gclk));
	jor g1410(.dina(n1710),.dinb(w_n1698_0[0]),.dout(n1711),.clk(gclk));
	jand g1411(.dina(w_n1674_0[0]),.dinb(w_G1691_1[2]),.dout(n1712),.clk(gclk));
	jand g1412(.dina(w_n1679_0[0]),.dinb(w_n1008_1[1]),.dout(n1713),.clk(gclk));
	jor g1413(.dina(n1713),.dinb(w_G1694_0[1]),.dout(n1714),.clk(gclk));
	jor g1414(.dina(n1714),.dinb(w_dff_B_MI2lEjEz8_1),.dout(n1715),.clk(gclk));
	jand g1415(.dina(n1715),.dinb(w_dff_B_ccUhAJav5_1),.dout(n1716),.clk(gclk));
	jand g1416(.dina(n1716),.dinb(w_dff_B_xIkb5FXp4_1),.dout(n1717),.clk(gclk));
	jor g1417(.dina(n1717),.dinb(w_n1694_0[0]),.dout(G690),.clk(gclk));
	buf g1418(.din(w_G141_1[0]),.dout(w_dff_A_KBaZDOHP1_1));
	buf g1419(.din(w_G293_0[0]),.dout(w_dff_A_4s92yFbR3_1));
	buf g1420(.din(w_G3173_0[0]),.dout(w_dff_A_nC4ucAtV8_1));
	jnot g1421(.din(w_G545_0[1]),.dout(w_dff_A_RRZ9uML84_1),.clk(gclk));
	jnot g1422(.din(w_G545_0[0]),.dout(w_dff_A_xFbNgCE53_1),.clk(gclk));
	buf g1423(.din(w_G137_3[0]),.dout(w_dff_A_89syVh4x7_1));
	buf g1424(.din(w_G141_0[2]),.dout(w_dff_A_Djl8qfsF2_1));
	buf g1425(.din(w_G1_2[0]),.dout(w_dff_A_yjWZdSrI8_1));
	buf g1426(.din(w_G549_0[1]),.dout(w_dff_A_qN7P6uT37_1));
	buf g1427(.din(w_G299_0[1]),.dout(w_dff_A_PSsXJ15W0_1));
	jnot g1428(.din(w_G549_0[0]),.dout(w_dff_A_qEhQ7mZt4_1),.clk(gclk));
	buf g1429(.din(w_G1_1[2]),.dout(w_dff_A_Jr8Poux14_1));
	buf g1430(.din(w_G1_1[1]),.dout(w_dff_A_5qB1Wwgm5_1));
	buf g1431(.din(w_G1_1[0]),.dout(w_dff_A_6PibwFQP0_1));
	buf g1432(.din(w_G1_0[2]),.dout(w_dff_A_qMdRBAAX3_1));
	buf g1433(.din(w_G299_0[0]),.dout(w_dff_A_Zz1Li1Zx3_1));
	jor g1434(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(w_dff_A_2DKLk9un4_2),.clk(gclk));
	jand g1435(.dina(w_n661_0[0]),.dinb(w_n641_0[1]),.dout(w_dff_A_Bq7pFif89_2),.clk(gclk));
	jand g1436(.dina(w_n611_0[0]),.dinb(w_n588_0[1]),.dout(w_dff_A_evdjIyls0_2),.clk(gclk));
	jor g1437(.dina(w_n717_0[0]),.dinb(w_n704_0[0]),.dout(w_dff_A_QcszTcHB2_2),.clk(gclk));
	jor g1438(.dina(w_n747_0[0]),.dinb(w_n738_0[0]),.dout(w_dff_A_wQ8OfEWM6_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_dff_A_Mo9sV4jz4_1),.doutc(w_G4_0[2]),.din(w_dff_B_UYB3ZrXN6_3));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(G11));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(G14));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(w_dff_B_kXvSSlQq3_2));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(w_dff_B_2S5587Jz0_2));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(w_dff_B_lHCNbdw67_2));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(w_dff_B_t85foF892_2));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(G43));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(G46));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(w_dff_B_BpkAsc1y6_2));
	jspl3 jspl3_w_G54_0(.douta(w_dff_A_TB7xn0HS8_0),.doutb(w_dff_A_Q3jqABZ76_1),.doutc(w_G54_0[2]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(w_dff_B_D334u1qO2_2));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(w_dff_B_elWrQJ4U4_2));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(G67));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(w_dff_B_OdJBfi1i5_2));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(G73));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(G76));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(G91));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(G100));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(w_dff_B_BGVVzNqh7_2));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(w_dff_B_613TrTLX7_2));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(G109));
	jspl jspl_w_G123_0(.douta(w_dff_A_tVjet4u93_0),.doutb(w_G123_0[1]),.din(G123));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_x4dZmg6f6_0),.doutb(w_dff_A_tQnXJQLk8_1),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_tDErR2Fk5_0),.doutb(w_dff_A_BlHPAdPJ1_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_D5l59Qyj7_0),.doutb(w_dff_A_5YLdQIJG0_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_dff_A_ggIDazgF3_2),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_dff_A_7MpZfYVu0_0),.doutb(w_dff_A_twaGs9Zc4_1),.doutc(w_G137_4[2]),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_dff_A_yx0qjRcw3_0),.doutb(w_G137_5[1]),.doutc(w_G137_5[2]),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_f5mbHDtI7_0),.doutb(w_dff_A_9zUtyW7p6_1),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_rpRPwpt80_1),.doutc(w_dff_A_kkjYvLWy1_2),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_G137_8[0]),.doutb(w_G137_8[1]),.doutc(w_dff_A_RkhToDx10_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_G137_9[0]),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_4zGRtotu7_1),.doutc(w_dff_A_TccOO6vn9_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_QsBAZN6D1_0),.doutb(w_dff_A_4zSc1LyP2_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(w_dff_B_TqW49frs3_2));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(w_dff_B_dil3UexK9_2));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(w_dff_B_1lHDzU4e3_2));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(w_dff_B_D4nHgDTr3_2));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(w_dff_B_focYSCPh7_2));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(w_dff_B_Gd68TiCk6_2));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(w_dff_B_ZtJzWLSh7_2));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(w_dff_B_neZGfiL07_2));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(w_dff_B_33vZx0Wk4_2));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(w_dff_B_YqnsoghZ2_2));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(w_dff_B_4NfCGkbl4_2));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(w_dff_B_eZ8BiIdW9_2));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(w_dff_B_bLSBvltT6_2));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(w_dff_B_tFRk1qYy6_2));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(w_dff_B_TFS1KFt26_2));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(w_dff_B_F37cIesD2_2));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(w_dff_B_Z7RccH1E0_2));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(w_dff_B_nk58Ujfl0_2));
	jspl3 jspl3_w_G206_0(.douta(w_G206_0[0]),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G206_1(.douta(w_dff_A_qKmwbaOo2_0),.doutb(w_G206_1[1]),.doutc(w_G206_1[2]),.din(w_G206_0[0]));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_dff_A_kvwfYG590_2),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_G210_1[1]),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl jspl_w_G210_2(.douta(w_dff_A_YTqdcaIL5_0),.doutb(w_G210_2[1]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_dff_A_5T6fR9mq7_0),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl jspl_w_G218_2(.douta(w_dff_A_9Ucm2QPV0_0),.doutb(w_G218_2[1]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_dff_A_L2otT6Jw9_2),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_G226_1[0]),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl jspl_w_G226_2(.douta(w_dff_A_Jv4JdZ5u5_0),.doutb(w_G226_2[1]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_dff_A_2Fs1iHVf5_2),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_dff_A_6W7MCHnj4_0),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_dff_A_l8cnWHa37_1),.doutc(w_dff_A_USw4L3wP5_2),.din(G242));
	jspl jspl_w_G242_1(.douta(w_dff_A_ZPs6zkcb8_0),.doutb(w_G242_1[1]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_dff_A_h3X8GGaS8_0),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_dff_A_clY56xZi9_2),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl3 jspl3_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.doutc(w_G248_5[2]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_dff_A_kUArhjPR1_1),.doutc(w_dff_A_1XgLJ2H39_2),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_dff_A_EgLqHu1D1_0),.doutb(w_G251_1[1]),.doutc(w_dff_A_fN7vApHP4_2),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_G251_4[1]),.doutc(w_G251_4[2]),.din(w_G251_1[0]));
	jspl jspl_w_G251_5(.douta(w_dff_A_T83XRwcv4_0),.doutb(w_G251_5[1]),.din(w_G251_1[1]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl jspl_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_dff_A_I6WA4MZP3_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_G257_1[0]),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl jspl_w_G257_2(.douta(w_dff_A_m2EfBMWh9_0),.doutb(w_G257_2[1]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_dff_A_GWO37M1N8_2),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_dff_A_HdWVF1nR3_1),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_dff_A_wwkj1LBC5_2),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_dff_A_2Rh94nuT9_1),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl jspl_w_G273_2(.douta(w_dff_A_q5DKJWwU8_0),.doutb(w_G273_2[1]),.din(w_G273_0[1]));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_dff_A_iLESAI844_2),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_dff_A_4sti3Suj9_0),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_G289_0[0]),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_dff_A_G0NBzf615_1),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_dff_A_AHXN0R4U7_0),.doutb(w_dff_A_mio5KJpD3_1),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_dff_A_cCAn80oG9_0),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_dff_A_6KzOBrkF1_2),.din(G316));
	jspl jspl_w_G316_1(.douta(w_G316_1[0]),.doutb(w_G316_1[1]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_G324_0[1]),.doutc(w_dff_A_ws0VB4db8_2),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_dff_A_UNfn2Mjz9_1),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_dff_A_1BDoj2j67_1),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_dff_A_MtyJ4roH9_1),.doutc(w_G332_1[2]),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_dff_A_X7X2iXnx4_0),.doutb(w_G332_2[1]),.doutc(w_dff_A_z476YpM93_2),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_G332_3[0]),.doutb(w_G332_3[1]),.doutc(w_G332_3[2]),.din(w_G332_0[2]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl jspl_w_G338_0(.douta(w_dff_A_IPcIksHL9_0),.doutb(w_G338_0[1]),.din(G338));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_dff_A_E8mdAG5M9_2),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_dff_A_XoUV0c5b2_1),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_dff_A_FIfD5XyQ4_0),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_dff_A_mPKOD2o62_2),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_G351_1[0]),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_dff_A_3iL9ABnu6_1),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_dff_A_4Jm7U9iH9_0),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_G361_0[1]),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G361_1(.douta(w_dff_A_iuRPSOYI0_0),.doutb(w_G361_1[1]),.din(w_G361_0[0]));
	jspl jspl_w_G366_0(.douta(w_dff_A_zCn3yGKH3_0),.doutb(w_G366_0[1]),.din(G366));
	jspl jspl_w_G369_0(.douta(w_G369_0[0]),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_G374_0[0]),.doutb(w_dff_A_Dw0DhlT63_1),.doutc(w_dff_A_k06UHQ5A1_2),.din(G374));
	jspl3 jspl3_w_G374_1(.douta(w_dff_A_n93wh5bo2_0),.doutb(w_dff_A_Gn4kNrmx8_1),.doutc(w_G374_1[2]),.din(w_G374_0[0]));
	jspl3 jspl3_w_G389_0(.douta(w_G389_0[0]),.doutb(w_dff_A_GQKc1rbV2_1),.doutc(w_dff_A_Mr0oGODM8_2),.din(G389));
	jspl3 jspl3_w_G389_1(.douta(w_dff_A_Lc2dYLdb9_0),.doutb(w_dff_A_21gc5b9b6_1),.doutc(w_G389_1[2]),.din(w_G389_0[0]));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_dff_A_8feY9c7F4_1),.doutc(w_dff_A_TNgrttFd5_2),.din(G400));
	jspl3 jspl3_w_G400_1(.douta(w_dff_A_PqVa93ns6_0),.doutb(w_dff_A_sAN6ISD43_1),.doutc(w_G400_1[2]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_dff_A_ug8P8f0F0_0),.doutb(w_G411_0[1]),.doutc(w_dff_A_ai55PT6o1_2),.din(G411));
	jspl3 jspl3_w_G411_1(.douta(w_G411_1[0]),.doutb(w_G411_1[1]),.doutc(w_G411_1[2]),.din(w_G411_0[0]));
	jspl jspl_w_G411_2(.douta(w_dff_A_TnqCR82Q3_0),.doutb(w_G411_2[1]),.din(w_G411_0[1]));
	jspl3 jspl3_w_G422_0(.douta(w_G422_0[0]),.doutb(w_dff_A_V3QMQZlU8_1),.doutc(w_dff_A_6SJLGo5A5_2),.din(G422));
	jspl jspl_w_G422_1(.douta(w_dff_A_Y8ywuaNP0_0),.doutb(w_G422_1[1]),.din(w_G422_0[0]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_dff_A_Ien8KOZI6_1),.doutc(w_dff_A_fMLuO8Bl6_2),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_dff_A_hBJWfctI0_0),.doutb(w_dff_A_Lb2WQcSu6_1),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_dff_A_J674rONt9_1),.doutc(w_dff_A_f02csFex8_2),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_dff_A_VNw9zwzH9_0),.doutb(w_dff_A_Bt3PYd0s2_1),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_G457_0[0]),.doutb(w_dff_A_oskN5ta20_1),.doutc(w_dff_A_2y2w50oe2_2),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_dff_A_5NXR3OFP8_0),.doutb(w_dff_A_U8qclugG4_1),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_dff_A_CBiKKZIS9_1),.doutc(w_dff_A_iNfwLSLT6_2),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_dff_A_YYWsJkFt2_0),.doutb(w_dff_A_7boYskag2_1),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_dff_A_HdGKWoCy4_0),.doutb(w_dff_A_DMdqylml7_1),.doutc(w_G479_0[2]),.din(G479));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_dff_A_zutWcC9k7_1),.doutc(w_dff_A_ZvPz6YQa3_2),.din(G490));
	jspl jspl_w_G490_1(.douta(w_dff_A_Knhhl1uN2_0),.doutb(w_G490_1[1]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_dff_A_zj7BXK0S0_0),.doutb(w_G503_0[1]),.doutc(w_dff_A_tnwJ9HxF4_2),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_G503_1[0]),.doutb(w_G503_1[1]),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl jspl_w_G503_2(.douta(w_dff_A_c0cF66of2_0),.doutb(w_G503_2[1]),.din(w_G503_0[1]));
	jspl3 jspl3_w_G514_0(.douta(w_dff_A_4vW2gdeH9_0),.doutb(w_G514_0[1]),.doutc(w_dff_A_QJgWHiKz1_2),.din(G514));
	jspl3 jspl3_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.doutc(w_G514_1[2]),.din(w_G514_0[0]));
	jspl jspl_w_G514_2(.douta(w_G514_2[0]),.doutb(w_G514_2[1]),.din(w_G514_0[1]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_dff_A_06pQuPHL0_1),.doutc(w_dff_A_vVYz0nIU7_2),.din(G523));
	jspl3 jspl3_w_G523_1(.douta(w_dff_A_a1pkJkDq3_0),.doutb(w_dff_A_5Ds71fVU2_1),.doutc(w_G523_1[2]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_dff_A_zizoQuCR7_0),.doutb(w_G534_0[1]),.doutc(w_dff_A_OxQjbA5L0_2),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_G534_1[0]),.doutb(w_G534_1[1]),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl jspl_w_G534_2(.douta(w_dff_A_jEfd3TcK5_0),.doutb(w_G534_2[1]),.din(w_G534_0[1]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_dff_A_2cTOs3ML8_0),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_dff_A_ezjoubcI2_0),.doutb(w_dff_A_EP0AG1Mv3_1),.doutc(w_G1497_0[2]),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_dff_A_71Hv8wWq6_1),.doutc(w_dff_A_MHwIKS9y3_2),.din(G1689));
	jspl3 jspl3_w_G1689_1(.douta(w_dff_A_SXzeJC4S4_0),.doutb(w_G1689_1[1]),.doutc(w_dff_A_KG0OdvOF6_2),.din(w_G1689_0[0]));
	jspl3 jspl3_w_G1689_2(.douta(w_dff_A_6wDgPfXN7_0),.doutb(w_G1689_2[1]),.doutc(w_dff_A_aNM8e70a3_2),.din(w_G1689_0[1]));
	jspl3 jspl3_w_G1689_3(.douta(w_dff_A_wZh9lAPx0_0),.doutb(w_dff_A_logOGiod7_1),.doutc(w_G1689_3[2]),.din(w_G1689_0[2]));
	jspl3 jspl3_w_G1689_4(.douta(w_dff_A_QuEJt7JU6_0),.doutb(w_dff_A_90mI8wQY7_1),.doutc(w_G1689_4[2]),.din(w_G1689_1[0]));
	jspl jspl_w_G1689_5(.douta(w_G1689_5[0]),.doutb(w_G1689_5[1]),.din(w_G1689_1[1]));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_dff_A_WFpyXQE98_1),.doutc(w_G1690_0[2]),.din(G1690));
	jspl jspl_w_G1690_1(.douta(w_G1690_1[0]),.doutb(w_dff_A_7MZiC1pn7_1),.din(w_G1690_0[0]));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_dff_A_1UZ6pyuM0_1),.doutc(w_dff_A_vIIwWw7D2_2),.din(G1691));
	jspl3 jspl3_w_G1691_1(.douta(w_G1691_1[0]),.doutb(w_G1691_1[1]),.doutc(w_dff_A_qR4PjBAd9_2),.din(w_G1691_0[0]));
	jspl3 jspl3_w_G1691_2(.douta(w_dff_A_OnstN0Yx8_0),.doutb(w_G1691_2[1]),.doutc(w_dff_A_T3jpC6XO6_2),.din(w_G1691_0[1]));
	jspl3 jspl3_w_G1691_3(.douta(w_dff_A_Txew2Vfp7_0),.doutb(w_dff_A_dUMO3B2W6_1),.doutc(w_G1691_3[2]),.din(w_G1691_0[2]));
	jspl3 jspl3_w_G1691_4(.douta(w_dff_A_9EMamk5B2_0),.doutb(w_dff_A_gA8plgWv0_1),.doutc(w_G1691_4[2]),.din(w_G1691_1[0]));
	jspl jspl_w_G1691_5(.douta(w_G1691_5[0]),.doutb(w_dff_A_RC3RjUy58_1),.din(w_G1691_1[1]));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_dff_A_MVuEkKuY4_1),.doutc(w_dff_A_VuDmMeGV7_2),.din(G1694));
	jspl jspl_w_G1694_1(.douta(w_G1694_1[0]),.doutb(w_G1694_1[1]),.din(w_G1694_0[0]));
	jspl3 jspl3_w_G2174_0(.douta(w_dff_A_iO8l3Xcp1_0),.doutb(w_dff_A_inQvp69a0_1),.doutc(w_G2174_0[2]),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_dff_A_sfF8rck74_0),.doutb(w_dff_A_LxfFmvmr5_1),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(w_dff_B_whIVPNaU5_3));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_dff_A_5vksmMD30_0),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_G3724_0[0]),.doutb(w_G3724_0[1]),.doutc(w_dff_A_HSDjMAYL4_2),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_dff_A_q6Ybc1Cz7_1),.doutc(w_dff_A_xUOYB4Xr8_2),.din(G4087));
	jspl3 jspl3_w_G4087_1(.douta(w_G4087_1[0]),.doutb(w_dff_A_Qd0zoQ9U3_1),.doutc(w_dff_A_huOUs4Y20_2),.din(w_G4087_0[0]));
	jspl3 jspl3_w_G4087_2(.douta(w_G4087_2[0]),.doutb(w_G4087_2[1]),.doutc(w_G4087_2[2]),.din(w_G4087_0[1]));
	jspl3 jspl3_w_G4087_3(.douta(w_G4087_3[0]),.doutb(w_G4087_3[1]),.doutc(w_G4087_3[2]),.din(w_G4087_0[2]));
	jspl3 jspl3_w_G4087_4(.douta(w_dff_A_QYL6DxgV9_0),.doutb(w_dff_A_OfrUFjPQ7_1),.doutc(w_G4087_4[2]),.din(w_G4087_1[0]));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_G4088_0[2]),.din(G4088));
	jspl3 jspl3_w_G4088_1(.douta(w_G4088_1[0]),.doutb(w_G4088_1[1]),.doutc(w_G4088_1[2]),.din(w_G4088_0[0]));
	jspl3 jspl3_w_G4088_2(.douta(w_G4088_2[0]),.doutb(w_G4088_2[1]),.doutc(w_G4088_2[2]),.din(w_G4088_0[1]));
	jspl3 jspl3_w_G4088_3(.douta(w_dff_A_kH3PP8cX2_0),.doutb(w_G4088_3[1]),.doutc(w_G4088_3[2]),.din(w_G4088_0[2]));
	jspl3 jspl3_w_G4088_4(.douta(w_dff_A_n56Cg8U79_0),.doutb(w_G4088_4[1]),.doutc(w_dff_A_3MTawk6p2_2),.din(w_G4088_1[0]));
	jspl3 jspl3_w_G4088_5(.douta(w_G4088_5[0]),.doutb(w_dff_A_cNzuEArp5_1),.doutc(w_G4088_5[2]),.din(w_G4088_1[1]));
	jspl3 jspl3_w_G4088_6(.douta(w_dff_A_DnGrOMJs5_0),.doutb(w_G4088_6[1]),.doutc(w_dff_A_wDrieCip9_2),.din(w_G4088_1[2]));
	jspl3 jspl3_w_G4088_7(.douta(w_G4088_7[0]),.doutb(w_dff_A_SGXCpmyO5_1),.doutc(w_G4088_7[2]),.din(w_G4088_2[0]));
	jspl3 jspl3_w_G4088_8(.douta(w_dff_A_neKuS7Eu8_0),.doutb(w_G4088_8[1]),.doutc(w_dff_A_zDaWfg2a1_2),.din(w_G4088_2[1]));
	jspl3 jspl3_w_G4088_9(.douta(w_G4088_9[0]),.doutb(w_dff_A_8wb7EXNr3_1),.doutc(w_G4088_9[2]),.din(w_G4088_2[2]));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_G4089_0[2]),.din(G4089));
	jspl3 jspl3_w_G4089_1(.douta(w_G4089_1[0]),.doutb(w_G4089_1[1]),.doutc(w_G4089_1[2]),.din(w_G4089_0[0]));
	jspl3 jspl3_w_G4089_2(.douta(w_G4089_2[0]),.doutb(w_G4089_2[1]),.doutc(w_G4089_2[2]),.din(w_G4089_0[1]));
	jspl3 jspl3_w_G4089_3(.douta(w_dff_A_EoOpLKUe9_0),.doutb(w_G4089_3[1]),.doutc(w_G4089_3[2]),.din(w_G4089_0[2]));
	jspl3 jspl3_w_G4089_4(.douta(w_dff_A_KR9zwP2a9_0),.doutb(w_G4089_4[1]),.doutc(w_dff_A_u9j9nshs9_2),.din(w_G4089_1[0]));
	jspl3 jspl3_w_G4089_5(.douta(w_G4089_5[0]),.doutb(w_dff_A_AZUk2N372_1),.doutc(w_dff_A_4PPCRYOm0_2),.din(w_G4089_1[1]));
	jspl3 jspl3_w_G4089_6(.douta(w_G4089_6[0]),.doutb(w_G4089_6[1]),.doutc(w_dff_A_Uy0iffnN3_2),.din(w_G4089_1[2]));
	jspl3 jspl3_w_G4089_7(.douta(w_dff_A_ttTEApFA6_0),.doutb(w_G4089_7[1]),.doutc(w_dff_A_AtGQZzA59_2),.din(w_G4089_2[0]));
	jspl3 jspl3_w_G4089_8(.douta(w_G4089_8[0]),.doutb(w_dff_A_WeY6qbfv3_1),.doutc(w_G4089_8[2]),.din(w_G4089_2[1]));
	jspl3 jspl3_w_G4089_9(.douta(w_G4089_9[0]),.doutb(w_dff_A_I5dEYBgk2_1),.doutc(w_G4089_9[2]),.din(w_G4089_2[2]));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_dff_A_BYXvFlgx9_1),.doutc(w_dff_A_f0KPsERX4_2),.din(G4090));
	jspl3 jspl3_w_G4090_1(.douta(w_G4090_1[0]),.doutb(w_dff_A_ksc0atqM3_1),.doutc(w_dff_A_sRvNW2HZ1_2),.din(w_G4090_0[0]));
	jspl3 jspl3_w_G4090_2(.douta(w_G4090_2[0]),.doutb(w_G4090_2[1]),.doutc(w_dff_A_uRkmLDwz7_2),.din(w_G4090_0[1]));
	jspl3 jspl3_w_G4090_3(.douta(w_G4090_3[0]),.doutb(w_dff_A_klxH40F92_1),.doutc(w_dff_A_7JjJKAlK5_2),.din(w_G4090_0[2]));
	jspl3 jspl3_w_G4090_4(.douta(w_dff_A_8kpK9Msz0_0),.doutb(w_dff_A_26cKSgzW0_1),.doutc(w_G4090_4[2]),.din(w_G4090_1[0]));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_dff_A_TYG55EF44_1),.doutc(w_dff_A_4Hx3joJk7_2),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_dff_A_hln36Jja8_0),.doutb(w_dff_A_0NTHthet9_1),.doutc(w_G4091_1[2]),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_dff_A_Biw7FZMg8_0),.doutb(w_dff_A_mOsICq916_1),.doutc(w_G4091_2[2]),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4091_3(.douta(w_G4091_3[0]),.doutb(w_dff_A_hjTmyCYm9_1),.doutc(w_dff_A_1d6GvdyF2_2),.din(w_G4091_0[2]));
	jspl3 jspl3_w_G4091_4(.douta(w_dff_A_wEzJNpno8_0),.doutb(w_G4091_4[1]),.doutc(w_dff_A_ZzP2sz4o8_2),.din(w_G4091_1[0]));
	jspl3 jspl3_w_G4091_5(.douta(w_dff_A_FZrxiTix6_0),.doutb(w_G4091_5[1]),.doutc(w_dff_A_awc91F4R1_2),.din(w_G4091_1[1]));
	jspl jspl_w_G4091_6(.douta(w_dff_A_7ltQG4E96_0),.doutb(w_G4091_6[1]),.din(w_G4091_1[2]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_dff_A_TPiTsZpu7_1),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_dff_A_B5jVEXVJ8_0),.doutb(w_G4092_1[1]),.doutc(w_dff_A_MqQyiEH24_2),.din(w_G4092_0[0]));
	jspl3 jspl3_w_G4092_2(.douta(w_dff_A_UQCIH12x2_0),.doutb(w_dff_A_tnyGzhZ58_1),.doutc(w_G4092_2[2]),.din(w_G4092_0[1]));
	jspl3 jspl3_w_G4092_3(.douta(w_G4092_3[0]),.doutb(w_G4092_3[1]),.doutc(w_dff_A_MOuVyOFp9_2),.din(w_G4092_0[2]));
	jspl3 jspl3_w_G4092_4(.douta(w_dff_A_8XkyozXV8_0),.doutb(w_G4092_4[1]),.doutc(w_G4092_4[2]),.din(w_G4092_1[0]));
	jspl3 jspl3_w_G4092_5(.douta(w_dff_A_AOhrr9dn7_0),.doutb(w_dff_A_lB8jkucz9_1),.doutc(w_G4092_5[2]),.din(w_G4092_1[1]));
	jspl3 jspl3_w_G4092_6(.douta(w_G4092_6[0]),.doutb(w_dff_A_1qyT3Zbc1_1),.doutc(w_dff_A_bqRP7G405_2),.din(w_G4092_1[2]));
	jspl3 jspl3_w_G4092_7(.douta(w_G4092_7[0]),.doutb(w_G4092_7[1]),.doutc(w_dff_A_sXs48mAJ2_2),.din(w_G4092_2[0]));
	jspl3 jspl3_w_G4092_8(.douta(w_G4092_8[0]),.doutb(w_dff_A_aIHJe3SX5_1),.doutc(w_dff_A_fsG94DFF4_2),.din(w_G4092_2[1]));
	jspl3 jspl3_w_G4092_9(.douta(w_dff_A_OQJ74M3V3_0),.doutb(w_dff_A_Nuq3dACF0_1),.doutc(w_G4092_9[2]),.din(w_G4092_2[2]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(w_dff_A_vVTXHN0Y8_1),.din(G599_fa_));
	jspl jspl_w_G601_0(.douta(w_G601_0),.doutb(w_dff_A_vJT8vmhz2_1),.din(G601_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(w_dff_A_ICrsPWT71_1),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_G809_1[0]),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_G809_2[2]),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_G809_3[0]),.doutb(w_G809_3[1]),.doutc(w_dff_A_CwjD3V1R2_2),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(w_dff_A_AujOhDyB6_1),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(w_dff_A_JwnIrGQk0_1),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(w_dff_A_VFIEsrzx7_1),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(w_dff_A_ZyftNr317_1),.din(G861_fa_));
	jspl jspl_w_G623_0(.douta(w_G623_0),.doutb(w_dff_A_mtoJbP4h4_1),.din(G623_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(w_dff_A_0TreeCMY9_1),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(w_dff_A_aRP8PpQw1_1),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(w_dff_A_cWVz6Ubw9_1),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(w_dff_A_Xcf1pYNP1_1),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(w_dff_A_4fYXhbSz2_1),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(w_dff_A_cecI00zW2_1),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(w_dff_A_j4wRy3eY7_1),.din(G877_fa_));
	jspl jspl_w_G998_0(.douta(w_G998_0),.doutb(w_dff_A_LDVmy6xf9_1),.din(G998_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(w_dff_A_rvkGvTDO1_1),.din(G830_fa_));
	jspl jspl_w_G865_0(.douta(w_G865_0),.doutb(w_dff_A_6AWDkRJl7_1),.din(G865_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(w_dff_A_XkPdcrtq8_1),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(w_dff_B_uZZ3q6Nx0_2));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.doutc(w_n369_0[2]),.din(n369));
	jspl3 jspl3_w_n369_1(.douta(w_n369_1[0]),.doutb(w_n369_1[1]),.doutc(w_n369_1[2]),.din(w_n369_0[0]));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl3 jspl3_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.doutc(w_n374_0[2]),.din(n374));
	jspl jspl_w_n374_1(.douta(w_n374_1[0]),.doutb(w_n374_1[1]),.din(w_n374_0[0]));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl3 jspl3_w_n375_1(.douta(w_n375_1[0]),.doutb(w_n375_1[1]),.doutc(w_n375_1[2]),.din(w_n375_0[0]));
	jspl3 jspl3_w_n375_2(.douta(w_n375_2[0]),.doutb(w_n375_2[1]),.doutc(w_n375_2[2]),.din(w_n375_0[1]));
	jspl3 jspl3_w_n375_3(.douta(w_n375_3[0]),.doutb(w_n375_3[1]),.doutc(w_n375_3[2]),.din(w_n375_0[2]));
	jspl3 jspl3_w_n375_4(.douta(w_n375_4[0]),.doutb(w_n375_4[1]),.doutc(w_n375_4[2]),.din(w_n375_1[0]));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_dff_A_ITtg9bl70_2),.din(w_dff_B_XnDd9siy9_3));
	jspl jspl_w_n377_1(.douta(w_dff_A_NcYLiKqL2_0),.doutb(w_n377_1[1]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.doutc(w_n378_0[2]),.din(n378));
	jspl3 jspl3_w_n378_1(.douta(w_n378_1[0]),.doutb(w_n378_1[1]),.doutc(w_n378_1[2]),.din(w_n378_0[0]));
	jspl3 jspl3_w_n378_2(.douta(w_n378_2[0]),.doutb(w_n378_2[1]),.doutc(w_n378_2[2]),.din(w_n378_0[1]));
	jspl3 jspl3_w_n378_3(.douta(w_n378_3[0]),.doutb(w_n378_3[1]),.doutc(w_n378_3[2]),.din(w_n378_0[2]));
	jspl3 jspl3_w_n378_4(.douta(w_n378_4[0]),.doutb(w_n378_4[1]),.doutc(w_n378_4[2]),.din(w_n378_1[0]));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_dff_A_xx4rnksF6_2),.din(w_dff_B_5144iDOd1_3));
	jspl jspl_w_n389_1(.douta(w_dff_A_DrDwCHlH4_0),.doutb(w_n389_1[1]),.din(w_n389_0[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n401_0(.douta(w_dff_A_Mpz7Wox11_0),.doutb(w_n401_0[1]),.din(w_dff_B_4XfIYN468_2));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.doutc(w_n406_0[2]),.din(n406));
	jspl3 jspl3_w_n406_1(.douta(w_n406_1[0]),.doutb(w_n406_1[1]),.doutc(w_n406_1[2]),.din(w_n406_0[0]));
	jspl3 jspl3_w_n406_2(.douta(w_n406_2[0]),.doutb(w_n406_2[1]),.doutc(w_n406_2[2]),.din(w_n406_0[1]));
	jspl3 jspl3_w_n406_3(.douta(w_n406_3[0]),.doutb(w_n406_3[1]),.doutc(w_n406_3[2]),.din(w_n406_0[2]));
	jspl3 jspl3_w_n406_4(.douta(w_n406_4[0]),.doutb(w_n406_4[1]),.doutc(w_n406_4[2]),.din(w_n406_1[0]));
	jspl jspl_w_n406_5(.douta(w_n406_5[0]),.doutb(w_n406_5[1]),.din(w_n406_1[1]));
	jspl3 jspl3_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.doutc(w_n408_0[2]),.din(n408));
	jspl3 jspl3_w_n408_1(.douta(w_n408_1[0]),.doutb(w_n408_1[1]),.doutc(w_n408_1[2]),.din(w_n408_0[0]));
	jspl3 jspl3_w_n408_2(.douta(w_n408_2[0]),.doutb(w_n408_2[1]),.doutc(w_n408_2[2]),.din(w_n408_0[1]));
	jspl3 jspl3_w_n408_3(.douta(w_n408_3[0]),.doutb(w_n408_3[1]),.doutc(w_n408_3[2]),.din(w_n408_0[2]));
	jspl3 jspl3_w_n408_4(.douta(w_n408_4[0]),.doutb(w_n408_4[1]),.doutc(w_n408_4[2]),.din(w_n408_1[0]));
	jspl3 jspl3_w_n408_5(.douta(w_n408_5[0]),.doutb(w_n408_5[1]),.doutc(w_n408_5[2]),.din(w_n408_1[1]));
	jspl3 jspl3_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.doutc(w_n412_0[2]),.din(n412));
	jspl jspl_w_n414_0(.douta(w_dff_A_VNOLxWZW2_0),.doutb(w_n414_0[1]),.din(w_dff_B_ONHJmS7E4_2));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl3 jspl3_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.doutc(w_n423_0[2]),.din(n423));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_n425_0[2]),.din(n425));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_dff_A_H8tCWae42_1),.doutc(w_n428_0[2]),.din(n428));
	jspl jspl_w_n428_1(.douta(w_n428_1[0]),.doutb(w_dff_A_KNKfWtxB6_1),.din(w_n428_0[0]));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl3 jspl3_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.doutc(w_n433_0[2]),.din(n433));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl jspl_w_n435_2(.douta(w_n435_2[0]),.doutb(w_n435_2[1]),.din(w_n435_0[1]));
	jspl jspl_w_n437_0(.douta(w_dff_A_Unoy0Uw58_0),.doutb(w_n437_0[1]),.din(w_dff_B_FbiuPYQL1_2));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_dff_A_N1aipDxO8_1),.doutc(w_n451_0[2]),.din(w_dff_B_MEJV5t838_3));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_dff_A_WtRAsExu8_1),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_JEmkZMiG7_1),.doutc(w_n462_0[2]),.din(w_dff_B_MdGS8fv19_3));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl3 jspl3_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.doutc(w_n471_1[2]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_dff_A_AAJrBaP18_1),.doutc(w_dff_A_4IPrpr5s0_2),.din(w_dff_B_7icCghZd5_3));
	jspl jspl_w_n473_1(.douta(w_n473_1[0]),.doutb(w_n473_1[1]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.doutc(w_n483_0[2]),.din(n483));
	jspl3 jspl3_w_n483_1(.douta(w_n483_1[0]),.doutb(w_n483_1[1]),.doutc(w_n483_1[2]),.din(w_n483_0[0]));
	jspl jspl_w_n483_2(.douta(w_n483_2[0]),.doutb(w_n483_2[1]),.din(w_n483_0[1]));
	jspl3 jspl3_w_n485_0(.douta(w_n485_0[0]),.doutb(w_dff_A_iRVMvfNT1_1),.doutc(w_dff_A_DxScrfm78_2),.din(w_dff_B_Kg99jZtm0_3));
	jspl jspl_w_n485_1(.douta(w_dff_A_PEoHeZnd2_0),.doutb(w_n485_1[1]),.din(w_n485_0[0]));
	jspl jspl_w_n493_0(.douta(w_n493_0[0]),.doutb(w_n493_0[1]),.din(n493));
	jspl3 jspl3_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.doutc(w_n494_0[2]),.din(n494));
	jspl3 jspl3_w_n494_1(.douta(w_n494_1[0]),.doutb(w_n494_1[1]),.doutc(w_n494_1[2]),.din(w_n494_0[0]));
	jspl3 jspl3_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.doutc(w_dff_A_cKTpejlu2_2),.din(w_dff_B_sAWPCcwN2_3));
	jspl jspl_w_n496_1(.douta(w_dff_A_07Q4LIuX7_0),.doutb(w_n496_1[1]),.din(w_n496_0[0]));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl3 jspl3_w_n509_0(.douta(w_dff_A_6Kekg5Mn7_0),.doutb(w_dff_A_T9ZByXAe4_1),.doutc(w_n509_0[2]),.din(w_dff_B_tNG1fmo45_3));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl3 jspl3_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.doutc(w_n518_1[2]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n520_0(.douta(w_n520_0[0]),.doutb(w_dff_A_1JaE5bQI8_1),.doutc(w_n520_0[2]),.din(w_dff_B_rPXNYChq5_3));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl3 jspl3_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.doutc(w_n530_1[2]),.din(w_n530_0[0]));
	jspl3 jspl3_w_n532_0(.douta(w_n532_0[0]),.doutb(w_dff_A_7c7731Fg5_1),.doutc(w_dff_A_toLIV1WJ6_2),.din(w_dff_B_AdYaPkP42_3));
	jspl jspl_w_n532_1(.douta(w_n532_1[0]),.doutb(w_n532_1[1]),.din(w_n532_0[0]));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.doutc(w_n551_0[2]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl3 jspl3_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.doutc(w_n556_5[2]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n556_6(.douta(w_n556_6[0]),.doutb(w_n556_6[1]),.doutc(w_n556_6[2]),.din(w_n556_1[2]));
	jspl3 jspl3_w_n556_7(.douta(w_n556_7[0]),.doutb(w_n556_7[1]),.doutc(w_n556_7[2]),.din(w_n556_2[0]));
	jspl jspl_w_n556_8(.douta(w_n556_8[0]),.doutb(w_n556_8[1]),.din(w_n556_2[1]));
	jspl jspl_w_n557_0(.douta(w_dff_A_IWEv4cNs6_0),.doutb(w_n557_0[1]),.din(n557));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_dff_A_TQ7VFzdl0_1),.din(n559));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n561_1(.douta(w_n561_1[0]),.doutb(w_n561_1[1]),.din(w_n561_0[0]));
	jspl jspl_w_n562_0(.douta(w_dff_A_ASeZkNt49_0),.doutb(w_n562_0[1]),.din(n562));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_jlXW2jXy4_1),.din(n564));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n569_0(.douta(w_dff_A_UsLowW160_0),.doutb(w_n569_0[1]),.din(n569));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_dff_A_ehmpgBWb6_1),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_dff_A_3SbmSsG54_0),.doutb(w_dff_A_0hLVK2JU2_1),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_dff_A_iC3wlEyD1_1),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.doutc(w_n578_0[2]),.din(n578));
	jspl jspl_w_n578_1(.douta(w_n578_1[0]),.doutb(w_n578_1[1]),.din(w_n578_0[0]));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_dff_A_rxH08Yi38_1),.doutc(w_dff_A_1OUAiVoj1_2),.din(n579));
	jspl jspl_w_n579_1(.douta(w_n579_1[0]),.doutb(w_dff_A_E7y64BeT8_1),.din(w_n579_0[0]));
	jspl jspl_w_n581_0(.douta(w_dff_A_wABGtHPL5_0),.doutb(w_n581_0[1]),.din(n581));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n586_1(.douta(w_n586_1[0]),.doutb(w_n586_1[1]),.din(w_n586_0[0]));
	jspl jspl_w_n587_0(.douta(w_n587_0[0]),.doutb(w_dff_A_LMNkz2cr9_1),.din(n587));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_dff_A_7ToaC0wk1_2),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.doutc(w_n591_0[2]),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_dff_A_hBJz7Zz76_0),.doutb(w_n592_0[1]),.doutc(w_dff_A_aRbml7jY4_2),.din(n592));
	jspl3 jspl3_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl jspl_w_n596_1(.douta(w_n596_1[0]),.doutb(w_n596_1[1]),.din(w_n596_0[0]));
	jspl3 jspl3_w_n597_0(.douta(w_dff_A_ExtVVazX9_0),.doutb(w_n597_0[1]),.doutc(w_n597_0[2]),.din(n597));
	jspl3 jspl3_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.doutc(w_n601_0[2]),.din(n601));
	jspl jspl_w_n601_1(.douta(w_n601_1[0]),.doutb(w_n601_1[1]),.din(w_n601_0[0]));
	jspl3 jspl3_w_n602_0(.douta(w_dff_A_soHz0zdW4_0),.doutb(w_n602_0[1]),.doutc(w_n602_0[2]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n607_1(.douta(w_n607_1[0]),.doutb(w_n607_1[1]),.din(w_n607_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_dff_A_RpA6Tcj95_1),.doutc(w_dff_A_T3e2k0WO5_2),.din(n608));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_dff_A_Jx6W1WJ93_1),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n611_0(.douta(w_n611_0[0]),.doutb(w_dff_A_wK0ga2Vk4_1),.doutc(w_n611_0[2]),.din(w_dff_B_Y78scTpD4_3));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.doutc(w_n613_1[2]),.din(w_n613_0[0]));
	jspl3 jspl3_w_n613_2(.douta(w_n613_2[0]),.doutb(w_n613_2[1]),.doutc(w_n613_2[2]),.din(w_n613_0[1]));
	jspl3 jspl3_w_n613_3(.douta(w_n613_3[0]),.doutb(w_n613_3[1]),.doutc(w_n613_3[2]),.din(w_n613_0[2]));
	jspl3 jspl3_w_n613_4(.douta(w_n613_4[0]),.doutb(w_n613_4[1]),.doutc(w_n613_4[2]),.din(w_n613_1[0]));
	jspl3 jspl3_w_n613_5(.douta(w_n613_5[0]),.doutb(w_n613_5[1]),.doutc(w_n613_5[2]),.din(w_n613_1[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_dff_A_4U3jWDXQ1_1),.doutc(w_dff_A_qMHXqdRa3_2),.din(n618));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_dff_A_Q12d3uM86_1),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n619_1(.douta(w_n619_1[0]),.doutb(w_n619_1[1]),.doutc(w_n619_1[2]),.din(w_n619_0[0]));
	jspl3 jspl3_w_n620_0(.douta(w_n620_0[0]),.doutb(w_dff_A_NKahmuzI0_1),.doutc(w_dff_A_igeem2lH7_2),.din(n620));
	jspl jspl_w_n620_1(.douta(w_n620_1[0]),.doutb(w_dff_A_QSN4LlY07_1),.din(w_n620_0[0]));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_dff_A_ckaHTcbS1_1),.din(n621));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_dff_A_UsjWnzyx7_0),.doutb(w_dff_A_Zmwi3UTf3_1),.doutc(w_n624_0[2]),.din(w_dff_B_4iQ1YXwM3_3));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_dff_A_2JWxP9z98_1),.din(n625));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl jspl_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n628_0(.douta(w_dff_A_uudzYH4a6_0),.doutb(w_n628_0[1]),.doutc(w_dff_A_DIDKx7dg3_2),.din(n628));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_dff_A_vKyo0vsz3_1),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n635_1(.douta(w_dff_A_GtdLA4qw5_0),.doutb(w_n635_1[1]),.din(w_n635_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.doutc(w_n637_0[2]),.din(n637));
	jspl jspl_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.din(n638));
	jspl3 jspl3_w_n639_0(.douta(w_dff_A_9qjiZtE58_0),.doutb(w_n639_0[1]),.doutc(w_n639_0[2]),.din(n639));
	jspl jspl_w_n640_0(.douta(w_dff_A_ZlM4TwFe9_0),.doutb(w_n640_0[1]),.din(n640));
	jspl3 jspl3_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.doutc(w_dff_A_ZBOaviyN3_2),.din(n641));
	jspl3 jspl3_w_n641_1(.douta(w_n641_1[0]),.doutb(w_n641_1[1]),.doutc(w_n641_1[2]),.din(w_n641_0[0]));
	jspl3 jspl3_w_n644_0(.douta(w_dff_A_908jh8XE2_0),.doutb(w_n644_0[1]),.doutc(w_dff_A_zyvbQmbi4_2),.din(n644));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_dff_A_Pdohg5pg3_1),.doutc(w_dff_A_z5GEAU9j4_2),.din(n648));
	jspl jspl_w_n648_1(.douta(w_n648_1[0]),.doutb(w_n648_1[1]),.din(w_n648_0[0]));
	jspl jspl_w_n649_0(.douta(w_dff_A_RofdZU6q4_0),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n653_0(.douta(w_dff_A_HWxL4K037_0),.doutb(w_n653_0[1]),.doutc(w_n653_0[2]),.din(n653));
	jspl3 jspl3_w_n654_0(.douta(w_dff_A_v3GcPNiR7_0),.doutb(w_n654_0[1]),.doutc(w_n654_0[2]),.din(w_dff_B_vw3vRAA64_3));
	jspl3 jspl3_w_n654_1(.douta(w_n654_1[0]),.doutb(w_dff_A_b3hINvNF7_1),.doutc(w_n654_1[2]),.din(w_n654_0[0]));
	jspl3 jspl3_w_n654_2(.douta(w_dff_A_dQzCsD9g8_0),.doutb(w_n654_2[1]),.doutc(w_n654_2[2]),.din(w_n654_0[1]));
	jspl3 jspl3_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.doutc(w_n658_0[2]),.din(n658));
	jspl jspl_w_n658_1(.douta(w_n658_1[0]),.doutb(w_n658_1[1]),.din(w_n658_0[0]));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_dff_A_lpXRusux6_2),.din(n660));
	jspl jspl_w_n660_1(.douta(w_dff_A_q7uSuu5a5_0),.doutb(w_n660_1[1]),.din(w_n660_0[0]));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(w_dff_B_fOGWVeyJ0_2));
	jspl jspl_w_n670_0(.douta(w_n670_0[0]),.doutb(w_n670_0[1]),.din(n670));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl3 jspl3_w_n682_0(.douta(w_n682_0[0]),.doutb(w_dff_A_5USy8GVJ0_1),.doutc(w_dff_A_5VPYhO5W0_2),.din(n682));
	jspl jspl_w_n684_0(.douta(w_dff_A_N5RCJTb54_0),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_dff_A_m5S8r6zo1_0),.doutb(w_n685_0[1]),.din(w_dff_B_FTkfTvPN9_2));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_dff_A_1VkHJzJt5_1),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_dff_A_64xSURsP6_1),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_dff_A_VXalCOdH3_0),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n692_0(.douta(w_dff_A_FyyMCPEK9_0),.doutb(w_n692_0[1]),.din(n692));
	jspl3 jspl3_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.doutc(w_n694_0[2]),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_dff_A_OMQ6DNjv3_0),.doutb(w_dff_A_YkubTpUK1_1),.doutc(w_n695_0[2]),.din(n695));
	jspl3 jspl3_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.doutc(w_n699_0[2]),.din(n699));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_dff_A_Bq7f18HZ2_1),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_dff_A_Hkcjyptd3_1),.din(n709));
	jspl jspl_w_n710_0(.douta(w_dff_A_UVhmSwRi2_0),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_dff_A_vvtsNuvE8_0),.doutb(w_n711_0[1]),.din(n711));
	jspl3 jspl3_w_n713_0(.douta(w_n713_0[0]),.doutb(w_dff_A_fNtva72h0_1),.doutc(w_n713_0[2]),.din(n713));
	jspl3 jspl3_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.doutc(w_n715_0[2]),.din(n715));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(w_dff_B_HaW6KD374_2));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_dff_A_UnSMDFQx4_1),.din(n719));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_dff_A_qoh4vhNv1_1),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_dff_A_ysBaB5zn3_1),.din(n721));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_dff_A_dMeO5M2X8_1),.din(n722));
	jspl3 jspl3_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.doutc(w_n725_0[2]),.din(n725));
	jspl jspl_w_n726_0(.douta(w_dff_A_X7ZMSWaE8_0),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.doutc(w_n733_0[2]),.din(n733));
	jspl3 jspl3_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.doutc(w_n735_0[2]),.din(n735));
	jspl3 jspl3_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl jspl_w_n737_1(.douta(w_n737_1[0]),.doutb(w_n737_1[1]),.din(w_n737_0[0]));
	jspl jspl_w_n738_0(.douta(w_n738_0[0]),.doutb(w_n738_0[1]),.din(n738));
	jspl3 jspl3_w_n742_0(.douta(w_n742_0[0]),.doutb(w_dff_A_h2ENW0g59_1),.doutc(w_n742_0[2]),.din(n742));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_dff_A_AGM8M7Sv0_1),.doutc(w_n746_0[2]),.din(n746));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(w_dff_B_59QTf0HI5_2));
	jspl3 jspl3_w_n749_0(.douta(w_n749_0[0]),.doutb(w_dff_A_wjIhlaw92_1),.doutc(w_dff_A_UxkExz4G1_2),.din(n749));
	jspl3 jspl3_w_n749_1(.douta(w_n749_1[0]),.doutb(w_dff_A_XjrQOuP52_1),.doutc(w_dff_A_Dq9oZTdE6_2),.din(w_n749_0[0]));
	jspl3 jspl3_w_n749_2(.douta(w_dff_A_fScvVv0S0_0),.doutb(w_dff_A_NtPI2eCN5_1),.doutc(w_n749_2[2]),.din(w_n749_0[1]));
	jspl3 jspl3_w_n749_3(.douta(w_dff_A_sGjd8nTr1_0),.doutb(w_n749_3[1]),.doutc(w_dff_A_K6riXqK07_2),.din(w_n749_0[2]));
	jspl3 jspl3_w_n749_4(.douta(w_n749_4[0]),.doutb(w_dff_A_BR90ggWF7_1),.doutc(w_dff_A_l3hale7f1_2),.din(w_n749_1[0]));
	jspl3 jspl3_w_n749_5(.douta(w_dff_A_2mXuuQ4Y2_0),.doutb(w_dff_A_0Z3Tn8FY6_1),.doutc(w_n749_5[2]),.din(w_n749_1[1]));
	jspl3 jspl3_w_n749_6(.douta(w_dff_A_9QojdME74_0),.doutb(w_n749_6[1]),.doutc(w_n749_6[2]),.din(w_n749_1[2]));
	jspl3 jspl3_w_n749_7(.douta(w_dff_A_7x2yeONB8_0),.doutb(w_n749_7[1]),.doutc(w_n749_7[2]),.din(w_n749_2[0]));
	jspl3 jspl3_w_n749_8(.douta(w_n749_8[0]),.doutb(w_dff_A_dIDY0ASi7_1),.doutc(w_dff_A_tTXFHE0C8_2),.din(w_n749_2[1]));
	jspl3 jspl3_w_n749_9(.douta(w_dff_A_Xjp4Fyrw4_0),.doutb(w_n749_9[1]),.doutc(w_dff_A_4cKtydrZ2_2),.din(w_n749_2[2]));
	jspl3 jspl3_w_n749_10(.douta(w_n749_10[0]),.doutb(w_n749_10[1]),.doutc(w_n749_10[2]),.din(w_n749_3[0]));
	jspl3 jspl3_w_n749_11(.douta(w_dff_A_YBRV6JoW0_0),.doutb(w_dff_A_wmEkHaAt4_1),.doutc(w_n749_11[2]),.din(w_n749_3[1]));
	jspl3 jspl3_w_n749_12(.douta(w_n749_12[0]),.doutb(w_n749_12[1]),.doutc(w_n749_12[2]),.din(w_n749_3[2]));
	jspl jspl_w_n749_13(.douta(w_dff_A_xnnPnaiM2_0),.doutb(w_n749_13[1]),.din(w_n749_4[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.doutc(w_n750_0[2]),.din(n750));
	jspl3 jspl3_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.doutc(w_n750_1[2]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n750_2(.douta(w_n750_2[0]),.doutb(w_n750_2[1]),.doutc(w_n750_2[2]),.din(w_n750_0[1]));
	jspl3 jspl3_w_n750_3(.douta(w_n750_3[0]),.doutb(w_n750_3[1]),.doutc(w_n750_3[2]),.din(w_n750_0[2]));
	jspl3 jspl3_w_n750_4(.douta(w_n750_4[0]),.doutb(w_n750_4[1]),.doutc(w_n750_4[2]),.din(w_n750_1[0]));
	jspl3 jspl3_w_n750_5(.douta(w_n750_5[0]),.doutb(w_n750_5[1]),.doutc(w_n750_5[2]),.din(w_n750_1[1]));
	jspl3 jspl3_w_n750_6(.douta(w_n750_6[0]),.doutb(w_n750_6[1]),.doutc(w_n750_6[2]),.din(w_n750_1[2]));
	jspl3 jspl3_w_n750_7(.douta(w_n750_7[0]),.doutb(w_n750_7[1]),.doutc(w_n750_7[2]),.din(w_n750_2[0]));
	jspl3 jspl3_w_n750_8(.douta(w_n750_8[0]),.doutb(w_n750_8[1]),.doutc(w_n750_8[2]),.din(w_n750_2[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_dff_A_butyZvEC9_1),.doutc(w_dff_A_wBk3dmqZ4_2),.din(w_dff_B_CabbYQKU6_3));
	jspl jspl_w_n753_1(.douta(w_dff_A_OFptFf4R2_0),.doutb(w_n753_1[1]),.din(w_n753_0[0]));
	jspl jspl_w_n755_0(.douta(w_dff_A_YzDgD4NE9_0),.doutb(w_n755_0[1]),.din(n755));
	jspl3 jspl3_w_n763_0(.douta(w_dff_A_pxtAKnMq3_0),.doutb(w_n763_0[1]),.doutc(w_n763_0[2]),.din(n763));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl jspl_w_n779_0(.douta(w_dff_A_QmtQyr2u7_0),.doutb(w_n779_0[1]),.din(n779));
	jspl3 jspl3_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.doutc(w_n786_0[2]),.din(n786));
	jspl3 jspl3_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.doutc(w_n788_0[2]),.din(n788));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_dff_A_VwbmPG1e6_1),.doutc(w_n790_0[2]),.din(n790));
	jspl3 jspl3_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.doutc(w_dff_A_H7atk1yL6_2),.din(n792));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_n797_1[1]),.doutc(w_n797_1[2]),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_n797_2[2]),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_dff_A_wZ31z6lw8_0),.doutb(w_n797_3[1]),.doutc(w_n797_3[2]),.din(w_n797_0[2]));
	jspl3 jspl3_w_n797_4(.douta(w_dff_A_0PAbTmFU7_0),.doutb(w_n797_4[1]),.doutc(w_dff_A_qOvYg6Ov9_2),.din(w_n797_1[0]));
	jspl3 jspl3_w_n797_5(.douta(w_n797_5[0]),.doutb(w_dff_A_bxqxQOu92_1),.doutc(w_n797_5[2]),.din(w_n797_1[1]));
	jspl3 jspl3_w_n797_6(.douta(w_dff_A_e2azE1u77_0),.doutb(w_n797_6[1]),.doutc(w_dff_A_yraG014I1_2),.din(w_n797_1[2]));
	jspl3 jspl3_w_n797_7(.douta(w_n797_7[0]),.doutb(w_dff_A_ktRA898b1_1),.doutc(w_n797_7[2]),.din(w_n797_2[0]));
	jspl3 jspl3_w_n797_8(.douta(w_dff_A_WkEANbXK0_0),.doutb(w_n797_8[1]),.doutc(w_dff_A_DhSM3jhv1_2),.din(w_n797_2[1]));
	jspl jspl_w_n797_9(.douta(w_n797_9[0]),.doutb(w_dff_A_jwufuSU28_1),.din(w_n797_2[2]));
	jspl3 jspl3_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.doutc(w_n798_0[2]),.din(n798));
	jspl jspl_w_n798_1(.douta(w_n798_1[0]),.doutb(w_n798_1[1]),.din(w_n798_0[0]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_dff_A_a9eq3c733_1),.doutc(w_dff_A_aolLGTMm4_2),.din(w_dff_B_x66oaevu3_3));
	jspl3 jspl3_w_n800_1(.douta(w_n800_1[0]),.doutb(w_dff_A_twRL69CU3_1),.doutc(w_dff_A_llbMoU9z6_2),.din(w_n800_0[0]));
	jspl3 jspl3_w_n800_2(.douta(w_n800_2[0]),.doutb(w_n800_2[1]),.doutc(w_dff_A_F6kEEoLb0_2),.din(w_n800_0[1]));
	jspl3 jspl3_w_n800_3(.douta(w_dff_A_nbDlv0sp1_0),.doutb(w_n800_3[1]),.doutc(w_dff_A_LYsHmIKq1_2),.din(w_n800_0[2]));
	jspl jspl_w_n800_4(.douta(w_dff_A_7SbTxlr39_0),.doutb(w_n800_4[1]),.din(w_n800_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl jspl_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n814_0(.douta(w_dff_A_ci6v7xUY3_0),.doutb(w_dff_A_qUeNlPd81_1),.doutc(w_n814_0[2]),.din(n814));
	jspl3 jspl3_w_n819_0(.douta(w_n819_0[0]),.doutb(w_dff_A_hZ5D2cD50_1),.doutc(w_n819_0[2]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_dff_A_iSB1yla53_1),.din(n821));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n836_0(.douta(w_dff_A_hFWOoDh04_0),.doutb(w_n836_0[1]),.din(n836));
	jspl jspl_w_n847_0(.douta(w_dff_A_QodupDsy5_0),.doutb(w_n847_0[1]),.din(n847));
	jspl3 jspl3_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.doutc(w_n852_0[2]),.din(n852));
	jspl3 jspl3_w_n852_1(.douta(w_n852_1[0]),.doutb(w_n852_1[1]),.doutc(w_n852_1[2]),.din(w_n852_0[0]));
	jspl3 jspl3_w_n852_2(.douta(w_n852_2[0]),.doutb(w_n852_2[1]),.doutc(w_n852_2[2]),.din(w_n852_0[1]));
	jspl3 jspl3_w_n852_3(.douta(w_dff_A_9DvEUrSW2_0),.doutb(w_n852_3[1]),.doutc(w_n852_3[2]),.din(w_n852_0[2]));
	jspl3 jspl3_w_n852_4(.douta(w_dff_A_fxyaCb5N2_0),.doutb(w_n852_4[1]),.doutc(w_dff_A_HFOfGJ697_2),.din(w_n852_1[0]));
	jspl3 jspl3_w_n852_5(.douta(w_n852_5[0]),.doutb(w_dff_A_bn9BiymC4_1),.doutc(w_dff_A_l7yjVuJE0_2),.din(w_n852_1[1]));
	jspl3 jspl3_w_n852_6(.douta(w_n852_6[0]),.doutb(w_n852_6[1]),.doutc(w_dff_A_KgpDjXJt6_2),.din(w_n852_1[2]));
	jspl3 jspl3_w_n852_7(.douta(w_dff_A_VSekOTg48_0),.doutb(w_n852_7[1]),.doutc(w_dff_A_gQ0ePflD6_2),.din(w_n852_2[0]));
	jspl3 jspl3_w_n852_8(.douta(w_n852_8[0]),.doutb(w_dff_A_fbZ2eGkt8_1),.doutc(w_n852_8[2]),.din(w_n852_2[1]));
	jspl jspl_w_n852_9(.douta(w_n852_9[0]),.doutb(w_dff_A_nQHq9kuD5_1),.din(w_n852_2[2]));
	jspl3 jspl3_w_n854_0(.douta(w_n854_0[0]),.doutb(w_dff_A_M28Bwhdm8_1),.doutc(w_dff_A_sm2eBv348_2),.din(w_dff_B_x6sYVZQl0_3));
	jspl3 jspl3_w_n854_1(.douta(w_n854_1[0]),.doutb(w_dff_A_VXwxUIU01_1),.doutc(w_dff_A_nkBS7BN47_2),.din(w_n854_0[0]));
	jspl3 jspl3_w_n854_2(.douta(w_n854_2[0]),.doutb(w_n854_2[1]),.doutc(w_n854_2[2]),.din(w_n854_0[1]));
	jspl3 jspl3_w_n854_3(.douta(w_n854_3[0]),.doutb(w_n854_3[1]),.doutc(w_dff_A_tfvNvX5W5_2),.din(w_n854_0[2]));
	jspl jspl_w_n854_4(.douta(w_dff_A_Y9uM1MYt2_0),.doutb(w_n854_4[1]),.din(w_n854_1[0]));
	jspl3 jspl3_w_n865_0(.douta(w_dff_A_PPDwXgPR8_0),.doutb(w_n865_0[1]),.doutc(w_dff_A_oJqkeyL69_2),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n868_0(.douta(w_n868_0[0]),.doutb(w_n868_0[1]),.din(n868));
	jspl jspl_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.din(n870));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl jspl_w_n880_0(.douta(w_dff_A_UqfCelNO3_0),.doutb(w_n880_0[1]),.din(n880));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(n890));
	jspl jspl_w_n901_0(.douta(w_dff_A_S3xNVy6Y3_0),.doutb(w_n901_0[1]),.din(n901));
	jspl3 jspl3_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.doutc(w_n923_0[2]),.din(n923));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl3 jspl3_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.doutc(w_dff_A_BN6ZpJxo8_2),.din(n938));
	jspl3 jspl3_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.doutc(w_n940_0[2]),.din(n940));
	jspl jspl_w_n940_1(.douta(w_n940_1[0]),.doutb(w_n940_1[1]),.din(w_n940_0[0]));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(n944));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_dff_A_DN6DoIr47_1),.din(n949));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl3 jspl3_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.doutc(w_dff_A_ccdkAcaE8_2),.din(n954));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_dff_A_m7ftWT6w2_1),.din(w_dff_B_85atRmAC4_2));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl3 jspl3_w_n977_0(.douta(w_n977_0[0]),.doutb(w_n977_0[1]),.doutc(w_n977_0[2]),.din(n977));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_dff_A_NWcfJXEZ4_1),.din(n989));
	jspl3 jspl3_w_n993_0(.douta(w_n993_0[0]),.doutb(w_dff_A_yLxDTtHx7_1),.doutc(w_dff_A_7HUVL1Pp0_2),.din(n993));
	jspl3 jspl3_w_n993_1(.douta(w_n993_1[0]),.doutb(w_dff_A_4fDZu6Ro7_1),.doutc(w_dff_A_0ShZnwgW3_2),.din(w_n993_0[0]));
	jspl3 jspl3_w_n993_2(.douta(w_dff_A_UJV9MCdP1_0),.doutb(w_dff_A_LZMJYExx1_1),.doutc(w_n993_2[2]),.din(w_n993_0[1]));
	jspl3 jspl3_w_n993_3(.douta(w_dff_A_IhOTjENe3_0),.doutb(w_dff_A_qCkbwAAw0_1),.doutc(w_n993_3[2]),.din(w_n993_0[2]));
	jspl3 jspl3_w_n993_4(.douta(w_dff_A_RiCzsvby6_0),.doutb(w_dff_A_svDBm8Jc3_1),.doutc(w_n993_4[2]),.din(w_n993_1[0]));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n994_1(.douta(w_n994_1[0]),.doutb(w_n994_1[1]),.doutc(w_n994_1[2]),.din(w_n994_0[0]));
	jspl3 jspl3_w_n994_2(.douta(w_n994_2[0]),.doutb(w_n994_2[1]),.doutc(w_n994_2[2]),.din(w_n994_0[1]));
	jspl3 jspl3_w_n994_3(.douta(w_n994_3[0]),.doutb(w_n994_3[1]),.doutc(w_n994_3[2]),.din(w_n994_0[2]));
	jspl jspl_w_n994_4(.douta(w_n994_4[0]),.doutb(w_n994_4[1]),.din(w_n994_1[0]));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl3 jspl3_w_n996_1(.douta(w_n996_1[0]),.doutb(w_n996_1[1]),.doutc(w_n996_1[2]),.din(w_n996_0[0]));
	jspl3 jspl3_w_n996_2(.douta(w_n996_2[0]),.doutb(w_n996_2[1]),.doutc(w_n996_2[2]),.din(w_n996_0[1]));
	jspl3 jspl3_w_n996_3(.douta(w_n996_3[0]),.doutb(w_n996_3[1]),.doutc(w_n996_3[2]),.din(w_n996_0[2]));
	jspl jspl_w_n996_4(.douta(w_n996_4[0]),.doutb(w_n996_4[1]),.din(w_n996_1[0]));
	jspl3 jspl3_w_n999_0(.douta(w_dff_A_icU0pCwP7_0),.doutb(w_dff_A_aU4vB9mg4_1),.doutc(w_n999_0[2]),.din(w_dff_B_p5mSOc3W6_3));
	jspl3 jspl3_w_n999_1(.douta(w_dff_A_lDSczqec3_0),.doutb(w_dff_A_50ph0ZCE3_1),.doutc(w_n999_1[2]),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_dff_A_ofsuAHg40_0),.doutb(w_dff_A_BCdCY5Bq5_1),.doutc(w_n999_2[2]),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_dff_A_iItlQ5sG3_0),.doutb(w_dff_A_CZiGEFGF6_1),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl3 jspl3_w_n1007_0(.douta(w_dff_A_UbutgT4e4_0),.doutb(w_dff_A_xDJ80oeC7_1),.doutc(w_n1007_0[2]),.din(w_dff_B_Oqq6t7dM4_3));
	jspl3 jspl3_w_n1007_1(.douta(w_n1007_1[0]),.doutb(w_n1007_1[1]),.doutc(w_dff_A_DhcTfbY66_2),.din(w_n1007_0[0]));
	jspl3 jspl3_w_n1007_2(.douta(w_dff_A_aQU1CCTB6_0),.doutb(w_dff_A_VvUbhN3i4_1),.doutc(w_n1007_2[2]),.din(w_n1007_0[1]));
	jspl3 jspl3_w_n1007_3(.douta(w_dff_A_jx8wBfJg7_0),.doutb(w_dff_A_0UNvS99k5_1),.doutc(w_n1007_3[2]),.din(w_n1007_0[2]));
	jspl3 jspl3_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_dff_A_pkIOg8DR5_1),.doutc(w_dff_A_d18Xh9zG0_2),.din(n1008));
	jspl3 jspl3_w_n1008_1(.douta(w_n1008_1[0]),.doutb(w_dff_A_nvVPJzbg4_1),.doutc(w_dff_A_zLTOu8JK5_2),.din(w_n1008_0[0]));
	jspl3 jspl3_w_n1008_2(.douta(w_dff_A_gg4BFt0t4_0),.doutb(w_dff_A_4itjFJvj8_1),.doutc(w_n1008_2[2]),.din(w_n1008_0[1]));
	jspl3 jspl3_w_n1008_3(.douta(w_dff_A_KBPGaox53_0),.doutb(w_dff_A_7kP6WV9w4_1),.doutc(w_n1008_3[2]),.din(w_n1008_0[2]));
	jspl3 jspl3_w_n1008_4(.douta(w_dff_A_9DaxWcVe5_0),.doutb(w_n1008_4[1]),.doutc(w_dff_A_wdof90BC0_2),.din(w_n1008_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl3 jspl3_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.doutc(w_n1012_1[2]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1012_2(.douta(w_n1012_2[0]),.doutb(w_n1012_2[1]),.doutc(w_n1012_2[2]),.din(w_n1012_0[1]));
	jspl3 jspl3_w_n1012_3(.douta(w_n1012_3[0]),.doutb(w_n1012_3[1]),.doutc(w_n1012_3[2]),.din(w_n1012_0[2]));
	jspl jspl_w_n1012_4(.douta(w_n1012_4[0]),.doutb(w_n1012_4[1]),.din(w_n1012_1[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl3 jspl3_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.doutc(w_n1014_1[2]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1014_2(.douta(w_n1014_2[0]),.doutb(w_n1014_2[1]),.doutc(w_n1014_2[2]),.din(w_n1014_0[1]));
	jspl3 jspl3_w_n1014_3(.douta(w_n1014_3[0]),.doutb(w_n1014_3[1]),.doutc(w_n1014_3[2]),.din(w_n1014_0[2]));
	jspl jspl_w_n1014_4(.douta(w_n1014_4[0]),.doutb(w_n1014_4[1]),.din(w_n1014_1[0]));
	jspl3 jspl3_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.doutc(w_n1019_0[2]),.din(n1019));
	jspl jspl_w_n1019_1(.douta(w_n1019_1[0]),.doutb(w_n1019_1[1]),.din(w_n1019_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl3 jspl3_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.doutc(w_n1043_0[2]),.din(n1043));
	jspl jspl_w_n1043_1(.douta(w_n1043_1[0]),.doutb(w_n1043_1[1]),.din(w_n1043_0[0]));
	jspl3 jspl3_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.doutc(w_n1052_0[2]),.din(n1052));
	jspl jspl_w_n1052_1(.douta(w_n1052_1[0]),.doutb(w_n1052_1[1]),.din(w_n1052_0[0]));
	jspl3 jspl3_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.doutc(w_n1054_0[2]),.din(n1054));
	jspl jspl_w_n1054_1(.douta(w_n1054_1[0]),.doutb(w_n1054_1[1]),.din(w_n1054_0[0]));
	jspl jspl_w_n1177_0(.douta(w_dff_A_64TXrpuB7_0),.doutb(w_n1177_0[1]),.din(w_dff_B_504jPPon2_2));
	jspl jspl_w_n1179_0(.douta(w_dff_A_5GDr8oCN8_0),.doutb(w_n1179_0[1]),.din(n1179));
	jspl3 jspl3_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.doutc(w_n1196_0[2]),.din(n1196));
	jspl3 jspl3_w_n1196_1(.douta(w_n1196_1[0]),.doutb(w_n1196_1[1]),.doutc(w_n1196_1[2]),.din(w_n1196_0[0]));
	jspl3 jspl3_w_n1201_0(.douta(w_dff_A_9yjaLKeD7_0),.doutb(w_dff_A_t9wquEM91_1),.doutc(w_n1201_0[2]),.din(w_dff_B_6JI8y1nQ3_3));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.doutc(w_n1213_0[2]),.din(n1213));
	jspl3 jspl3_w_n1213_1(.douta(w_n1213_1[0]),.doutb(w_n1213_1[1]),.doutc(w_n1213_1[2]),.din(w_n1213_0[0]));
	jspl3 jspl3_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.doutc(w_n1236_0[2]),.din(n1236));
	jspl3 jspl3_w_n1236_1(.douta(w_n1236_1[0]),.doutb(w_n1236_1[1]),.doutc(w_n1236_1[2]),.din(w_n1236_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl3 jspl3_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.doutc(w_n1251_1[2]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.doutc(w_n1279_0[2]),.din(n1279));
	jspl jspl_w_n1279_1(.douta(w_n1279_1[0]),.doutb(w_n1279_1[1]),.din(w_n1279_0[0]));
	jspl3 jspl3_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.doutc(w_n1297_0[2]),.din(n1297));
	jspl jspl_w_n1297_1(.douta(w_n1297_1[0]),.doutb(w_n1297_1[1]),.din(w_n1297_0[0]));
	jspl3 jspl3_w_n1299_0(.douta(w_n1299_0[0]),.doutb(w_n1299_0[1]),.doutc(w_n1299_0[2]),.din(n1299));
	jspl jspl_w_n1299_1(.douta(w_n1299_1[0]),.doutb(w_n1299_1[1]),.din(w_n1299_0[0]));
	jspl3 jspl3_w_n1410_0(.douta(w_dff_A_FPsJvK3N9_0),.doutb(w_n1410_0[1]),.doutc(w_n1410_0[2]),.din(n1410));
	jspl3 jspl3_w_n1412_0(.douta(w_n1412_0[0]),.doutb(w_dff_A_gOqqgfa46_1),.doutc(w_dff_A_DisGo5P51_2),.din(w_dff_B_X9d1K3tK5_3));
	jspl jspl_w_n1416_0(.douta(w_n1416_0[0]),.doutb(w_n1416_0[1]),.din(n1416));
	jspl jspl_w_n1422_0(.douta(w_dff_A_pph0MgxZ3_0),.doutb(w_n1422_0[1]),.din(n1422));
	jspl jspl_w_n1425_0(.douta(w_dff_A_w7MUFPIP6_0),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(n1428));
	jspl jspl_w_n1429_0(.douta(w_dff_A_4tImIQIC6_0),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1451_0(.douta(w_dff_A_ABbQpe6u2_0),.doutb(w_n1451_0[1]),.din(n1451));
	jspl jspl_w_n1503_0(.douta(w_n1503_0[0]),.doutb(w_n1503_0[1]),.din(n1503));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1592_0(.douta(w_n1592_0[0]),.doutb(w_n1592_0[1]),.din(n1592));
	jspl jspl_w_n1593_0(.douta(w_n1593_0[0]),.doutb(w_n1593_0[1]),.din(n1593));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1599_0(.douta(w_dff_A_8aoAnBKr2_0),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_n1603_0[1]),.din(n1603));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl3 jspl3_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.doutc(w_n1611_0[2]),.din(n1611));
	jspl jspl_w_n1613_0(.douta(w_dff_A_FcJRNiM37_0),.doutb(w_n1613_0[1]),.din(n1613));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(n1615));
	jspl jspl_w_n1618_0(.douta(w_dff_A_pDMn4PWS6_0),.doutb(w_n1618_0[1]),.din(w_dff_B_r7JxUxaj9_2));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(w_dff_B_bA6fv7q99_2));
	jspl jspl_w_n1637_0(.douta(w_dff_A_ufo0E6sZ2_0),.doutb(w_n1637_0[1]),.din(w_dff_B_Y8KYvAO46_2));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(n1643));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_dff_A_P4SEEAWN6_1),.din(n1652));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl3 jspl3_w_n1674_0(.douta(w_n1674_0[0]),.doutb(w_n1674_0[1]),.doutc(w_n1674_0[2]),.din(n1674));
	jspl jspl_w_n1675_0(.douta(w_n1675_0[0]),.doutb(w_n1675_0[1]),.din(n1675));
	jspl3 jspl3_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.doutc(w_n1679_0[2]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(w_dff_B_njf0WG6e3_2));
	jspl jspl_w_n1695_0(.douta(w_n1695_0[0]),.doutb(w_n1695_0[1]),.din(w_dff_B_poQPHa3h8_2));
	jspl jspl_w_n1698_0(.douta(w_n1698_0[0]),.doutb(w_n1698_0[1]),.din(w_dff_B_dv0Sk1rx6_2));
	jdff dff_B_5pseY3ze5_1(.din(G136),.dout(w_dff_B_5pseY3ze5_1),.clk(gclk));
	jdff dff_B_5d0LIbSn2_0(.din(G2824),.dout(w_dff_B_5d0LIbSn2_0),.clk(gclk));
	jdff dff_B_gZLfCesE0_1(.din(n320),.dout(w_dff_B_gZLfCesE0_1),.clk(gclk));
	jdff dff_B_XXGaiOMy4_1(.din(n327),.dout(w_dff_B_XXGaiOMy4_1),.clk(gclk));
	jdff dff_B_uZZ3q6Nx0_2(.din(n333),.dout(w_dff_B_uZZ3q6Nx0_2),.clk(gclk));
	jdff dff_B_3l13xEUy4_1(.din(n338),.dout(w_dff_B_3l13xEUy4_1),.clk(gclk));
	jdff dff_B_uWMWTVN67_1(.din(n340),.dout(w_dff_B_uWMWTVN67_1),.clk(gclk));
	jdff dff_B_0UaRHFHX3_0(.din(n341),.dout(w_dff_B_0UaRHFHX3_0),.clk(gclk));
	jdff dff_B_1gs4QHJx1_1(.din(G24),.dout(w_dff_B_1gs4QHJx1_1),.clk(gclk));
	jdff dff_B_rtRIxOw27_1(.din(n345),.dout(w_dff_B_rtRIxOw27_1),.clk(gclk));
	jdff dff_B_fcKXeWTj0_0(.din(n346),.dout(w_dff_B_fcKXeWTj0_0),.clk(gclk));
	jdff dff_B_U8XNJdiR0_1(.din(G26),.dout(w_dff_B_U8XNJdiR0_1),.clk(gclk));
	jdff dff_A_QQ8poydE2_0(.dout(w_G141_2[0]),.din(w_dff_A_QQ8poydE2_0),.clk(gclk));
	jdff dff_A_Vom0CuN06_0(.dout(w_dff_A_QQ8poydE2_0),.din(w_dff_A_Vom0CuN06_0),.clk(gclk));
	jdff dff_A_nxHYnxi72_0(.dout(w_dff_A_Vom0CuN06_0),.din(w_dff_A_nxHYnxi72_0),.clk(gclk));
	jdff dff_A_QsBAZN6D1_0(.dout(w_dff_A_nxHYnxi72_0),.din(w_dff_A_QsBAZN6D1_0),.clk(gclk));
	jdff dff_A_p77QdkLy9_1(.dout(w_G141_2[1]),.din(w_dff_A_p77QdkLy9_1),.clk(gclk));
	jdff dff_A_XtZe12Jn2_1(.dout(w_dff_A_p77QdkLy9_1),.din(w_dff_A_XtZe12Jn2_1),.clk(gclk));
	jdff dff_A_nZjOPtI04_1(.dout(w_dff_A_XtZe12Jn2_1),.din(w_dff_A_nZjOPtI04_1),.clk(gclk));
	jdff dff_A_4zSc1LyP2_1(.dout(w_dff_A_nZjOPtI04_1),.din(w_dff_A_4zSc1LyP2_1),.clk(gclk));
	jdff dff_B_49CQMAWp8_1(.din(n350),.dout(w_dff_B_49CQMAWp8_1),.clk(gclk));
	jdff dff_B_mV6sOTPV5_0(.din(n351),.dout(w_dff_B_mV6sOTPV5_0),.clk(gclk));
	jdff dff_B_dxVJs3kJ3_1(.din(G79),.dout(w_dff_B_dxVJs3kJ3_1),.clk(gclk));
	jdff dff_B_JNlV6HdC8_1(.din(n355),.dout(w_dff_B_JNlV6HdC8_1),.clk(gclk));
	jdff dff_B_24q7TdUc7_1(.din(w_dff_B_JNlV6HdC8_1),.dout(w_dff_B_24q7TdUc7_1),.clk(gclk));
	jdff dff_B_TonoSrvx8_1(.din(G82),.dout(w_dff_B_TonoSrvx8_1),.clk(gclk));
	jdff dff_A_sfF8rck74_0(.dout(w_G2358_2[0]),.din(w_dff_A_sfF8rck74_0),.clk(gclk));
	jdff dff_A_LxfFmvmr5_1(.dout(w_G2358_2[1]),.din(w_dff_A_LxfFmvmr5_1),.clk(gclk));
	jdff dff_A_RnnwGZJ82_1(.dout(w_G141_1[1]),.din(w_dff_A_RnnwGZJ82_1),.clk(gclk));
	jdff dff_A_wf2fsBPP2_1(.dout(w_dff_A_RnnwGZJ82_1),.din(w_dff_A_wf2fsBPP2_1),.clk(gclk));
	jdff dff_A_x0BvDMD32_1(.dout(w_dff_A_wf2fsBPP2_1),.din(w_dff_A_x0BvDMD32_1),.clk(gclk));
	jdff dff_A_4zGRtotu7_1(.dout(w_dff_A_x0BvDMD32_1),.din(w_dff_A_4zGRtotu7_1),.clk(gclk));
	jdff dff_A_LO9HR7Du4_2(.dout(w_G141_1[2]),.din(w_dff_A_LO9HR7Du4_2),.clk(gclk));
	jdff dff_A_9sIB7H2L7_2(.dout(w_dff_A_LO9HR7Du4_2),.din(w_dff_A_9sIB7H2L7_2),.clk(gclk));
	jdff dff_A_LAtJFuWb8_2(.dout(w_dff_A_9sIB7H2L7_2),.din(w_dff_A_LAtJFuWb8_2),.clk(gclk));
	jdff dff_A_TccOO6vn9_2(.dout(w_dff_A_LAtJFuWb8_2),.din(w_dff_A_TccOO6vn9_2),.clk(gclk));
	jdff dff_B_JiQHGNmO2_1(.din(n373),.dout(w_dff_B_JiQHGNmO2_1),.clk(gclk));
	jdff dff_B_hKIdI6aE7_2(.din(n661),.dout(w_dff_B_hKIdI6aE7_2),.clk(gclk));
	jdff dff_B_fOGWVeyJ0_2(.din(w_dff_B_hKIdI6aE7_2),.dout(w_dff_B_fOGWVeyJ0_2),.clk(gclk));
	jdff dff_B_Apk4W4Cq7_2(.din(n717),.dout(w_dff_B_Apk4W4Cq7_2),.clk(gclk));
	jdff dff_B_HaW6KD374_2(.din(w_dff_B_Apk4W4Cq7_2),.dout(w_dff_B_HaW6KD374_2),.clk(gclk));
	jdff dff_B_5scfG8PG4_1(.din(n705),.dout(w_dff_B_5scfG8PG4_1),.clk(gclk));
	jdff dff_B_C0HkSu132_1(.din(w_dff_B_5scfG8PG4_1),.dout(w_dff_B_C0HkSu132_1),.clk(gclk));
	jdff dff_B_OtJkf61N6_1(.din(w_dff_B_C0HkSu132_1),.dout(w_dff_B_OtJkf61N6_1),.clk(gclk));
	jdff dff_B_lNqwqNLr0_1(.din(w_dff_B_OtJkf61N6_1),.dout(w_dff_B_lNqwqNLr0_1),.clk(gclk));
	jdff dff_B_t2G5m4Xl0_1(.din(w_dff_B_lNqwqNLr0_1),.dout(w_dff_B_t2G5m4Xl0_1),.clk(gclk));
	jdff dff_B_9A2iSTBK3_1(.din(w_dff_B_t2G5m4Xl0_1),.dout(w_dff_B_9A2iSTBK3_1),.clk(gclk));
	jdff dff_B_gcvUXHpN5_1(.din(n706),.dout(w_dff_B_gcvUXHpN5_1),.clk(gclk));
	jdff dff_B_dM0hsl3E7_1(.din(w_dff_B_gcvUXHpN5_1),.dout(w_dff_B_dM0hsl3E7_1),.clk(gclk));
	jdff dff_B_kovXpwa96_1(.din(w_dff_B_dM0hsl3E7_1),.dout(w_dff_B_kovXpwa96_1),.clk(gclk));
	jdff dff_B_v9eAHOge7_1(.din(w_dff_B_kovXpwa96_1),.dout(w_dff_B_v9eAHOge7_1),.clk(gclk));
	jdff dff_B_cb2UIZEQ3_1(.din(w_dff_B_v9eAHOge7_1),.dout(w_dff_B_cb2UIZEQ3_1),.clk(gclk));
	jdff dff_A_TBJLgtFH8_1(.dout(w_n611_0[1]),.din(w_dff_A_TBJLgtFH8_1),.clk(gclk));
	jdff dff_A_wK0ga2Vk4_1(.dout(w_dff_A_TBJLgtFH8_1),.din(w_dff_A_wK0ga2Vk4_1),.clk(gclk));
	jdff dff_B_Y78scTpD4_3(.din(n611),.dout(w_dff_B_Y78scTpD4_3),.clk(gclk));
	jdff dff_B_7f7BGebr2_2(.din(n747),.dout(w_dff_B_7f7BGebr2_2),.clk(gclk));
	jdff dff_B_59QTf0HI5_2(.din(w_dff_B_7f7BGebr2_2),.dout(w_dff_B_59QTf0HI5_2),.clk(gclk));
	jdff dff_B_ip4JU1t60_1(.din(n739),.dout(w_dff_B_ip4JU1t60_1),.clk(gclk));
	jdff dff_B_lgf4lBax9_1(.din(w_dff_B_ip4JU1t60_1),.dout(w_dff_B_lgf4lBax9_1),.clk(gclk));
	jdff dff_A_h1J2x2Ra4_0(.dout(w_n660_1[0]),.din(w_dff_A_h1J2x2Ra4_0),.clk(gclk));
	jdff dff_A_75yJteUV9_0(.dout(w_dff_A_h1J2x2Ra4_0),.din(w_dff_A_75yJteUV9_0),.clk(gclk));
	jdff dff_A_1nYH5uZI8_0(.dout(w_dff_A_75yJteUV9_0),.din(w_dff_A_1nYH5uZI8_0),.clk(gclk));
	jdff dff_A_szz1ylTx7_0(.dout(w_dff_A_1nYH5uZI8_0),.din(w_dff_A_szz1ylTx7_0),.clk(gclk));
	jdff dff_A_q7uSuu5a5_0(.dout(w_dff_A_szz1ylTx7_0),.din(w_dff_A_q7uSuu5a5_0),.clk(gclk));
	jdff dff_B_OW6jf2Sd3_0(.din(n808),.dout(w_dff_B_OW6jf2Sd3_0),.clk(gclk));
	jdff dff_B_WgOLK0H23_0(.din(w_dff_B_OW6jf2Sd3_0),.dout(w_dff_B_WgOLK0H23_0),.clk(gclk));
	jdff dff_B_cEH97czM1_0(.din(w_dff_B_WgOLK0H23_0),.dout(w_dff_B_cEH97czM1_0),.clk(gclk));
	jdff dff_B_dJCb12AO3_0(.din(w_dff_B_cEH97czM1_0),.dout(w_dff_B_dJCb12AO3_0),.clk(gclk));
	jdff dff_B_r7lcnJvL4_0(.din(w_dff_B_dJCb12AO3_0),.dout(w_dff_B_r7lcnJvL4_0),.clk(gclk));
	jdff dff_B_7vEWjXbf7_0(.din(w_dff_B_r7lcnJvL4_0),.dout(w_dff_B_7vEWjXbf7_0),.clk(gclk));
	jdff dff_B_pjcJhtvT5_0(.din(w_dff_B_7vEWjXbf7_0),.dout(w_dff_B_pjcJhtvT5_0),.clk(gclk));
	jdff dff_B_9Z1qVH0j7_0(.din(w_dff_B_pjcJhtvT5_0),.dout(w_dff_B_9Z1qVH0j7_0),.clk(gclk));
	jdff dff_B_aCMTOUZe0_0(.din(w_dff_B_9Z1qVH0j7_0),.dout(w_dff_B_aCMTOUZe0_0),.clk(gclk));
	jdff dff_B_YQx7uU1H6_0(.din(w_dff_B_aCMTOUZe0_0),.dout(w_dff_B_YQx7uU1H6_0),.clk(gclk));
	jdff dff_B_6UaTBp6x0_0(.din(n803),.dout(w_dff_B_6UaTBp6x0_0),.clk(gclk));
	jdff dff_A_yvkTFnJ01_1(.dout(w_n797_9[1]),.din(w_dff_A_yvkTFnJ01_1),.clk(gclk));
	jdff dff_A_QbrgWKe19_1(.dout(w_dff_A_yvkTFnJ01_1),.din(w_dff_A_QbrgWKe19_1),.clk(gclk));
	jdff dff_A_cRhSMklw6_1(.dout(w_dff_A_QbrgWKe19_1),.din(w_dff_A_cRhSMklw6_1),.clk(gclk));
	jdff dff_A_Hmk375zk1_1(.dout(w_dff_A_cRhSMklw6_1),.din(w_dff_A_Hmk375zk1_1),.clk(gclk));
	jdff dff_A_XS65W3Tb0_1(.dout(w_dff_A_Hmk375zk1_1),.din(w_dff_A_XS65W3Tb0_1),.clk(gclk));
	jdff dff_A_XLu2d7qV7_1(.dout(w_dff_A_XS65W3Tb0_1),.din(w_dff_A_XLu2d7qV7_1),.clk(gclk));
	jdff dff_A_ffpR4mWY8_1(.dout(w_dff_A_XLu2d7qV7_1),.din(w_dff_A_ffpR4mWY8_1),.clk(gclk));
	jdff dff_A_hfbZ9uG27_1(.dout(w_dff_A_ffpR4mWY8_1),.din(w_dff_A_hfbZ9uG27_1),.clk(gclk));
	jdff dff_A_NKHrKRDb4_1(.dout(w_dff_A_hfbZ9uG27_1),.din(w_dff_A_NKHrKRDb4_1),.clk(gclk));
	jdff dff_A_jwufuSU28_1(.dout(w_dff_A_NKHrKRDb4_1),.din(w_dff_A_jwufuSU28_1),.clk(gclk));
	jdff dff_B_dxadoulk7_0(.din(n861),.dout(w_dff_B_dxadoulk7_0),.clk(gclk));
	jdff dff_B_nflMTdIG9_0(.din(w_dff_B_dxadoulk7_0),.dout(w_dff_B_nflMTdIG9_0),.clk(gclk));
	jdff dff_B_xvDPDxmy0_0(.din(w_dff_B_nflMTdIG9_0),.dout(w_dff_B_xvDPDxmy0_0),.clk(gclk));
	jdff dff_B_o0ptTId29_0(.din(w_dff_B_xvDPDxmy0_0),.dout(w_dff_B_o0ptTId29_0),.clk(gclk));
	jdff dff_B_qOKjY7rs7_0(.din(w_dff_B_o0ptTId29_0),.dout(w_dff_B_qOKjY7rs7_0),.clk(gclk));
	jdff dff_B_yVBOucxr8_0(.din(w_dff_B_qOKjY7rs7_0),.dout(w_dff_B_yVBOucxr8_0),.clk(gclk));
	jdff dff_B_AYQD91Uo5_0(.din(w_dff_B_yVBOucxr8_0),.dout(w_dff_B_AYQD91Uo5_0),.clk(gclk));
	jdff dff_B_uhReZfBD9_0(.din(w_dff_B_AYQD91Uo5_0),.dout(w_dff_B_uhReZfBD9_0),.clk(gclk));
	jdff dff_B_adVclcQ96_0(.din(w_dff_B_uhReZfBD9_0),.dout(w_dff_B_adVclcQ96_0),.clk(gclk));
	jdff dff_B_9jj3DoR38_0(.din(w_dff_B_adVclcQ96_0),.dout(w_dff_B_9jj3DoR38_0),.clk(gclk));
	jdff dff_B_D334u1qO2_2(.din(G61),.dout(w_dff_B_D334u1qO2_2),.clk(gclk));
	jdff dff_B_0IFzQppa9_0(.din(n856),.dout(w_dff_B_0IFzQppa9_0),.clk(gclk));
	jdff dff_A_BM69SWUv2_1(.dout(w_n852_9[1]),.din(w_dff_A_BM69SWUv2_1),.clk(gclk));
	jdff dff_A_M8Q9Df9q4_1(.dout(w_dff_A_BM69SWUv2_1),.din(w_dff_A_M8Q9Df9q4_1),.clk(gclk));
	jdff dff_A_ASZC6nE61_1(.dout(w_dff_A_M8Q9Df9q4_1),.din(w_dff_A_ASZC6nE61_1),.clk(gclk));
	jdff dff_A_NASzT5FX1_1(.dout(w_dff_A_ASZC6nE61_1),.din(w_dff_A_NASzT5FX1_1),.clk(gclk));
	jdff dff_A_ATEQW8G72_1(.dout(w_dff_A_NASzT5FX1_1),.din(w_dff_A_ATEQW8G72_1),.clk(gclk));
	jdff dff_A_1GaqXvWj0_1(.dout(w_dff_A_ATEQW8G72_1),.din(w_dff_A_1GaqXvWj0_1),.clk(gclk));
	jdff dff_A_IvliJj7m2_1(.dout(w_dff_A_1GaqXvWj0_1),.din(w_dff_A_IvliJj7m2_1),.clk(gclk));
	jdff dff_A_1jJHwIJK8_1(.dout(w_dff_A_IvliJj7m2_1),.din(w_dff_A_1jJHwIJK8_1),.clk(gclk));
	jdff dff_A_4MVfoLgo8_1(.dout(w_dff_A_1jJHwIJK8_1),.din(w_dff_A_4MVfoLgo8_1),.clk(gclk));
	jdff dff_A_nQHq9kuD5_1(.dout(w_dff_A_4MVfoLgo8_1),.din(w_dff_A_nQHq9kuD5_1),.clk(gclk));
	jdff dff_B_QIMtgdLF5_0(.din(n967),.dout(w_dff_B_QIMtgdLF5_0),.clk(gclk));
	jdff dff_B_MCoew3nT4_1(.din(n961),.dout(w_dff_B_MCoew3nT4_1),.clk(gclk));
	jdff dff_B_KbbBnvZI2_1(.din(w_dff_B_MCoew3nT4_1),.dout(w_dff_B_KbbBnvZI2_1),.clk(gclk));
	jdff dff_B_RH5sCLMh0_1(.din(w_dff_B_KbbBnvZI2_1),.dout(w_dff_B_RH5sCLMh0_1),.clk(gclk));
	jdff dff_B_LNKh3xgB8_0(.din(n960),.dout(w_dff_B_LNKh3xgB8_0),.clk(gclk));
	jdff dff_B_MsSxupwE8_1(.din(n975),.dout(w_dff_B_MsSxupwE8_1),.clk(gclk));
	jdff dff_B_gwZZCsGf6_1(.din(w_dff_B_MsSxupwE8_1),.dout(w_dff_B_gwZZCsGf6_1),.clk(gclk));
	jdff dff_B_xUjzgfDb8_1(.din(w_dff_B_gwZZCsGf6_1),.dout(w_dff_B_xUjzgfDb8_1),.clk(gclk));
	jdff dff_B_AG9aNpSz3_1(.din(w_dff_B_xUjzgfDb8_1),.dout(w_dff_B_AG9aNpSz3_1),.clk(gclk));
	jdff dff_B_cA5UtwHA5_1(.din(w_dff_B_AG9aNpSz3_1),.dout(w_dff_B_cA5UtwHA5_1),.clk(gclk));
	jdff dff_B_hTywLHFX4_1(.din(n971),.dout(w_dff_B_hTywLHFX4_1),.clk(gclk));
	jdff dff_B_AUY7s4db5_1(.din(w_dff_B_hTywLHFX4_1),.dout(w_dff_B_AUY7s4db5_1),.clk(gclk));
	jdff dff_B_Qya5qyKF1_1(.din(n995),.dout(w_dff_B_Qya5qyKF1_1),.clk(gclk));
	jdff dff_B_EN9kUsYt2_1(.din(w_dff_B_Qya5qyKF1_1),.dout(w_dff_B_EN9kUsYt2_1),.clk(gclk));
	jdff dff_B_LGtJH1MA6_1(.din(w_dff_B_EN9kUsYt2_1),.dout(w_dff_B_LGtJH1MA6_1),.clk(gclk));
	jdff dff_B_rLse5twH7_1(.din(w_dff_B_LGtJH1MA6_1),.dout(w_dff_B_rLse5twH7_1),.clk(gclk));
	jdff dff_B_dyr2GmnC0_1(.din(w_dff_B_rLse5twH7_1),.dout(w_dff_B_dyr2GmnC0_1),.clk(gclk));
	jdff dff_B_QOBSfU5f1_1(.din(w_dff_B_dyr2GmnC0_1),.dout(w_dff_B_QOBSfU5f1_1),.clk(gclk));
	jdff dff_B_WGGjwLHl1_1(.din(w_dff_B_QOBSfU5f1_1),.dout(w_dff_B_WGGjwLHl1_1),.clk(gclk));
	jdff dff_B_oNDzFxhm3_1(.din(w_dff_B_WGGjwLHl1_1),.dout(w_dff_B_oNDzFxhm3_1),.clk(gclk));
	jdff dff_B_1dDUVuTi6_1(.din(w_dff_B_oNDzFxhm3_1),.dout(w_dff_B_1dDUVuTi6_1),.clk(gclk));
	jdff dff_B_Ynynngap4_1(.din(w_dff_B_1dDUVuTi6_1),.dout(w_dff_B_Ynynngap4_1),.clk(gclk));
	jdff dff_B_96gCK1kk3_1(.din(w_dff_B_Ynynngap4_1),.dout(w_dff_B_96gCK1kk3_1),.clk(gclk));
	jdff dff_B_Bj8SxTbY3_1(.din(n997),.dout(w_dff_B_Bj8SxTbY3_1),.clk(gclk));
	jdff dff_B_OHythTkV1_1(.din(w_dff_B_Bj8SxTbY3_1),.dout(w_dff_B_OHythTkV1_1),.clk(gclk));
	jdff dff_B_E5dUUKBX6_1(.din(w_dff_B_OHythTkV1_1),.dout(w_dff_B_E5dUUKBX6_1),.clk(gclk));
	jdff dff_B_SGWjoghx5_1(.din(w_dff_B_E5dUUKBX6_1),.dout(w_dff_B_SGWjoghx5_1),.clk(gclk));
	jdff dff_B_8CAnK0on1_1(.din(w_dff_B_SGWjoghx5_1),.dout(w_dff_B_8CAnK0on1_1),.clk(gclk));
	jdff dff_B_atnPbo0f4_1(.din(w_dff_B_8CAnK0on1_1),.dout(w_dff_B_atnPbo0f4_1),.clk(gclk));
	jdff dff_B_L1Ma3WVe6_1(.din(w_dff_B_atnPbo0f4_1),.dout(w_dff_B_L1Ma3WVe6_1),.clk(gclk));
	jdff dff_B_j6UYEdby3_1(.din(w_dff_B_L1Ma3WVe6_1),.dout(w_dff_B_j6UYEdby3_1),.clk(gclk));
	jdff dff_B_2ozp6x2H3_1(.din(w_dff_B_j6UYEdby3_1),.dout(w_dff_B_2ozp6x2H3_1),.clk(gclk));
	jdff dff_B_zHVZMFQC0_1(.din(w_dff_B_2ozp6x2H3_1),.dout(w_dff_B_zHVZMFQC0_1),.clk(gclk));
	jdff dff_B_wixnft3X6_1(.din(w_dff_B_zHVZMFQC0_1),.dout(w_dff_B_wixnft3X6_1),.clk(gclk));
	jdff dff_B_LB8GxHHJ9_0(.din(n1001),.dout(w_dff_B_LB8GxHHJ9_0),.clk(gclk));
	jdff dff_B_umFULM2S3_0(.din(n1016),.dout(w_dff_B_umFULM2S3_0),.clk(gclk));
	jdff dff_B_xcyEfhkz8_0(.din(w_dff_B_umFULM2S3_0),.dout(w_dff_B_xcyEfhkz8_0),.clk(gclk));
	jdff dff_B_IHGACzIj0_0(.din(w_dff_B_xcyEfhkz8_0),.dout(w_dff_B_IHGACzIj0_0),.clk(gclk));
	jdff dff_B_kshCvsy17_0(.din(w_dff_B_IHGACzIj0_0),.dout(w_dff_B_kshCvsy17_0),.clk(gclk));
	jdff dff_B_2T2lo8qZ5_0(.din(w_dff_B_kshCvsy17_0),.dout(w_dff_B_2T2lo8qZ5_0),.clk(gclk));
	jdff dff_B_iakkHnI28_0(.din(w_dff_B_2T2lo8qZ5_0),.dout(w_dff_B_iakkHnI28_0),.clk(gclk));
	jdff dff_B_pGe9HiPR0_0(.din(w_dff_B_iakkHnI28_0),.dout(w_dff_B_pGe9HiPR0_0),.clk(gclk));
	jdff dff_B_wnqpi1zG9_0(.din(w_dff_B_pGe9HiPR0_0),.dout(w_dff_B_wnqpi1zG9_0),.clk(gclk));
	jdff dff_B_dzUXXO4t5_0(.din(w_dff_B_wnqpi1zG9_0),.dout(w_dff_B_dzUXXO4t5_0),.clk(gclk));
	jdff dff_B_jYwc0CJA9_0(.din(w_dff_B_dzUXXO4t5_0),.dout(w_dff_B_jYwc0CJA9_0),.clk(gclk));
	jdff dff_B_Er9MKswT7_1(.din(n1013),.dout(w_dff_B_Er9MKswT7_1),.clk(gclk));
	jdff dff_B_QwwoiTRd0_2(.din(G182),.dout(w_dff_B_QwwoiTRd0_2),.clk(gclk));
	jdff dff_B_4NfCGkbl4_2(.din(w_dff_B_QwwoiTRd0_2),.dout(w_dff_B_4NfCGkbl4_2),.clk(gclk));
	jdff dff_B_eZ8BiIdW9_2(.din(G185),.dout(w_dff_B_eZ8BiIdW9_2),.clk(gclk));
	jdff dff_B_hG0UErfk8_1(.din(n1006),.dout(w_dff_B_hG0UErfk8_1),.clk(gclk));
	jdff dff_B_SaMigYhO5_1(.din(w_dff_B_hG0UErfk8_1),.dout(w_dff_B_SaMigYhO5_1),.clk(gclk));
	jdff dff_B_sObn9bEK3_1(.din(w_dff_B_SaMigYhO5_1),.dout(w_dff_B_sObn9bEK3_1),.clk(gclk));
	jdff dff_B_zUVC3qY25_1(.din(n777),.dout(w_dff_B_zUVC3qY25_1),.clk(gclk));
	jdff dff_B_tcmkMNDz8_1(.din(w_dff_B_zUVC3qY25_1),.dout(w_dff_B_tcmkMNDz8_1),.clk(gclk));
	jdff dff_B_n1ABL9mY3_1(.din(w_dff_B_tcmkMNDz8_1),.dout(w_dff_B_n1ABL9mY3_1),.clk(gclk));
	jdff dff_B_dyaOGlLv3_1(.din(w_dff_B_n1ABL9mY3_1),.dout(w_dff_B_dyaOGlLv3_1),.clk(gclk));
	jdff dff_B_8ZKG8dxr1_1(.din(w_dff_B_dyaOGlLv3_1),.dout(w_dff_B_8ZKG8dxr1_1),.clk(gclk));
	jdff dff_B_zK5ZTSk17_0(.din(n782),.dout(w_dff_B_zK5ZTSk17_0),.clk(gclk));
	jdff dff_B_QgSZRQ2D7_1(.din(n536),.dout(w_dff_B_QgSZRQ2D7_1),.clk(gclk));
	jdff dff_B_vfk6ABnv7_1(.din(n531),.dout(w_dff_B_vfk6ABnv7_1),.clk(gclk));
	jdff dff_A_rnixLMeT4_0(.dout(w_n779_0[0]),.din(w_dff_A_rnixLMeT4_0),.clk(gclk));
	jdff dff_A_QmtQyr2u7_0(.dout(w_dff_A_rnixLMeT4_0),.din(w_dff_A_QmtQyr2u7_0),.clk(gclk));
	jdff dff_B_fSWHe2016_1(.din(G117),.dout(w_dff_B_fSWHe2016_1),.clk(gclk));
	jdff dff_B_6cjba8ES8_1(.din(w_dff_B_fSWHe2016_1),.dout(w_dff_B_6cjba8ES8_1),.clk(gclk));
	jdff dff_B_412dZbzB8_1(.din(n752),.dout(w_dff_B_412dZbzB8_1),.clk(gclk));
	jdff dff_B_Evl6tKCs9_1(.din(w_dff_B_412dZbzB8_1),.dout(w_dff_B_Evl6tKCs9_1),.clk(gclk));
	jdff dff_B_9CjPmnQA1_1(.din(w_dff_B_Evl6tKCs9_1),.dout(w_dff_B_9CjPmnQA1_1),.clk(gclk));
	jdff dff_A_7iOJvDjX4_0(.dout(w_n755_0[0]),.din(w_dff_A_7iOJvDjX4_0),.clk(gclk));
	jdff dff_A_vRVddJJz5_0(.dout(w_dff_A_7iOJvDjX4_0),.din(w_dff_A_vRVddJJz5_0),.clk(gclk));
	jdff dff_A_CxBDqyPT0_0(.dout(w_dff_A_vRVddJJz5_0),.din(w_dff_A_CxBDqyPT0_0),.clk(gclk));
	jdff dff_A_jdCE27XT0_0(.dout(w_dff_A_CxBDqyPT0_0),.din(w_dff_A_jdCE27XT0_0),.clk(gclk));
	jdff dff_A_u4v0WMYu4_0(.dout(w_dff_A_jdCE27XT0_0),.din(w_dff_A_u4v0WMYu4_0),.clk(gclk));
	jdff dff_A_ZXn6SsW18_0(.dout(w_dff_A_u4v0WMYu4_0),.din(w_dff_A_ZXn6SsW18_0),.clk(gclk));
	jdff dff_A_HOGXNGNK0_0(.dout(w_dff_A_ZXn6SsW18_0),.din(w_dff_A_HOGXNGNK0_0),.clk(gclk));
	jdff dff_A_jeVpKP5m4_0(.dout(w_dff_A_HOGXNGNK0_0),.din(w_dff_A_jeVpKP5m4_0),.clk(gclk));
	jdff dff_A_AVD6DKrQ3_0(.dout(w_dff_A_jeVpKP5m4_0),.din(w_dff_A_AVD6DKrQ3_0),.clk(gclk));
	jdff dff_A_XotcTJEI5_0(.dout(w_dff_A_AVD6DKrQ3_0),.din(w_dff_A_XotcTJEI5_0),.clk(gclk));
	jdff dff_A_YzDgD4NE9_0(.dout(w_dff_A_XotcTJEI5_0),.din(w_dff_A_YzDgD4NE9_0),.clk(gclk));
	jdff dff_B_tNxFShYp2_1(.din(G131),.dout(w_dff_B_tNxFShYp2_1),.clk(gclk));
	jdff dff_B_QCr6Roxr9_1(.din(w_dff_B_tNxFShYp2_1),.dout(w_dff_B_QCr6Roxr9_1),.clk(gclk));
	jdff dff_B_hem3m85J9_0(.din(n1028),.dout(w_dff_B_hem3m85J9_0),.clk(gclk));
	jdff dff_B_jB9kaDXI6_0(.din(w_dff_B_hem3m85J9_0),.dout(w_dff_B_jB9kaDXI6_0),.clk(gclk));
	jdff dff_B_imStMAos3_0(.din(w_dff_B_jB9kaDXI6_0),.dout(w_dff_B_imStMAos3_0),.clk(gclk));
	jdff dff_B_qpRosqnp9_0(.din(w_dff_B_imStMAos3_0),.dout(w_dff_B_qpRosqnp9_0),.clk(gclk));
	jdff dff_B_lPeYGUcP2_0(.din(w_dff_B_qpRosqnp9_0),.dout(w_dff_B_lPeYGUcP2_0),.clk(gclk));
	jdff dff_B_xLM2x2TL0_0(.din(w_dff_B_lPeYGUcP2_0),.dout(w_dff_B_xLM2x2TL0_0),.clk(gclk));
	jdff dff_B_afLguixQ7_0(.din(w_dff_B_xLM2x2TL0_0),.dout(w_dff_B_afLguixQ7_0),.clk(gclk));
	jdff dff_B_J8SFRSD43_0(.din(w_dff_B_afLguixQ7_0),.dout(w_dff_B_J8SFRSD43_0),.clk(gclk));
	jdff dff_B_TWNIPGHf4_0(.din(w_dff_B_J8SFRSD43_0),.dout(w_dff_B_TWNIPGHf4_0),.clk(gclk));
	jdff dff_B_G0CDObb12_0(.din(w_dff_B_TWNIPGHf4_0),.dout(w_dff_B_G0CDObb12_0),.clk(gclk));
	jdff dff_B_6GrgtVyM6_0(.din(w_dff_B_G0CDObb12_0),.dout(w_dff_B_6GrgtVyM6_0),.clk(gclk));
	jdff dff_B_Lb0MexbC2_0(.din(w_dff_B_6GrgtVyM6_0),.dout(w_dff_B_Lb0MexbC2_0),.clk(gclk));
	jdff dff_B_Yw796fOH8_0(.din(w_dff_B_Lb0MexbC2_0),.dout(w_dff_B_Yw796fOH8_0),.clk(gclk));
	jdff dff_B_DUIetwC06_0(.din(w_dff_B_Yw796fOH8_0),.dout(w_dff_B_DUIetwC06_0),.clk(gclk));
	jdff dff_B_sfwCod1Y0_0(.din(w_dff_B_DUIetwC06_0),.dout(w_dff_B_sfwCod1Y0_0),.clk(gclk));
	jdff dff_B_XbfJ5Bvn5_0(.din(w_dff_B_sfwCod1Y0_0),.dout(w_dff_B_XbfJ5Bvn5_0),.clk(gclk));
	jdff dff_B_0j02iMEa7_1(.din(n1020),.dout(w_dff_B_0j02iMEa7_1),.clk(gclk));
	jdff dff_A_vdnHW2mK9_0(.dout(w_n800_4[0]),.din(w_dff_A_vdnHW2mK9_0),.clk(gclk));
	jdff dff_A_CNfTMicX7_0(.dout(w_dff_A_vdnHW2mK9_0),.din(w_dff_A_CNfTMicX7_0),.clk(gclk));
	jdff dff_A_DiHdsEXo0_0(.dout(w_dff_A_CNfTMicX7_0),.din(w_dff_A_DiHdsEXo0_0),.clk(gclk));
	jdff dff_A_eCkujpTU6_0(.dout(w_dff_A_DiHdsEXo0_0),.din(w_dff_A_eCkujpTU6_0),.clk(gclk));
	jdff dff_A_KOlomuab5_0(.dout(w_dff_A_eCkujpTU6_0),.din(w_dff_A_KOlomuab5_0),.clk(gclk));
	jdff dff_A_HjnkrWBB2_0(.dout(w_dff_A_KOlomuab5_0),.din(w_dff_A_HjnkrWBB2_0),.clk(gclk));
	jdff dff_A_7SbTxlr39_0(.dout(w_dff_A_HjnkrWBB2_0),.din(w_dff_A_7SbTxlr39_0),.clk(gclk));
	jdff dff_B_aZnhjJwS1_0(.din(n1039),.dout(w_dff_B_aZnhjJwS1_0),.clk(gclk));
	jdff dff_B_HGXdE1JU2_0(.din(w_dff_B_aZnhjJwS1_0),.dout(w_dff_B_HGXdE1JU2_0),.clk(gclk));
	jdff dff_B_wbHK1kru7_0(.din(w_dff_B_HGXdE1JU2_0),.dout(w_dff_B_wbHK1kru7_0),.clk(gclk));
	jdff dff_B_1ORWIEv39_0(.din(w_dff_B_wbHK1kru7_0),.dout(w_dff_B_1ORWIEv39_0),.clk(gclk));
	jdff dff_B_whN8cBP94_0(.din(w_dff_B_1ORWIEv39_0),.dout(w_dff_B_whN8cBP94_0),.clk(gclk));
	jdff dff_B_JmR7KTY56_0(.din(w_dff_B_whN8cBP94_0),.dout(w_dff_B_JmR7KTY56_0),.clk(gclk));
	jdff dff_B_Xzul8GGG7_0(.din(w_dff_B_JmR7KTY56_0),.dout(w_dff_B_Xzul8GGG7_0),.clk(gclk));
	jdff dff_B_ezuhTk814_0(.din(w_dff_B_Xzul8GGG7_0),.dout(w_dff_B_ezuhTk814_0),.clk(gclk));
	jdff dff_B_dnpunXcO3_0(.din(w_dff_B_ezuhTk814_0),.dout(w_dff_B_dnpunXcO3_0),.clk(gclk));
	jdff dff_B_xCa9bdv23_0(.din(w_dff_B_dnpunXcO3_0),.dout(w_dff_B_xCa9bdv23_0),.clk(gclk));
	jdff dff_B_kQjoGtDh7_0(.din(w_dff_B_xCa9bdv23_0),.dout(w_dff_B_kQjoGtDh7_0),.clk(gclk));
	jdff dff_B_EO0LESZg7_0(.din(w_dff_B_kQjoGtDh7_0),.dout(w_dff_B_EO0LESZg7_0),.clk(gclk));
	jdff dff_B_8LpmW8yO4_0(.din(w_dff_B_EO0LESZg7_0),.dout(w_dff_B_8LpmW8yO4_0),.clk(gclk));
	jdff dff_B_CE7e9NrA5_0(.din(w_dff_B_8LpmW8yO4_0),.dout(w_dff_B_CE7e9NrA5_0),.clk(gclk));
	jdff dff_B_MzogfC1j1_0(.din(w_dff_B_CE7e9NrA5_0),.dout(w_dff_B_MzogfC1j1_0),.clk(gclk));
	jdff dff_B_ewZDUYYX1_1(.din(n1031),.dout(w_dff_B_ewZDUYYX1_1),.clk(gclk));
	jdff dff_B_Hp4BtsS16_1(.din(w_dff_B_ewZDUYYX1_1),.dout(w_dff_B_Hp4BtsS16_1),.clk(gclk));
	jdff dff_A_1SidvPKG3_0(.dout(w_G4088_8[0]),.din(w_dff_A_1SidvPKG3_0),.clk(gclk));
	jdff dff_A_gQlOEQWk7_0(.dout(w_dff_A_1SidvPKG3_0),.din(w_dff_A_gQlOEQWk7_0),.clk(gclk));
	jdff dff_A_FoGlKVWx7_0(.dout(w_dff_A_gQlOEQWk7_0),.din(w_dff_A_FoGlKVWx7_0),.clk(gclk));
	jdff dff_A_VSuBAylf6_0(.dout(w_dff_A_FoGlKVWx7_0),.din(w_dff_A_VSuBAylf6_0),.clk(gclk));
	jdff dff_A_9Pp4vPt31_0(.dout(w_dff_A_VSuBAylf6_0),.din(w_dff_A_9Pp4vPt31_0),.clk(gclk));
	jdff dff_A_fweZvjD31_0(.dout(w_dff_A_9Pp4vPt31_0),.din(w_dff_A_fweZvjD31_0),.clk(gclk));
	jdff dff_A_qZRtGKRU3_0(.dout(w_dff_A_fweZvjD31_0),.din(w_dff_A_qZRtGKRU3_0),.clk(gclk));
	jdff dff_A_MuP6YyT31_0(.dout(w_dff_A_qZRtGKRU3_0),.din(w_dff_A_MuP6YyT31_0),.clk(gclk));
	jdff dff_A_pP6kBUgi0_0(.dout(w_dff_A_MuP6YyT31_0),.din(w_dff_A_pP6kBUgi0_0),.clk(gclk));
	jdff dff_A_EEv23slt9_0(.dout(w_dff_A_pP6kBUgi0_0),.din(w_dff_A_EEv23slt9_0),.clk(gclk));
	jdff dff_A_ok7JKiik8_0(.dout(w_dff_A_EEv23slt9_0),.din(w_dff_A_ok7JKiik8_0),.clk(gclk));
	jdff dff_A_Jftb7nTX1_0(.dout(w_dff_A_ok7JKiik8_0),.din(w_dff_A_Jftb7nTX1_0),.clk(gclk));
	jdff dff_A_m5XKEMfx7_0(.dout(w_dff_A_Jftb7nTX1_0),.din(w_dff_A_m5XKEMfx7_0),.clk(gclk));
	jdff dff_A_JjJ0bDPt0_0(.dout(w_dff_A_m5XKEMfx7_0),.din(w_dff_A_JjJ0bDPt0_0),.clk(gclk));
	jdff dff_A_neKuS7Eu8_0(.dout(w_dff_A_JjJ0bDPt0_0),.din(w_dff_A_neKuS7Eu8_0),.clk(gclk));
	jdff dff_A_9iDDQStT0_2(.dout(w_G4088_8[2]),.din(w_dff_A_9iDDQStT0_2),.clk(gclk));
	jdff dff_A_aaEC14nC7_2(.dout(w_dff_A_9iDDQStT0_2),.din(w_dff_A_aaEC14nC7_2),.clk(gclk));
	jdff dff_A_zWgHIMGW7_2(.dout(w_dff_A_aaEC14nC7_2),.din(w_dff_A_zWgHIMGW7_2),.clk(gclk));
	jdff dff_A_LPEzXf2q2_2(.dout(w_dff_A_zWgHIMGW7_2),.din(w_dff_A_LPEzXf2q2_2),.clk(gclk));
	jdff dff_A_jAa0sGrV2_2(.dout(w_dff_A_LPEzXf2q2_2),.din(w_dff_A_jAa0sGrV2_2),.clk(gclk));
	jdff dff_A_KdxEX8AO0_2(.dout(w_dff_A_jAa0sGrV2_2),.din(w_dff_A_KdxEX8AO0_2),.clk(gclk));
	jdff dff_A_XHQqgWwY6_2(.dout(w_dff_A_KdxEX8AO0_2),.din(w_dff_A_XHQqgWwY6_2),.clk(gclk));
	jdff dff_A_fpgmwc9O5_2(.dout(w_dff_A_XHQqgWwY6_2),.din(w_dff_A_fpgmwc9O5_2),.clk(gclk));
	jdff dff_A_xEIdpfM55_2(.dout(w_dff_A_fpgmwc9O5_2),.din(w_dff_A_xEIdpfM55_2),.clk(gclk));
	jdff dff_A_rjsII0Je5_2(.dout(w_dff_A_xEIdpfM55_2),.din(w_dff_A_rjsII0Je5_2),.clk(gclk));
	jdff dff_A_MOpea18H8_2(.dout(w_dff_A_rjsII0Je5_2),.din(w_dff_A_MOpea18H8_2),.clk(gclk));
	jdff dff_A_oe67f4Qu4_2(.dout(w_dff_A_MOpea18H8_2),.din(w_dff_A_oe67f4Qu4_2),.clk(gclk));
	jdff dff_A_01MzUA0w5_2(.dout(w_dff_A_oe67f4Qu4_2),.din(w_dff_A_01MzUA0w5_2),.clk(gclk));
	jdff dff_A_jNCimEpT6_2(.dout(w_dff_A_01MzUA0w5_2),.din(w_dff_A_jNCimEpT6_2),.clk(gclk));
	jdff dff_A_3ssK2ygp8_2(.dout(w_dff_A_jNCimEpT6_2),.din(w_dff_A_3ssK2ygp8_2),.clk(gclk));
	jdff dff_A_zDaWfg2a1_2(.dout(w_dff_A_3ssK2ygp8_2),.din(w_dff_A_zDaWfg2a1_2),.clk(gclk));
	jdff dff_A_ZAGSIkLI4_0(.dout(w_n797_8[0]),.din(w_dff_A_ZAGSIkLI4_0),.clk(gclk));
	jdff dff_A_v4x7lXO91_0(.dout(w_dff_A_ZAGSIkLI4_0),.din(w_dff_A_v4x7lXO91_0),.clk(gclk));
	jdff dff_A_FdnfLvON5_0(.dout(w_dff_A_v4x7lXO91_0),.din(w_dff_A_FdnfLvON5_0),.clk(gclk));
	jdff dff_A_CpOhPon59_0(.dout(w_dff_A_FdnfLvON5_0),.din(w_dff_A_CpOhPon59_0),.clk(gclk));
	jdff dff_A_Qfb5vhqN4_0(.dout(w_dff_A_CpOhPon59_0),.din(w_dff_A_Qfb5vhqN4_0),.clk(gclk));
	jdff dff_A_gEPDidKX5_0(.dout(w_dff_A_Qfb5vhqN4_0),.din(w_dff_A_gEPDidKX5_0),.clk(gclk));
	jdff dff_A_Ppaf1Vnl2_0(.dout(w_dff_A_gEPDidKX5_0),.din(w_dff_A_Ppaf1Vnl2_0),.clk(gclk));
	jdff dff_A_jeZCQKRq0_0(.dout(w_dff_A_Ppaf1Vnl2_0),.din(w_dff_A_jeZCQKRq0_0),.clk(gclk));
	jdff dff_A_6QQgHyQG6_0(.dout(w_dff_A_jeZCQKRq0_0),.din(w_dff_A_6QQgHyQG6_0),.clk(gclk));
	jdff dff_A_ZqnhYi1e2_0(.dout(w_dff_A_6QQgHyQG6_0),.din(w_dff_A_ZqnhYi1e2_0),.clk(gclk));
	jdff dff_A_mwdqPnKb4_0(.dout(w_dff_A_ZqnhYi1e2_0),.din(w_dff_A_mwdqPnKb4_0),.clk(gclk));
	jdff dff_A_bKBLcDTV3_0(.dout(w_dff_A_mwdqPnKb4_0),.din(w_dff_A_bKBLcDTV3_0),.clk(gclk));
	jdff dff_A_WkEANbXK0_0(.dout(w_dff_A_bKBLcDTV3_0),.din(w_dff_A_WkEANbXK0_0),.clk(gclk));
	jdff dff_A_ou2QQ6fy9_2(.dout(w_n797_8[2]),.din(w_dff_A_ou2QQ6fy9_2),.clk(gclk));
	jdff dff_A_c5Dp73J89_2(.dout(w_dff_A_ou2QQ6fy9_2),.din(w_dff_A_c5Dp73J89_2),.clk(gclk));
	jdff dff_A_Hix2Sr1j7_2(.dout(w_dff_A_c5Dp73J89_2),.din(w_dff_A_Hix2Sr1j7_2),.clk(gclk));
	jdff dff_A_RlbRqm319_2(.dout(w_dff_A_Hix2Sr1j7_2),.din(w_dff_A_RlbRqm319_2),.clk(gclk));
	jdff dff_A_SIXkhWH32_2(.dout(w_dff_A_RlbRqm319_2),.din(w_dff_A_SIXkhWH32_2),.clk(gclk));
	jdff dff_A_kOVtR4pq6_2(.dout(w_dff_A_SIXkhWH32_2),.din(w_dff_A_kOVtR4pq6_2),.clk(gclk));
	jdff dff_A_REWzpq9E4_2(.dout(w_dff_A_kOVtR4pq6_2),.din(w_dff_A_REWzpq9E4_2),.clk(gclk));
	jdff dff_A_UlP05Wkw8_2(.dout(w_dff_A_REWzpq9E4_2),.din(w_dff_A_UlP05Wkw8_2),.clk(gclk));
	jdff dff_A_RGWDA76O5_2(.dout(w_dff_A_UlP05Wkw8_2),.din(w_dff_A_RGWDA76O5_2),.clk(gclk));
	jdff dff_A_HrUtZ42O6_2(.dout(w_dff_A_RGWDA76O5_2),.din(w_dff_A_HrUtZ42O6_2),.clk(gclk));
	jdff dff_A_7vAGRxiF9_2(.dout(w_dff_A_HrUtZ42O6_2),.din(w_dff_A_7vAGRxiF9_2),.clk(gclk));
	jdff dff_A_PThipe6u7_2(.dout(w_dff_A_7vAGRxiF9_2),.din(w_dff_A_PThipe6u7_2),.clk(gclk));
	jdff dff_A_ydXySLI27_2(.dout(w_dff_A_PThipe6u7_2),.din(w_dff_A_ydXySLI27_2),.clk(gclk));
	jdff dff_A_dpNgruTi0_2(.dout(w_dff_A_ydXySLI27_2),.din(w_dff_A_dpNgruTi0_2),.clk(gclk));
	jdff dff_A_DhSM3jhv1_2(.dout(w_dff_A_dpNgruTi0_2),.din(w_dff_A_DhSM3jhv1_2),.clk(gclk));
	jdff dff_B_PpPZ4mCF7_0(.din(n1050),.dout(w_dff_B_PpPZ4mCF7_0),.clk(gclk));
	jdff dff_B_buytFbIi2_0(.din(w_dff_B_PpPZ4mCF7_0),.dout(w_dff_B_buytFbIi2_0),.clk(gclk));
	jdff dff_B_SUfuZQEe8_0(.din(w_dff_B_buytFbIi2_0),.dout(w_dff_B_SUfuZQEe8_0),.clk(gclk));
	jdff dff_B_d4GLyjtf2_0(.din(w_dff_B_SUfuZQEe8_0),.dout(w_dff_B_d4GLyjtf2_0),.clk(gclk));
	jdff dff_B_crnmLoxB9_0(.din(w_dff_B_d4GLyjtf2_0),.dout(w_dff_B_crnmLoxB9_0),.clk(gclk));
	jdff dff_B_Zv9QWa687_0(.din(w_dff_B_crnmLoxB9_0),.dout(w_dff_B_Zv9QWa687_0),.clk(gclk));
	jdff dff_B_SnANx2NB0_0(.din(w_dff_B_Zv9QWa687_0),.dout(w_dff_B_SnANx2NB0_0),.clk(gclk));
	jdff dff_B_mhTozrtV2_0(.din(w_dff_B_SnANx2NB0_0),.dout(w_dff_B_mhTozrtV2_0),.clk(gclk));
	jdff dff_B_dsIZujJ90_0(.din(w_dff_B_mhTozrtV2_0),.dout(w_dff_B_dsIZujJ90_0),.clk(gclk));
	jdff dff_B_xhMl4xgP7_0(.din(w_dff_B_dsIZujJ90_0),.dout(w_dff_B_xhMl4xgP7_0),.clk(gclk));
	jdff dff_B_mkGZjtUB5_0(.din(w_dff_B_xhMl4xgP7_0),.dout(w_dff_B_mkGZjtUB5_0),.clk(gclk));
	jdff dff_B_3nORkulA1_0(.din(w_dff_B_mkGZjtUB5_0),.dout(w_dff_B_3nORkulA1_0),.clk(gclk));
	jdff dff_B_Yerqif9U3_0(.din(w_dff_B_3nORkulA1_0),.dout(w_dff_B_Yerqif9U3_0),.clk(gclk));
	jdff dff_B_GSF4OTTx6_1(.din(n1042),.dout(w_dff_B_GSF4OTTx6_1),.clk(gclk));
	jdff dff_A_n29bVcSe6_1(.dout(w_n797_7[1]),.din(w_dff_A_n29bVcSe6_1),.clk(gclk));
	jdff dff_A_bJHrf9zj4_1(.dout(w_dff_A_n29bVcSe6_1),.din(w_dff_A_bJHrf9zj4_1),.clk(gclk));
	jdff dff_A_bXIbCL2N4_1(.dout(w_dff_A_bJHrf9zj4_1),.din(w_dff_A_bXIbCL2N4_1),.clk(gclk));
	jdff dff_A_PnZuGu2T4_1(.dout(w_dff_A_bXIbCL2N4_1),.din(w_dff_A_PnZuGu2T4_1),.clk(gclk));
	jdff dff_A_puB3p0UK8_1(.dout(w_dff_A_PnZuGu2T4_1),.din(w_dff_A_puB3p0UK8_1),.clk(gclk));
	jdff dff_A_g03S2BFt7_1(.dout(w_dff_A_puB3p0UK8_1),.din(w_dff_A_g03S2BFt7_1),.clk(gclk));
	jdff dff_A_m6QhEtQX8_1(.dout(w_dff_A_g03S2BFt7_1),.din(w_dff_A_m6QhEtQX8_1),.clk(gclk));
	jdff dff_A_zmH8t6tw7_1(.dout(w_dff_A_m6QhEtQX8_1),.din(w_dff_A_zmH8t6tw7_1),.clk(gclk));
	jdff dff_A_B5ruK8Uz3_1(.dout(w_dff_A_zmH8t6tw7_1),.din(w_dff_A_B5ruK8Uz3_1),.clk(gclk));
	jdff dff_A_fxnPmKbg2_1(.dout(w_dff_A_B5ruK8Uz3_1),.din(w_dff_A_fxnPmKbg2_1),.clk(gclk));
	jdff dff_A_VFQbVcPE5_1(.dout(w_dff_A_fxnPmKbg2_1),.din(w_dff_A_VFQbVcPE5_1),.clk(gclk));
	jdff dff_A_ktRA898b1_1(.dout(w_dff_A_VFQbVcPE5_1),.din(w_dff_A_ktRA898b1_1),.clk(gclk));
	jdff dff_A_axkdoY4Q0_1(.dout(w_G4088_7[1]),.din(w_dff_A_axkdoY4Q0_1),.clk(gclk));
	jdff dff_A_7M0IHwGm2_1(.dout(w_dff_A_axkdoY4Q0_1),.din(w_dff_A_7M0IHwGm2_1),.clk(gclk));
	jdff dff_A_bxoWGViU6_1(.dout(w_dff_A_7M0IHwGm2_1),.din(w_dff_A_bxoWGViU6_1),.clk(gclk));
	jdff dff_A_01JYIkab4_1(.dout(w_dff_A_bxoWGViU6_1),.din(w_dff_A_01JYIkab4_1),.clk(gclk));
	jdff dff_A_UUIxNnyx7_1(.dout(w_dff_A_01JYIkab4_1),.din(w_dff_A_UUIxNnyx7_1),.clk(gclk));
	jdff dff_A_gvF91yLG1_1(.dout(w_dff_A_UUIxNnyx7_1),.din(w_dff_A_gvF91yLG1_1),.clk(gclk));
	jdff dff_A_veiMbtOw5_1(.dout(w_dff_A_gvF91yLG1_1),.din(w_dff_A_veiMbtOw5_1),.clk(gclk));
	jdff dff_A_wBADW5Wd7_1(.dout(w_dff_A_veiMbtOw5_1),.din(w_dff_A_wBADW5Wd7_1),.clk(gclk));
	jdff dff_A_n1dyIVjz4_1(.dout(w_dff_A_wBADW5Wd7_1),.din(w_dff_A_n1dyIVjz4_1),.clk(gclk));
	jdff dff_A_25f27IqB4_1(.dout(w_dff_A_n1dyIVjz4_1),.din(w_dff_A_25f27IqB4_1),.clk(gclk));
	jdff dff_A_c8QfGWm31_1(.dout(w_dff_A_25f27IqB4_1),.din(w_dff_A_c8QfGWm31_1),.clk(gclk));
	jdff dff_A_9sSALoD26_1(.dout(w_dff_A_c8QfGWm31_1),.din(w_dff_A_9sSALoD26_1),.clk(gclk));
	jdff dff_A_SGXCpmyO5_1(.dout(w_dff_A_9sSALoD26_1),.din(w_dff_A_SGXCpmyO5_1),.clk(gclk));
	jdff dff_B_dYn8RS1x1_0(.din(n1061),.dout(w_dff_B_dYn8RS1x1_0),.clk(gclk));
	jdff dff_B_lH2NefW04_0(.din(w_dff_B_dYn8RS1x1_0),.dout(w_dff_B_lH2NefW04_0),.clk(gclk));
	jdff dff_B_eQRB0NKi3_0(.din(w_dff_B_lH2NefW04_0),.dout(w_dff_B_eQRB0NKi3_0),.clk(gclk));
	jdff dff_B_wsr3lvtj0_0(.din(w_dff_B_eQRB0NKi3_0),.dout(w_dff_B_wsr3lvtj0_0),.clk(gclk));
	jdff dff_B_rTMxEox44_0(.din(w_dff_B_wsr3lvtj0_0),.dout(w_dff_B_rTMxEox44_0),.clk(gclk));
	jdff dff_B_rAXi5MGZ2_0(.din(w_dff_B_rTMxEox44_0),.dout(w_dff_B_rAXi5MGZ2_0),.clk(gclk));
	jdff dff_B_f3Ordk8G1_0(.din(w_dff_B_rAXi5MGZ2_0),.dout(w_dff_B_f3Ordk8G1_0),.clk(gclk));
	jdff dff_B_4cf75ATx5_0(.din(w_dff_B_f3Ordk8G1_0),.dout(w_dff_B_4cf75ATx5_0),.clk(gclk));
	jdff dff_B_qtS4LE9L9_0(.din(w_dff_B_4cf75ATx5_0),.dout(w_dff_B_qtS4LE9L9_0),.clk(gclk));
	jdff dff_B_6e6VC4629_0(.din(w_dff_B_qtS4LE9L9_0),.dout(w_dff_B_6e6VC4629_0),.clk(gclk));
	jdff dff_B_1bNeTI3B4_0(.din(w_dff_B_6e6VC4629_0),.dout(w_dff_B_1bNeTI3B4_0),.clk(gclk));
	jdff dff_B_cmGXKS7h8_0(.din(w_dff_B_1bNeTI3B4_0),.dout(w_dff_B_cmGXKS7h8_0),.clk(gclk));
	jdff dff_B_2ufFjAIS4_0(.din(w_dff_B_cmGXKS7h8_0),.dout(w_dff_B_2ufFjAIS4_0),.clk(gclk));
	jdff dff_B_NXlOkNV54_0(.din(w_dff_B_2ufFjAIS4_0),.dout(w_dff_B_NXlOkNV54_0),.clk(gclk));
	jdff dff_B_Vs09V1U34_1(.din(n1053),.dout(w_dff_B_Vs09V1U34_1),.clk(gclk));
	jdff dff_B_OVdatxwx6_1(.din(w_dff_B_Vs09V1U34_1),.dout(w_dff_B_OVdatxwx6_1),.clk(gclk));
	jdff dff_B_XPkTXUtv3_1(.din(w_dff_B_OVdatxwx6_1),.dout(w_dff_B_XPkTXUtv3_1),.clk(gclk));
	jdff dff_A_nbDlv0sp1_0(.dout(w_n800_3[0]),.din(w_dff_A_nbDlv0sp1_0),.clk(gclk));
	jdff dff_A_UWVHTOkT5_2(.dout(w_n800_3[2]),.din(w_dff_A_UWVHTOkT5_2),.clk(gclk));
	jdff dff_A_LYsHmIKq1_2(.dout(w_dff_A_UWVHTOkT5_2),.din(w_dff_A_LYsHmIKq1_2),.clk(gclk));
	jdff dff_B_Vok9Jdl50_1(.din(n1066),.dout(w_dff_B_Vok9Jdl50_1),.clk(gclk));
	jdff dff_B_pbBmfKE70_1(.din(w_dff_B_Vok9Jdl50_1),.dout(w_dff_B_pbBmfKE70_1),.clk(gclk));
	jdff dff_B_cm38cG3f5_1(.din(w_dff_B_pbBmfKE70_1),.dout(w_dff_B_cm38cG3f5_1),.clk(gclk));
	jdff dff_B_VnpyObGo1_1(.din(w_dff_B_cm38cG3f5_1),.dout(w_dff_B_VnpyObGo1_1),.clk(gclk));
	jdff dff_B_PCmAm8xV7_1(.din(w_dff_B_VnpyObGo1_1),.dout(w_dff_B_PCmAm8xV7_1),.clk(gclk));
	jdff dff_B_RPERlSfS4_1(.din(w_dff_B_PCmAm8xV7_1),.dout(w_dff_B_RPERlSfS4_1),.clk(gclk));
	jdff dff_B_wlMOJKNq7_1(.din(w_dff_B_RPERlSfS4_1),.dout(w_dff_B_wlMOJKNq7_1),.clk(gclk));
	jdff dff_B_GSrExPpn2_1(.din(w_dff_B_wlMOJKNq7_1),.dout(w_dff_B_GSrExPpn2_1),.clk(gclk));
	jdff dff_B_fmHxdKZr7_1(.din(w_dff_B_GSrExPpn2_1),.dout(w_dff_B_fmHxdKZr7_1),.clk(gclk));
	jdff dff_B_TpOQrr2C8_1(.din(w_dff_B_fmHxdKZr7_1),.dout(w_dff_B_TpOQrr2C8_1),.clk(gclk));
	jdff dff_B_XXZ18Gv14_1(.din(w_dff_B_TpOQrr2C8_1),.dout(w_dff_B_XXZ18Gv14_1),.clk(gclk));
	jdff dff_B_WXInNCAx2_1(.din(w_dff_B_XXZ18Gv14_1),.dout(w_dff_B_WXInNCAx2_1),.clk(gclk));
	jdff dff_B_shGYiVLn1_1(.din(w_dff_B_WXInNCAx2_1),.dout(w_dff_B_shGYiVLn1_1),.clk(gclk));
	jdff dff_B_WBzlmFzL0_1(.din(w_dff_B_shGYiVLn1_1),.dout(w_dff_B_WBzlmFzL0_1),.clk(gclk));
	jdff dff_B_IZm3Gvzd0_1(.din(w_dff_B_WBzlmFzL0_1),.dout(w_dff_B_IZm3Gvzd0_1),.clk(gclk));
	jdff dff_A_VW3jl7Ex2_0(.dout(w_n854_4[0]),.din(w_dff_A_VW3jl7Ex2_0),.clk(gclk));
	jdff dff_A_79Oez01Q9_0(.dout(w_dff_A_VW3jl7Ex2_0),.din(w_dff_A_79Oez01Q9_0),.clk(gclk));
	jdff dff_A_D2NTLLU55_0(.dout(w_dff_A_79Oez01Q9_0),.din(w_dff_A_D2NTLLU55_0),.clk(gclk));
	jdff dff_A_eYo1lnmW7_0(.dout(w_dff_A_D2NTLLU55_0),.din(w_dff_A_eYo1lnmW7_0),.clk(gclk));
	jdff dff_A_6JZNvong7_0(.dout(w_dff_A_eYo1lnmW7_0),.din(w_dff_A_6JZNvong7_0),.clk(gclk));
	jdff dff_A_CiWSb2bP5_0(.dout(w_dff_A_6JZNvong7_0),.din(w_dff_A_CiWSb2bP5_0),.clk(gclk));
	jdff dff_A_1AhnXBIo2_0(.dout(w_dff_A_CiWSb2bP5_0),.din(w_dff_A_1AhnXBIo2_0),.clk(gclk));
	jdff dff_A_Y9uM1MYt2_0(.dout(w_dff_A_1AhnXBIo2_0),.din(w_dff_A_Y9uM1MYt2_0),.clk(gclk));
	jdff dff_B_7alQrAGz6_1(.din(n1063),.dout(w_dff_B_7alQrAGz6_1),.clk(gclk));
	jdff dff_B_JwnPyo986_1(.din(w_dff_B_7alQrAGz6_1),.dout(w_dff_B_JwnPyo986_1),.clk(gclk));
	jdff dff_B_lHCNbdw67_2(.din(G37),.dout(w_dff_B_lHCNbdw67_2),.clk(gclk));
	jdff dff_B_Or7ieCL40_1(.din(n1075),.dout(w_dff_B_Or7ieCL40_1),.clk(gclk));
	jdff dff_B_jyW51YLO6_1(.din(w_dff_B_Or7ieCL40_1),.dout(w_dff_B_jyW51YLO6_1),.clk(gclk));
	jdff dff_B_Ti1HaDSO1_1(.din(w_dff_B_jyW51YLO6_1),.dout(w_dff_B_Ti1HaDSO1_1),.clk(gclk));
	jdff dff_B_VK6F6Gs06_1(.din(w_dff_B_Ti1HaDSO1_1),.dout(w_dff_B_VK6F6Gs06_1),.clk(gclk));
	jdff dff_B_LqmTnlO72_1(.din(w_dff_B_VK6F6Gs06_1),.dout(w_dff_B_LqmTnlO72_1),.clk(gclk));
	jdff dff_B_6kmkD8AC8_1(.din(w_dff_B_LqmTnlO72_1),.dout(w_dff_B_6kmkD8AC8_1),.clk(gclk));
	jdff dff_B_n506kiGD5_1(.din(w_dff_B_6kmkD8AC8_1),.dout(w_dff_B_n506kiGD5_1),.clk(gclk));
	jdff dff_B_xL2ZF1gM3_1(.din(w_dff_B_n506kiGD5_1),.dout(w_dff_B_xL2ZF1gM3_1),.clk(gclk));
	jdff dff_B_ZH1SJDAf2_1(.din(w_dff_B_xL2ZF1gM3_1),.dout(w_dff_B_ZH1SJDAf2_1),.clk(gclk));
	jdff dff_B_dpwT5ush0_1(.din(w_dff_B_ZH1SJDAf2_1),.dout(w_dff_B_dpwT5ush0_1),.clk(gclk));
	jdff dff_B_uu52JJP23_1(.din(w_dff_B_dpwT5ush0_1),.dout(w_dff_B_uu52JJP23_1),.clk(gclk));
	jdff dff_B_ke0txx4M7_1(.din(w_dff_B_uu52JJP23_1),.dout(w_dff_B_ke0txx4M7_1),.clk(gclk));
	jdff dff_B_BaNWfyXH9_1(.din(w_dff_B_ke0txx4M7_1),.dout(w_dff_B_BaNWfyXH9_1),.clk(gclk));
	jdff dff_B_3PqhCcif5_1(.din(w_dff_B_BaNWfyXH9_1),.dout(w_dff_B_3PqhCcif5_1),.clk(gclk));
	jdff dff_B_OTTsIfBA1_0(.din(n1077),.dout(w_dff_B_OTTsIfBA1_0),.clk(gclk));
	jdff dff_B_O6sgrkC04_1(.din(n1072),.dout(w_dff_B_O6sgrkC04_1),.clk(gclk));
	jdff dff_B_z2wmbyYC3_1(.din(w_dff_B_O6sgrkC04_1),.dout(w_dff_B_z2wmbyYC3_1),.clk(gclk));
	jdff dff_A_6ugtbfPB3_1(.dout(w_n852_8[1]),.din(w_dff_A_6ugtbfPB3_1),.clk(gclk));
	jdff dff_A_oh1lAM2o7_1(.dout(w_dff_A_6ugtbfPB3_1),.din(w_dff_A_oh1lAM2o7_1),.clk(gclk));
	jdff dff_A_u3l2NVtL2_1(.dout(w_dff_A_oh1lAM2o7_1),.din(w_dff_A_u3l2NVtL2_1),.clk(gclk));
	jdff dff_A_s6fVlPWS9_1(.dout(w_dff_A_u3l2NVtL2_1),.din(w_dff_A_s6fVlPWS9_1),.clk(gclk));
	jdff dff_A_qweThpfB5_1(.dout(w_dff_A_s6fVlPWS9_1),.din(w_dff_A_qweThpfB5_1),.clk(gclk));
	jdff dff_A_OU2kOwBn0_1(.dout(w_dff_A_qweThpfB5_1),.din(w_dff_A_OU2kOwBn0_1),.clk(gclk));
	jdff dff_A_zPAMdFSs7_1(.dout(w_dff_A_OU2kOwBn0_1),.din(w_dff_A_zPAMdFSs7_1),.clk(gclk));
	jdff dff_A_yCh42Enh1_1(.dout(w_dff_A_zPAMdFSs7_1),.din(w_dff_A_yCh42Enh1_1),.clk(gclk));
	jdff dff_A_gdzIDZF52_1(.dout(w_dff_A_yCh42Enh1_1),.din(w_dff_A_gdzIDZF52_1),.clk(gclk));
	jdff dff_A_mTP01M8b7_1(.dout(w_dff_A_gdzIDZF52_1),.din(w_dff_A_mTP01M8b7_1),.clk(gclk));
	jdff dff_A_hwpktazI0_1(.dout(w_dff_A_mTP01M8b7_1),.din(w_dff_A_hwpktazI0_1),.clk(gclk));
	jdff dff_A_bEnidND31_1(.dout(w_dff_A_hwpktazI0_1),.din(w_dff_A_bEnidND31_1),.clk(gclk));
	jdff dff_A_wMdmBG4W9_1(.dout(w_dff_A_bEnidND31_1),.din(w_dff_A_wMdmBG4W9_1),.clk(gclk));
	jdff dff_A_PgdRUJlY1_1(.dout(w_dff_A_wMdmBG4W9_1),.din(w_dff_A_PgdRUJlY1_1),.clk(gclk));
	jdff dff_A_fbZ2eGkt8_1(.dout(w_dff_A_PgdRUJlY1_1),.din(w_dff_A_fbZ2eGkt8_1),.clk(gclk));
	jdff dff_B_2S5587Jz0_2(.din(G20),.dout(w_dff_B_2S5587Jz0_2),.clk(gclk));
	jdff dff_A_z3IMOOoq7_1(.dout(w_G4089_8[1]),.din(w_dff_A_z3IMOOoq7_1),.clk(gclk));
	jdff dff_A_a4w9YAAH5_1(.dout(w_dff_A_z3IMOOoq7_1),.din(w_dff_A_a4w9YAAH5_1),.clk(gclk));
	jdff dff_A_tzjLVKs71_1(.dout(w_dff_A_a4w9YAAH5_1),.din(w_dff_A_tzjLVKs71_1),.clk(gclk));
	jdff dff_A_IaYJB8XB0_1(.dout(w_dff_A_tzjLVKs71_1),.din(w_dff_A_IaYJB8XB0_1),.clk(gclk));
	jdff dff_A_yWUBgGhE0_1(.dout(w_dff_A_IaYJB8XB0_1),.din(w_dff_A_yWUBgGhE0_1),.clk(gclk));
	jdff dff_A_U3azGVav7_1(.dout(w_dff_A_yWUBgGhE0_1),.din(w_dff_A_U3azGVav7_1),.clk(gclk));
	jdff dff_A_34zAk1gL3_1(.dout(w_dff_A_U3azGVav7_1),.din(w_dff_A_34zAk1gL3_1),.clk(gclk));
	jdff dff_A_aQsWuZ0H7_1(.dout(w_dff_A_34zAk1gL3_1),.din(w_dff_A_aQsWuZ0H7_1),.clk(gclk));
	jdff dff_A_oK0W2Tqd0_1(.dout(w_dff_A_aQsWuZ0H7_1),.din(w_dff_A_oK0W2Tqd0_1),.clk(gclk));
	jdff dff_A_8Y5jKg274_1(.dout(w_dff_A_oK0W2Tqd0_1),.din(w_dff_A_8Y5jKg274_1),.clk(gclk));
	jdff dff_A_r9bJ7dDD4_1(.dout(w_dff_A_8Y5jKg274_1),.din(w_dff_A_r9bJ7dDD4_1),.clk(gclk));
	jdff dff_A_xNCVyGLH7_1(.dout(w_dff_A_r9bJ7dDD4_1),.din(w_dff_A_xNCVyGLH7_1),.clk(gclk));
	jdff dff_A_lIpPLIlz4_1(.dout(w_dff_A_xNCVyGLH7_1),.din(w_dff_A_lIpPLIlz4_1),.clk(gclk));
	jdff dff_A_PJktRTXK0_1(.dout(w_dff_A_lIpPLIlz4_1),.din(w_dff_A_PJktRTXK0_1),.clk(gclk));
	jdff dff_A_wbLq5Ln62_1(.dout(w_dff_A_PJktRTXK0_1),.din(w_dff_A_wbLq5Ln62_1),.clk(gclk));
	jdff dff_A_WeY6qbfv3_1(.dout(w_dff_A_wbLq5Ln62_1),.din(w_dff_A_WeY6qbfv3_1),.clk(gclk));
	jdff dff_B_XLnPo97s6_1(.din(n1084),.dout(w_dff_B_XLnPo97s6_1),.clk(gclk));
	jdff dff_B_9Hi7TPf16_1(.din(w_dff_B_XLnPo97s6_1),.dout(w_dff_B_9Hi7TPf16_1),.clk(gclk));
	jdff dff_B_nx7no1rL6_1(.din(w_dff_B_9Hi7TPf16_1),.dout(w_dff_B_nx7no1rL6_1),.clk(gclk));
	jdff dff_B_B6MzBm4y3_1(.din(w_dff_B_nx7no1rL6_1),.dout(w_dff_B_B6MzBm4y3_1),.clk(gclk));
	jdff dff_B_2Oqfe33G1_1(.din(w_dff_B_B6MzBm4y3_1),.dout(w_dff_B_2Oqfe33G1_1),.clk(gclk));
	jdff dff_B_9lMLVFMa8_1(.din(w_dff_B_2Oqfe33G1_1),.dout(w_dff_B_9lMLVFMa8_1),.clk(gclk));
	jdff dff_B_2GOZwkDz6_1(.din(w_dff_B_9lMLVFMa8_1),.dout(w_dff_B_2GOZwkDz6_1),.clk(gclk));
	jdff dff_B_CvbipimJ4_1(.din(w_dff_B_2GOZwkDz6_1),.dout(w_dff_B_CvbipimJ4_1),.clk(gclk));
	jdff dff_B_1UWSti0X0_1(.din(w_dff_B_CvbipimJ4_1),.dout(w_dff_B_1UWSti0X0_1),.clk(gclk));
	jdff dff_B_TzLFqooJ8_1(.din(w_dff_B_1UWSti0X0_1),.dout(w_dff_B_TzLFqooJ8_1),.clk(gclk));
	jdff dff_B_iadIqWnp5_1(.din(w_dff_B_TzLFqooJ8_1),.dout(w_dff_B_iadIqWnp5_1),.clk(gclk));
	jdff dff_B_CMFnyfac9_1(.din(w_dff_B_iadIqWnp5_1),.dout(w_dff_B_CMFnyfac9_1),.clk(gclk));
	jdff dff_B_1pUSJGLJ6_1(.din(n1081),.dout(w_dff_B_1pUSJGLJ6_1),.clk(gclk));
	jdff dff_B_f9HXrqET1_1(.din(w_dff_B_1pUSJGLJ6_1),.dout(w_dff_B_f9HXrqET1_1),.clk(gclk));
	jdff dff_A_QIGa4Vxw0_0(.dout(w_n852_7[0]),.din(w_dff_A_QIGa4Vxw0_0),.clk(gclk));
	jdff dff_A_jR5m4kYB0_0(.dout(w_dff_A_QIGa4Vxw0_0),.din(w_dff_A_jR5m4kYB0_0),.clk(gclk));
	jdff dff_A_YBwAHMoQ3_0(.dout(w_dff_A_jR5m4kYB0_0),.din(w_dff_A_YBwAHMoQ3_0),.clk(gclk));
	jdff dff_A_VUc2TGVB7_0(.dout(w_dff_A_YBwAHMoQ3_0),.din(w_dff_A_VUc2TGVB7_0),.clk(gclk));
	jdff dff_A_M4JBrh589_0(.dout(w_dff_A_VUc2TGVB7_0),.din(w_dff_A_M4JBrh589_0),.clk(gclk));
	jdff dff_A_XTX7mUEQ6_0(.dout(w_dff_A_M4JBrh589_0),.din(w_dff_A_XTX7mUEQ6_0),.clk(gclk));
	jdff dff_A_JkH3f71n7_0(.dout(w_dff_A_XTX7mUEQ6_0),.din(w_dff_A_JkH3f71n7_0),.clk(gclk));
	jdff dff_A_0xeiQsgV3_0(.dout(w_dff_A_JkH3f71n7_0),.din(w_dff_A_0xeiQsgV3_0),.clk(gclk));
	jdff dff_A_zgYvJxwK8_0(.dout(w_dff_A_0xeiQsgV3_0),.din(w_dff_A_zgYvJxwK8_0),.clk(gclk));
	jdff dff_A_8Y89BlU08_0(.dout(w_dff_A_zgYvJxwK8_0),.din(w_dff_A_8Y89BlU08_0),.clk(gclk));
	jdff dff_A_TPAe0JcF3_0(.dout(w_dff_A_8Y89BlU08_0),.din(w_dff_A_TPAe0JcF3_0),.clk(gclk));
	jdff dff_A_VSekOTg48_0(.dout(w_dff_A_TPAe0JcF3_0),.din(w_dff_A_VSekOTg48_0),.clk(gclk));
	jdff dff_A_jcig5Us53_2(.dout(w_n852_7[2]),.din(w_dff_A_jcig5Us53_2),.clk(gclk));
	jdff dff_A_D6EBUCPr5_2(.dout(w_dff_A_jcig5Us53_2),.din(w_dff_A_D6EBUCPr5_2),.clk(gclk));
	jdff dff_A_KeX40C7E4_2(.dout(w_dff_A_D6EBUCPr5_2),.din(w_dff_A_KeX40C7E4_2),.clk(gclk));
	jdff dff_A_Nx206cUP8_2(.dout(w_dff_A_KeX40C7E4_2),.din(w_dff_A_Nx206cUP8_2),.clk(gclk));
	jdff dff_A_2iImcXw27_2(.dout(w_dff_A_Nx206cUP8_2),.din(w_dff_A_2iImcXw27_2),.clk(gclk));
	jdff dff_A_T0lbkzxz2_2(.dout(w_dff_A_2iImcXw27_2),.din(w_dff_A_T0lbkzxz2_2),.clk(gclk));
	jdff dff_A_XFKTu5Ma0_2(.dout(w_dff_A_T0lbkzxz2_2),.din(w_dff_A_XFKTu5Ma0_2),.clk(gclk));
	jdff dff_A_wWADclJz7_2(.dout(w_dff_A_XFKTu5Ma0_2),.din(w_dff_A_wWADclJz7_2),.clk(gclk));
	jdff dff_A_r2F5r87r9_2(.dout(w_dff_A_wWADclJz7_2),.din(w_dff_A_r2F5r87r9_2),.clk(gclk));
	jdff dff_A_0nm2xijW1_2(.dout(w_dff_A_r2F5r87r9_2),.din(w_dff_A_0nm2xijW1_2),.clk(gclk));
	jdff dff_A_x0KPSQ9a9_2(.dout(w_dff_A_0nm2xijW1_2),.din(w_dff_A_x0KPSQ9a9_2),.clk(gclk));
	jdff dff_A_pqzAX0Kb3_2(.dout(w_dff_A_x0KPSQ9a9_2),.din(w_dff_A_pqzAX0Kb3_2),.clk(gclk));
	jdff dff_A_gQ0ePflD6_2(.dout(w_dff_A_pqzAX0Kb3_2),.din(w_dff_A_gQ0ePflD6_2),.clk(gclk));
	jdff dff_B_kXvSSlQq3_2(.din(G17),.dout(w_dff_B_kXvSSlQq3_2),.clk(gclk));
	jdff dff_A_EVSU5lyt1_0(.dout(w_G4089_7[0]),.din(w_dff_A_EVSU5lyt1_0),.clk(gclk));
	jdff dff_A_9dcVJLK39_0(.dout(w_dff_A_EVSU5lyt1_0),.din(w_dff_A_9dcVJLK39_0),.clk(gclk));
	jdff dff_A_ScFoQiCK6_0(.dout(w_dff_A_9dcVJLK39_0),.din(w_dff_A_ScFoQiCK6_0),.clk(gclk));
	jdff dff_A_UaGggClO3_0(.dout(w_dff_A_ScFoQiCK6_0),.din(w_dff_A_UaGggClO3_0),.clk(gclk));
	jdff dff_A_ODBnUjcP9_0(.dout(w_dff_A_UaGggClO3_0),.din(w_dff_A_ODBnUjcP9_0),.clk(gclk));
	jdff dff_A_aq99JOlU2_0(.dout(w_dff_A_ODBnUjcP9_0),.din(w_dff_A_aq99JOlU2_0),.clk(gclk));
	jdff dff_A_WdATVlpF8_0(.dout(w_dff_A_aq99JOlU2_0),.din(w_dff_A_WdATVlpF8_0),.clk(gclk));
	jdff dff_A_U8WVisHU5_0(.dout(w_dff_A_WdATVlpF8_0),.din(w_dff_A_U8WVisHU5_0),.clk(gclk));
	jdff dff_A_6ZccGNd50_0(.dout(w_dff_A_U8WVisHU5_0),.din(w_dff_A_6ZccGNd50_0),.clk(gclk));
	jdff dff_A_uCiFszMf5_0(.dout(w_dff_A_6ZccGNd50_0),.din(w_dff_A_uCiFszMf5_0),.clk(gclk));
	jdff dff_A_vsvynI6l4_0(.dout(w_dff_A_uCiFszMf5_0),.din(w_dff_A_vsvynI6l4_0),.clk(gclk));
	jdff dff_A_Cq8pswRj8_0(.dout(w_dff_A_vsvynI6l4_0),.din(w_dff_A_Cq8pswRj8_0),.clk(gclk));
	jdff dff_A_ttTEApFA6_0(.dout(w_dff_A_Cq8pswRj8_0),.din(w_dff_A_ttTEApFA6_0),.clk(gclk));
	jdff dff_A_ljERb6es5_2(.dout(w_G4089_7[2]),.din(w_dff_A_ljERb6es5_2),.clk(gclk));
	jdff dff_A_pDi6sdYw2_2(.dout(w_dff_A_ljERb6es5_2),.din(w_dff_A_pDi6sdYw2_2),.clk(gclk));
	jdff dff_A_4GRQRVfW1_2(.dout(w_dff_A_pDi6sdYw2_2),.din(w_dff_A_4GRQRVfW1_2),.clk(gclk));
	jdff dff_A_Zf8PCDGj7_2(.dout(w_dff_A_4GRQRVfW1_2),.din(w_dff_A_Zf8PCDGj7_2),.clk(gclk));
	jdff dff_A_dcOF4l9u1_2(.dout(w_dff_A_Zf8PCDGj7_2),.din(w_dff_A_dcOF4l9u1_2),.clk(gclk));
	jdff dff_A_blIdSm9Z9_2(.dout(w_dff_A_dcOF4l9u1_2),.din(w_dff_A_blIdSm9Z9_2),.clk(gclk));
	jdff dff_A_njF9yI397_2(.dout(w_dff_A_blIdSm9Z9_2),.din(w_dff_A_njF9yI397_2),.clk(gclk));
	jdff dff_A_hKxsYyVD2_2(.dout(w_dff_A_njF9yI397_2),.din(w_dff_A_hKxsYyVD2_2),.clk(gclk));
	jdff dff_A_Dd0CuaQU7_2(.dout(w_dff_A_hKxsYyVD2_2),.din(w_dff_A_Dd0CuaQU7_2),.clk(gclk));
	jdff dff_A_MfHzTLBw5_2(.dout(w_dff_A_Dd0CuaQU7_2),.din(w_dff_A_MfHzTLBw5_2),.clk(gclk));
	jdff dff_A_bUuxeHB43_2(.dout(w_dff_A_MfHzTLBw5_2),.din(w_dff_A_bUuxeHB43_2),.clk(gclk));
	jdff dff_A_X0pE9JoL7_2(.dout(w_dff_A_bUuxeHB43_2),.din(w_dff_A_X0pE9JoL7_2),.clk(gclk));
	jdff dff_A_pdByMsJz9_2(.dout(w_dff_A_X0pE9JoL7_2),.din(w_dff_A_pdByMsJz9_2),.clk(gclk));
	jdff dff_A_D48t4b391_2(.dout(w_dff_A_pdByMsJz9_2),.din(w_dff_A_D48t4b391_2),.clk(gclk));
	jdff dff_A_AtGQZzA59_2(.dout(w_dff_A_D48t4b391_2),.din(w_dff_A_AtGQZzA59_2),.clk(gclk));
	jdff dff_B_jTMkOXTe0_0(.din(n1097),.dout(w_dff_B_jTMkOXTe0_0),.clk(gclk));
	jdff dff_B_AnWszdc59_0(.din(w_dff_B_jTMkOXTe0_0),.dout(w_dff_B_AnWszdc59_0),.clk(gclk));
	jdff dff_B_nDCKo3bF5_0(.din(w_dff_B_AnWszdc59_0),.dout(w_dff_B_nDCKo3bF5_0),.clk(gclk));
	jdff dff_B_rFulOtJ36_0(.din(w_dff_B_nDCKo3bF5_0),.dout(w_dff_B_rFulOtJ36_0),.clk(gclk));
	jdff dff_B_0rAR0gjE5_0(.din(w_dff_B_rFulOtJ36_0),.dout(w_dff_B_0rAR0gjE5_0),.clk(gclk));
	jdff dff_B_jBCxrajO0_0(.din(w_dff_B_0rAR0gjE5_0),.dout(w_dff_B_jBCxrajO0_0),.clk(gclk));
	jdff dff_B_PZTJQhVQ7_0(.din(w_dff_B_jBCxrajO0_0),.dout(w_dff_B_PZTJQhVQ7_0),.clk(gclk));
	jdff dff_B_smqajFHb2_0(.din(w_dff_B_PZTJQhVQ7_0),.dout(w_dff_B_smqajFHb2_0),.clk(gclk));
	jdff dff_B_BANfFmOR9_0(.din(w_dff_B_smqajFHb2_0),.dout(w_dff_B_BANfFmOR9_0),.clk(gclk));
	jdff dff_B_8MOYsacq3_0(.din(w_dff_B_BANfFmOR9_0),.dout(w_dff_B_8MOYsacq3_0),.clk(gclk));
	jdff dff_B_15W2sopy9_0(.din(w_dff_B_8MOYsacq3_0),.dout(w_dff_B_15W2sopy9_0),.clk(gclk));
	jdff dff_B_3yet1Eid8_0(.din(w_dff_B_15W2sopy9_0),.dout(w_dff_B_3yet1Eid8_0),.clk(gclk));
	jdff dff_B_bccQQaUr7_0(.din(w_dff_B_3yet1Eid8_0),.dout(w_dff_B_bccQQaUr7_0),.clk(gclk));
	jdff dff_B_LKSFC2wQ7_0(.din(w_dff_B_bccQQaUr7_0),.dout(w_dff_B_LKSFC2wQ7_0),.clk(gclk));
	jdff dff_A_klxH40F92_1(.dout(w_G4090_3[1]),.din(w_dff_A_klxH40F92_1),.clk(gclk));
	jdff dff_A_7JjJKAlK5_2(.dout(w_G4090_3[2]),.din(w_dff_A_7JjJKAlK5_2),.clk(gclk));
	jdff dff_B_OdJBfi1i5_2(.din(G70),.dout(w_dff_B_OdJBfi1i5_2),.clk(gclk));
	jdff dff_B_VgSWLDu21_1(.din(n1090),.dout(w_dff_B_VgSWLDu21_1),.clk(gclk));
	jdff dff_B_X2FQN6vl5_1(.din(w_dff_B_VgSWLDu21_1),.dout(w_dff_B_X2FQN6vl5_1),.clk(gclk));
	jdff dff_B_e1PvzZF09_1(.din(w_dff_B_X2FQN6vl5_1),.dout(w_dff_B_e1PvzZF09_1),.clk(gclk));
	jdff dff_A_PJpeYuDT6_2(.dout(w_n854_3[2]),.din(w_dff_A_PJpeYuDT6_2),.clk(gclk));
	jdff dff_A_tfvNvX5W5_2(.dout(w_dff_A_PJpeYuDT6_2),.din(w_dff_A_tfvNvX5W5_2),.clk(gclk));
	jdff dff_B_ASjmq8333_0(.din(n1105),.dout(w_dff_B_ASjmq8333_0),.clk(gclk));
	jdff dff_B_Hj3oGY198_0(.din(w_dff_B_ASjmq8333_0),.dout(w_dff_B_Hj3oGY198_0),.clk(gclk));
	jdff dff_B_rDbHduqH3_0(.din(w_dff_B_Hj3oGY198_0),.dout(w_dff_B_rDbHduqH3_0),.clk(gclk));
	jdff dff_B_nBDadRNt4_0(.din(w_dff_B_rDbHduqH3_0),.dout(w_dff_B_nBDadRNt4_0),.clk(gclk));
	jdff dff_B_jggZGPEQ4_0(.din(w_dff_B_nBDadRNt4_0),.dout(w_dff_B_jggZGPEQ4_0),.clk(gclk));
	jdff dff_B_HsfYJFYe5_0(.din(w_dff_B_jggZGPEQ4_0),.dout(w_dff_B_HsfYJFYe5_0),.clk(gclk));
	jdff dff_B_Lk9noBZP0_0(.din(w_dff_B_HsfYJFYe5_0),.dout(w_dff_B_Lk9noBZP0_0),.clk(gclk));
	jdff dff_B_EIfO8b2u0_0(.din(w_dff_B_Lk9noBZP0_0),.dout(w_dff_B_EIfO8b2u0_0),.clk(gclk));
	jdff dff_B_xPAqGxKl7_0(.din(w_dff_B_EIfO8b2u0_0),.dout(w_dff_B_xPAqGxKl7_0),.clk(gclk));
	jdff dff_B_JOPDo2TI9_0(.din(w_dff_B_xPAqGxKl7_0),.dout(w_dff_B_JOPDo2TI9_0),.clk(gclk));
	jdff dff_B_ipUpO3rW9_0(.din(w_dff_B_JOPDo2TI9_0),.dout(w_dff_B_ipUpO3rW9_0),.clk(gclk));
	jdff dff_B_aDUJAUWH2_0(.din(w_dff_B_ipUpO3rW9_0),.dout(w_dff_B_aDUJAUWH2_0),.clk(gclk));
	jdff dff_B_Fjx6FOmC5_0(.din(w_dff_B_aDUJAUWH2_0),.dout(w_dff_B_Fjx6FOmC5_0),.clk(gclk));
	jdff dff_B_mH6hBIym7_0(.din(w_dff_B_Fjx6FOmC5_0),.dout(w_dff_B_mH6hBIym7_0),.clk(gclk));
	jdff dff_B_URYxDwxI2_0(.din(w_dff_B_mH6hBIym7_0),.dout(w_dff_B_URYxDwxI2_0),.clk(gclk));
	jdff dff_B_BcTWHefg0_0(.din(n1104),.dout(w_dff_B_BcTWHefg0_0),.clk(gclk));
	jdff dff_B_JeJ532NP3_1(.din(n1099),.dout(w_dff_B_JeJ532NP3_1),.clk(gclk));
	jdff dff_B_KfFW1Fkk3_0(.din(n1114),.dout(w_dff_B_KfFW1Fkk3_0),.clk(gclk));
	jdff dff_B_ywbCWTgM4_0(.din(w_dff_B_KfFW1Fkk3_0),.dout(w_dff_B_ywbCWTgM4_0),.clk(gclk));
	jdff dff_B_prB4rSPH2_0(.din(w_dff_B_ywbCWTgM4_0),.dout(w_dff_B_prB4rSPH2_0),.clk(gclk));
	jdff dff_B_4TUwwte84_0(.din(w_dff_B_prB4rSPH2_0),.dout(w_dff_B_4TUwwte84_0),.clk(gclk));
	jdff dff_B_GIcoci6S0_0(.din(w_dff_B_4TUwwte84_0),.dout(w_dff_B_GIcoci6S0_0),.clk(gclk));
	jdff dff_B_PYiQKGSz9_0(.din(w_dff_B_GIcoci6S0_0),.dout(w_dff_B_PYiQKGSz9_0),.clk(gclk));
	jdff dff_B_Pr2RB04Y5_0(.din(w_dff_B_PYiQKGSz9_0),.dout(w_dff_B_Pr2RB04Y5_0),.clk(gclk));
	jdff dff_B_5TMt0c0u6_0(.din(w_dff_B_Pr2RB04Y5_0),.dout(w_dff_B_5TMt0c0u6_0),.clk(gclk));
	jdff dff_B_S8q2Y4OC4_0(.din(w_dff_B_5TMt0c0u6_0),.dout(w_dff_B_S8q2Y4OC4_0),.clk(gclk));
	jdff dff_B_HnqMlbLq3_0(.din(w_dff_B_S8q2Y4OC4_0),.dout(w_dff_B_HnqMlbLq3_0),.clk(gclk));
	jdff dff_B_G7x6S2a65_0(.din(w_dff_B_HnqMlbLq3_0),.dout(w_dff_B_G7x6S2a65_0),.clk(gclk));
	jdff dff_B_VxYJZoC49_0(.din(w_dff_B_G7x6S2a65_0),.dout(w_dff_B_VxYJZoC49_0),.clk(gclk));
	jdff dff_B_ZTwiHh5O9_0(.din(n1113),.dout(w_dff_B_ZTwiHh5O9_0),.clk(gclk));
	jdff dff_B_YAFkuvKh2_0(.din(n1110),.dout(w_dff_B_YAFkuvKh2_0),.clk(gclk));
	jdff dff_A_Ni8pVGn12_0(.dout(w_n999_3[0]),.din(w_dff_A_Ni8pVGn12_0),.clk(gclk));
	jdff dff_A_EFk0UZYV1_0(.dout(w_dff_A_Ni8pVGn12_0),.din(w_dff_A_EFk0UZYV1_0),.clk(gclk));
	jdff dff_A_iItlQ5sG3_0(.dout(w_dff_A_EFk0UZYV1_0),.din(w_dff_A_iItlQ5sG3_0),.clk(gclk));
	jdff dff_A_sZ7qQDgD8_1(.dout(w_n999_3[1]),.din(w_dff_A_sZ7qQDgD8_1),.clk(gclk));
	jdff dff_A_O9LgnZvy7_1(.dout(w_dff_A_sZ7qQDgD8_1),.din(w_dff_A_O9LgnZvy7_1),.clk(gclk));
	jdff dff_A_jLVWflxl8_1(.dout(w_dff_A_O9LgnZvy7_1),.din(w_dff_A_jLVWflxl8_1),.clk(gclk));
	jdff dff_A_2d3zzqSu0_1(.dout(w_dff_A_jLVWflxl8_1),.din(w_dff_A_2d3zzqSu0_1),.clk(gclk));
	jdff dff_A_o7fd8FI87_1(.dout(w_dff_A_2d3zzqSu0_1),.din(w_dff_A_o7fd8FI87_1),.clk(gclk));
	jdff dff_A_WjqiIhQa3_1(.dout(w_dff_A_o7fd8FI87_1),.din(w_dff_A_WjqiIhQa3_1),.clk(gclk));
	jdff dff_A_CZiGEFGF6_1(.dout(w_dff_A_WjqiIhQa3_1),.din(w_dff_A_CZiGEFGF6_1),.clk(gclk));
	jdff dff_A_zBqjoj2v6_0(.dout(w_G1689_4[0]),.din(w_dff_A_zBqjoj2v6_0),.clk(gclk));
	jdff dff_A_O75CPJQW1_0(.dout(w_dff_A_zBqjoj2v6_0),.din(w_dff_A_O75CPJQW1_0),.clk(gclk));
	jdff dff_A_PDtPIIxj8_0(.dout(w_dff_A_O75CPJQW1_0),.din(w_dff_A_PDtPIIxj8_0),.clk(gclk));
	jdff dff_A_sPNwTG3r6_0(.dout(w_dff_A_PDtPIIxj8_0),.din(w_dff_A_sPNwTG3r6_0),.clk(gclk));
	jdff dff_A_QuEJt7JU6_0(.dout(w_dff_A_sPNwTG3r6_0),.din(w_dff_A_QuEJt7JU6_0),.clk(gclk));
	jdff dff_A_m4anppy54_1(.dout(w_G1689_4[1]),.din(w_dff_A_m4anppy54_1),.clk(gclk));
	jdff dff_A_mWAL1dEc8_1(.dout(w_dff_A_m4anppy54_1),.din(w_dff_A_mWAL1dEc8_1),.clk(gclk));
	jdff dff_A_pe7FpfbB5_1(.dout(w_dff_A_mWAL1dEc8_1),.din(w_dff_A_pe7FpfbB5_1),.clk(gclk));
	jdff dff_A_UK5h9lDg4_1(.dout(w_dff_A_pe7FpfbB5_1),.din(w_dff_A_UK5h9lDg4_1),.clk(gclk));
	jdff dff_A_umvdPpb11_1(.dout(w_dff_A_UK5h9lDg4_1),.din(w_dff_A_umvdPpb11_1),.clk(gclk));
	jdff dff_A_9ya0V2IF3_1(.dout(w_dff_A_umvdPpb11_1),.din(w_dff_A_9ya0V2IF3_1),.clk(gclk));
	jdff dff_A_90mI8wQY7_1(.dout(w_dff_A_9ya0V2IF3_1),.din(w_dff_A_90mI8wQY7_1),.clk(gclk));
	jdff dff_B_WgLtXsRa3_0(.din(n1123),.dout(w_dff_B_WgLtXsRa3_0),.clk(gclk));
	jdff dff_B_dpcbcZS22_0(.din(w_dff_B_WgLtXsRa3_0),.dout(w_dff_B_dpcbcZS22_0),.clk(gclk));
	jdff dff_B_FXWbEvUQ8_0(.din(w_dff_B_dpcbcZS22_0),.dout(w_dff_B_FXWbEvUQ8_0),.clk(gclk));
	jdff dff_B_IwjpEjEa5_0(.din(w_dff_B_FXWbEvUQ8_0),.dout(w_dff_B_IwjpEjEa5_0),.clk(gclk));
	jdff dff_B_yvqEcoX00_0(.din(w_dff_B_IwjpEjEa5_0),.dout(w_dff_B_yvqEcoX00_0),.clk(gclk));
	jdff dff_B_hi1waNrn4_0(.din(w_dff_B_yvqEcoX00_0),.dout(w_dff_B_hi1waNrn4_0),.clk(gclk));
	jdff dff_B_UvOcAHl45_0(.din(w_dff_B_hi1waNrn4_0),.dout(w_dff_B_UvOcAHl45_0),.clk(gclk));
	jdff dff_B_PzumL7cK2_0(.din(w_dff_B_UvOcAHl45_0),.dout(w_dff_B_PzumL7cK2_0),.clk(gclk));
	jdff dff_B_uvcy7Fap1_0(.din(w_dff_B_PzumL7cK2_0),.dout(w_dff_B_uvcy7Fap1_0),.clk(gclk));
	jdff dff_B_qhTRHxet7_0(.din(w_dff_B_uvcy7Fap1_0),.dout(w_dff_B_qhTRHxet7_0),.clk(gclk));
	jdff dff_B_823xxaS29_0(.din(w_dff_B_qhTRHxet7_0),.dout(w_dff_B_823xxaS29_0),.clk(gclk));
	jdff dff_B_93Pkxbgz0_0(.din(w_dff_B_823xxaS29_0),.dout(w_dff_B_93Pkxbgz0_0),.clk(gclk));
	jdff dff_B_qeCi42wT9_0(.din(n1122),.dout(w_dff_B_qeCi42wT9_0),.clk(gclk));
	jdff dff_B_3QEbJYIQ0_1(.din(n1117),.dout(w_dff_B_3QEbJYIQ0_1),.clk(gclk));
	jdff dff_A_GqhGK6Ko6_2(.dout(w_G137_8[2]),.din(w_dff_A_GqhGK6Ko6_2),.clk(gclk));
	jdff dff_A_iozQxqyE8_2(.dout(w_dff_A_GqhGK6Ko6_2),.din(w_dff_A_iozQxqyE8_2),.clk(gclk));
	jdff dff_A_RkhToDx10_2(.dout(w_dff_A_iozQxqyE8_2),.din(w_dff_A_RkhToDx10_2),.clk(gclk));
	jdff dff_B_kqndtGmv5_0(.din(n1132),.dout(w_dff_B_kqndtGmv5_0),.clk(gclk));
	jdff dff_B_becFu0ta7_0(.din(w_dff_B_kqndtGmv5_0),.dout(w_dff_B_becFu0ta7_0),.clk(gclk));
	jdff dff_B_WoZs7mQy0_0(.din(w_dff_B_becFu0ta7_0),.dout(w_dff_B_WoZs7mQy0_0),.clk(gclk));
	jdff dff_B_rCpMffo45_0(.din(w_dff_B_WoZs7mQy0_0),.dout(w_dff_B_rCpMffo45_0),.clk(gclk));
	jdff dff_B_l0rf3xqv1_0(.din(w_dff_B_rCpMffo45_0),.dout(w_dff_B_l0rf3xqv1_0),.clk(gclk));
	jdff dff_B_GkCLHMos6_0(.din(w_dff_B_l0rf3xqv1_0),.dout(w_dff_B_GkCLHMos6_0),.clk(gclk));
	jdff dff_B_jJdAtBfJ7_0(.din(w_dff_B_GkCLHMos6_0),.dout(w_dff_B_jJdAtBfJ7_0),.clk(gclk));
	jdff dff_B_H8GxjWtT6_0(.din(w_dff_B_jJdAtBfJ7_0),.dout(w_dff_B_H8GxjWtT6_0),.clk(gclk));
	jdff dff_B_Z2I8Q26F6_0(.din(w_dff_B_H8GxjWtT6_0),.dout(w_dff_B_Z2I8Q26F6_0),.clk(gclk));
	jdff dff_B_qb0oIRn35_0(.din(w_dff_B_Z2I8Q26F6_0),.dout(w_dff_B_qb0oIRn35_0),.clk(gclk));
	jdff dff_B_llJ7JzUh5_0(.din(w_dff_B_qb0oIRn35_0),.dout(w_dff_B_llJ7JzUh5_0),.clk(gclk));
	jdff dff_B_EcZf0wcu0_0(.din(w_dff_B_llJ7JzUh5_0),.dout(w_dff_B_EcZf0wcu0_0),.clk(gclk));
	jdff dff_B_Zp7KqYat4_0(.din(w_dff_B_EcZf0wcu0_0),.dout(w_dff_B_Zp7KqYat4_0),.clk(gclk));
	jdff dff_B_P8C265hN7_0(.din(n1131),.dout(w_dff_B_P8C265hN7_0),.clk(gclk));
	jdff dff_A_TGCFqqnx8_0(.dout(w_n993_3[0]),.din(w_dff_A_TGCFqqnx8_0),.clk(gclk));
	jdff dff_A_IhOTjENe3_0(.dout(w_dff_A_TGCFqqnx8_0),.din(w_dff_A_IhOTjENe3_0),.clk(gclk));
	jdff dff_A_qCkbwAAw0_1(.dout(w_n993_3[1]),.din(w_dff_A_qCkbwAAw0_1),.clk(gclk));
	jdff dff_B_Mg9EJ5kz0_1(.din(n1135),.dout(w_dff_B_Mg9EJ5kz0_1),.clk(gclk));
	jdff dff_B_LLmtF0zo3_1(.din(w_dff_B_Mg9EJ5kz0_1),.dout(w_dff_B_LLmtF0zo3_1),.clk(gclk));
	jdff dff_B_qJu1NlfA0_1(.din(w_dff_B_LLmtF0zo3_1),.dout(w_dff_B_qJu1NlfA0_1),.clk(gclk));
	jdff dff_B_rvQOjbCt1_1(.din(w_dff_B_qJu1NlfA0_1),.dout(w_dff_B_rvQOjbCt1_1),.clk(gclk));
	jdff dff_B_Svymtap50_1(.din(w_dff_B_rvQOjbCt1_1),.dout(w_dff_B_Svymtap50_1),.clk(gclk));
	jdff dff_B_4tNpsCiz0_1(.din(w_dff_B_Svymtap50_1),.dout(w_dff_B_4tNpsCiz0_1),.clk(gclk));
	jdff dff_B_Zk5OPS667_1(.din(w_dff_B_4tNpsCiz0_1),.dout(w_dff_B_Zk5OPS667_1),.clk(gclk));
	jdff dff_B_EKj1OGyS0_1(.din(w_dff_B_Zk5OPS667_1),.dout(w_dff_B_EKj1OGyS0_1),.clk(gclk));
	jdff dff_B_JPxczKMH0_1(.din(w_dff_B_EKj1OGyS0_1),.dout(w_dff_B_JPxczKMH0_1),.clk(gclk));
	jdff dff_B_lihhcyfF2_1(.din(w_dff_B_JPxczKMH0_1),.dout(w_dff_B_lihhcyfF2_1),.clk(gclk));
	jdff dff_B_nTKZW1Cr2_1(.din(w_dff_B_lihhcyfF2_1),.dout(w_dff_B_nTKZW1Cr2_1),.clk(gclk));
	jdff dff_B_0Qevwsqk0_1(.din(w_dff_B_nTKZW1Cr2_1),.dout(w_dff_B_0Qevwsqk0_1),.clk(gclk));
	jdff dff_B_v8txGR5D8_1(.din(w_dff_B_0Qevwsqk0_1),.dout(w_dff_B_v8txGR5D8_1),.clk(gclk));
	jdff dff_B_OGJYKypv5_1(.din(w_dff_B_v8txGR5D8_1),.dout(w_dff_B_OGJYKypv5_1),.clk(gclk));
	jdff dff_B_Jum9HHgx3_1(.din(w_dff_B_OGJYKypv5_1),.dout(w_dff_B_Jum9HHgx3_1),.clk(gclk));
	jdff dff_B_34ILIyfT2_1(.din(w_dff_B_Jum9HHgx3_1),.dout(w_dff_B_34ILIyfT2_1),.clk(gclk));
	jdff dff_B_YPte2gEs3_1(.din(w_dff_B_34ILIyfT2_1),.dout(w_dff_B_YPte2gEs3_1),.clk(gclk));
	jdff dff_B_EA3HTJ9z4_1(.din(n1136),.dout(w_dff_B_EA3HTJ9z4_1),.clk(gclk));
	jdff dff_B_vx3EQJt79_1(.din(w_dff_B_EA3HTJ9z4_1),.dout(w_dff_B_vx3EQJt79_1),.clk(gclk));
	jdff dff_B_3sRK3wxY0_1(.din(w_dff_B_vx3EQJt79_1),.dout(w_dff_B_3sRK3wxY0_1),.clk(gclk));
	jdff dff_B_YlHWyepJ5_1(.din(w_dff_B_3sRK3wxY0_1),.dout(w_dff_B_YlHWyepJ5_1),.clk(gclk));
	jdff dff_B_5iW68SO90_1(.din(w_dff_B_YlHWyepJ5_1),.dout(w_dff_B_5iW68SO90_1),.clk(gclk));
	jdff dff_B_gXd6knBH9_1(.din(w_dff_B_5iW68SO90_1),.dout(w_dff_B_gXd6knBH9_1),.clk(gclk));
	jdff dff_B_ZTf8MQTh6_1(.din(w_dff_B_gXd6knBH9_1),.dout(w_dff_B_ZTf8MQTh6_1),.clk(gclk));
	jdff dff_B_EEeSmgZ44_1(.din(w_dff_B_ZTf8MQTh6_1),.dout(w_dff_B_EEeSmgZ44_1),.clk(gclk));
	jdff dff_B_FfwXozkg9_1(.din(w_dff_B_EEeSmgZ44_1),.dout(w_dff_B_FfwXozkg9_1),.clk(gclk));
	jdff dff_B_kSkScJmV4_1(.din(w_dff_B_FfwXozkg9_1),.dout(w_dff_B_kSkScJmV4_1),.clk(gclk));
	jdff dff_B_UQrUsxZJ0_1(.din(w_dff_B_kSkScJmV4_1),.dout(w_dff_B_UQrUsxZJ0_1),.clk(gclk));
	jdff dff_B_APgQFSPT5_1(.din(w_dff_B_UQrUsxZJ0_1),.dout(w_dff_B_APgQFSPT5_1),.clk(gclk));
	jdff dff_B_Ddu4rOUr7_1(.din(w_dff_B_APgQFSPT5_1),.dout(w_dff_B_Ddu4rOUr7_1),.clk(gclk));
	jdff dff_B_UWwOies06_1(.din(w_dff_B_Ddu4rOUr7_1),.dout(w_dff_B_UWwOies06_1),.clk(gclk));
	jdff dff_B_FamlHe4h4_1(.din(w_dff_B_UWwOies06_1),.dout(w_dff_B_FamlHe4h4_1),.clk(gclk));
	jdff dff_B_M5ccVy9N4_1(.din(w_dff_B_FamlHe4h4_1),.dout(w_dff_B_M5ccVy9N4_1),.clk(gclk));
	jdff dff_B_b0B1pIhC7_1(.din(w_dff_B_M5ccVy9N4_1),.dout(w_dff_B_b0B1pIhC7_1),.clk(gclk));
	jdff dff_B_ZFXfjuh32_1(.din(n811),.dout(w_dff_B_ZFXfjuh32_1),.clk(gclk));
	jdff dff_B_auqaRaO50_1(.din(w_dff_B_ZFXfjuh32_1),.dout(w_dff_B_auqaRaO50_1),.clk(gclk));
	jdff dff_B_8hmBxek14_1(.din(w_dff_B_auqaRaO50_1),.dout(w_dff_B_8hmBxek14_1),.clk(gclk));
	jdff dff_B_N33P6Y9g5_1(.din(w_dff_B_8hmBxek14_1),.dout(w_dff_B_N33P6Y9g5_1),.clk(gclk));
	jdff dff_B_7EHHcQ7p9_1(.din(w_dff_B_N33P6Y9g5_1),.dout(w_dff_B_7EHHcQ7p9_1),.clk(gclk));
	jdff dff_B_RUU5PmNh1_1(.din(w_dff_B_7EHHcQ7p9_1),.dout(w_dff_B_RUU5PmNh1_1),.clk(gclk));
	jdff dff_B_60Q6r02i0_1(.din(w_dff_B_RUU5PmNh1_1),.dout(w_dff_B_60Q6r02i0_1),.clk(gclk));
	jdff dff_B_VBLEOHd63_1(.din(w_dff_B_60Q6r02i0_1),.dout(w_dff_B_VBLEOHd63_1),.clk(gclk));
	jdff dff_B_dDaX9vin5_1(.din(w_dff_B_VBLEOHd63_1),.dout(w_dff_B_dDaX9vin5_1),.clk(gclk));
	jdff dff_B_bvhI34cd3_1(.din(w_dff_B_dDaX9vin5_1),.dout(w_dff_B_bvhI34cd3_1),.clk(gclk));
	jdff dff_B_L8i3cC3X1_0(.din(n830),.dout(w_dff_B_L8i3cC3X1_0),.clk(gclk));
	jdff dff_B_VhaICDBA5_0(.din(w_dff_B_L8i3cC3X1_0),.dout(w_dff_B_VhaICDBA5_0),.clk(gclk));
	jdff dff_B_Vj2hRPJ01_0(.din(w_dff_B_VhaICDBA5_0),.dout(w_dff_B_Vj2hRPJ01_0),.clk(gclk));
	jdff dff_B_Xsa2AxOe3_0(.din(w_dff_B_Vj2hRPJ01_0),.dout(w_dff_B_Xsa2AxOe3_0),.clk(gclk));
	jdff dff_B_9QOCPZyK3_0(.din(w_dff_B_Xsa2AxOe3_0),.dout(w_dff_B_9QOCPZyK3_0),.clk(gclk));
	jdff dff_B_qH1jI7nu0_0(.din(w_dff_B_9QOCPZyK3_0),.dout(w_dff_B_qH1jI7nu0_0),.clk(gclk));
	jdff dff_B_HCIzJQ130_1(.din(n441),.dout(w_dff_B_HCIzJQ130_1),.clk(gclk));
	jdff dff_B_6jRaOUUu8_1(.din(n436),.dout(w_dff_B_6jRaOUUu8_1),.clk(gclk));
	jdff dff_B_ha0atSkg5_1(.din(n822),.dout(w_dff_B_ha0atSkg5_1),.clk(gclk));
	jdff dff_B_l2sgmT7n1_1(.din(w_dff_B_ha0atSkg5_1),.dout(w_dff_B_l2sgmT7n1_1),.clk(gclk));
	jdff dff_B_9llXinuz3_1(.din(w_dff_B_l2sgmT7n1_1),.dout(w_dff_B_9llXinuz3_1),.clk(gclk));
	jdff dff_B_w1vflgpN3_1(.din(w_dff_B_9llXinuz3_1),.dout(w_dff_B_w1vflgpN3_1),.clk(gclk));
	jdff dff_B_DbDIyK689_1(.din(w_dff_B_w1vflgpN3_1),.dout(w_dff_B_DbDIyK689_1),.clk(gclk));
	jdff dff_B_7lpTNgCX8_1(.din(G52),.dout(w_dff_B_7lpTNgCX8_1),.clk(gclk));
	jdff dff_B_PiyvcPOW4_1(.din(w_dff_B_7lpTNgCX8_1),.dout(w_dff_B_PiyvcPOW4_1),.clk(gclk));
	jdff dff_B_JgNojHL90_1(.din(n864),.dout(w_dff_B_JgNojHL90_1),.clk(gclk));
	jdff dff_B_YBylxNfk1_1(.din(w_dff_B_JgNojHL90_1),.dout(w_dff_B_YBylxNfk1_1),.clk(gclk));
	jdff dff_B_AO4fSm5S0_1(.din(w_dff_B_YBylxNfk1_1),.dout(w_dff_B_AO4fSm5S0_1),.clk(gclk));
	jdff dff_B_iQuXzvXk5_1(.din(w_dff_B_AO4fSm5S0_1),.dout(w_dff_B_iQuXzvXk5_1),.clk(gclk));
	jdff dff_B_3Z7GaG621_1(.din(w_dff_B_iQuXzvXk5_1),.dout(w_dff_B_3Z7GaG621_1),.clk(gclk));
	jdff dff_B_wyxXsqek5_1(.din(w_dff_B_3Z7GaG621_1),.dout(w_dff_B_wyxXsqek5_1),.clk(gclk));
	jdff dff_B_Zoh1sYfm8_1(.din(w_dff_B_wyxXsqek5_1),.dout(w_dff_B_Zoh1sYfm8_1),.clk(gclk));
	jdff dff_B_qcUKq5av0_1(.din(w_dff_B_Zoh1sYfm8_1),.dout(w_dff_B_qcUKq5av0_1),.clk(gclk));
	jdff dff_B_DowEpmwH5_1(.din(w_dff_B_qcUKq5av0_1),.dout(w_dff_B_DowEpmwH5_1),.clk(gclk));
	jdff dff_B_WwJ0NSWx1_1(.din(w_dff_B_DowEpmwH5_1),.dout(w_dff_B_WwJ0NSWx1_1),.clk(gclk));
	jdff dff_B_JfwrxIuU8_0(.din(n874),.dout(w_dff_B_JfwrxIuU8_0),.clk(gclk));
	jdff dff_B_RXLcMShc3_0(.din(w_dff_B_JfwrxIuU8_0),.dout(w_dff_B_RXLcMShc3_0),.clk(gclk));
	jdff dff_B_ZNulepyy7_0(.din(w_dff_B_RXLcMShc3_0),.dout(w_dff_B_ZNulepyy7_0),.clk(gclk));
	jdff dff_B_9p04cYS64_0(.din(w_dff_B_ZNulepyy7_0),.dout(w_dff_B_9p04cYS64_0),.clk(gclk));
	jdff dff_B_9wyuRh0q9_0(.din(w_dff_B_9p04cYS64_0),.dout(w_dff_B_9wyuRh0q9_0),.clk(gclk));
	jdff dff_B_mXSWqqI47_0(.din(w_dff_B_9wyuRh0q9_0),.dout(w_dff_B_mXSWqqI47_0),.clk(gclk));
	jdff dff_B_iLPynGW98_1(.din(n466),.dout(w_dff_B_iLPynGW98_1),.clk(gclk));
	jdff dff_B_Xl5HX38I0_1(.din(n461),.dout(w_dff_B_Xl5HX38I0_1),.clk(gclk));
	jdff dff_B_1sVHQLs98_1(.din(G122),.dout(w_dff_B_1sVHQLs98_1),.clk(gclk));
	jdff dff_B_qakfyPmS7_1(.din(w_dff_B_1sVHQLs98_1),.dout(w_dff_B_qakfyPmS7_1),.clk(gclk));
	jdff dff_B_33vZx0Wk4_2(.din(G170),.dout(w_dff_B_33vZx0Wk4_2),.clk(gclk));
	jdff dff_B_nOEfcpdq6_2(.din(G200),.dout(w_dff_B_nOEfcpdq6_2),.clk(gclk));
	jdff dff_B_Z7RccH1E0_2(.din(w_dff_B_nOEfcpdq6_2),.dout(w_dff_B_Z7RccH1E0_2),.clk(gclk));
	jdff dff_B_2uabgvoB1_0(.din(n1150),.dout(w_dff_B_2uabgvoB1_0),.clk(gclk));
	jdff dff_B_6yuWUfCZ6_0(.din(w_dff_B_2uabgvoB1_0),.dout(w_dff_B_6yuWUfCZ6_0),.clk(gclk));
	jdff dff_B_GoDZdDgy7_0(.din(w_dff_B_6yuWUfCZ6_0),.dout(w_dff_B_GoDZdDgy7_0),.clk(gclk));
	jdff dff_B_YLSk5S105_0(.din(w_dff_B_GoDZdDgy7_0),.dout(w_dff_B_YLSk5S105_0),.clk(gclk));
	jdff dff_B_x8W7rtEd7_0(.din(w_dff_B_YLSk5S105_0),.dout(w_dff_B_x8W7rtEd7_0),.clk(gclk));
	jdff dff_B_caJdmGw79_0(.din(w_dff_B_x8W7rtEd7_0),.dout(w_dff_B_caJdmGw79_0),.clk(gclk));
	jdff dff_B_Mpn6ZRof5_0(.din(w_dff_B_caJdmGw79_0),.dout(w_dff_B_Mpn6ZRof5_0),.clk(gclk));
	jdff dff_B_fssDAQDr5_0(.din(w_dff_B_Mpn6ZRof5_0),.dout(w_dff_B_fssDAQDr5_0),.clk(gclk));
	jdff dff_B_I09pJjqL9_0(.din(w_dff_B_fssDAQDr5_0),.dout(w_dff_B_I09pJjqL9_0),.clk(gclk));
	jdff dff_B_K7L63pMg9_0(.din(w_dff_B_I09pJjqL9_0),.dout(w_dff_B_K7L63pMg9_0),.clk(gclk));
	jdff dff_B_9pBGq7fL8_0(.din(w_dff_B_K7L63pMg9_0),.dout(w_dff_B_9pBGq7fL8_0),.clk(gclk));
	jdff dff_B_0mHdEneZ3_0(.din(w_dff_B_9pBGq7fL8_0),.dout(w_dff_B_0mHdEneZ3_0),.clk(gclk));
	jdff dff_B_KoFZQHj32_0(.din(n1149),.dout(w_dff_B_KoFZQHj32_0),.clk(gclk));
	jdff dff_B_focYSCPh7_2(.din(G158),.dout(w_dff_B_focYSCPh7_2),.clk(gclk));
	jdff dff_B_y55UpSa60_2(.din(G188),.dout(w_dff_B_y55UpSa60_2),.clk(gclk));
	jdff dff_B_bLSBvltT6_2(.din(w_dff_B_y55UpSa60_2),.dout(w_dff_B_bLSBvltT6_2),.clk(gclk));
	jdff dff_B_WevrzoMI7_0(.din(n1146),.dout(w_dff_B_WevrzoMI7_0),.clk(gclk));
	jdff dff_B_fCcYb1HK3_1(.din(n897),.dout(w_dff_B_fCcYb1HK3_1),.clk(gclk));
	jdff dff_B_u3X9cDNy1_1(.din(w_dff_B_fCcYb1HK3_1),.dout(w_dff_B_u3X9cDNy1_1),.clk(gclk));
	jdff dff_B_K1lhKfP65_1(.din(w_dff_B_u3X9cDNy1_1),.dout(w_dff_B_K1lhKfP65_1),.clk(gclk));
	jdff dff_B_170aO85v8_1(.din(w_dff_B_K1lhKfP65_1),.dout(w_dff_B_170aO85v8_1),.clk(gclk));
	jdff dff_B_cpKPO1eC0_1(.din(w_dff_B_170aO85v8_1),.dout(w_dff_B_cpKPO1eC0_1),.clk(gclk));
	jdff dff_B_4xRmqUBc3_1(.din(w_dff_B_cpKPO1eC0_1),.dout(w_dff_B_4xRmqUBc3_1),.clk(gclk));
	jdff dff_B_Zo5UtX9N0_0(.din(n904),.dout(w_dff_B_Zo5UtX9N0_0),.clk(gclk));
	jdff dff_B_PgKBBWqC0_0(.din(w_dff_B_Zo5UtX9N0_0),.dout(w_dff_B_PgKBBWqC0_0),.clk(gclk));
	jdff dff_B_3XH3aMG67_1(.din(n477),.dout(w_dff_B_3XH3aMG67_1),.clk(gclk));
	jdff dff_B_aQUqQRTG7_1(.din(n472),.dout(w_dff_B_aQUqQRTG7_1),.clk(gclk));
	jdff dff_A_Fpaig06N3_0(.dout(w_n901_0[0]),.din(w_dff_A_Fpaig06N3_0),.clk(gclk));
	jdff dff_A_S3xNVy6Y3_0(.dout(w_dff_A_Fpaig06N3_0),.din(w_dff_A_S3xNVy6Y3_0),.clk(gclk));
	jdff dff_B_Bm6FwsJ27_1(.din(n898),.dout(w_dff_B_Bm6FwsJ27_1),.clk(gclk));
	jdff dff_B_et0bOagX2_1(.din(G126),.dout(w_dff_B_et0bOagX2_1),.clk(gclk));
	jdff dff_B_yaRqtMlG8_1(.din(w_dff_B_et0bOagX2_1),.dout(w_dff_B_yaRqtMlG8_1),.clk(gclk));
	jdff dff_A_jx8wBfJg7_0(.dout(w_n1007_3[0]),.din(w_dff_A_jx8wBfJg7_0),.clk(gclk));
	jdff dff_A_GPrWgRHY4_1(.dout(w_n1007_3[1]),.din(w_dff_A_GPrWgRHY4_1),.clk(gclk));
	jdff dff_A_W3h0h3592_1(.dout(w_dff_A_GPrWgRHY4_1),.din(w_dff_A_W3h0h3592_1),.clk(gclk));
	jdff dff_A_b6OH5gk64_1(.dout(w_dff_A_W3h0h3592_1),.din(w_dff_A_b6OH5gk64_1),.clk(gclk));
	jdff dff_A_3lodQBnn5_1(.dout(w_dff_A_b6OH5gk64_1),.din(w_dff_A_3lodQBnn5_1),.clk(gclk));
	jdff dff_A_IIYIDKfM5_1(.dout(w_dff_A_3lodQBnn5_1),.din(w_dff_A_IIYIDKfM5_1),.clk(gclk));
	jdff dff_A_0UNvS99k5_1(.dout(w_dff_A_IIYIDKfM5_1),.din(w_dff_A_0UNvS99k5_1),.clk(gclk));
	jdff dff_B_HH3jiI268_1(.din(n762),.dout(w_dff_B_HH3jiI268_1),.clk(gclk));
	jdff dff_B_uEG2tnnx6_1(.din(w_dff_B_HH3jiI268_1),.dout(w_dff_B_uEG2tnnx6_1),.clk(gclk));
	jdff dff_B_gT9CoaJA8_1(.din(w_dff_B_uEG2tnnx6_1),.dout(w_dff_B_gT9CoaJA8_1),.clk(gclk));
	jdff dff_B_PVwQTJdm6_1(.din(w_dff_B_gT9CoaJA8_1),.dout(w_dff_B_PVwQTJdm6_1),.clk(gclk));
	jdff dff_B_e3NDGQlq6_1(.din(w_dff_B_PVwQTJdm6_1),.dout(w_dff_B_e3NDGQlq6_1),.clk(gclk));
	jdff dff_B_Cy1N3WdK5_1(.din(w_dff_B_e3NDGQlq6_1),.dout(w_dff_B_Cy1N3WdK5_1),.clk(gclk));
	jdff dff_B_IwJouphq5_1(.din(w_dff_B_Cy1N3WdK5_1),.dout(w_dff_B_IwJouphq5_1),.clk(gclk));
	jdff dff_B_W86gbJTr4_1(.din(w_dff_B_IwJouphq5_1),.dout(w_dff_B_W86gbJTr4_1),.clk(gclk));
	jdff dff_B_OhH9u7m70_0(.din(n773),.dout(w_dff_B_OhH9u7m70_0),.clk(gclk));
	jdff dff_B_eMz8smkY6_0(.din(w_dff_B_OhH9u7m70_0),.dout(w_dff_B_eMz8smkY6_0),.clk(gclk));
	jdff dff_B_zszzuhX94_0(.din(w_dff_B_eMz8smkY6_0),.dout(w_dff_B_zszzuhX94_0),.clk(gclk));
	jdff dff_B_5OSjEKub0_0(.din(w_dff_B_zszzuhX94_0),.dout(w_dff_B_5OSjEKub0_0),.clk(gclk));
	jdff dff_B_ndtQ8J8A2_1(.din(n382),.dout(w_dff_B_ndtQ8J8A2_1),.clk(gclk));
	jdff dff_B_1zB6cnra8_1(.din(n376),.dout(w_dff_B_1zB6cnra8_1),.clk(gclk));
	jdff dff_B_6ggxj0f47_0(.din(n769),.dout(w_dff_B_6ggxj0f47_0),.clk(gclk));
	jdff dff_B_bXxiS1Vt8_0(.din(w_dff_B_6ggxj0f47_0),.dout(w_dff_B_bXxiS1Vt8_0),.clk(gclk));
	jdff dff_B_gIJJEWgu0_0(.din(w_dff_B_bXxiS1Vt8_0),.dout(w_dff_B_gIJJEWgu0_0),.clk(gclk));
	jdff dff_B_xI1S3T0I1_0(.din(w_dff_B_gIJJEWgu0_0),.dout(w_dff_B_xI1S3T0I1_0),.clk(gclk));
	jdff dff_A_A1X0X5sl5_0(.dout(w_n753_1[0]),.din(w_dff_A_A1X0X5sl5_0),.clk(gclk));
	jdff dff_A_r1D25C2M4_0(.dout(w_dff_A_A1X0X5sl5_0),.din(w_dff_A_r1D25C2M4_0),.clk(gclk));
	jdff dff_A_gUq2Ekrx3_0(.dout(w_dff_A_r1D25C2M4_0),.din(w_dff_A_gUq2Ekrx3_0),.clk(gclk));
	jdff dff_A_dCKwEEz49_0(.dout(w_dff_A_gUq2Ekrx3_0),.din(w_dff_A_dCKwEEz49_0),.clk(gclk));
	jdff dff_A_OFptFf4R2_0(.dout(w_dff_A_dCKwEEz49_0),.din(w_dff_A_OFptFf4R2_0),.clk(gclk));
	jdff dff_A_rRRegyjH1_0(.dout(w_G4091_5[0]),.din(w_dff_A_rRRegyjH1_0),.clk(gclk));
	jdff dff_A_LHqCxxok4_0(.dout(w_dff_A_rRRegyjH1_0),.din(w_dff_A_LHqCxxok4_0),.clk(gclk));
	jdff dff_A_ggZuIP4t4_0(.dout(w_dff_A_LHqCxxok4_0),.din(w_dff_A_ggZuIP4t4_0),.clk(gclk));
	jdff dff_A_aEzecLA27_0(.dout(w_dff_A_ggZuIP4t4_0),.din(w_dff_A_aEzecLA27_0),.clk(gclk));
	jdff dff_A_FZrxiTix6_0(.dout(w_dff_A_aEzecLA27_0),.din(w_dff_A_FZrxiTix6_0),.clk(gclk));
	jdff dff_A_jxpmN3le4_2(.dout(w_G4091_5[2]),.din(w_dff_A_jxpmN3le4_2),.clk(gclk));
	jdff dff_A_2ievJ18M9_2(.dout(w_dff_A_jxpmN3le4_2),.din(w_dff_A_2ievJ18M9_2),.clk(gclk));
	jdff dff_A_awc91F4R1_2(.dout(w_dff_A_2ievJ18M9_2),.din(w_dff_A_awc91F4R1_2),.clk(gclk));
	jdff dff_B_ueIeBsUt2_1(.din(G129),.dout(w_dff_B_ueIeBsUt2_1),.clk(gclk));
	jdff dff_B_3PWJPcsw6_1(.din(w_dff_B_ueIeBsUt2_1),.dout(w_dff_B_3PWJPcsw6_1),.clk(gclk));
	jdff dff_A_bW5mP7gb9_1(.dout(w_G137_7[1]),.din(w_dff_A_bW5mP7gb9_1),.clk(gclk));
	jdff dff_A_2FQneTPi2_1(.dout(w_dff_A_bW5mP7gb9_1),.din(w_dff_A_2FQneTPi2_1),.clk(gclk));
	jdff dff_A_HsfrBfd07_1(.dout(w_dff_A_2FQneTPi2_1),.din(w_dff_A_HsfrBfd07_1),.clk(gclk));
	jdff dff_A_rpRPwpt80_1(.dout(w_dff_A_HsfrBfd07_1),.din(w_dff_A_rpRPwpt80_1),.clk(gclk));
	jdff dff_A_kkjYvLWy1_2(.dout(w_G137_7[2]),.din(w_dff_A_kkjYvLWy1_2),.clk(gclk));
	jdff dff_A_BkSHWRxp6_0(.dout(w_G137_2[0]),.din(w_dff_A_BkSHWRxp6_0),.clk(gclk));
	jdff dff_A_D5l59Qyj7_0(.dout(w_dff_A_BkSHWRxp6_0),.din(w_dff_A_D5l59Qyj7_0),.clk(gclk));
	jdff dff_A_a8XZ43Js4_1(.dout(w_G137_2[1]),.din(w_dff_A_a8XZ43Js4_1),.clk(gclk));
	jdff dff_A_5YLdQIJG0_1(.dout(w_dff_A_a8XZ43Js4_1),.din(w_dff_A_5YLdQIJG0_1),.clk(gclk));
	jdff dff_B_WkgTgB8s2_0(.din(n1159),.dout(w_dff_B_WkgTgB8s2_0),.clk(gclk));
	jdff dff_B_jj7QTbvu5_0(.din(w_dff_B_WkgTgB8s2_0),.dout(w_dff_B_jj7QTbvu5_0),.clk(gclk));
	jdff dff_B_G8YWFHHL2_0(.din(w_dff_B_jj7QTbvu5_0),.dout(w_dff_B_G8YWFHHL2_0),.clk(gclk));
	jdff dff_B_X7tN8g4a7_0(.din(w_dff_B_G8YWFHHL2_0),.dout(w_dff_B_X7tN8g4a7_0),.clk(gclk));
	jdff dff_B_Q3toTGed4_0(.din(w_dff_B_X7tN8g4a7_0),.dout(w_dff_B_Q3toTGed4_0),.clk(gclk));
	jdff dff_B_RTKBsLD81_0(.din(w_dff_B_Q3toTGed4_0),.dout(w_dff_B_RTKBsLD81_0),.clk(gclk));
	jdff dff_B_OTbKmBll2_0(.din(w_dff_B_RTKBsLD81_0),.dout(w_dff_B_OTbKmBll2_0),.clk(gclk));
	jdff dff_B_0strUoqp1_0(.din(w_dff_B_OTbKmBll2_0),.dout(w_dff_B_0strUoqp1_0),.clk(gclk));
	jdff dff_B_gHsL6Q9M2_0(.din(w_dff_B_0strUoqp1_0),.dout(w_dff_B_gHsL6Q9M2_0),.clk(gclk));
	jdff dff_B_hAveu1Gn1_0(.din(w_dff_B_gHsL6Q9M2_0),.dout(w_dff_B_hAveu1Gn1_0),.clk(gclk));
	jdff dff_B_4O5FlavO8_0(.din(w_dff_B_hAveu1Gn1_0),.dout(w_dff_B_4O5FlavO8_0),.clk(gclk));
	jdff dff_B_2iqz4Qca6_0(.din(w_dff_B_4O5FlavO8_0),.dout(w_dff_B_2iqz4Qca6_0),.clk(gclk));
	jdff dff_B_hrPZbIHP1_0(.din(n1158),.dout(w_dff_B_hrPZbIHP1_0),.clk(gclk));
	jdff dff_B_1lHDzU4e3_2(.din(G152),.dout(w_dff_B_1lHDzU4e3_2),.clk(gclk));
	jdff dff_B_iSPI2NTX6_2(.din(G155),.dout(w_dff_B_iSPI2NTX6_2),.clk(gclk));
	jdff dff_B_D4nHgDTr3_2(.din(w_dff_B_iSPI2NTX6_2),.dout(w_dff_B_D4nHgDTr3_2),.clk(gclk));
	jdff dff_B_SMMNfKzr1_1(.din(n1153),.dout(w_dff_B_SMMNfKzr1_1),.clk(gclk));
	jdff dff_B_fqoEoEid8_1(.din(n887),.dout(w_dff_B_fqoEoEid8_1),.clk(gclk));
	jdff dff_B_u34MmkyJ4_1(.din(w_dff_B_fqoEoEid8_1),.dout(w_dff_B_u34MmkyJ4_1),.clk(gclk));
	jdff dff_B_n9ADeJyW6_1(.din(w_dff_B_u34MmkyJ4_1),.dout(w_dff_B_n9ADeJyW6_1),.clk(gclk));
	jdff dff_B_loUnZsCX4_1(.din(w_dff_B_n9ADeJyW6_1),.dout(w_dff_B_loUnZsCX4_1),.clk(gclk));
	jdff dff_B_LGSufPLq9_1(.din(w_dff_B_loUnZsCX4_1),.dout(w_dff_B_LGSufPLq9_1),.clk(gclk));
	jdff dff_B_aDsq1VDI1_1(.din(w_dff_B_LGSufPLq9_1),.dout(w_dff_B_aDsq1VDI1_1),.clk(gclk));
	jdff dff_B_zJDkO5pI3_1(.din(w_dff_B_aDsq1VDI1_1),.dout(w_dff_B_zJDkO5pI3_1),.clk(gclk));
	jdff dff_B_G7gUarwH4_0(.din(n893),.dout(w_dff_B_G7gUarwH4_0),.clk(gclk));
	jdff dff_B_mBbYEeAf7_0(.din(w_dff_B_G7gUarwH4_0),.dout(w_dff_B_mBbYEeAf7_0),.clk(gclk));
	jdff dff_B_tjkDXg8y1_0(.din(w_dff_B_mBbYEeAf7_0),.dout(w_dff_B_tjkDXg8y1_0),.clk(gclk));
	jdff dff_B_ebyXWjon0_1(.din(n489),.dout(w_dff_B_ebyXWjon0_1),.clk(gclk));
	jdff dff_B_u09SE55u4_1(.din(n484),.dout(w_dff_B_u09SE55u4_1),.clk(gclk));
	jdff dff_B_L7NYPyV12_1(.din(G127),.dout(w_dff_B_L7NYPyV12_1),.clk(gclk));
	jdff dff_B_x4PZrSTy0_1(.din(w_dff_B_L7NYPyV12_1),.dout(w_dff_B_x4PZrSTy0_1),.clk(gclk));
	jdff dff_B_shPkzRl94_1(.din(n843),.dout(w_dff_B_shPkzRl94_1),.clk(gclk));
	jdff dff_B_whuvM3Q51_1(.din(w_dff_B_shPkzRl94_1),.dout(w_dff_B_whuvM3Q51_1),.clk(gclk));
	jdff dff_B_Q531J5yL6_1(.din(w_dff_B_whuvM3Q51_1),.dout(w_dff_B_Q531J5yL6_1),.clk(gclk));
	jdff dff_B_oUFeRytN2_1(.din(w_dff_B_Q531J5yL6_1),.dout(w_dff_B_oUFeRytN2_1),.clk(gclk));
	jdff dff_B_w8b7rGUl0_1(.din(w_dff_B_oUFeRytN2_1),.dout(w_dff_B_w8b7rGUl0_1),.clk(gclk));
	jdff dff_B_EOjIbgGb2_1(.din(w_dff_B_w8b7rGUl0_1),.dout(w_dff_B_EOjIbgGb2_1),.clk(gclk));
	jdff dff_B_vS45smQj3_1(.din(w_dff_B_EOjIbgGb2_1),.dout(w_dff_B_vS45smQj3_1),.clk(gclk));
	jdff dff_B_2qKPxEwx7_1(.din(n844),.dout(w_dff_B_2qKPxEwx7_1),.clk(gclk));
	jdff dff_B_KthAG3j72_1(.din(w_dff_B_2qKPxEwx7_1),.dout(w_dff_B_KthAG3j72_1),.clk(gclk));
	jdff dff_B_UygP64ca7_1(.din(w_dff_B_KthAG3j72_1),.dout(w_dff_B_UygP64ca7_1),.clk(gclk));
	jdff dff_B_vO0YA87X3_1(.din(w_dff_B_UygP64ca7_1),.dout(w_dff_B_vO0YA87X3_1),.clk(gclk));
	jdff dff_A_BkmynQCa8_0(.dout(w_n847_0[0]),.din(w_dff_A_BkmynQCa8_0),.clk(gclk));
	jdff dff_A_L7OWDQXr2_0(.dout(w_dff_A_BkmynQCa8_0),.din(w_dff_A_L7OWDQXr2_0),.clk(gclk));
	jdff dff_A_8dO28ARF5_0(.dout(w_dff_A_L7OWDQXr2_0),.din(w_dff_A_8dO28ARF5_0),.clk(gclk));
	jdff dff_A_6yGPh6Yv3_0(.dout(w_dff_A_8dO28ARF5_0),.din(w_dff_A_6yGPh6Yv3_0),.clk(gclk));
	jdff dff_A_QodupDsy5_0(.dout(w_dff_A_6yGPh6Yv3_0),.din(w_dff_A_QodupDsy5_0),.clk(gclk));
	jdff dff_B_6pT1L4yy1_1(.din(n393),.dout(w_dff_B_6pT1L4yy1_1),.clk(gclk));
	jdff dff_B_6bDH561l7_1(.din(n388),.dout(w_dff_B_6bDH561l7_1),.clk(gclk));
	jdff dff_B_kbMravUl7_1(.din(G119),.dout(w_dff_B_kbMravUl7_1),.clk(gclk));
	jdff dff_B_gzn3ppYX3_1(.din(w_dff_B_kbMravUl7_1),.dout(w_dff_B_gzn3ppYX3_1),.clk(gclk));
	jdff dff_B_L5gyn8Za0_0(.din(n1168),.dout(w_dff_B_L5gyn8Za0_0),.clk(gclk));
	jdff dff_B_ofQbNUbt5_0(.din(w_dff_B_L5gyn8Za0_0),.dout(w_dff_B_ofQbNUbt5_0),.clk(gclk));
	jdff dff_B_XBsHMG8d2_0(.din(w_dff_B_ofQbNUbt5_0),.dout(w_dff_B_XBsHMG8d2_0),.clk(gclk));
	jdff dff_B_qHGkKn6b1_0(.din(w_dff_B_XBsHMG8d2_0),.dout(w_dff_B_qHGkKn6b1_0),.clk(gclk));
	jdff dff_B_NPBVLA1n1_0(.din(w_dff_B_qHGkKn6b1_0),.dout(w_dff_B_NPBVLA1n1_0),.clk(gclk));
	jdff dff_B_r5x4ks831_0(.din(w_dff_B_NPBVLA1n1_0),.dout(w_dff_B_r5x4ks831_0),.clk(gclk));
	jdff dff_B_n4OzFfxW7_0(.din(w_dff_B_r5x4ks831_0),.dout(w_dff_B_n4OzFfxW7_0),.clk(gclk));
	jdff dff_B_RXu676aU5_0(.din(w_dff_B_n4OzFfxW7_0),.dout(w_dff_B_RXu676aU5_0),.clk(gclk));
	jdff dff_B_ykUVoXwi4_0(.din(w_dff_B_RXu676aU5_0),.dout(w_dff_B_ykUVoXwi4_0),.clk(gclk));
	jdff dff_B_AmiUrmva0_0(.din(w_dff_B_ykUVoXwi4_0),.dout(w_dff_B_AmiUrmva0_0),.clk(gclk));
	jdff dff_B_l9L4pKaY8_0(.din(w_dff_B_AmiUrmva0_0),.dout(w_dff_B_l9L4pKaY8_0),.clk(gclk));
	jdff dff_B_JJ9BEM7M2_0(.din(w_dff_B_l9L4pKaY8_0),.dout(w_dff_B_JJ9BEM7M2_0),.clk(gclk));
	jdff dff_B_yHemKvBF0_0(.din(w_dff_B_JJ9BEM7M2_0),.dout(w_dff_B_yHemKvBF0_0),.clk(gclk));
	jdff dff_B_zBKxwZd23_0(.din(n1167),.dout(w_dff_B_zBKxwZd23_0),.clk(gclk));
	jdff dff_B_TqW49frs3_2(.din(G146),.dout(w_dff_B_TqW49frs3_2),.clk(gclk));
	jdff dff_B_jiFN7tWL0_2(.din(G149),.dout(w_dff_B_jiFN7tWL0_2),.clk(gclk));
	jdff dff_B_dil3UexK9_2(.din(w_dff_B_jiFN7tWL0_2),.dout(w_dff_B_dil3UexK9_2),.clk(gclk));
	jdff dff_B_enXgUU5g4_1(.din(n878),.dout(w_dff_B_enXgUU5g4_1),.clk(gclk));
	jdff dff_B_sF91ZaHz1_1(.din(w_dff_B_enXgUU5g4_1),.dout(w_dff_B_sF91ZaHz1_1),.clk(gclk));
	jdff dff_B_KuakVzVa2_1(.din(w_dff_B_sF91ZaHz1_1),.dout(w_dff_B_KuakVzVa2_1),.clk(gclk));
	jdff dff_B_Kp0eYmnF7_1(.din(w_dff_B_KuakVzVa2_1),.dout(w_dff_B_Kp0eYmnF7_1),.clk(gclk));
	jdff dff_B_AbMsTt9T4_1(.din(w_dff_B_Kp0eYmnF7_1),.dout(w_dff_B_AbMsTt9T4_1),.clk(gclk));
	jdff dff_B_feve4orU4_1(.din(w_dff_B_AbMsTt9T4_1),.dout(w_dff_B_feve4orU4_1),.clk(gclk));
	jdff dff_B_vzEfQoki3_1(.din(w_dff_B_feve4orU4_1),.dout(w_dff_B_vzEfQoki3_1),.clk(gclk));
	jdff dff_B_EMjRTHoL2_1(.din(w_dff_B_vzEfQoki3_1),.dout(w_dff_B_EMjRTHoL2_1),.clk(gclk));
	jdff dff_B_5HsUXeEf0_0(.din(n883),.dout(w_dff_B_5HsUXeEf0_0),.clk(gclk));
	jdff dff_B_yefxkvvk1_0(.din(w_dff_B_5HsUXeEf0_0),.dout(w_dff_B_yefxkvvk1_0),.clk(gclk));
	jdff dff_B_u4BizK8s4_0(.din(w_dff_B_yefxkvvk1_0),.dout(w_dff_B_u4BizK8s4_0),.clk(gclk));
	jdff dff_B_fte8Gnki9_0(.din(w_dff_B_u4BizK8s4_0),.dout(w_dff_B_fte8Gnki9_0),.clk(gclk));
	jdff dff_B_4tWlY9bq3_1(.din(n524),.dout(w_dff_B_4tWlY9bq3_1),.clk(gclk));
	jdff dff_B_Icuqqmhk5_1(.din(n519),.dout(w_dff_B_Icuqqmhk5_1),.clk(gclk));
	jdff dff_A_ToPV5wHw3_2(.dout(w_G4092_7[2]),.din(w_dff_A_ToPV5wHw3_2),.clk(gclk));
	jdff dff_A_2Ag8oVJY1_2(.dout(w_dff_A_ToPV5wHw3_2),.din(w_dff_A_2Ag8oVJY1_2),.clk(gclk));
	jdff dff_A_sXs48mAJ2_2(.dout(w_dff_A_2Ag8oVJY1_2),.din(w_dff_A_sXs48mAJ2_2),.clk(gclk));
	jdff dff_A_pkrpol0q8_0(.dout(w_n880_0[0]),.din(w_dff_A_pkrpol0q8_0),.clk(gclk));
	jdff dff_A_Rc4alZ5s4_0(.dout(w_dff_A_pkrpol0q8_0),.din(w_dff_A_Rc4alZ5s4_0),.clk(gclk));
	jdff dff_A_nZHAwGjk1_0(.dout(w_dff_A_Rc4alZ5s4_0),.din(w_dff_A_nZHAwGjk1_0),.clk(gclk));
	jdff dff_A_1awNcfCx8_0(.dout(w_dff_A_nZHAwGjk1_0),.din(w_dff_A_1awNcfCx8_0),.clk(gclk));
	jdff dff_A_UqfCelNO3_0(.dout(w_dff_A_1awNcfCx8_0),.din(w_dff_A_UqfCelNO3_0),.clk(gclk));
	jdff dff_A_hjTmyCYm9_1(.dout(w_G4091_3[1]),.din(w_dff_A_hjTmyCYm9_1),.clk(gclk));
	jdff dff_A_Q826vMP53_2(.dout(w_G4091_3[2]),.din(w_dff_A_Q826vMP53_2),.clk(gclk));
	jdff dff_A_1d6GvdyF2_2(.dout(w_dff_A_Q826vMP53_2),.din(w_dff_A_1d6GvdyF2_2),.clk(gclk));
	jdff dff_B_JKC03qpZ6_1(.din(G128),.dout(w_dff_B_JKC03qpZ6_1),.clk(gclk));
	jdff dff_B_I2URrG8P0_1(.din(w_dff_B_JKC03qpZ6_1),.dout(w_dff_B_I2URrG8P0_1),.clk(gclk));
	jdff dff_A_Xf4DBYUo9_0(.dout(w_n1008_3[0]),.din(w_dff_A_Xf4DBYUo9_0),.clk(gclk));
	jdff dff_A_KBPGaox53_0(.dout(w_dff_A_Xf4DBYUo9_0),.din(w_dff_A_KBPGaox53_0),.clk(gclk));
	jdff dff_A_7kP6WV9w4_1(.dout(w_n1008_3[1]),.din(w_dff_A_7kP6WV9w4_1),.clk(gclk));
	jdff dff_B_fDChoKtb0_1(.din(n834),.dout(w_dff_B_fDChoKtb0_1),.clk(gclk));
	jdff dff_B_x5qi5khF1_1(.din(w_dff_B_fDChoKtb0_1),.dout(w_dff_B_x5qi5khF1_1),.clk(gclk));
	jdff dff_B_GJS68R1O6_1(.din(w_dff_B_x5qi5khF1_1),.dout(w_dff_B_GJS68R1O6_1),.clk(gclk));
	jdff dff_B_iKAp5iwP1_1(.din(w_dff_B_GJS68R1O6_1),.dout(w_dff_B_iKAp5iwP1_1),.clk(gclk));
	jdff dff_B_ltgUwjIp9_1(.din(w_dff_B_iKAp5iwP1_1),.dout(w_dff_B_ltgUwjIp9_1),.clk(gclk));
	jdff dff_B_rbnADBru1_1(.din(w_dff_B_ltgUwjIp9_1),.dout(w_dff_B_rbnADBru1_1),.clk(gclk));
	jdff dff_B_ATgaZu0P8_1(.din(w_dff_B_rbnADBru1_1),.dout(w_dff_B_ATgaZu0P8_1),.clk(gclk));
	jdff dff_B_o9FCPZlq3_1(.din(w_dff_B_ATgaZu0P8_1),.dout(w_dff_B_o9FCPZlq3_1),.clk(gclk));
	jdff dff_B_lXbCqQiA8_1(.din(w_dff_B_o9FCPZlq3_1),.dout(w_dff_B_lXbCqQiA8_1),.clk(gclk));
	jdff dff_B_3xas6Zzu6_0(.din(n839),.dout(w_dff_B_3xas6Zzu6_0),.clk(gclk));
	jdff dff_B_qP4G1cQn3_0(.din(w_dff_B_3xas6Zzu6_0),.dout(w_dff_B_qP4G1cQn3_0),.clk(gclk));
	jdff dff_B_hqjbsfWB2_0(.din(w_dff_B_qP4G1cQn3_0),.dout(w_dff_B_hqjbsfWB2_0),.clk(gclk));
	jdff dff_B_XFTdOrUM3_0(.din(w_dff_B_hqjbsfWB2_0),.dout(w_dff_B_XFTdOrUM3_0),.clk(gclk));
	jdff dff_B_h26Tk7ao5_0(.din(w_dff_B_XFTdOrUM3_0),.dout(w_dff_B_h26Tk7ao5_0),.clk(gclk));
	jdff dff_B_YwyUonoH8_0(.din(w_dff_B_h26Tk7ao5_0),.dout(w_dff_B_YwyUonoH8_0),.clk(gclk));
	jdff dff_B_xP1DKWMQ0_1(.din(n360),.dout(w_dff_B_xP1DKWMQ0_1),.clk(gclk));
	jdff dff_A_YBRV6JoW0_0(.dout(w_n749_11[0]),.din(w_dff_A_YBRV6JoW0_0),.clk(gclk));
	jdff dff_A_wmEkHaAt4_1(.dout(w_n749_11[1]),.din(w_dff_A_wmEkHaAt4_1),.clk(gclk));
	jdff dff_A_sGjd8nTr1_0(.dout(w_n749_3[0]),.din(w_dff_A_sGjd8nTr1_0),.clk(gclk));
	jdff dff_A_K6riXqK07_2(.dout(w_n749_3[2]),.din(w_dff_A_K6riXqK07_2),.clk(gclk));
	jdff dff_A_aIHJe3SX5_1(.dout(w_G4092_8[1]),.din(w_dff_A_aIHJe3SX5_1),.clk(gclk));
	jdff dff_A_fsG94DFF4_2(.dout(w_G4092_8[2]),.din(w_dff_A_fsG94DFF4_2),.clk(gclk));
	jdff dff_A_Q8gasQY60_0(.dout(w_n836_0[0]),.din(w_dff_A_Q8gasQY60_0),.clk(gclk));
	jdff dff_A_oo1MVGZV9_0(.dout(w_dff_A_Q8gasQY60_0),.din(w_dff_A_oo1MVGZV9_0),.clk(gclk));
	jdff dff_A_n4GJO1j45_0(.dout(w_dff_A_oo1MVGZV9_0),.din(w_dff_A_n4GJO1j45_0),.clk(gclk));
	jdff dff_A_Vg2LN1cI2_0(.dout(w_dff_A_n4GJO1j45_0),.din(w_dff_A_Vg2LN1cI2_0),.clk(gclk));
	jdff dff_A_4YVVfOtG6_0(.dout(w_dff_A_Vg2LN1cI2_0),.din(w_dff_A_4YVVfOtG6_0),.clk(gclk));
	jdff dff_A_d0YTLvCK5_0(.dout(w_dff_A_4YVVfOtG6_0),.din(w_dff_A_d0YTLvCK5_0),.clk(gclk));
	jdff dff_A_hFWOoDh04_0(.dout(w_dff_A_d0YTLvCK5_0),.din(w_dff_A_hFWOoDh04_0),.clk(gclk));
	jdff dff_A_dG2T47mw8_1(.dout(w_n753_0[1]),.din(w_dff_A_dG2T47mw8_1),.clk(gclk));
	jdff dff_A_butyZvEC9_1(.dout(w_dff_A_dG2T47mw8_1),.din(w_dff_A_butyZvEC9_1),.clk(gclk));
	jdff dff_A_NhU4K2DY7_2(.dout(w_n753_0[2]),.din(w_dff_A_NhU4K2DY7_2),.clk(gclk));
	jdff dff_A_rAsnwgLK2_2(.dout(w_dff_A_NhU4K2DY7_2),.din(w_dff_A_rAsnwgLK2_2),.clk(gclk));
	jdff dff_A_wmGJVR450_2(.dout(w_dff_A_rAsnwgLK2_2),.din(w_dff_A_wmGJVR450_2),.clk(gclk));
	jdff dff_A_edRtoikW4_2(.dout(w_dff_A_wmGJVR450_2),.din(w_dff_A_edRtoikW4_2),.clk(gclk));
	jdff dff_A_wBk3dmqZ4_2(.dout(w_dff_A_edRtoikW4_2),.din(w_dff_A_wBk3dmqZ4_2),.clk(gclk));
	jdff dff_B_6WPuEnl14_3(.din(n753),.dout(w_dff_B_6WPuEnl14_3),.clk(gclk));
	jdff dff_B_CabbYQKU6_3(.din(w_dff_B_6WPuEnl14_3),.dout(w_dff_B_CabbYQKU6_3),.clk(gclk));
	jdff dff_A_3t32s8AQ0_0(.dout(w_G4091_4[0]),.din(w_dff_A_3t32s8AQ0_0),.clk(gclk));
	jdff dff_A_2vAXRqdl8_0(.dout(w_dff_A_3t32s8AQ0_0),.din(w_dff_A_2vAXRqdl8_0),.clk(gclk));
	jdff dff_A_KdetSORu4_0(.dout(w_dff_A_2vAXRqdl8_0),.din(w_dff_A_KdetSORu4_0),.clk(gclk));
	jdff dff_A_wEzJNpno8_0(.dout(w_dff_A_KdetSORu4_0),.din(w_dff_A_wEzJNpno8_0),.clk(gclk));
	jdff dff_A_Bi8XuIGL9_2(.dout(w_G4091_4[2]),.din(w_dff_A_Bi8XuIGL9_2),.clk(gclk));
	jdff dff_A_NzwxeOLa6_2(.dout(w_dff_A_Bi8XuIGL9_2),.din(w_dff_A_NzwxeOLa6_2),.clk(gclk));
	jdff dff_A_ZzP2sz4o8_2(.dout(w_dff_A_NzwxeOLa6_2),.din(w_dff_A_ZzP2sz4o8_2),.clk(gclk));
	jdff dff_B_UQ6NEMru6_1(.din(G130),.dout(w_dff_B_UQ6NEMru6_1),.clk(gclk));
	jdff dff_B_0QuqJQqF4_1(.din(w_dff_B_UQ6NEMru6_1),.dout(w_dff_B_0QuqJQqF4_1),.clk(gclk));
	jdff dff_B_q6jkLf9D4_1(.din(n1173),.dout(w_dff_B_q6jkLf9D4_1),.clk(gclk));
	jdff dff_B_gvWWt8179_1(.din(w_dff_B_q6jkLf9D4_1),.dout(w_dff_B_gvWWt8179_1),.clk(gclk));
	jdff dff_B_HCVvmeyx9_1(.din(w_dff_B_gvWWt8179_1),.dout(w_dff_B_HCVvmeyx9_1),.clk(gclk));
	jdff dff_B_Towb3JhV2_1(.din(w_dff_B_HCVvmeyx9_1),.dout(w_dff_B_Towb3JhV2_1),.clk(gclk));
	jdff dff_B_DvYmC1dl7_1(.din(w_dff_B_Towb3JhV2_1),.dout(w_dff_B_DvYmC1dl7_1),.clk(gclk));
	jdff dff_B_X4A99RoH5_1(.din(w_dff_B_DvYmC1dl7_1),.dout(w_dff_B_X4A99RoH5_1),.clk(gclk));
	jdff dff_B_JmXHJZjB7_1(.din(w_dff_B_X4A99RoH5_1),.dout(w_dff_B_JmXHJZjB7_1),.clk(gclk));
	jdff dff_B_iZKQKn2k8_1(.din(w_dff_B_JmXHJZjB7_1),.dout(w_dff_B_iZKQKn2k8_1),.clk(gclk));
	jdff dff_B_dlWD6ODR7_1(.din(w_dff_B_iZKQKn2k8_1),.dout(w_dff_B_dlWD6ODR7_1),.clk(gclk));
	jdff dff_B_mPyDFJ913_1(.din(w_dff_B_dlWD6ODR7_1),.dout(w_dff_B_mPyDFJ913_1),.clk(gclk));
	jdff dff_B_p2ZINNA54_1(.din(w_dff_B_mPyDFJ913_1),.dout(w_dff_B_p2ZINNA54_1),.clk(gclk));
	jdff dff_B_G3tm66WX3_1(.din(w_dff_B_p2ZINNA54_1),.dout(w_dff_B_G3tm66WX3_1),.clk(gclk));
	jdff dff_B_hH16Nipb3_1(.din(w_dff_B_G3tm66WX3_1),.dout(w_dff_B_hH16Nipb3_1),.clk(gclk));
	jdff dff_B_qmmAf7A57_1(.din(w_dff_B_hH16Nipb3_1),.dout(w_dff_B_qmmAf7A57_1),.clk(gclk));
	jdff dff_B_DjZx3B481_1(.din(w_dff_B_qmmAf7A57_1),.dout(w_dff_B_DjZx3B481_1),.clk(gclk));
	jdff dff_B_JpgqzGnk3_1(.din(w_dff_B_DjZx3B481_1),.dout(w_dff_B_JpgqzGnk3_1),.clk(gclk));
	jdff dff_B_xmQ7M9xF6_1(.din(w_dff_B_JpgqzGnk3_1),.dout(w_dff_B_xmQ7M9xF6_1),.clk(gclk));
	jdff dff_B_Ivd7VMH57_1(.din(w_dff_B_xmQ7M9xF6_1),.dout(w_dff_B_Ivd7VMH57_1),.clk(gclk));
	jdff dff_B_XhjxZbDM4_1(.din(n1182),.dout(w_dff_B_XhjxZbDM4_1),.clk(gclk));
	jdff dff_B_6mQgSj0s0_1(.din(w_dff_B_XhjxZbDM4_1),.dout(w_dff_B_6mQgSj0s0_1),.clk(gclk));
	jdff dff_B_Jc6CjSTS4_1(.din(w_dff_B_6mQgSj0s0_1),.dout(w_dff_B_Jc6CjSTS4_1),.clk(gclk));
	jdff dff_B_ZqqnOma20_1(.din(w_dff_B_Jc6CjSTS4_1),.dout(w_dff_B_ZqqnOma20_1),.clk(gclk));
	jdff dff_B_YH5U34AS3_1(.din(w_dff_B_ZqqnOma20_1),.dout(w_dff_B_YH5U34AS3_1),.clk(gclk));
	jdff dff_B_QU4SmOqC5_1(.din(w_dff_B_YH5U34AS3_1),.dout(w_dff_B_QU4SmOqC5_1),.clk(gclk));
	jdff dff_B_8DMwpq5A1_1(.din(w_dff_B_QU4SmOqC5_1),.dout(w_dff_B_8DMwpq5A1_1),.clk(gclk));
	jdff dff_B_AS9Mmiq39_1(.din(w_dff_B_8DMwpq5A1_1),.dout(w_dff_B_AS9Mmiq39_1),.clk(gclk));
	jdff dff_B_WW3sFcDx4_1(.din(w_dff_B_AS9Mmiq39_1),.dout(w_dff_B_WW3sFcDx4_1),.clk(gclk));
	jdff dff_B_Pzz3Wyd36_1(.din(w_dff_B_WW3sFcDx4_1),.dout(w_dff_B_Pzz3Wyd36_1),.clk(gclk));
	jdff dff_B_dIuZ8OO31_0(.din(n1185),.dout(w_dff_B_dIuZ8OO31_0),.clk(gclk));
	jdff dff_B_KFEIgUKM1_0(.din(w_dff_B_dIuZ8OO31_0),.dout(w_dff_B_KFEIgUKM1_0),.clk(gclk));
	jdff dff_B_fj5SL7Wz5_0(.din(w_dff_B_KFEIgUKM1_0),.dout(w_dff_B_fj5SL7Wz5_0),.clk(gclk));
	jdff dff_B_Noki1fYK8_0(.din(w_dff_B_fj5SL7Wz5_0),.dout(w_dff_B_Noki1fYK8_0),.clk(gclk));
	jdff dff_B_snpjvWNa3_0(.din(w_dff_B_Noki1fYK8_0),.dout(w_dff_B_snpjvWNa3_0),.clk(gclk));
	jdff dff_B_p2Syoab75_0(.din(w_dff_B_snpjvWNa3_0),.dout(w_dff_B_p2Syoab75_0),.clk(gclk));
	jdff dff_B_82ZWVWhY8_0(.din(w_dff_B_p2Syoab75_0),.dout(w_dff_B_82ZWVWhY8_0),.clk(gclk));
	jdff dff_B_f4vuB5h31_0(.din(w_dff_B_82ZWVWhY8_0),.dout(w_dff_B_f4vuB5h31_0),.clk(gclk));
	jdff dff_B_yqVOazlv2_0(.din(w_dff_B_f4vuB5h31_0),.dout(w_dff_B_yqVOazlv2_0),.clk(gclk));
	jdff dff_B_32nEx41T3_0(.din(w_dff_B_yqVOazlv2_0),.dout(w_dff_B_32nEx41T3_0),.clk(gclk));
	jdff dff_B_aCFUkeCV3_0(.din(w_dff_B_32nEx41T3_0),.dout(w_dff_B_aCFUkeCV3_0),.clk(gclk));
	jdff dff_B_Dm3ZAoIg6_0(.din(w_dff_B_aCFUkeCV3_0),.dout(w_dff_B_Dm3ZAoIg6_0),.clk(gclk));
	jdff dff_B_IdJBzlcj5_0(.din(w_dff_B_Dm3ZAoIg6_0),.dout(w_dff_B_IdJBzlcj5_0),.clk(gclk));
	jdff dff_B_yVH7W18P1_0(.din(w_dff_B_IdJBzlcj5_0),.dout(w_dff_B_yVH7W18P1_0),.clk(gclk));
	jdff dff_B_VC63psti9_0(.din(w_dff_B_yVH7W18P1_0),.dout(w_dff_B_VC63psti9_0),.clk(gclk));
	jdff dff_B_2fXFua545_0(.din(w_dff_B_VC63psti9_0),.dout(w_dff_B_2fXFua545_0),.clk(gclk));
	jdff dff_B_YBD5ZGiK7_1(.din(n1175),.dout(w_dff_B_YBD5ZGiK7_1),.clk(gclk));
	jdff dff_B_ueT7NGUG0_1(.din(w_dff_B_YBD5ZGiK7_1),.dout(w_dff_B_ueT7NGUG0_1),.clk(gclk));
	jdff dff_B_twTMpFZ06_1(.din(w_dff_B_ueT7NGUG0_1),.dout(w_dff_B_twTMpFZ06_1),.clk(gclk));
	jdff dff_B_n8RVwXTT6_1(.din(n1176),.dout(w_dff_B_n8RVwXTT6_1),.clk(gclk));
	jdff dff_B_d8bkvUs89_1(.din(w_dff_B_n8RVwXTT6_1),.dout(w_dff_B_d8bkvUs89_1),.clk(gclk));
	jdff dff_B_q9dJCnUC4_1(.din(w_dff_B_d8bkvUs89_1),.dout(w_dff_B_q9dJCnUC4_1),.clk(gclk));
	jdff dff_B_AsmfxMTM7_1(.din(w_dff_B_q9dJCnUC4_1),.dout(w_dff_B_AsmfxMTM7_1),.clk(gclk));
	jdff dff_B_MPqOTiqy8_1(.din(w_dff_B_AsmfxMTM7_1),.dout(w_dff_B_MPqOTiqy8_1),.clk(gclk));
	jdff dff_B_oO0itrCv6_1(.din(w_dff_B_MPqOTiqy8_1),.dout(w_dff_B_oO0itrCv6_1),.clk(gclk));
	jdff dff_A_frpBbFp05_0(.dout(w_n1177_0[0]),.din(w_dff_A_frpBbFp05_0),.clk(gclk));
	jdff dff_A_aitynTe77_0(.dout(w_dff_A_frpBbFp05_0),.din(w_dff_A_aitynTe77_0),.clk(gclk));
	jdff dff_A_LVeLffIQ7_0(.dout(w_dff_A_aitynTe77_0),.din(w_dff_A_LVeLffIQ7_0),.clk(gclk));
	jdff dff_A_aaGYHJJX7_0(.dout(w_dff_A_LVeLffIQ7_0),.din(w_dff_A_aaGYHJJX7_0),.clk(gclk));
	jdff dff_A_sXkJnJh31_0(.dout(w_dff_A_aaGYHJJX7_0),.din(w_dff_A_sXkJnJh31_0),.clk(gclk));
	jdff dff_A_W9KmvIw12_0(.dout(w_dff_A_sXkJnJh31_0),.din(w_dff_A_W9KmvIw12_0),.clk(gclk));
	jdff dff_A_Ed2tEucy6_0(.dout(w_dff_A_W9KmvIw12_0),.din(w_dff_A_Ed2tEucy6_0),.clk(gclk));
	jdff dff_A_IYpiv8BJ8_0(.dout(w_dff_A_Ed2tEucy6_0),.din(w_dff_A_IYpiv8BJ8_0),.clk(gclk));
	jdff dff_A_JJOQs7Wi4_0(.dout(w_dff_A_IYpiv8BJ8_0),.din(w_dff_A_JJOQs7Wi4_0),.clk(gclk));
	jdff dff_A_RqAIpejz8_0(.dout(w_dff_A_JJOQs7Wi4_0),.din(w_dff_A_RqAIpejz8_0),.clk(gclk));
	jdff dff_A_64TXrpuB7_0(.dout(w_dff_A_RqAIpejz8_0),.din(w_dff_A_64TXrpuB7_0),.clk(gclk));
	jdff dff_B_OOPdKPrC6_2(.din(n1177),.dout(w_dff_B_OOPdKPrC6_2),.clk(gclk));
	jdff dff_B_Y02DkMOs8_2(.din(w_dff_B_OOPdKPrC6_2),.dout(w_dff_B_Y02DkMOs8_2),.clk(gclk));
	jdff dff_B_BP0FHnd11_2(.din(w_dff_B_Y02DkMOs8_2),.dout(w_dff_B_BP0FHnd11_2),.clk(gclk));
	jdff dff_B_QLVd4Pmh4_2(.din(w_dff_B_BP0FHnd11_2),.dout(w_dff_B_QLVd4Pmh4_2),.clk(gclk));
	jdff dff_B_504jPPon2_2(.din(w_dff_B_QLVd4Pmh4_2),.dout(w_dff_B_504jPPon2_2),.clk(gclk));
	jdff dff_A_5vksmMD30_0(.dout(w_G3717_0[0]),.din(w_dff_A_5vksmMD30_0),.clk(gclk));
	jdff dff_A_KNKfWtxB6_1(.dout(w_n428_1[1]),.din(w_dff_A_KNKfWtxB6_1),.clk(gclk));
	jdff dff_A_tCh7tCAi7_2(.dout(w_G3724_0[2]),.din(w_dff_A_tCh7tCAi7_2),.clk(gclk));
	jdff dff_A_dKM9fRZC2_2(.dout(w_dff_A_tCh7tCAi7_2),.din(w_dff_A_dKM9fRZC2_2),.clk(gclk));
	jdff dff_A_w6FAsZmD5_2(.dout(w_dff_A_dKM9fRZC2_2),.din(w_dff_A_w6FAsZmD5_2),.clk(gclk));
	jdff dff_A_HSDjMAYL4_2(.dout(w_dff_A_w6FAsZmD5_2),.din(w_dff_A_HSDjMAYL4_2),.clk(gclk));
	jdff dff_A_KHTTcMNu5_0(.dout(w_n1179_0[0]),.din(w_dff_A_KHTTcMNu5_0),.clk(gclk));
	jdff dff_A_oPjllWo38_0(.dout(w_dff_A_KHTTcMNu5_0),.din(w_dff_A_oPjllWo38_0),.clk(gclk));
	jdff dff_A_EcjYyVXo1_0(.dout(w_dff_A_oPjllWo38_0),.din(w_dff_A_EcjYyVXo1_0),.clk(gclk));
	jdff dff_A_fTJeBMfM6_0(.dout(w_dff_A_EcjYyVXo1_0),.din(w_dff_A_fTJeBMfM6_0),.clk(gclk));
	jdff dff_A_1kcaw7ez7_0(.dout(w_dff_A_fTJeBMfM6_0),.din(w_dff_A_1kcaw7ez7_0),.clk(gclk));
	jdff dff_A_DnJ5DBzF1_0(.dout(w_dff_A_1kcaw7ez7_0),.din(w_dff_A_DnJ5DBzF1_0),.clk(gclk));
	jdff dff_A_faTBR8PZ7_0(.dout(w_dff_A_DnJ5DBzF1_0),.din(w_dff_A_faTBR8PZ7_0),.clk(gclk));
	jdff dff_A_aqGYU6qh7_0(.dout(w_dff_A_faTBR8PZ7_0),.din(w_dff_A_aqGYU6qh7_0),.clk(gclk));
	jdff dff_A_hF4QMVNa8_0(.dout(w_dff_A_aqGYU6qh7_0),.din(w_dff_A_hF4QMVNa8_0),.clk(gclk));
	jdff dff_A_EMneLXFc6_0(.dout(w_dff_A_hF4QMVNa8_0),.din(w_dff_A_EMneLXFc6_0),.clk(gclk));
	jdff dff_A_5GDr8oCN8_0(.dout(w_dff_A_EMneLXFc6_0),.din(w_dff_A_5GDr8oCN8_0),.clk(gclk));
	jdff dff_B_3ZtdagPq9_1(.din(G132),.dout(w_dff_B_3ZtdagPq9_1),.clk(gclk));
	jdff dff_B_u0WOS3Pc4_1(.din(w_dff_B_3ZtdagPq9_1),.dout(w_dff_B_u0WOS3Pc4_1),.clk(gclk));
	jdff dff_B_V53cg0X02_1(.din(w_dff_B_u0WOS3Pc4_1),.dout(w_dff_B_V53cg0X02_1),.clk(gclk));
	jdff dff_B_K8TahF035_1(.din(w_dff_B_V53cg0X02_1),.dout(w_dff_B_K8TahF035_1),.clk(gclk));
	jdff dff_B_btmOODy13_1(.din(n1223),.dout(w_dff_B_btmOODy13_1),.clk(gclk));
	jdff dff_B_qEQQpsKk5_0(.din(n1227),.dout(w_dff_B_qEQQpsKk5_0),.clk(gclk));
	jdff dff_B_r9MmtNCY7_0(.din(w_dff_B_qEQQpsKk5_0),.dout(w_dff_B_r9MmtNCY7_0),.clk(gclk));
	jdff dff_B_MS3xUnKy5_0(.din(w_dff_B_r9MmtNCY7_0),.dout(w_dff_B_MS3xUnKy5_0),.clk(gclk));
	jdff dff_B_xC81aw5z5_0(.din(w_dff_B_MS3xUnKy5_0),.dout(w_dff_B_xC81aw5z5_0),.clk(gclk));
	jdff dff_B_eh53O0zL0_0(.din(n1226),.dout(w_dff_B_eh53O0zL0_0),.clk(gclk));
	jdff dff_A_PcpneghQ7_0(.dout(w_G559_0[0]),.din(w_dff_A_PcpneghQ7_0),.clk(gclk));
	jdff dff_A_2cTOs3ML8_0(.dout(w_dff_A_PcpneghQ7_0),.din(w_dff_A_2cTOs3ML8_0),.clk(gclk));
	jdff dff_B_T9BYHnEv1_0(.din(n668),.dout(w_dff_B_T9BYHnEv1_0),.clk(gclk));
	jdff dff_B_6lPqW0NK3_1(.din(n663),.dout(w_dff_B_6lPqW0NK3_1),.clk(gclk));
	jdff dff_B_TJmzSrc90_1(.din(n916),.dout(w_dff_B_TJmzSrc90_1),.clk(gclk));
	jdff dff_B_odN55ZPf6_1(.din(n917),.dout(w_dff_B_odN55ZPf6_1),.clk(gclk));
	jdff dff_B_z8WZTYfZ4_0(.din(n915),.dout(w_dff_B_z8WZTYfZ4_0),.clk(gclk));
	jdff dff_B_qe1eSGki3_1(.din(n913),.dout(w_dff_B_qe1eSGki3_1),.clk(gclk));
	jdff dff_B_lJIOTZQH6_0(.din(G372),.dout(w_dff_B_lJIOTZQH6_0),.clk(gclk));
	jdff dff_B_4gwmfbNS1_1(.din(n909),.dout(w_dff_B_4gwmfbNS1_1),.clk(gclk));
	jdff dff_B_uu6sxKaR8_1(.din(n907),.dout(w_dff_B_uu6sxKaR8_1),.clk(gclk));
	jdff dff_B_7wKi2Shd7_1(.din(w_dff_B_uu6sxKaR8_1),.dout(w_dff_B_7wKi2Shd7_1),.clk(gclk));
	jdff dff_B_RV9gjbcG5_0(.din(n1222),.dout(w_dff_B_RV9gjbcG5_0),.clk(gclk));
	jdff dff_B_FcX5Hktv6_0(.din(w_dff_B_RV9gjbcG5_0),.dout(w_dff_B_FcX5Hktv6_0),.clk(gclk));
	jdff dff_B_2ri51vPv3_0(.din(w_dff_B_FcX5Hktv6_0),.dout(w_dff_B_2ri51vPv3_0),.clk(gclk));
	jdff dff_B_GktndBhK1_0(.din(n678),.dout(w_dff_B_GktndBhK1_0),.clk(gclk));
	jdff dff_B_fJLKRzUl4_1(.din(n672),.dout(w_dff_B_fJLKRzUl4_1),.clk(gclk));
	jdff dff_A_lNYH5L6n4_0(.dout(w_G245_0[0]),.din(w_dff_A_lNYH5L6n4_0),.clk(gclk));
	jdff dff_A_mwcxET8O5_0(.dout(w_dff_A_lNYH5L6n4_0),.din(w_dff_A_mwcxET8O5_0),.clk(gclk));
	jdff dff_A_yPcGyAXE4_0(.dout(w_dff_A_mwcxET8O5_0),.din(w_dff_A_yPcGyAXE4_0),.clk(gclk));
	jdff dff_A_h3X8GGaS8_0(.dout(w_dff_A_yPcGyAXE4_0),.din(w_dff_A_h3X8GGaS8_0),.clk(gclk));
	jdff dff_B_L0gb3Hkz2_1(.din(n926),.dout(w_dff_B_L0gb3Hkz2_1),.clk(gclk));
	jdff dff_B_yyP4thTY9_1(.din(n930),.dout(w_dff_B_yyP4thTY9_1),.clk(gclk));
	jdff dff_B_S0xTrdX29_1(.din(w_dff_B_yyP4thTY9_1),.dout(w_dff_B_S0xTrdX29_1),.clk(gclk));
	jdff dff_B_da3s2Xhl4_1(.din(n927),.dout(w_dff_B_da3s2Xhl4_1),.clk(gclk));
	jdff dff_B_LYANNG6m0_1(.din(G292),.dout(w_dff_B_LYANNG6m0_1),.clk(gclk));
	jdff dff_B_cS5Q11L10_1(.din(n1263),.dout(w_dff_B_cS5Q11L10_1),.clk(gclk));
	jdff dff_B_eeGo6B2W3_1(.din(w_dff_B_cS5Q11L10_1),.dout(w_dff_B_eeGo6B2W3_1),.clk(gclk));
	jdff dff_B_GjL4teN95_1(.din(w_dff_B_eeGo6B2W3_1),.dout(w_dff_B_GjL4teN95_1),.clk(gclk));
	jdff dff_B_zTLMdmw39_1(.din(w_dff_B_GjL4teN95_1),.dout(w_dff_B_zTLMdmw39_1),.clk(gclk));
	jdff dff_B_9ra4wDRl9_1(.din(w_dff_B_zTLMdmw39_1),.dout(w_dff_B_9ra4wDRl9_1),.clk(gclk));
	jdff dff_B_Fh2gQ6be0_1(.din(w_dff_B_9ra4wDRl9_1),.dout(w_dff_B_Fh2gQ6be0_1),.clk(gclk));
	jdff dff_B_Juy0Tt2p6_1(.din(w_dff_B_Fh2gQ6be0_1),.dout(w_dff_B_Juy0Tt2p6_1),.clk(gclk));
	jdff dff_B_PWnJhhAO2_1(.din(w_dff_B_Juy0Tt2p6_1),.dout(w_dff_B_PWnJhhAO2_1),.clk(gclk));
	jdff dff_B_vRy6dq1h5_1(.din(w_dff_B_PWnJhhAO2_1),.dout(w_dff_B_vRy6dq1h5_1),.clk(gclk));
	jdff dff_B_vSFtWIEC2_1(.din(w_dff_B_vRy6dq1h5_1),.dout(w_dff_B_vSFtWIEC2_1),.clk(gclk));
	jdff dff_B_1g47Foue8_1(.din(w_dff_B_vSFtWIEC2_1),.dout(w_dff_B_1g47Foue8_1),.clk(gclk));
	jdff dff_B_kAndRELX8_1(.din(w_dff_B_1g47Foue8_1),.dout(w_dff_B_kAndRELX8_1),.clk(gclk));
	jdff dff_B_6EBdFV0W8_1(.din(w_dff_B_kAndRELX8_1),.dout(w_dff_B_6EBdFV0W8_1),.clk(gclk));
	jdff dff_B_ziHDoDNs1_1(.din(w_dff_B_6EBdFV0W8_1),.dout(w_dff_B_ziHDoDNs1_1),.clk(gclk));
	jdff dff_B_xPNZux7h1_1(.din(w_dff_B_ziHDoDNs1_1),.dout(w_dff_B_xPNZux7h1_1),.clk(gclk));
	jdff dff_B_X36jGgTQ2_1(.din(w_dff_B_xPNZux7h1_1),.dout(w_dff_B_X36jGgTQ2_1),.clk(gclk));
	jdff dff_B_QrhlCgfN8_1(.din(w_dff_B_X36jGgTQ2_1),.dout(w_dff_B_QrhlCgfN8_1),.clk(gclk));
	jdff dff_B_eBNDRAH97_1(.din(w_dff_B_QrhlCgfN8_1),.dout(w_dff_B_eBNDRAH97_1),.clk(gclk));
	jdff dff_B_Oa4FPMrk7_1(.din(w_dff_B_eBNDRAH97_1),.dout(w_dff_B_Oa4FPMrk7_1),.clk(gclk));
	jdff dff_B_yXaaSN0r9_1(.din(n1260),.dout(w_dff_B_yXaaSN0r9_1),.clk(gclk));
	jdff dff_B_EllftlNr1_1(.din(w_dff_B_yXaaSN0r9_1),.dout(w_dff_B_EllftlNr1_1),.clk(gclk));
	jdff dff_A_E29owVpO8_2(.dout(w_n852_6[2]),.din(w_dff_A_E29owVpO8_2),.clk(gclk));
	jdff dff_A_fLvleYC64_2(.dout(w_dff_A_E29owVpO8_2),.din(w_dff_A_fLvleYC64_2),.clk(gclk));
	jdff dff_A_4caMF2zU4_2(.dout(w_dff_A_fLvleYC64_2),.din(w_dff_A_4caMF2zU4_2),.clk(gclk));
	jdff dff_A_vf3Gj3wd1_2(.dout(w_dff_A_4caMF2zU4_2),.din(w_dff_A_vf3Gj3wd1_2),.clk(gclk));
	jdff dff_A_jkbpH5wQ5_2(.dout(w_dff_A_vf3Gj3wd1_2),.din(w_dff_A_jkbpH5wQ5_2),.clk(gclk));
	jdff dff_A_KDIgANww9_2(.dout(w_dff_A_jkbpH5wQ5_2),.din(w_dff_A_KDIgANww9_2),.clk(gclk));
	jdff dff_A_RyklNXlN7_2(.dout(w_dff_A_KDIgANww9_2),.din(w_dff_A_RyklNXlN7_2),.clk(gclk));
	jdff dff_A_oOfK8kwV9_2(.dout(w_dff_A_RyklNXlN7_2),.din(w_dff_A_oOfK8kwV9_2),.clk(gclk));
	jdff dff_A_9shosCWL7_2(.dout(w_dff_A_oOfK8kwV9_2),.din(w_dff_A_9shosCWL7_2),.clk(gclk));
	jdff dff_A_s4vdH9qE5_2(.dout(w_dff_A_9shosCWL7_2),.din(w_dff_A_s4vdH9qE5_2),.clk(gclk));
	jdff dff_A_KgpDjXJt6_2(.dout(w_dff_A_s4vdH9qE5_2),.din(w_dff_A_KgpDjXJt6_2),.clk(gclk));
	jdff dff_A_dlwQqz3t3_2(.dout(w_G4089_6[2]),.din(w_dff_A_dlwQqz3t3_2),.clk(gclk));
	jdff dff_A_eJ7z3tGy4_2(.dout(w_dff_A_dlwQqz3t3_2),.din(w_dff_A_eJ7z3tGy4_2),.clk(gclk));
	jdff dff_A_VsuE2nZs8_2(.dout(w_dff_A_eJ7z3tGy4_2),.din(w_dff_A_VsuE2nZs8_2),.clk(gclk));
	jdff dff_A_C4BKBJs97_2(.dout(w_dff_A_VsuE2nZs8_2),.din(w_dff_A_C4BKBJs97_2),.clk(gclk));
	jdff dff_A_AlozjURd2_2(.dout(w_dff_A_C4BKBJs97_2),.din(w_dff_A_AlozjURd2_2),.clk(gclk));
	jdff dff_A_r60OqSVx4_2(.dout(w_dff_A_AlozjURd2_2),.din(w_dff_A_r60OqSVx4_2),.clk(gclk));
	jdff dff_A_VMaU69V91_2(.dout(w_dff_A_r60OqSVx4_2),.din(w_dff_A_VMaU69V91_2),.clk(gclk));
	jdff dff_A_aPSaX0Ac6_2(.dout(w_dff_A_VMaU69V91_2),.din(w_dff_A_aPSaX0Ac6_2),.clk(gclk));
	jdff dff_A_4OA7GnSW0_2(.dout(w_dff_A_aPSaX0Ac6_2),.din(w_dff_A_4OA7GnSW0_2),.clk(gclk));
	jdff dff_A_s9qkZEY39_2(.dout(w_dff_A_4OA7GnSW0_2),.din(w_dff_A_s9qkZEY39_2),.clk(gclk));
	jdff dff_A_N0O1RP3f7_2(.dout(w_dff_A_s9qkZEY39_2),.din(w_dff_A_N0O1RP3f7_2),.clk(gclk));
	jdff dff_A_6l7D93C82_2(.dout(w_dff_A_N0O1RP3f7_2),.din(w_dff_A_6l7D93C82_2),.clk(gclk));
	jdff dff_A_VDxF2ZcP8_2(.dout(w_dff_A_6l7D93C82_2),.din(w_dff_A_VDxF2ZcP8_2),.clk(gclk));
	jdff dff_A_Uy0iffnN3_2(.dout(w_dff_A_VDxF2ZcP8_2),.din(w_dff_A_Uy0iffnN3_2),.clk(gclk));
	jdff dff_B_ZRoBCCT49_0(.din(n1276),.dout(w_dff_B_ZRoBCCT49_0),.clk(gclk));
	jdff dff_B_fmSecLm54_0(.din(w_dff_B_ZRoBCCT49_0),.dout(w_dff_B_fmSecLm54_0),.clk(gclk));
	jdff dff_B_zgNCQm5D1_0(.din(w_dff_B_fmSecLm54_0),.dout(w_dff_B_zgNCQm5D1_0),.clk(gclk));
	jdff dff_B_FHmxkujZ1_0(.din(w_dff_B_zgNCQm5D1_0),.dout(w_dff_B_FHmxkujZ1_0),.clk(gclk));
	jdff dff_B_amlKhovH2_0(.din(w_dff_B_FHmxkujZ1_0),.dout(w_dff_B_amlKhovH2_0),.clk(gclk));
	jdff dff_B_ccDsk3zu6_0(.din(w_dff_B_amlKhovH2_0),.dout(w_dff_B_ccDsk3zu6_0),.clk(gclk));
	jdff dff_B_hn76hPMW8_0(.din(w_dff_B_ccDsk3zu6_0),.dout(w_dff_B_hn76hPMW8_0),.clk(gclk));
	jdff dff_B_0HX4qyA17_0(.din(w_dff_B_hn76hPMW8_0),.dout(w_dff_B_0HX4qyA17_0),.clk(gclk));
	jdff dff_B_wbCmYHaw6_0(.din(w_dff_B_0HX4qyA17_0),.dout(w_dff_B_wbCmYHaw6_0),.clk(gclk));
	jdff dff_B_BObX65gH8_0(.din(w_dff_B_wbCmYHaw6_0),.dout(w_dff_B_BObX65gH8_0),.clk(gclk));
	jdff dff_B_Rv7rYFht8_0(.din(w_dff_B_BObX65gH8_0),.dout(w_dff_B_Rv7rYFht8_0),.clk(gclk));
	jdff dff_B_4eeXoA0X8_0(.din(w_dff_B_Rv7rYFht8_0),.dout(w_dff_B_4eeXoA0X8_0),.clk(gclk));
	jdff dff_B_OA0MvQRM5_0(.din(w_dff_B_4eeXoA0X8_0),.dout(w_dff_B_OA0MvQRM5_0),.clk(gclk));
	jdff dff_B_qvNlr5RR8_0(.din(w_dff_B_OA0MvQRM5_0),.dout(w_dff_B_qvNlr5RR8_0),.clk(gclk));
	jdff dff_B_CGoMiKOQ9_0(.din(w_dff_B_qvNlr5RR8_0),.dout(w_dff_B_CGoMiKOQ9_0),.clk(gclk));
	jdff dff_B_YEdl7OfL6_0(.din(w_dff_B_CGoMiKOQ9_0),.dout(w_dff_B_YEdl7OfL6_0),.clk(gclk));
	jdff dff_B_yp8qlzjU5_0(.din(w_dff_B_YEdl7OfL6_0),.dout(w_dff_B_yp8qlzjU5_0),.clk(gclk));
	jdff dff_B_YQtkHUAk7_0(.din(w_dff_B_yp8qlzjU5_0),.dout(w_dff_B_YQtkHUAk7_0),.clk(gclk));
	jdff dff_B_Z9IXGwA60_0(.din(w_dff_B_YQtkHUAk7_0),.dout(w_dff_B_Z9IXGwA60_0),.clk(gclk));
	jdff dff_B_ipqgx8Tu0_0(.din(w_dff_B_Z9IXGwA60_0),.dout(w_dff_B_ipqgx8Tu0_0),.clk(gclk));
	jdff dff_B_Oc5FpvzU5_0(.din(w_dff_B_ipqgx8Tu0_0),.dout(w_dff_B_Oc5FpvzU5_0),.clk(gclk));
	jdff dff_B_613TrTLX7_2(.din(G106),.dout(w_dff_B_613TrTLX7_2),.clk(gclk));
	jdff dff_B_fVB9cpGC4_1(.din(n1269),.dout(w_dff_B_fVB9cpGC4_1),.clk(gclk));
	jdff dff_B_5kW2X1Jt1_1(.din(w_dff_B_fVB9cpGC4_1),.dout(w_dff_B_5kW2X1Jt1_1),.clk(gclk));
	jdff dff_A_vmu3grkC7_0(.dout(w_n797_6[0]),.din(w_dff_A_vmu3grkC7_0),.clk(gclk));
	jdff dff_A_P0qOsKlY4_0(.dout(w_dff_A_vmu3grkC7_0),.din(w_dff_A_P0qOsKlY4_0),.clk(gclk));
	jdff dff_A_DXKRFzAL8_0(.dout(w_dff_A_P0qOsKlY4_0),.din(w_dff_A_DXKRFzAL8_0),.clk(gclk));
	jdff dff_A_CyFPFsgZ5_0(.dout(w_dff_A_DXKRFzAL8_0),.din(w_dff_A_CyFPFsgZ5_0),.clk(gclk));
	jdff dff_A_Ak71Hu3n0_0(.dout(w_dff_A_CyFPFsgZ5_0),.din(w_dff_A_Ak71Hu3n0_0),.clk(gclk));
	jdff dff_A_1cpvF5ce9_0(.dout(w_dff_A_Ak71Hu3n0_0),.din(w_dff_A_1cpvF5ce9_0),.clk(gclk));
	jdff dff_A_mWPLGSTW8_0(.dout(w_dff_A_1cpvF5ce9_0),.din(w_dff_A_mWPLGSTW8_0),.clk(gclk));
	jdff dff_A_LYZ5Ozx56_0(.dout(w_dff_A_mWPLGSTW8_0),.din(w_dff_A_LYZ5Ozx56_0),.clk(gclk));
	jdff dff_A_N8kS113w0_0(.dout(w_dff_A_LYZ5Ozx56_0),.din(w_dff_A_N8kS113w0_0),.clk(gclk));
	jdff dff_A_Tz8aNJD11_0(.dout(w_dff_A_N8kS113w0_0),.din(w_dff_A_Tz8aNJD11_0),.clk(gclk));
	jdff dff_A_msNELFM06_0(.dout(w_dff_A_Tz8aNJD11_0),.din(w_dff_A_msNELFM06_0),.clk(gclk));
	jdff dff_A_gYhWE2PL5_0(.dout(w_dff_A_msNELFM06_0),.din(w_dff_A_gYhWE2PL5_0),.clk(gclk));
	jdff dff_A_ZOR8hdyJ7_0(.dout(w_dff_A_gYhWE2PL5_0),.din(w_dff_A_ZOR8hdyJ7_0),.clk(gclk));
	jdff dff_A_swTQvqRQ1_0(.dout(w_dff_A_ZOR8hdyJ7_0),.din(w_dff_A_swTQvqRQ1_0),.clk(gclk));
	jdff dff_A_UMTYZDQ84_0(.dout(w_dff_A_swTQvqRQ1_0),.din(w_dff_A_UMTYZDQ84_0),.clk(gclk));
	jdff dff_A_8dg1W2673_0(.dout(w_dff_A_UMTYZDQ84_0),.din(w_dff_A_8dg1W2673_0),.clk(gclk));
	jdff dff_A_3nVv4tEd8_0(.dout(w_dff_A_8dg1W2673_0),.din(w_dff_A_3nVv4tEd8_0),.clk(gclk));
	jdff dff_A_eiblXQ9W4_0(.dout(w_dff_A_3nVv4tEd8_0),.din(w_dff_A_eiblXQ9W4_0),.clk(gclk));
	jdff dff_A_Klmtffqm4_0(.dout(w_dff_A_eiblXQ9W4_0),.din(w_dff_A_Klmtffqm4_0),.clk(gclk));
	jdff dff_A_e2azE1u77_0(.dout(w_dff_A_Klmtffqm4_0),.din(w_dff_A_e2azE1u77_0),.clk(gclk));
	jdff dff_A_ilKoLCXX7_2(.dout(w_n797_6[2]),.din(w_dff_A_ilKoLCXX7_2),.clk(gclk));
	jdff dff_A_j9wGIjuJ3_2(.dout(w_dff_A_ilKoLCXX7_2),.din(w_dff_A_j9wGIjuJ3_2),.clk(gclk));
	jdff dff_A_iv4jWVui0_2(.dout(w_dff_A_j9wGIjuJ3_2),.din(w_dff_A_iv4jWVui0_2),.clk(gclk));
	jdff dff_A_slBwO6yM4_2(.dout(w_dff_A_iv4jWVui0_2),.din(w_dff_A_slBwO6yM4_2),.clk(gclk));
	jdff dff_A_m865teEJ0_2(.dout(w_dff_A_slBwO6yM4_2),.din(w_dff_A_m865teEJ0_2),.clk(gclk));
	jdff dff_A_cCAvu9o55_2(.dout(w_dff_A_m865teEJ0_2),.din(w_dff_A_cCAvu9o55_2),.clk(gclk));
	jdff dff_A_vz4vnveJ1_2(.dout(w_dff_A_cCAvu9o55_2),.din(w_dff_A_vz4vnveJ1_2),.clk(gclk));
	jdff dff_A_ndDbO4cl5_2(.dout(w_dff_A_vz4vnveJ1_2),.din(w_dff_A_ndDbO4cl5_2),.clk(gclk));
	jdff dff_A_hPePvWMc1_2(.dout(w_dff_A_ndDbO4cl5_2),.din(w_dff_A_hPePvWMc1_2),.clk(gclk));
	jdff dff_A_PBISrbJt7_2(.dout(w_dff_A_hPePvWMc1_2),.din(w_dff_A_PBISrbJt7_2),.clk(gclk));
	jdff dff_A_yraG014I1_2(.dout(w_dff_A_PBISrbJt7_2),.din(w_dff_A_yraG014I1_2),.clk(gclk));
	jdff dff_A_VTL4K4AN2_0(.dout(w_G4088_6[0]),.din(w_dff_A_VTL4K4AN2_0),.clk(gclk));
	jdff dff_A_cZycAh8e0_0(.dout(w_dff_A_VTL4K4AN2_0),.din(w_dff_A_cZycAh8e0_0),.clk(gclk));
	jdff dff_A_L2OUdAyE3_0(.dout(w_dff_A_cZycAh8e0_0),.din(w_dff_A_L2OUdAyE3_0),.clk(gclk));
	jdff dff_A_FHyPy2w78_0(.dout(w_dff_A_L2OUdAyE3_0),.din(w_dff_A_FHyPy2w78_0),.clk(gclk));
	jdff dff_A_H9OFNDI03_0(.dout(w_dff_A_FHyPy2w78_0),.din(w_dff_A_H9OFNDI03_0),.clk(gclk));
	jdff dff_A_6p5mLKqQ5_0(.dout(w_dff_A_H9OFNDI03_0),.din(w_dff_A_6p5mLKqQ5_0),.clk(gclk));
	jdff dff_A_XMqXqIrL6_0(.dout(w_dff_A_6p5mLKqQ5_0),.din(w_dff_A_XMqXqIrL6_0),.clk(gclk));
	jdff dff_A_hIqNW8aG6_0(.dout(w_dff_A_XMqXqIrL6_0),.din(w_dff_A_hIqNW8aG6_0),.clk(gclk));
	jdff dff_A_OH0nMXVi0_0(.dout(w_dff_A_hIqNW8aG6_0),.din(w_dff_A_OH0nMXVi0_0),.clk(gclk));
	jdff dff_A_YKE7TXah8_0(.dout(w_dff_A_OH0nMXVi0_0),.din(w_dff_A_YKE7TXah8_0),.clk(gclk));
	jdff dff_A_mRTnXCtn3_0(.dout(w_dff_A_YKE7TXah8_0),.din(w_dff_A_mRTnXCtn3_0),.clk(gclk));
	jdff dff_A_NUax58OZ8_0(.dout(w_dff_A_mRTnXCtn3_0),.din(w_dff_A_NUax58OZ8_0),.clk(gclk));
	jdff dff_A_IXgFBrHy9_0(.dout(w_dff_A_NUax58OZ8_0),.din(w_dff_A_IXgFBrHy9_0),.clk(gclk));
	jdff dff_A_ykhlCQX31_0(.dout(w_dff_A_IXgFBrHy9_0),.din(w_dff_A_ykhlCQX31_0),.clk(gclk));
	jdff dff_A_5aeUg1Co1_0(.dout(w_dff_A_ykhlCQX31_0),.din(w_dff_A_5aeUg1Co1_0),.clk(gclk));
	jdff dff_A_Yd56h4Yw5_0(.dout(w_dff_A_5aeUg1Co1_0),.din(w_dff_A_Yd56h4Yw5_0),.clk(gclk));
	jdff dff_A_A0EatiEj7_0(.dout(w_dff_A_Yd56h4Yw5_0),.din(w_dff_A_A0EatiEj7_0),.clk(gclk));
	jdff dff_A_2gT5xT5g5_0(.dout(w_dff_A_A0EatiEj7_0),.din(w_dff_A_2gT5xT5g5_0),.clk(gclk));
	jdff dff_A_rqTnFF352_0(.dout(w_dff_A_2gT5xT5g5_0),.din(w_dff_A_rqTnFF352_0),.clk(gclk));
	jdff dff_A_DnGrOMJs5_0(.dout(w_dff_A_rqTnFF352_0),.din(w_dff_A_DnGrOMJs5_0),.clk(gclk));
	jdff dff_A_mZPRQKzC3_2(.dout(w_G4088_6[2]),.din(w_dff_A_mZPRQKzC3_2),.clk(gclk));
	jdff dff_A_uDSmtvhE7_2(.dout(w_dff_A_mZPRQKzC3_2),.din(w_dff_A_uDSmtvhE7_2),.clk(gclk));
	jdff dff_A_0rz0RcBA5_2(.dout(w_dff_A_uDSmtvhE7_2),.din(w_dff_A_0rz0RcBA5_2),.clk(gclk));
	jdff dff_A_WwdrCMyo0_2(.dout(w_dff_A_0rz0RcBA5_2),.din(w_dff_A_WwdrCMyo0_2),.clk(gclk));
	jdff dff_A_P5KRAUwM4_2(.dout(w_dff_A_WwdrCMyo0_2),.din(w_dff_A_P5KRAUwM4_2),.clk(gclk));
	jdff dff_A_AV0x3rVB6_2(.dout(w_dff_A_P5KRAUwM4_2),.din(w_dff_A_AV0x3rVB6_2),.clk(gclk));
	jdff dff_A_uQ4ODTvv1_2(.dout(w_dff_A_AV0x3rVB6_2),.din(w_dff_A_uQ4ODTvv1_2),.clk(gclk));
	jdff dff_A_zep5KxRb6_2(.dout(w_dff_A_uQ4ODTvv1_2),.din(w_dff_A_zep5KxRb6_2),.clk(gclk));
	jdff dff_A_ldWFV7vf9_2(.dout(w_dff_A_zep5KxRb6_2),.din(w_dff_A_ldWFV7vf9_2),.clk(gclk));
	jdff dff_A_NZMNoHdR2_2(.dout(w_dff_A_ldWFV7vf9_2),.din(w_dff_A_NZMNoHdR2_2),.clk(gclk));
	jdff dff_A_m3suCFgq3_2(.dout(w_dff_A_NZMNoHdR2_2),.din(w_dff_A_m3suCFgq3_2),.clk(gclk));
	jdff dff_A_n8vnFEGM9_2(.dout(w_dff_A_m3suCFgq3_2),.din(w_dff_A_n8vnFEGM9_2),.clk(gclk));
	jdff dff_A_5gIW36ZP4_2(.dout(w_dff_A_n8vnFEGM9_2),.din(w_dff_A_5gIW36ZP4_2),.clk(gclk));
	jdff dff_A_wDrieCip9_2(.dout(w_dff_A_5gIW36ZP4_2),.din(w_dff_A_wDrieCip9_2),.clk(gclk));
	jdff dff_B_26vXIsBq6_0(.din(n1286),.dout(w_dff_B_26vXIsBq6_0),.clk(gclk));
	jdff dff_B_237LmwaP1_0(.din(w_dff_B_26vXIsBq6_0),.dout(w_dff_B_237LmwaP1_0),.clk(gclk));
	jdff dff_B_HYqnMS4b3_0(.din(w_dff_B_237LmwaP1_0),.dout(w_dff_B_HYqnMS4b3_0),.clk(gclk));
	jdff dff_B_KIlfmhqN7_0(.din(w_dff_B_HYqnMS4b3_0),.dout(w_dff_B_KIlfmhqN7_0),.clk(gclk));
	jdff dff_B_b0aBPuSw9_0(.din(w_dff_B_KIlfmhqN7_0),.dout(w_dff_B_b0aBPuSw9_0),.clk(gclk));
	jdff dff_B_Q9E1as2H0_0(.din(w_dff_B_b0aBPuSw9_0),.dout(w_dff_B_Q9E1as2H0_0),.clk(gclk));
	jdff dff_B_melxdjnz5_0(.din(w_dff_B_Q9E1as2H0_0),.dout(w_dff_B_melxdjnz5_0),.clk(gclk));
	jdff dff_B_NvLChvnn6_0(.din(w_dff_B_melxdjnz5_0),.dout(w_dff_B_NvLChvnn6_0),.clk(gclk));
	jdff dff_B_X4ZlOaTY1_0(.din(w_dff_B_NvLChvnn6_0),.dout(w_dff_B_X4ZlOaTY1_0),.clk(gclk));
	jdff dff_B_tybX5DEv3_0(.din(w_dff_B_X4ZlOaTY1_0),.dout(w_dff_B_tybX5DEv3_0),.clk(gclk));
	jdff dff_B_DqusuIoh6_0(.din(w_dff_B_tybX5DEv3_0),.dout(w_dff_B_DqusuIoh6_0),.clk(gclk));
	jdff dff_B_by69jzI17_0(.din(w_dff_B_DqusuIoh6_0),.dout(w_dff_B_by69jzI17_0),.clk(gclk));
	jdff dff_B_nvGFCjNw2_0(.din(w_dff_B_by69jzI17_0),.dout(w_dff_B_nvGFCjNw2_0),.clk(gclk));
	jdff dff_B_OVYSqZTJ5_0(.din(w_dff_B_nvGFCjNw2_0),.dout(w_dff_B_OVYSqZTJ5_0),.clk(gclk));
	jdff dff_B_JVYlG0v43_0(.din(w_dff_B_OVYSqZTJ5_0),.dout(w_dff_B_JVYlG0v43_0),.clk(gclk));
	jdff dff_B_4vBj07Vh5_0(.din(w_dff_B_JVYlG0v43_0),.dout(w_dff_B_4vBj07Vh5_0),.clk(gclk));
	jdff dff_B_2YsL8ecb2_0(.din(w_dff_B_4vBj07Vh5_0),.dout(w_dff_B_2YsL8ecb2_0),.clk(gclk));
	jdff dff_B_XRI0FZX86_0(.din(w_dff_B_2YsL8ecb2_0),.dout(w_dff_B_XRI0FZX86_0),.clk(gclk));
	jdff dff_B_0mBTJR4Q8_0(.din(w_dff_B_XRI0FZX86_0),.dout(w_dff_B_0mBTJR4Q8_0),.clk(gclk));
	jdff dff_B_ucBX0RAq0_0(.din(w_dff_B_0mBTJR4Q8_0),.dout(w_dff_B_ucBX0RAq0_0),.clk(gclk));
	jdff dff_B_Kldu5qHO6_1(.din(n1278),.dout(w_dff_B_Kldu5qHO6_1),.clk(gclk));
	jdff dff_B_gocFImUT3_1(.din(w_dff_B_Kldu5qHO6_1),.dout(w_dff_B_gocFImUT3_1),.clk(gclk));
	jdff dff_A_fW0wnGPG7_1(.dout(w_n797_5[1]),.din(w_dff_A_fW0wnGPG7_1),.clk(gclk));
	jdff dff_A_c2JOarfZ8_1(.dout(w_dff_A_fW0wnGPG7_1),.din(w_dff_A_c2JOarfZ8_1),.clk(gclk));
	jdff dff_A_f4wIRi5n4_1(.dout(w_dff_A_c2JOarfZ8_1),.din(w_dff_A_f4wIRi5n4_1),.clk(gclk));
	jdff dff_A_G7U2y4mg0_1(.dout(w_dff_A_f4wIRi5n4_1),.din(w_dff_A_G7U2y4mg0_1),.clk(gclk));
	jdff dff_A_eb5TBan76_1(.dout(w_dff_A_G7U2y4mg0_1),.din(w_dff_A_eb5TBan76_1),.clk(gclk));
	jdff dff_A_NaHnANhF3_1(.dout(w_dff_A_eb5TBan76_1),.din(w_dff_A_NaHnANhF3_1),.clk(gclk));
	jdff dff_A_AEMtDXUi3_1(.dout(w_dff_A_NaHnANhF3_1),.din(w_dff_A_AEMtDXUi3_1),.clk(gclk));
	jdff dff_A_CfQ9ro8Z8_1(.dout(w_dff_A_AEMtDXUi3_1),.din(w_dff_A_CfQ9ro8Z8_1),.clk(gclk));
	jdff dff_A_Kdko3opX3_1(.dout(w_dff_A_CfQ9ro8Z8_1),.din(w_dff_A_Kdko3opX3_1),.clk(gclk));
	jdff dff_A_JaJAejEe3_1(.dout(w_dff_A_Kdko3opX3_1),.din(w_dff_A_JaJAejEe3_1),.clk(gclk));
	jdff dff_A_OHDH7wRu3_1(.dout(w_dff_A_JaJAejEe3_1),.din(w_dff_A_OHDH7wRu3_1),.clk(gclk));
	jdff dff_A_Kx6c7k823_1(.dout(w_dff_A_OHDH7wRu3_1),.din(w_dff_A_Kx6c7k823_1),.clk(gclk));
	jdff dff_A_Epcwrcqr2_1(.dout(w_dff_A_Kx6c7k823_1),.din(w_dff_A_Epcwrcqr2_1),.clk(gclk));
	jdff dff_A_gnIEyZ3w4_1(.dout(w_dff_A_Epcwrcqr2_1),.din(w_dff_A_gnIEyZ3w4_1),.clk(gclk));
	jdff dff_A_FQO6eSNF1_1(.dout(w_dff_A_gnIEyZ3w4_1),.din(w_dff_A_FQO6eSNF1_1),.clk(gclk));
	jdff dff_A_4eWSPZKd2_1(.dout(w_dff_A_FQO6eSNF1_1),.din(w_dff_A_4eWSPZKd2_1),.clk(gclk));
	jdff dff_A_H6tcGR0p0_1(.dout(w_dff_A_4eWSPZKd2_1),.din(w_dff_A_H6tcGR0p0_1),.clk(gclk));
	jdff dff_A_Bc2Y3kNT6_1(.dout(w_dff_A_H6tcGR0p0_1),.din(w_dff_A_Bc2Y3kNT6_1),.clk(gclk));
	jdff dff_A_bxqxQOu92_1(.dout(w_dff_A_Bc2Y3kNT6_1),.din(w_dff_A_bxqxQOu92_1),.clk(gclk));
	jdff dff_A_qr1zaZfW9_1(.dout(w_G4088_5[1]),.din(w_dff_A_qr1zaZfW9_1),.clk(gclk));
	jdff dff_A_ouVm1GKL6_1(.dout(w_dff_A_qr1zaZfW9_1),.din(w_dff_A_ouVm1GKL6_1),.clk(gclk));
	jdff dff_A_Ddie4o278_1(.dout(w_dff_A_ouVm1GKL6_1),.din(w_dff_A_Ddie4o278_1),.clk(gclk));
	jdff dff_A_WnITRA3p3_1(.dout(w_dff_A_Ddie4o278_1),.din(w_dff_A_WnITRA3p3_1),.clk(gclk));
	jdff dff_A_96QPoJ9O4_1(.dout(w_dff_A_WnITRA3p3_1),.din(w_dff_A_96QPoJ9O4_1),.clk(gclk));
	jdff dff_A_6HbkPmG85_1(.dout(w_dff_A_96QPoJ9O4_1),.din(w_dff_A_6HbkPmG85_1),.clk(gclk));
	jdff dff_A_zhxWjCru4_1(.dout(w_dff_A_6HbkPmG85_1),.din(w_dff_A_zhxWjCru4_1),.clk(gclk));
	jdff dff_A_y4arpHE37_1(.dout(w_dff_A_zhxWjCru4_1),.din(w_dff_A_y4arpHE37_1),.clk(gclk));
	jdff dff_A_QlFPTUxj5_1(.dout(w_dff_A_y4arpHE37_1),.din(w_dff_A_QlFPTUxj5_1),.clk(gclk));
	jdff dff_A_WIEMXsFY3_1(.dout(w_dff_A_QlFPTUxj5_1),.din(w_dff_A_WIEMXsFY3_1),.clk(gclk));
	jdff dff_A_pDA50E2E5_1(.dout(w_dff_A_WIEMXsFY3_1),.din(w_dff_A_pDA50E2E5_1),.clk(gclk));
	jdff dff_A_8AnJhNNe4_1(.dout(w_dff_A_pDA50E2E5_1),.din(w_dff_A_8AnJhNNe4_1),.clk(gclk));
	jdff dff_A_ReZifjbl4_1(.dout(w_dff_A_8AnJhNNe4_1),.din(w_dff_A_ReZifjbl4_1),.clk(gclk));
	jdff dff_A_d5Cz99bG2_1(.dout(w_dff_A_ReZifjbl4_1),.din(w_dff_A_d5Cz99bG2_1),.clk(gclk));
	jdff dff_A_9ZZjS1ph8_1(.dout(w_dff_A_d5Cz99bG2_1),.din(w_dff_A_9ZZjS1ph8_1),.clk(gclk));
	jdff dff_A_lH7F1bdL0_1(.dout(w_dff_A_9ZZjS1ph8_1),.din(w_dff_A_lH7F1bdL0_1),.clk(gclk));
	jdff dff_A_oOFGgjiW7_1(.dout(w_dff_A_lH7F1bdL0_1),.din(w_dff_A_oOFGgjiW7_1),.clk(gclk));
	jdff dff_A_nrZt1lOM6_1(.dout(w_dff_A_oOFGgjiW7_1),.din(w_dff_A_nrZt1lOM6_1),.clk(gclk));
	jdff dff_A_cNzuEArp5_1(.dout(w_dff_A_nrZt1lOM6_1),.din(w_dff_A_cNzuEArp5_1),.clk(gclk));
	jdff dff_B_7UjudSZW9_0(.din(n1295),.dout(w_dff_B_7UjudSZW9_0),.clk(gclk));
	jdff dff_B_DcadDWTU5_0(.din(w_dff_B_7UjudSZW9_0),.dout(w_dff_B_DcadDWTU5_0),.clk(gclk));
	jdff dff_B_gX3TpLfj4_0(.din(w_dff_B_DcadDWTU5_0),.dout(w_dff_B_gX3TpLfj4_0),.clk(gclk));
	jdff dff_B_Vo5jpYLr7_0(.din(w_dff_B_gX3TpLfj4_0),.dout(w_dff_B_Vo5jpYLr7_0),.clk(gclk));
	jdff dff_B_tOna3Ym00_0(.din(w_dff_B_Vo5jpYLr7_0),.dout(w_dff_B_tOna3Ym00_0),.clk(gclk));
	jdff dff_B_tgNBYLqh4_0(.din(w_dff_B_tOna3Ym00_0),.dout(w_dff_B_tgNBYLqh4_0),.clk(gclk));
	jdff dff_B_7yaZaOhd8_0(.din(w_dff_B_tgNBYLqh4_0),.dout(w_dff_B_7yaZaOhd8_0),.clk(gclk));
	jdff dff_B_4vDqfosu3_0(.din(w_dff_B_7yaZaOhd8_0),.dout(w_dff_B_4vDqfosu3_0),.clk(gclk));
	jdff dff_B_mOLvacjo2_0(.din(w_dff_B_4vDqfosu3_0),.dout(w_dff_B_mOLvacjo2_0),.clk(gclk));
	jdff dff_B_2PpFbc1B8_0(.din(w_dff_B_mOLvacjo2_0),.dout(w_dff_B_2PpFbc1B8_0),.clk(gclk));
	jdff dff_B_WE21cq7c4_0(.din(w_dff_B_2PpFbc1B8_0),.dout(w_dff_B_WE21cq7c4_0),.clk(gclk));
	jdff dff_B_VflmCJ1O8_0(.din(w_dff_B_WE21cq7c4_0),.dout(w_dff_B_VflmCJ1O8_0),.clk(gclk));
	jdff dff_B_t6KdXIAc2_0(.din(w_dff_B_VflmCJ1O8_0),.dout(w_dff_B_t6KdXIAc2_0),.clk(gclk));
	jdff dff_B_Ea27ydjA8_0(.din(w_dff_B_t6KdXIAc2_0),.dout(w_dff_B_Ea27ydjA8_0),.clk(gclk));
	jdff dff_B_8mtSHyKK6_0(.din(w_dff_B_Ea27ydjA8_0),.dout(w_dff_B_8mtSHyKK6_0),.clk(gclk));
	jdff dff_B_VT34JV8y1_0(.din(w_dff_B_8mtSHyKK6_0),.dout(w_dff_B_VT34JV8y1_0),.clk(gclk));
	jdff dff_B_oZPXF36v3_0(.din(w_dff_B_VT34JV8y1_0),.dout(w_dff_B_oZPXF36v3_0),.clk(gclk));
	jdff dff_B_8pkK5WnP2_0(.din(w_dff_B_oZPXF36v3_0),.dout(w_dff_B_8pkK5WnP2_0),.clk(gclk));
	jdff dff_B_4ZDBi9CO4_0(.din(w_dff_B_8pkK5WnP2_0),.dout(w_dff_B_4ZDBi9CO4_0),.clk(gclk));
	jdff dff_B_ckn15Wxm8_0(.din(w_dff_B_4ZDBi9CO4_0),.dout(w_dff_B_ckn15Wxm8_0),.clk(gclk));
	jdff dff_B_0D6r4phK0_1(.din(n1288),.dout(w_dff_B_0D6r4phK0_1),.clk(gclk));
	jdff dff_A_F6kEEoLb0_2(.dout(w_n800_2[2]),.din(w_dff_A_F6kEEoLb0_2),.clk(gclk));
	jdff dff_B_vp73fETp6_0(.din(n1306),.dout(w_dff_B_vp73fETp6_0),.clk(gclk));
	jdff dff_B_tLVzxb7o8_0(.din(w_dff_B_vp73fETp6_0),.dout(w_dff_B_tLVzxb7o8_0),.clk(gclk));
	jdff dff_B_LnGzdbko1_0(.din(w_dff_B_tLVzxb7o8_0),.dout(w_dff_B_LnGzdbko1_0),.clk(gclk));
	jdff dff_B_OJeBpcXP6_0(.din(w_dff_B_LnGzdbko1_0),.dout(w_dff_B_OJeBpcXP6_0),.clk(gclk));
	jdff dff_B_ndmMawgf5_0(.din(w_dff_B_OJeBpcXP6_0),.dout(w_dff_B_ndmMawgf5_0),.clk(gclk));
	jdff dff_B_5LIcaxSZ6_0(.din(w_dff_B_ndmMawgf5_0),.dout(w_dff_B_5LIcaxSZ6_0),.clk(gclk));
	jdff dff_B_vjChEcSU9_0(.din(w_dff_B_5LIcaxSZ6_0),.dout(w_dff_B_vjChEcSU9_0),.clk(gclk));
	jdff dff_B_9LRB2zkL8_0(.din(w_dff_B_vjChEcSU9_0),.dout(w_dff_B_9LRB2zkL8_0),.clk(gclk));
	jdff dff_B_pGcqzuNM2_0(.din(w_dff_B_9LRB2zkL8_0),.dout(w_dff_B_pGcqzuNM2_0),.clk(gclk));
	jdff dff_B_CPZiW7jH9_0(.din(w_dff_B_pGcqzuNM2_0),.dout(w_dff_B_CPZiW7jH9_0),.clk(gclk));
	jdff dff_B_lcrO5USL6_0(.din(w_dff_B_CPZiW7jH9_0),.dout(w_dff_B_lcrO5USL6_0),.clk(gclk));
	jdff dff_B_drPAWo4y3_0(.din(w_dff_B_lcrO5USL6_0),.dout(w_dff_B_drPAWo4y3_0),.clk(gclk));
	jdff dff_B_uZW28TeO5_0(.din(w_dff_B_drPAWo4y3_0),.dout(w_dff_B_uZW28TeO5_0),.clk(gclk));
	jdff dff_B_L9wP2SIE6_0(.din(w_dff_B_uZW28TeO5_0),.dout(w_dff_B_L9wP2SIE6_0),.clk(gclk));
	jdff dff_B_6B1BSFVf9_0(.din(w_dff_B_L9wP2SIE6_0),.dout(w_dff_B_6B1BSFVf9_0),.clk(gclk));
	jdff dff_B_8LweTrcT8_0(.din(w_dff_B_6B1BSFVf9_0),.dout(w_dff_B_8LweTrcT8_0),.clk(gclk));
	jdff dff_B_zpWxDfUm7_0(.din(w_dff_B_8LweTrcT8_0),.dout(w_dff_B_zpWxDfUm7_0),.clk(gclk));
	jdff dff_B_ovcS07R84_0(.din(w_dff_B_zpWxDfUm7_0),.dout(w_dff_B_ovcS07R84_0),.clk(gclk));
	jdff dff_B_ZPD2HFVt2_0(.din(w_dff_B_ovcS07R84_0),.dout(w_dff_B_ZPD2HFVt2_0),.clk(gclk));
	jdff dff_B_gnu0io0Y0_1(.din(n1298),.dout(w_dff_B_gnu0io0Y0_1),.clk(gclk));
	jdff dff_B_Mguj03XS6_1(.din(w_dff_B_gnu0io0Y0_1),.dout(w_dff_B_Mguj03XS6_1),.clk(gclk));
	jdff dff_B_Y0iBS1MF6_1(.din(w_dff_B_Mguj03XS6_1),.dout(w_dff_B_Y0iBS1MF6_1),.clk(gclk));
	jdff dff_A_c8Kmh86T8_0(.dout(w_n797_4[0]),.din(w_dff_A_c8Kmh86T8_0),.clk(gclk));
	jdff dff_A_mcKseCPZ0_0(.dout(w_dff_A_c8Kmh86T8_0),.din(w_dff_A_mcKseCPZ0_0),.clk(gclk));
	jdff dff_A_gzFjyGFk8_0(.dout(w_dff_A_mcKseCPZ0_0),.din(w_dff_A_gzFjyGFk8_0),.clk(gclk));
	jdff dff_A_aTbMuSXF5_0(.dout(w_dff_A_gzFjyGFk8_0),.din(w_dff_A_aTbMuSXF5_0),.clk(gclk));
	jdff dff_A_dkModUv92_0(.dout(w_dff_A_aTbMuSXF5_0),.din(w_dff_A_dkModUv92_0),.clk(gclk));
	jdff dff_A_mmi0TJ2l1_0(.dout(w_dff_A_dkModUv92_0),.din(w_dff_A_mmi0TJ2l1_0),.clk(gclk));
	jdff dff_A_ZzFSyu8U7_0(.dout(w_dff_A_mmi0TJ2l1_0),.din(w_dff_A_ZzFSyu8U7_0),.clk(gclk));
	jdff dff_A_xJs2sFMc6_0(.dout(w_dff_A_ZzFSyu8U7_0),.din(w_dff_A_xJs2sFMc6_0),.clk(gclk));
	jdff dff_A_6TiupRoT3_0(.dout(w_dff_A_xJs2sFMc6_0),.din(w_dff_A_6TiupRoT3_0),.clk(gclk));
	jdff dff_A_hP8Luy1H1_0(.dout(w_dff_A_6TiupRoT3_0),.din(w_dff_A_hP8Luy1H1_0),.clk(gclk));
	jdff dff_A_WTS0IMSz4_0(.dout(w_dff_A_hP8Luy1H1_0),.din(w_dff_A_WTS0IMSz4_0),.clk(gclk));
	jdff dff_A_t9DcpFOp2_0(.dout(w_dff_A_WTS0IMSz4_0),.din(w_dff_A_t9DcpFOp2_0),.clk(gclk));
	jdff dff_A_4fcaJOul6_0(.dout(w_dff_A_t9DcpFOp2_0),.din(w_dff_A_4fcaJOul6_0),.clk(gclk));
	jdff dff_A_yxrj8M9C6_0(.dout(w_dff_A_4fcaJOul6_0),.din(w_dff_A_yxrj8M9C6_0),.clk(gclk));
	jdff dff_A_JQAb2F3x3_0(.dout(w_dff_A_yxrj8M9C6_0),.din(w_dff_A_JQAb2F3x3_0),.clk(gclk));
	jdff dff_A_OE3fPINj8_0(.dout(w_dff_A_JQAb2F3x3_0),.din(w_dff_A_OE3fPINj8_0),.clk(gclk));
	jdff dff_A_D21QqSyu6_0(.dout(w_dff_A_OE3fPINj8_0),.din(w_dff_A_D21QqSyu6_0),.clk(gclk));
	jdff dff_A_0PAbTmFU7_0(.dout(w_dff_A_D21QqSyu6_0),.din(w_dff_A_0PAbTmFU7_0),.clk(gclk));
	jdff dff_A_l5VQZLGs8_2(.dout(w_n797_4[2]),.din(w_dff_A_l5VQZLGs8_2),.clk(gclk));
	jdff dff_A_Wi8FS5Qf4_2(.dout(w_dff_A_l5VQZLGs8_2),.din(w_dff_A_Wi8FS5Qf4_2),.clk(gclk));
	jdff dff_A_MgFTMBNo6_2(.dout(w_dff_A_Wi8FS5Qf4_2),.din(w_dff_A_MgFTMBNo6_2),.clk(gclk));
	jdff dff_A_Zw79KdCA2_2(.dout(w_dff_A_MgFTMBNo6_2),.din(w_dff_A_Zw79KdCA2_2),.clk(gclk));
	jdff dff_A_gMiMV8FR9_2(.dout(w_dff_A_Zw79KdCA2_2),.din(w_dff_A_gMiMV8FR9_2),.clk(gclk));
	jdff dff_A_ix6r8cx42_2(.dout(w_dff_A_gMiMV8FR9_2),.din(w_dff_A_ix6r8cx42_2),.clk(gclk));
	jdff dff_A_8RyrBXgn9_2(.dout(w_dff_A_ix6r8cx42_2),.din(w_dff_A_8RyrBXgn9_2),.clk(gclk));
	jdff dff_A_4KYwUy5x1_2(.dout(w_dff_A_8RyrBXgn9_2),.din(w_dff_A_4KYwUy5x1_2),.clk(gclk));
	jdff dff_A_Dmet1Hgc7_2(.dout(w_dff_A_4KYwUy5x1_2),.din(w_dff_A_Dmet1Hgc7_2),.clk(gclk));
	jdff dff_A_MAyHAZ0z1_2(.dout(w_dff_A_Dmet1Hgc7_2),.din(w_dff_A_MAyHAZ0z1_2),.clk(gclk));
	jdff dff_A_b185gkc21_2(.dout(w_dff_A_MAyHAZ0z1_2),.din(w_dff_A_b185gkc21_2),.clk(gclk));
	jdff dff_A_aTCTlvJy2_2(.dout(w_dff_A_b185gkc21_2),.din(w_dff_A_aTCTlvJy2_2),.clk(gclk));
	jdff dff_A_2RMoAcWF9_2(.dout(w_dff_A_aTCTlvJy2_2),.din(w_dff_A_2RMoAcWF9_2),.clk(gclk));
	jdff dff_A_PiGyPitN2_2(.dout(w_dff_A_2RMoAcWF9_2),.din(w_dff_A_PiGyPitN2_2),.clk(gclk));
	jdff dff_A_MHh1cXZs6_2(.dout(w_dff_A_PiGyPitN2_2),.din(w_dff_A_MHh1cXZs6_2),.clk(gclk));
	jdff dff_A_l4R2yFE22_2(.dout(w_dff_A_MHh1cXZs6_2),.din(w_dff_A_l4R2yFE22_2),.clk(gclk));
	jdff dff_A_PJVQDKlL0_2(.dout(w_dff_A_l4R2yFE22_2),.din(w_dff_A_PJVQDKlL0_2),.clk(gclk));
	jdff dff_A_C4ifFUPk4_2(.dout(w_dff_A_PJVQDKlL0_2),.din(w_dff_A_C4ifFUPk4_2),.clk(gclk));
	jdff dff_A_qOvYg6Ov9_2(.dout(w_dff_A_C4ifFUPk4_2),.din(w_dff_A_qOvYg6Ov9_2),.clk(gclk));
	jdff dff_A_qESsbqie3_0(.dout(w_G4088_4[0]),.din(w_dff_A_qESsbqie3_0),.clk(gclk));
	jdff dff_A_YJTwBiIT3_0(.dout(w_dff_A_qESsbqie3_0),.din(w_dff_A_YJTwBiIT3_0),.clk(gclk));
	jdff dff_A_a3otgkqM4_0(.dout(w_dff_A_YJTwBiIT3_0),.din(w_dff_A_a3otgkqM4_0),.clk(gclk));
	jdff dff_A_fL0tGpx44_0(.dout(w_dff_A_a3otgkqM4_0),.din(w_dff_A_fL0tGpx44_0),.clk(gclk));
	jdff dff_A_Q93y5Iik5_0(.dout(w_dff_A_fL0tGpx44_0),.din(w_dff_A_Q93y5Iik5_0),.clk(gclk));
	jdff dff_A_45hqZKf57_0(.dout(w_dff_A_Q93y5Iik5_0),.din(w_dff_A_45hqZKf57_0),.clk(gclk));
	jdff dff_A_dQRPsQqf2_0(.dout(w_dff_A_45hqZKf57_0),.din(w_dff_A_dQRPsQqf2_0),.clk(gclk));
	jdff dff_A_OEbN8EXk5_0(.dout(w_dff_A_dQRPsQqf2_0),.din(w_dff_A_OEbN8EXk5_0),.clk(gclk));
	jdff dff_A_DRJflWKr9_0(.dout(w_dff_A_OEbN8EXk5_0),.din(w_dff_A_DRJflWKr9_0),.clk(gclk));
	jdff dff_A_gSLcyW3V2_0(.dout(w_dff_A_DRJflWKr9_0),.din(w_dff_A_gSLcyW3V2_0),.clk(gclk));
	jdff dff_A_Z3HRJwEi0_0(.dout(w_dff_A_gSLcyW3V2_0),.din(w_dff_A_Z3HRJwEi0_0),.clk(gclk));
	jdff dff_A_M5wqTL3w1_0(.dout(w_dff_A_Z3HRJwEi0_0),.din(w_dff_A_M5wqTL3w1_0),.clk(gclk));
	jdff dff_A_HyEHA1b12_0(.dout(w_dff_A_M5wqTL3w1_0),.din(w_dff_A_HyEHA1b12_0),.clk(gclk));
	jdff dff_A_z966KQDq9_0(.dout(w_dff_A_HyEHA1b12_0),.din(w_dff_A_z966KQDq9_0),.clk(gclk));
	jdff dff_A_Fa0uN8os5_0(.dout(w_dff_A_z966KQDq9_0),.din(w_dff_A_Fa0uN8os5_0),.clk(gclk));
	jdff dff_A_vH4D8Mmr4_0(.dout(w_dff_A_Fa0uN8os5_0),.din(w_dff_A_vH4D8Mmr4_0),.clk(gclk));
	jdff dff_A_n56Cg8U79_0(.dout(w_dff_A_vH4D8Mmr4_0),.din(w_dff_A_n56Cg8U79_0),.clk(gclk));
	jdff dff_A_g60qJbka0_2(.dout(w_G4088_4[2]),.din(w_dff_A_g60qJbka0_2),.clk(gclk));
	jdff dff_A_Z7AbxlRT4_2(.dout(w_dff_A_g60qJbka0_2),.din(w_dff_A_Z7AbxlRT4_2),.clk(gclk));
	jdff dff_A_sLlhvxc51_2(.dout(w_dff_A_Z7AbxlRT4_2),.din(w_dff_A_sLlhvxc51_2),.clk(gclk));
	jdff dff_A_nTKTtuIH6_2(.dout(w_dff_A_sLlhvxc51_2),.din(w_dff_A_nTKTtuIH6_2),.clk(gclk));
	jdff dff_A_1LACJbbj5_2(.dout(w_dff_A_nTKTtuIH6_2),.din(w_dff_A_1LACJbbj5_2),.clk(gclk));
	jdff dff_A_tGuooKm99_2(.dout(w_dff_A_1LACJbbj5_2),.din(w_dff_A_tGuooKm99_2),.clk(gclk));
	jdff dff_A_HMeDhRlP1_2(.dout(w_dff_A_tGuooKm99_2),.din(w_dff_A_HMeDhRlP1_2),.clk(gclk));
	jdff dff_A_Z9An5mDf6_2(.dout(w_dff_A_HMeDhRlP1_2),.din(w_dff_A_Z9An5mDf6_2),.clk(gclk));
	jdff dff_A_nwo6rMuK4_2(.dout(w_dff_A_Z9An5mDf6_2),.din(w_dff_A_nwo6rMuK4_2),.clk(gclk));
	jdff dff_A_GIRc0fds5_2(.dout(w_dff_A_nwo6rMuK4_2),.din(w_dff_A_GIRc0fds5_2),.clk(gclk));
	jdff dff_A_WNH877zU8_2(.dout(w_dff_A_GIRc0fds5_2),.din(w_dff_A_WNH877zU8_2),.clk(gclk));
	jdff dff_A_LkUCL5xp3_2(.dout(w_dff_A_WNH877zU8_2),.din(w_dff_A_LkUCL5xp3_2),.clk(gclk));
	jdff dff_A_CotZHC4G3_2(.dout(w_dff_A_LkUCL5xp3_2),.din(w_dff_A_CotZHC4G3_2),.clk(gclk));
	jdff dff_A_ubrXqq9h7_2(.dout(w_dff_A_CotZHC4G3_2),.din(w_dff_A_ubrXqq9h7_2),.clk(gclk));
	jdff dff_A_h6ODVTHe3_2(.dout(w_dff_A_ubrXqq9h7_2),.din(w_dff_A_h6ODVTHe3_2),.clk(gclk));
	jdff dff_A_Rkj2NQzS1_2(.dout(w_dff_A_h6ODVTHe3_2),.din(w_dff_A_Rkj2NQzS1_2),.clk(gclk));
	jdff dff_A_y4MCU1Or5_2(.dout(w_dff_A_Rkj2NQzS1_2),.din(w_dff_A_y4MCU1Or5_2),.clk(gclk));
	jdff dff_A_OGv8jIoD3_2(.dout(w_dff_A_y4MCU1Or5_2),.din(w_dff_A_OGv8jIoD3_2),.clk(gclk));
	jdff dff_A_GLLu1T570_2(.dout(w_dff_A_OGv8jIoD3_2),.din(w_dff_A_GLLu1T570_2),.clk(gclk));
	jdff dff_A_3MTawk6p2_2(.dout(w_dff_A_GLLu1T570_2),.din(w_dff_A_3MTawk6p2_2),.clk(gclk));
	jdff dff_B_sLQnThb07_0(.din(n1315),.dout(w_dff_B_sLQnThb07_0),.clk(gclk));
	jdff dff_B_FpPR17FD1_0(.din(w_dff_B_sLQnThb07_0),.dout(w_dff_B_FpPR17FD1_0),.clk(gclk));
	jdff dff_B_fDzXJuTr2_0(.din(w_dff_B_FpPR17FD1_0),.dout(w_dff_B_fDzXJuTr2_0),.clk(gclk));
	jdff dff_B_clEgHPOm1_0(.din(w_dff_B_fDzXJuTr2_0),.dout(w_dff_B_clEgHPOm1_0),.clk(gclk));
	jdff dff_B_huIMoZ791_0(.din(w_dff_B_clEgHPOm1_0),.dout(w_dff_B_huIMoZ791_0),.clk(gclk));
	jdff dff_B_4T6hSof15_0(.din(w_dff_B_huIMoZ791_0),.dout(w_dff_B_4T6hSof15_0),.clk(gclk));
	jdff dff_B_mP2gaJKY6_0(.din(w_dff_B_4T6hSof15_0),.dout(w_dff_B_mP2gaJKY6_0),.clk(gclk));
	jdff dff_B_ZFDINmTe2_0(.din(w_dff_B_mP2gaJKY6_0),.dout(w_dff_B_ZFDINmTe2_0),.clk(gclk));
	jdff dff_B_2f4Odfvv7_0(.din(w_dff_B_ZFDINmTe2_0),.dout(w_dff_B_2f4Odfvv7_0),.clk(gclk));
	jdff dff_B_1MX9Kp512_0(.din(w_dff_B_2f4Odfvv7_0),.dout(w_dff_B_1MX9Kp512_0),.clk(gclk));
	jdff dff_B_DzZl1J0C9_0(.din(w_dff_B_1MX9Kp512_0),.dout(w_dff_B_DzZl1J0C9_0),.clk(gclk));
	jdff dff_B_uLmsER0w4_0(.din(w_dff_B_DzZl1J0C9_0),.dout(w_dff_B_uLmsER0w4_0),.clk(gclk));
	jdff dff_B_HB9Uenv55_0(.din(w_dff_B_uLmsER0w4_0),.dout(w_dff_B_HB9Uenv55_0),.clk(gclk));
	jdff dff_B_0GPm6Bc90_0(.din(w_dff_B_HB9Uenv55_0),.dout(w_dff_B_0GPm6Bc90_0),.clk(gclk));
	jdff dff_B_99IbGpKN5_0(.din(w_dff_B_0GPm6Bc90_0),.dout(w_dff_B_99IbGpKN5_0),.clk(gclk));
	jdff dff_B_5cShaHcV2_0(.din(w_dff_B_99IbGpKN5_0),.dout(w_dff_B_5cShaHcV2_0),.clk(gclk));
	jdff dff_B_679P78Q55_0(.din(w_dff_B_5cShaHcV2_0),.dout(w_dff_B_679P78Q55_0),.clk(gclk));
	jdff dff_B_5zcaT43A4_0(.din(w_dff_B_679P78Q55_0),.dout(w_dff_B_5zcaT43A4_0),.clk(gclk));
	jdff dff_B_k5gzeLve0_0(.din(w_dff_B_5zcaT43A4_0),.dout(w_dff_B_k5gzeLve0_0),.clk(gclk));
	jdff dff_B_sS6HhTvr8_0(.din(w_dff_B_k5gzeLve0_0),.dout(w_dff_B_sS6HhTvr8_0),.clk(gclk));
	jdff dff_B_BpkAsc1y6_2(.din(G49),.dout(w_dff_B_BpkAsc1y6_2),.clk(gclk));
	jdff dff_B_tnKmZ8XB9_1(.din(n1308),.dout(w_dff_B_tnKmZ8XB9_1),.clk(gclk));
	jdff dff_B_Xq6EIfTl7_1(.din(w_dff_B_tnKmZ8XB9_1),.dout(w_dff_B_Xq6EIfTl7_1),.clk(gclk));
	jdff dff_A_YwCVStrG5_1(.dout(w_n852_5[1]),.din(w_dff_A_YwCVStrG5_1),.clk(gclk));
	jdff dff_A_iqM4HQ2X9_1(.dout(w_dff_A_YwCVStrG5_1),.din(w_dff_A_iqM4HQ2X9_1),.clk(gclk));
	jdff dff_A_3sqNHz3t1_1(.dout(w_dff_A_iqM4HQ2X9_1),.din(w_dff_A_3sqNHz3t1_1),.clk(gclk));
	jdff dff_A_CbzZsDXQ2_1(.dout(w_dff_A_3sqNHz3t1_1),.din(w_dff_A_CbzZsDXQ2_1),.clk(gclk));
	jdff dff_A_eaVJy22C3_1(.dout(w_dff_A_CbzZsDXQ2_1),.din(w_dff_A_eaVJy22C3_1),.clk(gclk));
	jdff dff_A_iQS3qMlv3_1(.dout(w_dff_A_eaVJy22C3_1),.din(w_dff_A_iQS3qMlv3_1),.clk(gclk));
	jdff dff_A_W1kud2fI7_1(.dout(w_dff_A_iQS3qMlv3_1),.din(w_dff_A_W1kud2fI7_1),.clk(gclk));
	jdff dff_A_F0ZOs3nt1_1(.dout(w_dff_A_W1kud2fI7_1),.din(w_dff_A_F0ZOs3nt1_1),.clk(gclk));
	jdff dff_A_8V78MCKm0_1(.dout(w_dff_A_F0ZOs3nt1_1),.din(w_dff_A_8V78MCKm0_1),.clk(gclk));
	jdff dff_A_R51gQHhk2_1(.dout(w_dff_A_8V78MCKm0_1),.din(w_dff_A_R51gQHhk2_1),.clk(gclk));
	jdff dff_A_UIZHmYXx2_1(.dout(w_dff_A_R51gQHhk2_1),.din(w_dff_A_UIZHmYXx2_1),.clk(gclk));
	jdff dff_A_QISS2oXA3_1(.dout(w_dff_A_UIZHmYXx2_1),.din(w_dff_A_QISS2oXA3_1),.clk(gclk));
	jdff dff_A_tBzkUQdT8_1(.dout(w_dff_A_QISS2oXA3_1),.din(w_dff_A_tBzkUQdT8_1),.clk(gclk));
	jdff dff_A_UBf3TArc6_1(.dout(w_dff_A_tBzkUQdT8_1),.din(w_dff_A_UBf3TArc6_1),.clk(gclk));
	jdff dff_A_5h51zdDZ3_1(.dout(w_dff_A_UBf3TArc6_1),.din(w_dff_A_5h51zdDZ3_1),.clk(gclk));
	jdff dff_A_6Lp0Fj9l6_1(.dout(w_dff_A_5h51zdDZ3_1),.din(w_dff_A_6Lp0Fj9l6_1),.clk(gclk));
	jdff dff_A_dzJ10lsn6_1(.dout(w_dff_A_6Lp0Fj9l6_1),.din(w_dff_A_dzJ10lsn6_1),.clk(gclk));
	jdff dff_A_DPVYKORw1_1(.dout(w_dff_A_dzJ10lsn6_1),.din(w_dff_A_DPVYKORw1_1),.clk(gclk));
	jdff dff_A_bn9BiymC4_1(.dout(w_dff_A_DPVYKORw1_1),.din(w_dff_A_bn9BiymC4_1),.clk(gclk));
	jdff dff_A_d0PDyUJm9_2(.dout(w_n852_5[2]),.din(w_dff_A_d0PDyUJm9_2),.clk(gclk));
	jdff dff_A_y2a2Dp8J0_2(.dout(w_dff_A_d0PDyUJm9_2),.din(w_dff_A_y2a2Dp8J0_2),.clk(gclk));
	jdff dff_A_LAJorAAD2_2(.dout(w_dff_A_y2a2Dp8J0_2),.din(w_dff_A_LAJorAAD2_2),.clk(gclk));
	jdff dff_A_vew6i1Ws8_2(.dout(w_dff_A_LAJorAAD2_2),.din(w_dff_A_vew6i1Ws8_2),.clk(gclk));
	jdff dff_A_nsPb19gP9_2(.dout(w_dff_A_vew6i1Ws8_2),.din(w_dff_A_nsPb19gP9_2),.clk(gclk));
	jdff dff_A_DvmywXrd9_2(.dout(w_dff_A_nsPb19gP9_2),.din(w_dff_A_DvmywXrd9_2),.clk(gclk));
	jdff dff_A_qoXdwmNy8_2(.dout(w_dff_A_DvmywXrd9_2),.din(w_dff_A_qoXdwmNy8_2),.clk(gclk));
	jdff dff_A_CISUJWI08_2(.dout(w_dff_A_qoXdwmNy8_2),.din(w_dff_A_CISUJWI08_2),.clk(gclk));
	jdff dff_A_LUfgd2Hd7_2(.dout(w_dff_A_CISUJWI08_2),.din(w_dff_A_LUfgd2Hd7_2),.clk(gclk));
	jdff dff_A_dEneHv9m8_2(.dout(w_dff_A_LUfgd2Hd7_2),.din(w_dff_A_dEneHv9m8_2),.clk(gclk));
	jdff dff_A_i0Yk1vAb5_2(.dout(w_dff_A_dEneHv9m8_2),.din(w_dff_A_i0Yk1vAb5_2),.clk(gclk));
	jdff dff_A_1rX1K71I0_2(.dout(w_dff_A_i0Yk1vAb5_2),.din(w_dff_A_1rX1K71I0_2),.clk(gclk));
	jdff dff_A_LrGycIDG9_2(.dout(w_dff_A_1rX1K71I0_2),.din(w_dff_A_LrGycIDG9_2),.clk(gclk));
	jdff dff_A_Snd94FQK2_2(.dout(w_dff_A_LrGycIDG9_2),.din(w_dff_A_Snd94FQK2_2),.clk(gclk));
	jdff dff_A_om8VqVgx9_2(.dout(w_dff_A_Snd94FQK2_2),.din(w_dff_A_om8VqVgx9_2),.clk(gclk));
	jdff dff_A_Az5eyil72_2(.dout(w_dff_A_om8VqVgx9_2),.din(w_dff_A_Az5eyil72_2),.clk(gclk));
	jdff dff_A_Js4HmcVz2_2(.dout(w_dff_A_Az5eyil72_2),.din(w_dff_A_Js4HmcVz2_2),.clk(gclk));
	jdff dff_A_Q2nWyxKH7_2(.dout(w_dff_A_Js4HmcVz2_2),.din(w_dff_A_Q2nWyxKH7_2),.clk(gclk));
	jdff dff_A_3Je4OfGt1_2(.dout(w_dff_A_Q2nWyxKH7_2),.din(w_dff_A_3Je4OfGt1_2),.clk(gclk));
	jdff dff_A_l7yjVuJE0_2(.dout(w_dff_A_3Je4OfGt1_2),.din(w_dff_A_l7yjVuJE0_2),.clk(gclk));
	jdff dff_A_YoMJhFeU5_1(.dout(w_G4089_5[1]),.din(w_dff_A_YoMJhFeU5_1),.clk(gclk));
	jdff dff_A_udvKaqGj0_1(.dout(w_dff_A_YoMJhFeU5_1),.din(w_dff_A_udvKaqGj0_1),.clk(gclk));
	jdff dff_A_gD303vOn0_1(.dout(w_dff_A_udvKaqGj0_1),.din(w_dff_A_gD303vOn0_1),.clk(gclk));
	jdff dff_A_wB0nvP2l9_1(.dout(w_dff_A_gD303vOn0_1),.din(w_dff_A_wB0nvP2l9_1),.clk(gclk));
	jdff dff_A_qDASnoKV9_1(.dout(w_dff_A_wB0nvP2l9_1),.din(w_dff_A_qDASnoKV9_1),.clk(gclk));
	jdff dff_A_qvhKjY1a3_1(.dout(w_dff_A_qDASnoKV9_1),.din(w_dff_A_qvhKjY1a3_1),.clk(gclk));
	jdff dff_A_xvay0Dri8_1(.dout(w_dff_A_qvhKjY1a3_1),.din(w_dff_A_xvay0Dri8_1),.clk(gclk));
	jdff dff_A_Gzin9HnS2_1(.dout(w_dff_A_xvay0Dri8_1),.din(w_dff_A_Gzin9HnS2_1),.clk(gclk));
	jdff dff_A_BzPsx90L0_1(.dout(w_dff_A_Gzin9HnS2_1),.din(w_dff_A_BzPsx90L0_1),.clk(gclk));
	jdff dff_A_jFyLk3b71_1(.dout(w_dff_A_BzPsx90L0_1),.din(w_dff_A_jFyLk3b71_1),.clk(gclk));
	jdff dff_A_7aNaPJP95_1(.dout(w_dff_A_jFyLk3b71_1),.din(w_dff_A_7aNaPJP95_1),.clk(gclk));
	jdff dff_A_SnlfO4Ny4_1(.dout(w_dff_A_7aNaPJP95_1),.din(w_dff_A_SnlfO4Ny4_1),.clk(gclk));
	jdff dff_A_Wxc2EWao9_1(.dout(w_dff_A_SnlfO4Ny4_1),.din(w_dff_A_Wxc2EWao9_1),.clk(gclk));
	jdff dff_A_vl56YY354_1(.dout(w_dff_A_Wxc2EWao9_1),.din(w_dff_A_vl56YY354_1),.clk(gclk));
	jdff dff_A_yFPcyPHm1_1(.dout(w_dff_A_vl56YY354_1),.din(w_dff_A_yFPcyPHm1_1),.clk(gclk));
	jdff dff_A_E9Ao7VvB8_1(.dout(w_dff_A_yFPcyPHm1_1),.din(w_dff_A_E9Ao7VvB8_1),.clk(gclk));
	jdff dff_A_gocVw8n22_1(.dout(w_dff_A_E9Ao7VvB8_1),.din(w_dff_A_gocVw8n22_1),.clk(gclk));
	jdff dff_A_epruyMLi0_1(.dout(w_dff_A_gocVw8n22_1),.din(w_dff_A_epruyMLi0_1),.clk(gclk));
	jdff dff_A_AZUk2N372_1(.dout(w_dff_A_epruyMLi0_1),.din(w_dff_A_AZUk2N372_1),.clk(gclk));
	jdff dff_A_sSo3SwRo0_2(.dout(w_G4089_5[2]),.din(w_dff_A_sSo3SwRo0_2),.clk(gclk));
	jdff dff_A_9qiF0ob89_2(.dout(w_dff_A_sSo3SwRo0_2),.din(w_dff_A_9qiF0ob89_2),.clk(gclk));
	jdff dff_A_G5sR4Sco4_2(.dout(w_dff_A_9qiF0ob89_2),.din(w_dff_A_G5sR4Sco4_2),.clk(gclk));
	jdff dff_A_Oedmlh5m1_2(.dout(w_dff_A_G5sR4Sco4_2),.din(w_dff_A_Oedmlh5m1_2),.clk(gclk));
	jdff dff_A_7kD2yT968_2(.dout(w_dff_A_Oedmlh5m1_2),.din(w_dff_A_7kD2yT968_2),.clk(gclk));
	jdff dff_A_hbjkuKhH9_2(.dout(w_dff_A_7kD2yT968_2),.din(w_dff_A_hbjkuKhH9_2),.clk(gclk));
	jdff dff_A_1avGh9X24_2(.dout(w_dff_A_hbjkuKhH9_2),.din(w_dff_A_1avGh9X24_2),.clk(gclk));
	jdff dff_A_q9DS2HfD8_2(.dout(w_dff_A_1avGh9X24_2),.din(w_dff_A_q9DS2HfD8_2),.clk(gclk));
	jdff dff_A_KSBaIyKx3_2(.dout(w_dff_A_q9DS2HfD8_2),.din(w_dff_A_KSBaIyKx3_2),.clk(gclk));
	jdff dff_A_00t9mj1C0_2(.dout(w_dff_A_KSBaIyKx3_2),.din(w_dff_A_00t9mj1C0_2),.clk(gclk));
	jdff dff_A_nr47YXuu8_2(.dout(w_dff_A_00t9mj1C0_2),.din(w_dff_A_nr47YXuu8_2),.clk(gclk));
	jdff dff_A_IRWHGHsC2_2(.dout(w_dff_A_nr47YXuu8_2),.din(w_dff_A_IRWHGHsC2_2),.clk(gclk));
	jdff dff_A_2HsNTUVT5_2(.dout(w_dff_A_IRWHGHsC2_2),.din(w_dff_A_2HsNTUVT5_2),.clk(gclk));
	jdff dff_A_hZw2nYKR1_2(.dout(w_dff_A_2HsNTUVT5_2),.din(w_dff_A_hZw2nYKR1_2),.clk(gclk));
	jdff dff_A_ePxzCj0Z4_2(.dout(w_dff_A_hZw2nYKR1_2),.din(w_dff_A_ePxzCj0Z4_2),.clk(gclk));
	jdff dff_A_0Z7jcUqa5_2(.dout(w_dff_A_ePxzCj0Z4_2),.din(w_dff_A_0Z7jcUqa5_2),.clk(gclk));
	jdff dff_A_SwmEI5h61_2(.dout(w_dff_A_0Z7jcUqa5_2),.din(w_dff_A_SwmEI5h61_2),.clk(gclk));
	jdff dff_A_EzcBz4r93_2(.dout(w_dff_A_SwmEI5h61_2),.din(w_dff_A_EzcBz4r93_2),.clk(gclk));
	jdff dff_A_hoBTjbXv9_2(.dout(w_dff_A_EzcBz4r93_2),.din(w_dff_A_hoBTjbXv9_2),.clk(gclk));
	jdff dff_A_4PPCRYOm0_2(.dout(w_dff_A_hoBTjbXv9_2),.din(w_dff_A_4PPCRYOm0_2),.clk(gclk));
	jdff dff_B_YIHEzFLr0_0(.din(n1324),.dout(w_dff_B_YIHEzFLr0_0),.clk(gclk));
	jdff dff_B_jdUK9P8A4_0(.din(w_dff_B_YIHEzFLr0_0),.dout(w_dff_B_jdUK9P8A4_0),.clk(gclk));
	jdff dff_B_8VbUnEOV0_0(.din(w_dff_B_jdUK9P8A4_0),.dout(w_dff_B_8VbUnEOV0_0),.clk(gclk));
	jdff dff_B_g9gjqgJv5_0(.din(w_dff_B_8VbUnEOV0_0),.dout(w_dff_B_g9gjqgJv5_0),.clk(gclk));
	jdff dff_B_iI5WRS1v9_0(.din(w_dff_B_g9gjqgJv5_0),.dout(w_dff_B_iI5WRS1v9_0),.clk(gclk));
	jdff dff_B_6JDFyqZo5_0(.din(w_dff_B_iI5WRS1v9_0),.dout(w_dff_B_6JDFyqZo5_0),.clk(gclk));
	jdff dff_B_GlVtUsFp6_0(.din(w_dff_B_6JDFyqZo5_0),.dout(w_dff_B_GlVtUsFp6_0),.clk(gclk));
	jdff dff_B_8ahMyhzz3_0(.din(w_dff_B_GlVtUsFp6_0),.dout(w_dff_B_8ahMyhzz3_0),.clk(gclk));
	jdff dff_B_mksuzE8m9_0(.din(w_dff_B_8ahMyhzz3_0),.dout(w_dff_B_mksuzE8m9_0),.clk(gclk));
	jdff dff_B_nqkE2MRd7_0(.din(w_dff_B_mksuzE8m9_0),.dout(w_dff_B_nqkE2MRd7_0),.clk(gclk));
	jdff dff_B_1xVD6u4R2_0(.din(w_dff_B_nqkE2MRd7_0),.dout(w_dff_B_1xVD6u4R2_0),.clk(gclk));
	jdff dff_B_MjtRJtDF1_0(.din(w_dff_B_1xVD6u4R2_0),.dout(w_dff_B_MjtRJtDF1_0),.clk(gclk));
	jdff dff_B_ryiqz1h99_0(.din(w_dff_B_MjtRJtDF1_0),.dout(w_dff_B_ryiqz1h99_0),.clk(gclk));
	jdff dff_B_HP1w4vLn7_0(.din(w_dff_B_ryiqz1h99_0),.dout(w_dff_B_HP1w4vLn7_0),.clk(gclk));
	jdff dff_B_sO7Fx42m4_0(.din(w_dff_B_HP1w4vLn7_0),.dout(w_dff_B_sO7Fx42m4_0),.clk(gclk));
	jdff dff_B_M9Muah9E5_0(.din(w_dff_B_sO7Fx42m4_0),.dout(w_dff_B_M9Muah9E5_0),.clk(gclk));
	jdff dff_B_af4HBjBw3_0(.din(w_dff_B_M9Muah9E5_0),.dout(w_dff_B_af4HBjBw3_0),.clk(gclk));
	jdff dff_B_28uQhLBD8_0(.din(w_dff_B_af4HBjBw3_0),.dout(w_dff_B_28uQhLBD8_0),.clk(gclk));
	jdff dff_B_O2kpaOd25_0(.din(w_dff_B_28uQhLBD8_0),.dout(w_dff_B_O2kpaOd25_0),.clk(gclk));
	jdff dff_B_KRwNmUJd6_0(.din(w_dff_B_O2kpaOd25_0),.dout(w_dff_B_KRwNmUJd6_0),.clk(gclk));
	jdff dff_A_uRkmLDwz7_2(.dout(w_G4090_2[2]),.din(w_dff_A_uRkmLDwz7_2),.clk(gclk));
	jdff dff_B_BGVVzNqh7_2(.din(G103),.dout(w_dff_B_BGVVzNqh7_2),.clk(gclk));
	jdff dff_B_VwyDH8wE1_1(.din(n1317),.dout(w_dff_B_VwyDH8wE1_1),.clk(gclk));
	jdff dff_B_XOjiSMhh1_0(.din(n1333),.dout(w_dff_B_XOjiSMhh1_0),.clk(gclk));
	jdff dff_B_Z8tTqNO08_0(.din(w_dff_B_XOjiSMhh1_0),.dout(w_dff_B_Z8tTqNO08_0),.clk(gclk));
	jdff dff_B_EPscGlBm4_0(.din(w_dff_B_Z8tTqNO08_0),.dout(w_dff_B_EPscGlBm4_0),.clk(gclk));
	jdff dff_B_ZSuExcoD5_0(.din(w_dff_B_EPscGlBm4_0),.dout(w_dff_B_ZSuExcoD5_0),.clk(gclk));
	jdff dff_B_Z9FwUdeg9_0(.din(w_dff_B_ZSuExcoD5_0),.dout(w_dff_B_Z9FwUdeg9_0),.clk(gclk));
	jdff dff_B_rxgoapfK8_0(.din(w_dff_B_Z9FwUdeg9_0),.dout(w_dff_B_rxgoapfK8_0),.clk(gclk));
	jdff dff_B_cg5CIlMC6_0(.din(w_dff_B_rxgoapfK8_0),.dout(w_dff_B_cg5CIlMC6_0),.clk(gclk));
	jdff dff_B_9CDAg0i09_0(.din(w_dff_B_cg5CIlMC6_0),.dout(w_dff_B_9CDAg0i09_0),.clk(gclk));
	jdff dff_B_ko5wrpcG1_0(.din(w_dff_B_9CDAg0i09_0),.dout(w_dff_B_ko5wrpcG1_0),.clk(gclk));
	jdff dff_B_eL2xxCXb3_0(.din(w_dff_B_ko5wrpcG1_0),.dout(w_dff_B_eL2xxCXb3_0),.clk(gclk));
	jdff dff_B_TdetwKw54_0(.din(w_dff_B_eL2xxCXb3_0),.dout(w_dff_B_TdetwKw54_0),.clk(gclk));
	jdff dff_B_it33mLoO2_0(.din(w_dff_B_TdetwKw54_0),.dout(w_dff_B_it33mLoO2_0),.clk(gclk));
	jdff dff_B_CgJk59Z23_0(.din(w_dff_B_it33mLoO2_0),.dout(w_dff_B_CgJk59Z23_0),.clk(gclk));
	jdff dff_B_DiUfPGgd6_0(.din(w_dff_B_CgJk59Z23_0),.dout(w_dff_B_DiUfPGgd6_0),.clk(gclk));
	jdff dff_B_zJalZ0Rc6_0(.din(w_dff_B_DiUfPGgd6_0),.dout(w_dff_B_zJalZ0Rc6_0),.clk(gclk));
	jdff dff_B_2Qzm5fIQ3_0(.din(w_dff_B_zJalZ0Rc6_0),.dout(w_dff_B_2Qzm5fIQ3_0),.clk(gclk));
	jdff dff_B_SZYu7Suh5_0(.din(w_dff_B_2Qzm5fIQ3_0),.dout(w_dff_B_SZYu7Suh5_0),.clk(gclk));
	jdff dff_B_P9BQJHRS3_0(.din(w_dff_B_SZYu7Suh5_0),.dout(w_dff_B_P9BQJHRS3_0),.clk(gclk));
	jdff dff_B_ZMLXcoSU6_0(.din(w_dff_B_P9BQJHRS3_0),.dout(w_dff_B_ZMLXcoSU6_0),.clk(gclk));
	jdff dff_B_t85foF892_2(.din(G40),.dout(w_dff_B_t85foF892_2),.clk(gclk));
	jdff dff_B_SitaWkjy3_1(.din(n1326),.dout(w_dff_B_SitaWkjy3_1),.clk(gclk));
	jdff dff_B_hOIKizSm7_1(.din(w_dff_B_SitaWkjy3_1),.dout(w_dff_B_hOIKizSm7_1),.clk(gclk));
	jdff dff_B_ZdDAzTRd3_1(.din(w_dff_B_hOIKizSm7_1),.dout(w_dff_B_ZdDAzTRd3_1),.clk(gclk));
	jdff dff_A_by2ZWpO37_0(.dout(w_n852_4[0]),.din(w_dff_A_by2ZWpO37_0),.clk(gclk));
	jdff dff_A_ie0b4jAk4_0(.dout(w_dff_A_by2ZWpO37_0),.din(w_dff_A_ie0b4jAk4_0),.clk(gclk));
	jdff dff_A_esGKByTC7_0(.dout(w_dff_A_ie0b4jAk4_0),.din(w_dff_A_esGKByTC7_0),.clk(gclk));
	jdff dff_A_hZs1WtX98_0(.dout(w_dff_A_esGKByTC7_0),.din(w_dff_A_hZs1WtX98_0),.clk(gclk));
	jdff dff_A_K1Rw60c30_0(.dout(w_dff_A_hZs1WtX98_0),.din(w_dff_A_K1Rw60c30_0),.clk(gclk));
	jdff dff_A_VF7lNyY25_0(.dout(w_dff_A_K1Rw60c30_0),.din(w_dff_A_VF7lNyY25_0),.clk(gclk));
	jdff dff_A_ILcIecHr3_0(.dout(w_dff_A_VF7lNyY25_0),.din(w_dff_A_ILcIecHr3_0),.clk(gclk));
	jdff dff_A_mQIQYFXF7_0(.dout(w_dff_A_ILcIecHr3_0),.din(w_dff_A_mQIQYFXF7_0),.clk(gclk));
	jdff dff_A_ahNcR6lG6_0(.dout(w_dff_A_mQIQYFXF7_0),.din(w_dff_A_ahNcR6lG6_0),.clk(gclk));
	jdff dff_A_2ayUgYl83_0(.dout(w_dff_A_ahNcR6lG6_0),.din(w_dff_A_2ayUgYl83_0),.clk(gclk));
	jdff dff_A_8yTjE47g1_0(.dout(w_dff_A_2ayUgYl83_0),.din(w_dff_A_8yTjE47g1_0),.clk(gclk));
	jdff dff_A_a3TyolLG8_0(.dout(w_dff_A_8yTjE47g1_0),.din(w_dff_A_a3TyolLG8_0),.clk(gclk));
	jdff dff_A_c4RUVjH83_0(.dout(w_dff_A_a3TyolLG8_0),.din(w_dff_A_c4RUVjH83_0),.clk(gclk));
	jdff dff_A_TaHuFmQ14_0(.dout(w_dff_A_c4RUVjH83_0),.din(w_dff_A_TaHuFmQ14_0),.clk(gclk));
	jdff dff_A_T8Pmqg4G4_0(.dout(w_dff_A_TaHuFmQ14_0),.din(w_dff_A_T8Pmqg4G4_0),.clk(gclk));
	jdff dff_A_KvoQN0Ve8_0(.dout(w_dff_A_T8Pmqg4G4_0),.din(w_dff_A_KvoQN0Ve8_0),.clk(gclk));
	jdff dff_A_LGZ0akvm4_0(.dout(w_dff_A_KvoQN0Ve8_0),.din(w_dff_A_LGZ0akvm4_0),.clk(gclk));
	jdff dff_A_fxyaCb5N2_0(.dout(w_dff_A_LGZ0akvm4_0),.din(w_dff_A_fxyaCb5N2_0),.clk(gclk));
	jdff dff_A_XbjMvyRI0_2(.dout(w_n852_4[2]),.din(w_dff_A_XbjMvyRI0_2),.clk(gclk));
	jdff dff_A_T2bA6jRM9_2(.dout(w_dff_A_XbjMvyRI0_2),.din(w_dff_A_T2bA6jRM9_2),.clk(gclk));
	jdff dff_A_AKOBf5E62_2(.dout(w_dff_A_T2bA6jRM9_2),.din(w_dff_A_AKOBf5E62_2),.clk(gclk));
	jdff dff_A_y8fZEZoG9_2(.dout(w_dff_A_AKOBf5E62_2),.din(w_dff_A_y8fZEZoG9_2),.clk(gclk));
	jdff dff_A_8l70AWw09_2(.dout(w_dff_A_y8fZEZoG9_2),.din(w_dff_A_8l70AWw09_2),.clk(gclk));
	jdff dff_A_8yeNDHZb9_2(.dout(w_dff_A_8l70AWw09_2),.din(w_dff_A_8yeNDHZb9_2),.clk(gclk));
	jdff dff_A_pTbMdTeW4_2(.dout(w_dff_A_8yeNDHZb9_2),.din(w_dff_A_pTbMdTeW4_2),.clk(gclk));
	jdff dff_A_DTl5ZaCh6_2(.dout(w_dff_A_pTbMdTeW4_2),.din(w_dff_A_DTl5ZaCh6_2),.clk(gclk));
	jdff dff_A_niERBPN88_2(.dout(w_dff_A_DTl5ZaCh6_2),.din(w_dff_A_niERBPN88_2),.clk(gclk));
	jdff dff_A_sHfpWgE41_2(.dout(w_dff_A_niERBPN88_2),.din(w_dff_A_sHfpWgE41_2),.clk(gclk));
	jdff dff_A_U0dCrpGY6_2(.dout(w_dff_A_sHfpWgE41_2),.din(w_dff_A_U0dCrpGY6_2),.clk(gclk));
	jdff dff_A_y4Ho3ifi1_2(.dout(w_dff_A_U0dCrpGY6_2),.din(w_dff_A_y4Ho3ifi1_2),.clk(gclk));
	jdff dff_A_olHhnR640_2(.dout(w_dff_A_y4Ho3ifi1_2),.din(w_dff_A_olHhnR640_2),.clk(gclk));
	jdff dff_A_wq7z9bw63_2(.dout(w_dff_A_olHhnR640_2),.din(w_dff_A_wq7z9bw63_2),.clk(gclk));
	jdff dff_A_jYAnm2Ef5_2(.dout(w_dff_A_wq7z9bw63_2),.din(w_dff_A_jYAnm2Ef5_2),.clk(gclk));
	jdff dff_A_idF6996p9_2(.dout(w_dff_A_jYAnm2Ef5_2),.din(w_dff_A_idF6996p9_2),.clk(gclk));
	jdff dff_A_TN4Wuusu5_2(.dout(w_dff_A_idF6996p9_2),.din(w_dff_A_TN4Wuusu5_2),.clk(gclk));
	jdff dff_A_uvaYWoK85_2(.dout(w_dff_A_TN4Wuusu5_2),.din(w_dff_A_uvaYWoK85_2),.clk(gclk));
	jdff dff_A_HFOfGJ697_2(.dout(w_dff_A_uvaYWoK85_2),.din(w_dff_A_HFOfGJ697_2),.clk(gclk));
	jdff dff_A_PbS1Dyty5_0(.dout(w_G4089_4[0]),.din(w_dff_A_PbS1Dyty5_0),.clk(gclk));
	jdff dff_A_qJUwRZle8_0(.dout(w_dff_A_PbS1Dyty5_0),.din(w_dff_A_qJUwRZle8_0),.clk(gclk));
	jdff dff_A_RXQT9YT18_0(.dout(w_dff_A_qJUwRZle8_0),.din(w_dff_A_RXQT9YT18_0),.clk(gclk));
	jdff dff_A_OtAELsg52_0(.dout(w_dff_A_RXQT9YT18_0),.din(w_dff_A_OtAELsg52_0),.clk(gclk));
	jdff dff_A_asBKpU700_0(.dout(w_dff_A_OtAELsg52_0),.din(w_dff_A_asBKpU700_0),.clk(gclk));
	jdff dff_A_7imHS2CW0_0(.dout(w_dff_A_asBKpU700_0),.din(w_dff_A_7imHS2CW0_0),.clk(gclk));
	jdff dff_A_z4Qm6UW55_0(.dout(w_dff_A_7imHS2CW0_0),.din(w_dff_A_z4Qm6UW55_0),.clk(gclk));
	jdff dff_A_Eg5EPzsk6_0(.dout(w_dff_A_z4Qm6UW55_0),.din(w_dff_A_Eg5EPzsk6_0),.clk(gclk));
	jdff dff_A_KIvcsf1l0_0(.dout(w_dff_A_Eg5EPzsk6_0),.din(w_dff_A_KIvcsf1l0_0),.clk(gclk));
	jdff dff_A_3hLwwdsr3_0(.dout(w_dff_A_KIvcsf1l0_0),.din(w_dff_A_3hLwwdsr3_0),.clk(gclk));
	jdff dff_A_rkMHbOso7_0(.dout(w_dff_A_3hLwwdsr3_0),.din(w_dff_A_rkMHbOso7_0),.clk(gclk));
	jdff dff_A_7jqmFCAY6_0(.dout(w_dff_A_rkMHbOso7_0),.din(w_dff_A_7jqmFCAY6_0),.clk(gclk));
	jdff dff_A_GIN3W9H24_0(.dout(w_dff_A_7jqmFCAY6_0),.din(w_dff_A_GIN3W9H24_0),.clk(gclk));
	jdff dff_A_QumNV0cR9_0(.dout(w_dff_A_GIN3W9H24_0),.din(w_dff_A_QumNV0cR9_0),.clk(gclk));
	jdff dff_A_2XITXUSG1_0(.dout(w_dff_A_QumNV0cR9_0),.din(w_dff_A_2XITXUSG1_0),.clk(gclk));
	jdff dff_A_D1Nz5B0M1_0(.dout(w_dff_A_2XITXUSG1_0),.din(w_dff_A_D1Nz5B0M1_0),.clk(gclk));
	jdff dff_A_KR9zwP2a9_0(.dout(w_dff_A_D1Nz5B0M1_0),.din(w_dff_A_KR9zwP2a9_0),.clk(gclk));
	jdff dff_A_ofsxSK8w5_2(.dout(w_G4089_4[2]),.din(w_dff_A_ofsxSK8w5_2),.clk(gclk));
	jdff dff_A_2eh89Xiw1_2(.dout(w_dff_A_ofsxSK8w5_2),.din(w_dff_A_2eh89Xiw1_2),.clk(gclk));
	jdff dff_A_FxuohrWp6_2(.dout(w_dff_A_2eh89Xiw1_2),.din(w_dff_A_FxuohrWp6_2),.clk(gclk));
	jdff dff_A_iCoN45B83_2(.dout(w_dff_A_FxuohrWp6_2),.din(w_dff_A_iCoN45B83_2),.clk(gclk));
	jdff dff_A_LTHvzbjP6_2(.dout(w_dff_A_iCoN45B83_2),.din(w_dff_A_LTHvzbjP6_2),.clk(gclk));
	jdff dff_A_6CLnFoqv8_2(.dout(w_dff_A_LTHvzbjP6_2),.din(w_dff_A_6CLnFoqv8_2),.clk(gclk));
	jdff dff_A_i9sVupR50_2(.dout(w_dff_A_6CLnFoqv8_2),.din(w_dff_A_i9sVupR50_2),.clk(gclk));
	jdff dff_A_klecAp9m1_2(.dout(w_dff_A_i9sVupR50_2),.din(w_dff_A_klecAp9m1_2),.clk(gclk));
	jdff dff_A_iUvccvH48_2(.dout(w_dff_A_klecAp9m1_2),.din(w_dff_A_iUvccvH48_2),.clk(gclk));
	jdff dff_A_3adhuu0b5_2(.dout(w_dff_A_iUvccvH48_2),.din(w_dff_A_3adhuu0b5_2),.clk(gclk));
	jdff dff_A_i3ApvijZ2_2(.dout(w_dff_A_3adhuu0b5_2),.din(w_dff_A_i3ApvijZ2_2),.clk(gclk));
	jdff dff_A_nU4ZQWXR0_2(.dout(w_dff_A_i3ApvijZ2_2),.din(w_dff_A_nU4ZQWXR0_2),.clk(gclk));
	jdff dff_A_p3UwHcrX3_2(.dout(w_dff_A_nU4ZQWXR0_2),.din(w_dff_A_p3UwHcrX3_2),.clk(gclk));
	jdff dff_A_OkLzUhR09_2(.dout(w_dff_A_p3UwHcrX3_2),.din(w_dff_A_OkLzUhR09_2),.clk(gclk));
	jdff dff_A_AWvzkvRJ0_2(.dout(w_dff_A_OkLzUhR09_2),.din(w_dff_A_AWvzkvRJ0_2),.clk(gclk));
	jdff dff_A_S61aay9x6_2(.dout(w_dff_A_AWvzkvRJ0_2),.din(w_dff_A_S61aay9x6_2),.clk(gclk));
	jdff dff_A_TttGYNRt5_2(.dout(w_dff_A_S61aay9x6_2),.din(w_dff_A_TttGYNRt5_2),.clk(gclk));
	jdff dff_A_lkiDT9Ip1_2(.dout(w_dff_A_TttGYNRt5_2),.din(w_dff_A_lkiDT9Ip1_2),.clk(gclk));
	jdff dff_A_QVJf2g3j8_2(.dout(w_dff_A_lkiDT9Ip1_2),.din(w_dff_A_QVJf2g3j8_2),.clk(gclk));
	jdff dff_A_u9j9nshs9_2(.dout(w_dff_A_QVJf2g3j8_2),.din(w_dff_A_u9j9nshs9_2),.clk(gclk));
	jdff dff_B_mshRwsy15_0(.din(n1341),.dout(w_dff_B_mshRwsy15_0),.clk(gclk));
	jdff dff_B_5OUtjts12_0(.din(w_dff_B_mshRwsy15_0),.dout(w_dff_B_5OUtjts12_0),.clk(gclk));
	jdff dff_B_VYbzqxtc2_0(.din(w_dff_B_5OUtjts12_0),.dout(w_dff_B_VYbzqxtc2_0),.clk(gclk));
	jdff dff_B_IU7kvnLJ1_0(.din(w_dff_B_VYbzqxtc2_0),.dout(w_dff_B_IU7kvnLJ1_0),.clk(gclk));
	jdff dff_B_YgT2FB157_0(.din(w_dff_B_IU7kvnLJ1_0),.dout(w_dff_B_YgT2FB157_0),.clk(gclk));
	jdff dff_B_3K9M6PQ34_0(.din(w_dff_B_YgT2FB157_0),.dout(w_dff_B_3K9M6PQ34_0),.clk(gclk));
	jdff dff_B_B6TgXyfQ6_0(.din(w_dff_B_3K9M6PQ34_0),.dout(w_dff_B_B6TgXyfQ6_0),.clk(gclk));
	jdff dff_B_HaxRkJZa8_0(.din(w_dff_B_B6TgXyfQ6_0),.dout(w_dff_B_HaxRkJZa8_0),.clk(gclk));
	jdff dff_B_w7AOvR1R4_0(.din(w_dff_B_HaxRkJZa8_0),.dout(w_dff_B_w7AOvR1R4_0),.clk(gclk));
	jdff dff_B_OF7SeKIn9_0(.din(w_dff_B_w7AOvR1R4_0),.dout(w_dff_B_OF7SeKIn9_0),.clk(gclk));
	jdff dff_B_MCjGfvfv8_0(.din(w_dff_B_OF7SeKIn9_0),.dout(w_dff_B_MCjGfvfv8_0),.clk(gclk));
	jdff dff_B_3nJ1XFp51_0(.din(w_dff_B_MCjGfvfv8_0),.dout(w_dff_B_3nJ1XFp51_0),.clk(gclk));
	jdff dff_B_bjWvK6MY7_0(.din(w_dff_B_3nJ1XFp51_0),.dout(w_dff_B_bjWvK6MY7_0),.clk(gclk));
	jdff dff_B_hfGImiBG3_0(.din(w_dff_B_bjWvK6MY7_0),.dout(w_dff_B_hfGImiBG3_0),.clk(gclk));
	jdff dff_B_3jmRfZ6H2_0(.din(w_dff_B_hfGImiBG3_0),.dout(w_dff_B_3jmRfZ6H2_0),.clk(gclk));
	jdff dff_B_oSGRjATN5_0(.din(w_dff_B_3jmRfZ6H2_0),.dout(w_dff_B_oSGRjATN5_0),.clk(gclk));
	jdff dff_B_Ds0udzs05_0(.din(w_dff_B_oSGRjATN5_0),.dout(w_dff_B_Ds0udzs05_0),.clk(gclk));
	jdff dff_B_eVq55WOs0_0(.din(w_dff_B_Ds0udzs05_0),.dout(w_dff_B_eVq55WOs0_0),.clk(gclk));
	jdff dff_B_ZwbUsRCP6_0(.din(n1340),.dout(w_dff_B_ZwbUsRCP6_0),.clk(gclk));
	jdff dff_B_G4jUsiup6_1(.din(n1335),.dout(w_dff_B_G4jUsiup6_1),.clk(gclk));
	jdff dff_B_4t4hdD2x4_1(.din(w_dff_B_G4jUsiup6_1),.dout(w_dff_B_4t4hdD2x4_1),.clk(gclk));
	jdff dff_B_iodepxmR8_1(.din(w_dff_B_4t4hdD2x4_1),.dout(w_dff_B_iodepxmR8_1),.clk(gclk));
	jdff dff_A_GSyRofOQ7_0(.dout(w_n999_2[0]),.din(w_dff_A_GSyRofOQ7_0),.clk(gclk));
	jdff dff_A_hgh9N07M2_0(.dout(w_dff_A_GSyRofOQ7_0),.din(w_dff_A_hgh9N07M2_0),.clk(gclk));
	jdff dff_A_u9sRUKwF3_0(.dout(w_dff_A_hgh9N07M2_0),.din(w_dff_A_u9sRUKwF3_0),.clk(gclk));
	jdff dff_A_Tyr7VT9b3_0(.dout(w_dff_A_u9sRUKwF3_0),.din(w_dff_A_Tyr7VT9b3_0),.clk(gclk));
	jdff dff_A_Q1yahVas4_0(.dout(w_dff_A_Tyr7VT9b3_0),.din(w_dff_A_Q1yahVas4_0),.clk(gclk));
	jdff dff_A_ofsuAHg40_0(.dout(w_dff_A_Q1yahVas4_0),.din(w_dff_A_ofsuAHg40_0),.clk(gclk));
	jdff dff_A_BCdCY5Bq5_1(.dout(w_n999_2[1]),.din(w_dff_A_BCdCY5Bq5_1),.clk(gclk));
	jdff dff_A_ECxU1y2h3_0(.dout(w_G1689_3[0]),.din(w_dff_A_ECxU1y2h3_0),.clk(gclk));
	jdff dff_A_4CVT1Hot5_0(.dout(w_dff_A_ECxU1y2h3_0),.din(w_dff_A_4CVT1Hot5_0),.clk(gclk));
	jdff dff_A_ctnCsLVJ4_0(.dout(w_dff_A_4CVT1Hot5_0),.din(w_dff_A_ctnCsLVJ4_0),.clk(gclk));
	jdff dff_A_wZh9lAPx0_0(.dout(w_dff_A_ctnCsLVJ4_0),.din(w_dff_A_wZh9lAPx0_0),.clk(gclk));
	jdff dff_A_8mUEnxPQ0_1(.dout(w_G1689_3[1]),.din(w_dff_A_8mUEnxPQ0_1),.clk(gclk));
	jdff dff_A_logOGiod7_1(.dout(w_dff_A_8mUEnxPQ0_1),.din(w_dff_A_logOGiod7_1),.clk(gclk));
	jdff dff_A_ifnZ00NC1_0(.dout(w_G137_6[0]),.din(w_dff_A_ifnZ00NC1_0),.clk(gclk));
	jdff dff_A_D1Ua89gJ3_0(.dout(w_dff_A_ifnZ00NC1_0),.din(w_dff_A_D1Ua89gJ3_0),.clk(gclk));
	jdff dff_A_k64mAtH56_0(.dout(w_dff_A_D1Ua89gJ3_0),.din(w_dff_A_k64mAtH56_0),.clk(gclk));
	jdff dff_A_SLZgQgE55_0(.dout(w_dff_A_k64mAtH56_0),.din(w_dff_A_SLZgQgE55_0),.clk(gclk));
	jdff dff_A_BwyTTUWD1_0(.dout(w_dff_A_SLZgQgE55_0),.din(w_dff_A_BwyTTUWD1_0),.clk(gclk));
	jdff dff_A_f5mbHDtI7_0(.dout(w_dff_A_BwyTTUWD1_0),.din(w_dff_A_f5mbHDtI7_0),.clk(gclk));
	jdff dff_A_9zUtyW7p6_1(.dout(w_G137_6[1]),.din(w_dff_A_9zUtyW7p6_1),.clk(gclk));
	jdff dff_B_XjaC9nKG1_0(.din(n1350),.dout(w_dff_B_XjaC9nKG1_0),.clk(gclk));
	jdff dff_B_ZEDC7mwH7_0(.din(w_dff_B_XjaC9nKG1_0),.dout(w_dff_B_ZEDC7mwH7_0),.clk(gclk));
	jdff dff_B_EkORrSbH4_0(.din(w_dff_B_ZEDC7mwH7_0),.dout(w_dff_B_EkORrSbH4_0),.clk(gclk));
	jdff dff_B_NvgGy6PA7_0(.din(w_dff_B_EkORrSbH4_0),.dout(w_dff_B_NvgGy6PA7_0),.clk(gclk));
	jdff dff_B_8tzfis8M8_0(.din(w_dff_B_NvgGy6PA7_0),.dout(w_dff_B_8tzfis8M8_0),.clk(gclk));
	jdff dff_B_0PaRI3PM5_0(.din(w_dff_B_8tzfis8M8_0),.dout(w_dff_B_0PaRI3PM5_0),.clk(gclk));
	jdff dff_B_JTsamusx0_0(.din(w_dff_B_0PaRI3PM5_0),.dout(w_dff_B_JTsamusx0_0),.clk(gclk));
	jdff dff_B_HjvntQIJ4_0(.din(w_dff_B_JTsamusx0_0),.dout(w_dff_B_HjvntQIJ4_0),.clk(gclk));
	jdff dff_B_wrYh4IKt1_0(.din(w_dff_B_HjvntQIJ4_0),.dout(w_dff_B_wrYh4IKt1_0),.clk(gclk));
	jdff dff_B_GOTQGqsC4_0(.din(w_dff_B_wrYh4IKt1_0),.dout(w_dff_B_GOTQGqsC4_0),.clk(gclk));
	jdff dff_B_5sRSuzAU3_0(.din(w_dff_B_GOTQGqsC4_0),.dout(w_dff_B_5sRSuzAU3_0),.clk(gclk));
	jdff dff_B_bB6CWHQR7_0(.din(w_dff_B_5sRSuzAU3_0),.dout(w_dff_B_bB6CWHQR7_0),.clk(gclk));
	jdff dff_B_f1w60ZHt1_0(.din(w_dff_B_bB6CWHQR7_0),.dout(w_dff_B_f1w60ZHt1_0),.clk(gclk));
	jdff dff_B_1f3yI4xk6_0(.din(w_dff_B_f1w60ZHt1_0),.dout(w_dff_B_1f3yI4xk6_0),.clk(gclk));
	jdff dff_B_FOvcNYLR7_0(.din(w_dff_B_1f3yI4xk6_0),.dout(w_dff_B_FOvcNYLR7_0),.clk(gclk));
	jdff dff_B_PKY53IIb3_0(.din(w_dff_B_FOvcNYLR7_0),.dout(w_dff_B_PKY53IIb3_0),.clk(gclk));
	jdff dff_B_TCGNstJk9_0(.din(w_dff_B_PKY53IIb3_0),.dout(w_dff_B_TCGNstJk9_0),.clk(gclk));
	jdff dff_B_RiYAOghw7_0(.din(w_dff_B_TCGNstJk9_0),.dout(w_dff_B_RiYAOghw7_0),.clk(gclk));
	jdff dff_B_MSnu5F2k2_0(.din(w_dff_B_RiYAOghw7_0),.dout(w_dff_B_MSnu5F2k2_0),.clk(gclk));
	jdff dff_B_A9RfTUUr4_0(.din(n1349),.dout(w_dff_B_A9RfTUUr4_0),.clk(gclk));
	jdff dff_B_pXPjkzqj2_1(.din(n1344),.dout(w_dff_B_pXPjkzqj2_1),.clk(gclk));
	jdff dff_B_rVKnJ34T9_1(.din(n1355),.dout(w_dff_B_rVKnJ34T9_1),.clk(gclk));
	jdff dff_B_Hkk4bdr51_1(.din(w_dff_B_rVKnJ34T9_1),.dout(w_dff_B_Hkk4bdr51_1),.clk(gclk));
	jdff dff_B_5SSN6Lbr9_1(.din(w_dff_B_Hkk4bdr51_1),.dout(w_dff_B_5SSN6Lbr9_1),.clk(gclk));
	jdff dff_B_B44k5oz26_1(.din(w_dff_B_5SSN6Lbr9_1),.dout(w_dff_B_B44k5oz26_1),.clk(gclk));
	jdff dff_B_Sl64ll7i0_1(.din(w_dff_B_B44k5oz26_1),.dout(w_dff_B_Sl64ll7i0_1),.clk(gclk));
	jdff dff_B_q7pKPDPL3_1(.din(w_dff_B_Sl64ll7i0_1),.dout(w_dff_B_q7pKPDPL3_1),.clk(gclk));
	jdff dff_B_HiWYwMmy0_1(.din(w_dff_B_q7pKPDPL3_1),.dout(w_dff_B_HiWYwMmy0_1),.clk(gclk));
	jdff dff_B_VptNvT6w3_1(.din(w_dff_B_HiWYwMmy0_1),.dout(w_dff_B_VptNvT6w3_1),.clk(gclk));
	jdff dff_B_O5t6VBUW4_1(.din(w_dff_B_VptNvT6w3_1),.dout(w_dff_B_O5t6VBUW4_1),.clk(gclk));
	jdff dff_B_R1GJTSVh0_1(.din(w_dff_B_O5t6VBUW4_1),.dout(w_dff_B_R1GJTSVh0_1),.clk(gclk));
	jdff dff_B_AeROLd9g8_1(.din(w_dff_B_R1GJTSVh0_1),.dout(w_dff_B_AeROLd9g8_1),.clk(gclk));
	jdff dff_B_OtN8yW254_1(.din(w_dff_B_AeROLd9g8_1),.dout(w_dff_B_OtN8yW254_1),.clk(gclk));
	jdff dff_B_xMoW2Dhx7_1(.din(w_dff_B_OtN8yW254_1),.dout(w_dff_B_xMoW2Dhx7_1),.clk(gclk));
	jdff dff_B_nc1BxIhm3_1(.din(w_dff_B_xMoW2Dhx7_1),.dout(w_dff_B_nc1BxIhm3_1),.clk(gclk));
	jdff dff_B_9OE8mQuF3_1(.din(w_dff_B_nc1BxIhm3_1),.dout(w_dff_B_9OE8mQuF3_1),.clk(gclk));
	jdff dff_B_2fhg3qiy4_1(.din(w_dff_B_9OE8mQuF3_1),.dout(w_dff_B_2fhg3qiy4_1),.clk(gclk));
	jdff dff_B_HvNa44bQ7_1(.din(w_dff_B_2fhg3qiy4_1),.dout(w_dff_B_HvNa44bQ7_1),.clk(gclk));
	jdff dff_B_62WZ5jra6_1(.din(w_dff_B_HvNa44bQ7_1),.dout(w_dff_B_62WZ5jra6_1),.clk(gclk));
	jdff dff_B_KUFA6Oyb8_1(.din(w_dff_B_62WZ5jra6_1),.dout(w_dff_B_KUFA6Oyb8_1),.clk(gclk));
	jdff dff_B_dzStsXEr1_1(.din(n1356),.dout(w_dff_B_dzStsXEr1_1),.clk(gclk));
	jdff dff_A_UJV9MCdP1_0(.dout(w_n993_2[0]),.din(w_dff_A_UJV9MCdP1_0),.clk(gclk));
	jdff dff_A_LZMJYExx1_1(.dout(w_n993_2[1]),.din(w_dff_A_LZMJYExx1_1),.clk(gclk));
	jdff dff_B_CWFOGWVM9_0(.din(n1354),.dout(w_dff_B_CWFOGWVM9_0),.clk(gclk));
	jdff dff_B_wh8zH6Xi6_1(.din(n1364),.dout(w_dff_B_wh8zH6Xi6_1),.clk(gclk));
	jdff dff_B_72Kzoy8E7_1(.din(w_dff_B_wh8zH6Xi6_1),.dout(w_dff_B_72Kzoy8E7_1),.clk(gclk));
	jdff dff_B_Q6iNnIcH9_1(.din(w_dff_B_72Kzoy8E7_1),.dout(w_dff_B_Q6iNnIcH9_1),.clk(gclk));
	jdff dff_B_ksA3Qrcc9_1(.din(w_dff_B_Q6iNnIcH9_1),.dout(w_dff_B_ksA3Qrcc9_1),.clk(gclk));
	jdff dff_B_wevj9OWe1_1(.din(w_dff_B_ksA3Qrcc9_1),.dout(w_dff_B_wevj9OWe1_1),.clk(gclk));
	jdff dff_B_Hyvlp0Q17_1(.din(w_dff_B_wevj9OWe1_1),.dout(w_dff_B_Hyvlp0Q17_1),.clk(gclk));
	jdff dff_B_VO9tCWRW9_1(.din(w_dff_B_Hyvlp0Q17_1),.dout(w_dff_B_VO9tCWRW9_1),.clk(gclk));
	jdff dff_B_6qWfUCn13_1(.din(w_dff_B_VO9tCWRW9_1),.dout(w_dff_B_6qWfUCn13_1),.clk(gclk));
	jdff dff_B_rF5XBp3F5_1(.din(w_dff_B_6qWfUCn13_1),.dout(w_dff_B_rF5XBp3F5_1),.clk(gclk));
	jdff dff_B_q2oX5MxI5_1(.din(w_dff_B_rF5XBp3F5_1),.dout(w_dff_B_q2oX5MxI5_1),.clk(gclk));
	jdff dff_B_Zf2qB9y65_1(.din(w_dff_B_q2oX5MxI5_1),.dout(w_dff_B_Zf2qB9y65_1),.clk(gclk));
	jdff dff_B_opxgwODg5_1(.din(w_dff_B_Zf2qB9y65_1),.dout(w_dff_B_opxgwODg5_1),.clk(gclk));
	jdff dff_B_2Qs9TehO5_1(.din(w_dff_B_opxgwODg5_1),.dout(w_dff_B_2Qs9TehO5_1),.clk(gclk));
	jdff dff_B_mkKF3TOm3_1(.din(w_dff_B_2Qs9TehO5_1),.dout(w_dff_B_mkKF3TOm3_1),.clk(gclk));
	jdff dff_B_CF0ODAgd0_1(.din(w_dff_B_mkKF3TOm3_1),.dout(w_dff_B_CF0ODAgd0_1),.clk(gclk));
	jdff dff_B_ITanyA184_1(.din(w_dff_B_CF0ODAgd0_1),.dout(w_dff_B_ITanyA184_1),.clk(gclk));
	jdff dff_B_TnTWAq0f1_1(.din(w_dff_B_ITanyA184_1),.dout(w_dff_B_TnTWAq0f1_1),.clk(gclk));
	jdff dff_B_avgwYtql8_1(.din(w_dff_B_TnTWAq0f1_1),.dout(w_dff_B_avgwYtql8_1),.clk(gclk));
	jdff dff_B_iOkN3Tgq2_1(.din(w_dff_B_avgwYtql8_1),.dout(w_dff_B_iOkN3Tgq2_1),.clk(gclk));
	jdff dff_B_uDgQeQAK7_1(.din(w_dff_B_iOkN3Tgq2_1),.dout(w_dff_B_uDgQeQAK7_1),.clk(gclk));
	jdff dff_B_7pe10V1S7_1(.din(n1365),.dout(w_dff_B_7pe10V1S7_1),.clk(gclk));
	jdff dff_A_6wDgPfXN7_0(.dout(w_G1689_2[0]),.din(w_dff_A_6wDgPfXN7_0),.clk(gclk));
	jdff dff_A_aNM8e70a3_2(.dout(w_G1689_2[2]),.din(w_dff_A_aNM8e70a3_2),.clk(gclk));
	jdff dff_A_qISB8Hi53_0(.dout(w_n999_1[0]),.din(w_dff_A_qISB8Hi53_0),.clk(gclk));
	jdff dff_A_lDSczqec3_0(.dout(w_dff_A_qISB8Hi53_0),.din(w_dff_A_lDSczqec3_0),.clk(gclk));
	jdff dff_A_50ph0ZCE3_1(.dout(w_n999_1[1]),.din(w_dff_A_50ph0ZCE3_1),.clk(gclk));
	jdff dff_A_WwQXQ3I17_0(.dout(w_n999_0[0]),.din(w_dff_A_WwQXQ3I17_0),.clk(gclk));
	jdff dff_A_eVmXohnV6_0(.dout(w_dff_A_WwQXQ3I17_0),.din(w_dff_A_eVmXohnV6_0),.clk(gclk));
	jdff dff_A_DbZeV6nr6_0(.dout(w_dff_A_eVmXohnV6_0),.din(w_dff_A_DbZeV6nr6_0),.clk(gclk));
	jdff dff_A_1etL4rPz1_0(.dout(w_dff_A_DbZeV6nr6_0),.din(w_dff_A_1etL4rPz1_0),.clk(gclk));
	jdff dff_A_bfifcuy50_0(.dout(w_dff_A_1etL4rPz1_0),.din(w_dff_A_bfifcuy50_0),.clk(gclk));
	jdff dff_A_VdkDATmk3_0(.dout(w_dff_A_bfifcuy50_0),.din(w_dff_A_VdkDATmk3_0),.clk(gclk));
	jdff dff_A_2kyhzeyN1_0(.dout(w_dff_A_VdkDATmk3_0),.din(w_dff_A_2kyhzeyN1_0),.clk(gclk));
	jdff dff_A_gPS5eRIT7_0(.dout(w_dff_A_2kyhzeyN1_0),.din(w_dff_A_gPS5eRIT7_0),.clk(gclk));
	jdff dff_A_SKtBkKNz4_0(.dout(w_dff_A_gPS5eRIT7_0),.din(w_dff_A_SKtBkKNz4_0),.clk(gclk));
	jdff dff_A_YWrBOHVH9_0(.dout(w_dff_A_SKtBkKNz4_0),.din(w_dff_A_YWrBOHVH9_0),.clk(gclk));
	jdff dff_A_icU0pCwP7_0(.dout(w_dff_A_YWrBOHVH9_0),.din(w_dff_A_icU0pCwP7_0),.clk(gclk));
	jdff dff_A_8I1dSzGc2_1(.dout(w_n999_0[1]),.din(w_dff_A_8I1dSzGc2_1),.clk(gclk));
	jdff dff_A_cTZ304fU9_1(.dout(w_dff_A_8I1dSzGc2_1),.din(w_dff_A_cTZ304fU9_1),.clk(gclk));
	jdff dff_A_vvxP8EPU3_1(.dout(w_dff_A_cTZ304fU9_1),.din(w_dff_A_vvxP8EPU3_1),.clk(gclk));
	jdff dff_A_aU4vB9mg4_1(.dout(w_dff_A_vvxP8EPU3_1),.din(w_dff_A_aU4vB9mg4_1),.clk(gclk));
	jdff dff_B_MiQC4BOV2_3(.din(n999),.dout(w_dff_B_MiQC4BOV2_3),.clk(gclk));
	jdff dff_B_j9vnrFtC6_3(.din(w_dff_B_MiQC4BOV2_3),.dout(w_dff_B_j9vnrFtC6_3),.clk(gclk));
	jdff dff_B_CHG1cYSZ7_3(.din(w_dff_B_j9vnrFtC6_3),.dout(w_dff_B_CHG1cYSZ7_3),.clk(gclk));
	jdff dff_B_43syjiHN9_3(.din(w_dff_B_CHG1cYSZ7_3),.dout(w_dff_B_43syjiHN9_3),.clk(gclk));
	jdff dff_B_qScJs4je2_3(.din(w_dff_B_43syjiHN9_3),.dout(w_dff_B_qScJs4je2_3),.clk(gclk));
	jdff dff_B_k72mfSlZ3_3(.din(w_dff_B_qScJs4je2_3),.dout(w_dff_B_k72mfSlZ3_3),.clk(gclk));
	jdff dff_B_GMYqfW2v4_3(.din(w_dff_B_k72mfSlZ3_3),.dout(w_dff_B_GMYqfW2v4_3),.clk(gclk));
	jdff dff_B_oSYOYOBo4_3(.din(w_dff_B_GMYqfW2v4_3),.dout(w_dff_B_oSYOYOBo4_3),.clk(gclk));
	jdff dff_B_p5mSOc3W6_3(.din(w_dff_B_oSYOYOBo4_3),.dout(w_dff_B_p5mSOc3W6_3),.clk(gclk));
	jdff dff_B_1G6woDmf7_0(.din(n1363),.dout(w_dff_B_1G6woDmf7_0),.clk(gclk));
	jdff dff_A_yx0qjRcw3_0(.dout(w_G137_5[0]),.din(w_dff_A_yx0qjRcw3_0),.clk(gclk));
	jdff dff_B_V96hvkE21_0(.din(n1377),.dout(w_dff_B_V96hvkE21_0),.clk(gclk));
	jdff dff_B_0ebIHGfR9_0(.din(w_dff_B_V96hvkE21_0),.dout(w_dff_B_0ebIHGfR9_0),.clk(gclk));
	jdff dff_B_JrInJpB18_0(.din(w_dff_B_0ebIHGfR9_0),.dout(w_dff_B_JrInJpB18_0),.clk(gclk));
	jdff dff_B_tJhIb1Y94_0(.din(w_dff_B_JrInJpB18_0),.dout(w_dff_B_tJhIb1Y94_0),.clk(gclk));
	jdff dff_B_iZd4IPhy2_0(.din(w_dff_B_tJhIb1Y94_0),.dout(w_dff_B_iZd4IPhy2_0),.clk(gclk));
	jdff dff_B_C8WdSPPp4_0(.din(w_dff_B_iZd4IPhy2_0),.dout(w_dff_B_C8WdSPPp4_0),.clk(gclk));
	jdff dff_B_2x7Nb5SJ0_0(.din(w_dff_B_C8WdSPPp4_0),.dout(w_dff_B_2x7Nb5SJ0_0),.clk(gclk));
	jdff dff_B_uxahMi3I1_0(.din(w_dff_B_2x7Nb5SJ0_0),.dout(w_dff_B_uxahMi3I1_0),.clk(gclk));
	jdff dff_B_MOWosIV59_0(.din(w_dff_B_uxahMi3I1_0),.dout(w_dff_B_MOWosIV59_0),.clk(gclk));
	jdff dff_B_RRjpjFhs7_0(.din(w_dff_B_MOWosIV59_0),.dout(w_dff_B_RRjpjFhs7_0),.clk(gclk));
	jdff dff_B_4yVWTyJK9_0(.din(w_dff_B_RRjpjFhs7_0),.dout(w_dff_B_4yVWTyJK9_0),.clk(gclk));
	jdff dff_B_EWZchb1d4_0(.din(w_dff_B_4yVWTyJK9_0),.dout(w_dff_B_EWZchb1d4_0),.clk(gclk));
	jdff dff_B_XQUCCKxY1_0(.din(w_dff_B_EWZchb1d4_0),.dout(w_dff_B_XQUCCKxY1_0),.clk(gclk));
	jdff dff_B_qhLkxiM24_0(.din(w_dff_B_XQUCCKxY1_0),.dout(w_dff_B_qhLkxiM24_0),.clk(gclk));
	jdff dff_B_Peuvko154_0(.din(w_dff_B_qhLkxiM24_0),.dout(w_dff_B_Peuvko154_0),.clk(gclk));
	jdff dff_B_2IsVHzDB9_0(.din(w_dff_B_Peuvko154_0),.dout(w_dff_B_2IsVHzDB9_0),.clk(gclk));
	jdff dff_B_v5HfP5tI9_0(.din(w_dff_B_2IsVHzDB9_0),.dout(w_dff_B_v5HfP5tI9_0),.clk(gclk));
	jdff dff_B_hE9dgaei3_0(.din(w_dff_B_v5HfP5tI9_0),.dout(w_dff_B_hE9dgaei3_0),.clk(gclk));
	jdff dff_B_uQVjHuL17_0(.din(n1376),.dout(w_dff_B_uQVjHuL17_0),.clk(gclk));
	jdff dff_B_YqnsoghZ2_2(.din(G173),.dout(w_dff_B_YqnsoghZ2_2),.clk(gclk));
	jdff dff_B_L9QBeQMZ4_2(.din(G203),.dout(w_dff_B_L9QBeQMZ4_2),.clk(gclk));
	jdff dff_B_nk58Ujfl0_2(.din(w_dff_B_L9QBeQMZ4_2),.dout(w_dff_B_nk58Ujfl0_2),.clk(gclk));
	jdff dff_B_9dwlTRPK6_1(.din(n1371),.dout(w_dff_B_9dwlTRPK6_1),.clk(gclk));
	jdff dff_B_PT7K2flI5_1(.din(w_dff_B_9dwlTRPK6_1),.dout(w_dff_B_PT7K2flI5_1),.clk(gclk));
	jdff dff_B_loIilNij4_1(.din(w_dff_B_PT7K2flI5_1),.dout(w_dff_B_loIilNij4_1),.clk(gclk));
	jdff dff_B_rjIiuDHl2_1(.din(n1254),.dout(w_dff_B_rjIiuDHl2_1),.clk(gclk));
	jdff dff_B_7TDxlIQa1_1(.din(w_dff_B_rjIiuDHl2_1),.dout(w_dff_B_7TDxlIQa1_1),.clk(gclk));
	jdff dff_B_5ihw5G2E1_1(.din(w_dff_B_7TDxlIQa1_1),.dout(w_dff_B_5ihw5G2E1_1),.clk(gclk));
	jdff dff_B_wviYuKru8_1(.din(w_dff_B_5ihw5G2E1_1),.dout(w_dff_B_wviYuKru8_1),.clk(gclk));
	jdff dff_B_zbm6UKsS6_1(.din(w_dff_B_wviYuKru8_1),.dout(w_dff_B_zbm6UKsS6_1),.clk(gclk));
	jdff dff_B_K3n1nNSV3_1(.din(w_dff_B_zbm6UKsS6_1),.dout(w_dff_B_K3n1nNSV3_1),.clk(gclk));
	jdff dff_B_ZcR4iINm1_1(.din(w_dff_B_K3n1nNSV3_1),.dout(w_dff_B_ZcR4iINm1_1),.clk(gclk));
	jdff dff_B_gMj0zf4J9_1(.din(w_dff_B_ZcR4iINm1_1),.dout(w_dff_B_gMj0zf4J9_1),.clk(gclk));
	jdff dff_B_zWezU6xw5_1(.din(w_dff_B_gMj0zf4J9_1),.dout(w_dff_B_zWezU6xw5_1),.clk(gclk));
	jdff dff_B_gWEPWpSj1_1(.din(w_dff_B_zWezU6xw5_1),.dout(w_dff_B_gWEPWpSj1_1),.clk(gclk));
	jdff dff_B_87kswRpq0_1(.din(w_dff_B_gWEPWpSj1_1),.dout(w_dff_B_87kswRpq0_1),.clk(gclk));
	jdff dff_B_Nemvtexz4_1(.din(w_dff_B_87kswRpq0_1),.dout(w_dff_B_Nemvtexz4_1),.clk(gclk));
	jdff dff_B_WgBFhtdP5_1(.din(w_dff_B_Nemvtexz4_1),.dout(w_dff_B_WgBFhtdP5_1),.clk(gclk));
	jdff dff_B_cZwe1DK44_0(.din(n1257),.dout(w_dff_B_cZwe1DK44_0),.clk(gclk));
	jdff dff_B_o9C2OPcf2_0(.din(w_dff_B_cZwe1DK44_0),.dout(w_dff_B_o9C2OPcf2_0),.clk(gclk));
	jdff dff_B_wLPm1KOO0_0(.din(w_dff_B_o9C2OPcf2_0),.dout(w_dff_B_wLPm1KOO0_0),.clk(gclk));
	jdff dff_B_nDHwnwGW7_0(.din(w_dff_B_wLPm1KOO0_0),.dout(w_dff_B_nDHwnwGW7_0),.clk(gclk));
	jdff dff_B_EYSEgImC0_0(.din(w_dff_B_nDHwnwGW7_0),.dout(w_dff_B_EYSEgImC0_0),.clk(gclk));
	jdff dff_B_bAtU5uxE1_0(.din(w_dff_B_EYSEgImC0_0),.dout(w_dff_B_bAtU5uxE1_0),.clk(gclk));
	jdff dff_B_w91Uzqrj3_0(.din(w_dff_B_bAtU5uxE1_0),.dout(w_dff_B_w91Uzqrj3_0),.clk(gclk));
	jdff dff_B_GLBNoV7e9_0(.din(w_dff_B_w91Uzqrj3_0),.dout(w_dff_B_GLBNoV7e9_0),.clk(gclk));
	jdff dff_B_hcrYth2O5_0(.din(w_dff_B_GLBNoV7e9_0),.dout(w_dff_B_hcrYth2O5_0),.clk(gclk));
	jdff dff_B_0aVBOMGB7_1(.din(n500),.dout(w_dff_B_0aVBOMGB7_1),.clk(gclk));
	jdff dff_B_NJkMpDqu5_1(.din(n495),.dout(w_dff_B_NJkMpDqu5_1),.clk(gclk));
	jdff dff_B_a8do0Dqr7_1(.din(G113),.dout(w_dff_B_a8do0Dqr7_1),.clk(gclk));
	jdff dff_B_Z0yc7H8z2_1(.din(w_dff_B_a8do0Dqr7_1),.dout(w_dff_B_Z0yc7H8z2_1),.clk(gclk));
	jdff dff_A_drOFPCxq5_0(.dout(w_n1007_2[0]),.din(w_dff_A_drOFPCxq5_0),.clk(gclk));
	jdff dff_A_8rLOe6ph0_0(.dout(w_dff_A_drOFPCxq5_0),.din(w_dff_A_8rLOe6ph0_0),.clk(gclk));
	jdff dff_A_2058o5338_0(.dout(w_dff_A_8rLOe6ph0_0),.din(w_dff_A_2058o5338_0),.clk(gclk));
	jdff dff_A_tWvOCbwQ7_0(.dout(w_dff_A_2058o5338_0),.din(w_dff_A_tWvOCbwQ7_0),.clk(gclk));
	jdff dff_A_hJmoriM15_0(.dout(w_dff_A_tWvOCbwQ7_0),.din(w_dff_A_hJmoriM15_0),.clk(gclk));
	jdff dff_A_aQU1CCTB6_0(.dout(w_dff_A_hJmoriM15_0),.din(w_dff_A_aQU1CCTB6_0),.clk(gclk));
	jdff dff_A_VvUbhN3i4_1(.dout(w_n1007_2[1]),.din(w_dff_A_VvUbhN3i4_1),.clk(gclk));
	jdff dff_B_0cT48kfH1_1(.din(n1216),.dout(w_dff_B_0cT48kfH1_1),.clk(gclk));
	jdff dff_B_YqWTLaJc9_1(.din(w_dff_B_0cT48kfH1_1),.dout(w_dff_B_YqWTLaJc9_1),.clk(gclk));
	jdff dff_B_2wtltuUq8_1(.din(w_dff_B_YqWTLaJc9_1),.dout(w_dff_B_2wtltuUq8_1),.clk(gclk));
	jdff dff_B_EiUttOfP5_1(.din(w_dff_B_2wtltuUq8_1),.dout(w_dff_B_EiUttOfP5_1),.clk(gclk));
	jdff dff_B_mzEKJfeg8_1(.din(w_dff_B_EiUttOfP5_1),.dout(w_dff_B_mzEKJfeg8_1),.clk(gclk));
	jdff dff_B_qfssFEbD9_1(.din(w_dff_B_mzEKJfeg8_1),.dout(w_dff_B_qfssFEbD9_1),.clk(gclk));
	jdff dff_B_crIQj7qM0_1(.din(w_dff_B_qfssFEbD9_1),.dout(w_dff_B_crIQj7qM0_1),.clk(gclk));
	jdff dff_B_o6X1Biji3_1(.din(w_dff_B_crIQj7qM0_1),.dout(w_dff_B_o6X1Biji3_1),.clk(gclk));
	jdff dff_B_plA96Sp41_1(.din(w_dff_B_o6X1Biji3_1),.dout(w_dff_B_plA96Sp41_1),.clk(gclk));
	jdff dff_B_wYcNF72E0_1(.din(w_dff_B_plA96Sp41_1),.dout(w_dff_B_wYcNF72E0_1),.clk(gclk));
	jdff dff_B_AJAIRTUo0_1(.din(w_dff_B_wYcNF72E0_1),.dout(w_dff_B_AJAIRTUo0_1),.clk(gclk));
	jdff dff_B_Yz38cpht3_0(.din(n1219),.dout(w_dff_B_Yz38cpht3_0),.clk(gclk));
	jdff dff_B_16grj9909_0(.din(w_dff_B_Yz38cpht3_0),.dout(w_dff_B_16grj9909_0),.clk(gclk));
	jdff dff_B_jMmVjyZ13_0(.din(w_dff_B_16grj9909_0),.dout(w_dff_B_jMmVjyZ13_0),.clk(gclk));
	jdff dff_B_kYUGtDk47_0(.din(w_dff_B_jMmVjyZ13_0),.dout(w_dff_B_kYUGtDk47_0),.clk(gclk));
	jdff dff_B_bRt2jkGY6_0(.din(w_dff_B_kYUGtDk47_0),.dout(w_dff_B_bRt2jkGY6_0),.clk(gclk));
	jdff dff_B_1D18vVm55_0(.din(w_dff_B_bRt2jkGY6_0),.dout(w_dff_B_1D18vVm55_0),.clk(gclk));
	jdff dff_B_gq1cU9fC3_0(.din(w_dff_B_1D18vVm55_0),.dout(w_dff_B_gq1cU9fC3_0),.clk(gclk));
	jdff dff_A_XuHGCyMi4_1(.dout(w_n989_0[1]),.din(w_dff_A_XuHGCyMi4_1),.clk(gclk));
	jdff dff_A_3UiLo4Hm1_1(.dout(w_dff_A_XuHGCyMi4_1),.din(w_dff_A_3UiLo4Hm1_1),.clk(gclk));
	jdff dff_A_j4GCz1dc7_1(.dout(w_dff_A_3UiLo4Hm1_1),.din(w_dff_A_j4GCz1dc7_1),.clk(gclk));
	jdff dff_A_Dd14Iau00_1(.dout(w_dff_A_j4GCz1dc7_1),.din(w_dff_A_Dd14Iau00_1),.clk(gclk));
	jdff dff_A_NWcfJXEZ4_1(.dout(w_dff_A_Dd14Iau00_1),.din(w_dff_A_NWcfJXEZ4_1),.clk(gclk));
	jdff dff_B_FXQfZfv44_1(.din(n988),.dout(w_dff_B_FXQfZfv44_1),.clk(gclk));
	jdff dff_B_ZkhZLG0U8_1(.din(w_dff_B_FXQfZfv44_1),.dout(w_dff_B_ZkhZLG0U8_1),.clk(gclk));
	jdff dff_B_6zUhAI5o8_1(.din(w_dff_B_ZkhZLG0U8_1),.dout(w_dff_B_6zUhAI5o8_1),.clk(gclk));
	jdff dff_B_NHWHS9m69_1(.din(w_dff_B_6zUhAI5o8_1),.dout(w_dff_B_NHWHS9m69_1),.clk(gclk));
	jdff dff_B_Yf1OiBcp7_1(.din(w_dff_B_NHWHS9m69_1),.dout(w_dff_B_Yf1OiBcp7_1),.clk(gclk));
	jdff dff_B_sfEVgNFW5_1(.din(w_dff_B_Yf1OiBcp7_1),.dout(w_dff_B_sfEVgNFW5_1),.clk(gclk));
	jdff dff_B_cI72lTST0_1(.din(G112),.dout(w_dff_B_cI72lTST0_1),.clk(gclk));
	jdff dff_B_a73Lzl8l8_1(.din(w_dff_B_cI72lTST0_1),.dout(w_dff_B_a73Lzl8l8_1),.clk(gclk));
	jdff dff_A_YUy9gswz0_0(.dout(w_G1691_3[0]),.din(w_dff_A_YUy9gswz0_0),.clk(gclk));
	jdff dff_A_wJ0rPfhU5_0(.dout(w_dff_A_YUy9gswz0_0),.din(w_dff_A_wJ0rPfhU5_0),.clk(gclk));
	jdff dff_A_IyJKfD3T3_0(.dout(w_dff_A_wJ0rPfhU5_0),.din(w_dff_A_IyJKfD3T3_0),.clk(gclk));
	jdff dff_A_Txew2Vfp7_0(.dout(w_dff_A_IyJKfD3T3_0),.din(w_dff_A_Txew2Vfp7_0),.clk(gclk));
	jdff dff_A_vQklMjXr9_1(.dout(w_G1691_3[1]),.din(w_dff_A_vQklMjXr9_1),.clk(gclk));
	jdff dff_A_dUMO3B2W6_1(.dout(w_dff_A_vQklMjXr9_1),.din(w_dff_A_dUMO3B2W6_1),.clk(gclk));
	jdff dff_B_oiWrOPgC5_1(.din(n1382),.dout(w_dff_B_oiWrOPgC5_1),.clk(gclk));
	jdff dff_B_uPoQbdIH4_1(.din(w_dff_B_oiWrOPgC5_1),.dout(w_dff_B_uPoQbdIH4_1),.clk(gclk));
	jdff dff_B_OBS3g2MD6_1(.din(w_dff_B_uPoQbdIH4_1),.dout(w_dff_B_OBS3g2MD6_1),.clk(gclk));
	jdff dff_B_vRpJerCc7_1(.din(w_dff_B_OBS3g2MD6_1),.dout(w_dff_B_vRpJerCc7_1),.clk(gclk));
	jdff dff_B_eEOFLAnR3_1(.din(w_dff_B_vRpJerCc7_1),.dout(w_dff_B_eEOFLAnR3_1),.clk(gclk));
	jdff dff_B_iG0hA9XB8_1(.din(w_dff_B_eEOFLAnR3_1),.dout(w_dff_B_iG0hA9XB8_1),.clk(gclk));
	jdff dff_B_bLBowyVr4_1(.din(w_dff_B_iG0hA9XB8_1),.dout(w_dff_B_bLBowyVr4_1),.clk(gclk));
	jdff dff_B_Vw1PNlQ50_1(.din(w_dff_B_bLBowyVr4_1),.dout(w_dff_B_Vw1PNlQ50_1),.clk(gclk));
	jdff dff_B_B1Drztfj2_1(.din(w_dff_B_Vw1PNlQ50_1),.dout(w_dff_B_B1Drztfj2_1),.clk(gclk));
	jdff dff_B_s33XO3VT3_1(.din(w_dff_B_B1Drztfj2_1),.dout(w_dff_B_s33XO3VT3_1),.clk(gclk));
	jdff dff_B_Hvj9p1CS1_1(.din(w_dff_B_s33XO3VT3_1),.dout(w_dff_B_Hvj9p1CS1_1),.clk(gclk));
	jdff dff_B_Z0FtxrQn2_1(.din(w_dff_B_Hvj9p1CS1_1),.dout(w_dff_B_Z0FtxrQn2_1),.clk(gclk));
	jdff dff_B_HzCBsusF0_1(.din(w_dff_B_Z0FtxrQn2_1),.dout(w_dff_B_HzCBsusF0_1),.clk(gclk));
	jdff dff_B_n8thrS4o6_1(.din(w_dff_B_HzCBsusF0_1),.dout(w_dff_B_n8thrS4o6_1),.clk(gclk));
	jdff dff_B_y3wcn8El9_1(.din(w_dff_B_n8thrS4o6_1),.dout(w_dff_B_y3wcn8El9_1),.clk(gclk));
	jdff dff_B_FLllfVbz0_1(.din(w_dff_B_y3wcn8El9_1),.dout(w_dff_B_FLllfVbz0_1),.clk(gclk));
	jdff dff_B_FhaLKTVj6_1(.din(w_dff_B_FLllfVbz0_1),.dout(w_dff_B_FhaLKTVj6_1),.clk(gclk));
	jdff dff_B_v0WGhzjX8_1(.din(w_dff_B_FhaLKTVj6_1),.dout(w_dff_B_v0WGhzjX8_1),.clk(gclk));
	jdff dff_B_bzeMK1fT3_1(.din(w_dff_B_v0WGhzjX8_1),.dout(w_dff_B_bzeMK1fT3_1),.clk(gclk));
	jdff dff_B_5IvycdOU8_1(.din(n1245),.dout(w_dff_B_5IvycdOU8_1),.clk(gclk));
	jdff dff_B_vUtVT9m51_1(.din(w_dff_B_5IvycdOU8_1),.dout(w_dff_B_vUtVT9m51_1),.clk(gclk));
	jdff dff_B_ihfIsuao4_1(.din(w_dff_B_vUtVT9m51_1),.dout(w_dff_B_ihfIsuao4_1),.clk(gclk));
	jdff dff_B_VWcK5Uf26_1(.din(w_dff_B_ihfIsuao4_1),.dout(w_dff_B_VWcK5Uf26_1),.clk(gclk));
	jdff dff_B_YyvVml4o9_1(.din(w_dff_B_VWcK5Uf26_1),.dout(w_dff_B_YyvVml4o9_1),.clk(gclk));
	jdff dff_B_Ox1teccs8_1(.din(w_dff_B_YyvVml4o9_1),.dout(w_dff_B_Ox1teccs8_1),.clk(gclk));
	jdff dff_B_IL0nLb354_1(.din(w_dff_B_Ox1teccs8_1),.dout(w_dff_B_IL0nLb354_1),.clk(gclk));
	jdff dff_B_xBqMGKt79_1(.din(w_dff_B_IL0nLb354_1),.dout(w_dff_B_xBqMGKt79_1),.clk(gclk));
	jdff dff_B_TyuQO03d8_1(.din(w_dff_B_xBqMGKt79_1),.dout(w_dff_B_TyuQO03d8_1),.clk(gclk));
	jdff dff_B_PmO4LLJt6_1(.din(w_dff_B_TyuQO03d8_1),.dout(w_dff_B_PmO4LLJt6_1),.clk(gclk));
	jdff dff_B_OH7RfCxk1_1(.din(w_dff_B_PmO4LLJt6_1),.dout(w_dff_B_OH7RfCxk1_1),.clk(gclk));
	jdff dff_B_TY5Sj4AG7_1(.din(w_dff_B_OH7RfCxk1_1),.dout(w_dff_B_TY5Sj4AG7_1),.clk(gclk));
	jdff dff_B_orCNM4oi7_1(.din(w_dff_B_TY5Sj4AG7_1),.dout(w_dff_B_orCNM4oi7_1),.clk(gclk));
	jdff dff_B_YQPpm5Ql9_1(.din(w_dff_B_orCNM4oi7_1),.dout(w_dff_B_YQPpm5Ql9_1),.clk(gclk));
	jdff dff_B_LDa2sPMR3_1(.din(w_dff_B_YQPpm5Ql9_1),.dout(w_dff_B_LDa2sPMR3_1),.clk(gclk));
	jdff dff_B_3gr4XNVP0_1(.din(w_dff_B_LDa2sPMR3_1),.dout(w_dff_B_3gr4XNVP0_1),.clk(gclk));
	jdff dff_B_1UIdvnZ30_1(.din(n1247),.dout(w_dff_B_1UIdvnZ30_1),.clk(gclk));
	jdff dff_B_0dAciVI05_1(.din(w_dff_B_1UIdvnZ30_1),.dout(w_dff_B_0dAciVI05_1),.clk(gclk));
	jdff dff_B_wL4MJtRq5_1(.din(w_dff_B_0dAciVI05_1),.dout(w_dff_B_wL4MJtRq5_1),.clk(gclk));
	jdff dff_B_CnZd14OF3_1(.din(w_dff_B_wL4MJtRq5_1),.dout(w_dff_B_CnZd14OF3_1),.clk(gclk));
	jdff dff_B_1GFeygu12_1(.din(w_dff_B_CnZd14OF3_1),.dout(w_dff_B_1GFeygu12_1),.clk(gclk));
	jdff dff_B_VbEgjxJI3_1(.din(w_dff_B_1GFeygu12_1),.dout(w_dff_B_VbEgjxJI3_1),.clk(gclk));
	jdff dff_B_iWrNKJ1q4_1(.din(w_dff_B_VbEgjxJI3_1),.dout(w_dff_B_iWrNKJ1q4_1),.clk(gclk));
	jdff dff_B_EoFMXOvM4_1(.din(w_dff_B_iWrNKJ1q4_1),.dout(w_dff_B_EoFMXOvM4_1),.clk(gclk));
	jdff dff_B_mecnd2lm6_1(.din(w_dff_B_EoFMXOvM4_1),.dout(w_dff_B_mecnd2lm6_1),.clk(gclk));
	jdff dff_B_pWooJQ6N1_1(.din(w_dff_B_mecnd2lm6_1),.dout(w_dff_B_pWooJQ6N1_1),.clk(gclk));
	jdff dff_B_SpJwA4xT9_1(.din(w_dff_B_pWooJQ6N1_1),.dout(w_dff_B_SpJwA4xT9_1),.clk(gclk));
	jdff dff_B_4aUXaKp82_1(.din(n951),.dout(w_dff_B_4aUXaKp82_1),.clk(gclk));
	jdff dff_B_NSWFAZke9_1(.din(w_dff_B_4aUXaKp82_1),.dout(w_dff_B_NSWFAZke9_1),.clk(gclk));
	jdff dff_B_9FWr1jvA3_1(.din(w_dff_B_NSWFAZke9_1),.dout(w_dff_B_9FWr1jvA3_1),.clk(gclk));
	jdff dff_B_LkMPGFUk7_1(.din(w_dff_B_9FWr1jvA3_1),.dout(w_dff_B_LkMPGFUk7_1),.clk(gclk));
	jdff dff_B_09uUXe1F4_1(.din(w_dff_B_LkMPGFUk7_1),.dout(w_dff_B_09uUXe1F4_1),.clk(gclk));
	jdff dff_B_6miQpeoH1_1(.din(w_dff_B_09uUXe1F4_1),.dout(w_dff_B_6miQpeoH1_1),.clk(gclk));
	jdff dff_B_SUQali7o2_1(.din(w_dff_B_6miQpeoH1_1),.dout(w_dff_B_SUQali7o2_1),.clk(gclk));
	jdff dff_B_TX8TZ7nS5_1(.din(w_dff_B_SUQali7o2_1),.dout(w_dff_B_TX8TZ7nS5_1),.clk(gclk));
	jdff dff_B_ml053Y7a4_1(.din(w_dff_B_TX8TZ7nS5_1),.dout(w_dff_B_ml053Y7a4_1),.clk(gclk));
	jdff dff_B_zM4vQe9H9_1(.din(n513),.dout(w_dff_B_zM4vQe9H9_1),.clk(gclk));
	jdff dff_B_NqMwqEwj1_1(.din(n508),.dout(w_dff_B_NqMwqEwj1_1),.clk(gclk));
	jdff dff_B_uDIAkuJh8_1(.din(G53),.dout(w_dff_B_uDIAkuJh8_1),.clk(gclk));
	jdff dff_B_4Ds4lwDP6_1(.din(w_dff_B_uDIAkuJh8_1),.dout(w_dff_B_4Ds4lwDP6_1),.clk(gclk));
	jdff dff_B_rugrNiAY1_1(.din(n1207),.dout(w_dff_B_rugrNiAY1_1),.clk(gclk));
	jdff dff_B_2GLPIZQU0_1(.din(w_dff_B_rugrNiAY1_1),.dout(w_dff_B_2GLPIZQU0_1),.clk(gclk));
	jdff dff_B_wmJzhUul9_1(.din(w_dff_B_2GLPIZQU0_1),.dout(w_dff_B_wmJzhUul9_1),.clk(gclk));
	jdff dff_B_6iZu3XYm1_1(.din(w_dff_B_wmJzhUul9_1),.dout(w_dff_B_6iZu3XYm1_1),.clk(gclk));
	jdff dff_B_36cErOhx8_1(.din(w_dff_B_6iZu3XYm1_1),.dout(w_dff_B_36cErOhx8_1),.clk(gclk));
	jdff dff_B_hdVA9NAc7_1(.din(w_dff_B_36cErOhx8_1),.dout(w_dff_B_hdVA9NAc7_1),.clk(gclk));
	jdff dff_B_YXFtEMAb1_1(.din(w_dff_B_hdVA9NAc7_1),.dout(w_dff_B_YXFtEMAb1_1),.clk(gclk));
	jdff dff_B_Mdvbhfnk6_1(.din(w_dff_B_YXFtEMAb1_1),.dout(w_dff_B_Mdvbhfnk6_1),.clk(gclk));
	jdff dff_B_BbWxzuR80_1(.din(w_dff_B_Mdvbhfnk6_1),.dout(w_dff_B_BbWxzuR80_1),.clk(gclk));
	jdff dff_B_Vn79ltD42_1(.din(w_dff_B_BbWxzuR80_1),.dout(w_dff_B_Vn79ltD42_1),.clk(gclk));
	jdff dff_B_6ozC2TyU9_1(.din(w_dff_B_Vn79ltD42_1),.dout(w_dff_B_6ozC2TyU9_1),.clk(gclk));
	jdff dff_B_4rAGShJn3_1(.din(w_dff_B_6ozC2TyU9_1),.dout(w_dff_B_4rAGShJn3_1),.clk(gclk));
	jdff dff_B_vlAIQwl63_1(.din(w_dff_B_4rAGShJn3_1),.dout(w_dff_B_vlAIQwl63_1),.clk(gclk));
	jdff dff_B_wMyLAZ3k7_1(.din(w_dff_B_vlAIQwl63_1),.dout(w_dff_B_wMyLAZ3k7_1),.clk(gclk));
	jdff dff_B_Q27boKAz4_1(.din(w_dff_B_wMyLAZ3k7_1),.dout(w_dff_B_Q27boKAz4_1),.clk(gclk));
	jdff dff_B_35MiG9rW5_1(.din(w_dff_B_Q27boKAz4_1),.dout(w_dff_B_35MiG9rW5_1),.clk(gclk));
	jdff dff_B_ir4hScXx5_0(.din(n1211),.dout(w_dff_B_ir4hScXx5_0),.clk(gclk));
	jdff dff_B_obby5ZU81_0(.din(w_dff_B_ir4hScXx5_0),.dout(w_dff_B_obby5ZU81_0),.clk(gclk));
	jdff dff_B_m85n1ZBn4_0(.din(w_dff_B_obby5ZU81_0),.dout(w_dff_B_m85n1ZBn4_0),.clk(gclk));
	jdff dff_B_b8kt6Wkf8_0(.din(w_dff_B_m85n1ZBn4_0),.dout(w_dff_B_b8kt6Wkf8_0),.clk(gclk));
	jdff dff_B_AKBW287S2_0(.din(w_dff_B_b8kt6Wkf8_0),.dout(w_dff_B_AKBW287S2_0),.clk(gclk));
	jdff dff_B_D5xZkAnS0_0(.din(w_dff_B_AKBW287S2_0),.dout(w_dff_B_D5xZkAnS0_0),.clk(gclk));
	jdff dff_B_7EN0PYJH2_0(.din(w_dff_B_D5xZkAnS0_0),.dout(w_dff_B_7EN0PYJH2_0),.clk(gclk));
	jdff dff_B_x5B54nql4_0(.din(w_dff_B_7EN0PYJH2_0),.dout(w_dff_B_x5B54nql4_0),.clk(gclk));
	jdff dff_B_a6DELSnI0_0(.din(w_dff_B_x5B54nql4_0),.dout(w_dff_B_a6DELSnI0_0),.clk(gclk));
	jdff dff_B_UTvvvdCC3_0(.din(w_dff_B_a6DELSnI0_0),.dout(w_dff_B_UTvvvdCC3_0),.clk(gclk));
	jdff dff_B_OAYKGmcQ1_1(.din(n978),.dout(w_dff_B_OAYKGmcQ1_1),.clk(gclk));
	jdff dff_B_CLR5woc61_1(.din(w_dff_B_OAYKGmcQ1_1),.dout(w_dff_B_CLR5woc61_1),.clk(gclk));
	jdff dff_B_XX0ct9dH3_1(.din(w_dff_B_CLR5woc61_1),.dout(w_dff_B_XX0ct9dH3_1),.clk(gclk));
	jdff dff_B_Y7CtRPxk3_1(.din(w_dff_B_XX0ct9dH3_1),.dout(w_dff_B_Y7CtRPxk3_1),.clk(gclk));
	jdff dff_B_KRGjoyy10_1(.din(w_dff_B_Y7CtRPxk3_1),.dout(w_dff_B_KRGjoyy10_1),.clk(gclk));
	jdff dff_B_0E93b3yT7_1(.din(w_dff_B_KRGjoyy10_1),.dout(w_dff_B_0E93b3yT7_1),.clk(gclk));
	jdff dff_B_LYFCAq8x0_1(.din(w_dff_B_0E93b3yT7_1),.dout(w_dff_B_LYFCAq8x0_1),.clk(gclk));
	jdff dff_B_x1Br0cAA6_1(.din(w_dff_B_LYFCAq8x0_1),.dout(w_dff_B_x1Br0cAA6_1),.clk(gclk));
	jdff dff_B_moZESCAc2_1(.din(w_dff_B_x1Br0cAA6_1),.dout(w_dff_B_moZESCAc2_1),.clk(gclk));
	jdff dff_B_u6qAhvxI0_1(.din(n982),.dout(w_dff_B_u6qAhvxI0_1),.clk(gclk));
	jdff dff_B_CqzsS1yo9_1(.din(n980),.dout(w_dff_B_CqzsS1yo9_1),.clk(gclk));
	jdff dff_B_LkPlro0g7_1(.din(w_dff_B_CqzsS1yo9_1),.dout(w_dff_B_LkPlro0g7_1),.clk(gclk));
	jdff dff_B_yOBdlYSZ5_1(.din(w_dff_B_LkPlro0g7_1),.dout(w_dff_B_yOBdlYSZ5_1),.clk(gclk));
	jdff dff_B_1V7xgzM43_1(.din(w_dff_B_yOBdlYSZ5_1),.dout(w_dff_B_1V7xgzM43_1),.clk(gclk));
	jdff dff_B_34l2otit6_1(.din(w_dff_B_1V7xgzM43_1),.dout(w_dff_B_34l2otit6_1),.clk(gclk));
	jdff dff_B_H0lVh1nh9_1(.din(G116),.dout(w_dff_B_H0lVh1nh9_1),.clk(gclk));
	jdff dff_B_QvouAMqL3_1(.din(w_dff_B_H0lVh1nh9_1),.dout(w_dff_B_QvouAMqL3_1),.clk(gclk));
	jdff dff_B_8OPEYJCD1_0(.din(n1381),.dout(w_dff_B_8OPEYJCD1_0),.clk(gclk));
	jdff dff_B_neZGfiL07_2(.din(G167),.dout(w_dff_B_neZGfiL07_2),.clk(gclk));
	jdff dff_B_ZnjI2Mea3_2(.din(G197),.dout(w_dff_B_ZnjI2Mea3_2),.clk(gclk));
	jdff dff_B_F37cIesD2_2(.din(w_dff_B_ZnjI2Mea3_2),.dout(w_dff_B_F37cIesD2_2),.clk(gclk));
	jdff dff_B_NJKycKug6_0(.din(n1395),.dout(w_dff_B_NJKycKug6_0),.clk(gclk));
	jdff dff_B_XaZ9PEMo0_0(.din(w_dff_B_NJKycKug6_0),.dout(w_dff_B_XaZ9PEMo0_0),.clk(gclk));
	jdff dff_B_XVgbybfh2_0(.din(w_dff_B_XaZ9PEMo0_0),.dout(w_dff_B_XVgbybfh2_0),.clk(gclk));
	jdff dff_B_GY20Zzwl9_0(.din(w_dff_B_XVgbybfh2_0),.dout(w_dff_B_GY20Zzwl9_0),.clk(gclk));
	jdff dff_B_12NrCWhL7_0(.din(w_dff_B_GY20Zzwl9_0),.dout(w_dff_B_12NrCWhL7_0),.clk(gclk));
	jdff dff_B_LIThVoW39_0(.din(w_dff_B_12NrCWhL7_0),.dout(w_dff_B_LIThVoW39_0),.clk(gclk));
	jdff dff_B_yV6ugsuj1_0(.din(w_dff_B_LIThVoW39_0),.dout(w_dff_B_yV6ugsuj1_0),.clk(gclk));
	jdff dff_B_xmSoYhIA3_0(.din(w_dff_B_yV6ugsuj1_0),.dout(w_dff_B_xmSoYhIA3_0),.clk(gclk));
	jdff dff_B_xIb444Sp1_0(.din(w_dff_B_xmSoYhIA3_0),.dout(w_dff_B_xIb444Sp1_0),.clk(gclk));
	jdff dff_B_w8M16BaX6_0(.din(w_dff_B_xIb444Sp1_0),.dout(w_dff_B_w8M16BaX6_0),.clk(gclk));
	jdff dff_B_ZP7sJByb6_0(.din(w_dff_B_w8M16BaX6_0),.dout(w_dff_B_ZP7sJByb6_0),.clk(gclk));
	jdff dff_B_mxeqjROu1_0(.din(w_dff_B_ZP7sJByb6_0),.dout(w_dff_B_mxeqjROu1_0),.clk(gclk));
	jdff dff_B_dR9Cj0wd5_0(.din(w_dff_B_mxeqjROu1_0),.dout(w_dff_B_dR9Cj0wd5_0),.clk(gclk));
	jdff dff_B_8R29XEmq1_0(.din(w_dff_B_dR9Cj0wd5_0),.dout(w_dff_B_8R29XEmq1_0),.clk(gclk));
	jdff dff_B_3t0ytUIN2_0(.din(w_dff_B_8R29XEmq1_0),.dout(w_dff_B_3t0ytUIN2_0),.clk(gclk));
	jdff dff_B_VdFA3uXc8_0(.din(w_dff_B_3t0ytUIN2_0),.dout(w_dff_B_VdFA3uXc8_0),.clk(gclk));
	jdff dff_B_zBOwiPRE2_0(.din(w_dff_B_VdFA3uXc8_0),.dout(w_dff_B_zBOwiPRE2_0),.clk(gclk));
	jdff dff_B_R9I2p3F84_0(.din(w_dff_B_zBOwiPRE2_0),.dout(w_dff_B_R9I2p3F84_0),.clk(gclk));
	jdff dff_B_c0egVQFZ4_0(.din(w_dff_B_R9I2p3F84_0),.dout(w_dff_B_c0egVQFZ4_0),.clk(gclk));
	jdff dff_B_fv6coIyT0_0(.din(n1394),.dout(w_dff_B_fv6coIyT0_0),.clk(gclk));
	jdff dff_B_ZtJzWLSh7_2(.din(G164),.dout(w_dff_B_ZtJzWLSh7_2),.clk(gclk));
	jdff dff_B_yNKzXfDQ4_2(.din(G194),.dout(w_dff_B_yNKzXfDQ4_2),.clk(gclk));
	jdff dff_B_TFS1KFt26_2(.din(w_dff_B_yNKzXfDQ4_2),.dout(w_dff_B_TFS1KFt26_2),.clk(gclk));
	jdff dff_B_5R8yb2h83_1(.din(n1389),.dout(w_dff_B_5R8yb2h83_1),.clk(gclk));
	jdff dff_B_MuWztHRc9_1(.din(w_dff_B_5R8yb2h83_1),.dout(w_dff_B_MuWztHRc9_1),.clk(gclk));
	jdff dff_B_47rOcSoE7_1(.din(n1239),.dout(w_dff_B_47rOcSoE7_1),.clk(gclk));
	jdff dff_B_2mtnGLZK5_1(.din(w_dff_B_47rOcSoE7_1),.dout(w_dff_B_2mtnGLZK5_1),.clk(gclk));
	jdff dff_B_BzZH3Vxg6_1(.din(w_dff_B_2mtnGLZK5_1),.dout(w_dff_B_BzZH3Vxg6_1),.clk(gclk));
	jdff dff_B_HIwuIvE63_1(.din(w_dff_B_BzZH3Vxg6_1),.dout(w_dff_B_HIwuIvE63_1),.clk(gclk));
	jdff dff_B_aTWj3rFY0_1(.din(w_dff_B_HIwuIvE63_1),.dout(w_dff_B_aTWj3rFY0_1),.clk(gclk));
	jdff dff_B_tU45p0v45_1(.din(w_dff_B_aTWj3rFY0_1),.dout(w_dff_B_tU45p0v45_1),.clk(gclk));
	jdff dff_B_thUqQi0U2_1(.din(w_dff_B_tU45p0v45_1),.dout(w_dff_B_thUqQi0U2_1),.clk(gclk));
	jdff dff_B_G6K8jEA21_1(.din(w_dff_B_thUqQi0U2_1),.dout(w_dff_B_G6K8jEA21_1),.clk(gclk));
	jdff dff_B_BFwHCQF72_1(.din(w_dff_B_G6K8jEA21_1),.dout(w_dff_B_BFwHCQF72_1),.clk(gclk));
	jdff dff_B_KcQfyADH8_1(.din(w_dff_B_BFwHCQF72_1),.dout(w_dff_B_KcQfyADH8_1),.clk(gclk));
	jdff dff_B_4WokPKmk0_1(.din(w_dff_B_KcQfyADH8_1),.dout(w_dff_B_4WokPKmk0_1),.clk(gclk));
	jdff dff_B_BUurbvki8_1(.din(w_dff_B_4WokPKmk0_1),.dout(w_dff_B_BUurbvki8_1),.clk(gclk));
	jdff dff_B_U2AdnZx40_1(.din(w_dff_B_BUurbvki8_1),.dout(w_dff_B_U2AdnZx40_1),.clk(gclk));
	jdff dff_B_6vS3LmRH4_1(.din(w_dff_B_U2AdnZx40_1),.dout(w_dff_B_6vS3LmRH4_1),.clk(gclk));
	jdff dff_B_4K2baa6I4_0(.din(n1242),.dout(w_dff_B_4K2baa6I4_0),.clk(gclk));
	jdff dff_B_EP8hHyTu6_0(.din(w_dff_B_4K2baa6I4_0),.dout(w_dff_B_EP8hHyTu6_0),.clk(gclk));
	jdff dff_B_9rBKJiMz1_0(.din(w_dff_B_EP8hHyTu6_0),.dout(w_dff_B_9rBKJiMz1_0),.clk(gclk));
	jdff dff_B_bKCYm0Lj0_0(.din(w_dff_B_9rBKJiMz1_0),.dout(w_dff_B_bKCYm0Lj0_0),.clk(gclk));
	jdff dff_B_ygQFlegl9_0(.din(w_dff_B_bKCYm0Lj0_0),.dout(w_dff_B_ygQFlegl9_0),.clk(gclk));
	jdff dff_B_qGnB5wcK3_0(.din(w_dff_B_ygQFlegl9_0),.dout(w_dff_B_qGnB5wcK3_0),.clk(gclk));
	jdff dff_B_FIvrXbRt6_0(.din(w_dff_B_qGnB5wcK3_0),.dout(w_dff_B_FIvrXbRt6_0),.clk(gclk));
	jdff dff_B_PWAiMeGW4_0(.din(w_dff_B_FIvrXbRt6_0),.dout(w_dff_B_PWAiMeGW4_0),.clk(gclk));
	jdff dff_B_GwYmBqHV9_0(.din(w_dff_B_PWAiMeGW4_0),.dout(w_dff_B_GwYmBqHV9_0),.clk(gclk));
	jdff dff_B_QRj5i3yC5_0(.din(w_dff_B_GwYmBqHV9_0),.dout(w_dff_B_QRj5i3yC5_0),.clk(gclk));
	jdff dff_A_jnYcwbEQ9_1(.dout(w_n459_0[1]),.din(w_dff_A_jnYcwbEQ9_1),.clk(gclk));
	jdff dff_A_EUTT2E089_1(.dout(w_dff_A_jnYcwbEQ9_1),.din(w_dff_A_EUTT2E089_1),.clk(gclk));
	jdff dff_A_WtRAsExu8_1(.dout(w_dff_A_EUTT2E089_1),.din(w_dff_A_WtRAsExu8_1),.clk(gclk));
	jdff dff_B_zSbUmewt1_1(.din(n455),.dout(w_dff_B_zSbUmewt1_1),.clk(gclk));
	jdff dff_B_whIVPNaU5_3(.din(G3548),.dout(w_dff_B_whIVPNaU5_3),.clk(gclk));
	jdff dff_B_19v3Jvts2_1(.din(n450),.dout(w_dff_B_19v3Jvts2_1),.clk(gclk));
	jdff dff_A_nlNa4cWH9_0(.dout(w_n749_6[0]),.din(w_dff_A_nlNa4cWH9_0),.clk(gclk));
	jdff dff_A_KMteQsiu9_0(.dout(w_dff_A_nlNa4cWH9_0),.din(w_dff_A_KMteQsiu9_0),.clk(gclk));
	jdff dff_A_okgQU3dp8_0(.dout(w_dff_A_KMteQsiu9_0),.din(w_dff_A_okgQU3dp8_0),.clk(gclk));
	jdff dff_A_qxrxUja80_0(.dout(w_dff_A_okgQU3dp8_0),.din(w_dff_A_qxrxUja80_0),.clk(gclk));
	jdff dff_A_kfHq47ow2_0(.dout(w_dff_A_qxrxUja80_0),.din(w_dff_A_kfHq47ow2_0),.clk(gclk));
	jdff dff_A_FNeIz5LM0_0(.dout(w_dff_A_kfHq47ow2_0),.din(w_dff_A_FNeIz5LM0_0),.clk(gclk));
	jdff dff_A_r2kxfEzD2_0(.dout(w_dff_A_FNeIz5LM0_0),.din(w_dff_A_r2kxfEzD2_0),.clk(gclk));
	jdff dff_A_k7px8ZIV7_0(.dout(w_dff_A_r2kxfEzD2_0),.din(w_dff_A_k7px8ZIV7_0),.clk(gclk));
	jdff dff_A_LtgjpQ8i8_0(.dout(w_dff_A_k7px8ZIV7_0),.din(w_dff_A_LtgjpQ8i8_0),.clk(gclk));
	jdff dff_A_U321d9H42_0(.dout(w_dff_A_LtgjpQ8i8_0),.din(w_dff_A_U321d9H42_0),.clk(gclk));
	jdff dff_A_9QojdME74_0(.dout(w_dff_A_U321d9H42_0),.din(w_dff_A_9QojdME74_0),.clk(gclk));
	jdff dff_A_nZtcsZiB6_1(.dout(w_n949_0[1]),.din(w_dff_A_nZtcsZiB6_1),.clk(gclk));
	jdff dff_A_DN6DoIr47_1(.dout(w_dff_A_nZtcsZiB6_1),.din(w_dff_A_DN6DoIr47_1),.clk(gclk));
	jdff dff_B_LI1JA4KH8_1(.din(n946),.dout(w_dff_B_LI1JA4KH8_1),.clk(gclk));
	jdff dff_B_2FIk3Z3e5_1(.din(w_dff_B_LI1JA4KH8_1),.dout(w_dff_B_2FIk3Z3e5_1),.clk(gclk));
	jdff dff_B_DTvxGPpS9_1(.din(w_dff_B_2FIk3Z3e5_1),.dout(w_dff_B_DTvxGPpS9_1),.clk(gclk));
	jdff dff_B_i6u3ojuc0_1(.din(w_dff_B_DTvxGPpS9_1),.dout(w_dff_B_i6u3ojuc0_1),.clk(gclk));
	jdff dff_B_mtLjG21W7_1(.din(w_dff_B_i6u3ojuc0_1),.dout(w_dff_B_mtLjG21W7_1),.clk(gclk));
	jdff dff_B_myCJoxAL4_1(.din(w_dff_B_mtLjG21W7_1),.dout(w_dff_B_myCJoxAL4_1),.clk(gclk));
	jdff dff_A_81UxL76d2_0(.dout(w_G4091_2[0]),.din(w_dff_A_81UxL76d2_0),.clk(gclk));
	jdff dff_A_Biw7FZMg8_0(.dout(w_dff_A_81UxL76d2_0),.din(w_dff_A_Biw7FZMg8_0),.clk(gclk));
	jdff dff_A_wZafjZe65_1(.dout(w_G4091_2[1]),.din(w_dff_A_wZafjZe65_1),.clk(gclk));
	jdff dff_A_PYSskl8b8_1(.dout(w_dff_A_wZafjZe65_1),.din(w_dff_A_PYSskl8b8_1),.clk(gclk));
	jdff dff_A_mOsICq916_1(.dout(w_dff_A_PYSskl8b8_1),.din(w_dff_A_mOsICq916_1),.clk(gclk));
	jdff dff_B_QHGv122k0_1(.din(G114),.dout(w_dff_B_QHGv122k0_1),.clk(gclk));
	jdff dff_B_vTfpB1Oo6_1(.din(w_dff_B_QHGv122k0_1),.dout(w_dff_B_vTfpB1Oo6_1),.clk(gclk));
	jdff dff_A_gg4BFt0t4_0(.dout(w_n1008_2[0]),.din(w_dff_A_gg4BFt0t4_0),.clk(gclk));
	jdff dff_A_4itjFJvj8_1(.dout(w_n1008_2[1]),.din(w_dff_A_4itjFJvj8_1),.clk(gclk));
	jdff dff_B_qUj5qikX1_1(.din(n1198),.dout(w_dff_B_qUj5qikX1_1),.clk(gclk));
	jdff dff_B_soXvq5cY5_1(.din(w_dff_B_qUj5qikX1_1),.dout(w_dff_B_soXvq5cY5_1),.clk(gclk));
	jdff dff_B_FA1bullw2_1(.din(w_dff_B_soXvq5cY5_1),.dout(w_dff_B_FA1bullw2_1),.clk(gclk));
	jdff dff_B_GB4S7wDx5_1(.din(w_dff_B_FA1bullw2_1),.dout(w_dff_B_GB4S7wDx5_1),.clk(gclk));
	jdff dff_B_yztnDgi42_1(.din(w_dff_B_GB4S7wDx5_1),.dout(w_dff_B_yztnDgi42_1),.clk(gclk));
	jdff dff_B_okmNacrg6_1(.din(w_dff_B_yztnDgi42_1),.dout(w_dff_B_okmNacrg6_1),.clk(gclk));
	jdff dff_B_BcDB7RYW2_1(.din(w_dff_B_okmNacrg6_1),.dout(w_dff_B_BcDB7RYW2_1),.clk(gclk));
	jdff dff_B_I5N7PxVN3_1(.din(w_dff_B_BcDB7RYW2_1),.dout(w_dff_B_I5N7PxVN3_1),.clk(gclk));
	jdff dff_B_YFyVXOaN4_1(.din(w_dff_B_I5N7PxVN3_1),.dout(w_dff_B_YFyVXOaN4_1),.clk(gclk));
	jdff dff_B_Ks4m6jrm6_1(.din(w_dff_B_YFyVXOaN4_1),.dout(w_dff_B_Ks4m6jrm6_1),.clk(gclk));
	jdff dff_B_YzEV7fZk4_1(.din(w_dff_B_Ks4m6jrm6_1),.dout(w_dff_B_YzEV7fZk4_1),.clk(gclk));
	jdff dff_B_6ciOveFz7_1(.din(w_dff_B_YzEV7fZk4_1),.dout(w_dff_B_6ciOveFz7_1),.clk(gclk));
	jdff dff_B_YGLLw1ly6_1(.din(w_dff_B_6ciOveFz7_1),.dout(w_dff_B_YGLLw1ly6_1),.clk(gclk));
	jdff dff_B_knVKXUQD9_1(.din(w_dff_B_YGLLw1ly6_1),.dout(w_dff_B_knVKXUQD9_1),.clk(gclk));
	jdff dff_B_JnMTqY8m2_1(.din(w_dff_B_knVKXUQD9_1),.dout(w_dff_B_JnMTqY8m2_1),.clk(gclk));
	jdff dff_B_hq34FAy57_1(.din(n1200),.dout(w_dff_B_hq34FAy57_1),.clk(gclk));
	jdff dff_B_s074vNxE3_1(.din(w_dff_B_hq34FAy57_1),.dout(w_dff_B_s074vNxE3_1),.clk(gclk));
	jdff dff_B_hrsDR4cm0_1(.din(w_dff_B_s074vNxE3_1),.dout(w_dff_B_hrsDR4cm0_1),.clk(gclk));
	jdff dff_B_TqwmG5rH1_1(.din(w_dff_B_hrsDR4cm0_1),.dout(w_dff_B_TqwmG5rH1_1),.clk(gclk));
	jdff dff_B_grEZ1lrA2_1(.din(w_dff_B_TqwmG5rH1_1),.dout(w_dff_B_grEZ1lrA2_1),.clk(gclk));
	jdff dff_B_xPtK0Ird3_1(.din(w_dff_B_grEZ1lrA2_1),.dout(w_dff_B_xPtK0Ird3_1),.clk(gclk));
	jdff dff_B_BbqvFFVD4_1(.din(w_dff_B_xPtK0Ird3_1),.dout(w_dff_B_BbqvFFVD4_1),.clk(gclk));
	jdff dff_B_PrYZA3Vf6_1(.din(w_dff_B_BbqvFFVD4_1),.dout(w_dff_B_PrYZA3Vf6_1),.clk(gclk));
	jdff dff_B_AGpDPeXA6_1(.din(w_dff_B_PrYZA3Vf6_1),.dout(w_dff_B_AGpDPeXA6_1),.clk(gclk));
	jdff dff_B_viVeim727_1(.din(w_dff_B_AGpDPeXA6_1),.dout(w_dff_B_viVeim727_1),.clk(gclk));
	jdff dff_B_n8YfteQh9_1(.din(w_dff_B_viVeim727_1),.dout(w_dff_B_n8YfteQh9_1),.clk(gclk));
	jdff dff_A_48Lg9FeE2_0(.dout(w_n649_0[0]),.din(w_dff_A_48Lg9FeE2_0),.clk(gclk));
	jdff dff_A_PmrJgT1l0_0(.dout(w_dff_A_48Lg9FeE2_0),.din(w_dff_A_PmrJgT1l0_0),.clk(gclk));
	jdff dff_A_OvYhlNeR9_0(.dout(w_dff_A_PmrJgT1l0_0),.din(w_dff_A_OvYhlNeR9_0),.clk(gclk));
	jdff dff_A_Ht6mC1u15_0(.dout(w_dff_A_OvYhlNeR9_0),.din(w_dff_A_Ht6mC1u15_0),.clk(gclk));
	jdff dff_A_CPPaZf2j7_0(.dout(w_dff_A_Ht6mC1u15_0),.din(w_dff_A_CPPaZf2j7_0),.clk(gclk));
	jdff dff_A_kD5OqBHZ5_0(.dout(w_dff_A_CPPaZf2j7_0),.din(w_dff_A_kD5OqBHZ5_0),.clk(gclk));
	jdff dff_A_HuO9a9D43_0(.dout(w_dff_A_kD5OqBHZ5_0),.din(w_dff_A_HuO9a9D43_0),.clk(gclk));
	jdff dff_A_VhgcBHLo4_0(.dout(w_dff_A_HuO9a9D43_0),.din(w_dff_A_VhgcBHLo4_0),.clk(gclk));
	jdff dff_A_RofdZU6q4_0(.dout(w_dff_A_VhgcBHLo4_0),.din(w_dff_A_RofdZU6q4_0),.clk(gclk));
	jdff dff_A_Z2uzUbwh6_1(.dout(w_n749_8[1]),.din(w_dff_A_Z2uzUbwh6_1),.clk(gclk));
	jdff dff_A_u4BSjaXN8_1(.dout(w_dff_A_Z2uzUbwh6_1),.din(w_dff_A_u4BSjaXN8_1),.clk(gclk));
	jdff dff_A_amWxjfOZ8_1(.dout(w_dff_A_u4BSjaXN8_1),.din(w_dff_A_amWxjfOZ8_1),.clk(gclk));
	jdff dff_A_JHdr3CR71_1(.dout(w_dff_A_amWxjfOZ8_1),.din(w_dff_A_JHdr3CR71_1),.clk(gclk));
	jdff dff_A_VlXlr4Zx1_1(.dout(w_dff_A_JHdr3CR71_1),.din(w_dff_A_VlXlr4Zx1_1),.clk(gclk));
	jdff dff_A_EKaufpOh9_1(.dout(w_dff_A_VlXlr4Zx1_1),.din(w_dff_A_EKaufpOh9_1),.clk(gclk));
	jdff dff_A_bz1X9iPL0_1(.dout(w_dff_A_EKaufpOh9_1),.din(w_dff_A_bz1X9iPL0_1),.clk(gclk));
	jdff dff_A_slPUXqXl0_1(.dout(w_dff_A_bz1X9iPL0_1),.din(w_dff_A_slPUXqXl0_1),.clk(gclk));
	jdff dff_A_p4crpk3Y4_1(.dout(w_dff_A_slPUXqXl0_1),.din(w_dff_A_p4crpk3Y4_1),.clk(gclk));
	jdff dff_A_2Aco52Z85_1(.dout(w_dff_A_p4crpk3Y4_1),.din(w_dff_A_2Aco52Z85_1),.clk(gclk));
	jdff dff_A_rCM9b6PR0_1(.dout(w_dff_A_2Aco52Z85_1),.din(w_dff_A_rCM9b6PR0_1),.clk(gclk));
	jdff dff_A_dIDY0ASi7_1(.dout(w_dff_A_rCM9b6PR0_1),.din(w_dff_A_dIDY0ASi7_1),.clk(gclk));
	jdff dff_A_QEtZXnjq8_2(.dout(w_n749_8[2]),.din(w_dff_A_QEtZXnjq8_2),.clk(gclk));
	jdff dff_A_nD2zMoYV7_2(.dout(w_dff_A_QEtZXnjq8_2),.din(w_dff_A_nD2zMoYV7_2),.clk(gclk));
	jdff dff_A_n9UM1KJa2_2(.dout(w_dff_A_nD2zMoYV7_2),.din(w_dff_A_n9UM1KJa2_2),.clk(gclk));
	jdff dff_A_XC1Ky63H8_2(.dout(w_dff_A_n9UM1KJa2_2),.din(w_dff_A_XC1Ky63H8_2),.clk(gclk));
	jdff dff_A_ahjHc97C7_2(.dout(w_dff_A_XC1Ky63H8_2),.din(w_dff_A_ahjHc97C7_2),.clk(gclk));
	jdff dff_A_eu1v8Eyz1_2(.dout(w_dff_A_ahjHc97C7_2),.din(w_dff_A_eu1v8Eyz1_2),.clk(gclk));
	jdff dff_A_AOUMzYVg1_2(.dout(w_dff_A_eu1v8Eyz1_2),.din(w_dff_A_AOUMzYVg1_2),.clk(gclk));
	jdff dff_A_bLirk2oD2_2(.dout(w_dff_A_AOUMzYVg1_2),.din(w_dff_A_bLirk2oD2_2),.clk(gclk));
	jdff dff_A_EJRghaxr4_2(.dout(w_dff_A_bLirk2oD2_2),.din(w_dff_A_EJRghaxr4_2),.clk(gclk));
	jdff dff_A_tTXFHE0C8_2(.dout(w_dff_A_EJRghaxr4_2),.din(w_dff_A_tTXFHE0C8_2),.clk(gclk));
	jdff dff_B_RxFp7TsG0_1(.din(G121),.dout(w_dff_B_RxFp7TsG0_1),.clk(gclk));
	jdff dff_B_znfhQR8X5_1(.din(w_dff_B_RxFp7TsG0_1),.dout(w_dff_B_znfhQR8X5_1),.clk(gclk));
	jdff dff_A_7MpZfYVu0_0(.dout(w_G137_4[0]),.din(w_dff_A_7MpZfYVu0_0),.clk(gclk));
	jdff dff_A_twaGs9Zc4_1(.dout(w_G137_4[1]),.din(w_dff_A_twaGs9Zc4_1),.clk(gclk));
	jdff dff_A_2ZJ92eYq8_0(.dout(w_G137_1[0]),.din(w_dff_A_2ZJ92eYq8_0),.clk(gclk));
	jdff dff_A_NEQHZNTm8_0(.dout(w_dff_A_2ZJ92eYq8_0),.din(w_dff_A_NEQHZNTm8_0),.clk(gclk));
	jdff dff_A_48O7lkU96_0(.dout(w_dff_A_NEQHZNTm8_0),.din(w_dff_A_48O7lkU96_0),.clk(gclk));
	jdff dff_A_7bQf64Kj1_0(.dout(w_dff_A_48O7lkU96_0),.din(w_dff_A_7bQf64Kj1_0),.clk(gclk));
	jdff dff_A_6P2fUvRx9_0(.dout(w_dff_A_7bQf64Kj1_0),.din(w_dff_A_6P2fUvRx9_0),.clk(gclk));
	jdff dff_A_tDErR2Fk5_0(.dout(w_dff_A_6P2fUvRx9_0),.din(w_dff_A_tDErR2Fk5_0),.clk(gclk));
	jdff dff_A_LdXCM8TE3_1(.dout(w_G137_1[1]),.din(w_dff_A_LdXCM8TE3_1),.clk(gclk));
	jdff dff_A_5pjFRJaM5_1(.dout(w_dff_A_LdXCM8TE3_1),.din(w_dff_A_5pjFRJaM5_1),.clk(gclk));
	jdff dff_A_LFNYy1Rz5_1(.dout(w_dff_A_5pjFRJaM5_1),.din(w_dff_A_LFNYy1Rz5_1),.clk(gclk));
	jdff dff_A_J5bUeEfp8_1(.dout(w_dff_A_LFNYy1Rz5_1),.din(w_dff_A_J5bUeEfp8_1),.clk(gclk));
	jdff dff_A_x9SmHMpY2_1(.dout(w_dff_A_J5bUeEfp8_1),.din(w_dff_A_x9SmHMpY2_1),.clk(gclk));
	jdff dff_A_E2TeOGMc6_1(.dout(w_dff_A_x9SmHMpY2_1),.din(w_dff_A_E2TeOGMc6_1),.clk(gclk));
	jdff dff_A_BlHPAdPJ1_1(.dout(w_dff_A_E2TeOGMc6_1),.din(w_dff_A_BlHPAdPJ1_1),.clk(gclk));
	jdff dff_B_cxjMtlJw8_0(.din(n1404),.dout(w_dff_B_cxjMtlJw8_0),.clk(gclk));
	jdff dff_B_bZ5cU1fT1_0(.din(w_dff_B_cxjMtlJw8_0),.dout(w_dff_B_bZ5cU1fT1_0),.clk(gclk));
	jdff dff_B_tsEXBXId4_0(.din(w_dff_B_bZ5cU1fT1_0),.dout(w_dff_B_tsEXBXId4_0),.clk(gclk));
	jdff dff_B_ffqNDHdl9_0(.din(w_dff_B_tsEXBXId4_0),.dout(w_dff_B_ffqNDHdl9_0),.clk(gclk));
	jdff dff_B_ckBadHMd5_0(.din(w_dff_B_ffqNDHdl9_0),.dout(w_dff_B_ckBadHMd5_0),.clk(gclk));
	jdff dff_B_hib07Wuo9_0(.din(w_dff_B_ckBadHMd5_0),.dout(w_dff_B_hib07Wuo9_0),.clk(gclk));
	jdff dff_B_lFNrILTE4_0(.din(w_dff_B_hib07Wuo9_0),.dout(w_dff_B_lFNrILTE4_0),.clk(gclk));
	jdff dff_B_rl3MElyJ5_0(.din(w_dff_B_lFNrILTE4_0),.dout(w_dff_B_rl3MElyJ5_0),.clk(gclk));
	jdff dff_B_6dzn9GO70_0(.din(w_dff_B_rl3MElyJ5_0),.dout(w_dff_B_6dzn9GO70_0),.clk(gclk));
	jdff dff_B_bZRkqF2K7_0(.din(w_dff_B_6dzn9GO70_0),.dout(w_dff_B_bZRkqF2K7_0),.clk(gclk));
	jdff dff_B_GR5fnkDR0_0(.din(w_dff_B_bZRkqF2K7_0),.dout(w_dff_B_GR5fnkDR0_0),.clk(gclk));
	jdff dff_B_Tz2X3wya2_0(.din(w_dff_B_GR5fnkDR0_0),.dout(w_dff_B_Tz2X3wya2_0),.clk(gclk));
	jdff dff_B_33A2G5uo7_0(.din(w_dff_B_Tz2X3wya2_0),.dout(w_dff_B_33A2G5uo7_0),.clk(gclk));
	jdff dff_B_XoFoH3AL8_0(.din(w_dff_B_33A2G5uo7_0),.dout(w_dff_B_XoFoH3AL8_0),.clk(gclk));
	jdff dff_B_ZS5T9I4M9_0(.din(w_dff_B_XoFoH3AL8_0),.dout(w_dff_B_ZS5T9I4M9_0),.clk(gclk));
	jdff dff_B_TO8jWDqr6_0(.din(w_dff_B_ZS5T9I4M9_0),.dout(w_dff_B_TO8jWDqr6_0),.clk(gclk));
	jdff dff_B_wvWJ9g7h6_0(.din(w_dff_B_TO8jWDqr6_0),.dout(w_dff_B_wvWJ9g7h6_0),.clk(gclk));
	jdff dff_B_m3ss79Mj7_0(.din(w_dff_B_wvWJ9g7h6_0),.dout(w_dff_B_m3ss79Mj7_0),.clk(gclk));
	jdff dff_B_pD1sRVPu5_0(.din(w_dff_B_m3ss79Mj7_0),.dout(w_dff_B_pD1sRVPu5_0),.clk(gclk));
	jdff dff_B_Q00mXVOW6_0(.din(n1403),.dout(w_dff_B_Q00mXVOW6_0),.clk(gclk));
	jdff dff_B_Gd68TiCk6_2(.din(G161),.dout(w_dff_B_Gd68TiCk6_2),.clk(gclk));
	jdff dff_B_O0W6fqH48_2(.din(G191),.dout(w_dff_B_O0W6fqH48_2),.clk(gclk));
	jdff dff_B_tFRk1qYy6_2(.din(w_dff_B_O0W6fqH48_2),.dout(w_dff_B_tFRk1qYy6_2),.clk(gclk));
	jdff dff_B_qYaEM9A89_1(.din(n1190),.dout(w_dff_B_qYaEM9A89_1),.clk(gclk));
	jdff dff_B_HcIJJcHd9_1(.din(w_dff_B_qYaEM9A89_1),.dout(w_dff_B_HcIJJcHd9_1),.clk(gclk));
	jdff dff_B_O0DIQGRk2_1(.din(w_dff_B_HcIJJcHd9_1),.dout(w_dff_B_O0DIQGRk2_1),.clk(gclk));
	jdff dff_B_yld60UzA6_1(.din(w_dff_B_O0DIQGRk2_1),.dout(w_dff_B_yld60UzA6_1),.clk(gclk));
	jdff dff_B_3IgSQrui5_1(.din(w_dff_B_yld60UzA6_1),.dout(w_dff_B_3IgSQrui5_1),.clk(gclk));
	jdff dff_B_qiOAYz3y8_1(.din(w_dff_B_3IgSQrui5_1),.dout(w_dff_B_qiOAYz3y8_1),.clk(gclk));
	jdff dff_B_WlieLL8S0_1(.din(w_dff_B_qiOAYz3y8_1),.dout(w_dff_B_WlieLL8S0_1),.clk(gclk));
	jdff dff_B_NpWqOmwQ7_1(.din(w_dff_B_WlieLL8S0_1),.dout(w_dff_B_NpWqOmwQ7_1),.clk(gclk));
	jdff dff_B_ASSwQiPh3_1(.din(w_dff_B_NpWqOmwQ7_1),.dout(w_dff_B_ASSwQiPh3_1),.clk(gclk));
	jdff dff_B_38TLV40j6_1(.din(w_dff_B_ASSwQiPh3_1),.dout(w_dff_B_38TLV40j6_1),.clk(gclk));
	jdff dff_B_lzFDADZH4_1(.din(w_dff_B_38TLV40j6_1),.dout(w_dff_B_lzFDADZH4_1),.clk(gclk));
	jdff dff_B_PDh3NrwN4_1(.din(w_dff_B_lzFDADZH4_1),.dout(w_dff_B_PDh3NrwN4_1),.clk(gclk));
	jdff dff_B_4G2NvpMz1_1(.din(w_dff_B_PDh3NrwN4_1),.dout(w_dff_B_4G2NvpMz1_1),.clk(gclk));
	jdff dff_B_u6HFsEeJ0_1(.din(w_dff_B_4G2NvpMz1_1),.dout(w_dff_B_u6HFsEeJ0_1),.clk(gclk));
	jdff dff_B_HwXft9pr8_1(.din(w_dff_B_u6HFsEeJ0_1),.dout(w_dff_B_HwXft9pr8_1),.clk(gclk));
	jdff dff_B_AMKwCWI48_1(.din(w_dff_B_HwXft9pr8_1),.dout(w_dff_B_AMKwCWI48_1),.clk(gclk));
	jdff dff_B_sN7HnCoS3_0(.din(n1194),.dout(w_dff_B_sN7HnCoS3_0),.clk(gclk));
	jdff dff_B_dztaGO7m3_0(.din(w_dff_B_sN7HnCoS3_0),.dout(w_dff_B_dztaGO7m3_0),.clk(gclk));
	jdff dff_B_vRp4HNDj0_0(.din(w_dff_B_dztaGO7m3_0),.dout(w_dff_B_vRp4HNDj0_0),.clk(gclk));
	jdff dff_B_sAM8TalL7_0(.din(w_dff_B_vRp4HNDj0_0),.dout(w_dff_B_sAM8TalL7_0),.clk(gclk));
	jdff dff_B_EorSIbqx9_0(.din(w_dff_B_sAM8TalL7_0),.dout(w_dff_B_EorSIbqx9_0),.clk(gclk));
	jdff dff_B_5XM3uvJJ3_0(.din(w_dff_B_EorSIbqx9_0),.dout(w_dff_B_5XM3uvJJ3_0),.clk(gclk));
	jdff dff_B_zOyDH3mQ8_0(.din(w_dff_B_5XM3uvJJ3_0),.dout(w_dff_B_zOyDH3mQ8_0),.clk(gclk));
	jdff dff_B_mldHocTn9_0(.din(w_dff_B_zOyDH3mQ8_0),.dout(w_dff_B_mldHocTn9_0),.clk(gclk));
	jdff dff_B_pHvw4bJ66_0(.din(w_dff_B_mldHocTn9_0),.dout(w_dff_B_pHvw4bJ66_0),.clk(gclk));
	jdff dff_B_QqSS2F190_0(.din(w_dff_B_pHvw4bJ66_0),.dout(w_dff_B_QqSS2F190_0),.clk(gclk));
	jdff dff_B_qLenSkaw9_0(.din(w_dff_B_QqSS2F190_0),.dout(w_dff_B_qLenSkaw9_0),.clk(gclk));
	jdff dff_B_0MzYLJRa4_0(.din(w_dff_B_qLenSkaw9_0),.dout(w_dff_B_0MzYLJRa4_0),.clk(gclk));
	jdff dff_A_SG3G3CBN4_1(.dout(w_G4092_6[1]),.din(w_dff_A_SG3G3CBN4_1),.clk(gclk));
	jdff dff_A_1qyT3Zbc1_1(.dout(w_dff_A_SG3G3CBN4_1),.din(w_dff_A_1qyT3Zbc1_1),.clk(gclk));
	jdff dff_A_HFuQmKcx2_2(.dout(w_G4092_6[2]),.din(w_dff_A_HFuQmKcx2_2),.clk(gclk));
	jdff dff_A_bqRP7G405_2(.dout(w_dff_A_HFuQmKcx2_2),.din(w_dff_A_bqRP7G405_2),.clk(gclk));
	jdff dff_B_teBg1fcI7_0(.din(n794),.dout(w_dff_B_teBg1fcI7_0),.clk(gclk));
	jdff dff_B_JsXWV9FB2_0(.din(n785),.dout(w_dff_B_JsXWV9FB2_0),.clk(gclk));
	jdff dff_A_h5ADyBn98_0(.dout(w_G54_0[0]),.din(w_dff_A_h5ADyBn98_0),.clk(gclk));
	jdff dff_A_bourfFbx5_0(.dout(w_dff_A_h5ADyBn98_0),.din(w_dff_A_bourfFbx5_0),.clk(gclk));
	jdff dff_A_sCcRFz7k0_0(.dout(w_dff_A_bourfFbx5_0),.din(w_dff_A_sCcRFz7k0_0),.clk(gclk));
	jdff dff_A_sJYbWsjZ4_0(.dout(w_dff_A_sCcRFz7k0_0),.din(w_dff_A_sJYbWsjZ4_0),.clk(gclk));
	jdff dff_A_SBP5Ix5F2_0(.dout(w_dff_A_sJYbWsjZ4_0),.din(w_dff_A_SBP5Ix5F2_0),.clk(gclk));
	jdff dff_A_BCdrsiL09_0(.dout(w_dff_A_SBP5Ix5F2_0),.din(w_dff_A_BCdrsiL09_0),.clk(gclk));
	jdff dff_A_mTjCCKB56_0(.dout(w_dff_A_BCdrsiL09_0),.din(w_dff_A_mTjCCKB56_0),.clk(gclk));
	jdff dff_A_yP8gDsbq5_0(.dout(w_dff_A_mTjCCKB56_0),.din(w_dff_A_yP8gDsbq5_0),.clk(gclk));
	jdff dff_A_TB7xn0HS8_0(.dout(w_dff_A_yP8gDsbq5_0),.din(w_dff_A_TB7xn0HS8_0),.clk(gclk));
	jdff dff_A_IaFBTQD19_1(.dout(w_G54_0[1]),.din(w_dff_A_IaFBTQD19_1),.clk(gclk));
	jdff dff_A_4JUUZQCO5_1(.dout(w_dff_A_IaFBTQD19_1),.din(w_dff_A_4JUUZQCO5_1),.clk(gclk));
	jdff dff_A_04xqFnmw4_1(.dout(w_dff_A_4JUUZQCO5_1),.din(w_dff_A_04xqFnmw4_1),.clk(gclk));
	jdff dff_A_Q3jqABZ76_1(.dout(w_dff_A_04xqFnmw4_1),.din(w_dff_A_Q3jqABZ76_1),.clk(gclk));
	jdff dff_A_Xjp4Fyrw4_0(.dout(w_n749_9[0]),.din(w_dff_A_Xjp4Fyrw4_0),.clk(gclk));
	jdff dff_A_Ia90jEnu5_2(.dout(w_n749_9[2]),.din(w_dff_A_Ia90jEnu5_2),.clk(gclk));
	jdff dff_A_rM0uCabR7_2(.dout(w_dff_A_Ia90jEnu5_2),.din(w_dff_A_rM0uCabR7_2),.clk(gclk));
	jdff dff_A_1CM9AJNo4_2(.dout(w_dff_A_rM0uCabR7_2),.din(w_dff_A_1CM9AJNo4_2),.clk(gclk));
	jdff dff_A_UBpo4WQX6_2(.dout(w_dff_A_1CM9AJNo4_2),.din(w_dff_A_UBpo4WQX6_2),.clk(gclk));
	jdff dff_A_hh5e29xM8_2(.dout(w_dff_A_UBpo4WQX6_2),.din(w_dff_A_hh5e29xM8_2),.clk(gclk));
	jdff dff_A_M33o1OnK1_2(.dout(w_dff_A_hh5e29xM8_2),.din(w_dff_A_M33o1OnK1_2),.clk(gclk));
	jdff dff_A_psOYotzO8_2(.dout(w_dff_A_M33o1OnK1_2),.din(w_dff_A_psOYotzO8_2),.clk(gclk));
	jdff dff_A_TL9SRI464_2(.dout(w_dff_A_psOYotzO8_2),.din(w_dff_A_TL9SRI464_2),.clk(gclk));
	jdff dff_A_GUynjsb18_2(.dout(w_dff_A_TL9SRI464_2),.din(w_dff_A_GUynjsb18_2),.clk(gclk));
	jdff dff_A_DBT6MTiZ9_2(.dout(w_dff_A_GUynjsb18_2),.din(w_dff_A_DBT6MTiZ9_2),.clk(gclk));
	jdff dff_A_M4lVm0cV4_2(.dout(w_dff_A_DBT6MTiZ9_2),.din(w_dff_A_M4lVm0cV4_2),.clk(gclk));
	jdff dff_A_dOIPu4iG2_2(.dout(w_dff_A_M4lVm0cV4_2),.din(w_dff_A_dOIPu4iG2_2),.clk(gclk));
	jdff dff_A_TKAGjbmO2_2(.dout(w_dff_A_dOIPu4iG2_2),.din(w_dff_A_TKAGjbmO2_2),.clk(gclk));
	jdff dff_A_4cKtydrZ2_2(.dout(w_dff_A_TKAGjbmO2_2),.din(w_dff_A_4cKtydrZ2_2),.clk(gclk));
	jdff dff_A_rIPRvKlC4_0(.dout(w_G123_0[0]),.din(w_dff_A_rIPRvKlC4_0),.clk(gclk));
	jdff dff_A_tVjet4u93_0(.dout(w_dff_A_rIPRvKlC4_0),.din(w_dff_A_tVjet4u93_0),.clk(gclk));
	jdff dff_A_OnstN0Yx8_0(.dout(w_G1691_2[0]),.din(w_dff_A_OnstN0Yx8_0),.clk(gclk));
	jdff dff_A_T3jpC6XO6_2(.dout(w_G1691_2[2]),.din(w_dff_A_T3jpC6XO6_2),.clk(gclk));
	jdff dff_A_DhcTfbY66_2(.dout(w_n1007_1[2]),.din(w_dff_A_DhcTfbY66_2),.clk(gclk));
	jdff dff_A_yRoGyYAK2_0(.dout(w_n1007_0[0]),.din(w_dff_A_yRoGyYAK2_0),.clk(gclk));
	jdff dff_A_sXry6PBj4_0(.dout(w_dff_A_yRoGyYAK2_0),.din(w_dff_A_sXry6PBj4_0),.clk(gclk));
	jdff dff_A_46GWPNeP7_0(.dout(w_dff_A_sXry6PBj4_0),.din(w_dff_A_46GWPNeP7_0),.clk(gclk));
	jdff dff_A_hKkU8OVO1_0(.dout(w_dff_A_46GWPNeP7_0),.din(w_dff_A_hKkU8OVO1_0),.clk(gclk));
	jdff dff_A_wf6cAqmr3_0(.dout(w_dff_A_hKkU8OVO1_0),.din(w_dff_A_wf6cAqmr3_0),.clk(gclk));
	jdff dff_A_8EA8ujsr5_0(.dout(w_dff_A_wf6cAqmr3_0),.din(w_dff_A_8EA8ujsr5_0),.clk(gclk));
	jdff dff_A_Tsv6D9am1_0(.dout(w_dff_A_8EA8ujsr5_0),.din(w_dff_A_Tsv6D9am1_0),.clk(gclk));
	jdff dff_A_klfcE5ZW5_0(.dout(w_dff_A_Tsv6D9am1_0),.din(w_dff_A_klfcE5ZW5_0),.clk(gclk));
	jdff dff_A_UbutgT4e4_0(.dout(w_dff_A_klfcE5ZW5_0),.din(w_dff_A_UbutgT4e4_0),.clk(gclk));
	jdff dff_A_XT0ifyt51_1(.dout(w_n1007_0[1]),.din(w_dff_A_XT0ifyt51_1),.clk(gclk));
	jdff dff_A_xDJ80oeC7_1(.dout(w_dff_A_XT0ifyt51_1),.din(w_dff_A_xDJ80oeC7_1),.clk(gclk));
	jdff dff_B_IyTF2DcU4_3(.din(n1007),.dout(w_dff_B_IyTF2DcU4_3),.clk(gclk));
	jdff dff_B_WHkje4zU7_3(.din(w_dff_B_IyTF2DcU4_3),.dout(w_dff_B_WHkje4zU7_3),.clk(gclk));
	jdff dff_B_vyq0mpfB3_3(.din(w_dff_B_WHkje4zU7_3),.dout(w_dff_B_vyq0mpfB3_3),.clk(gclk));
	jdff dff_B_N1nOxGne4_3(.din(w_dff_B_vyq0mpfB3_3),.dout(w_dff_B_N1nOxGne4_3),.clk(gclk));
	jdff dff_B_c1AparXY2_3(.din(w_dff_B_N1nOxGne4_3),.dout(w_dff_B_c1AparXY2_3),.clk(gclk));
	jdff dff_B_0dlJOkYq9_3(.din(w_dff_B_c1AparXY2_3),.dout(w_dff_B_0dlJOkYq9_3),.clk(gclk));
	jdff dff_B_rtLfTblU3_3(.din(w_dff_B_0dlJOkYq9_3),.dout(w_dff_B_rtLfTblU3_3),.clk(gclk));
	jdff dff_B_FJNAxe5d6_3(.din(w_dff_B_rtLfTblU3_3),.dout(w_dff_B_FJNAxe5d6_3),.clk(gclk));
	jdff dff_B_V0fEmAEL9_3(.din(w_dff_B_FJNAxe5d6_3),.dout(w_dff_B_V0fEmAEL9_3),.clk(gclk));
	jdff dff_B_eebWSicJ6_3(.din(w_dff_B_V0fEmAEL9_3),.dout(w_dff_B_eebWSicJ6_3),.clk(gclk));
	jdff dff_B_Oqq6t7dM4_3(.din(w_dff_B_eebWSicJ6_3),.dout(w_dff_B_Oqq6t7dM4_3),.clk(gclk));
	jdff dff_B_x6DPUGDY8_1(.din(n1230),.dout(w_dff_B_x6DPUGDY8_1),.clk(gclk));
	jdff dff_B_DZn4P6eY6_1(.din(w_dff_B_x6DPUGDY8_1),.dout(w_dff_B_DZn4P6eY6_1),.clk(gclk));
	jdff dff_B_JqBHtfFn8_1(.din(w_dff_B_DZn4P6eY6_1),.dout(w_dff_B_JqBHtfFn8_1),.clk(gclk));
	jdff dff_B_Y8deJoUJ1_1(.din(w_dff_B_JqBHtfFn8_1),.dout(w_dff_B_Y8deJoUJ1_1),.clk(gclk));
	jdff dff_B_T1WueL0q9_1(.din(w_dff_B_Y8deJoUJ1_1),.dout(w_dff_B_T1WueL0q9_1),.clk(gclk));
	jdff dff_B_fhEtG3S93_1(.din(w_dff_B_T1WueL0q9_1),.dout(w_dff_B_fhEtG3S93_1),.clk(gclk));
	jdff dff_B_sPtZDwYz6_1(.din(w_dff_B_fhEtG3S93_1),.dout(w_dff_B_sPtZDwYz6_1),.clk(gclk));
	jdff dff_B_vTuHdIBO3_1(.din(w_dff_B_sPtZDwYz6_1),.dout(w_dff_B_vTuHdIBO3_1),.clk(gclk));
	jdff dff_B_Y7hqqX3B0_1(.din(w_dff_B_vTuHdIBO3_1),.dout(w_dff_B_Y7hqqX3B0_1),.clk(gclk));
	jdff dff_B_nZyru5xd0_1(.din(w_dff_B_Y7hqqX3B0_1),.dout(w_dff_B_nZyru5xd0_1),.clk(gclk));
	jdff dff_B_uY9k2vfD6_1(.din(w_dff_B_nZyru5xd0_1),.dout(w_dff_B_uY9k2vfD6_1),.clk(gclk));
	jdff dff_B_mdCuGgsK5_1(.din(w_dff_B_uY9k2vfD6_1),.dout(w_dff_B_mdCuGgsK5_1),.clk(gclk));
	jdff dff_B_dGYrlCKi3_1(.din(w_dff_B_mdCuGgsK5_1),.dout(w_dff_B_dGYrlCKi3_1),.clk(gclk));
	jdff dff_B_6Wyove6d3_1(.din(w_dff_B_dGYrlCKi3_1),.dout(w_dff_B_6Wyove6d3_1),.clk(gclk));
	jdff dff_B_HiWT2w0S7_1(.din(w_dff_B_6Wyove6d3_1),.dout(w_dff_B_HiWT2w0S7_1),.clk(gclk));
	jdff dff_B_KjJlP0Ik6_1(.din(w_dff_B_HiWT2w0S7_1),.dout(w_dff_B_KjJlP0Ik6_1),.clk(gclk));
	jdff dff_B_xBbinTII5_1(.din(w_dff_B_KjJlP0Ik6_1),.dout(w_dff_B_xBbinTII5_1),.clk(gclk));
	jdff dff_B_U1VjBKb27_1(.din(n1232),.dout(w_dff_B_U1VjBKb27_1),.clk(gclk));
	jdff dff_B_WcuDG3Rh0_1(.din(w_dff_B_U1VjBKb27_1),.dout(w_dff_B_WcuDG3Rh0_1),.clk(gclk));
	jdff dff_B_MZHgArMs4_1(.din(w_dff_B_WcuDG3Rh0_1),.dout(w_dff_B_MZHgArMs4_1),.clk(gclk));
	jdff dff_B_PQVlnszt2_1(.din(w_dff_B_MZHgArMs4_1),.dout(w_dff_B_PQVlnszt2_1),.clk(gclk));
	jdff dff_B_RkINFyKm2_1(.din(w_dff_B_PQVlnszt2_1),.dout(w_dff_B_RkINFyKm2_1),.clk(gclk));
	jdff dff_B_QJgowWFx3_1(.din(w_dff_B_RkINFyKm2_1),.dout(w_dff_B_QJgowWFx3_1),.clk(gclk));
	jdff dff_B_pW2uDacm8_1(.din(w_dff_B_QJgowWFx3_1),.dout(w_dff_B_pW2uDacm8_1),.clk(gclk));
	jdff dff_B_aanXl7Ko2_1(.din(w_dff_B_pW2uDacm8_1),.dout(w_dff_B_aanXl7Ko2_1),.clk(gclk));
	jdff dff_B_AbRIiNki4_1(.din(w_dff_B_aanXl7Ko2_1),.dout(w_dff_B_AbRIiNki4_1),.clk(gclk));
	jdff dff_B_2xpmdX743_1(.din(w_dff_B_AbRIiNki4_1),.dout(w_dff_B_2xpmdX743_1),.clk(gclk));
	jdff dff_B_ME5vetwx8_1(.din(w_dff_B_2xpmdX743_1),.dout(w_dff_B_ME5vetwx8_1),.clk(gclk));
	jdff dff_B_GtU33t4T5_1(.din(w_dff_B_ME5vetwx8_1),.dout(w_dff_B_GtU33t4T5_1),.clk(gclk));
	jdff dff_B_xrdT1GMN5_1(.din(n937),.dout(w_dff_B_xrdT1GMN5_1),.clk(gclk));
	jdff dff_B_zXT6ynzD3_1(.din(w_dff_B_xrdT1GMN5_1),.dout(w_dff_B_zXT6ynzD3_1),.clk(gclk));
	jdff dff_B_0HBF12dA9_1(.din(w_dff_B_zXT6ynzD3_1),.dout(w_dff_B_0HBF12dA9_1),.clk(gclk));
	jdff dff_B_M8VSGcPA7_1(.din(w_dff_B_0HBF12dA9_1),.dout(w_dff_B_M8VSGcPA7_1),.clk(gclk));
	jdff dff_B_Xfnlr1HJ1_1(.din(w_dff_B_M8VSGcPA7_1),.dout(w_dff_B_Xfnlr1HJ1_1),.clk(gclk));
	jdff dff_B_3WgbZ8Dl5_1(.din(w_dff_B_Xfnlr1HJ1_1),.dout(w_dff_B_3WgbZ8Dl5_1),.clk(gclk));
	jdff dff_B_m9iJzj4t6_1(.din(w_dff_B_3WgbZ8Dl5_1),.dout(w_dff_B_m9iJzj4t6_1),.clk(gclk));
	jdff dff_B_WIqywlki5_1(.din(w_dff_B_m9iJzj4t6_1),.dout(w_dff_B_WIqywlki5_1),.clk(gclk));
	jdff dff_B_VxkkGQO10_1(.din(w_dff_B_WIqywlki5_1),.dout(w_dff_B_VxkkGQO10_1),.clk(gclk));
	jdff dff_B_PvmQsIGm0_1(.din(w_dff_B_VxkkGQO10_1),.dout(w_dff_B_PvmQsIGm0_1),.clk(gclk));
	jdff dff_B_Gyu7mPT03_1(.din(w_dff_B_PvmQsIGm0_1),.dout(w_dff_B_Gyu7mPT03_1),.clk(gclk));
	jdff dff_B_zzQxdAZy6_0(.din(n869),.dout(w_dff_B_zzQxdAZy6_0),.clk(gclk));
	jdff dff_B_IKO5kJGV8_1(.din(n866),.dout(w_dff_B_IKO5kJGV8_1),.clk(gclk));
	jdff dff_B_Hm0NnoUi5_1(.din(w_dff_B_IKO5kJGV8_1),.dout(w_dff_B_Hm0NnoUi5_1),.clk(gclk));
	jdff dff_A_Mo9sV4jz4_1(.dout(w_G4_0[1]),.din(w_dff_A_Mo9sV4jz4_1),.clk(gclk));
	jdff dff_B_naccYboo1_3(.din(G4),.dout(w_dff_B_naccYboo1_3),.clk(gclk));
	jdff dff_B_8MPEj8T95_3(.din(w_dff_B_naccYboo1_3),.dout(w_dff_B_8MPEj8T95_3),.clk(gclk));
	jdff dff_B_LILldglh2_3(.din(w_dff_B_8MPEj8T95_3),.dout(w_dff_B_LILldglh2_3),.clk(gclk));
	jdff dff_B_aOff08097_3(.din(w_dff_B_LILldglh2_3),.dout(w_dff_B_aOff08097_3),.clk(gclk));
	jdff dff_B_UYB3ZrXN6_3(.din(w_dff_B_aOff08097_3),.dout(w_dff_B_UYB3ZrXN6_3),.clk(gclk));
	jdff dff_A_9yjaLKeD7_0(.dout(w_n1201_0[0]),.din(w_dff_A_9yjaLKeD7_0),.clk(gclk));
	jdff dff_A_IBBWSIUp1_1(.dout(w_n1201_0[1]),.din(w_dff_A_IBBWSIUp1_1),.clk(gclk));
	jdff dff_A_t9wquEM91_1(.dout(w_dff_A_IBBWSIUp1_1),.din(w_dff_A_t9wquEM91_1),.clk(gclk));
	jdff dff_B_PqvOZdZ71_3(.din(n1201),.dout(w_dff_B_PqvOZdZ71_3),.clk(gclk));
	jdff dff_B_efUeAKq74_3(.din(w_dff_B_PqvOZdZ71_3),.dout(w_dff_B_efUeAKq74_3),.clk(gclk));
	jdff dff_B_kFqFvyp07_3(.din(w_dff_B_efUeAKq74_3),.dout(w_dff_B_kFqFvyp07_3),.clk(gclk));
	jdff dff_B_se4LDacT7_3(.din(w_dff_B_kFqFvyp07_3),.dout(w_dff_B_se4LDacT7_3),.clk(gclk));
	jdff dff_B_zzah0dQD8_3(.din(w_dff_B_se4LDacT7_3),.dout(w_dff_B_zzah0dQD8_3),.clk(gclk));
	jdff dff_B_B5S7AWBv8_3(.din(w_dff_B_zzah0dQD8_3),.dout(w_dff_B_B5S7AWBv8_3),.clk(gclk));
	jdff dff_B_gpdwNBUO6_3(.din(w_dff_B_B5S7AWBv8_3),.dout(w_dff_B_gpdwNBUO6_3),.clk(gclk));
	jdff dff_B_JjLzSQoQ5_3(.din(w_dff_B_gpdwNBUO6_3),.dout(w_dff_B_JjLzSQoQ5_3),.clk(gclk));
	jdff dff_B_dCJ9NGDw9_3(.din(w_dff_B_JjLzSQoQ5_3),.dout(w_dff_B_dCJ9NGDw9_3),.clk(gclk));
	jdff dff_B_kIrk9FHa7_3(.din(w_dff_B_dCJ9NGDw9_3),.dout(w_dff_B_kIrk9FHa7_3),.clk(gclk));
	jdff dff_B_xpHjaMtT7_3(.din(w_dff_B_kIrk9FHa7_3),.dout(w_dff_B_xpHjaMtT7_3),.clk(gclk));
	jdff dff_B_LeEQJQeX5_3(.din(w_dff_B_xpHjaMtT7_3),.dout(w_dff_B_LeEQJQeX5_3),.clk(gclk));
	jdff dff_B_o7daRyHo8_3(.din(w_dff_B_LeEQJQeX5_3),.dout(w_dff_B_o7daRyHo8_3),.clk(gclk));
	jdff dff_B_20QxDwqu1_3(.din(w_dff_B_o7daRyHo8_3),.dout(w_dff_B_20QxDwqu1_3),.clk(gclk));
	jdff dff_B_6JI8y1nQ3_3(.din(w_dff_B_20QxDwqu1_3),.dout(w_dff_B_6JI8y1nQ3_3),.clk(gclk));
	jdff dff_A_0LASztWG5_0(.dout(w_G4092_5[0]),.din(w_dff_A_0LASztWG5_0),.clk(gclk));
	jdff dff_A_Mli2ce8Q1_0(.dout(w_dff_A_0LASztWG5_0),.din(w_dff_A_Mli2ce8Q1_0),.clk(gclk));
	jdff dff_A_VRkDdy4a7_0(.dout(w_dff_A_Mli2ce8Q1_0),.din(w_dff_A_VRkDdy4a7_0),.clk(gclk));
	jdff dff_A_ZM5H8oma0_0(.dout(w_dff_A_VRkDdy4a7_0),.din(w_dff_A_ZM5H8oma0_0),.clk(gclk));
	jdff dff_A_TNMG6spc9_0(.dout(w_dff_A_ZM5H8oma0_0),.din(w_dff_A_TNMG6spc9_0),.clk(gclk));
	jdff dff_A_AOhrr9dn7_0(.dout(w_dff_A_TNMG6spc9_0),.din(w_dff_A_AOhrr9dn7_0),.clk(gclk));
	jdff dff_A_5zR3yP6r9_1(.dout(w_G4092_5[1]),.din(w_dff_A_5zR3yP6r9_1),.clk(gclk));
	jdff dff_A_9HxEik9S3_1(.dout(w_dff_A_5zR3yP6r9_1),.din(w_dff_A_9HxEik9S3_1),.clk(gclk));
	jdff dff_A_uRsiHsta8_1(.dout(w_dff_A_9HxEik9S3_1),.din(w_dff_A_uRsiHsta8_1),.clk(gclk));
	jdff dff_A_OJRTFFqW7_1(.dout(w_dff_A_uRsiHsta8_1),.din(w_dff_A_OJRTFFqW7_1),.clk(gclk));
	jdff dff_A_2CQVESU27_1(.dout(w_dff_A_OJRTFFqW7_1),.din(w_dff_A_2CQVESU27_1),.clk(gclk));
	jdff dff_A_lB8jkucz9_1(.dout(w_dff_A_2CQVESU27_1),.din(w_dff_A_lB8jkucz9_1),.clk(gclk));
	jdff dff_A_CclZyRgt7_0(.dout(w_n749_7[0]),.din(w_dff_A_CclZyRgt7_0),.clk(gclk));
	jdff dff_A_sHnMweYL9_0(.dout(w_dff_A_CclZyRgt7_0),.din(w_dff_A_sHnMweYL9_0),.clk(gclk));
	jdff dff_A_RzxkQFGd9_0(.dout(w_dff_A_sHnMweYL9_0),.din(w_dff_A_RzxkQFGd9_0),.clk(gclk));
	jdff dff_A_VuzFRFpJ3_0(.dout(w_dff_A_RzxkQFGd9_0),.din(w_dff_A_VuzFRFpJ3_0),.clk(gclk));
	jdff dff_A_oHcayFwH2_0(.dout(w_dff_A_VuzFRFpJ3_0),.din(w_dff_A_oHcayFwH2_0),.clk(gclk));
	jdff dff_A_wbv0D6hL1_0(.dout(w_dff_A_oHcayFwH2_0),.din(w_dff_A_wbv0D6hL1_0),.clk(gclk));
	jdff dff_A_jqeDkZhf1_0(.dout(w_dff_A_wbv0D6hL1_0),.din(w_dff_A_jqeDkZhf1_0),.clk(gclk));
	jdff dff_A_VeGW5vE50_0(.dout(w_dff_A_jqeDkZhf1_0),.din(w_dff_A_VeGW5vE50_0),.clk(gclk));
	jdff dff_A_WzB4BH967_0(.dout(w_dff_A_VeGW5vE50_0),.din(w_dff_A_WzB4BH967_0),.clk(gclk));
	jdff dff_A_HOVFvIwm8_0(.dout(w_dff_A_WzB4BH967_0),.din(w_dff_A_HOVFvIwm8_0),.clk(gclk));
	jdff dff_A_JO9RWGma1_0(.dout(w_dff_A_HOVFvIwm8_0),.din(w_dff_A_JO9RWGma1_0),.clk(gclk));
	jdff dff_A_7x2yeONB8_0(.dout(w_dff_A_JO9RWGma1_0),.din(w_dff_A_7x2yeONB8_0),.clk(gclk));
	jdff dff_A_Etcec46M3_0(.dout(w_n749_2[0]),.din(w_dff_A_Etcec46M3_0),.clk(gclk));
	jdff dff_A_fScvVv0S0_0(.dout(w_dff_A_Etcec46M3_0),.din(w_dff_A_fScvVv0S0_0),.clk(gclk));
	jdff dff_A_poGi5q4w6_1(.dout(w_n749_2[1]),.din(w_dff_A_poGi5q4w6_1),.clk(gclk));
	jdff dff_A_NtPI2eCN5_1(.dout(w_dff_A_poGi5q4w6_1),.din(w_dff_A_NtPI2eCN5_1),.clk(gclk));
	jdff dff_B_6wMq7sdz6_1(.din(G115),.dout(w_dff_B_6wMq7sdz6_1),.clk(gclk));
	jdff dff_B_OUybV2HC1_1(.din(w_dff_B_6wMq7sdz6_1),.dout(w_dff_B_OUybV2HC1_1),.clk(gclk));
	jdff dff_B_Dpc3eSHg5_0(.din(n1505),.dout(w_dff_B_Dpc3eSHg5_0),.clk(gclk));
	jdff dff_B_33XXtlKC0_0(.din(w_dff_B_Dpc3eSHg5_0),.dout(w_dff_B_33XXtlKC0_0),.clk(gclk));
	jdff dff_B_xPQrDetT7_0(.din(w_dff_B_33XXtlKC0_0),.dout(w_dff_B_xPQrDetT7_0),.clk(gclk));
	jdff dff_B_VjUnHcXl1_0(.din(w_dff_B_xPQrDetT7_0),.dout(w_dff_B_VjUnHcXl1_0),.clk(gclk));
	jdff dff_B_NyYosQTj0_0(.din(w_dff_B_VjUnHcXl1_0),.dout(w_dff_B_NyYosQTj0_0),.clk(gclk));
	jdff dff_B_6GiQMakZ3_0(.din(w_dff_B_NyYosQTj0_0),.dout(w_dff_B_6GiQMakZ3_0),.clk(gclk));
	jdff dff_B_xDIgkjsQ7_0(.din(w_dff_B_6GiQMakZ3_0),.dout(w_dff_B_xDIgkjsQ7_0),.clk(gclk));
	jdff dff_B_Vn6DWYu36_0(.din(w_dff_B_xDIgkjsQ7_0),.dout(w_dff_B_Vn6DWYu36_0),.clk(gclk));
	jdff dff_B_Xy6Pan1d4_0(.din(w_dff_B_Vn6DWYu36_0),.dout(w_dff_B_Xy6Pan1d4_0),.clk(gclk));
	jdff dff_B_E3XKDFEP0_0(.din(w_dff_B_Xy6Pan1d4_0),.dout(w_dff_B_E3XKDFEP0_0),.clk(gclk));
	jdff dff_B_RGuPtAUl9_0(.din(w_dff_B_E3XKDFEP0_0),.dout(w_dff_B_RGuPtAUl9_0),.clk(gclk));
	jdff dff_B_HsBGya5a5_0(.din(w_dff_B_RGuPtAUl9_0),.dout(w_dff_B_HsBGya5a5_0),.clk(gclk));
	jdff dff_B_FFNl50ZA3_0(.din(w_dff_B_HsBGya5a5_0),.dout(w_dff_B_FFNl50ZA3_0),.clk(gclk));
	jdff dff_B_LfUUAna41_0(.din(w_dff_B_FFNl50ZA3_0),.dout(w_dff_B_LfUUAna41_0),.clk(gclk));
	jdff dff_B_9jbclwIf6_0(.din(w_dff_B_LfUUAna41_0),.dout(w_dff_B_9jbclwIf6_0),.clk(gclk));
	jdff dff_B_54sFbtbX3_0(.din(w_dff_B_9jbclwIf6_0),.dout(w_dff_B_54sFbtbX3_0),.clk(gclk));
	jdff dff_B_bBgJxmY12_0(.din(w_dff_B_54sFbtbX3_0),.dout(w_dff_B_bBgJxmY12_0),.clk(gclk));
	jdff dff_B_LssX4v2H2_1(.din(G120),.dout(w_dff_B_LssX4v2H2_1),.clk(gclk));
	jdff dff_B_aybXx0cm8_1(.din(w_dff_B_LssX4v2H2_1),.dout(w_dff_B_aybXx0cm8_1),.clk(gclk));
	jdff dff_B_yIyzP5Yo3_1(.din(w_dff_B_aybXx0cm8_1),.dout(w_dff_B_yIyzP5Yo3_1),.clk(gclk));
	jdff dff_B_AQMrhbqO2_0(.din(n1666),.dout(w_dff_B_AQMrhbqO2_0),.clk(gclk));
	jdff dff_B_639ljYov0_0(.din(w_dff_B_AQMrhbqO2_0),.dout(w_dff_B_639ljYov0_0),.clk(gclk));
	jdff dff_B_HlDp2aqp3_0(.din(w_dff_B_639ljYov0_0),.dout(w_dff_B_HlDp2aqp3_0),.clk(gclk));
	jdff dff_B_6RcG2bXo2_0(.din(w_dff_B_HlDp2aqp3_0),.dout(w_dff_B_6RcG2bXo2_0),.clk(gclk));
	jdff dff_B_i48s8PXH0_0(.din(w_dff_B_6RcG2bXo2_0),.dout(w_dff_B_i48s8PXH0_0),.clk(gclk));
	jdff dff_B_nx1Xqc5Y0_0(.din(w_dff_B_i48s8PXH0_0),.dout(w_dff_B_nx1Xqc5Y0_0),.clk(gclk));
	jdff dff_B_SDKdmsel8_0(.din(w_dff_B_nx1Xqc5Y0_0),.dout(w_dff_B_SDKdmsel8_0),.clk(gclk));
	jdff dff_B_QWJZBtDZ5_0(.din(w_dff_B_SDKdmsel8_0),.dout(w_dff_B_QWJZBtDZ5_0),.clk(gclk));
	jdff dff_B_RX0gvrzg4_0(.din(w_dff_B_QWJZBtDZ5_0),.dout(w_dff_B_RX0gvrzg4_0),.clk(gclk));
	jdff dff_B_YPJ1XIzA3_0(.din(w_dff_B_RX0gvrzg4_0),.dout(w_dff_B_YPJ1XIzA3_0),.clk(gclk));
	jdff dff_B_e0xHLQmV3_0(.din(w_dff_B_YPJ1XIzA3_0),.dout(w_dff_B_e0xHLQmV3_0),.clk(gclk));
	jdff dff_B_4lCDyEm47_0(.din(w_dff_B_e0xHLQmV3_0),.dout(w_dff_B_4lCDyEm47_0),.clk(gclk));
	jdff dff_B_3JJNPPks3_0(.din(w_dff_B_4lCDyEm47_0),.dout(w_dff_B_3JJNPPks3_0),.clk(gclk));
	jdff dff_B_SNRbhPRA2_0(.din(w_dff_B_3JJNPPks3_0),.dout(w_dff_B_SNRbhPRA2_0),.clk(gclk));
	jdff dff_B_56tIiNrx0_0(.din(w_dff_B_SNRbhPRA2_0),.dout(w_dff_B_56tIiNrx0_0),.clk(gclk));
	jdff dff_B_UF81N8mv8_0(.din(w_dff_B_56tIiNrx0_0),.dout(w_dff_B_UF81N8mv8_0),.clk(gclk));
	jdff dff_B_ivEnXF2Z0_0(.din(w_dff_B_UF81N8mv8_0),.dout(w_dff_B_ivEnXF2Z0_0),.clk(gclk));
	jdff dff_B_R8WvSjL46_1(.din(G118),.dout(w_dff_B_R8WvSjL46_1),.clk(gclk));
	jdff dff_B_0jJGfgzu4_1(.din(w_dff_B_R8WvSjL46_1),.dout(w_dff_B_0jJGfgzu4_1),.clk(gclk));
	jdff dff_B_kALI9UUy4_1(.din(w_dff_B_0jJGfgzu4_1),.dout(w_dff_B_kALI9UUy4_1),.clk(gclk));
	jdff dff_A_s6k4vIgb7_0(.dout(w_G4092_9[0]),.din(w_dff_A_s6k4vIgb7_0),.clk(gclk));
	jdff dff_A_TGt0vwSs9_0(.dout(w_dff_A_s6k4vIgb7_0),.din(w_dff_A_TGt0vwSs9_0),.clk(gclk));
	jdff dff_A_X5Ahz7o40_0(.dout(w_dff_A_TGt0vwSs9_0),.din(w_dff_A_X5Ahz7o40_0),.clk(gclk));
	jdff dff_A_tot8P65E9_0(.dout(w_dff_A_X5Ahz7o40_0),.din(w_dff_A_tot8P65E9_0),.clk(gclk));
	jdff dff_A_OQJ74M3V3_0(.dout(w_dff_A_tot8P65E9_0),.din(w_dff_A_OQJ74M3V3_0),.clk(gclk));
	jdff dff_A_4XETqUAy6_1(.dout(w_G4092_9[1]),.din(w_dff_A_4XETqUAy6_1),.clk(gclk));
	jdff dff_A_t69nBHlN1_1(.dout(w_dff_A_4XETqUAy6_1),.din(w_dff_A_t69nBHlN1_1),.clk(gclk));
	jdff dff_A_de7GXQsn2_1(.dout(w_dff_A_t69nBHlN1_1),.din(w_dff_A_de7GXQsn2_1),.clk(gclk));
	jdff dff_A_Nuq3dACF0_1(.dout(w_dff_A_de7GXQsn2_1),.din(w_dff_A_Nuq3dACF0_1),.clk(gclk));
	jdff dff_A_diLxcyc94_0(.dout(w_G4092_2[0]),.din(w_dff_A_diLxcyc94_0),.clk(gclk));
	jdff dff_A_FdR8LCEy3_0(.dout(w_dff_A_diLxcyc94_0),.din(w_dff_A_FdR8LCEy3_0),.clk(gclk));
	jdff dff_A_Y34mV9nf4_0(.dout(w_dff_A_FdR8LCEy3_0),.din(w_dff_A_Y34mV9nf4_0),.clk(gclk));
	jdff dff_A_IzyPLtpV7_0(.dout(w_dff_A_Y34mV9nf4_0),.din(w_dff_A_IzyPLtpV7_0),.clk(gclk));
	jdff dff_A_UQCIH12x2_0(.dout(w_dff_A_IzyPLtpV7_0),.din(w_dff_A_UQCIH12x2_0),.clk(gclk));
	jdff dff_A_4nQMsEJZ0_1(.dout(w_G4092_2[1]),.din(w_dff_A_4nQMsEJZ0_1),.clk(gclk));
	jdff dff_A_sEYg9hlu1_1(.dout(w_dff_A_4nQMsEJZ0_1),.din(w_dff_A_sEYg9hlu1_1),.clk(gclk));
	jdff dff_A_mSesgIDu5_1(.dout(w_dff_A_sEYg9hlu1_1),.din(w_dff_A_mSesgIDu5_1),.clk(gclk));
	jdff dff_A_tnyGzhZ58_1(.dout(w_dff_A_mSesgIDu5_1),.din(w_dff_A_tnyGzhZ58_1),.clk(gclk));
	jdff dff_A_qyUmYJxd1_0(.dout(w_n749_13[0]),.din(w_dff_A_qyUmYJxd1_0),.clk(gclk));
	jdff dff_A_e5nWRFdM4_0(.dout(w_dff_A_qyUmYJxd1_0),.din(w_dff_A_e5nWRFdM4_0),.clk(gclk));
	jdff dff_A_xnnPnaiM2_0(.dout(w_dff_A_e5nWRFdM4_0),.din(w_dff_A_xnnPnaiM2_0),.clk(gclk));
	jdff dff_B_KpTvdyl23_1(.din(n1671),.dout(w_dff_B_KpTvdyl23_1),.clk(gclk));
	jdff dff_B_afC9Rhzc5_1(.din(w_dff_B_KpTvdyl23_1),.dout(w_dff_B_afC9Rhzc5_1),.clk(gclk));
	jdff dff_B_1ovAACwt8_1(.din(w_dff_B_afC9Rhzc5_1),.dout(w_dff_B_1ovAACwt8_1),.clk(gclk));
	jdff dff_B_956HnWuz3_1(.din(w_dff_B_1ovAACwt8_1),.dout(w_dff_B_956HnWuz3_1),.clk(gclk));
	jdff dff_B_xc1ZUklw0_1(.din(w_dff_B_956HnWuz3_1),.dout(w_dff_B_xc1ZUklw0_1),.clk(gclk));
	jdff dff_B_kpz4Wosn0_1(.din(w_dff_B_xc1ZUklw0_1),.dout(w_dff_B_kpz4Wosn0_1),.clk(gclk));
	jdff dff_B_8nsS6u1d7_1(.din(w_dff_B_kpz4Wosn0_1),.dout(w_dff_B_8nsS6u1d7_1),.clk(gclk));
	jdff dff_B_5uEH2ZZq8_1(.din(w_dff_B_8nsS6u1d7_1),.dout(w_dff_B_5uEH2ZZq8_1),.clk(gclk));
	jdff dff_B_S2ZwWOyy1_1(.din(w_dff_B_5uEH2ZZq8_1),.dout(w_dff_B_S2ZwWOyy1_1),.clk(gclk));
	jdff dff_B_dH5pHsAD8_1(.din(w_dff_B_S2ZwWOyy1_1),.dout(w_dff_B_dH5pHsAD8_1),.clk(gclk));
	jdff dff_B_1D23wk9X7_1(.din(w_dff_B_dH5pHsAD8_1),.dout(w_dff_B_1D23wk9X7_1),.clk(gclk));
	jdff dff_B_2qVySc086_1(.din(w_dff_B_1D23wk9X7_1),.dout(w_dff_B_2qVySc086_1),.clk(gclk));
	jdff dff_B_FN6Y1TDz0_1(.din(w_dff_B_2qVySc086_1),.dout(w_dff_B_FN6Y1TDz0_1),.clk(gclk));
	jdff dff_B_9Z9xNBnA7_1(.din(w_dff_B_FN6Y1TDz0_1),.dout(w_dff_B_9Z9xNBnA7_1),.clk(gclk));
	jdff dff_B_JYRFyvTf1_1(.din(w_dff_B_9Z9xNBnA7_1),.dout(w_dff_B_JYRFyvTf1_1),.clk(gclk));
	jdff dff_B_2u7nNcwk6_1(.din(w_dff_B_JYRFyvTf1_1),.dout(w_dff_B_2u7nNcwk6_1),.clk(gclk));
	jdff dff_B_Hdw1ig2D4_1(.din(w_dff_B_2u7nNcwk6_1),.dout(w_dff_B_Hdw1ig2D4_1),.clk(gclk));
	jdff dff_B_k6vZVOWm4_1(.din(w_dff_B_Hdw1ig2D4_1),.dout(w_dff_B_k6vZVOWm4_1),.clk(gclk));
	jdff dff_B_EzSnGYyx7_1(.din(w_dff_B_k6vZVOWm4_1),.dout(w_dff_B_EzSnGYyx7_1),.clk(gclk));
	jdff dff_B_Y3yrwssN7_1(.din(w_dff_B_EzSnGYyx7_1),.dout(w_dff_B_Y3yrwssN7_1),.clk(gclk));
	jdff dff_B_df65VDdF6_1(.din(w_dff_B_Y3yrwssN7_1),.dout(w_dff_B_df65VDdF6_1),.clk(gclk));
	jdff dff_B_Dzxeri387_1(.din(w_dff_B_df65VDdF6_1),.dout(w_dff_B_Dzxeri387_1),.clk(gclk));
	jdff dff_B_z0n0vzl45_1(.din(n1676),.dout(w_dff_B_z0n0vzl45_1),.clk(gclk));
	jdff dff_A_BIiek8Bj7_1(.dout(w_n800_1[1]),.din(w_dff_A_BIiek8Bj7_1),.clk(gclk));
	jdff dff_A_RptDZlU53_1(.dout(w_dff_A_BIiek8Bj7_1),.din(w_dff_A_RptDZlU53_1),.clk(gclk));
	jdff dff_A_NcSppiiC5_1(.dout(w_dff_A_RptDZlU53_1),.din(w_dff_A_NcSppiiC5_1),.clk(gclk));
	jdff dff_A_uOwvCTMW1_1(.dout(w_dff_A_NcSppiiC5_1),.din(w_dff_A_uOwvCTMW1_1),.clk(gclk));
	jdff dff_A_ILyyk1Ts0_1(.dout(w_dff_A_uOwvCTMW1_1),.din(w_dff_A_ILyyk1Ts0_1),.clk(gclk));
	jdff dff_A_8sxACelC8_1(.dout(w_dff_A_ILyyk1Ts0_1),.din(w_dff_A_8sxACelC8_1),.clk(gclk));
	jdff dff_A_rII7vRHv4_1(.dout(w_dff_A_8sxACelC8_1),.din(w_dff_A_rII7vRHv4_1),.clk(gclk));
	jdff dff_A_6TnomH5k7_1(.dout(w_dff_A_rII7vRHv4_1),.din(w_dff_A_6TnomH5k7_1),.clk(gclk));
	jdff dff_A_iF88Yg0d9_1(.dout(w_dff_A_6TnomH5k7_1),.din(w_dff_A_iF88Yg0d9_1),.clk(gclk));
	jdff dff_A_bKu8rEoc6_1(.dout(w_dff_A_iF88Yg0d9_1),.din(w_dff_A_bKu8rEoc6_1),.clk(gclk));
	jdff dff_A_K30UDXMw2_1(.dout(w_dff_A_bKu8rEoc6_1),.din(w_dff_A_K30UDXMw2_1),.clk(gclk));
	jdff dff_A_QPyYg0kv1_1(.dout(w_dff_A_K30UDXMw2_1),.din(w_dff_A_QPyYg0kv1_1),.clk(gclk));
	jdff dff_A_v386zVsG1_1(.dout(w_dff_A_QPyYg0kv1_1),.din(w_dff_A_v386zVsG1_1),.clk(gclk));
	jdff dff_A_twRL69CU3_1(.dout(w_dff_A_v386zVsG1_1),.din(w_dff_A_twRL69CU3_1),.clk(gclk));
	jdff dff_A_8NNw33gg1_2(.dout(w_n800_1[2]),.din(w_dff_A_8NNw33gg1_2),.clk(gclk));
	jdff dff_A_0sGD3zE15_2(.dout(w_dff_A_8NNw33gg1_2),.din(w_dff_A_0sGD3zE15_2),.clk(gclk));
	jdff dff_A_cLpzrqEb4_2(.dout(w_dff_A_0sGD3zE15_2),.din(w_dff_A_cLpzrqEb4_2),.clk(gclk));
	jdff dff_A_mpZKO8EQ1_2(.dout(w_dff_A_cLpzrqEb4_2),.din(w_dff_A_mpZKO8EQ1_2),.clk(gclk));
	jdff dff_A_CAhSMrq20_2(.dout(w_dff_A_mpZKO8EQ1_2),.din(w_dff_A_CAhSMrq20_2),.clk(gclk));
	jdff dff_A_DI3kWwgr6_2(.dout(w_dff_A_CAhSMrq20_2),.din(w_dff_A_DI3kWwgr6_2),.clk(gclk));
	jdff dff_A_uxVazMlK0_2(.dout(w_dff_A_DI3kWwgr6_2),.din(w_dff_A_uxVazMlK0_2),.clk(gclk));
	jdff dff_A_L7vU8Fzk1_2(.dout(w_dff_A_uxVazMlK0_2),.din(w_dff_A_L7vU8Fzk1_2),.clk(gclk));
	jdff dff_A_pdF860xr3_2(.dout(w_dff_A_L7vU8Fzk1_2),.din(w_dff_A_pdF860xr3_2),.clk(gclk));
	jdff dff_A_llbMoU9z6_2(.dout(w_dff_A_pdF860xr3_2),.din(w_dff_A_llbMoU9z6_2),.clk(gclk));
	jdff dff_A_V54IQlgl9_1(.dout(w_n800_0[1]),.din(w_dff_A_V54IQlgl9_1),.clk(gclk));
	jdff dff_A_9fu9BnWB3_1(.dout(w_dff_A_V54IQlgl9_1),.din(w_dff_A_9fu9BnWB3_1),.clk(gclk));
	jdff dff_A_u89riaRk0_1(.dout(w_dff_A_9fu9BnWB3_1),.din(w_dff_A_u89riaRk0_1),.clk(gclk));
	jdff dff_A_QZvFthX22_1(.dout(w_dff_A_u89riaRk0_1),.din(w_dff_A_QZvFthX22_1),.clk(gclk));
	jdff dff_A_GJWRm6WC3_1(.dout(w_dff_A_QZvFthX22_1),.din(w_dff_A_GJWRm6WC3_1),.clk(gclk));
	jdff dff_A_HRt0K5jK9_1(.dout(w_dff_A_GJWRm6WC3_1),.din(w_dff_A_HRt0K5jK9_1),.clk(gclk));
	jdff dff_A_mAJinRlJ0_1(.dout(w_dff_A_HRt0K5jK9_1),.din(w_dff_A_mAJinRlJ0_1),.clk(gclk));
	jdff dff_A_AVlTkWD56_1(.dout(w_dff_A_mAJinRlJ0_1),.din(w_dff_A_AVlTkWD56_1),.clk(gclk));
	jdff dff_A_Q0LnOjhy7_1(.dout(w_dff_A_AVlTkWD56_1),.din(w_dff_A_Q0LnOjhy7_1),.clk(gclk));
	jdff dff_A_h6pbmVRJ9_1(.dout(w_dff_A_Q0LnOjhy7_1),.din(w_dff_A_h6pbmVRJ9_1),.clk(gclk));
	jdff dff_A_a9eq3c733_1(.dout(w_dff_A_h6pbmVRJ9_1),.din(w_dff_A_a9eq3c733_1),.clk(gclk));
	jdff dff_A_lIbZN6lz7_2(.dout(w_n800_0[2]),.din(w_dff_A_lIbZN6lz7_2),.clk(gclk));
	jdff dff_A_9QX48GXi0_2(.dout(w_dff_A_lIbZN6lz7_2),.din(w_dff_A_9QX48GXi0_2),.clk(gclk));
	jdff dff_A_Zdz5MnjK3_2(.dout(w_dff_A_9QX48GXi0_2),.din(w_dff_A_Zdz5MnjK3_2),.clk(gclk));
	jdff dff_A_aolLGTMm4_2(.dout(w_dff_A_Zdz5MnjK3_2),.din(w_dff_A_aolLGTMm4_2),.clk(gclk));
	jdff dff_B_d9uxW4Ca2_3(.din(n800),.dout(w_dff_B_d9uxW4Ca2_3),.clk(gclk));
	jdff dff_B_aYP5Hrdf1_3(.din(w_dff_B_d9uxW4Ca2_3),.dout(w_dff_B_aYP5Hrdf1_3),.clk(gclk));
	jdff dff_B_ie2B6lhi7_3(.din(w_dff_B_aYP5Hrdf1_3),.dout(w_dff_B_ie2B6lhi7_3),.clk(gclk));
	jdff dff_B_7oGvw9J40_3(.din(w_dff_B_ie2B6lhi7_3),.dout(w_dff_B_7oGvw9J40_3),.clk(gclk));
	jdff dff_B_TRdCt46c9_3(.din(w_dff_B_7oGvw9J40_3),.dout(w_dff_B_TRdCt46c9_3),.clk(gclk));
	jdff dff_B_867Gc1Oh4_3(.din(w_dff_B_TRdCt46c9_3),.dout(w_dff_B_867Gc1Oh4_3),.clk(gclk));
	jdff dff_B_GptRj8EL6_3(.din(w_dff_B_867Gc1Oh4_3),.dout(w_dff_B_GptRj8EL6_3),.clk(gclk));
	jdff dff_B_YkdDG63U7_3(.din(w_dff_B_GptRj8EL6_3),.dout(w_dff_B_YkdDG63U7_3),.clk(gclk));
	jdff dff_B_x66oaevu3_3(.din(w_dff_B_YkdDG63U7_3),.dout(w_dff_B_x66oaevu3_3),.clk(gclk));
	jdff dff_A_QYL6DxgV9_0(.dout(w_G4087_4[0]),.din(w_dff_A_QYL6DxgV9_0),.clk(gclk));
	jdff dff_A_OfrUFjPQ7_1(.dout(w_G4087_4[1]),.din(w_dff_A_OfrUFjPQ7_1),.clk(gclk));
	jdff dff_B_A8hND6lq2_1(.din(n1668),.dout(w_dff_B_A8hND6lq2_1),.clk(gclk));
	jdff dff_B_hkA2TYSN3_1(.din(w_dff_B_A8hND6lq2_1),.dout(w_dff_B_hkA2TYSN3_1),.clk(gclk));
	jdff dff_A_ouJpcfxc9_0(.dout(w_n797_3[0]),.din(w_dff_A_ouJpcfxc9_0),.clk(gclk));
	jdff dff_A_12LU00iM3_0(.dout(w_dff_A_ouJpcfxc9_0),.din(w_dff_A_12LU00iM3_0),.clk(gclk));
	jdff dff_A_hSL1wZhs8_0(.dout(w_dff_A_12LU00iM3_0),.din(w_dff_A_hSL1wZhs8_0),.clk(gclk));
	jdff dff_A_HJpLEwt92_0(.dout(w_dff_A_hSL1wZhs8_0),.din(w_dff_A_HJpLEwt92_0),.clk(gclk));
	jdff dff_A_sdQo5WV29_0(.dout(w_dff_A_HJpLEwt92_0),.din(w_dff_A_sdQo5WV29_0),.clk(gclk));
	jdff dff_A_RJoqGr2d3_0(.dout(w_dff_A_sdQo5WV29_0),.din(w_dff_A_RJoqGr2d3_0),.clk(gclk));
	jdff dff_A_9ty7zU8L3_0(.dout(w_dff_A_RJoqGr2d3_0),.din(w_dff_A_9ty7zU8L3_0),.clk(gclk));
	jdff dff_A_7szxLVo21_0(.dout(w_dff_A_9ty7zU8L3_0),.din(w_dff_A_7szxLVo21_0),.clk(gclk));
	jdff dff_A_EnKdrWTh2_0(.dout(w_dff_A_7szxLVo21_0),.din(w_dff_A_EnKdrWTh2_0),.clk(gclk));
	jdff dff_A_ADFmU96c5_0(.dout(w_dff_A_EnKdrWTh2_0),.din(w_dff_A_ADFmU96c5_0),.clk(gclk));
	jdff dff_A_BizjAxo16_0(.dout(w_dff_A_ADFmU96c5_0),.din(w_dff_A_BizjAxo16_0),.clk(gclk));
	jdff dff_A_NFeBwL6s4_0(.dout(w_dff_A_BizjAxo16_0),.din(w_dff_A_NFeBwL6s4_0),.clk(gclk));
	jdff dff_A_iFHkitDq1_0(.dout(w_dff_A_NFeBwL6s4_0),.din(w_dff_A_iFHkitDq1_0),.clk(gclk));
	jdff dff_A_elFdEM5y3_0(.dout(w_dff_A_iFHkitDq1_0),.din(w_dff_A_elFdEM5y3_0),.clk(gclk));
	jdff dff_A_zfcyOCwO3_0(.dout(w_dff_A_elFdEM5y3_0),.din(w_dff_A_zfcyOCwO3_0),.clk(gclk));
	jdff dff_A_sNyB5mEX0_0(.dout(w_dff_A_zfcyOCwO3_0),.din(w_dff_A_sNyB5mEX0_0),.clk(gclk));
	jdff dff_A_bOSgJ2gc0_0(.dout(w_dff_A_sNyB5mEX0_0),.din(w_dff_A_bOSgJ2gc0_0),.clk(gclk));
	jdff dff_A_hJMWeikJ5_0(.dout(w_dff_A_bOSgJ2gc0_0),.din(w_dff_A_hJMWeikJ5_0),.clk(gclk));
	jdff dff_A_bNfrraTM5_0(.dout(w_dff_A_hJMWeikJ5_0),.din(w_dff_A_bNfrraTM5_0),.clk(gclk));
	jdff dff_A_Suo2QwC29_0(.dout(w_dff_A_bNfrraTM5_0),.din(w_dff_A_Suo2QwC29_0),.clk(gclk));
	jdff dff_A_7JHi7eg18_0(.dout(w_dff_A_Suo2QwC29_0),.din(w_dff_A_7JHi7eg18_0),.clk(gclk));
	jdff dff_A_wZ31z6lw8_0(.dout(w_dff_A_7JHi7eg18_0),.din(w_dff_A_wZ31z6lw8_0),.clk(gclk));
	jdff dff_A_F9pE1UfG6_1(.dout(w_G4088_9[1]),.din(w_dff_A_F9pE1UfG6_1),.clk(gclk));
	jdff dff_A_KghyqK1q7_1(.dout(w_dff_A_F9pE1UfG6_1),.din(w_dff_A_KghyqK1q7_1),.clk(gclk));
	jdff dff_A_Hm9r92oa5_1(.dout(w_dff_A_KghyqK1q7_1),.din(w_dff_A_Hm9r92oa5_1),.clk(gclk));
	jdff dff_A_WZAZvzlb7_1(.dout(w_dff_A_Hm9r92oa5_1),.din(w_dff_A_WZAZvzlb7_1),.clk(gclk));
	jdff dff_A_gvhV625k2_1(.dout(w_dff_A_WZAZvzlb7_1),.din(w_dff_A_gvhV625k2_1),.clk(gclk));
	jdff dff_A_sOYq1amW1_1(.dout(w_dff_A_gvhV625k2_1),.din(w_dff_A_sOYq1amW1_1),.clk(gclk));
	jdff dff_A_N7iJ4y353_1(.dout(w_dff_A_sOYq1amW1_1),.din(w_dff_A_N7iJ4y353_1),.clk(gclk));
	jdff dff_A_sZcA6URo5_1(.dout(w_dff_A_N7iJ4y353_1),.din(w_dff_A_sZcA6URo5_1),.clk(gclk));
	jdff dff_A_8wb7EXNr3_1(.dout(w_dff_A_sZcA6URo5_1),.din(w_dff_A_8wb7EXNr3_1),.clk(gclk));
	jdff dff_A_xmdQFswB1_1(.dout(w_G4087_1[1]),.din(w_dff_A_xmdQFswB1_1),.clk(gclk));
	jdff dff_A_Qd0zoQ9U3_1(.dout(w_dff_A_xmdQFswB1_1),.din(w_dff_A_Qd0zoQ9U3_1),.clk(gclk));
	jdff dff_A_huOUs4Y20_2(.dout(w_G4087_1[2]),.din(w_dff_A_huOUs4Y20_2),.clk(gclk));
	jdff dff_A_q6Ybc1Cz7_1(.dout(w_G4087_0[1]),.din(w_dff_A_q6Ybc1Cz7_1),.clk(gclk));
	jdff dff_A_xUOYB4Xr8_2(.dout(w_G4087_0[2]),.din(w_dff_A_xUOYB4Xr8_2),.clk(gclk));
	jdff dff_A_brdJO78o5_0(.dout(w_G4088_3[0]),.din(w_dff_A_brdJO78o5_0),.clk(gclk));
	jdff dff_A_y2a0ACGn3_0(.dout(w_dff_A_brdJO78o5_0),.din(w_dff_A_y2a0ACGn3_0),.clk(gclk));
	jdff dff_A_DSonxTwS0_0(.dout(w_dff_A_y2a0ACGn3_0),.din(w_dff_A_DSonxTwS0_0),.clk(gclk));
	jdff dff_A_5jmEpHNJ9_0(.dout(w_dff_A_DSonxTwS0_0),.din(w_dff_A_5jmEpHNJ9_0),.clk(gclk));
	jdff dff_A_n5eK6xO55_0(.dout(w_dff_A_5jmEpHNJ9_0),.din(w_dff_A_n5eK6xO55_0),.clk(gclk));
	jdff dff_A_AMhzHlyw1_0(.dout(w_dff_A_n5eK6xO55_0),.din(w_dff_A_AMhzHlyw1_0),.clk(gclk));
	jdff dff_A_LM9O3iq19_0(.dout(w_dff_A_AMhzHlyw1_0),.din(w_dff_A_LM9O3iq19_0),.clk(gclk));
	jdff dff_A_yGc5cONx6_0(.dout(w_dff_A_LM9O3iq19_0),.din(w_dff_A_yGc5cONx6_0),.clk(gclk));
	jdff dff_A_nWVBq4qJ2_0(.dout(w_dff_A_yGc5cONx6_0),.din(w_dff_A_nWVBq4qJ2_0),.clk(gclk));
	jdff dff_A_w73qp5rs8_0(.dout(w_dff_A_nWVBq4qJ2_0),.din(w_dff_A_w73qp5rs8_0),.clk(gclk));
	jdff dff_A_tL4Et7y13_0(.dout(w_dff_A_w73qp5rs8_0),.din(w_dff_A_tL4Et7y13_0),.clk(gclk));
	jdff dff_A_4CjAXStS3_0(.dout(w_dff_A_tL4Et7y13_0),.din(w_dff_A_4CjAXStS3_0),.clk(gclk));
	jdff dff_A_MIxjJF3f0_0(.dout(w_dff_A_4CjAXStS3_0),.din(w_dff_A_MIxjJF3f0_0),.clk(gclk));
	jdff dff_A_4VSsuf7r8_0(.dout(w_dff_A_MIxjJF3f0_0),.din(w_dff_A_4VSsuf7r8_0),.clk(gclk));
	jdff dff_A_Jg3el3Hr4_0(.dout(w_dff_A_4VSsuf7r8_0),.din(w_dff_A_Jg3el3Hr4_0),.clk(gclk));
	jdff dff_A_oBrtqtPF7_0(.dout(w_dff_A_Jg3el3Hr4_0),.din(w_dff_A_oBrtqtPF7_0),.clk(gclk));
	jdff dff_A_bV8ocIrG5_0(.dout(w_dff_A_oBrtqtPF7_0),.din(w_dff_A_bV8ocIrG5_0),.clk(gclk));
	jdff dff_A_4vUaiIPe2_0(.dout(w_dff_A_bV8ocIrG5_0),.din(w_dff_A_4vUaiIPe2_0),.clk(gclk));
	jdff dff_A_FdsMZ58L2_0(.dout(w_dff_A_4vUaiIPe2_0),.din(w_dff_A_FdsMZ58L2_0),.clk(gclk));
	jdff dff_A_gYL0V17u2_0(.dout(w_dff_A_FdsMZ58L2_0),.din(w_dff_A_gYL0V17u2_0),.clk(gclk));
	jdff dff_A_v39QAdSF2_0(.dout(w_dff_A_gYL0V17u2_0),.din(w_dff_A_v39QAdSF2_0),.clk(gclk));
	jdff dff_A_SrMSNxNn8_0(.dout(w_dff_A_v39QAdSF2_0),.din(w_dff_A_SrMSNxNn8_0),.clk(gclk));
	jdff dff_A_kH3PP8cX2_0(.dout(w_dff_A_SrMSNxNn8_0),.din(w_dff_A_kH3PP8cX2_0),.clk(gclk));
	jdff dff_B_wWgEURmU6_1(.din(n1688),.dout(w_dff_B_wWgEURmU6_1),.clk(gclk));
	jdff dff_B_6RbDTDSY8_1(.din(w_dff_B_wWgEURmU6_1),.dout(w_dff_B_6RbDTDSY8_1),.clk(gclk));
	jdff dff_B_sjHsPvrq4_1(.din(w_dff_B_6RbDTDSY8_1),.dout(w_dff_B_sjHsPvrq4_1),.clk(gclk));
	jdff dff_B_TylWqUZJ8_1(.din(w_dff_B_sjHsPvrq4_1),.dout(w_dff_B_TylWqUZJ8_1),.clk(gclk));
	jdff dff_B_WMB2ssSy3_1(.din(w_dff_B_TylWqUZJ8_1),.dout(w_dff_B_WMB2ssSy3_1),.clk(gclk));
	jdff dff_B_deotQdSc1_1(.din(w_dff_B_WMB2ssSy3_1),.dout(w_dff_B_deotQdSc1_1),.clk(gclk));
	jdff dff_B_prHKaGzT1_1(.din(w_dff_B_deotQdSc1_1),.dout(w_dff_B_prHKaGzT1_1),.clk(gclk));
	jdff dff_B_cmoVJNVd4_1(.din(w_dff_B_prHKaGzT1_1),.dout(w_dff_B_cmoVJNVd4_1),.clk(gclk));
	jdff dff_B_ECow2kHo5_1(.din(w_dff_B_cmoVJNVd4_1),.dout(w_dff_B_ECow2kHo5_1),.clk(gclk));
	jdff dff_B_UrhRL9iy3_1(.din(w_dff_B_ECow2kHo5_1),.dout(w_dff_B_UrhRL9iy3_1),.clk(gclk));
	jdff dff_B_Drpq8IWm2_1(.din(w_dff_B_UrhRL9iy3_1),.dout(w_dff_B_Drpq8IWm2_1),.clk(gclk));
	jdff dff_B_VbuI1Wgc4_1(.din(w_dff_B_Drpq8IWm2_1),.dout(w_dff_B_VbuI1Wgc4_1),.clk(gclk));
	jdff dff_B_u7BCC4MM6_1(.din(w_dff_B_VbuI1Wgc4_1),.dout(w_dff_B_u7BCC4MM6_1),.clk(gclk));
	jdff dff_B_ggCWKT6J9_1(.din(w_dff_B_u7BCC4MM6_1),.dout(w_dff_B_ggCWKT6J9_1),.clk(gclk));
	jdff dff_B_K72oyMdX8_1(.din(w_dff_B_ggCWKT6J9_1),.dout(w_dff_B_K72oyMdX8_1),.clk(gclk));
	jdff dff_B_nBpREnqN9_1(.din(w_dff_B_K72oyMdX8_1),.dout(w_dff_B_nBpREnqN9_1),.clk(gclk));
	jdff dff_B_HTK439Wq1_1(.din(w_dff_B_nBpREnqN9_1),.dout(w_dff_B_HTK439Wq1_1),.clk(gclk));
	jdff dff_B_mQkpyUbh2_1(.din(w_dff_B_HTK439Wq1_1),.dout(w_dff_B_mQkpyUbh2_1),.clk(gclk));
	jdff dff_B_nakUJG386_1(.din(w_dff_B_mQkpyUbh2_1),.dout(w_dff_B_nakUJG386_1),.clk(gclk));
	jdff dff_B_6UeAQqf66_1(.din(w_dff_B_nakUJG386_1),.dout(w_dff_B_6UeAQqf66_1),.clk(gclk));
	jdff dff_B_xEScLYl45_1(.din(w_dff_B_6UeAQqf66_1),.dout(w_dff_B_xEScLYl45_1),.clk(gclk));
	jdff dff_B_KXlTl6Of8_1(.din(w_dff_B_xEScLYl45_1),.dout(w_dff_B_KXlTl6Of8_1),.clk(gclk));
	jdff dff_B_mpBfkQmG0_1(.din(n1689),.dout(w_dff_B_mpBfkQmG0_1),.clk(gclk));
	jdff dff_A_8CO2i2n78_1(.dout(w_n854_1[1]),.din(w_dff_A_8CO2i2n78_1),.clk(gclk));
	jdff dff_A_m0qmgwmF4_1(.dout(w_dff_A_8CO2i2n78_1),.din(w_dff_A_m0qmgwmF4_1),.clk(gclk));
	jdff dff_A_GABnNBn65_1(.dout(w_dff_A_m0qmgwmF4_1),.din(w_dff_A_GABnNBn65_1),.clk(gclk));
	jdff dff_A_dMeydbTF0_1(.dout(w_dff_A_GABnNBn65_1),.din(w_dff_A_dMeydbTF0_1),.clk(gclk));
	jdff dff_A_XCxnLEyM4_1(.dout(w_dff_A_dMeydbTF0_1),.din(w_dff_A_XCxnLEyM4_1),.clk(gclk));
	jdff dff_A_o0KZ2Ry60_1(.dout(w_dff_A_XCxnLEyM4_1),.din(w_dff_A_o0KZ2Ry60_1),.clk(gclk));
	jdff dff_A_5iQzyDiR2_1(.dout(w_dff_A_o0KZ2Ry60_1),.din(w_dff_A_5iQzyDiR2_1),.clk(gclk));
	jdff dff_A_nv6Uky7c9_1(.dout(w_dff_A_5iQzyDiR2_1),.din(w_dff_A_nv6Uky7c9_1),.clk(gclk));
	jdff dff_A_OhRSnYM09_1(.dout(w_dff_A_nv6Uky7c9_1),.din(w_dff_A_OhRSnYM09_1),.clk(gclk));
	jdff dff_A_eHUfQdXt0_1(.dout(w_dff_A_OhRSnYM09_1),.din(w_dff_A_eHUfQdXt0_1),.clk(gclk));
	jdff dff_A_1EjJS5qT2_1(.dout(w_dff_A_eHUfQdXt0_1),.din(w_dff_A_1EjJS5qT2_1),.clk(gclk));
	jdff dff_A_SBtYyH3t3_1(.dout(w_dff_A_1EjJS5qT2_1),.din(w_dff_A_SBtYyH3t3_1),.clk(gclk));
	jdff dff_A_o5DxYfoU2_1(.dout(w_dff_A_SBtYyH3t3_1),.din(w_dff_A_o5DxYfoU2_1),.clk(gclk));
	jdff dff_A_VXwxUIU01_1(.dout(w_dff_A_o5DxYfoU2_1),.din(w_dff_A_VXwxUIU01_1),.clk(gclk));
	jdff dff_A_IqYpwzBl4_2(.dout(w_n854_1[2]),.din(w_dff_A_IqYpwzBl4_2),.clk(gclk));
	jdff dff_A_owqyUvqg6_2(.dout(w_dff_A_IqYpwzBl4_2),.din(w_dff_A_owqyUvqg6_2),.clk(gclk));
	jdff dff_A_FxL2PiIP3_2(.dout(w_dff_A_owqyUvqg6_2),.din(w_dff_A_FxL2PiIP3_2),.clk(gclk));
	jdff dff_A_oPiS4LRt9_2(.dout(w_dff_A_FxL2PiIP3_2),.din(w_dff_A_oPiS4LRt9_2),.clk(gclk));
	jdff dff_A_diyjyDMc6_2(.dout(w_dff_A_oPiS4LRt9_2),.din(w_dff_A_diyjyDMc6_2),.clk(gclk));
	jdff dff_A_BGpPLwCp0_2(.dout(w_dff_A_diyjyDMc6_2),.din(w_dff_A_BGpPLwCp0_2),.clk(gclk));
	jdff dff_A_2oeB6MbB8_2(.dout(w_dff_A_BGpPLwCp0_2),.din(w_dff_A_2oeB6MbB8_2),.clk(gclk));
	jdff dff_A_8p5hOO8r7_2(.dout(w_dff_A_2oeB6MbB8_2),.din(w_dff_A_8p5hOO8r7_2),.clk(gclk));
	jdff dff_A_UHVhXrBV7_2(.dout(w_dff_A_8p5hOO8r7_2),.din(w_dff_A_UHVhXrBV7_2),.clk(gclk));
	jdff dff_A_nkBS7BN47_2(.dout(w_dff_A_UHVhXrBV7_2),.din(w_dff_A_nkBS7BN47_2),.clk(gclk));
	jdff dff_A_DaTcnhiw0_1(.dout(w_n854_0[1]),.din(w_dff_A_DaTcnhiw0_1),.clk(gclk));
	jdff dff_A_KOZClzYI2_1(.dout(w_dff_A_DaTcnhiw0_1),.din(w_dff_A_KOZClzYI2_1),.clk(gclk));
	jdff dff_A_43adTSv83_1(.dout(w_dff_A_KOZClzYI2_1),.din(w_dff_A_43adTSv83_1),.clk(gclk));
	jdff dff_A_Tk4bY1Up4_1(.dout(w_dff_A_43adTSv83_1),.din(w_dff_A_Tk4bY1Up4_1),.clk(gclk));
	jdff dff_A_r54mcXYe8_1(.dout(w_dff_A_Tk4bY1Up4_1),.din(w_dff_A_r54mcXYe8_1),.clk(gclk));
	jdff dff_A_trPqvmZV0_1(.dout(w_dff_A_r54mcXYe8_1),.din(w_dff_A_trPqvmZV0_1),.clk(gclk));
	jdff dff_A_OJ9QNloY1_1(.dout(w_dff_A_trPqvmZV0_1),.din(w_dff_A_OJ9QNloY1_1),.clk(gclk));
	jdff dff_A_KibaWw0P6_1(.dout(w_dff_A_OJ9QNloY1_1),.din(w_dff_A_KibaWw0P6_1),.clk(gclk));
	jdff dff_A_Wrm4RB169_1(.dout(w_dff_A_KibaWw0P6_1),.din(w_dff_A_Wrm4RB169_1),.clk(gclk));
	jdff dff_A_QXVvkGMr7_1(.dout(w_dff_A_Wrm4RB169_1),.din(w_dff_A_QXVvkGMr7_1),.clk(gclk));
	jdff dff_A_M28Bwhdm8_1(.dout(w_dff_A_QXVvkGMr7_1),.din(w_dff_A_M28Bwhdm8_1),.clk(gclk));
	jdff dff_A_rl4KCP451_2(.dout(w_n854_0[2]),.din(w_dff_A_rl4KCP451_2),.clk(gclk));
	jdff dff_A_6D0AXka91_2(.dout(w_dff_A_rl4KCP451_2),.din(w_dff_A_6D0AXka91_2),.clk(gclk));
	jdff dff_A_tvVAPV5y0_2(.dout(w_dff_A_6D0AXka91_2),.din(w_dff_A_tvVAPV5y0_2),.clk(gclk));
	jdff dff_A_ot9sPm6n9_2(.dout(w_dff_A_tvVAPV5y0_2),.din(w_dff_A_ot9sPm6n9_2),.clk(gclk));
	jdff dff_A_sm2eBv348_2(.dout(w_dff_A_ot9sPm6n9_2),.din(w_dff_A_sm2eBv348_2),.clk(gclk));
	jdff dff_B_0qH55en87_3(.din(n854),.dout(w_dff_B_0qH55en87_3),.clk(gclk));
	jdff dff_B_fIOicQFV5_3(.din(w_dff_B_0qH55en87_3),.dout(w_dff_B_fIOicQFV5_3),.clk(gclk));
	jdff dff_B_CTQbOwnL9_3(.din(w_dff_B_fIOicQFV5_3),.dout(w_dff_B_CTQbOwnL9_3),.clk(gclk));
	jdff dff_B_yXMAhMSb3_3(.din(w_dff_B_CTQbOwnL9_3),.dout(w_dff_B_yXMAhMSb3_3),.clk(gclk));
	jdff dff_B_vHJR4ZOj0_3(.din(w_dff_B_yXMAhMSb3_3),.dout(w_dff_B_vHJR4ZOj0_3),.clk(gclk));
	jdff dff_B_yHu6d2yL6_3(.din(w_dff_B_vHJR4ZOj0_3),.dout(w_dff_B_yHu6d2yL6_3),.clk(gclk));
	jdff dff_B_38IArHka8_3(.din(w_dff_B_yHu6d2yL6_3),.dout(w_dff_B_38IArHka8_3),.clk(gclk));
	jdff dff_B_6H7KQBPs7_3(.din(w_dff_B_38IArHka8_3),.dout(w_dff_B_6H7KQBPs7_3),.clk(gclk));
	jdff dff_B_x6sYVZQl0_3(.din(w_dff_B_6H7KQBPs7_3),.dout(w_dff_B_x6sYVZQl0_3),.clk(gclk));
	jdff dff_A_Ha3cWrG17_0(.dout(w_G4090_4[0]),.din(w_dff_A_Ha3cWrG17_0),.clk(gclk));
	jdff dff_A_8kpK9Msz0_0(.dout(w_dff_A_Ha3cWrG17_0),.din(w_dff_A_8kpK9Msz0_0),.clk(gclk));
	jdff dff_A_26cKSgzW0_1(.dout(w_G4090_4[1]),.din(w_dff_A_26cKSgzW0_1),.clk(gclk));
	jdff dff_B_XPvaKtdg5_1(.din(n1685),.dout(w_dff_B_XPvaKtdg5_1),.clk(gclk));
	jdff dff_B_BTPIfn9Y7_1(.din(w_dff_B_XPvaKtdg5_1),.dout(w_dff_B_BTPIfn9Y7_1),.clk(gclk));
	jdff dff_A_1kJQdAkM7_0(.dout(w_n852_3[0]),.din(w_dff_A_1kJQdAkM7_0),.clk(gclk));
	jdff dff_A_xtTjGC7B2_0(.dout(w_dff_A_1kJQdAkM7_0),.din(w_dff_A_xtTjGC7B2_0),.clk(gclk));
	jdff dff_A_tumRi2mC0_0(.dout(w_dff_A_xtTjGC7B2_0),.din(w_dff_A_tumRi2mC0_0),.clk(gclk));
	jdff dff_A_5d8H4D965_0(.dout(w_dff_A_tumRi2mC0_0),.din(w_dff_A_5d8H4D965_0),.clk(gclk));
	jdff dff_A_t4LOqunI9_0(.dout(w_dff_A_5d8H4D965_0),.din(w_dff_A_t4LOqunI9_0),.clk(gclk));
	jdff dff_A_lvXE7poB5_0(.dout(w_dff_A_t4LOqunI9_0),.din(w_dff_A_lvXE7poB5_0),.clk(gclk));
	jdff dff_A_JrSzFae68_0(.dout(w_dff_A_lvXE7poB5_0),.din(w_dff_A_JrSzFae68_0),.clk(gclk));
	jdff dff_A_wl3A6yNu6_0(.dout(w_dff_A_JrSzFae68_0),.din(w_dff_A_wl3A6yNu6_0),.clk(gclk));
	jdff dff_A_e2NVKZAD3_0(.dout(w_dff_A_wl3A6yNu6_0),.din(w_dff_A_e2NVKZAD3_0),.clk(gclk));
	jdff dff_A_30FZuT7V4_0(.dout(w_dff_A_e2NVKZAD3_0),.din(w_dff_A_30FZuT7V4_0),.clk(gclk));
	jdff dff_A_VFU3y2Mj3_0(.dout(w_dff_A_30FZuT7V4_0),.din(w_dff_A_VFU3y2Mj3_0),.clk(gclk));
	jdff dff_A_yYh1NV9p7_0(.dout(w_dff_A_VFU3y2Mj3_0),.din(w_dff_A_yYh1NV9p7_0),.clk(gclk));
	jdff dff_A_fUWMkXjP4_0(.dout(w_dff_A_yYh1NV9p7_0),.din(w_dff_A_fUWMkXjP4_0),.clk(gclk));
	jdff dff_A_50TLP7jU3_0(.dout(w_dff_A_fUWMkXjP4_0),.din(w_dff_A_50TLP7jU3_0),.clk(gclk));
	jdff dff_A_EZxFsrWR7_0(.dout(w_dff_A_50TLP7jU3_0),.din(w_dff_A_EZxFsrWR7_0),.clk(gclk));
	jdff dff_A_zCOHU7d92_0(.dout(w_dff_A_EZxFsrWR7_0),.din(w_dff_A_zCOHU7d92_0),.clk(gclk));
	jdff dff_A_ZEJQY0ik1_0(.dout(w_dff_A_zCOHU7d92_0),.din(w_dff_A_ZEJQY0ik1_0),.clk(gclk));
	jdff dff_A_mfdDrOci0_0(.dout(w_dff_A_ZEJQY0ik1_0),.din(w_dff_A_mfdDrOci0_0),.clk(gclk));
	jdff dff_A_knC7x9lC2_0(.dout(w_dff_A_mfdDrOci0_0),.din(w_dff_A_knC7x9lC2_0),.clk(gclk));
	jdff dff_A_VHtaA9oV7_0(.dout(w_dff_A_knC7x9lC2_0),.din(w_dff_A_VHtaA9oV7_0),.clk(gclk));
	jdff dff_A_mL9wRMd47_0(.dout(w_dff_A_VHtaA9oV7_0),.din(w_dff_A_mL9wRMd47_0),.clk(gclk));
	jdff dff_A_9DvEUrSW2_0(.dout(w_dff_A_mL9wRMd47_0),.din(w_dff_A_9DvEUrSW2_0),.clk(gclk));
	jdff dff_A_hbAMZKfq7_1(.dout(w_G4089_9[1]),.din(w_dff_A_hbAMZKfq7_1),.clk(gclk));
	jdff dff_A_vmjKJRSN1_1(.dout(w_dff_A_hbAMZKfq7_1),.din(w_dff_A_vmjKJRSN1_1),.clk(gclk));
	jdff dff_A_Tiajxx3A1_1(.dout(w_dff_A_vmjKJRSN1_1),.din(w_dff_A_Tiajxx3A1_1),.clk(gclk));
	jdff dff_A_oWsllihA0_1(.dout(w_dff_A_Tiajxx3A1_1),.din(w_dff_A_oWsllihA0_1),.clk(gclk));
	jdff dff_A_5YVu1MZ45_1(.dout(w_dff_A_oWsllihA0_1),.din(w_dff_A_5YVu1MZ45_1),.clk(gclk));
	jdff dff_A_g70oY7j37_1(.dout(w_dff_A_5YVu1MZ45_1),.din(w_dff_A_g70oY7j37_1),.clk(gclk));
	jdff dff_A_du8J4sTC8_1(.dout(w_dff_A_g70oY7j37_1),.din(w_dff_A_du8J4sTC8_1),.clk(gclk));
	jdff dff_A_p6eEK0KJ2_1(.dout(w_dff_A_du8J4sTC8_1),.din(w_dff_A_p6eEK0KJ2_1),.clk(gclk));
	jdff dff_A_I5dEYBgk2_1(.dout(w_dff_A_p6eEK0KJ2_1),.din(w_dff_A_I5dEYBgk2_1),.clk(gclk));
	jdff dff_B_elWrQJ4U4_2(.din(G64),.dout(w_dff_B_elWrQJ4U4_2),.clk(gclk));
	jdff dff_A_J7W1hXpk2_1(.dout(w_G4090_1[1]),.din(w_dff_A_J7W1hXpk2_1),.clk(gclk));
	jdff dff_A_ksc0atqM3_1(.dout(w_dff_A_J7W1hXpk2_1),.din(w_dff_A_ksc0atqM3_1),.clk(gclk));
	jdff dff_A_sRvNW2HZ1_2(.dout(w_G4090_1[2]),.din(w_dff_A_sRvNW2HZ1_2),.clk(gclk));
	jdff dff_A_BYXvFlgx9_1(.dout(w_G4090_0[1]),.din(w_dff_A_BYXvFlgx9_1),.clk(gclk));
	jdff dff_A_f0KPsERX4_2(.dout(w_G4090_0[2]),.din(w_dff_A_f0KPsERX4_2),.clk(gclk));
	jdff dff_A_5bHnMgvO1_0(.dout(w_G4089_3[0]),.din(w_dff_A_5bHnMgvO1_0),.clk(gclk));
	jdff dff_A_NcOI8saR6_0(.dout(w_dff_A_5bHnMgvO1_0),.din(w_dff_A_NcOI8saR6_0),.clk(gclk));
	jdff dff_A_AAY4v8W08_0(.dout(w_dff_A_NcOI8saR6_0),.din(w_dff_A_AAY4v8W08_0),.clk(gclk));
	jdff dff_A_Y2CJTJSH4_0(.dout(w_dff_A_AAY4v8W08_0),.din(w_dff_A_Y2CJTJSH4_0),.clk(gclk));
	jdff dff_A_WXvvYtay2_0(.dout(w_dff_A_Y2CJTJSH4_0),.din(w_dff_A_WXvvYtay2_0),.clk(gclk));
	jdff dff_A_sRvXD0DF0_0(.dout(w_dff_A_WXvvYtay2_0),.din(w_dff_A_sRvXD0DF0_0),.clk(gclk));
	jdff dff_A_rYlRiy2b1_0(.dout(w_dff_A_sRvXD0DF0_0),.din(w_dff_A_rYlRiy2b1_0),.clk(gclk));
	jdff dff_A_gDuGQ8eQ2_0(.dout(w_dff_A_rYlRiy2b1_0),.din(w_dff_A_gDuGQ8eQ2_0),.clk(gclk));
	jdff dff_A_x3ZlMNPZ7_0(.dout(w_dff_A_gDuGQ8eQ2_0),.din(w_dff_A_x3ZlMNPZ7_0),.clk(gclk));
	jdff dff_A_xZ2iOT8N9_0(.dout(w_dff_A_x3ZlMNPZ7_0),.din(w_dff_A_xZ2iOT8N9_0),.clk(gclk));
	jdff dff_A_YuXCB6yR0_0(.dout(w_dff_A_xZ2iOT8N9_0),.din(w_dff_A_YuXCB6yR0_0),.clk(gclk));
	jdff dff_A_5SncczX37_0(.dout(w_dff_A_YuXCB6yR0_0),.din(w_dff_A_5SncczX37_0),.clk(gclk));
	jdff dff_A_xctXUhwh6_0(.dout(w_dff_A_5SncczX37_0),.din(w_dff_A_xctXUhwh6_0),.clk(gclk));
	jdff dff_A_OiIq1dkr0_0(.dout(w_dff_A_xctXUhwh6_0),.din(w_dff_A_OiIq1dkr0_0),.clk(gclk));
	jdff dff_A_07BlpJUB8_0(.dout(w_dff_A_OiIq1dkr0_0),.din(w_dff_A_07BlpJUB8_0),.clk(gclk));
	jdff dff_A_WcGox2sJ8_0(.dout(w_dff_A_07BlpJUB8_0),.din(w_dff_A_WcGox2sJ8_0),.clk(gclk));
	jdff dff_A_ra6KoJbO5_0(.dout(w_dff_A_WcGox2sJ8_0),.din(w_dff_A_ra6KoJbO5_0),.clk(gclk));
	jdff dff_A_7Qshy0Zq4_0(.dout(w_dff_A_ra6KoJbO5_0),.din(w_dff_A_7Qshy0Zq4_0),.clk(gclk));
	jdff dff_A_NtQSdMAy2_0(.dout(w_dff_A_7Qshy0Zq4_0),.din(w_dff_A_NtQSdMAy2_0),.clk(gclk));
	jdff dff_A_lm9sZBkW6_0(.dout(w_dff_A_NtQSdMAy2_0),.din(w_dff_A_lm9sZBkW6_0),.clk(gclk));
	jdff dff_A_r609rUzY5_0(.dout(w_dff_A_lm9sZBkW6_0),.din(w_dff_A_r609rUzY5_0),.clk(gclk));
	jdff dff_A_r2wKOvRB6_0(.dout(w_dff_A_r609rUzY5_0),.din(w_dff_A_r2wKOvRB6_0),.clk(gclk));
	jdff dff_A_EoOpLKUe9_0(.dout(w_dff_A_r2wKOvRB6_0),.din(w_dff_A_EoOpLKUe9_0),.clk(gclk));
	jdff dff_B_11fBWxV75_1(.din(n1697),.dout(w_dff_B_11fBWxV75_1),.clk(gclk));
	jdff dff_B_FXIPiwZP5_1(.din(w_dff_B_11fBWxV75_1),.dout(w_dff_B_FXIPiwZP5_1),.clk(gclk));
	jdff dff_B_S06WoP7R8_1(.din(w_dff_B_FXIPiwZP5_1),.dout(w_dff_B_S06WoP7R8_1),.clk(gclk));
	jdff dff_B_btFqaB1x0_1(.din(w_dff_B_S06WoP7R8_1),.dout(w_dff_B_btFqaB1x0_1),.clk(gclk));
	jdff dff_B_OrAOC1Ty0_1(.din(w_dff_B_btFqaB1x0_1),.dout(w_dff_B_OrAOC1Ty0_1),.clk(gclk));
	jdff dff_B_CJRag0Yy6_1(.din(w_dff_B_OrAOC1Ty0_1),.dout(w_dff_B_CJRag0Yy6_1),.clk(gclk));
	jdff dff_B_oyELLvTh7_1(.din(w_dff_B_CJRag0Yy6_1),.dout(w_dff_B_oyELLvTh7_1),.clk(gclk));
	jdff dff_B_SYYQl30m5_1(.din(w_dff_B_oyELLvTh7_1),.dout(w_dff_B_SYYQl30m5_1),.clk(gclk));
	jdff dff_B_3FIhqHQg4_1(.din(w_dff_B_SYYQl30m5_1),.dout(w_dff_B_3FIhqHQg4_1),.clk(gclk));
	jdff dff_B_TxWDfSME5_1(.din(w_dff_B_3FIhqHQg4_1),.dout(w_dff_B_TxWDfSME5_1),.clk(gclk));
	jdff dff_B_c0yzu0w89_1(.din(w_dff_B_TxWDfSME5_1),.dout(w_dff_B_c0yzu0w89_1),.clk(gclk));
	jdff dff_B_XdpeJQ4V3_1(.din(w_dff_B_c0yzu0w89_1),.dout(w_dff_B_XdpeJQ4V3_1),.clk(gclk));
	jdff dff_B_AcwP5iZV3_1(.din(w_dff_B_XdpeJQ4V3_1),.dout(w_dff_B_AcwP5iZV3_1),.clk(gclk));
	jdff dff_B_VHsBF9nZ9_1(.din(w_dff_B_AcwP5iZV3_1),.dout(w_dff_B_VHsBF9nZ9_1),.clk(gclk));
	jdff dff_B_qesynLFK6_1(.din(w_dff_B_VHsBF9nZ9_1),.dout(w_dff_B_qesynLFK6_1),.clk(gclk));
	jdff dff_B_A5gozeRD2_1(.din(w_dff_B_qesynLFK6_1),.dout(w_dff_B_A5gozeRD2_1),.clk(gclk));
	jdff dff_B_7V00o5xe1_1(.din(w_dff_B_A5gozeRD2_1),.dout(w_dff_B_7V00o5xe1_1),.clk(gclk));
	jdff dff_B_otCXgSgC8_1(.din(w_dff_B_7V00o5xe1_1),.dout(w_dff_B_otCXgSgC8_1),.clk(gclk));
	jdff dff_B_0hJ2ADGE9_1(.din(w_dff_B_otCXgSgC8_1),.dout(w_dff_B_0hJ2ADGE9_1),.clk(gclk));
	jdff dff_B_QRkYaDOT7_1(.din(w_dff_B_0hJ2ADGE9_1),.dout(w_dff_B_QRkYaDOT7_1),.clk(gclk));
	jdff dff_B_8i9nuOTJ5_1(.din(w_dff_B_QRkYaDOT7_1),.dout(w_dff_B_8i9nuOTJ5_1),.clk(gclk));
	jdff dff_B_7IEUh2D10_1(.din(w_dff_B_8i9nuOTJ5_1),.dout(w_dff_B_7IEUh2D10_1),.clk(gclk));
	jdff dff_B_e9Ghi6we9_1(.din(w_dff_B_7IEUh2D10_1),.dout(w_dff_B_e9Ghi6we9_1),.clk(gclk));
	jdff dff_B_qvliIxqM3_1(.din(n1700),.dout(w_dff_B_qvliIxqM3_1),.clk(gclk));
	jdff dff_B_9Zn9xc292_1(.din(w_dff_B_qvliIxqM3_1),.dout(w_dff_B_9Zn9xc292_1),.clk(gclk));
	jdff dff_B_KjZ2BQb95_1(.din(w_dff_B_9Zn9xc292_1),.dout(w_dff_B_KjZ2BQb95_1),.clk(gclk));
	jdff dff_B_4KVRDxTW8_1(.din(w_dff_B_KjZ2BQb95_1),.dout(w_dff_B_4KVRDxTW8_1),.clk(gclk));
	jdff dff_B_ZWqa6y3m1_1(.din(w_dff_B_4KVRDxTW8_1),.dout(w_dff_B_ZWqa6y3m1_1),.clk(gclk));
	jdff dff_B_lJcCMNJ15_1(.din(w_dff_B_ZWqa6y3m1_1),.dout(w_dff_B_lJcCMNJ15_1),.clk(gclk));
	jdff dff_B_C4rCKfyl7_1(.din(w_dff_B_lJcCMNJ15_1),.dout(w_dff_B_C4rCKfyl7_1),.clk(gclk));
	jdff dff_B_E5hECoeZ3_1(.din(w_dff_B_C4rCKfyl7_1),.dout(w_dff_B_E5hECoeZ3_1),.clk(gclk));
	jdff dff_B_gXlz2jwY6_1(.din(w_dff_B_E5hECoeZ3_1),.dout(w_dff_B_gXlz2jwY6_1),.clk(gclk));
	jdff dff_B_6VLSEagO9_1(.din(w_dff_B_gXlz2jwY6_1),.dout(w_dff_B_6VLSEagO9_1),.clk(gclk));
	jdff dff_B_cym21weM8_1(.din(w_dff_B_6VLSEagO9_1),.dout(w_dff_B_cym21weM8_1),.clk(gclk));
	jdff dff_B_paNP8PIy2_1(.din(w_dff_B_cym21weM8_1),.dout(w_dff_B_paNP8PIy2_1),.clk(gclk));
	jdff dff_B_GaLW9uUh6_1(.din(w_dff_B_paNP8PIy2_1),.dout(w_dff_B_GaLW9uUh6_1),.clk(gclk));
	jdff dff_B_QZiAHxv07_1(.din(w_dff_B_GaLW9uUh6_1),.dout(w_dff_B_QZiAHxv07_1),.clk(gclk));
	jdff dff_B_uP6EeV9O2_1(.din(w_dff_B_QZiAHxv07_1),.dout(w_dff_B_uP6EeV9O2_1),.clk(gclk));
	jdff dff_B_7HbNEO788_1(.din(w_dff_B_uP6EeV9O2_1),.dout(w_dff_B_7HbNEO788_1),.clk(gclk));
	jdff dff_B_1OTuK1qe0_1(.din(w_dff_B_7HbNEO788_1),.dout(w_dff_B_1OTuK1qe0_1),.clk(gclk));
	jdff dff_B_TPuzgZuV2_1(.din(w_dff_B_1OTuK1qe0_1),.dout(w_dff_B_TPuzgZuV2_1),.clk(gclk));
	jdff dff_B_cvKNrSBj8_1(.din(w_dff_B_TPuzgZuV2_1),.dout(w_dff_B_cvKNrSBj8_1),.clk(gclk));
	jdff dff_B_btY59Hp39_1(.din(w_dff_B_cvKNrSBj8_1),.dout(w_dff_B_btY59Hp39_1),.clk(gclk));
	jdff dff_B_67NfPwbU8_1(.din(w_dff_B_btY59Hp39_1),.dout(w_dff_B_67NfPwbU8_1),.clk(gclk));
	jdff dff_B_yJssm8oz1_1(.din(n1701),.dout(w_dff_B_yJssm8oz1_1),.clk(gclk));
	jdff dff_A_TRNTqb8g7_0(.dout(w_n993_4[0]),.din(w_dff_A_TRNTqb8g7_0),.clk(gclk));
	jdff dff_A_X5YbrzOk1_0(.dout(w_dff_A_TRNTqb8g7_0),.din(w_dff_A_X5YbrzOk1_0),.clk(gclk));
	jdff dff_A_IDWv58Lr6_0(.dout(w_dff_A_X5YbrzOk1_0),.din(w_dff_A_IDWv58Lr6_0),.clk(gclk));
	jdff dff_A_ZfHDAFS63_0(.dout(w_dff_A_IDWv58Lr6_0),.din(w_dff_A_ZfHDAFS63_0),.clk(gclk));
	jdff dff_A_iQJ7qmd52_0(.dout(w_dff_A_ZfHDAFS63_0),.din(w_dff_A_iQJ7qmd52_0),.clk(gclk));
	jdff dff_A_Y3WZuILJ2_0(.dout(w_dff_A_iQJ7qmd52_0),.din(w_dff_A_Y3WZuILJ2_0),.clk(gclk));
	jdff dff_A_XpehRAJP9_0(.dout(w_dff_A_Y3WZuILJ2_0),.din(w_dff_A_XpehRAJP9_0),.clk(gclk));
	jdff dff_A_zjPyLzpi2_0(.dout(w_dff_A_XpehRAJP9_0),.din(w_dff_A_zjPyLzpi2_0),.clk(gclk));
	jdff dff_A_3NQp8nO86_0(.dout(w_dff_A_zjPyLzpi2_0),.din(w_dff_A_3NQp8nO86_0),.clk(gclk));
	jdff dff_A_LwYGzmdy1_0(.dout(w_dff_A_3NQp8nO86_0),.din(w_dff_A_LwYGzmdy1_0),.clk(gclk));
	jdff dff_A_S5FsDPRN0_0(.dout(w_dff_A_LwYGzmdy1_0),.din(w_dff_A_S5FsDPRN0_0),.clk(gclk));
	jdff dff_A_5uSh1v011_0(.dout(w_dff_A_S5FsDPRN0_0),.din(w_dff_A_5uSh1v011_0),.clk(gclk));
	jdff dff_A_yAi5FUeR2_0(.dout(w_dff_A_5uSh1v011_0),.din(w_dff_A_yAi5FUeR2_0),.clk(gclk));
	jdff dff_A_Ti2KgWbf0_0(.dout(w_dff_A_yAi5FUeR2_0),.din(w_dff_A_Ti2KgWbf0_0),.clk(gclk));
	jdff dff_A_RiCzsvby6_0(.dout(w_dff_A_Ti2KgWbf0_0),.din(w_dff_A_RiCzsvby6_0),.clk(gclk));
	jdff dff_A_Q4yZm4bD6_1(.dout(w_n993_4[1]),.din(w_dff_A_Q4yZm4bD6_1),.clk(gclk));
	jdff dff_A_g2SDyqyM2_1(.dout(w_dff_A_Q4yZm4bD6_1),.din(w_dff_A_g2SDyqyM2_1),.clk(gclk));
	jdff dff_A_oMrIZnTf2_1(.dout(w_dff_A_g2SDyqyM2_1),.din(w_dff_A_oMrIZnTf2_1),.clk(gclk));
	jdff dff_A_RPm7PPa61_1(.dout(w_dff_A_oMrIZnTf2_1),.din(w_dff_A_RPm7PPa61_1),.clk(gclk));
	jdff dff_A_5QFWDxTx5_1(.dout(w_dff_A_RPm7PPa61_1),.din(w_dff_A_5QFWDxTx5_1),.clk(gclk));
	jdff dff_A_wKAjSvf32_1(.dout(w_dff_A_5QFWDxTx5_1),.din(w_dff_A_wKAjSvf32_1),.clk(gclk));
	jdff dff_A_Ndw55JCg7_1(.dout(w_dff_A_wKAjSvf32_1),.din(w_dff_A_Ndw55JCg7_1),.clk(gclk));
	jdff dff_A_wZ1L0jbV0_1(.dout(w_dff_A_Ndw55JCg7_1),.din(w_dff_A_wZ1L0jbV0_1),.clk(gclk));
	jdff dff_A_eoxyatnW6_1(.dout(w_dff_A_wZ1L0jbV0_1),.din(w_dff_A_eoxyatnW6_1),.clk(gclk));
	jdff dff_A_svDBm8Jc3_1(.dout(w_dff_A_eoxyatnW6_1),.din(w_dff_A_svDBm8Jc3_1),.clk(gclk));
	jdff dff_A_8LsS5AGs9_1(.dout(w_n993_1[1]),.din(w_dff_A_8LsS5AGs9_1),.clk(gclk));
	jdff dff_A_Hzv45t1J9_1(.dout(w_dff_A_8LsS5AGs9_1),.din(w_dff_A_Hzv45t1J9_1),.clk(gclk));
	jdff dff_A_l0mfcFzJ7_1(.dout(w_dff_A_Hzv45t1J9_1),.din(w_dff_A_l0mfcFzJ7_1),.clk(gclk));
	jdff dff_A_mpCLWfXX3_1(.dout(w_dff_A_l0mfcFzJ7_1),.din(w_dff_A_mpCLWfXX3_1),.clk(gclk));
	jdff dff_A_k114UFWy1_1(.dout(w_dff_A_mpCLWfXX3_1),.din(w_dff_A_k114UFWy1_1),.clk(gclk));
	jdff dff_A_isexrxmM3_1(.dout(w_dff_A_k114UFWy1_1),.din(w_dff_A_isexrxmM3_1),.clk(gclk));
	jdff dff_A_GUbHTYic0_1(.dout(w_dff_A_isexrxmM3_1),.din(w_dff_A_GUbHTYic0_1),.clk(gclk));
	jdff dff_A_YxFsmCUO9_1(.dout(w_dff_A_GUbHTYic0_1),.din(w_dff_A_YxFsmCUO9_1),.clk(gclk));
	jdff dff_A_7WzjAGkN5_1(.dout(w_dff_A_YxFsmCUO9_1),.din(w_dff_A_7WzjAGkN5_1),.clk(gclk));
	jdff dff_A_Cfa3sRpq4_1(.dout(w_dff_A_7WzjAGkN5_1),.din(w_dff_A_Cfa3sRpq4_1),.clk(gclk));
	jdff dff_A_pJUeIIJh9_1(.dout(w_dff_A_Cfa3sRpq4_1),.din(w_dff_A_pJUeIIJh9_1),.clk(gclk));
	jdff dff_A_g3NAHuLU2_1(.dout(w_dff_A_pJUeIIJh9_1),.din(w_dff_A_g3NAHuLU2_1),.clk(gclk));
	jdff dff_A_L9QpcrDr6_1(.dout(w_dff_A_g3NAHuLU2_1),.din(w_dff_A_L9QpcrDr6_1),.clk(gclk));
	jdff dff_A_X4UDypwM9_1(.dout(w_dff_A_L9QpcrDr6_1),.din(w_dff_A_X4UDypwM9_1),.clk(gclk));
	jdff dff_A_BBPxCpfw1_1(.dout(w_dff_A_X4UDypwM9_1),.din(w_dff_A_BBPxCpfw1_1),.clk(gclk));
	jdff dff_A_fyusDvm38_1(.dout(w_dff_A_BBPxCpfw1_1),.din(w_dff_A_fyusDvm38_1),.clk(gclk));
	jdff dff_A_r8gYdgL39_1(.dout(w_dff_A_fyusDvm38_1),.din(w_dff_A_r8gYdgL39_1),.clk(gclk));
	jdff dff_A_0uuR7mHC8_1(.dout(w_dff_A_r8gYdgL39_1),.din(w_dff_A_0uuR7mHC8_1),.clk(gclk));
	jdff dff_A_pHuy2eHG2_1(.dout(w_dff_A_0uuR7mHC8_1),.din(w_dff_A_pHuy2eHG2_1),.clk(gclk));
	jdff dff_A_79esEI9F5_1(.dout(w_dff_A_pHuy2eHG2_1),.din(w_dff_A_79esEI9F5_1),.clk(gclk));
	jdff dff_A_4fDZu6Ro7_1(.dout(w_dff_A_79esEI9F5_1),.din(w_dff_A_4fDZu6Ro7_1),.clk(gclk));
	jdff dff_A_bhHgnIga9_2(.dout(w_n993_1[2]),.din(w_dff_A_bhHgnIga9_2),.clk(gclk));
	jdff dff_A_2ZpLNvk60_2(.dout(w_dff_A_bhHgnIga9_2),.din(w_dff_A_2ZpLNvk60_2),.clk(gclk));
	jdff dff_A_w41nB2O55_2(.dout(w_dff_A_2ZpLNvk60_2),.din(w_dff_A_w41nB2O55_2),.clk(gclk));
	jdff dff_A_TbQbsKlG1_2(.dout(w_dff_A_w41nB2O55_2),.din(w_dff_A_TbQbsKlG1_2),.clk(gclk));
	jdff dff_A_dTJhylH06_2(.dout(w_dff_A_TbQbsKlG1_2),.din(w_dff_A_dTJhylH06_2),.clk(gclk));
	jdff dff_A_36FRNv1h1_2(.dout(w_dff_A_dTJhylH06_2),.din(w_dff_A_36FRNv1h1_2),.clk(gclk));
	jdff dff_A_T3dr5okc6_2(.dout(w_dff_A_36FRNv1h1_2),.din(w_dff_A_T3dr5okc6_2),.clk(gclk));
	jdff dff_A_xxeHe6pM4_2(.dout(w_dff_A_T3dr5okc6_2),.din(w_dff_A_xxeHe6pM4_2),.clk(gclk));
	jdff dff_A_2IVIVj9N2_2(.dout(w_dff_A_xxeHe6pM4_2),.din(w_dff_A_2IVIVj9N2_2),.clk(gclk));
	jdff dff_A_BxGFoL9k0_2(.dout(w_dff_A_2IVIVj9N2_2),.din(w_dff_A_BxGFoL9k0_2),.clk(gclk));
	jdff dff_A_jtMf4PbW9_2(.dout(w_dff_A_BxGFoL9k0_2),.din(w_dff_A_jtMf4PbW9_2),.clk(gclk));
	jdff dff_A_S2GKDEcz2_2(.dout(w_dff_A_jtMf4PbW9_2),.din(w_dff_A_S2GKDEcz2_2),.clk(gclk));
	jdff dff_A_WDIrb1ft6_2(.dout(w_dff_A_S2GKDEcz2_2),.din(w_dff_A_WDIrb1ft6_2),.clk(gclk));
	jdff dff_A_mJwO8NvT9_2(.dout(w_dff_A_WDIrb1ft6_2),.din(w_dff_A_mJwO8NvT9_2),.clk(gclk));
	jdff dff_A_RkUI6C059_2(.dout(w_dff_A_mJwO8NvT9_2),.din(w_dff_A_RkUI6C059_2),.clk(gclk));
	jdff dff_A_vHeYE6ai7_2(.dout(w_dff_A_RkUI6C059_2),.din(w_dff_A_vHeYE6ai7_2),.clk(gclk));
	jdff dff_A_4k2iyqIT3_2(.dout(w_dff_A_vHeYE6ai7_2),.din(w_dff_A_4k2iyqIT3_2),.clk(gclk));
	jdff dff_A_aCnRQ2sd0_2(.dout(w_dff_A_4k2iyqIT3_2),.din(w_dff_A_aCnRQ2sd0_2),.clk(gclk));
	jdff dff_A_EHXd7r9L3_2(.dout(w_dff_A_aCnRQ2sd0_2),.din(w_dff_A_EHXd7r9L3_2),.clk(gclk));
	jdff dff_A_0ShZnwgW3_2(.dout(w_dff_A_EHXd7r9L3_2),.din(w_dff_A_0ShZnwgW3_2),.clk(gclk));
	jdff dff_A_Ts5ejSxw1_1(.dout(w_n993_0[1]),.din(w_dff_A_Ts5ejSxw1_1),.clk(gclk));
	jdff dff_A_CDe73UGK4_1(.dout(w_dff_A_Ts5ejSxw1_1),.din(w_dff_A_CDe73UGK4_1),.clk(gclk));
	jdff dff_A_bByk705m9_1(.dout(w_dff_A_CDe73UGK4_1),.din(w_dff_A_bByk705m9_1),.clk(gclk));
	jdff dff_A_GfZmk5934_1(.dout(w_dff_A_bByk705m9_1),.din(w_dff_A_GfZmk5934_1),.clk(gclk));
	jdff dff_A_3DGBthFm8_1(.dout(w_dff_A_GfZmk5934_1),.din(w_dff_A_3DGBthFm8_1),.clk(gclk));
	jdff dff_A_7nPDNg0F7_1(.dout(w_dff_A_3DGBthFm8_1),.din(w_dff_A_7nPDNg0F7_1),.clk(gclk));
	jdff dff_A_kzEOtdX72_1(.dout(w_dff_A_7nPDNg0F7_1),.din(w_dff_A_kzEOtdX72_1),.clk(gclk));
	jdff dff_A_CfeLAbC85_1(.dout(w_dff_A_kzEOtdX72_1),.din(w_dff_A_CfeLAbC85_1),.clk(gclk));
	jdff dff_A_AbLKmgaf6_1(.dout(w_dff_A_CfeLAbC85_1),.din(w_dff_A_AbLKmgaf6_1),.clk(gclk));
	jdff dff_A_juyqQyl61_1(.dout(w_dff_A_AbLKmgaf6_1),.din(w_dff_A_juyqQyl61_1),.clk(gclk));
	jdff dff_A_lPnI40po1_1(.dout(w_dff_A_juyqQyl61_1),.din(w_dff_A_lPnI40po1_1),.clk(gclk));
	jdff dff_A_a38Z7zQv2_1(.dout(w_dff_A_lPnI40po1_1),.din(w_dff_A_a38Z7zQv2_1),.clk(gclk));
	jdff dff_A_PVQH0J5H3_1(.dout(w_dff_A_a38Z7zQv2_1),.din(w_dff_A_PVQH0J5H3_1),.clk(gclk));
	jdff dff_A_vDD9AvLr0_1(.dout(w_dff_A_PVQH0J5H3_1),.din(w_dff_A_vDD9AvLr0_1),.clk(gclk));
	jdff dff_A_fxnYGVro0_1(.dout(w_dff_A_vDD9AvLr0_1),.din(w_dff_A_fxnYGVro0_1),.clk(gclk));
	jdff dff_A_55eL2Zly2_1(.dout(w_dff_A_fxnYGVro0_1),.din(w_dff_A_55eL2Zly2_1),.clk(gclk));
	jdff dff_A_2bvKdXBt2_1(.dout(w_dff_A_55eL2Zly2_1),.din(w_dff_A_2bvKdXBt2_1),.clk(gclk));
	jdff dff_A_yLxDTtHx7_1(.dout(w_dff_A_2bvKdXBt2_1),.din(w_dff_A_yLxDTtHx7_1),.clk(gclk));
	jdff dff_A_QDnuycIy2_2(.dout(w_n993_0[2]),.din(w_dff_A_QDnuycIy2_2),.clk(gclk));
	jdff dff_A_nVY3kyfG2_2(.dout(w_dff_A_QDnuycIy2_2),.din(w_dff_A_nVY3kyfG2_2),.clk(gclk));
	jdff dff_A_4uFGPOqR0_2(.dout(w_dff_A_nVY3kyfG2_2),.din(w_dff_A_4uFGPOqR0_2),.clk(gclk));
	jdff dff_A_qV0CoZK13_2(.dout(w_dff_A_4uFGPOqR0_2),.din(w_dff_A_qV0CoZK13_2),.clk(gclk));
	jdff dff_A_7ZCWIkBK5_2(.dout(w_dff_A_qV0CoZK13_2),.din(w_dff_A_7ZCWIkBK5_2),.clk(gclk));
	jdff dff_A_dXpnKGlN6_2(.dout(w_dff_A_7ZCWIkBK5_2),.din(w_dff_A_dXpnKGlN6_2),.clk(gclk));
	jdff dff_A_O3hIAkMv6_2(.dout(w_dff_A_dXpnKGlN6_2),.din(w_dff_A_O3hIAkMv6_2),.clk(gclk));
	jdff dff_A_XPplqGCX4_2(.dout(w_dff_A_O3hIAkMv6_2),.din(w_dff_A_XPplqGCX4_2),.clk(gclk));
	jdff dff_A_h47oQwxH6_2(.dout(w_dff_A_XPplqGCX4_2),.din(w_dff_A_h47oQwxH6_2),.clk(gclk));
	jdff dff_A_9MANMymo8_2(.dout(w_dff_A_h47oQwxH6_2),.din(w_dff_A_9MANMymo8_2),.clk(gclk));
	jdff dff_A_7HUVL1Pp0_2(.dout(w_dff_A_9MANMymo8_2),.din(w_dff_A_7HUVL1Pp0_2),.clk(gclk));
	jdff dff_A_7MZiC1pn7_1(.dout(w_G1690_1[1]),.din(w_dff_A_7MZiC1pn7_1),.clk(gclk));
	jdff dff_A_CozOhow45_1(.dout(w_G1690_0[1]),.din(w_dff_A_CozOhow45_1),.clk(gclk));
	jdff dff_A_KNoEf7Di6_1(.dout(w_dff_A_CozOhow45_1),.din(w_dff_A_KNoEf7Di6_1),.clk(gclk));
	jdff dff_A_iDD1DUjj3_1(.dout(w_dff_A_KNoEf7Di6_1),.din(w_dff_A_iDD1DUjj3_1),.clk(gclk));
	jdff dff_A_fJZFzTZc2_1(.dout(w_dff_A_iDD1DUjj3_1),.din(w_dff_A_fJZFzTZc2_1),.clk(gclk));
	jdff dff_A_svg15Zt01_1(.dout(w_dff_A_fJZFzTZc2_1),.din(w_dff_A_svg15Zt01_1),.clk(gclk));
	jdff dff_A_1IzpDqem3_1(.dout(w_dff_A_svg15Zt01_1),.din(w_dff_A_1IzpDqem3_1),.clk(gclk));
	jdff dff_A_OBV2Z7rV0_1(.dout(w_dff_A_1IzpDqem3_1),.din(w_dff_A_OBV2Z7rV0_1),.clk(gclk));
	jdff dff_A_LvLFPvna1_1(.dout(w_dff_A_OBV2Z7rV0_1),.din(w_dff_A_LvLFPvna1_1),.clk(gclk));
	jdff dff_A_XlGW3R8C5_1(.dout(w_dff_A_LvLFPvna1_1),.din(w_dff_A_XlGW3R8C5_1),.clk(gclk));
	jdff dff_A_Hr0t9hil2_1(.dout(w_dff_A_XlGW3R8C5_1),.din(w_dff_A_Hr0t9hil2_1),.clk(gclk));
	jdff dff_A_ycKLrXAJ5_1(.dout(w_dff_A_Hr0t9hil2_1),.din(w_dff_A_ycKLrXAJ5_1),.clk(gclk));
	jdff dff_A_4Xxacixz3_1(.dout(w_dff_A_ycKLrXAJ5_1),.din(w_dff_A_4Xxacixz3_1),.clk(gclk));
	jdff dff_A_PIjAaaZW0_1(.dout(w_dff_A_4Xxacixz3_1),.din(w_dff_A_PIjAaaZW0_1),.clk(gclk));
	jdff dff_A_57glIP3i7_1(.dout(w_dff_A_PIjAaaZW0_1),.din(w_dff_A_57glIP3i7_1),.clk(gclk));
	jdff dff_A_YxmSF84j0_1(.dout(w_dff_A_57glIP3i7_1),.din(w_dff_A_YxmSF84j0_1),.clk(gclk));
	jdff dff_A_jhMcZnbt2_1(.dout(w_dff_A_YxmSF84j0_1),.din(w_dff_A_jhMcZnbt2_1),.clk(gclk));
	jdff dff_A_DnaIkzaT3_1(.dout(w_dff_A_jhMcZnbt2_1),.din(w_dff_A_DnaIkzaT3_1),.clk(gclk));
	jdff dff_A_imHxDDda9_1(.dout(w_dff_A_DnaIkzaT3_1),.din(w_dff_A_imHxDDda9_1),.clk(gclk));
	jdff dff_A_6hVWXkjQ6_1(.dout(w_dff_A_imHxDDda9_1),.din(w_dff_A_6hVWXkjQ6_1),.clk(gclk));
	jdff dff_A_xTtnHCis9_1(.dout(w_dff_A_6hVWXkjQ6_1),.din(w_dff_A_xTtnHCis9_1),.clk(gclk));
	jdff dff_A_DKnsmow48_1(.dout(w_dff_A_xTtnHCis9_1),.din(w_dff_A_DKnsmow48_1),.clk(gclk));
	jdff dff_A_vfyF6Ycp1_1(.dout(w_dff_A_DKnsmow48_1),.din(w_dff_A_vfyF6Ycp1_1),.clk(gclk));
	jdff dff_A_WFpyXQE98_1(.dout(w_dff_A_vfyF6Ycp1_1),.din(w_dff_A_WFpyXQE98_1),.clk(gclk));
	jdff dff_A_aMDjTctL1_0(.dout(w_G1689_1[0]),.din(w_dff_A_aMDjTctL1_0),.clk(gclk));
	jdff dff_A_BwJs6p1G3_0(.dout(w_dff_A_aMDjTctL1_0),.din(w_dff_A_BwJs6p1G3_0),.clk(gclk));
	jdff dff_A_zbC3LCll8_0(.dout(w_dff_A_BwJs6p1G3_0),.din(w_dff_A_zbC3LCll8_0),.clk(gclk));
	jdff dff_A_ejgauGLC4_0(.dout(w_dff_A_zbC3LCll8_0),.din(w_dff_A_ejgauGLC4_0),.clk(gclk));
	jdff dff_A_Kw3svK8O4_0(.dout(w_dff_A_ejgauGLC4_0),.din(w_dff_A_Kw3svK8O4_0),.clk(gclk));
	jdff dff_A_mEdP1J3l8_0(.dout(w_dff_A_Kw3svK8O4_0),.din(w_dff_A_mEdP1J3l8_0),.clk(gclk));
	jdff dff_A_IfJ6Ji1l7_0(.dout(w_dff_A_mEdP1J3l8_0),.din(w_dff_A_IfJ6Ji1l7_0),.clk(gclk));
	jdff dff_A_0FwZ7po26_0(.dout(w_dff_A_IfJ6Ji1l7_0),.din(w_dff_A_0FwZ7po26_0),.clk(gclk));
	jdff dff_A_SXzeJC4S4_0(.dout(w_dff_A_0FwZ7po26_0),.din(w_dff_A_SXzeJC4S4_0),.clk(gclk));
	jdff dff_A_mDWta6TW9_2(.dout(w_G1689_1[2]),.din(w_dff_A_mDWta6TW9_2),.clk(gclk));
	jdff dff_A_hHzCmzeS4_2(.dout(w_dff_A_mDWta6TW9_2),.din(w_dff_A_hHzCmzeS4_2),.clk(gclk));
	jdff dff_A_TtGEkeY89_2(.dout(w_dff_A_hHzCmzeS4_2),.din(w_dff_A_TtGEkeY89_2),.clk(gclk));
	jdff dff_A_K1x60O0N4_2(.dout(w_dff_A_TtGEkeY89_2),.din(w_dff_A_K1x60O0N4_2),.clk(gclk));
	jdff dff_A_Uarh9PFV1_2(.dout(w_dff_A_K1x60O0N4_2),.din(w_dff_A_Uarh9PFV1_2),.clk(gclk));
	jdff dff_A_gj7lFmNP8_2(.dout(w_dff_A_Uarh9PFV1_2),.din(w_dff_A_gj7lFmNP8_2),.clk(gclk));
	jdff dff_A_RwD8JSBg5_2(.dout(w_dff_A_gj7lFmNP8_2),.din(w_dff_A_RwD8JSBg5_2),.clk(gclk));
	jdff dff_A_wT8289un0_2(.dout(w_dff_A_RwD8JSBg5_2),.din(w_dff_A_wT8289un0_2),.clk(gclk));
	jdff dff_A_Xr0Kvv8Y5_2(.dout(w_dff_A_wT8289un0_2),.din(w_dff_A_Xr0Kvv8Y5_2),.clk(gclk));
	jdff dff_A_OP52JwfC9_2(.dout(w_dff_A_Xr0Kvv8Y5_2),.din(w_dff_A_OP52JwfC9_2),.clk(gclk));
	jdff dff_A_Y6gUf3oU0_2(.dout(w_dff_A_OP52JwfC9_2),.din(w_dff_A_Y6gUf3oU0_2),.clk(gclk));
	jdff dff_A_9AAW29E89_2(.dout(w_dff_A_Y6gUf3oU0_2),.din(w_dff_A_9AAW29E89_2),.clk(gclk));
	jdff dff_A_6P32KFym1_2(.dout(w_dff_A_9AAW29E89_2),.din(w_dff_A_6P32KFym1_2),.clk(gclk));
	jdff dff_A_3TKcNZZK1_2(.dout(w_dff_A_6P32KFym1_2),.din(w_dff_A_3TKcNZZK1_2),.clk(gclk));
	jdff dff_A_D8gzYsni2_2(.dout(w_dff_A_3TKcNZZK1_2),.din(w_dff_A_D8gzYsni2_2),.clk(gclk));
	jdff dff_A_8ITYveoI6_2(.dout(w_dff_A_D8gzYsni2_2),.din(w_dff_A_8ITYveoI6_2),.clk(gclk));
	jdff dff_A_2D84yOlR5_2(.dout(w_dff_A_8ITYveoI6_2),.din(w_dff_A_2D84yOlR5_2),.clk(gclk));
	jdff dff_A_wc0xcGdp5_2(.dout(w_dff_A_2D84yOlR5_2),.din(w_dff_A_wc0xcGdp5_2),.clk(gclk));
	jdff dff_A_MJEHKelT9_2(.dout(w_dff_A_wc0xcGdp5_2),.din(w_dff_A_MJEHKelT9_2),.clk(gclk));
	jdff dff_A_TpLGOVxJ3_2(.dout(w_dff_A_MJEHKelT9_2),.din(w_dff_A_TpLGOVxJ3_2),.clk(gclk));
	jdff dff_A_Sn4d4rc53_2(.dout(w_dff_A_TpLGOVxJ3_2),.din(w_dff_A_Sn4d4rc53_2),.clk(gclk));
	jdff dff_A_KG0OdvOF6_2(.dout(w_dff_A_Sn4d4rc53_2),.din(w_dff_A_KG0OdvOF6_2),.clk(gclk));
	jdff dff_A_kxet5FjL6_1(.dout(w_G1689_0[1]),.din(w_dff_A_kxet5FjL6_1),.clk(gclk));
	jdff dff_A_o5CGr2Xd1_1(.dout(w_dff_A_kxet5FjL6_1),.din(w_dff_A_o5CGr2Xd1_1),.clk(gclk));
	jdff dff_A_3Pv0tZvA9_1(.dout(w_dff_A_o5CGr2Xd1_1),.din(w_dff_A_3Pv0tZvA9_1),.clk(gclk));
	jdff dff_A_Luggkojh2_1(.dout(w_dff_A_3Pv0tZvA9_1),.din(w_dff_A_Luggkojh2_1),.clk(gclk));
	jdff dff_A_bNAwkg675_1(.dout(w_dff_A_Luggkojh2_1),.din(w_dff_A_bNAwkg675_1),.clk(gclk));
	jdff dff_A_EU1Dvvx85_1(.dout(w_dff_A_bNAwkg675_1),.din(w_dff_A_EU1Dvvx85_1),.clk(gclk));
	jdff dff_A_VNq02SJX2_1(.dout(w_dff_A_EU1Dvvx85_1),.din(w_dff_A_VNq02SJX2_1),.clk(gclk));
	jdff dff_A_0403zIP21_1(.dout(w_dff_A_VNq02SJX2_1),.din(w_dff_A_0403zIP21_1),.clk(gclk));
	jdff dff_A_7vdJej4w7_1(.dout(w_dff_A_0403zIP21_1),.din(w_dff_A_7vdJej4w7_1),.clk(gclk));
	jdff dff_A_ILyRnmIo6_1(.dout(w_dff_A_7vdJej4w7_1),.din(w_dff_A_ILyRnmIo6_1),.clk(gclk));
	jdff dff_A_1FParwAR7_1(.dout(w_dff_A_ILyRnmIo6_1),.din(w_dff_A_1FParwAR7_1),.clk(gclk));
	jdff dff_A_MxY3InuG6_1(.dout(w_dff_A_1FParwAR7_1),.din(w_dff_A_MxY3InuG6_1),.clk(gclk));
	jdff dff_A_MjDO53oV9_1(.dout(w_dff_A_MxY3InuG6_1),.din(w_dff_A_MjDO53oV9_1),.clk(gclk));
	jdff dff_A_TzqSrlq20_1(.dout(w_dff_A_MjDO53oV9_1),.din(w_dff_A_TzqSrlq20_1),.clk(gclk));
	jdff dff_A_6gXZQCVX2_1(.dout(w_dff_A_TzqSrlq20_1),.din(w_dff_A_6gXZQCVX2_1),.clk(gclk));
	jdff dff_A_8kdbvXo36_1(.dout(w_dff_A_6gXZQCVX2_1),.din(w_dff_A_8kdbvXo36_1),.clk(gclk));
	jdff dff_A_rBj5yH7m2_1(.dout(w_dff_A_8kdbvXo36_1),.din(w_dff_A_rBj5yH7m2_1),.clk(gclk));
	jdff dff_A_c2wt0MIR8_1(.dout(w_dff_A_rBj5yH7m2_1),.din(w_dff_A_c2wt0MIR8_1),.clk(gclk));
	jdff dff_A_71Hv8wWq6_1(.dout(w_dff_A_c2wt0MIR8_1),.din(w_dff_A_71Hv8wWq6_1),.clk(gclk));
	jdff dff_A_PgFreHKh6_2(.dout(w_G1689_0[2]),.din(w_dff_A_PgFreHKh6_2),.clk(gclk));
	jdff dff_A_xafjBsPZ9_2(.dout(w_dff_A_PgFreHKh6_2),.din(w_dff_A_xafjBsPZ9_2),.clk(gclk));
	jdff dff_A_CQU9iPEY5_2(.dout(w_dff_A_xafjBsPZ9_2),.din(w_dff_A_CQU9iPEY5_2),.clk(gclk));
	jdff dff_A_DbsFcYV09_2(.dout(w_dff_A_CQU9iPEY5_2),.din(w_dff_A_DbsFcYV09_2),.clk(gclk));
	jdff dff_A_qiPvhrsf0_2(.dout(w_dff_A_DbsFcYV09_2),.din(w_dff_A_qiPvhrsf0_2),.clk(gclk));
	jdff dff_A_LUvOHpZi3_2(.dout(w_dff_A_qiPvhrsf0_2),.din(w_dff_A_LUvOHpZi3_2),.clk(gclk));
	jdff dff_A_OlIIpLag3_2(.dout(w_dff_A_LUvOHpZi3_2),.din(w_dff_A_OlIIpLag3_2),.clk(gclk));
	jdff dff_A_EHiiTA7u0_2(.dout(w_dff_A_OlIIpLag3_2),.din(w_dff_A_EHiiTA7u0_2),.clk(gclk));
	jdff dff_A_hgA0ILHc4_2(.dout(w_dff_A_EHiiTA7u0_2),.din(w_dff_A_hgA0ILHc4_2),.clk(gclk));
	jdff dff_A_y04p6kf26_2(.dout(w_dff_A_hgA0ILHc4_2),.din(w_dff_A_y04p6kf26_2),.clk(gclk));
	jdff dff_A_2D4206v07_2(.dout(w_dff_A_y04p6kf26_2),.din(w_dff_A_2D4206v07_2),.clk(gclk));
	jdff dff_A_Pfca8OpW5_2(.dout(w_dff_A_2D4206v07_2),.din(w_dff_A_Pfca8OpW5_2),.clk(gclk));
	jdff dff_A_MHwIKS9y3_2(.dout(w_dff_A_Pfca8OpW5_2),.din(w_dff_A_MHwIKS9y3_2),.clk(gclk));
	jdff dff_B_GcMdmMVM2_1(.din(n1709),.dout(w_dff_B_GcMdmMVM2_1),.clk(gclk));
	jdff dff_B_zMZMUDlf5_1(.din(w_dff_B_GcMdmMVM2_1),.dout(w_dff_B_zMZMUDlf5_1),.clk(gclk));
	jdff dff_B_RhyuXJLF6_1(.din(w_dff_B_zMZMUDlf5_1),.dout(w_dff_B_RhyuXJLF6_1),.clk(gclk));
	jdff dff_B_WGARJiUp5_1(.din(w_dff_B_RhyuXJLF6_1),.dout(w_dff_B_WGARJiUp5_1),.clk(gclk));
	jdff dff_B_BvxJ2Mm64_1(.din(w_dff_B_WGARJiUp5_1),.dout(w_dff_B_BvxJ2Mm64_1),.clk(gclk));
	jdff dff_B_pLeBhFNz9_1(.din(w_dff_B_BvxJ2Mm64_1),.dout(w_dff_B_pLeBhFNz9_1),.clk(gclk));
	jdff dff_B_nqh3MVxB1_1(.din(w_dff_B_pLeBhFNz9_1),.dout(w_dff_B_nqh3MVxB1_1),.clk(gclk));
	jdff dff_B_dV5BTFhk1_1(.din(w_dff_B_nqh3MVxB1_1),.dout(w_dff_B_dV5BTFhk1_1),.clk(gclk));
	jdff dff_B_P2lTB8rS3_1(.din(w_dff_B_dV5BTFhk1_1),.dout(w_dff_B_P2lTB8rS3_1),.clk(gclk));
	jdff dff_B_s9tCs7Ub1_1(.din(w_dff_B_P2lTB8rS3_1),.dout(w_dff_B_s9tCs7Ub1_1),.clk(gclk));
	jdff dff_B_3Y0mdJ9U4_1(.din(w_dff_B_s9tCs7Ub1_1),.dout(w_dff_B_3Y0mdJ9U4_1),.clk(gclk));
	jdff dff_B_0eWqvDC76_1(.din(w_dff_B_3Y0mdJ9U4_1),.dout(w_dff_B_0eWqvDC76_1),.clk(gclk));
	jdff dff_B_0vl2vCaa8_1(.din(w_dff_B_0eWqvDC76_1),.dout(w_dff_B_0vl2vCaa8_1),.clk(gclk));
	jdff dff_B_lPlH5lt62_1(.din(w_dff_B_0vl2vCaa8_1),.dout(w_dff_B_lPlH5lt62_1),.clk(gclk));
	jdff dff_B_unJ015bL8_1(.din(w_dff_B_lPlH5lt62_1),.dout(w_dff_B_unJ015bL8_1),.clk(gclk));
	jdff dff_B_O2eDBG042_1(.din(w_dff_B_unJ015bL8_1),.dout(w_dff_B_O2eDBG042_1),.clk(gclk));
	jdff dff_B_BCbxBWk33_1(.din(w_dff_B_O2eDBG042_1),.dout(w_dff_B_BCbxBWk33_1),.clk(gclk));
	jdff dff_B_nUzOZrMs5_1(.din(w_dff_B_BCbxBWk33_1),.dout(w_dff_B_nUzOZrMs5_1),.clk(gclk));
	jdff dff_B_nPxXPHIc5_1(.din(w_dff_B_nUzOZrMs5_1),.dout(w_dff_B_nPxXPHIc5_1),.clk(gclk));
	jdff dff_B_YTIhUTTB4_1(.din(w_dff_B_nPxXPHIc5_1),.dout(w_dff_B_YTIhUTTB4_1),.clk(gclk));
	jdff dff_B_NOp2b5xe5_1(.din(w_dff_B_YTIhUTTB4_1),.dout(w_dff_B_NOp2b5xe5_1),.clk(gclk));
	jdff dff_B_OMqhVrpM7_1(.din(w_dff_B_NOp2b5xe5_1),.dout(w_dff_B_OMqhVrpM7_1),.clk(gclk));
	jdff dff_B_xIkb5FXp4_1(.din(w_dff_B_OMqhVrpM7_1),.dout(w_dff_B_xIkb5FXp4_1),.clk(gclk));
	jdff dff_B_B6rP9bDy7_1(.din(n1711),.dout(w_dff_B_B6rP9bDy7_1),.clk(gclk));
	jdff dff_B_JVohYFZe8_1(.din(w_dff_B_B6rP9bDy7_1),.dout(w_dff_B_JVohYFZe8_1),.clk(gclk));
	jdff dff_B_XL1w188B3_1(.din(w_dff_B_JVohYFZe8_1),.dout(w_dff_B_XL1w188B3_1),.clk(gclk));
	jdff dff_B_T7AklfjQ6_1(.din(w_dff_B_XL1w188B3_1),.dout(w_dff_B_T7AklfjQ6_1),.clk(gclk));
	jdff dff_B_N8Qk7xNi3_1(.din(w_dff_B_T7AklfjQ6_1),.dout(w_dff_B_N8Qk7xNi3_1),.clk(gclk));
	jdff dff_B_0EcG2cvJ4_1(.din(w_dff_B_N8Qk7xNi3_1),.dout(w_dff_B_0EcG2cvJ4_1),.clk(gclk));
	jdff dff_B_ng0t5frc6_1(.din(w_dff_B_0EcG2cvJ4_1),.dout(w_dff_B_ng0t5frc6_1),.clk(gclk));
	jdff dff_B_FXUugAvv8_1(.din(w_dff_B_ng0t5frc6_1),.dout(w_dff_B_FXUugAvv8_1),.clk(gclk));
	jdff dff_B_Bt6acUxp3_1(.din(w_dff_B_FXUugAvv8_1),.dout(w_dff_B_Bt6acUxp3_1),.clk(gclk));
	jdff dff_B_Iv9TBwiM1_1(.din(w_dff_B_Bt6acUxp3_1),.dout(w_dff_B_Iv9TBwiM1_1),.clk(gclk));
	jdff dff_B_R82TuCAp8_1(.din(w_dff_B_Iv9TBwiM1_1),.dout(w_dff_B_R82TuCAp8_1),.clk(gclk));
	jdff dff_B_jFKLyiBR8_1(.din(w_dff_B_R82TuCAp8_1),.dout(w_dff_B_jFKLyiBR8_1),.clk(gclk));
	jdff dff_B_r52Jz6kg4_1(.din(w_dff_B_jFKLyiBR8_1),.dout(w_dff_B_r52Jz6kg4_1),.clk(gclk));
	jdff dff_B_6CDC7SuT2_1(.din(w_dff_B_r52Jz6kg4_1),.dout(w_dff_B_6CDC7SuT2_1),.clk(gclk));
	jdff dff_B_GNiAnel13_1(.din(w_dff_B_6CDC7SuT2_1),.dout(w_dff_B_GNiAnel13_1),.clk(gclk));
	jdff dff_B_bH3FXHlC6_1(.din(w_dff_B_GNiAnel13_1),.dout(w_dff_B_bH3FXHlC6_1),.clk(gclk));
	jdff dff_B_FOs56RDq4_1(.din(w_dff_B_bH3FXHlC6_1),.dout(w_dff_B_FOs56RDq4_1),.clk(gclk));
	jdff dff_B_W4xFd2Mv8_1(.din(w_dff_B_FOs56RDq4_1),.dout(w_dff_B_W4xFd2Mv8_1),.clk(gclk));
	jdff dff_B_DWwOLS1p7_1(.din(w_dff_B_W4xFd2Mv8_1),.dout(w_dff_B_DWwOLS1p7_1),.clk(gclk));
	jdff dff_B_tB2tv4WR3_1(.din(w_dff_B_DWwOLS1p7_1),.dout(w_dff_B_tB2tv4WR3_1),.clk(gclk));
	jdff dff_B_ccUhAJav5_1(.din(w_dff_B_tB2tv4WR3_1),.dout(w_dff_B_ccUhAJav5_1),.clk(gclk));
	jdff dff_B_MI2lEjEz8_1(.din(n1712),.dout(w_dff_B_MI2lEjEz8_1),.clk(gclk));
	jdff dff_B_CpST3Fer2_0(.din(n1678),.dout(w_dff_B_CpST3Fer2_0),.clk(gclk));
	jdff dff_B_LxWmpUSM6_0(.din(w_dff_B_CpST3Fer2_0),.dout(w_dff_B_LxWmpUSM6_0),.clk(gclk));
	jdff dff_B_pZcb0Kqh3_0(.din(w_dff_B_LxWmpUSM6_0),.dout(w_dff_B_pZcb0Kqh3_0),.clk(gclk));
	jdff dff_B_q5nww98O8_0(.din(w_dff_B_pZcb0Kqh3_0),.dout(w_dff_B_q5nww98O8_0),.clk(gclk));
	jdff dff_B_vqc6fzrr5_0(.din(w_dff_B_q5nww98O8_0),.dout(w_dff_B_vqc6fzrr5_0),.clk(gclk));
	jdff dff_B_OeVZYOW70_0(.din(w_dff_B_vqc6fzrr5_0),.dout(w_dff_B_OeVZYOW70_0),.clk(gclk));
	jdff dff_B_SdjibiUX6_0(.din(w_dff_B_OeVZYOW70_0),.dout(w_dff_B_SdjibiUX6_0),.clk(gclk));
	jdff dff_B_iqEsNM4v1_0(.din(w_dff_B_SdjibiUX6_0),.dout(w_dff_B_iqEsNM4v1_0),.clk(gclk));
	jdff dff_B_MTRkLikJ2_0(.din(w_dff_B_iqEsNM4v1_0),.dout(w_dff_B_MTRkLikJ2_0),.clk(gclk));
	jdff dff_B_ofABOZhb3_0(.din(w_dff_B_MTRkLikJ2_0),.dout(w_dff_B_ofABOZhb3_0),.clk(gclk));
	jdff dff_B_fvXc74ma0_0(.din(w_dff_B_ofABOZhb3_0),.dout(w_dff_B_fvXc74ma0_0),.clk(gclk));
	jdff dff_B_AQRQ9Uxa9_0(.din(w_dff_B_fvXc74ma0_0),.dout(w_dff_B_AQRQ9Uxa9_0),.clk(gclk));
	jdff dff_B_HGhr1ADv1_0(.din(w_dff_B_AQRQ9Uxa9_0),.dout(w_dff_B_HGhr1ADv1_0),.clk(gclk));
	jdff dff_B_MGkbql5G1_0(.din(w_dff_B_HGhr1ADv1_0),.dout(w_dff_B_MGkbql5G1_0),.clk(gclk));
	jdff dff_B_mN4fDTrq4_0(.din(w_dff_B_MGkbql5G1_0),.dout(w_dff_B_mN4fDTrq4_0),.clk(gclk));
	jdff dff_B_Azu6K8Sc3_0(.din(w_dff_B_mN4fDTrq4_0),.dout(w_dff_B_Azu6K8Sc3_0),.clk(gclk));
	jdff dff_B_7pOQs7l51_0(.din(w_dff_B_Azu6K8Sc3_0),.dout(w_dff_B_7pOQs7l51_0),.clk(gclk));
	jdff dff_B_GpEUyCfx2_0(.din(w_dff_B_7pOQs7l51_0),.dout(w_dff_B_GpEUyCfx2_0),.clk(gclk));
	jdff dff_B_g7SLLSYW6_0(.din(w_dff_B_GpEUyCfx2_0),.dout(w_dff_B_g7SLLSYW6_0),.clk(gclk));
	jdff dff_B_eSIga0pe3_0(.din(n1501),.dout(w_dff_B_eSIga0pe3_0),.clk(gclk));
	jdff dff_B_IrUnlNG80_0(.din(w_dff_B_eSIga0pe3_0),.dout(w_dff_B_IrUnlNG80_0),.clk(gclk));
	jdff dff_B_gMDbBuhw1_0(.din(w_dff_B_IrUnlNG80_0),.dout(w_dff_B_gMDbBuhw1_0),.clk(gclk));
	jdff dff_B_eDYGrcpj3_0(.din(w_dff_B_gMDbBuhw1_0),.dout(w_dff_B_eDYGrcpj3_0),.clk(gclk));
	jdff dff_B_ryH6SxkN9_0(.din(w_dff_B_eDYGrcpj3_0),.dout(w_dff_B_ryH6SxkN9_0),.clk(gclk));
	jdff dff_B_r5rBMJ1U1_0(.din(w_dff_B_ryH6SxkN9_0),.dout(w_dff_B_r5rBMJ1U1_0),.clk(gclk));
	jdff dff_B_oL51l6mP4_0(.din(w_dff_B_r5rBMJ1U1_0),.dout(w_dff_B_oL51l6mP4_0),.clk(gclk));
	jdff dff_B_wySAC3OF1_0(.din(w_dff_B_oL51l6mP4_0),.dout(w_dff_B_wySAC3OF1_0),.clk(gclk));
	jdff dff_B_Z6XkuS7b3_0(.din(w_dff_B_wySAC3OF1_0),.dout(w_dff_B_Z6XkuS7b3_0),.clk(gclk));
	jdff dff_B_zU9xVylp3_1(.din(n1496),.dout(w_dff_B_zU9xVylp3_1),.clk(gclk));
	jdff dff_B_3bQpT2b02_1(.din(n413),.dout(w_dff_B_3bQpT2b02_1),.clk(gclk));
	jdff dff_B_h6IJkdMG1_1(.din(w_dff_B_3bQpT2b02_1),.dout(w_dff_B_h6IJkdMG1_1),.clk(gclk));
	jdff dff_A_cCAn80oG9_0(.dout(w_G308_1[0]),.din(w_dff_A_cCAn80oG9_0),.clk(gclk));
	jdff dff_B_wFu7iZoY4_1(.din(n400),.dout(w_dff_B_wFu7iZoY4_1),.clk(gclk));
	jdff dff_B_fbBXViZA9_1(.din(w_dff_B_wFu7iZoY4_1),.dout(w_dff_B_fbBXViZA9_1),.clk(gclk));
	jdff dff_A_H8tCWae42_1(.dout(w_n428_0[1]),.din(w_dff_A_H8tCWae42_1),.clk(gclk));
	jdff dff_B_JZ7huyEY5_0(.din(n1493),.dout(w_dff_B_JZ7huyEY5_0),.clk(gclk));
	jdff dff_A_iuRPSOYI0_0(.dout(w_G361_1[0]),.din(w_dff_A_iuRPSOYI0_0),.clk(gclk));
	jdff dff_B_29o6Iq4y3_1(.din(n1485),.dout(w_dff_B_29o6Iq4y3_1),.clk(gclk));
	jdff dff_A_Unoy0Uw58_0(.dout(w_n437_0[0]),.din(w_dff_A_Unoy0Uw58_0),.clk(gclk));
	jdff dff_B_FbiuPYQL1_2(.din(n437),.dout(w_dff_B_FbiuPYQL1_2),.clk(gclk));
	jdff dff_A_N3JHm29S7_0(.dout(w_G503_2[0]),.din(w_dff_A_N3JHm29S7_0),.clk(gclk));
	jdff dff_A_GPJO0iP97_0(.dout(w_dff_A_N3JHm29S7_0),.din(w_dff_A_GPJO0iP97_0),.clk(gclk));
	jdff dff_A_c0cF66of2_0(.dout(w_dff_A_GPJO0iP97_0),.din(w_dff_A_c0cF66of2_0),.clk(gclk));
	jdff dff_B_KuVIetra4_1(.din(n1481),.dout(w_dff_B_KuVIetra4_1),.clk(gclk));
	jdff dff_B_OkaoFZ6D5_1(.din(n1471),.dout(w_dff_B_OkaoFZ6D5_1),.clk(gclk));
	jdff dff_B_qItMzJlr6_1(.din(w_dff_B_OkaoFZ6D5_1),.dout(w_dff_B_qItMzJlr6_1),.clk(gclk));
	jdff dff_A_XoUV0c5b2_1(.dout(w_G341_2[1]),.din(w_dff_A_XoUV0c5b2_1),.clk(gclk));
	jdff dff_B_U9CtPUDe4_1(.din(n1462),.dout(w_dff_B_U9CtPUDe4_1),.clk(gclk));
	jdff dff_B_eFO82afY2_1(.din(w_dff_B_U9CtPUDe4_1),.dout(w_dff_B_eFO82afY2_1),.clk(gclk));
	jdff dff_A_3iL9ABnu6_1(.dout(w_G351_2[1]),.din(w_dff_A_3iL9ABnu6_1),.clk(gclk));
	jdff dff_B_nmS8vhuX1_1(.din(n1453),.dout(w_dff_B_nmS8vhuX1_1),.clk(gclk));
	jdff dff_A_pcFGW0Pn6_0(.dout(w_n749_5[0]),.din(w_dff_A_pcFGW0Pn6_0),.clk(gclk));
	jdff dff_A_Laqa2d835_0(.dout(w_dff_A_pcFGW0Pn6_0),.din(w_dff_A_Laqa2d835_0),.clk(gclk));
	jdff dff_A_2mXuuQ4Y2_0(.dout(w_dff_A_Laqa2d835_0),.din(w_dff_A_2mXuuQ4Y2_0),.clk(gclk));
	jdff dff_A_2g984dOy4_1(.dout(w_n749_5[1]),.din(w_dff_A_2g984dOy4_1),.clk(gclk));
	jdff dff_A_ufLtg2qa8_1(.dout(w_dff_A_2g984dOy4_1),.din(w_dff_A_ufLtg2qa8_1),.clk(gclk));
	jdff dff_A_9GU07UWk6_1(.dout(w_dff_A_ufLtg2qa8_1),.din(w_dff_A_9GU07UWk6_1),.clk(gclk));
	jdff dff_A_vrKrY8cu5_1(.dout(w_dff_A_9GU07UWk6_1),.din(w_dff_A_vrKrY8cu5_1),.clk(gclk));
	jdff dff_A_i6YE0F3L3_1(.dout(w_dff_A_vrKrY8cu5_1),.din(w_dff_A_i6YE0F3L3_1),.clk(gclk));
	jdff dff_A_G2mtEQOr2_1(.dout(w_dff_A_i6YE0F3L3_1),.din(w_dff_A_G2mtEQOr2_1),.clk(gclk));
	jdff dff_A_U2mXfd1S2_1(.dout(w_dff_A_G2mtEQOr2_1),.din(w_dff_A_U2mXfd1S2_1),.clk(gclk));
	jdff dff_A_8fGymNBb2_1(.dout(w_dff_A_U2mXfd1S2_1),.din(w_dff_A_8fGymNBb2_1),.clk(gclk));
	jdff dff_A_ECjd5M5B9_1(.dout(w_dff_A_8fGymNBb2_1),.din(w_dff_A_ECjd5M5B9_1),.clk(gclk));
	jdff dff_A_Q38jjBbW6_1(.dout(w_dff_A_ECjd5M5B9_1),.din(w_dff_A_Q38jjBbW6_1),.clk(gclk));
	jdff dff_A_8i6JpYol0_1(.dout(w_dff_A_Q38jjBbW6_1),.din(w_dff_A_8i6JpYol0_1),.clk(gclk));
	jdff dff_A_0Z3Tn8FY6_1(.dout(w_dff_A_8i6JpYol0_1),.din(w_dff_A_0Z3Tn8FY6_1),.clk(gclk));
	jdff dff_B_oJvbEFDl0_0(.din(n1452),.dout(w_dff_B_oJvbEFDl0_0),.clk(gclk));
	jdff dff_A_JPKQlNbV4_0(.dout(w_n1451_0[0]),.din(w_dff_A_JPKQlNbV4_0),.clk(gclk));
	jdff dff_A_ABbQpe6u2_0(.dout(w_dff_A_JPKQlNbV4_0),.din(w_dff_A_ABbQpe6u2_0),.clk(gclk));
	jdff dff_B_6FG4Q1yi3_0(.din(n1450),.dout(w_dff_B_6FG4Q1yi3_0),.clk(gclk));
	jdff dff_B_6rVycu836_0(.din(w_dff_B_6FG4Q1yi3_0),.dout(w_dff_B_6rVycu836_0),.clk(gclk));
	jdff dff_B_YUJFSNRH8_0(.din(w_dff_B_6rVycu836_0),.dout(w_dff_B_YUJFSNRH8_0),.clk(gclk));
	jdff dff_B_IsU0fbo28_1(.din(n1448),.dout(w_dff_B_IsU0fbo28_1),.clk(gclk));
	jdff dff_B_jVmOc66Q0_1(.din(w_dff_B_IsU0fbo28_1),.dout(w_dff_B_jVmOc66Q0_1),.clk(gclk));
	jdff dff_B_rQR8s6aN8_1(.din(w_dff_B_jVmOc66Q0_1),.dout(w_dff_B_rQR8s6aN8_1),.clk(gclk));
	jdff dff_A_N6FBxErh3_0(.dout(w_n763_0[0]),.din(w_dff_A_N6FBxErh3_0),.clk(gclk));
	jdff dff_A_khXuzogl9_0(.dout(w_dff_A_N6FBxErh3_0),.din(w_dff_A_khXuzogl9_0),.clk(gclk));
	jdff dff_A_c21A9dki1_0(.dout(w_dff_A_khXuzogl9_0),.din(w_dff_A_c21A9dki1_0),.clk(gclk));
	jdff dff_A_5Foc6wzG5_0(.dout(w_dff_A_c21A9dki1_0),.din(w_dff_A_5Foc6wzG5_0),.clk(gclk));
	jdff dff_A_srcgfnHl6_0(.dout(w_dff_A_5Foc6wzG5_0),.din(w_dff_A_srcgfnHl6_0),.clk(gclk));
	jdff dff_A_cpKxORtp9_0(.dout(w_dff_A_srcgfnHl6_0),.din(w_dff_A_cpKxORtp9_0),.clk(gclk));
	jdff dff_A_9PnZh8QN7_0(.dout(w_dff_A_cpKxORtp9_0),.din(w_dff_A_9PnZh8QN7_0),.clk(gclk));
	jdff dff_A_pxtAKnMq3_0(.dout(w_dff_A_9PnZh8QN7_0),.din(w_dff_A_pxtAKnMq3_0),.clk(gclk));
	jdff dff_B_Pwwn9wzk7_1(.din(n1439),.dout(w_dff_B_Pwwn9wzk7_1),.clk(gclk));
	jdff dff_B_GQA8Bv4Z2_1(.din(n1441),.dout(w_dff_B_GQA8Bv4Z2_1),.clk(gclk));
	jdff dff_B_68DvjMJx9_0(.din(n1437),.dout(w_dff_B_68DvjMJx9_0),.clk(gclk));
	jdff dff_B_94lpjmqD7_0(.din(n1436),.dout(w_dff_B_94lpjmqD7_0),.clk(gclk));
	jdff dff_A_4tImIQIC6_0(.dout(w_n1429_0[0]),.din(w_dff_A_4tImIQIC6_0),.clk(gclk));
	jdff dff_B_ZdQHdSHF7_1(.din(n1427),.dout(w_dff_B_ZdQHdSHF7_1),.clk(gclk));
	jdff dff_A_rJLsUqjl8_2(.dout(w_n641_0[2]),.din(w_dff_A_rJLsUqjl8_2),.clk(gclk));
	jdff dff_A_ZBOaviyN3_2(.dout(w_dff_A_rJLsUqjl8_2),.din(w_dff_A_ZBOaviyN3_2),.clk(gclk));
	jdff dff_A_ZlM4TwFe9_0(.dout(w_n640_0[0]),.din(w_dff_A_ZlM4TwFe9_0),.clk(gclk));
	jdff dff_A_9qjiZtE58_0(.dout(w_n639_0[0]),.din(w_dff_A_9qjiZtE58_0),.clk(gclk));
	jdff dff_A_0UXFHcve6_0(.dout(w_n624_0[0]),.din(w_dff_A_0UXFHcve6_0),.clk(gclk));
	jdff dff_A_UsjWnzyx7_0(.dout(w_dff_A_0UXFHcve6_0),.din(w_dff_A_UsjWnzyx7_0),.clk(gclk));
	jdff dff_A_Zmwi3UTf3_1(.dout(w_n624_0[1]),.din(w_dff_A_Zmwi3UTf3_1),.clk(gclk));
	jdff dff_B_YcEiYVfb1_3(.din(n624),.dout(w_dff_B_YcEiYVfb1_3),.clk(gclk));
	jdff dff_B_4iQ1YXwM3_3(.din(w_dff_B_YcEiYVfb1_3),.dout(w_dff_B_4iQ1YXwM3_3),.clk(gclk));
	jdff dff_A_CMqfPapT7_1(.dout(w_n620_1[1]),.din(w_dff_A_CMqfPapT7_1),.clk(gclk));
	jdff dff_A_9olhZSYh5_1(.dout(w_dff_A_CMqfPapT7_1),.din(w_dff_A_9olhZSYh5_1),.clk(gclk));
	jdff dff_A_fr8kjHLB5_1(.dout(w_dff_A_9olhZSYh5_1),.din(w_dff_A_fr8kjHLB5_1),.clk(gclk));
	jdff dff_A_QSN4LlY07_1(.dout(w_dff_A_fr8kjHLB5_1),.din(w_dff_A_QSN4LlY07_1),.clk(gclk));
	jdff dff_A_UsqvMGoB4_1(.dout(w_n620_0[1]),.din(w_dff_A_UsqvMGoB4_1),.clk(gclk));
	jdff dff_A_NKahmuzI0_1(.dout(w_dff_A_UsqvMGoB4_1),.din(w_dff_A_NKahmuzI0_1),.clk(gclk));
	jdff dff_A_qWlyI1sH6_2(.dout(w_n620_0[2]),.din(w_dff_A_qWlyI1sH6_2),.clk(gclk));
	jdff dff_A_mGAL2BkJ7_2(.dout(w_dff_A_qWlyI1sH6_2),.din(w_dff_A_mGAL2BkJ7_2),.clk(gclk));
	jdff dff_A_A9HHPL6c9_2(.dout(w_dff_A_mGAL2BkJ7_2),.din(w_dff_A_A9HHPL6c9_2),.clk(gclk));
	jdff dff_A_9ogfngCa2_2(.dout(w_dff_A_A9HHPL6c9_2),.din(w_dff_A_9ogfngCa2_2),.clk(gclk));
	jdff dff_A_XVAy8ZRa0_2(.dout(w_dff_A_9ogfngCa2_2),.din(w_dff_A_XVAy8ZRa0_2),.clk(gclk));
	jdff dff_A_FRIHcNj08_2(.dout(w_dff_A_XVAy8ZRa0_2),.din(w_dff_A_FRIHcNj08_2),.clk(gclk));
	jdff dff_A_igeem2lH7_2(.dout(w_dff_A_FRIHcNj08_2),.din(w_dff_A_igeem2lH7_2),.clk(gclk));
	jdff dff_A_3JeCS0Rb0_1(.dout(w_n618_0[1]),.din(w_dff_A_3JeCS0Rb0_1),.clk(gclk));
	jdff dff_A_tGz2ldo26_1(.dout(w_dff_A_3JeCS0Rb0_1),.din(w_dff_A_tGz2ldo26_1),.clk(gclk));
	jdff dff_A_Aj2wo3kE8_1(.dout(w_dff_A_tGz2ldo26_1),.din(w_dff_A_Aj2wo3kE8_1),.clk(gclk));
	jdff dff_A_uNBldFdh9_1(.dout(w_dff_A_Aj2wo3kE8_1),.din(w_dff_A_uNBldFdh9_1),.clk(gclk));
	jdff dff_A_jWl5fsZ09_1(.dout(w_dff_A_uNBldFdh9_1),.din(w_dff_A_jWl5fsZ09_1),.clk(gclk));
	jdff dff_A_4U3jWDXQ1_1(.dout(w_dff_A_jWl5fsZ09_1),.din(w_dff_A_4U3jWDXQ1_1),.clk(gclk));
	jdff dff_A_sFUW312X0_2(.dout(w_n618_0[2]),.din(w_dff_A_sFUW312X0_2),.clk(gclk));
	jdff dff_A_fdxC9CnN2_2(.dout(w_dff_A_sFUW312X0_2),.din(w_dff_A_fdxC9CnN2_2),.clk(gclk));
	jdff dff_A_qMHXqdRa3_2(.dout(w_dff_A_fdxC9CnN2_2),.din(w_dff_A_qMHXqdRa3_2),.clk(gclk));
	jdff dff_A_w7MUFPIP6_0(.dout(w_n1425_0[0]),.din(w_dff_A_w7MUFPIP6_0),.clk(gclk));
	jdff dff_B_rGgM8vH17_1(.din(n1411),.dout(w_dff_B_rGgM8vH17_1),.clk(gclk));
	jdff dff_A_pph0MgxZ3_0(.dout(w_n1422_0[0]),.din(w_dff_A_pph0MgxZ3_0),.clk(gclk));
	jdff dff_B_aMolQQ517_1(.din(n1418),.dout(w_dff_B_aMolQQ517_1),.clk(gclk));
	jdff dff_B_HoeLbVlP7_1(.din(w_dff_B_aMolQQ517_1),.dout(w_dff_B_HoeLbVlP7_1),.clk(gclk));
	jdff dff_B_gjHkMSii5_1(.din(w_dff_B_HoeLbVlP7_1),.dout(w_dff_B_gjHkMSii5_1),.clk(gclk));
	jdff dff_B_WS7nlbgh7_1(.din(n1419),.dout(w_dff_B_WS7nlbgh7_1),.clk(gclk));
	jdff dff_B_EPT7mUVs7_1(.din(w_dff_B_WS7nlbgh7_1),.dout(w_dff_B_EPT7mUVs7_1),.clk(gclk));
	jdff dff_A_IotwBgAe4_2(.dout(w_n660_0[2]),.din(w_dff_A_IotwBgAe4_2),.clk(gclk));
	jdff dff_A_fIBMuMh99_2(.dout(w_dff_A_IotwBgAe4_2),.din(w_dff_A_fIBMuMh99_2),.clk(gclk));
	jdff dff_A_FbaP9dS96_2(.dout(w_dff_A_fIBMuMh99_2),.din(w_dff_A_FbaP9dS96_2),.clk(gclk));
	jdff dff_A_j6HjCMk69_2(.dout(w_dff_A_FbaP9dS96_2),.din(w_dff_A_j6HjCMk69_2),.clk(gclk));
	jdff dff_A_tSJb9xXv4_2(.dout(w_dff_A_j6HjCMk69_2),.din(w_dff_A_tSJb9xXv4_2),.clk(gclk));
	jdff dff_A_lpXRusux6_2(.dout(w_dff_A_tSJb9xXv4_2),.din(w_dff_A_lpXRusux6_2),.clk(gclk));
	jdff dff_A_Z1cv1RsF6_2(.dout(w_n792_0[2]),.din(w_dff_A_Z1cv1RsF6_2),.clk(gclk));
	jdff dff_A_VJ4feSW02_2(.dout(w_dff_A_Z1cv1RsF6_2),.din(w_dff_A_VJ4feSW02_2),.clk(gclk));
	jdff dff_A_oZ9B3eiY8_2(.dout(w_dff_A_VJ4feSW02_2),.din(w_dff_A_oZ9B3eiY8_2),.clk(gclk));
	jdff dff_A_amKvZqLm9_2(.dout(w_dff_A_oZ9B3eiY8_2),.din(w_dff_A_amKvZqLm9_2),.clk(gclk));
	jdff dff_A_fb2ZOYWl2_2(.dout(w_dff_A_amKvZqLm9_2),.din(w_dff_A_fb2ZOYWl2_2),.clk(gclk));
	jdff dff_A_TOnJGDtJ1_2(.dout(w_dff_A_fb2ZOYWl2_2),.din(w_dff_A_TOnJGDtJ1_2),.clk(gclk));
	jdff dff_A_Fi3ptPpt7_2(.dout(w_dff_A_TOnJGDtJ1_2),.din(w_dff_A_Fi3ptPpt7_2),.clk(gclk));
	jdff dff_A_fh4gxAWV4_2(.dout(w_dff_A_Fi3ptPpt7_2),.din(w_dff_A_fh4gxAWV4_2),.clk(gclk));
	jdff dff_A_H7atk1yL6_2(.dout(w_dff_A_fh4gxAWV4_2),.din(w_dff_A_H7atk1yL6_2),.clk(gclk));
	jdff dff_A_p6IIo7T53_1(.dout(w_n790_0[1]),.din(w_dff_A_p6IIo7T53_1),.clk(gclk));
	jdff dff_A_ZuXyQCnJ5_1(.dout(w_dff_A_p6IIo7T53_1),.din(w_dff_A_ZuXyQCnJ5_1),.clk(gclk));
	jdff dff_A_eKvoSu1N5_1(.dout(w_dff_A_ZuXyQCnJ5_1),.din(w_dff_A_eKvoSu1N5_1),.clk(gclk));
	jdff dff_A_KKEvQSj34_1(.dout(w_dff_A_eKvoSu1N5_1),.din(w_dff_A_KKEvQSj34_1),.clk(gclk));
	jdff dff_A_D4pdAtop8_1(.dout(w_dff_A_KKEvQSj34_1),.din(w_dff_A_D4pdAtop8_1),.clk(gclk));
	jdff dff_A_FJSxXbdl7_1(.dout(w_dff_A_D4pdAtop8_1),.din(w_dff_A_FJSxXbdl7_1),.clk(gclk));
	jdff dff_A_xpvPGOKX5_1(.dout(w_dff_A_FJSxXbdl7_1),.din(w_dff_A_xpvPGOKX5_1),.clk(gclk));
	jdff dff_A_D3jclvVg1_1(.dout(w_dff_A_xpvPGOKX5_1),.din(w_dff_A_D3jclvVg1_1),.clk(gclk));
	jdff dff_A_HyqSYiZF9_1(.dout(w_dff_A_D3jclvVg1_1),.din(w_dff_A_HyqSYiZF9_1),.clk(gclk));
	jdff dff_A_VwbmPG1e6_1(.dout(w_dff_A_HyqSYiZF9_1),.din(w_dff_A_VwbmPG1e6_1),.clk(gclk));
	jdff dff_B_9fuAt7GB5_1(.din(n1413),.dout(w_dff_B_9fuAt7GB5_1),.clk(gclk));
	jdff dff_B_lUK1UlOm6_1(.din(w_dff_B_9fuAt7GB5_1),.dout(w_dff_B_lUK1UlOm6_1),.clk(gclk));
	jdff dff_B_WPPJIrq28_1(.din(w_dff_B_lUK1UlOm6_1),.dout(w_dff_B_WPPJIrq28_1),.clk(gclk));
	jdff dff_B_qr4C19tO9_1(.din(w_dff_B_WPPJIrq28_1),.dout(w_dff_B_qr4C19tO9_1),.clk(gclk));
	jdff dff_B_GRuNwgC55_1(.din(n1414),.dout(w_dff_B_GRuNwgC55_1),.clk(gclk));
	jdff dff_B_NrtkYxHm3_1(.din(w_dff_B_GRuNwgC55_1),.dout(w_dff_B_NrtkYxHm3_1),.clk(gclk));
	jdff dff_B_2IxeBqju2_1(.din(w_dff_B_NrtkYxHm3_1),.dout(w_dff_B_2IxeBqju2_1),.clk(gclk));
	jdff dff_A_iSB1yla53_1(.dout(w_n821_0[1]),.din(w_dff_A_iSB1yla53_1),.clk(gclk));
	jdff dff_B_SRgyzuye7_1(.din(n812),.dout(w_dff_B_SRgyzuye7_1),.clk(gclk));
	jdff dff_B_B3B9hQjx5_1(.din(w_dff_B_SRgyzuye7_1),.dout(w_dff_B_B3B9hQjx5_1),.clk(gclk));
	jdff dff_B_6y5gUE284_1(.din(w_dff_B_B3B9hQjx5_1),.dout(w_dff_B_6y5gUE284_1),.clk(gclk));
	jdff dff_B_hrLyDgLw7_1(.din(w_dff_B_6y5gUE284_1),.dout(w_dff_B_hrLyDgLw7_1),.clk(gclk));
	jdff dff_B_IFUxW3UB8_1(.din(n813),.dout(w_dff_B_IFUxW3UB8_1),.clk(gclk));
	jdff dff_B_NeZtH99f4_1(.din(w_dff_B_IFUxW3UB8_1),.dout(w_dff_B_NeZtH99f4_1),.clk(gclk));
	jdff dff_B_PzqaW83H4_1(.din(w_dff_B_NeZtH99f4_1),.dout(w_dff_B_PzqaW83H4_1),.clk(gclk));
	jdff dff_A_9EaeI22C0_1(.dout(w_n819_0[1]),.din(w_dff_A_9EaeI22C0_1),.clk(gclk));
	jdff dff_A_hZ5D2cD50_1(.dout(w_dff_A_9EaeI22C0_1),.din(w_dff_A_hZ5D2cD50_1),.clk(gclk));
	jdff dff_A_NcYLiKqL2_0(.dout(w_n377_1[0]),.din(w_dff_A_NcYLiKqL2_0),.clk(gclk));
	jdff dff_A_ANjvwgwf4_0(.dout(w_n814_0[0]),.din(w_dff_A_ANjvwgwf4_0),.clk(gclk));
	jdff dff_A_mxHttHXo8_0(.dout(w_dff_A_ANjvwgwf4_0),.din(w_dff_A_mxHttHXo8_0),.clk(gclk));
	jdff dff_A_ci6v7xUY3_0(.dout(w_dff_A_mxHttHXo8_0),.din(w_dff_A_ci6v7xUY3_0),.clk(gclk));
	jdff dff_A_yEJUWmDc9_1(.dout(w_n814_0[1]),.din(w_dff_A_yEJUWmDc9_1),.clk(gclk));
	jdff dff_A_qUeNlPd81_1(.dout(w_dff_A_yEJUWmDc9_1),.din(w_dff_A_qUeNlPd81_1),.clk(gclk));
	jdff dff_A_ITtg9bl70_2(.dout(w_n377_0[2]),.din(w_dff_A_ITtg9bl70_2),.clk(gclk));
	jdff dff_B_XnDd9siy9_3(.din(n377),.dout(w_dff_B_XnDd9siy9_3),.clk(gclk));
	jdff dff_A_vnwryK2G1_0(.dout(w_G534_2[0]),.din(w_dff_A_vnwryK2G1_0),.clk(gclk));
	jdff dff_A_hAlFR93x7_0(.dout(w_dff_A_vnwryK2G1_0),.din(w_dff_A_hAlFR93x7_0),.clk(gclk));
	jdff dff_A_jEfd3TcK5_0(.dout(w_dff_A_hAlFR93x7_0),.din(w_dff_A_jEfd3TcK5_0),.clk(gclk));
	jdff dff_A_YX2znO8M5_1(.dout(w_n1412_0[1]),.din(w_dff_A_YX2znO8M5_1),.clk(gclk));
	jdff dff_A_gOqqgfa46_1(.dout(w_dff_A_YX2znO8M5_1),.din(w_dff_A_gOqqgfa46_1),.clk(gclk));
	jdff dff_A_DisGo5P51_2(.dout(w_n1412_0[2]),.din(w_dff_A_DisGo5P51_2),.clk(gclk));
	jdff dff_B_8Q3FfvoL7_3(.din(n1412),.dout(w_dff_B_8Q3FfvoL7_3),.clk(gclk));
	jdff dff_B_pbMff5Cz1_3(.din(w_dff_B_8Q3FfvoL7_3),.dout(w_dff_B_pbMff5Cz1_3),.clk(gclk));
	jdff dff_B_POX1SfP90_3(.din(w_dff_B_pbMff5Cz1_3),.dout(w_dff_B_POX1SfP90_3),.clk(gclk));
	jdff dff_B_VnSme4hm7_3(.din(w_dff_B_POX1SfP90_3),.dout(w_dff_B_VnSme4hm7_3),.clk(gclk));
	jdff dff_B_80wDeluw5_3(.din(w_dff_B_VnSme4hm7_3),.dout(w_dff_B_80wDeluw5_3),.clk(gclk));
	jdff dff_B_BoJPt3mV0_3(.din(w_dff_B_80wDeluw5_3),.dout(w_dff_B_BoJPt3mV0_3),.clk(gclk));
	jdff dff_B_zcciXxZc3_3(.din(w_dff_B_BoJPt3mV0_3),.dout(w_dff_B_zcciXxZc3_3),.clk(gclk));
	jdff dff_B_4vv7aUqS2_3(.din(w_dff_B_zcciXxZc3_3),.dout(w_dff_B_4vv7aUqS2_3),.clk(gclk));
	jdff dff_B_bPFowCxE0_3(.din(w_dff_B_4vv7aUqS2_3),.dout(w_dff_B_bPFowCxE0_3),.clk(gclk));
	jdff dff_B_X9d1K3tK5_3(.din(w_dff_B_bPFowCxE0_3),.dout(w_dff_B_X9d1K3tK5_3),.clk(gclk));
	jdff dff_A_eJBzFm3K3_0(.dout(w_G2174_0[0]),.din(w_dff_A_eJBzFm3K3_0),.clk(gclk));
	jdff dff_A_1fyaFBeA8_0(.dout(w_dff_A_eJBzFm3K3_0),.din(w_dff_A_1fyaFBeA8_0),.clk(gclk));
	jdff dff_A_5UZS9S6D2_0(.dout(w_dff_A_1fyaFBeA8_0),.din(w_dff_A_5UZS9S6D2_0),.clk(gclk));
	jdff dff_A_n2wbnxKo6_0(.dout(w_dff_A_5UZS9S6D2_0),.din(w_dff_A_n2wbnxKo6_0),.clk(gclk));
	jdff dff_A_1dsQ5K8h8_0(.dout(w_dff_A_n2wbnxKo6_0),.din(w_dff_A_1dsQ5K8h8_0),.clk(gclk));
	jdff dff_A_riFO6sSa8_0(.dout(w_dff_A_1dsQ5K8h8_0),.din(w_dff_A_riFO6sSa8_0),.clk(gclk));
	jdff dff_A_N3lgVb1j0_0(.dout(w_dff_A_riFO6sSa8_0),.din(w_dff_A_N3lgVb1j0_0),.clk(gclk));
	jdff dff_A_fWXMmo2N7_0(.dout(w_dff_A_N3lgVb1j0_0),.din(w_dff_A_fWXMmo2N7_0),.clk(gclk));
	jdff dff_A_DaPhHxza4_0(.dout(w_dff_A_fWXMmo2N7_0),.din(w_dff_A_DaPhHxza4_0),.clk(gclk));
	jdff dff_A_13B4Nrks8_0(.dout(w_dff_A_DaPhHxza4_0),.din(w_dff_A_13B4Nrks8_0),.clk(gclk));
	jdff dff_A_gZ5FYZpZ7_0(.dout(w_dff_A_13B4Nrks8_0),.din(w_dff_A_gZ5FYZpZ7_0),.clk(gclk));
	jdff dff_A_YPSpdvYW5_0(.dout(w_dff_A_gZ5FYZpZ7_0),.din(w_dff_A_YPSpdvYW5_0),.clk(gclk));
	jdff dff_A_iO8l3Xcp1_0(.dout(w_dff_A_YPSpdvYW5_0),.din(w_dff_A_iO8l3Xcp1_0),.clk(gclk));
	jdff dff_A_2wygWxmI5_1(.dout(w_G2174_0[1]),.din(w_dff_A_2wygWxmI5_1),.clk(gclk));
	jdff dff_A_eY4OjLz98_1(.dout(w_dff_A_2wygWxmI5_1),.din(w_dff_A_eY4OjLz98_1),.clk(gclk));
	jdff dff_A_tr02KA827_1(.dout(w_dff_A_eY4OjLz98_1),.din(w_dff_A_tr02KA827_1),.clk(gclk));
	jdff dff_A_hXEBdvMU1_1(.dout(w_dff_A_tr02KA827_1),.din(w_dff_A_hXEBdvMU1_1),.clk(gclk));
	jdff dff_A_XdB1QHq36_1(.dout(w_dff_A_hXEBdvMU1_1),.din(w_dff_A_XdB1QHq36_1),.clk(gclk));
	jdff dff_A_kTLuUohm9_1(.dout(w_dff_A_XdB1QHq36_1),.din(w_dff_A_kTLuUohm9_1),.clk(gclk));
	jdff dff_A_ntI7QtOM7_1(.dout(w_dff_A_kTLuUohm9_1),.din(w_dff_A_ntI7QtOM7_1),.clk(gclk));
	jdff dff_A_DtcriHOY9_1(.dout(w_dff_A_ntI7QtOM7_1),.din(w_dff_A_DtcriHOY9_1),.clk(gclk));
	jdff dff_A_eAAHlm9e9_1(.dout(w_dff_A_DtcriHOY9_1),.din(w_dff_A_eAAHlm9e9_1),.clk(gclk));
	jdff dff_A_inQvp69a0_1(.dout(w_dff_A_eAAHlm9e9_1),.din(w_dff_A_inQvp69a0_1),.clk(gclk));
	jdff dff_A_FPsJvK3N9_0(.dout(w_n1410_0[0]),.din(w_dff_A_FPsJvK3N9_0),.clk(gclk));
	jdff dff_B_sagk3Rbh6_0(.din(n1409),.dout(w_dff_B_sagk3Rbh6_0),.clk(gclk));
	jdff dff_B_JPQ5n1MR2_0(.din(w_dff_B_sagk3Rbh6_0),.dout(w_dff_B_JPQ5n1MR2_0),.clk(gclk));
	jdff dff_A_VjKBCpmZ8_0(.dout(w_n401_0[0]),.din(w_dff_A_VjKBCpmZ8_0),.clk(gclk));
	jdff dff_A_1mMfmRST8_0(.dout(w_dff_A_VjKBCpmZ8_0),.din(w_dff_A_1mMfmRST8_0),.clk(gclk));
	jdff dff_A_Mpz7Wox11_0(.dout(w_dff_A_1mMfmRST8_0),.din(w_dff_A_Mpz7Wox11_0),.clk(gclk));
	jdff dff_B_4XfIYN468_2(.din(n401),.dout(w_dff_B_4XfIYN468_2),.clk(gclk));
	jdff dff_A_lLMQcsDI1_0(.dout(w_G490_1[0]),.din(w_dff_A_lLMQcsDI1_0),.clk(gclk));
	jdff dff_A_mYnJAxXX6_0(.dout(w_dff_A_lLMQcsDI1_0),.din(w_dff_A_mYnJAxXX6_0),.clk(gclk));
	jdff dff_A_Knhhl1uN2_0(.dout(w_dff_A_mYnJAxXX6_0),.din(w_dff_A_Knhhl1uN2_0),.clk(gclk));
	jdff dff_A_HEhayoAF5_1(.dout(w_n654_1[1]),.din(w_dff_A_HEhayoAF5_1),.clk(gclk));
	jdff dff_A_Mm1K6Wtr8_1(.dout(w_dff_A_HEhayoAF5_1),.din(w_dff_A_Mm1K6Wtr8_1),.clk(gclk));
	jdff dff_A_9nVqtLlm0_1(.dout(w_dff_A_Mm1K6Wtr8_1),.din(w_dff_A_9nVqtLlm0_1),.clk(gclk));
	jdff dff_A_HIQsbQFI5_1(.dout(w_dff_A_9nVqtLlm0_1),.din(w_dff_A_HIQsbQFI5_1),.clk(gclk));
	jdff dff_A_5s9HAUx73_1(.dout(w_dff_A_HIQsbQFI5_1),.din(w_dff_A_5s9HAUx73_1),.clk(gclk));
	jdff dff_A_aWOUgwhr9_1(.dout(w_dff_A_5s9HAUx73_1),.din(w_dff_A_aWOUgwhr9_1),.clk(gclk));
	jdff dff_A_TLALxBQU3_1(.dout(w_dff_A_aWOUgwhr9_1),.din(w_dff_A_TLALxBQU3_1),.clk(gclk));
	jdff dff_A_b3hINvNF7_1(.dout(w_dff_A_TLALxBQU3_1),.din(w_dff_A_b3hINvNF7_1),.clk(gclk));
	jdff dff_A_q5eO7kLE9_0(.dout(w_n644_0[0]),.din(w_dff_A_q5eO7kLE9_0),.clk(gclk));
	jdff dff_A_nnT4j9Jv7_0(.dout(w_dff_A_q5eO7kLE9_0),.din(w_dff_A_nnT4j9Jv7_0),.clk(gclk));
	jdff dff_A_AL058DZw2_0(.dout(w_dff_A_nnT4j9Jv7_0),.din(w_dff_A_AL058DZw2_0),.clk(gclk));
	jdff dff_A_908jh8XE2_0(.dout(w_dff_A_AL058DZw2_0),.din(w_dff_A_908jh8XE2_0),.clk(gclk));
	jdff dff_A_IIOM7Qkz1_2(.dout(w_n644_0[2]),.din(w_dff_A_IIOM7Qkz1_2),.clk(gclk));
	jdff dff_A_zyvbQmbi4_2(.dout(w_dff_A_IIOM7Qkz1_2),.din(w_dff_A_zyvbQmbi4_2),.clk(gclk));
	jdff dff_A_G0NBzf615_1(.dout(w_G293_0[1]),.din(w_dff_A_G0NBzf615_1),.clk(gclk));
	jdff dff_A_suv6ryfC7_1(.dout(w_n746_0[1]),.din(w_dff_A_suv6ryfC7_1),.clk(gclk));
	jdff dff_A_YnTQFQCz7_1(.dout(w_dff_A_suv6ryfC7_1),.din(w_dff_A_YnTQFQCz7_1),.clk(gclk));
	jdff dff_A_KJtXCf6k5_1(.dout(w_dff_A_YnTQFQCz7_1),.din(w_dff_A_KJtXCf6k5_1),.clk(gclk));
	jdff dff_A_AGM8M7Sv0_1(.dout(w_dff_A_KJtXCf6k5_1),.din(w_dff_A_AGM8M7Sv0_1),.clk(gclk));
	jdff dff_B_jb0y8H540_1(.din(n741),.dout(w_dff_B_jb0y8H540_1),.clk(gclk));
	jdff dff_B_w5V504Yr2_1(.din(w_dff_B_jb0y8H540_1),.dout(w_dff_B_w5V504Yr2_1),.clk(gclk));
	jdff dff_A_plH1km8d8_1(.dout(w_n742_0[1]),.din(w_dff_A_plH1km8d8_1),.clk(gclk));
	jdff dff_A_RWh6EijB0_1(.dout(w_dff_A_plH1km8d8_1),.din(w_dff_A_RWh6EijB0_1),.clk(gclk));
	jdff dff_A_KxjkrfVe2_1(.dout(w_dff_A_RWh6EijB0_1),.din(w_dff_A_KxjkrfVe2_1),.clk(gclk));
	jdff dff_A_wBrxynoD4_1(.dout(w_dff_A_KxjkrfVe2_1),.din(w_dff_A_wBrxynoD4_1),.clk(gclk));
	jdff dff_A_sWBYShcs2_1(.dout(w_dff_A_wBrxynoD4_1),.din(w_dff_A_sWBYShcs2_1),.clk(gclk));
	jdff dff_A_sztsfTGm4_1(.dout(w_dff_A_sWBYShcs2_1),.din(w_dff_A_sztsfTGm4_1),.clk(gclk));
	jdff dff_A_h2ENW0g59_1(.dout(w_dff_A_sztsfTGm4_1),.din(w_dff_A_h2ENW0g59_1),.clk(gclk));
	jdff dff_B_yFdrxyFS0_0(.din(n657),.dout(w_dff_B_yFdrxyFS0_0),.clk(gclk));
	jdff dff_B_jWYeyIKN8_1(.din(G323),.dout(w_dff_B_jWYeyIKN8_1),.clk(gclk));
	jdff dff_A_6KzOBrkF1_2(.dout(w_G316_0[2]),.din(w_dff_A_6KzOBrkF1_2),.clk(gclk));
	jdff dff_A_UgdAQFHI9_1(.dout(w_G490_0[1]),.din(w_dff_A_UgdAQFHI9_1),.clk(gclk));
	jdff dff_A_nWJxO2Ho7_1(.dout(w_dff_A_UgdAQFHI9_1),.din(w_dff_A_nWJxO2Ho7_1),.clk(gclk));
	jdff dff_A_mbyb7jcW9_1(.dout(w_dff_A_nWJxO2Ho7_1),.din(w_dff_A_mbyb7jcW9_1),.clk(gclk));
	jdff dff_A_zutWcC9k7_1(.dout(w_dff_A_mbyb7jcW9_1),.din(w_dff_A_zutWcC9k7_1),.clk(gclk));
	jdff dff_A_rKzJjZLt6_2(.dout(w_G490_0[2]),.din(w_dff_A_rKzJjZLt6_2),.clk(gclk));
	jdff dff_A_aD3rUtgm9_2(.dout(w_dff_A_rKzJjZLt6_2),.din(w_dff_A_aD3rUtgm9_2),.clk(gclk));
	jdff dff_A_fIw77XNS0_2(.dout(w_dff_A_aD3rUtgm9_2),.din(w_dff_A_fIw77XNS0_2),.clk(gclk));
	jdff dff_A_ZvPz6YQa3_2(.dout(w_dff_A_fIw77XNS0_2),.din(w_dff_A_ZvPz6YQa3_2),.clk(gclk));
	jdff dff_A_dQzCsD9g8_0(.dout(w_n654_2[0]),.din(w_dff_A_dQzCsD9g8_0),.clk(gclk));
	jdff dff_A_v3GcPNiR7_0(.dout(w_n654_0[0]),.din(w_dff_A_v3GcPNiR7_0),.clk(gclk));
	jdff dff_B_vw3vRAA64_3(.din(n654),.dout(w_dff_B_vw3vRAA64_3),.clk(gclk));
	jdff dff_A_HWxL4K037_0(.dout(w_n653_0[0]),.din(w_dff_A_HWxL4K037_0),.clk(gclk));
	jdff dff_B_4pBthudu4_1(.din(n651),.dout(w_dff_B_4pBthudu4_1),.clk(gclk));
	jdff dff_B_TkDvYJKb3_1(.din(G315),.dout(w_dff_B_TkDvYJKb3_1),.clk(gclk));
	jdff dff_A_CRbXyWah2_0(.dout(w_n414_0[0]),.din(w_dff_A_CRbXyWah2_0),.clk(gclk));
	jdff dff_A_VNOLxWZW2_0(.dout(w_dff_A_CRbXyWah2_0),.din(w_dff_A_VNOLxWZW2_0),.clk(gclk));
	jdff dff_B_ONHJmS7E4_2(.din(n414),.dout(w_dff_B_ONHJmS7E4_2),.clk(gclk));
	jdff dff_A_FXZqEKHe9_0(.dout(w_G479_0[0]),.din(w_dff_A_FXZqEKHe9_0),.clk(gclk));
	jdff dff_A_GmEHFD3f9_0(.dout(w_dff_A_FXZqEKHe9_0),.din(w_dff_A_GmEHFD3f9_0),.clk(gclk));
	jdff dff_A_HdGKWoCy4_0(.dout(w_dff_A_GmEHFD3f9_0),.din(w_dff_A_HdGKWoCy4_0),.clk(gclk));
	jdff dff_A_77MecEph4_1(.dout(w_G479_0[1]),.din(w_dff_A_77MecEph4_1),.clk(gclk));
	jdff dff_A_W8er2Mim7_1(.dout(w_dff_A_77MecEph4_1),.din(w_dff_A_W8er2Mim7_1),.clk(gclk));
	jdff dff_A_DMdqylml7_1(.dout(w_dff_A_W8er2Mim7_1),.din(w_dff_A_DMdqylml7_1),.clk(gclk));
	jdff dff_A_aYMbA9d67_1(.dout(w_n648_0[1]),.din(w_dff_A_aYMbA9d67_1),.clk(gclk));
	jdff dff_A_xJZG6co13_1(.dout(w_dff_A_aYMbA9d67_1),.din(w_dff_A_xJZG6co13_1),.clk(gclk));
	jdff dff_A_ltIQVsce8_1(.dout(w_dff_A_xJZG6co13_1),.din(w_dff_A_ltIQVsce8_1),.clk(gclk));
	jdff dff_A_Pdohg5pg3_1(.dout(w_dff_A_ltIQVsce8_1),.din(w_dff_A_Pdohg5pg3_1),.clk(gclk));
	jdff dff_A_K3cruJ2w0_2(.dout(w_n648_0[2]),.din(w_dff_A_K3cruJ2w0_2),.clk(gclk));
	jdff dff_A_DI0ckUu57_2(.dout(w_dff_A_K3cruJ2w0_2),.din(w_dff_A_DI0ckUu57_2),.clk(gclk));
	jdff dff_A_qpfmLGMv9_2(.dout(w_dff_A_DI0ckUu57_2),.din(w_dff_A_qpfmLGMv9_2),.clk(gclk));
	jdff dff_A_Azp1elas1_2(.dout(w_dff_A_qpfmLGMv9_2),.din(w_dff_A_Azp1elas1_2),.clk(gclk));
	jdff dff_A_z5GEAU9j4_2(.dout(w_dff_A_Azp1elas1_2),.din(w_dff_A_z5GEAU9j4_2),.clk(gclk));
	jdff dff_B_LqUkf7YI2_0(.din(n647),.dout(w_dff_B_LqUkf7YI2_0),.clk(gclk));
	jdff dff_B_TZ9GQanc9_1(.din(G307),.dout(w_dff_B_TZ9GQanc9_1),.clk(gclk));
	jdff dff_A_AHXN0R4U7_0(.dout(w_G302_0[0]),.din(w_dff_A_AHXN0R4U7_0),.clk(gclk));
	jdff dff_A_mio5KJpD3_1(.dout(w_G302_0[1]),.din(w_dff_A_mio5KJpD3_1),.clk(gclk));
	jdff dff_B_sQM3zmHS5_1(.din(n727),.dout(w_dff_B_sQM3zmHS5_1),.clk(gclk));
	jdff dff_A_GtdLA4qw5_0(.dout(w_n635_1[0]),.din(w_dff_A_GtdLA4qw5_0),.clk(gclk));
	jdff dff_A_ShosyFsw9_1(.dout(w_n635_0[1]),.din(w_dff_A_ShosyFsw9_1),.clk(gclk));
	jdff dff_A_vKyo0vsz3_1(.dout(w_dff_A_ShosyFsw9_1),.din(w_dff_A_vKyo0vsz3_1),.clk(gclk));
	jdff dff_B_D4YMhMGO0_1(.din(n633),.dout(w_dff_B_D4YMhMGO0_1),.clk(gclk));
	jdff dff_A_zCn3yGKH3_0(.dout(w_G366_0[0]),.din(w_dff_A_zCn3yGKH3_0),.clk(gclk));
	jdff dff_A_X7X2iXnx4_0(.dout(w_G332_2[0]),.din(w_dff_A_X7X2iXnx4_0),.clk(gclk));
	jdff dff_A_z476YpM93_2(.dout(w_G332_2[2]),.din(w_dff_A_z476YpM93_2),.clk(gclk));
	jdff dff_A_Dy7yROMc0_0(.dout(w_n628_0[0]),.din(w_dff_A_Dy7yROMc0_0),.clk(gclk));
	jdff dff_A_IJzczlmd7_0(.dout(w_dff_A_Dy7yROMc0_0),.din(w_dff_A_IJzczlmd7_0),.clk(gclk));
	jdff dff_A_uudzYH4a6_0(.dout(w_dff_A_IJzczlmd7_0),.din(w_dff_A_uudzYH4a6_0),.clk(gclk));
	jdff dff_A_DIDKx7dg3_2(.dout(w_n628_0[2]),.din(w_dff_A_DIDKx7dg3_2),.clk(gclk));
	jdff dff_A_4Jm7U9iH9_0(.dout(w_G358_0[0]),.din(w_dff_A_4Jm7U9iH9_0),.clk(gclk));
	jdff dff_A_2JWxP9z98_1(.dout(w_n625_0[1]),.din(w_dff_A_2JWxP9z98_1),.clk(gclk));
	jdff dff_A_mPKOD2o62_2(.dout(w_G351_0[2]),.din(w_dff_A_mPKOD2o62_2),.clk(gclk));
	jdff dff_A_RsPkIsbe4_0(.dout(w_G534_0[0]),.din(w_dff_A_RsPkIsbe4_0),.clk(gclk));
	jdff dff_A_LADkelDj8_0(.dout(w_dff_A_RsPkIsbe4_0),.din(w_dff_A_LADkelDj8_0),.clk(gclk));
	jdff dff_A_zizoQuCR7_0(.dout(w_dff_A_LADkelDj8_0),.din(w_dff_A_zizoQuCR7_0),.clk(gclk));
	jdff dff_A_DMbad3hU7_2(.dout(w_G534_0[2]),.din(w_dff_A_DMbad3hU7_2),.clk(gclk));
	jdff dff_A_JGbEjWLn7_2(.dout(w_dff_A_DMbad3hU7_2),.din(w_dff_A_JGbEjWLn7_2),.clk(gclk));
	jdff dff_A_OxQjbA5L0_2(.dout(w_dff_A_JGbEjWLn7_2),.din(w_dff_A_OxQjbA5L0_2),.clk(gclk));
	jdff dff_A_BDpeNNmD2_0(.dout(w_n726_0[0]),.din(w_dff_A_BDpeNNmD2_0),.clk(gclk));
	jdff dff_A_X7ZMSWaE8_0(.dout(w_dff_A_BDpeNNmD2_0),.din(w_dff_A_X7ZMSWaE8_0),.clk(gclk));
	jdff dff_A_FIfD5XyQ4_0(.dout(w_G348_0[0]),.din(w_dff_A_FIfD5XyQ4_0),.clk(gclk));
	jdff dff_A_MtyJ4roH9_1(.dout(w_G332_1[1]),.din(w_dff_A_MtyJ4roH9_1),.clk(gclk));
	jdff dff_A_ckaHTcbS1_1(.dout(w_n621_0[1]),.din(w_dff_A_ckaHTcbS1_1),.clk(gclk));
	jdff dff_A_E8mdAG5M9_2(.dout(w_G341_0[2]),.din(w_dff_A_E8mdAG5M9_2),.clk(gclk));
	jdff dff_A_DrDwCHlH4_0(.dout(w_n389_1[0]),.din(w_dff_A_DrDwCHlH4_0),.clk(gclk));
	jdff dff_A_xx4rnksF6_2(.dout(w_n389_0[2]),.din(w_dff_A_xx4rnksF6_2),.clk(gclk));
	jdff dff_B_5144iDOd1_3(.din(n389),.dout(w_dff_B_5144iDOd1_3),.clk(gclk));
	jdff dff_A_0RiWWR2i3_0(.dout(w_G523_1[0]),.din(w_dff_A_0RiWWR2i3_0),.clk(gclk));
	jdff dff_A_nwJKUgmw2_0(.dout(w_dff_A_0RiWWR2i3_0),.din(w_dff_A_nwJKUgmw2_0),.clk(gclk));
	jdff dff_A_a1pkJkDq3_0(.dout(w_dff_A_nwJKUgmw2_0),.din(w_dff_A_a1pkJkDq3_0),.clk(gclk));
	jdff dff_A_cCHYyOHs7_1(.dout(w_G523_1[1]),.din(w_dff_A_cCHYyOHs7_1),.clk(gclk));
	jdff dff_A_VpVhB3k29_1(.dout(w_dff_A_cCHYyOHs7_1),.din(w_dff_A_VpVhB3k29_1),.clk(gclk));
	jdff dff_A_5Ds71fVU2_1(.dout(w_dff_A_VpVhB3k29_1),.din(w_dff_A_5Ds71fVU2_1),.clk(gclk));
	jdff dff_A_hrEhE4iP4_1(.dout(w_G523_0[1]),.din(w_dff_A_hrEhE4iP4_1),.clk(gclk));
	jdff dff_A_zh3jNfwi9_1(.dout(w_dff_A_hrEhE4iP4_1),.din(w_dff_A_zh3jNfwi9_1),.clk(gclk));
	jdff dff_A_06pQuPHL0_1(.dout(w_dff_A_zh3jNfwi9_1),.din(w_dff_A_06pQuPHL0_1),.clk(gclk));
	jdff dff_A_6DzUmaNR4_2(.dout(w_G523_0[2]),.din(w_dff_A_6DzUmaNR4_2),.clk(gclk));
	jdff dff_A_X3m6gHGT3_2(.dout(w_dff_A_6DzUmaNR4_2),.din(w_dff_A_X3m6gHGT3_2),.clk(gclk));
	jdff dff_A_vVYz0nIU7_2(.dout(w_dff_A_X3m6gHGT3_2),.din(w_dff_A_vVYz0nIU7_2),.clk(gclk));
	jdff dff_A_j7HvhEyZ8_1(.dout(w_n722_0[1]),.din(w_dff_A_j7HvhEyZ8_1),.clk(gclk));
	jdff dff_A_ezuIGCO32_1(.dout(w_dff_A_j7HvhEyZ8_1),.din(w_dff_A_ezuIGCO32_1),.clk(gclk));
	jdff dff_A_62MADGjn5_1(.dout(w_dff_A_ezuIGCO32_1),.din(w_dff_A_62MADGjn5_1),.clk(gclk));
	jdff dff_A_dMeO5M2X8_1(.dout(w_dff_A_62MADGjn5_1),.din(w_dff_A_dMeO5M2X8_1),.clk(gclk));
	jdff dff_A_mqI9zWK44_1(.dout(w_n721_0[1]),.din(w_dff_A_mqI9zWK44_1),.clk(gclk));
	jdff dff_A_77yJpoSn1_1(.dout(w_dff_A_mqI9zWK44_1),.din(w_dff_A_77yJpoSn1_1),.clk(gclk));
	jdff dff_A_Hcj920qD0_1(.dout(w_dff_A_77yJpoSn1_1),.din(w_dff_A_Hcj920qD0_1),.clk(gclk));
	jdff dff_A_qZvNo7G69_1(.dout(w_dff_A_Hcj920qD0_1),.din(w_dff_A_qZvNo7G69_1),.clk(gclk));
	jdff dff_A_ysBaB5zn3_1(.dout(w_dff_A_qZvNo7G69_1),.din(w_dff_A_ysBaB5zn3_1),.clk(gclk));
	jdff dff_A_Su4vCRfa8_1(.dout(w_n619_0[1]),.din(w_dff_A_Su4vCRfa8_1),.clk(gclk));
	jdff dff_A_Q12d3uM86_1(.dout(w_dff_A_Su4vCRfa8_1),.din(w_dff_A_Q12d3uM86_1),.clk(gclk));
	jdff dff_A_IPcIksHL9_0(.dout(w_G338_0[0]),.din(w_dff_A_IPcIksHL9_0),.clk(gclk));
	jdff dff_A_ffhFOXib9_0(.dout(w_G514_0[0]),.din(w_dff_A_ffhFOXib9_0),.clk(gclk));
	jdff dff_A_4vW2gdeH9_0(.dout(w_dff_A_ffhFOXib9_0),.din(w_dff_A_4vW2gdeH9_0),.clk(gclk));
	jdff dff_A_QJgWHiKz1_2(.dout(w_G514_0[2]),.din(w_dff_A_QJgWHiKz1_2),.clk(gclk));
	jdff dff_A_rAA9UwGv7_1(.dout(w_n720_0[1]),.din(w_dff_A_rAA9UwGv7_1),.clk(gclk));
	jdff dff_A_SXdVppZN2_1(.dout(w_dff_A_rAA9UwGv7_1),.din(w_dff_A_SXdVppZN2_1),.clk(gclk));
	jdff dff_A_RkwJ56zm0_1(.dout(w_dff_A_SXdVppZN2_1),.din(w_dff_A_RkwJ56zm0_1),.clk(gclk));
	jdff dff_A_qoh4vhNv1_1(.dout(w_dff_A_RkwJ56zm0_1),.din(w_dff_A_qoh4vhNv1_1),.clk(gclk));
	jdff dff_A_nh51Fih91_1(.dout(w_n719_0[1]),.din(w_dff_A_nh51Fih91_1),.clk(gclk));
	jdff dff_A_y7muOgyZ4_1(.dout(w_dff_A_nh51Fih91_1),.din(w_dff_A_y7muOgyZ4_1),.clk(gclk));
	jdff dff_A_3DNjikiI9_1(.dout(w_dff_A_y7muOgyZ4_1),.din(w_dff_A_3DNjikiI9_1),.clk(gclk));
	jdff dff_A_QZDGlfHh3_1(.dout(w_dff_A_3DNjikiI9_1),.din(w_dff_A_QZDGlfHh3_1),.clk(gclk));
	jdff dff_A_UnSMDFQx4_1(.dout(w_dff_A_QZDGlfHh3_1),.din(w_dff_A_UnSMDFQx4_1),.clk(gclk));
	jdff dff_B_XT6WQqUp7_0(.din(n616),.dout(w_dff_B_XT6WQqUp7_0),.clk(gclk));
	jdff dff_A_1BDoj2j67_1(.dout(w_G331_0[1]),.din(w_dff_A_1BDoj2j67_1),.clk(gclk));
	jdff dff_A_UNfn2Mjz9_1(.dout(w_G324_1[1]),.din(w_dff_A_UNfn2Mjz9_1),.clk(gclk));
	jdff dff_A_ws0VB4db8_2(.dout(w_G324_0[2]),.din(w_dff_A_ws0VB4db8_2),.clk(gclk));
	jdff dff_A_804CLJld9_0(.dout(w_G503_0[0]),.din(w_dff_A_804CLJld9_0),.clk(gclk));
	jdff dff_A_qAHGF4p58_0(.dout(w_dff_A_804CLJld9_0),.din(w_dff_A_qAHGF4p58_0),.clk(gclk));
	jdff dff_A_Zje9Avjg1_0(.dout(w_dff_A_qAHGF4p58_0),.din(w_dff_A_Zje9Avjg1_0),.clk(gclk));
	jdff dff_A_zj7BXK0S0_0(.dout(w_dff_A_Zje9Avjg1_0),.din(w_dff_A_zj7BXK0S0_0),.clk(gclk));
	jdff dff_A_yshMyeTV6_2(.dout(w_G503_0[2]),.din(w_dff_A_yshMyeTV6_2),.clk(gclk));
	jdff dff_A_tnwJ9HxF4_2(.dout(w_dff_A_yshMyeTV6_2),.din(w_dff_A_tnwJ9HxF4_2),.clk(gclk));
	jdff dff_A_zPkn3j5y7_0(.dout(w_G4092_4[0]),.din(w_dff_A_zPkn3j5y7_0),.clk(gclk));
	jdff dff_A_fpMLpCsI5_0(.dout(w_dff_A_zPkn3j5y7_0),.din(w_dff_A_fpMLpCsI5_0),.clk(gclk));
	jdff dff_A_eybolzBm1_0(.dout(w_dff_A_fpMLpCsI5_0),.din(w_dff_A_eybolzBm1_0),.clk(gclk));
	jdff dff_A_9yck677m1_0(.dout(w_dff_A_eybolzBm1_0),.din(w_dff_A_9yck677m1_0),.clk(gclk));
	jdff dff_A_ipuRDokf7_0(.dout(w_dff_A_9yck677m1_0),.din(w_dff_A_ipuRDokf7_0),.clk(gclk));
	jdff dff_A_h0ySRBKO7_0(.dout(w_dff_A_ipuRDokf7_0),.din(w_dff_A_h0ySRBKO7_0),.clk(gclk));
	jdff dff_A_snFo9xDQ4_0(.dout(w_dff_A_h0ySRBKO7_0),.din(w_dff_A_snFo9xDQ4_0),.clk(gclk));
	jdff dff_A_8BKRwdoV7_0(.dout(w_dff_A_snFo9xDQ4_0),.din(w_dff_A_8BKRwdoV7_0),.clk(gclk));
	jdff dff_A_gBj7XBNV9_0(.dout(w_dff_A_8BKRwdoV7_0),.din(w_dff_A_gBj7XBNV9_0),.clk(gclk));
	jdff dff_A_La1cuWoT6_0(.dout(w_dff_A_gBj7XBNV9_0),.din(w_dff_A_La1cuWoT6_0),.clk(gclk));
	jdff dff_A_hhz5Finv0_0(.dout(w_dff_A_La1cuWoT6_0),.din(w_dff_A_hhz5Finv0_0),.clk(gclk));
	jdff dff_A_um0Y8Tlh3_0(.dout(w_dff_A_hhz5Finv0_0),.din(w_dff_A_um0Y8Tlh3_0),.clk(gclk));
	jdff dff_A_dXCQTO4B1_0(.dout(w_dff_A_um0Y8Tlh3_0),.din(w_dff_A_dXCQTO4B1_0),.clk(gclk));
	jdff dff_A_8XkyozXV8_0(.dout(w_dff_A_dXCQTO4B1_0),.din(w_dff_A_8XkyozXV8_0),.clk(gclk));
	jdff dff_A_5AjmUA0r5_0(.dout(w_G4092_1[0]),.din(w_dff_A_5AjmUA0r5_0),.clk(gclk));
	jdff dff_A_8cAvl1RM6_0(.dout(w_dff_A_5AjmUA0r5_0),.din(w_dff_A_8cAvl1RM6_0),.clk(gclk));
	jdff dff_A_6FZFw8Wn2_0(.dout(w_dff_A_8cAvl1RM6_0),.din(w_dff_A_6FZFw8Wn2_0),.clk(gclk));
	jdff dff_A_UMb2lxUr7_0(.dout(w_dff_A_6FZFw8Wn2_0),.din(w_dff_A_UMb2lxUr7_0),.clk(gclk));
	jdff dff_A_UThKjtyT3_0(.dout(w_dff_A_UMb2lxUr7_0),.din(w_dff_A_UThKjtyT3_0),.clk(gclk));
	jdff dff_A_B5jVEXVJ8_0(.dout(w_dff_A_UThKjtyT3_0),.din(w_dff_A_B5jVEXVJ8_0),.clk(gclk));
	jdff dff_A_IyFtmgwg1_2(.dout(w_G4092_1[2]),.din(w_dff_A_IyFtmgwg1_2),.clk(gclk));
	jdff dff_A_93sZyrYH7_2(.dout(w_dff_A_IyFtmgwg1_2),.din(w_dff_A_93sZyrYH7_2),.clk(gclk));
	jdff dff_A_vwpPry2y5_2(.dout(w_dff_A_93sZyrYH7_2),.din(w_dff_A_vwpPry2y5_2),.clk(gclk));
	jdff dff_A_MqQyiEH24_2(.dout(w_dff_A_vwpPry2y5_2),.din(w_dff_A_MqQyiEH24_2),.clk(gclk));
	jdff dff_B_BkxlJdZ46_0(.din(n1673),.dout(w_dff_B_BkxlJdZ46_0),.clk(gclk));
	jdff dff_B_O0ZUx5wi3_0(.din(w_dff_B_BkxlJdZ46_0),.dout(w_dff_B_O0ZUx5wi3_0),.clk(gclk));
	jdff dff_B_WxdPq4aF7_0(.din(w_dff_B_O0ZUx5wi3_0),.dout(w_dff_B_WxdPq4aF7_0),.clk(gclk));
	jdff dff_B_NHCck5hr7_0(.din(w_dff_B_WxdPq4aF7_0),.dout(w_dff_B_NHCck5hr7_0),.clk(gclk));
	jdff dff_B_C8rDAqsc1_0(.din(w_dff_B_NHCck5hr7_0),.dout(w_dff_B_C8rDAqsc1_0),.clk(gclk));
	jdff dff_B_0ap6VvY94_0(.din(w_dff_B_C8rDAqsc1_0),.dout(w_dff_B_0ap6VvY94_0),.clk(gclk));
	jdff dff_B_YK1nnchb2_0(.din(w_dff_B_0ap6VvY94_0),.dout(w_dff_B_YK1nnchb2_0),.clk(gclk));
	jdff dff_B_vX0LSfgT8_0(.din(w_dff_B_YK1nnchb2_0),.dout(w_dff_B_vX0LSfgT8_0),.clk(gclk));
	jdff dff_B_6kJ1aIoB0_0(.din(w_dff_B_vX0LSfgT8_0),.dout(w_dff_B_6kJ1aIoB0_0),.clk(gclk));
	jdff dff_B_WPfkaipq5_0(.din(w_dff_B_6kJ1aIoB0_0),.dout(w_dff_B_WPfkaipq5_0),.clk(gclk));
	jdff dff_B_gGWEjK925_0(.din(w_dff_B_WPfkaipq5_0),.dout(w_dff_B_gGWEjK925_0),.clk(gclk));
	jdff dff_B_KOiFVQEN6_0(.din(w_dff_B_gGWEjK925_0),.dout(w_dff_B_KOiFVQEN6_0),.clk(gclk));
	jdff dff_B_0wk7J7iX9_0(.din(w_dff_B_KOiFVQEN6_0),.dout(w_dff_B_0wk7J7iX9_0),.clk(gclk));
	jdff dff_B_sZlIW0VD8_0(.din(w_dff_B_0wk7J7iX9_0),.dout(w_dff_B_sZlIW0VD8_0),.clk(gclk));
	jdff dff_B_j3rZniwi8_0(.din(w_dff_B_sZlIW0VD8_0),.dout(w_dff_B_j3rZniwi8_0),.clk(gclk));
	jdff dff_B_uq0MPfYp7_0(.din(w_dff_B_j3rZniwi8_0),.dout(w_dff_B_uq0MPfYp7_0),.clk(gclk));
	jdff dff_B_vDw7soEk5_0(.din(w_dff_B_uq0MPfYp7_0),.dout(w_dff_B_vDw7soEk5_0),.clk(gclk));
	jdff dff_B_vZOAtpMZ1_0(.din(w_dff_B_vDw7soEk5_0),.dout(w_dff_B_vZOAtpMZ1_0),.clk(gclk));
	jdff dff_B_d5vIGQs41_0(.din(w_dff_B_vZOAtpMZ1_0),.dout(w_dff_B_d5vIGQs41_0),.clk(gclk));
	jdff dff_B_ZqXl24ZW1_1(.din(n1588),.dout(w_dff_B_ZqXl24ZW1_1),.clk(gclk));
	jdff dff_B_uC3bIeM93_1(.din(w_dff_B_ZqXl24ZW1_1),.dout(w_dff_B_uC3bIeM93_1),.clk(gclk));
	jdff dff_B_MWJj8SXT8_1(.din(w_dff_B_uC3bIeM93_1),.dout(w_dff_B_MWJj8SXT8_1),.clk(gclk));
	jdff dff_B_XZAIPmcT9_1(.din(w_dff_B_MWJj8SXT8_1),.dout(w_dff_B_XZAIPmcT9_1),.clk(gclk));
	jdff dff_B_xleXgPAa7_1(.din(w_dff_B_XZAIPmcT9_1),.dout(w_dff_B_xleXgPAa7_1),.clk(gclk));
	jdff dff_B_lMMR4Cfn6_1(.din(w_dff_B_xleXgPAa7_1),.dout(w_dff_B_lMMR4Cfn6_1),.clk(gclk));
	jdff dff_B_CFUSpfow9_1(.din(w_dff_B_lMMR4Cfn6_1),.dout(w_dff_B_CFUSpfow9_1),.clk(gclk));
	jdff dff_B_tiupQjuw9_1(.din(w_dff_B_CFUSpfow9_1),.dout(w_dff_B_tiupQjuw9_1),.clk(gclk));
	jdff dff_B_bScsnL8T1_1(.din(n1655),.dout(w_dff_B_bScsnL8T1_1),.clk(gclk));
	jdff dff_B_ibd6MUij4_1(.din(w_dff_B_bScsnL8T1_1),.dout(w_dff_B_ibd6MUij4_1),.clk(gclk));
	jdff dff_A_5n6wNkML4_2(.dout(w_n588_0[2]),.din(w_dff_A_5n6wNkML4_2),.clk(gclk));
	jdff dff_A_7ToaC0wk1_2(.dout(w_dff_A_5n6wNkML4_2),.din(w_dff_A_7ToaC0wk1_2),.clk(gclk));
	jdff dff_A_P4SEEAWN6_1(.dout(w_n1652_0[1]),.din(w_dff_A_P4SEEAWN6_1),.clk(gclk));
	jdff dff_B_CIh7LDlr1_0(.din(n1649),.dout(w_dff_B_CIh7LDlr1_0),.clk(gclk));
	jdff dff_B_FsANhX6v6_1(.din(n1645),.dout(w_dff_B_FsANhX6v6_1),.clk(gclk));
	jdff dff_B_K0LZ4egM2_1(.din(w_dff_B_FsANhX6v6_1),.dout(w_dff_B_K0LZ4egM2_1),.clk(gclk));
	jdff dff_B_DnPGAQ225_1(.din(w_dff_B_K0LZ4egM2_1),.dout(w_dff_B_DnPGAQ225_1),.clk(gclk));
	jdff dff_B_QfmQDYsv4_1(.din(w_dff_B_DnPGAQ225_1),.dout(w_dff_B_QfmQDYsv4_1),.clk(gclk));
	jdff dff_B_HtBxJ4xT0_1(.din(w_dff_B_QfmQDYsv4_1),.dout(w_dff_B_HtBxJ4xT0_1),.clk(gclk));
	jdff dff_B_mlib1XFp3_1(.din(n1638),.dout(w_dff_B_mlib1XFp3_1),.clk(gclk));
	jdff dff_B_cWMUahs32_1(.din(w_dff_B_mlib1XFp3_1),.dout(w_dff_B_cWMUahs32_1),.clk(gclk));
	jdff dff_B_LNpshacK4_0(.din(n1641),.dout(w_dff_B_LNpshacK4_0),.clk(gclk));
	jdff dff_B_d5zF6k0X1_0(.din(n1640),.dout(w_dff_B_d5zF6k0X1_0),.clk(gclk));
	jdff dff_A_psAXok7z0_1(.dout(w_n609_0[1]),.din(w_dff_A_psAXok7z0_1),.clk(gclk));
	jdff dff_A_GAH6Qt1h4_1(.dout(w_dff_A_psAXok7z0_1),.din(w_dff_A_GAH6Qt1h4_1),.clk(gclk));
	jdff dff_A_F8gxj0VY4_1(.dout(w_dff_A_GAH6Qt1h4_1),.din(w_dff_A_F8gxj0VY4_1),.clk(gclk));
	jdff dff_A_WSsWGxBs5_1(.dout(w_dff_A_F8gxj0VY4_1),.din(w_dff_A_WSsWGxBs5_1),.clk(gclk));
	jdff dff_A_hEztNyTD8_1(.dout(w_dff_A_WSsWGxBs5_1),.din(w_dff_A_hEztNyTD8_1),.clk(gclk));
	jdff dff_A_CXmnyfZQ8_1(.dout(w_dff_A_hEztNyTD8_1),.din(w_dff_A_CXmnyfZQ8_1),.clk(gclk));
	jdff dff_A_Jx6W1WJ93_1(.dout(w_dff_A_CXmnyfZQ8_1),.din(w_dff_A_Jx6W1WJ93_1),.clk(gclk));
	jdff dff_A_zLeIUgkS0_1(.dout(w_n962_0[1]),.din(w_dff_A_zLeIUgkS0_1),.clk(gclk));
	jdff dff_A_NN3yA7u52_1(.dout(w_dff_A_zLeIUgkS0_1),.din(w_dff_A_NN3yA7u52_1),.clk(gclk));
	jdff dff_A_eDMU0LZO7_1(.dout(w_dff_A_NN3yA7u52_1),.din(w_dff_A_eDMU0LZO7_1),.clk(gclk));
	jdff dff_A_xBIqZVoy4_1(.dout(w_dff_A_eDMU0LZO7_1),.din(w_dff_A_xBIqZVoy4_1),.clk(gclk));
	jdff dff_A_HOxDukn92_1(.dout(w_dff_A_xBIqZVoy4_1),.din(w_dff_A_HOxDukn92_1),.clk(gclk));
	jdff dff_A_m7ftWT6w2_1(.dout(w_dff_A_HOxDukn92_1),.din(w_dff_A_m7ftWT6w2_1),.clk(gclk));
	jdff dff_B_85atRmAC4_2(.din(n962),.dout(w_dff_B_85atRmAC4_2),.clk(gclk));
	jdff dff_A_wMsnKMJ88_2(.dout(w_n938_0[2]),.din(w_dff_A_wMsnKMJ88_2),.clk(gclk));
	jdff dff_A_uoeP3skZ5_2(.dout(w_dff_A_wMsnKMJ88_2),.din(w_dff_A_uoeP3skZ5_2),.clk(gclk));
	jdff dff_A_yNVUy8E48_2(.dout(w_dff_A_uoeP3skZ5_2),.din(w_dff_A_yNVUy8E48_2),.clk(gclk));
	jdff dff_A_WbG1ljAS0_2(.dout(w_dff_A_yNVUy8E48_2),.din(w_dff_A_WbG1ljAS0_2),.clk(gclk));
	jdff dff_A_BN6ZpJxo8_2(.dout(w_dff_A_WbG1ljAS0_2),.din(w_dff_A_BN6ZpJxo8_2),.clk(gclk));
	jdff dff_B_Geu16LN10_1(.din(n707),.dout(w_dff_B_Geu16LN10_1),.clk(gclk));
	jdff dff_B_A6Ci5U740_1(.din(w_dff_B_Geu16LN10_1),.dout(w_dff_B_A6Ci5U740_1),.clk(gclk));
	jdff dff_B_18LzI1ED4_1(.din(w_dff_B_A6Ci5U740_1),.dout(w_dff_B_18LzI1ED4_1),.clk(gclk));
	jdff dff_B_ZWyfy5xQ9_1(.din(n708),.dout(w_dff_B_ZWyfy5xQ9_1),.clk(gclk));
	jdff dff_B_6oCEeYCx3_1(.din(w_dff_B_ZWyfy5xQ9_1),.dout(w_dff_B_6oCEeYCx3_1),.clk(gclk));
	jdff dff_A_gGvEFFCe5_1(.dout(w_n713_0[1]),.din(w_dff_A_gGvEFFCe5_1),.clk(gclk));
	jdff dff_A_i3QuapY35_1(.dout(w_dff_A_gGvEFFCe5_1),.din(w_dff_A_i3QuapY35_1),.clk(gclk));
	jdff dff_A_rfj2WLJI8_1(.dout(w_dff_A_i3QuapY35_1),.din(w_dff_A_rfj2WLJI8_1),.clk(gclk));
	jdff dff_A_ROlElPWS5_1(.dout(w_dff_A_rfj2WLJI8_1),.din(w_dff_A_ROlElPWS5_1),.clk(gclk));
	jdff dff_A_RQf5Tvz91_1(.dout(w_dff_A_ROlElPWS5_1),.din(w_dff_A_RQf5Tvz91_1),.clk(gclk));
	jdff dff_A_kLRNieab5_1(.dout(w_dff_A_RQf5Tvz91_1),.din(w_dff_A_kLRNieab5_1),.clk(gclk));
	jdff dff_A_fNtva72h0_1(.dout(w_dff_A_kLRNieab5_1),.din(w_dff_A_fNtva72h0_1),.clk(gclk));
	jdff dff_A_aglSFw1X4_0(.dout(w_n710_0[0]),.din(w_dff_A_aglSFw1X4_0),.clk(gclk));
	jdff dff_A_tCBNZm7E8_0(.dout(w_dff_A_aglSFw1X4_0),.din(w_dff_A_tCBNZm7E8_0),.clk(gclk));
	jdff dff_A_HHfVC22M3_0(.dout(w_dff_A_tCBNZm7E8_0),.din(w_dff_A_HHfVC22M3_0),.clk(gclk));
	jdff dff_A_066BfeTR1_0(.dout(w_dff_A_HHfVC22M3_0),.din(w_dff_A_066BfeTR1_0),.clk(gclk));
	jdff dff_A_Z1WB7ngR6_0(.dout(w_dff_A_066BfeTR1_0),.din(w_dff_A_Z1WB7ngR6_0),.clk(gclk));
	jdff dff_A_RyoELTp12_0(.dout(w_dff_A_Z1WB7ngR6_0),.din(w_dff_A_RyoELTp12_0),.clk(gclk));
	jdff dff_A_ZML9gGz17_0(.dout(w_dff_A_RyoELTp12_0),.din(w_dff_A_ZML9gGz17_0),.clk(gclk));
	jdff dff_A_UVhmSwRi2_0(.dout(w_dff_A_ZML9gGz17_0),.din(w_dff_A_UVhmSwRi2_0),.clk(gclk));
	jdff dff_A_zw6mIUv48_0(.dout(w_n597_0[0]),.din(w_dff_A_zw6mIUv48_0),.clk(gclk));
	jdff dff_A_4TkgQVI47_0(.dout(w_dff_A_zw6mIUv48_0),.din(w_dff_A_4TkgQVI47_0),.clk(gclk));
	jdff dff_A_W8pUR8FL8_0(.dout(w_dff_A_4TkgQVI47_0),.din(w_dff_A_W8pUR8FL8_0),.clk(gclk));
	jdff dff_A_AcJYINxx4_0(.dout(w_dff_A_W8pUR8FL8_0),.din(w_dff_A_AcJYINxx4_0),.clk(gclk));
	jdff dff_A_ExtVVazX9_0(.dout(w_dff_A_AcJYINxx4_0),.din(w_dff_A_ExtVVazX9_0),.clk(gclk));
	jdff dff_A_GFxP12ni9_0(.dout(w_n496_1[0]),.din(w_dff_A_GFxP12ni9_0),.clk(gclk));
	jdff dff_A_07Q4LIuX7_0(.dout(w_dff_A_GFxP12ni9_0),.din(w_dff_A_07Q4LIuX7_0),.clk(gclk));
	jdff dff_A_1LHGQENa9_0(.dout(w_n1637_0[0]),.din(w_dff_A_1LHGQENa9_0),.clk(gclk));
	jdff dff_A_ufo0E6sZ2_0(.dout(w_dff_A_1LHGQENa9_0),.din(w_dff_A_ufo0E6sZ2_0),.clk(gclk));
	jdff dff_B_FpG3zss28_2(.din(n1637),.dout(w_dff_B_FpG3zss28_2),.clk(gclk));
	jdff dff_B_Y8KYvAO46_2(.din(w_dff_B_FpG3zss28_2),.dout(w_dff_B_Y8KYvAO46_2),.clk(gclk));
	jdff dff_A_bZFrhxba1_1(.dout(w_n608_0[1]),.din(w_dff_A_bZFrhxba1_1),.clk(gclk));
	jdff dff_A_ieECgFmf2_1(.dout(w_dff_A_bZFrhxba1_1),.din(w_dff_A_ieECgFmf2_1),.clk(gclk));
	jdff dff_A_aiAFb0Bb7_1(.dout(w_dff_A_ieECgFmf2_1),.din(w_dff_A_aiAFb0Bb7_1),.clk(gclk));
	jdff dff_A_WU2MSFyF2_1(.dout(w_dff_A_aiAFb0Bb7_1),.din(w_dff_A_WU2MSFyF2_1),.clk(gclk));
	jdff dff_A_OCMk77wF2_1(.dout(w_dff_A_WU2MSFyF2_1),.din(w_dff_A_OCMk77wF2_1),.clk(gclk));
	jdff dff_A_DpDS1xpR7_1(.dout(w_dff_A_OCMk77wF2_1),.din(w_dff_A_DpDS1xpR7_1),.clk(gclk));
	jdff dff_A_tMLLDGjh3_1(.dout(w_dff_A_DpDS1xpR7_1),.din(w_dff_A_tMLLDGjh3_1),.clk(gclk));
	jdff dff_A_DcebTOye1_1(.dout(w_dff_A_tMLLDGjh3_1),.din(w_dff_A_DcebTOye1_1),.clk(gclk));
	jdff dff_A_LtRWGmHs8_1(.dout(w_dff_A_DcebTOye1_1),.din(w_dff_A_LtRWGmHs8_1),.clk(gclk));
	jdff dff_A_RpA6Tcj95_1(.dout(w_dff_A_LtRWGmHs8_1),.din(w_dff_A_RpA6Tcj95_1),.clk(gclk));
	jdff dff_A_T3e2k0WO5_2(.dout(w_n608_0[2]),.din(w_dff_A_T3e2k0WO5_2),.clk(gclk));
	jdff dff_B_D4fOFHL32_0(.din(n606),.dout(w_dff_B_D4fOFHL32_0),.clk(gclk));
	jdff dff_B_WRS1WKld4_1(.din(G217),.dout(w_dff_B_WRS1WKld4_1),.clk(gclk));
	jdff dff_A_hBJz7Zz76_0(.dout(w_n592_0[0]),.din(w_dff_A_hBJz7Zz76_0),.clk(gclk));
	jdff dff_A_eLuM00936_2(.dout(w_n592_0[2]),.din(w_dff_A_eLuM00936_2),.clk(gclk));
	jdff dff_A_SvbF4Bdf8_2(.dout(w_dff_A_eLuM00936_2),.din(w_dff_A_SvbF4Bdf8_2),.clk(gclk));
	jdff dff_A_1NICf9Y90_2(.dout(w_dff_A_SvbF4Bdf8_2),.din(w_dff_A_1NICf9Y90_2),.clk(gclk));
	jdff dff_A_aRbml7jY4_2(.dout(w_dff_A_1NICf9Y90_2),.din(w_dff_A_aRbml7jY4_2),.clk(gclk));
	jdff dff_B_KjkXO6uF3_1(.din(n589),.dout(w_dff_B_KjkXO6uF3_1),.clk(gclk));
	jdff dff_B_2HPg2p4d3_1(.din(G209),.dout(w_dff_B_2HPg2p4d3_1),.clk(gclk));
	jdff dff_A_soHz0zdW4_0(.dout(w_n602_0[0]),.din(w_dff_A_soHz0zdW4_0),.clk(gclk));
	jdff dff_A_BuuBg4Y98_0(.dout(w_n711_0[0]),.din(w_dff_A_BuuBg4Y98_0),.clk(gclk));
	jdff dff_A_vvtsNuvE8_0(.dout(w_dff_A_BuuBg4Y98_0),.din(w_dff_A_vvtsNuvE8_0),.clk(gclk));
	jdff dff_A_tHGNU3MT1_2(.dout(w_n954_0[2]),.din(w_dff_A_tHGNU3MT1_2),.clk(gclk));
	jdff dff_A_aGjrNP4F6_2(.dout(w_dff_A_tHGNU3MT1_2),.din(w_dff_A_aGjrNP4F6_2),.clk(gclk));
	jdff dff_A_MmMhsMmR4_2(.dout(w_dff_A_aGjrNP4F6_2),.din(w_dff_A_MmMhsMmR4_2),.clk(gclk));
	jdff dff_A_1zbcjddR5_2(.dout(w_dff_A_MmMhsMmR4_2),.din(w_dff_A_1zbcjddR5_2),.clk(gclk));
	jdff dff_A_aMve6OvM1_2(.dout(w_dff_A_1zbcjddR5_2),.din(w_dff_A_aMve6OvM1_2),.clk(gclk));
	jdff dff_A_ZZpAA2XQ4_2(.dout(w_dff_A_aMve6OvM1_2),.din(w_dff_A_ZZpAA2XQ4_2),.clk(gclk));
	jdff dff_A_ccdkAcaE8_2(.dout(w_dff_A_ZZpAA2XQ4_2),.din(w_dff_A_ccdkAcaE8_2),.clk(gclk));
	jdff dff_B_bA6fv7q99_2(.din(n1633),.dout(w_dff_B_bA6fv7q99_2),.clk(gclk));
	jdff dff_A_Hkcjyptd3_1(.dout(w_n709_0[1]),.din(w_dff_A_Hkcjyptd3_1),.clk(gclk));
	jdff dff_B_4gpgBaTR1_0(.din(n600),.dout(w_dff_B_4gpgBaTR1_0),.clk(gclk));
	jdff dff_B_RwubvhTj3_1(.din(G225),.dout(w_dff_B_RwubvhTj3_1),.clk(gclk));
	jdff dff_B_vL2FhdQC8_0(.din(n595),.dout(w_dff_B_vL2FhdQC8_0),.clk(gclk));
	jdff dff_B_cgsVAW2z9_1(.din(G233),.dout(w_dff_B_cgsVAW2z9_1),.clk(gclk));
	jdff dff_A_Bq7f18HZ2_1(.dout(w_n703_0[1]),.din(w_dff_A_Bq7f18HZ2_1),.clk(gclk));
	jdff dff_A_mHZ70Jib2_0(.dout(w_n685_0[0]),.din(w_dff_A_mHZ70Jib2_0),.clk(gclk));
	jdff dff_A_m5S8r6zo1_0(.dout(w_dff_A_mHZ70Jib2_0),.din(w_dff_A_m5S8r6zo1_0),.clk(gclk));
	jdff dff_B_DMsN892w7_2(.din(n685),.dout(w_dff_B_DMsN892w7_2),.clk(gclk));
	jdff dff_B_xHtQRvQv8_2(.din(w_dff_B_DMsN892w7_2),.dout(w_dff_B_xHtQRvQv8_2),.clk(gclk));
	jdff dff_B_FTkfTvPN9_2(.din(w_dff_B_xHtQRvQv8_2),.dout(w_dff_B_FTkfTvPN9_2),.clk(gclk));
	jdff dff_A_kz7MEoVC4_0(.dout(w_n684_0[0]),.din(w_dff_A_kz7MEoVC4_0),.clk(gclk));
	jdff dff_A_nvuB8LKZ9_0(.dout(w_dff_A_kz7MEoVC4_0),.din(w_dff_A_nvuB8LKZ9_0),.clk(gclk));
	jdff dff_A_0oBK8ZAp0_0(.dout(w_dff_A_nvuB8LKZ9_0),.din(w_dff_A_0oBK8ZAp0_0),.clk(gclk));
	jdff dff_A_N5RCJTb54_0(.dout(w_dff_A_0oBK8ZAp0_0),.din(w_dff_A_N5RCJTb54_0),.clk(gclk));
	jdff dff_A_URK2xtwG4_1(.dout(w_n682_0[1]),.din(w_dff_A_URK2xtwG4_1),.clk(gclk));
	jdff dff_A_rEhQI14U6_1(.dout(w_dff_A_URK2xtwG4_1),.din(w_dff_A_rEhQI14U6_1),.clk(gclk));
	jdff dff_A_LxSrrlcH4_1(.dout(w_dff_A_rEhQI14U6_1),.din(w_dff_A_LxSrrlcH4_1),.clk(gclk));
	jdff dff_A_KeuITP3b5_1(.dout(w_dff_A_LxSrrlcH4_1),.din(w_dff_A_KeuITP3b5_1),.clk(gclk));
	jdff dff_A_qF7txXay8_1(.dout(w_dff_A_KeuITP3b5_1),.din(w_dff_A_qF7txXay8_1),.clk(gclk));
	jdff dff_A_5USy8GVJ0_1(.dout(w_dff_A_qF7txXay8_1),.din(w_dff_A_5USy8GVJ0_1),.clk(gclk));
	jdff dff_A_lJZaxkb85_2(.dout(w_n682_0[2]),.din(w_dff_A_lJZaxkb85_2),.clk(gclk));
	jdff dff_A_xW9fUiXb0_2(.dout(w_dff_A_lJZaxkb85_2),.din(w_dff_A_xW9fUiXb0_2),.clk(gclk));
	jdff dff_A_QPI551Ni1_2(.dout(w_dff_A_xW9fUiXb0_2),.din(w_dff_A_QPI551Ni1_2),.clk(gclk));
	jdff dff_A_rfz3GYIR9_2(.dout(w_dff_A_QPI551Ni1_2),.din(w_dff_A_rfz3GYIR9_2),.clk(gclk));
	jdff dff_A_olY8EaMS8_2(.dout(w_dff_A_rfz3GYIR9_2),.din(w_dff_A_olY8EaMS8_2),.clk(gclk));
	jdff dff_A_5VPYhO5W0_2(.dout(w_dff_A_olY8EaMS8_2),.din(w_dff_A_5VPYhO5W0_2),.clk(gclk));
	jdff dff_B_nyBQTdjM8_0(.din(n1630),.dout(w_dff_B_nyBQTdjM8_0),.clk(gclk));
	jdff dff_B_6PRfqFmm3_0(.din(w_dff_B_nyBQTdjM8_0),.dout(w_dff_B_6PRfqFmm3_0),.clk(gclk));
	jdff dff_B_E2p7tr5q6_0(.din(w_dff_B_6PRfqFmm3_0),.dout(w_dff_B_E2p7tr5q6_0),.clk(gclk));
	jdff dff_B_nbXMw3Mw3_0(.din(w_dff_B_E2p7tr5q6_0),.dout(w_dff_B_nbXMw3Mw3_0),.clk(gclk));
	jdff dff_B_2cukDi5m9_0(.din(w_dff_B_nbXMw3Mw3_0),.dout(w_dff_B_2cukDi5m9_0),.clk(gclk));
	jdff dff_B_9tz4d4xd9_0(.din(w_dff_B_2cukDi5m9_0),.dout(w_dff_B_9tz4d4xd9_0),.clk(gclk));
	jdff dff_B_tBGgbLg64_0(.din(w_dff_B_9tz4d4xd9_0),.dout(w_dff_B_tBGgbLg64_0),.clk(gclk));
	jdff dff_B_SOO4Pp8b8_0(.din(w_dff_B_tBGgbLg64_0),.dout(w_dff_B_SOO4Pp8b8_0),.clk(gclk));
	jdff dff_B_Kf66Vzf82_0(.din(w_dff_B_SOO4Pp8b8_0),.dout(w_dff_B_Kf66Vzf82_0),.clk(gclk));
	jdff dff_B_2psLhj9J6_0(.din(n1628),.dout(w_dff_B_2psLhj9J6_0),.clk(gclk));
	jdff dff_B_saGac2ra0_0(.din(w_dff_B_2psLhj9J6_0),.dout(w_dff_B_saGac2ra0_0),.clk(gclk));
	jdff dff_B_UNIAtMf36_1(.din(n1625),.dout(w_dff_B_UNIAtMf36_1),.clk(gclk));
	jdff dff_B_9OsZINS98_1(.din(n1623),.dout(w_dff_B_9OsZINS98_1),.clk(gclk));
	jdff dff_B_7lVXvREL6_1(.din(w_dff_B_9OsZINS98_1),.dout(w_dff_B_7lVXvREL6_1),.clk(gclk));
	jdff dff_A_iKgtqary5_0(.dout(w_n1618_0[0]),.din(w_dff_A_iKgtqary5_0),.clk(gclk));
	jdff dff_A_pDMn4PWS6_0(.dout(w_dff_A_iKgtqary5_0),.din(w_dff_A_pDMn4PWS6_0),.clk(gclk));
	jdff dff_B_TGZRu1Wg8_2(.din(n1618),.dout(w_dff_B_TGZRu1Wg8_2),.clk(gclk));
	jdff dff_B_9t6qxJNc1_2(.din(w_dff_B_TGZRu1Wg8_2),.dout(w_dff_B_9t6qxJNc1_2),.clk(gclk));
	jdff dff_B_rrJ8SN4V1_2(.din(w_dff_B_9t6qxJNc1_2),.dout(w_dff_B_rrJ8SN4V1_2),.clk(gclk));
	jdff dff_B_GDBc4ZsU0_2(.din(w_dff_B_rrJ8SN4V1_2),.dout(w_dff_B_GDBc4ZsU0_2),.clk(gclk));
	jdff dff_B_X4yL09Gx8_2(.din(w_dff_B_GDBc4ZsU0_2),.dout(w_dff_B_X4yL09Gx8_2),.clk(gclk));
	jdff dff_B_uYtmjByw1_2(.din(w_dff_B_X4yL09Gx8_2),.dout(w_dff_B_uYtmjByw1_2),.clk(gclk));
	jdff dff_B_nXFOZ9vY9_2(.din(w_dff_B_uYtmjByw1_2),.dout(w_dff_B_nXFOZ9vY9_2),.clk(gclk));
	jdff dff_B_MLAzN9QG9_2(.din(w_dff_B_nXFOZ9vY9_2),.dout(w_dff_B_MLAzN9QG9_2),.clk(gclk));
	jdff dff_B_Z8maTnec1_2(.din(w_dff_B_MLAzN9QG9_2),.dout(w_dff_B_Z8maTnec1_2),.clk(gclk));
	jdff dff_B_eMhbkInQ9_2(.din(w_dff_B_Z8maTnec1_2),.dout(w_dff_B_eMhbkInQ9_2),.clk(gclk));
	jdff dff_B_4180wa9x2_2(.din(w_dff_B_eMhbkInQ9_2),.dout(w_dff_B_4180wa9x2_2),.clk(gclk));
	jdff dff_B_r7JxUxaj9_2(.din(w_dff_B_4180wa9x2_2),.dout(w_dff_B_r7JxUxaj9_2),.clk(gclk));
	jdff dff_A_4uMTWYY66_0(.dout(w_G1497_0[0]),.din(w_dff_A_4uMTWYY66_0),.clk(gclk));
	jdff dff_A_teNYVAXO2_0(.dout(w_dff_A_4uMTWYY66_0),.din(w_dff_A_teNYVAXO2_0),.clk(gclk));
	jdff dff_A_85z2pYkP1_0(.dout(w_dff_A_teNYVAXO2_0),.din(w_dff_A_85z2pYkP1_0),.clk(gclk));
	jdff dff_A_Zur9GXe36_0(.dout(w_dff_A_85z2pYkP1_0),.din(w_dff_A_Zur9GXe36_0),.clk(gclk));
	jdff dff_A_skKNapTl4_0(.dout(w_dff_A_Zur9GXe36_0),.din(w_dff_A_skKNapTl4_0),.clk(gclk));
	jdff dff_A_UBVNAlgo3_0(.dout(w_dff_A_skKNapTl4_0),.din(w_dff_A_UBVNAlgo3_0),.clk(gclk));
	jdff dff_A_N8BJuBMI5_0(.dout(w_dff_A_UBVNAlgo3_0),.din(w_dff_A_N8BJuBMI5_0),.clk(gclk));
	jdff dff_A_Yrw8BFI23_0(.dout(w_dff_A_N8BJuBMI5_0),.din(w_dff_A_Yrw8BFI23_0),.clk(gclk));
	jdff dff_A_gqBH0egq3_0(.dout(w_dff_A_Yrw8BFI23_0),.din(w_dff_A_gqBH0egq3_0),.clk(gclk));
	jdff dff_A_83IIzFRi1_0(.dout(w_dff_A_gqBH0egq3_0),.din(w_dff_A_83IIzFRi1_0),.clk(gclk));
	jdff dff_A_mfaNR6rt2_0(.dout(w_dff_A_83IIzFRi1_0),.din(w_dff_A_mfaNR6rt2_0),.clk(gclk));
	jdff dff_A_TEOkXkTo7_0(.dout(w_dff_A_mfaNR6rt2_0),.din(w_dff_A_TEOkXkTo7_0),.clk(gclk));
	jdff dff_A_h9CeMrqq8_0(.dout(w_dff_A_TEOkXkTo7_0),.din(w_dff_A_h9CeMrqq8_0),.clk(gclk));
	jdff dff_A_0lGGwlJU3_0(.dout(w_dff_A_h9CeMrqq8_0),.din(w_dff_A_0lGGwlJU3_0),.clk(gclk));
	jdff dff_A_ezjoubcI2_0(.dout(w_dff_A_0lGGwlJU3_0),.din(w_dff_A_ezjoubcI2_0),.clk(gclk));
	jdff dff_A_cPARA59N3_1(.dout(w_G1497_0[1]),.din(w_dff_A_cPARA59N3_1),.clk(gclk));
	jdff dff_A_R1FXdyIR7_1(.dout(w_dff_A_cPARA59N3_1),.din(w_dff_A_R1FXdyIR7_1),.clk(gclk));
	jdff dff_A_1njxCRKP6_1(.dout(w_dff_A_R1FXdyIR7_1),.din(w_dff_A_1njxCRKP6_1),.clk(gclk));
	jdff dff_A_p9fMp0Yu5_1(.dout(w_dff_A_1njxCRKP6_1),.din(w_dff_A_p9fMp0Yu5_1),.clk(gclk));
	jdff dff_A_98tYvckP5_1(.dout(w_dff_A_p9fMp0Yu5_1),.din(w_dff_A_98tYvckP5_1),.clk(gclk));
	jdff dff_A_rkkqxecX0_1(.dout(w_dff_A_98tYvckP5_1),.din(w_dff_A_rkkqxecX0_1),.clk(gclk));
	jdff dff_A_wEkh6VZ99_1(.dout(w_dff_A_rkkqxecX0_1),.din(w_dff_A_wEkh6VZ99_1),.clk(gclk));
	jdff dff_A_pv1zHmMR5_1(.dout(w_dff_A_wEkh6VZ99_1),.din(w_dff_A_pv1zHmMR5_1),.clk(gclk));
	jdff dff_A_qmZQARQv9_1(.dout(w_dff_A_pv1zHmMR5_1),.din(w_dff_A_qmZQARQv9_1),.clk(gclk));
	jdff dff_A_kOZ4e30O9_1(.dout(w_dff_A_qmZQARQv9_1),.din(w_dff_A_kOZ4e30O9_1),.clk(gclk));
	jdff dff_A_HGOM2LJm0_1(.dout(w_dff_A_kOZ4e30O9_1),.din(w_dff_A_HGOM2LJm0_1),.clk(gclk));
	jdff dff_A_EP0AG1Mv3_1(.dout(w_dff_A_HGOM2LJm0_1),.din(w_dff_A_EP0AG1Mv3_1),.clk(gclk));
	jdff dff_B_1UoxQOPg5_1(.din(n1600),.dout(w_dff_B_1UoxQOPg5_1),.clk(gclk));
	jdff dff_B_gjBGjyHe4_1(.din(w_dff_B_1UoxQOPg5_1),.dout(w_dff_B_gjBGjyHe4_1),.clk(gclk));
	jdff dff_B_3qSVlTZF9_0(.din(n1614),.dout(w_dff_B_3qSVlTZF9_0),.clk(gclk));
	jdff dff_B_H6WJMbzw8_0(.din(w_dff_B_3qSVlTZF9_0),.dout(w_dff_B_H6WJMbzw8_0),.clk(gclk));
	jdff dff_B_1WSuVNJs3_0(.din(w_dff_B_H6WJMbzw8_0),.dout(w_dff_B_1WSuVNJs3_0),.clk(gclk));
	jdff dff_B_s5FvmlJb1_0(.din(w_dff_B_1WSuVNJs3_0),.dout(w_dff_B_s5FvmlJb1_0),.clk(gclk));
	jdff dff_A_jRI9t6sW0_0(.dout(w_n1613_0[0]),.din(w_dff_A_jRI9t6sW0_0),.clk(gclk));
	jdff dff_A_FcJRNiM37_0(.dout(w_dff_A_jRI9t6sW0_0),.din(w_dff_A_FcJRNiM37_0),.clk(gclk));
	jdff dff_A_pY7wjSMf9_0(.dout(w_n865_0[0]),.din(w_dff_A_pY7wjSMf9_0),.clk(gclk));
	jdff dff_A_xpLZ6p1m0_0(.dout(w_dff_A_pY7wjSMf9_0),.din(w_dff_A_xpLZ6p1m0_0),.clk(gclk));
	jdff dff_A_NENDBLe24_0(.dout(w_dff_A_xpLZ6p1m0_0),.din(w_dff_A_NENDBLe24_0),.clk(gclk));
	jdff dff_A_PPDwXgPR8_0(.dout(w_dff_A_NENDBLe24_0),.din(w_dff_A_PPDwXgPR8_0),.clk(gclk));
	jdff dff_A_hfb1qTpJ0_2(.dout(w_n865_0[2]),.din(w_dff_A_hfb1qTpJ0_2),.clk(gclk));
	jdff dff_A_yIo3iudj5_2(.dout(w_dff_A_hfb1qTpJ0_2),.din(w_dff_A_yIo3iudj5_2),.clk(gclk));
	jdff dff_A_VkK6Io6I5_2(.dout(w_dff_A_yIo3iudj5_2),.din(w_dff_A_VkK6Io6I5_2),.clk(gclk));
	jdff dff_A_WL1htVC61_2(.dout(w_dff_A_VkK6Io6I5_2),.din(w_dff_A_WL1htVC61_2),.clk(gclk));
	jdff dff_A_oJqkeyL69_2(.dout(w_dff_A_WL1htVC61_2),.din(w_dff_A_oJqkeyL69_2),.clk(gclk));
	jdff dff_A_SdP4WpJM4_1(.dout(w_n587_0[1]),.din(w_dff_A_SdP4WpJM4_1),.clk(gclk));
	jdff dff_A_0XO0nWKt9_1(.dout(w_dff_A_SdP4WpJM4_1),.din(w_dff_A_0XO0nWKt9_1),.clk(gclk));
	jdff dff_A_2M7lTDwp8_1(.dout(w_dff_A_0XO0nWKt9_1),.din(w_dff_A_2M7lTDwp8_1),.clk(gclk));
	jdff dff_A_LMNkz2cr9_1(.dout(w_dff_A_2M7lTDwp8_1),.din(w_dff_A_LMNkz2cr9_1),.clk(gclk));
	jdff dff_B_fmvCkGY62_0(.din(n585),.dout(w_dff_B_fmvCkGY62_0),.clk(gclk));
	jdff dff_B_X5fR3mvU3_1(.din(G241),.dout(w_dff_B_X5fR3mvU3_1),.clk(gclk));
	jdff dff_B_GBYNEvny9_1(.din(n1601),.dout(w_dff_B_GBYNEvny9_1),.clk(gclk));
	jdff dff_B_fTIeKDWs3_1(.din(w_dff_B_GBYNEvny9_1),.dout(w_dff_B_fTIeKDWs3_1),.clk(gclk));
	jdff dff_B_SkzEZ1708_1(.din(w_dff_B_fTIeKDWs3_1),.dout(w_dff_B_SkzEZ1708_1),.clk(gclk));
	jdff dff_B_W85vc1fY2_1(.din(n1602),.dout(w_dff_B_W85vc1fY2_1),.clk(gclk));
	jdff dff_B_bYjTbIzm8_1(.din(w_dff_B_W85vc1fY2_1),.dout(w_dff_B_bYjTbIzm8_1),.clk(gclk));
	jdff dff_A_xnNU7dEY7_1(.dout(w_n687_0[1]),.din(w_dff_A_xnNU7dEY7_1),.clk(gclk));
	jdff dff_A_dSuVNv8h2_1(.dout(w_dff_A_xnNU7dEY7_1),.din(w_dff_A_dSuVNv8h2_1),.clk(gclk));
	jdff dff_A_64xSURsP6_1(.dout(w_dff_A_dSuVNv8h2_1),.din(w_dff_A_64xSURsP6_1),.clk(gclk));
	jdff dff_A_TvANIoqV8_1(.dout(w_n686_0[1]),.din(w_dff_A_TvANIoqV8_1),.clk(gclk));
	jdff dff_A_yyqZ9IIT8_1(.dout(w_dff_A_TvANIoqV8_1),.din(w_dff_A_yyqZ9IIT8_1),.clk(gclk));
	jdff dff_A_wgGvhUbi2_1(.dout(w_dff_A_yyqZ9IIT8_1),.din(w_dff_A_wgGvhUbi2_1),.clk(gclk));
	jdff dff_A_1VkHJzJt5_1(.dout(w_dff_A_wgGvhUbi2_1),.din(w_dff_A_1VkHJzJt5_1),.clk(gclk));
	jdff dff_A_O9Os1Fyr6_0(.dout(w_n581_0[0]),.din(w_dff_A_O9Os1Fyr6_0),.clk(gclk));
	jdff dff_A_wABGtHPL5_0(.dout(w_dff_A_O9Os1Fyr6_0),.din(w_dff_A_wABGtHPL5_0),.clk(gclk));
	jdff dff_A_E7y64BeT8_1(.dout(w_n579_1[1]),.din(w_dff_A_E7y64BeT8_1),.clk(gclk));
	jdff dff_A_rxH08Yi38_1(.dout(w_n579_0[1]),.din(w_dff_A_rxH08Yi38_1),.clk(gclk));
	jdff dff_A_jnfhIwPP8_2(.dout(w_n579_0[2]),.din(w_dff_A_jnfhIwPP8_2),.clk(gclk));
	jdff dff_A_KwXpfViK5_2(.dout(w_dff_A_jnfhIwPP8_2),.din(w_dff_A_KwXpfViK5_2),.clk(gclk));
	jdff dff_A_kTB2hiAI9_2(.dout(w_dff_A_KwXpfViK5_2),.din(w_dff_A_kTB2hiAI9_2),.clk(gclk));
	jdff dff_A_1OUAiVoj1_2(.dout(w_dff_A_kTB2hiAI9_2),.din(w_dff_A_1OUAiVoj1_2),.clk(gclk));
	jdff dff_B_U3UaKWHr1_0(.din(n577),.dout(w_dff_B_U3UaKWHr1_0),.clk(gclk));
	jdff dff_B_7BuA7NsW1_1(.din(G264),.dout(w_dff_B_7BuA7NsW1_1),.clk(gclk));
	jdff dff_A_2vTjOU3w6_1(.dout(w_n574_0[1]),.din(w_dff_A_2vTjOU3w6_1),.clk(gclk));
	jdff dff_A_iC3wlEyD1_1(.dout(w_dff_A_2vTjOU3w6_1),.din(w_dff_A_iC3wlEyD1_1),.clk(gclk));
	jdff dff_A_RRDptfXs3_0(.dout(w_n1599_0[0]),.din(w_dff_A_RRDptfXs3_0),.clk(gclk));
	jdff dff_A_8aoAnBKr2_0(.dout(w_dff_A_RRDptfXs3_0),.din(w_dff_A_8aoAnBKr2_0),.clk(gclk));
	jdff dff_B_90XiUeBv2_0(.din(n1598),.dout(w_dff_B_90XiUeBv2_0),.clk(gclk));
	jdff dff_B_7FjASU305_0(.din(n1597),.dout(w_dff_B_7FjASU305_0),.clk(gclk));
	jdff dff_B_xFYDrjga7_0(.din(n1589),.dout(w_dff_B_xFYDrjga7_0),.clk(gclk));
	jdff dff_A_3SbmSsG54_0(.dout(w_n573_0[0]),.din(w_dff_A_3SbmSsG54_0),.clk(gclk));
	jdff dff_A_iThb78dO1_1(.dout(w_n573_0[1]),.din(w_dff_A_iThb78dO1_1),.clk(gclk));
	jdff dff_A_0hLVK2JU2_1(.dout(w_dff_A_iThb78dO1_1),.din(w_dff_A_0hLVK2JU2_1),.clk(gclk));
	jdff dff_B_ZNUr6u3F5_1(.din(n691),.dout(w_dff_B_ZNUr6u3F5_1),.clk(gclk));
	jdff dff_A_OMQ6DNjv3_0(.dout(w_n695_0[0]),.din(w_dff_A_OMQ6DNjv3_0),.clk(gclk));
	jdff dff_A_YkubTpUK1_1(.dout(w_n695_0[1]),.din(w_dff_A_YkubTpUK1_1),.clk(gclk));
	jdff dff_A_jlXW2jXy4_1(.dout(w_n564_0[1]),.din(w_dff_A_jlXW2jXy4_1),.clk(gclk));
	jdff dff_B_2qOmZ1NT3_1(.din(G280),.dout(w_dff_B_2qOmZ1NT3_1),.clk(gclk));
	jdff dff_A_ASeZkNt49_0(.dout(w_n562_0[0]),.din(w_dff_A_ASeZkNt49_0),.clk(gclk));
	jdff dff_A_FyyMCPEK9_0(.dout(w_n692_0[0]),.din(w_dff_A_FyyMCPEK9_0),.clk(gclk));
	jdff dff_A_TQ7VFzdl0_1(.dout(w_n559_0[1]),.din(w_dff_A_TQ7VFzdl0_1),.clk(gclk));
	jdff dff_B_npbHaFo88_1(.din(G288),.dout(w_dff_B_npbHaFo88_1),.clk(gclk));
	jdff dff_A_IWEv4cNs6_0(.dout(w_n557_0[0]),.din(w_dff_A_IWEv4cNs6_0),.clk(gclk));
	jdff dff_A_U0oiwZ160_0(.dout(w_n690_0[0]),.din(w_dff_A_U0oiwZ160_0),.clk(gclk));
	jdff dff_A_VXalCOdH3_0(.dout(w_dff_A_U0oiwZ160_0),.din(w_dff_A_VXalCOdH3_0),.clk(gclk));
	jdff dff_A_ehmpgBWb6_1(.dout(w_n571_0[1]),.din(w_dff_A_ehmpgBWb6_1),.clk(gclk));
	jdff dff_B_5xHzJPFB5_1(.din(G272),.dout(w_dff_B_5xHzJPFB5_1),.clk(gclk));
	jdff dff_A_UsLowW160_0(.dout(w_n569_0[0]),.din(w_dff_A_UsLowW160_0),.clk(gclk));
	jdff dff_A_7TY8sx288_0(.dout(w_n485_1[0]),.din(w_dff_A_7TY8sx288_0),.clk(gclk));
	jdff dff_A_PEoHeZnd2_0(.dout(w_dff_A_7TY8sx288_0),.din(w_dff_A_PEoHeZnd2_0),.clk(gclk));
	jdff dff_B_9vqikBI63_0(.din(n1585),.dout(w_dff_B_9vqikBI63_0),.clk(gclk));
	jdff dff_B_qcI4xhpd3_1(.din(n1575),.dout(w_dff_B_qcI4xhpd3_1),.clk(gclk));
	jdff dff_B_1M5Qhs089_1(.din(w_dff_B_qcI4xhpd3_1),.dout(w_dff_B_1M5Qhs089_1),.clk(gclk));
	jdff dff_A_YTqdcaIL5_0(.dout(w_G210_2[0]),.din(w_dff_A_YTqdcaIL5_0),.clk(gclk));
	jdff dff_A_pNIdrQYI2_1(.dout(w_n451_0[1]),.din(w_dff_A_pNIdrQYI2_1),.clk(gclk));
	jdff dff_A_N1aipDxO8_1(.dout(w_dff_A_pNIdrQYI2_1),.din(w_dff_A_N1aipDxO8_1),.clk(gclk));
	jdff dff_B_MEJV5t838_3(.din(n451),.dout(w_dff_B_MEJV5t838_3),.clk(gclk));
	jdff dff_A_akd0nIm96_0(.dout(w_G457_1[0]),.din(w_dff_A_akd0nIm96_0),.clk(gclk));
	jdff dff_A_D4p2fYwl0_0(.dout(w_dff_A_akd0nIm96_0),.din(w_dff_A_D4p2fYwl0_0),.clk(gclk));
	jdff dff_A_HIrzIPQQ3_0(.dout(w_dff_A_D4p2fYwl0_0),.din(w_dff_A_HIrzIPQQ3_0),.clk(gclk));
	jdff dff_A_5NXR3OFP8_0(.dout(w_dff_A_HIrzIPQQ3_0),.din(w_dff_A_5NXR3OFP8_0),.clk(gclk));
	jdff dff_A_TT2Fd5ad6_1(.dout(w_G457_1[1]),.din(w_dff_A_TT2Fd5ad6_1),.clk(gclk));
	jdff dff_A_05JR57BF6_1(.dout(w_dff_A_TT2Fd5ad6_1),.din(w_dff_A_05JR57BF6_1),.clk(gclk));
	jdff dff_A_U8qclugG4_1(.dout(w_dff_A_05JR57BF6_1),.din(w_dff_A_U8qclugG4_1),.clk(gclk));
	jdff dff_A_92iJuFfX5_1(.dout(w_G457_0[1]),.din(w_dff_A_92iJuFfX5_1),.clk(gclk));
	jdff dff_A_dUzOfJsY5_1(.dout(w_dff_A_92iJuFfX5_1),.din(w_dff_A_dUzOfJsY5_1),.clk(gclk));
	jdff dff_A_oskN5ta20_1(.dout(w_dff_A_dUzOfJsY5_1),.din(w_dff_A_oskN5ta20_1),.clk(gclk));
	jdff dff_A_IGdw9cT14_2(.dout(w_G457_0[2]),.din(w_dff_A_IGdw9cT14_2),.clk(gclk));
	jdff dff_A_ie5uQqXi4_2(.dout(w_dff_A_IGdw9cT14_2),.din(w_dff_A_ie5uQqXi4_2),.clk(gclk));
	jdff dff_A_atSMxOPA5_2(.dout(w_dff_A_ie5uQqXi4_2),.din(w_dff_A_atSMxOPA5_2),.clk(gclk));
	jdff dff_A_2y2w50oe2_2(.dout(w_dff_A_atSMxOPA5_2),.din(w_dff_A_2y2w50oe2_2),.clk(gclk));
	jdff dff_A_kvwfYG590_2(.dout(w_G210_0[2]),.din(w_dff_A_kvwfYG590_2),.clk(gclk));
	jdff dff_B_9Ce1NkLg6_1(.din(n1570),.dout(w_dff_B_9Ce1NkLg6_1),.clk(gclk));
	jdff dff_A_6Kekg5Mn7_0(.dout(w_n509_0[0]),.din(w_dff_A_6Kekg5Mn7_0),.clk(gclk));
	jdff dff_A_ZABLnUU79_1(.dout(w_n509_0[1]),.din(w_dff_A_ZABLnUU79_1),.clk(gclk));
	jdff dff_A_T9ZByXAe4_1(.dout(w_dff_A_ZABLnUU79_1),.din(w_dff_A_T9ZByXAe4_1),.clk(gclk));
	jdff dff_B_tNG1fmo45_3(.din(n509),.dout(w_dff_B_tNG1fmo45_3),.clk(gclk));
	jdff dff_A_vk3DHFRB9_0(.dout(w_G468_1[0]),.din(w_dff_A_vk3DHFRB9_0),.clk(gclk));
	jdff dff_A_KrTo8HK52_0(.dout(w_dff_A_vk3DHFRB9_0),.din(w_dff_A_KrTo8HK52_0),.clk(gclk));
	jdff dff_A_3EyJadJB5_0(.dout(w_dff_A_KrTo8HK52_0),.din(w_dff_A_3EyJadJB5_0),.clk(gclk));
	jdff dff_A_YYWsJkFt2_0(.dout(w_dff_A_3EyJadJB5_0),.din(w_dff_A_YYWsJkFt2_0),.clk(gclk));
	jdff dff_A_CAtbH0kG3_1(.dout(w_G468_1[1]),.din(w_dff_A_CAtbH0kG3_1),.clk(gclk));
	jdff dff_A_UDKg6Xpi4_1(.dout(w_dff_A_CAtbH0kG3_1),.din(w_dff_A_UDKg6Xpi4_1),.clk(gclk));
	jdff dff_A_7boYskag2_1(.dout(w_dff_A_UDKg6Xpi4_1),.din(w_dff_A_7boYskag2_1),.clk(gclk));
	jdff dff_B_Uu9M7lfg3_1(.din(n1566),.dout(w_dff_B_Uu9M7lfg3_1),.clk(gclk));
	jdff dff_A_5T6fR9mq7_0(.dout(w_G218_1[0]),.din(w_dff_A_5T6fR9mq7_0),.clk(gclk));
	jdff dff_A_V2kTa9Hc7_1(.dout(w_G468_0[1]),.din(w_dff_A_V2kTa9Hc7_1),.clk(gclk));
	jdff dff_A_CBiKKZIS9_1(.dout(w_dff_A_V2kTa9Hc7_1),.din(w_dff_A_CBiKKZIS9_1),.clk(gclk));
	jdff dff_A_m63lOlLZ0_2(.dout(w_G468_0[2]),.din(w_dff_A_m63lOlLZ0_2),.clk(gclk));
	jdff dff_A_RCuN0zd90_2(.dout(w_dff_A_m63lOlLZ0_2),.din(w_dff_A_RCuN0zd90_2),.clk(gclk));
	jdff dff_A_ceAiW7Ji5_2(.dout(w_dff_A_RCuN0zd90_2),.din(w_dff_A_ceAiW7Ji5_2),.clk(gclk));
	jdff dff_A_iNfwLSLT6_2(.dout(w_dff_A_ceAiW7Ji5_2),.din(w_dff_A_iNfwLSLT6_2),.clk(gclk));
	jdff dff_A_9Ucm2QPV0_0(.dout(w_G218_2[0]),.din(w_dff_A_9Ucm2QPV0_0),.clk(gclk));
	jdff dff_B_ylgvBcdh8_1(.din(n1556),.dout(w_dff_B_ylgvBcdh8_1),.clk(gclk));
	jdff dff_B_StMgBiOW8_1(.din(w_dff_B_ylgvBcdh8_1),.dout(w_dff_B_StMgBiOW8_1),.clk(gclk));
	jdff dff_A_Jv4JdZ5u5_0(.dout(w_G226_2[0]),.din(w_dff_A_Jv4JdZ5u5_0),.clk(gclk));
	jdff dff_A_bObf0x0p0_2(.dout(w_n496_0[2]),.din(w_dff_A_bObf0x0p0_2),.clk(gclk));
	jdff dff_A_QUtchzXp5_2(.dout(w_dff_A_bObf0x0p0_2),.din(w_dff_A_QUtchzXp5_2),.clk(gclk));
	jdff dff_A_cKTpejlu2_2(.dout(w_dff_A_QUtchzXp5_2),.din(w_dff_A_cKTpejlu2_2),.clk(gclk));
	jdff dff_B_sAWPCcwN2_3(.din(n496),.dout(w_dff_B_sAWPCcwN2_3),.clk(gclk));
	jdff dff_A_LiPYbX3r1_0(.dout(w_G422_1[0]),.din(w_dff_A_LiPYbX3r1_0),.clk(gclk));
	jdff dff_A_h8wzHYHy1_0(.dout(w_dff_A_LiPYbX3r1_0),.din(w_dff_A_h8wzHYHy1_0),.clk(gclk));
	jdff dff_A_Y8ywuaNP0_0(.dout(w_dff_A_h8wzHYHy1_0),.din(w_dff_A_Y8ywuaNP0_0),.clk(gclk));
	jdff dff_A_n7tyjkY01_1(.dout(w_G422_0[1]),.din(w_dff_A_n7tyjkY01_1),.clk(gclk));
	jdff dff_A_t0O7mI4e6_1(.dout(w_dff_A_n7tyjkY01_1),.din(w_dff_A_t0O7mI4e6_1),.clk(gclk));
	jdff dff_A_V3QMQZlU8_1(.dout(w_dff_A_t0O7mI4e6_1),.din(w_dff_A_V3QMQZlU8_1),.clk(gclk));
	jdff dff_A_Aw4CuAdT5_2(.dout(w_G422_0[2]),.din(w_dff_A_Aw4CuAdT5_2),.clk(gclk));
	jdff dff_A_fy8QgxEM9_2(.dout(w_dff_A_Aw4CuAdT5_2),.din(w_dff_A_fy8QgxEM9_2),.clk(gclk));
	jdff dff_A_TqHrAkxw9_2(.dout(w_dff_A_fy8QgxEM9_2),.din(w_dff_A_TqHrAkxw9_2),.clk(gclk));
	jdff dff_A_6SJLGo5A5_2(.dout(w_dff_A_TqHrAkxw9_2),.din(w_dff_A_6SJLGo5A5_2),.clk(gclk));
	jdff dff_A_L2otT6Jw9_2(.dout(w_G226_0[2]),.din(w_dff_A_L2otT6Jw9_2),.clk(gclk));
	jdff dff_B_PlhzTukc7_1(.din(n541),.dout(w_dff_B_PlhzTukc7_1),.clk(gclk));
	jdff dff_B_z34FMFxU3_1(.din(w_dff_B_PlhzTukc7_1),.dout(w_dff_B_z34FMFxU3_1),.clk(gclk));
	jdff dff_B_urOdmBcw5_1(.din(n542),.dout(w_dff_B_urOdmBcw5_1),.clk(gclk));
	jdff dff_A_zDVZzJHB6_0(.dout(w_G446_1[0]),.din(w_dff_A_zDVZzJHB6_0),.clk(gclk));
	jdff dff_A_h0CDLY6r9_0(.dout(w_dff_A_zDVZzJHB6_0),.din(w_dff_A_h0CDLY6r9_0),.clk(gclk));
	jdff dff_A_VNw9zwzH9_0(.dout(w_dff_A_h0CDLY6r9_0),.din(w_dff_A_VNw9zwzH9_0),.clk(gclk));
	jdff dff_A_8WUE9jgd9_1(.dout(w_G446_1[1]),.din(w_dff_A_8WUE9jgd9_1),.clk(gclk));
	jdff dff_A_xzteHJPG2_1(.dout(w_dff_A_8WUE9jgd9_1),.din(w_dff_A_xzteHJPG2_1),.clk(gclk));
	jdff dff_A_Bt3PYd0s2_1(.dout(w_dff_A_xzteHJPG2_1),.din(w_dff_A_Bt3PYd0s2_1),.clk(gclk));
	jdff dff_A_lHGUgZ8b5_1(.dout(w_G446_0[1]),.din(w_dff_A_lHGUgZ8b5_1),.clk(gclk));
	jdff dff_A_soqt4kU63_1(.dout(w_dff_A_lHGUgZ8b5_1),.din(w_dff_A_soqt4kU63_1),.clk(gclk));
	jdff dff_A_J674rONt9_1(.dout(w_dff_A_soqt4kU63_1),.din(w_dff_A_J674rONt9_1),.clk(gclk));
	jdff dff_A_5IPRpY9Y5_2(.dout(w_G446_0[2]),.din(w_dff_A_5IPRpY9Y5_2),.clk(gclk));
	jdff dff_A_hO3uPZj88_2(.dout(w_dff_A_5IPRpY9Y5_2),.din(w_dff_A_hO3uPZj88_2),.clk(gclk));
	jdff dff_A_f02csFex8_2(.dout(w_dff_A_hO3uPZj88_2),.din(w_dff_A_f02csFex8_2),.clk(gclk));
	jdff dff_A_qKmwbaOo2_0(.dout(w_G206_1[0]),.din(w_dff_A_qKmwbaOo2_0),.clk(gclk));
	jdff dff_B_kI5zuntE0_1(.din(n1525),.dout(w_dff_B_kI5zuntE0_1),.clk(gclk));
	jdff dff_B_nIieNhIp4_1(.din(n1534),.dout(w_dff_B_nIieNhIp4_1),.clk(gclk));
	jdff dff_B_sAsxMiBZ5_1(.din(n1544),.dout(w_dff_B_sAsxMiBZ5_1),.clk(gclk));
	jdff dff_B_LRLQwiRy6_1(.din(w_dff_B_sAsxMiBZ5_1),.dout(w_dff_B_LRLQwiRy6_1),.clk(gclk));
	jdff dff_A_6W7MCHnj4_0(.dout(w_G234_2[0]),.din(w_dff_A_6W7MCHnj4_0),.clk(gclk));
	jdff dff_A_Dsae1irt7_1(.dout(w_n462_0[1]),.din(w_dff_A_Dsae1irt7_1),.clk(gclk));
	jdff dff_A_d1Rk1TxE4_1(.dout(w_dff_A_Dsae1irt7_1),.din(w_dff_A_d1Rk1TxE4_1),.clk(gclk));
	jdff dff_A_JEmkZMiG7_1(.dout(w_dff_A_d1Rk1TxE4_1),.din(w_dff_A_JEmkZMiG7_1),.clk(gclk));
	jdff dff_B_MdGS8fv19_3(.din(n462),.dout(w_dff_B_MdGS8fv19_3),.clk(gclk));
	jdff dff_A_M6dwSquL8_0(.dout(w_G435_1[0]),.din(w_dff_A_M6dwSquL8_0),.clk(gclk));
	jdff dff_A_6mWxIoI89_0(.dout(w_dff_A_M6dwSquL8_0),.din(w_dff_A_6mWxIoI89_0),.clk(gclk));
	jdff dff_A_eW6SjnNt7_0(.dout(w_dff_A_6mWxIoI89_0),.din(w_dff_A_eW6SjnNt7_0),.clk(gclk));
	jdff dff_A_hBJWfctI0_0(.dout(w_dff_A_eW6SjnNt7_0),.din(w_dff_A_hBJWfctI0_0),.clk(gclk));
	jdff dff_A_oei47RLu4_1(.dout(w_G435_1[1]),.din(w_dff_A_oei47RLu4_1),.clk(gclk));
	jdff dff_A_DcZGlTqU3_1(.dout(w_dff_A_oei47RLu4_1),.din(w_dff_A_DcZGlTqU3_1),.clk(gclk));
	jdff dff_A_Lb2WQcSu6_1(.dout(w_dff_A_DcZGlTqU3_1),.din(w_dff_A_Lb2WQcSu6_1),.clk(gclk));
	jdff dff_A_yApM7iip3_1(.dout(w_G435_0[1]),.din(w_dff_A_yApM7iip3_1),.clk(gclk));
	jdff dff_A_chyFBETF2_1(.dout(w_dff_A_yApM7iip3_1),.din(w_dff_A_chyFBETF2_1),.clk(gclk));
	jdff dff_A_Ien8KOZI6_1(.dout(w_dff_A_chyFBETF2_1),.din(w_dff_A_Ien8KOZI6_1),.clk(gclk));
	jdff dff_A_neKV7vsi6_2(.dout(w_G435_0[2]),.din(w_dff_A_neKV7vsi6_2),.clk(gclk));
	jdff dff_A_zOuC35UD9_2(.dout(w_dff_A_neKV7vsi6_2),.din(w_dff_A_zOuC35UD9_2),.clk(gclk));
	jdff dff_A_nAihT9iC1_2(.dout(w_dff_A_zOuC35UD9_2),.din(w_dff_A_nAihT9iC1_2),.clk(gclk));
	jdff dff_A_fMLuO8Bl6_2(.dout(w_dff_A_nAihT9iC1_2),.din(w_dff_A_fMLuO8Bl6_2),.clk(gclk));
	jdff dff_A_2Fs1iHVf5_2(.dout(w_G234_0[2]),.din(w_dff_A_2Fs1iHVf5_2),.clk(gclk));
	jdff dff_B_9PHn1ibD1_1(.din(n1535),.dout(w_dff_B_9PHn1ibD1_1),.clk(gclk));
	jdff dff_B_4dGYIH7l0_1(.din(w_dff_B_9PHn1ibD1_1),.dout(w_dff_B_4dGYIH7l0_1),.clk(gclk));
	jdff dff_A_m2EfBMWh9_0(.dout(w_G257_2[0]),.din(w_dff_A_m2EfBMWh9_0),.clk(gclk));
	jdff dff_A_lyM7So0B9_1(.dout(w_n520_0[1]),.din(w_dff_A_lyM7So0B9_1),.clk(gclk));
	jdff dff_A_1JaE5bQI8_1(.dout(w_dff_A_lyM7So0B9_1),.din(w_dff_A_1JaE5bQI8_1),.clk(gclk));
	jdff dff_B_rPXNYChq5_3(.din(n520),.dout(w_dff_B_rPXNYChq5_3),.clk(gclk));
	jdff dff_A_AkSqn7jB1_0(.dout(w_G389_1[0]),.din(w_dff_A_AkSqn7jB1_0),.clk(gclk));
	jdff dff_A_7evdrxR06_0(.dout(w_dff_A_AkSqn7jB1_0),.din(w_dff_A_7evdrxR06_0),.clk(gclk));
	jdff dff_A_wHxj0fRF9_0(.dout(w_dff_A_7evdrxR06_0),.din(w_dff_A_wHxj0fRF9_0),.clk(gclk));
	jdff dff_A_Lc2dYLdb9_0(.dout(w_dff_A_wHxj0fRF9_0),.din(w_dff_A_Lc2dYLdb9_0),.clk(gclk));
	jdff dff_A_R3XFGVbj1_1(.dout(w_G389_1[1]),.din(w_dff_A_R3XFGVbj1_1),.clk(gclk));
	jdff dff_A_sbI6OpWy7_1(.dout(w_dff_A_R3XFGVbj1_1),.din(w_dff_A_sbI6OpWy7_1),.clk(gclk));
	jdff dff_A_21gc5b9b6_1(.dout(w_dff_A_sbI6OpWy7_1),.din(w_dff_A_21gc5b9b6_1),.clk(gclk));
	jdff dff_A_ESqOpbAI9_1(.dout(w_G389_0[1]),.din(w_dff_A_ESqOpbAI9_1),.clk(gclk));
	jdff dff_A_WiOLTzjr3_1(.dout(w_dff_A_ESqOpbAI9_1),.din(w_dff_A_WiOLTzjr3_1),.clk(gclk));
	jdff dff_A_GQKc1rbV2_1(.dout(w_dff_A_WiOLTzjr3_1),.din(w_dff_A_GQKc1rbV2_1),.clk(gclk));
	jdff dff_A_IgQAQ7Lt9_2(.dout(w_G389_0[2]),.din(w_dff_A_IgQAQ7Lt9_2),.clk(gclk));
	jdff dff_A_KfzvHsFa9_2(.dout(w_dff_A_IgQAQ7Lt9_2),.din(w_dff_A_KfzvHsFa9_2),.clk(gclk));
	jdff dff_A_c3nhZ7hv3_2(.dout(w_dff_A_KfzvHsFa9_2),.din(w_dff_A_c3nhZ7hv3_2),.clk(gclk));
	jdff dff_A_Mr0oGODM8_2(.dout(w_dff_A_c3nhZ7hv3_2),.din(w_dff_A_Mr0oGODM8_2),.clk(gclk));
	jdff dff_A_I6WA4MZP3_2(.dout(w_G257_0[2]),.din(w_dff_A_I6WA4MZP3_2),.clk(gclk));
	jdff dff_B_XtCAGJFa0_1(.din(n1530),.dout(w_dff_B_XtCAGJFa0_1),.clk(gclk));
	jdff dff_A_ZS8Xkajg5_1(.dout(w_n485_0[1]),.din(w_dff_A_ZS8Xkajg5_1),.clk(gclk));
	jdff dff_A_iRVMvfNT1_1(.dout(w_dff_A_ZS8Xkajg5_1),.din(w_dff_A_iRVMvfNT1_1),.clk(gclk));
	jdff dff_A_DxScrfm78_2(.dout(w_n485_0[2]),.din(w_dff_A_DxScrfm78_2),.clk(gclk));
	jdff dff_B_Kg99jZtm0_3(.din(n485),.dout(w_dff_B_Kg99jZtm0_3),.clk(gclk));
	jdff dff_A_WG9HIbrZ6_0(.dout(w_G400_1[0]),.din(w_dff_A_WG9HIbrZ6_0),.clk(gclk));
	jdff dff_A_6smh6VMm0_0(.dout(w_dff_A_WG9HIbrZ6_0),.din(w_dff_A_6smh6VMm0_0),.clk(gclk));
	jdff dff_A_tiMkaR712_0(.dout(w_dff_A_6smh6VMm0_0),.din(w_dff_A_tiMkaR712_0),.clk(gclk));
	jdff dff_A_PqVa93ns6_0(.dout(w_dff_A_tiMkaR712_0),.din(w_dff_A_PqVa93ns6_0),.clk(gclk));
	jdff dff_A_TlxaThbe6_1(.dout(w_G400_1[1]),.din(w_dff_A_TlxaThbe6_1),.clk(gclk));
	jdff dff_A_Hh6tT1RF8_1(.dout(w_dff_A_TlxaThbe6_1),.din(w_dff_A_Hh6tT1RF8_1),.clk(gclk));
	jdff dff_A_sAN6ISD43_1(.dout(w_dff_A_Hh6tT1RF8_1),.din(w_dff_A_sAN6ISD43_1),.clk(gclk));
	jdff dff_B_qOYXn8xu5_1(.din(n1526),.dout(w_dff_B_qOYXn8xu5_1),.clk(gclk));
	jdff dff_A_T83XRwcv4_0(.dout(w_G251_5[0]),.din(w_dff_A_T83XRwcv4_0),.clk(gclk));
	jdff dff_A_EgLqHu1D1_0(.dout(w_G251_1[0]),.din(w_dff_A_EgLqHu1D1_0),.clk(gclk));
	jdff dff_A_fN7vApHP4_2(.dout(w_G251_1[2]),.din(w_dff_A_fN7vApHP4_2),.clk(gclk));
	jdff dff_A_JpespLa43_1(.dout(w_G400_0[1]),.din(w_dff_A_JpespLa43_1),.clk(gclk));
	jdff dff_A_8feY9c7F4_1(.dout(w_dff_A_JpespLa43_1),.din(w_dff_A_8feY9c7F4_1),.clk(gclk));
	jdff dff_A_8Lh2rrkD9_2(.dout(w_G400_0[2]),.din(w_dff_A_8Lh2rrkD9_2),.clk(gclk));
	jdff dff_A_1vRxJY3l1_2(.dout(w_dff_A_8Lh2rrkD9_2),.din(w_dff_A_1vRxJY3l1_2),.clk(gclk));
	jdff dff_A_43WpCtLJ3_2(.dout(w_dff_A_1vRxJY3l1_2),.din(w_dff_A_43WpCtLJ3_2),.clk(gclk));
	jdff dff_A_TNgrttFd5_2(.dout(w_dff_A_43WpCtLJ3_2),.din(w_dff_A_TNgrttFd5_2),.clk(gclk));
	jdff dff_A_HdWVF1nR3_1(.dout(w_G265_1[1]),.din(w_dff_A_HdWVF1nR3_1),.clk(gclk));
	jdff dff_A_GWO37M1N8_2(.dout(w_G265_0[2]),.din(w_dff_A_GWO37M1N8_2),.clk(gclk));
	jdff dff_B_6xNAJWZH8_1(.din(n1516),.dout(w_dff_B_6xNAJWZH8_1),.clk(gclk));
	jdff dff_B_w3oQLA3K1_1(.din(w_dff_B_6xNAJWZH8_1),.dout(w_dff_B_w3oQLA3K1_1),.clk(gclk));
	jdff dff_A_4sti3Suj9_0(.dout(w_G281_2[0]),.din(w_dff_A_4sti3Suj9_0),.clk(gclk));
	jdff dff_A_eXonkdlb7_1(.dout(w_n532_0[1]),.din(w_dff_A_eXonkdlb7_1),.clk(gclk));
	jdff dff_A_7c7731Fg5_1(.dout(w_dff_A_eXonkdlb7_1),.din(w_dff_A_7c7731Fg5_1),.clk(gclk));
	jdff dff_A_pdvO5LkK8_2(.dout(w_n532_0[2]),.din(w_dff_A_pdvO5LkK8_2),.clk(gclk));
	jdff dff_A_toLIV1WJ6_2(.dout(w_dff_A_pdvO5LkK8_2),.din(w_dff_A_toLIV1WJ6_2),.clk(gclk));
	jdff dff_B_AdYaPkP42_3(.din(n532),.dout(w_dff_B_AdYaPkP42_3),.clk(gclk));
	jdff dff_A_VSZtUZ2U3_0(.dout(w_G374_1[0]),.din(w_dff_A_VSZtUZ2U3_0),.clk(gclk));
	jdff dff_A_8iuV7Q6Y6_0(.dout(w_dff_A_VSZtUZ2U3_0),.din(w_dff_A_8iuV7Q6Y6_0),.clk(gclk));
	jdff dff_A_aRqKwDbl9_0(.dout(w_dff_A_8iuV7Q6Y6_0),.din(w_dff_A_aRqKwDbl9_0),.clk(gclk));
	jdff dff_A_n93wh5bo2_0(.dout(w_dff_A_aRqKwDbl9_0),.din(w_dff_A_n93wh5bo2_0),.clk(gclk));
	jdff dff_A_Qh7Wzjfr2_1(.dout(w_G374_1[1]),.din(w_dff_A_Qh7Wzjfr2_1),.clk(gclk));
	jdff dff_A_Ix1uHo1p1_1(.dout(w_dff_A_Qh7Wzjfr2_1),.din(w_dff_A_Ix1uHo1p1_1),.clk(gclk));
	jdff dff_A_Gn4kNrmx8_1(.dout(w_dff_A_Ix1uHo1p1_1),.din(w_dff_A_Gn4kNrmx8_1),.clk(gclk));
	jdff dff_A_BO4uaQtK5_1(.dout(w_G374_0[1]),.din(w_dff_A_BO4uaQtK5_1),.clk(gclk));
	jdff dff_A_zeXCtxqQ1_1(.dout(w_dff_A_BO4uaQtK5_1),.din(w_dff_A_zeXCtxqQ1_1),.clk(gclk));
	jdff dff_A_Dw0DhlT63_1(.dout(w_dff_A_zeXCtxqQ1_1),.din(w_dff_A_Dw0DhlT63_1),.clk(gclk));
	jdff dff_A_9wZqrTU88_2(.dout(w_G374_0[2]),.din(w_dff_A_9wZqrTU88_2),.clk(gclk));
	jdff dff_A_TK5xeshE4_2(.dout(w_dff_A_9wZqrTU88_2),.din(w_dff_A_TK5xeshE4_2),.clk(gclk));
	jdff dff_A_bvrIgDs56_2(.dout(w_dff_A_TK5xeshE4_2),.din(w_dff_A_bvrIgDs56_2),.clk(gclk));
	jdff dff_A_k06UHQ5A1_2(.dout(w_dff_A_bvrIgDs56_2),.din(w_dff_A_k06UHQ5A1_2),.clk(gclk));
	jdff dff_A_iLESAI844_2(.dout(w_G281_0[2]),.din(w_dff_A_iLESAI844_2),.clk(gclk));
	jdff dff_A_ZPs6zkcb8_0(.dout(w_G242_1[0]),.din(w_dff_A_ZPs6zkcb8_0),.clk(gclk));
	jdff dff_A_l8cnWHa37_1(.dout(w_G242_0[1]),.din(w_dff_A_l8cnWHa37_1),.clk(gclk));
	jdff dff_A_USw4L3wP5_2(.dout(w_G242_0[2]),.din(w_dff_A_USw4L3wP5_2),.clk(gclk));
	jdff dff_B_Ql6raKPb3_1(.din(n1507),.dout(w_dff_B_Ql6raKPb3_1),.clk(gclk));
	jdff dff_B_6uWvkJM58_1(.din(w_dff_B_Ql6raKPb3_1),.dout(w_dff_B_6uWvkJM58_1),.clk(gclk));
	jdff dff_A_q5DKJWwU8_0(.dout(w_G273_2[0]),.din(w_dff_A_q5DKJWwU8_0),.clk(gclk));
	jdff dff_A_kUArhjPR1_1(.dout(w_G251_0[1]),.din(w_dff_A_kUArhjPR1_1),.clk(gclk));
	jdff dff_A_1XgLJ2H39_2(.dout(w_G251_0[2]),.din(w_dff_A_1XgLJ2H39_2),.clk(gclk));
	jdff dff_A_zHIQzKii4_1(.dout(w_n473_0[1]),.din(w_dff_A_zHIQzKii4_1),.clk(gclk));
	jdff dff_A_AAJrBaP18_1(.dout(w_dff_A_zHIQzKii4_1),.din(w_dff_A_AAJrBaP18_1),.clk(gclk));
	jdff dff_A_Q9KvcXOf2_2(.dout(w_n473_0[2]),.din(w_dff_A_Q9KvcXOf2_2),.clk(gclk));
	jdff dff_A_4IPrpr5s0_2(.dout(w_dff_A_Q9KvcXOf2_2),.din(w_dff_A_4IPrpr5s0_2),.clk(gclk));
	jdff dff_B_7icCghZd5_3(.din(n473),.dout(w_dff_B_7icCghZd5_3),.clk(gclk));
	jdff dff_A_VCgnQjQ24_0(.dout(w_G411_2[0]),.din(w_dff_A_VCgnQjQ24_0),.clk(gclk));
	jdff dff_A_1bSRuFLQ6_0(.dout(w_dff_A_VCgnQjQ24_0),.din(w_dff_A_1bSRuFLQ6_0),.clk(gclk));
	jdff dff_A_TnqCR82Q3_0(.dout(w_dff_A_1bSRuFLQ6_0),.din(w_dff_A_TnqCR82Q3_0),.clk(gclk));
	jdff dff_A_brC3Vu6C4_0(.dout(w_G411_0[0]),.din(w_dff_A_brC3Vu6C4_0),.clk(gclk));
	jdff dff_A_8ZqrcTiy8_0(.dout(w_dff_A_brC3Vu6C4_0),.din(w_dff_A_8ZqrcTiy8_0),.clk(gclk));
	jdff dff_A_ltWXsAXG3_0(.dout(w_dff_A_8ZqrcTiy8_0),.din(w_dff_A_ltWXsAXG3_0),.clk(gclk));
	jdff dff_A_ug8P8f0F0_0(.dout(w_dff_A_ltWXsAXG3_0),.din(w_dff_A_ug8P8f0F0_0),.clk(gclk));
	jdff dff_A_BJ7UxRqH7_2(.dout(w_G411_0[2]),.din(w_dff_A_BJ7UxRqH7_2),.clk(gclk));
	jdff dff_A_UccuB1zX9_2(.dout(w_dff_A_BJ7UxRqH7_2),.din(w_dff_A_UccuB1zX9_2),.clk(gclk));
	jdff dff_A_ai55PT6o1_2(.dout(w_dff_A_UccuB1zX9_2),.din(w_dff_A_ai55PT6o1_2),.clk(gclk));
	jdff dff_A_2Rh94nuT9_1(.dout(w_G273_1[1]),.din(w_dff_A_2Rh94nuT9_1),.clk(gclk));
	jdff dff_A_wwkj1LBC5_2(.dout(w_G273_0[2]),.din(w_dff_A_wwkj1LBC5_2),.clk(gclk));
	jdff dff_A_clY56xZi9_2(.dout(w_G248_3[2]),.din(w_dff_A_clY56xZi9_2),.clk(gclk));
	jdff dff_A_4BjCnYsa4_1(.dout(w_n749_4[1]),.din(w_dff_A_4BjCnYsa4_1),.clk(gclk));
	jdff dff_A_njzoyN1m1_1(.dout(w_dff_A_4BjCnYsa4_1),.din(w_dff_A_njzoyN1m1_1),.clk(gclk));
	jdff dff_A_TXctprQw6_1(.dout(w_dff_A_njzoyN1m1_1),.din(w_dff_A_TXctprQw6_1),.clk(gclk));
	jdff dff_A_TZQPaEs70_1(.dout(w_dff_A_TXctprQw6_1),.din(w_dff_A_TZQPaEs70_1),.clk(gclk));
	jdff dff_A_wzyPVgss4_1(.dout(w_dff_A_TZQPaEs70_1),.din(w_dff_A_wzyPVgss4_1),.clk(gclk));
	jdff dff_A_Q2uzrKly3_1(.dout(w_dff_A_wzyPVgss4_1),.din(w_dff_A_Q2uzrKly3_1),.clk(gclk));
	jdff dff_A_jtu5VeW96_1(.dout(w_dff_A_Q2uzrKly3_1),.din(w_dff_A_jtu5VeW96_1),.clk(gclk));
	jdff dff_A_c7aqkdPO9_1(.dout(w_dff_A_jtu5VeW96_1),.din(w_dff_A_c7aqkdPO9_1),.clk(gclk));
	jdff dff_A_gjXtJhIe4_1(.dout(w_dff_A_c7aqkdPO9_1),.din(w_dff_A_gjXtJhIe4_1),.clk(gclk));
	jdff dff_A_uNcQqXEt9_1(.dout(w_dff_A_gjXtJhIe4_1),.din(w_dff_A_uNcQqXEt9_1),.clk(gclk));
	jdff dff_A_lzXJE4H84_1(.dout(w_dff_A_uNcQqXEt9_1),.din(w_dff_A_lzXJE4H84_1),.clk(gclk));
	jdff dff_A_OYGfwP1Z3_1(.dout(w_dff_A_lzXJE4H84_1),.din(w_dff_A_OYGfwP1Z3_1),.clk(gclk));
	jdff dff_A_Vng23Yzf7_1(.dout(w_dff_A_OYGfwP1Z3_1),.din(w_dff_A_Vng23Yzf7_1),.clk(gclk));
	jdff dff_A_KmbM6YnM1_1(.dout(w_dff_A_Vng23Yzf7_1),.din(w_dff_A_KmbM6YnM1_1),.clk(gclk));
	jdff dff_A_7jCuN2SO5_1(.dout(w_dff_A_KmbM6YnM1_1),.din(w_dff_A_7jCuN2SO5_1),.clk(gclk));
	jdff dff_A_B0JxwjqZ0_1(.dout(w_dff_A_7jCuN2SO5_1),.din(w_dff_A_B0JxwjqZ0_1),.clk(gclk));
	jdff dff_A_BR90ggWF7_1(.dout(w_dff_A_B0JxwjqZ0_1),.din(w_dff_A_BR90ggWF7_1),.clk(gclk));
	jdff dff_A_TwZAxml05_2(.dout(w_n749_4[2]),.din(w_dff_A_TwZAxml05_2),.clk(gclk));
	jdff dff_A_CAfVWKOV4_2(.dout(w_dff_A_TwZAxml05_2),.din(w_dff_A_CAfVWKOV4_2),.clk(gclk));
	jdff dff_A_IO2PFiQm1_2(.dout(w_dff_A_CAfVWKOV4_2),.din(w_dff_A_IO2PFiQm1_2),.clk(gclk));
	jdff dff_A_d7PL8Z2r4_2(.dout(w_dff_A_IO2PFiQm1_2),.din(w_dff_A_d7PL8Z2r4_2),.clk(gclk));
	jdff dff_A_0HITXgMS0_2(.dout(w_dff_A_d7PL8Z2r4_2),.din(w_dff_A_0HITXgMS0_2),.clk(gclk));
	jdff dff_A_Roh18i988_2(.dout(w_dff_A_0HITXgMS0_2),.din(w_dff_A_Roh18i988_2),.clk(gclk));
	jdff dff_A_jfhLXF6C8_2(.dout(w_dff_A_Roh18i988_2),.din(w_dff_A_jfhLXF6C8_2),.clk(gclk));
	jdff dff_A_l3hale7f1_2(.dout(w_dff_A_jfhLXF6C8_2),.din(w_dff_A_l3hale7f1_2),.clk(gclk));
	jdff dff_A_3vhr76GN0_1(.dout(w_n749_1[1]),.din(w_dff_A_3vhr76GN0_1),.clk(gclk));
	jdff dff_A_WtPchuSZ3_1(.dout(w_dff_A_3vhr76GN0_1),.din(w_dff_A_WtPchuSZ3_1),.clk(gclk));
	jdff dff_A_AP2UQUWH2_1(.dout(w_dff_A_WtPchuSZ3_1),.din(w_dff_A_AP2UQUWH2_1),.clk(gclk));
	jdff dff_A_XjrQOuP52_1(.dout(w_dff_A_AP2UQUWH2_1),.din(w_dff_A_XjrQOuP52_1),.clk(gclk));
	jdff dff_A_R3CgJ9rL2_2(.dout(w_n749_1[2]),.din(w_dff_A_R3CgJ9rL2_2),.clk(gclk));
	jdff dff_A_s3CCG6I42_2(.dout(w_dff_A_R3CgJ9rL2_2),.din(w_dff_A_s3CCG6I42_2),.clk(gclk));
	jdff dff_A_j0w5OR4N7_2(.dout(w_dff_A_s3CCG6I42_2),.din(w_dff_A_j0w5OR4N7_2),.clk(gclk));
	jdff dff_A_Dq9oZTdE6_2(.dout(w_dff_A_j0w5OR4N7_2),.din(w_dff_A_Dq9oZTdE6_2),.clk(gclk));
	jdff dff_A_z1Hfe0YB5_1(.dout(w_n749_0[1]),.din(w_dff_A_z1Hfe0YB5_1),.clk(gclk));
	jdff dff_A_wjIhlaw92_1(.dout(w_dff_A_z1Hfe0YB5_1),.din(w_dff_A_wjIhlaw92_1),.clk(gclk));
	jdff dff_A_HcshvQVC3_2(.dout(w_n749_0[2]),.din(w_dff_A_HcshvQVC3_2),.clk(gclk));
	jdff dff_A_g0hCcZSf8_2(.dout(w_dff_A_HcshvQVC3_2),.din(w_dff_A_g0hCcZSf8_2),.clk(gclk));
	jdff dff_A_UxkExz4G1_2(.dout(w_dff_A_g0hCcZSf8_2),.din(w_dff_A_UxkExz4G1_2),.clk(gclk));
	jdff dff_A_IOgCYga15_0(.dout(w_G4091_6[0]),.din(w_dff_A_IOgCYga15_0),.clk(gclk));
	jdff dff_A_86Kd2LNp4_0(.dout(w_dff_A_IOgCYga15_0),.din(w_dff_A_86Kd2LNp4_0),.clk(gclk));
	jdff dff_A_GN6xquat4_0(.dout(w_dff_A_86Kd2LNp4_0),.din(w_dff_A_GN6xquat4_0),.clk(gclk));
	jdff dff_A_14eD1Mxq5_0(.dout(w_dff_A_GN6xquat4_0),.din(w_dff_A_14eD1Mxq5_0),.clk(gclk));
	jdff dff_A_7ltQG4E96_0(.dout(w_dff_A_14eD1Mxq5_0),.din(w_dff_A_7ltQG4E96_0),.clk(gclk));
	jdff dff_A_gLWajmgg3_0(.dout(w_G4091_1[0]),.din(w_dff_A_gLWajmgg3_0),.clk(gclk));
	jdff dff_A_n6tz4ecN4_0(.dout(w_dff_A_gLWajmgg3_0),.din(w_dff_A_n6tz4ecN4_0),.clk(gclk));
	jdff dff_A_sHtRfTck5_0(.dout(w_dff_A_n6tz4ecN4_0),.din(w_dff_A_sHtRfTck5_0),.clk(gclk));
	jdff dff_A_wS8O3pQt5_0(.dout(w_dff_A_sHtRfTck5_0),.din(w_dff_A_wS8O3pQt5_0),.clk(gclk));
	jdff dff_A_K1oLFTwL1_0(.dout(w_dff_A_wS8O3pQt5_0),.din(w_dff_A_K1oLFTwL1_0),.clk(gclk));
	jdff dff_A_lQ52r2gm2_0(.dout(w_dff_A_K1oLFTwL1_0),.din(w_dff_A_lQ52r2gm2_0),.clk(gclk));
	jdff dff_A_8eESOUSb4_0(.dout(w_dff_A_lQ52r2gm2_0),.din(w_dff_A_8eESOUSb4_0),.clk(gclk));
	jdff dff_A_hln36Jja8_0(.dout(w_dff_A_8eESOUSb4_0),.din(w_dff_A_hln36Jja8_0),.clk(gclk));
	jdff dff_A_yr91NgLu6_1(.dout(w_G4091_1[1]),.din(w_dff_A_yr91NgLu6_1),.clk(gclk));
	jdff dff_A_mR1OWuD16_1(.dout(w_dff_A_yr91NgLu6_1),.din(w_dff_A_mR1OWuD16_1),.clk(gclk));
	jdff dff_A_4J4jjHV49_1(.dout(w_dff_A_mR1OWuD16_1),.din(w_dff_A_4J4jjHV49_1),.clk(gclk));
	jdff dff_A_PDU8dyMk8_1(.dout(w_dff_A_4J4jjHV49_1),.din(w_dff_A_PDU8dyMk8_1),.clk(gclk));
	jdff dff_A_7GFOFje68_1(.dout(w_dff_A_PDU8dyMk8_1),.din(w_dff_A_7GFOFje68_1),.clk(gclk));
	jdff dff_A_OVOQANxh2_1(.dout(w_dff_A_7GFOFje68_1),.din(w_dff_A_OVOQANxh2_1),.clk(gclk));
	jdff dff_A_0NTHthet9_1(.dout(w_dff_A_OVOQANxh2_1),.din(w_dff_A_0NTHthet9_1),.clk(gclk));
	jdff dff_A_zonUQtxB9_1(.dout(w_G4091_0[1]),.din(w_dff_A_zonUQtxB9_1),.clk(gclk));
	jdff dff_A_GLtjp44R2_1(.dout(w_dff_A_zonUQtxB9_1),.din(w_dff_A_GLtjp44R2_1),.clk(gclk));
	jdff dff_A_LTlLwcGZ3_1(.dout(w_dff_A_GLtjp44R2_1),.din(w_dff_A_LTlLwcGZ3_1),.clk(gclk));
	jdff dff_A_pVlcDcYX3_1(.dout(w_dff_A_LTlLwcGZ3_1),.din(w_dff_A_pVlcDcYX3_1),.clk(gclk));
	jdff dff_A_0cskcqzx9_1(.dout(w_dff_A_pVlcDcYX3_1),.din(w_dff_A_0cskcqzx9_1),.clk(gclk));
	jdff dff_A_0YbbMCGp7_1(.dout(w_dff_A_0cskcqzx9_1),.din(w_dff_A_0YbbMCGp7_1),.clk(gclk));
	jdff dff_A_VZTMw77M2_1(.dout(w_dff_A_0YbbMCGp7_1),.din(w_dff_A_VZTMw77M2_1),.clk(gclk));
	jdff dff_A_fGYA6cGq5_1(.dout(w_dff_A_VZTMw77M2_1),.din(w_dff_A_fGYA6cGq5_1),.clk(gclk));
	jdff dff_A_rkY8ZJQK5_1(.dout(w_dff_A_fGYA6cGq5_1),.din(w_dff_A_rkY8ZJQK5_1),.clk(gclk));
	jdff dff_A_WSYn5Wlw5_1(.dout(w_dff_A_rkY8ZJQK5_1),.din(w_dff_A_WSYn5Wlw5_1),.clk(gclk));
	jdff dff_A_JKDn27689_1(.dout(w_dff_A_WSYn5Wlw5_1),.din(w_dff_A_JKDn27689_1),.clk(gclk));
	jdff dff_A_yCTbubjL7_1(.dout(w_dff_A_JKDn27689_1),.din(w_dff_A_yCTbubjL7_1),.clk(gclk));
	jdff dff_A_TYG55EF44_1(.dout(w_dff_A_yCTbubjL7_1),.din(w_dff_A_TYG55EF44_1),.clk(gclk));
	jdff dff_A_LyDSgra93_2(.dout(w_G4091_0[2]),.din(w_dff_A_LyDSgra93_2),.clk(gclk));
	jdff dff_A_ngEZdzKZ3_2(.dout(w_dff_A_LyDSgra93_2),.din(w_dff_A_ngEZdzKZ3_2),.clk(gclk));
	jdff dff_A_JhkqXMBe3_2(.dout(w_dff_A_ngEZdzKZ3_2),.din(w_dff_A_JhkqXMBe3_2),.clk(gclk));
	jdff dff_A_ERXfpw1o9_2(.dout(w_dff_A_JhkqXMBe3_2),.din(w_dff_A_ERXfpw1o9_2),.clk(gclk));
	jdff dff_A_GYFs6pbO1_2(.dout(w_dff_A_ERXfpw1o9_2),.din(w_dff_A_GYFs6pbO1_2),.clk(gclk));
	jdff dff_A_LCeujrmB4_2(.dout(w_dff_A_GYFs6pbO1_2),.din(w_dff_A_LCeujrmB4_2),.clk(gclk));
	jdff dff_A_fcMhHoWx4_2(.dout(w_dff_A_LCeujrmB4_2),.din(w_dff_A_fcMhHoWx4_2),.clk(gclk));
	jdff dff_A_4Hx3joJk7_2(.dout(w_dff_A_fcMhHoWx4_2),.din(w_dff_A_4Hx3joJk7_2),.clk(gclk));
	jdff dff_A_8YGmmi2j1_2(.dout(w_G4092_3[2]),.din(w_dff_A_8YGmmi2j1_2),.clk(gclk));
	jdff dff_A_iGCt53WG4_2(.dout(w_dff_A_8YGmmi2j1_2),.din(w_dff_A_iGCt53WG4_2),.clk(gclk));
	jdff dff_A_C3JoLAx09_2(.dout(w_dff_A_iGCt53WG4_2),.din(w_dff_A_C3JoLAx09_2),.clk(gclk));
	jdff dff_A_3XBG0hhS1_2(.dout(w_dff_A_C3JoLAx09_2),.din(w_dff_A_3XBG0hhS1_2),.clk(gclk));
	jdff dff_A_fwdwVIQH1_2(.dout(w_dff_A_3XBG0hhS1_2),.din(w_dff_A_fwdwVIQH1_2),.clk(gclk));
	jdff dff_A_zvli0YFL3_2(.dout(w_dff_A_fwdwVIQH1_2),.din(w_dff_A_zvli0YFL3_2),.clk(gclk));
	jdff dff_A_ZT65vYE69_2(.dout(w_dff_A_zvli0YFL3_2),.din(w_dff_A_ZT65vYE69_2),.clk(gclk));
	jdff dff_A_HTHRu8sE3_2(.dout(w_dff_A_ZT65vYE69_2),.din(w_dff_A_HTHRu8sE3_2),.clk(gclk));
	jdff dff_A_SlmKESRw3_2(.dout(w_dff_A_HTHRu8sE3_2),.din(w_dff_A_SlmKESRw3_2),.clk(gclk));
	jdff dff_A_y64vHxzW0_2(.dout(w_dff_A_SlmKESRw3_2),.din(w_dff_A_y64vHxzW0_2),.clk(gclk));
	jdff dff_A_bIjzEVme5_2(.dout(w_dff_A_y64vHxzW0_2),.din(w_dff_A_bIjzEVme5_2),.clk(gclk));
	jdff dff_A_b2zXDVxs2_2(.dout(w_dff_A_bIjzEVme5_2),.din(w_dff_A_b2zXDVxs2_2),.clk(gclk));
	jdff dff_A_4QIAdU0v9_2(.dout(w_dff_A_b2zXDVxs2_2),.din(w_dff_A_4QIAdU0v9_2),.clk(gclk));
	jdff dff_A_w1dqKSWk9_2(.dout(w_dff_A_4QIAdU0v9_2),.din(w_dff_A_w1dqKSWk9_2),.clk(gclk));
	jdff dff_A_CW0nffzh6_2(.dout(w_dff_A_w1dqKSWk9_2),.din(w_dff_A_CW0nffzh6_2),.clk(gclk));
	jdff dff_A_NqbDsvmf2_2(.dout(w_dff_A_CW0nffzh6_2),.din(w_dff_A_NqbDsvmf2_2),.clk(gclk));
	jdff dff_A_QjbnviA39_2(.dout(w_dff_A_NqbDsvmf2_2),.din(w_dff_A_QjbnviA39_2),.clk(gclk));
	jdff dff_A_LP9E1LB19_2(.dout(w_dff_A_QjbnviA39_2),.din(w_dff_A_LP9E1LB19_2),.clk(gclk));
	jdff dff_A_5YG3Ifyi2_2(.dout(w_dff_A_LP9E1LB19_2),.din(w_dff_A_5YG3Ifyi2_2),.clk(gclk));
	jdff dff_A_MOuVyOFp9_2(.dout(w_dff_A_5YG3Ifyi2_2),.din(w_dff_A_MOuVyOFp9_2),.clk(gclk));
	jdff dff_A_TPiTsZpu7_1(.dout(w_G4092_0[1]),.din(w_dff_A_TPiTsZpu7_1),.clk(gclk));
	jdff dff_A_hwZAhzoJ4_0(.dout(w_n1008_4[0]),.din(w_dff_A_hwZAhzoJ4_0),.clk(gclk));
	jdff dff_A_8hWr8K4g5_0(.dout(w_dff_A_hwZAhzoJ4_0),.din(w_dff_A_8hWr8K4g5_0),.clk(gclk));
	jdff dff_A_IW0G3zbl3_0(.dout(w_dff_A_8hWr8K4g5_0),.din(w_dff_A_IW0G3zbl3_0),.clk(gclk));
	jdff dff_A_SFV9tUrV6_0(.dout(w_dff_A_IW0G3zbl3_0),.din(w_dff_A_SFV9tUrV6_0),.clk(gclk));
	jdff dff_A_V2XmpVEJ7_0(.dout(w_dff_A_SFV9tUrV6_0),.din(w_dff_A_V2XmpVEJ7_0),.clk(gclk));
	jdff dff_A_tYF0k17L9_0(.dout(w_dff_A_V2XmpVEJ7_0),.din(w_dff_A_tYF0k17L9_0),.clk(gclk));
	jdff dff_A_4Kl91n3z9_0(.dout(w_dff_A_tYF0k17L9_0),.din(w_dff_A_4Kl91n3z9_0),.clk(gclk));
	jdff dff_A_D4IbTBJh3_0(.dout(w_dff_A_4Kl91n3z9_0),.din(w_dff_A_D4IbTBJh3_0),.clk(gclk));
	jdff dff_A_idSQuNNg4_0(.dout(w_dff_A_D4IbTBJh3_0),.din(w_dff_A_idSQuNNg4_0),.clk(gclk));
	jdff dff_A_u0Q7WlNR5_0(.dout(w_dff_A_idSQuNNg4_0),.din(w_dff_A_u0Q7WlNR5_0),.clk(gclk));
	jdff dff_A_wh87OkOv4_0(.dout(w_dff_A_u0Q7WlNR5_0),.din(w_dff_A_wh87OkOv4_0),.clk(gclk));
	jdff dff_A_6IdwTX7I1_0(.dout(w_dff_A_wh87OkOv4_0),.din(w_dff_A_6IdwTX7I1_0),.clk(gclk));
	jdff dff_A_0eu9l9GI7_0(.dout(w_dff_A_6IdwTX7I1_0),.din(w_dff_A_0eu9l9GI7_0),.clk(gclk));
	jdff dff_A_Fr2NndvB0_0(.dout(w_dff_A_0eu9l9GI7_0),.din(w_dff_A_Fr2NndvB0_0),.clk(gclk));
	jdff dff_A_9DaxWcVe5_0(.dout(w_dff_A_Fr2NndvB0_0),.din(w_dff_A_9DaxWcVe5_0),.clk(gclk));
	jdff dff_A_sEoFq9KD7_2(.dout(w_n1008_4[2]),.din(w_dff_A_sEoFq9KD7_2),.clk(gclk));
	jdff dff_A_fdHghczS2_2(.dout(w_dff_A_sEoFq9KD7_2),.din(w_dff_A_fdHghczS2_2),.clk(gclk));
	jdff dff_A_qQcbAbSF7_2(.dout(w_dff_A_fdHghczS2_2),.din(w_dff_A_qQcbAbSF7_2),.clk(gclk));
	jdff dff_A_YoyrKpu44_2(.dout(w_dff_A_qQcbAbSF7_2),.din(w_dff_A_YoyrKpu44_2),.clk(gclk));
	jdff dff_A_BKE3x8si3_2(.dout(w_dff_A_YoyrKpu44_2),.din(w_dff_A_BKE3x8si3_2),.clk(gclk));
	jdff dff_A_I1FDdZFv7_2(.dout(w_dff_A_BKE3x8si3_2),.din(w_dff_A_I1FDdZFv7_2),.clk(gclk));
	jdff dff_A_Ck1vgoxk8_2(.dout(w_dff_A_I1FDdZFv7_2),.din(w_dff_A_Ck1vgoxk8_2),.clk(gclk));
	jdff dff_A_DBsxoXEE2_2(.dout(w_dff_A_Ck1vgoxk8_2),.din(w_dff_A_DBsxoXEE2_2),.clk(gclk));
	jdff dff_A_vtwLbDZy9_2(.dout(w_dff_A_DBsxoXEE2_2),.din(w_dff_A_vtwLbDZy9_2),.clk(gclk));
	jdff dff_A_wdof90BC0_2(.dout(w_dff_A_vtwLbDZy9_2),.din(w_dff_A_wdof90BC0_2),.clk(gclk));
	jdff dff_A_4EUYFJ4L3_1(.dout(w_n1008_1[1]),.din(w_dff_A_4EUYFJ4L3_1),.clk(gclk));
	jdff dff_A_ouFZAQwf3_1(.dout(w_dff_A_4EUYFJ4L3_1),.din(w_dff_A_ouFZAQwf3_1),.clk(gclk));
	jdff dff_A_I6UTQ0tw0_1(.dout(w_dff_A_ouFZAQwf3_1),.din(w_dff_A_I6UTQ0tw0_1),.clk(gclk));
	jdff dff_A_3o6uXX6Y4_1(.dout(w_dff_A_I6UTQ0tw0_1),.din(w_dff_A_3o6uXX6Y4_1),.clk(gclk));
	jdff dff_A_eQ2Nzjiz0_1(.dout(w_dff_A_3o6uXX6Y4_1),.din(w_dff_A_eQ2Nzjiz0_1),.clk(gclk));
	jdff dff_A_wEBWTMQW0_1(.dout(w_dff_A_eQ2Nzjiz0_1),.din(w_dff_A_wEBWTMQW0_1),.clk(gclk));
	jdff dff_A_JOMmBiyi7_1(.dout(w_dff_A_wEBWTMQW0_1),.din(w_dff_A_JOMmBiyi7_1),.clk(gclk));
	jdff dff_A_ypNZPoWa5_1(.dout(w_dff_A_JOMmBiyi7_1),.din(w_dff_A_ypNZPoWa5_1),.clk(gclk));
	jdff dff_A_Q05xcyJb8_1(.dout(w_dff_A_ypNZPoWa5_1),.din(w_dff_A_Q05xcyJb8_1),.clk(gclk));
	jdff dff_A_GQQrUn1Z3_1(.dout(w_dff_A_Q05xcyJb8_1),.din(w_dff_A_GQQrUn1Z3_1),.clk(gclk));
	jdff dff_A_DIcUxRg03_1(.dout(w_dff_A_GQQrUn1Z3_1),.din(w_dff_A_DIcUxRg03_1),.clk(gclk));
	jdff dff_A_sS5DdR5W9_1(.dout(w_dff_A_DIcUxRg03_1),.din(w_dff_A_sS5DdR5W9_1),.clk(gclk));
	jdff dff_A_RcDW4DBp8_1(.dout(w_dff_A_sS5DdR5W9_1),.din(w_dff_A_RcDW4DBp8_1),.clk(gclk));
	jdff dff_A_Q5T4PhPy6_1(.dout(w_dff_A_RcDW4DBp8_1),.din(w_dff_A_Q5T4PhPy6_1),.clk(gclk));
	jdff dff_A_wZLdBuM37_1(.dout(w_dff_A_Q5T4PhPy6_1),.din(w_dff_A_wZLdBuM37_1),.clk(gclk));
	jdff dff_A_DTuIgggF4_1(.dout(w_dff_A_wZLdBuM37_1),.din(w_dff_A_DTuIgggF4_1),.clk(gclk));
	jdff dff_A_4s07I5ZL8_1(.dout(w_dff_A_DTuIgggF4_1),.din(w_dff_A_4s07I5ZL8_1),.clk(gclk));
	jdff dff_A_XXMmGeEz2_1(.dout(w_dff_A_4s07I5ZL8_1),.din(w_dff_A_XXMmGeEz2_1),.clk(gclk));
	jdff dff_A_LAjly4nG4_1(.dout(w_dff_A_XXMmGeEz2_1),.din(w_dff_A_LAjly4nG4_1),.clk(gclk));
	jdff dff_A_asQoPrAi2_1(.dout(w_dff_A_LAjly4nG4_1),.din(w_dff_A_asQoPrAi2_1),.clk(gclk));
	jdff dff_A_nvVPJzbg4_1(.dout(w_dff_A_asQoPrAi2_1),.din(w_dff_A_nvVPJzbg4_1),.clk(gclk));
	jdff dff_A_L6992mk66_2(.dout(w_n1008_1[2]),.din(w_dff_A_L6992mk66_2),.clk(gclk));
	jdff dff_A_s5BfF6w16_2(.dout(w_dff_A_L6992mk66_2),.din(w_dff_A_s5BfF6w16_2),.clk(gclk));
	jdff dff_A_n6dlcIh69_2(.dout(w_dff_A_s5BfF6w16_2),.din(w_dff_A_n6dlcIh69_2),.clk(gclk));
	jdff dff_A_BGSjREbP3_2(.dout(w_dff_A_n6dlcIh69_2),.din(w_dff_A_BGSjREbP3_2),.clk(gclk));
	jdff dff_A_t0rquWFF1_2(.dout(w_dff_A_BGSjREbP3_2),.din(w_dff_A_t0rquWFF1_2),.clk(gclk));
	jdff dff_A_y5xFEzsz2_2(.dout(w_dff_A_t0rquWFF1_2),.din(w_dff_A_y5xFEzsz2_2),.clk(gclk));
	jdff dff_A_2ZlucQDn5_2(.dout(w_dff_A_y5xFEzsz2_2),.din(w_dff_A_2ZlucQDn5_2),.clk(gclk));
	jdff dff_A_KXEVUhWT2_2(.dout(w_dff_A_2ZlucQDn5_2),.din(w_dff_A_KXEVUhWT2_2),.clk(gclk));
	jdff dff_A_HlvbUxnE9_2(.dout(w_dff_A_KXEVUhWT2_2),.din(w_dff_A_HlvbUxnE9_2),.clk(gclk));
	jdff dff_A_SKyEw6Pd4_2(.dout(w_dff_A_HlvbUxnE9_2),.din(w_dff_A_SKyEw6Pd4_2),.clk(gclk));
	jdff dff_A_ByH6PFG89_2(.dout(w_dff_A_SKyEw6Pd4_2),.din(w_dff_A_ByH6PFG89_2),.clk(gclk));
	jdff dff_A_Z28xNWPq5_2(.dout(w_dff_A_ByH6PFG89_2),.din(w_dff_A_Z28xNWPq5_2),.clk(gclk));
	jdff dff_A_OZOfdAdC6_2(.dout(w_dff_A_Z28xNWPq5_2),.din(w_dff_A_OZOfdAdC6_2),.clk(gclk));
	jdff dff_A_Lxo8zdzp5_2(.dout(w_dff_A_OZOfdAdC6_2),.din(w_dff_A_Lxo8zdzp5_2),.clk(gclk));
	jdff dff_A_MCd0vN6K2_2(.dout(w_dff_A_Lxo8zdzp5_2),.din(w_dff_A_MCd0vN6K2_2),.clk(gclk));
	jdff dff_A_23t6YQOa0_2(.dout(w_dff_A_MCd0vN6K2_2),.din(w_dff_A_23t6YQOa0_2),.clk(gclk));
	jdff dff_A_pmVLIJvz9_2(.dout(w_dff_A_23t6YQOa0_2),.din(w_dff_A_pmVLIJvz9_2),.clk(gclk));
	jdff dff_A_PisEcUlx9_2(.dout(w_dff_A_pmVLIJvz9_2),.din(w_dff_A_PisEcUlx9_2),.clk(gclk));
	jdff dff_A_bxTVlKjW6_2(.dout(w_dff_A_PisEcUlx9_2),.din(w_dff_A_bxTVlKjW6_2),.clk(gclk));
	jdff dff_A_zLTOu8JK5_2(.dout(w_dff_A_bxTVlKjW6_2),.din(w_dff_A_zLTOu8JK5_2),.clk(gclk));
	jdff dff_A_mpLRE0Je6_1(.dout(w_n1008_0[1]),.din(w_dff_A_mpLRE0Je6_1),.clk(gclk));
	jdff dff_A_am7yIxmf3_1(.dout(w_dff_A_mpLRE0Je6_1),.din(w_dff_A_am7yIxmf3_1),.clk(gclk));
	jdff dff_A_rzsCQKzX1_1(.dout(w_dff_A_am7yIxmf3_1),.din(w_dff_A_rzsCQKzX1_1),.clk(gclk));
	jdff dff_A_egFPZ24v2_1(.dout(w_dff_A_rzsCQKzX1_1),.din(w_dff_A_egFPZ24v2_1),.clk(gclk));
	jdff dff_A_vzNTSyJY8_1(.dout(w_dff_A_egFPZ24v2_1),.din(w_dff_A_vzNTSyJY8_1),.clk(gclk));
	jdff dff_A_1pgYDBut5_1(.dout(w_dff_A_vzNTSyJY8_1),.din(w_dff_A_1pgYDBut5_1),.clk(gclk));
	jdff dff_A_FBWrHvsX9_1(.dout(w_dff_A_1pgYDBut5_1),.din(w_dff_A_FBWrHvsX9_1),.clk(gclk));
	jdff dff_A_8cEyKX9r7_1(.dout(w_dff_A_FBWrHvsX9_1),.din(w_dff_A_8cEyKX9r7_1),.clk(gclk));
	jdff dff_A_u2oM8zTL1_1(.dout(w_dff_A_8cEyKX9r7_1),.din(w_dff_A_u2oM8zTL1_1),.clk(gclk));
	jdff dff_A_kPBZg1MM1_1(.dout(w_dff_A_u2oM8zTL1_1),.din(w_dff_A_kPBZg1MM1_1),.clk(gclk));
	jdff dff_A_xr7TWG8s3_1(.dout(w_dff_A_kPBZg1MM1_1),.din(w_dff_A_xr7TWG8s3_1),.clk(gclk));
	jdff dff_A_MypX9fp29_1(.dout(w_dff_A_xr7TWG8s3_1),.din(w_dff_A_MypX9fp29_1),.clk(gclk));
	jdff dff_A_ePr8cnFI4_1(.dout(w_dff_A_MypX9fp29_1),.din(w_dff_A_ePr8cnFI4_1),.clk(gclk));
	jdff dff_A_WpdWctLV6_1(.dout(w_dff_A_ePr8cnFI4_1),.din(w_dff_A_WpdWctLV6_1),.clk(gclk));
	jdff dff_A_ZQuJxd5R4_1(.dout(w_dff_A_WpdWctLV6_1),.din(w_dff_A_ZQuJxd5R4_1),.clk(gclk));
	jdff dff_A_yuy19z7y0_1(.dout(w_dff_A_ZQuJxd5R4_1),.din(w_dff_A_yuy19z7y0_1),.clk(gclk));
	jdff dff_A_bOMjcM938_1(.dout(w_dff_A_yuy19z7y0_1),.din(w_dff_A_bOMjcM938_1),.clk(gclk));
	jdff dff_A_pkIOg8DR5_1(.dout(w_dff_A_bOMjcM938_1),.din(w_dff_A_pkIOg8DR5_1),.clk(gclk));
	jdff dff_A_VxFFKIej9_2(.dout(w_n1008_0[2]),.din(w_dff_A_VxFFKIej9_2),.clk(gclk));
	jdff dff_A_HqDQvGCU4_2(.dout(w_dff_A_VxFFKIej9_2),.din(w_dff_A_HqDQvGCU4_2),.clk(gclk));
	jdff dff_A_55ETpfEB6_2(.dout(w_dff_A_HqDQvGCU4_2),.din(w_dff_A_55ETpfEB6_2),.clk(gclk));
	jdff dff_A_9nnvYlqY6_2(.dout(w_dff_A_55ETpfEB6_2),.din(w_dff_A_9nnvYlqY6_2),.clk(gclk));
	jdff dff_A_BFUe0ssz2_2(.dout(w_dff_A_9nnvYlqY6_2),.din(w_dff_A_BFUe0ssz2_2),.clk(gclk));
	jdff dff_A_ez6mDYfh9_2(.dout(w_dff_A_BFUe0ssz2_2),.din(w_dff_A_ez6mDYfh9_2),.clk(gclk));
	jdff dff_A_XzE95zm61_2(.dout(w_dff_A_ez6mDYfh9_2),.din(w_dff_A_XzE95zm61_2),.clk(gclk));
	jdff dff_A_XhWeXWgj3_2(.dout(w_dff_A_XzE95zm61_2),.din(w_dff_A_XhWeXWgj3_2),.clk(gclk));
	jdff dff_A_uV4raij88_2(.dout(w_dff_A_XhWeXWgj3_2),.din(w_dff_A_uV4raij88_2),.clk(gclk));
	jdff dff_A_8EB01zUN2_2(.dout(w_dff_A_uV4raij88_2),.din(w_dff_A_8EB01zUN2_2),.clk(gclk));
	jdff dff_A_d18Xh9zG0_2(.dout(w_dff_A_8EB01zUN2_2),.din(w_dff_A_d18Xh9zG0_2),.clk(gclk));
	jdff dff_A_4E7c0JBK7_1(.dout(w_G1691_5[1]),.din(w_dff_A_4E7c0JBK7_1),.clk(gclk));
	jdff dff_A_WLJRdjkR5_1(.dout(w_dff_A_4E7c0JBK7_1),.din(w_dff_A_WLJRdjkR5_1),.clk(gclk));
	jdff dff_A_JQwaCszr1_1(.dout(w_dff_A_WLJRdjkR5_1),.din(w_dff_A_JQwaCszr1_1),.clk(gclk));
	jdff dff_A_GbYZZhVE4_1(.dout(w_dff_A_JQwaCszr1_1),.din(w_dff_A_GbYZZhVE4_1),.clk(gclk));
	jdff dff_A_OkmxD4018_1(.dout(w_dff_A_GbYZZhVE4_1),.din(w_dff_A_OkmxD4018_1),.clk(gclk));
	jdff dff_A_gdG4XFfr2_1(.dout(w_dff_A_OkmxD4018_1),.din(w_dff_A_gdG4XFfr2_1),.clk(gclk));
	jdff dff_A_WnK7dBLg2_1(.dout(w_dff_A_gdG4XFfr2_1),.din(w_dff_A_WnK7dBLg2_1),.clk(gclk));
	jdff dff_A_kORXSVfs4_1(.dout(w_dff_A_WnK7dBLg2_1),.din(w_dff_A_kORXSVfs4_1),.clk(gclk));
	jdff dff_A_RC3RjUy58_1(.dout(w_dff_A_kORXSVfs4_1),.din(w_dff_A_RC3RjUy58_1),.clk(gclk));
	jdff dff_B_vYP787lz7_2(.din(n1698),.dout(w_dff_B_vYP787lz7_2),.clk(gclk));
	jdff dff_B_dv0Sk1rx6_2(.din(w_dff_B_vYP787lz7_2),.dout(w_dff_B_dv0Sk1rx6_2),.clk(gclk));
	jdff dff_A_JyTimGTZ8_1(.dout(w_G1694_0[1]),.din(w_dff_A_JyTimGTZ8_1),.clk(gclk));
	jdff dff_A_tgSDKJZS0_1(.dout(w_dff_A_JyTimGTZ8_1),.din(w_dff_A_tgSDKJZS0_1),.clk(gclk));
	jdff dff_A_2FMNP6gm3_1(.dout(w_dff_A_tgSDKJZS0_1),.din(w_dff_A_2FMNP6gm3_1),.clk(gclk));
	jdff dff_A_SlXD9Zaz1_1(.dout(w_dff_A_2FMNP6gm3_1),.din(w_dff_A_SlXD9Zaz1_1),.clk(gclk));
	jdff dff_A_4YxIrAtO3_1(.dout(w_dff_A_SlXD9Zaz1_1),.din(w_dff_A_4YxIrAtO3_1),.clk(gclk));
	jdff dff_A_DR8HT2Cz2_1(.dout(w_dff_A_4YxIrAtO3_1),.din(w_dff_A_DR8HT2Cz2_1),.clk(gclk));
	jdff dff_A_UqXC2gA67_1(.dout(w_dff_A_DR8HT2Cz2_1),.din(w_dff_A_UqXC2gA67_1),.clk(gclk));
	jdff dff_A_7Aw2yds87_1(.dout(w_dff_A_UqXC2gA67_1),.din(w_dff_A_7Aw2yds87_1),.clk(gclk));
	jdff dff_A_BSpXy12l8_1(.dout(w_dff_A_7Aw2yds87_1),.din(w_dff_A_BSpXy12l8_1),.clk(gclk));
	jdff dff_A_bxIaF5Z25_1(.dout(w_dff_A_BSpXy12l8_1),.din(w_dff_A_bxIaF5Z25_1),.clk(gclk));
	jdff dff_A_ol4IIpzV2_1(.dout(w_dff_A_bxIaF5Z25_1),.din(w_dff_A_ol4IIpzV2_1),.clk(gclk));
	jdff dff_A_K6JfdkhC0_1(.dout(w_dff_A_ol4IIpzV2_1),.din(w_dff_A_K6JfdkhC0_1),.clk(gclk));
	jdff dff_A_9A60RQXf2_1(.dout(w_dff_A_K6JfdkhC0_1),.din(w_dff_A_9A60RQXf2_1),.clk(gclk));
	jdff dff_A_OMbpm80E8_1(.dout(w_dff_A_9A60RQXf2_1),.din(w_dff_A_OMbpm80E8_1),.clk(gclk));
	jdff dff_A_i55synqN9_1(.dout(w_dff_A_OMbpm80E8_1),.din(w_dff_A_i55synqN9_1),.clk(gclk));
	jdff dff_A_QmNlyXPh1_1(.dout(w_dff_A_i55synqN9_1),.din(w_dff_A_QmNlyXPh1_1),.clk(gclk));
	jdff dff_A_PIsCQWs12_1(.dout(w_dff_A_QmNlyXPh1_1),.din(w_dff_A_PIsCQWs12_1),.clk(gclk));
	jdff dff_A_9iITZDPc3_1(.dout(w_dff_A_PIsCQWs12_1),.din(w_dff_A_9iITZDPc3_1),.clk(gclk));
	jdff dff_A_aaRdwr1T9_1(.dout(w_dff_A_9iITZDPc3_1),.din(w_dff_A_aaRdwr1T9_1),.clk(gclk));
	jdff dff_A_5zpX7mQT5_1(.dout(w_dff_A_aaRdwr1T9_1),.din(w_dff_A_5zpX7mQT5_1),.clk(gclk));
	jdff dff_A_MCoDUxPh8_1(.dout(w_dff_A_5zpX7mQT5_1),.din(w_dff_A_MCoDUxPh8_1),.clk(gclk));
	jdff dff_A_4JolZxLh1_1(.dout(w_dff_A_MCoDUxPh8_1),.din(w_dff_A_4JolZxLh1_1),.clk(gclk));
	jdff dff_A_MVuEkKuY4_1(.dout(w_dff_A_4JolZxLh1_1),.din(w_dff_A_MVuEkKuY4_1),.clk(gclk));
	jdff dff_A_VuDmMeGV7_2(.dout(w_G1694_0[2]),.din(w_dff_A_VuDmMeGV7_2),.clk(gclk));
	jdff dff_A_Jk7SZmKU1_0(.dout(w_G1691_4[0]),.din(w_dff_A_Jk7SZmKU1_0),.clk(gclk));
	jdff dff_A_FKs06vOf6_0(.dout(w_dff_A_Jk7SZmKU1_0),.din(w_dff_A_FKs06vOf6_0),.clk(gclk));
	jdff dff_A_m97GAm8A1_0(.dout(w_dff_A_FKs06vOf6_0),.din(w_dff_A_m97GAm8A1_0),.clk(gclk));
	jdff dff_A_jc7UkP114_0(.dout(w_dff_A_m97GAm8A1_0),.din(w_dff_A_jc7UkP114_0),.clk(gclk));
	jdff dff_A_caH9ZvRL1_0(.dout(w_dff_A_jc7UkP114_0),.din(w_dff_A_caH9ZvRL1_0),.clk(gclk));
	jdff dff_A_kElsjG2o5_0(.dout(w_dff_A_caH9ZvRL1_0),.din(w_dff_A_kElsjG2o5_0),.clk(gclk));
	jdff dff_A_ryM8UOrg9_0(.dout(w_dff_A_kElsjG2o5_0),.din(w_dff_A_ryM8UOrg9_0),.clk(gclk));
	jdff dff_A_DU3H0pKq2_0(.dout(w_dff_A_ryM8UOrg9_0),.din(w_dff_A_DU3H0pKq2_0),.clk(gclk));
	jdff dff_A_Zw2VpOzO0_0(.dout(w_dff_A_DU3H0pKq2_0),.din(w_dff_A_Zw2VpOzO0_0),.clk(gclk));
	jdff dff_A_ZSJKYVm82_0(.dout(w_dff_A_Zw2VpOzO0_0),.din(w_dff_A_ZSJKYVm82_0),.clk(gclk));
	jdff dff_A_hjgvEmeW6_0(.dout(w_dff_A_ZSJKYVm82_0),.din(w_dff_A_hjgvEmeW6_0),.clk(gclk));
	jdff dff_A_azay8LDz1_0(.dout(w_dff_A_hjgvEmeW6_0),.din(w_dff_A_azay8LDz1_0),.clk(gclk));
	jdff dff_A_AK73ZF6E9_0(.dout(w_dff_A_azay8LDz1_0),.din(w_dff_A_AK73ZF6E9_0),.clk(gclk));
	jdff dff_A_9EMamk5B2_0(.dout(w_dff_A_AK73ZF6E9_0),.din(w_dff_A_9EMamk5B2_0),.clk(gclk));
	jdff dff_A_7P1JnGap3_1(.dout(w_G1691_4[1]),.din(w_dff_A_7P1JnGap3_1),.clk(gclk));
	jdff dff_A_VA0e6dU49_1(.dout(w_dff_A_7P1JnGap3_1),.din(w_dff_A_VA0e6dU49_1),.clk(gclk));
	jdff dff_A_3gBVCCOo6_1(.dout(w_dff_A_VA0e6dU49_1),.din(w_dff_A_3gBVCCOo6_1),.clk(gclk));
	jdff dff_A_En2PdWcd5_1(.dout(w_dff_A_3gBVCCOo6_1),.din(w_dff_A_En2PdWcd5_1),.clk(gclk));
	jdff dff_A_cDENqyZV9_1(.dout(w_dff_A_En2PdWcd5_1),.din(w_dff_A_cDENqyZV9_1),.clk(gclk));
	jdff dff_A_QmRFrdBT0_1(.dout(w_dff_A_cDENqyZV9_1),.din(w_dff_A_QmRFrdBT0_1),.clk(gclk));
	jdff dff_A_zukXn5n45_1(.dout(w_dff_A_QmRFrdBT0_1),.din(w_dff_A_zukXn5n45_1),.clk(gclk));
	jdff dff_A_THYbqjPJ2_1(.dout(w_dff_A_zukXn5n45_1),.din(w_dff_A_THYbqjPJ2_1),.clk(gclk));
	jdff dff_A_6kFmL9K90_1(.dout(w_dff_A_THYbqjPJ2_1),.din(w_dff_A_6kFmL9K90_1),.clk(gclk));
	jdff dff_A_MDqysnyc5_1(.dout(w_dff_A_6kFmL9K90_1),.din(w_dff_A_MDqysnyc5_1),.clk(gclk));
	jdff dff_A_jJf4eWaU4_1(.dout(w_dff_A_MDqysnyc5_1),.din(w_dff_A_jJf4eWaU4_1),.clk(gclk));
	jdff dff_A_eKR2wk7F9_1(.dout(w_dff_A_jJf4eWaU4_1),.din(w_dff_A_eKR2wk7F9_1),.clk(gclk));
	jdff dff_A_4PRyniVS0_1(.dout(w_dff_A_eKR2wk7F9_1),.din(w_dff_A_4PRyniVS0_1),.clk(gclk));
	jdff dff_A_oc9mtfTm5_1(.dout(w_dff_A_4PRyniVS0_1),.din(w_dff_A_oc9mtfTm5_1),.clk(gclk));
	jdff dff_A_SRXyEb8c0_1(.dout(w_dff_A_oc9mtfTm5_1),.din(w_dff_A_SRXyEb8c0_1),.clk(gclk));
	jdff dff_A_gA8plgWv0_1(.dout(w_dff_A_SRXyEb8c0_1),.din(w_dff_A_gA8plgWv0_1),.clk(gclk));
	jdff dff_A_nAlCE6Zu1_2(.dout(w_G1691_1[2]),.din(w_dff_A_nAlCE6Zu1_2),.clk(gclk));
	jdff dff_A_tONs35pE1_2(.dout(w_dff_A_nAlCE6Zu1_2),.din(w_dff_A_tONs35pE1_2),.clk(gclk));
	jdff dff_A_H0ENVOgR9_2(.dout(w_dff_A_tONs35pE1_2),.din(w_dff_A_H0ENVOgR9_2),.clk(gclk));
	jdff dff_A_OYPEqwMm4_2(.dout(w_dff_A_H0ENVOgR9_2),.din(w_dff_A_OYPEqwMm4_2),.clk(gclk));
	jdff dff_A_8z4UllSI9_2(.dout(w_dff_A_OYPEqwMm4_2),.din(w_dff_A_8z4UllSI9_2),.clk(gclk));
	jdff dff_A_ttefBYj68_2(.dout(w_dff_A_8z4UllSI9_2),.din(w_dff_A_ttefBYj68_2),.clk(gclk));
	jdff dff_A_XtqX9Khd7_2(.dout(w_dff_A_ttefBYj68_2),.din(w_dff_A_XtqX9Khd7_2),.clk(gclk));
	jdff dff_A_Qy9KWbIF1_2(.dout(w_dff_A_XtqX9Khd7_2),.din(w_dff_A_Qy9KWbIF1_2),.clk(gclk));
	jdff dff_A_nKzJime58_2(.dout(w_dff_A_Qy9KWbIF1_2),.din(w_dff_A_nKzJime58_2),.clk(gclk));
	jdff dff_A_s8CsorvS4_2(.dout(w_dff_A_nKzJime58_2),.din(w_dff_A_s8CsorvS4_2),.clk(gclk));
	jdff dff_A_0DJTXydb5_2(.dout(w_dff_A_s8CsorvS4_2),.din(w_dff_A_0DJTXydb5_2),.clk(gclk));
	jdff dff_A_HxUoWY1V0_2(.dout(w_dff_A_0DJTXydb5_2),.din(w_dff_A_HxUoWY1V0_2),.clk(gclk));
	jdff dff_A_r4M3zkXA1_2(.dout(w_dff_A_HxUoWY1V0_2),.din(w_dff_A_r4M3zkXA1_2),.clk(gclk));
	jdff dff_A_TMOLMh414_2(.dout(w_dff_A_r4M3zkXA1_2),.din(w_dff_A_TMOLMh414_2),.clk(gclk));
	jdff dff_A_YaTrhLx00_2(.dout(w_dff_A_TMOLMh414_2),.din(w_dff_A_YaTrhLx00_2),.clk(gclk));
	jdff dff_A_Cw34PnhY4_2(.dout(w_dff_A_YaTrhLx00_2),.din(w_dff_A_Cw34PnhY4_2),.clk(gclk));
	jdff dff_A_jtW2qP6v7_2(.dout(w_dff_A_Cw34PnhY4_2),.din(w_dff_A_jtW2qP6v7_2),.clk(gclk));
	jdff dff_A_bQxer46m5_2(.dout(w_dff_A_jtW2qP6v7_2),.din(w_dff_A_bQxer46m5_2),.clk(gclk));
	jdff dff_A_3n4sw47y0_2(.dout(w_dff_A_bQxer46m5_2),.din(w_dff_A_3n4sw47y0_2),.clk(gclk));
	jdff dff_A_2udhEhhk6_2(.dout(w_dff_A_3n4sw47y0_2),.din(w_dff_A_2udhEhhk6_2),.clk(gclk));
	jdff dff_A_ZGOI0Qfx5_2(.dout(w_dff_A_2udhEhhk6_2),.din(w_dff_A_ZGOI0Qfx5_2),.clk(gclk));
	jdff dff_A_qR4PjBAd9_2(.dout(w_dff_A_ZGOI0Qfx5_2),.din(w_dff_A_qR4PjBAd9_2),.clk(gclk));
	jdff dff_A_PSVaiqWh9_1(.dout(w_G1691_0[1]),.din(w_dff_A_PSVaiqWh9_1),.clk(gclk));
	jdff dff_A_Q0BsbUps8_1(.dout(w_dff_A_PSVaiqWh9_1),.din(w_dff_A_Q0BsbUps8_1),.clk(gclk));
	jdff dff_A_bHyQFTVD8_1(.dout(w_dff_A_Q0BsbUps8_1),.din(w_dff_A_bHyQFTVD8_1),.clk(gclk));
	jdff dff_A_tSy389Iw5_1(.dout(w_dff_A_bHyQFTVD8_1),.din(w_dff_A_tSy389Iw5_1),.clk(gclk));
	jdff dff_A_ZdkB8XYl8_1(.dout(w_dff_A_tSy389Iw5_1),.din(w_dff_A_ZdkB8XYl8_1),.clk(gclk));
	jdff dff_A_a2PHSSgC0_1(.dout(w_dff_A_ZdkB8XYl8_1),.din(w_dff_A_a2PHSSgC0_1),.clk(gclk));
	jdff dff_A_4y1WoQs30_1(.dout(w_dff_A_a2PHSSgC0_1),.din(w_dff_A_4y1WoQs30_1),.clk(gclk));
	jdff dff_A_u1wMxsoM7_1(.dout(w_dff_A_4y1WoQs30_1),.din(w_dff_A_u1wMxsoM7_1),.clk(gclk));
	jdff dff_A_RnSWeJMG5_1(.dout(w_dff_A_u1wMxsoM7_1),.din(w_dff_A_RnSWeJMG5_1),.clk(gclk));
	jdff dff_A_ZFfkZLAp9_1(.dout(w_dff_A_RnSWeJMG5_1),.din(w_dff_A_ZFfkZLAp9_1),.clk(gclk));
	jdff dff_A_CINpUQmP2_1(.dout(w_dff_A_ZFfkZLAp9_1),.din(w_dff_A_CINpUQmP2_1),.clk(gclk));
	jdff dff_A_wfKobEfZ0_1(.dout(w_dff_A_CINpUQmP2_1),.din(w_dff_A_wfKobEfZ0_1),.clk(gclk));
	jdff dff_A_xOC9gKt38_1(.dout(w_dff_A_wfKobEfZ0_1),.din(w_dff_A_xOC9gKt38_1),.clk(gclk));
	jdff dff_A_QzWa2Z5n5_1(.dout(w_dff_A_xOC9gKt38_1),.din(w_dff_A_QzWa2Z5n5_1),.clk(gclk));
	jdff dff_A_ZjwBPAsB1_1(.dout(w_dff_A_QzWa2Z5n5_1),.din(w_dff_A_ZjwBPAsB1_1),.clk(gclk));
	jdff dff_A_9Fnp6qaA7_1(.dout(w_dff_A_ZjwBPAsB1_1),.din(w_dff_A_9Fnp6qaA7_1),.clk(gclk));
	jdff dff_A_CGO9D06C0_1(.dout(w_dff_A_9Fnp6qaA7_1),.din(w_dff_A_CGO9D06C0_1),.clk(gclk));
	jdff dff_A_S1zFmDVS4_1(.dout(w_dff_A_CGO9D06C0_1),.din(w_dff_A_S1zFmDVS4_1),.clk(gclk));
	jdff dff_A_1UZ6pyuM0_1(.dout(w_dff_A_S1zFmDVS4_1),.din(w_dff_A_1UZ6pyuM0_1),.clk(gclk));
	jdff dff_A_OZQKo4iO6_2(.dout(w_G1691_0[2]),.din(w_dff_A_OZQKo4iO6_2),.clk(gclk));
	jdff dff_A_c1b1bM6v6_2(.dout(w_dff_A_OZQKo4iO6_2),.din(w_dff_A_c1b1bM6v6_2),.clk(gclk));
	jdff dff_A_N5q6kPc40_2(.dout(w_dff_A_c1b1bM6v6_2),.din(w_dff_A_N5q6kPc40_2),.clk(gclk));
	jdff dff_A_UxubReMS9_2(.dout(w_dff_A_N5q6kPc40_2),.din(w_dff_A_UxubReMS9_2),.clk(gclk));
	jdff dff_A_pgvIfkwn4_2(.dout(w_dff_A_UxubReMS9_2),.din(w_dff_A_pgvIfkwn4_2),.clk(gclk));
	jdff dff_A_8tNVIIbT6_2(.dout(w_dff_A_pgvIfkwn4_2),.din(w_dff_A_8tNVIIbT6_2),.clk(gclk));
	jdff dff_A_uuwaA6sV0_2(.dout(w_dff_A_8tNVIIbT6_2),.din(w_dff_A_uuwaA6sV0_2),.clk(gclk));
	jdff dff_A_ZQsuTpCw2_2(.dout(w_dff_A_uuwaA6sV0_2),.din(w_dff_A_ZQsuTpCw2_2),.clk(gclk));
	jdff dff_A_A5cFD2H06_2(.dout(w_dff_A_ZQsuTpCw2_2),.din(w_dff_A_A5cFD2H06_2),.clk(gclk));
	jdff dff_A_HXPeOfLY2_2(.dout(w_dff_A_A5cFD2H06_2),.din(w_dff_A_HXPeOfLY2_2),.clk(gclk));
	jdff dff_A_REPLKCAk0_2(.dout(w_dff_A_HXPeOfLY2_2),.din(w_dff_A_REPLKCAk0_2),.clk(gclk));
	jdff dff_A_s6N5LyGp7_2(.dout(w_dff_A_REPLKCAk0_2),.din(w_dff_A_s6N5LyGp7_2),.clk(gclk));
	jdff dff_A_vIIwWw7D2_2(.dout(w_dff_A_s6N5LyGp7_2),.din(w_dff_A_vIIwWw7D2_2),.clk(gclk));
	jdff dff_B_poQPHa3h8_2(.din(n1695),.dout(w_dff_B_poQPHa3h8_2),.clk(gclk));
	jdff dff_B_9f5pCFcU7_2(.din(n1694),.dout(w_dff_B_9f5pCFcU7_2),.clk(gclk));
	jdff dff_B_YVCPnw5W1_2(.din(w_dff_B_9f5pCFcU7_2),.dout(w_dff_B_YVCPnw5W1_2),.clk(gclk));
	jdff dff_B_03d0JNAd2_2(.din(w_dff_B_YVCPnw5W1_2),.dout(w_dff_B_03d0JNAd2_2),.clk(gclk));
	jdff dff_B_wxCaaXBG2_2(.din(w_dff_B_03d0JNAd2_2),.dout(w_dff_B_wxCaaXBG2_2),.clk(gclk));
	jdff dff_B_cTF7mqUj3_2(.din(w_dff_B_wxCaaXBG2_2),.dout(w_dff_B_cTF7mqUj3_2),.clk(gclk));
	jdff dff_B_3Z9z2qyF9_2(.din(w_dff_B_cTF7mqUj3_2),.dout(w_dff_B_3Z9z2qyF9_2),.clk(gclk));
	jdff dff_B_WO8yaWsY6_2(.din(w_dff_B_3Z9z2qyF9_2),.dout(w_dff_B_WO8yaWsY6_2),.clk(gclk));
	jdff dff_B_G7S84XVG2_2(.din(w_dff_B_WO8yaWsY6_2),.dout(w_dff_B_G7S84XVG2_2),.clk(gclk));
	jdff dff_B_F4ejeGlL8_2(.din(w_dff_B_G7S84XVG2_2),.dout(w_dff_B_F4ejeGlL8_2),.clk(gclk));
	jdff dff_B_gAbkvH4z9_2(.din(w_dff_B_F4ejeGlL8_2),.dout(w_dff_B_gAbkvH4z9_2),.clk(gclk));
	jdff dff_B_lzassceA1_2(.din(w_dff_B_gAbkvH4z9_2),.dout(w_dff_B_lzassceA1_2),.clk(gclk));
	jdff dff_B_prZSGH047_2(.din(w_dff_B_lzassceA1_2),.dout(w_dff_B_prZSGH047_2),.clk(gclk));
	jdff dff_B_YpQaawxc3_2(.din(w_dff_B_prZSGH047_2),.dout(w_dff_B_YpQaawxc3_2),.clk(gclk));
	jdff dff_B_touOMwKo6_2(.din(w_dff_B_YpQaawxc3_2),.dout(w_dff_B_touOMwKo6_2),.clk(gclk));
	jdff dff_B_I22Xh09X7_2(.din(w_dff_B_touOMwKo6_2),.dout(w_dff_B_I22Xh09X7_2),.clk(gclk));
	jdff dff_B_UnqBlSJv9_2(.din(w_dff_B_I22Xh09X7_2),.dout(w_dff_B_UnqBlSJv9_2),.clk(gclk));
	jdff dff_B_UUV3vhOh6_2(.din(w_dff_B_UnqBlSJv9_2),.dout(w_dff_B_UUV3vhOh6_2),.clk(gclk));
	jdff dff_B_ocsGrU6Y3_2(.din(w_dff_B_UUV3vhOh6_2),.dout(w_dff_B_ocsGrU6Y3_2),.clk(gclk));
	jdff dff_B_T64IbHBO2_2(.din(w_dff_B_ocsGrU6Y3_2),.dout(w_dff_B_T64IbHBO2_2),.clk(gclk));
	jdff dff_B_N35Ki1o12_2(.din(w_dff_B_T64IbHBO2_2),.dout(w_dff_B_N35Ki1o12_2),.clk(gclk));
	jdff dff_B_eI2nSmHx0_2(.din(w_dff_B_N35Ki1o12_2),.dout(w_dff_B_eI2nSmHx0_2),.clk(gclk));
	jdff dff_B_oJDt5xgE5_2(.din(w_dff_B_eI2nSmHx0_2),.dout(w_dff_B_oJDt5xgE5_2),.clk(gclk));
	jdff dff_B_ieX59DMA8_2(.din(w_dff_B_oJDt5xgE5_2),.dout(w_dff_B_ieX59DMA8_2),.clk(gclk));
	jdff dff_B_LB8SAABg1_2(.din(w_dff_B_ieX59DMA8_2),.dout(w_dff_B_LB8SAABg1_2),.clk(gclk));
	jdff dff_B_I3xFUquT7_2(.din(w_dff_B_LB8SAABg1_2),.dout(w_dff_B_I3xFUquT7_2),.clk(gclk));
	jdff dff_B_njf0WG6e3_2(.din(w_dff_B_I3xFUquT7_2),.dout(w_dff_B_njf0WG6e3_2),.clk(gclk));
	jdff dff_A_5643B7op6_2(.dout(w_G137_3[2]),.din(w_dff_A_5643B7op6_2),.clk(gclk));
	jdff dff_A_1Mm6hNVS3_2(.dout(w_dff_A_5643B7op6_2),.din(w_dff_A_1Mm6hNVS3_2),.clk(gclk));
	jdff dff_A_QFt1YS2g4_2(.dout(w_dff_A_1Mm6hNVS3_2),.din(w_dff_A_QFt1YS2g4_2),.clk(gclk));
	jdff dff_A_qLNO8SMa7_2(.dout(w_dff_A_QFt1YS2g4_2),.din(w_dff_A_qLNO8SMa7_2),.clk(gclk));
	jdff dff_A_6wQ9wlX69_2(.dout(w_dff_A_qLNO8SMa7_2),.din(w_dff_A_6wQ9wlX69_2),.clk(gclk));
	jdff dff_A_rh9CCW4X3_2(.dout(w_dff_A_6wQ9wlX69_2),.din(w_dff_A_rh9CCW4X3_2),.clk(gclk));
	jdff dff_A_HY8txvO21_2(.dout(w_dff_A_rh9CCW4X3_2),.din(w_dff_A_HY8txvO21_2),.clk(gclk));
	jdff dff_A_azKJV0qw6_2(.dout(w_dff_A_HY8txvO21_2),.din(w_dff_A_azKJV0qw6_2),.clk(gclk));
	jdff dff_A_OyQiFhFZ3_2(.dout(w_dff_A_azKJV0qw6_2),.din(w_dff_A_OyQiFhFZ3_2),.clk(gclk));
	jdff dff_A_J24N0Do60_2(.dout(w_dff_A_OyQiFhFZ3_2),.din(w_dff_A_J24N0Do60_2),.clk(gclk));
	jdff dff_A_5KMFeiJ76_2(.dout(w_dff_A_J24N0Do60_2),.din(w_dff_A_5KMFeiJ76_2),.clk(gclk));
	jdff dff_A_WuSZRG9k6_2(.dout(w_dff_A_5KMFeiJ76_2),.din(w_dff_A_WuSZRG9k6_2),.clk(gclk));
	jdff dff_A_7FYlEURy4_2(.dout(w_dff_A_WuSZRG9k6_2),.din(w_dff_A_7FYlEURy4_2),.clk(gclk));
	jdff dff_A_5pDfpnE62_2(.dout(w_dff_A_7FYlEURy4_2),.din(w_dff_A_5pDfpnE62_2),.clk(gclk));
	jdff dff_A_scV9Pi6d3_2(.dout(w_dff_A_5pDfpnE62_2),.din(w_dff_A_scV9Pi6d3_2),.clk(gclk));
	jdff dff_A_4JKI4OUM2_2(.dout(w_dff_A_scV9Pi6d3_2),.din(w_dff_A_4JKI4OUM2_2),.clk(gclk));
	jdff dff_A_aG4fRHmC3_2(.dout(w_dff_A_4JKI4OUM2_2),.din(w_dff_A_aG4fRHmC3_2),.clk(gclk));
	jdff dff_A_Ddc85VlV1_2(.dout(w_dff_A_aG4fRHmC3_2),.din(w_dff_A_Ddc85VlV1_2),.clk(gclk));
	jdff dff_A_ZnZQwgwF9_2(.dout(w_dff_A_Ddc85VlV1_2),.din(w_dff_A_ZnZQwgwF9_2),.clk(gclk));
	jdff dff_A_Md0HSSz69_2(.dout(w_dff_A_ZnZQwgwF9_2),.din(w_dff_A_Md0HSSz69_2),.clk(gclk));
	jdff dff_A_POH6v1gU4_2(.dout(w_dff_A_Md0HSSz69_2),.din(w_dff_A_POH6v1gU4_2),.clk(gclk));
	jdff dff_A_nMEdVV4X7_2(.dout(w_dff_A_POH6v1gU4_2),.din(w_dff_A_nMEdVV4X7_2),.clk(gclk));
	jdff dff_A_6fVhreec5_2(.dout(w_dff_A_nMEdVV4X7_2),.din(w_dff_A_6fVhreec5_2),.clk(gclk));
	jdff dff_A_ggIDazgF3_2(.dout(w_dff_A_6fVhreec5_2),.din(w_dff_A_ggIDazgF3_2),.clk(gclk));
	jdff dff_A_MDteAlzh1_0(.dout(w_G137_0[0]),.din(w_dff_A_MDteAlzh1_0),.clk(gclk));
	jdff dff_A_OjM5MU2Y3_0(.dout(w_dff_A_MDteAlzh1_0),.din(w_dff_A_OjM5MU2Y3_0),.clk(gclk));
	jdff dff_A_r64M6Z4L3_0(.dout(w_dff_A_OjM5MU2Y3_0),.din(w_dff_A_r64M6Z4L3_0),.clk(gclk));
	jdff dff_A_b6XHtIlt2_0(.dout(w_dff_A_r64M6Z4L3_0),.din(w_dff_A_b6XHtIlt2_0),.clk(gclk));
	jdff dff_A_vWktkhc98_0(.dout(w_dff_A_b6XHtIlt2_0),.din(w_dff_A_vWktkhc98_0),.clk(gclk));
	jdff dff_A_jzLh2cW58_0(.dout(w_dff_A_vWktkhc98_0),.din(w_dff_A_jzLh2cW58_0),.clk(gclk));
	jdff dff_A_crX2azFC6_0(.dout(w_dff_A_jzLh2cW58_0),.din(w_dff_A_crX2azFC6_0),.clk(gclk));
	jdff dff_A_yOE54uKE6_0(.dout(w_dff_A_crX2azFC6_0),.din(w_dff_A_yOE54uKE6_0),.clk(gclk));
	jdff dff_A_Rv8TeEZj6_0(.dout(w_dff_A_yOE54uKE6_0),.din(w_dff_A_Rv8TeEZj6_0),.clk(gclk));
	jdff dff_A_sw2wXDE82_0(.dout(w_dff_A_Rv8TeEZj6_0),.din(w_dff_A_sw2wXDE82_0),.clk(gclk));
	jdff dff_A_9V0ji26O5_0(.dout(w_dff_A_sw2wXDE82_0),.din(w_dff_A_9V0ji26O5_0),.clk(gclk));
	jdff dff_A_lMp6oV2H2_0(.dout(w_dff_A_9V0ji26O5_0),.din(w_dff_A_lMp6oV2H2_0),.clk(gclk));
	jdff dff_A_mI4bnq797_0(.dout(w_dff_A_lMp6oV2H2_0),.din(w_dff_A_mI4bnq797_0),.clk(gclk));
	jdff dff_A_8PRL8ZI45_0(.dout(w_dff_A_mI4bnq797_0),.din(w_dff_A_8PRL8ZI45_0),.clk(gclk));
	jdff dff_A_JlWSIpyw7_0(.dout(w_dff_A_8PRL8ZI45_0),.din(w_dff_A_JlWSIpyw7_0),.clk(gclk));
	jdff dff_A_5bAthwJX1_0(.dout(w_dff_A_JlWSIpyw7_0),.din(w_dff_A_5bAthwJX1_0),.clk(gclk));
	jdff dff_A_x4dZmg6f6_0(.dout(w_dff_A_5bAthwJX1_0),.din(w_dff_A_x4dZmg6f6_0),.clk(gclk));
	jdff dff_A_nQdMsAbm8_1(.dout(w_G137_0[1]),.din(w_dff_A_nQdMsAbm8_1),.clk(gclk));
	jdff dff_A_XX5yG7cJ0_1(.dout(w_dff_A_nQdMsAbm8_1),.din(w_dff_A_XX5yG7cJ0_1),.clk(gclk));
	jdff dff_A_zuaPrjdN7_1(.dout(w_dff_A_XX5yG7cJ0_1),.din(w_dff_A_zuaPrjdN7_1),.clk(gclk));
	jdff dff_A_QHhwW1gN1_1(.dout(w_dff_A_zuaPrjdN7_1),.din(w_dff_A_QHhwW1gN1_1),.clk(gclk));
	jdff dff_A_SJG7vEhs8_1(.dout(w_dff_A_QHhwW1gN1_1),.din(w_dff_A_SJG7vEhs8_1),.clk(gclk));
	jdff dff_A_gKQP4ugM2_1(.dout(w_dff_A_SJG7vEhs8_1),.din(w_dff_A_gKQP4ugM2_1),.clk(gclk));
	jdff dff_A_9JUSLCV17_1(.dout(w_dff_A_gKQP4ugM2_1),.din(w_dff_A_9JUSLCV17_1),.clk(gclk));
	jdff dff_A_wkBd0UsZ7_1(.dout(w_dff_A_9JUSLCV17_1),.din(w_dff_A_wkBd0UsZ7_1),.clk(gclk));
	jdff dff_A_cibIhkzl2_1(.dout(w_dff_A_wkBd0UsZ7_1),.din(w_dff_A_cibIhkzl2_1),.clk(gclk));
	jdff dff_A_khUFWdNW0_1(.dout(w_dff_A_cibIhkzl2_1),.din(w_dff_A_khUFWdNW0_1),.clk(gclk));
	jdff dff_A_HLjqzoFC3_1(.dout(w_dff_A_khUFWdNW0_1),.din(w_dff_A_HLjqzoFC3_1),.clk(gclk));
	jdff dff_A_j4YTQQb54_1(.dout(w_dff_A_HLjqzoFC3_1),.din(w_dff_A_j4YTQQb54_1),.clk(gclk));
	jdff dff_A_c02mr9Nj5_1(.dout(w_dff_A_j4YTQQb54_1),.din(w_dff_A_c02mr9Nj5_1),.clk(gclk));
	jdff dff_A_BpFCaTCQ1_1(.dout(w_dff_A_c02mr9Nj5_1),.din(w_dff_A_BpFCaTCQ1_1),.clk(gclk));
	jdff dff_A_tQnXJQLk8_1(.dout(w_dff_A_BpFCaTCQ1_1),.din(w_dff_A_tQnXJQLk8_1),.clk(gclk));
	jdff dff_A_KBaZDOHP1_1(.dout(w_dff_A_O55q3XcK7_0),.din(w_dff_A_KBaZDOHP1_1),.clk(gclk));
	jdff dff_A_O55q3XcK7_0(.dout(w_dff_A_w1WlN4AI1_0),.din(w_dff_A_O55q3XcK7_0),.clk(gclk));
	jdff dff_A_w1WlN4AI1_0(.dout(w_dff_A_d39dEwf79_0),.din(w_dff_A_w1WlN4AI1_0),.clk(gclk));
	jdff dff_A_d39dEwf79_0(.dout(w_dff_A_iRFpg1AX9_0),.din(w_dff_A_d39dEwf79_0),.clk(gclk));
	jdff dff_A_iRFpg1AX9_0(.dout(w_dff_A_gE5dWq0S1_0),.din(w_dff_A_iRFpg1AX9_0),.clk(gclk));
	jdff dff_A_gE5dWq0S1_0(.dout(w_dff_A_ZsBMiGr98_0),.din(w_dff_A_gE5dWq0S1_0),.clk(gclk));
	jdff dff_A_ZsBMiGr98_0(.dout(w_dff_A_nwvxDHjX7_0),.din(w_dff_A_ZsBMiGr98_0),.clk(gclk));
	jdff dff_A_nwvxDHjX7_0(.dout(w_dff_A_aO9mcUsK9_0),.din(w_dff_A_nwvxDHjX7_0),.clk(gclk));
	jdff dff_A_aO9mcUsK9_0(.dout(w_dff_A_n17gOZIr2_0),.din(w_dff_A_aO9mcUsK9_0),.clk(gclk));
	jdff dff_A_n17gOZIr2_0(.dout(w_dff_A_YFNalbol9_0),.din(w_dff_A_n17gOZIr2_0),.clk(gclk));
	jdff dff_A_YFNalbol9_0(.dout(w_dff_A_YG0sqLTW2_0),.din(w_dff_A_YFNalbol9_0),.clk(gclk));
	jdff dff_A_YG0sqLTW2_0(.dout(w_dff_A_YpF1Lz788_0),.din(w_dff_A_YG0sqLTW2_0),.clk(gclk));
	jdff dff_A_YpF1Lz788_0(.dout(w_dff_A_JAwS5IiX2_0),.din(w_dff_A_YpF1Lz788_0),.clk(gclk));
	jdff dff_A_JAwS5IiX2_0(.dout(w_dff_A_CXTW5kwL9_0),.din(w_dff_A_JAwS5IiX2_0),.clk(gclk));
	jdff dff_A_CXTW5kwL9_0(.dout(w_dff_A_BH73yURA2_0),.din(w_dff_A_CXTW5kwL9_0),.clk(gclk));
	jdff dff_A_BH73yURA2_0(.dout(w_dff_A_vk5O05BE9_0),.din(w_dff_A_BH73yURA2_0),.clk(gclk));
	jdff dff_A_vk5O05BE9_0(.dout(w_dff_A_Sdq6fSR90_0),.din(w_dff_A_vk5O05BE9_0),.clk(gclk));
	jdff dff_A_Sdq6fSR90_0(.dout(w_dff_A_uBjr6PJN0_0),.din(w_dff_A_Sdq6fSR90_0),.clk(gclk));
	jdff dff_A_uBjr6PJN0_0(.dout(w_dff_A_oSINyjGd2_0),.din(w_dff_A_uBjr6PJN0_0),.clk(gclk));
	jdff dff_A_oSINyjGd2_0(.dout(w_dff_A_scs8vgnV1_0),.din(w_dff_A_oSINyjGd2_0),.clk(gclk));
	jdff dff_A_scs8vgnV1_0(.dout(w_dff_A_DVBqqvXa1_0),.din(w_dff_A_scs8vgnV1_0),.clk(gclk));
	jdff dff_A_DVBqqvXa1_0(.dout(w_dff_A_ZhkqUzOK5_0),.din(w_dff_A_DVBqqvXa1_0),.clk(gclk));
	jdff dff_A_ZhkqUzOK5_0(.dout(w_dff_A_fiDNaUrJ2_0),.din(w_dff_A_ZhkqUzOK5_0),.clk(gclk));
	jdff dff_A_fiDNaUrJ2_0(.dout(w_dff_A_wAivC2bE7_0),.din(w_dff_A_fiDNaUrJ2_0),.clk(gclk));
	jdff dff_A_wAivC2bE7_0(.dout(w_dff_A_9d6KjivI6_0),.din(w_dff_A_wAivC2bE7_0),.clk(gclk));
	jdff dff_A_9d6KjivI6_0(.dout(w_dff_A_qDCk6K6o9_0),.din(w_dff_A_9d6KjivI6_0),.clk(gclk));
	jdff dff_A_qDCk6K6o9_0(.dout(w_dff_A_sQ8TdCZo1_0),.din(w_dff_A_qDCk6K6o9_0),.clk(gclk));
	jdff dff_A_sQ8TdCZo1_0(.dout(G144),.din(w_dff_A_sQ8TdCZo1_0),.clk(gclk));
	jdff dff_A_4s92yFbR3_1(.dout(w_dff_A_iaNi7GL72_0),.din(w_dff_A_4s92yFbR3_1),.clk(gclk));
	jdff dff_A_iaNi7GL72_0(.dout(w_dff_A_jeeHocm09_0),.din(w_dff_A_iaNi7GL72_0),.clk(gclk));
	jdff dff_A_jeeHocm09_0(.dout(w_dff_A_iEpSj3AB0_0),.din(w_dff_A_jeeHocm09_0),.clk(gclk));
	jdff dff_A_iEpSj3AB0_0(.dout(w_dff_A_wQ5QBoUP2_0),.din(w_dff_A_iEpSj3AB0_0),.clk(gclk));
	jdff dff_A_wQ5QBoUP2_0(.dout(w_dff_A_ACyjzPfS1_0),.din(w_dff_A_wQ5QBoUP2_0),.clk(gclk));
	jdff dff_A_ACyjzPfS1_0(.dout(w_dff_A_Du8rORXL4_0),.din(w_dff_A_ACyjzPfS1_0),.clk(gclk));
	jdff dff_A_Du8rORXL4_0(.dout(w_dff_A_HCIvCoYX1_0),.din(w_dff_A_Du8rORXL4_0),.clk(gclk));
	jdff dff_A_HCIvCoYX1_0(.dout(w_dff_A_Fs8KLIcd3_0),.din(w_dff_A_HCIvCoYX1_0),.clk(gclk));
	jdff dff_A_Fs8KLIcd3_0(.dout(w_dff_A_Evrcr3Cn2_0),.din(w_dff_A_Fs8KLIcd3_0),.clk(gclk));
	jdff dff_A_Evrcr3Cn2_0(.dout(w_dff_A_SYf1JhFY3_0),.din(w_dff_A_Evrcr3Cn2_0),.clk(gclk));
	jdff dff_A_SYf1JhFY3_0(.dout(w_dff_A_4dNXf1YS2_0),.din(w_dff_A_SYf1JhFY3_0),.clk(gclk));
	jdff dff_A_4dNXf1YS2_0(.dout(w_dff_A_l9JSuQe12_0),.din(w_dff_A_4dNXf1YS2_0),.clk(gclk));
	jdff dff_A_l9JSuQe12_0(.dout(w_dff_A_V4cbptXz5_0),.din(w_dff_A_l9JSuQe12_0),.clk(gclk));
	jdff dff_A_V4cbptXz5_0(.dout(w_dff_A_heYE8yQO8_0),.din(w_dff_A_V4cbptXz5_0),.clk(gclk));
	jdff dff_A_heYE8yQO8_0(.dout(w_dff_A_owQF4Orj7_0),.din(w_dff_A_heYE8yQO8_0),.clk(gclk));
	jdff dff_A_owQF4Orj7_0(.dout(w_dff_A_gmbncTAf6_0),.din(w_dff_A_owQF4Orj7_0),.clk(gclk));
	jdff dff_A_gmbncTAf6_0(.dout(w_dff_A_p0EEFjqn4_0),.din(w_dff_A_gmbncTAf6_0),.clk(gclk));
	jdff dff_A_p0EEFjqn4_0(.dout(w_dff_A_c79ofdHL9_0),.din(w_dff_A_p0EEFjqn4_0),.clk(gclk));
	jdff dff_A_c79ofdHL9_0(.dout(w_dff_A_BsmwsAGq7_0),.din(w_dff_A_c79ofdHL9_0),.clk(gclk));
	jdff dff_A_BsmwsAGq7_0(.dout(w_dff_A_81mxqh3e1_0),.din(w_dff_A_BsmwsAGq7_0),.clk(gclk));
	jdff dff_A_81mxqh3e1_0(.dout(w_dff_A_f28vrxeI8_0),.din(w_dff_A_81mxqh3e1_0),.clk(gclk));
	jdff dff_A_f28vrxeI8_0(.dout(w_dff_A_FMJuHK8E2_0),.din(w_dff_A_f28vrxeI8_0),.clk(gclk));
	jdff dff_A_FMJuHK8E2_0(.dout(w_dff_A_aSCv58Ye4_0),.din(w_dff_A_FMJuHK8E2_0),.clk(gclk));
	jdff dff_A_aSCv58Ye4_0(.dout(w_dff_A_Vfi4Qppj4_0),.din(w_dff_A_aSCv58Ye4_0),.clk(gclk));
	jdff dff_A_Vfi4Qppj4_0(.dout(w_dff_A_t1JBGe2o0_0),.din(w_dff_A_Vfi4Qppj4_0),.clk(gclk));
	jdff dff_A_t1JBGe2o0_0(.dout(w_dff_A_QtudEZHd5_0),.din(w_dff_A_t1JBGe2o0_0),.clk(gclk));
	jdff dff_A_QtudEZHd5_0(.dout(w_dff_A_1lI57vtL8_0),.din(w_dff_A_QtudEZHd5_0),.clk(gclk));
	jdff dff_A_1lI57vtL8_0(.dout(G298),.din(w_dff_A_1lI57vtL8_0),.clk(gclk));
	jdff dff_A_nC4ucAtV8_1(.dout(w_dff_A_yj1mftS23_0),.din(w_dff_A_nC4ucAtV8_1),.clk(gclk));
	jdff dff_A_yj1mftS23_0(.dout(w_dff_A_C808ufh08_0),.din(w_dff_A_yj1mftS23_0),.clk(gclk));
	jdff dff_A_C808ufh08_0(.dout(w_dff_A_Sk05vxiE6_0),.din(w_dff_A_C808ufh08_0),.clk(gclk));
	jdff dff_A_Sk05vxiE6_0(.dout(w_dff_A_tT5h57D99_0),.din(w_dff_A_Sk05vxiE6_0),.clk(gclk));
	jdff dff_A_tT5h57D99_0(.dout(w_dff_A_Ut2HIQPJ1_0),.din(w_dff_A_tT5h57D99_0),.clk(gclk));
	jdff dff_A_Ut2HIQPJ1_0(.dout(w_dff_A_kBa65aPK7_0),.din(w_dff_A_Ut2HIQPJ1_0),.clk(gclk));
	jdff dff_A_kBa65aPK7_0(.dout(w_dff_A_Lda4FzC81_0),.din(w_dff_A_kBa65aPK7_0),.clk(gclk));
	jdff dff_A_Lda4FzC81_0(.dout(w_dff_A_0KLFGTHZ8_0),.din(w_dff_A_Lda4FzC81_0),.clk(gclk));
	jdff dff_A_0KLFGTHZ8_0(.dout(w_dff_A_BD20nFcH8_0),.din(w_dff_A_0KLFGTHZ8_0),.clk(gclk));
	jdff dff_A_BD20nFcH8_0(.dout(w_dff_A_TixNXhdh6_0),.din(w_dff_A_BD20nFcH8_0),.clk(gclk));
	jdff dff_A_TixNXhdh6_0(.dout(w_dff_A_9C3qfpFN7_0),.din(w_dff_A_TixNXhdh6_0),.clk(gclk));
	jdff dff_A_9C3qfpFN7_0(.dout(w_dff_A_QLk8oJKB1_0),.din(w_dff_A_9C3qfpFN7_0),.clk(gclk));
	jdff dff_A_QLk8oJKB1_0(.dout(w_dff_A_OBdxKKiw8_0),.din(w_dff_A_QLk8oJKB1_0),.clk(gclk));
	jdff dff_A_OBdxKKiw8_0(.dout(w_dff_A_xBXelP438_0),.din(w_dff_A_OBdxKKiw8_0),.clk(gclk));
	jdff dff_A_xBXelP438_0(.dout(w_dff_A_glkSImVQ6_0),.din(w_dff_A_xBXelP438_0),.clk(gclk));
	jdff dff_A_glkSImVQ6_0(.dout(w_dff_A_qFRBqL0F8_0),.din(w_dff_A_glkSImVQ6_0),.clk(gclk));
	jdff dff_A_qFRBqL0F8_0(.dout(w_dff_A_kDerP2dF3_0),.din(w_dff_A_qFRBqL0F8_0),.clk(gclk));
	jdff dff_A_kDerP2dF3_0(.dout(w_dff_A_7vWTjxYE3_0),.din(w_dff_A_kDerP2dF3_0),.clk(gclk));
	jdff dff_A_7vWTjxYE3_0(.dout(w_dff_A_NF90MJWc2_0),.din(w_dff_A_7vWTjxYE3_0),.clk(gclk));
	jdff dff_A_NF90MJWc2_0(.dout(w_dff_A_wLf5JT0f0_0),.din(w_dff_A_NF90MJWc2_0),.clk(gclk));
	jdff dff_A_wLf5JT0f0_0(.dout(w_dff_A_czaFwE1w0_0),.din(w_dff_A_wLf5JT0f0_0),.clk(gclk));
	jdff dff_A_czaFwE1w0_0(.dout(w_dff_A_VAl9tb9u1_0),.din(w_dff_A_czaFwE1w0_0),.clk(gclk));
	jdff dff_A_VAl9tb9u1_0(.dout(w_dff_A_45WW4B4c5_0),.din(w_dff_A_VAl9tb9u1_0),.clk(gclk));
	jdff dff_A_45WW4B4c5_0(.dout(w_dff_A_fwYGUm3D2_0),.din(w_dff_A_45WW4B4c5_0),.clk(gclk));
	jdff dff_A_fwYGUm3D2_0(.dout(w_dff_A_iiHRlj2M3_0),.din(w_dff_A_fwYGUm3D2_0),.clk(gclk));
	jdff dff_A_iiHRlj2M3_0(.dout(w_dff_A_w7a0VZHC3_0),.din(w_dff_A_iiHRlj2M3_0),.clk(gclk));
	jdff dff_A_w7a0VZHC3_0(.dout(w_dff_A_5mOEKxsL9_0),.din(w_dff_A_w7a0VZHC3_0),.clk(gclk));
	jdff dff_A_5mOEKxsL9_0(.dout(G973),.din(w_dff_A_5mOEKxsL9_0),.clk(gclk));
	jdff dff_A_ep1FTgkM5_1(.dout(w_dff_A_sG5fiiKG3_0),.din(w_dff_A_ep1FTgkM5_1),.clk(gclk));
	jdff dff_A_sG5fiiKG3_0(.dout(w_dff_A_8mLk11gH5_0),.din(w_dff_A_sG5fiiKG3_0),.clk(gclk));
	jdff dff_A_8mLk11gH5_0(.dout(w_dff_A_gEGTZFFE5_0),.din(w_dff_A_8mLk11gH5_0),.clk(gclk));
	jdff dff_A_gEGTZFFE5_0(.dout(w_dff_A_Ex4zNjTg9_0),.din(w_dff_A_gEGTZFFE5_0),.clk(gclk));
	jdff dff_A_Ex4zNjTg9_0(.dout(w_dff_A_50WgwozR5_0),.din(w_dff_A_Ex4zNjTg9_0),.clk(gclk));
	jdff dff_A_50WgwozR5_0(.dout(w_dff_A_v9fQoIi61_0),.din(w_dff_A_50WgwozR5_0),.clk(gclk));
	jdff dff_A_v9fQoIi61_0(.dout(w_dff_A_jMuvNS7h7_0),.din(w_dff_A_v9fQoIi61_0),.clk(gclk));
	jdff dff_A_jMuvNS7h7_0(.dout(w_dff_A_8RCay6Fk4_0),.din(w_dff_A_jMuvNS7h7_0),.clk(gclk));
	jdff dff_A_8RCay6Fk4_0(.dout(w_dff_A_pudPBWr98_0),.din(w_dff_A_8RCay6Fk4_0),.clk(gclk));
	jdff dff_A_pudPBWr98_0(.dout(w_dff_A_8jl9caJj3_0),.din(w_dff_A_pudPBWr98_0),.clk(gclk));
	jdff dff_A_8jl9caJj3_0(.dout(w_dff_A_KDPIP7dV9_0),.din(w_dff_A_8jl9caJj3_0),.clk(gclk));
	jdff dff_A_KDPIP7dV9_0(.dout(w_dff_A_8I1KSjuQ0_0),.din(w_dff_A_KDPIP7dV9_0),.clk(gclk));
	jdff dff_A_8I1KSjuQ0_0(.dout(w_dff_A_tW4BgmE30_0),.din(w_dff_A_8I1KSjuQ0_0),.clk(gclk));
	jdff dff_A_tW4BgmE30_0(.dout(w_dff_A_CEMWlLdu1_0),.din(w_dff_A_tW4BgmE30_0),.clk(gclk));
	jdff dff_A_CEMWlLdu1_0(.dout(w_dff_A_A1QkQi018_0),.din(w_dff_A_CEMWlLdu1_0),.clk(gclk));
	jdff dff_A_A1QkQi018_0(.dout(w_dff_A_FqUWZ8wB4_0),.din(w_dff_A_A1QkQi018_0),.clk(gclk));
	jdff dff_A_FqUWZ8wB4_0(.dout(w_dff_A_wmIzeUMo4_0),.din(w_dff_A_FqUWZ8wB4_0),.clk(gclk));
	jdff dff_A_wmIzeUMo4_0(.dout(w_dff_A_Ai5N5ciN2_0),.din(w_dff_A_wmIzeUMo4_0),.clk(gclk));
	jdff dff_A_Ai5N5ciN2_0(.dout(w_dff_A_xqazbTIo7_0),.din(w_dff_A_Ai5N5ciN2_0),.clk(gclk));
	jdff dff_A_xqazbTIo7_0(.dout(w_dff_A_nswAEyaX7_0),.din(w_dff_A_xqazbTIo7_0),.clk(gclk));
	jdff dff_A_nswAEyaX7_0(.dout(w_dff_A_zlEdpTdk9_0),.din(w_dff_A_nswAEyaX7_0),.clk(gclk));
	jdff dff_A_zlEdpTdk9_0(.dout(w_dff_A_M3qfnjbV0_0),.din(w_dff_A_zlEdpTdk9_0),.clk(gclk));
	jdff dff_A_M3qfnjbV0_0(.dout(w_dff_A_wzzMYBWz1_0),.din(w_dff_A_M3qfnjbV0_0),.clk(gclk));
	jdff dff_A_wzzMYBWz1_0(.dout(w_dff_A_Ig5Xr1RJ6_0),.din(w_dff_A_wzzMYBWz1_0),.clk(gclk));
	jdff dff_A_Ig5Xr1RJ6_0(.dout(w_dff_A_JbWVN4om8_0),.din(w_dff_A_Ig5Xr1RJ6_0),.clk(gclk));
	jdff dff_A_JbWVN4om8_0(.dout(w_dff_A_shGbW1mx5_0),.din(w_dff_A_JbWVN4om8_0),.clk(gclk));
	jdff dff_A_shGbW1mx5_0(.dout(G594),.din(w_dff_A_shGbW1mx5_0),.clk(gclk));
	jdff dff_A_vVTXHN0Y8_1(.dout(w_dff_A_T7qej8Wr6_0),.din(w_dff_A_vVTXHN0Y8_1),.clk(gclk));
	jdff dff_A_T7qej8Wr6_0(.dout(w_dff_A_00lGSYGk9_0),.din(w_dff_A_T7qej8Wr6_0),.clk(gclk));
	jdff dff_A_00lGSYGk9_0(.dout(w_dff_A_o3xTl1vp0_0),.din(w_dff_A_00lGSYGk9_0),.clk(gclk));
	jdff dff_A_o3xTl1vp0_0(.dout(w_dff_A_61azdeHC7_0),.din(w_dff_A_o3xTl1vp0_0),.clk(gclk));
	jdff dff_A_61azdeHC7_0(.dout(w_dff_A_7lUkVmbZ0_0),.din(w_dff_A_61azdeHC7_0),.clk(gclk));
	jdff dff_A_7lUkVmbZ0_0(.dout(w_dff_A_NqiOp5g87_0),.din(w_dff_A_7lUkVmbZ0_0),.clk(gclk));
	jdff dff_A_NqiOp5g87_0(.dout(w_dff_A_PFBfGFmI6_0),.din(w_dff_A_NqiOp5g87_0),.clk(gclk));
	jdff dff_A_PFBfGFmI6_0(.dout(w_dff_A_tgKKQzvn0_0),.din(w_dff_A_PFBfGFmI6_0),.clk(gclk));
	jdff dff_A_tgKKQzvn0_0(.dout(w_dff_A_HsB2ReTN3_0),.din(w_dff_A_tgKKQzvn0_0),.clk(gclk));
	jdff dff_A_HsB2ReTN3_0(.dout(w_dff_A_amEKxW6y8_0),.din(w_dff_A_HsB2ReTN3_0),.clk(gclk));
	jdff dff_A_amEKxW6y8_0(.dout(w_dff_A_cbTfVXzF2_0),.din(w_dff_A_amEKxW6y8_0),.clk(gclk));
	jdff dff_A_cbTfVXzF2_0(.dout(w_dff_A_AFQXmTym4_0),.din(w_dff_A_cbTfVXzF2_0),.clk(gclk));
	jdff dff_A_AFQXmTym4_0(.dout(w_dff_A_Y2LEw09O5_0),.din(w_dff_A_AFQXmTym4_0),.clk(gclk));
	jdff dff_A_Y2LEw09O5_0(.dout(w_dff_A_qXAZ85gj6_0),.din(w_dff_A_Y2LEw09O5_0),.clk(gclk));
	jdff dff_A_qXAZ85gj6_0(.dout(w_dff_A_jHVNiXGu0_0),.din(w_dff_A_qXAZ85gj6_0),.clk(gclk));
	jdff dff_A_jHVNiXGu0_0(.dout(w_dff_A_Ah5OEZOB8_0),.din(w_dff_A_jHVNiXGu0_0),.clk(gclk));
	jdff dff_A_Ah5OEZOB8_0(.dout(w_dff_A_Gr2rXtPe2_0),.din(w_dff_A_Ah5OEZOB8_0),.clk(gclk));
	jdff dff_A_Gr2rXtPe2_0(.dout(w_dff_A_2ZorcICg0_0),.din(w_dff_A_Gr2rXtPe2_0),.clk(gclk));
	jdff dff_A_2ZorcICg0_0(.dout(w_dff_A_Ec6mxR3J3_0),.din(w_dff_A_2ZorcICg0_0),.clk(gclk));
	jdff dff_A_Ec6mxR3J3_0(.dout(w_dff_A_NfA4Wpet6_0),.din(w_dff_A_Ec6mxR3J3_0),.clk(gclk));
	jdff dff_A_NfA4Wpet6_0(.dout(w_dff_A_2WIERxJT2_0),.din(w_dff_A_NfA4Wpet6_0),.clk(gclk));
	jdff dff_A_2WIERxJT2_0(.dout(w_dff_A_prNjylbA6_0),.din(w_dff_A_2WIERxJT2_0),.clk(gclk));
	jdff dff_A_prNjylbA6_0(.dout(w_dff_A_gszMv0ZJ1_0),.din(w_dff_A_prNjylbA6_0),.clk(gclk));
	jdff dff_A_gszMv0ZJ1_0(.dout(w_dff_A_c2GUCEwU2_0),.din(w_dff_A_gszMv0ZJ1_0),.clk(gclk));
	jdff dff_A_c2GUCEwU2_0(.dout(w_dff_A_QPI9oVNu0_0),.din(w_dff_A_c2GUCEwU2_0),.clk(gclk));
	jdff dff_A_QPI9oVNu0_0(.dout(w_dff_A_ayQKAA0n6_0),.din(w_dff_A_QPI9oVNu0_0),.clk(gclk));
	jdff dff_A_ayQKAA0n6_0(.dout(G599),.din(w_dff_A_ayQKAA0n6_0),.clk(gclk));
	jdff dff_A_3AcVMzYK5_1(.dout(w_dff_A_0j5bfoEz0_0),.din(w_dff_A_3AcVMzYK5_1),.clk(gclk));
	jdff dff_A_0j5bfoEz0_0(.dout(w_dff_A_5msFLLaZ2_0),.din(w_dff_A_0j5bfoEz0_0),.clk(gclk));
	jdff dff_A_5msFLLaZ2_0(.dout(w_dff_A_HQ7EyUs90_0),.din(w_dff_A_5msFLLaZ2_0),.clk(gclk));
	jdff dff_A_HQ7EyUs90_0(.dout(w_dff_A_tVzeAobB4_0),.din(w_dff_A_HQ7EyUs90_0),.clk(gclk));
	jdff dff_A_tVzeAobB4_0(.dout(w_dff_A_46BXZkeF5_0),.din(w_dff_A_tVzeAobB4_0),.clk(gclk));
	jdff dff_A_46BXZkeF5_0(.dout(w_dff_A_pKa5FU5T1_0),.din(w_dff_A_46BXZkeF5_0),.clk(gclk));
	jdff dff_A_pKa5FU5T1_0(.dout(w_dff_A_ktA3ajId1_0),.din(w_dff_A_pKa5FU5T1_0),.clk(gclk));
	jdff dff_A_ktA3ajId1_0(.dout(w_dff_A_sVJ62UAT1_0),.din(w_dff_A_ktA3ajId1_0),.clk(gclk));
	jdff dff_A_sVJ62UAT1_0(.dout(w_dff_A_6dTh5qJ81_0),.din(w_dff_A_sVJ62UAT1_0),.clk(gclk));
	jdff dff_A_6dTh5qJ81_0(.dout(w_dff_A_tPGzkkzL1_0),.din(w_dff_A_6dTh5qJ81_0),.clk(gclk));
	jdff dff_A_tPGzkkzL1_0(.dout(w_dff_A_IA5TMtTJ8_0),.din(w_dff_A_tPGzkkzL1_0),.clk(gclk));
	jdff dff_A_IA5TMtTJ8_0(.dout(w_dff_A_pOyCgSsE2_0),.din(w_dff_A_IA5TMtTJ8_0),.clk(gclk));
	jdff dff_A_pOyCgSsE2_0(.dout(w_dff_A_4hUIvpAP3_0),.din(w_dff_A_pOyCgSsE2_0),.clk(gclk));
	jdff dff_A_4hUIvpAP3_0(.dout(w_dff_A_0O0QB71m9_0),.din(w_dff_A_4hUIvpAP3_0),.clk(gclk));
	jdff dff_A_0O0QB71m9_0(.dout(w_dff_A_vn66pJ4c5_0),.din(w_dff_A_0O0QB71m9_0),.clk(gclk));
	jdff dff_A_vn66pJ4c5_0(.dout(w_dff_A_xHGnSItg4_0),.din(w_dff_A_vn66pJ4c5_0),.clk(gclk));
	jdff dff_A_xHGnSItg4_0(.dout(w_dff_A_IqmN4zcM3_0),.din(w_dff_A_xHGnSItg4_0),.clk(gclk));
	jdff dff_A_IqmN4zcM3_0(.dout(w_dff_A_pUTUQbj52_0),.din(w_dff_A_IqmN4zcM3_0),.clk(gclk));
	jdff dff_A_pUTUQbj52_0(.dout(w_dff_A_WeKdg6F09_0),.din(w_dff_A_pUTUQbj52_0),.clk(gclk));
	jdff dff_A_WeKdg6F09_0(.dout(w_dff_A_EI9YwJ1u6_0),.din(w_dff_A_WeKdg6F09_0),.clk(gclk));
	jdff dff_A_EI9YwJ1u6_0(.dout(w_dff_A_bo3gmzBx1_0),.din(w_dff_A_EI9YwJ1u6_0),.clk(gclk));
	jdff dff_A_bo3gmzBx1_0(.dout(w_dff_A_u698IDfd9_0),.din(w_dff_A_bo3gmzBx1_0),.clk(gclk));
	jdff dff_A_u698IDfd9_0(.dout(w_dff_A_KZA8eMev8_0),.din(w_dff_A_u698IDfd9_0),.clk(gclk));
	jdff dff_A_KZA8eMev8_0(.dout(w_dff_A_Q0hFrD3t4_0),.din(w_dff_A_KZA8eMev8_0),.clk(gclk));
	jdff dff_A_Q0hFrD3t4_0(.dout(w_dff_A_DBz8CL4e2_0),.din(w_dff_A_Q0hFrD3t4_0),.clk(gclk));
	jdff dff_A_DBz8CL4e2_0(.dout(w_dff_A_ey8ymUK49_0),.din(w_dff_A_DBz8CL4e2_0),.clk(gclk));
	jdff dff_A_ey8ymUK49_0(.dout(G600),.din(w_dff_A_ey8ymUK49_0),.clk(gclk));
	jdff dff_A_vJT8vmhz2_1(.dout(w_dff_A_npcMJPQN3_0),.din(w_dff_A_vJT8vmhz2_1),.clk(gclk));
	jdff dff_A_npcMJPQN3_0(.dout(w_dff_A_M1pwvoLi1_0),.din(w_dff_A_npcMJPQN3_0),.clk(gclk));
	jdff dff_A_M1pwvoLi1_0(.dout(w_dff_A_kkReI27O4_0),.din(w_dff_A_M1pwvoLi1_0),.clk(gclk));
	jdff dff_A_kkReI27O4_0(.dout(w_dff_A_Nv32qHlP3_0),.din(w_dff_A_kkReI27O4_0),.clk(gclk));
	jdff dff_A_Nv32qHlP3_0(.dout(w_dff_A_Q3zV6DgZ0_0),.din(w_dff_A_Nv32qHlP3_0),.clk(gclk));
	jdff dff_A_Q3zV6DgZ0_0(.dout(w_dff_A_PS7bCVib4_0),.din(w_dff_A_Q3zV6DgZ0_0),.clk(gclk));
	jdff dff_A_PS7bCVib4_0(.dout(w_dff_A_pHzQrpJB6_0),.din(w_dff_A_PS7bCVib4_0),.clk(gclk));
	jdff dff_A_pHzQrpJB6_0(.dout(w_dff_A_BIzqZff30_0),.din(w_dff_A_pHzQrpJB6_0),.clk(gclk));
	jdff dff_A_BIzqZff30_0(.dout(w_dff_A_xTc5dEBV1_0),.din(w_dff_A_BIzqZff30_0),.clk(gclk));
	jdff dff_A_xTc5dEBV1_0(.dout(w_dff_A_fdQWXOgn6_0),.din(w_dff_A_xTc5dEBV1_0),.clk(gclk));
	jdff dff_A_fdQWXOgn6_0(.dout(w_dff_A_ZuCcz3uN6_0),.din(w_dff_A_fdQWXOgn6_0),.clk(gclk));
	jdff dff_A_ZuCcz3uN6_0(.dout(w_dff_A_CacUs3Gb8_0),.din(w_dff_A_ZuCcz3uN6_0),.clk(gclk));
	jdff dff_A_CacUs3Gb8_0(.dout(w_dff_A_uvgeC17M7_0),.din(w_dff_A_CacUs3Gb8_0),.clk(gclk));
	jdff dff_A_uvgeC17M7_0(.dout(w_dff_A_XhEB0sUY4_0),.din(w_dff_A_uvgeC17M7_0),.clk(gclk));
	jdff dff_A_XhEB0sUY4_0(.dout(w_dff_A_ZLfHUCVs8_0),.din(w_dff_A_XhEB0sUY4_0),.clk(gclk));
	jdff dff_A_ZLfHUCVs8_0(.dout(w_dff_A_H4CR3XYo6_0),.din(w_dff_A_ZLfHUCVs8_0),.clk(gclk));
	jdff dff_A_H4CR3XYo6_0(.dout(w_dff_A_1LnKWEV83_0),.din(w_dff_A_H4CR3XYo6_0),.clk(gclk));
	jdff dff_A_1LnKWEV83_0(.dout(w_dff_A_PzdUgxQs7_0),.din(w_dff_A_1LnKWEV83_0),.clk(gclk));
	jdff dff_A_PzdUgxQs7_0(.dout(w_dff_A_UsPgI78c7_0),.din(w_dff_A_PzdUgxQs7_0),.clk(gclk));
	jdff dff_A_UsPgI78c7_0(.dout(w_dff_A_Dj1o5tiA7_0),.din(w_dff_A_UsPgI78c7_0),.clk(gclk));
	jdff dff_A_Dj1o5tiA7_0(.dout(w_dff_A_dWu8hV7i1_0),.din(w_dff_A_Dj1o5tiA7_0),.clk(gclk));
	jdff dff_A_dWu8hV7i1_0(.dout(w_dff_A_A3g2c3Ur5_0),.din(w_dff_A_dWu8hV7i1_0),.clk(gclk));
	jdff dff_A_A3g2c3Ur5_0(.dout(w_dff_A_hHr3EZtt5_0),.din(w_dff_A_A3g2c3Ur5_0),.clk(gclk));
	jdff dff_A_hHr3EZtt5_0(.dout(w_dff_A_k9SaaSDn3_0),.din(w_dff_A_hHr3EZtt5_0),.clk(gclk));
	jdff dff_A_k9SaaSDn3_0(.dout(w_dff_A_qMPiwV2W2_0),.din(w_dff_A_k9SaaSDn3_0),.clk(gclk));
	jdff dff_A_qMPiwV2W2_0(.dout(w_dff_A_DW3x1vES3_0),.din(w_dff_A_qMPiwV2W2_0),.clk(gclk));
	jdff dff_A_DW3x1vES3_0(.dout(G601),.din(w_dff_A_DW3x1vES3_0),.clk(gclk));
	jdff dff_A_izx8mPSq2_1(.dout(w_dff_A_LX1UfqQN8_0),.din(w_dff_A_izx8mPSq2_1),.clk(gclk));
	jdff dff_A_LX1UfqQN8_0(.dout(w_dff_A_nDs8iTmV8_0),.din(w_dff_A_LX1UfqQN8_0),.clk(gclk));
	jdff dff_A_nDs8iTmV8_0(.dout(w_dff_A_Xdeug0Jp0_0),.din(w_dff_A_nDs8iTmV8_0),.clk(gclk));
	jdff dff_A_Xdeug0Jp0_0(.dout(w_dff_A_BtBvgrzV4_0),.din(w_dff_A_Xdeug0Jp0_0),.clk(gclk));
	jdff dff_A_BtBvgrzV4_0(.dout(w_dff_A_QMA8XHCb9_0),.din(w_dff_A_BtBvgrzV4_0),.clk(gclk));
	jdff dff_A_QMA8XHCb9_0(.dout(w_dff_A_iWmqhsGu4_0),.din(w_dff_A_QMA8XHCb9_0),.clk(gclk));
	jdff dff_A_iWmqhsGu4_0(.dout(w_dff_A_GaADXKXM5_0),.din(w_dff_A_iWmqhsGu4_0),.clk(gclk));
	jdff dff_A_GaADXKXM5_0(.dout(w_dff_A_aiYxBukP0_0),.din(w_dff_A_GaADXKXM5_0),.clk(gclk));
	jdff dff_A_aiYxBukP0_0(.dout(w_dff_A_cvbiK8eE6_0),.din(w_dff_A_aiYxBukP0_0),.clk(gclk));
	jdff dff_A_cvbiK8eE6_0(.dout(w_dff_A_7QoaRM451_0),.din(w_dff_A_cvbiK8eE6_0),.clk(gclk));
	jdff dff_A_7QoaRM451_0(.dout(w_dff_A_WVOGs99W8_0),.din(w_dff_A_7QoaRM451_0),.clk(gclk));
	jdff dff_A_WVOGs99W8_0(.dout(w_dff_A_Ar65qGqw4_0),.din(w_dff_A_WVOGs99W8_0),.clk(gclk));
	jdff dff_A_Ar65qGqw4_0(.dout(w_dff_A_C6Wsa84o6_0),.din(w_dff_A_Ar65qGqw4_0),.clk(gclk));
	jdff dff_A_C6Wsa84o6_0(.dout(w_dff_A_7FZ4qnfn4_0),.din(w_dff_A_C6Wsa84o6_0),.clk(gclk));
	jdff dff_A_7FZ4qnfn4_0(.dout(w_dff_A_WomVql2A1_0),.din(w_dff_A_7FZ4qnfn4_0),.clk(gclk));
	jdff dff_A_WomVql2A1_0(.dout(w_dff_A_XWfPtfUX1_0),.din(w_dff_A_WomVql2A1_0),.clk(gclk));
	jdff dff_A_XWfPtfUX1_0(.dout(w_dff_A_wNg1G72Z6_0),.din(w_dff_A_XWfPtfUX1_0),.clk(gclk));
	jdff dff_A_wNg1G72Z6_0(.dout(w_dff_A_zBoW7lHC5_0),.din(w_dff_A_wNg1G72Z6_0),.clk(gclk));
	jdff dff_A_zBoW7lHC5_0(.dout(w_dff_A_El2akflr1_0),.din(w_dff_A_zBoW7lHC5_0),.clk(gclk));
	jdff dff_A_El2akflr1_0(.dout(w_dff_A_PYo80HcF8_0),.din(w_dff_A_El2akflr1_0),.clk(gclk));
	jdff dff_A_PYo80HcF8_0(.dout(w_dff_A_pF6sYABj2_0),.din(w_dff_A_PYo80HcF8_0),.clk(gclk));
	jdff dff_A_pF6sYABj2_0(.dout(w_dff_A_LO29noL97_0),.din(w_dff_A_pF6sYABj2_0),.clk(gclk));
	jdff dff_A_LO29noL97_0(.dout(w_dff_A_6vS7HMc92_0),.din(w_dff_A_LO29noL97_0),.clk(gclk));
	jdff dff_A_6vS7HMc92_0(.dout(w_dff_A_ZncOYlGO8_0),.din(w_dff_A_6vS7HMc92_0),.clk(gclk));
	jdff dff_A_ZncOYlGO8_0(.dout(w_dff_A_cYqjTFUI8_0),.din(w_dff_A_ZncOYlGO8_0),.clk(gclk));
	jdff dff_A_cYqjTFUI8_0(.dout(w_dff_A_SpSsRYeB7_0),.din(w_dff_A_cYqjTFUI8_0),.clk(gclk));
	jdff dff_A_SpSsRYeB7_0(.dout(G602),.din(w_dff_A_SpSsRYeB7_0),.clk(gclk));
	jdff dff_A_RRZ9uML84_1(.dout(w_dff_A_6EptrX162_0),.din(w_dff_A_RRZ9uML84_1),.clk(gclk));
	jdff dff_A_6EptrX162_0(.dout(w_dff_A_G1Od5GP96_0),.din(w_dff_A_6EptrX162_0),.clk(gclk));
	jdff dff_A_G1Od5GP96_0(.dout(w_dff_A_ww2wX3W68_0),.din(w_dff_A_G1Od5GP96_0),.clk(gclk));
	jdff dff_A_ww2wX3W68_0(.dout(w_dff_A_eUpFYx1Q4_0),.din(w_dff_A_ww2wX3W68_0),.clk(gclk));
	jdff dff_A_eUpFYx1Q4_0(.dout(w_dff_A_9jyRWsz84_0),.din(w_dff_A_eUpFYx1Q4_0),.clk(gclk));
	jdff dff_A_9jyRWsz84_0(.dout(w_dff_A_cEOuKijU0_0),.din(w_dff_A_9jyRWsz84_0),.clk(gclk));
	jdff dff_A_cEOuKijU0_0(.dout(w_dff_A_U1dLwSpL4_0),.din(w_dff_A_cEOuKijU0_0),.clk(gclk));
	jdff dff_A_U1dLwSpL4_0(.dout(w_dff_A_qJrjx8857_0),.din(w_dff_A_U1dLwSpL4_0),.clk(gclk));
	jdff dff_A_qJrjx8857_0(.dout(w_dff_A_6YM9uwZO4_0),.din(w_dff_A_qJrjx8857_0),.clk(gclk));
	jdff dff_A_6YM9uwZO4_0(.dout(w_dff_A_bMHsJKsV9_0),.din(w_dff_A_6YM9uwZO4_0),.clk(gclk));
	jdff dff_A_bMHsJKsV9_0(.dout(w_dff_A_l7qQ59Ii4_0),.din(w_dff_A_bMHsJKsV9_0),.clk(gclk));
	jdff dff_A_l7qQ59Ii4_0(.dout(w_dff_A_85XxBP1b8_0),.din(w_dff_A_l7qQ59Ii4_0),.clk(gclk));
	jdff dff_A_85XxBP1b8_0(.dout(w_dff_A_SMiNRLFk5_0),.din(w_dff_A_85XxBP1b8_0),.clk(gclk));
	jdff dff_A_SMiNRLFk5_0(.dout(w_dff_A_0aw2phkN3_0),.din(w_dff_A_SMiNRLFk5_0),.clk(gclk));
	jdff dff_A_0aw2phkN3_0(.dout(w_dff_A_4MAuS9uP6_0),.din(w_dff_A_0aw2phkN3_0),.clk(gclk));
	jdff dff_A_4MAuS9uP6_0(.dout(w_dff_A_eqCk8I1c9_0),.din(w_dff_A_4MAuS9uP6_0),.clk(gclk));
	jdff dff_A_eqCk8I1c9_0(.dout(w_dff_A_zQJHRcpS0_0),.din(w_dff_A_eqCk8I1c9_0),.clk(gclk));
	jdff dff_A_zQJHRcpS0_0(.dout(w_dff_A_F4v23b1g8_0),.din(w_dff_A_zQJHRcpS0_0),.clk(gclk));
	jdff dff_A_F4v23b1g8_0(.dout(w_dff_A_ONfuArJk5_0),.din(w_dff_A_F4v23b1g8_0),.clk(gclk));
	jdff dff_A_ONfuArJk5_0(.dout(w_dff_A_B31WohRv9_0),.din(w_dff_A_ONfuArJk5_0),.clk(gclk));
	jdff dff_A_B31WohRv9_0(.dout(w_dff_A_56J56wQp5_0),.din(w_dff_A_B31WohRv9_0),.clk(gclk));
	jdff dff_A_56J56wQp5_0(.dout(w_dff_A_M4bXR5LO2_0),.din(w_dff_A_56J56wQp5_0),.clk(gclk));
	jdff dff_A_M4bXR5LO2_0(.dout(w_dff_A_cSeaWL8f3_0),.din(w_dff_A_M4bXR5LO2_0),.clk(gclk));
	jdff dff_A_cSeaWL8f3_0(.dout(w_dff_A_tXdSZS8I1_0),.din(w_dff_A_cSeaWL8f3_0),.clk(gclk));
	jdff dff_A_tXdSZS8I1_0(.dout(w_dff_A_ZTusLnzd9_0),.din(w_dff_A_tXdSZS8I1_0),.clk(gclk));
	jdff dff_A_ZTusLnzd9_0(.dout(w_dff_A_niCrNmJs9_0),.din(w_dff_A_ZTusLnzd9_0),.clk(gclk));
	jdff dff_A_niCrNmJs9_0(.dout(G603),.din(w_dff_A_niCrNmJs9_0),.clk(gclk));
	jdff dff_A_xFbNgCE53_1(.dout(w_dff_A_5893aecq4_0),.din(w_dff_A_xFbNgCE53_1),.clk(gclk));
	jdff dff_A_5893aecq4_0(.dout(w_dff_A_GIAAGkXz9_0),.din(w_dff_A_5893aecq4_0),.clk(gclk));
	jdff dff_A_GIAAGkXz9_0(.dout(w_dff_A_UwzRAMYG4_0),.din(w_dff_A_GIAAGkXz9_0),.clk(gclk));
	jdff dff_A_UwzRAMYG4_0(.dout(w_dff_A_SDc5B45W1_0),.din(w_dff_A_UwzRAMYG4_0),.clk(gclk));
	jdff dff_A_SDc5B45W1_0(.dout(w_dff_A_r0iswRXw1_0),.din(w_dff_A_SDc5B45W1_0),.clk(gclk));
	jdff dff_A_r0iswRXw1_0(.dout(w_dff_A_yVCieAOq5_0),.din(w_dff_A_r0iswRXw1_0),.clk(gclk));
	jdff dff_A_yVCieAOq5_0(.dout(w_dff_A_3WVmII6p7_0),.din(w_dff_A_yVCieAOq5_0),.clk(gclk));
	jdff dff_A_3WVmII6p7_0(.dout(w_dff_A_uUYAF0u26_0),.din(w_dff_A_3WVmII6p7_0),.clk(gclk));
	jdff dff_A_uUYAF0u26_0(.dout(w_dff_A_14UI74mt7_0),.din(w_dff_A_uUYAF0u26_0),.clk(gclk));
	jdff dff_A_14UI74mt7_0(.dout(w_dff_A_99ogk7Wt1_0),.din(w_dff_A_14UI74mt7_0),.clk(gclk));
	jdff dff_A_99ogk7Wt1_0(.dout(w_dff_A_QlvLiMzP3_0),.din(w_dff_A_99ogk7Wt1_0),.clk(gclk));
	jdff dff_A_QlvLiMzP3_0(.dout(w_dff_A_6jDRWn8f6_0),.din(w_dff_A_QlvLiMzP3_0),.clk(gclk));
	jdff dff_A_6jDRWn8f6_0(.dout(w_dff_A_iDhn2Ez91_0),.din(w_dff_A_6jDRWn8f6_0),.clk(gclk));
	jdff dff_A_iDhn2Ez91_0(.dout(w_dff_A_2L4os6hZ9_0),.din(w_dff_A_iDhn2Ez91_0),.clk(gclk));
	jdff dff_A_2L4os6hZ9_0(.dout(w_dff_A_bJeOn2mx4_0),.din(w_dff_A_2L4os6hZ9_0),.clk(gclk));
	jdff dff_A_bJeOn2mx4_0(.dout(w_dff_A_5RDOpVQg8_0),.din(w_dff_A_bJeOn2mx4_0),.clk(gclk));
	jdff dff_A_5RDOpVQg8_0(.dout(w_dff_A_Nw4UiyEO0_0),.din(w_dff_A_5RDOpVQg8_0),.clk(gclk));
	jdff dff_A_Nw4UiyEO0_0(.dout(w_dff_A_TiAHNh6O2_0),.din(w_dff_A_Nw4UiyEO0_0),.clk(gclk));
	jdff dff_A_TiAHNh6O2_0(.dout(w_dff_A_1SWJcjHW5_0),.din(w_dff_A_TiAHNh6O2_0),.clk(gclk));
	jdff dff_A_1SWJcjHW5_0(.dout(w_dff_A_8GAHJglx9_0),.din(w_dff_A_1SWJcjHW5_0),.clk(gclk));
	jdff dff_A_8GAHJglx9_0(.dout(w_dff_A_AETZv4DY2_0),.din(w_dff_A_8GAHJglx9_0),.clk(gclk));
	jdff dff_A_AETZv4DY2_0(.dout(w_dff_A_5dYYkKEV6_0),.din(w_dff_A_AETZv4DY2_0),.clk(gclk));
	jdff dff_A_5dYYkKEV6_0(.dout(w_dff_A_12FzcyT90_0),.din(w_dff_A_5dYYkKEV6_0),.clk(gclk));
	jdff dff_A_12FzcyT90_0(.dout(w_dff_A_ub9PuNV94_0),.din(w_dff_A_12FzcyT90_0),.clk(gclk));
	jdff dff_A_ub9PuNV94_0(.dout(w_dff_A_1VprEJfk0_0),.din(w_dff_A_ub9PuNV94_0),.clk(gclk));
	jdff dff_A_1VprEJfk0_0(.dout(w_dff_A_Rx9e6H5w5_0),.din(w_dff_A_1VprEJfk0_0),.clk(gclk));
	jdff dff_A_Rx9e6H5w5_0(.dout(G604),.din(w_dff_A_Rx9e6H5w5_0),.clk(gclk));
	jdff dff_A_myx6F0wm9_1(.dout(w_dff_A_UPbPSexA2_0),.din(w_dff_A_myx6F0wm9_1),.clk(gclk));
	jdff dff_A_UPbPSexA2_0(.dout(w_dff_A_SKSuOZ973_0),.din(w_dff_A_UPbPSexA2_0),.clk(gclk));
	jdff dff_A_SKSuOZ973_0(.dout(w_dff_A_bC6iMBGw3_0),.din(w_dff_A_SKSuOZ973_0),.clk(gclk));
	jdff dff_A_bC6iMBGw3_0(.dout(w_dff_A_QORnzm0y5_0),.din(w_dff_A_bC6iMBGw3_0),.clk(gclk));
	jdff dff_A_QORnzm0y5_0(.dout(w_dff_A_OWgtybLQ2_0),.din(w_dff_A_QORnzm0y5_0),.clk(gclk));
	jdff dff_A_OWgtybLQ2_0(.dout(w_dff_A_shekAVmn9_0),.din(w_dff_A_OWgtybLQ2_0),.clk(gclk));
	jdff dff_A_shekAVmn9_0(.dout(w_dff_A_BlVWxxaJ9_0),.din(w_dff_A_shekAVmn9_0),.clk(gclk));
	jdff dff_A_BlVWxxaJ9_0(.dout(w_dff_A_ttLcXXNe3_0),.din(w_dff_A_BlVWxxaJ9_0),.clk(gclk));
	jdff dff_A_ttLcXXNe3_0(.dout(w_dff_A_2zaXesmB2_0),.din(w_dff_A_ttLcXXNe3_0),.clk(gclk));
	jdff dff_A_2zaXesmB2_0(.dout(w_dff_A_17yAvfwv3_0),.din(w_dff_A_2zaXesmB2_0),.clk(gclk));
	jdff dff_A_17yAvfwv3_0(.dout(w_dff_A_7zb7YPEd1_0),.din(w_dff_A_17yAvfwv3_0),.clk(gclk));
	jdff dff_A_7zb7YPEd1_0(.dout(w_dff_A_JnvVGCU53_0),.din(w_dff_A_7zb7YPEd1_0),.clk(gclk));
	jdff dff_A_JnvVGCU53_0(.dout(w_dff_A_MR65cec07_0),.din(w_dff_A_JnvVGCU53_0),.clk(gclk));
	jdff dff_A_MR65cec07_0(.dout(w_dff_A_GUMvMTUg2_0),.din(w_dff_A_MR65cec07_0),.clk(gclk));
	jdff dff_A_GUMvMTUg2_0(.dout(w_dff_A_q1ryTd3G0_0),.din(w_dff_A_GUMvMTUg2_0),.clk(gclk));
	jdff dff_A_q1ryTd3G0_0(.dout(w_dff_A_r1NabILy2_0),.din(w_dff_A_q1ryTd3G0_0),.clk(gclk));
	jdff dff_A_r1NabILy2_0(.dout(w_dff_A_yNOMKLxZ6_0),.din(w_dff_A_r1NabILy2_0),.clk(gclk));
	jdff dff_A_yNOMKLxZ6_0(.dout(w_dff_A_iZ4HgfDc1_0),.din(w_dff_A_yNOMKLxZ6_0),.clk(gclk));
	jdff dff_A_iZ4HgfDc1_0(.dout(w_dff_A_nV6Otl9y6_0),.din(w_dff_A_iZ4HgfDc1_0),.clk(gclk));
	jdff dff_A_nV6Otl9y6_0(.dout(w_dff_A_Ow890cCz1_0),.din(w_dff_A_nV6Otl9y6_0),.clk(gclk));
	jdff dff_A_Ow890cCz1_0(.dout(w_dff_A_S2SnoV9C1_0),.din(w_dff_A_Ow890cCz1_0),.clk(gclk));
	jdff dff_A_S2SnoV9C1_0(.dout(w_dff_A_UFtKd3I17_0),.din(w_dff_A_S2SnoV9C1_0),.clk(gclk));
	jdff dff_A_UFtKd3I17_0(.dout(w_dff_A_RtH6a8AC7_0),.din(w_dff_A_UFtKd3I17_0),.clk(gclk));
	jdff dff_A_RtH6a8AC7_0(.dout(w_dff_A_xkoRBOk70_0),.din(w_dff_A_RtH6a8AC7_0),.clk(gclk));
	jdff dff_A_xkoRBOk70_0(.dout(w_dff_A_Ip0SWz022_0),.din(w_dff_A_xkoRBOk70_0),.clk(gclk));
	jdff dff_A_Ip0SWz022_0(.dout(w_dff_A_F2VHMPQ78_0),.din(w_dff_A_Ip0SWz022_0),.clk(gclk));
	jdff dff_A_F2VHMPQ78_0(.dout(G611),.din(w_dff_A_F2VHMPQ78_0),.clk(gclk));
	jdff dff_A_ICrsPWT71_1(.dout(w_dff_A_PwUBf2Dt3_0),.din(w_dff_A_ICrsPWT71_1),.clk(gclk));
	jdff dff_A_PwUBf2Dt3_0(.dout(w_dff_A_ejEYJ2y29_0),.din(w_dff_A_PwUBf2Dt3_0),.clk(gclk));
	jdff dff_A_ejEYJ2y29_0(.dout(w_dff_A_zUDYgoom1_0),.din(w_dff_A_ejEYJ2y29_0),.clk(gclk));
	jdff dff_A_zUDYgoom1_0(.dout(w_dff_A_mmYMCBTp6_0),.din(w_dff_A_zUDYgoom1_0),.clk(gclk));
	jdff dff_A_mmYMCBTp6_0(.dout(w_dff_A_hKYDvdL87_0),.din(w_dff_A_mmYMCBTp6_0),.clk(gclk));
	jdff dff_A_hKYDvdL87_0(.dout(w_dff_A_iJoOZddR5_0),.din(w_dff_A_hKYDvdL87_0),.clk(gclk));
	jdff dff_A_iJoOZddR5_0(.dout(w_dff_A_mMv9XXRP0_0),.din(w_dff_A_iJoOZddR5_0),.clk(gclk));
	jdff dff_A_mMv9XXRP0_0(.dout(w_dff_A_1lJy1rlA8_0),.din(w_dff_A_mMv9XXRP0_0),.clk(gclk));
	jdff dff_A_1lJy1rlA8_0(.dout(w_dff_A_Ek8V9XCu6_0),.din(w_dff_A_1lJy1rlA8_0),.clk(gclk));
	jdff dff_A_Ek8V9XCu6_0(.dout(w_dff_A_za8WoKtK7_0),.din(w_dff_A_Ek8V9XCu6_0),.clk(gclk));
	jdff dff_A_za8WoKtK7_0(.dout(w_dff_A_jgz879Xc9_0),.din(w_dff_A_za8WoKtK7_0),.clk(gclk));
	jdff dff_A_jgz879Xc9_0(.dout(w_dff_A_3YbwhwE11_0),.din(w_dff_A_jgz879Xc9_0),.clk(gclk));
	jdff dff_A_3YbwhwE11_0(.dout(w_dff_A_ags6rIIn5_0),.din(w_dff_A_3YbwhwE11_0),.clk(gclk));
	jdff dff_A_ags6rIIn5_0(.dout(w_dff_A_kFUpKGHf1_0),.din(w_dff_A_ags6rIIn5_0),.clk(gclk));
	jdff dff_A_kFUpKGHf1_0(.dout(w_dff_A_pDtrcHpW6_0),.din(w_dff_A_kFUpKGHf1_0),.clk(gclk));
	jdff dff_A_pDtrcHpW6_0(.dout(w_dff_A_MnISrHh18_0),.din(w_dff_A_pDtrcHpW6_0),.clk(gclk));
	jdff dff_A_MnISrHh18_0(.dout(w_dff_A_QRIQjPyF8_0),.din(w_dff_A_MnISrHh18_0),.clk(gclk));
	jdff dff_A_QRIQjPyF8_0(.dout(w_dff_A_sWlWgiQ21_0),.din(w_dff_A_QRIQjPyF8_0),.clk(gclk));
	jdff dff_A_sWlWgiQ21_0(.dout(w_dff_A_Tbd5q3mP1_0),.din(w_dff_A_sWlWgiQ21_0),.clk(gclk));
	jdff dff_A_Tbd5q3mP1_0(.dout(w_dff_A_Af1WBMLx1_0),.din(w_dff_A_Tbd5q3mP1_0),.clk(gclk));
	jdff dff_A_Af1WBMLx1_0(.dout(w_dff_A_lqXiPWlu4_0),.din(w_dff_A_Af1WBMLx1_0),.clk(gclk));
	jdff dff_A_lqXiPWlu4_0(.dout(w_dff_A_pmC392pt7_0),.din(w_dff_A_lqXiPWlu4_0),.clk(gclk));
	jdff dff_A_pmC392pt7_0(.dout(w_dff_A_D3CK5Nub1_0),.din(w_dff_A_pmC392pt7_0),.clk(gclk));
	jdff dff_A_D3CK5Nub1_0(.dout(w_dff_A_HiEfJDVg9_0),.din(w_dff_A_D3CK5Nub1_0),.clk(gclk));
	jdff dff_A_HiEfJDVg9_0(.dout(w_dff_A_WzXcBO7K7_0),.din(w_dff_A_HiEfJDVg9_0),.clk(gclk));
	jdff dff_A_WzXcBO7K7_0(.dout(w_dff_A_Js0F6f5W7_0),.din(w_dff_A_WzXcBO7K7_0),.clk(gclk));
	jdff dff_A_Js0F6f5W7_0(.dout(G612),.din(w_dff_A_Js0F6f5W7_0),.clk(gclk));
	jdff dff_A_7QTZeYzo7_2(.dout(w_dff_A_GKPCB9Sa5_0),.din(w_dff_A_7QTZeYzo7_2),.clk(gclk));
	jdff dff_A_GKPCB9Sa5_0(.dout(w_dff_A_hPEAL11N7_0),.din(w_dff_A_GKPCB9Sa5_0),.clk(gclk));
	jdff dff_A_hPEAL11N7_0(.dout(w_dff_A_l86Jl5LI4_0),.din(w_dff_A_hPEAL11N7_0),.clk(gclk));
	jdff dff_A_l86Jl5LI4_0(.dout(w_dff_A_iJg4hL9o0_0),.din(w_dff_A_l86Jl5LI4_0),.clk(gclk));
	jdff dff_A_iJg4hL9o0_0(.dout(w_dff_A_3NxsMPhs9_0),.din(w_dff_A_iJg4hL9o0_0),.clk(gclk));
	jdff dff_A_3NxsMPhs9_0(.dout(w_dff_A_LTz9gH5m4_0),.din(w_dff_A_3NxsMPhs9_0),.clk(gclk));
	jdff dff_A_LTz9gH5m4_0(.dout(w_dff_A_iIf1YJl75_0),.din(w_dff_A_LTz9gH5m4_0),.clk(gclk));
	jdff dff_A_iIf1YJl75_0(.dout(w_dff_A_2wgJWx869_0),.din(w_dff_A_iIf1YJl75_0),.clk(gclk));
	jdff dff_A_2wgJWx869_0(.dout(w_dff_A_i1KxliVk9_0),.din(w_dff_A_2wgJWx869_0),.clk(gclk));
	jdff dff_A_i1KxliVk9_0(.dout(w_dff_A_qbU5CQJt0_0),.din(w_dff_A_i1KxliVk9_0),.clk(gclk));
	jdff dff_A_qbU5CQJt0_0(.dout(w_dff_A_qAV053ju7_0),.din(w_dff_A_qbU5CQJt0_0),.clk(gclk));
	jdff dff_A_qAV053ju7_0(.dout(w_dff_A_tN3hkU5U5_0),.din(w_dff_A_qAV053ju7_0),.clk(gclk));
	jdff dff_A_tN3hkU5U5_0(.dout(w_dff_A_0IpKMhuG4_0),.din(w_dff_A_tN3hkU5U5_0),.clk(gclk));
	jdff dff_A_0IpKMhuG4_0(.dout(w_dff_A_H8Soonyh7_0),.din(w_dff_A_0IpKMhuG4_0),.clk(gclk));
	jdff dff_A_H8Soonyh7_0(.dout(w_dff_A_I9015LC60_0),.din(w_dff_A_H8Soonyh7_0),.clk(gclk));
	jdff dff_A_I9015LC60_0(.dout(w_dff_A_Pdyd3hMk8_0),.din(w_dff_A_I9015LC60_0),.clk(gclk));
	jdff dff_A_Pdyd3hMk8_0(.dout(w_dff_A_JSPV5HPF4_0),.din(w_dff_A_Pdyd3hMk8_0),.clk(gclk));
	jdff dff_A_JSPV5HPF4_0(.dout(w_dff_A_kGL9ChU40_0),.din(w_dff_A_JSPV5HPF4_0),.clk(gclk));
	jdff dff_A_kGL9ChU40_0(.dout(w_dff_A_UGxOMLY81_0),.din(w_dff_A_kGL9ChU40_0),.clk(gclk));
	jdff dff_A_UGxOMLY81_0(.dout(w_dff_A_ZN6s2Yu81_0),.din(w_dff_A_UGxOMLY81_0),.clk(gclk));
	jdff dff_A_ZN6s2Yu81_0(.dout(w_dff_A_uDXdqO9o8_0),.din(w_dff_A_ZN6s2Yu81_0),.clk(gclk));
	jdff dff_A_uDXdqO9o8_0(.dout(w_dff_A_0I6ypgUF7_0),.din(w_dff_A_uDXdqO9o8_0),.clk(gclk));
	jdff dff_A_0I6ypgUF7_0(.dout(w_dff_A_7avwLBt46_0),.din(w_dff_A_0I6ypgUF7_0),.clk(gclk));
	jdff dff_A_7avwLBt46_0(.dout(w_dff_A_YrTK3Fc87_0),.din(w_dff_A_7avwLBt46_0),.clk(gclk));
	jdff dff_A_YrTK3Fc87_0(.dout(w_dff_A_1hjW2mnA6_0),.din(w_dff_A_YrTK3Fc87_0),.clk(gclk));
	jdff dff_A_1hjW2mnA6_0(.dout(w_dff_A_C6jLwmaC6_0),.din(w_dff_A_1hjW2mnA6_0),.clk(gclk));
	jdff dff_A_C6jLwmaC6_0(.dout(G810),.din(w_dff_A_C6jLwmaC6_0),.clk(gclk));
	jdff dff_A_aACQTVri0_1(.dout(w_dff_A_LwA9mG537_0),.din(w_dff_A_aACQTVri0_1),.clk(gclk));
	jdff dff_A_LwA9mG537_0(.dout(w_dff_A_jGHiufHt5_0),.din(w_dff_A_LwA9mG537_0),.clk(gclk));
	jdff dff_A_jGHiufHt5_0(.dout(w_dff_A_dQu7MDDI8_0),.din(w_dff_A_jGHiufHt5_0),.clk(gclk));
	jdff dff_A_dQu7MDDI8_0(.dout(w_dff_A_pxAoMv8v9_0),.din(w_dff_A_dQu7MDDI8_0),.clk(gclk));
	jdff dff_A_pxAoMv8v9_0(.dout(w_dff_A_fwb8saOd2_0),.din(w_dff_A_pxAoMv8v9_0),.clk(gclk));
	jdff dff_A_fwb8saOd2_0(.dout(w_dff_A_K7AggtN31_0),.din(w_dff_A_fwb8saOd2_0),.clk(gclk));
	jdff dff_A_K7AggtN31_0(.dout(w_dff_A_cbt7OtFF1_0),.din(w_dff_A_K7AggtN31_0),.clk(gclk));
	jdff dff_A_cbt7OtFF1_0(.dout(w_dff_A_LFJ0a3Ok5_0),.din(w_dff_A_cbt7OtFF1_0),.clk(gclk));
	jdff dff_A_LFJ0a3Ok5_0(.dout(w_dff_A_JgF2gRN58_0),.din(w_dff_A_LFJ0a3Ok5_0),.clk(gclk));
	jdff dff_A_JgF2gRN58_0(.dout(w_dff_A_pmc21HvS8_0),.din(w_dff_A_JgF2gRN58_0),.clk(gclk));
	jdff dff_A_pmc21HvS8_0(.dout(w_dff_A_GdlUhXSt2_0),.din(w_dff_A_pmc21HvS8_0),.clk(gclk));
	jdff dff_A_GdlUhXSt2_0(.dout(w_dff_A_ruJevEXR0_0),.din(w_dff_A_GdlUhXSt2_0),.clk(gclk));
	jdff dff_A_ruJevEXR0_0(.dout(w_dff_A_McHwuMQ00_0),.din(w_dff_A_ruJevEXR0_0),.clk(gclk));
	jdff dff_A_McHwuMQ00_0(.dout(w_dff_A_Akw6YEm68_0),.din(w_dff_A_McHwuMQ00_0),.clk(gclk));
	jdff dff_A_Akw6YEm68_0(.dout(w_dff_A_3X7OKRyH5_0),.din(w_dff_A_Akw6YEm68_0),.clk(gclk));
	jdff dff_A_3X7OKRyH5_0(.dout(w_dff_A_PO5r0l5i0_0),.din(w_dff_A_3X7OKRyH5_0),.clk(gclk));
	jdff dff_A_PO5r0l5i0_0(.dout(w_dff_A_sgOvqIYj5_0),.din(w_dff_A_PO5r0l5i0_0),.clk(gclk));
	jdff dff_A_sgOvqIYj5_0(.dout(w_dff_A_Sb7svTrN6_0),.din(w_dff_A_sgOvqIYj5_0),.clk(gclk));
	jdff dff_A_Sb7svTrN6_0(.dout(w_dff_A_MRVGfrX30_0),.din(w_dff_A_Sb7svTrN6_0),.clk(gclk));
	jdff dff_A_MRVGfrX30_0(.dout(w_dff_A_SMApoT755_0),.din(w_dff_A_MRVGfrX30_0),.clk(gclk));
	jdff dff_A_SMApoT755_0(.dout(w_dff_A_yFe9BGHJ4_0),.din(w_dff_A_SMApoT755_0),.clk(gclk));
	jdff dff_A_yFe9BGHJ4_0(.dout(w_dff_A_1SmvKHDK6_0),.din(w_dff_A_yFe9BGHJ4_0),.clk(gclk));
	jdff dff_A_1SmvKHDK6_0(.dout(w_dff_A_XYOhwMu25_0),.din(w_dff_A_1SmvKHDK6_0),.clk(gclk));
	jdff dff_A_XYOhwMu25_0(.dout(w_dff_A_IjEbgNNA6_0),.din(w_dff_A_XYOhwMu25_0),.clk(gclk));
	jdff dff_A_IjEbgNNA6_0(.dout(w_dff_A_9bt5RQ0b4_0),.din(w_dff_A_IjEbgNNA6_0),.clk(gclk));
	jdff dff_A_9bt5RQ0b4_0(.dout(w_dff_A_j8wplm9r5_0),.din(w_dff_A_9bt5RQ0b4_0),.clk(gclk));
	jdff dff_A_j8wplm9r5_0(.dout(G848),.din(w_dff_A_j8wplm9r5_0),.clk(gclk));
	jdff dff_A_GGl98Dw74_1(.dout(w_dff_A_7fjAglrO2_0),.din(w_dff_A_GGl98Dw74_1),.clk(gclk));
	jdff dff_A_7fjAglrO2_0(.dout(w_dff_A_XThLXVq02_0),.din(w_dff_A_7fjAglrO2_0),.clk(gclk));
	jdff dff_A_XThLXVq02_0(.dout(w_dff_A_guqdJuRK9_0),.din(w_dff_A_XThLXVq02_0),.clk(gclk));
	jdff dff_A_guqdJuRK9_0(.dout(w_dff_A_1SwR83JX8_0),.din(w_dff_A_guqdJuRK9_0),.clk(gclk));
	jdff dff_A_1SwR83JX8_0(.dout(w_dff_A_A19UkKn51_0),.din(w_dff_A_1SwR83JX8_0),.clk(gclk));
	jdff dff_A_A19UkKn51_0(.dout(w_dff_A_YQL2e9g54_0),.din(w_dff_A_A19UkKn51_0),.clk(gclk));
	jdff dff_A_YQL2e9g54_0(.dout(w_dff_A_GcbbKzAH6_0),.din(w_dff_A_YQL2e9g54_0),.clk(gclk));
	jdff dff_A_GcbbKzAH6_0(.dout(w_dff_A_wgZzcywv2_0),.din(w_dff_A_GcbbKzAH6_0),.clk(gclk));
	jdff dff_A_wgZzcywv2_0(.dout(w_dff_A_PldWPQ5A2_0),.din(w_dff_A_wgZzcywv2_0),.clk(gclk));
	jdff dff_A_PldWPQ5A2_0(.dout(w_dff_A_Y92iBXCG4_0),.din(w_dff_A_PldWPQ5A2_0),.clk(gclk));
	jdff dff_A_Y92iBXCG4_0(.dout(w_dff_A_XMUZeDWV4_0),.din(w_dff_A_Y92iBXCG4_0),.clk(gclk));
	jdff dff_A_XMUZeDWV4_0(.dout(w_dff_A_u3W0J0Um6_0),.din(w_dff_A_XMUZeDWV4_0),.clk(gclk));
	jdff dff_A_u3W0J0Um6_0(.dout(w_dff_A_dlgQr5Jj5_0),.din(w_dff_A_u3W0J0Um6_0),.clk(gclk));
	jdff dff_A_dlgQr5Jj5_0(.dout(w_dff_A_iZUt9QcP7_0),.din(w_dff_A_dlgQr5Jj5_0),.clk(gclk));
	jdff dff_A_iZUt9QcP7_0(.dout(w_dff_A_ddDbZ63u6_0),.din(w_dff_A_iZUt9QcP7_0),.clk(gclk));
	jdff dff_A_ddDbZ63u6_0(.dout(w_dff_A_kBNOjV2F0_0),.din(w_dff_A_ddDbZ63u6_0),.clk(gclk));
	jdff dff_A_kBNOjV2F0_0(.dout(w_dff_A_hXM72C1y1_0),.din(w_dff_A_kBNOjV2F0_0),.clk(gclk));
	jdff dff_A_hXM72C1y1_0(.dout(w_dff_A_runAglZL5_0),.din(w_dff_A_hXM72C1y1_0),.clk(gclk));
	jdff dff_A_runAglZL5_0(.dout(w_dff_A_PeYKnPUy0_0),.din(w_dff_A_runAglZL5_0),.clk(gclk));
	jdff dff_A_PeYKnPUy0_0(.dout(w_dff_A_kLpdds3F5_0),.din(w_dff_A_PeYKnPUy0_0),.clk(gclk));
	jdff dff_A_kLpdds3F5_0(.dout(w_dff_A_F2BeMjGk0_0),.din(w_dff_A_kLpdds3F5_0),.clk(gclk));
	jdff dff_A_F2BeMjGk0_0(.dout(w_dff_A_fu3FUC8D8_0),.din(w_dff_A_F2BeMjGk0_0),.clk(gclk));
	jdff dff_A_fu3FUC8D8_0(.dout(w_dff_A_NKnQs0Ww5_0),.din(w_dff_A_fu3FUC8D8_0),.clk(gclk));
	jdff dff_A_NKnQs0Ww5_0(.dout(w_dff_A_rJjBTX8p7_0),.din(w_dff_A_NKnQs0Ww5_0),.clk(gclk));
	jdff dff_A_rJjBTX8p7_0(.dout(w_dff_A_I6nzBz4j0_0),.din(w_dff_A_rJjBTX8p7_0),.clk(gclk));
	jdff dff_A_I6nzBz4j0_0(.dout(w_dff_A_BPa1Y1LR5_0),.din(w_dff_A_I6nzBz4j0_0),.clk(gclk));
	jdff dff_A_BPa1Y1LR5_0(.dout(G849),.din(w_dff_A_BPa1Y1LR5_0),.clk(gclk));
	jdff dff_A_SSAqx4n50_1(.dout(w_dff_A_cr9RgTlP6_0),.din(w_dff_A_SSAqx4n50_1),.clk(gclk));
	jdff dff_A_cr9RgTlP6_0(.dout(w_dff_A_FB44OejC9_0),.din(w_dff_A_cr9RgTlP6_0),.clk(gclk));
	jdff dff_A_FB44OejC9_0(.dout(w_dff_A_SnEljJZ02_0),.din(w_dff_A_FB44OejC9_0),.clk(gclk));
	jdff dff_A_SnEljJZ02_0(.dout(w_dff_A_TMteaZIn9_0),.din(w_dff_A_SnEljJZ02_0),.clk(gclk));
	jdff dff_A_TMteaZIn9_0(.dout(w_dff_A_qevtscPe9_0),.din(w_dff_A_TMteaZIn9_0),.clk(gclk));
	jdff dff_A_qevtscPe9_0(.dout(w_dff_A_8ZexlqBd3_0),.din(w_dff_A_qevtscPe9_0),.clk(gclk));
	jdff dff_A_8ZexlqBd3_0(.dout(w_dff_A_NWHFzZc57_0),.din(w_dff_A_8ZexlqBd3_0),.clk(gclk));
	jdff dff_A_NWHFzZc57_0(.dout(w_dff_A_TIoK4kMv6_0),.din(w_dff_A_NWHFzZc57_0),.clk(gclk));
	jdff dff_A_TIoK4kMv6_0(.dout(w_dff_A_Yi6o9clo9_0),.din(w_dff_A_TIoK4kMv6_0),.clk(gclk));
	jdff dff_A_Yi6o9clo9_0(.dout(w_dff_A_dbWxIeWy7_0),.din(w_dff_A_Yi6o9clo9_0),.clk(gclk));
	jdff dff_A_dbWxIeWy7_0(.dout(w_dff_A_w29kXXER8_0),.din(w_dff_A_dbWxIeWy7_0),.clk(gclk));
	jdff dff_A_w29kXXER8_0(.dout(w_dff_A_tfZsEWzc3_0),.din(w_dff_A_w29kXXER8_0),.clk(gclk));
	jdff dff_A_tfZsEWzc3_0(.dout(w_dff_A_C2vpX75T4_0),.din(w_dff_A_tfZsEWzc3_0),.clk(gclk));
	jdff dff_A_C2vpX75T4_0(.dout(w_dff_A_GwFpnkWH7_0),.din(w_dff_A_C2vpX75T4_0),.clk(gclk));
	jdff dff_A_GwFpnkWH7_0(.dout(w_dff_A_wUciIsyg1_0),.din(w_dff_A_GwFpnkWH7_0),.clk(gclk));
	jdff dff_A_wUciIsyg1_0(.dout(w_dff_A_GFDUZido9_0),.din(w_dff_A_wUciIsyg1_0),.clk(gclk));
	jdff dff_A_GFDUZido9_0(.dout(w_dff_A_iuXFaMRO5_0),.din(w_dff_A_GFDUZido9_0),.clk(gclk));
	jdff dff_A_iuXFaMRO5_0(.dout(w_dff_A_050FeFT91_0),.din(w_dff_A_iuXFaMRO5_0),.clk(gclk));
	jdff dff_A_050FeFT91_0(.dout(w_dff_A_wqbvMCEV7_0),.din(w_dff_A_050FeFT91_0),.clk(gclk));
	jdff dff_A_wqbvMCEV7_0(.dout(w_dff_A_aKzwPIWl6_0),.din(w_dff_A_wqbvMCEV7_0),.clk(gclk));
	jdff dff_A_aKzwPIWl6_0(.dout(w_dff_A_YoYnhh8B7_0),.din(w_dff_A_aKzwPIWl6_0),.clk(gclk));
	jdff dff_A_YoYnhh8B7_0(.dout(w_dff_A_Djp167xu6_0),.din(w_dff_A_YoYnhh8B7_0),.clk(gclk));
	jdff dff_A_Djp167xu6_0(.dout(w_dff_A_O62PEz0Z7_0),.din(w_dff_A_Djp167xu6_0),.clk(gclk));
	jdff dff_A_O62PEz0Z7_0(.dout(w_dff_A_jipahLvn4_0),.din(w_dff_A_O62PEz0Z7_0),.clk(gclk));
	jdff dff_A_jipahLvn4_0(.dout(w_dff_A_gNCqqYGt2_0),.din(w_dff_A_jipahLvn4_0),.clk(gclk));
	jdff dff_A_gNCqqYGt2_0(.dout(w_dff_A_H6SLc7GP5_0),.din(w_dff_A_gNCqqYGt2_0),.clk(gclk));
	jdff dff_A_H6SLc7GP5_0(.dout(G850),.din(w_dff_A_H6SLc7GP5_0),.clk(gclk));
	jdff dff_A_DYNjfypZ7_1(.dout(w_dff_A_SXllwUeB1_0),.din(w_dff_A_DYNjfypZ7_1),.clk(gclk));
	jdff dff_A_SXllwUeB1_0(.dout(w_dff_A_k5Ibsu3p7_0),.din(w_dff_A_SXllwUeB1_0),.clk(gclk));
	jdff dff_A_k5Ibsu3p7_0(.dout(w_dff_A_biIsWMuc3_0),.din(w_dff_A_k5Ibsu3p7_0),.clk(gclk));
	jdff dff_A_biIsWMuc3_0(.dout(w_dff_A_Kr1aarx15_0),.din(w_dff_A_biIsWMuc3_0),.clk(gclk));
	jdff dff_A_Kr1aarx15_0(.dout(w_dff_A_DkJhcVR97_0),.din(w_dff_A_Kr1aarx15_0),.clk(gclk));
	jdff dff_A_DkJhcVR97_0(.dout(w_dff_A_jTgN8fta8_0),.din(w_dff_A_DkJhcVR97_0),.clk(gclk));
	jdff dff_A_jTgN8fta8_0(.dout(w_dff_A_iML8XhOG3_0),.din(w_dff_A_jTgN8fta8_0),.clk(gclk));
	jdff dff_A_iML8XhOG3_0(.dout(w_dff_A_8Aet4vXu4_0),.din(w_dff_A_iML8XhOG3_0),.clk(gclk));
	jdff dff_A_8Aet4vXu4_0(.dout(w_dff_A_Js5oazjZ3_0),.din(w_dff_A_8Aet4vXu4_0),.clk(gclk));
	jdff dff_A_Js5oazjZ3_0(.dout(w_dff_A_BOCHaZHH5_0),.din(w_dff_A_Js5oazjZ3_0),.clk(gclk));
	jdff dff_A_BOCHaZHH5_0(.dout(w_dff_A_6wdpodPw6_0),.din(w_dff_A_BOCHaZHH5_0),.clk(gclk));
	jdff dff_A_6wdpodPw6_0(.dout(w_dff_A_zDEwES4z6_0),.din(w_dff_A_6wdpodPw6_0),.clk(gclk));
	jdff dff_A_zDEwES4z6_0(.dout(w_dff_A_yEzLuGhL0_0),.din(w_dff_A_zDEwES4z6_0),.clk(gclk));
	jdff dff_A_yEzLuGhL0_0(.dout(w_dff_A_Qq2DYUyR9_0),.din(w_dff_A_yEzLuGhL0_0),.clk(gclk));
	jdff dff_A_Qq2DYUyR9_0(.dout(w_dff_A_T7ZlTZ0P5_0),.din(w_dff_A_Qq2DYUyR9_0),.clk(gclk));
	jdff dff_A_T7ZlTZ0P5_0(.dout(w_dff_A_vgb0VQIe9_0),.din(w_dff_A_T7ZlTZ0P5_0),.clk(gclk));
	jdff dff_A_vgb0VQIe9_0(.dout(w_dff_A_LjnDNZyK1_0),.din(w_dff_A_vgb0VQIe9_0),.clk(gclk));
	jdff dff_A_LjnDNZyK1_0(.dout(w_dff_A_OQarA5w44_0),.din(w_dff_A_LjnDNZyK1_0),.clk(gclk));
	jdff dff_A_OQarA5w44_0(.dout(w_dff_A_GBG7CNlC0_0),.din(w_dff_A_OQarA5w44_0),.clk(gclk));
	jdff dff_A_GBG7CNlC0_0(.dout(w_dff_A_KTNGYh7P9_0),.din(w_dff_A_GBG7CNlC0_0),.clk(gclk));
	jdff dff_A_KTNGYh7P9_0(.dout(w_dff_A_aUv6D9Ez0_0),.din(w_dff_A_KTNGYh7P9_0),.clk(gclk));
	jdff dff_A_aUv6D9Ez0_0(.dout(w_dff_A_4Uh8XPLD4_0),.din(w_dff_A_aUv6D9Ez0_0),.clk(gclk));
	jdff dff_A_4Uh8XPLD4_0(.dout(w_dff_A_8oc1e8s20_0),.din(w_dff_A_4Uh8XPLD4_0),.clk(gclk));
	jdff dff_A_8oc1e8s20_0(.dout(w_dff_A_WjdJYfX37_0),.din(w_dff_A_8oc1e8s20_0),.clk(gclk));
	jdff dff_A_WjdJYfX37_0(.dout(w_dff_A_bLIr58ez0_0),.din(w_dff_A_WjdJYfX37_0),.clk(gclk));
	jdff dff_A_bLIr58ez0_0(.dout(w_dff_A_wej7VxvF9_0),.din(w_dff_A_bLIr58ez0_0),.clk(gclk));
	jdff dff_A_wej7VxvF9_0(.dout(G851),.din(w_dff_A_wej7VxvF9_0),.clk(gclk));
	jdff dff_A_z8qnRYpc3_2(.dout(w_dff_A_KSXl4TP58_0),.din(w_dff_A_z8qnRYpc3_2),.clk(gclk));
	jdff dff_A_KSXl4TP58_0(.dout(w_dff_A_4kRIGyic3_0),.din(w_dff_A_KSXl4TP58_0),.clk(gclk));
	jdff dff_A_4kRIGyic3_0(.dout(w_dff_A_6Mk5wrQW2_0),.din(w_dff_A_4kRIGyic3_0),.clk(gclk));
	jdff dff_A_6Mk5wrQW2_0(.dout(w_dff_A_2ri2mYmV2_0),.din(w_dff_A_6Mk5wrQW2_0),.clk(gclk));
	jdff dff_A_2ri2mYmV2_0(.dout(w_dff_A_PbMBeDGo4_0),.din(w_dff_A_2ri2mYmV2_0),.clk(gclk));
	jdff dff_A_PbMBeDGo4_0(.dout(w_dff_A_id4IJGMU3_0),.din(w_dff_A_PbMBeDGo4_0),.clk(gclk));
	jdff dff_A_id4IJGMU3_0(.dout(w_dff_A_ZDbmA7uH5_0),.din(w_dff_A_id4IJGMU3_0),.clk(gclk));
	jdff dff_A_ZDbmA7uH5_0(.dout(w_dff_A_nPJVA8tO1_0),.din(w_dff_A_ZDbmA7uH5_0),.clk(gclk));
	jdff dff_A_nPJVA8tO1_0(.dout(w_dff_A_7DhbAVRD6_0),.din(w_dff_A_nPJVA8tO1_0),.clk(gclk));
	jdff dff_A_7DhbAVRD6_0(.dout(w_dff_A_Hx3PPjQL0_0),.din(w_dff_A_7DhbAVRD6_0),.clk(gclk));
	jdff dff_A_Hx3PPjQL0_0(.dout(w_dff_A_AhdqAkx50_0),.din(w_dff_A_Hx3PPjQL0_0),.clk(gclk));
	jdff dff_A_AhdqAkx50_0(.dout(w_dff_A_9fliU4jh0_0),.din(w_dff_A_AhdqAkx50_0),.clk(gclk));
	jdff dff_A_9fliU4jh0_0(.dout(w_dff_A_pgZXVOqW9_0),.din(w_dff_A_9fliU4jh0_0),.clk(gclk));
	jdff dff_A_pgZXVOqW9_0(.dout(w_dff_A_pBgHZpUf1_0),.din(w_dff_A_pgZXVOqW9_0),.clk(gclk));
	jdff dff_A_pBgHZpUf1_0(.dout(w_dff_A_YenyigRT8_0),.din(w_dff_A_pBgHZpUf1_0),.clk(gclk));
	jdff dff_A_YenyigRT8_0(.dout(w_dff_A_EU6A3Fsr0_0),.din(w_dff_A_YenyigRT8_0),.clk(gclk));
	jdff dff_A_EU6A3Fsr0_0(.dout(w_dff_A_BZr8u2Y53_0),.din(w_dff_A_EU6A3Fsr0_0),.clk(gclk));
	jdff dff_A_BZr8u2Y53_0(.dout(w_dff_A_r6Jbh0ju9_0),.din(w_dff_A_BZr8u2Y53_0),.clk(gclk));
	jdff dff_A_r6Jbh0ju9_0(.dout(w_dff_A_080Svrp25_0),.din(w_dff_A_r6Jbh0ju9_0),.clk(gclk));
	jdff dff_A_080Svrp25_0(.dout(w_dff_A_zelzBhZh2_0),.din(w_dff_A_080Svrp25_0),.clk(gclk));
	jdff dff_A_zelzBhZh2_0(.dout(w_dff_A_tePGh3O03_0),.din(w_dff_A_zelzBhZh2_0),.clk(gclk));
	jdff dff_A_tePGh3O03_0(.dout(w_dff_A_WpEobw7u0_0),.din(w_dff_A_tePGh3O03_0),.clk(gclk));
	jdff dff_A_WpEobw7u0_0(.dout(w_dff_A_Hc1wxwZ89_0),.din(w_dff_A_WpEobw7u0_0),.clk(gclk));
	jdff dff_A_Hc1wxwZ89_0(.dout(w_dff_A_SXGBn3E45_0),.din(w_dff_A_Hc1wxwZ89_0),.clk(gclk));
	jdff dff_A_SXGBn3E45_0(.dout(w_dff_A_Pb3eeLyY6_0),.din(w_dff_A_SXGBn3E45_0),.clk(gclk));
	jdff dff_A_Pb3eeLyY6_0(.dout(w_dff_A_jzOhX75Q6_0),.din(w_dff_A_Pb3eeLyY6_0),.clk(gclk));
	jdff dff_A_jzOhX75Q6_0(.dout(G634),.din(w_dff_A_jzOhX75Q6_0),.clk(gclk));
	jdff dff_A_OH6Zh5AK0_2(.dout(w_dff_A_N2KEKsvI8_0),.din(w_dff_A_OH6Zh5AK0_2),.clk(gclk));
	jdff dff_A_N2KEKsvI8_0(.dout(w_dff_A_MIMUbMn05_0),.din(w_dff_A_N2KEKsvI8_0),.clk(gclk));
	jdff dff_A_MIMUbMn05_0(.dout(w_dff_A_kxJNJilI8_0),.din(w_dff_A_MIMUbMn05_0),.clk(gclk));
	jdff dff_A_kxJNJilI8_0(.dout(w_dff_A_quTJmNWY2_0),.din(w_dff_A_kxJNJilI8_0),.clk(gclk));
	jdff dff_A_quTJmNWY2_0(.dout(w_dff_A_5hsWFbi39_0),.din(w_dff_A_quTJmNWY2_0),.clk(gclk));
	jdff dff_A_5hsWFbi39_0(.dout(w_dff_A_IfMazg3J2_0),.din(w_dff_A_5hsWFbi39_0),.clk(gclk));
	jdff dff_A_IfMazg3J2_0(.dout(w_dff_A_4ElZgcsd8_0),.din(w_dff_A_IfMazg3J2_0),.clk(gclk));
	jdff dff_A_4ElZgcsd8_0(.dout(w_dff_A_TEvPyqf50_0),.din(w_dff_A_4ElZgcsd8_0),.clk(gclk));
	jdff dff_A_TEvPyqf50_0(.dout(w_dff_A_pTX8Lrj61_0),.din(w_dff_A_TEvPyqf50_0),.clk(gclk));
	jdff dff_A_pTX8Lrj61_0(.dout(w_dff_A_0RrTwjxH4_0),.din(w_dff_A_pTX8Lrj61_0),.clk(gclk));
	jdff dff_A_0RrTwjxH4_0(.dout(w_dff_A_H0GP8xz22_0),.din(w_dff_A_0RrTwjxH4_0),.clk(gclk));
	jdff dff_A_H0GP8xz22_0(.dout(w_dff_A_ePVgpfCd9_0),.din(w_dff_A_H0GP8xz22_0),.clk(gclk));
	jdff dff_A_ePVgpfCd9_0(.dout(w_dff_A_eiHZuPqO9_0),.din(w_dff_A_ePVgpfCd9_0),.clk(gclk));
	jdff dff_A_eiHZuPqO9_0(.dout(w_dff_A_fnOeO3MS8_0),.din(w_dff_A_eiHZuPqO9_0),.clk(gclk));
	jdff dff_A_fnOeO3MS8_0(.dout(w_dff_A_L9fLYnFc6_0),.din(w_dff_A_fnOeO3MS8_0),.clk(gclk));
	jdff dff_A_L9fLYnFc6_0(.dout(w_dff_A_I2pDEBjq2_0),.din(w_dff_A_L9fLYnFc6_0),.clk(gclk));
	jdff dff_A_I2pDEBjq2_0(.dout(w_dff_A_yKFCD9rK7_0),.din(w_dff_A_I2pDEBjq2_0),.clk(gclk));
	jdff dff_A_yKFCD9rK7_0(.dout(w_dff_A_iUXtmZsD8_0),.din(w_dff_A_yKFCD9rK7_0),.clk(gclk));
	jdff dff_A_iUXtmZsD8_0(.dout(w_dff_A_z8lBlD5z9_0),.din(w_dff_A_iUXtmZsD8_0),.clk(gclk));
	jdff dff_A_z8lBlD5z9_0(.dout(w_dff_A_sfhm1jSA3_0),.din(w_dff_A_z8lBlD5z9_0),.clk(gclk));
	jdff dff_A_sfhm1jSA3_0(.dout(w_dff_A_tGGJOsZT3_0),.din(w_dff_A_sfhm1jSA3_0),.clk(gclk));
	jdff dff_A_tGGJOsZT3_0(.dout(w_dff_A_9DxYxE720_0),.din(w_dff_A_tGGJOsZT3_0),.clk(gclk));
	jdff dff_A_9DxYxE720_0(.dout(w_dff_A_T5KojIuZ8_0),.din(w_dff_A_9DxYxE720_0),.clk(gclk));
	jdff dff_A_T5KojIuZ8_0(.dout(w_dff_A_qK0KQUEf0_0),.din(w_dff_A_T5KojIuZ8_0),.clk(gclk));
	jdff dff_A_qK0KQUEf0_0(.dout(w_dff_A_C9JJiO8j7_0),.din(w_dff_A_qK0KQUEf0_0),.clk(gclk));
	jdff dff_A_C9JJiO8j7_0(.dout(G815),.din(w_dff_A_C9JJiO8j7_0),.clk(gclk));
	jdff dff_A_VhL8a7Hi2_2(.dout(w_dff_A_lmDI3Xpy0_0),.din(w_dff_A_VhL8a7Hi2_2),.clk(gclk));
	jdff dff_A_lmDI3Xpy0_0(.dout(w_dff_A_xmJYH3i71_0),.din(w_dff_A_lmDI3Xpy0_0),.clk(gclk));
	jdff dff_A_xmJYH3i71_0(.dout(w_dff_A_X4bah6s66_0),.din(w_dff_A_xmJYH3i71_0),.clk(gclk));
	jdff dff_A_X4bah6s66_0(.dout(w_dff_A_GG8xJHLR0_0),.din(w_dff_A_X4bah6s66_0),.clk(gclk));
	jdff dff_A_GG8xJHLR0_0(.dout(w_dff_A_Am0rr8ia6_0),.din(w_dff_A_GG8xJHLR0_0),.clk(gclk));
	jdff dff_A_Am0rr8ia6_0(.dout(w_dff_A_ziniP1yg0_0),.din(w_dff_A_Am0rr8ia6_0),.clk(gclk));
	jdff dff_A_ziniP1yg0_0(.dout(w_dff_A_0QqbKVWN2_0),.din(w_dff_A_ziniP1yg0_0),.clk(gclk));
	jdff dff_A_0QqbKVWN2_0(.dout(w_dff_A_qNiaCk008_0),.din(w_dff_A_0QqbKVWN2_0),.clk(gclk));
	jdff dff_A_qNiaCk008_0(.dout(w_dff_A_B8eWEI7M4_0),.din(w_dff_A_qNiaCk008_0),.clk(gclk));
	jdff dff_A_B8eWEI7M4_0(.dout(w_dff_A_Tmn3B10n1_0),.din(w_dff_A_B8eWEI7M4_0),.clk(gclk));
	jdff dff_A_Tmn3B10n1_0(.dout(w_dff_A_AdqvXExo8_0),.din(w_dff_A_Tmn3B10n1_0),.clk(gclk));
	jdff dff_A_AdqvXExo8_0(.dout(w_dff_A_IZIvzXdC9_0),.din(w_dff_A_AdqvXExo8_0),.clk(gclk));
	jdff dff_A_IZIvzXdC9_0(.dout(w_dff_A_I6cozvEI7_0),.din(w_dff_A_IZIvzXdC9_0),.clk(gclk));
	jdff dff_A_I6cozvEI7_0(.dout(w_dff_A_aVQFqvYm5_0),.din(w_dff_A_I6cozvEI7_0),.clk(gclk));
	jdff dff_A_aVQFqvYm5_0(.dout(w_dff_A_42X3hUSL4_0),.din(w_dff_A_aVQFqvYm5_0),.clk(gclk));
	jdff dff_A_42X3hUSL4_0(.dout(w_dff_A_mnsE0i5h7_0),.din(w_dff_A_42X3hUSL4_0),.clk(gclk));
	jdff dff_A_mnsE0i5h7_0(.dout(w_dff_A_08ZjJ4CS0_0),.din(w_dff_A_mnsE0i5h7_0),.clk(gclk));
	jdff dff_A_08ZjJ4CS0_0(.dout(w_dff_A_ddxzzvO39_0),.din(w_dff_A_08ZjJ4CS0_0),.clk(gclk));
	jdff dff_A_ddxzzvO39_0(.dout(w_dff_A_w7YCfT897_0),.din(w_dff_A_ddxzzvO39_0),.clk(gclk));
	jdff dff_A_w7YCfT897_0(.dout(w_dff_A_JZ6UktA11_0),.din(w_dff_A_w7YCfT897_0),.clk(gclk));
	jdff dff_A_JZ6UktA11_0(.dout(w_dff_A_2J2pDMNO7_0),.din(w_dff_A_JZ6UktA11_0),.clk(gclk));
	jdff dff_A_2J2pDMNO7_0(.dout(w_dff_A_pQCXdcjM9_0),.din(w_dff_A_2J2pDMNO7_0),.clk(gclk));
	jdff dff_A_pQCXdcjM9_0(.dout(w_dff_A_os0MY85t2_0),.din(w_dff_A_pQCXdcjM9_0),.clk(gclk));
	jdff dff_A_os0MY85t2_0(.dout(w_dff_A_FxIb3VD82_0),.din(w_dff_A_os0MY85t2_0),.clk(gclk));
	jdff dff_A_FxIb3VD82_0(.dout(w_dff_A_DBAqT5CM5_0),.din(w_dff_A_FxIb3VD82_0),.clk(gclk));
	jdff dff_A_DBAqT5CM5_0(.dout(G845),.din(w_dff_A_DBAqT5CM5_0),.clk(gclk));
	jdff dff_A_bVnKpyJe2_1(.dout(w_dff_A_sNMes2xq3_0),.din(w_dff_A_bVnKpyJe2_1),.clk(gclk));
	jdff dff_A_sNMes2xq3_0(.dout(w_dff_A_gcwI9eLp5_0),.din(w_dff_A_sNMes2xq3_0),.clk(gclk));
	jdff dff_A_gcwI9eLp5_0(.dout(w_dff_A_DhLlgaSN6_0),.din(w_dff_A_gcwI9eLp5_0),.clk(gclk));
	jdff dff_A_DhLlgaSN6_0(.dout(w_dff_A_j0Lu4hRI0_0),.din(w_dff_A_DhLlgaSN6_0),.clk(gclk));
	jdff dff_A_j0Lu4hRI0_0(.dout(w_dff_A_xbCIpbPw8_0),.din(w_dff_A_j0Lu4hRI0_0),.clk(gclk));
	jdff dff_A_xbCIpbPw8_0(.dout(w_dff_A_VVOeO6qV9_0),.din(w_dff_A_xbCIpbPw8_0),.clk(gclk));
	jdff dff_A_VVOeO6qV9_0(.dout(w_dff_A_AMPNKxgC4_0),.din(w_dff_A_VVOeO6qV9_0),.clk(gclk));
	jdff dff_A_AMPNKxgC4_0(.dout(w_dff_A_5vUqcwrY2_0),.din(w_dff_A_AMPNKxgC4_0),.clk(gclk));
	jdff dff_A_5vUqcwrY2_0(.dout(w_dff_A_X2FJdbXX2_0),.din(w_dff_A_5vUqcwrY2_0),.clk(gclk));
	jdff dff_A_X2FJdbXX2_0(.dout(w_dff_A_J4CyiKpG1_0),.din(w_dff_A_X2FJdbXX2_0),.clk(gclk));
	jdff dff_A_J4CyiKpG1_0(.dout(w_dff_A_0GBY2gXW5_0),.din(w_dff_A_J4CyiKpG1_0),.clk(gclk));
	jdff dff_A_0GBY2gXW5_0(.dout(w_dff_A_LZiyji1t2_0),.din(w_dff_A_0GBY2gXW5_0),.clk(gclk));
	jdff dff_A_LZiyji1t2_0(.dout(w_dff_A_WG8yMshn7_0),.din(w_dff_A_LZiyji1t2_0),.clk(gclk));
	jdff dff_A_WG8yMshn7_0(.dout(w_dff_A_kpnAInKq8_0),.din(w_dff_A_WG8yMshn7_0),.clk(gclk));
	jdff dff_A_kpnAInKq8_0(.dout(w_dff_A_fb6p92pT0_0),.din(w_dff_A_kpnAInKq8_0),.clk(gclk));
	jdff dff_A_fb6p92pT0_0(.dout(w_dff_A_9CbOgmPp7_0),.din(w_dff_A_fb6p92pT0_0),.clk(gclk));
	jdff dff_A_9CbOgmPp7_0(.dout(w_dff_A_H7bL1R8s8_0),.din(w_dff_A_9CbOgmPp7_0),.clk(gclk));
	jdff dff_A_H7bL1R8s8_0(.dout(w_dff_A_FS1QuHnS5_0),.din(w_dff_A_H7bL1R8s8_0),.clk(gclk));
	jdff dff_A_FS1QuHnS5_0(.dout(w_dff_A_wYxCKXSC5_0),.din(w_dff_A_FS1QuHnS5_0),.clk(gclk));
	jdff dff_A_wYxCKXSC5_0(.dout(w_dff_A_ByRSjIIX1_0),.din(w_dff_A_wYxCKXSC5_0),.clk(gclk));
	jdff dff_A_ByRSjIIX1_0(.dout(w_dff_A_mdZ8LgLo8_0),.din(w_dff_A_ByRSjIIX1_0),.clk(gclk));
	jdff dff_A_mdZ8LgLo8_0(.dout(w_dff_A_1o1MSxgE0_0),.din(w_dff_A_mdZ8LgLo8_0),.clk(gclk));
	jdff dff_A_1o1MSxgE0_0(.dout(w_dff_A_xgltJCvw2_0),.din(w_dff_A_1o1MSxgE0_0),.clk(gclk));
	jdff dff_A_xgltJCvw2_0(.dout(w_dff_A_rcFxavpJ4_0),.din(w_dff_A_xgltJCvw2_0),.clk(gclk));
	jdff dff_A_rcFxavpJ4_0(.dout(w_dff_A_pbKwJ33I5_0),.din(w_dff_A_rcFxavpJ4_0),.clk(gclk));
	jdff dff_A_pbKwJ33I5_0(.dout(G847),.din(w_dff_A_pbKwJ33I5_0),.clk(gclk));
	jdff dff_A_89syVh4x7_1(.dout(w_dff_A_1uvbwhDw4_0),.din(w_dff_A_89syVh4x7_1),.clk(gclk));
	jdff dff_A_1uvbwhDw4_0(.dout(w_dff_A_38iV7vhd5_0),.din(w_dff_A_1uvbwhDw4_0),.clk(gclk));
	jdff dff_A_38iV7vhd5_0(.dout(w_dff_A_NLaJEFPh8_0),.din(w_dff_A_38iV7vhd5_0),.clk(gclk));
	jdff dff_A_NLaJEFPh8_0(.dout(w_dff_A_0pXMRSfR2_0),.din(w_dff_A_NLaJEFPh8_0),.clk(gclk));
	jdff dff_A_0pXMRSfR2_0(.dout(w_dff_A_s5o6lvEh9_0),.din(w_dff_A_0pXMRSfR2_0),.clk(gclk));
	jdff dff_A_s5o6lvEh9_0(.dout(w_dff_A_NATKnATn3_0),.din(w_dff_A_s5o6lvEh9_0),.clk(gclk));
	jdff dff_A_NATKnATn3_0(.dout(w_dff_A_MHlUP8Er2_0),.din(w_dff_A_NATKnATn3_0),.clk(gclk));
	jdff dff_A_MHlUP8Er2_0(.dout(w_dff_A_kS1BFII74_0),.din(w_dff_A_MHlUP8Er2_0),.clk(gclk));
	jdff dff_A_kS1BFII74_0(.dout(w_dff_A_J3185Slh8_0),.din(w_dff_A_kS1BFII74_0),.clk(gclk));
	jdff dff_A_J3185Slh8_0(.dout(w_dff_A_K0N75OsA6_0),.din(w_dff_A_J3185Slh8_0),.clk(gclk));
	jdff dff_A_K0N75OsA6_0(.dout(w_dff_A_EYyHNL9i5_0),.din(w_dff_A_K0N75OsA6_0),.clk(gclk));
	jdff dff_A_EYyHNL9i5_0(.dout(w_dff_A_i1k7lZIg6_0),.din(w_dff_A_EYyHNL9i5_0),.clk(gclk));
	jdff dff_A_i1k7lZIg6_0(.dout(w_dff_A_EPBu9JjM2_0),.din(w_dff_A_i1k7lZIg6_0),.clk(gclk));
	jdff dff_A_EPBu9JjM2_0(.dout(w_dff_A_bakxyuKq1_0),.din(w_dff_A_EPBu9JjM2_0),.clk(gclk));
	jdff dff_A_bakxyuKq1_0(.dout(w_dff_A_xJfYTcoW5_0),.din(w_dff_A_bakxyuKq1_0),.clk(gclk));
	jdff dff_A_xJfYTcoW5_0(.dout(w_dff_A_Ti61som40_0),.din(w_dff_A_xJfYTcoW5_0),.clk(gclk));
	jdff dff_A_Ti61som40_0(.dout(w_dff_A_OrvTgNDg2_0),.din(w_dff_A_Ti61som40_0),.clk(gclk));
	jdff dff_A_OrvTgNDg2_0(.dout(w_dff_A_W8zT1ZWT0_0),.din(w_dff_A_OrvTgNDg2_0),.clk(gclk));
	jdff dff_A_W8zT1ZWT0_0(.dout(w_dff_A_r0tORCi30_0),.din(w_dff_A_W8zT1ZWT0_0),.clk(gclk));
	jdff dff_A_r0tORCi30_0(.dout(w_dff_A_5ieYbjB38_0),.din(w_dff_A_r0tORCi30_0),.clk(gclk));
	jdff dff_A_5ieYbjB38_0(.dout(w_dff_A_yjf03Y5Q5_0),.din(w_dff_A_5ieYbjB38_0),.clk(gclk));
	jdff dff_A_yjf03Y5Q5_0(.dout(w_dff_A_7AIEKMpy6_0),.din(w_dff_A_yjf03Y5Q5_0),.clk(gclk));
	jdff dff_A_7AIEKMpy6_0(.dout(w_dff_A_kl2cAbLN1_0),.din(w_dff_A_7AIEKMpy6_0),.clk(gclk));
	jdff dff_A_kl2cAbLN1_0(.dout(w_dff_A_cIFvpTN56_0),.din(w_dff_A_kl2cAbLN1_0),.clk(gclk));
	jdff dff_A_cIFvpTN56_0(.dout(w_dff_A_RB8vrvXz7_0),.din(w_dff_A_cIFvpTN56_0),.clk(gclk));
	jdff dff_A_RB8vrvXz7_0(.dout(w_dff_A_TrrcuXLq7_0),.din(w_dff_A_RB8vrvXz7_0),.clk(gclk));
	jdff dff_A_TrrcuXLq7_0(.dout(w_dff_A_gx8JxHGs8_0),.din(w_dff_A_TrrcuXLq7_0),.clk(gclk));
	jdff dff_A_gx8JxHGs8_0(.dout(G926),.din(w_dff_A_gx8JxHGs8_0),.clk(gclk));
	jdff dff_A_Djl8qfsF2_1(.dout(w_dff_A_uHwNA8uP4_0),.din(w_dff_A_Djl8qfsF2_1),.clk(gclk));
	jdff dff_A_uHwNA8uP4_0(.dout(w_dff_A_DdyKhmnY6_0),.din(w_dff_A_uHwNA8uP4_0),.clk(gclk));
	jdff dff_A_DdyKhmnY6_0(.dout(w_dff_A_o8HuD9hM3_0),.din(w_dff_A_DdyKhmnY6_0),.clk(gclk));
	jdff dff_A_o8HuD9hM3_0(.dout(w_dff_A_FTFAQXl47_0),.din(w_dff_A_o8HuD9hM3_0),.clk(gclk));
	jdff dff_A_FTFAQXl47_0(.dout(w_dff_A_cbB2SOQa6_0),.din(w_dff_A_FTFAQXl47_0),.clk(gclk));
	jdff dff_A_cbB2SOQa6_0(.dout(w_dff_A_ptTRaTXg6_0),.din(w_dff_A_cbB2SOQa6_0),.clk(gclk));
	jdff dff_A_ptTRaTXg6_0(.dout(w_dff_A_f3TOpIVJ4_0),.din(w_dff_A_ptTRaTXg6_0),.clk(gclk));
	jdff dff_A_f3TOpIVJ4_0(.dout(w_dff_A_NDvHUJmN6_0),.din(w_dff_A_f3TOpIVJ4_0),.clk(gclk));
	jdff dff_A_NDvHUJmN6_0(.dout(w_dff_A_ydJy0zww6_0),.din(w_dff_A_NDvHUJmN6_0),.clk(gclk));
	jdff dff_A_ydJy0zww6_0(.dout(w_dff_A_OrkTTjHp0_0),.din(w_dff_A_ydJy0zww6_0),.clk(gclk));
	jdff dff_A_OrkTTjHp0_0(.dout(w_dff_A_pbXFo8wI0_0),.din(w_dff_A_OrkTTjHp0_0),.clk(gclk));
	jdff dff_A_pbXFo8wI0_0(.dout(w_dff_A_FAcIb2ZA9_0),.din(w_dff_A_pbXFo8wI0_0),.clk(gclk));
	jdff dff_A_FAcIb2ZA9_0(.dout(w_dff_A_DuVQZ8Zp5_0),.din(w_dff_A_FAcIb2ZA9_0),.clk(gclk));
	jdff dff_A_DuVQZ8Zp5_0(.dout(w_dff_A_qCYSapFb8_0),.din(w_dff_A_DuVQZ8Zp5_0),.clk(gclk));
	jdff dff_A_qCYSapFb8_0(.dout(w_dff_A_Ce3eQfKm3_0),.din(w_dff_A_qCYSapFb8_0),.clk(gclk));
	jdff dff_A_Ce3eQfKm3_0(.dout(w_dff_A_5yqLeVTs9_0),.din(w_dff_A_Ce3eQfKm3_0),.clk(gclk));
	jdff dff_A_5yqLeVTs9_0(.dout(w_dff_A_X4Dd6mIJ0_0),.din(w_dff_A_5yqLeVTs9_0),.clk(gclk));
	jdff dff_A_X4Dd6mIJ0_0(.dout(w_dff_A_Xsg4b4qM0_0),.din(w_dff_A_X4Dd6mIJ0_0),.clk(gclk));
	jdff dff_A_Xsg4b4qM0_0(.dout(w_dff_A_y0Q2HcCC9_0),.din(w_dff_A_Xsg4b4qM0_0),.clk(gclk));
	jdff dff_A_y0Q2HcCC9_0(.dout(w_dff_A_vswiE9ur9_0),.din(w_dff_A_y0Q2HcCC9_0),.clk(gclk));
	jdff dff_A_vswiE9ur9_0(.dout(w_dff_A_mkWQvSHp5_0),.din(w_dff_A_vswiE9ur9_0),.clk(gclk));
	jdff dff_A_mkWQvSHp5_0(.dout(w_dff_A_1ysOx7qy7_0),.din(w_dff_A_mkWQvSHp5_0),.clk(gclk));
	jdff dff_A_1ysOx7qy7_0(.dout(w_dff_A_iYMq4zli7_0),.din(w_dff_A_1ysOx7qy7_0),.clk(gclk));
	jdff dff_A_iYMq4zli7_0(.dout(w_dff_A_V9FvTsy90_0),.din(w_dff_A_iYMq4zli7_0),.clk(gclk));
	jdff dff_A_V9FvTsy90_0(.dout(w_dff_A_78Xgc0hA2_0),.din(w_dff_A_V9FvTsy90_0),.clk(gclk));
	jdff dff_A_78Xgc0hA2_0(.dout(w_dff_A_bK7AZ3K36_0),.din(w_dff_A_78Xgc0hA2_0),.clk(gclk));
	jdff dff_A_bK7AZ3K36_0(.dout(w_dff_A_EDnwvmV64_0),.din(w_dff_A_bK7AZ3K36_0),.clk(gclk));
	jdff dff_A_EDnwvmV64_0(.dout(G923),.din(w_dff_A_EDnwvmV64_0),.clk(gclk));
	jdff dff_A_yjWZdSrI8_1(.dout(w_dff_A_ms8Ogwvj0_0),.din(w_dff_A_yjWZdSrI8_1),.clk(gclk));
	jdff dff_A_ms8Ogwvj0_0(.dout(w_dff_A_83jEZO4Q4_0),.din(w_dff_A_ms8Ogwvj0_0),.clk(gclk));
	jdff dff_A_83jEZO4Q4_0(.dout(w_dff_A_simhCqkU3_0),.din(w_dff_A_83jEZO4Q4_0),.clk(gclk));
	jdff dff_A_simhCqkU3_0(.dout(w_dff_A_z7IpTcvV0_0),.din(w_dff_A_simhCqkU3_0),.clk(gclk));
	jdff dff_A_z7IpTcvV0_0(.dout(w_dff_A_YLrRpXNn3_0),.din(w_dff_A_z7IpTcvV0_0),.clk(gclk));
	jdff dff_A_YLrRpXNn3_0(.dout(w_dff_A_9MUSjGPC7_0),.din(w_dff_A_YLrRpXNn3_0),.clk(gclk));
	jdff dff_A_9MUSjGPC7_0(.dout(w_dff_A_2V62cTiC1_0),.din(w_dff_A_9MUSjGPC7_0),.clk(gclk));
	jdff dff_A_2V62cTiC1_0(.dout(w_dff_A_P2XWxGm99_0),.din(w_dff_A_2V62cTiC1_0),.clk(gclk));
	jdff dff_A_P2XWxGm99_0(.dout(w_dff_A_fCJR7X7t6_0),.din(w_dff_A_P2XWxGm99_0),.clk(gclk));
	jdff dff_A_fCJR7X7t6_0(.dout(w_dff_A_OrE62XP96_0),.din(w_dff_A_fCJR7X7t6_0),.clk(gclk));
	jdff dff_A_OrE62XP96_0(.dout(w_dff_A_YbgL1t2N4_0),.din(w_dff_A_OrE62XP96_0),.clk(gclk));
	jdff dff_A_YbgL1t2N4_0(.dout(w_dff_A_IKaVbsgN3_0),.din(w_dff_A_YbgL1t2N4_0),.clk(gclk));
	jdff dff_A_IKaVbsgN3_0(.dout(w_dff_A_XaXi0i4v6_0),.din(w_dff_A_IKaVbsgN3_0),.clk(gclk));
	jdff dff_A_XaXi0i4v6_0(.dout(w_dff_A_dPhcw7DX7_0),.din(w_dff_A_XaXi0i4v6_0),.clk(gclk));
	jdff dff_A_dPhcw7DX7_0(.dout(w_dff_A_5SrttqCL2_0),.din(w_dff_A_dPhcw7DX7_0),.clk(gclk));
	jdff dff_A_5SrttqCL2_0(.dout(w_dff_A_Dmy6ELkT9_0),.din(w_dff_A_5SrttqCL2_0),.clk(gclk));
	jdff dff_A_Dmy6ELkT9_0(.dout(w_dff_A_fO7YP6j59_0),.din(w_dff_A_Dmy6ELkT9_0),.clk(gclk));
	jdff dff_A_fO7YP6j59_0(.dout(w_dff_A_zbgsl6pe4_0),.din(w_dff_A_fO7YP6j59_0),.clk(gclk));
	jdff dff_A_zbgsl6pe4_0(.dout(w_dff_A_KAM6vUaN3_0),.din(w_dff_A_zbgsl6pe4_0),.clk(gclk));
	jdff dff_A_KAM6vUaN3_0(.dout(w_dff_A_2DWTLcxA1_0),.din(w_dff_A_KAM6vUaN3_0),.clk(gclk));
	jdff dff_A_2DWTLcxA1_0(.dout(w_dff_A_Rg5ZErBR2_0),.din(w_dff_A_2DWTLcxA1_0),.clk(gclk));
	jdff dff_A_Rg5ZErBR2_0(.dout(w_dff_A_CvJIUbm24_0),.din(w_dff_A_Rg5ZErBR2_0),.clk(gclk));
	jdff dff_A_CvJIUbm24_0(.dout(w_dff_A_ay0qS0rU1_0),.din(w_dff_A_CvJIUbm24_0),.clk(gclk));
	jdff dff_A_ay0qS0rU1_0(.dout(w_dff_A_NS0MKecF1_0),.din(w_dff_A_ay0qS0rU1_0),.clk(gclk));
	jdff dff_A_NS0MKecF1_0(.dout(w_dff_A_Y3YPvJS25_0),.din(w_dff_A_NS0MKecF1_0),.clk(gclk));
	jdff dff_A_Y3YPvJS25_0(.dout(w_dff_A_6vBVRovC8_0),.din(w_dff_A_Y3YPvJS25_0),.clk(gclk));
	jdff dff_A_6vBVRovC8_0(.dout(w_dff_A_IY6SMMSa5_0),.din(w_dff_A_6vBVRovC8_0),.clk(gclk));
	jdff dff_A_IY6SMMSa5_0(.dout(G921),.din(w_dff_A_IY6SMMSa5_0),.clk(gclk));
	jdff dff_A_qN7P6uT37_1(.dout(w_dff_A_TGX3X0lo1_0),.din(w_dff_A_qN7P6uT37_1),.clk(gclk));
	jdff dff_A_TGX3X0lo1_0(.dout(w_dff_A_aTTNi7kC6_0),.din(w_dff_A_TGX3X0lo1_0),.clk(gclk));
	jdff dff_A_aTTNi7kC6_0(.dout(w_dff_A_yoUPXft99_0),.din(w_dff_A_aTTNi7kC6_0),.clk(gclk));
	jdff dff_A_yoUPXft99_0(.dout(w_dff_A_k5TYflGb8_0),.din(w_dff_A_yoUPXft99_0),.clk(gclk));
	jdff dff_A_k5TYflGb8_0(.dout(w_dff_A_GGgCHdBl1_0),.din(w_dff_A_k5TYflGb8_0),.clk(gclk));
	jdff dff_A_GGgCHdBl1_0(.dout(w_dff_A_p9ZBD0Ij4_0),.din(w_dff_A_GGgCHdBl1_0),.clk(gclk));
	jdff dff_A_p9ZBD0Ij4_0(.dout(w_dff_A_qWaDCNBU8_0),.din(w_dff_A_p9ZBD0Ij4_0),.clk(gclk));
	jdff dff_A_qWaDCNBU8_0(.dout(w_dff_A_LAUJW3rj5_0),.din(w_dff_A_qWaDCNBU8_0),.clk(gclk));
	jdff dff_A_LAUJW3rj5_0(.dout(w_dff_A_spjQNx6D8_0),.din(w_dff_A_LAUJW3rj5_0),.clk(gclk));
	jdff dff_A_spjQNx6D8_0(.dout(w_dff_A_newntnSS8_0),.din(w_dff_A_spjQNx6D8_0),.clk(gclk));
	jdff dff_A_newntnSS8_0(.dout(w_dff_A_R6nLkOSR2_0),.din(w_dff_A_newntnSS8_0),.clk(gclk));
	jdff dff_A_R6nLkOSR2_0(.dout(w_dff_A_350XQWaM0_0),.din(w_dff_A_R6nLkOSR2_0),.clk(gclk));
	jdff dff_A_350XQWaM0_0(.dout(w_dff_A_LFiiiwHC7_0),.din(w_dff_A_350XQWaM0_0),.clk(gclk));
	jdff dff_A_LFiiiwHC7_0(.dout(w_dff_A_kqEd3cFC5_0),.din(w_dff_A_LFiiiwHC7_0),.clk(gclk));
	jdff dff_A_kqEd3cFC5_0(.dout(w_dff_A_VAHWTEKF6_0),.din(w_dff_A_kqEd3cFC5_0),.clk(gclk));
	jdff dff_A_VAHWTEKF6_0(.dout(w_dff_A_CCjeenWr3_0),.din(w_dff_A_VAHWTEKF6_0),.clk(gclk));
	jdff dff_A_CCjeenWr3_0(.dout(w_dff_A_yPlqqW1x7_0),.din(w_dff_A_CCjeenWr3_0),.clk(gclk));
	jdff dff_A_yPlqqW1x7_0(.dout(w_dff_A_vEnxif705_0),.din(w_dff_A_yPlqqW1x7_0),.clk(gclk));
	jdff dff_A_vEnxif705_0(.dout(w_dff_A_jMyqDxfU2_0),.din(w_dff_A_vEnxif705_0),.clk(gclk));
	jdff dff_A_jMyqDxfU2_0(.dout(w_dff_A_nq7ZcTK26_0),.din(w_dff_A_jMyqDxfU2_0),.clk(gclk));
	jdff dff_A_nq7ZcTK26_0(.dout(w_dff_A_oSAov2VM7_0),.din(w_dff_A_nq7ZcTK26_0),.clk(gclk));
	jdff dff_A_oSAov2VM7_0(.dout(w_dff_A_FLyvadE44_0),.din(w_dff_A_oSAov2VM7_0),.clk(gclk));
	jdff dff_A_FLyvadE44_0(.dout(w_dff_A_g1VTKuQY6_0),.din(w_dff_A_FLyvadE44_0),.clk(gclk));
	jdff dff_A_g1VTKuQY6_0(.dout(w_dff_A_7Xl50UlW7_0),.din(w_dff_A_g1VTKuQY6_0),.clk(gclk));
	jdff dff_A_7Xl50UlW7_0(.dout(w_dff_A_NPqMWFeW8_0),.din(w_dff_A_7Xl50UlW7_0),.clk(gclk));
	jdff dff_A_NPqMWFeW8_0(.dout(w_dff_A_xPevfiNR4_0),.din(w_dff_A_NPqMWFeW8_0),.clk(gclk));
	jdff dff_A_xPevfiNR4_0(.dout(w_dff_A_QSkIBtqJ1_0),.din(w_dff_A_xPevfiNR4_0),.clk(gclk));
	jdff dff_A_QSkIBtqJ1_0(.dout(G892),.din(w_dff_A_QSkIBtqJ1_0),.clk(gclk));
	jdff dff_A_PSsXJ15W0_1(.dout(w_dff_A_Ug2BgSzk9_0),.din(w_dff_A_PSsXJ15W0_1),.clk(gclk));
	jdff dff_A_Ug2BgSzk9_0(.dout(w_dff_A_BBu9EIOM9_0),.din(w_dff_A_Ug2BgSzk9_0),.clk(gclk));
	jdff dff_A_BBu9EIOM9_0(.dout(w_dff_A_ZMFkfpbE7_0),.din(w_dff_A_BBu9EIOM9_0),.clk(gclk));
	jdff dff_A_ZMFkfpbE7_0(.dout(w_dff_A_qI1Ph0Ky6_0),.din(w_dff_A_ZMFkfpbE7_0),.clk(gclk));
	jdff dff_A_qI1Ph0Ky6_0(.dout(w_dff_A_qDukArh07_0),.din(w_dff_A_qI1Ph0Ky6_0),.clk(gclk));
	jdff dff_A_qDukArh07_0(.dout(w_dff_A_9U8MbDxN4_0),.din(w_dff_A_qDukArh07_0),.clk(gclk));
	jdff dff_A_9U8MbDxN4_0(.dout(w_dff_A_895ieqmJ4_0),.din(w_dff_A_9U8MbDxN4_0),.clk(gclk));
	jdff dff_A_895ieqmJ4_0(.dout(w_dff_A_uryfAE3j1_0),.din(w_dff_A_895ieqmJ4_0),.clk(gclk));
	jdff dff_A_uryfAE3j1_0(.dout(w_dff_A_NpFoXssA1_0),.din(w_dff_A_uryfAE3j1_0),.clk(gclk));
	jdff dff_A_NpFoXssA1_0(.dout(w_dff_A_HJGLyjP44_0),.din(w_dff_A_NpFoXssA1_0),.clk(gclk));
	jdff dff_A_HJGLyjP44_0(.dout(w_dff_A_OzFBeN273_0),.din(w_dff_A_HJGLyjP44_0),.clk(gclk));
	jdff dff_A_OzFBeN273_0(.dout(w_dff_A_MC5kieKL0_0),.din(w_dff_A_OzFBeN273_0),.clk(gclk));
	jdff dff_A_MC5kieKL0_0(.dout(w_dff_A_Q58p9H0s4_0),.din(w_dff_A_MC5kieKL0_0),.clk(gclk));
	jdff dff_A_Q58p9H0s4_0(.dout(w_dff_A_agzX51c82_0),.din(w_dff_A_Q58p9H0s4_0),.clk(gclk));
	jdff dff_A_agzX51c82_0(.dout(w_dff_A_RLXXXLze6_0),.din(w_dff_A_agzX51c82_0),.clk(gclk));
	jdff dff_A_RLXXXLze6_0(.dout(w_dff_A_5EE25wH68_0),.din(w_dff_A_RLXXXLze6_0),.clk(gclk));
	jdff dff_A_5EE25wH68_0(.dout(w_dff_A_ylk7N2wh6_0),.din(w_dff_A_5EE25wH68_0),.clk(gclk));
	jdff dff_A_ylk7N2wh6_0(.dout(w_dff_A_pTINlDbJ7_0),.din(w_dff_A_ylk7N2wh6_0),.clk(gclk));
	jdff dff_A_pTINlDbJ7_0(.dout(w_dff_A_tAIuwWch8_0),.din(w_dff_A_pTINlDbJ7_0),.clk(gclk));
	jdff dff_A_tAIuwWch8_0(.dout(w_dff_A_Y2dLup4P3_0),.din(w_dff_A_tAIuwWch8_0),.clk(gclk));
	jdff dff_A_Y2dLup4P3_0(.dout(w_dff_A_C8dXU2ed3_0),.din(w_dff_A_Y2dLup4P3_0),.clk(gclk));
	jdff dff_A_C8dXU2ed3_0(.dout(w_dff_A_aZdJrW847_0),.din(w_dff_A_C8dXU2ed3_0),.clk(gclk));
	jdff dff_A_aZdJrW847_0(.dout(w_dff_A_EHyLl6oL0_0),.din(w_dff_A_aZdJrW847_0),.clk(gclk));
	jdff dff_A_EHyLl6oL0_0(.dout(w_dff_A_wdukhdF37_0),.din(w_dff_A_EHyLl6oL0_0),.clk(gclk));
	jdff dff_A_wdukhdF37_0(.dout(w_dff_A_jR4NHXAp0_0),.din(w_dff_A_wdukhdF37_0),.clk(gclk));
	jdff dff_A_jR4NHXAp0_0(.dout(w_dff_A_6466RNsy0_0),.din(w_dff_A_jR4NHXAp0_0),.clk(gclk));
	jdff dff_A_6466RNsy0_0(.dout(w_dff_A_05582kQs1_0),.din(w_dff_A_6466RNsy0_0),.clk(gclk));
	jdff dff_A_05582kQs1_0(.dout(G887),.din(w_dff_A_05582kQs1_0),.clk(gclk));
	jdff dff_A_qEhQ7mZt4_1(.dout(w_dff_A_VYiq91BK4_0),.din(w_dff_A_qEhQ7mZt4_1),.clk(gclk));
	jdff dff_A_VYiq91BK4_0(.dout(w_dff_A_Id3VjDEr4_0),.din(w_dff_A_VYiq91BK4_0),.clk(gclk));
	jdff dff_A_Id3VjDEr4_0(.dout(w_dff_A_r7VL3lMI1_0),.din(w_dff_A_Id3VjDEr4_0),.clk(gclk));
	jdff dff_A_r7VL3lMI1_0(.dout(w_dff_A_oQmAHtLq9_0),.din(w_dff_A_r7VL3lMI1_0),.clk(gclk));
	jdff dff_A_oQmAHtLq9_0(.dout(w_dff_A_6nHge9MI2_0),.din(w_dff_A_oQmAHtLq9_0),.clk(gclk));
	jdff dff_A_6nHge9MI2_0(.dout(w_dff_A_4tdLart07_0),.din(w_dff_A_6nHge9MI2_0),.clk(gclk));
	jdff dff_A_4tdLart07_0(.dout(w_dff_A_bMz4h6uN1_0),.din(w_dff_A_4tdLart07_0),.clk(gclk));
	jdff dff_A_bMz4h6uN1_0(.dout(w_dff_A_sb8KNqAg8_0),.din(w_dff_A_bMz4h6uN1_0),.clk(gclk));
	jdff dff_A_sb8KNqAg8_0(.dout(w_dff_A_cyFhwre65_0),.din(w_dff_A_sb8KNqAg8_0),.clk(gclk));
	jdff dff_A_cyFhwre65_0(.dout(w_dff_A_yVQM5J398_0),.din(w_dff_A_cyFhwre65_0),.clk(gclk));
	jdff dff_A_yVQM5J398_0(.dout(w_dff_A_COp3oKn32_0),.din(w_dff_A_yVQM5J398_0),.clk(gclk));
	jdff dff_A_COp3oKn32_0(.dout(w_dff_A_CXY1px9e1_0),.din(w_dff_A_COp3oKn32_0),.clk(gclk));
	jdff dff_A_CXY1px9e1_0(.dout(w_dff_A_PegklGeu8_0),.din(w_dff_A_CXY1px9e1_0),.clk(gclk));
	jdff dff_A_PegklGeu8_0(.dout(w_dff_A_kXDuMQTE0_0),.din(w_dff_A_PegklGeu8_0),.clk(gclk));
	jdff dff_A_kXDuMQTE0_0(.dout(w_dff_A_w6Oqor3X4_0),.din(w_dff_A_kXDuMQTE0_0),.clk(gclk));
	jdff dff_A_w6Oqor3X4_0(.dout(w_dff_A_ualuFDsY8_0),.din(w_dff_A_w6Oqor3X4_0),.clk(gclk));
	jdff dff_A_ualuFDsY8_0(.dout(w_dff_A_ObytXB1X9_0),.din(w_dff_A_ualuFDsY8_0),.clk(gclk));
	jdff dff_A_ObytXB1X9_0(.dout(w_dff_A_ACsoLH0A7_0),.din(w_dff_A_ObytXB1X9_0),.clk(gclk));
	jdff dff_A_ACsoLH0A7_0(.dout(w_dff_A_tAq5Jsva7_0),.din(w_dff_A_ACsoLH0A7_0),.clk(gclk));
	jdff dff_A_tAq5Jsva7_0(.dout(w_dff_A_bysvXtS30_0),.din(w_dff_A_tAq5Jsva7_0),.clk(gclk));
	jdff dff_A_bysvXtS30_0(.dout(w_dff_A_9JVwg8Y61_0),.din(w_dff_A_bysvXtS30_0),.clk(gclk));
	jdff dff_A_9JVwg8Y61_0(.dout(w_dff_A_M5BuBABE1_0),.din(w_dff_A_9JVwg8Y61_0),.clk(gclk));
	jdff dff_A_M5BuBABE1_0(.dout(w_dff_A_tjDV1YYa0_0),.din(w_dff_A_M5BuBABE1_0),.clk(gclk));
	jdff dff_A_tjDV1YYa0_0(.dout(w_dff_A_iolEBKst5_0),.din(w_dff_A_tjDV1YYa0_0),.clk(gclk));
	jdff dff_A_iolEBKst5_0(.dout(w_dff_A_pJdVrf4L0_0),.din(w_dff_A_iolEBKst5_0),.clk(gclk));
	jdff dff_A_pJdVrf4L0_0(.dout(w_dff_A_du2bENbP6_0),.din(w_dff_A_pJdVrf4L0_0),.clk(gclk));
	jdff dff_A_du2bENbP6_0(.dout(G606),.din(w_dff_A_du2bENbP6_0),.clk(gclk));
	jdff dff_A_oqcc29e21_2(.dout(w_dff_A_Yqimw46x8_0),.din(w_dff_A_oqcc29e21_2),.clk(gclk));
	jdff dff_A_Yqimw46x8_0(.dout(w_dff_A_t5B54jkc1_0),.din(w_dff_A_Yqimw46x8_0),.clk(gclk));
	jdff dff_A_t5B54jkc1_0(.dout(w_dff_A_u9HB3Ruf2_0),.din(w_dff_A_t5B54jkc1_0),.clk(gclk));
	jdff dff_A_u9HB3Ruf2_0(.dout(w_dff_A_v32F4mKa2_0),.din(w_dff_A_u9HB3Ruf2_0),.clk(gclk));
	jdff dff_A_v32F4mKa2_0(.dout(w_dff_A_QVtkJ8h12_0),.din(w_dff_A_v32F4mKa2_0),.clk(gclk));
	jdff dff_A_QVtkJ8h12_0(.dout(w_dff_A_mas9Mo8i8_0),.din(w_dff_A_QVtkJ8h12_0),.clk(gclk));
	jdff dff_A_mas9Mo8i8_0(.dout(w_dff_A_1QJItDNs2_0),.din(w_dff_A_mas9Mo8i8_0),.clk(gclk));
	jdff dff_A_1QJItDNs2_0(.dout(w_dff_A_U6lWPRgU2_0),.din(w_dff_A_1QJItDNs2_0),.clk(gclk));
	jdff dff_A_U6lWPRgU2_0(.dout(w_dff_A_5PelUQCX2_0),.din(w_dff_A_U6lWPRgU2_0),.clk(gclk));
	jdff dff_A_5PelUQCX2_0(.dout(w_dff_A_0AEkfg3q1_0),.din(w_dff_A_5PelUQCX2_0),.clk(gclk));
	jdff dff_A_0AEkfg3q1_0(.dout(w_dff_A_xTN3EjxV8_0),.din(w_dff_A_0AEkfg3q1_0),.clk(gclk));
	jdff dff_A_xTN3EjxV8_0(.dout(w_dff_A_ZOHblKiH6_0),.din(w_dff_A_xTN3EjxV8_0),.clk(gclk));
	jdff dff_A_ZOHblKiH6_0(.dout(w_dff_A_0kqwJ3S26_0),.din(w_dff_A_ZOHblKiH6_0),.clk(gclk));
	jdff dff_A_0kqwJ3S26_0(.dout(w_dff_A_Q3AYVYiL7_0),.din(w_dff_A_0kqwJ3S26_0),.clk(gclk));
	jdff dff_A_Q3AYVYiL7_0(.dout(w_dff_A_XOSBnFRT1_0),.din(w_dff_A_Q3AYVYiL7_0),.clk(gclk));
	jdff dff_A_XOSBnFRT1_0(.dout(w_dff_A_c9tAdXBx3_0),.din(w_dff_A_XOSBnFRT1_0),.clk(gclk));
	jdff dff_A_c9tAdXBx3_0(.dout(w_dff_A_WnqdlrYJ9_0),.din(w_dff_A_c9tAdXBx3_0),.clk(gclk));
	jdff dff_A_WnqdlrYJ9_0(.dout(w_dff_A_fdPuh2TP5_0),.din(w_dff_A_WnqdlrYJ9_0),.clk(gclk));
	jdff dff_A_fdPuh2TP5_0(.dout(w_dff_A_O0VEYkna8_0),.din(w_dff_A_fdPuh2TP5_0),.clk(gclk));
	jdff dff_A_O0VEYkna8_0(.dout(w_dff_A_4Zq9FWId0_0),.din(w_dff_A_O0VEYkna8_0),.clk(gclk));
	jdff dff_A_4Zq9FWId0_0(.dout(w_dff_A_juj8VRgE0_0),.din(w_dff_A_4Zq9FWId0_0),.clk(gclk));
	jdff dff_A_juj8VRgE0_0(.dout(w_dff_A_MvIbOGo68_0),.din(w_dff_A_juj8VRgE0_0),.clk(gclk));
	jdff dff_A_MvIbOGo68_0(.dout(w_dff_A_WDNapyno5_0),.din(w_dff_A_MvIbOGo68_0),.clk(gclk));
	jdff dff_A_WDNapyno5_0(.dout(w_dff_A_XJ2fTZCO6_0),.din(w_dff_A_WDNapyno5_0),.clk(gclk));
	jdff dff_A_XJ2fTZCO6_0(.dout(G656),.din(w_dff_A_XJ2fTZCO6_0),.clk(gclk));
	jdff dff_A_CwjD3V1R2_2(.dout(w_dff_A_DS5EGWgg1_0),.din(w_dff_A_CwjD3V1R2_2),.clk(gclk));
	jdff dff_A_DS5EGWgg1_0(.dout(w_dff_A_GFwzC6XV8_0),.din(w_dff_A_DS5EGWgg1_0),.clk(gclk));
	jdff dff_A_GFwzC6XV8_0(.dout(w_dff_A_aPHB6ZpI6_0),.din(w_dff_A_GFwzC6XV8_0),.clk(gclk));
	jdff dff_A_aPHB6ZpI6_0(.dout(w_dff_A_rF5evuqK8_0),.din(w_dff_A_aPHB6ZpI6_0),.clk(gclk));
	jdff dff_A_rF5evuqK8_0(.dout(w_dff_A_NdI6BpDJ8_0),.din(w_dff_A_rF5evuqK8_0),.clk(gclk));
	jdff dff_A_NdI6BpDJ8_0(.dout(w_dff_A_MDggdN5e4_0),.din(w_dff_A_NdI6BpDJ8_0),.clk(gclk));
	jdff dff_A_MDggdN5e4_0(.dout(w_dff_A_TPIh1QrY3_0),.din(w_dff_A_MDggdN5e4_0),.clk(gclk));
	jdff dff_A_TPIh1QrY3_0(.dout(w_dff_A_Gkcfn5RK4_0),.din(w_dff_A_TPIh1QrY3_0),.clk(gclk));
	jdff dff_A_Gkcfn5RK4_0(.dout(w_dff_A_D9V4I86y1_0),.din(w_dff_A_Gkcfn5RK4_0),.clk(gclk));
	jdff dff_A_D9V4I86y1_0(.dout(w_dff_A_BJIcDcHs5_0),.din(w_dff_A_D9V4I86y1_0),.clk(gclk));
	jdff dff_A_BJIcDcHs5_0(.dout(w_dff_A_ttLtsfud7_0),.din(w_dff_A_BJIcDcHs5_0),.clk(gclk));
	jdff dff_A_ttLtsfud7_0(.dout(w_dff_A_0UDfAeTo2_0),.din(w_dff_A_ttLtsfud7_0),.clk(gclk));
	jdff dff_A_0UDfAeTo2_0(.dout(w_dff_A_XbXavE0S9_0),.din(w_dff_A_0UDfAeTo2_0),.clk(gclk));
	jdff dff_A_XbXavE0S9_0(.dout(w_dff_A_TSVMNdIC4_0),.din(w_dff_A_XbXavE0S9_0),.clk(gclk));
	jdff dff_A_TSVMNdIC4_0(.dout(w_dff_A_CI6NKT2n6_0),.din(w_dff_A_TSVMNdIC4_0),.clk(gclk));
	jdff dff_A_CI6NKT2n6_0(.dout(w_dff_A_0kPwUYkb7_0),.din(w_dff_A_CI6NKT2n6_0),.clk(gclk));
	jdff dff_A_0kPwUYkb7_0(.dout(w_dff_A_Ww5aTARl9_0),.din(w_dff_A_0kPwUYkb7_0),.clk(gclk));
	jdff dff_A_Ww5aTARl9_0(.dout(w_dff_A_ye4Yh7GD0_0),.din(w_dff_A_Ww5aTARl9_0),.clk(gclk));
	jdff dff_A_ye4Yh7GD0_0(.dout(w_dff_A_5w0oXtj81_0),.din(w_dff_A_ye4Yh7GD0_0),.clk(gclk));
	jdff dff_A_5w0oXtj81_0(.dout(w_dff_A_WHCClyld9_0),.din(w_dff_A_5w0oXtj81_0),.clk(gclk));
	jdff dff_A_WHCClyld9_0(.dout(w_dff_A_7VwZvmNA6_0),.din(w_dff_A_WHCClyld9_0),.clk(gclk));
	jdff dff_A_7VwZvmNA6_0(.dout(w_dff_A_Ka95FIKu8_0),.din(w_dff_A_7VwZvmNA6_0),.clk(gclk));
	jdff dff_A_Ka95FIKu8_0(.dout(w_dff_A_5GR9xbYu7_0),.din(w_dff_A_Ka95FIKu8_0),.clk(gclk));
	jdff dff_A_5GR9xbYu7_0(.dout(w_dff_A_jqBiUilE3_0),.din(w_dff_A_5GR9xbYu7_0),.clk(gclk));
	jdff dff_A_jqBiUilE3_0(.dout(w_dff_A_y50DGCjn9_0),.din(w_dff_A_jqBiUilE3_0),.clk(gclk));
	jdff dff_A_y50DGCjn9_0(.dout(G809),.din(w_dff_A_y50DGCjn9_0),.clk(gclk));
	jdff dff_A_Jr8Poux14_1(.dout(w_dff_A_F8bSBTaH3_0),.din(w_dff_A_Jr8Poux14_1),.clk(gclk));
	jdff dff_A_F8bSBTaH3_0(.dout(w_dff_A_o3dv0q6f5_0),.din(w_dff_A_F8bSBTaH3_0),.clk(gclk));
	jdff dff_A_o3dv0q6f5_0(.dout(w_dff_A_cx2ZOHkk1_0),.din(w_dff_A_o3dv0q6f5_0),.clk(gclk));
	jdff dff_A_cx2ZOHkk1_0(.dout(w_dff_A_qZhtsyp25_0),.din(w_dff_A_cx2ZOHkk1_0),.clk(gclk));
	jdff dff_A_qZhtsyp25_0(.dout(w_dff_A_oAEqgSbh1_0),.din(w_dff_A_qZhtsyp25_0),.clk(gclk));
	jdff dff_A_oAEqgSbh1_0(.dout(w_dff_A_dKSe6A4v2_0),.din(w_dff_A_oAEqgSbh1_0),.clk(gclk));
	jdff dff_A_dKSe6A4v2_0(.dout(w_dff_A_AfOoE4qC9_0),.din(w_dff_A_dKSe6A4v2_0),.clk(gclk));
	jdff dff_A_AfOoE4qC9_0(.dout(w_dff_A_S5GWcIcB5_0),.din(w_dff_A_AfOoE4qC9_0),.clk(gclk));
	jdff dff_A_S5GWcIcB5_0(.dout(w_dff_A_h9cYaEAZ0_0),.din(w_dff_A_S5GWcIcB5_0),.clk(gclk));
	jdff dff_A_h9cYaEAZ0_0(.dout(w_dff_A_4Zxeq7Up4_0),.din(w_dff_A_h9cYaEAZ0_0),.clk(gclk));
	jdff dff_A_4Zxeq7Up4_0(.dout(w_dff_A_eH7dVURb0_0),.din(w_dff_A_4Zxeq7Up4_0),.clk(gclk));
	jdff dff_A_eH7dVURb0_0(.dout(w_dff_A_8HFsyjQs2_0),.din(w_dff_A_eH7dVURb0_0),.clk(gclk));
	jdff dff_A_8HFsyjQs2_0(.dout(w_dff_A_RIZedcK41_0),.din(w_dff_A_8HFsyjQs2_0),.clk(gclk));
	jdff dff_A_RIZedcK41_0(.dout(w_dff_A_1anNgPut1_0),.din(w_dff_A_RIZedcK41_0),.clk(gclk));
	jdff dff_A_1anNgPut1_0(.dout(w_dff_A_tpO0IO2S8_0),.din(w_dff_A_1anNgPut1_0),.clk(gclk));
	jdff dff_A_tpO0IO2S8_0(.dout(w_dff_A_GHavWRYA0_0),.din(w_dff_A_tpO0IO2S8_0),.clk(gclk));
	jdff dff_A_GHavWRYA0_0(.dout(w_dff_A_b16INpQS9_0),.din(w_dff_A_GHavWRYA0_0),.clk(gclk));
	jdff dff_A_b16INpQS9_0(.dout(w_dff_A_pcgwPvLI0_0),.din(w_dff_A_b16INpQS9_0),.clk(gclk));
	jdff dff_A_pcgwPvLI0_0(.dout(w_dff_A_5UoSz9aN1_0),.din(w_dff_A_pcgwPvLI0_0),.clk(gclk));
	jdff dff_A_5UoSz9aN1_0(.dout(w_dff_A_1teGdIhy7_0),.din(w_dff_A_5UoSz9aN1_0),.clk(gclk));
	jdff dff_A_1teGdIhy7_0(.dout(w_dff_A_8z1PV1PL9_0),.din(w_dff_A_1teGdIhy7_0),.clk(gclk));
	jdff dff_A_8z1PV1PL9_0(.dout(w_dff_A_E7ikNyBW4_0),.din(w_dff_A_8z1PV1PL9_0),.clk(gclk));
	jdff dff_A_E7ikNyBW4_0(.dout(w_dff_A_Hd6RFwKU0_0),.din(w_dff_A_E7ikNyBW4_0),.clk(gclk));
	jdff dff_A_Hd6RFwKU0_0(.dout(w_dff_A_GZxFGRy99_0),.din(w_dff_A_Hd6RFwKU0_0),.clk(gclk));
	jdff dff_A_GZxFGRy99_0(.dout(w_dff_A_XYlrOvK51_0),.din(w_dff_A_GZxFGRy99_0),.clk(gclk));
	jdff dff_A_XYlrOvK51_0(.dout(w_dff_A_7l2rTrJ02_0),.din(w_dff_A_XYlrOvK51_0),.clk(gclk));
	jdff dff_A_7l2rTrJ02_0(.dout(w_dff_A_0pxxqC283_0),.din(w_dff_A_7l2rTrJ02_0),.clk(gclk));
	jdff dff_A_0pxxqC283_0(.dout(G993),.din(w_dff_A_0pxxqC283_0),.clk(gclk));
	jdff dff_A_5qB1Wwgm5_1(.dout(w_dff_A_QiFcPK1d2_0),.din(w_dff_A_5qB1Wwgm5_1),.clk(gclk));
	jdff dff_A_QiFcPK1d2_0(.dout(w_dff_A_KcNW2Nji3_0),.din(w_dff_A_QiFcPK1d2_0),.clk(gclk));
	jdff dff_A_KcNW2Nji3_0(.dout(w_dff_A_mY0YDJSm5_0),.din(w_dff_A_KcNW2Nji3_0),.clk(gclk));
	jdff dff_A_mY0YDJSm5_0(.dout(w_dff_A_Pai1qV8N2_0),.din(w_dff_A_mY0YDJSm5_0),.clk(gclk));
	jdff dff_A_Pai1qV8N2_0(.dout(w_dff_A_YECSUc3l7_0),.din(w_dff_A_Pai1qV8N2_0),.clk(gclk));
	jdff dff_A_YECSUc3l7_0(.dout(w_dff_A_NiFIqM7g0_0),.din(w_dff_A_YECSUc3l7_0),.clk(gclk));
	jdff dff_A_NiFIqM7g0_0(.dout(w_dff_A_aTPMHJjz4_0),.din(w_dff_A_NiFIqM7g0_0),.clk(gclk));
	jdff dff_A_aTPMHJjz4_0(.dout(w_dff_A_vZP94e7T5_0),.din(w_dff_A_aTPMHJjz4_0),.clk(gclk));
	jdff dff_A_vZP94e7T5_0(.dout(w_dff_A_c5hovwXG6_0),.din(w_dff_A_vZP94e7T5_0),.clk(gclk));
	jdff dff_A_c5hovwXG6_0(.dout(w_dff_A_LTrnyG2e6_0),.din(w_dff_A_c5hovwXG6_0),.clk(gclk));
	jdff dff_A_LTrnyG2e6_0(.dout(w_dff_A_pJ4DMt4b8_0),.din(w_dff_A_LTrnyG2e6_0),.clk(gclk));
	jdff dff_A_pJ4DMt4b8_0(.dout(w_dff_A_my9kqod26_0),.din(w_dff_A_pJ4DMt4b8_0),.clk(gclk));
	jdff dff_A_my9kqod26_0(.dout(w_dff_A_z4148bWO6_0),.din(w_dff_A_my9kqod26_0),.clk(gclk));
	jdff dff_A_z4148bWO6_0(.dout(w_dff_A_oebE02oE6_0),.din(w_dff_A_z4148bWO6_0),.clk(gclk));
	jdff dff_A_oebE02oE6_0(.dout(w_dff_A_sidP7CfN8_0),.din(w_dff_A_oebE02oE6_0),.clk(gclk));
	jdff dff_A_sidP7CfN8_0(.dout(w_dff_A_5QARFbBz1_0),.din(w_dff_A_sidP7CfN8_0),.clk(gclk));
	jdff dff_A_5QARFbBz1_0(.dout(w_dff_A_qM7MkbBq3_0),.din(w_dff_A_5QARFbBz1_0),.clk(gclk));
	jdff dff_A_qM7MkbBq3_0(.dout(w_dff_A_9hJpMHN12_0),.din(w_dff_A_qM7MkbBq3_0),.clk(gclk));
	jdff dff_A_9hJpMHN12_0(.dout(w_dff_A_PHmR1R8v3_0),.din(w_dff_A_9hJpMHN12_0),.clk(gclk));
	jdff dff_A_PHmR1R8v3_0(.dout(w_dff_A_xE7gTKhy9_0),.din(w_dff_A_PHmR1R8v3_0),.clk(gclk));
	jdff dff_A_xE7gTKhy9_0(.dout(w_dff_A_MdGHM0hg4_0),.din(w_dff_A_xE7gTKhy9_0),.clk(gclk));
	jdff dff_A_MdGHM0hg4_0(.dout(w_dff_A_BW4Rz7Wx0_0),.din(w_dff_A_MdGHM0hg4_0),.clk(gclk));
	jdff dff_A_BW4Rz7Wx0_0(.dout(w_dff_A_iPTIjNHM8_0),.din(w_dff_A_BW4Rz7Wx0_0),.clk(gclk));
	jdff dff_A_iPTIjNHM8_0(.dout(w_dff_A_gaaf1wZa8_0),.din(w_dff_A_iPTIjNHM8_0),.clk(gclk));
	jdff dff_A_gaaf1wZa8_0(.dout(w_dff_A_77sej2RW2_0),.din(w_dff_A_gaaf1wZa8_0),.clk(gclk));
	jdff dff_A_77sej2RW2_0(.dout(w_dff_A_Wjmm5db44_0),.din(w_dff_A_77sej2RW2_0),.clk(gclk));
	jdff dff_A_Wjmm5db44_0(.dout(w_dff_A_Dyi2xxG79_0),.din(w_dff_A_Wjmm5db44_0),.clk(gclk));
	jdff dff_A_Dyi2xxG79_0(.dout(G978),.din(w_dff_A_Dyi2xxG79_0),.clk(gclk));
	jdff dff_A_6PibwFQP0_1(.dout(w_dff_A_NAr0nbiS0_0),.din(w_dff_A_6PibwFQP0_1),.clk(gclk));
	jdff dff_A_NAr0nbiS0_0(.dout(w_dff_A_7vcpugSA5_0),.din(w_dff_A_NAr0nbiS0_0),.clk(gclk));
	jdff dff_A_7vcpugSA5_0(.dout(w_dff_A_PMuoWas64_0),.din(w_dff_A_7vcpugSA5_0),.clk(gclk));
	jdff dff_A_PMuoWas64_0(.dout(w_dff_A_9mjG3KIa4_0),.din(w_dff_A_PMuoWas64_0),.clk(gclk));
	jdff dff_A_9mjG3KIa4_0(.dout(w_dff_A_WGFi5evy5_0),.din(w_dff_A_9mjG3KIa4_0),.clk(gclk));
	jdff dff_A_WGFi5evy5_0(.dout(w_dff_A_raik2fwo0_0),.din(w_dff_A_WGFi5evy5_0),.clk(gclk));
	jdff dff_A_raik2fwo0_0(.dout(w_dff_A_G1ZFgysv0_0),.din(w_dff_A_raik2fwo0_0),.clk(gclk));
	jdff dff_A_G1ZFgysv0_0(.dout(w_dff_A_yk23dkXe0_0),.din(w_dff_A_G1ZFgysv0_0),.clk(gclk));
	jdff dff_A_yk23dkXe0_0(.dout(w_dff_A_oxQ6hHQa2_0),.din(w_dff_A_yk23dkXe0_0),.clk(gclk));
	jdff dff_A_oxQ6hHQa2_0(.dout(w_dff_A_NM7hZlOk6_0),.din(w_dff_A_oxQ6hHQa2_0),.clk(gclk));
	jdff dff_A_NM7hZlOk6_0(.dout(w_dff_A_RURjXBRE1_0),.din(w_dff_A_NM7hZlOk6_0),.clk(gclk));
	jdff dff_A_RURjXBRE1_0(.dout(w_dff_A_NEPMgGSQ6_0),.din(w_dff_A_RURjXBRE1_0),.clk(gclk));
	jdff dff_A_NEPMgGSQ6_0(.dout(w_dff_A_D3rzod2Y8_0),.din(w_dff_A_NEPMgGSQ6_0),.clk(gclk));
	jdff dff_A_D3rzod2Y8_0(.dout(w_dff_A_CHiL6nAq2_0),.din(w_dff_A_D3rzod2Y8_0),.clk(gclk));
	jdff dff_A_CHiL6nAq2_0(.dout(w_dff_A_fVNyg9GQ7_0),.din(w_dff_A_CHiL6nAq2_0),.clk(gclk));
	jdff dff_A_fVNyg9GQ7_0(.dout(w_dff_A_HV1qglns7_0),.din(w_dff_A_fVNyg9GQ7_0),.clk(gclk));
	jdff dff_A_HV1qglns7_0(.dout(w_dff_A_gQdVYz3g4_0),.din(w_dff_A_HV1qglns7_0),.clk(gclk));
	jdff dff_A_gQdVYz3g4_0(.dout(w_dff_A_GGZ1bkbJ2_0),.din(w_dff_A_gQdVYz3g4_0),.clk(gclk));
	jdff dff_A_GGZ1bkbJ2_0(.dout(w_dff_A_48b1dG4j4_0),.din(w_dff_A_GGZ1bkbJ2_0),.clk(gclk));
	jdff dff_A_48b1dG4j4_0(.dout(w_dff_A_NX0Mbq458_0),.din(w_dff_A_48b1dG4j4_0),.clk(gclk));
	jdff dff_A_NX0Mbq458_0(.dout(w_dff_A_lBLOVfDg7_0),.din(w_dff_A_NX0Mbq458_0),.clk(gclk));
	jdff dff_A_lBLOVfDg7_0(.dout(w_dff_A_LqqgSHtT6_0),.din(w_dff_A_lBLOVfDg7_0),.clk(gclk));
	jdff dff_A_LqqgSHtT6_0(.dout(w_dff_A_qjoztbQ95_0),.din(w_dff_A_LqqgSHtT6_0),.clk(gclk));
	jdff dff_A_qjoztbQ95_0(.dout(w_dff_A_x7PphQwi2_0),.din(w_dff_A_qjoztbQ95_0),.clk(gclk));
	jdff dff_A_x7PphQwi2_0(.dout(w_dff_A_jpb0fABL6_0),.din(w_dff_A_x7PphQwi2_0),.clk(gclk));
	jdff dff_A_jpb0fABL6_0(.dout(w_dff_A_5gaDKYYD1_0),.din(w_dff_A_jpb0fABL6_0),.clk(gclk));
	jdff dff_A_5gaDKYYD1_0(.dout(w_dff_A_KRlEvn7Q5_0),.din(w_dff_A_5gaDKYYD1_0),.clk(gclk));
	jdff dff_A_KRlEvn7Q5_0(.dout(G949),.din(w_dff_A_KRlEvn7Q5_0),.clk(gclk));
	jdff dff_A_qMdRBAAX3_1(.dout(w_dff_A_PbAy1E7j9_0),.din(w_dff_A_qMdRBAAX3_1),.clk(gclk));
	jdff dff_A_PbAy1E7j9_0(.dout(w_dff_A_VP7Yuk048_0),.din(w_dff_A_PbAy1E7j9_0),.clk(gclk));
	jdff dff_A_VP7Yuk048_0(.dout(w_dff_A_9JWn5wmt9_0),.din(w_dff_A_VP7Yuk048_0),.clk(gclk));
	jdff dff_A_9JWn5wmt9_0(.dout(w_dff_A_OytqGTUF2_0),.din(w_dff_A_9JWn5wmt9_0),.clk(gclk));
	jdff dff_A_OytqGTUF2_0(.dout(w_dff_A_iYOkjqJI0_0),.din(w_dff_A_OytqGTUF2_0),.clk(gclk));
	jdff dff_A_iYOkjqJI0_0(.dout(w_dff_A_ngq5qNrN9_0),.din(w_dff_A_iYOkjqJI0_0),.clk(gclk));
	jdff dff_A_ngq5qNrN9_0(.dout(w_dff_A_mdTBWsOS5_0),.din(w_dff_A_ngq5qNrN9_0),.clk(gclk));
	jdff dff_A_mdTBWsOS5_0(.dout(w_dff_A_hNF3nORq8_0),.din(w_dff_A_mdTBWsOS5_0),.clk(gclk));
	jdff dff_A_hNF3nORq8_0(.dout(w_dff_A_c9pQJQ6f5_0),.din(w_dff_A_hNF3nORq8_0),.clk(gclk));
	jdff dff_A_c9pQJQ6f5_0(.dout(w_dff_A_CxOK3SWi6_0),.din(w_dff_A_c9pQJQ6f5_0),.clk(gclk));
	jdff dff_A_CxOK3SWi6_0(.dout(w_dff_A_V1rAConY6_0),.din(w_dff_A_CxOK3SWi6_0),.clk(gclk));
	jdff dff_A_V1rAConY6_0(.dout(w_dff_A_Rb6VoArY3_0),.din(w_dff_A_V1rAConY6_0),.clk(gclk));
	jdff dff_A_Rb6VoArY3_0(.dout(w_dff_A_TyodUl2B5_0),.din(w_dff_A_Rb6VoArY3_0),.clk(gclk));
	jdff dff_A_TyodUl2B5_0(.dout(w_dff_A_kwjCYwuU4_0),.din(w_dff_A_TyodUl2B5_0),.clk(gclk));
	jdff dff_A_kwjCYwuU4_0(.dout(w_dff_A_Gxen4T7b6_0),.din(w_dff_A_kwjCYwuU4_0),.clk(gclk));
	jdff dff_A_Gxen4T7b6_0(.dout(w_dff_A_QkFChoAe0_0),.din(w_dff_A_Gxen4T7b6_0),.clk(gclk));
	jdff dff_A_QkFChoAe0_0(.dout(w_dff_A_PrRUgtQT1_0),.din(w_dff_A_QkFChoAe0_0),.clk(gclk));
	jdff dff_A_PrRUgtQT1_0(.dout(w_dff_A_jflovsba6_0),.din(w_dff_A_PrRUgtQT1_0),.clk(gclk));
	jdff dff_A_jflovsba6_0(.dout(w_dff_A_TOa7h5G44_0),.din(w_dff_A_jflovsba6_0),.clk(gclk));
	jdff dff_A_TOa7h5G44_0(.dout(w_dff_A_oG70jydl1_0),.din(w_dff_A_TOa7h5G44_0),.clk(gclk));
	jdff dff_A_oG70jydl1_0(.dout(w_dff_A_SECA2VR75_0),.din(w_dff_A_oG70jydl1_0),.clk(gclk));
	jdff dff_A_SECA2VR75_0(.dout(w_dff_A_bQp0DKEC5_0),.din(w_dff_A_SECA2VR75_0),.clk(gclk));
	jdff dff_A_bQp0DKEC5_0(.dout(w_dff_A_HPPl2pon6_0),.din(w_dff_A_bQp0DKEC5_0),.clk(gclk));
	jdff dff_A_HPPl2pon6_0(.dout(w_dff_A_4c3i4UQN2_0),.din(w_dff_A_HPPl2pon6_0),.clk(gclk));
	jdff dff_A_4c3i4UQN2_0(.dout(w_dff_A_KWNXN5WD7_0),.din(w_dff_A_4c3i4UQN2_0),.clk(gclk));
	jdff dff_A_KWNXN5WD7_0(.dout(w_dff_A_WeWgc0Ks3_0),.din(w_dff_A_KWNXN5WD7_0),.clk(gclk));
	jdff dff_A_WeWgc0Ks3_0(.dout(w_dff_A_cBoqA3M19_0),.din(w_dff_A_WeWgc0Ks3_0),.clk(gclk));
	jdff dff_A_cBoqA3M19_0(.dout(G939),.din(w_dff_A_cBoqA3M19_0),.clk(gclk));
	jdff dff_A_Zz1Li1Zx3_1(.dout(w_dff_A_cCR9KJWS9_0),.din(w_dff_A_Zz1Li1Zx3_1),.clk(gclk));
	jdff dff_A_cCR9KJWS9_0(.dout(w_dff_A_IqOjfl9g1_0),.din(w_dff_A_cCR9KJWS9_0),.clk(gclk));
	jdff dff_A_IqOjfl9g1_0(.dout(w_dff_A_pK0WH2ev0_0),.din(w_dff_A_IqOjfl9g1_0),.clk(gclk));
	jdff dff_A_pK0WH2ev0_0(.dout(w_dff_A_DUvRX0o68_0),.din(w_dff_A_pK0WH2ev0_0),.clk(gclk));
	jdff dff_A_DUvRX0o68_0(.dout(w_dff_A_0ADnCMfh8_0),.din(w_dff_A_DUvRX0o68_0),.clk(gclk));
	jdff dff_A_0ADnCMfh8_0(.dout(w_dff_A_3RaMxQkp4_0),.din(w_dff_A_0ADnCMfh8_0),.clk(gclk));
	jdff dff_A_3RaMxQkp4_0(.dout(w_dff_A_ArgoCyNb1_0),.din(w_dff_A_3RaMxQkp4_0),.clk(gclk));
	jdff dff_A_ArgoCyNb1_0(.dout(w_dff_A_HDwlHXnf4_0),.din(w_dff_A_ArgoCyNb1_0),.clk(gclk));
	jdff dff_A_HDwlHXnf4_0(.dout(w_dff_A_Z6I7FigU6_0),.din(w_dff_A_HDwlHXnf4_0),.clk(gclk));
	jdff dff_A_Z6I7FigU6_0(.dout(w_dff_A_pWvkJEzi8_0),.din(w_dff_A_Z6I7FigU6_0),.clk(gclk));
	jdff dff_A_pWvkJEzi8_0(.dout(w_dff_A_BdFtLRAU6_0),.din(w_dff_A_pWvkJEzi8_0),.clk(gclk));
	jdff dff_A_BdFtLRAU6_0(.dout(w_dff_A_eNYZQxEt5_0),.din(w_dff_A_BdFtLRAU6_0),.clk(gclk));
	jdff dff_A_eNYZQxEt5_0(.dout(w_dff_A_IZnJYaqC9_0),.din(w_dff_A_eNYZQxEt5_0),.clk(gclk));
	jdff dff_A_IZnJYaqC9_0(.dout(w_dff_A_ICqH0h6V2_0),.din(w_dff_A_IZnJYaqC9_0),.clk(gclk));
	jdff dff_A_ICqH0h6V2_0(.dout(w_dff_A_FwWfb5WH2_0),.din(w_dff_A_ICqH0h6V2_0),.clk(gclk));
	jdff dff_A_FwWfb5WH2_0(.dout(w_dff_A_8yEdFNwL8_0),.din(w_dff_A_FwWfb5WH2_0),.clk(gclk));
	jdff dff_A_8yEdFNwL8_0(.dout(w_dff_A_Z4A7ykqo3_0),.din(w_dff_A_8yEdFNwL8_0),.clk(gclk));
	jdff dff_A_Z4A7ykqo3_0(.dout(w_dff_A_KEw0JQQO1_0),.din(w_dff_A_Z4A7ykqo3_0),.clk(gclk));
	jdff dff_A_KEw0JQQO1_0(.dout(w_dff_A_vyWxBQaY6_0),.din(w_dff_A_KEw0JQQO1_0),.clk(gclk));
	jdff dff_A_vyWxBQaY6_0(.dout(w_dff_A_6FoVjSK19_0),.din(w_dff_A_vyWxBQaY6_0),.clk(gclk));
	jdff dff_A_6FoVjSK19_0(.dout(w_dff_A_dSgNEWpI3_0),.din(w_dff_A_6FoVjSK19_0),.clk(gclk));
	jdff dff_A_dSgNEWpI3_0(.dout(w_dff_A_66KyrKr42_0),.din(w_dff_A_dSgNEWpI3_0),.clk(gclk));
	jdff dff_A_66KyrKr42_0(.dout(w_dff_A_tz0oaOhV2_0),.din(w_dff_A_66KyrKr42_0),.clk(gclk));
	jdff dff_A_tz0oaOhV2_0(.dout(w_dff_A_UZ1tRybF8_0),.din(w_dff_A_tz0oaOhV2_0),.clk(gclk));
	jdff dff_A_UZ1tRybF8_0(.dout(w_dff_A_0bfURztX9_0),.din(w_dff_A_UZ1tRybF8_0),.clk(gclk));
	jdff dff_A_0bfURztX9_0(.dout(w_dff_A_WsJHWIyI8_0),.din(w_dff_A_0bfURztX9_0),.clk(gclk));
	jdff dff_A_WsJHWIyI8_0(.dout(w_dff_A_sVE4msgX6_0),.din(w_dff_A_WsJHWIyI8_0),.clk(gclk));
	jdff dff_A_sVE4msgX6_0(.dout(G889),.din(w_dff_A_sVE4msgX6_0),.clk(gclk));
	jdff dff_A_AujOhDyB6_1(.dout(w_dff_A_TaYAKsDG3_0),.din(w_dff_A_AujOhDyB6_1),.clk(gclk));
	jdff dff_A_TaYAKsDG3_0(.dout(w_dff_A_CvY2WmNa8_0),.din(w_dff_A_TaYAKsDG3_0),.clk(gclk));
	jdff dff_A_CvY2WmNa8_0(.dout(w_dff_A_IWtdi0Qj8_0),.din(w_dff_A_CvY2WmNa8_0),.clk(gclk));
	jdff dff_A_IWtdi0Qj8_0(.dout(w_dff_A_NELiMDpj0_0),.din(w_dff_A_IWtdi0Qj8_0),.clk(gclk));
	jdff dff_A_NELiMDpj0_0(.dout(w_dff_A_ZPHDB9T20_0),.din(w_dff_A_NELiMDpj0_0),.clk(gclk));
	jdff dff_A_ZPHDB9T20_0(.dout(w_dff_A_4DPSxF180_0),.din(w_dff_A_ZPHDB9T20_0),.clk(gclk));
	jdff dff_A_4DPSxF180_0(.dout(w_dff_A_1gPRKQvg4_0),.din(w_dff_A_4DPSxF180_0),.clk(gclk));
	jdff dff_A_1gPRKQvg4_0(.dout(w_dff_A_w3qxbbPi0_0),.din(w_dff_A_1gPRKQvg4_0),.clk(gclk));
	jdff dff_A_w3qxbbPi0_0(.dout(w_dff_A_RDwaEHnY7_0),.din(w_dff_A_w3qxbbPi0_0),.clk(gclk));
	jdff dff_A_RDwaEHnY7_0(.dout(w_dff_A_6eApylkC4_0),.din(w_dff_A_RDwaEHnY7_0),.clk(gclk));
	jdff dff_A_6eApylkC4_0(.dout(w_dff_A_J2IOZki74_0),.din(w_dff_A_6eApylkC4_0),.clk(gclk));
	jdff dff_A_J2IOZki74_0(.dout(w_dff_A_V4V9GpGs7_0),.din(w_dff_A_J2IOZki74_0),.clk(gclk));
	jdff dff_A_V4V9GpGs7_0(.dout(w_dff_A_8OiKwdFj1_0),.din(w_dff_A_V4V9GpGs7_0),.clk(gclk));
	jdff dff_A_8OiKwdFj1_0(.dout(w_dff_A_LPupaLFz1_0),.din(w_dff_A_8OiKwdFj1_0),.clk(gclk));
	jdff dff_A_LPupaLFz1_0(.dout(w_dff_A_TikIZPQr3_0),.din(w_dff_A_LPupaLFz1_0),.clk(gclk));
	jdff dff_A_TikIZPQr3_0(.dout(w_dff_A_HCWY5qnu1_0),.din(w_dff_A_TikIZPQr3_0),.clk(gclk));
	jdff dff_A_HCWY5qnu1_0(.dout(w_dff_A_8ixV8VVE1_0),.din(w_dff_A_HCWY5qnu1_0),.clk(gclk));
	jdff dff_A_8ixV8VVE1_0(.dout(w_dff_A_jBRbCC2h8_0),.din(w_dff_A_8ixV8VVE1_0),.clk(gclk));
	jdff dff_A_jBRbCC2h8_0(.dout(w_dff_A_iB7WVXaT5_0),.din(w_dff_A_jBRbCC2h8_0),.clk(gclk));
	jdff dff_A_iB7WVXaT5_0(.dout(w_dff_A_f0K8BVYe9_0),.din(w_dff_A_iB7WVXaT5_0),.clk(gclk));
	jdff dff_A_f0K8BVYe9_0(.dout(w_dff_A_SKy5dBIu3_0),.din(w_dff_A_f0K8BVYe9_0),.clk(gclk));
	jdff dff_A_SKy5dBIu3_0(.dout(w_dff_A_wcQfNUWc9_0),.din(w_dff_A_SKy5dBIu3_0),.clk(gclk));
	jdff dff_A_wcQfNUWc9_0(.dout(w_dff_A_xv2Ejnxx7_0),.din(w_dff_A_wcQfNUWc9_0),.clk(gclk));
	jdff dff_A_xv2Ejnxx7_0(.dout(w_dff_A_qbXzBuoM0_0),.din(w_dff_A_xv2Ejnxx7_0),.clk(gclk));
	jdff dff_A_qbXzBuoM0_0(.dout(w_dff_A_HiDj1bum9_0),.din(w_dff_A_qbXzBuoM0_0),.clk(gclk));
	jdff dff_A_HiDj1bum9_0(.dout(w_dff_A_IQzfYfcm2_0),.din(w_dff_A_HiDj1bum9_0),.clk(gclk));
	jdff dff_A_IQzfYfcm2_0(.dout(G593),.din(w_dff_A_IQzfYfcm2_0),.clk(gclk));
	jdff dff_A_pWrd5YD36_2(.dout(w_dff_A_jOtAdkIz7_0),.din(w_dff_A_pWrd5YD36_2),.clk(gclk));
	jdff dff_A_jOtAdkIz7_0(.dout(w_dff_A_PfJ98FuH0_0),.din(w_dff_A_jOtAdkIz7_0),.clk(gclk));
	jdff dff_A_PfJ98FuH0_0(.dout(w_dff_A_mgKKCepW8_0),.din(w_dff_A_PfJ98FuH0_0),.clk(gclk));
	jdff dff_A_mgKKCepW8_0(.dout(w_dff_A_Jzpmppu41_0),.din(w_dff_A_mgKKCepW8_0),.clk(gclk));
	jdff dff_A_Jzpmppu41_0(.dout(w_dff_A_ph7FrcEQ1_0),.din(w_dff_A_Jzpmppu41_0),.clk(gclk));
	jdff dff_A_ph7FrcEQ1_0(.dout(w_dff_A_k9shR9gN6_0),.din(w_dff_A_ph7FrcEQ1_0),.clk(gclk));
	jdff dff_A_k9shR9gN6_0(.dout(w_dff_A_PBJVTjTi4_0),.din(w_dff_A_k9shR9gN6_0),.clk(gclk));
	jdff dff_A_PBJVTjTi4_0(.dout(w_dff_A_KKnSm9h82_0),.din(w_dff_A_PBJVTjTi4_0),.clk(gclk));
	jdff dff_A_KKnSm9h82_0(.dout(w_dff_A_FtoURUJU1_0),.din(w_dff_A_KKnSm9h82_0),.clk(gclk));
	jdff dff_A_FtoURUJU1_0(.dout(w_dff_A_ZYYQSpt12_0),.din(w_dff_A_FtoURUJU1_0),.clk(gclk));
	jdff dff_A_ZYYQSpt12_0(.dout(w_dff_A_CyfyQaoC9_0),.din(w_dff_A_ZYYQSpt12_0),.clk(gclk));
	jdff dff_A_CyfyQaoC9_0(.dout(w_dff_A_N3WZ1PBY1_0),.din(w_dff_A_CyfyQaoC9_0),.clk(gclk));
	jdff dff_A_N3WZ1PBY1_0(.dout(w_dff_A_SW35YDbg5_0),.din(w_dff_A_N3WZ1PBY1_0),.clk(gclk));
	jdff dff_A_SW35YDbg5_0(.dout(w_dff_A_HI8RGUM81_0),.din(w_dff_A_SW35YDbg5_0),.clk(gclk));
	jdff dff_A_HI8RGUM81_0(.dout(w_dff_A_J9v79Wsf9_0),.din(w_dff_A_HI8RGUM81_0),.clk(gclk));
	jdff dff_A_J9v79Wsf9_0(.dout(w_dff_A_HzN4Au3a0_0),.din(w_dff_A_J9v79Wsf9_0),.clk(gclk));
	jdff dff_A_HzN4Au3a0_0(.dout(w_dff_A_lnQSdueK3_0),.din(w_dff_A_HzN4Au3a0_0),.clk(gclk));
	jdff dff_A_lnQSdueK3_0(.dout(w_dff_A_v5lUbtTR4_0),.din(w_dff_A_lnQSdueK3_0),.clk(gclk));
	jdff dff_A_v5lUbtTR4_0(.dout(w_dff_A_siiUskm97_0),.din(w_dff_A_v5lUbtTR4_0),.clk(gclk));
	jdff dff_A_siiUskm97_0(.dout(w_dff_A_ucsfF0rl3_0),.din(w_dff_A_siiUskm97_0),.clk(gclk));
	jdff dff_A_ucsfF0rl3_0(.dout(w_dff_A_vpalG9se3_0),.din(w_dff_A_ucsfF0rl3_0),.clk(gclk));
	jdff dff_A_vpalG9se3_0(.dout(w_dff_A_kjjs7I8w5_0),.din(w_dff_A_vpalG9se3_0),.clk(gclk));
	jdff dff_A_kjjs7I8w5_0(.dout(w_dff_A_B9rike742_0),.din(w_dff_A_kjjs7I8w5_0),.clk(gclk));
	jdff dff_A_B9rike742_0(.dout(G636),.din(w_dff_A_B9rike742_0),.clk(gclk));
	jdff dff_A_N46YAxsg6_2(.dout(w_dff_A_8TcrshsE6_0),.din(w_dff_A_N46YAxsg6_2),.clk(gclk));
	jdff dff_A_8TcrshsE6_0(.dout(w_dff_A_3374SqzC3_0),.din(w_dff_A_8TcrshsE6_0),.clk(gclk));
	jdff dff_A_3374SqzC3_0(.dout(w_dff_A_rfb9R1XU1_0),.din(w_dff_A_3374SqzC3_0),.clk(gclk));
	jdff dff_A_rfb9R1XU1_0(.dout(w_dff_A_25gbLvOf5_0),.din(w_dff_A_rfb9R1XU1_0),.clk(gclk));
	jdff dff_A_25gbLvOf5_0(.dout(w_dff_A_7w2yytWT2_0),.din(w_dff_A_25gbLvOf5_0),.clk(gclk));
	jdff dff_A_7w2yytWT2_0(.dout(w_dff_A_JJuSxVmI3_0),.din(w_dff_A_7w2yytWT2_0),.clk(gclk));
	jdff dff_A_JJuSxVmI3_0(.dout(w_dff_A_mMtFRIlC6_0),.din(w_dff_A_JJuSxVmI3_0),.clk(gclk));
	jdff dff_A_mMtFRIlC6_0(.dout(w_dff_A_81ut6cuy9_0),.din(w_dff_A_mMtFRIlC6_0),.clk(gclk));
	jdff dff_A_81ut6cuy9_0(.dout(w_dff_A_TcAigBwB3_0),.din(w_dff_A_81ut6cuy9_0),.clk(gclk));
	jdff dff_A_TcAigBwB3_0(.dout(w_dff_A_cxziEPDK9_0),.din(w_dff_A_TcAigBwB3_0),.clk(gclk));
	jdff dff_A_cxziEPDK9_0(.dout(w_dff_A_P3xiG4970_0),.din(w_dff_A_cxziEPDK9_0),.clk(gclk));
	jdff dff_A_P3xiG4970_0(.dout(w_dff_A_Ok59sxxA5_0),.din(w_dff_A_P3xiG4970_0),.clk(gclk));
	jdff dff_A_Ok59sxxA5_0(.dout(w_dff_A_qkfIa3ib4_0),.din(w_dff_A_Ok59sxxA5_0),.clk(gclk));
	jdff dff_A_qkfIa3ib4_0(.dout(w_dff_A_vQnTcW883_0),.din(w_dff_A_qkfIa3ib4_0),.clk(gclk));
	jdff dff_A_vQnTcW883_0(.dout(w_dff_A_GNqKwT5m5_0),.din(w_dff_A_vQnTcW883_0),.clk(gclk));
	jdff dff_A_GNqKwT5m5_0(.dout(w_dff_A_MpB9vjwZ8_0),.din(w_dff_A_GNqKwT5m5_0),.clk(gclk));
	jdff dff_A_MpB9vjwZ8_0(.dout(w_dff_A_Ib0P5ISv5_0),.din(w_dff_A_MpB9vjwZ8_0),.clk(gclk));
	jdff dff_A_Ib0P5ISv5_0(.dout(w_dff_A_J5G9ejAb0_0),.din(w_dff_A_Ib0P5ISv5_0),.clk(gclk));
	jdff dff_A_J5G9ejAb0_0(.dout(w_dff_A_VV0ccLqg3_0),.din(w_dff_A_J5G9ejAb0_0),.clk(gclk));
	jdff dff_A_VV0ccLqg3_0(.dout(w_dff_A_fhZ0wCzH2_0),.din(w_dff_A_VV0ccLqg3_0),.clk(gclk));
	jdff dff_A_fhZ0wCzH2_0(.dout(w_dff_A_rUEVe7jm1_0),.din(w_dff_A_fhZ0wCzH2_0),.clk(gclk));
	jdff dff_A_rUEVe7jm1_0(.dout(w_dff_A_n9aOoSr31_0),.din(w_dff_A_rUEVe7jm1_0),.clk(gclk));
	jdff dff_A_n9aOoSr31_0(.dout(w_dff_A_OisW3IkR8_0),.din(w_dff_A_n9aOoSr31_0),.clk(gclk));
	jdff dff_A_OisW3IkR8_0(.dout(G704),.din(w_dff_A_OisW3IkR8_0),.clk(gclk));
	jdff dff_A_2DKLk9un4_2(.dout(w_dff_A_JgRWRyUM9_0),.din(w_dff_A_2DKLk9un4_2),.clk(gclk));
	jdff dff_A_JgRWRyUM9_0(.dout(w_dff_A_sRsUIoki6_0),.din(w_dff_A_JgRWRyUM9_0),.clk(gclk));
	jdff dff_A_sRsUIoki6_0(.dout(w_dff_A_cLNbfYRR9_0),.din(w_dff_A_sRsUIoki6_0),.clk(gclk));
	jdff dff_A_cLNbfYRR9_0(.dout(w_dff_A_CzXinyke2_0),.din(w_dff_A_cLNbfYRR9_0),.clk(gclk));
	jdff dff_A_CzXinyke2_0(.dout(w_dff_A_jlDt2KvY0_0),.din(w_dff_A_CzXinyke2_0),.clk(gclk));
	jdff dff_A_jlDt2KvY0_0(.dout(w_dff_A_lHKAmdl23_0),.din(w_dff_A_jlDt2KvY0_0),.clk(gclk));
	jdff dff_A_lHKAmdl23_0(.dout(w_dff_A_meSPHwYE2_0),.din(w_dff_A_lHKAmdl23_0),.clk(gclk));
	jdff dff_A_meSPHwYE2_0(.dout(w_dff_A_5qWV42Zh4_0),.din(w_dff_A_meSPHwYE2_0),.clk(gclk));
	jdff dff_A_5qWV42Zh4_0(.dout(w_dff_A_qbs43c601_0),.din(w_dff_A_5qWV42Zh4_0),.clk(gclk));
	jdff dff_A_qbs43c601_0(.dout(w_dff_A_M8ughsjL8_0),.din(w_dff_A_qbs43c601_0),.clk(gclk));
	jdff dff_A_M8ughsjL8_0(.dout(w_dff_A_1zvoTGZW5_0),.din(w_dff_A_M8ughsjL8_0),.clk(gclk));
	jdff dff_A_1zvoTGZW5_0(.dout(w_dff_A_EEj56grY2_0),.din(w_dff_A_1zvoTGZW5_0),.clk(gclk));
	jdff dff_A_EEj56grY2_0(.dout(w_dff_A_JEWybB8X1_0),.din(w_dff_A_EEj56grY2_0),.clk(gclk));
	jdff dff_A_JEWybB8X1_0(.dout(w_dff_A_ZifTnYWB5_0),.din(w_dff_A_JEWybB8X1_0),.clk(gclk));
	jdff dff_A_ZifTnYWB5_0(.dout(w_dff_A_zYfBxUM84_0),.din(w_dff_A_ZifTnYWB5_0),.clk(gclk));
	jdff dff_A_zYfBxUM84_0(.dout(w_dff_A_LieJn0700_0),.din(w_dff_A_zYfBxUM84_0),.clk(gclk));
	jdff dff_A_LieJn0700_0(.dout(w_dff_A_gmSlfClF6_0),.din(w_dff_A_LieJn0700_0),.clk(gclk));
	jdff dff_A_gmSlfClF6_0(.dout(w_dff_A_o8esnD4y7_0),.din(w_dff_A_gmSlfClF6_0),.clk(gclk));
	jdff dff_A_o8esnD4y7_0(.dout(w_dff_A_6MMOqSuP1_0),.din(w_dff_A_o8esnD4y7_0),.clk(gclk));
	jdff dff_A_6MMOqSuP1_0(.dout(w_dff_A_IIoEG4Ic0_0),.din(w_dff_A_6MMOqSuP1_0),.clk(gclk));
	jdff dff_A_IIoEG4Ic0_0(.dout(w_dff_A_j7QSh7pg8_0),.din(w_dff_A_IIoEG4Ic0_0),.clk(gclk));
	jdff dff_A_j7QSh7pg8_0(.dout(w_dff_A_DZvvssdZ8_0),.din(w_dff_A_j7QSh7pg8_0),.clk(gclk));
	jdff dff_A_DZvvssdZ8_0(.dout(w_dff_A_605ik9r09_0),.din(w_dff_A_DZvvssdZ8_0),.clk(gclk));
	jdff dff_A_605ik9r09_0(.dout(G717),.din(w_dff_A_605ik9r09_0),.clk(gclk));
	jdff dff_A_u4ojv5bs3_2(.dout(w_dff_A_16KvtlDM5_0),.din(w_dff_A_u4ojv5bs3_2),.clk(gclk));
	jdff dff_A_16KvtlDM5_0(.dout(w_dff_A_AE1V1d4u8_0),.din(w_dff_A_16KvtlDM5_0),.clk(gclk));
	jdff dff_A_AE1V1d4u8_0(.dout(w_dff_A_5JZE5UhL5_0),.din(w_dff_A_AE1V1d4u8_0),.clk(gclk));
	jdff dff_A_5JZE5UhL5_0(.dout(w_dff_A_BFqDstg08_0),.din(w_dff_A_5JZE5UhL5_0),.clk(gclk));
	jdff dff_A_BFqDstg08_0(.dout(w_dff_A_Baqx0k3F7_0),.din(w_dff_A_BFqDstg08_0),.clk(gclk));
	jdff dff_A_Baqx0k3F7_0(.dout(w_dff_A_wvgErWK60_0),.din(w_dff_A_Baqx0k3F7_0),.clk(gclk));
	jdff dff_A_wvgErWK60_0(.dout(w_dff_A_SWFk9gmT3_0),.din(w_dff_A_wvgErWK60_0),.clk(gclk));
	jdff dff_A_SWFk9gmT3_0(.dout(w_dff_A_CQR9DwNd3_0),.din(w_dff_A_SWFk9gmT3_0),.clk(gclk));
	jdff dff_A_CQR9DwNd3_0(.dout(w_dff_A_D41rGFeQ3_0),.din(w_dff_A_CQR9DwNd3_0),.clk(gclk));
	jdff dff_A_D41rGFeQ3_0(.dout(w_dff_A_ntIYE8CX3_0),.din(w_dff_A_D41rGFeQ3_0),.clk(gclk));
	jdff dff_A_ntIYE8CX3_0(.dout(w_dff_A_HLx8Hkqy9_0),.din(w_dff_A_ntIYE8CX3_0),.clk(gclk));
	jdff dff_A_HLx8Hkqy9_0(.dout(w_dff_A_wq140oL94_0),.din(w_dff_A_HLx8Hkqy9_0),.clk(gclk));
	jdff dff_A_wq140oL94_0(.dout(w_dff_A_kBVz0q0L4_0),.din(w_dff_A_wq140oL94_0),.clk(gclk));
	jdff dff_A_kBVz0q0L4_0(.dout(w_dff_A_vPg3e92w8_0),.din(w_dff_A_kBVz0q0L4_0),.clk(gclk));
	jdff dff_A_vPg3e92w8_0(.dout(w_dff_A_2pZdvSAW8_0),.din(w_dff_A_vPg3e92w8_0),.clk(gclk));
	jdff dff_A_2pZdvSAW8_0(.dout(w_dff_A_BfJvqf762_0),.din(w_dff_A_2pZdvSAW8_0),.clk(gclk));
	jdff dff_A_BfJvqf762_0(.dout(w_dff_A_b5crP4Yu0_0),.din(w_dff_A_BfJvqf762_0),.clk(gclk));
	jdff dff_A_b5crP4Yu0_0(.dout(w_dff_A_MgVB2XwL9_0),.din(w_dff_A_b5crP4Yu0_0),.clk(gclk));
	jdff dff_A_MgVB2XwL9_0(.dout(w_dff_A_4iW5KogW8_0),.din(w_dff_A_MgVB2XwL9_0),.clk(gclk));
	jdff dff_A_4iW5KogW8_0(.dout(w_dff_A_DJNjM5wY4_0),.din(w_dff_A_4iW5KogW8_0),.clk(gclk));
	jdff dff_A_DJNjM5wY4_0(.dout(w_dff_A_r4NeWXKY5_0),.din(w_dff_A_DJNjM5wY4_0),.clk(gclk));
	jdff dff_A_r4NeWXKY5_0(.dout(w_dff_A_l70H96972_0),.din(w_dff_A_r4NeWXKY5_0),.clk(gclk));
	jdff dff_A_l70H96972_0(.dout(w_dff_A_i06YsaSI0_0),.din(w_dff_A_l70H96972_0),.clk(gclk));
	jdff dff_A_i06YsaSI0_0(.dout(w_dff_A_epPjhTZb9_0),.din(w_dff_A_i06YsaSI0_0),.clk(gclk));
	jdff dff_A_epPjhTZb9_0(.dout(G820),.din(w_dff_A_epPjhTZb9_0),.clk(gclk));
	jdff dff_A_bFJAJXPe1_2(.dout(w_dff_A_HRxkIp9o4_0),.din(w_dff_A_bFJAJXPe1_2),.clk(gclk));
	jdff dff_A_HRxkIp9o4_0(.dout(w_dff_A_brxhaajo8_0),.din(w_dff_A_HRxkIp9o4_0),.clk(gclk));
	jdff dff_A_brxhaajo8_0(.dout(w_dff_A_rqEgMzgx2_0),.din(w_dff_A_brxhaajo8_0),.clk(gclk));
	jdff dff_A_rqEgMzgx2_0(.dout(w_dff_A_xtmTGpx37_0),.din(w_dff_A_rqEgMzgx2_0),.clk(gclk));
	jdff dff_A_xtmTGpx37_0(.dout(w_dff_A_j9YDmjJY6_0),.din(w_dff_A_xtmTGpx37_0),.clk(gclk));
	jdff dff_A_j9YDmjJY6_0(.dout(w_dff_A_qFNuSUng6_0),.din(w_dff_A_j9YDmjJY6_0),.clk(gclk));
	jdff dff_A_qFNuSUng6_0(.dout(w_dff_A_jDpHhVf28_0),.din(w_dff_A_qFNuSUng6_0),.clk(gclk));
	jdff dff_A_jDpHhVf28_0(.dout(w_dff_A_SXcJ6NHi3_0),.din(w_dff_A_jDpHhVf28_0),.clk(gclk));
	jdff dff_A_SXcJ6NHi3_0(.dout(w_dff_A_iv66C4Kf9_0),.din(w_dff_A_SXcJ6NHi3_0),.clk(gclk));
	jdff dff_A_iv66C4Kf9_0(.dout(w_dff_A_mXKibCkS0_0),.din(w_dff_A_iv66C4Kf9_0),.clk(gclk));
	jdff dff_A_mXKibCkS0_0(.dout(w_dff_A_0Z5jUYvR1_0),.din(w_dff_A_mXKibCkS0_0),.clk(gclk));
	jdff dff_A_0Z5jUYvR1_0(.dout(w_dff_A_lNvV7wTx0_0),.din(w_dff_A_0Z5jUYvR1_0),.clk(gclk));
	jdff dff_A_lNvV7wTx0_0(.dout(w_dff_A_nuiuHEdQ2_0),.din(w_dff_A_lNvV7wTx0_0),.clk(gclk));
	jdff dff_A_nuiuHEdQ2_0(.dout(w_dff_A_LSOREHcD1_0),.din(w_dff_A_nuiuHEdQ2_0),.clk(gclk));
	jdff dff_A_LSOREHcD1_0(.dout(w_dff_A_0zWs6Ish4_0),.din(w_dff_A_LSOREHcD1_0),.clk(gclk));
	jdff dff_A_0zWs6Ish4_0(.dout(w_dff_A_AchSd57e2_0),.din(w_dff_A_0zWs6Ish4_0),.clk(gclk));
	jdff dff_A_AchSd57e2_0(.dout(w_dff_A_isLWvKQ74_0),.din(w_dff_A_AchSd57e2_0),.clk(gclk));
	jdff dff_A_isLWvKQ74_0(.dout(w_dff_A_2YAx5rET6_0),.din(w_dff_A_isLWvKQ74_0),.clk(gclk));
	jdff dff_A_2YAx5rET6_0(.dout(w_dff_A_XD4Wiv597_0),.din(w_dff_A_2YAx5rET6_0),.clk(gclk));
	jdff dff_A_XD4Wiv597_0(.dout(w_dff_A_93AyXj409_0),.din(w_dff_A_XD4Wiv597_0),.clk(gclk));
	jdff dff_A_93AyXj409_0(.dout(w_dff_A_Y0BA1O5Y9_0),.din(w_dff_A_93AyXj409_0),.clk(gclk));
	jdff dff_A_Y0BA1O5Y9_0(.dout(w_dff_A_BForkMmX6_0),.din(w_dff_A_Y0BA1O5Y9_0),.clk(gclk));
	jdff dff_A_BForkMmX6_0(.dout(G639),.din(w_dff_A_BForkMmX6_0),.clk(gclk));
	jdff dff_A_toTyowSq4_2(.dout(w_dff_A_huRvzYvG5_0),.din(w_dff_A_toTyowSq4_2),.clk(gclk));
	jdff dff_A_huRvzYvG5_0(.dout(w_dff_A_mrisWpg32_0),.din(w_dff_A_huRvzYvG5_0),.clk(gclk));
	jdff dff_A_mrisWpg32_0(.dout(w_dff_A_bneBZArb2_0),.din(w_dff_A_mrisWpg32_0),.clk(gclk));
	jdff dff_A_bneBZArb2_0(.dout(w_dff_A_bHtGCzG00_0),.din(w_dff_A_bneBZArb2_0),.clk(gclk));
	jdff dff_A_bHtGCzG00_0(.dout(w_dff_A_smvkZ8QC9_0),.din(w_dff_A_bHtGCzG00_0),.clk(gclk));
	jdff dff_A_smvkZ8QC9_0(.dout(w_dff_A_FIShRQMh4_0),.din(w_dff_A_smvkZ8QC9_0),.clk(gclk));
	jdff dff_A_FIShRQMh4_0(.dout(w_dff_A_ZHW6TmRm9_0),.din(w_dff_A_FIShRQMh4_0),.clk(gclk));
	jdff dff_A_ZHW6TmRm9_0(.dout(w_dff_A_Qx4k9JMK7_0),.din(w_dff_A_ZHW6TmRm9_0),.clk(gclk));
	jdff dff_A_Qx4k9JMK7_0(.dout(w_dff_A_4LjNqzSN8_0),.din(w_dff_A_Qx4k9JMK7_0),.clk(gclk));
	jdff dff_A_4LjNqzSN8_0(.dout(w_dff_A_87ywqVwj9_0),.din(w_dff_A_4LjNqzSN8_0),.clk(gclk));
	jdff dff_A_87ywqVwj9_0(.dout(w_dff_A_IgpJrgJ06_0),.din(w_dff_A_87ywqVwj9_0),.clk(gclk));
	jdff dff_A_IgpJrgJ06_0(.dout(w_dff_A_J0E4AVTD5_0),.din(w_dff_A_IgpJrgJ06_0),.clk(gclk));
	jdff dff_A_J0E4AVTD5_0(.dout(w_dff_A_5Ltba8tL6_0),.din(w_dff_A_J0E4AVTD5_0),.clk(gclk));
	jdff dff_A_5Ltba8tL6_0(.dout(w_dff_A_R86nVaq74_0),.din(w_dff_A_5Ltba8tL6_0),.clk(gclk));
	jdff dff_A_R86nVaq74_0(.dout(w_dff_A_eXhXKr1I6_0),.din(w_dff_A_R86nVaq74_0),.clk(gclk));
	jdff dff_A_eXhXKr1I6_0(.dout(w_dff_A_2t9xbKcH2_0),.din(w_dff_A_eXhXKr1I6_0),.clk(gclk));
	jdff dff_A_2t9xbKcH2_0(.dout(w_dff_A_tJcF31Fj1_0),.din(w_dff_A_2t9xbKcH2_0),.clk(gclk));
	jdff dff_A_tJcF31Fj1_0(.dout(w_dff_A_nl8SbuXr2_0),.din(w_dff_A_tJcF31Fj1_0),.clk(gclk));
	jdff dff_A_nl8SbuXr2_0(.dout(w_dff_A_waSge6q12_0),.din(w_dff_A_nl8SbuXr2_0),.clk(gclk));
	jdff dff_A_waSge6q12_0(.dout(w_dff_A_OJPwxRea2_0),.din(w_dff_A_waSge6q12_0),.clk(gclk));
	jdff dff_A_OJPwxRea2_0(.dout(w_dff_A_yxwC9F1D4_0),.din(w_dff_A_OJPwxRea2_0),.clk(gclk));
	jdff dff_A_yxwC9F1D4_0(.dout(w_dff_A_xDV7McIN4_0),.din(w_dff_A_yxwC9F1D4_0),.clk(gclk));
	jdff dff_A_xDV7McIN4_0(.dout(G673),.din(w_dff_A_xDV7McIN4_0),.clk(gclk));
	jdff dff_A_OVjaSAb91_2(.dout(w_dff_A_Y9m4OCJQ8_0),.din(w_dff_A_OVjaSAb91_2),.clk(gclk));
	jdff dff_A_Y9m4OCJQ8_0(.dout(w_dff_A_d3en3JWA3_0),.din(w_dff_A_Y9m4OCJQ8_0),.clk(gclk));
	jdff dff_A_d3en3JWA3_0(.dout(w_dff_A_8tjISI2k2_0),.din(w_dff_A_d3en3JWA3_0),.clk(gclk));
	jdff dff_A_8tjISI2k2_0(.dout(w_dff_A_Jk1Oclct9_0),.din(w_dff_A_8tjISI2k2_0),.clk(gclk));
	jdff dff_A_Jk1Oclct9_0(.dout(w_dff_A_f8fnUCoo8_0),.din(w_dff_A_Jk1Oclct9_0),.clk(gclk));
	jdff dff_A_f8fnUCoo8_0(.dout(w_dff_A_S0CLXpMb0_0),.din(w_dff_A_f8fnUCoo8_0),.clk(gclk));
	jdff dff_A_S0CLXpMb0_0(.dout(w_dff_A_IGTgyIzK7_0),.din(w_dff_A_S0CLXpMb0_0),.clk(gclk));
	jdff dff_A_IGTgyIzK7_0(.dout(w_dff_A_aicJM0Jc2_0),.din(w_dff_A_IGTgyIzK7_0),.clk(gclk));
	jdff dff_A_aicJM0Jc2_0(.dout(w_dff_A_ognLfPum9_0),.din(w_dff_A_aicJM0Jc2_0),.clk(gclk));
	jdff dff_A_ognLfPum9_0(.dout(w_dff_A_lzdKMGrs7_0),.din(w_dff_A_ognLfPum9_0),.clk(gclk));
	jdff dff_A_lzdKMGrs7_0(.dout(w_dff_A_sx8U9IIE6_0),.din(w_dff_A_lzdKMGrs7_0),.clk(gclk));
	jdff dff_A_sx8U9IIE6_0(.dout(w_dff_A_JDAyKZwk6_0),.din(w_dff_A_sx8U9IIE6_0),.clk(gclk));
	jdff dff_A_JDAyKZwk6_0(.dout(w_dff_A_kjLfUmyf6_0),.din(w_dff_A_JDAyKZwk6_0),.clk(gclk));
	jdff dff_A_kjLfUmyf6_0(.dout(w_dff_A_w7y70Prj3_0),.din(w_dff_A_kjLfUmyf6_0),.clk(gclk));
	jdff dff_A_w7y70Prj3_0(.dout(w_dff_A_Y7Tzjf2d9_0),.din(w_dff_A_w7y70Prj3_0),.clk(gclk));
	jdff dff_A_Y7Tzjf2d9_0(.dout(w_dff_A_ObMxRUlg5_0),.din(w_dff_A_Y7Tzjf2d9_0),.clk(gclk));
	jdff dff_A_ObMxRUlg5_0(.dout(w_dff_A_iaQv0iVY3_0),.din(w_dff_A_ObMxRUlg5_0),.clk(gclk));
	jdff dff_A_iaQv0iVY3_0(.dout(w_dff_A_FR42bIRy8_0),.din(w_dff_A_iaQv0iVY3_0),.clk(gclk));
	jdff dff_A_FR42bIRy8_0(.dout(w_dff_A_Z3XH0dUe1_0),.din(w_dff_A_FR42bIRy8_0),.clk(gclk));
	jdff dff_A_Z3XH0dUe1_0(.dout(w_dff_A_zjRU8IB00_0),.din(w_dff_A_Z3XH0dUe1_0),.clk(gclk));
	jdff dff_A_zjRU8IB00_0(.dout(w_dff_A_NzFuA0gO8_0),.din(w_dff_A_zjRU8IB00_0),.clk(gclk));
	jdff dff_A_NzFuA0gO8_0(.dout(w_dff_A_1wTxoZSx7_0),.din(w_dff_A_NzFuA0gO8_0),.clk(gclk));
	jdff dff_A_1wTxoZSx7_0(.dout(G707),.din(w_dff_A_1wTxoZSx7_0),.clk(gclk));
	jdff dff_A_YdWlFp8S9_2(.dout(w_dff_A_KCdz1AxZ4_0),.din(w_dff_A_YdWlFp8S9_2),.clk(gclk));
	jdff dff_A_KCdz1AxZ4_0(.dout(w_dff_A_9bUfZwSh9_0),.din(w_dff_A_KCdz1AxZ4_0),.clk(gclk));
	jdff dff_A_9bUfZwSh9_0(.dout(w_dff_A_DbnKsDVZ5_0),.din(w_dff_A_9bUfZwSh9_0),.clk(gclk));
	jdff dff_A_DbnKsDVZ5_0(.dout(w_dff_A_JLStcglA9_0),.din(w_dff_A_DbnKsDVZ5_0),.clk(gclk));
	jdff dff_A_JLStcglA9_0(.dout(w_dff_A_IHmy4y6X4_0),.din(w_dff_A_JLStcglA9_0),.clk(gclk));
	jdff dff_A_IHmy4y6X4_0(.dout(w_dff_A_z405AW0f4_0),.din(w_dff_A_IHmy4y6X4_0),.clk(gclk));
	jdff dff_A_z405AW0f4_0(.dout(w_dff_A_5D34Nn9Z9_0),.din(w_dff_A_z405AW0f4_0),.clk(gclk));
	jdff dff_A_5D34Nn9Z9_0(.dout(w_dff_A_7wpAMKDJ5_0),.din(w_dff_A_5D34Nn9Z9_0),.clk(gclk));
	jdff dff_A_7wpAMKDJ5_0(.dout(w_dff_A_7sdL923o5_0),.din(w_dff_A_7wpAMKDJ5_0),.clk(gclk));
	jdff dff_A_7sdL923o5_0(.dout(w_dff_A_hZszDikc8_0),.din(w_dff_A_7sdL923o5_0),.clk(gclk));
	jdff dff_A_hZszDikc8_0(.dout(w_dff_A_XHtnOvIV4_0),.din(w_dff_A_hZszDikc8_0),.clk(gclk));
	jdff dff_A_XHtnOvIV4_0(.dout(w_dff_A_l2TqMT775_0),.din(w_dff_A_XHtnOvIV4_0),.clk(gclk));
	jdff dff_A_l2TqMT775_0(.dout(w_dff_A_WtjTUU7V3_0),.din(w_dff_A_l2TqMT775_0),.clk(gclk));
	jdff dff_A_WtjTUU7V3_0(.dout(w_dff_A_bGyd42oc7_0),.din(w_dff_A_WtjTUU7V3_0),.clk(gclk));
	jdff dff_A_bGyd42oc7_0(.dout(w_dff_A_boebuFR06_0),.din(w_dff_A_bGyd42oc7_0),.clk(gclk));
	jdff dff_A_boebuFR06_0(.dout(w_dff_A_ilrHZdo72_0),.din(w_dff_A_boebuFR06_0),.clk(gclk));
	jdff dff_A_ilrHZdo72_0(.dout(w_dff_A_xps0psrB4_0),.din(w_dff_A_ilrHZdo72_0),.clk(gclk));
	jdff dff_A_xps0psrB4_0(.dout(w_dff_A_ADz86t9A8_0),.din(w_dff_A_xps0psrB4_0),.clk(gclk));
	jdff dff_A_ADz86t9A8_0(.dout(w_dff_A_JassX8VE4_0),.din(w_dff_A_ADz86t9A8_0),.clk(gclk));
	jdff dff_A_JassX8VE4_0(.dout(w_dff_A_clyvudyc4_0),.din(w_dff_A_JassX8VE4_0),.clk(gclk));
	jdff dff_A_clyvudyc4_0(.dout(w_dff_A_PiTLjypD1_0),.din(w_dff_A_clyvudyc4_0),.clk(gclk));
	jdff dff_A_PiTLjypD1_0(.dout(w_dff_A_PRaWv27G2_0),.din(w_dff_A_PiTLjypD1_0),.clk(gclk));
	jdff dff_A_PRaWv27G2_0(.dout(G715),.din(w_dff_A_PRaWv27G2_0),.clk(gclk));
	jdff dff_A_Cd9m9dFW8_2(.dout(w_dff_A_x1CFo4sI0_0),.din(w_dff_A_Cd9m9dFW8_2),.clk(gclk));
	jdff dff_A_x1CFo4sI0_0(.dout(w_dff_A_ZO2M8zcj7_0),.din(w_dff_A_x1CFo4sI0_0),.clk(gclk));
	jdff dff_A_ZO2M8zcj7_0(.dout(w_dff_A_TApE9Qia4_0),.din(w_dff_A_ZO2M8zcj7_0),.clk(gclk));
	jdff dff_A_TApE9Qia4_0(.dout(w_dff_A_cvEC4Gjj9_0),.din(w_dff_A_TApE9Qia4_0),.clk(gclk));
	jdff dff_A_cvEC4Gjj9_0(.dout(w_dff_A_69kCW8C87_0),.din(w_dff_A_cvEC4Gjj9_0),.clk(gclk));
	jdff dff_A_69kCW8C87_0(.dout(w_dff_A_GGNGD3Ei0_0),.din(w_dff_A_69kCW8C87_0),.clk(gclk));
	jdff dff_A_GGNGD3Ei0_0(.dout(w_dff_A_itbBHohL7_0),.din(w_dff_A_GGNGD3Ei0_0),.clk(gclk));
	jdff dff_A_itbBHohL7_0(.dout(w_dff_A_P0SKdzAc4_0),.din(w_dff_A_itbBHohL7_0),.clk(gclk));
	jdff dff_A_P0SKdzAc4_0(.dout(w_dff_A_0xQlZc8H7_0),.din(w_dff_A_P0SKdzAc4_0),.clk(gclk));
	jdff dff_A_0xQlZc8H7_0(.dout(w_dff_A_r6cAHvdX3_0),.din(w_dff_A_0xQlZc8H7_0),.clk(gclk));
	jdff dff_A_r6cAHvdX3_0(.dout(w_dff_A_W8Qf7Pa14_0),.din(w_dff_A_r6cAHvdX3_0),.clk(gclk));
	jdff dff_A_W8Qf7Pa14_0(.dout(w_dff_A_bn5LFuq27_0),.din(w_dff_A_W8Qf7Pa14_0),.clk(gclk));
	jdff dff_A_bn5LFuq27_0(.dout(w_dff_A_Ni8FRK3D5_0),.din(w_dff_A_bn5LFuq27_0),.clk(gclk));
	jdff dff_A_Ni8FRK3D5_0(.dout(w_dff_A_4GroKpjZ2_0),.din(w_dff_A_Ni8FRK3D5_0),.clk(gclk));
	jdff dff_A_4GroKpjZ2_0(.dout(w_dff_A_HZFcZRWK7_0),.din(w_dff_A_4GroKpjZ2_0),.clk(gclk));
	jdff dff_A_HZFcZRWK7_0(.dout(w_dff_A_3hiyNlRf6_0),.din(w_dff_A_HZFcZRWK7_0),.clk(gclk));
	jdff dff_A_3hiyNlRf6_0(.dout(w_dff_A_dvsqEEWl7_0),.din(w_dff_A_3hiyNlRf6_0),.clk(gclk));
	jdff dff_A_dvsqEEWl7_0(.dout(w_dff_A_jD9Sw1kX4_0),.din(w_dff_A_dvsqEEWl7_0),.clk(gclk));
	jdff dff_A_jD9Sw1kX4_0(.dout(w_dff_A_r4sKjRsk2_0),.din(w_dff_A_jD9Sw1kX4_0),.clk(gclk));
	jdff dff_A_r4sKjRsk2_0(.dout(G598),.din(w_dff_A_r4sKjRsk2_0),.clk(gclk));
	jdff dff_A_ZvM57l6Z2_2(.dout(w_dff_A_WdJboYY90_0),.din(w_dff_A_ZvM57l6Z2_2),.clk(gclk));
	jdff dff_A_WdJboYY90_0(.dout(w_dff_A_6kOSiZz19_0),.din(w_dff_A_WdJboYY90_0),.clk(gclk));
	jdff dff_A_6kOSiZz19_0(.dout(w_dff_A_RG1W8S5X7_0),.din(w_dff_A_6kOSiZz19_0),.clk(gclk));
	jdff dff_A_RG1W8S5X7_0(.dout(w_dff_A_RMyvq1En7_0),.din(w_dff_A_RG1W8S5X7_0),.clk(gclk));
	jdff dff_A_RMyvq1En7_0(.dout(w_dff_A_qCi5ix938_0),.din(w_dff_A_RMyvq1En7_0),.clk(gclk));
	jdff dff_A_qCi5ix938_0(.dout(w_dff_A_eeraTqlt9_0),.din(w_dff_A_qCi5ix938_0),.clk(gclk));
	jdff dff_A_eeraTqlt9_0(.dout(w_dff_A_IPY8snXA5_0),.din(w_dff_A_eeraTqlt9_0),.clk(gclk));
	jdff dff_A_IPY8snXA5_0(.dout(w_dff_A_NIAZ5XQd5_0),.din(w_dff_A_IPY8snXA5_0),.clk(gclk));
	jdff dff_A_NIAZ5XQd5_0(.dout(w_dff_A_QGNLrBLj6_0),.din(w_dff_A_NIAZ5XQd5_0),.clk(gclk));
	jdff dff_A_QGNLrBLj6_0(.dout(w_dff_A_2LWrXZGn6_0),.din(w_dff_A_QGNLrBLj6_0),.clk(gclk));
	jdff dff_A_2LWrXZGn6_0(.dout(w_dff_A_5tWQYmJe0_0),.din(w_dff_A_2LWrXZGn6_0),.clk(gclk));
	jdff dff_A_5tWQYmJe0_0(.dout(w_dff_A_utghDYRT6_0),.din(w_dff_A_5tWQYmJe0_0),.clk(gclk));
	jdff dff_A_utghDYRT6_0(.dout(w_dff_A_2p0QNLZG3_0),.din(w_dff_A_utghDYRT6_0),.clk(gclk));
	jdff dff_A_2p0QNLZG3_0(.dout(w_dff_A_EDWWRofg9_0),.din(w_dff_A_2p0QNLZG3_0),.clk(gclk));
	jdff dff_A_EDWWRofg9_0(.dout(w_dff_A_n3ScF3jt9_0),.din(w_dff_A_EDWWRofg9_0),.clk(gclk));
	jdff dff_A_n3ScF3jt9_0(.dout(w_dff_A_PiVqCAeu7_0),.din(w_dff_A_n3ScF3jt9_0),.clk(gclk));
	jdff dff_A_PiVqCAeu7_0(.dout(w_dff_A_oKIJQUEf6_0),.din(w_dff_A_PiVqCAeu7_0),.clk(gclk));
	jdff dff_A_oKIJQUEf6_0(.dout(w_dff_A_S5A92AwA3_0),.din(w_dff_A_oKIJQUEf6_0),.clk(gclk));
	jdff dff_A_S5A92AwA3_0(.dout(G610),.din(w_dff_A_S5A92AwA3_0),.clk(gclk));
	jdff dff_A_NVY0g9Mn7_2(.dout(w_dff_A_te31V8tb8_0),.din(w_dff_A_NVY0g9Mn7_2),.clk(gclk));
	jdff dff_A_te31V8tb8_0(.dout(w_dff_A_7PSFedEB8_0),.din(w_dff_A_te31V8tb8_0),.clk(gclk));
	jdff dff_A_7PSFedEB8_0(.dout(w_dff_A_cSiEQ6Tz3_0),.din(w_dff_A_7PSFedEB8_0),.clk(gclk));
	jdff dff_A_cSiEQ6Tz3_0(.dout(w_dff_A_9wrg9FnJ0_0),.din(w_dff_A_cSiEQ6Tz3_0),.clk(gclk));
	jdff dff_A_9wrg9FnJ0_0(.dout(w_dff_A_MtM22qNV1_0),.din(w_dff_A_9wrg9FnJ0_0),.clk(gclk));
	jdff dff_A_MtM22qNV1_0(.dout(w_dff_A_xyOHZi835_0),.din(w_dff_A_MtM22qNV1_0),.clk(gclk));
	jdff dff_A_xyOHZi835_0(.dout(w_dff_A_gynlntUb3_0),.din(w_dff_A_xyOHZi835_0),.clk(gclk));
	jdff dff_A_gynlntUb3_0(.dout(w_dff_A_xFQm1ZIx9_0),.din(w_dff_A_gynlntUb3_0),.clk(gclk));
	jdff dff_A_xFQm1ZIx9_0(.dout(w_dff_A_acEaxo339_0),.din(w_dff_A_xFQm1ZIx9_0),.clk(gclk));
	jdff dff_A_acEaxo339_0(.dout(w_dff_A_phwkpT6u2_0),.din(w_dff_A_acEaxo339_0),.clk(gclk));
	jdff dff_A_phwkpT6u2_0(.dout(w_dff_A_3kII0ws02_0),.din(w_dff_A_phwkpT6u2_0),.clk(gclk));
	jdff dff_A_3kII0ws02_0(.dout(w_dff_A_MNbb10fD7_0),.din(w_dff_A_3kII0ws02_0),.clk(gclk));
	jdff dff_A_MNbb10fD7_0(.dout(w_dff_A_9iz9nXQX7_0),.din(w_dff_A_MNbb10fD7_0),.clk(gclk));
	jdff dff_A_9iz9nXQX7_0(.dout(w_dff_A_ILKO7dgF6_0),.din(w_dff_A_9iz9nXQX7_0),.clk(gclk));
	jdff dff_A_ILKO7dgF6_0(.dout(w_dff_A_atIJreu34_0),.din(w_dff_A_ILKO7dgF6_0),.clk(gclk));
	jdff dff_A_atIJreu34_0(.dout(w_dff_A_3WiXZ4bC9_0),.din(w_dff_A_atIJreu34_0),.clk(gclk));
	jdff dff_A_3WiXZ4bC9_0(.dout(G588),.din(w_dff_A_3WiXZ4bC9_0),.clk(gclk));
	jdff dff_A_mk7Y1tBd1_2(.dout(w_dff_A_XWkYgDBl3_0),.din(w_dff_A_mk7Y1tBd1_2),.clk(gclk));
	jdff dff_A_XWkYgDBl3_0(.dout(w_dff_A_MYYB1R0X3_0),.din(w_dff_A_XWkYgDBl3_0),.clk(gclk));
	jdff dff_A_MYYB1R0X3_0(.dout(w_dff_A_EEHsWfuj6_0),.din(w_dff_A_MYYB1R0X3_0),.clk(gclk));
	jdff dff_A_EEHsWfuj6_0(.dout(w_dff_A_VrCn3CYH3_0),.din(w_dff_A_EEHsWfuj6_0),.clk(gclk));
	jdff dff_A_VrCn3CYH3_0(.dout(w_dff_A_4WCah3Wi3_0),.din(w_dff_A_VrCn3CYH3_0),.clk(gclk));
	jdff dff_A_4WCah3Wi3_0(.dout(w_dff_A_6bc9hTeH8_0),.din(w_dff_A_4WCah3Wi3_0),.clk(gclk));
	jdff dff_A_6bc9hTeH8_0(.dout(w_dff_A_AUrJXpFU8_0),.din(w_dff_A_6bc9hTeH8_0),.clk(gclk));
	jdff dff_A_AUrJXpFU8_0(.dout(w_dff_A_1Nuf7zd55_0),.din(w_dff_A_AUrJXpFU8_0),.clk(gclk));
	jdff dff_A_1Nuf7zd55_0(.dout(w_dff_A_RRrW0xeS8_0),.din(w_dff_A_1Nuf7zd55_0),.clk(gclk));
	jdff dff_A_RRrW0xeS8_0(.dout(w_dff_A_4t3pMGx94_0),.din(w_dff_A_RRrW0xeS8_0),.clk(gclk));
	jdff dff_A_4t3pMGx94_0(.dout(w_dff_A_A1kuQrvv4_0),.din(w_dff_A_4t3pMGx94_0),.clk(gclk));
	jdff dff_A_A1kuQrvv4_0(.dout(w_dff_A_Sg7zNRAK4_0),.din(w_dff_A_A1kuQrvv4_0),.clk(gclk));
	jdff dff_A_Sg7zNRAK4_0(.dout(w_dff_A_nyCrfboS4_0),.din(w_dff_A_Sg7zNRAK4_0),.clk(gclk));
	jdff dff_A_nyCrfboS4_0(.dout(w_dff_A_GrVukXrF5_0),.din(w_dff_A_nyCrfboS4_0),.clk(gclk));
	jdff dff_A_GrVukXrF5_0(.dout(w_dff_A_m6xzbOsq9_0),.din(w_dff_A_GrVukXrF5_0),.clk(gclk));
	jdff dff_A_m6xzbOsq9_0(.dout(w_dff_A_ZUlGVPQ64_0),.din(w_dff_A_m6xzbOsq9_0),.clk(gclk));
	jdff dff_A_ZUlGVPQ64_0(.dout(w_dff_A_Csz3Tef33_0),.din(w_dff_A_ZUlGVPQ64_0),.clk(gclk));
	jdff dff_A_Csz3Tef33_0(.dout(G615),.din(w_dff_A_Csz3Tef33_0),.clk(gclk));
	jdff dff_A_Bq7pFif89_2(.dout(w_dff_A_NyBMqd4Z6_0),.din(w_dff_A_Bq7pFif89_2),.clk(gclk));
	jdff dff_A_NyBMqd4Z6_0(.dout(w_dff_A_qcNk22lr4_0),.din(w_dff_A_NyBMqd4Z6_0),.clk(gclk));
	jdff dff_A_qcNk22lr4_0(.dout(w_dff_A_I8yrylqY5_0),.din(w_dff_A_qcNk22lr4_0),.clk(gclk));
	jdff dff_A_I8yrylqY5_0(.dout(w_dff_A_WeN5lfva2_0),.din(w_dff_A_I8yrylqY5_0),.clk(gclk));
	jdff dff_A_WeN5lfva2_0(.dout(w_dff_A_eeV7OZKH9_0),.din(w_dff_A_WeN5lfva2_0),.clk(gclk));
	jdff dff_A_eeV7OZKH9_0(.dout(w_dff_A_Q1SYxoPh1_0),.din(w_dff_A_eeV7OZKH9_0),.clk(gclk));
	jdff dff_A_Q1SYxoPh1_0(.dout(w_dff_A_1MwazopU0_0),.din(w_dff_A_Q1SYxoPh1_0),.clk(gclk));
	jdff dff_A_1MwazopU0_0(.dout(w_dff_A_gcK41StV0_0),.din(w_dff_A_1MwazopU0_0),.clk(gclk));
	jdff dff_A_gcK41StV0_0(.dout(w_dff_A_ohIOO6na6_0),.din(w_dff_A_gcK41StV0_0),.clk(gclk));
	jdff dff_A_ohIOO6na6_0(.dout(w_dff_A_9E7vaMOn9_0),.din(w_dff_A_ohIOO6na6_0),.clk(gclk));
	jdff dff_A_9E7vaMOn9_0(.dout(w_dff_A_gO7jvR3r9_0),.din(w_dff_A_9E7vaMOn9_0),.clk(gclk));
	jdff dff_A_gO7jvR3r9_0(.dout(w_dff_A_3rtWMCxk3_0),.din(w_dff_A_gO7jvR3r9_0),.clk(gclk));
	jdff dff_A_3rtWMCxk3_0(.dout(w_dff_A_iOEkgF5u4_0),.din(w_dff_A_3rtWMCxk3_0),.clk(gclk));
	jdff dff_A_iOEkgF5u4_0(.dout(w_dff_A_8k6WEvqe0_0),.din(w_dff_A_iOEkgF5u4_0),.clk(gclk));
	jdff dff_A_8k6WEvqe0_0(.dout(w_dff_A_0dsAzb7T7_0),.din(w_dff_A_8k6WEvqe0_0),.clk(gclk));
	jdff dff_A_0dsAzb7T7_0(.dout(w_dff_A_fxjTDloC7_0),.din(w_dff_A_0dsAzb7T7_0),.clk(gclk));
	jdff dff_A_fxjTDloC7_0(.dout(w_dff_A_NoDo0o8j6_0),.din(w_dff_A_fxjTDloC7_0),.clk(gclk));
	jdff dff_A_NoDo0o8j6_0(.dout(G626),.din(w_dff_A_NoDo0o8j6_0),.clk(gclk));
	jdff dff_A_evdjIyls0_2(.dout(w_dff_A_jzBkylD54_0),.din(w_dff_A_evdjIyls0_2),.clk(gclk));
	jdff dff_A_jzBkylD54_0(.dout(w_dff_A_dOvZoZQW8_0),.din(w_dff_A_jzBkylD54_0),.clk(gclk));
	jdff dff_A_dOvZoZQW8_0(.dout(w_dff_A_flU1OcbQ4_0),.din(w_dff_A_dOvZoZQW8_0),.clk(gclk));
	jdff dff_A_flU1OcbQ4_0(.dout(w_dff_A_IaCaBPG70_0),.din(w_dff_A_flU1OcbQ4_0),.clk(gclk));
	jdff dff_A_IaCaBPG70_0(.dout(w_dff_A_MNscD1Yw7_0),.din(w_dff_A_IaCaBPG70_0),.clk(gclk));
	jdff dff_A_MNscD1Yw7_0(.dout(w_dff_A_qCZCqPYK8_0),.din(w_dff_A_MNscD1Yw7_0),.clk(gclk));
	jdff dff_A_qCZCqPYK8_0(.dout(w_dff_A_RutWYGiw4_0),.din(w_dff_A_qCZCqPYK8_0),.clk(gclk));
	jdff dff_A_RutWYGiw4_0(.dout(w_dff_A_LINAJobM1_0),.din(w_dff_A_RutWYGiw4_0),.clk(gclk));
	jdff dff_A_LINAJobM1_0(.dout(w_dff_A_Enp72iWw3_0),.din(w_dff_A_LINAJobM1_0),.clk(gclk));
	jdff dff_A_Enp72iWw3_0(.dout(w_dff_A_7Xzq3iC61_0),.din(w_dff_A_Enp72iWw3_0),.clk(gclk));
	jdff dff_A_7Xzq3iC61_0(.dout(w_dff_A_t84mrXfC6_0),.din(w_dff_A_7Xzq3iC61_0),.clk(gclk));
	jdff dff_A_t84mrXfC6_0(.dout(w_dff_A_WQLg3pm16_0),.din(w_dff_A_t84mrXfC6_0),.clk(gclk));
	jdff dff_A_WQLg3pm16_0(.dout(w_dff_A_llFN5Ogb6_0),.din(w_dff_A_WQLg3pm16_0),.clk(gclk));
	jdff dff_A_llFN5Ogb6_0(.dout(w_dff_A_IFpwLAmU4_0),.din(w_dff_A_llFN5Ogb6_0),.clk(gclk));
	jdff dff_A_IFpwLAmU4_0(.dout(w_dff_A_xc9BbSpL5_0),.din(w_dff_A_IFpwLAmU4_0),.clk(gclk));
	jdff dff_A_xc9BbSpL5_0(.dout(w_dff_A_TOOwjg3q4_0),.din(w_dff_A_xc9BbSpL5_0),.clk(gclk));
	jdff dff_A_TOOwjg3q4_0(.dout(G632),.din(w_dff_A_TOOwjg3q4_0),.clk(gclk));
	jdff dff_A_jptqbv0j0_1(.dout(w_dff_A_FtqcvtRC6_0),.din(w_dff_A_jptqbv0j0_1),.clk(gclk));
	jdff dff_A_FtqcvtRC6_0(.dout(w_dff_A_3LSHXnf81_0),.din(w_dff_A_FtqcvtRC6_0),.clk(gclk));
	jdff dff_A_3LSHXnf81_0(.dout(w_dff_A_gp9y5sWh5_0),.din(w_dff_A_3LSHXnf81_0),.clk(gclk));
	jdff dff_A_gp9y5sWh5_0(.dout(w_dff_A_pYAb7dtf3_0),.din(w_dff_A_gp9y5sWh5_0),.clk(gclk));
	jdff dff_A_pYAb7dtf3_0(.dout(w_dff_A_VCTACPVm4_0),.din(w_dff_A_pYAb7dtf3_0),.clk(gclk));
	jdff dff_A_VCTACPVm4_0(.dout(w_dff_A_DqzWFCu97_0),.din(w_dff_A_VCTACPVm4_0),.clk(gclk));
	jdff dff_A_DqzWFCu97_0(.dout(w_dff_A_mbaUhdEn2_0),.din(w_dff_A_DqzWFCu97_0),.clk(gclk));
	jdff dff_A_mbaUhdEn2_0(.dout(w_dff_A_8PlfjvkJ0_0),.din(w_dff_A_mbaUhdEn2_0),.clk(gclk));
	jdff dff_A_8PlfjvkJ0_0(.dout(w_dff_A_AmAi9hWm9_0),.din(w_dff_A_8PlfjvkJ0_0),.clk(gclk));
	jdff dff_A_AmAi9hWm9_0(.dout(w_dff_A_Dfn5Cc469_0),.din(w_dff_A_AmAi9hWm9_0),.clk(gclk));
	jdff dff_A_Dfn5Cc469_0(.dout(w_dff_A_7Wt5ohOY3_0),.din(w_dff_A_Dfn5Cc469_0),.clk(gclk));
	jdff dff_A_7Wt5ohOY3_0(.dout(w_dff_A_gE6SrsAq3_0),.din(w_dff_A_7Wt5ohOY3_0),.clk(gclk));
	jdff dff_A_gE6SrsAq3_0(.dout(w_dff_A_HAroxZOP3_0),.din(w_dff_A_gE6SrsAq3_0),.clk(gclk));
	jdff dff_A_HAroxZOP3_0(.dout(w_dff_A_tZoFuRcZ1_0),.din(w_dff_A_HAroxZOP3_0),.clk(gclk));
	jdff dff_A_tZoFuRcZ1_0(.dout(w_dff_A_GEJ6F2ho5_0),.din(w_dff_A_tZoFuRcZ1_0),.clk(gclk));
	jdff dff_A_GEJ6F2ho5_0(.dout(w_dff_A_i5tlMJ861_0),.din(w_dff_A_GEJ6F2ho5_0),.clk(gclk));
	jdff dff_A_i5tlMJ861_0(.dout(w_dff_A_p4bE12gd5_0),.din(w_dff_A_i5tlMJ861_0),.clk(gclk));
	jdff dff_A_p4bE12gd5_0(.dout(w_dff_A_4uzXs4RZ7_0),.din(w_dff_A_p4bE12gd5_0),.clk(gclk));
	jdff dff_A_4uzXs4RZ7_0(.dout(w_dff_A_7mdSQPoi2_0),.din(w_dff_A_4uzXs4RZ7_0),.clk(gclk));
	jdff dff_A_7mdSQPoi2_0(.dout(w_dff_A_51ifvy761_0),.din(w_dff_A_7mdSQPoi2_0),.clk(gclk));
	jdff dff_A_51ifvy761_0(.dout(w_dff_A_c0AQma3q7_0),.din(w_dff_A_51ifvy761_0),.clk(gclk));
	jdff dff_A_c0AQma3q7_0(.dout(w_dff_A_Ict1Uw3T0_0),.din(w_dff_A_c0AQma3q7_0),.clk(gclk));
	jdff dff_A_Ict1Uw3T0_0(.dout(G1002),.din(w_dff_A_Ict1Uw3T0_0),.clk(gclk));
	jdff dff_A_Pd8CgEzt0_1(.dout(w_dff_A_v7Pd294j0_0),.din(w_dff_A_Pd8CgEzt0_1),.clk(gclk));
	jdff dff_A_v7Pd294j0_0(.dout(w_dff_A_2S2kANZ27_0),.din(w_dff_A_v7Pd294j0_0),.clk(gclk));
	jdff dff_A_2S2kANZ27_0(.dout(w_dff_A_hC0YtMyi8_0),.din(w_dff_A_2S2kANZ27_0),.clk(gclk));
	jdff dff_A_hC0YtMyi8_0(.dout(w_dff_A_YYD5lvIl2_0),.din(w_dff_A_hC0YtMyi8_0),.clk(gclk));
	jdff dff_A_YYD5lvIl2_0(.dout(w_dff_A_XLHXkMNy9_0),.din(w_dff_A_YYD5lvIl2_0),.clk(gclk));
	jdff dff_A_XLHXkMNy9_0(.dout(w_dff_A_wC4oP5EB6_0),.din(w_dff_A_XLHXkMNy9_0),.clk(gclk));
	jdff dff_A_wC4oP5EB6_0(.dout(w_dff_A_cHdSX8lB0_0),.din(w_dff_A_wC4oP5EB6_0),.clk(gclk));
	jdff dff_A_cHdSX8lB0_0(.dout(w_dff_A_OPyH4G9c4_0),.din(w_dff_A_cHdSX8lB0_0),.clk(gclk));
	jdff dff_A_OPyH4G9c4_0(.dout(w_dff_A_Nnbs9u3D5_0),.din(w_dff_A_OPyH4G9c4_0),.clk(gclk));
	jdff dff_A_Nnbs9u3D5_0(.dout(w_dff_A_UHG6XuRY9_0),.din(w_dff_A_Nnbs9u3D5_0),.clk(gclk));
	jdff dff_A_UHG6XuRY9_0(.dout(w_dff_A_YlzH4YUg0_0),.din(w_dff_A_UHG6XuRY9_0),.clk(gclk));
	jdff dff_A_YlzH4YUg0_0(.dout(w_dff_A_Cd08q5VN0_0),.din(w_dff_A_YlzH4YUg0_0),.clk(gclk));
	jdff dff_A_Cd08q5VN0_0(.dout(w_dff_A_PUGdYKYd2_0),.din(w_dff_A_Cd08q5VN0_0),.clk(gclk));
	jdff dff_A_PUGdYKYd2_0(.dout(w_dff_A_C5C7xX8N9_0),.din(w_dff_A_PUGdYKYd2_0),.clk(gclk));
	jdff dff_A_C5C7xX8N9_0(.dout(w_dff_A_OJ08mxmH9_0),.din(w_dff_A_C5C7xX8N9_0),.clk(gclk));
	jdff dff_A_OJ08mxmH9_0(.dout(w_dff_A_U0S7q3rb6_0),.din(w_dff_A_OJ08mxmH9_0),.clk(gclk));
	jdff dff_A_U0S7q3rb6_0(.dout(w_dff_A_4EP3LCcU4_0),.din(w_dff_A_U0S7q3rb6_0),.clk(gclk));
	jdff dff_A_4EP3LCcU4_0(.dout(w_dff_A_nqM6Xfxs1_0),.din(w_dff_A_4EP3LCcU4_0),.clk(gclk));
	jdff dff_A_nqM6Xfxs1_0(.dout(w_dff_A_y6gvat6o4_0),.din(w_dff_A_nqM6Xfxs1_0),.clk(gclk));
	jdff dff_A_y6gvat6o4_0(.dout(w_dff_A_rIVKxv6q7_0),.din(w_dff_A_y6gvat6o4_0),.clk(gclk));
	jdff dff_A_rIVKxv6q7_0(.dout(w_dff_A_2VdlY8Fw0_0),.din(w_dff_A_rIVKxv6q7_0),.clk(gclk));
	jdff dff_A_2VdlY8Fw0_0(.dout(w_dff_A_RldWZnr82_0),.din(w_dff_A_2VdlY8Fw0_0),.clk(gclk));
	jdff dff_A_RldWZnr82_0(.dout(G1004),.din(w_dff_A_RldWZnr82_0),.clk(gclk));
	jdff dff_A_q1kryMCV0_2(.dout(w_dff_A_aRU6WpdG5_0),.din(w_dff_A_q1kryMCV0_2),.clk(gclk));
	jdff dff_A_aRU6WpdG5_0(.dout(w_dff_A_neWwQV9V9_0),.din(w_dff_A_aRU6WpdG5_0),.clk(gclk));
	jdff dff_A_neWwQV9V9_0(.dout(w_dff_A_ZCBEazSx6_0),.din(w_dff_A_neWwQV9V9_0),.clk(gclk));
	jdff dff_A_ZCBEazSx6_0(.dout(w_dff_A_gZXIM8G05_0),.din(w_dff_A_ZCBEazSx6_0),.clk(gclk));
	jdff dff_A_gZXIM8G05_0(.dout(w_dff_A_LT7T9m3H3_0),.din(w_dff_A_gZXIM8G05_0),.clk(gclk));
	jdff dff_A_LT7T9m3H3_0(.dout(w_dff_A_3nXPjOxT4_0),.din(w_dff_A_LT7T9m3H3_0),.clk(gclk));
	jdff dff_A_3nXPjOxT4_0(.dout(w_dff_A_TVwHny2S3_0),.din(w_dff_A_3nXPjOxT4_0),.clk(gclk));
	jdff dff_A_TVwHny2S3_0(.dout(w_dff_A_8aftCEWg1_0),.din(w_dff_A_TVwHny2S3_0),.clk(gclk));
	jdff dff_A_8aftCEWg1_0(.dout(w_dff_A_JKR21ULp9_0),.din(w_dff_A_8aftCEWg1_0),.clk(gclk));
	jdff dff_A_JKR21ULp9_0(.dout(w_dff_A_qH4se6w52_0),.din(w_dff_A_JKR21ULp9_0),.clk(gclk));
	jdff dff_A_qH4se6w52_0(.dout(w_dff_A_wEQxfWDP6_0),.din(w_dff_A_qH4se6w52_0),.clk(gclk));
	jdff dff_A_wEQxfWDP6_0(.dout(w_dff_A_mlub69cP0_0),.din(w_dff_A_wEQxfWDP6_0),.clk(gclk));
	jdff dff_A_mlub69cP0_0(.dout(w_dff_A_APahAb4G9_0),.din(w_dff_A_mlub69cP0_0),.clk(gclk));
	jdff dff_A_APahAb4G9_0(.dout(G591),.din(w_dff_A_APahAb4G9_0),.clk(gclk));
	jdff dff_A_LaQp9IAo6_2(.dout(w_dff_A_PgdewXPo4_0),.din(w_dff_A_LaQp9IAo6_2),.clk(gclk));
	jdff dff_A_PgdewXPo4_0(.dout(w_dff_A_0JXjAOFx6_0),.din(w_dff_A_PgdewXPo4_0),.clk(gclk));
	jdff dff_A_0JXjAOFx6_0(.dout(w_dff_A_z9jSVDB27_0),.din(w_dff_A_0JXjAOFx6_0),.clk(gclk));
	jdff dff_A_z9jSVDB27_0(.dout(w_dff_A_66Et3iiE7_0),.din(w_dff_A_z9jSVDB27_0),.clk(gclk));
	jdff dff_A_66Et3iiE7_0(.dout(w_dff_A_CjumOJ5r8_0),.din(w_dff_A_66Et3iiE7_0),.clk(gclk));
	jdff dff_A_CjumOJ5r8_0(.dout(w_dff_A_Si0UQOSo6_0),.din(w_dff_A_CjumOJ5r8_0),.clk(gclk));
	jdff dff_A_Si0UQOSo6_0(.dout(w_dff_A_oYrTmP3u3_0),.din(w_dff_A_Si0UQOSo6_0),.clk(gclk));
	jdff dff_A_oYrTmP3u3_0(.dout(w_dff_A_8QS1SAlJ2_0),.din(w_dff_A_oYrTmP3u3_0),.clk(gclk));
	jdff dff_A_8QS1SAlJ2_0(.dout(w_dff_A_65bIpZYP5_0),.din(w_dff_A_8QS1SAlJ2_0),.clk(gclk));
	jdff dff_A_65bIpZYP5_0(.dout(w_dff_A_ZhJTY5Jk0_0),.din(w_dff_A_65bIpZYP5_0),.clk(gclk));
	jdff dff_A_ZhJTY5Jk0_0(.dout(w_dff_A_N8mTUgdb1_0),.din(w_dff_A_ZhJTY5Jk0_0),.clk(gclk));
	jdff dff_A_N8mTUgdb1_0(.dout(w_dff_A_Zrs1DhXz5_0),.din(w_dff_A_N8mTUgdb1_0),.clk(gclk));
	jdff dff_A_Zrs1DhXz5_0(.dout(w_dff_A_dQPZa2Kn0_0),.din(w_dff_A_Zrs1DhXz5_0),.clk(gclk));
	jdff dff_A_dQPZa2Kn0_0(.dout(w_dff_A_Z1WTcebV0_0),.din(w_dff_A_dQPZa2Kn0_0),.clk(gclk));
	jdff dff_A_Z1WTcebV0_0(.dout(G618),.din(w_dff_A_Z1WTcebV0_0),.clk(gclk));
	jdff dff_A_QcszTcHB2_2(.dout(w_dff_A_pIDMkYQ89_0),.din(w_dff_A_QcszTcHB2_2),.clk(gclk));
	jdff dff_A_pIDMkYQ89_0(.dout(w_dff_A_cOkzL3up4_0),.din(w_dff_A_pIDMkYQ89_0),.clk(gclk));
	jdff dff_A_cOkzL3up4_0(.dout(w_dff_A_u9CK4Sxx0_0),.din(w_dff_A_cOkzL3up4_0),.clk(gclk));
	jdff dff_A_u9CK4Sxx0_0(.dout(w_dff_A_PsOa3JsT8_0),.din(w_dff_A_u9CK4Sxx0_0),.clk(gclk));
	jdff dff_A_PsOa3JsT8_0(.dout(w_dff_A_TsbGEXhh5_0),.din(w_dff_A_PsOa3JsT8_0),.clk(gclk));
	jdff dff_A_TsbGEXhh5_0(.dout(w_dff_A_3dlKoi9A8_0),.din(w_dff_A_TsbGEXhh5_0),.clk(gclk));
	jdff dff_A_3dlKoi9A8_0(.dout(w_dff_A_MSz5598y0_0),.din(w_dff_A_3dlKoi9A8_0),.clk(gclk));
	jdff dff_A_MSz5598y0_0(.dout(w_dff_A_18B72YHQ9_0),.din(w_dff_A_MSz5598y0_0),.clk(gclk));
	jdff dff_A_18B72YHQ9_0(.dout(w_dff_A_r3B5LYTP4_0),.din(w_dff_A_18B72YHQ9_0),.clk(gclk));
	jdff dff_A_r3B5LYTP4_0(.dout(w_dff_A_mvRDQt976_0),.din(w_dff_A_r3B5LYTP4_0),.clk(gclk));
	jdff dff_A_mvRDQt976_0(.dout(w_dff_A_nFHU9ngs0_0),.din(w_dff_A_mvRDQt976_0),.clk(gclk));
	jdff dff_A_nFHU9ngs0_0(.dout(w_dff_A_Y8YY6d2j0_0),.din(w_dff_A_nFHU9ngs0_0),.clk(gclk));
	jdff dff_A_Y8YY6d2j0_0(.dout(w_dff_A_eHysdSF98_0),.din(w_dff_A_Y8YY6d2j0_0),.clk(gclk));
	jdff dff_A_eHysdSF98_0(.dout(G621),.din(w_dff_A_eHysdSF98_0),.clk(gclk));
	jdff dff_A_wQ8OfEWM6_2(.dout(w_dff_A_aELJTW9w2_0),.din(w_dff_A_wQ8OfEWM6_2),.clk(gclk));
	jdff dff_A_aELJTW9w2_0(.dout(w_dff_A_pE0RVzCB1_0),.din(w_dff_A_aELJTW9w2_0),.clk(gclk));
	jdff dff_A_pE0RVzCB1_0(.dout(w_dff_A_biQdVpgB5_0),.din(w_dff_A_pE0RVzCB1_0),.clk(gclk));
	jdff dff_A_biQdVpgB5_0(.dout(w_dff_A_ZkOG7nRf2_0),.din(w_dff_A_biQdVpgB5_0),.clk(gclk));
	jdff dff_A_ZkOG7nRf2_0(.dout(w_dff_A_FAMRmQsz3_0),.din(w_dff_A_ZkOG7nRf2_0),.clk(gclk));
	jdff dff_A_FAMRmQsz3_0(.dout(w_dff_A_w7XM9guO7_0),.din(w_dff_A_FAMRmQsz3_0),.clk(gclk));
	jdff dff_A_w7XM9guO7_0(.dout(w_dff_A_pHhItWgi0_0),.din(w_dff_A_w7XM9guO7_0),.clk(gclk));
	jdff dff_A_pHhItWgi0_0(.dout(w_dff_A_AU7jaCK34_0),.din(w_dff_A_pHhItWgi0_0),.clk(gclk));
	jdff dff_A_AU7jaCK34_0(.dout(w_dff_A_0WpNeB0Z9_0),.din(w_dff_A_AU7jaCK34_0),.clk(gclk));
	jdff dff_A_0WpNeB0Z9_0(.dout(w_dff_A_PC8ItbCz1_0),.din(w_dff_A_0WpNeB0Z9_0),.clk(gclk));
	jdff dff_A_PC8ItbCz1_0(.dout(w_dff_A_btSCVhcQ1_0),.din(w_dff_A_PC8ItbCz1_0),.clk(gclk));
	jdff dff_A_btSCVhcQ1_0(.dout(w_dff_A_6S4bjSJH8_0),.din(w_dff_A_btSCVhcQ1_0),.clk(gclk));
	jdff dff_A_6S4bjSJH8_0(.dout(w_dff_A_v3qbmY2d3_0),.din(w_dff_A_6S4bjSJH8_0),.clk(gclk));
	jdff dff_A_v3qbmY2d3_0(.dout(w_dff_A_Z2ObU6dd2_0),.din(w_dff_A_v3qbmY2d3_0),.clk(gclk));
	jdff dff_A_Z2ObU6dd2_0(.dout(G629),.din(w_dff_A_Z2ObU6dd2_0),.clk(gclk));
	jdff dff_A_JwnIrGQk0_1(.dout(w_dff_A_C4xH7tVi7_0),.din(w_dff_A_JwnIrGQk0_1),.clk(gclk));
	jdff dff_A_C4xH7tVi7_0(.dout(w_dff_A_OcGXpt8Z9_0),.din(w_dff_A_C4xH7tVi7_0),.clk(gclk));
	jdff dff_A_OcGXpt8Z9_0(.dout(w_dff_A_n91V6SEJ8_0),.din(w_dff_A_OcGXpt8Z9_0),.clk(gclk));
	jdff dff_A_n91V6SEJ8_0(.dout(w_dff_A_tynL68rk3_0),.din(w_dff_A_n91V6SEJ8_0),.clk(gclk));
	jdff dff_A_tynL68rk3_0(.dout(w_dff_A_hGwbCVo08_0),.din(w_dff_A_tynL68rk3_0),.clk(gclk));
	jdff dff_A_hGwbCVo08_0(.dout(w_dff_A_8nc4jCvo7_0),.din(w_dff_A_hGwbCVo08_0),.clk(gclk));
	jdff dff_A_8nc4jCvo7_0(.dout(w_dff_A_IKyIqu9h2_0),.din(w_dff_A_8nc4jCvo7_0),.clk(gclk));
	jdff dff_A_IKyIqu9h2_0(.dout(w_dff_A_3Ky37lAy2_0),.din(w_dff_A_IKyIqu9h2_0),.clk(gclk));
	jdff dff_A_3Ky37lAy2_0(.dout(w_dff_A_vvi2pJoo8_0),.din(w_dff_A_3Ky37lAy2_0),.clk(gclk));
	jdff dff_A_vvi2pJoo8_0(.dout(w_dff_A_2zdUVoqD6_0),.din(w_dff_A_vvi2pJoo8_0),.clk(gclk));
	jdff dff_A_2zdUVoqD6_0(.dout(w_dff_A_1CsSKF3k1_0),.din(w_dff_A_2zdUVoqD6_0),.clk(gclk));
	jdff dff_A_1CsSKF3k1_0(.dout(w_dff_A_KmtHVL3c2_0),.din(w_dff_A_1CsSKF3k1_0),.clk(gclk));
	jdff dff_A_KmtHVL3c2_0(.dout(w_dff_A_GjFEdSDm0_0),.din(w_dff_A_KmtHVL3c2_0),.clk(gclk));
	jdff dff_A_GjFEdSDm0_0(.dout(w_dff_A_QAetyHhr6_0),.din(w_dff_A_GjFEdSDm0_0),.clk(gclk));
	jdff dff_A_QAetyHhr6_0(.dout(w_dff_A_VwPCmeLr2_0),.din(w_dff_A_QAetyHhr6_0),.clk(gclk));
	jdff dff_A_VwPCmeLr2_0(.dout(w_dff_A_0MA9bC231_0),.din(w_dff_A_VwPCmeLr2_0),.clk(gclk));
	jdff dff_A_0MA9bC231_0(.dout(w_dff_A_aswn5hTa0_0),.din(w_dff_A_0MA9bC231_0),.clk(gclk));
	jdff dff_A_aswn5hTa0_0(.dout(w_dff_A_8e8HGB357_0),.din(w_dff_A_aswn5hTa0_0),.clk(gclk));
	jdff dff_A_8e8HGB357_0(.dout(w_dff_A_dKqdSLq24_0),.din(w_dff_A_8e8HGB357_0),.clk(gclk));
	jdff dff_A_dKqdSLq24_0(.dout(G822),.din(w_dff_A_dKqdSLq24_0),.clk(gclk));
	jdff dff_A_VFIEsrzx7_1(.dout(w_dff_A_Kk1amslp4_0),.din(w_dff_A_VFIEsrzx7_1),.clk(gclk));
	jdff dff_A_Kk1amslp4_0(.dout(w_dff_A_ctHwxDA26_0),.din(w_dff_A_Kk1amslp4_0),.clk(gclk));
	jdff dff_A_ctHwxDA26_0(.dout(w_dff_A_fL1uaJKE5_0),.din(w_dff_A_ctHwxDA26_0),.clk(gclk));
	jdff dff_A_fL1uaJKE5_0(.dout(w_dff_A_sgJBLYAJ9_0),.din(w_dff_A_fL1uaJKE5_0),.clk(gclk));
	jdff dff_A_sgJBLYAJ9_0(.dout(w_dff_A_DKCyW6pd8_0),.din(w_dff_A_sgJBLYAJ9_0),.clk(gclk));
	jdff dff_A_DKCyW6pd8_0(.dout(w_dff_A_8vlTKZo39_0),.din(w_dff_A_DKCyW6pd8_0),.clk(gclk));
	jdff dff_A_8vlTKZo39_0(.dout(w_dff_A_Vb3Fqu1d0_0),.din(w_dff_A_8vlTKZo39_0),.clk(gclk));
	jdff dff_A_Vb3Fqu1d0_0(.dout(w_dff_A_4mvlN60C0_0),.din(w_dff_A_Vb3Fqu1d0_0),.clk(gclk));
	jdff dff_A_4mvlN60C0_0(.dout(w_dff_A_9QQMqnPi6_0),.din(w_dff_A_4mvlN60C0_0),.clk(gclk));
	jdff dff_A_9QQMqnPi6_0(.dout(w_dff_A_XN0SEcMI0_0),.din(w_dff_A_9QQMqnPi6_0),.clk(gclk));
	jdff dff_A_XN0SEcMI0_0(.dout(w_dff_A_L97a1K454_0),.din(w_dff_A_XN0SEcMI0_0),.clk(gclk));
	jdff dff_A_L97a1K454_0(.dout(w_dff_A_azqoZSDg4_0),.din(w_dff_A_L97a1K454_0),.clk(gclk));
	jdff dff_A_azqoZSDg4_0(.dout(w_dff_A_VpMHyHyO1_0),.din(w_dff_A_azqoZSDg4_0),.clk(gclk));
	jdff dff_A_VpMHyHyO1_0(.dout(w_dff_A_LMHIKbp41_0),.din(w_dff_A_VpMHyHyO1_0),.clk(gclk));
	jdff dff_A_LMHIKbp41_0(.dout(G838),.din(w_dff_A_LMHIKbp41_0),.clk(gclk));
	jdff dff_A_ZyftNr317_1(.dout(w_dff_A_3untLjXb5_0),.din(w_dff_A_ZyftNr317_1),.clk(gclk));
	jdff dff_A_3untLjXb5_0(.dout(w_dff_A_SqPFw5wX7_0),.din(w_dff_A_3untLjXb5_0),.clk(gclk));
	jdff dff_A_SqPFw5wX7_0(.dout(w_dff_A_0IjxmDpF6_0),.din(w_dff_A_SqPFw5wX7_0),.clk(gclk));
	jdff dff_A_0IjxmDpF6_0(.dout(w_dff_A_wlmcdczE0_0),.din(w_dff_A_0IjxmDpF6_0),.clk(gclk));
	jdff dff_A_wlmcdczE0_0(.dout(w_dff_A_v0pAfD2J4_0),.din(w_dff_A_wlmcdczE0_0),.clk(gclk));
	jdff dff_A_v0pAfD2J4_0(.dout(w_dff_A_tAOAqvb11_0),.din(w_dff_A_v0pAfD2J4_0),.clk(gclk));
	jdff dff_A_tAOAqvb11_0(.dout(w_dff_A_cFNv92mf3_0),.din(w_dff_A_tAOAqvb11_0),.clk(gclk));
	jdff dff_A_cFNv92mf3_0(.dout(w_dff_A_h0Tjdrh89_0),.din(w_dff_A_cFNv92mf3_0),.clk(gclk));
	jdff dff_A_h0Tjdrh89_0(.dout(w_dff_A_serLEDNa0_0),.din(w_dff_A_h0Tjdrh89_0),.clk(gclk));
	jdff dff_A_serLEDNa0_0(.dout(w_dff_A_1IB063gI7_0),.din(w_dff_A_serLEDNa0_0),.clk(gclk));
	jdff dff_A_1IB063gI7_0(.dout(w_dff_A_WGlETsiS5_0),.din(w_dff_A_1IB063gI7_0),.clk(gclk));
	jdff dff_A_WGlETsiS5_0(.dout(w_dff_A_UPp9Vnop8_0),.din(w_dff_A_WGlETsiS5_0),.clk(gclk));
	jdff dff_A_UPp9Vnop8_0(.dout(w_dff_A_MeRrixpo5_0),.din(w_dff_A_UPp9Vnop8_0),.clk(gclk));
	jdff dff_A_MeRrixpo5_0(.dout(w_dff_A_7vHO491q0_0),.din(w_dff_A_MeRrixpo5_0),.clk(gclk));
	jdff dff_A_7vHO491q0_0(.dout(w_dff_A_1TnEsA7g0_0),.din(w_dff_A_7vHO491q0_0),.clk(gclk));
	jdff dff_A_1TnEsA7g0_0(.dout(w_dff_A_1grLQ4el5_0),.din(w_dff_A_1TnEsA7g0_0),.clk(gclk));
	jdff dff_A_1grLQ4el5_0(.dout(w_dff_A_6IdK8xAF1_0),.din(w_dff_A_1grLQ4el5_0),.clk(gclk));
	jdff dff_A_6IdK8xAF1_0(.dout(G861),.din(w_dff_A_6IdK8xAF1_0),.clk(gclk));
	jdff dff_A_mtoJbP4h4_1(.dout(w_dff_A_nvCzGaTf6_0),.din(w_dff_A_mtoJbP4h4_1),.clk(gclk));
	jdff dff_A_nvCzGaTf6_0(.dout(w_dff_A_9EtarGos9_0),.din(w_dff_A_nvCzGaTf6_0),.clk(gclk));
	jdff dff_A_9EtarGos9_0(.dout(w_dff_A_VEDWxJV33_0),.din(w_dff_A_9EtarGos9_0),.clk(gclk));
	jdff dff_A_VEDWxJV33_0(.dout(w_dff_A_vhvYq4SF9_0),.din(w_dff_A_VEDWxJV33_0),.clk(gclk));
	jdff dff_A_vhvYq4SF9_0(.dout(w_dff_A_SkpyfsEZ7_0),.din(w_dff_A_vhvYq4SF9_0),.clk(gclk));
	jdff dff_A_SkpyfsEZ7_0(.dout(w_dff_A_7ngbVZOH2_0),.din(w_dff_A_SkpyfsEZ7_0),.clk(gclk));
	jdff dff_A_7ngbVZOH2_0(.dout(w_dff_A_gQkpQBel8_0),.din(w_dff_A_7ngbVZOH2_0),.clk(gclk));
	jdff dff_A_gQkpQBel8_0(.dout(w_dff_A_nf7oNB5I5_0),.din(w_dff_A_gQkpQBel8_0),.clk(gclk));
	jdff dff_A_nf7oNB5I5_0(.dout(w_dff_A_Kism8BVd5_0),.din(w_dff_A_nf7oNB5I5_0),.clk(gclk));
	jdff dff_A_Kism8BVd5_0(.dout(G623),.din(w_dff_A_Kism8BVd5_0),.clk(gclk));
	jdff dff_A_CgLAglrU8_2(.dout(w_dff_A_LXK5wWH77_0),.din(w_dff_A_CgLAglrU8_2),.clk(gclk));
	jdff dff_A_LXK5wWH77_0(.dout(w_dff_A_79ufvbh97_0),.din(w_dff_A_LXK5wWH77_0),.clk(gclk));
	jdff dff_A_79ufvbh97_0(.dout(w_dff_A_RZAVZjJD8_0),.din(w_dff_A_79ufvbh97_0),.clk(gclk));
	jdff dff_A_RZAVZjJD8_0(.dout(w_dff_A_kqVTFC2E8_0),.din(w_dff_A_RZAVZjJD8_0),.clk(gclk));
	jdff dff_A_kqVTFC2E8_0(.dout(w_dff_A_8jBoo9gs0_0),.din(w_dff_A_kqVTFC2E8_0),.clk(gclk));
	jdff dff_A_8jBoo9gs0_0(.dout(w_dff_A_kwk7g0yc3_0),.din(w_dff_A_8jBoo9gs0_0),.clk(gclk));
	jdff dff_A_kwk7g0yc3_0(.dout(w_dff_A_0jQu3geu3_0),.din(w_dff_A_kwk7g0yc3_0),.clk(gclk));
	jdff dff_A_0jQu3geu3_0(.dout(w_dff_A_JerQidNt3_0),.din(w_dff_A_0jQu3geu3_0),.clk(gclk));
	jdff dff_A_JerQidNt3_0(.dout(w_dff_A_PV84EtTp6_0),.din(w_dff_A_JerQidNt3_0),.clk(gclk));
	jdff dff_A_PV84EtTp6_0(.dout(w_dff_A_dedbp4CL7_0),.din(w_dff_A_PV84EtTp6_0),.clk(gclk));
	jdff dff_A_dedbp4CL7_0(.dout(w_dff_A_dXcX4MYR2_0),.din(w_dff_A_dedbp4CL7_0),.clk(gclk));
	jdff dff_A_dXcX4MYR2_0(.dout(w_dff_A_IyEev7oO5_0),.din(w_dff_A_dXcX4MYR2_0),.clk(gclk));
	jdff dff_A_IyEev7oO5_0(.dout(w_dff_A_Pk0pOnrI0_0),.din(w_dff_A_IyEev7oO5_0),.clk(gclk));
	jdff dff_A_Pk0pOnrI0_0(.dout(G722),.din(w_dff_A_Pk0pOnrI0_0),.clk(gclk));
	jdff dff_A_0TreeCMY9_1(.dout(w_dff_A_jCdOdkov6_0),.din(w_dff_A_0TreeCMY9_1),.clk(gclk));
	jdff dff_A_jCdOdkov6_0(.dout(w_dff_A_mu3R57fZ9_0),.din(w_dff_A_jCdOdkov6_0),.clk(gclk));
	jdff dff_A_mu3R57fZ9_0(.dout(w_dff_A_5kOFeQuL7_0),.din(w_dff_A_mu3R57fZ9_0),.clk(gclk));
	jdff dff_A_5kOFeQuL7_0(.dout(w_dff_A_g44jRxw19_0),.din(w_dff_A_5kOFeQuL7_0),.clk(gclk));
	jdff dff_A_g44jRxw19_0(.dout(w_dff_A_3WNorKJD9_0),.din(w_dff_A_g44jRxw19_0),.clk(gclk));
	jdff dff_A_3WNorKJD9_0(.dout(w_dff_A_HDw7VX9D5_0),.din(w_dff_A_3WNorKJD9_0),.clk(gclk));
	jdff dff_A_HDw7VX9D5_0(.dout(w_dff_A_mK8JQec03_0),.din(w_dff_A_HDw7VX9D5_0),.clk(gclk));
	jdff dff_A_mK8JQec03_0(.dout(w_dff_A_T5qYpt4V1_0),.din(w_dff_A_mK8JQec03_0),.clk(gclk));
	jdff dff_A_T5qYpt4V1_0(.dout(w_dff_A_fOoMB7R01_0),.din(w_dff_A_T5qYpt4V1_0),.clk(gclk));
	jdff dff_A_fOoMB7R01_0(.dout(w_dff_A_i4N3sXmR0_0),.din(w_dff_A_fOoMB7R01_0),.clk(gclk));
	jdff dff_A_i4N3sXmR0_0(.dout(w_dff_A_tqhg0jtD8_0),.din(w_dff_A_i4N3sXmR0_0),.clk(gclk));
	jdff dff_A_tqhg0jtD8_0(.dout(w_dff_A_bJ2UM7v22_0),.din(w_dff_A_tqhg0jtD8_0),.clk(gclk));
	jdff dff_A_bJ2UM7v22_0(.dout(G832),.din(w_dff_A_bJ2UM7v22_0),.clk(gclk));
	jdff dff_A_aRP8PpQw1_1(.dout(w_dff_A_xoxA61ev1_0),.din(w_dff_A_aRP8PpQw1_1),.clk(gclk));
	jdff dff_A_xoxA61ev1_0(.dout(w_dff_A_l8BlxnMc0_0),.din(w_dff_A_xoxA61ev1_0),.clk(gclk));
	jdff dff_A_l8BlxnMc0_0(.dout(w_dff_A_8Wb5QN4C9_0),.din(w_dff_A_l8BlxnMc0_0),.clk(gclk));
	jdff dff_A_8Wb5QN4C9_0(.dout(w_dff_A_imF7gaFM1_0),.din(w_dff_A_8Wb5QN4C9_0),.clk(gclk));
	jdff dff_A_imF7gaFM1_0(.dout(w_dff_A_sc6v5Ou48_0),.din(w_dff_A_imF7gaFM1_0),.clk(gclk));
	jdff dff_A_sc6v5Ou48_0(.dout(w_dff_A_t9rMzcAm4_0),.din(w_dff_A_sc6v5Ou48_0),.clk(gclk));
	jdff dff_A_t9rMzcAm4_0(.dout(w_dff_A_5b7lwdYk7_0),.din(w_dff_A_t9rMzcAm4_0),.clk(gclk));
	jdff dff_A_5b7lwdYk7_0(.dout(w_dff_A_5857ocSk5_0),.din(w_dff_A_5b7lwdYk7_0),.clk(gclk));
	jdff dff_A_5857ocSk5_0(.dout(w_dff_A_rNpGfDUn0_0),.din(w_dff_A_5857ocSk5_0),.clk(gclk));
	jdff dff_A_rNpGfDUn0_0(.dout(w_dff_A_yIjaXRsn3_0),.din(w_dff_A_rNpGfDUn0_0),.clk(gclk));
	jdff dff_A_yIjaXRsn3_0(.dout(w_dff_A_5i0K9DG29_0),.din(w_dff_A_yIjaXRsn3_0),.clk(gclk));
	jdff dff_A_5i0K9DG29_0(.dout(w_dff_A_rNxl7Uz86_0),.din(w_dff_A_5i0K9DG29_0),.clk(gclk));
	jdff dff_A_rNxl7Uz86_0(.dout(w_dff_A_O7iZCGfN9_0),.din(w_dff_A_rNxl7Uz86_0),.clk(gclk));
	jdff dff_A_O7iZCGfN9_0(.dout(G834),.din(w_dff_A_O7iZCGfN9_0),.clk(gclk));
	jdff dff_A_cWVz6Ubw9_1(.dout(w_dff_A_gwtc3gQh9_0),.din(w_dff_A_cWVz6Ubw9_1),.clk(gclk));
	jdff dff_A_gwtc3gQh9_0(.dout(w_dff_A_1Yob8p3J1_0),.din(w_dff_A_gwtc3gQh9_0),.clk(gclk));
	jdff dff_A_1Yob8p3J1_0(.dout(w_dff_A_NDy6gCHK4_0),.din(w_dff_A_1Yob8p3J1_0),.clk(gclk));
	jdff dff_A_NDy6gCHK4_0(.dout(w_dff_A_yxZRWfcC9_0),.din(w_dff_A_NDy6gCHK4_0),.clk(gclk));
	jdff dff_A_yxZRWfcC9_0(.dout(w_dff_A_b2IEnacL4_0),.din(w_dff_A_yxZRWfcC9_0),.clk(gclk));
	jdff dff_A_b2IEnacL4_0(.dout(w_dff_A_DItqIM3H4_0),.din(w_dff_A_b2IEnacL4_0),.clk(gclk));
	jdff dff_A_DItqIM3H4_0(.dout(w_dff_A_fVD7jDbe1_0),.din(w_dff_A_DItqIM3H4_0),.clk(gclk));
	jdff dff_A_fVD7jDbe1_0(.dout(w_dff_A_AdOfJN4w4_0),.din(w_dff_A_fVD7jDbe1_0),.clk(gclk));
	jdff dff_A_AdOfJN4w4_0(.dout(w_dff_A_JfhjMLSu2_0),.din(w_dff_A_AdOfJN4w4_0),.clk(gclk));
	jdff dff_A_JfhjMLSu2_0(.dout(w_dff_A_KasOH0KW7_0),.din(w_dff_A_JfhjMLSu2_0),.clk(gclk));
	jdff dff_A_KasOH0KW7_0(.dout(w_dff_A_CcgIE2kV6_0),.din(w_dff_A_KasOH0KW7_0),.clk(gclk));
	jdff dff_A_CcgIE2kV6_0(.dout(w_dff_A_ROHbMZeR3_0),.din(w_dff_A_CcgIE2kV6_0),.clk(gclk));
	jdff dff_A_ROHbMZeR3_0(.dout(w_dff_A_q01qvI1b7_0),.din(w_dff_A_ROHbMZeR3_0),.clk(gclk));
	jdff dff_A_q01qvI1b7_0(.dout(w_dff_A_oAAEG4Qb2_0),.din(w_dff_A_q01qvI1b7_0),.clk(gclk));
	jdff dff_A_oAAEG4Qb2_0(.dout(w_dff_A_eB7LN01l1_0),.din(w_dff_A_oAAEG4Qb2_0),.clk(gclk));
	jdff dff_A_eB7LN01l1_0(.dout(G836),.din(w_dff_A_eB7LN01l1_0),.clk(gclk));
	jdff dff_A_WzDV50rL1_2(.dout(w_dff_A_1WQqNT460_0),.din(w_dff_A_WzDV50rL1_2),.clk(gclk));
	jdff dff_A_1WQqNT460_0(.dout(w_dff_A_SgEYbjjc6_0),.din(w_dff_A_1WQqNT460_0),.clk(gclk));
	jdff dff_A_SgEYbjjc6_0(.dout(w_dff_A_FZ8QYBHj0_0),.din(w_dff_A_SgEYbjjc6_0),.clk(gclk));
	jdff dff_A_FZ8QYBHj0_0(.dout(w_dff_A_xl0ZOeH14_0),.din(w_dff_A_FZ8QYBHj0_0),.clk(gclk));
	jdff dff_A_xl0ZOeH14_0(.dout(w_dff_A_zasEgTdG2_0),.din(w_dff_A_xl0ZOeH14_0),.clk(gclk));
	jdff dff_A_zasEgTdG2_0(.dout(w_dff_A_n72n2s850_0),.din(w_dff_A_zasEgTdG2_0),.clk(gclk));
	jdff dff_A_n72n2s850_0(.dout(w_dff_A_rHA126FP0_0),.din(w_dff_A_n72n2s850_0),.clk(gclk));
	jdff dff_A_rHA126FP0_0(.dout(w_dff_A_tb6ca8a54_0),.din(w_dff_A_rHA126FP0_0),.clk(gclk));
	jdff dff_A_tb6ca8a54_0(.dout(w_dff_A_vwET7jYv4_0),.din(w_dff_A_tb6ca8a54_0),.clk(gclk));
	jdff dff_A_vwET7jYv4_0(.dout(w_dff_A_xQ3aBGyg2_0),.din(w_dff_A_vwET7jYv4_0),.clk(gclk));
	jdff dff_A_xQ3aBGyg2_0(.dout(w_dff_A_NACuYeNd7_0),.din(w_dff_A_xQ3aBGyg2_0),.clk(gclk));
	jdff dff_A_NACuYeNd7_0(.dout(w_dff_A_MPnZkezm8_0),.din(w_dff_A_NACuYeNd7_0),.clk(gclk));
	jdff dff_A_MPnZkezm8_0(.dout(w_dff_A_PL5MABKR8_0),.din(w_dff_A_MPnZkezm8_0),.clk(gclk));
	jdff dff_A_PL5MABKR8_0(.dout(G859),.din(w_dff_A_PL5MABKR8_0),.clk(gclk));
	jdff dff_A_Xcf1pYNP1_1(.dout(w_dff_A_Xfb3PSfA2_0),.din(w_dff_A_Xcf1pYNP1_1),.clk(gclk));
	jdff dff_A_Xfb3PSfA2_0(.dout(w_dff_A_v0HqC36K5_0),.din(w_dff_A_Xfb3PSfA2_0),.clk(gclk));
	jdff dff_A_v0HqC36K5_0(.dout(w_dff_A_LQ0IBVtq5_0),.din(w_dff_A_v0HqC36K5_0),.clk(gclk));
	jdff dff_A_LQ0IBVtq5_0(.dout(w_dff_A_StdEhPuv8_0),.din(w_dff_A_LQ0IBVtq5_0),.clk(gclk));
	jdff dff_A_StdEhPuv8_0(.dout(w_dff_A_xxsUecIf7_0),.din(w_dff_A_StdEhPuv8_0),.clk(gclk));
	jdff dff_A_xxsUecIf7_0(.dout(w_dff_A_ydwbPhue5_0),.din(w_dff_A_xxsUecIf7_0),.clk(gclk));
	jdff dff_A_ydwbPhue5_0(.dout(w_dff_A_AsFgkaCG4_0),.din(w_dff_A_ydwbPhue5_0),.clk(gclk));
	jdff dff_A_AsFgkaCG4_0(.dout(w_dff_A_Vq00UK2h0_0),.din(w_dff_A_AsFgkaCG4_0),.clk(gclk));
	jdff dff_A_Vq00UK2h0_0(.dout(w_dff_A_ZG74mYlJ4_0),.din(w_dff_A_Vq00UK2h0_0),.clk(gclk));
	jdff dff_A_ZG74mYlJ4_0(.dout(w_dff_A_UH5QMYWn8_0),.din(w_dff_A_ZG74mYlJ4_0),.clk(gclk));
	jdff dff_A_UH5QMYWn8_0(.dout(w_dff_A_TmxGSpUR0_0),.din(w_dff_A_UH5QMYWn8_0),.clk(gclk));
	jdff dff_A_TmxGSpUR0_0(.dout(w_dff_A_kFOPrfOa3_0),.din(w_dff_A_TmxGSpUR0_0),.clk(gclk));
	jdff dff_A_kFOPrfOa3_0(.dout(G871),.din(w_dff_A_kFOPrfOa3_0),.clk(gclk));
	jdff dff_A_4fYXhbSz2_1(.dout(w_dff_A_4s2xqPvZ1_0),.din(w_dff_A_4fYXhbSz2_1),.clk(gclk));
	jdff dff_A_4s2xqPvZ1_0(.dout(w_dff_A_alSrChwX5_0),.din(w_dff_A_4s2xqPvZ1_0),.clk(gclk));
	jdff dff_A_alSrChwX5_0(.dout(w_dff_A_xKfg0DK49_0),.din(w_dff_A_alSrChwX5_0),.clk(gclk));
	jdff dff_A_xKfg0DK49_0(.dout(w_dff_A_CiNnPCiG6_0),.din(w_dff_A_xKfg0DK49_0),.clk(gclk));
	jdff dff_A_CiNnPCiG6_0(.dout(w_dff_A_w1ALeF1X6_0),.din(w_dff_A_CiNnPCiG6_0),.clk(gclk));
	jdff dff_A_w1ALeF1X6_0(.dout(w_dff_A_SDXx9UyQ6_0),.din(w_dff_A_w1ALeF1X6_0),.clk(gclk));
	jdff dff_A_SDXx9UyQ6_0(.dout(w_dff_A_FQLZYEwQ5_0),.din(w_dff_A_SDXx9UyQ6_0),.clk(gclk));
	jdff dff_A_FQLZYEwQ5_0(.dout(w_dff_A_7xFGPKkV4_0),.din(w_dff_A_FQLZYEwQ5_0),.clk(gclk));
	jdff dff_A_7xFGPKkV4_0(.dout(w_dff_A_H0OqcpjM6_0),.din(w_dff_A_7xFGPKkV4_0),.clk(gclk));
	jdff dff_A_H0OqcpjM6_0(.dout(w_dff_A_kDAT9Psb4_0),.din(w_dff_A_H0OqcpjM6_0),.clk(gclk));
	jdff dff_A_kDAT9Psb4_0(.dout(w_dff_A_WkFCRsQT1_0),.din(w_dff_A_kDAT9Psb4_0),.clk(gclk));
	jdff dff_A_WkFCRsQT1_0(.dout(w_dff_A_Rq35Tq8u4_0),.din(w_dff_A_WkFCRsQT1_0),.clk(gclk));
	jdff dff_A_Rq35Tq8u4_0(.dout(w_dff_A_5VGOjIgQ6_0),.din(w_dff_A_Rq35Tq8u4_0),.clk(gclk));
	jdff dff_A_5VGOjIgQ6_0(.dout(w_dff_A_uA1xalqg8_0),.din(w_dff_A_5VGOjIgQ6_0),.clk(gclk));
	jdff dff_A_uA1xalqg8_0(.dout(G873),.din(w_dff_A_uA1xalqg8_0),.clk(gclk));
	jdff dff_A_cecI00zW2_1(.dout(w_dff_A_a2OhQGic0_0),.din(w_dff_A_cecI00zW2_1),.clk(gclk));
	jdff dff_A_a2OhQGic0_0(.dout(w_dff_A_iiVW7oig7_0),.din(w_dff_A_a2OhQGic0_0),.clk(gclk));
	jdff dff_A_iiVW7oig7_0(.dout(w_dff_A_AR3vXfHt2_0),.din(w_dff_A_iiVW7oig7_0),.clk(gclk));
	jdff dff_A_AR3vXfHt2_0(.dout(w_dff_A_tIxfdXRJ4_0),.din(w_dff_A_AR3vXfHt2_0),.clk(gclk));
	jdff dff_A_tIxfdXRJ4_0(.dout(w_dff_A_QJIVTP0M3_0),.din(w_dff_A_tIxfdXRJ4_0),.clk(gclk));
	jdff dff_A_QJIVTP0M3_0(.dout(w_dff_A_sqkYLEe03_0),.din(w_dff_A_QJIVTP0M3_0),.clk(gclk));
	jdff dff_A_sqkYLEe03_0(.dout(w_dff_A_VO3EppYI0_0),.din(w_dff_A_sqkYLEe03_0),.clk(gclk));
	jdff dff_A_VO3EppYI0_0(.dout(w_dff_A_t097MXi33_0),.din(w_dff_A_VO3EppYI0_0),.clk(gclk));
	jdff dff_A_t097MXi33_0(.dout(w_dff_A_8tUlZekN8_0),.din(w_dff_A_t097MXi33_0),.clk(gclk));
	jdff dff_A_8tUlZekN8_0(.dout(w_dff_A_oXRdMPiV4_0),.din(w_dff_A_8tUlZekN8_0),.clk(gclk));
	jdff dff_A_oXRdMPiV4_0(.dout(w_dff_A_r8uGsviM5_0),.din(w_dff_A_oXRdMPiV4_0),.clk(gclk));
	jdff dff_A_r8uGsviM5_0(.dout(w_dff_A_HSH9YHwR7_0),.din(w_dff_A_r8uGsviM5_0),.clk(gclk));
	jdff dff_A_HSH9YHwR7_0(.dout(w_dff_A_yT8r4ESN7_0),.din(w_dff_A_HSH9YHwR7_0),.clk(gclk));
	jdff dff_A_yT8r4ESN7_0(.dout(w_dff_A_hoIEO0MO1_0),.din(w_dff_A_yT8r4ESN7_0),.clk(gclk));
	jdff dff_A_hoIEO0MO1_0(.dout(w_dff_A_5JvVsRDQ2_0),.din(w_dff_A_hoIEO0MO1_0),.clk(gclk));
	jdff dff_A_5JvVsRDQ2_0(.dout(G875),.din(w_dff_A_5JvVsRDQ2_0),.clk(gclk));
	jdff dff_A_j4wRy3eY7_1(.dout(w_dff_A_whizhFCe3_0),.din(w_dff_A_j4wRy3eY7_1),.clk(gclk));
	jdff dff_A_whizhFCe3_0(.dout(w_dff_A_32kIXURn1_0),.din(w_dff_A_whizhFCe3_0),.clk(gclk));
	jdff dff_A_32kIXURn1_0(.dout(w_dff_A_hBA4Sey01_0),.din(w_dff_A_32kIXURn1_0),.clk(gclk));
	jdff dff_A_hBA4Sey01_0(.dout(w_dff_A_obbFt1O36_0),.din(w_dff_A_hBA4Sey01_0),.clk(gclk));
	jdff dff_A_obbFt1O36_0(.dout(w_dff_A_VCaAMLQt7_0),.din(w_dff_A_obbFt1O36_0),.clk(gclk));
	jdff dff_A_VCaAMLQt7_0(.dout(w_dff_A_o6UflteS0_0),.din(w_dff_A_VCaAMLQt7_0),.clk(gclk));
	jdff dff_A_o6UflteS0_0(.dout(w_dff_A_X5EEzZRu3_0),.din(w_dff_A_o6UflteS0_0),.clk(gclk));
	jdff dff_A_X5EEzZRu3_0(.dout(w_dff_A_ThuzIoiq5_0),.din(w_dff_A_X5EEzZRu3_0),.clk(gclk));
	jdff dff_A_ThuzIoiq5_0(.dout(w_dff_A_hvssTaIL6_0),.din(w_dff_A_ThuzIoiq5_0),.clk(gclk));
	jdff dff_A_hvssTaIL6_0(.dout(w_dff_A_LGr9TRnY2_0),.din(w_dff_A_hvssTaIL6_0),.clk(gclk));
	jdff dff_A_LGr9TRnY2_0(.dout(w_dff_A_8zm7Iq9E2_0),.din(w_dff_A_LGr9TRnY2_0),.clk(gclk));
	jdff dff_A_8zm7Iq9E2_0(.dout(w_dff_A_7yQz3Z012_0),.din(w_dff_A_8zm7Iq9E2_0),.clk(gclk));
	jdff dff_A_7yQz3Z012_0(.dout(w_dff_A_vngx1fyN1_0),.din(w_dff_A_7yQz3Z012_0),.clk(gclk));
	jdff dff_A_vngx1fyN1_0(.dout(w_dff_A_YADLfDM62_0),.din(w_dff_A_vngx1fyN1_0),.clk(gclk));
	jdff dff_A_YADLfDM62_0(.dout(w_dff_A_tFxjjqFZ0_0),.din(w_dff_A_YADLfDM62_0),.clk(gclk));
	jdff dff_A_tFxjjqFZ0_0(.dout(w_dff_A_4uw0WhNL4_0),.din(w_dff_A_tFxjjqFZ0_0),.clk(gclk));
	jdff dff_A_4uw0WhNL4_0(.dout(G877),.din(w_dff_A_4uw0WhNL4_0),.clk(gclk));
	jdff dff_A_LDVmy6xf9_1(.dout(w_dff_A_DNhCCQWP5_0),.din(w_dff_A_LDVmy6xf9_1),.clk(gclk));
	jdff dff_A_DNhCCQWP5_0(.dout(w_dff_A_hHg4PhMJ7_0),.din(w_dff_A_DNhCCQWP5_0),.clk(gclk));
	jdff dff_A_hHg4PhMJ7_0(.dout(w_dff_A_Yki2C0eC2_0),.din(w_dff_A_hHg4PhMJ7_0),.clk(gclk));
	jdff dff_A_Yki2C0eC2_0(.dout(w_dff_A_DF6MiZSk7_0),.din(w_dff_A_Yki2C0eC2_0),.clk(gclk));
	jdff dff_A_DF6MiZSk7_0(.dout(w_dff_A_1DpJCtoK7_0),.din(w_dff_A_DF6MiZSk7_0),.clk(gclk));
	jdff dff_A_1DpJCtoK7_0(.dout(w_dff_A_UHiBLZ2m6_0),.din(w_dff_A_1DpJCtoK7_0),.clk(gclk));
	jdff dff_A_UHiBLZ2m6_0(.dout(w_dff_A_ohLDOpWV4_0),.din(w_dff_A_UHiBLZ2m6_0),.clk(gclk));
	jdff dff_A_ohLDOpWV4_0(.dout(w_dff_A_O7xkq8va3_0),.din(w_dff_A_ohLDOpWV4_0),.clk(gclk));
	jdff dff_A_O7xkq8va3_0(.dout(w_dff_A_VjHFoiEg1_0),.din(w_dff_A_O7xkq8va3_0),.clk(gclk));
	jdff dff_A_VjHFoiEg1_0(.dout(w_dff_A_Bu9c7gBV1_0),.din(w_dff_A_VjHFoiEg1_0),.clk(gclk));
	jdff dff_A_Bu9c7gBV1_0(.dout(w_dff_A_I3ofLbNy3_0),.din(w_dff_A_Bu9c7gBV1_0),.clk(gclk));
	jdff dff_A_I3ofLbNy3_0(.dout(w_dff_A_Df5wHkPL5_0),.din(w_dff_A_I3ofLbNy3_0),.clk(gclk));
	jdff dff_A_Df5wHkPL5_0(.dout(w_dff_A_s3xTOZCM8_0),.din(w_dff_A_Df5wHkPL5_0),.clk(gclk));
	jdff dff_A_s3xTOZCM8_0(.dout(w_dff_A_5lTxik1F7_0),.din(w_dff_A_s3xTOZCM8_0),.clk(gclk));
	jdff dff_A_5lTxik1F7_0(.dout(w_dff_A_0oScPgZE3_0),.din(w_dff_A_5lTxik1F7_0),.clk(gclk));
	jdff dff_A_0oScPgZE3_0(.dout(w_dff_A_os7iufY74_0),.din(w_dff_A_0oScPgZE3_0),.clk(gclk));
	jdff dff_A_os7iufY74_0(.dout(w_dff_A_zgFimIi60_0),.din(w_dff_A_os7iufY74_0),.clk(gclk));
	jdff dff_A_zgFimIi60_0(.dout(w_dff_A_5Omzibjx3_0),.din(w_dff_A_zgFimIi60_0),.clk(gclk));
	jdff dff_A_5Omzibjx3_0(.dout(w_dff_A_NDhWr5cn3_0),.din(w_dff_A_5Omzibjx3_0),.clk(gclk));
	jdff dff_A_NDhWr5cn3_0(.dout(G998),.din(w_dff_A_NDhWr5cn3_0),.clk(gclk));
	jdff dff_A_XFSPDDuF1_1(.dout(w_dff_A_Gyv3mvEr2_0),.din(w_dff_A_XFSPDDuF1_1),.clk(gclk));
	jdff dff_A_Gyv3mvEr2_0(.dout(w_dff_A_WPysNjOK6_0),.din(w_dff_A_Gyv3mvEr2_0),.clk(gclk));
	jdff dff_A_WPysNjOK6_0(.dout(w_dff_A_LJ2FMCiX4_0),.din(w_dff_A_WPysNjOK6_0),.clk(gclk));
	jdff dff_A_LJ2FMCiX4_0(.dout(w_dff_A_qalRgpAi5_0),.din(w_dff_A_LJ2FMCiX4_0),.clk(gclk));
	jdff dff_A_qalRgpAi5_0(.dout(w_dff_A_lRdXNXv91_0),.din(w_dff_A_qalRgpAi5_0),.clk(gclk));
	jdff dff_A_lRdXNXv91_0(.dout(w_dff_A_BhnySF2a4_0),.din(w_dff_A_lRdXNXv91_0),.clk(gclk));
	jdff dff_A_BhnySF2a4_0(.dout(w_dff_A_2KhPCSam7_0),.din(w_dff_A_BhnySF2a4_0),.clk(gclk));
	jdff dff_A_2KhPCSam7_0(.dout(w_dff_A_VpwJHiuj2_0),.din(w_dff_A_2KhPCSam7_0),.clk(gclk));
	jdff dff_A_VpwJHiuj2_0(.dout(w_dff_A_JwwS0Ze11_0),.din(w_dff_A_VpwJHiuj2_0),.clk(gclk));
	jdff dff_A_JwwS0Ze11_0(.dout(w_dff_A_rWcrur6b6_0),.din(w_dff_A_JwwS0Ze11_0),.clk(gclk));
	jdff dff_A_rWcrur6b6_0(.dout(w_dff_A_MvCoxQho3_0),.din(w_dff_A_rWcrur6b6_0),.clk(gclk));
	jdff dff_A_MvCoxQho3_0(.dout(w_dff_A_0lz9rzBO6_0),.din(w_dff_A_MvCoxQho3_0),.clk(gclk));
	jdff dff_A_0lz9rzBO6_0(.dout(w_dff_A_iariGLAp4_0),.din(w_dff_A_0lz9rzBO6_0),.clk(gclk));
	jdff dff_A_iariGLAp4_0(.dout(w_dff_A_sNCdhDWI2_0),.din(w_dff_A_iariGLAp4_0),.clk(gclk));
	jdff dff_A_sNCdhDWI2_0(.dout(w_dff_A_5OZwGQr93_0),.din(w_dff_A_sNCdhDWI2_0),.clk(gclk));
	jdff dff_A_5OZwGQr93_0(.dout(w_dff_A_90VmhJ6N4_0),.din(w_dff_A_5OZwGQr93_0),.clk(gclk));
	jdff dff_A_90VmhJ6N4_0(.dout(w_dff_A_rwzH8ctH0_0),.din(w_dff_A_90VmhJ6N4_0),.clk(gclk));
	jdff dff_A_rwzH8ctH0_0(.dout(w_dff_A_RYcuxKUY6_0),.din(w_dff_A_rwzH8ctH0_0),.clk(gclk));
	jdff dff_A_RYcuxKUY6_0(.dout(G1000),.din(w_dff_A_RYcuxKUY6_0),.clk(gclk));
	jdff dff_A_LojQ4O6a8_2(.dout(w_dff_A_fhRTsr0g6_0),.din(w_dff_A_LojQ4O6a8_2),.clk(gclk));
	jdff dff_A_fhRTsr0g6_0(.dout(w_dff_A_Qav62Bm62_0),.din(w_dff_A_fhRTsr0g6_0),.clk(gclk));
	jdff dff_A_Qav62Bm62_0(.dout(w_dff_A_choGXKAM6_0),.din(w_dff_A_Qav62Bm62_0),.clk(gclk));
	jdff dff_A_choGXKAM6_0(.dout(w_dff_A_cM2HiBzD5_0),.din(w_dff_A_choGXKAM6_0),.clk(gclk));
	jdff dff_A_cM2HiBzD5_0(.dout(w_dff_A_lD4PhfTP5_0),.din(w_dff_A_cM2HiBzD5_0),.clk(gclk));
	jdff dff_A_lD4PhfTP5_0(.dout(w_dff_A_aGlRU6By9_0),.din(w_dff_A_lD4PhfTP5_0),.clk(gclk));
	jdff dff_A_aGlRU6By9_0(.dout(w_dff_A_3qAT6j0y8_0),.din(w_dff_A_aGlRU6By9_0),.clk(gclk));
	jdff dff_A_3qAT6j0y8_0(.dout(G575),.din(w_dff_A_3qAT6j0y8_0),.clk(gclk));
	jdff dff_A_ifO26XYC5_2(.dout(w_dff_A_Ga7U7ueu8_0),.din(w_dff_A_ifO26XYC5_2),.clk(gclk));
	jdff dff_A_Ga7U7ueu8_0(.dout(w_dff_A_iADms8vr3_0),.din(w_dff_A_Ga7U7ueu8_0),.clk(gclk));
	jdff dff_A_iADms8vr3_0(.dout(w_dff_A_FI0QRrNN2_0),.din(w_dff_A_iADms8vr3_0),.clk(gclk));
	jdff dff_A_FI0QRrNN2_0(.dout(w_dff_A_kJ5MLS4y0_0),.din(w_dff_A_FI0QRrNN2_0),.clk(gclk));
	jdff dff_A_kJ5MLS4y0_0(.dout(w_dff_A_gP10RLMl1_0),.din(w_dff_A_kJ5MLS4y0_0),.clk(gclk));
	jdff dff_A_gP10RLMl1_0(.dout(w_dff_A_05DtLBpD9_0),.din(w_dff_A_gP10RLMl1_0),.clk(gclk));
	jdff dff_A_05DtLBpD9_0(.dout(G585),.din(w_dff_A_05DtLBpD9_0),.clk(gclk));
	jdff dff_A_FG5x9kcg6_2(.dout(w_dff_A_3KjLJqhc3_0),.din(w_dff_A_FG5x9kcg6_2),.clk(gclk));
	jdff dff_A_3KjLJqhc3_0(.dout(w_dff_A_pHWukCto8_0),.din(w_dff_A_3KjLJqhc3_0),.clk(gclk));
	jdff dff_A_pHWukCto8_0(.dout(w_dff_A_7wbJbWma3_0),.din(w_dff_A_pHWukCto8_0),.clk(gclk));
	jdff dff_A_7wbJbWma3_0(.dout(w_dff_A_tVUV7PH33_0),.din(w_dff_A_7wbJbWma3_0),.clk(gclk));
	jdff dff_A_tVUV7PH33_0(.dout(w_dff_A_369qkXKi3_0),.din(w_dff_A_tVUV7PH33_0),.clk(gclk));
	jdff dff_A_369qkXKi3_0(.dout(w_dff_A_aPrPoqpV4_0),.din(w_dff_A_369qkXKi3_0),.clk(gclk));
	jdff dff_A_aPrPoqpV4_0(.dout(w_dff_A_W9Vo4v9l8_0),.din(w_dff_A_aPrPoqpV4_0),.clk(gclk));
	jdff dff_A_W9Vo4v9l8_0(.dout(w_dff_A_saKgwT7n1_0),.din(w_dff_A_W9Vo4v9l8_0),.clk(gclk));
	jdff dff_A_saKgwT7n1_0(.dout(w_dff_A_WwXd2Wx76_0),.din(w_dff_A_saKgwT7n1_0),.clk(gclk));
	jdff dff_A_WwXd2Wx76_0(.dout(w_dff_A_HS5fnaWm6_0),.din(w_dff_A_WwXd2Wx76_0),.clk(gclk));
	jdff dff_A_HS5fnaWm6_0(.dout(w_dff_A_z5rDJbAn4_0),.din(w_dff_A_HS5fnaWm6_0),.clk(gclk));
	jdff dff_A_z5rDJbAn4_0(.dout(G661),.din(w_dff_A_z5rDJbAn4_0),.clk(gclk));
	jdff dff_A_JOmnUMds0_2(.dout(w_dff_A_ThLxdI1c2_0),.din(w_dff_A_JOmnUMds0_2),.clk(gclk));
	jdff dff_A_ThLxdI1c2_0(.dout(w_dff_A_CNOC1cE41_0),.din(w_dff_A_ThLxdI1c2_0),.clk(gclk));
	jdff dff_A_CNOC1cE41_0(.dout(w_dff_A_0FJgxq9G5_0),.din(w_dff_A_CNOC1cE41_0),.clk(gclk));
	jdff dff_A_0FJgxq9G5_0(.dout(w_dff_A_xdblaibq2_0),.din(w_dff_A_0FJgxq9G5_0),.clk(gclk));
	jdff dff_A_xdblaibq2_0(.dout(w_dff_A_o9EvYuQR7_0),.din(w_dff_A_xdblaibq2_0),.clk(gclk));
	jdff dff_A_o9EvYuQR7_0(.dout(w_dff_A_3SdChd5U6_0),.din(w_dff_A_o9EvYuQR7_0),.clk(gclk));
	jdff dff_A_3SdChd5U6_0(.dout(w_dff_A_ZP9E1GS63_0),.din(w_dff_A_3SdChd5U6_0),.clk(gclk));
	jdff dff_A_ZP9E1GS63_0(.dout(w_dff_A_6k6qiJuN0_0),.din(w_dff_A_ZP9E1GS63_0),.clk(gclk));
	jdff dff_A_6k6qiJuN0_0(.dout(w_dff_A_S8u6oNdq2_0),.din(w_dff_A_6k6qiJuN0_0),.clk(gclk));
	jdff dff_A_S8u6oNdq2_0(.dout(w_dff_A_REeoh9Ix1_0),.din(w_dff_A_S8u6oNdq2_0),.clk(gclk));
	jdff dff_A_REeoh9Ix1_0(.dout(w_dff_A_yZz67w788_0),.din(w_dff_A_REeoh9Ix1_0),.clk(gclk));
	jdff dff_A_yZz67w788_0(.dout(G693),.din(w_dff_A_yZz67w788_0),.clk(gclk));
	jdff dff_A_jqIyVt3z5_2(.dout(w_dff_A_a6w4mOZa7_0),.din(w_dff_A_jqIyVt3z5_2),.clk(gclk));
	jdff dff_A_a6w4mOZa7_0(.dout(w_dff_A_SU9TATiq3_0),.din(w_dff_A_a6w4mOZa7_0),.clk(gclk));
	jdff dff_A_SU9TATiq3_0(.dout(w_dff_A_os4xKN308_0),.din(w_dff_A_SU9TATiq3_0),.clk(gclk));
	jdff dff_A_os4xKN308_0(.dout(w_dff_A_7GXsRNkE0_0),.din(w_dff_A_os4xKN308_0),.clk(gclk));
	jdff dff_A_7GXsRNkE0_0(.dout(w_dff_A_6xhTyW7e6_0),.din(w_dff_A_7GXsRNkE0_0),.clk(gclk));
	jdff dff_A_6xhTyW7e6_0(.dout(w_dff_A_lWPPiM2p9_0),.din(w_dff_A_6xhTyW7e6_0),.clk(gclk));
	jdff dff_A_lWPPiM2p9_0(.dout(w_dff_A_PKe6noIS6_0),.din(w_dff_A_lWPPiM2p9_0),.clk(gclk));
	jdff dff_A_PKe6noIS6_0(.dout(G747),.din(w_dff_A_PKe6noIS6_0),.clk(gclk));
	jdff dff_A_BPQdP7vV4_2(.dout(w_dff_A_pV3GcW802_0),.din(w_dff_A_BPQdP7vV4_2),.clk(gclk));
	jdff dff_A_pV3GcW802_0(.dout(w_dff_A_aQaJ0lxD2_0),.din(w_dff_A_pV3GcW802_0),.clk(gclk));
	jdff dff_A_aQaJ0lxD2_0(.dout(w_dff_A_HOTC0lbI8_0),.din(w_dff_A_aQaJ0lxD2_0),.clk(gclk));
	jdff dff_A_HOTC0lbI8_0(.dout(w_dff_A_wC1FHTSu7_0),.din(w_dff_A_HOTC0lbI8_0),.clk(gclk));
	jdff dff_A_wC1FHTSu7_0(.dout(w_dff_A_AGE81Mej8_0),.din(w_dff_A_wC1FHTSu7_0),.clk(gclk));
	jdff dff_A_AGE81Mej8_0(.dout(w_dff_A_fmaFpMg28_0),.din(w_dff_A_AGE81Mej8_0),.clk(gclk));
	jdff dff_A_fmaFpMg28_0(.dout(w_dff_A_75YbuoFO9_0),.din(w_dff_A_fmaFpMg28_0),.clk(gclk));
	jdff dff_A_75YbuoFO9_0(.dout(w_dff_A_JZqJ9of82_0),.din(w_dff_A_75YbuoFO9_0),.clk(gclk));
	jdff dff_A_JZqJ9of82_0(.dout(G752),.din(w_dff_A_JZqJ9of82_0),.clk(gclk));
	jdff dff_A_D2cceXBm3_2(.dout(w_dff_A_aVQSBQqr3_0),.din(w_dff_A_D2cceXBm3_2),.clk(gclk));
	jdff dff_A_aVQSBQqr3_0(.dout(w_dff_A_ekpLxEU60_0),.din(w_dff_A_aVQSBQqr3_0),.clk(gclk));
	jdff dff_A_ekpLxEU60_0(.dout(w_dff_A_oXiNrvFE7_0),.din(w_dff_A_ekpLxEU60_0),.clk(gclk));
	jdff dff_A_oXiNrvFE7_0(.dout(w_dff_A_gztFXmxf0_0),.din(w_dff_A_oXiNrvFE7_0),.clk(gclk));
	jdff dff_A_gztFXmxf0_0(.dout(w_dff_A_ISA4hZLw1_0),.din(w_dff_A_gztFXmxf0_0),.clk(gclk));
	jdff dff_A_ISA4hZLw1_0(.dout(w_dff_A_cE3UymY29_0),.din(w_dff_A_ISA4hZLw1_0),.clk(gclk));
	jdff dff_A_cE3UymY29_0(.dout(w_dff_A_B0TYGzQ58_0),.din(w_dff_A_cE3UymY29_0),.clk(gclk));
	jdff dff_A_B0TYGzQ58_0(.dout(w_dff_A_ZpEqsrB63_0),.din(w_dff_A_B0TYGzQ58_0),.clk(gclk));
	jdff dff_A_ZpEqsrB63_0(.dout(w_dff_A_RmBYI8wY6_0),.din(w_dff_A_ZpEqsrB63_0),.clk(gclk));
	jdff dff_A_RmBYI8wY6_0(.dout(w_dff_A_Y6QgWCFW9_0),.din(w_dff_A_RmBYI8wY6_0),.clk(gclk));
	jdff dff_A_Y6QgWCFW9_0(.dout(G757),.din(w_dff_A_Y6QgWCFW9_0),.clk(gclk));
	jdff dff_A_AEoA2Y3E4_2(.dout(w_dff_A_GDke7ttV5_0),.din(w_dff_A_AEoA2Y3E4_2),.clk(gclk));
	jdff dff_A_GDke7ttV5_0(.dout(w_dff_A_O2XduvVY3_0),.din(w_dff_A_GDke7ttV5_0),.clk(gclk));
	jdff dff_A_O2XduvVY3_0(.dout(w_dff_A_GWzhwAwj9_0),.din(w_dff_A_O2XduvVY3_0),.clk(gclk));
	jdff dff_A_GWzhwAwj9_0(.dout(w_dff_A_yVCUwG0X9_0),.din(w_dff_A_GWzhwAwj9_0),.clk(gclk));
	jdff dff_A_yVCUwG0X9_0(.dout(w_dff_A_lrXr0hMv8_0),.din(w_dff_A_yVCUwG0X9_0),.clk(gclk));
	jdff dff_A_lrXr0hMv8_0(.dout(w_dff_A_GVenb3qR0_0),.din(w_dff_A_lrXr0hMv8_0),.clk(gclk));
	jdff dff_A_GVenb3qR0_0(.dout(w_dff_A_1OVXuacQ4_0),.din(w_dff_A_GVenb3qR0_0),.clk(gclk));
	jdff dff_A_1OVXuacQ4_0(.dout(w_dff_A_iAcPN2iP0_0),.din(w_dff_A_1OVXuacQ4_0),.clk(gclk));
	jdff dff_A_iAcPN2iP0_0(.dout(w_dff_A_5nsuGzt59_0),.din(w_dff_A_iAcPN2iP0_0),.clk(gclk));
	jdff dff_A_5nsuGzt59_0(.dout(G762),.din(w_dff_A_5nsuGzt59_0),.clk(gclk));
	jdff dff_A_0GA9B52D4_2(.dout(w_dff_A_7OUcHV2K3_0),.din(w_dff_A_0GA9B52D4_2),.clk(gclk));
	jdff dff_A_7OUcHV2K3_0(.dout(w_dff_A_SoXXNMqx1_0),.din(w_dff_A_7OUcHV2K3_0),.clk(gclk));
	jdff dff_A_SoXXNMqx1_0(.dout(w_dff_A_PWbcLNIh1_0),.din(w_dff_A_SoXXNMqx1_0),.clk(gclk));
	jdff dff_A_PWbcLNIh1_0(.dout(w_dff_A_zVF2CYju0_0),.din(w_dff_A_PWbcLNIh1_0),.clk(gclk));
	jdff dff_A_zVF2CYju0_0(.dout(w_dff_A_hIXASEkO7_0),.din(w_dff_A_zVF2CYju0_0),.clk(gclk));
	jdff dff_A_hIXASEkO7_0(.dout(w_dff_A_nSZhUOqs9_0),.din(w_dff_A_hIXASEkO7_0),.clk(gclk));
	jdff dff_A_nSZhUOqs9_0(.dout(w_dff_A_8ooaBXL27_0),.din(w_dff_A_nSZhUOqs9_0),.clk(gclk));
	jdff dff_A_8ooaBXL27_0(.dout(G787),.din(w_dff_A_8ooaBXL27_0),.clk(gclk));
	jdff dff_A_PIbZeKxV2_2(.dout(w_dff_A_UeU8kFsv7_0),.din(w_dff_A_PIbZeKxV2_2),.clk(gclk));
	jdff dff_A_UeU8kFsv7_0(.dout(w_dff_A_ANrpXbpp0_0),.din(w_dff_A_UeU8kFsv7_0),.clk(gclk));
	jdff dff_A_ANrpXbpp0_0(.dout(w_dff_A_nmSiswmL9_0),.din(w_dff_A_ANrpXbpp0_0),.clk(gclk));
	jdff dff_A_nmSiswmL9_0(.dout(w_dff_A_cbSy4NbF0_0),.din(w_dff_A_nmSiswmL9_0),.clk(gclk));
	jdff dff_A_cbSy4NbF0_0(.dout(w_dff_A_JbQS280h0_0),.din(w_dff_A_cbSy4NbF0_0),.clk(gclk));
	jdff dff_A_JbQS280h0_0(.dout(w_dff_A_GJdXwLX77_0),.din(w_dff_A_JbQS280h0_0),.clk(gclk));
	jdff dff_A_GJdXwLX77_0(.dout(w_dff_A_0p93KERt6_0),.din(w_dff_A_GJdXwLX77_0),.clk(gclk));
	jdff dff_A_0p93KERt6_0(.dout(w_dff_A_im0l4GSm8_0),.din(w_dff_A_0p93KERt6_0),.clk(gclk));
	jdff dff_A_im0l4GSm8_0(.dout(G792),.din(w_dff_A_im0l4GSm8_0),.clk(gclk));
	jdff dff_A_ARx0zPuV9_2(.dout(w_dff_A_3oykOsDX5_0),.din(w_dff_A_ARx0zPuV9_2),.clk(gclk));
	jdff dff_A_3oykOsDX5_0(.dout(w_dff_A_4aWo7xLC6_0),.din(w_dff_A_3oykOsDX5_0),.clk(gclk));
	jdff dff_A_4aWo7xLC6_0(.dout(w_dff_A_KLBQhzhK4_0),.din(w_dff_A_4aWo7xLC6_0),.clk(gclk));
	jdff dff_A_KLBQhzhK4_0(.dout(w_dff_A_pNQ4GnV84_0),.din(w_dff_A_KLBQhzhK4_0),.clk(gclk));
	jdff dff_A_pNQ4GnV84_0(.dout(w_dff_A_VI5K4YOW2_0),.din(w_dff_A_pNQ4GnV84_0),.clk(gclk));
	jdff dff_A_VI5K4YOW2_0(.dout(w_dff_A_Tr6O11BU3_0),.din(w_dff_A_VI5K4YOW2_0),.clk(gclk));
	jdff dff_A_Tr6O11BU3_0(.dout(w_dff_A_sCvOXCik8_0),.din(w_dff_A_Tr6O11BU3_0),.clk(gclk));
	jdff dff_A_sCvOXCik8_0(.dout(w_dff_A_xWsBFvJe6_0),.din(w_dff_A_sCvOXCik8_0),.clk(gclk));
	jdff dff_A_xWsBFvJe6_0(.dout(w_dff_A_eyJRHqdw6_0),.din(w_dff_A_xWsBFvJe6_0),.clk(gclk));
	jdff dff_A_eyJRHqdw6_0(.dout(w_dff_A_cf8GP5E74_0),.din(w_dff_A_eyJRHqdw6_0),.clk(gclk));
	jdff dff_A_cf8GP5E74_0(.dout(G797),.din(w_dff_A_cf8GP5E74_0),.clk(gclk));
	jdff dff_A_ViDIITJZ5_2(.dout(w_dff_A_7BmhX4q84_0),.din(w_dff_A_ViDIITJZ5_2),.clk(gclk));
	jdff dff_A_7BmhX4q84_0(.dout(w_dff_A_VQQhsHgK0_0),.din(w_dff_A_7BmhX4q84_0),.clk(gclk));
	jdff dff_A_VQQhsHgK0_0(.dout(w_dff_A_xXm3HKaJ6_0),.din(w_dff_A_VQQhsHgK0_0),.clk(gclk));
	jdff dff_A_xXm3HKaJ6_0(.dout(w_dff_A_G9QnRSkN4_0),.din(w_dff_A_xXm3HKaJ6_0),.clk(gclk));
	jdff dff_A_G9QnRSkN4_0(.dout(w_dff_A_nu3dZDVW2_0),.din(w_dff_A_G9QnRSkN4_0),.clk(gclk));
	jdff dff_A_nu3dZDVW2_0(.dout(w_dff_A_q10fcxTz1_0),.din(w_dff_A_nu3dZDVW2_0),.clk(gclk));
	jdff dff_A_q10fcxTz1_0(.dout(w_dff_A_TPVfqmyn0_0),.din(w_dff_A_q10fcxTz1_0),.clk(gclk));
	jdff dff_A_TPVfqmyn0_0(.dout(w_dff_A_W7Q6ycmE1_0),.din(w_dff_A_TPVfqmyn0_0),.clk(gclk));
	jdff dff_A_W7Q6ycmE1_0(.dout(w_dff_A_1RimJmaU4_0),.din(w_dff_A_W7Q6ycmE1_0),.clk(gclk));
	jdff dff_A_1RimJmaU4_0(.dout(G802),.din(w_dff_A_1RimJmaU4_0),.clk(gclk));
	jdff dff_A_WJMGnPZm5_2(.dout(w_dff_A_jNVhEOKB2_0),.din(w_dff_A_WJMGnPZm5_2),.clk(gclk));
	jdff dff_A_jNVhEOKB2_0(.dout(w_dff_A_9twF5CGM4_0),.din(w_dff_A_jNVhEOKB2_0),.clk(gclk));
	jdff dff_A_9twF5CGM4_0(.dout(w_dff_A_GkN6wtgT7_0),.din(w_dff_A_9twF5CGM4_0),.clk(gclk));
	jdff dff_A_GkN6wtgT7_0(.dout(w_dff_A_aSumYti10_0),.din(w_dff_A_GkN6wtgT7_0),.clk(gclk));
	jdff dff_A_aSumYti10_0(.dout(w_dff_A_KcoZXFZX4_0),.din(w_dff_A_aSumYti10_0),.clk(gclk));
	jdff dff_A_KcoZXFZX4_0(.dout(w_dff_A_SSNmn5mZ1_0),.din(w_dff_A_KcoZXFZX4_0),.clk(gclk));
	jdff dff_A_SSNmn5mZ1_0(.dout(G642),.din(w_dff_A_SSNmn5mZ1_0),.clk(gclk));
	jdff dff_A_3gh9jhrR8_2(.dout(w_dff_A_rygam42w0_0),.din(w_dff_A_3gh9jhrR8_2),.clk(gclk));
	jdff dff_A_rygam42w0_0(.dout(w_dff_A_d0Tv3I3B3_0),.din(w_dff_A_rygam42w0_0),.clk(gclk));
	jdff dff_A_d0Tv3I3B3_0(.dout(w_dff_A_KsLV205o3_0),.din(w_dff_A_d0Tv3I3B3_0),.clk(gclk));
	jdff dff_A_KsLV205o3_0(.dout(w_dff_A_Ks4nR7gK1_0),.din(w_dff_A_KsLV205o3_0),.clk(gclk));
	jdff dff_A_Ks4nR7gK1_0(.dout(w_dff_A_3roPNQ8t0_0),.din(w_dff_A_Ks4nR7gK1_0),.clk(gclk));
	jdff dff_A_3roPNQ8t0_0(.dout(w_dff_A_8lQwb43X2_0),.din(w_dff_A_3roPNQ8t0_0),.clk(gclk));
	jdff dff_A_8lQwb43X2_0(.dout(w_dff_A_1VW3DmDd3_0),.din(w_dff_A_8lQwb43X2_0),.clk(gclk));
	jdff dff_A_1VW3DmDd3_0(.dout(w_dff_A_swGinSef6_0),.din(w_dff_A_1VW3DmDd3_0),.clk(gclk));
	jdff dff_A_swGinSef6_0(.dout(w_dff_A_1uBpjeJa9_0),.din(w_dff_A_swGinSef6_0),.clk(gclk));
	jdff dff_A_1uBpjeJa9_0(.dout(G664),.din(w_dff_A_1uBpjeJa9_0),.clk(gclk));
	jdff dff_A_JYKdF5A27_2(.dout(w_dff_A_criGi8qa7_0),.din(w_dff_A_JYKdF5A27_2),.clk(gclk));
	jdff dff_A_criGi8qa7_0(.dout(w_dff_A_qGQ1eYVr5_0),.din(w_dff_A_criGi8qa7_0),.clk(gclk));
	jdff dff_A_qGQ1eYVr5_0(.dout(w_dff_A_UnQd9nmp9_0),.din(w_dff_A_qGQ1eYVr5_0),.clk(gclk));
	jdff dff_A_UnQd9nmp9_0(.dout(w_dff_A_2da2ZqQE7_0),.din(w_dff_A_UnQd9nmp9_0),.clk(gclk));
	jdff dff_A_2da2ZqQE7_0(.dout(w_dff_A_2c9eMvlY4_0),.din(w_dff_A_2da2ZqQE7_0),.clk(gclk));
	jdff dff_A_2c9eMvlY4_0(.dout(w_dff_A_3oWSqGQX5_0),.din(w_dff_A_2c9eMvlY4_0),.clk(gclk));
	jdff dff_A_3oWSqGQX5_0(.dout(w_dff_A_a0QAE0996_0),.din(w_dff_A_3oWSqGQX5_0),.clk(gclk));
	jdff dff_A_a0QAE0996_0(.dout(w_dff_A_TipkdRtq8_0),.din(w_dff_A_a0QAE0996_0),.clk(gclk));
	jdff dff_A_TipkdRtq8_0(.dout(w_dff_A_F4nNpyMV2_0),.din(w_dff_A_TipkdRtq8_0),.clk(gclk));
	jdff dff_A_F4nNpyMV2_0(.dout(G667),.din(w_dff_A_F4nNpyMV2_0),.clk(gclk));
	jdff dff_A_N23fx6Y26_2(.dout(w_dff_A_MZIpwCEs1_0),.din(w_dff_A_N23fx6Y26_2),.clk(gclk));
	jdff dff_A_MZIpwCEs1_0(.dout(w_dff_A_4i2XggU13_0),.din(w_dff_A_MZIpwCEs1_0),.clk(gclk));
	jdff dff_A_4i2XggU13_0(.dout(w_dff_A_DqHzC5t82_0),.din(w_dff_A_4i2XggU13_0),.clk(gclk));
	jdff dff_A_DqHzC5t82_0(.dout(w_dff_A_yKAQ5gaz3_0),.din(w_dff_A_DqHzC5t82_0),.clk(gclk));
	jdff dff_A_yKAQ5gaz3_0(.dout(w_dff_A_xjGl09qk2_0),.din(w_dff_A_yKAQ5gaz3_0),.clk(gclk));
	jdff dff_A_xjGl09qk2_0(.dout(w_dff_A_nNcdRbdL0_0),.din(w_dff_A_xjGl09qk2_0),.clk(gclk));
	jdff dff_A_nNcdRbdL0_0(.dout(w_dff_A_KQ3abjVD8_0),.din(w_dff_A_nNcdRbdL0_0),.clk(gclk));
	jdff dff_A_KQ3abjVD8_0(.dout(w_dff_A_DbzolyGj5_0),.din(w_dff_A_KQ3abjVD8_0),.clk(gclk));
	jdff dff_A_DbzolyGj5_0(.dout(G670),.din(w_dff_A_DbzolyGj5_0),.clk(gclk));
	jdff dff_A_1W05j3Ma7_2(.dout(w_dff_A_HczZGVG62_0),.din(w_dff_A_1W05j3Ma7_2),.clk(gclk));
	jdff dff_A_HczZGVG62_0(.dout(w_dff_A_ypFB5xwd2_0),.din(w_dff_A_HczZGVG62_0),.clk(gclk));
	jdff dff_A_ypFB5xwd2_0(.dout(w_dff_A_VJxtsCrL3_0),.din(w_dff_A_ypFB5xwd2_0),.clk(gclk));
	jdff dff_A_VJxtsCrL3_0(.dout(w_dff_A_eEbU4kSa5_0),.din(w_dff_A_VJxtsCrL3_0),.clk(gclk));
	jdff dff_A_eEbU4kSa5_0(.dout(w_dff_A_RnW1Otv69_0),.din(w_dff_A_eEbU4kSa5_0),.clk(gclk));
	jdff dff_A_RnW1Otv69_0(.dout(G676),.din(w_dff_A_RnW1Otv69_0),.clk(gclk));
	jdff dff_A_vTDZFZYD2_2(.dout(w_dff_A_dzXYR51q2_0),.din(w_dff_A_vTDZFZYD2_2),.clk(gclk));
	jdff dff_A_dzXYR51q2_0(.dout(w_dff_A_ntbpoAp36_0),.din(w_dff_A_dzXYR51q2_0),.clk(gclk));
	jdff dff_A_ntbpoAp36_0(.dout(w_dff_A_niYem8mS4_0),.din(w_dff_A_ntbpoAp36_0),.clk(gclk));
	jdff dff_A_niYem8mS4_0(.dout(w_dff_A_V0cwFGeF1_0),.din(w_dff_A_niYem8mS4_0),.clk(gclk));
	jdff dff_A_V0cwFGeF1_0(.dout(w_dff_A_y6GK1rNB0_0),.din(w_dff_A_V0cwFGeF1_0),.clk(gclk));
	jdff dff_A_y6GK1rNB0_0(.dout(w_dff_A_omhyUGMP0_0),.din(w_dff_A_y6GK1rNB0_0),.clk(gclk));
	jdff dff_A_omhyUGMP0_0(.dout(w_dff_A_DnkTZt5R7_0),.din(w_dff_A_omhyUGMP0_0),.clk(gclk));
	jdff dff_A_DnkTZt5R7_0(.dout(w_dff_A_xzw6bPNm8_0),.din(w_dff_A_DnkTZt5R7_0),.clk(gclk));
	jdff dff_A_xzw6bPNm8_0(.dout(w_dff_A_MJBaLzfO8_0),.din(w_dff_A_xzw6bPNm8_0),.clk(gclk));
	jdff dff_A_MJBaLzfO8_0(.dout(G696),.din(w_dff_A_MJBaLzfO8_0),.clk(gclk));
	jdff dff_A_AjepxUwp4_2(.dout(w_dff_A_XCQr6ENL5_0),.din(w_dff_A_AjepxUwp4_2),.clk(gclk));
	jdff dff_A_XCQr6ENL5_0(.dout(w_dff_A_4iUBItTP6_0),.din(w_dff_A_XCQr6ENL5_0),.clk(gclk));
	jdff dff_A_4iUBItTP6_0(.dout(w_dff_A_5fy59RcD7_0),.din(w_dff_A_4iUBItTP6_0),.clk(gclk));
	jdff dff_A_5fy59RcD7_0(.dout(w_dff_A_KEY2srag6_0),.din(w_dff_A_5fy59RcD7_0),.clk(gclk));
	jdff dff_A_KEY2srag6_0(.dout(w_dff_A_mjtU9AHk4_0),.din(w_dff_A_KEY2srag6_0),.clk(gclk));
	jdff dff_A_mjtU9AHk4_0(.dout(w_dff_A_orjcsuiy3_0),.din(w_dff_A_mjtU9AHk4_0),.clk(gclk));
	jdff dff_A_orjcsuiy3_0(.dout(w_dff_A_pdsxLkeO1_0),.din(w_dff_A_orjcsuiy3_0),.clk(gclk));
	jdff dff_A_pdsxLkeO1_0(.dout(w_dff_A_Jy8wTgxs7_0),.din(w_dff_A_pdsxLkeO1_0),.clk(gclk));
	jdff dff_A_Jy8wTgxs7_0(.dout(w_dff_A_ljOFfVkY1_0),.din(w_dff_A_Jy8wTgxs7_0),.clk(gclk));
	jdff dff_A_ljOFfVkY1_0(.dout(G699),.din(w_dff_A_ljOFfVkY1_0),.clk(gclk));
	jdff dff_A_YYfSZWDj9_2(.dout(w_dff_A_lUhqxXJL7_0),.din(w_dff_A_YYfSZWDj9_2),.clk(gclk));
	jdff dff_A_lUhqxXJL7_0(.dout(w_dff_A_YMjM2Ud85_0),.din(w_dff_A_lUhqxXJL7_0),.clk(gclk));
	jdff dff_A_YMjM2Ud85_0(.dout(w_dff_A_0UB1Df464_0),.din(w_dff_A_YMjM2Ud85_0),.clk(gclk));
	jdff dff_A_0UB1Df464_0(.dout(w_dff_A_9jfZYRcd1_0),.din(w_dff_A_0UB1Df464_0),.clk(gclk));
	jdff dff_A_9jfZYRcd1_0(.dout(w_dff_A_PdQpDT420_0),.din(w_dff_A_9jfZYRcd1_0),.clk(gclk));
	jdff dff_A_PdQpDT420_0(.dout(w_dff_A_E0S89ySh4_0),.din(w_dff_A_PdQpDT420_0),.clk(gclk));
	jdff dff_A_E0S89ySh4_0(.dout(w_dff_A_BHXCaqFf0_0),.din(w_dff_A_E0S89ySh4_0),.clk(gclk));
	jdff dff_A_BHXCaqFf0_0(.dout(w_dff_A_noQDTBnq8_0),.din(w_dff_A_BHXCaqFf0_0),.clk(gclk));
	jdff dff_A_noQDTBnq8_0(.dout(G702),.din(w_dff_A_noQDTBnq8_0),.clk(gclk));
	jdff dff_A_NtujIeyr1_2(.dout(w_dff_A_3GEXZkbc4_0),.din(w_dff_A_NtujIeyr1_2),.clk(gclk));
	jdff dff_A_3GEXZkbc4_0(.dout(w_dff_A_5uzGkFqz9_0),.din(w_dff_A_3GEXZkbc4_0),.clk(gclk));
	jdff dff_A_5uzGkFqz9_0(.dout(w_dff_A_XYPAskFG3_0),.din(w_dff_A_5uzGkFqz9_0),.clk(gclk));
	jdff dff_A_XYPAskFG3_0(.dout(w_dff_A_fHltWVbY3_0),.din(w_dff_A_XYPAskFG3_0),.clk(gclk));
	jdff dff_A_fHltWVbY3_0(.dout(w_dff_A_JuACqhWv4_0),.din(w_dff_A_fHltWVbY3_0),.clk(gclk));
	jdff dff_A_JuACqhWv4_0(.dout(w_dff_A_aKGtkH7S1_0),.din(w_dff_A_JuACqhWv4_0),.clk(gclk));
	jdff dff_A_aKGtkH7S1_0(.dout(G818),.din(w_dff_A_aKGtkH7S1_0),.clk(gclk));
	jdff dff_A_bLgQBZ9M2_2(.dout(w_dff_A_Ry7IyVw57_0),.din(w_dff_A_bLgQBZ9M2_2),.clk(gclk));
	jdff dff_A_Ry7IyVw57_0(.dout(w_dff_A_zKt59K149_0),.din(w_dff_A_Ry7IyVw57_0),.clk(gclk));
	jdff dff_A_zKt59K149_0(.dout(w_dff_A_NSdd7evn8_0),.din(w_dff_A_zKt59K149_0),.clk(gclk));
	jdff dff_A_NSdd7evn8_0(.dout(w_dff_A_yCH3Lclx7_0),.din(w_dff_A_NSdd7evn8_0),.clk(gclk));
	jdff dff_A_yCH3Lclx7_0(.dout(w_dff_A_yW12xv8D7_0),.din(w_dff_A_yCH3Lclx7_0),.clk(gclk));
	jdff dff_A_yW12xv8D7_0(.dout(w_dff_A_ZmWFKoF42_0),.din(w_dff_A_yW12xv8D7_0),.clk(gclk));
	jdff dff_A_ZmWFKoF42_0(.dout(w_dff_A_6j1meksg1_0),.din(w_dff_A_ZmWFKoF42_0),.clk(gclk));
	jdff dff_A_6j1meksg1_0(.dout(w_dff_A_N7k9uy9l9_0),.din(w_dff_A_6j1meksg1_0),.clk(gclk));
	jdff dff_A_N7k9uy9l9_0(.dout(w_dff_A_HFyqO3fr6_0),.din(w_dff_A_N7k9uy9l9_0),.clk(gclk));
	jdff dff_A_HFyqO3fr6_0(.dout(G813),.din(w_dff_A_HFyqO3fr6_0),.clk(gclk));
	jdff dff_A_IwSzkPSy1_1(.dout(w_dff_A_xmLRzduV5_0),.din(w_dff_A_IwSzkPSy1_1),.clk(gclk));
	jdff dff_A_xmLRzduV5_0(.dout(w_dff_A_M57NM7Aw3_0),.din(w_dff_A_xmLRzduV5_0),.clk(gclk));
	jdff dff_A_M57NM7Aw3_0(.dout(w_dff_A_SPCSwg5j3_0),.din(w_dff_A_M57NM7Aw3_0),.clk(gclk));
	jdff dff_A_SPCSwg5j3_0(.dout(w_dff_A_vGuKqxff8_0),.din(w_dff_A_SPCSwg5j3_0),.clk(gclk));
	jdff dff_A_vGuKqxff8_0(.dout(w_dff_A_11Clv3lA0_0),.din(w_dff_A_vGuKqxff8_0),.clk(gclk));
	jdff dff_A_11Clv3lA0_0(.dout(w_dff_A_7dPYPCaj9_0),.din(w_dff_A_11Clv3lA0_0),.clk(gclk));
	jdff dff_A_7dPYPCaj9_0(.dout(G824),.din(w_dff_A_7dPYPCaj9_0),.clk(gclk));
	jdff dff_A_LBerTre86_1(.dout(w_dff_A_7glTpZaY8_0),.din(w_dff_A_LBerTre86_1),.clk(gclk));
	jdff dff_A_7glTpZaY8_0(.dout(w_dff_A_sOEkLcEg6_0),.din(w_dff_A_7glTpZaY8_0),.clk(gclk));
	jdff dff_A_sOEkLcEg6_0(.dout(w_dff_A_Dklo9zPs0_0),.din(w_dff_A_sOEkLcEg6_0),.clk(gclk));
	jdff dff_A_Dklo9zPs0_0(.dout(w_dff_A_3YWx98ka9_0),.din(w_dff_A_Dklo9zPs0_0),.clk(gclk));
	jdff dff_A_3YWx98ka9_0(.dout(w_dff_A_3jdzWI766_0),.din(w_dff_A_3YWx98ka9_0),.clk(gclk));
	jdff dff_A_3jdzWI766_0(.dout(w_dff_A_fKuXXjJx4_0),.din(w_dff_A_3jdzWI766_0),.clk(gclk));
	jdff dff_A_fKuXXjJx4_0(.dout(w_dff_A_rmyDQuBi2_0),.din(w_dff_A_fKuXXjJx4_0),.clk(gclk));
	jdff dff_A_rmyDQuBi2_0(.dout(G826),.din(w_dff_A_rmyDQuBi2_0),.clk(gclk));
	jdff dff_A_2FsCfOkF2_1(.dout(w_dff_A_KlbY66Mt6_0),.din(w_dff_A_2FsCfOkF2_1),.clk(gclk));
	jdff dff_A_KlbY66Mt6_0(.dout(w_dff_A_ocCd8uyj8_0),.din(w_dff_A_KlbY66Mt6_0),.clk(gclk));
	jdff dff_A_ocCd8uyj8_0(.dout(w_dff_A_fls6G7XE8_0),.din(w_dff_A_ocCd8uyj8_0),.clk(gclk));
	jdff dff_A_fls6G7XE8_0(.dout(w_dff_A_OkihA47d8_0),.din(w_dff_A_fls6G7XE8_0),.clk(gclk));
	jdff dff_A_OkihA47d8_0(.dout(w_dff_A_1fDItDbd7_0),.din(w_dff_A_OkihA47d8_0),.clk(gclk));
	jdff dff_A_1fDItDbd7_0(.dout(w_dff_A_i6pwenAP1_0),.din(w_dff_A_1fDItDbd7_0),.clk(gclk));
	jdff dff_A_i6pwenAP1_0(.dout(G828),.din(w_dff_A_i6pwenAP1_0),.clk(gclk));
	jdff dff_A_rvkGvTDO1_1(.dout(w_dff_A_6Cpsv1q82_0),.din(w_dff_A_rvkGvTDO1_1),.clk(gclk));
	jdff dff_A_6Cpsv1q82_0(.dout(w_dff_A_MErzE5j98_0),.din(w_dff_A_6Cpsv1q82_0),.clk(gclk));
	jdff dff_A_MErzE5j98_0(.dout(w_dff_A_Wqgza2RQ9_0),.din(w_dff_A_MErzE5j98_0),.clk(gclk));
	jdff dff_A_Wqgza2RQ9_0(.dout(w_dff_A_hWOZ5pYt5_0),.din(w_dff_A_Wqgza2RQ9_0),.clk(gclk));
	jdff dff_A_hWOZ5pYt5_0(.dout(w_dff_A_p9EJNKVZ2_0),.din(w_dff_A_hWOZ5pYt5_0),.clk(gclk));
	jdff dff_A_p9EJNKVZ2_0(.dout(w_dff_A_nhz6DzGj1_0),.din(w_dff_A_p9EJNKVZ2_0),.clk(gclk));
	jdff dff_A_nhz6DzGj1_0(.dout(w_dff_A_hTYwL6zP1_0),.din(w_dff_A_nhz6DzGj1_0),.clk(gclk));
	jdff dff_A_hTYwL6zP1_0(.dout(w_dff_A_06RPFrg26_0),.din(w_dff_A_hTYwL6zP1_0),.clk(gclk));
	jdff dff_A_06RPFrg26_0(.dout(w_dff_A_e0hzDGeR8_0),.din(w_dff_A_06RPFrg26_0),.clk(gclk));
	jdff dff_A_e0hzDGeR8_0(.dout(w_dff_A_hdaSVyk01_0),.din(w_dff_A_e0hzDGeR8_0),.clk(gclk));
	jdff dff_A_hdaSVyk01_0(.dout(w_dff_A_C1ao7ope7_0),.din(w_dff_A_hdaSVyk01_0),.clk(gclk));
	jdff dff_A_C1ao7ope7_0(.dout(G830),.din(w_dff_A_C1ao7ope7_0),.clk(gclk));
	jdff dff_A_GCA5ODBX8_2(.dout(w_dff_A_E1qSkLM86_0),.din(w_dff_A_GCA5ODBX8_2),.clk(gclk));
	jdff dff_A_E1qSkLM86_0(.dout(w_dff_A_1QYWHjkS6_0),.din(w_dff_A_E1qSkLM86_0),.clk(gclk));
	jdff dff_A_1QYWHjkS6_0(.dout(w_dff_A_Il36ld8O1_0),.din(w_dff_A_1QYWHjkS6_0),.clk(gclk));
	jdff dff_A_Il36ld8O1_0(.dout(w_dff_A_vW0gvt8x0_0),.din(w_dff_A_Il36ld8O1_0),.clk(gclk));
	jdff dff_A_vW0gvt8x0_0(.dout(w_dff_A_rBtOGuzq8_0),.din(w_dff_A_vW0gvt8x0_0),.clk(gclk));
	jdff dff_A_rBtOGuzq8_0(.dout(w_dff_A_nswSbyau4_0),.din(w_dff_A_rBtOGuzq8_0),.clk(gclk));
	jdff dff_A_nswSbyau4_0(.dout(w_dff_A_4R1SgZ0V5_0),.din(w_dff_A_nswSbyau4_0),.clk(gclk));
	jdff dff_A_4R1SgZ0V5_0(.dout(w_dff_A_Bk3R6bQQ2_0),.din(w_dff_A_4R1SgZ0V5_0),.clk(gclk));
	jdff dff_A_Bk3R6bQQ2_0(.dout(w_dff_A_NVyKeG0k4_0),.din(w_dff_A_Bk3R6bQQ2_0),.clk(gclk));
	jdff dff_A_NVyKeG0k4_0(.dout(w_dff_A_4dm6cnJD6_0),.din(w_dff_A_NVyKeG0k4_0),.clk(gclk));
	jdff dff_A_4dm6cnJD6_0(.dout(w_dff_A_krqCzVYp3_0),.din(w_dff_A_4dm6cnJD6_0),.clk(gclk));
	jdff dff_A_krqCzVYp3_0(.dout(w_dff_A_iGMB3ghD4_0),.din(w_dff_A_krqCzVYp3_0),.clk(gclk));
	jdff dff_A_iGMB3ghD4_0(.dout(w_dff_A_RmCZmxKB9_0),.din(w_dff_A_iGMB3ghD4_0),.clk(gclk));
	jdff dff_A_RmCZmxKB9_0(.dout(w_dff_A_6q9Z6IT89_0),.din(w_dff_A_RmCZmxKB9_0),.clk(gclk));
	jdff dff_A_6q9Z6IT89_0(.dout(w_dff_A_OqgYmzyH3_0),.din(w_dff_A_6q9Z6IT89_0),.clk(gclk));
	jdff dff_A_OqgYmzyH3_0(.dout(w_dff_A_6H9zuHzz1_0),.din(w_dff_A_OqgYmzyH3_0),.clk(gclk));
	jdff dff_A_6H9zuHzz1_0(.dout(G854),.din(w_dff_A_6H9zuHzz1_0),.clk(gclk));
	jdff dff_A_17s6VL7c5_1(.dout(w_dff_A_xJX52c8s6_0),.din(w_dff_A_17s6VL7c5_1),.clk(gclk));
	jdff dff_A_xJX52c8s6_0(.dout(w_dff_A_c4goXiz96_0),.din(w_dff_A_xJX52c8s6_0),.clk(gclk));
	jdff dff_A_c4goXiz96_0(.dout(w_dff_A_rgA4Rmsz0_0),.din(w_dff_A_c4goXiz96_0),.clk(gclk));
	jdff dff_A_rgA4Rmsz0_0(.dout(w_dff_A_2HcFLX1g2_0),.din(w_dff_A_rgA4Rmsz0_0),.clk(gclk));
	jdff dff_A_2HcFLX1g2_0(.dout(w_dff_A_ogovuXZC5_0),.din(w_dff_A_2HcFLX1g2_0),.clk(gclk));
	jdff dff_A_ogovuXZC5_0(.dout(G863),.din(w_dff_A_ogovuXZC5_0),.clk(gclk));
	jdff dff_A_6AWDkRJl7_1(.dout(w_dff_A_CMvyFcM13_0),.din(w_dff_A_6AWDkRJl7_1),.clk(gclk));
	jdff dff_A_CMvyFcM13_0(.dout(w_dff_A_KzUiaDeT1_0),.din(w_dff_A_CMvyFcM13_0),.clk(gclk));
	jdff dff_A_KzUiaDeT1_0(.dout(w_dff_A_DzyFzZU60_0),.din(w_dff_A_KzUiaDeT1_0),.clk(gclk));
	jdff dff_A_DzyFzZU60_0(.dout(w_dff_A_fOCbuJSH7_0),.din(w_dff_A_DzyFzZU60_0),.clk(gclk));
	jdff dff_A_fOCbuJSH7_0(.dout(w_dff_A_xbFWoSHn1_0),.din(w_dff_A_fOCbuJSH7_0),.clk(gclk));
	jdff dff_A_xbFWoSHn1_0(.dout(w_dff_A_WDtBrpU84_0),.din(w_dff_A_xbFWoSHn1_0),.clk(gclk));
	jdff dff_A_WDtBrpU84_0(.dout(w_dff_A_rndAmwxd1_0),.din(w_dff_A_WDtBrpU84_0),.clk(gclk));
	jdff dff_A_rndAmwxd1_0(.dout(w_dff_A_3FCjCRUX7_0),.din(w_dff_A_rndAmwxd1_0),.clk(gclk));
	jdff dff_A_3FCjCRUX7_0(.dout(G865),.din(w_dff_A_3FCjCRUX7_0),.clk(gclk));
	jdff dff_A_RDGMn0975_1(.dout(w_dff_A_BO6oQZSM1_0),.din(w_dff_A_RDGMn0975_1),.clk(gclk));
	jdff dff_A_BO6oQZSM1_0(.dout(w_dff_A_7mTk3Ov96_0),.din(w_dff_A_BO6oQZSM1_0),.clk(gclk));
	jdff dff_A_7mTk3Ov96_0(.dout(w_dff_A_79c8EDKn7_0),.din(w_dff_A_7mTk3Ov96_0),.clk(gclk));
	jdff dff_A_79c8EDKn7_0(.dout(w_dff_A_WASfQaS48_0),.din(w_dff_A_79c8EDKn7_0),.clk(gclk));
	jdff dff_A_WASfQaS48_0(.dout(w_dff_A_q32xcWwK2_0),.din(w_dff_A_WASfQaS48_0),.clk(gclk));
	jdff dff_A_q32xcWwK2_0(.dout(w_dff_A_kfyGwrzl8_0),.din(w_dff_A_q32xcWwK2_0),.clk(gclk));
	jdff dff_A_kfyGwrzl8_0(.dout(G867),.din(w_dff_A_kfyGwrzl8_0),.clk(gclk));
	jdff dff_A_XkPdcrtq8_1(.dout(w_dff_A_gzDeM6uj5_0),.din(w_dff_A_XkPdcrtq8_1),.clk(gclk));
	jdff dff_A_gzDeM6uj5_0(.dout(w_dff_A_20ru1FE20_0),.din(w_dff_A_gzDeM6uj5_0),.clk(gclk));
	jdff dff_A_20ru1FE20_0(.dout(w_dff_A_L0fqvtNV9_0),.din(w_dff_A_20ru1FE20_0),.clk(gclk));
	jdff dff_A_L0fqvtNV9_0(.dout(w_dff_A_D6KCyxOu2_0),.din(w_dff_A_L0fqvtNV9_0),.clk(gclk));
	jdff dff_A_D6KCyxOu2_0(.dout(w_dff_A_1nW2iSBe6_0),.din(w_dff_A_D6KCyxOu2_0),.clk(gclk));
	jdff dff_A_1nW2iSBe6_0(.dout(w_dff_A_gNwfsd558_0),.din(w_dff_A_1nW2iSBe6_0),.clk(gclk));
	jdff dff_A_gNwfsd558_0(.dout(w_dff_A_iQi5mYeG0_0),.din(w_dff_A_gNwfsd558_0),.clk(gclk));
	jdff dff_A_iQi5mYeG0_0(.dout(w_dff_A_EnVzPwhT1_0),.din(w_dff_A_iQi5mYeG0_0),.clk(gclk));
	jdff dff_A_EnVzPwhT1_0(.dout(w_dff_A_dunK0EDY6_0),.din(w_dff_A_EnVzPwhT1_0),.clk(gclk));
	jdff dff_A_dunK0EDY6_0(.dout(G869),.din(w_dff_A_dunK0EDY6_0),.clk(gclk));
	jdff dff_A_e2RZ5Gl43_2(.dout(w_dff_A_bG2uJ3eV1_0),.din(w_dff_A_e2RZ5Gl43_2),.clk(gclk));
	jdff dff_A_bG2uJ3eV1_0(.dout(w_dff_A_xVvOH0tH8_0),.din(w_dff_A_bG2uJ3eV1_0),.clk(gclk));
	jdff dff_A_xVvOH0tH8_0(.dout(w_dff_A_lS0zHRg66_0),.din(w_dff_A_xVvOH0tH8_0),.clk(gclk));
	jdff dff_A_lS0zHRg66_0(.dout(G712),.din(w_dff_A_lS0zHRg66_0),.clk(gclk));
	jdff dff_A_FqM4NOCB0_2(.dout(w_dff_A_4DvjwDJx3_0),.din(w_dff_A_FqM4NOCB0_2),.clk(gclk));
	jdff dff_A_4DvjwDJx3_0(.dout(w_dff_A_DeZOut8m1_0),.din(w_dff_A_4DvjwDJx3_0),.clk(gclk));
	jdff dff_A_DeZOut8m1_0(.dout(G727),.din(w_dff_A_DeZOut8m1_0),.clk(gclk));
	jdff dff_A_lz8TOsR45_2(.dout(w_dff_A_T7GgUKXY0_0),.din(w_dff_A_lz8TOsR45_2),.clk(gclk));
	jdff dff_A_T7GgUKXY0_0(.dout(w_dff_A_PmtGzS3m3_0),.din(w_dff_A_T7GgUKXY0_0),.clk(gclk));
	jdff dff_A_PmtGzS3m3_0(.dout(w_dff_A_sgYWj5mX7_0),.din(w_dff_A_PmtGzS3m3_0),.clk(gclk));
	jdff dff_A_sgYWj5mX7_0(.dout(G732),.din(w_dff_A_sgYWj5mX7_0),.clk(gclk));
	jdff dff_A_WIFa6DUd8_2(.dout(w_dff_A_IGZem14g4_0),.din(w_dff_A_WIFa6DUd8_2),.clk(gclk));
	jdff dff_A_IGZem14g4_0(.dout(w_dff_A_0hmhzQZq2_0),.din(w_dff_A_IGZem14g4_0),.clk(gclk));
	jdff dff_A_0hmhzQZq2_0(.dout(w_dff_A_lqFU7hcd2_0),.din(w_dff_A_0hmhzQZq2_0),.clk(gclk));
	jdff dff_A_lqFU7hcd2_0(.dout(G737),.din(w_dff_A_lqFU7hcd2_0),.clk(gclk));
	jdff dff_A_qzcfvnFP9_2(.dout(w_dff_A_EaHqP5YT5_0),.din(w_dff_A_qzcfvnFP9_2),.clk(gclk));
	jdff dff_A_EaHqP5YT5_0(.dout(w_dff_A_GL5Omq3X5_0),.din(w_dff_A_EaHqP5YT5_0),.clk(gclk));
	jdff dff_A_GL5Omq3X5_0(.dout(w_dff_A_OEgS7cZX5_0),.din(w_dff_A_GL5Omq3X5_0),.clk(gclk));
	jdff dff_A_OEgS7cZX5_0(.dout(w_dff_A_YP9pzYy54_0),.din(w_dff_A_OEgS7cZX5_0),.clk(gclk));
	jdff dff_A_YP9pzYy54_0(.dout(G742),.din(w_dff_A_YP9pzYy54_0),.clk(gclk));
	jdff dff_A_OWe3VifZ2_2(.dout(w_dff_A_aUeO30zP0_0),.din(w_dff_A_OWe3VifZ2_2),.clk(gclk));
	jdff dff_A_aUeO30zP0_0(.dout(w_dff_A_XIo6DZ1C0_0),.din(w_dff_A_aUeO30zP0_0),.clk(gclk));
	jdff dff_A_XIo6DZ1C0_0(.dout(w_dff_A_FRUnh6fN7_0),.din(w_dff_A_XIo6DZ1C0_0),.clk(gclk));
	jdff dff_A_FRUnh6fN7_0(.dout(G772),.din(w_dff_A_FRUnh6fN7_0),.clk(gclk));
	jdff dff_A_SnzgluzA6_2(.dout(w_dff_A_HV3vwFJI0_0),.din(w_dff_A_SnzgluzA6_2),.clk(gclk));
	jdff dff_A_HV3vwFJI0_0(.dout(w_dff_A_2k0MkZu08_0),.din(w_dff_A_HV3vwFJI0_0),.clk(gclk));
	jdff dff_A_2k0MkZu08_0(.dout(w_dff_A_tiNEzIGs1_0),.din(w_dff_A_2k0MkZu08_0),.clk(gclk));
	jdff dff_A_tiNEzIGs1_0(.dout(G777),.din(w_dff_A_tiNEzIGs1_0),.clk(gclk));
	jdff dff_A_xWOXwuxG9_2(.dout(w_dff_A_RMXMFMqp9_0),.din(w_dff_A_xWOXwuxG9_2),.clk(gclk));
	jdff dff_A_RMXMFMqp9_0(.dout(w_dff_A_eHIQODzU2_0),.din(w_dff_A_RMXMFMqp9_0),.clk(gclk));
	jdff dff_A_eHIQODzU2_0(.dout(w_dff_A_qKI4RqgR6_0),.din(w_dff_A_eHIQODzU2_0),.clk(gclk));
	jdff dff_A_qKI4RqgR6_0(.dout(w_dff_A_W9aXYAXe0_0),.din(w_dff_A_qKI4RqgR6_0),.clk(gclk));
	jdff dff_A_W9aXYAXe0_0(.dout(G782),.din(w_dff_A_W9aXYAXe0_0),.clk(gclk));
	jdff dff_A_XEra2e6U0_2(.dout(w_dff_A_zqQ1hpHe8_0),.din(w_dff_A_XEra2e6U0_2),.clk(gclk));
	jdff dff_A_zqQ1hpHe8_0(.dout(w_dff_A_gZvxIxvA7_0),.din(w_dff_A_zqQ1hpHe8_0),.clk(gclk));
	jdff dff_A_gZvxIxvA7_0(.dout(w_dff_A_1gmJbbnx5_0),.din(w_dff_A_gZvxIxvA7_0),.clk(gclk));
	jdff dff_A_1gmJbbnx5_0(.dout(G645),.din(w_dff_A_1gmJbbnx5_0),.clk(gclk));
	jdff dff_A_nhdDMIc41_2(.dout(w_dff_A_c9kVy9Yk9_0),.din(w_dff_A_nhdDMIc41_2),.clk(gclk));
	jdff dff_A_c9kVy9Yk9_0(.dout(w_dff_A_iEsytF7y2_0),.din(w_dff_A_c9kVy9Yk9_0),.clk(gclk));
	jdff dff_A_iEsytF7y2_0(.dout(G648),.din(w_dff_A_iEsytF7y2_0),.clk(gclk));
	jdff dff_A_8corv2mp0_2(.dout(w_dff_A_IQ7GLwJM3_0),.din(w_dff_A_8corv2mp0_2),.clk(gclk));
	jdff dff_A_IQ7GLwJM3_0(.dout(w_dff_A_T1bIQLwm5_0),.din(w_dff_A_IQ7GLwJM3_0),.clk(gclk));
	jdff dff_A_T1bIQLwm5_0(.dout(G651),.din(w_dff_A_T1bIQLwm5_0),.clk(gclk));
	jdff dff_A_8CLLA1Vs8_2(.dout(w_dff_A_M2kpsJKY0_0),.din(w_dff_A_8CLLA1Vs8_2),.clk(gclk));
	jdff dff_A_M2kpsJKY0_0(.dout(G654),.din(w_dff_A_M2kpsJKY0_0),.clk(gclk));
	jdff dff_A_DYPsKfAw4_2(.dout(w_dff_A_EIWhP4VZ5_0),.din(w_dff_A_DYPsKfAw4_2),.clk(gclk));
	jdff dff_A_EIWhP4VZ5_0(.dout(w_dff_A_KEz0mcUa8_0),.din(w_dff_A_EIWhP4VZ5_0),.clk(gclk));
	jdff dff_A_KEz0mcUa8_0(.dout(w_dff_A_TC8wh8Mq3_0),.din(w_dff_A_KEz0mcUa8_0),.clk(gclk));
	jdff dff_A_TC8wh8Mq3_0(.dout(G679),.din(w_dff_A_TC8wh8Mq3_0),.clk(gclk));
	jdff dff_A_atPMyXnW8_2(.dout(w_dff_A_1TS8HJWG3_0),.din(w_dff_A_atPMyXnW8_2),.clk(gclk));
	jdff dff_A_1TS8HJWG3_0(.dout(w_dff_A_BoJpPChj2_0),.din(w_dff_A_1TS8HJWG3_0),.clk(gclk));
	jdff dff_A_BoJpPChj2_0(.dout(G682),.din(w_dff_A_BoJpPChj2_0),.clk(gclk));
	jdff dff_A_7Un7AyR00_2(.dout(w_dff_A_e2zYwXgF4_0),.din(w_dff_A_7Un7AyR00_2),.clk(gclk));
	jdff dff_A_e2zYwXgF4_0(.dout(w_dff_A_A9ssMPdF2_0),.din(w_dff_A_e2zYwXgF4_0),.clk(gclk));
	jdff dff_A_A9ssMPdF2_0(.dout(G685),.din(w_dff_A_A9ssMPdF2_0),.clk(gclk));
	jdff dff_A_JgJF4PTq7_2(.dout(w_dff_A_uQqnHAwU1_0),.din(w_dff_A_JgJF4PTq7_2),.clk(gclk));
	jdff dff_A_uQqnHAwU1_0(.dout(w_dff_A_PlcUNtY39_0),.din(w_dff_A_uQqnHAwU1_0),.clk(gclk));
	jdff dff_A_PlcUNtY39_0(.dout(G688),.din(w_dff_A_PlcUNtY39_0),.clk(gclk));
	jdff dff_A_UlPKT5TM8_2(.dout(w_dff_A_PM5GHO3P3_0),.din(w_dff_A_UlPKT5TM8_2),.clk(gclk));
	jdff dff_A_PM5GHO3P3_0(.dout(w_dff_A_qwxGPqp95_0),.din(w_dff_A_PM5GHO3P3_0),.clk(gclk));
	jdff dff_A_qwxGPqp95_0(.dout(w_dff_A_aueYEHx92_0),.din(w_dff_A_qwxGPqp95_0),.clk(gclk));
	jdff dff_A_aueYEHx92_0(.dout(w_dff_A_vETPxkNk9_0),.din(w_dff_A_aueYEHx92_0),.clk(gclk));
	jdff dff_A_vETPxkNk9_0(.dout(w_dff_A_JBFDhhb70_0),.din(w_dff_A_vETPxkNk9_0),.clk(gclk));
	jdff dff_A_JBFDhhb70_0(.dout(G843),.din(w_dff_A_JBFDhhb70_0),.clk(gclk));
	jdff dff_A_7huooCbl2_2(.dout(w_dff_A_A6z6T7NX4_0),.din(w_dff_A_7huooCbl2_2),.clk(gclk));
	jdff dff_A_A6z6T7NX4_0(.dout(w_dff_A_kKt2Q9X98_0),.din(w_dff_A_A6z6T7NX4_0),.clk(gclk));
	jdff dff_A_kKt2Q9X98_0(.dout(w_dff_A_qQ9eMm2M7_0),.din(w_dff_A_kKt2Q9X98_0),.clk(gclk));
	jdff dff_A_qQ9eMm2M7_0(.dout(w_dff_A_v3AVm0XO2_0),.din(w_dff_A_qQ9eMm2M7_0),.clk(gclk));
	jdff dff_A_v3AVm0XO2_0(.dout(w_dff_A_yp9N7ak12_0),.din(w_dff_A_v3AVm0XO2_0),.clk(gclk));
	jdff dff_A_yp9N7ak12_0(.dout(G882),.din(w_dff_A_yp9N7ak12_0),.clk(gclk));
	jdff dff_A_8I5o8ymm2_2(.dout(G767),.din(w_dff_A_8I5o8ymm2_2),.clk(gclk));
	jdff dff_A_fkiBKvyy9_2(.dout(G807),.din(w_dff_A_fkiBKvyy9_2),.clk(gclk));
endmodule

