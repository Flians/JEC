/*
gf_c3540:
	jxor: 52
	jspl: 225
	jspl3: 338
	jnot: 188
	jdff: 2183
	jand: 525
	jor: 352

Summary:
	jxor: 52
	jspl: 225
	jspl3: 338
	jnot: 188
	jdff: 2183
	jand: 525
	jor: 352

The maximum logic level gap of any gate:
	gf_c3540: 26
*/

module gf_c3540(gclk, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402);
	input gclk;
	input G1;
	input G13;
	input G20;
	input G33;
	input G41;
	input G45;
	input G50;
	input G58;
	input G68;
	input G77;
	input G87;
	input G97;
	input G107;
	input G116;
	input G124;
	input G125;
	input G128;
	input G132;
	input G137;
	input G143;
	input G150;
	input G159;
	input G169;
	input G179;
	input G190;
	input G200;
	input G213;
	input G222;
	input G223;
	input G226;
	input G232;
	input G238;
	input G244;
	input G250;
	input G257;
	input G264;
	input G270;
	input G274;
	input G283;
	input G294;
	input G303;
	input G311;
	input G317;
	input G322;
	input G326;
	input G329;
	input G330;
	input G343;
	input G1698;
	input G2897;
	output G353;
	output G355;
	output G361;
	output G358;
	output G351;
	output G372;
	output G369;
	output G399;
	output G364;
	output G396;
	output G384;
	output G367;
	output G387;
	output G393;
	output G390;
	output G378;
	output G375;
	output G381;
	output G407;
	output G409;
	output G405;
	output G402;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [1:0] w_G1_2;
	wire [2:0] w_G13_0;
	wire [2:0] w_G13_1;
	wire [1:0] w_G13_2;
	wire [2:0] w_G20_0;
	wire [2:0] w_G20_1;
	wire [2:0] w_G20_2;
	wire [2:0] w_G20_3;
	wire [2:0] w_G20_4;
	wire [2:0] w_G20_5;
	wire [2:0] w_G20_6;
	wire [2:0] w_G33_0;
	wire [2:0] w_G33_1;
	wire [2:0] w_G33_2;
	wire [2:0] w_G33_3;
	wire [2:0] w_G33_4;
	wire [2:0] w_G33_5;
	wire [2:0] w_G33_6;
	wire [2:0] w_G33_7;
	wire [2:0] w_G33_8;
	wire [2:0] w_G33_9;
	wire [2:0] w_G33_10;
	wire [2:0] w_G33_11;
	wire [2:0] w_G33_12;
	wire [2:0] w_G41_0;
	wire [2:0] w_G45_0;
	wire [1:0] w_G45_1;
	wire [2:0] w_G50_0;
	wire [2:0] w_G50_1;
	wire [2:0] w_G50_2;
	wire [2:0] w_G50_3;
	wire [2:0] w_G50_4;
	wire [2:0] w_G50_5;
	wire [2:0] w_G58_0;
	wire [2:0] w_G58_1;
	wire [2:0] w_G58_2;
	wire [2:0] w_G58_3;
	wire [2:0] w_G58_4;
	wire [2:0] w_G58_5;
	wire [2:0] w_G68_0;
	wire [2:0] w_G68_1;
	wire [2:0] w_G68_2;
	wire [2:0] w_G68_3;
	wire [2:0] w_G68_4;
	wire [2:0] w_G68_5;
	wire [2:0] w_G77_0;
	wire [2:0] w_G77_1;
	wire [2:0] w_G77_2;
	wire [2:0] w_G77_3;
	wire [2:0] w_G77_4;
	wire [2:0] w_G87_0;
	wire [2:0] w_G87_1;
	wire [2:0] w_G87_2;
	wire [2:0] w_G87_3;
	wire [2:0] w_G97_0;
	wire [2:0] w_G97_1;
	wire [2:0] w_G97_2;
	wire [2:0] w_G97_3;
	wire [2:0] w_G97_4;
	wire [2:0] w_G107_0;
	wire [2:0] w_G107_1;
	wire [2:0] w_G107_2;
	wire [2:0] w_G107_3;
	wire [1:0] w_G107_4;
	wire [2:0] w_G116_0;
	wire [2:0] w_G116_1;
	wire [2:0] w_G116_2;
	wire [2:0] w_G116_3;
	wire [2:0] w_G116_4;
	wire [2:0] w_G116_5;
	wire [1:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [2:0] w_G132_0;
	wire [1:0] w_G132_1;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G143_0;
	wire [2:0] w_G143_1;
	wire [1:0] w_G143_2;
	wire [2:0] w_G150_0;
	wire [2:0] w_G150_1;
	wire [2:0] w_G150_2;
	wire [1:0] w_G150_3;
	wire [2:0] w_G159_0;
	wire [2:0] w_G159_1;
	wire [2:0] w_G159_2;
	wire [2:0] w_G159_3;
	wire [2:0] w_G169_0;
	wire [2:0] w_G169_1;
	wire [2:0] w_G169_2;
	wire [1:0] w_G169_3;
	wire [2:0] w_G179_0;
	wire [2:0] w_G179_1;
	wire [2:0] w_G179_2;
	wire [2:0] w_G190_0;
	wire [2:0] w_G190_1;
	wire [2:0] w_G190_2;
	wire [2:0] w_G190_3;
	wire [2:0] w_G190_4;
	wire [2:0] w_G200_0;
	wire [2:0] w_G200_1;
	wire [2:0] w_G200_2;
	wire [1:0] w_G200_3;
	wire [2:0] w_G213_0;
	wire [1:0] w_G223_0;
	wire [2:0] w_G226_0;
	wire [2:0] w_G226_1;
	wire [2:0] w_G232_0;
	wire [2:0] w_G232_1;
	wire [2:0] w_G238_0;
	wire [2:0] w_G244_0;
	wire [1:0] w_G244_1;
	wire [2:0] w_G250_0;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [2:0] w_G264_0;
	wire [2:0] w_G270_0;
	wire [2:0] w_G274_0;
	wire [2:0] w_G283_0;
	wire [2:0] w_G283_1;
	wire [2:0] w_G283_2;
	wire [2:0] w_G283_3;
	wire [2:0] w_G294_0;
	wire [2:0] w_G294_1;
	wire [2:0] w_G294_2;
	wire [1:0] w_G294_3;
	wire [2:0] w_G303_0;
	wire [2:0] w_G303_1;
	wire [2:0] w_G303_2;
	wire [2:0] w_G311_0;
	wire [2:0] w_G311_1;
	wire [2:0] w_G317_0;
	wire [1:0] w_G317_1;
	wire [2:0] w_G322_0;
	wire [1:0] w_G326_0;
	wire [2:0] w_G330_0;
	wire [1:0] w_G343_0;
	wire [2:0] w_G1698_0;
	wire w_G355_0;
	wire G355_fa_;
	wire w_G396_0;
	wire G396_fa_;
	wire w_G384_0;
	wire G384_fa_;
	wire [2:0] w_n72_0;
	wire [2:0] w_n72_1;
	wire [2:0] w_n73_0;
	wire [2:0] w_n73_1;
	wire [2:0] w_n73_2;
	wire [2:0] w_n74_0;
	wire [2:0] w_n74_1;
	wire [1:0] w_n74_2;
	wire [2:0] w_n75_0;
	wire [2:0] w_n75_1;
	wire [1:0] w_n75_2;
	wire [1:0] w_n76_0;
	wire [1:0] w_n77_0;
	wire [2:0] w_n79_0;
	wire [2:0] w_n79_1;
	wire [2:0] w_n80_0;
	wire [2:0] w_n80_1;
	wire [2:0] w_n81_0;
	wire [2:0] w_n81_1;
	wire [1:0] w_n81_2;
	wire [2:0] w_n84_0;
	wire [2:0] w_n84_1;
	wire [1:0] w_n85_0;
	wire [2:0] w_n86_0;
	wire [1:0] w_n89_0;
	wire [2:0] w_n90_0;
	wire [2:0] w_n91_0;
	wire [2:0] w_n91_1;
	wire [2:0] w_n94_0;
	wire [2:0] w_n96_0;
	wire [2:0] w_n105_0;
	wire [1:0] w_n105_1;
	wire [2:0] w_n111_0;
	wire [1:0] w_n112_0;
	wire [2:0] w_n118_0;
	wire [1:0] w_n120_0;
	wire [1:0] w_n126_0;
	wire [1:0] w_n130_0;
	wire [1:0] w_n134_0;
	wire [1:0] w_n137_0;
	wire [2:0] w_n139_0;
	wire [2:0] w_n139_1;
	wire [1:0] w_n140_0;
	wire [2:0] w_n141_0;
	wire [2:0] w_n141_1;
	wire [2:0] w_n141_2;
	wire [1:0] w_n141_3;
	wire [2:0] w_n142_0;
	wire [2:0] w_n142_1;
	wire [1:0] w_n142_2;
	wire [1:0] w_n143_0;
	wire [2:0] w_n144_0;
	wire [2:0] w_n144_1;
	wire [1:0] w_n144_2;
	wire [2:0] w_n147_0;
	wire [1:0] w_n148_0;
	wire [2:0] w_n151_0;
	wire [2:0] w_n151_1;
	wire [2:0] w_n151_2;
	wire [2:0] w_n151_3;
	wire [2:0] w_n151_4;
	wire [2:0] w_n151_5;
	wire [1:0] w_n151_6;
	wire [2:0] w_n152_0;
	wire [2:0] w_n153_0;
	wire [2:0] w_n153_1;
	wire [2:0] w_n153_2;
	wire [2:0] w_n153_3;
	wire [2:0] w_n153_4;
	wire [2:0] w_n153_5;
	wire [2:0] w_n153_6;
	wire [2:0] w_n153_7;
	wire [1:0] w_n153_8;
	wire [2:0] w_n161_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n163_1;
	wire [2:0] w_n164_0;
	wire [1:0] w_n165_0;
	wire [1:0] w_n167_0;
	wire [2:0] w_n168_0;
	wire [2:0] w_n168_1;
	wire [2:0] w_n168_2;
	wire [2:0] w_n168_3;
	wire [2:0] w_n168_4;
	wire [1:0] w_n168_5;
	wire [1:0] w_n169_0;
	wire [2:0] w_n170_0;
	wire [2:0] w_n172_0;
	wire [2:0] w_n172_1;
	wire [2:0] w_n172_2;
	wire [2:0] w_n172_3;
	wire [2:0] w_n172_4;
	wire [2:0] w_n173_0;
	wire [2:0] w_n173_1;
	wire [2:0] w_n173_2;
	wire [1:0] w_n173_3;
	wire [1:0] w_n176_0;
	wire [2:0] w_n177_0;
	wire [2:0] w_n177_1;
	wire [2:0] w_n182_0;
	wire [1:0] w_n182_1;
	wire [2:0] w_n186_0;
	wire [2:0] w_n186_1;
	wire [2:0] w_n189_0;
	wire [2:0] w_n189_1;
	wire [2:0] w_n189_2;
	wire [1:0] w_n190_0;
	wire [2:0] w_n192_0;
	wire [2:0] w_n198_0;
	wire [2:0] w_n199_0;
	wire [1:0] w_n201_0;
	wire [1:0] w_n202_0;
	wire [2:0] w_n205_0;
	wire [1:0] w_n205_1;
	wire [1:0] w_n207_0;
	wire [2:0] w_n212_0;
	wire [1:0] w_n212_1;
	wire [1:0] w_n213_0;
	wire [1:0] w_n215_0;
	wire [1:0] w_n218_0;
	wire [2:0] w_n224_0;
	wire [1:0] w_n224_1;
	wire [1:0] w_n225_0;
	wire [1:0] w_n229_0;
	wire [2:0] w_n234_0;
	wire [1:0] w_n234_1;
	wire [2:0] w_n237_0;
	wire [1:0] w_n238_0;
	wire [2:0] w_n242_0;
	wire [1:0] w_n243_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n250_0;
	wire [1:0] w_n251_0;
	wire [2:0] w_n255_0;
	wire [1:0] w_n255_1;
	wire [1:0] w_n256_0;
	wire [1:0] w_n257_0;
	wire [1:0] w_n259_0;
	wire [1:0] w_n260_0;
	wire [2:0] w_n261_0;
	wire [2:0] w_n261_1;
	wire [2:0] w_n262_0;
	wire [1:0] w_n269_0;
	wire [1:0] w_n272_0;
	wire [2:0] w_n279_0;
	wire [1:0] w_n279_1;
	wire [1:0] w_n282_0;
	wire [1:0] w_n283_0;
	wire [2:0] w_n292_0;
	wire [1:0] w_n298_0;
	wire [2:0] w_n308_0;
	wire [2:0] w_n308_1;
	wire [1:0] w_n309_0;
	wire [1:0] w_n310_0;
	wire [1:0] w_n312_0;
	wire [1:0] w_n313_0;
	wire [2:0] w_n315_0;
	wire [1:0] w_n321_0;
	wire [2:0] w_n323_0;
	wire [2:0] w_n330_0;
	wire [1:0] w_n333_0;
	wire [1:0] w_n334_0;
	wire [1:0] w_n344_0;
	wire [1:0] w_n347_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n349_0;
	wire [1:0] w_n350_0;
	wire [1:0] w_n351_0;
	wire [2:0] w_n352_0;
	wire [1:0] w_n352_1;
	wire [2:0] w_n354_0;
	wire [1:0] w_n354_1;
	wire [1:0] w_n355_0;
	wire [2:0] w_n356_0;
	wire [1:0] w_n356_1;
	wire [1:0] w_n357_0;
	wire [2:0] w_n367_0;
	wire [1:0] w_n367_1;
	wire [1:0] w_n370_0;
	wire [1:0] w_n375_0;
	wire [1:0] w_n378_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n387_0;
	wire [2:0] w_n388_0;
	wire [2:0] w_n388_1;
	wire [1:0] w_n388_2;
	wire [1:0] w_n394_0;
	wire [1:0] w_n395_0;
	wire [2:0] w_n404_0;
	wire [1:0] w_n405_0;
	wire [1:0] w_n407_0;
	wire [2:0] w_n414_0;
	wire [2:0] w_n417_0;
	wire [1:0] w_n420_0;
	wire [1:0] w_n425_0;
	wire [1:0] w_n426_0;
	wire [1:0] w_n428_0;
	wire [1:0] w_n430_0;
	wire [1:0] w_n435_0;
	wire [2:0] w_n439_0;
	wire [1:0] w_n441_0;
	wire [1:0] w_n445_0;
	wire [1:0] w_n450_0;
	wire [1:0] w_n452_0;
	wire [1:0] w_n456_0;
	wire [1:0] w_n457_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n472_0;
	wire [1:0] w_n473_0;
	wire [2:0] w_n482_0;
	wire [1:0] w_n483_0;
	wire [1:0] w_n494_0;
	wire [1:0] w_n499_0;
	wire [1:0] w_n500_0;
	wire [2:0] w_n503_0;
	wire [2:0] w_n507_0;
	wire [2:0] w_n507_1;
	wire [1:0] w_n507_2;
	wire [1:0] w_n511_0;
	wire [1:0] w_n512_0;
	wire [2:0] w_n514_0;
	wire [1:0] w_n514_1;
	wire [1:0] w_n520_0;
	wire [1:0] w_n533_0;
	wire [1:0] w_n534_0;
	wire [1:0] w_n541_0;
	wire [1:0] w_n542_0;
	wire [1:0] w_n543_0;
	wire [1:0] w_n544_0;
	wire [1:0] w_n548_0;
	wire [1:0] w_n550_0;
	wire [1:0] w_n551_0;
	wire [1:0] w_n559_0;
	wire [1:0] w_n562_0;
	wire [2:0] w_n566_0;
	wire [1:0] w_n566_1;
	wire [2:0] w_n567_0;
	wire [2:0] w_n567_1;
	wire [2:0] w_n567_2;
	wire [2:0] w_n567_3;
	wire [2:0] w_n567_4;
	wire [1:0] w_n567_5;
	wire [1:0] w_n569_0;
	wire [1:0] w_n570_0;
	wire [2:0] w_n571_0;
	wire [2:0] w_n571_1;
	wire [1:0] w_n571_2;
	wire [2:0] w_n572_0;
	wire [1:0] w_n573_0;
	wire [1:0] w_n574_0;
	wire [2:0] w_n576_0;
	wire [1:0] w_n577_0;
	wire [2:0] w_n579_0;
	wire [1:0] w_n579_1;
	wire [2:0] w_n580_0;
	wire [1:0] w_n582_0;
	wire [1:0] w_n584_0;
	wire [1:0] w_n598_0;
	wire [2:0] w_n600_0;
	wire [2:0] w_n600_1;
	wire [2:0] w_n601_0;
	wire [1:0] w_n602_0;
	wire [2:0] w_n604_0;
	wire [2:0] w_n604_1;
	wire [2:0] w_n604_2;
	wire [2:0] w_n605_0;
	wire [2:0] w_n613_0;
	wire [2:0] w_n613_1;
	wire [2:0] w_n614_0;
	wire [2:0] w_n614_1;
	wire [2:0] w_n614_2;
	wire [2:0] w_n614_3;
	wire [2:0] w_n614_4;
	wire [1:0] w_n614_5;
	wire [2:0] w_n618_0;
	wire [2:0] w_n618_1;
	wire [1:0] w_n618_2;
	wire [2:0] w_n619_0;
	wire [2:0] w_n620_0;
	wire [1:0] w_n622_0;
	wire [1:0] w_n624_0;
	wire [2:0] w_n626_0;
	wire [1:0] w_n628_0;
	wire [2:0] w_n629_0;
	wire [2:0] w_n629_1;
	wire [2:0] w_n629_2;
	wire [2:0] w_n629_3;
	wire [2:0] w_n629_4;
	wire [1:0] w_n629_5;
	wire [1:0] w_n630_0;
	wire [1:0] w_n632_0;
	wire [2:0] w_n633_0;
	wire [2:0] w_n633_1;
	wire [2:0] w_n633_2;
	wire [2:0] w_n633_3;
	wire [2:0] w_n633_4;
	wire [2:0] w_n633_5;
	wire [1:0] w_n633_6;
	wire [1:0] w_n634_0;
	wire [1:0] w_n637_0;
	wire [2:0] w_n638_0;
	wire [2:0] w_n638_1;
	wire [2:0] w_n638_2;
	wire [2:0] w_n638_3;
	wire [2:0] w_n638_4;
	wire [2:0] w_n638_5;
	wire [2:0] w_n638_6;
	wire [1:0] w_n638_7;
	wire [2:0] w_n640_0;
	wire [2:0] w_n640_1;
	wire [2:0] w_n640_2;
	wire [2:0] w_n640_3;
	wire [2:0] w_n640_4;
	wire [2:0] w_n640_5;
	wire [2:0] w_n640_6;
	wire [1:0] w_n640_7;
	wire [2:0] w_n646_0;
	wire [2:0] w_n646_1;
	wire [2:0] w_n646_2;
	wire [2:0] w_n646_3;
	wire [2:0] w_n646_4;
	wire [2:0] w_n646_5;
	wire [2:0] w_n646_6;
	wire [1:0] w_n646_7;
	wire [2:0] w_n648_0;
	wire [2:0] w_n648_1;
	wire [2:0] w_n648_2;
	wire [2:0] w_n648_3;
	wire [1:0] w_n648_4;
	wire [1:0] w_n649_0;
	wire [1:0] w_n650_0;
	wire [2:0] w_n651_0;
	wire [2:0] w_n651_1;
	wire [2:0] w_n651_2;
	wire [2:0] w_n651_3;
	wire [2:0] w_n651_4;
	wire [2:0] w_n651_5;
	wire [2:0] w_n651_6;
	wire [1:0] w_n651_7;
	wire [2:0] w_n653_0;
	wire [2:0] w_n653_1;
	wire [2:0] w_n653_2;
	wire [2:0] w_n653_3;
	wire [2:0] w_n653_4;
	wire [2:0] w_n653_5;
	wire [2:0] w_n653_6;
	wire [1:0] w_n653_7;
	wire [2:0] w_n680_0;
	wire [2:0] w_n680_1;
	wire [2:0] w_n680_2;
	wire [2:0] w_n680_3;
	wire [1:0] w_n680_4;
	wire [1:0] w_n682_0;
	wire [2:0] w_n684_0;
	wire [1:0] w_n685_0;
	wire [2:0] w_n690_0;
	wire [1:0] w_n690_1;
	wire [1:0] w_n692_0;
	wire [2:0] w_n703_0;
	wire [1:0] w_n703_1;
	wire [1:0] w_n704_0;
	wire [1:0] w_n718_0;
	wire [1:0] w_n733_0;
	wire [2:0] w_n741_0;
	wire [1:0] w_n741_1;
	wire [1:0] w_n748_0;
	wire [1:0] w_n754_0;
	wire [1:0] w_n759_0;
	wire [1:0] w_n766_0;
	wire [2:0] w_n767_0;
	wire [1:0] w_n767_1;
	wire [2:0] w_n771_0;
	wire [1:0] w_n771_1;
	wire [1:0] w_n772_0;
	wire [1:0] w_n773_0;
	wire [1:0] w_n775_0;
	wire [1:0] w_n777_0;
	wire [1:0] w_n782_0;
	wire [1:0] w_n798_0;
	wire [2:0] w_n802_0;
	wire [1:0] w_n817_0;
	wire [1:0] w_n830_0;
	wire [1:0] w_n833_0;
	wire [2:0] w_n845_0;
	wire [1:0] w_n855_0;
	wire [1:0] w_n860_0;
	wire [1:0] w_n861_0;
	wire [2:0] w_n863_0;
	wire [2:0] w_n869_0;
	wire [1:0] w_n873_0;
	wire [1:0] w_n875_0;
	wire [1:0] w_n884_0;
	wire [1:0] w_n887_0;
	wire [2:0] w_n937_0;
	wire [1:0] w_n959_0;
	wire [2:0] w_n987_0;
	wire [2:0] w_n1029_0;
	wire [1:0] w_n1033_0;
	wire [1:0] w_n1036_0;
	wire [1:0] w_n1039_0;
	wire [1:0] w_n1040_0;
	wire [1:0] w_n1041_0;
	wire [1:0] w_n1043_0;
	wire [1:0] w_n1044_0;
	wire [1:0] w_n1045_0;
	wire [1:0] w_n1048_0;
	wire [2:0] w_n1053_0;
	wire [1:0] w_n1056_0;
	wire [1:0] w_n1062_0;
	wire [1:0] w_n1091_0;
	wire [2:0] w_n1114_0;
	wire [2:0] w_n1159_0;
	wire [1:0] w_n1161_0;
	wire [1:0] w_n1164_0;
	wire [1:0] w_n1168_0;
	wire [1:0] w_n1170_0;
	wire [1:0] w_n1177_0;
	wire [1:0] w_n1178_0;
	wire [1:0] w_n1179_0;
	wire [1:0] w_n1184_0;
	wire w_dff_B_ynZ5YnHd1_1;
	wire w_dff_B_xrbgYCPy3_1;
	wire w_dff_B_Pb9h1aHH6_1;
	wire w_dff_B_q71j2OGx8_0;
	wire w_dff_B_udMr7RwF5_0;
	wire w_dff_B_9z3KwyPI0_1;
	wire w_dff_B_hbZGDMrg3_1;
	wire w_dff_B_zCONiVVC8_0;
	wire w_dff_B_WG4S1uzv0_1;
	wire w_dff_B_e4hfOEbK7_1;
	wire w_dff_B_ZbTG51FI0_1;
	wire w_dff_B_t6YLDsJf6_1;
	wire w_dff_B_JHWAjE433_1;
	wire w_dff_B_Ws5GYjEw0_1;
	wire w_dff_B_xB1RSBq43_1;
	wire w_dff_B_rpt2txpk2_1;
	wire w_dff_B_CXcfAsYh9_1;
	wire w_dff_B_8FKXV26O9_1;
	wire w_dff_B_N9BGqFE76_1;
	wire w_dff_B_VtB1sIV48_1;
	wire w_dff_B_mL75RmLX6_1;
	wire w_dff_B_N6Lw2OXO1_1;
	wire w_dff_B_S51GjHWv7_1;
	wire w_dff_B_prADZb7W6_1;
	wire w_dff_B_fHOwcBxf0_0;
	wire w_dff_B_Jvtvvq538_0;
	wire w_dff_B_3M27IcLs1_0;
	wire w_dff_B_I7gb4k2j7_0;
	wire w_dff_B_Q0OU1C3u7_0;
	wire w_dff_B_cFVEODNb8_0;
	wire w_dff_B_jOwdAJi95_0;
	wire w_dff_B_1m3mqAGi7_0;
	wire w_dff_B_jnU9okez8_0;
	wire w_dff_B_oyimtRpZ0_0;
	wire w_dff_B_EAroxufK9_0;
	wire w_dff_B_0OMFfL6U4_0;
	wire w_dff_B_kUcR5PsM8_0;
	wire w_dff_B_mOPif1fF3_0;
	wire w_dff_B_bLAKcHKe6_0;
	wire w_dff_B_SPiR5Gfq0_0;
	wire w_dff_B_40lhxiL72_0;
	wire w_dff_B_U7NvSjUt8_0;
	wire w_dff_B_c7m59G2O8_0;
	wire w_dff_B_lUWwwYmu7_0;
	wire w_dff_B_H9wIZlfo4_0;
	wire w_dff_B_1EC4mkL36_0;
	wire w_dff_B_sNMgBzfb4_0;
	wire w_dff_B_dYU2wWJk4_0;
	wire w_dff_B_KCoETwj26_0;
	wire w_dff_B_347UTkUS3_0;
	wire w_dff_B_6RgXlCOo7_0;
	wire w_dff_B_huhjNFeY1_0;
	wire w_dff_B_1TU4w3Jl0_0;
	wire w_dff_B_fHVw0UMH6_0;
	wire w_dff_B_eyzArHIQ3_0;
	wire w_dff_B_sq671Pcx0_0;
	wire w_dff_A_rwvnvfyK3_1;
	wire w_dff_A_Gv04fcjb4_1;
	wire w_dff_A_fqJ0YkIr5_1;
	wire w_dff_B_AVjPnWhX9_0;
	wire w_dff_B_KpnIjPAZ5_1;
	wire w_dff_B_TwPIIMOM4_1;
	wire w_dff_B_cYnRrgGN4_1;
	wire w_dff_B_QsOWg22Z7_1;
	wire w_dff_B_9puWg91t9_1;
	wire w_dff_B_pdUogo6x0_1;
	wire w_dff_B_7P58rKmj8_1;
	wire w_dff_B_k6DQEmqy0_1;
	wire w_dff_B_KAQ6kGp86_1;
	wire w_dff_B_mfgfwltP7_1;
	wire w_dff_B_IiyhBUHa3_1;
	wire w_dff_B_xGeWlfHP1_1;
	wire w_dff_B_F7txf4wl7_1;
	wire w_dff_B_FMWNkpb43_1;
	wire w_dff_B_rDYpXZLK3_1;
	wire w_dff_B_F6XMW7zK9_1;
	wire w_dff_B_mCBbpt9J8_1;
	wire w_dff_B_mirvIYcZ8_1;
	wire w_dff_B_NNpb1PAP1_0;
	wire w_dff_A_VV0G5Xfi3_0;
	wire w_dff_B_MOGcl5UV4_1;
	wire w_dff_B_pLHv3hyp7_1;
	wire w_dff_B_HfCFKUce9_1;
	wire w_dff_B_oUye4lm36_1;
	wire w_dff_B_ccCmc88O3_1;
	wire w_dff_B_Oyyhcu7R7_1;
	wire w_dff_B_3yH9xtxp0_1;
	wire w_dff_B_fVa69rRd2_1;
	wire w_dff_B_ISIuAwLU4_1;
	wire w_dff_B_MiPcuc7d1_1;
	wire w_dff_B_i56ZNTFD4_1;
	wire w_dff_B_Yg9QwWVa5_1;
	wire w_dff_B_uh65DdRn2_1;
	wire w_dff_B_lkpLCRPL1_1;
	wire w_dff_B_OHSAB6HG1_1;
	wire w_dff_B_j1VOoZqi5_1;
	wire w_dff_B_LFokzkIg5_1;
	wire w_dff_B_GcFzOQHz3_1;
	wire w_dff_B_CP8Qiqn29_1;
	wire w_dff_B_ZhLnKxlj9_1;
	wire w_dff_B_CE4hUIpS1_1;
	wire w_dff_B_yqcq7O9G2_1;
	wire w_dff_B_FoniNyag2_1;
	wire w_dff_B_1tFGnpYG7_1;
	wire w_dff_B_iQ6wkzeT9_1;
	wire w_dff_B_bFmJ5DuS4_1;
	wire w_dff_B_HkKtItOb4_1;
	wire w_dff_B_LvvcfnQ51_1;
	wire w_dff_B_9RlCuJE84_1;
	wire w_dff_B_jy3F7UiK7_1;
	wire w_dff_B_NZyNgzld3_0;
	wire w_dff_B_HSI4VBVl1_0;
	wire w_dff_A_NlX6DN6V3_1;
	wire w_dff_B_4Jva4wWJ7_1;
	wire w_dff_B_Yp126YZE0_1;
	wire w_dff_B_WjTJ54NR6_1;
	wire w_dff_B_KxS9j7Ct8_1;
	wire w_dff_B_ooJVhPtl4_1;
	wire w_dff_B_Swa2GdbL7_1;
	wire w_dff_B_Gp7nP9S90_1;
	wire w_dff_B_XY1pnQ3s1_1;
	wire w_dff_B_JRXFOd4X2_1;
	wire w_dff_B_VWEfQuec5_1;
	wire w_dff_B_hkHyVgjx6_1;
	wire w_dff_B_ElenyalL8_1;
	wire w_dff_B_LL1UC17n5_1;
	wire w_dff_B_onvbfAJl0_1;
	wire w_dff_B_7GqXLUBk4_1;
	wire w_dff_B_TJrrlA0t2_1;
	wire w_dff_B_QJSsaXGL6_1;
	wire w_dff_B_AvtvG76D6_1;
	wire w_dff_B_4YD8iW2l7_1;
	wire w_dff_B_EZATfHu78_1;
	wire w_dff_B_rPPpTlqc4_1;
	wire w_dff_B_YTkb88oz0_1;
	wire w_dff_B_hRMMJKQr8_1;
	wire w_dff_B_0ug2eyZl8_1;
	wire w_dff_B_ep09lUf91_1;
	wire w_dff_B_tCTyTYsZ1_1;
	wire w_dff_B_nNZ0GruW3_1;
	wire w_dff_B_Sb1jYBl36_1;
	wire w_dff_B_FoKlvykA8_1;
	wire w_dff_B_92NfxHvE5_1;
	wire w_dff_B_akcrgVn10_1;
	wire w_dff_B_LkkgUbfh9_1;
	wire w_dff_B_DdU91plB6_1;
	wire w_dff_B_NkrRuS4v6_1;
	wire w_dff_B_kGzofVkP0_1;
	wire w_dff_B_FkDjUroM5_1;
	wire w_dff_B_a5qsdpPl0_1;
	wire w_dff_B_geszqRin9_1;
	wire w_dff_B_XPPkmska3_1;
	wire w_dff_B_q6xrlLHy0_1;
	wire w_dff_B_u4YvyHno2_1;
	wire w_dff_B_oiUAum5a2_1;
	wire w_dff_B_Dj4EA9br3_1;
	wire w_dff_B_AVlSSToM7_1;
	wire w_dff_B_2wh4DxzF3_1;
	wire w_dff_B_kqcm35Et6_1;
	wire w_dff_B_9Lneeevi3_1;
	wire w_dff_B_SccqQPVF0_1;
	wire w_dff_B_DpKEq05N3_1;
	wire w_dff_B_CkLQh78X3_1;
	wire w_dff_B_UM0Lkz9K1_1;
	wire w_dff_B_PsF3JsDJ6_1;
	wire w_dff_A_ILeDfsuw7_1;
	wire w_dff_A_pxawqQ3a3_1;
	wire w_dff_A_D2wsoZKF9_1;
	wire w_dff_A_Inn18rz07_1;
	wire w_dff_A_FXi9Q7wi5_1;
	wire w_dff_A_AIxfc44U1_1;
	wire w_dff_A_iS0tUClF8_1;
	wire w_dff_A_OXTVixPV4_1;
	wire w_dff_A_kx9jF2yE1_1;
	wire w_dff_A_f5EBb4x37_1;
	wire w_dff_A_KaqR2Yu58_1;
	wire w_dff_A_pEQqklk58_1;
	wire w_dff_A_PLmr5Ubr7_1;
	wire w_dff_A_fApyZn363_1;
	wire w_dff_A_sTXFaWHj3_1;
	wire w_dff_A_OmsWeqas0_1;
	wire w_dff_A_KKksWgzY0_1;
	wire w_dff_A_hFSP9obF9_1;
	wire w_dff_A_YzSysODz5_1;
	wire w_dff_A_YGXs8kLG2_1;
	wire w_dff_A_Q9MBdEoW4_1;
	wire w_dff_A_oiDLfZe90_1;
	wire w_dff_A_FqziWXfs7_1;
	wire w_dff_A_ZZi18SpG5_1;
	wire w_dff_A_HODbHNBK8_1;
	wire w_dff_A_cebzNpmp2_1;
	wire w_dff_A_5IgX0xir6_1;
	wire w_dff_A_vyPi09V38_1;
	wire w_dff_A_9BDr473e2_1;
	wire w_dff_A_5ynAQ5FP8_1;
	wire w_dff_A_3QWOje9G8_1;
	wire w_dff_A_Dw1jRvsm7_1;
	wire w_dff_A_rYyvzy0h3_1;
	wire w_dff_A_CK34gOZr6_1;
	wire w_dff_A_JoU1LoiZ6_1;
	wire w_dff_A_348Mxk9U0_1;
	wire w_dff_A_WvnTDaGw9_1;
	wire w_dff_A_Y29Mh8P43_1;
	wire w_dff_A_34Hh8ZaC5_1;
	wire w_dff_A_6j09Spgg0_1;
	wire w_dff_A_ksMFUMwP3_1;
	wire w_dff_A_MagO818t6_1;
	wire w_dff_A_VdYA3Qjv1_1;
	wire w_dff_A_mRX1fxRK9_1;
	wire w_dff_A_Zm5e9g7P5_1;
	wire w_dff_A_O5r1H6216_1;
	wire w_dff_A_1gOiWsKn6_1;
	wire w_dff_A_3dzdKn6K9_1;
	wire w_dff_A_agWKvC6d4_1;
	wire w_dff_A_6kZ25O5i0_1;
	wire w_dff_A_pKK2AQ8o9_1;
	wire w_dff_A_WWo1OGan9_1;
	wire w_dff_B_9IOKiBPx3_0;
	wire w_dff_B_AmBrGIhR0_0;
	wire w_dff_B_M6ZwTmD70_0;
	wire w_dff_B_8kcLwFOF0_0;
	wire w_dff_B_FXcr77hx2_0;
	wire w_dff_B_yGoT3d7y9_0;
	wire w_dff_B_yX29Iaal8_0;
	wire w_dff_B_2PGtm2bd1_0;
	wire w_dff_B_b2c5cbPb0_0;
	wire w_dff_B_etvtQCR71_0;
	wire w_dff_B_xIkmAwaF3_0;
	wire w_dff_B_14GPHnhZ5_0;
	wire w_dff_B_1bzYNzPb2_0;
	wire w_dff_B_LpNv12ZK0_0;
	wire w_dff_B_2YJIO6bP1_1;
	wire w_dff_B_TVj34eH45_1;
	wire w_dff_B_a2suvZFA7_1;
	wire w_dff_B_vCoqdJZO5_1;
	wire w_dff_B_qwclzErK5_1;
	wire w_dff_B_fmH78Oyd7_1;
	wire w_dff_B_WQ2yBKPr1_1;
	wire w_dff_B_jY1lzMXy0_1;
	wire w_dff_B_AgLcT7f60_1;
	wire w_dff_B_UcePQ7nO9_1;
	wire w_dff_B_6p2TD6t02_1;
	wire w_dff_B_vIG23IUk8_0;
	wire w_dff_B_PAQIdhXW3_1;
	wire w_dff_B_seMa3UNg8_1;
	wire w_dff_B_SRmOgYXh7_0;
	wire w_dff_B_q2JofDlD2_1;
	wire w_dff_B_TdsIXP264_0;
	wire w_dff_B_7SvklPTh7_1;
	wire w_dff_B_eqVYmkLb8_1;
	wire w_dff_B_sDZ488Y14_1;
	wire w_dff_B_C7SLVvkC7_1;
	wire w_dff_B_dfAUOGxt2_1;
	wire w_dff_B_Vn3lvBwj6_0;
	wire w_dff_B_f72n7whF8_0;
	wire w_dff_B_dIaU5zlH8_0;
	wire w_dff_B_jIOqZmB33_1;
	wire w_dff_A_AQjdfNJy3_1;
	wire w_dff_A_RYql7SpD6_1;
	wire w_dff_A_M7cIU7oP7_1;
	wire w_dff_A_g66tHovf5_1;
	wire w_dff_A_OD4kqRMI8_1;
	wire w_dff_A_gBPuj7GC2_1;
	wire w_dff_A_4E3ZfTzQ6_1;
	wire w_dff_A_NvbC047F9_1;
	wire w_dff_B_t3YZ9YNv1_0;
	wire w_dff_B_QnLRwrnw8_0;
	wire w_dff_B_nCJnhmBj5_1;
	wire w_dff_B_6uSLkFyL4_1;
	wire w_dff_B_vXSWPy6C5_1;
	wire w_dff_B_SfkCUuyu4_1;
	wire w_dff_B_E6LEHatv5_1;
	wire w_dff_B_9mUJs9TO4_1;
	wire w_dff_B_uCU5BhTa0_1;
	wire w_dff_B_4HRWX6FB9_1;
	wire w_dff_A_Iys6T4A83_1;
	wire w_dff_A_i2Gbulu39_1;
	wire w_dff_A_JEo4JplL4_1;
	wire w_dff_B_MzbukCNK4_0;
	wire w_dff_B_s8dXbXUQ9_0;
	wire w_dff_B_qQRl7ORa8_0;
	wire w_dff_B_6xmW4B3f8_0;
	wire w_dff_B_mDHgUgxZ7_0;
	wire w_dff_B_uxtRcIsy7_0;
	wire w_dff_B_XZ06BLZb3_0;
	wire w_dff_B_soZKWZSH9_1;
	wire w_dff_B_DVJbvddl0_1;
	wire w_dff_B_t14mZ7Wt6_1;
	wire w_dff_B_TKIzkszB4_1;
	wire w_dff_B_YmC8U9uy1_1;
	wire w_dff_B_NEDV5Qq39_1;
	wire w_dff_B_O181L9ZS5_1;
	wire w_dff_B_4uF57oCj4_1;
	wire w_dff_B_1N7T31AP7_0;
	wire w_dff_A_L99Ypaxn3_1;
	wire w_dff_A_qSzqW1xY9_1;
	wire w_dff_B_Go0Z7t8Q7_1;
	wire w_dff_B_ED5gFEA37_1;
	wire w_dff_A_vvtvW8iE0_1;
	wire w_dff_A_XTyFZhMw1_1;
	wire w_dff_A_PocpNMT54_1;
	wire w_dff_A_Mo2Sva0V8_1;
	wire w_dff_A_Ney4EExm3_1;
	wire w_dff_A_ggCuepbO8_2;
	wire w_dff_A_mAfW15vs4_2;
	wire w_dff_A_z0M12BCP9_2;
	wire w_dff_B_nasyWk486_3;
	wire w_dff_B_p5X6eS3F5_3;
	wire w_dff_A_pXjCxg399_1;
	wire w_dff_B_B2gUorcj5_0;
	wire w_dff_B_6UKKzey64_0;
	wire w_dff_B_8GJiAsB33_0;
	wire w_dff_B_ELkhX7KN4_0;
	wire w_dff_B_t3fUfV9F2_0;
	wire w_dff_B_QKTeOl1e3_0;
	wire w_dff_B_m88xIWPw1_1;
	wire w_dff_B_8gPGC0Fu6_1;
	wire w_dff_B_AaXitViX9_0;
	wire w_dff_B_Jp6T2fN52_1;
	wire w_dff_B_CLm81odN6_1;
	wire w_dff_B_CkUcccqP4_1;
	wire w_dff_B_eEs0hkWs3_1;
	wire w_dff_B_4qBjV5F97_1;
	wire w_dff_B_8UkSvFVL7_1;
	wire w_dff_B_0ccWCGf52_1;
	wire w_dff_B_mpEZYCdW1_1;
	wire w_dff_B_qpyT6lIT2_0;
	wire w_dff_B_MemRcEoA6_1;
	wire w_dff_A_6fwpVXDc5_1;
	wire w_dff_B_kYAY9cCE3_2;
	wire w_dff_B_DvAMv9hV5_2;
	wire w_dff_B_osGoo7l30_2;
	wire w_dff_A_ctnulHmK7_0;
	wire w_dff_A_wsO9wAL21_0;
	wire w_dff_A_peMkkoOB8_0;
	wire w_dff_A_lBHOKvxP8_1;
	wire w_dff_A_lN4oWSO32_1;
	wire w_dff_A_zJXLAHkh2_1;
	wire w_dff_A_6XkRdgC42_1;
	wire w_dff_A_UPHyR0D85_1;
	wire w_dff_A_IId9JDG40_1;
	wire w_dff_A_8vlSL97B9_1;
	wire w_dff_A_TkQ626Ep1_1;
	wire w_dff_A_Eq3uJins8_1;
	wire w_dff_A_e0sy6Ty21_1;
	wire w_dff_A_gps9NreM1_1;
	wire w_dff_B_kwjGrP3X0_0;
	wire w_dff_B_pgpnDPot6_0;
	wire w_dff_B_bbDuC9hg5_1;
	wire w_dff_B_tofmwiV27_1;
	wire w_dff_B_O2CbvBPK1_1;
	wire w_dff_B_Q26YwzAT5_1;
	wire w_dff_B_zb8rwFO40_1;
	wire w_dff_B_aPConhyT7_1;
	wire w_dff_B_DuplOqxG0_0;
	wire w_dff_B_wko8F1q72_1;
	wire w_dff_B_zOWbBvLs7_0;
	wire w_dff_A_obDpq9Wc4_0;
	wire w_dff_A_KtaDcr6o2_1;
	wire w_dff_A_YS7cNnUb6_1;
	wire w_dff_A_76GUKfTK9_2;
	wire w_dff_A_6ypzyubQ1_2;
	wire w_dff_A_Vep6fdi22_0;
	wire w_dff_B_codiG89P1_1;
	wire w_dff_B_a6D3DV1K1_1;
	wire w_dff_B_Xsm9xh5N4_1;
	wire w_dff_B_3wtckWVD5_1;
	wire w_dff_B_K3A7R6M86_1;
	wire w_dff_B_GHDibozC2_1;
	wire w_dff_A_vSDsysS30_0;
	wire w_dff_B_gWM7VLxp7_1;
	wire w_dff_A_W5Ogq3VP7_1;
	wire w_dff_A_I33LFH801_1;
	wire w_dff_A_JrOA0bvg9_1;
	wire w_dff_A_jLEg05hM1_1;
	wire w_dff_A_0KyCEXJH5_1;
	wire w_dff_A_JEG8Zf214_1;
	wire w_dff_A_196A7o9u3_2;
	wire w_dff_A_XwUXAtVT4_2;
	wire w_dff_A_jI0YuI4j5_2;
	wire w_dff_A_uPxZXOvn9_0;
	wire w_dff_B_eapyrZRK4_1;
	wire w_dff_B_s7xqtnNw8_1;
	wire w_dff_B_fPSynR9i2_1;
	wire w_dff_B_mDqj1ljP3_1;
	wire w_dff_B_IOgjobww9_1;
	wire w_dff_B_GY5YBRnb7_1;
	wire w_dff_B_uAVr2jzw7_1;
	wire w_dff_B_G3EgqqmC4_1;
	wire w_dff_A_n48ZFbuf3_1;
	wire w_dff_A_NLrLty692_0;
	wire w_dff_B_OKK6X1Xx9_1;
	wire w_dff_A_ETyHwJZZ6_0;
	wire w_dff_A_5GUiSh0H6_0;
	wire w_dff_A_0l8nIW9H9_0;
	wire w_dff_A_o7WcTBV71_2;
	wire w_dff_A_kLHkaF9J4_2;
	wire w_dff_A_PzhApn8n0_2;
	wire w_dff_B_HPDhHTvl3_1;
	wire w_dff_A_Zh3LZqwt0_1;
	wire w_dff_A_Cqut5Hol2_0;
	wire w_dff_B_QuYqfTew0_2;
	wire w_dff_B_zdMtXarI8_2;
	wire w_dff_A_nzPHUKnK0_0;
	wire w_dff_A_UbfmXpYv9_0;
	wire w_dff_A_MpttRNvE6_0;
	wire w_dff_A_VvKWeSn83_0;
	wire w_dff_B_IF4NufHq0_2;
	wire w_dff_A_UUzuMJy37_1;
	wire w_dff_A_FtBHihML4_0;
	wire w_dff_A_D96Dk9uZ6_0;
	wire w_dff_A_Z55c4btw4_0;
	wire w_dff_A_aZSTRNcR3_0;
	wire w_dff_A_Fv85uBtG6_0;
	wire w_dff_A_M6D2HWEZ2_0;
	wire w_dff_A_EPTeD56R1_0;
	wire w_dff_B_wMi9uOsJ9_0;
	wire w_dff_B_4ZkfhsuZ8_0;
	wire w_dff_B_Uz0lf2br0_0;
	wire w_dff_B_CrutxyLd1_0;
	wire w_dff_B_kSpOWxbn2_0;
	wire w_dff_B_pgnI3aQB0_0;
	wire w_dff_B_PQ6gA8B69_0;
	wire w_dff_B_EGXmiC7J3_0;
	wire w_dff_B_kfpXk8sW5_0;
	wire w_dff_B_hFunX7DE5_0;
	wire w_dff_B_Alqur92y5_0;
	wire w_dff_B_mz2u4UQD9_1;
	wire w_dff_B_UeGz7vFO4_1;
	wire w_dff_B_VI8urFpX0_1;
	wire w_dff_B_qI34WO6Q9_1;
	wire w_dff_B_WtBCHLNl5_1;
	wire w_dff_B_I96gKeLI7_1;
	wire w_dff_B_OckltRcT2_1;
	wire w_dff_B_cBcHvVMM1_1;
	wire w_dff_B_c4620I9v0_1;
	wire w_dff_B_PXEpW0aS6_1;
	wire w_dff_B_KZ9JUhvf0_1;
	wire w_dff_A_YWRtBQ7V5_0;
	wire w_dff_B_W3iuT2RV1_3;
	wire w_dff_B_8O9yucme6_3;
	wire w_dff_B_aXjaDQ4M0_3;
	wire w_dff_A_5O647Yik4_0;
	wire w_dff_A_2F2Oudh08_1;
	wire w_dff_A_XtQxDIXw9_1;
	wire w_dff_A_LOuZt1hJ2_1;
	wire w_dff_A_90HwEfKC6_1;
	wire w_dff_B_FptpMnwi7_1;
	wire w_dff_B_JeNg2Ljz2_1;
	wire w_dff_A_0yyXrzMH2_0;
	wire w_dff_A_JIa7x4XB8_1;
	wire w_dff_A_oAPZEv3J5_2;
	wire w_dff_B_YPROuvuL0_1;
	wire w_dff_B_JxhsXLS99_1;
	wire w_dff_A_bvHEwYPn0_1;
	wire w_dff_A_NcO9Sjbo1_2;
	wire w_dff_A_6eiINvJZ3_2;
	wire w_dff_A_mdZgBqlb2_2;
	wire w_dff_A_TJwIehfe4_2;
	wire w_dff_B_5c9wZdRa0_0;
	wire w_dff_B_IWopkhLh1_0;
	wire w_dff_B_ZNbHQtQH4_0;
	wire w_dff_B_hQIfFVma4_0;
	wire w_dff_A_FcdkyXoc5_1;
	wire w_dff_A_Oh91G41R4_1;
	wire w_dff_A_SKxkA4gY1_2;
	wire w_dff_B_9sgztSk90_1;
	wire w_dff_B_bH0fzxpY2_1;
	wire w_dff_B_mqMdDvCO3_1;
	wire w_dff_B_BhPBEMs71_1;
	wire w_dff_A_MchgcMM65_0;
	wire w_dff_A_vb2mpHcf6_0;
	wire w_dff_A_SfnC8UI12_2;
	wire w_dff_A_0msoXEw23_2;
	wire w_dff_A_IMx4AmGF3_2;
	wire w_dff_A_gwvRXqe98_2;
	wire w_dff_A_OE7sgIuQ1_2;
	wire w_dff_B_lrgl6soP5_0;
	wire w_dff_A_xc49V2yN9_1;
	wire w_dff_B_Vz7Z6xjQ8_1;
	wire w_dff_B_947c0t5M6_1;
	wire w_dff_B_EwVOvqLO1_1;
	wire w_dff_A_ZrygzSyX5_0;
	wire w_dff_A_9QBz8RYs5_0;
	wire w_dff_A_e5E483ow0_0;
	wire w_dff_A_Q2U1rWYC3_0;
	wire w_dff_A_UDsUAlsV2_0;
	wire w_dff_A_g5xzbAJs4_0;
	wire w_dff_A_vgLnRoeq5_0;
	wire w_dff_A_UydSEI1R7_0;
	wire w_dff_A_akZQpuOp2_0;
	wire w_dff_B_rh4QLE558_1;
	wire w_dff_B_WE9fOSRN4_1;
	wire w_dff_B_UcjOiyLY9_0;
	wire w_dff_B_7B0RoYiB7_1;
	wire w_dff_A_EmMFb6Ux0_0;
	wire w_dff_A_zDloW7fa1_0;
	wire w_dff_A_YTi8Dgu26_0;
	wire w_dff_B_hVfg89iI1_0;
	wire w_dff_B_yiifLGK53_0;
	wire w_dff_B_vhBtoQwU7_0;
	wire w_dff_B_iNYb9PqW3_0;
	wire w_dff_B_6axqDvYD6_0;
	wire w_dff_B_a4VQMPiO2_0;
	wire w_dff_B_yOlpVy2k4_0;
	wire w_dff_B_vaDBoLY89_0;
	wire w_dff_B_QeiMDT8I5_1;
	wire w_dff_A_czxibepF3_0;
	wire w_dff_A_YimUmIaL6_0;
	wire w_dff_A_40nzIkoe9_0;
	wire w_dff_A_yXd4Uuu18_0;
	wire w_dff_A_YXZheSm79_0;
	wire w_dff_A_D0lwcCld0_0;
	wire w_dff_A_QGPlReu91_0;
	wire w_dff_A_82kfVSlJ5_0;
	wire w_dff_A_vqqHyQld4_0;
	wire w_dff_A_SCvhVDYY6_0;
	wire w_dff_A_vp9rvH7c9_0;
	wire w_dff_A_xgxKAMrc7_1;
	wire w_dff_A_W6tDfEn78_1;
	wire w_dff_A_sWjbEFMw4_1;
	wire w_dff_A_3WDz4osr6_1;
	wire w_dff_A_xlixRGKu3_1;
	wire w_dff_A_VM8dThXw0_1;
	wire w_dff_A_pOrw0prw5_1;
	wire w_dff_A_eWucBi366_1;
	wire w_dff_A_u5hNhmDB3_1;
	wire w_dff_A_Dz7BMP8p7_1;
	wire w_dff_A_om1uan588_1;
	wire w_dff_B_OhgEfmRx3_0;
	wire w_dff_B_c4JQbR9H5_0;
	wire w_dff_B_Qgk1zIAq1_1;
	wire w_dff_B_oCrH7Lgx0_1;
	wire w_dff_B_LPi0uogA1_1;
	wire w_dff_A_n5GY4sdo6_0;
	wire w_dff_A_9ipMDwCo7_0;
	wire w_dff_A_1uyzNcr30_0;
	wire w_dff_A_tpD3wjjN6_0;
	wire w_dff_B_5UdxwxRG3_2;
	wire w_dff_B_l3j8OZvY8_1;
	wire w_dff_A_97lxGxD29_1;
	wire w_dff_B_WfF5hDW57_3;
	wire w_dff_B_wPFcyzwI9_3;
	wire w_dff_B_EDPlRGQZ8_3;
	wire w_dff_B_yO4odglo3_1;
	wire w_dff_B_CsOHDHJM3_1;
	wire w_dff_B_0YsiHeIC6_0;
	wire w_dff_A_nbkZK3gz7_0;
	wire w_dff_A_226JHW4E9_0;
	wire w_dff_A_JH3Amltv7_0;
	wire w_dff_A_TXIsUPNy8_0;
	wire w_dff_A_39XrxDvY6_0;
	wire w_dff_A_iOdcPdRN2_0;
	wire w_dff_A_mjcIPlYI2_1;
	wire w_dff_A_W95K5KKG3_1;
	wire w_dff_A_ByPGuawY7_1;
	wire w_dff_A_qHvtVqkT7_2;
	wire w_dff_B_vI1890VH2_0;
	wire w_dff_B_gmxxOQzu0_0;
	wire w_dff_B_tIvO4YzW4_0;
	wire w_dff_B_oEGQHARh0_0;
	wire w_dff_B_LzxIiMpc8_0;
	wire w_dff_A_sdMQGsvz6_0;
	wire w_dff_A_ruwX4sgZ3_1;
	wire w_dff_A_wWlgZZ4S2_1;
	wire w_dff_A_RLsYC9xP9_1;
	wire w_dff_A_t9pnQjqb7_1;
	wire w_dff_A_1cZgT8FT3_1;
	wire w_dff_A_aYTPkeyl4_1;
	wire w_dff_A_dTjGelrD5_1;
	wire w_dff_A_LR5W7OFQ5_1;
	wire w_dff_B_qhibm7nF7_1;
	wire w_dff_B_IAH45NQo8_1;
	wire w_dff_A_UZ27vMAF8_1;
	wire w_dff_A_GdC3iBAj1_1;
	wire w_dff_A_PSySrwr68_1;
	wire w_dff_B_2DwCmg7O1_1;
	wire w_dff_B_2c83vRPV0_0;
	wire w_dff_B_aEtb0mcV1_1;
	wire w_dff_A_pgfK9uma1_0;
	wire w_dff_A_34WEawZK6_0;
	wire w_dff_B_gHQTSLrz0_2;
	wire w_dff_B_jLV0ghFw1_0;
	wire w_dff_B_pGicBI5G6_1;
	wire w_dff_A_jxVQlUsh1_1;
	wire w_dff_A_u0zShoW77_1;
	wire w_dff_A_Mi458JfJ5_0;
	wire w_dff_A_LB2BJLy78_1;
	wire w_dff_A_CwoR9y7N7_2;
	wire w_dff_A_uEuoVxFA7_0;
	wire w_dff_A_NDct26XZ8_1;
	wire w_dff_A_zzA9gOhC2_2;
	wire w_dff_A_7H2DEj1c7_1;
	wire w_dff_A_Lz3Y5PGp7_1;
	wire w_dff_B_hpwzkZhz7_2;
	wire w_dff_B_Dq2Xk9Zs5_2;
	wire w_dff_B_cRQ7BKJr4_1;
	wire w_dff_B_76G1R80I7_1;
	wire w_dff_B_MW8Bjtcc4_0;
	wire w_dff_B_EEa8Na864_0;
	wire w_dff_B_lnQ8HUb74_0;
	wire w_dff_B_L79gYsFG0_0;
	wire w_dff_B_JC0CyPB34_0;
	wire w_dff_B_gNQYeVZj1_0;
	wire w_dff_B_Og2VNfOO6_0;
	wire w_dff_B_Q6ihH8472_1;
	wire w_dff_B_p0uyDgDK6_1;
	wire w_dff_B_LpW2euEs6_1;
	wire w_dff_B_7g4tZBYO7_1;
	wire w_dff_B_7whsfyG25_1;
	wire w_dff_B_Y3pctb3y9_1;
	wire w_dff_A_cUW9NY2e1_2;
	wire w_dff_B_QGb6dHNc8_1;
	wire w_dff_A_p726uaCi3_1;
	wire w_dff_B_oesYkrT41_1;
	wire w_dff_B_1o1k8E266_1;
	wire w_dff_B_2fzj4tTD7_1;
	wire w_dff_B_00tOmlcV1_1;
	wire w_dff_B_yRAbqoPj3_1;
	wire w_dff_B_3538W6Se4_1;
	wire w_dff_A_n1qPfFTw9_0;
	wire w_dff_A_ceXLqub56_0;
	wire w_dff_A_AvSlXyCe7_0;
	wire w_dff_A_0FXdgbTT2_2;
	wire w_dff_A_Fweb03Sm6_1;
	wire w_dff_A_zkS5FPqg8_1;
	wire w_dff_A_N4Y2Mr3N2_1;
	wire w_dff_A_0JtXnC2e8_2;
	wire w_dff_A_q93wIPSs7_2;
	wire w_dff_A_nLJPHWsy8_2;
	wire w_dff_B_lm0hFwU34_1;
	wire w_dff_B_LY7bYntw8_1;
	wire w_dff_B_AwPZqyvy3_0;
	wire w_dff_A_NxLNoeNl9_0;
	wire w_dff_B_DZJ2aS4s0_0;
	wire w_dff_B_bmkZyDxZ1_1;
	wire w_dff_B_JvjjaOGR2_1;
	wire w_dff_B_P5QO7Brl0_1;
	wire w_dff_B_wnA5m0lB7_1;
	wire w_dff_B_vujsMn4w8_1;
	wire w_dff_B_pMhcoQm33_1;
	wire w_dff_B_u5krdrV44_1;
	wire w_dff_B_vSBWEpvC8_1;
	wire w_dff_B_DrZ5NFFL2_1;
	wire w_dff_B_EYZKU5ko9_1;
	wire w_dff_B_2qZ3BbhQ9_0;
	wire w_dff_A_ufV6lJRQ8_0;
	wire w_dff_A_oowgKUsw6_0;
	wire w_dff_A_lbuSIHpA8_0;
	wire w_dff_A_gfTtQOA63_2;
	wire w_dff_B_YAk8KxDc6_1;
	wire w_dff_B_FRUsGpKl3_1;
	wire w_dff_B_500HLwzz0_1;
	wire w_dff_B_8phYCkmE0_1;
	wire w_dff_B_ZAfep1yA9_1;
	wire w_dff_B_drb9tgyI3_0;
	wire w_dff_A_6SXdzCnI2_1;
	wire w_dff_A_WfzRtcFC0_1;
	wire w_dff_A_CrFou7NL0_0;
	wire w_dff_A_AcbZ4Tay0_0;
	wire w_dff_A_JS0Y1SzS9_0;
	wire w_dff_B_tascgUPq3_0;
	wire w_dff_B_olPxfAgE5_0;
	wire w_dff_A_zBDMi8J16_1;
	wire w_dff_A_41v9qUwg2_1;
	wire w_dff_A_jsVmobp23_1;
	wire w_dff_A_OG8upKwM1_1;
	wire w_dff_B_tDkrTTgd8_0;
	wire w_dff_B_XrN8ujoq0_0;
	wire w_dff_B_JiavlIFh1_0;
	wire w_dff_A_yxo8XTQb4_1;
	wire w_dff_A_nBTj7VM28_1;
	wire w_dff_B_reR9chzK7_0;
	wire w_dff_B_lryXG1jZ6_1;
	wire w_dff_B_dnmNCXeR4_1;
	wire w_dff_B_tbPUkQaw0_1;
	wire w_dff_B_3oQ96Ro83_1;
	wire w_dff_B_PwACYx4m9_1;
	wire w_dff_B_wcfSg0N25_1;
	wire w_dff_B_RxJFYEeT9_1;
	wire w_dff_B_evK5ALlS6_0;
	wire w_dff_A_1gSwhNQf5_0;
	wire w_dff_B_xumulVta2_1;
	wire w_dff_A_RooK4Q3D0_0;
	wire w_dff_A_bG2djZ6W8_0;
	wire w_dff_A_QDZZMnUA1_0;
	wire w_dff_A_YJiz5Z9H3_2;
	wire w_dff_A_3ZEmc1Qq4_2;
	wire w_dff_A_GR0woiLp9_2;
	wire w_dff_A_ziTFnVBC9_2;
	wire w_dff_B_OSTqnc9o9_3;
	wire w_dff_B_yZBK22iS5_3;
	wire w_dff_B_2fQBAMhR4_3;
	wire w_dff_B_J4G9mpnt1_1;
	wire w_dff_A_8cGpDfv52_1;
	wire w_dff_B_3A6t9QDM7_3;
	wire w_dff_B_Ux9afbeq9_3;
	wire w_dff_B_24faEiGY7_3;
	wire w_dff_B_Pa7mNo931_1;
	wire w_dff_B_E0lqSfHI1_1;
	wire w_dff_B_ITBo9cRh8_1;
	wire w_dff_B_tBpgZeHR6_1;
	wire w_dff_B_IcFqzFcb4_1;
	wire w_dff_A_GugwOcEI1_1;
	wire w_dff_B_ORF3evCs4_1;
	wire w_dff_A_s7wx6l3t2_0;
	wire w_dff_A_Hn3xa1Rf4_0;
	wire w_dff_A_HKxft28O8_0;
	wire w_dff_A_TQ8QPLsV9_0;
	wire w_dff_A_oyhoAt5v5_0;
	wire w_dff_A_XaaQSeDR1_0;
	wire w_dff_A_GbYdWwlj5_0;
	wire w_dff_A_UNfPpoSj7_2;
	wire w_dff_A_xDs9WJzV1_2;
	wire w_dff_A_JMSQkLdp9_2;
	wire w_dff_A_1xwARsnp4_2;
	wire w_dff_A_n8K1NTCA0_2;
	wire w_dff_A_JmyOfB7B1_2;
	wire w_dff_B_3EdAInlv4_1;
	wire w_dff_B_9kC6cd7E5_1;
	wire w_dff_B_jHdHPdUh9_0;
	wire w_dff_A_oZ09gIbv8_0;
	wire w_dff_B_PHRg72GV4_0;
	wire w_dff_A_f2O2TfQE2_1;
	wire w_dff_A_ROk1wMdd7_1;
	wire w_dff_A_O1iMba9j5_1;
	wire w_dff_A_N5L1lzpW5_1;
	wire w_dff_A_QjXIX3JX3_1;
	wire w_dff_A_q4424rMo6_1;
	wire w_dff_A_qQHdypN76_1;
	wire w_dff_A_p8ELpzs83_1;
	wire w_dff_A_NPPMvooM8_1;
	wire w_dff_A_zsDmacJB5_1;
	wire w_dff_A_7SMRNitG2_1;
	wire w_dff_A_aBqoN1gC4_1;
	wire w_dff_A_rhnNNtjf9_2;
	wire w_dff_A_TuA7yQBL6_2;
	wire w_dff_A_U4G2hbYB4_2;
	wire w_dff_A_VZajrdVB7_2;
	wire w_dff_A_FNF8GtI49_0;
	wire w_dff_A_cda3Ibtk0_0;
	wire w_dff_A_ZoqZzlTJ5_0;
	wire w_dff_A_PY053j2E3_0;
	wire w_dff_A_NWjxawI12_0;
	wire w_dff_B_aw7lozyC2_0;
	wire w_dff_B_n68jINf37_0;
	wire w_dff_A_CsKIKhNk8_2;
	wire w_dff_A_6ClywbqX8_2;
	wire w_dff_A_yv9RxOo11_2;
	wire w_dff_A_oCgTu8PU1_2;
	wire w_dff_A_om3QB3IG7_2;
	wire w_dff_A_kIFH2Ysa1_2;
	wire w_dff_A_b1lHgAcI0_2;
	wire w_dff_A_OKjBty4r9_2;
	wire w_dff_A_RsAMSWpq3_2;
	wire w_dff_B_mBIfwTu57_0;
	wire w_dff_B_HxCQNKHB7_0;
	wire w_dff_B_Qes4Prln1_0;
	wire w_dff_B_9gG2pNCA3_0;
	wire w_dff_B_jlxAK9nM9_0;
	wire w_dff_B_9cMgXHwX2_0;
	wire w_dff_B_t2YV5ulg4_0;
	wire w_dff_B_RF4hpguR9_1;
	wire w_dff_B_A3jLiNuo4_1;
	wire w_dff_B_BNt8wNsu8_1;
	wire w_dff_B_tyQKaLlA7_0;
	wire w_dff_B_KdZ70WhS7_0;
	wire w_dff_B_7ESZrZng0_0;
	wire w_dff_A_8psWY8rS6_1;
	wire w_dff_A_YyiYAuhi0_1;
	wire w_dff_A_XMNBXna95_2;
	wire w_dff_A_6uaoxXlx0_2;
	wire w_dff_A_DSLseczh2_2;
	wire w_dff_A_FadPCto76_2;
	wire w_dff_A_4iOF6mXk2_2;
	wire w_dff_A_Sd7ZNSfY2_2;
	wire w_dff_A_CVp4pTp89_2;
	wire w_dff_A_8fctjVtq2_2;
	wire w_dff_B_6MfxNJ1F1_0;
	wire w_dff_B_Q4nvGl6c1_0;
	wire w_dff_A_K5y6vMox0_1;
	wire w_dff_B_3f5k93LL3_0;
	wire w_dff_A_iXiu8ig33_0;
	wire w_dff_A_40PAzvkt0_0;
	wire w_dff_A_rNztm4fG1_1;
	wire w_dff_A_De6k9eKv4_1;
	wire w_dff_A_5mpRZrMx0_1;
	wire w_dff_A_PfoVU7vB4_2;
	wire w_dff_A_rGcJMBIj6_2;
	wire w_dff_A_WPNxCxhU7_0;
	wire w_dff_A_wBv5RdHQ9_0;
	wire w_dff_A_OHByhVgl2_1;
	wire w_dff_A_8DaOgCE19_1;
	wire w_dff_A_Sn8UzVX90_2;
	wire w_dff_A_AEw2G3VR6_2;
	wire w_dff_A_cOKP08oN6_2;
	wire w_dff_A_e6d3Dqpr7_1;
	wire w_dff_A_fJHbRvmw7_1;
	wire w_dff_A_gH7AkekS8_1;
	wire w_dff_A_eiDE24Oq2_1;
	wire w_dff_B_LDgdsH4j0_0;
	wire w_dff_B_mJyPI1ZB7_0;
	wire w_dff_B_K0aRBr5x9_1;
	wire w_dff_B_TGNX02BM7_1;
	wire w_dff_B_XsJZ1J8F9_1;
	wire w_dff_B_gNEDBGez0_1;
	wire w_dff_B_USA1XYU61_0;
	wire w_dff_A_JHKb9dFG7_1;
	wire w_dff_A_aPMWqlyr2_1;
	wire w_dff_A_AszVSaBX6_1;
	wire w_dff_A_qFW8mvb81_1;
	wire w_dff_A_tsGL62uo6_1;
	wire w_dff_A_yoJMUpJN0_2;
	wire w_dff_A_x9FcaIIF3_2;
	wire w_dff_B_ITkbkyJf1_1;
	wire w_dff_B_uJOhXaQ34_1;
	wire w_dff_A_XgHMaMKJ0_1;
	wire w_dff_B_PERCOOkK4_1;
	wire w_dff_B_h4qqhYoZ3_1;
	wire w_dff_B_O3Odp1da0_0;
	wire w_dff_B_v9iNmF707_0;
	wire w_dff_B_RwoL5VWu8_1;
	wire w_dff_A_sDiaw4jP0_1;
	wire w_dff_A_xY4JYrGU6_0;
	wire w_dff_A_fhwY2GGF7_1;
	wire w_dff_B_lOVN20O51_3;
	wire w_dff_B_rVxBzmCT4_3;
	wire w_dff_A_CxId2X4p1_0;
	wire w_dff_A_YeNUUbk43_0;
	wire w_dff_A_Yq1g9EbF9_0;
	wire w_dff_A_QovUWjK44_1;
	wire w_dff_A_PCgw152I9_1;
	wire w_dff_A_W5vhrWtU2_1;
	wire w_dff_A_xR7b1os08_1;
	wire w_dff_A_PcNxiZVX6_0;
	wire w_dff_A_IIsPcozW7_1;
	wire w_dff_A_O0UPS0rg6_1;
	wire w_dff_A_u3LkBAgE3_2;
	wire w_dff_B_UF5t5H872_1;
	wire w_dff_B_8Vywqy5C4_1;
	wire w_dff_A_C1qcDK9h2_1;
	wire w_dff_A_vSeCGvWH5_1;
	wire w_dff_A_xOXKEPir9_1;
	wire w_dff_A_A5yn995E5_2;
	wire w_dff_A_5zADzc499_2;
	wire w_dff_A_8LkxneID7_2;
	wire w_dff_A_V27RGjLX5_2;
	wire w_dff_A_jZ8bFWoo9_1;
	wire w_dff_A_YnKQKoVh5_1;
	wire w_dff_A_MzxxoxCA9_1;
	wire w_dff_A_DVdKI9wv2_1;
	wire w_dff_A_yuAZQRgU4_1;
	wire w_dff_A_ef7BMETH9_0;
	wire w_dff_A_tuXdhDwY1_0;
	wire w_dff_A_Ipm7vSBl0_2;
	wire w_dff_A_bAIyhmRv0_2;
	wire w_dff_A_JvW1s6wj8_0;
	wire w_dff_A_U5NGfB3C5_0;
	wire w_dff_A_4jPOWda36_2;
	wire w_dff_A_VXiDgnTl0_2;
	wire w_dff_A_mQ5PH6K54_2;
	wire w_dff_A_BZKHOI4D0_1;
	wire w_dff_A_w0RmUAOp6_1;
	wire w_dff_A_qcIAzvu09_1;
	wire w_dff_A_uhmDajlO9_1;
	wire w_dff_A_dHVanQTw5_2;
	wire w_dff_A_Nyew7vER2_2;
	wire w_dff_A_wqkhJfN54_2;
	wire w_dff_A_Zi7TV5ts4_2;
	wire w_dff_A_hwu55APx7_2;
	wire w_dff_A_K1yCmZ129_2;
	wire w_dff_A_FmQ1WqRS3_2;
	wire w_dff_A_nkb3mWIg6_2;
	wire w_dff_A_XOHknlG88_2;
	wire w_dff_A_Lq4xPcLF3_1;
	wire w_dff_A_GsUCtSeh1_1;
	wire w_dff_A_rV0vbByL7_0;
	wire w_dff_A_mUoU2YLO5_1;
	wire w_dff_A_wN72twRj6_1;
	wire w_dff_B_STIrPms96_0;
	wire w_dff_A_psZ4pvPn6_0;
	wire w_dff_A_mGCpcx5X1_0;
	wire w_dff_A_xy45DvJ30_1;
	wire w_dff_A_D6gbvKTe2_1;
	wire w_dff_A_dcoKiQBF6_1;
	wire w_dff_A_BlOSIGtz5_1;
	wire w_dff_A_UDYrwmQr2_1;
	wire w_dff_B_vcISusnL7_0;
	wire w_dff_B_rBoAC2sS8_0;
	wire w_dff_A_WW3mbcMB1_1;
	wire w_dff_A_fFhQYuH08_1;
	wire w_dff_A_I6SmfvYh6_1;
	wire w_dff_A_I6R4qOpr9_1;
	wire w_dff_A_CwkCNF3L1_1;
	wire w_dff_A_IvJ5Yk489_0;
	wire w_dff_B_OrLSHVmi8_1;
	wire w_dff_B_azq4YLDP6_1;
	wire w_dff_B_acPEU2UT6_1;
	wire w_dff_A_8l4yuvmS0_1;
	wire w_dff_A_BhmWJ5Xk8_2;
	wire w_dff_B_L6k4xnL21_1;
	wire w_dff_B_RxrF3lmL5_1;
	wire w_dff_A_CJmQAE0W4_2;
	wire w_dff_A_uBod4A164_1;
	wire w_dff_A_6qfkpFnA6_2;
	wire w_dff_A_VOUHRpC53_0;
	wire w_dff_A_iYvogae46_0;
	wire w_dff_A_gaaqrNnu9_0;
	wire w_dff_A_myzdZv9H0_1;
	wire w_dff_A_CZyKlEfI8_1;
	wire w_dff_B_vGb3QaKr3_0;
	wire w_dff_A_UH2mw9IG9_1;
	wire w_dff_A_v6Kexx641_1;
	wire w_dff_B_aDt2lZxg4_1;
	wire w_dff_A_lGjIW0tb1_2;
	wire w_dff_A_ZVkHsFxW5_2;
	wire w_dff_A_Wn6G64x50_1;
	wire w_dff_A_P5CCnnsY7_1;
	wire w_dff_A_vIN32VZI0_1;
	wire w_dff_A_UjcH846S9_1;
	wire w_dff_A_ugurzdDE3_2;
	wire w_dff_A_AOrGp42Y8_2;
	wire w_dff_A_4IRxXou16_0;
	wire w_dff_A_4u1g0nRA4_0;
	wire w_dff_A_c0kaHqI69_2;
	wire w_dff_A_sABhtlWN3_2;
	wire w_dff_A_ugfSWE8Z0_1;
	wire w_dff_A_S3P8vT1S3_0;
	wire w_dff_A_hyYF8zgZ9_0;
	wire w_dff_A_PoKWS1oL5_0;
	wire w_dff_A_4f98VY5J0_0;
	wire w_dff_A_r52exDBL5_0;
	wire w_dff_A_UL17uMyz6_1;
	wire w_dff_A_lCjPuVzC0_1;
	wire w_dff_A_zQqKriJB3_0;
	wire w_dff_A_KOZBvQqa7_0;
	wire w_dff_A_2fVsdO4y2_0;
	wire w_dff_A_DBtIjgyf7_0;
	wire w_dff_A_T04A5Jm83_0;
	wire w_dff_A_09glOBoH0_0;
	wire w_dff_A_EW6FVQyj1_0;
	wire w_dff_A_pI5UWDYu8_0;
	wire w_dff_A_K3q8J32N3_1;
	wire w_dff_A_rkfMiR059_1;
	wire w_dff_A_Gm4CyLtF8_1;
	wire w_dff_A_V6jSsjcw7_1;
	wire w_dff_B_zLrZuBmg2_0;
	wire w_dff_B_0yChTZMT8_1;
	wire w_dff_A_WruRIkvC8_0;
	wire w_dff_A_Maqp9vwT3_1;
	wire w_dff_A_7UT1Tdcn2_1;
	wire w_dff_A_IAiOz3ZI6_2;
	wire w_dff_A_FZAOHU4A3_2;
	wire w_dff_A_HKxjezPj9_1;
	wire w_dff_A_0C1uqOXc6_0;
	wire w_dff_A_ojfbe8eC4_2;
	wire w_dff_A_aIBsKakw8_2;
	wire w_dff_A_Q4Evzbr60_0;
	wire w_dff_A_ZNRnTKv70_0;
	wire w_dff_A_s9hBFqu00_0;
	wire w_dff_A_HmUdrO5U0_0;
	wire w_dff_A_cu6nqP592_1;
	wire w_dff_A_jIEF3LPd4_1;
	wire w_dff_A_LFqTsjbc6_0;
	wire w_dff_A_YBop4ogN4_1;
	wire w_dff_A_d4Ac9V5o7_1;
	wire w_dff_A_Mk9d0q7l7_1;
	wire w_dff_A_ptBuZUVv8_2;
	wire w_dff_A_bzBoME3G6_2;
	wire w_dff_A_Q2RwdHnB6_1;
	wire w_dff_A_y6QJ2NYk0_1;
	wire w_dff_A_LKGd0RP57_0;
	wire w_dff_A_5pvZ8Iej6_1;
	wire w_dff_A_jJRwyNRU9_1;
	wire w_dff_A_VMpsqkN26_0;
	wire w_dff_A_MgaHJqQP3_0;
	wire w_dff_A_WGcIau8i4_0;
	wire w_dff_A_kslexxj42_1;
	wire w_dff_A_vm0PmMfd2_1;
	wire w_dff_A_lUeRqMzZ6_0;
	wire w_dff_A_Lyne1nuA5_1;
	wire w_dff_A_xBgHXuCO4_1;
	wire w_dff_A_Yh9u04z25_2;
	wire w_dff_A_a4qbyPcr0_2;
	wire w_dff_A_ONNWueaN8_1;
	wire w_dff_A_JHn4h5fV4_2;
	wire w_dff_A_JoHpLu1U0_2;
	wire w_dff_A_xbHy7meL8_0;
	wire w_dff_A_SqJOrxYE3_0;
	wire w_dff_A_h97w8Uuz8_0;
	wire w_dff_A_q04uKjDl0_0;
	wire w_dff_A_XbByAM9Z5_1;
	wire w_dff_A_VK0Jemwn8_1;
	wire w_dff_A_lk2PBJq41_0;
	wire w_dff_B_Fsh1G4pF3_0;
	wire w_dff_A_4EkeUj953_2;
	wire w_dff_B_7izUGPf87_0;
	wire w_dff_B_7kdH1aLg2_0;
	wire w_dff_B_YHsPo9ub3_0;
	wire w_dff_A_pyvMT0dW7_0;
	wire w_dff_A_ubAFFJDR1_0;
	wire w_dff_A_eNjzWxfS2_1;
	wire w_dff_A_0YNUmbHB5_1;
	wire w_dff_A_BeM6e52w4_2;
	wire w_dff_A_tA6eYaIu4_2;
	wire w_dff_B_FCYgFZDb8_3;
	wire w_dff_B_Dgf2wMUK4_3;
	wire w_dff_B_0mSZYAmZ8_3;
	wire w_dff_B_leZnMZJz3_3;
	wire w_dff_B_fj0fuCCv9_3;
	wire w_dff_A_C6mqboJQ1_1;
	wire w_dff_A_yg7TGh7s4_1;
	wire w_dff_A_dMFM4oPT9_1;
	wire w_dff_A_0v9d9oYZ3_1;
	wire w_dff_A_Nbk5Aqs47_1;
	wire w_dff_A_fRorsgP65_1;
	wire w_dff_A_b8cO9g9e4_0;
	wire w_dff_A_Gva2bMP27_1;
	wire w_dff_A_MeHRTeA34_1;
	wire w_dff_A_tCXveOjQ6_2;
	wire w_dff_A_pbCCveUn4_1;
	wire w_dff_A_UM007gqd4_1;
	wire w_dff_A_1H4g7aOH3_1;
	wire w_dff_A_sSWuGHby9_1;
	wire w_dff_A_KXepKQry7_1;
	wire w_dff_A_Bc6Smvon8_1;
	wire w_dff_B_H5DWbEEY9_1;
	wire w_dff_A_ehyGtSRL7_1;
	wire w_dff_B_l6ynPKtQ1_1;
	wire w_dff_B_vjIuho306_1;
	wire w_dff_A_m0U3yfr82_0;
	wire w_dff_A_t9qhoLV72_2;
	wire w_dff_B_3956jpsI0_0;
	wire w_dff_B_v4umk7t39_1;
	wire w_dff_A_jTypQ46G6_1;
	wire w_dff_A_y5iOTmpa2_0;
	wire w_dff_B_b6QY8yMK0_0;
	wire w_dff_A_wpDTwxvd2_0;
	wire w_dff_A_hlo8UFjr6_1;
	wire w_dff_A_E0X6eWJ73_1;
	wire w_dff_A_BlTCyyYc9_1;
	wire w_dff_A_bViPQEmR9_0;
	wire w_dff_A_JqIje15q7_2;
	wire w_dff_A_4Z7QsvPG7_1;
	wire w_dff_A_9Zcfe4AD1_2;
	wire w_dff_A_XtgaX3F38_0;
	wire w_dff_A_UifMbqcT0_0;
	wire w_dff_A_eQ84Agja2_1;
	wire w_dff_A_GS59ELfG3_1;
	wire w_dff_A_smOwfoRH9_1;
	wire w_dff_A_dZlq84rC4_0;
	wire w_dff_A_ezplO8FG1_0;
	wire w_dff_A_9GkQ8nxk7_1;
	wire w_dff_A_UT5E5WLW6_1;
	wire w_dff_A_zwpxlafl6_0;
	wire w_dff_A_mCUAmSWn7_0;
	wire w_dff_A_kq9R0Hx92_0;
	wire w_dff_A_d9JyWCYQ8_2;
	wire w_dff_B_1o0b1wRq7_3;
	wire w_dff_B_2fIvKTzI6_3;
	wire w_dff_B_n66BveGg3_3;
	wire w_dff_B_dQmmLHRO0_3;
	wire w_dff_B_kMTbtHbg6_3;
	wire w_dff_B_ffUfftvl6_3;
	wire w_dff_A_2TRl5kqn1_0;
	wire w_dff_A_f3ju7Xvn3_0;
	wire w_dff_B_iXyxHpsb3_2;
	wire w_dff_B_mXIarFpT2_2;
	wire w_dff_B_CnME2FJ40_2;
	wire w_dff_B_W7UKalJt1_2;
	wire w_dff_B_7dexFQRr4_1;
	wire w_dff_B_3KsAx5iO0_0;
	wire w_dff_B_hoiOK8je7_0;
	wire w_dff_B_eIU6FKJH2_0;
	wire w_dff_B_H2ok2CHD2_0;
	wire w_dff_B_2uiw1TE68_0;
	wire w_dff_A_Icil9oyk6_0;
	wire w_dff_A_HV5MqwNv4_0;
	wire w_dff_A_wCY4BIU75_0;
	wire w_dff_A_FJXwIsoD3_0;
	wire w_dff_A_B099aipu7_0;
	wire w_dff_A_I9OoPHr58_0;
	wire w_dff_A_3RdTVT158_0;
	wire w_dff_A_0mHxmi5c9_1;
	wire w_dff_A_prntjCou7_1;
	wire w_dff_A_YJ7N1I1O6_1;
	wire w_dff_A_u93sXQNP5_1;
	wire w_dff_A_zIyt1ZDW7_1;
	wire w_dff_A_2tQIXM091_0;
	wire w_dff_A_BXp19r1I9_2;
	wire w_dff_A_Gtl4BAO57_2;
	wire w_dff_A_NKXy33Zt9_2;
	wire w_dff_A_FSrO6w4K0_0;
	wire w_dff_A_bZCkoJDo6_0;
	wire w_dff_A_6VTTiOdz4_0;
	wire w_dff_A_Y0dcH6Gw9_0;
	wire w_dff_A_DcO9EYeb0_0;
	wire w_dff_A_ieJJYPRg7_0;
	wire w_dff_A_VBAT3ybe9_1;
	wire w_dff_A_2Ub4ESG99_1;
	wire w_dff_A_6ineyHI54_1;
	wire w_dff_A_zThGJpvx2_2;
	wire w_dff_A_diHCYZvR4_2;
	wire w_dff_A_AfTxsI4D4_2;
	wire w_dff_A_ZqrpNP8R5_1;
	wire w_dff_A_sukh36C02_1;
	wire w_dff_A_uCHG4j7O2_2;
	wire w_dff_A_hrCraXZX3_2;
	wire w_dff_A_D9v8rz468_2;
	wire w_dff_A_pK4nazjv8_2;
	wire w_dff_A_AUfBtQ1c5_0;
	wire w_dff_A_PPGohfHm8_0;
	wire w_dff_A_Ib35Ox4U7_0;
	wire w_dff_A_OFeyg3eT2_0;
	wire w_dff_A_PRuOSv1q6_2;
	wire w_dff_A_pJD95jjG5_1;
	wire w_dff_A_N68nDtWQ1_1;
	wire w_dff_A_FMuI1CcA8_0;
	wire w_dff_B_g2BUHUmX1_1;
	wire w_dff_B_AroFzrwl4_1;
	wire w_dff_B_EOO2UkWM2_1;
	wire w_dff_B_zs0to0HM6_1;
	wire w_dff_A_JrF3vsGJ7_2;
	wire w_dff_A_Gul787wf1_2;
	wire w_dff_A_N1DAoVzM8_2;
	wire w_dff_A_Evudwhde2_2;
	wire w_dff_A_KpwcKUwN2_2;
	wire w_dff_A_gusQRcRR1_2;
	wire w_dff_A_Pgt8R5mk2_2;
	wire w_dff_A_Q82G0qZs0_2;
	wire w_dff_A_xSsMCRBr7_0;
	wire w_dff_A_lW4jTWas2_0;
	wire w_dff_A_3elhcIgK5_0;
	wire w_dff_A_Qz9JojIl6_0;
	wire w_dff_A_FvVptbhJ6_0;
	wire w_dff_A_tvZyrkCr1_0;
	wire w_dff_A_SprqBrJ81_1;
	wire w_dff_A_jlWWod3j4_1;
	wire w_dff_A_4ED3xgM51_1;
	wire w_dff_A_iVZsRrpd7_0;
	wire w_dff_A_2SGy3vXE7_0;
	wire w_dff_A_UfpkqPRw4_1;
	wire w_dff_A_iCkZqIXJ7_1;
	wire w_dff_A_IfmgPiJs5_1;
	wire w_dff_A_66Lb5xL71_0;
	wire w_dff_A_kk3grUL39_1;
	wire w_dff_A_DLOvlq2Y9_1;
	wire w_dff_A_U3yMFeo12_1;
	wire w_dff_A_t101vT8I6_1;
	wire w_dff_A_GYNZU5xm9_0;
	wire w_dff_A_Z5goGDQd7_2;
	wire w_dff_A_ywlBQ1Eu4_2;
	wire w_dff_A_atCkOc2f6_2;
	wire w_dff_A_4T2OBKU75_0;
	wire w_dff_A_uevzUhaB9_1;
	wire w_dff_A_YHrPatvI4_1;
	wire w_dff_A_5FfXtKws4_1;
	wire w_dff_A_Ur4fGXuz7_0;
	wire w_dff_A_tvIXBdGs1_1;
	wire w_dff_A_Om6iWjaW9_1;
	wire w_dff_A_skZTG5Uq4_1;
	wire w_dff_A_l5QVFNa52_1;
	wire w_dff_A_3kGape6e9_2;
	wire w_dff_A_Igq2p78F1_2;
	wire w_dff_A_OVOzVEbJ0_2;
	wire w_dff_A_HR4uFf1G5_1;
	wire w_dff_A_jvgRanVX8_1;
	wire w_dff_A_W5TRT1jw1_1;
	wire w_dff_A_sHAus9Hg6_1;
	wire w_dff_A_6lkBff8a2_1;
	wire w_dff_A_r3xTgCrX5_1;
	wire w_dff_A_cHLg8j5i1_1;
	wire w_dff_A_KxzTbend0_1;
	wire w_dff_A_L1OUvBOX5_1;
	wire w_dff_A_gLdsm9MT0_1;
	wire w_dff_A_vOdaRpIR9_1;
	wire w_dff_A_wVzkdJBF7_1;
	wire w_dff_A_WB1iM4RD7_1;
	wire w_dff_A_HlhaDl444_1;
	wire w_dff_A_bUjDrnwq9_1;
	wire w_dff_A_Uld5ZWv42_1;
	wire w_dff_A_pB17JVLV8_1;
	wire w_dff_A_RYyAyxtK4_1;
	wire w_dff_A_AieAZqdi9_1;
	wire w_dff_A_3UeoD8xh0_1;
	wire w_dff_A_mJel1wGl0_1;
	wire w_dff_A_iTbNsJcu3_1;
	wire w_dff_A_VLgwlKXU5_1;
	wire w_dff_A_sQCRFlbg1_1;
	wire w_dff_A_pilupIAD1_1;
	wire w_dff_A_LlXQbDvJ1_1;
	wire w_dff_A_3QuVspq13_1;
	wire w_dff_A_qabvBadO0_1;
	wire w_dff_A_vBIy6OKn2_1;
	wire w_dff_A_Zq0Bc14H4_1;
	wire w_dff_A_S1Gy7Grj3_2;
	wire w_dff_A_oXYJQoHw7_2;
	wire w_dff_A_PVds1BQh4_2;
	wire w_dff_A_VG8jbie57_2;
	wire w_dff_A_Eibqprn34_2;
	wire w_dff_A_abaKJPaS9_2;
	wire w_dff_A_huDPOu0W6_2;
	wire w_dff_A_n08iQj1A2_2;
	wire w_dff_A_NOo5No7a1_1;
	wire w_dff_A_ja4D9moc2_1;
	wire w_dff_A_4MwNiXOn4_1;
	wire w_dff_B_epnIwufb4_0;
	wire w_dff_B_IPXw9dON6_0;
	wire w_dff_B_zQEgkBVr2_1;
	wire w_dff_B_SI3vpvEF0_1;
	wire w_dff_B_duIrmeBB7_1;
	wire w_dff_B_2WX1sdRp1_1;
	wire w_dff_B_PGB7mGTc7_0;
	wire w_dff_A_wFVyREYN6_0;
	wire w_dff_B_15zbGLLk8_3;
	wire w_dff_B_PFBmPIhI2_3;
	wire w_dff_B_aZT4eAIR2_3;
	wire w_dff_A_FduAQ6k65_1;
	wire w_dff_B_YFWQiIGl2_3;
	wire w_dff_B_b8tum4Cb1_3;
	wire w_dff_B_DleL7hkB5_3;
	wire w_dff_B_Qoi6h4hS8_1;
	wire w_dff_B_MkNT7zZD7_1;
	wire w_dff_B_hpPNEX8y4_1;
	wire w_dff_B_U5SKTSDO0_1;
	wire w_dff_B_s0siIhop1_0;
	wire w_dff_B_Xa6NuVoZ9_0;
	wire w_dff_A_UAHBuC8a9_0;
	wire w_dff_B_ctEQa78R7_2;
	wire w_dff_B_uWuWFUxP0_2;
	wire w_dff_B_3IYLQbVv5_2;
	wire w_dff_B_MdHqP3XU9_1;
	wire w_dff_A_RvwD4hSX8_0;
	wire w_dff_A_HFE3nYvt1_0;
	wire w_dff_A_InUxnsUw6_0;
	wire w_dff_A_7KXAvexG1_0;
	wire w_dff_A_nCtp9fmY5_0;
	wire w_dff_A_imFC1NFv1_0;
	wire w_dff_A_M8PDc24u2_0;
	wire w_dff_A_dfPF7vOD9_1;
	wire w_dff_A_XA49QrCj3_1;
	wire w_dff_A_UGB6UDPz6_1;
	wire w_dff_A_IgwH6UHi3_0;
	wire w_dff_B_nT9B3m7w1_3;
	wire w_dff_B_DuNi19WN8_3;
	wire w_dff_B_76RyYuVJ5_3;
	wire w_dff_B_XZYEa8my8_0;
	wire w_dff_B_ZpGwgD9l5_1;
	wire w_dff_B_WwaOHHlo8_1;
	wire w_dff_A_Rpv7GXwZ4_1;
	wire w_dff_A_gkhyvNus0_1;
	wire w_dff_A_99bYBXMd5_2;
	wire w_dff_A_YbKn54312_2;
	wire w_dff_A_hIy1Evbj3_2;
	wire w_dff_A_Lvr95I756_0;
	wire w_dff_A_myzgEm6o4_0;
	wire w_dff_A_bPu9byLN0_1;
	wire w_dff_A_IatAuJ4D8_1;
	wire w_dff_A_uRXQAEmO4_0;
	wire w_dff_A_TYmLuvgm0_2;
	wire w_dff_A_iPQOF0Vq4_2;
	wire w_dff_A_PLpIwZTf2_2;
	wire w_dff_A_TfYO4oLX8_2;
	wire w_dff_A_BaM0tXbx0_1;
	wire w_dff_A_rwpDjkM27_0;
	wire w_dff_A_u7tOXK7N1_0;
	wire w_dff_A_1053Xzse9_0;
	wire w_dff_A_PSu8SQtN0_1;
	wire w_dff_A_mLeTIMsk2_1;
	wire w_dff_A_JOflgydm7_1;
	wire w_dff_A_lbRvUuZh2_0;
	wire w_dff_A_GjeJFaG75_0;
	wire w_dff_A_JDcLtCSU8_0;
	wire w_dff_A_jcmTerpl0_2;
	wire w_dff_A_ga0eICyE4_2;
	wire w_dff_A_S2EvNYYq9_2;
	wire w_dff_A_a8oYTciW2_2;
	wire w_dff_A_oDEU0Bbw2_2;
	wire w_dff_A_ID44LOwM4_1;
	wire w_dff_B_cx0kmtJb8_1;
	wire w_dff_B_cTi4cvda5_1;
	wire w_dff_A_Ud0i2WQE0_0;
	wire w_dff_A_LySYsfzo0_0;
	wire w_dff_A_uCHVmEAR2_0;
	wire w_dff_A_RRvMJjBr1_1;
	wire w_dff_A_easMpTaD7_1;
	wire w_dff_A_wBMgzwlS3_1;
	wire w_dff_A_OjRpaYTH3_1;
	wire w_dff_A_jPZB0Uh39_0;
	wire w_dff_A_fgpOljVt1_0;
	wire w_dff_A_gTmJHqmw8_0;
	wire w_dff_A_BoUr2vNR5_1;
	wire w_dff_A_7aLUCqxE7_1;
	wire w_dff_A_02gL5xdu7_1;
	wire w_dff_A_FNTuUT801_0;
	wire w_dff_A_HTBDeNDf9_0;
	wire w_dff_A_VJu7bfcK9_0;
	wire w_dff_A_rJbWsbZI0_0;
	wire w_dff_A_dhPSkfWg5_0;
	wire w_dff_A_hvqDGvPG2_0;
	wire w_dff_A_0DNBLfcy6_1;
	wire w_dff_A_roSSWwob9_1;
	wire w_dff_A_Gn1Ngk807_1;
	wire w_dff_A_wRJmGnUW9_1;
	wire w_dff_A_nEejx1Yk7_1;
	wire w_dff_A_eFTL9DI97_1;
	wire w_dff_A_5ZUteJJl5_1;
	wire w_dff_A_OVgrBv1T6_1;
	wire w_dff_A_CtOhJ50s6_1;
	wire w_dff_A_NnTjfPfF4_1;
	wire w_dff_A_Z8NYjraw5_1;
	wire w_dff_A_VaIGOAew9_1;
	wire w_dff_A_cNXzxi6f5_1;
	wire w_dff_A_9LhzQicR2_1;
	wire w_dff_A_JVEiqZj74_1;
	wire w_dff_A_juqI9PiX2_2;
	wire w_dff_A_dv0y0SBw3_2;
	wire w_dff_A_uf482u1O4_2;
	wire w_dff_A_ZGUTahiJ3_2;
	wire w_dff_A_9gTQKhFJ3_2;
	wire w_dff_A_ddD7f9Uq0_2;
	wire w_dff_A_RuwTxlmp4_2;
	wire w_dff_A_7bb0sUTJ1_0;
	wire w_dff_A_50Fg1vgp4_0;
	wire w_dff_A_RnLehcsx9_0;
	wire w_dff_A_i9CGDgPG3_2;
	wire w_dff_A_MlJChBlm4_2;
	wire w_dff_A_6R5e6Vpw8_2;
	wire w_dff_A_H00ab9SS9_1;
	wire w_dff_A_TlHlMIDS6_1;
	wire w_dff_A_WHNRDtKO3_0;
	wire w_dff_A_QzjSqOyr6_0;
	wire w_dff_A_iZdiPAK29_0;
	wire w_dff_A_i9Y28Gpo5_0;
	wire w_dff_A_eH5pr1Dt4_0;
	wire w_dff_A_KAokJYo86_0;
	wire w_dff_A_awdv05eE1_1;
	wire w_dff_B_HSexzlMl6_0;
	wire w_dff_A_f6htjZ0h2_0;
	wire w_dff_A_ctYTbV0I7_0;
	wire w_dff_A_lb8DHTMQ0_0;
	wire w_dff_A_2w6f3LV65_1;
	wire w_dff_A_8vQCB9x34_1;
	wire w_dff_A_sCFfnYDW2_1;
	wire w_dff_A_1cN0h2PT2_0;
	wire w_dff_A_gV5tDO9v0_0;
	wire w_dff_A_tP0ttjuI6_0;
	wire w_dff_A_WuJdh9tN4_0;
	wire w_dff_A_2SLOiQmU2_2;
	wire w_dff_A_JTPDVDkf9_2;
	wire w_dff_A_5qPkdKiB1_2;
	wire w_dff_A_oMVEQn4J3_2;
	wire w_dff_A_naVGPcSL9_2;
	wire w_dff_A_jcyD8gAL9_2;
	wire w_dff_A_tyIazhTB1_2;
	wire w_dff_A_qJJ0psJq6_2;
	wire w_dff_A_LNnhatrx2_0;
	wire w_dff_A_EdOHaFaB2_0;
	wire w_dff_A_HegGS2qX4_1;
	wire w_dff_A_aJvojiDY3_1;
	wire w_dff_A_NSxwuF543_1;
	wire w_dff_A_EgUzCAux4_1;
	wire w_dff_A_UZiJZi3v3_1;
	wire w_dff_A_yLXqfWQo9_1;
	wire w_dff_A_qdkzIen67_1;
	wire w_dff_A_kt9eReKY6_2;
	wire w_dff_A_U5zeaEBP4_0;
	wire w_dff_A_mj3y81XF0_0;
	wire w_dff_A_CirbFGOI2_2;
	wire w_dff_A_G1XrAQAe4_2;
	wire w_dff_A_kwMSiL5q6_2;
	wire w_dff_A_VbPXRntC0_2;
	wire w_dff_A_QiMpmbzV4_2;
	wire w_dff_A_ggKQXFRs6_2;
	wire w_dff_A_wOdYPzuO0_2;
	wire w_dff_A_exnGLAXE9_2;
	wire w_dff_A_Za5J4EeW1_2;
	wire w_dff_A_uAnlLjrn6_0;
	wire w_dff_A_uhWG3V3B0_0;
	wire w_dff_A_bKjz2g4f0_0;
	wire w_dff_A_P9BlaCSh4_0;
	wire w_dff_A_SdTEQVUl4_0;
	wire w_dff_A_EuxU2Int0_0;
	wire w_dff_A_tmBL4v1l1_0;
	wire w_dff_A_SZgxCPfN6_0;
	wire w_dff_A_2QJJym2f7_0;
	wire w_dff_A_AiEo29PQ1_0;
	wire w_dff_A_Gqltzonz4_0;
	wire w_dff_A_6RJezA6N7_0;
	wire w_dff_A_cLTLoYju5_0;
	wire w_dff_A_xbB1niDx1_2;
	wire w_dff_A_HzjUXLGv1_2;
	wire w_dff_A_uX9FTeu49_2;
	wire w_dff_A_xm2zcuXS4_2;
	wire w_dff_A_z9eqSGSK2_2;
	wire w_dff_A_6U9VqsfF3_2;
	wire w_dff_A_sH8FbVQ41_2;
	wire w_dff_A_ejUtGVit9_2;
	wire w_dff_A_hh3UPOJj3_2;
	wire w_dff_A_M3oKymkX0_2;
	wire w_dff_A_pAH16aaE0_0;
	wire w_dff_A_EhRKcNdn1_0;
	wire w_dff_A_kbRTm1KI5_0;
	wire w_dff_A_3F6v94TU0_0;
	wire w_dff_A_jiZw6dXz8_0;
	wire w_dff_A_gyGu27sC8_0;
	wire w_dff_A_HzuVDqZY0_0;
	wire w_dff_A_5ahwCGFI4_0;
	wire w_dff_A_pNIealtt9_0;
	wire w_dff_A_gUS2zuK58_0;
	wire w_dff_A_FigNKfxo7_1;
	wire w_dff_A_260bEBTC6_1;
	wire w_dff_A_VEn8q4z92_1;
	wire w_dff_A_msprWaCP2_1;
	wire w_dff_A_zdJ6DOrn3_1;
	wire w_dff_A_2mkDxWwO8_1;
	wire w_dff_A_XVHiTYCN8_1;
	wire w_dff_A_Gr4gVzGG9_1;
	wire w_dff_A_pRUa8Ttq1_1;
	wire w_dff_A_zJ3ZWgMV1_0;
	wire w_dff_A_4yptJBWd6_0;
	wire w_dff_A_yjrrCu7o5_0;
	wire w_dff_A_ibZVVIeY2_0;
	wire w_dff_A_DuypDAPN2_0;
	wire w_dff_A_2kPYGMWC2_0;
	wire w_dff_A_35poXltV8_0;
	wire w_dff_A_TwCJsRjF2_0;
	wire w_dff_A_SgxLCfYC5_0;
	wire w_dff_A_tFbVVaAs8_0;
	wire w_dff_A_oUZrYATW0_0;
	wire w_dff_A_QFvgbUU20_0;
	wire w_dff_A_8kOfjuPP0_0;
	wire w_dff_A_k7wsKiL36_2;
	wire w_dff_A_xf7JuvVR3_2;
	wire w_dff_A_qemMsgKK9_2;
	wire w_dff_A_HYhoACAY5_2;
	wire w_dff_A_w3mQjxe81_2;
	wire w_dff_A_zCGulpcr7_2;
	wire w_dff_A_0NDY6e3v0_2;
	wire w_dff_A_W0WBHR8e2_2;
	wire w_dff_A_K0Pad6Ns8_2;
	wire w_dff_A_4kzqbnWJ8_2;
	wire w_dff_A_yjipZPyy5_2;
	wire w_dff_A_V5rlJOz46_2;
	wire w_dff_A_I9dstlAO9_0;
	wire w_dff_A_JEtBTcVc0_0;
	wire w_dff_A_xWn1uct69_0;
	wire w_dff_A_uk6JKueg4_0;
	wire w_dff_A_cj41HD791_0;
	wire w_dff_A_RNoxb2dK4_0;
	wire w_dff_B_w3v2F4oM6_1;
	wire w_dff_B_HIhbgpsC2_1;
	wire w_dff_B_mV0nW1Tm9_1;
	wire w_dff_B_60ChBBxI3_1;
	wire w_dff_B_FKThuiyb9_1;
	wire w_dff_B_Od5Gk1gw0_1;
	wire w_dff_B_B3u4cSBY8_1;
	wire w_dff_B_q8k9MOuf7_1;
	wire w_dff_B_KvJ7e3XT4_0;
	wire w_dff_B_0Vssa9tt8_0;
	wire w_dff_B_7xDTL5ru8_0;
	wire w_dff_B_jvbrpiFg4_0;
	wire w_dff_A_m7ctGy0p4_0;
	wire w_dff_A_QGRxRHqV0_0;
	wire w_dff_A_NClwg5zS3_0;
	wire w_dff_A_28EEJ0Sn8_0;
	wire w_dff_A_3rZZEYLc6_0;
	wire w_dff_A_MEGH1NvO4_0;
	wire w_dff_A_uCmTs7TH7_0;
	wire w_dff_A_6TImLwIf6_0;
	wire w_dff_A_kYHBqgOM8_0;
	wire w_dff_A_VWP2JInt9_0;
	wire w_dff_A_H10i0gnZ4_0;
	wire w_dff_A_UdIxKefW1_2;
	wire w_dff_A_RFYth3pu9_2;
	wire w_dff_A_O7ydR7cm8_2;
	wire w_dff_A_OV09zMKu6_2;
	wire w_dff_A_0HMKhCxd2_2;
	wire w_dff_A_393srodo3_2;
	wire w_dff_A_LTo0MXWQ5_2;
	wire w_dff_A_BovatdL55_2;
	wire w_dff_A_icapLlXC4_2;
	wire w_dff_A_hqzJ7BUz0_2;
	wire w_dff_A_zyQLVVjd6_1;
	wire w_dff_A_Oye7c9t85_1;
	wire w_dff_A_AaWsLxke0_1;
	wire w_dff_A_cByZCHFb3_2;
	wire w_dff_A_MzwhkeoN1_2;
	wire w_dff_A_VwmtA1gA7_1;
	wire w_dff_A_Z2XBsqBC9_1;
	wire w_dff_A_AfCrQjjM0_1;
	wire w_dff_A_PuTXQgIf1_1;
	wire w_dff_A_az5jMjMD1_1;
	wire w_dff_A_q0CypoSz6_2;
	wire w_dff_A_QXZO0qHl4_2;
	wire w_dff_A_IHj1ibR70_2;
	wire w_dff_A_JJmQXtTo5_2;
	wire w_dff_A_00kALzpj4_2;
	wire w_dff_A_lJ5nagS34_0;
	wire w_dff_A_fFX9Wa6W5_2;
	wire w_dff_A_raF79JIE4_2;
	wire w_dff_A_5xFSuWWJ2_1;
	wire w_dff_A_VH4fbc1h7_1;
	wire w_dff_A_mLMEhh1X3_1;
	wire w_dff_A_aA2Efb6n2_1;
	wire w_dff_A_PyGxFW0l7_2;
	wire w_dff_B_GES3CfPU6_1;
	wire w_dff_B_tISGEVh33_1;
	wire w_dff_A_3jLZoVp15_1;
	wire w_dff_A_ZmYTtGjP7_2;
	wire w_dff_A_hxtQ4qkq4_2;
	wire w_dff_A_eXXOSfVr4_0;
	wire w_dff_A_pg2YfUI82_0;
	wire w_dff_A_gKdiZiIb8_0;
	wire w_dff_A_25PEjoF99_0;
	wire w_dff_A_e7aAggJJ6_0;
	wire w_dff_A_oUdYKSkV9_0;
	wire w_dff_A_AOAazSbn8_0;
	wire w_dff_A_268u0N709_2;
	wire w_dff_A_KUBNllBB7_2;
	wire w_dff_A_ZC8WDYmo0_2;
	wire w_dff_A_mrfJpwXB4_2;
	wire w_dff_A_WrRtgUhA4_2;
	wire w_dff_A_Xcuel7Tg7_2;
	wire w_dff_A_TufCRslF2_2;
	wire w_dff_A_iPX7Z4Cu9_2;
	wire w_dff_A_VefTAxdH1_2;
	wire w_dff_A_cXO4wwz39_2;
	wire w_dff_A_Ldn2NI1j8_2;
	wire w_dff_A_ttA7cKY37_2;
	wire w_dff_A_jOAji8bc1_2;
	wire w_dff_A_8rxErzIf8_2;
	wire w_dff_A_7TIFVRkI6_2;
	wire w_dff_A_NUfNMVn58_1;
	wire w_dff_A_oAfHk9in3_1;
	wire w_dff_B_2RLYosgE9_1;
	wire w_dff_B_4iA5VZ472_1;
	wire w_dff_A_Uw9rA5Q79_1;
	wire w_dff_A_maUN2Flg6_1;
	wire w_dff_A_gb7dweU23_2;
	wire w_dff_A_PeA8ptfg2_0;
	wire w_dff_A_VNirrpwN2_0;
	wire w_dff_A_50kHApfg2_0;
	wire w_dff_A_o4b01Lh21_0;
	wire w_dff_A_Ji9HKJb18_0;
	wire w_dff_A_oKT7Ez0f7_0;
	wire w_dff_A_xpS69ZrS3_1;
	wire w_dff_A_yJts9i7G6_1;
	wire w_dff_A_2yzE9Y8S6_1;
	wire w_dff_A_eM4pA4l30_1;
	wire w_dff_A_vn0SLuPI6_1;
	wire w_dff_A_FPx0BJSn6_1;
	wire w_dff_A_UFx35RBF0_0;
	wire w_dff_A_uVC9z8PY3_0;
	wire w_dff_A_HS9Rn81n8_0;
	wire w_dff_A_bSnjeapd9_0;
	wire w_dff_A_Gbdxrt8p0_0;
	wire w_dff_A_jzvCaJzW7_0;
	wire w_dff_A_W5jceAN66_0;
	wire w_dff_A_adNHm5Ts5_0;
	wire w_dff_A_VNW6KaN29_1;
	wire w_dff_A_Pncs4or61_1;
	wire w_dff_A_cQgTutSB9_1;
	wire w_dff_A_n8LNq6bN8_1;
	wire w_dff_A_JGeeLpHH8_1;
	wire w_dff_A_6CZSu0Gw2_1;
	wire w_dff_A_zdPn62Q54_1;
	wire w_dff_A_C1uqPPe31_1;
	wire w_dff_A_9CGFR2918_0;
	wire w_dff_A_cB6r0kEd9_0;
	wire w_dff_A_PJ0ANXx23_0;
	wire w_dff_A_d28yZRUN3_0;
	wire w_dff_A_8qmwtbr90_0;
	wire w_dff_A_dJhGqiUZ6_0;
	wire w_dff_A_RyIK6iYs2_0;
	wire w_dff_A_kBLVlvFw4_0;
	wire w_dff_A_SyzkO7SL4_1;
	wire w_dff_B_GcnqWhjj5_0;
	wire w_dff_A_21LTCwyy0_0;
	wire w_dff_A_5Os4Co0L7_0;
	wire w_dff_A_D30XsiAm4_0;
	wire w_dff_A_AYEVyLfQ3_1;
	wire w_dff_B_dI5peQw07_1;
	wire w_dff_B_SJl0iTHM2_1;
	wire w_dff_B_BgZDjfnJ5_1;
	wire w_dff_A_Yay1H0sT4_0;
	wire w_dff_A_XjVZ48HX4_0;
	wire w_dff_A_8O7tS3tU4_1;
	wire w_dff_A_axQXsGFK3_1;
	wire w_dff_A_LseBYIOK8_1;
	wire w_dff_A_DwDyRc4z4_2;
	wire w_dff_A_TGsmLIqQ6_2;
	wire w_dff_A_sAjQKnIV0_0;
	wire w_dff_A_25Ixg5Bz5_0;
	wire w_dff_A_hMpawB0o6_0;
	wire w_dff_A_J7DcwswV9_1;
	wire w_dff_A_VvwDY8HE4_1;
	wire w_dff_A_Z1eKN7YO8_1;
	wire w_dff_A_tA4WwVps9_0;
	wire w_dff_A_MY4gmzcB6_0;
	wire w_dff_A_5em3aR5A7_0;
	wire w_dff_A_Yu7uDWyd5_2;
	wire w_dff_A_jhzE4bo43_2;
	wire w_dff_A_K6oeFYj22_2;
	wire w_dff_A_qt1GiljN0_2;
	wire w_dff_A_rzrEgui05_2;
	wire w_dff_A_m34ss2Ex2_0;
	wire w_dff_A_2kBUp0gP7_0;
	wire w_dff_A_B212phLv9_0;
	wire w_dff_A_iK7dFzir4_1;
	wire w_dff_A_ahXSG8UL4_1;
	wire w_dff_A_ceBD7C2p2_1;
	wire w_dff_A_re8iwzaB9_1;
	wire w_dff_A_GVkq5jlA9_2;
	wire w_dff_A_qhl06zxv1_2;
	wire w_dff_A_XKjLqvyA4_1;
	wire w_dff_A_NwQFKoZl5_1;
	wire w_dff_A_bW7EyHf57_2;
	wire w_dff_A_dZmAmqcr4_2;
	wire w_dff_A_MW926Uyt6_1;
	wire w_dff_A_a7OroNKR0_1;
	wire w_dff_A_4NqUh69t6_2;
	wire w_dff_A_rPcvYyJw0_2;
	wire w_dff_A_YJlh3oE04_2;
	wire w_dff_B_j1gpmBTM4_3;
	wire w_dff_A_XTFGpIVr3_1;
	wire w_dff_A_yD4Oi5hU0_0;
	wire w_dff_A_u6jQZWCN8_0;
	wire w_dff_A_NSZ2h9dl9_2;
	wire w_dff_A_03ahk3n16_2;
	wire w_dff_A_GSO5PdCL6_2;
	wire w_dff_A_kNaDVNSq3_1;
	wire w_dff_A_gIp1idMr6_1;
	wire w_dff_A_jjyOFsE86_0;
	wire w_dff_A_NeFbVxgv6_0;
	wire w_dff_A_MncSweYv9_0;
	wire w_dff_A_gw5ysKeH9_0;
	wire w_dff_A_pLAuYhxD6_0;
	wire w_dff_A_xCWnU4zI3_0;
	wire w_dff_A_duVIurAX0_0;
	wire w_dff_A_H7Vs399g6_0;
	wire w_dff_A_8yMCUGnd6_0;
	wire w_dff_A_ei1SxWmQ4_0;
	wire w_dff_A_XdMqc9jc1_0;
	wire w_dff_A_fqjEorEV0_0;
	wire w_dff_A_4moNnSnd2_0;
	wire w_dff_A_p9d7fzAb5_0;
	wire w_dff_A_DdA5je7k2_0;
	wire w_dff_A_LwCLSk4Q9_0;
	wire w_dff_A_F2uvRqSV5_0;
	wire w_dff_A_RfddQYn10_0;
	wire w_dff_A_Ehupaxh00_1;
	wire w_dff_A_XM8BCtkG6_1;
	wire w_dff_A_BVNBrHJ22_1;
	wire w_dff_A_SFIRQzNx1_1;
	wire w_dff_A_wP7iAD9G9_1;
	wire w_dff_A_9MtHASw25_1;
	wire w_dff_A_OEB2aHrV7_1;
	wire w_dff_A_WrA9bOyU1_1;
	wire w_dff_A_53LigxUI3_1;
	wire w_dff_A_GBIGJCYs5_0;
	wire w_dff_A_QgG4Hyin7_1;
	wire w_dff_A_lQQRhe7H8_1;
	wire w_dff_A_yt34euw66_1;
	wire w_dff_A_ON8lIAsy5_1;
	wire w_dff_A_iyrgdOn12_1;
	wire w_dff_A_Zd6KN2l20_1;
	wire w_dff_A_Gi5qJDve0_1;
	wire w_dff_A_N0M2Dwtu1_1;
	wire w_dff_A_agZidya10_1;
	wire w_dff_B_izbAE8qO7_0;
	wire w_dff_B_M2hcu2Iu9_0;
	wire w_dff_A_wyilZyJB0_0;
	wire w_dff_A_qgWVCfvQ1_0;
	wire w_dff_A_awxo882Y8_1;
	wire w_dff_A_AzWh0D143_1;
	wire w_dff_A_TB5hfQ0o8_1;
	wire w_dff_A_6gcDyPwH1_2;
	wire w_dff_A_p1Lv5tZs8_2;
	wire w_dff_B_ZZIFyYAI8_1;
	wire w_dff_B_FzHTR9pu7_1;
	wire w_dff_B_QKp3wjYK2_1;
	wire w_dff_A_sDaQeqU74_0;
	wire w_dff_A_WKeEDn6S5_1;
	wire w_dff_A_CueYVveM3_1;
	wire w_dff_A_l8TPzBcC4_1;
	wire w_dff_A_Yg7is76d4_2;
	wire w_dff_A_xewqMdmD6_2;
	wire w_dff_A_6yYBYou13_2;
	wire w_dff_A_jbusTZln6_1;
	wire w_dff_A_0EFK6krm0_1;
	wire w_dff_A_ytpqUgnf0_1;
	wire w_dff_A_p63nj3rN5_2;
	wire w_dff_A_wGwwfJCx9_2;
	wire w_dff_A_hPOLBwJu3_2;
	wire w_dff_A_dZAaiECU3_2;
	wire w_dff_A_Xo8Car738_2;
	wire w_dff_A_tJ7Qxpoe3_2;
	wire w_dff_A_y8uCNX1z9_2;
	wire w_dff_A_9ngiHv6q8_0;
	wire w_dff_A_oJeBx24G4_0;
	wire w_dff_A_UWfbyl1h1_2;
	wire w_dff_A_bxpFVpxw1_0;
	wire w_dff_A_DcWhLFiX8_0;
	wire w_dff_A_UMyuYaC41_0;
	wire w_dff_A_VPcXu3Td2_1;
	wire w_dff_A_0daeuNOR1_1;
	wire w_dff_A_OcKfnYpe3_1;
	wire w_dff_A_NqqpT5bS4_0;
	wire w_dff_A_DXX6RVdY6_0;
	wire w_dff_A_G7tY3cCa7_0;
	wire w_dff_A_raukKi4E5_1;
	wire w_dff_A_W7JmUWlk9_1;
	wire w_dff_A_IrXp32UJ4_1;
	wire w_dff_A_lypYdccR6_0;
	wire w_dff_A_QoYS69xf0_1;
	wire w_dff_A_rMTa615l0_2;
	wire w_dff_A_J6xfLXCV2_2;
	wire w_dff_A_rB8oE75a0_0;
	wire w_dff_A_rrN7MSkv5_0;
	wire w_dff_A_aCfmhJLD5_0;
	wire w_dff_B_myevPPDS9_0;
	wire w_dff_B_TWpw5Lkn9_0;
	wire w_dff_A_1QcmdyLC6_0;
	wire w_dff_A_H7EoIeNt4_0;
	wire w_dff_A_4G19A59n2_1;
	wire w_dff_A_6UMkh2iw9_2;
	wire w_dff_A_JUyi6zAp5_0;
	wire w_dff_A_7hmPxE388_0;
	wire w_dff_A_Fe2KaN991_0;
	wire w_dff_A_4m3fVzqZ7_0;
	wire w_dff_A_Xf56kWhH1_2;
	wire w_dff_A_TYwDA2GO3_0;
	wire w_dff_A_a2pL4i4R6_0;
	wire w_dff_A_DU8SRIU89_1;
	wire w_dff_A_XtbjMlao6_0;
	wire w_dff_A_fBrIb4Yj7_0;
	wire w_dff_A_t1IPvC8r1_0;
	wire w_dff_A_ksJxD0uI3_0;
	wire w_dff_A_Y9rTJxB16_0;
	wire w_dff_A_cIXMQj1C0_0;
	wire w_dff_A_VKaiihHm3_1;
	wire w_dff_A_AhkhnfD37_2;
	wire w_dff_A_FPq6sE740_2;
	wire w_dff_A_7FnPaeON8_2;
	wire w_dff_A_1mvVggJS4_1;
	wire w_dff_A_wYohYmHl8_1;
	wire w_dff_A_6Jnib6tG3_1;
	wire w_dff_A_v6Tm0TTV7_2;
	wire w_dff_A_OWUQhYUJ5_2;
	wire w_dff_A_7SiU0GIE8_2;
	wire w_dff_A_92WyQHFf7_0;
	wire w_dff_A_2LB4S6lL1_2;
	wire w_dff_B_KJmYe58O5_3;
	wire w_dff_B_ni0jTr7x7_3;
	wire w_dff_B_6bk3x7n79_3;
	wire w_dff_B_rHPmGMoo8_3;
	wire w_dff_B_90HfVKk17_3;
	wire w_dff_B_5gC5FILO3_3;
	wire w_dff_B_qbxsD1Wv8_3;
	wire w_dff_B_MahJQJth5_3;
	wire w_dff_B_3lrWq1ZZ2_3;
	wire w_dff_B_9VXUoVH00_3;
	wire w_dff_B_D5Bx6L4k1_3;
	wire w_dff_B_XISZZfl35_3;
	wire w_dff_B_LllyakdK2_3;
	wire w_dff_A_EIouoLnc5_0;
	wire w_dff_A_QGN3FYtA1_0;
	wire w_dff_A_VPZDvZ3B7_0;
	wire w_dff_A_tOSKmY9K7_0;
	wire w_dff_A_tYyIqU8I4_0;
	wire w_dff_A_PednxCB11_0;
	wire w_dff_A_yc5yqWwW4_0;
	wire w_dff_A_nMsuSsbP8_0;
	wire w_dff_A_Rnhv3WZw1_0;
	wire w_dff_A_uHCxWV2a9_0;
	wire w_dff_A_pe4VyM901_0;
	wire w_dff_A_ax2aeJKe0_0;
	wire w_dff_A_riJUsCaV4_2;
	wire w_dff_A_NtHf2mZN3_2;
	wire w_dff_A_8c6wB8ym4_2;
	wire w_dff_A_fOXKGzIH2_2;
	wire w_dff_A_ZWk61n8A7_2;
	wire w_dff_A_NgFE8Z6K9_2;
	wire w_dff_A_lWijELjg8_2;
	wire w_dff_A_sucSOSwM4_2;
	wire w_dff_A_gidrEGX38_2;
	wire w_dff_A_2eUFjgy66_2;
	wire w_dff_A_OF6GhCY34_2;
	wire w_dff_A_LJbc8UgO7_1;
	wire w_dff_A_1ETxCsuV3_1;
	wire w_dff_A_L1rxmO587_1;
	wire w_dff_A_dRxpiVZy0_1;
	wire w_dff_A_X7aHFhnq1_1;
	wire w_dff_A_8v5wyk799_1;
	wire w_dff_A_TQSST8xv0_1;
	wire w_dff_A_fp8UZbm02_2;
	wire w_dff_A_qshZv7hQ7_2;
	wire w_dff_A_FcQcbM5U6_2;
	wire w_dff_A_fOMhSwhw7_2;
	wire w_dff_A_pMifdcYw3_2;
	wire w_dff_A_9O5Nxu9W0_0;
	wire w_dff_A_eOOd4Wzs3_0;
	wire w_dff_A_sfT8hdn89_0;
	wire w_dff_A_AelXYhZ19_0;
	wire w_dff_A_s2AiT7Rh9_0;
	wire w_dff_A_8AQttcRs1_0;
	wire w_dff_A_NnUSno4B3_0;
	wire w_dff_A_n64U0nQk4_0;
	wire w_dff_A_OkecXknK2_0;
	wire w_dff_A_TpMP28h14_0;
	wire w_dff_A_MyorrT4o6_0;
	wire w_dff_A_6cth4LiG5_0;
	wire w_dff_A_5zyMBQ4e6_0;
	wire w_dff_A_WPwKHGLe3_0;
	wire w_dff_A_aSvgI4nP6_1;
	wire w_dff_A_tFYi5S421_1;
	wire w_dff_A_C23dacP67_1;
	wire w_dff_A_x3oAx41T3_1;
	wire w_dff_A_DlW4a4Wk7_1;
	wire w_dff_A_r1h7pgr00_1;
	wire w_dff_A_eUW2J06r9_1;
	wire w_dff_A_9Coo9IHi9_1;
	wire w_dff_A_GY1MIUoT5_1;
	wire w_dff_A_VaePAUu87_1;
	wire w_dff_A_iVqHq4Hr1_1;
	wire w_dff_A_QF5aFoH61_1;
	wire w_dff_A_9VP9IOha1_1;
	wire w_dff_A_zKqqXszk4_1;
	wire w_dff_A_wuQD9Hzj0_1;
	wire w_dff_A_VIhe6DUA7_1;
	wire w_dff_A_WbCy81H91_1;
	wire w_dff_A_V4OFxZ083_1;
	wire w_dff_A_tkGJ9t5y6_1;
	wire w_dff_A_DQGtUc2l6_1;
	wire w_dff_A_vfWf3gR25_1;
	wire w_dff_A_nqPUHYk00_1;
	wire w_dff_A_x1s2U30T8_1;
	wire w_dff_A_CtcEoa8n2_1;
	wire w_dff_A_v9xiFeg96_1;
	wire w_dff_A_5C1hva4C5_1;
	wire w_dff_A_2x6djRsS9_1;
	wire w_dff_A_KoqiKnEX4_1;
	wire w_dff_A_e63nU98t4_1;
	wire w_dff_A_kFe3LRGZ8_2;
	wire w_dff_A_wA86aAFS4_2;
	wire w_dff_A_d4rvyG4T9_2;
	wire w_dff_A_0wVrAMwP3_2;
	wire w_dff_A_496hTPo42_2;
	wire w_dff_A_fOGu7ZWA5_2;
	wire w_dff_A_0CweugFC8_2;
	wire w_dff_A_4DpscUuV9_2;
	wire w_dff_A_GsdaWvN54_2;
	wire w_dff_A_IHTSHDyC1_2;
	wire w_dff_A_M8HdTe4Q8_2;
	wire w_dff_A_VrYoCOTw7_2;
	wire w_dff_A_AJeI4UoQ8_2;
	wire w_dff_A_4G8okOjd0_2;
	wire w_dff_A_JXIXWcGo8_2;
	wire w_dff_A_Rj63iQgT8_2;
	wire w_dff_A_qEGBsBzK4_2;
	wire w_dff_B_ZKL3QDgj6_3;
	wire w_dff_A_egaZa6cr5_1;
	wire w_dff_A_JMvy7szU2_1;
	wire w_dff_A_aZAttY8G0_1;
	wire w_dff_A_6jCIhLww4_0;
	wire w_dff_A_XHe6xMWF4_2;
	wire w_dff_A_0bioxm1z1_2;
	wire w_dff_A_S8Ex2UsS9_0;
	wire w_dff_A_VsLbwrtO3_2;
	wire w_dff_A_yAMMVBFC6_0;
	wire w_dff_A_N5jP9i6U3_0;
	wire w_dff_A_qSKEbZh49_0;
	wire w_dff_A_H35nGzRP5_0;
	wire w_dff_A_aI1RUtP61_0;
	wire w_dff_A_F7ERN3hQ1_0;
	wire w_dff_A_iVRRV7Sw1_0;
	wire w_dff_A_cWYLC7ju0_0;
	wire w_dff_A_ywYiSN8k3_0;
	wire w_dff_A_YTEdMcQC8_0;
	wire w_dff_A_wEp1EegM7_0;
	wire w_dff_A_AX1G0bb44_0;
	wire w_dff_A_1qPTpA1q6_0;
	wire w_dff_A_79mn2xNf3_0;
	wire w_dff_A_HDp4Rv4b7_0;
	wire w_dff_A_InXusHiD4_0;
	wire w_dff_A_2J4xUV9f5_0;
	wire w_dff_A_wmUZLzCh4_0;
	wire w_dff_A_p3nTqZD10_0;
	wire w_dff_A_wQHYfsYp4_0;
	wire w_dff_A_RHuUdByJ7_0;
	wire w_dff_A_Abwx3fK25_0;
	wire w_dff_A_taupPDeH9_0;
	wire w_dff_A_Tszw1cSD1_0;
	wire w_dff_A_96EuYVYl3_0;
	wire w_dff_A_WDZpszBJ8_0;
	wire w_dff_A_1aQXot4l1_0;
	wire w_dff_A_61jEzgoa0_0;
	wire w_dff_A_PUd3i7Rp2_0;
	wire w_dff_A_0NHp2NW70_0;
	wire w_dff_A_3cnhfRbG6_2;
	wire w_dff_A_2noCDfoW2_2;
	wire w_dff_A_NQJiFtDC4_2;
	wire w_dff_A_j50Xlt662_2;
	wire w_dff_A_hTCvXI2g6_2;
	wire w_dff_A_N1HLg4Qb8_2;
	wire w_dff_A_isP7eMnG7_2;
	wire w_dff_A_G9GbJgRh8_2;
	wire w_dff_A_obwNyN3M3_2;
	wire w_dff_A_dUxOj9k29_2;
	wire w_dff_A_dyi1Gi8L2_2;
	wire w_dff_A_ezUndS1G2_2;
	wire w_dff_A_XeLfyT332_2;
	wire w_dff_A_4RapG7jq9_2;
	wire w_dff_A_wDowTD480_2;
	wire w_dff_A_guTVlD6N5_2;
	wire w_dff_A_e3s8cSwM6_0;
	wire w_dff_A_aAR6pYCz9_1;
	wire w_dff_A_NOPU9yVk7_2;
	wire w_dff_A_5tQGUpOt2_2;
	wire w_dff_A_rq0kkRTd8_2;
	wire w_dff_A_Z3J2hJSb1_2;
	wire w_dff_A_8ZETPY5M4_0;
	wire w_dff_A_4naE8Tex9_0;
	wire w_dff_A_K1JJceJN9_2;
	wire w_dff_A_WDaLdjET0_2;
	wire w_dff_A_umfdCvHV8_0;
	wire w_dff_A_4X5ktXLG6_2;
	wire w_dff_A_kTSf2yCF4_1;
	wire w_dff_A_qD6GtDDf0_1;
	wire w_dff_A_skFdznOb0_1;
	wire w_dff_A_xir4isHr5_1;
	wire w_dff_A_jkhOXIw50_1;
	wire w_dff_A_4vkk07dQ3_1;
	wire w_dff_A_T1y13SqN0_1;
	wire w_dff_A_DGZgzgEp6_1;
	wire w_dff_A_cY9hvLqp3_1;
	wire w_dff_A_RBGcIbgw2_1;
	wire w_dff_A_Ug09h26b1_1;
	wire w_dff_A_nTFcBRwC5_2;
	wire w_dff_A_jIXxqQBl5_2;
	wire w_dff_A_Ai93AJFG8_2;
	wire w_dff_A_8wK8UJoV2_0;
	wire w_dff_A_6BjZhAeX9_0;
	wire w_dff_A_S5KM9Trm0_0;
	wire w_dff_A_c8gsiFJd5_0;
	wire w_dff_A_SOvO5oUh8_0;
	wire w_dff_A_tz7QtjWd6_0;
	wire w_dff_A_AVbjljYj0_0;
	wire w_dff_A_bzLOMo5p2_0;
	wire w_dff_A_EuImGtAL1_0;
	wire w_dff_A_il6Dvlg90_0;
	wire w_dff_A_ICHD9OEJ4_0;
	wire w_dff_A_ugjitDbz9_0;
	wire w_dff_A_Vpq56JlK0_0;
	wire w_dff_A_MFrcOJQK7_0;
	wire w_dff_A_jn2ogL1S9_0;
	wire w_dff_A_bC1ONhvq0_0;
	wire w_dff_A_USFsF0Q75_0;
	wire w_dff_A_eOJ13Mva0_0;
	wire w_dff_A_Q01RmBgn9_0;
	wire w_dff_A_QyRcSd7n2_0;
	wire w_dff_A_jOVPISwb2_0;
	wire w_dff_A_IRyFOeZM1_0;
	wire w_dff_A_xiulzJwB2_0;
	wire w_dff_A_3NHEjUHK0_0;
	wire w_dff_A_E6yqJQNg3_0;
	wire w_dff_A_kWSj6xz52_0;
	wire w_dff_A_heHbqSsj6_1;
	wire w_dff_A_6FpreaDL9_0;
	wire w_dff_A_oBlulQxO4_0;
	wire w_dff_A_zSHMdOlg5_0;
	wire w_dff_A_3ouQPzKh8_0;
	wire w_dff_A_4Z0zJ60r3_0;
	wire w_dff_A_BM61Geu76_0;
	wire w_dff_A_P98P93Vo1_0;
	wire w_dff_A_1bFkcBog0_0;
	wire w_dff_A_C5vjGe879_0;
	wire w_dff_A_fxx806kt2_0;
	wire w_dff_A_nRxvoZy43_0;
	wire w_dff_A_T1Ru8qFm5_0;
	wire w_dff_A_ZTSJahtc0_0;
	wire w_dff_A_CqozIHur5_0;
	wire w_dff_A_VQDCUjM34_0;
	wire w_dff_A_O3bEJz710_0;
	wire w_dff_A_1GVJ6AsH9_0;
	wire w_dff_A_N0on1wpE3_0;
	wire w_dff_A_mknWWI8a5_0;
	wire w_dff_A_7zuE67D02_0;
	wire w_dff_A_rmUqLk1b0_0;
	wire w_dff_A_p1L3MV9H0_0;
	wire w_dff_A_WhhtPLAe0_0;
	wire w_dff_A_8mTF0rtj6_0;
	wire w_dff_A_mE5NcZom7_0;
	wire w_dff_A_09oKH6DA8_0;
	wire w_dff_A_MhNMV9bW1_0;
	wire w_dff_A_dcDQDPxH8_2;
	wire w_dff_A_2JWF9wm07_0;
	wire w_dff_A_eOMG95CX1_0;
	wire w_dff_A_2tAQ40B94_0;
	wire w_dff_A_k3cg0RrP9_0;
	wire w_dff_A_OKX3pUMK6_0;
	wire w_dff_A_8qzrIc9S6_0;
	wire w_dff_A_zWpc0EmV8_0;
	wire w_dff_A_xeiXKon84_0;
	wire w_dff_A_WMmrDgGo0_0;
	wire w_dff_A_fXDVISIz7_0;
	wire w_dff_A_5KRr7hOJ1_0;
	wire w_dff_A_wNyduM9r0_0;
	wire w_dff_A_TWoDI0xq5_0;
	wire w_dff_A_mVa35RVi0_0;
	wire w_dff_A_5iZI7iGb1_0;
	wire w_dff_A_MLO4bTuK9_0;
	wire w_dff_A_eylU7JFY2_0;
	wire w_dff_A_SJifkAxx4_0;
	wire w_dff_A_ADLAh3eJ8_0;
	wire w_dff_A_MiEXD3jG9_0;
	wire w_dff_A_S8FkLZxb3_0;
	wire w_dff_A_1F2vq7cY6_0;
	wire w_dff_A_LguSs9EC9_2;
	wire w_dff_A_CFNiCZF28_0;
	wire w_dff_A_SxW2B5cl0_0;
	wire w_dff_A_viKuLYhm9_0;
	wire w_dff_A_cK1OG4ZC5_0;
	wire w_dff_A_mRQio0LQ0_0;
	wire w_dff_A_6xS7V23c1_0;
	wire w_dff_A_dHku9i8q2_0;
	wire w_dff_A_qUW0RoQM1_0;
	wire w_dff_A_Nihax5y29_0;
	wire w_dff_A_UAe7Fu759_0;
	wire w_dff_A_vqd355fq0_0;
	wire w_dff_A_fhGLWfSZ6_0;
	wire w_dff_A_AGd7AVLH3_0;
	wire w_dff_A_uzyAGsou2_0;
	wire w_dff_A_VyaPxz1f2_0;
	wire w_dff_A_8RHrabNL8_0;
	wire w_dff_A_UFIMXzq03_0;
	wire w_dff_A_RToiNRdE6_0;
	wire w_dff_A_mvxanOFS4_0;
	wire w_dff_A_Y3Md220M2_0;
	wire w_dff_A_K9ynOQIK4_0;
	wire w_dff_A_qRv3Kthb3_0;
	wire w_dff_A_QrDGQSQd8_0;
	wire w_dff_A_qiXxe7Fc9_0;
	wire w_dff_A_q1pa0OsA6_0;
	wire w_dff_A_jxO7Gb1E1_2;
	wire w_dff_A_2lCTvU9h2_0;
	wire w_dff_A_sMhKaenh0_0;
	wire w_dff_A_tJd3NBRk9_0;
	wire w_dff_A_k5TFpQE33_0;
	wire w_dff_A_qjN0MhyM1_0;
	wire w_dff_A_8mzykBEF3_0;
	wire w_dff_A_O5cozlGr7_0;
	wire w_dff_A_kMvDyWg85_0;
	wire w_dff_A_xGH5Ivs95_0;
	wire w_dff_A_ueyEnQai1_0;
	wire w_dff_A_1csAG2rb0_0;
	wire w_dff_A_YmqN1DgV8_0;
	wire w_dff_A_Ojk52XmW4_0;
	wire w_dff_A_j1ky04Bg4_0;
	wire w_dff_A_AJaRT1qj2_0;
	wire w_dff_A_QmxGzTpy0_0;
	wire w_dff_A_HdJhXA425_0;
	wire w_dff_A_MoOazLC59_0;
	wire w_dff_A_946hA4991_0;
	wire w_dff_A_9FAkzqTC5_0;
	wire w_dff_A_qP85N9KR9_0;
	wire w_dff_A_Cq8yWShR4_0;
	wire w_dff_A_meWnGMiq9_0;
	wire w_dff_A_cmSYvPGX9_0;
	wire w_dff_A_HbUE7IYu9_0;
	wire w_dff_A_HJpBciPx2_0;
	wire w_dff_A_JAByGg7B5_2;
	wire w_dff_A_EoICxVBu2_0;
	wire w_dff_A_gjrpNmAA2_0;
	wire w_dff_A_FAjOD6Oi6_0;
	wire w_dff_A_d6sMEsnZ6_0;
	wire w_dff_A_85CUouSP3_0;
	wire w_dff_A_lFczkg4K6_0;
	wire w_dff_A_VmKEePlN2_0;
	wire w_dff_A_XzLmBfRQ1_0;
	wire w_dff_A_urGzhT8P2_0;
	wire w_dff_A_4gVZ4j902_0;
	wire w_dff_A_C4EbJt2q8_0;
	wire w_dff_A_iCJ2GGev6_0;
	wire w_dff_A_S4Ge7OwR4_0;
	wire w_dff_A_qRdAfI1F8_2;
	wire w_dff_A_OyvXMKs59_0;
	wire w_dff_A_c0es5wGK8_0;
	wire w_dff_A_7Zfn1xMY5_0;
	wire w_dff_A_fknHQfj16_0;
	wire w_dff_A_85QK85lL7_0;
	wire w_dff_A_5GmK2co63_0;
	wire w_dff_A_oEKfbMSB8_0;
	wire w_dff_A_a4QoQGjb7_0;
	wire w_dff_A_FFSEMvOO7_0;
	wire w_dff_A_o8MDBcjX5_0;
	wire w_dff_A_4m1UV7fw5_0;
	wire w_dff_A_UHzT0RaE1_2;
	wire w_dff_A_KjTc5jEp4_0;
	wire w_dff_A_BN5PaiSn9_0;
	wire w_dff_A_ZLF4pp3d5_0;
	wire w_dff_A_lgoO7Orz8_0;
	wire w_dff_A_ZVNovf346_0;
	wire w_dff_A_m3L8a7Bg5_0;
	wire w_dff_A_6yVs5rtw8_0;
	wire w_dff_A_hok2NpAF2_0;
	wire w_dff_A_EdHWmoz13_0;
	wire w_dff_A_s7KFIQBH1_0;
	wire w_dff_A_e250Ta4u5_0;
	wire w_dff_A_cDq0uFlu5_0;
	wire w_dff_A_Q2ojPoe65_0;
	wire w_dff_A_PHITdRC31_2;
	wire w_dff_A_Mib1ZxWW6_0;
	wire w_dff_A_GkwRoEH73_0;
	wire w_dff_A_GDYQeMP93_0;
	wire w_dff_A_KRnIQjkJ0_0;
	wire w_dff_A_s9buAJxf5_0;
	wire w_dff_A_izzAIYDC1_0;
	wire w_dff_A_aDbrixL86_0;
	wire w_dff_A_qFi8lNVn2_0;
	wire w_dff_A_0XfjDTOX8_1;
	wire w_dff_A_OFpUOMpJ2_0;
	wire w_dff_A_gpCErC2J7_0;
	wire w_dff_A_1XaNwXtd4_0;
	wire w_dff_A_zaFEr2Qo4_0;
	wire w_dff_A_fjYciVHo3_0;
	wire w_dff_A_2mzac4AP3_0;
	wire w_dff_A_xToQ7eE15_0;
	wire w_dff_A_C3fHhtX00_0;
	wire w_dff_A_B1rZOdhm8_0;
	wire w_dff_A_RWQgGR7b9_0;
	wire w_dff_A_TJTCX4ic6_0;
	wire w_dff_A_pYpDbVvt6_0;
	wire w_dff_A_w0ospIK34_1;
	wire w_dff_A_s3gw2Kpf0_0;
	wire w_dff_A_OsULOYGU0_0;
	wire w_dff_A_Hs7YH4XS1_0;
	wire w_dff_A_kxVVvueZ2_0;
	wire w_dff_A_zwwGGmF66_0;
	wire w_dff_A_Qw83aOJF4_0;
	wire w_dff_A_iP8xR4Dp5_0;
	wire w_dff_A_s1BWpEPJ7_2;
	wire w_dff_A_xIPw46ed7_0;
	wire w_dff_A_Za09WhNt1_0;
	wire w_dff_A_KKwkaz148_0;
	wire w_dff_A_Egy2GMK16_0;
	wire w_dff_A_hKoYBXx60_0;
	wire w_dff_A_L68NbBTi7_0;
	wire w_dff_A_9T1uPaDL7_1;
	wire w_dff_A_Bt9wVzTt8_0;
	wire w_dff_A_XsprfBTq5_0;
	wire w_dff_A_BPJNqi4P9_0;
	wire w_dff_A_2VS1HYFM1_0;
	wire w_dff_A_ebIqPRx40_0;
	wire w_dff_A_AxGVX6TL1_1;
	wire w_dff_A_P9xmPpsY4_0;
	wire w_dff_A_bEHImB6t9_0;
	wire w_dff_A_cdgl24GK6_0;
	wire w_dff_A_P1VdzwAK9_0;
	wire w_dff_A_21LJ38qi8_0;
	wire w_dff_A_Jq6zQMHU6_0;
	wire w_dff_A_4z7A7QZb0_1;
	wire w_dff_A_70oyHGSA9_0;
	wire w_dff_A_K8cjy4tB5_0;
	wire w_dff_A_wsfjiJc34_0;
	wire w_dff_A_DlL4fp6E6_0;
	wire w_dff_A_C38MetWn2_0;
	wire w_dff_A_lKt9RnS31_1;
	wire w_dff_A_eOvyUM789_0;
	wire w_dff_A_zrE6ZEQR2_0;
	wire w_dff_A_Tyi4ypDL0_0;
	wire w_dff_A_1rpzyvbw3_1;
	wire w_dff_A_0f7I85Sz6_0;
	wire w_dff_A_ZtU3tyDA1_0;
	wire w_dff_A_OFjJ8rbw8_0;
	wire w_dff_A_ZFDj4KzA8_1;
	wire w_dff_A_GLrwuIti6_0;
	wire w_dff_A_ntiPQ6aK5_0;
	wire w_dff_A_Pr5W43mi1_0;
	wire w_dff_A_U9Dhhxdh2_1;
	wire w_dff_A_nMRnQXEZ3_2;
	wire w_dff_A_c0IRpd548_0;
	jnot g0000(.din(w_G77_4[2]),.dout(n72),.clk(gclk));
	jnot g0001(.din(w_G50_5[2]),.dout(n73),.clk(gclk));
	jnot g0002(.din(w_G58_5[2]),.dout(n74),.clk(gclk));
	jnot g0003(.din(w_G68_5[2]),.dout(n75),.clk(gclk));
	jand g0004(.dina(w_n75_2[1]),.dinb(w_n74_2[1]),.dout(n76),.clk(gclk));
	jand g0005(.dina(w_n76_0[1]),.dinb(w_n73_2[2]),.dout(n77),.clk(gclk));
	jand g0006(.dina(w_n77_0[1]),.dinb(w_n72_1[2]),.dout(w_dff_A_Ai93AJFG8_2),.clk(gclk));
	jnot g0007(.din(w_G87_3[2]),.dout(n79),.clk(gclk));
	jnot g0008(.din(w_G97_4[2]),.dout(n80),.clk(gclk));
	jnot g0009(.din(w_G107_4[1]),.dout(n81),.clk(gclk));
	jand g0010(.dina(w_n81_2[1]),.dinb(w_n80_1[2]),.dout(n82),.clk(gclk));
	jor g0011(.dina(n82),.dinb(w_n79_1[2]),.dout(G355_fa_),.clk(gclk));
	jnot g0012(.din(w_G250_0[2]),.dout(n84),.clk(gclk));
	jnot g0013(.din(w_G257_1[2]),.dout(n85),.clk(gclk));
	jnot g0014(.din(w_G264_0[2]),.dout(n86),.clk(gclk));
	jand g0015(.dina(w_n86_0[2]),.dinb(w_n85_0[1]),.dout(n87),.clk(gclk));
	jor g0016(.dina(n87),.dinb(w_n84_1[2]),.dout(n88),.clk(gclk));
	jnot g0017(.din(w_G13_2[1]),.dout(n89),.clk(gclk));
	jand g0018(.dina(w_n89_0[1]),.dinb(w_G1_2[1]),.dout(n90),.clk(gclk));
	jand g0019(.dina(w_n90_0[2]),.dinb(w_G20_6[2]),.dout(n91),.clk(gclk));
	jand g0020(.dina(w_n91_1[2]),.dinb(n88),.dout(n92),.clk(gclk));
	jor g0021(.dina(w_n85_0[0]),.dinb(w_n80_1[1]),.dout(n93),.clk(gclk));
	jnot g0022(.din(w_G244_1[1]),.dout(n94),.clk(gclk));
	jor g0023(.dina(w_n94_0[2]),.dinb(w_n72_1[1]),.dout(n95),.clk(gclk));
	jnot g0024(.din(w_G238_0[2]),.dout(n96),.clk(gclk));
	jor g0025(.dina(w_n96_0[2]),.dinb(w_n75_2[0]),.dout(n97),.clk(gclk));
	jand g0026(.dina(n97),.dinb(n95),.dout(n98),.clk(gclk));
	jnot g0027(.din(w_G226_1[2]),.dout(n99),.clk(gclk));
	jor g0028(.dina(n99),.dinb(w_n73_2[1]),.dout(n100),.clk(gclk));
	jand g0029(.dina(w_dff_B_zCONiVVC8_0),.dinb(n98),.dout(n101),.clk(gclk));
	jand g0030(.dina(n101),.dinb(w_dff_B_hbZGDMrg3_1),.dout(n102),.clk(gclk));
	jnot g0031(.din(w_G232_1[2]),.dout(n103),.clk(gclk));
	jor g0032(.dina(n103),.dinb(w_n74_2[0]),.dout(n104),.clk(gclk));
	jnot g0033(.din(w_G116_5[2]),.dout(n105),.clk(gclk));
	jnot g0034(.din(w_G270_0[2]),.dout(n106),.clk(gclk));
	jor g0035(.dina(n106),.dinb(w_n105_1[1]),.dout(n107),.clk(gclk));
	jand g0036(.dina(n107),.dinb(n104),.dout(n108),.clk(gclk));
	jor g0037(.dina(w_n86_0[1]),.dinb(w_n81_2[0]),.dout(n109),.clk(gclk));
	jand g0038(.dina(w_dff_B_udMr7RwF5_0),.dinb(n108),.dout(n110),.clk(gclk));
	jand g0039(.dina(w_G20_6[1]),.dinb(w_G1_2[0]),.dout(n111),.clk(gclk));
	jnot g0040(.din(w_n111_0[2]),.dout(n112),.clk(gclk));
	jor g0041(.dina(w_n84_1[1]),.dinb(w_n79_1[1]),.dout(n113),.clk(gclk));
	jand g0042(.dina(n113),.dinb(w_n112_0[1]),.dout(n114),.clk(gclk));
	jand g0043(.dina(w_dff_B_q71j2OGx8_0),.dinb(n110),.dout(n115),.clk(gclk));
	jand g0044(.dina(n115),.dinb(n102),.dout(n116),.clk(gclk));
	jnot g0045(.din(w_n76_0[0]),.dout(n117),.clk(gclk));
	jand g0046(.dina(n117),.dinb(w_G50_5[1]),.dout(n118),.clk(gclk));
	jnot g0047(.din(w_n118_0[2]),.dout(n119),.clk(gclk));
	jand g0048(.dina(w_n111_0[1]),.dinb(w_G13_2[0]),.dout(n120),.clk(gclk));
	jand g0049(.dina(w_n120_0[1]),.dinb(n119),.dout(n121),.clk(gclk));
	jor g0050(.dina(n121),.dinb(n116),.dout(n122),.clk(gclk));
	jor g0051(.dina(n122),.dinb(w_dff_B_Pb9h1aHH6_1),.dout(w_dff_A_dcDQDPxH8_2),.clk(gclk));
	jxor g0052(.dina(w_G270_0[1]),.dinb(w_n86_0[0]),.dout(n124),.clk(gclk));
	jxor g0053(.dina(w_G257_1[1]),.dinb(w_G250_0[1]),.dout(n125),.clk(gclk));
	jxor g0054(.dina(w_dff_B_PHRg72GV4_0),.dinb(n124),.dout(n126),.clk(gclk));
	jnot g0055(.din(w_n126_0[1]),.dout(n127),.clk(gclk));
	jxor g0056(.dina(w_G244_1[0]),.dinb(w_n96_0[1]),.dout(n128),.clk(gclk));
	jxor g0057(.dina(w_G232_1[1]),.dinb(w_G226_1[1]),.dout(n129),.clk(gclk));
	jxor g0058(.dina(w_dff_B_3f5k93LL3_0),.dinb(n128),.dout(n130),.clk(gclk));
	jxor g0059(.dina(w_n130_0[1]),.dinb(n127),.dout(w_dff_A_LguSs9EC9_2),.clk(gclk));
	jxor g0060(.dina(w_G58_5[1]),.dinb(w_G50_5[0]),.dout(n132),.clk(gclk));
	jxor g0061(.dina(w_G77_4[1]),.dinb(w_G68_5[1]),.dout(n133),.clk(gclk));
	jxor g0062(.dina(n133),.dinb(n132),.dout(n134),.clk(gclk));
	jxor g0063(.dina(w_G116_5[1]),.dinb(w_n81_1[2]),.dout(n135),.clk(gclk));
	jxor g0064(.dina(w_G97_4[1]),.dinb(w_G87_3[1]),.dout(n136),.clk(gclk));
	jxor g0065(.dina(w_dff_B_DZJ2aS4s0_0),.dinb(n135),.dout(n137),.clk(gclk));
	jxor g0066(.dina(w_n137_0[1]),.dinb(w_n134_0[1]),.dout(w_dff_A_jxO7Gb1E1_2),.clk(gclk));
	jand g0067(.dina(w_G13_1[2]),.dinb(w_G1_1[2]),.dout(n139),.clk(gclk));
	jand g0068(.dina(w_n111_0[0]),.dinb(w_G33_12[2]),.dout(n140),.clk(gclk));
	jor g0069(.dina(w_n140_0[1]),.dinb(w_n139_1[2]),.dout(n141),.clk(gclk));
	jnot g0070(.din(w_G1_1[1]),.dout(n142),.clk(gclk));
	jand g0071(.dina(w_G13_1[1]),.dinb(w_n142_2[1]),.dout(n143),.clk(gclk));
	jand g0072(.dina(w_n143_0[1]),.dinb(w_G20_6[0]),.dout(n144),.clk(gclk));
	jor g0073(.dina(w_n144_2[1]),.dinb(w_n141_3[1]),.dout(n145),.clk(gclk));
	jand g0074(.dina(w_G33_12[1]),.dinb(w_n142_2[0]),.dout(n146),.clk(gclk));
	jor g0075(.dina(w_dff_B_TWpw5Lkn9_0),.dinb(n145),.dout(n147),.clk(gclk));
	jnot g0076(.din(w_n147_0[2]),.dout(n148),.clk(gclk));
	jand g0077(.dina(w_n148_0[1]),.dinb(w_G116_5[0]),.dout(n149),.clk(gclk));
	jand g0078(.dina(w_G116_4[2]),.dinb(w_G20_5[2]),.dout(n150),.clk(gclk));
	jnot g0079(.din(w_G20_5[1]),.dout(n151),.clk(gclk));
	jand g0080(.dina(w_G283_3[2]),.dinb(w_G33_12[0]),.dout(n152),.clk(gclk));
	jnot g0081(.din(w_G33_11[2]),.dout(n153),.clk(gclk));
	jand g0082(.dina(w_G97_4[0]),.dinb(w_n153_8[1]),.dout(n154),.clk(gclk));
	jor g0083(.dina(n154),.dinb(w_n152_0[2]),.dout(n155),.clk(gclk));
	jand g0084(.dina(n155),.dinb(w_n151_6[1]),.dout(n156),.clk(gclk));
	jor g0085(.dina(n156),.dinb(w_dff_B_QKp3wjYK2_1),.dout(n157),.clk(gclk));
	jand g0086(.dina(n157),.dinb(w_n141_3[0]),.dout(n158),.clk(gclk));
	jand g0087(.dina(w_n144_2[0]),.dinb(w_n105_1[0]),.dout(n159),.clk(gclk));
	jor g0088(.dina(w_dff_B_M2hcu2Iu9_0),.dinb(n158),.dout(n160),.clk(gclk));
	jor g0089(.dina(n160),.dinb(n149),.dout(n161),.clk(gclk));
	jnot g0090(.din(w_n161_0[2]),.dout(n162),.clk(gclk));
	jnot g0091(.din(w_G41_0[2]),.dout(n163),.clk(gclk));
	jand g0092(.dina(w_G45_1[1]),.dinb(w_n142_1[2]),.dout(n164),.clk(gclk));
	jand g0093(.dina(w_n164_0[2]),.dinb(w_n163_1[1]),.dout(n165),.clk(gclk));
	jnot g0094(.din(w_n139_1[1]),.dout(n166),.clk(gclk));
	jand g0095(.dina(w_G41_0[1]),.dinb(w_G33_11[1]),.dout(n167),.clk(gclk));
	jor g0096(.dina(w_n167_0[1]),.dinb(n166),.dout(n168),.clk(gclk));
	jand g0097(.dina(w_n168_5[1]),.dinb(w_G274_0[2]),.dout(n169),.clk(gclk));
	jand g0098(.dina(w_n169_0[1]),.dinb(w_n165_0[1]),.dout(n170),.clk(gclk));
	jnot g0099(.din(w_n167_0[0]),.dout(n171),.clk(gclk));
	jand g0100(.dina(n171),.dinb(w_n139_1[0]),.dout(n172),.clk(gclk));
	jand g0101(.dina(w_G1698_0[2]),.dinb(w_n153_8[0]),.dout(n173),.clk(gclk));
	jand g0102(.dina(w_n173_3[1]),.dinb(w_G264_0[1]),.dout(n174),.clk(gclk));
	jand g0103(.dina(w_G303_2[2]),.dinb(w_G33_11[0]),.dout(n175),.clk(gclk));
	jnot g0104(.din(w_G1698_0[1]),.dout(n176),.clk(gclk));
	jand g0105(.dina(w_n176_0[1]),.dinb(w_n153_7[2]),.dout(n177),.clk(gclk));
	jand g0106(.dina(w_n177_1[2]),.dinb(w_G257_1[0]),.dout(n178),.clk(gclk));
	jor g0107(.dina(n178),.dinb(w_dff_B_BgZDjfnJ5_1),.dout(n179),.clk(gclk));
	jor g0108(.dina(n179),.dinb(w_dff_B_dI5peQw07_1),.dout(n180),.clk(gclk));
	jand g0109(.dina(n180),.dinb(w_n172_4[2]),.dout(n181),.clk(gclk));
	jnot g0110(.din(w_n165_0[0]),.dout(n182),.clk(gclk));
	jand g0111(.dina(w_n168_5[0]),.dinb(w_G270_0[0]),.dout(n183),.clk(gclk));
	jand g0112(.dina(n183),.dinb(w_n182_1[1]),.dout(n184),.clk(gclk));
	jor g0113(.dina(w_dff_B_GcnqWhjj5_0),.dinb(n181),.dout(n185),.clk(gclk));
	jor g0114(.dina(n185),.dinb(w_n170_0[2]),.dout(n186),.clk(gclk));
	jand g0115(.dina(w_n186_1[2]),.dinb(w_G169_3[1]),.dout(n187),.clk(gclk));
	jnot g0116(.din(n187),.dout(n188),.clk(gclk));
	jnot g0117(.din(w_G179_2[2]),.dout(n189),.clk(gclk));
	jor g0118(.dina(w_n186_1[1]),.dinb(w_n189_2[2]),.dout(n190),.clk(gclk));
	jand g0119(.dina(w_n190_0[1]),.dinb(n188),.dout(n191),.clk(gclk));
	jor g0120(.dina(n191),.dinb(w_dff_B_4iA5VZ472_1),.dout(n192),.clk(gclk));
	jand g0121(.dina(w_n186_1[0]),.dinb(w_G200_3[1]),.dout(n193),.clk(gclk));
	jnot g0122(.din(w_n186_0[2]),.dout(n194),.clk(gclk));
	jand g0123(.dina(n194),.dinb(w_G190_4[2]),.dout(n195),.clk(gclk));
	jor g0124(.dina(n195),.dinb(w_n161_0[1]),.dout(n196),.clk(gclk));
	jor g0125(.dina(n196),.dinb(w_dff_B_tISGEVh33_1),.dout(n197),.clk(gclk));
	jand g0126(.dina(n197),.dinb(w_n192_0[2]),.dout(n198),.clk(gclk));
	jnot g0127(.din(w_G169_3[0]),.dout(n199),.clk(gclk));
	jand g0128(.dina(w_n168_4[2]),.dinb(w_G264_0[0]),.dout(n200),.clk(gclk));
	jand g0129(.dina(n200),.dinb(w_n182_1[0]),.dout(n201),.clk(gclk));
	jand g0130(.dina(w_n173_3[0]),.dinb(w_G257_0[2]),.dout(n202),.clk(gclk));
	jand g0131(.dina(w_G294_3[1]),.dinb(w_G33_10[2]),.dout(n203),.clk(gclk));
	jnot g0132(.din(n203),.dout(n204),.clk(gclk));
	jor g0133(.dina(w_G1698_0[0]),.dinb(w_G33_10[1]),.dout(n205),.clk(gclk));
	jor g0134(.dina(w_n205_1[1]),.dinb(w_n84_1[0]),.dout(n206),.clk(gclk));
	jand g0135(.dina(n206),.dinb(n204),.dout(n207),.clk(gclk));
	jnot g0136(.din(w_n207_0[1]),.dout(n208),.clk(gclk));
	jor g0137(.dina(n208),.dinb(w_n202_0[1]),.dout(n209),.clk(gclk));
	jand g0138(.dina(n209),.dinb(w_n172_4[1]),.dout(n210),.clk(gclk));
	jor g0139(.dina(n210),.dinb(w_n170_0[1]),.dout(n211),.clk(gclk));
	jor g0140(.dina(n211),.dinb(w_n201_0[1]),.dout(n212),.clk(gclk));
	jand g0141(.dina(w_n212_1[1]),.dinb(w_n199_0[2]),.dout(n213),.clk(gclk));
	jand g0142(.dina(w_n148_0[0]),.dinb(w_G107_4[0]),.dout(n214),.clk(gclk));
	jor g0143(.dina(w_n140_0[0]),.dinb(w_G13_1[0]),.dout(n215),.clk(gclk));
	jand g0144(.dina(w_n81_1[1]),.dinb(w_G20_5[0]),.dout(n216),.clk(gclk));
	jand g0145(.dina(w_dff_B_b6QY8yMK0_0),.dinb(w_n215_0[1]),.dout(n217),.clk(gclk));
	jand g0146(.dina(w_G116_4[1]),.dinb(w_G33_10[0]),.dout(n218),.clk(gclk));
	jand g0147(.dina(w_G87_3[0]),.dinb(w_n153_7[1]),.dout(n219),.clk(gclk));
	jor g0148(.dina(n219),.dinb(w_n218_0[1]),.dout(n220),.clk(gclk));
	jand g0149(.dina(n220),.dinb(w_n141_2[2]),.dout(n221),.clk(gclk));
	jand g0150(.dina(n221),.dinb(w_n151_6[0]),.dout(n222),.clk(gclk));
	jor g0151(.dina(n222),.dinb(w_dff_B_v4umk7t39_1),.dout(n223),.clk(gclk));
	jor g0152(.dina(w_dff_B_3956jpsI0_0),.dinb(n214),.dout(n224),.clk(gclk));
	jnot g0153(.din(w_n224_1[1]),.dout(n225),.clk(gclk));
	jnot g0154(.din(w_n201_0[0]),.dout(n226),.clk(gclk));
	jnot g0155(.din(w_G274_0[1]),.dout(n227),.clk(gclk));
	jor g0156(.dina(w_n172_4[0]),.dinb(w_dff_B_vjIuho306_1),.dout(n228),.clk(gclk));
	jor g0157(.dina(n228),.dinb(w_n182_0[2]),.dout(n229),.clk(gclk));
	jnot g0158(.din(w_n202_0[0]),.dout(n230),.clk(gclk));
	jand g0159(.dina(w_n207_0[0]),.dinb(n230),.dout(n231),.clk(gclk));
	jor g0160(.dina(n231),.dinb(w_n168_4[1]),.dout(n232),.clk(gclk));
	jand g0161(.dina(n232),.dinb(w_n229_0[1]),.dout(n233),.clk(gclk));
	jand g0162(.dina(n233),.dinb(w_dff_B_H5DWbEEY9_1),.dout(n234),.clk(gclk));
	jand g0163(.dina(w_n234_1[1]),.dinb(w_n189_2[1]),.dout(n235),.clk(gclk));
	jor g0164(.dina(n235),.dinb(w_n225_0[1]),.dout(n236),.clk(gclk));
	jor g0165(.dina(n236),.dinb(w_n213_0[1]),.dout(n237),.clk(gclk));
	jand g0166(.dina(w_n234_1[0]),.dinb(w_G190_4[1]),.dout(n238),.clk(gclk));
	jand g0167(.dina(w_n212_1[0]),.dinb(w_G200_3[0]),.dout(n239),.clk(gclk));
	jor g0168(.dina(n239),.dinb(w_n224_1[0]),.dout(n240),.clk(gclk));
	jor g0169(.dina(n240),.dinb(w_n238_0[1]),.dout(n241),.clk(gclk));
	jand g0170(.dina(n241),.dinb(w_n237_0[2]),.dout(n242),.clk(gclk));
	jand g0171(.dina(w_n173_2[2]),.dinb(w_G244_0[2]),.dout(n243),.clk(gclk));
	jnot g0172(.din(w_n243_0[1]),.dout(n244),.clk(gclk));
	jnot g0173(.din(w_n218_0[0]),.dout(n245),.clk(gclk));
	jor g0174(.dina(w_n205_1[0]),.dinb(w_n96_0[0]),.dout(n246),.clk(gclk));
	jand g0175(.dina(n246),.dinb(n245),.dout(n247),.clk(gclk));
	jand g0176(.dina(w_n247_0[1]),.dinb(n244),.dout(n248),.clk(gclk));
	jand g0177(.dina(n248),.dinb(w_n172_3[2]),.dout(n249),.clk(gclk));
	jor g0178(.dina(w_n164_0[1]),.dinb(w_n84_0[2]),.dout(n250),.clk(gclk));
	jand g0179(.dina(w_n164_0[0]),.dinb(w_G274_0[0]),.dout(n251),.clk(gclk));
	jnot g0180(.din(w_n251_0[1]),.dout(n252),.clk(gclk));
	jand g0181(.dina(n252),.dinb(w_n250_0[1]),.dout(n253),.clk(gclk));
	jand g0182(.dina(n253),.dinb(w_n168_4[0]),.dout(n254),.clk(gclk));
	jor g0183(.dina(n254),.dinb(n249),.dout(n255),.clk(gclk));
	jand g0184(.dina(w_n255_1[1]),.dinb(w_n189_2[0]),.dout(n256),.clk(gclk));
	jor g0185(.dina(w_n147_0[1]),.dinb(w_n79_1[0]),.dout(n257),.clk(gclk));
	jand g0186(.dina(w_n80_1[0]),.dinb(w_n79_0[2]),.dout(n258),.clk(gclk));
	jand g0187(.dina(n258),.dinb(w_n81_1[0]),.dout(n259),.clk(gclk));
	jand g0188(.dina(w_n259_0[1]),.dinb(w_G20_4[2]),.dout(n260),.clk(gclk));
	jnot g0189(.din(w_n141_2[1]),.dout(n261),.clk(gclk));
	jand g0190(.dina(w_G97_3[2]),.dinb(w_G33_9[2]),.dout(n262),.clk(gclk));
	jnot g0191(.din(w_n262_0[2]),.dout(n263),.clk(gclk));
	jor g0192(.dina(w_n75_1[2]),.dinb(w_G33_9[1]),.dout(n264),.clk(gclk));
	jand g0193(.dina(n264),.dinb(w_n151_5[2]),.dout(n265),.clk(gclk));
	jand g0194(.dina(n265),.dinb(w_dff_B_0yChTZMT8_1),.dout(n266),.clk(gclk));
	jor g0195(.dina(n266),.dinb(w_n261_1[2]),.dout(n267),.clk(gclk));
	jor g0196(.dina(n267),.dinb(w_n260_0[1]),.dout(n268),.clk(gclk));
	jand g0197(.dina(w_n144_1[2]),.dinb(w_n79_0[1]),.dout(n269),.clk(gclk));
	jnot g0198(.din(w_n269_0[1]),.dout(n270),.clk(gclk));
	jand g0199(.dina(w_dff_B_zLrZuBmg2_0),.dinb(n268),.dout(n271),.clk(gclk));
	jand g0200(.dina(n271),.dinb(w_n257_0[1]),.dout(n272),.clk(gclk));
	jnot g0201(.din(w_n247_0[0]),.dout(n273),.clk(gclk));
	jor g0202(.dina(n273),.dinb(w_n243_0[0]),.dout(n274),.clk(gclk));
	jor g0203(.dina(n274),.dinb(w_n168_3[2]),.dout(n275),.clk(gclk));
	jnot g0204(.din(w_n250_0[0]),.dout(n276),.clk(gclk));
	jor g0205(.dina(w_n251_0[0]),.dinb(n276),.dout(n277),.clk(gclk));
	jor g0206(.dina(n277),.dinb(w_n172_3[1]),.dout(n278),.clk(gclk));
	jand g0207(.dina(n278),.dinb(n275),.dout(n279),.clk(gclk));
	jand g0208(.dina(w_n279_1[1]),.dinb(w_n199_0[1]),.dout(n280),.clk(gclk));
	jor g0209(.dina(n280),.dinb(w_n272_0[1]),.dout(n281),.clk(gclk));
	jor g0210(.dina(n281),.dinb(w_n256_0[1]),.dout(n282),.clk(gclk));
	jand g0211(.dina(w_n279_1[0]),.dinb(w_G200_2[2]),.dout(n283),.clk(gclk));
	jnot g0212(.din(w_n257_0[0]),.dout(n284),.clk(gclk));
	jnot g0213(.din(w_n260_0[0]),.dout(n285),.clk(gclk));
	jand g0214(.dina(w_G68_5[0]),.dinb(w_n153_7[0]),.dout(n286),.clk(gclk));
	jor g0215(.dina(n286),.dinb(w_G20_4[1]),.dout(n287),.clk(gclk));
	jor g0216(.dina(n287),.dinb(w_n262_0[1]),.dout(n288),.clk(gclk));
	jand g0217(.dina(n288),.dinb(w_n141_2[0]),.dout(n289),.clk(gclk));
	jand g0218(.dina(n289),.dinb(n285),.dout(n290),.clk(gclk));
	jor g0219(.dina(w_n269_0[0]),.dinb(n290),.dout(n291),.clk(gclk));
	jor g0220(.dina(n291),.dinb(n284),.dout(n292),.clk(gclk));
	jand g0221(.dina(w_n255_1[0]),.dinb(w_G190_4[0]),.dout(n293),.clk(gclk));
	jor g0222(.dina(n293),.dinb(w_n292_0[2]),.dout(n294),.clk(gclk));
	jor g0223(.dina(n294),.dinb(w_n283_0[1]),.dout(n295),.clk(gclk));
	jand g0224(.dina(n295),.dinb(w_n282_0[1]),.dout(n296),.clk(gclk));
	jand g0225(.dina(w_n168_3[1]),.dinb(w_G257_0[1]),.dout(n297),.clk(gclk));
	jand g0226(.dina(n297),.dinb(w_n182_0[1]),.dout(n298),.clk(gclk));
	jnot g0227(.din(w_n298_0[1]),.dout(n299),.clk(gclk));
	jor g0228(.dina(w_n176_0[0]),.dinb(w_G33_9[0]),.dout(n300),.clk(gclk));
	jor g0229(.dina(n300),.dinb(w_n84_0[1]),.dout(n301),.clk(gclk));
	jnot g0230(.din(w_n152_0[1]),.dout(n302),.clk(gclk));
	jor g0231(.dina(w_n205_0[2]),.dinb(w_n94_0[1]),.dout(n303),.clk(gclk));
	jand g0232(.dina(n303),.dinb(n302),.dout(n304),.clk(gclk));
	jand g0233(.dina(n304),.dinb(n301),.dout(n305),.clk(gclk));
	jor g0234(.dina(n305),.dinb(w_n168_3[0]),.dout(n306),.clk(gclk));
	jand g0235(.dina(n306),.dinb(w_n229_0[0]),.dout(n307),.clk(gclk));
	jand g0236(.dina(n307),.dinb(n299),.dout(n308),.clk(gclk));
	jand g0237(.dina(w_n308_1[2]),.dinb(w_G190_3[2]),.dout(n309),.clk(gclk));
	jor g0238(.dina(w_n147_0[0]),.dinb(w_n80_0[2]),.dout(n310),.clk(gclk));
	jnot g0239(.din(w_n310_0[1]),.dout(n311),.clk(gclk));
	jxor g0240(.dina(w_G107_3[2]),.dinb(w_G97_3[1]),.dout(n312),.clk(gclk));
	jand g0241(.dina(w_n312_0[1]),.dinb(w_G20_4[0]),.dout(n313),.clk(gclk));
	jnot g0242(.din(w_n313_0[1]),.dout(n314),.clk(gclk));
	jand g0243(.dina(w_G107_3[1]),.dinb(w_G33_8[2]),.dout(n315),.clk(gclk));
	jand g0244(.dina(w_G77_4[0]),.dinb(w_n153_6[2]),.dout(n316),.clk(gclk));
	jor g0245(.dina(n316),.dinb(w_G20_3[2]),.dout(n317),.clk(gclk));
	jor g0246(.dina(n317),.dinb(w_n315_0[2]),.dout(n318),.clk(gclk));
	jand g0247(.dina(n318),.dinb(w_n141_1[2]),.dout(n319),.clk(gclk));
	jand g0248(.dina(n319),.dinb(w_dff_B_RxrF3lmL5_1),.dout(n320),.clk(gclk));
	jand g0249(.dina(w_n144_1[1]),.dinb(w_n80_0[1]),.dout(n321),.clk(gclk));
	jor g0250(.dina(w_n321_0[1]),.dinb(n320),.dout(n322),.clk(gclk));
	jor g0251(.dina(n322),.dinb(n311),.dout(n323),.clk(gclk));
	jand g0252(.dina(w_n173_2[1]),.dinb(w_G250_0[0]),.dout(n324),.clk(gclk));
	jand g0253(.dina(w_n177_1[1]),.dinb(w_G244_0[1]),.dout(n325),.clk(gclk));
	jor g0254(.dina(n325),.dinb(w_n152_0[0]),.dout(n326),.clk(gclk));
	jor g0255(.dina(n326),.dinb(w_dff_B_acPEU2UT6_1),.dout(n327),.clk(gclk));
	jand g0256(.dina(n327),.dinb(w_n172_3[0]),.dout(n328),.clk(gclk));
	jor g0257(.dina(n328),.dinb(w_n170_0[0]),.dout(n329),.clk(gclk));
	jor g0258(.dina(n329),.dinb(w_n298_0[0]),.dout(n330),.clk(gclk));
	jand g0259(.dina(w_n330_0[2]),.dinb(w_G200_2[1]),.dout(n331),.clk(gclk));
	jor g0260(.dina(n331),.dinb(w_n323_0[2]),.dout(n332),.clk(gclk));
	jor g0261(.dina(n332),.dinb(w_n309_0[1]),.dout(n333),.clk(gclk));
	jor g0262(.dina(w_n308_1[1]),.dinb(w_G169_2[2]),.dout(n334),.clk(gclk));
	jnot g0263(.din(w_n334_0[1]),.dout(n335),.clk(gclk));
	jnot g0264(.din(w_n315_0[1]),.dout(n336),.clk(gclk));
	jor g0265(.dina(w_n72_1[0]),.dinb(w_G33_8[1]),.dout(n337),.clk(gclk));
	jand g0266(.dina(n337),.dinb(w_n151_5[1]),.dout(n338),.clk(gclk));
	jand g0267(.dina(n338),.dinb(w_dff_B_aDt2lZxg4_1),.dout(n339),.clk(gclk));
	jor g0268(.dina(n339),.dinb(w_n261_1[1]),.dout(n340),.clk(gclk));
	jor g0269(.dina(n340),.dinb(w_n313_0[0]),.dout(n341),.clk(gclk));
	jnot g0270(.din(w_n321_0[0]),.dout(n342),.clk(gclk));
	jand g0271(.dina(w_dff_B_vGb3QaKr3_0),.dinb(n341),.dout(n343),.clk(gclk));
	jand g0272(.dina(n343),.dinb(w_n310_0[0]),.dout(n344),.clk(gclk));
	jand g0273(.dina(w_n308_1[0]),.dinb(w_n189_1[2]),.dout(n345),.clk(gclk));
	jor g0274(.dina(n345),.dinb(w_n344_0[1]),.dout(n346),.clk(gclk));
	jor g0275(.dina(n346),.dinb(n335),.dout(n347),.clk(gclk));
	jand g0276(.dina(w_n347_0[1]),.dinb(w_n333_0[1]),.dout(n348),.clk(gclk));
	jand g0277(.dina(w_n348_0[1]),.dinb(w_dff_B_7B0RoYiB7_1),.dout(n349),.clk(gclk));
	jand g0278(.dina(w_n349_0[1]),.dinb(w_n242_0[2]),.dout(n350),.clk(gclk));
	jand g0279(.dina(w_n350_0[1]),.dinb(w_n198_0[2]),.dout(n351),.clk(gclk));
	jnot g0280(.din(w_G45_1[0]),.dout(n352),.clk(gclk));
	jand g0281(.dina(w_n352_1[1]),.dinb(w_n163_1[0]),.dout(n353),.clk(gclk));
	jor g0282(.dina(n353),.dinb(w_G1_1[0]),.dout(n354),.clk(gclk));
	jnot g0283(.din(w_n354_1[1]),.dout(n355),.clk(gclk));
	jand g0284(.dina(w_n355_0[1]),.dinb(w_n169_0[0]),.dout(n356),.clk(gclk));
	jnot g0285(.din(w_n356_1[1]),.dout(n357),.clk(gclk));
	jand g0286(.dina(w_n173_2[0]),.dinb(w_G238_0[1]),.dout(n358),.clk(gclk));
	jand g0287(.dina(w_n177_1[0]),.dinb(w_G232_1[0]),.dout(n359),.clk(gclk));
	jor g0288(.dina(n359),.dinb(w_n315_0[0]),.dout(n360),.clk(gclk));
	jor g0289(.dina(n360),.dinb(w_dff_B_pGicBI5G6_1),.dout(n361),.clk(gclk));
	jand g0290(.dina(n361),.dinb(w_n172_2[2]),.dout(n362),.clk(gclk));
	jnot g0291(.din(n362),.dout(n363),.clk(gclk));
	jor g0292(.dina(w_n355_0[0]),.dinb(w_n94_0[0]),.dout(n364),.clk(gclk));
	jor g0293(.dina(n364),.dinb(w_n172_2[1]),.dout(n365),.clk(gclk));
	jand g0294(.dina(w_dff_B_jLV0ghFw1_0),.dinb(n363),.dout(n366),.clk(gclk));
	jand g0295(.dina(n366),.dinb(w_n357_0[1]),.dout(n367),.clk(gclk));
	jnot g0296(.din(w_n367_1[1]),.dout(n368),.clk(gclk));
	jand g0297(.dina(n368),.dinb(w_n199_0[0]),.dout(n369),.clk(gclk));
	jand g0298(.dina(w_G87_2[2]),.dinb(w_G33_8[0]),.dout(n370),.clk(gclk));
	jand g0299(.dina(w_G58_5[0]),.dinb(w_n153_6[1]),.dout(n371),.clk(gclk));
	jor g0300(.dina(n371),.dinb(w_n370_0[1]),.dout(n372),.clk(gclk));
	jand g0301(.dina(n372),.dinb(w_n151_5[0]),.dout(n373),.clk(gclk));
	jand g0302(.dina(n373),.dinb(w_n141_1[1]),.dout(n374),.clk(gclk));
	jand g0303(.dina(w_n139_0[2]),.dinb(w_n151_4[2]),.dout(n375),.clk(gclk));
	jnot g0304(.din(w_n375_0[1]),.dout(n376),.clk(gclk));
	jand g0305(.dina(w_G20_3[1]),.dinb(w_n142_1[1]),.dout(n377),.clk(gclk));
	jnot g0306(.din(n377),.dout(n378),.clk(gclk));
	jand g0307(.dina(w_n378_0[1]),.dinb(w_G77_3[2]),.dout(n379),.clk(gclk));
	jand g0308(.dina(n379),.dinb(w_dff_B_aEtb0mcV1_1),.dout(n380),.clk(gclk));
	jand g0309(.dina(w_n144_1[0]),.dinb(w_n72_0[2]),.dout(n381),.clk(gclk));
	jor g0310(.dina(w_dff_B_2c83vRPV0_0),.dinb(n380),.dout(n382),.clk(gclk));
	jor g0311(.dina(n382),.dinb(w_dff_B_2DwCmg7O1_1),.dout(n383),.clk(gclk));
	jnot g0312(.din(w_n383_0[2]),.dout(n384),.clk(gclk));
	jand g0313(.dina(w_n367_1[0]),.dinb(w_n189_1[1]),.dout(n385),.clk(gclk));
	jor g0314(.dina(n385),.dinb(w_dff_B_IAH45NQo8_1),.dout(n386),.clk(gclk));
	jor g0315(.dina(n386),.dinb(n369),.dout(n387),.clk(gclk));
	jnot g0316(.din(w_G200_2[0]),.dout(n388),.clk(gclk));
	jor g0317(.dina(w_n367_0[2]),.dinb(w_n388_2[1]),.dout(n389),.clk(gclk));
	jnot g0318(.din(n389),.dout(n390),.clk(gclk));
	jand g0319(.dina(w_n367_0[1]),.dinb(w_G190_3[1]),.dout(n391),.clk(gclk));
	jor g0320(.dina(n391),.dinb(w_n383_0[1]),.dout(n392),.clk(gclk));
	jor g0321(.dina(n392),.dinb(n390),.dout(n393),.clk(gclk));
	jand g0322(.dina(n393),.dinb(w_n387_0[2]),.dout(n394),.clk(gclk));
	jnot g0323(.din(w_n394_0[1]),.dout(n395),.clk(gclk));
	jand g0324(.dina(w_n168_2[2]),.dinb(w_G238_0[0]),.dout(n396),.clk(gclk));
	jand g0325(.dina(n396),.dinb(w_n354_1[0]),.dout(n397),.clk(gclk));
	jand g0326(.dina(w_n173_1[2]),.dinb(w_G232_0[2]),.dout(n398),.clk(gclk));
	jand g0327(.dina(w_n177_0[2]),.dinb(w_G226_1[0]),.dout(n399),.clk(gclk));
	jor g0328(.dina(n399),.dinb(w_n262_0[0]),.dout(n400),.clk(gclk));
	jor g0329(.dina(n400),.dinb(w_dff_B_EwVOvqLO1_1),.dout(n401),.clk(gclk));
	jand g0330(.dina(n401),.dinb(w_n172_2[0]),.dout(n402),.clk(gclk));
	jor g0331(.dina(n402),.dinb(w_n356_1[0]),.dout(n403),.clk(gclk));
	jor g0332(.dina(n403),.dinb(w_dff_B_947c0t5M6_1),.dout(n404),.clk(gclk));
	jnot g0333(.din(w_n404_0[2]),.dout(n405),.clk(gclk));
	jor g0334(.dina(w_n405_0[1]),.dinb(w_G169_2[1]),.dout(n406),.clk(gclk));
	jand g0335(.dina(w_G77_3[1]),.dinb(w_G33_7[2]),.dout(n407),.clk(gclk));
	jand g0336(.dina(w_G50_4[2]),.dinb(w_n153_6[0]),.dout(n408),.clk(gclk));
	jor g0337(.dina(n408),.dinb(w_n407_0[1]),.dout(n409),.clk(gclk));
	jand g0338(.dina(n409),.dinb(w_n141_1[0]),.dout(n410),.clk(gclk));
	jand g0339(.dina(n410),.dinb(w_n151_4[1]),.dout(n411),.clk(gclk));
	jand g0340(.dina(w_n75_1[1]),.dinb(w_G20_3[0]),.dout(n412),.clk(gclk));
	jand g0341(.dina(w_dff_B_lrgl6soP5_0),.dinb(w_n215_0[0]),.dout(n413),.clk(gclk));
	jand g0342(.dina(w_n378_0[0]),.dinb(w_n261_1[0]),.dout(n414),.clk(gclk));
	jand g0343(.dina(w_n414_0[2]),.dinb(w_G68_4[2]),.dout(n415),.clk(gclk));
	jor g0344(.dina(n415),.dinb(w_dff_B_BhPBEMs71_1),.dout(n416),.clk(gclk));
	jor g0345(.dina(n416),.dinb(w_dff_B_bH0fzxpY2_1),.dout(n417),.clk(gclk));
	jor g0346(.dina(w_n404_0[1]),.dinb(w_G179_2[1]),.dout(n418),.clk(gclk));
	jand g0347(.dina(n418),.dinb(w_n417_0[2]),.dout(n419),.clk(gclk));
	jand g0348(.dina(n419),.dinb(n406),.dout(n420),.clk(gclk));
	jand g0349(.dina(w_n405_0[0]),.dinb(w_G190_3[0]),.dout(n421),.clk(gclk));
	jand g0350(.dina(w_n404_0[0]),.dinb(w_G200_1[2]),.dout(n422),.clk(gclk));
	jor g0351(.dina(n422),.dinb(w_n417_0[1]),.dout(n423),.clk(gclk));
	jor g0352(.dina(n423),.dinb(n421),.dout(n424),.clk(gclk));
	jnot g0353(.din(n424),.dout(n425),.clk(gclk));
	jor g0354(.dina(w_n425_0[1]),.dinb(w_n420_0[1]),.dout(n426),.clk(gclk));
	jand g0355(.dina(w_n168_2[1]),.dinb(w_G226_0[2]),.dout(n427),.clk(gclk));
	jand g0356(.dina(n427),.dinb(w_n354_0[2]),.dout(n428),.clk(gclk));
	jnot g0357(.din(w_n428_0[1]),.dout(n429),.clk(gclk));
	jand g0358(.dina(w_n173_1[1]),.dinb(w_G223_0[1]),.dout(n430),.clk(gclk));
	jnot g0359(.din(w_n430_0[1]),.dout(n431),.clk(gclk));
	jnot g0360(.din(w_n407_0[0]),.dout(n432),.clk(gclk));
	jnot g0361(.din(G222),.dout(n433),.clk(gclk));
	jor g0362(.dina(w_n205_0[1]),.dinb(n433),.dout(n434),.clk(gclk));
	jand g0363(.dina(n434),.dinb(n432),.dout(n435),.clk(gclk));
	jand g0364(.dina(w_n435_0[1]),.dinb(n431),.dout(n436),.clk(gclk));
	jor g0365(.dina(n436),.dinb(w_n168_2[0]),.dout(n437),.clk(gclk));
	jand g0366(.dina(n437),.dinb(w_n357_0[0]),.dout(n438),.clk(gclk));
	jand g0367(.dina(n438),.dinb(w_dff_B_HPDhHTvl3_1),.dout(n439),.clk(gclk));
	jor g0368(.dina(w_n439_0[2]),.dinb(w_G169_2[0]),.dout(n440),.clk(gclk));
	jand g0369(.dina(w_G33_7[1]),.dinb(w_n151_4[0]),.dout(n441),.clk(gclk));
	jand g0370(.dina(w_n441_0[1]),.dinb(w_G58_4[2]),.dout(n442),.clk(gclk));
	jnot g0371(.din(n442),.dout(n443),.clk(gclk));
	jor g0372(.dina(w_n77_0[0]),.dinb(w_n151_3[2]),.dout(n444),.clk(gclk));
	jand g0373(.dina(w_n153_5[2]),.dinb(w_n151_3[1]),.dout(n445),.clk(gclk));
	jand g0374(.dina(w_n445_0[1]),.dinb(w_G150_3[1]),.dout(n446),.clk(gclk));
	jnot g0375(.din(n446),.dout(n447),.clk(gclk));
	jand g0376(.dina(n447),.dinb(n444),.dout(n448),.clk(gclk));
	jand g0377(.dina(n448),.dinb(w_dff_B_OKK6X1Xx9_1),.dout(n449),.clk(gclk));
	jor g0378(.dina(n449),.dinb(w_n261_0[2]),.dout(n450),.clk(gclk));
	jnot g0379(.din(w_n450_0[1]),.dout(n451),.clk(gclk));
	jnot g0380(.din(w_n144_0[2]),.dout(n452),.clk(gclk));
	jand g0381(.dina(w_n452_0[1]),.dinb(w_n73_2[0]),.dout(n453),.clk(gclk));
	jnot g0382(.din(n453),.dout(n454),.clk(gclk));
	jor g0383(.dina(w_n414_0[1]),.dinb(w_n73_1[2]),.dout(n455),.clk(gclk));
	jand g0384(.dina(n455),.dinb(n454),.dout(n456),.clk(gclk));
	jor g0385(.dina(w_n456_0[1]),.dinb(n451),.dout(n457),.clk(gclk));
	jnot g0386(.din(w_n435_0[0]),.dout(n458),.clk(gclk));
	jor g0387(.dina(n458),.dinb(w_n430_0[0]),.dout(n459),.clk(gclk));
	jand g0388(.dina(n459),.dinb(w_n172_1[2]),.dout(n460),.clk(gclk));
	jor g0389(.dina(n460),.dinb(w_n356_0[2]),.dout(n461),.clk(gclk));
	jor g0390(.dina(n461),.dinb(w_n428_0[0]),.dout(n462),.clk(gclk));
	jor g0391(.dina(n462),.dinb(w_G179_2[0]),.dout(n463),.clk(gclk));
	jand g0392(.dina(n463),.dinb(w_n457_0[1]),.dout(n464),.clk(gclk));
	jand g0393(.dina(n464),.dinb(w_dff_B_gWM7VLxp7_1),.dout(n465),.clk(gclk));
	jand g0394(.dina(w_n439_0[1]),.dinb(w_G190_2[2]),.dout(n466),.clk(gclk));
	jnot g0395(.din(n466),.dout(n467),.clk(gclk));
	jnot g0396(.din(w_n456_0[0]),.dout(n468),.clk(gclk));
	jand g0397(.dina(n468),.dinb(w_n450_0[0]),.dout(n469),.clk(gclk));
	jor g0398(.dina(w_n439_0[0]),.dinb(w_n388_2[0]),.dout(n470),.clk(gclk));
	jand g0399(.dina(n470),.dinb(n469),.dout(n471),.clk(gclk));
	jand g0400(.dina(n471),.dinb(n467),.dout(n472),.clk(gclk));
	jor g0401(.dina(w_n472_0[1]),.dinb(w_n465_0[1]),.dout(n473),.clk(gclk));
	jand g0402(.dina(w_n168_1[2]),.dinb(w_G232_0[1]),.dout(n474),.clk(gclk));
	jand g0403(.dina(n474),.dinb(w_n354_0[1]),.dout(n475),.clk(gclk));
	jand g0404(.dina(w_n173_1[0]),.dinb(w_G226_0[1]),.dout(n476),.clk(gclk));
	jand g0405(.dina(w_n177_0[1]),.dinb(w_G223_0[0]),.dout(n477),.clk(gclk));
	jor g0406(.dina(n477),.dinb(w_n370_0[0]),.dout(n478),.clk(gclk));
	jor g0407(.dina(n478),.dinb(w_dff_B_G3EgqqmC4_1),.dout(n479),.clk(gclk));
	jand g0408(.dina(n479),.dinb(w_n172_1[1]),.dout(n480),.clk(gclk));
	jor g0409(.dina(n480),.dinb(w_n356_0[1]),.dout(n481),.clk(gclk));
	jor g0410(.dina(n481),.dinb(w_dff_B_uAVr2jzw7_1),.dout(n482),.clk(gclk));
	jnot g0411(.din(w_n482_0[2]),.dout(n483),.clk(gclk));
	jor g0412(.dina(w_n483_0[1]),.dinb(w_G169_1[2]),.dout(n484),.clk(gclk));
	jnot g0413(.din(w_G159_3[2]),.dout(n485),.clk(gclk));
	jnot g0414(.din(w_n445_0[0]),.dout(n486),.clk(gclk));
	jor g0415(.dina(n486),.dinb(w_dff_B_IOgjobww9_1),.dout(n487),.clk(gclk));
	jxor g0416(.dina(w_G68_4[1]),.dinb(w_G58_4[1]),.dout(n488),.clk(gclk));
	jor g0417(.dina(n488),.dinb(w_n151_3[0]),.dout(n489),.clk(gclk));
	jand g0418(.dina(w_n441_0[0]),.dinb(w_G68_4[0]),.dout(n490),.clk(gclk));
	jnot g0419(.din(n490),.dout(n491),.clk(gclk));
	jand g0420(.dina(n491),.dinb(w_dff_B_fPSynR9i2_1),.dout(n492),.clk(gclk));
	jand g0421(.dina(n492),.dinb(w_dff_B_eapyrZRK4_1),.dout(n493),.clk(gclk));
	jor g0422(.dina(n493),.dinb(w_n261_0[1]),.dout(n494),.clk(gclk));
	jnot g0423(.din(w_n494_0[1]),.dout(n495),.clk(gclk));
	jand g0424(.dina(w_n452_0[0]),.dinb(w_n74_1[2]),.dout(n496),.clk(gclk));
	jnot g0425(.din(n496),.dout(n497),.clk(gclk));
	jor g0426(.dina(w_n414_0[0]),.dinb(w_n74_1[1]),.dout(n498),.clk(gclk));
	jand g0427(.dina(n498),.dinb(n497),.dout(n499),.clk(gclk));
	jor g0428(.dina(w_n499_0[1]),.dinb(n495),.dout(n500),.clk(gclk));
	jor g0429(.dina(w_n482_0[1]),.dinb(w_G179_1[2]),.dout(n501),.clk(gclk));
	jand g0430(.dina(n501),.dinb(w_n500_0[1]),.dout(n502),.clk(gclk));
	jand g0431(.dina(n502),.dinb(n484),.dout(n503),.clk(gclk));
	jor g0432(.dina(w_n483_0[0]),.dinb(w_n388_1[2]),.dout(n504),.clk(gclk));
	jnot g0433(.din(w_n499_0[0]),.dout(n505),.clk(gclk));
	jand g0434(.dina(n505),.dinb(w_n494_0[0]),.dout(n506),.clk(gclk));
	jnot g0435(.din(w_G190_2[1]),.dout(n507),.clk(gclk));
	jor g0436(.dina(w_n482_0[0]),.dinb(w_n507_2[1]),.dout(n508),.clk(gclk));
	jand g0437(.dina(n508),.dinb(n506),.dout(n509),.clk(gclk));
	jand g0438(.dina(n509),.dinb(n504),.dout(n510),.clk(gclk));
	jor g0439(.dina(n510),.dinb(w_n503_0[2]),.dout(n511),.clk(gclk));
	jor g0440(.dina(w_n511_0[1]),.dinb(w_n473_0[1]),.dout(n512),.clk(gclk));
	jor g0441(.dina(w_n512_0[1]),.dinb(w_n426_0[1]),.dout(n513),.clk(gclk));
	jor g0442(.dina(n513),.dinb(w_n395_0[1]),.dout(n514),.clk(gclk));
	jnot g0443(.din(w_n514_1[1]),.dout(n515),.clk(gclk));
	jand g0444(.dina(n515),.dinb(w_n351_0[1]),.dout(w_dff_A_JAByGg7B5_2),.clk(gclk));
	jnot g0445(.din(w_n213_0[0]),.dout(n517),.clk(gclk));
	jor g0446(.dina(w_n212_0[2]),.dinb(w_G179_1[1]),.dout(n518),.clk(gclk));
	jand g0447(.dina(n518),.dinb(w_n224_0[2]),.dout(n519),.clk(gclk));
	jand g0448(.dina(n519),.dinb(n517),.dout(n520),.clk(gclk));
	jnot g0449(.din(w_n238_0[0]),.dout(n521),.clk(gclk));
	jor g0450(.dina(w_n234_0[2]),.dinb(w_n388_1[1]),.dout(n522),.clk(gclk));
	jand g0451(.dina(n522),.dinb(w_n225_0[0]),.dout(n523),.clk(gclk));
	jand g0452(.dina(n523),.dinb(n521),.dout(n524),.clk(gclk));
	jor g0453(.dina(n524),.dinb(w_n520_0[1]),.dout(n525),.clk(gclk));
	jnot g0454(.din(w_n256_0[0]),.dout(n526),.clk(gclk));
	jor g0455(.dina(w_n255_0[2]),.dinb(w_G169_1[1]),.dout(n527),.clk(gclk));
	jand g0456(.dina(n527),.dinb(w_n292_0[1]),.dout(n528),.clk(gclk));
	jand g0457(.dina(n528),.dinb(n526),.dout(n529),.clk(gclk));
	jnot g0458(.din(w_n283_0[0]),.dout(n530),.clk(gclk));
	jor g0459(.dina(w_n279_0[2]),.dinb(w_n507_2[0]),.dout(n531),.clk(gclk));
	jand g0460(.dina(n531),.dinb(w_n272_0[0]),.dout(n532),.clk(gclk));
	jand g0461(.dina(n532),.dinb(n530),.dout(n533),.clk(gclk));
	jor g0462(.dina(w_n533_0[1]),.dinb(n529),.dout(n534),.clk(gclk));
	jnot g0463(.din(w_n309_0[0]),.dout(n535),.clk(gclk));
	jor g0464(.dina(w_n308_0[2]),.dinb(w_n388_1[0]),.dout(n536),.clk(gclk));
	jand g0465(.dina(n536),.dinb(w_n344_0[0]),.dout(n537),.clk(gclk));
	jand g0466(.dina(n537),.dinb(n535),.dout(n538),.clk(gclk));
	jor g0467(.dina(w_n330_0[1]),.dinb(w_G179_1[0]),.dout(n539),.clk(gclk));
	jand g0468(.dina(n539),.dinb(w_n323_0[1]),.dout(n540),.clk(gclk));
	jand g0469(.dina(n540),.dinb(w_n334_0[0]),.dout(n541),.clk(gclk));
	jor g0470(.dina(w_n541_0[1]),.dinb(w_dff_B_azq4YLDP6_1),.dout(n542),.clk(gclk));
	jor g0471(.dina(w_n542_0[1]),.dinb(w_n534_0[1]),.dout(n543),.clk(gclk));
	jor g0472(.dina(w_n543_0[1]),.dinb(w_dff_B_OrLSHVmi8_1),.dout(n544),.clk(gclk));
	jor g0473(.dina(w_n544_0[1]),.dinb(w_n192_0[1]),.dout(n545),.clk(gclk));
	jor g0474(.dina(w_n543_0[0]),.dinb(w_n237_0[1]),.dout(n546),.clk(gclk));
	jor g0475(.dina(w_n347_0[0]),.dinb(w_n533_0[0]),.dout(n547),.clk(gclk));
	jand g0476(.dina(n547),.dinb(w_n282_0[0]),.dout(n548),.clk(gclk));
	jand g0477(.dina(w_n548_0[1]),.dinb(n546),.dout(n549),.clk(gclk));
	jand g0478(.dina(n549),.dinb(n545),.dout(n550),.clk(gclk));
	jor g0479(.dina(w_n550_0[1]),.dinb(w_n514_1[0]),.dout(n551),.clk(gclk));
	jnot g0480(.din(w_n551_0[1]),.dout(n552),.clk(gclk));
	jnot g0481(.din(w_n472_0[0]),.dout(n553),.clk(gclk));
	jand g0482(.dina(w_n503_0[1]),.dinb(n553),.dout(n554),.clk(gclk));
	jnot g0483(.din(n554),.dout(n555),.clk(gclk));
	jnot g0484(.din(w_n465_0[0]),.dout(n556),.clk(gclk));
	jnot g0485(.din(w_n420_0[0]),.dout(n557),.clk(gclk));
	jor g0486(.dina(w_n425_0[0]),.dinb(w_n387_0[1]),.dout(n558),.clk(gclk));
	jand g0487(.dina(n558),.dinb(w_dff_B_GHDibozC2_1),.dout(n559),.clk(gclk));
	jor g0488(.dina(w_n559_0[1]),.dinb(w_n512_0[0]),.dout(n560),.clk(gclk));
	jand g0489(.dina(n560),.dinb(w_dff_B_K3A7R6M86_1),.dout(n561),.clk(gclk));
	jand g0490(.dina(n561),.dinb(w_dff_B_a6D3DV1K1_1),.dout(n562),.clk(gclk));
	jnot g0491(.din(w_n562_0[1]),.dout(n563),.clk(gclk));
	jor g0492(.dina(n563),.dinb(n552),.dout(w_dff_A_qRdAfI1F8_2),.clk(gclk));
	jand g0493(.dina(w_n143_0[0]),.dinb(w_G213_0[2]),.dout(n565),.clk(gclk));
	jand g0494(.dina(n565),.dinb(w_n151_2[2]),.dout(n566),.clk(gclk));
	jand g0495(.dina(w_n566_1[1]),.dinb(w_G343_0[1]),.dout(n567),.clk(gclk));
	jor g0496(.dina(w_n567_5[1]),.dinb(w_n237_0[0]),.dout(n568),.clk(gclk));
	jnot g0497(.din(n568),.dout(n569),.clk(gclk));
	jnot g0498(.din(w_n192_0[0]),.dout(n570),.clk(gclk));
	jnot g0499(.din(w_n567_5[0]),.dout(n571),.clk(gclk));
	jand g0500(.dina(w_n571_2[1]),.dinb(w_n570_0[1]),.dout(n572),.clk(gclk));
	jand g0501(.dina(w_n572_0[2]),.dinb(w_n242_0[1]),.dout(n573),.clk(gclk));
	jor g0502(.dina(w_n573_0[1]),.dinb(w_n569_0[1]),.dout(n574),.clk(gclk));
	jand g0503(.dina(w_n567_4[2]),.dinb(w_n161_0[0]),.dout(n575),.clk(gclk));
	jxor g0504(.dina(w_dff_B_jvbrpiFg4_0),.dinb(w_n198_0[1]),.dout(n576),.clk(gclk));
	jand g0505(.dina(w_n576_0[2]),.dinb(w_G330_0[2]),.dout(n577),.clk(gclk));
	jand g0506(.dina(w_n567_4[1]),.dinb(w_n224_0[1]),.dout(n578),.clk(gclk));
	jxor g0507(.dina(w_dff_B_YHsPo9ub3_0),.dinb(w_n242_0[0]),.dout(n579),.clk(gclk));
	jand g0508(.dina(w_n579_1[1]),.dinb(w_n577_0[1]),.dout(n580),.clk(gclk));
	jor g0509(.dina(w_n580_0[2]),.dinb(w_n574_0[1]),.dout(w_dff_A_UHzT0RaE1_2),.clk(gclk));
	jand g0510(.dina(w_n91_1[1]),.dinb(w_n163_0[2]),.dout(n582),.clk(gclk));
	jand g0511(.dina(w_n582_0[1]),.dinb(w_n118_0[1]),.dout(n583),.clk(gclk));
	jor g0512(.dina(w_n567_4[0]),.dinb(w_n550_0[0]),.dout(n584),.clk(gclk));
	jnot g0513(.din(w_n198_0[0]),.dout(n585),.clk(gclk));
	jor g0514(.dina(w_n544_0[0]),.dinb(n585),.dout(n586),.clk(gclk));
	jand g0515(.dina(w_n571_2[0]),.dinb(n586),.dout(n587),.clk(gclk));
	jnot g0516(.din(w_n190_0[0]),.dout(n588),.clk(gclk));
	jand g0517(.dina(w_n308_0[1]),.dinb(w_n255_0[1]),.dout(n589),.clk(gclk));
	jand g0518(.dina(w_dff_B_rBoAC2sS8_0),.dinb(n588),.dout(n590),.clk(gclk));
	jand g0519(.dina(n590),.dinb(w_n234_0[1]),.dout(n591),.clk(gclk));
	jand g0520(.dina(w_n279_0[1]),.dinb(w_n189_1[0]),.dout(n592),.clk(gclk));
	jand g0521(.dina(n592),.dinb(w_n330_0[0]),.dout(n593),.clk(gclk));
	jand g0522(.dina(n593),.dinb(w_n186_0[1]),.dout(n594),.clk(gclk));
	jand g0523(.dina(n594),.dinb(w_n212_0[1]),.dout(n595),.clk(gclk));
	jor g0524(.dina(n595),.dinb(w_n571_1[2]),.dout(n596),.clk(gclk));
	jor g0525(.dina(n596),.dinb(n591),.dout(n597),.clk(gclk));
	jand g0526(.dina(n597),.dinb(w_G330_0[1]),.dout(n598),.clk(gclk));
	jnot g0527(.din(w_n598_0[1]),.dout(n599),.clk(gclk));
	jor g0528(.dina(w_dff_B_STIrPms96_0),.dinb(n587),.dout(n600),.clk(gclk));
	jand g0529(.dina(w_n600_1[2]),.dinb(w_n584_0[1]),.dout(n601),.clk(gclk));
	jnot g0530(.din(w_n601_0[2]),.dout(n602),.clk(gclk));
	jand g0531(.dina(w_n602_0[1]),.dinb(w_n142_1[0]),.dout(n603),.clk(gclk));
	jnot g0532(.din(w_n582_0[0]),.dout(n604),.clk(gclk));
	jand g0533(.dina(w_n259_0[0]),.dinb(w_n105_0[2]),.dout(n605),.clk(gclk));
	jand g0534(.dina(w_n605_0[2]),.dinb(w_G1_0[2]),.dout(n606),.clk(gclk));
	jand g0535(.dina(n606),.dinb(w_n604_2[2]),.dout(n607),.clk(gclk));
	jor g0536(.dina(w_dff_B_mOPif1fF3_0),.dinb(n603),.dout(n608),.clk(gclk));
	jor g0537(.dina(n608),.dinb(w_dff_B_prADZb7W6_1),.dout(w_dff_A_PHITdRC31_2),.clk(gclk));
	jand g0538(.dina(w_G45_0[2]),.dinb(w_G13_0[2]),.dout(n610),.clk(gclk));
	jand g0539(.dina(n610),.dinb(w_n151_2[1]),.dout(n611),.clk(gclk));
	jor g0540(.dina(n611),.dinb(w_n142_0[2]),.dout(n612),.clk(gclk));
	jnot g0541(.din(n612),.dout(n613),.clk(gclk));
	jand g0542(.dina(w_n613_1[2]),.dinb(w_n604_2[1]),.dout(n614),.clk(gclk));
	jnot g0543(.din(w_n614_5[1]),.dout(n615),.clk(gclk));
	jxor g0544(.dina(w_n576_0[1]),.dinb(w_G330_0[0]),.dout(n616),.clk(gclk));
	jand g0545(.dina(n616),.dinb(w_dff_B_q8k9MOuf7_1),.dout(n617),.clk(gclk));
	jand g0546(.dina(w_n153_5[1]),.dinb(w_n89_0[0]),.dout(n618),.clk(gclk));
	jand g0547(.dina(w_n618_2[1]),.dinb(w_n151_2[0]),.dout(n619),.clk(gclk));
	jnot g0548(.din(w_n619_0[2]),.dout(n620),.clk(gclk));
	jor g0549(.dina(w_n620_0[2]),.dinb(w_n576_0[0]),.dout(n621),.clk(gclk));
	jand g0550(.dina(w_n507_1[2]),.dinb(w_G20_2[2]),.dout(n622),.clk(gclk));
	jnot g0551(.din(w_n622_0[1]),.dout(n623),.clk(gclk));
	jand g0552(.dina(w_G200_1[1]),.dinb(w_G20_2[1]),.dout(n624),.clk(gclk));
	jnot g0553(.din(w_n624_0[1]),.dout(n625),.clk(gclk));
	jand g0554(.dina(w_G179_0[2]),.dinb(w_G20_2[0]),.dout(n626),.clk(gclk));
	jnot g0555(.din(w_n626_0[2]),.dout(n627),.clk(gclk));
	jand g0556(.dina(n627),.dinb(n625),.dout(n628),.clk(gclk));
	jand g0557(.dina(w_n628_0[1]),.dinb(n623),.dout(n629),.clk(gclk));
	jand g0558(.dina(w_n629_5[1]),.dinb(w_G97_3[0]),.dout(n630),.clk(gclk));
	jnot g0559(.din(w_n630_0[1]),.dout(n631),.clk(gclk));
	jand g0560(.dina(w_n624_0[0]),.dinb(w_n189_0[2]),.dout(n632),.clk(gclk));
	jand g0561(.dina(w_n632_0[1]),.dinb(w_G190_2[0]),.dout(n633),.clk(gclk));
	jand g0562(.dina(w_n633_6[1]),.dinb(w_G87_2[1]),.dout(n634),.clk(gclk));
	jnot g0563(.din(w_n634_0[1]),.dout(n635),.clk(gclk));
	jand g0564(.dina(w_dff_B_HSexzlMl6_0),.dinb(n631),.dout(n636),.clk(gclk));
	jand g0565(.dina(w_n626_0[1]),.dinb(w_n388_0[2]),.dout(n637),.clk(gclk));
	jand g0566(.dina(w_n637_0[1]),.dinb(w_n507_1[1]),.dout(n638),.clk(gclk));
	jand g0567(.dina(w_n638_7[1]),.dinb(w_G77_3[0]),.dout(n639),.clk(gclk));
	jand g0568(.dina(w_n628_0[0]),.dinb(w_n622_0[0]),.dout(n640),.clk(gclk));
	jand g0569(.dina(w_n640_7[1]),.dinb(w_G159_3[1]),.dout(n641),.clk(gclk));
	jor g0570(.dina(n641),.dinb(w_dff_B_cTi4cvda5_1),.dout(n642),.clk(gclk));
	jor g0571(.dina(n642),.dinb(w_G33_7[0]),.dout(n643),.clk(gclk));
	jnot g0572(.din(n643),.dout(n644),.clk(gclk));
	jand g0573(.dina(n644),.dinb(w_dff_B_cx0kmtJb8_1),.dout(n645),.clk(gclk));
	jand g0574(.dina(w_n637_0[0]),.dinb(w_G190_1[2]),.dout(n646),.clk(gclk));
	jand g0575(.dina(w_n646_7[1]),.dinb(w_G58_4[0]),.dout(n647),.clk(gclk));
	jand g0576(.dina(w_n632_0[0]),.dinb(w_n507_1[0]),.dout(n648),.clk(gclk));
	jand g0577(.dina(w_n648_4[1]),.dinb(w_G107_3[0]),.dout(n649),.clk(gclk));
	jand g0578(.dina(w_n626_0[0]),.dinb(w_G200_1[0]),.dout(n650),.clk(gclk));
	jand g0579(.dina(w_n650_0[1]),.dinb(w_G190_1[1]),.dout(n651),.clk(gclk));
	jand g0580(.dina(w_n651_7[1]),.dinb(w_G50_4[1]),.dout(n652),.clk(gclk));
	jand g0581(.dina(w_n650_0[0]),.dinb(w_n507_0[2]),.dout(n653),.clk(gclk));
	jand g0582(.dina(w_n653_7[1]),.dinb(w_G68_3[2]),.dout(n654),.clk(gclk));
	jor g0583(.dina(n654),.dinb(n652),.dout(n655),.clk(gclk));
	jor g0584(.dina(n655),.dinb(w_n649_0[1]),.dout(n656),.clk(gclk));
	jor g0585(.dina(n656),.dinb(w_dff_B_WwaOHHlo8_1),.dout(n657),.clk(gclk));
	jnot g0586(.din(n657),.dout(n658),.clk(gclk));
	jand g0587(.dina(w_dff_B_XZYEa8my8_0),.dinb(n645),.dout(n659),.clk(gclk));
	jnot g0588(.din(n659),.dout(n660),.clk(gclk));
	jand g0589(.dina(w_n646_7[0]),.dinb(w_G322_0[2]),.dout(n661),.clk(gclk));
	jand g0590(.dina(w_n633_6[0]),.dinb(w_G303_2[1]),.dout(n662),.clk(gclk));
	jand g0591(.dina(w_n629_5[0]),.dinb(w_G294_3[0]),.dout(n663),.clk(gclk));
	jor g0592(.dina(n663),.dinb(w_dff_B_MdHqP3XU9_1),.dout(n664),.clk(gclk));
	jand g0593(.dina(w_n651_7[0]),.dinb(w_G326_0[1]),.dout(n665),.clk(gclk));
	jor g0594(.dina(w_dff_B_Xa6NuVoZ9_0),.dinb(n664),.dout(n666),.clk(gclk));
	jand g0595(.dina(w_n640_7[0]),.dinb(w_dff_B_U5SKTSDO0_1),.dout(n667),.clk(gclk));
	jor g0596(.dina(n667),.dinb(w_n153_5[0]),.dout(n668),.clk(gclk));
	jand g0597(.dina(w_n638_7[0]),.dinb(w_G311_1[2]),.dout(n669),.clk(gclk));
	jand g0598(.dina(w_n653_7[0]),.dinb(w_G317_1[1]),.dout(n670),.clk(gclk));
	jor g0599(.dina(n670),.dinb(n669),.dout(n671),.clk(gclk));
	jand g0600(.dina(w_n648_4[0]),.dinb(w_G283_3[1]),.dout(n672),.clk(gclk));
	jor g0601(.dina(w_dff_B_PGB7mGTc7_0),.dinb(n671),.dout(n673),.clk(gclk));
	jor g0602(.dina(n673),.dinb(n668),.dout(n674),.clk(gclk));
	jor g0603(.dina(n674),.dinb(n666),.dout(n675),.clk(gclk));
	jor g0604(.dina(n675),.dinb(w_dff_B_2WX1sdRp1_1),.dout(n676),.clk(gclk));
	jand g0605(.dina(w_dff_B_IPXw9dON6_0),.dinb(n660),.dout(n677),.clk(gclk));
	jand g0606(.dina(w_n139_0[1]),.dinb(w_G169_1[0]),.dout(n678),.clk(gclk));
	jor g0607(.dina(n678),.dinb(w_n375_0[0]),.dout(n679),.clk(gclk));
	jnot g0608(.din(n679),.dout(n680),.clk(gclk));
	jor g0609(.dina(w_n680_4[1]),.dinb(n677),.dout(n681),.clk(gclk));
	jand g0610(.dina(w_n680_4[0]),.dinb(w_n620_0[1]),.dout(n682),.clk(gclk));
	jor g0611(.dina(w_n134_0[0]),.dinb(w_n352_1[0]),.dout(n683),.clk(gclk));
	jand g0612(.dina(w_n91_1[0]),.dinb(w_G33_6[2]),.dout(n684),.clk(gclk));
	jnot g0613(.din(w_n684_0[2]),.dout(n685),.clk(gclk));
	jand g0614(.dina(w_n118_0[0]),.dinb(w_n352_0[2]),.dout(n686),.clk(gclk));
	jor g0615(.dina(n686),.dinb(w_n685_0[1]),.dout(n687),.clk(gclk));
	jnot g0616(.din(n687),.dout(n688),.clk(gclk));
	jand g0617(.dina(n688),.dinb(w_dff_B_zs0to0HM6_1),.dout(n689),.clk(gclk));
	jnot g0618(.din(w_n91_0[2]),.dout(n690),.clk(gclk));
	jand g0619(.dina(w_n690_1[1]),.dinb(w_n105_0[1]),.dout(n691),.clk(gclk));
	jand g0620(.dina(w_n91_0[1]),.dinb(w_n153_4[2]),.dout(n692),.clk(gclk));
	jand g0621(.dina(w_n692_0[1]),.dinb(w_G355_0),.dout(n693),.clk(gclk));
	jor g0622(.dina(n693),.dinb(n691),.dout(n694),.clk(gclk));
	jor g0623(.dina(w_dff_B_2uiw1TE68_0),.dinb(n689),.dout(n695),.clk(gclk));
	jand g0624(.dina(n695),.dinb(w_n682_0[1]),.dout(n696),.clk(gclk));
	jnot g0625(.din(n696),.dout(n697),.clk(gclk));
	jand g0626(.dina(w_dff_B_eIU6FKJH2_0),.dinb(n681),.dout(n698),.clk(gclk));
	jand g0627(.dina(w_dff_B_3KsAx5iO0_0),.dinb(n621),.dout(n699),.clk(gclk));
	jand g0628(.dina(n699),.dinb(w_n614_5[0]),.dout(n700),.clk(gclk));
	jor g0629(.dina(n700),.dinb(w_dff_B_7dexFQRr4_1),.dout(G396_fa_),.clk(gclk));
	jand g0630(.dina(w_n567_3[2]),.dinb(w_n383_0[0]),.dout(n702),.clk(gclk));
	jxor g0631(.dina(w_dff_B_LzxIiMpc8_0),.dinb(w_n394_0[0]),.dout(n703),.clk(gclk));
	jnot g0632(.din(w_n703_1[1]),.dout(n704),.clk(gclk));
	jand g0633(.dina(w_n704_0[1]),.dinb(w_n618_2[0]),.dout(n705),.clk(gclk));
	jnot g0634(.din(n705),.dout(n706),.clk(gclk));
	jand g0635(.dina(w_n653_6[2]),.dinb(w_G150_3[0]),.dout(n707),.clk(gclk));
	jand g0636(.dina(w_n651_6[2]),.dinb(w_G137_1[2]),.dout(n708),.clk(gclk));
	jand g0637(.dina(w_n633_5[2]),.dinb(w_G50_4[0]),.dout(n709),.clk(gclk));
	jor g0638(.dina(n709),.dinb(n708),.dout(n710),.clk(gclk));
	jand g0639(.dina(w_n646_6[2]),.dinb(w_G143_2[1]),.dout(n711),.clk(gclk));
	jor g0640(.dina(w_dff_B_0YsiHeIC6_0),.dinb(n710),.dout(n712),.clk(gclk));
	jor g0641(.dina(n712),.dinb(w_dff_B_CsOHDHJM3_1),.dout(n713),.clk(gclk));
	jand g0642(.dina(w_n638_6[2]),.dinb(w_G159_3[0]),.dout(n714),.clk(gclk));
	jand g0643(.dina(w_n640_6[2]),.dinb(w_G132_1[1]),.dout(n715),.clk(gclk));
	jor g0644(.dina(n715),.dinb(w_dff_B_l3j8OZvY8_1),.dout(n716),.clk(gclk));
	jand g0645(.dina(w_n629_4[2]),.dinb(w_G58_3[2]),.dout(n717),.clk(gclk));
	jand g0646(.dina(w_n648_3[2]),.dinb(w_G68_3[1]),.dout(n718),.clk(gclk));
	jor g0647(.dina(w_n718_0[1]),.dinb(n717),.dout(n719),.clk(gclk));
	jor g0648(.dina(n719),.dinb(w_G33_6[1]),.dout(n720),.clk(gclk));
	jor g0649(.dina(n720),.dinb(w_dff_B_LPi0uogA1_1),.dout(n721),.clk(gclk));
	jor g0650(.dina(n721),.dinb(w_dff_B_oCrH7Lgx0_1),.dout(n722),.clk(gclk));
	jand g0651(.dina(w_n653_6[1]),.dinb(w_G283_3[0]),.dout(n723),.clk(gclk));
	jand g0652(.dina(w_n640_6[1]),.dinb(w_G311_1[1]),.dout(n724),.clk(gclk));
	jor g0653(.dina(n724),.dinb(w_dff_B_Qgk1zIAq1_1),.dout(n725),.clk(gclk));
	jand g0654(.dina(w_n633_5[1]),.dinb(w_G107_2[2]),.dout(n726),.clk(gclk));
	jor g0655(.dina(w_dff_B_c4JQbR9H5_0),.dinb(w_n630_0[0]),.dout(n727),.clk(gclk));
	jor g0656(.dina(n727),.dinb(n725),.dout(n728),.clk(gclk));
	jand g0657(.dina(w_n646_6[1]),.dinb(w_G294_2[2]),.dout(n729),.clk(gclk));
	jand g0658(.dina(w_n638_6[1]),.dinb(w_G116_4[0]),.dout(n730),.clk(gclk));
	jor g0659(.dina(n730),.dinb(n729),.dout(n731),.clk(gclk));
	jand g0660(.dina(w_n651_6[1]),.dinb(w_G303_2[0]),.dout(n732),.clk(gclk));
	jand g0661(.dina(w_n648_3[1]),.dinb(w_G87_2[0]),.dout(n733),.clk(gclk));
	jor g0662(.dina(w_n733_0[1]),.dinb(n732),.dout(n734),.clk(gclk));
	jor g0663(.dina(n734),.dinb(n731),.dout(n735),.clk(gclk));
	jor g0664(.dina(w_dff_B_OhgEfmRx3_0),.dinb(n728),.dout(n736),.clk(gclk));
	jor g0665(.dina(n736),.dinb(w_n153_4[1]),.dout(n737),.clk(gclk));
	jand g0666(.dina(n737),.dinb(n722),.dout(n738),.clk(gclk));
	jor g0667(.dina(n738),.dinb(w_n680_3[2]),.dout(n739),.clk(gclk));
	jnot g0668(.din(w_n618_1[2]),.dout(n740),.clk(gclk));
	jand g0669(.dina(w_n680_3[1]),.dinb(w_dff_B_QeiMDT8I5_1),.dout(n741),.clk(gclk));
	jand g0670(.dina(w_n741_1[1]),.dinb(w_n72_0[1]),.dout(n742),.clk(gclk));
	jnot g0671(.din(n742),.dout(n743),.clk(gclk));
	jand g0672(.dina(w_dff_B_vaDBoLY89_0),.dinb(n739),.dout(n744),.clk(gclk));
	jand g0673(.dina(n744),.dinb(w_n614_4[2]),.dout(n745),.clk(gclk));
	jand g0674(.dina(w_dff_B_iNYb9PqW3_0),.dinb(n706),.dout(n746),.clk(gclk));
	jnot g0675(.din(n746),.dout(n747),.clk(gclk));
	jor g0676(.dina(w_n584_0[0]),.dinb(w_n395_0[0]),.dout(n748),.clk(gclk));
	jand g0677(.dina(w_n350_0[0]),.dinb(w_n570_0[0]),.dout(n749),.clk(gclk));
	jand g0678(.dina(w_n349_0[0]),.dinb(w_n520_0[0]),.dout(n750),.clk(gclk));
	jnot g0679(.din(w_n548_0[0]),.dout(n751),.clk(gclk));
	jor g0680(.dina(w_dff_B_UcjOiyLY9_0),.dinb(n750),.dout(n752),.clk(gclk));
	jor g0681(.dina(n752),.dinb(n749),.dout(n753),.clk(gclk));
	jand g0682(.dina(w_n571_1[1]),.dinb(n753),.dout(n754),.clk(gclk));
	jor g0683(.dina(w_n703_1[0]),.dinb(w_n754_0[1]),.dout(n755),.clk(gclk));
	jand g0684(.dina(n755),.dinb(w_n748_0[1]),.dout(n756),.clk(gclk));
	jxor g0685(.dina(n756),.dinb(w_n600_1[1]),.dout(n757),.clk(gclk));
	jor g0686(.dina(n757),.dinb(w_n614_4[1]),.dout(n758),.clk(gclk));
	jand g0687(.dina(n758),.dinb(w_dff_B_WE9fOSRN4_1),.dout(n759),.clk(gclk));
	jnot g0688(.din(w_n759_0[1]),.dout(G384_fa_),.clk(gclk));
	jnot g0689(.din(w_n90_0[1]),.dout(n761),.clk(gclk));
	jand g0690(.dina(w_n112_0[0]),.dinb(n761),.dout(n762),.clk(gclk));
	jnot g0691(.din(w_n566_1[0]),.dout(n763),.clk(gclk));
	jand g0692(.dina(w_dff_B_uxtRcIsy7_0),.dinb(w_n503_0[0]),.dout(n764),.clk(gclk));
	jand g0693(.dina(w_n566_0[2]),.dinb(w_n500_0[0]),.dout(n765),.clk(gclk));
	jxor g0694(.dina(w_dff_B_pgpnDPot6_0),.dinb(w_n511_0[0]),.dout(n766),.clk(gclk));
	jnot g0695(.din(w_n766_0[1]),.dout(n767),.clk(gclk));
	jor g0696(.dina(w_n567_3[1]),.dinb(w_n559_0[0]),.dout(n768),.clk(gclk));
	jnot g0697(.din(n768),.dout(n769),.clk(gclk));
	jand g0698(.dina(w_n567_3[0]),.dinb(w_n417_0[0]),.dout(n770),.clk(gclk));
	jxor g0699(.dina(w_dff_B_hQIfFVma4_0),.dinb(w_n426_0[0]),.dout(n771),.clk(gclk));
	jnot g0700(.din(w_n771_1[1]),.dout(n772),.clk(gclk));
	jand g0701(.dina(w_n772_0[1]),.dinb(w_n703_0[2]),.dout(n773),.clk(gclk));
	jand g0702(.dina(w_n773_0[1]),.dinb(w_n754_0[0]),.dout(n774),.clk(gclk));
	jor g0703(.dina(n774),.dinb(w_dff_B_ED5gFEA37_1),.dout(n775),.clk(gclk));
	jand g0704(.dina(w_n775_0[1]),.dinb(w_n767_1[1]),.dout(n776),.clk(gclk));
	jor g0705(.dina(n776),.dinb(w_dff_B_4HRWX6FB9_1),.dout(n777),.clk(gclk));
	jand g0706(.dina(w_n773_0[0]),.dinb(w_n767_1[0]),.dout(n778),.clk(gclk));
	jxor g0707(.dina(n778),.dinb(w_n514_0[2]),.dout(n779),.clk(gclk));
	jor g0708(.dina(n779),.dinb(w_n600_1[0]),.dout(n780),.clk(gclk));
	jor g0709(.dina(w_n567_2[2]),.dinb(w_n551_0[0]),.dout(n781),.clk(gclk));
	jand g0710(.dina(n781),.dinb(w_n562_0[0]),.dout(n782),.clk(gclk));
	jxor g0711(.dina(w_n782_0[1]),.dinb(n780),.dout(n783),.clk(gclk));
	jxor g0712(.dina(w_dff_B_NNpb1PAP1_0),.dinb(w_n777_0[1]),.dout(n784),.clk(gclk));
	jand g0713(.dina(n784),.dinb(w_dff_B_mirvIYcZ8_1),.dout(n785),.clk(gclk));
	jor g0714(.dina(w_n75_1[0]),.dinb(w_n74_1[0]),.dout(n786),.clk(gclk));
	jand g0715(.dina(n786),.dinb(w_G77_2[2]),.dout(n787),.clk(gclk));
	jor g0716(.dina(n787),.dinb(w_n73_1[1]),.dout(n788),.clk(gclk));
	jand g0717(.dina(w_G58_3[1]),.dinb(w_G50_3[2]),.dout(n789),.clk(gclk));
	jor g0718(.dina(n789),.dinb(w_G68_3[0]),.dout(n790),.clk(gclk));
	jand g0719(.dina(n790),.dinb(w_n90_0[0]),.dout(n791),.clk(gclk));
	jand g0720(.dina(w_dff_B_AVjPnWhX9_0),.dinb(n788),.dout(n792),.clk(gclk));
	jand g0721(.dina(w_n312_0[0]),.dinb(w_n120_0[0]),.dout(n793),.clk(gclk));
	jand g0722(.dina(n793),.dinb(w_G116_3[2]),.dout(n794),.clk(gclk));
	jor g0723(.dina(w_dff_B_sq671Pcx0_0),.dinb(n792),.dout(n795),.clk(gclk));
	jor g0724(.dina(w_dff_B_eyzArHIQ3_0),.dinb(n785),.dout(w_dff_A_s1BWpEPJ7_2),.clk(gclk));
	jand g0725(.dina(w_n567_2[1]),.dinb(w_n292_0[0]),.dout(n797),.clk(gclk));
	jxor g0726(.dina(w_dff_B_n68jINf37_0),.dinb(w_n534_0[0]),.dout(n798),.clk(gclk));
	jand g0727(.dina(w_n798_0[1]),.dinb(w_n619_0[1]),.dout(n799),.clk(gclk));
	jnot g0728(.din(n799),.dout(n800),.clk(gclk));
	jand g0729(.dina(w_n684_0[1]),.dinb(w_n126_0[0]),.dout(n801),.clk(gclk));
	jnot g0730(.din(w_n682_0[0]),.dout(n802),.clk(gclk));
	jand g0731(.dina(w_n690_1[0]),.dinb(w_G87_1[2]),.dout(n803),.clk(gclk));
	jor g0732(.dina(w_dff_B_jHdHPdUh9_0),.dinb(w_n802_0[2]),.dout(n804),.clk(gclk));
	jor g0733(.dina(n804),.dinb(w_dff_B_9kC6cd7E5_1),.dout(n805),.clk(gclk));
	jand g0734(.dina(n805),.dinb(w_n614_4[0]),.dout(n806),.clk(gclk));
	jand g0735(.dina(w_n646_6[0]),.dinb(w_G303_1[2]),.dout(n807),.clk(gclk));
	jand g0736(.dina(w_n638_6[0]),.dinb(w_G283_2[2]),.dout(n808),.clk(gclk));
	jor g0737(.dina(n808),.dinb(n807),.dout(n809),.clk(gclk));
	jand g0738(.dina(w_n651_6[0]),.dinb(w_G311_1[0]),.dout(n810),.clk(gclk));
	jand g0739(.dina(w_n633_5[0]),.dinb(w_G116_3[1]),.dout(n811),.clk(gclk));
	jor g0740(.dina(n811),.dinb(n810),.dout(n812),.clk(gclk));
	jand g0741(.dina(w_n653_6[0]),.dinb(w_G294_2[1]),.dout(n813),.clk(gclk));
	jand g0742(.dina(w_n640_6[0]),.dinb(w_G317_1[0]),.dout(n814),.clk(gclk));
	jor g0743(.dina(n814),.dinb(w_dff_B_ORF3evCs4_1),.dout(n815),.clk(gclk));
	jand g0744(.dina(w_n629_4[1]),.dinb(w_G107_2[1]),.dout(n816),.clk(gclk));
	jand g0745(.dina(w_n648_3[0]),.dinb(w_G97_2[2]),.dout(n817),.clk(gclk));
	jor g0746(.dina(w_n817_0[1]),.dinb(n816),.dout(n818),.clk(gclk));
	jor g0747(.dina(n818),.dinb(n815),.dout(n819),.clk(gclk));
	jor g0748(.dina(n819),.dinb(w_dff_B_IcFqzFcb4_1),.dout(n820),.clk(gclk));
	jor g0749(.dina(n820),.dinb(w_dff_B_ITBo9cRh8_1),.dout(n821),.clk(gclk));
	jand g0750(.dina(n821),.dinb(w_G33_6[0]),.dout(n822),.clk(gclk));
	jand g0751(.dina(w_n638_5[2]),.dinb(w_G50_3[1]),.dout(n823),.clk(gclk));
	jand g0752(.dina(w_n640_5[2]),.dinb(w_G137_1[1]),.dout(n824),.clk(gclk));
	jor g0753(.dina(n824),.dinb(w_dff_B_J4G9mpnt1_1),.dout(n825),.clk(gclk));
	jand g0754(.dina(w_n651_5[2]),.dinb(w_G143_2[0]),.dout(n826),.clk(gclk));
	jand g0755(.dina(w_n653_5[2]),.dinb(w_G159_2[2]),.dout(n827),.clk(gclk));
	jor g0756(.dina(n827),.dinb(n826),.dout(n828),.clk(gclk));
	jand g0757(.dina(w_n633_4[2]),.dinb(w_G58_3[0]),.dout(n829),.clk(gclk));
	jand g0758(.dina(w_n629_4[0]),.dinb(w_G68_2[2]),.dout(n830),.clk(gclk));
	jor g0759(.dina(w_n830_0[1]),.dinb(w_dff_B_xumulVta2_1),.dout(n831),.clk(gclk));
	jand g0760(.dina(w_n646_5[2]),.dinb(w_G150_2[2]),.dout(n832),.clk(gclk));
	jand g0761(.dina(w_n648_2[2]),.dinb(w_G77_2[1]),.dout(n833),.clk(gclk));
	jor g0762(.dina(w_n833_0[1]),.dinb(n832),.dout(n834),.clk(gclk));
	jor g0763(.dina(w_dff_B_evK5ALlS6_0),.dinb(n831),.dout(n835),.clk(gclk));
	jor g0764(.dina(n835),.dinb(w_dff_B_RxJFYEeT9_1),.dout(n836),.clk(gclk));
	jor g0765(.dina(n836),.dinb(w_dff_B_PwACYx4m9_1),.dout(n837),.clk(gclk));
	jand g0766(.dina(n837),.dinb(w_n153_4[0]),.dout(n838),.clk(gclk));
	jor g0767(.dina(n838),.dinb(n822),.dout(n839),.clk(gclk));
	jor g0768(.dina(n839),.dinb(w_n680_3[0]),.dout(n840),.clk(gclk));
	jand g0769(.dina(n840),.dinb(w_dff_B_tbPUkQaw0_1),.dout(n841),.clk(gclk));
	jand g0770(.dina(w_dff_B_reR9chzK7_0),.dinb(n800),.dout(n842),.clk(gclk));
	jnot g0771(.din(n842),.dout(n843),.clk(gclk));
	jand g0772(.dina(w_n567_2[0]),.dinb(w_n323_0[0]),.dout(n844),.clk(gclk));
	jxor g0773(.dina(w_dff_B_JiavlIFh1_0),.dinb(w_n542_0[0]),.dout(n845),.clk(gclk));
	jnot g0774(.din(w_n845_0[2]),.dout(n846),.clk(gclk));
	jand g0775(.dina(w_dff_B_olPxfAgE5_0),.dinb(w_n580_0[1]),.dout(n847),.clk(gclk));
	jand g0776(.dina(w_n571_1[0]),.dinb(w_n541_0[0]),.dout(n848),.clk(gclk));
	jand g0777(.dina(w_n579_1[0]),.dinb(w_n348_0[0]),.dout(n849),.clk(gclk));
	jand g0778(.dina(n849),.dinb(w_n572_0[1]),.dout(n850),.clk(gclk));
	jand g0779(.dina(w_n569_0[0]),.dinb(w_n333_0[0]),.dout(n851),.clk(gclk));
	jor g0780(.dina(w_dff_B_drb9tgyI3_0),.dinb(n850),.dout(n852),.clk(gclk));
	jor g0781(.dina(n852),.dinb(w_dff_B_ZAfep1yA9_1),.dout(n853),.clk(gclk));
	jxor g0782(.dina(n853),.dinb(w_n798_0[0]),.dout(n854),.clk(gclk));
	jxor g0783(.dina(n854),.dinb(w_dff_B_YAk8KxDc6_1),.dout(n855),.clk(gclk));
	jor g0784(.dina(w_n855_0[1]),.dinb(w_n613_1[1]),.dout(n856),.clk(gclk));
	jnot g0785(.din(w_n573_0[0]),.dout(n857),.clk(gclk));
	jor g0786(.dina(w_n579_0[2]),.dinb(w_n572_0[0]),.dout(n858),.clk(gclk));
	jand g0787(.dina(w_dff_B_Fsh1G4pF3_0),.dinb(n857),.dout(n859),.clk(gclk));
	jxor g0788(.dina(n859),.dinb(w_n577_0[0]),.dout(n860),.clk(gclk));
	jnot g0789(.din(w_n860_0[1]),.dout(n861),.clk(gclk));
	jxor g0790(.dina(w_n580_0[0]),.dinb(w_n574_0[0]),.dout(n862),.clk(gclk));
	jxor g0791(.dina(n862),.dinb(w_n845_0[1]),.dout(n863),.clk(gclk));
	jor g0792(.dina(w_n863_0[2]),.dinb(w_n861_0[1]),.dout(n864),.clk(gclk));
	jand g0793(.dina(n864),.dinb(w_n601_0[1]),.dout(n865),.clk(gclk));
	jor g0794(.dina(w_n855_0[0]),.dinb(w_n604_2[0]),.dout(n866),.clk(gclk));
	jor g0795(.dina(w_dff_B_2qZ3BbhQ9_0),.dinb(n865),.dout(n867),.clk(gclk));
	jand g0796(.dina(n867),.dinb(w_dff_B_EYZKU5ko9_1),.dout(n868),.clk(gclk));
	jand g0797(.dina(n868),.dinb(w_dff_B_vSBWEpvC8_1),.dout(n869),.clk(gclk));
	jnot g0798(.din(w_n869_0[2]),.dout(w_dff_A_9T1uPaDL7_1),.clk(gclk));
	jor g0799(.dina(w_n602_0[0]),.dinb(w_n604_1[2]),.dout(n871),.clk(gclk));
	jand g0800(.dina(n871),.dinb(w_n861_0[0]),.dout(n872),.clk(gclk));
	jand g0801(.dina(w_n860_0[0]),.dinb(w_n601_0[0]),.dout(n873),.clk(gclk));
	jand g0802(.dina(w_n873_0[1]),.dinb(w_n613_1[0]),.dout(n874),.clk(gclk));
	jor g0803(.dina(n874),.dinb(w_n614_3[2]),.dout(n875),.clk(gclk));
	jor g0804(.dina(w_n875_0[1]),.dinb(n872),.dout(n876),.clk(gclk));
	jor g0805(.dina(w_n620_0[0]),.dinb(w_n579_0[1]),.dout(n877),.clk(gclk));
	jand g0806(.dina(w_n653_5[1]),.dinb(w_G58_2[2]),.dout(n878),.clk(gclk));
	jand g0807(.dina(w_n638_5[1]),.dinb(w_G68_2[1]),.dout(n879),.clk(gclk));
	jor g0808(.dina(n879),.dinb(w_n817_0[0]),.dout(n880),.clk(gclk));
	jor g0809(.dina(n880),.dinb(w_G33_5[2]),.dout(n881),.clk(gclk));
	jor g0810(.dina(n881),.dinb(w_dff_B_8Vywqy5C4_1),.dout(n882),.clk(gclk));
	jnot g0811(.din(n882),.dout(n883),.clk(gclk));
	jand g0812(.dina(w_n629_3[2]),.dinb(w_G87_1[1]),.dout(n884),.clk(gclk));
	jnot g0813(.din(w_n884_0[1]),.dout(n885),.clk(gclk));
	jand g0814(.dina(w_n633_4[1]),.dinb(w_G77_2[0]),.dout(n886),.clk(gclk));
	jnot g0815(.din(n886),.dout(n887),.clk(gclk));
	jand g0816(.dina(w_n887_0[1]),.dinb(n885),.dout(n888),.clk(gclk));
	jand g0817(.dina(w_n646_5[1]),.dinb(w_G50_3[0]),.dout(n889),.clk(gclk));
	jand g0818(.dina(w_n640_5[1]),.dinb(w_G150_2[1]),.dout(n890),.clk(gclk));
	jor g0819(.dina(n890),.dinb(w_dff_B_RwoL5VWu8_1),.dout(n891),.clk(gclk));
	jand g0820(.dina(w_n651_5[1]),.dinb(w_G159_2[1]),.dout(n892),.clk(gclk));
	jor g0821(.dina(w_dff_B_v9iNmF707_0),.dinb(n891),.dout(n893),.clk(gclk));
	jnot g0822(.din(n893),.dout(n894),.clk(gclk));
	jand g0823(.dina(n894),.dinb(w_dff_B_h4qqhYoZ3_1),.dout(n895),.clk(gclk));
	jand g0824(.dina(n895),.dinb(w_dff_B_PERCOOkK4_1),.dout(n896),.clk(gclk));
	jnot g0825(.din(n896),.dout(n897),.clk(gclk));
	jand g0826(.dina(w_n653_5[0]),.dinb(w_G311_0[2]),.dout(n898),.clk(gclk));
	jand g0827(.dina(w_n633_4[0]),.dinb(w_G294_2[0]),.dout(n899),.clk(gclk));
	jand g0828(.dina(w_n629_3[1]),.dinb(w_G283_2[1]),.dout(n900),.clk(gclk));
	jor g0829(.dina(n900),.dinb(w_dff_B_uJOhXaQ34_1),.dout(n901),.clk(gclk));
	jand g0830(.dina(w_n651_5[0]),.dinb(w_G322_0[1]),.dout(n902),.clk(gclk));
	jand g0831(.dina(w_n640_5[0]),.dinb(w_G326_0[0]),.dout(n903),.clk(gclk));
	jor g0832(.dina(n903),.dinb(w_dff_B_ITkbkyJf1_1),.dout(n904),.clk(gclk));
	jor g0833(.dina(n904),.dinb(n901),.dout(n905),.clk(gclk));
	jand g0834(.dina(w_n638_5[0]),.dinb(w_G303_1[1]),.dout(n906),.clk(gclk));
	jand g0835(.dina(w_n648_2[1]),.dinb(w_G116_3[0]),.dout(n907),.clk(gclk));
	jor g0836(.dina(n907),.dinb(n906),.dout(n908),.clk(gclk));
	jand g0837(.dina(w_n646_5[0]),.dinb(w_G317_0[2]),.dout(n909),.clk(gclk));
	jor g0838(.dina(w_dff_B_USA1XYU61_0),.dinb(n908),.dout(n910),.clk(gclk));
	jor g0839(.dina(n910),.dinb(w_n153_3[2]),.dout(n911),.clk(gclk));
	jor g0840(.dina(n911),.dinb(n905),.dout(n912),.clk(gclk));
	jor g0841(.dina(n912),.dinb(w_dff_B_gNEDBGez0_1),.dout(n913),.clk(gclk));
	jand g0842(.dina(w_dff_B_mJyPI1ZB7_0),.dinb(n897),.dout(n914),.clk(gclk));
	jor g0843(.dina(n914),.dinb(w_n680_2[2]),.dout(n915),.clk(gclk));
	jand g0844(.dina(w_n690_0[2]),.dinb(w_n81_0[2]),.dout(n916),.clk(gclk));
	jnot g0845(.din(n916),.dout(n917),.clk(gclk));
	jnot g0846(.din(w_n605_0[1]),.dout(n918),.clk(gclk));
	jand g0847(.dina(w_n692_0[0]),.dinb(n918),.dout(n919),.clk(gclk));
	jnot g0848(.din(n919),.dout(n920),.clk(gclk));
	jand g0849(.dina(w_n130_0[0]),.dinb(w_G45_0[1]),.dout(n921),.clk(gclk));
	jor g0850(.dina(w_dff_B_Q4nvGl6c1_0),.dinb(w_n685_0[0]),.dout(n922),.clk(gclk));
	jand g0851(.dina(w_dff_B_6MfxNJ1F1_0),.dinb(n920),.dout(n923),.clk(gclk));
	jand g0852(.dina(w_G77_1[2]),.dinb(w_G68_2[0]),.dout(n924),.clk(gclk));
	jnot g0853(.din(n924),.dout(n925),.clk(gclk));
	jand g0854(.dina(w_G58_2[1]),.dinb(w_n73_1[0]),.dout(n926),.clk(gclk));
	jand g0855(.dina(n926),.dinb(n925),.dout(n927),.clk(gclk));
	jand g0856(.dina(w_dff_B_7ESZrZng0_0),.dinb(w_n605_0[0]),.dout(n928),.clk(gclk));
	jand g0857(.dina(n928),.dinb(w_n352_0[1]),.dout(n929),.clk(gclk));
	jor g0858(.dina(w_dff_B_KdZ70WhS7_0),.dinb(n923),.dout(n930),.clk(gclk));
	jand g0859(.dina(n930),.dinb(w_dff_B_BNt8wNsu8_1),.dout(n931),.clk(gclk));
	jor g0860(.dina(n931),.dinb(w_n802_0[1]),.dout(n932),.clk(gclk));
	jand g0861(.dina(w_dff_B_t2YV5ulg4_0),.dinb(n915),.dout(n933),.clk(gclk));
	jand g0862(.dina(n933),.dinb(n877),.dout(n934),.clk(gclk));
	jand g0863(.dina(n934),.dinb(w_n614_3[1]),.dout(n935),.clk(gclk));
	jnot g0864(.din(n935),.dout(n936),.clk(gclk));
	jand g0865(.dina(w_dff_B_jlxAK9nM9_0),.dinb(n876),.dout(n937),.clk(gclk));
	jnot g0866(.din(w_n937_0[2]),.dout(w_dff_A_AxGVX6TL1_1),.clk(gclk));
	jnot g0867(.din(w_n863_0[1]),.dout(n939),.clk(gclk));
	jnot g0868(.din(w_n873_0[0]),.dout(n940),.clk(gclk));
	jor g0869(.dina(n940),.dinb(w_dff_B_bmkZyDxZ1_1),.dout(n941),.clk(gclk));
	jor g0870(.dina(n941),.dinb(w_n604_1[1]),.dout(n942),.clk(gclk));
	jor g0871(.dina(w_n875_0[0]),.dinb(w_n863_0[0]),.dout(n943),.clk(gclk));
	jand g0872(.dina(w_n845_0[0]),.dinb(w_n619_0[0]),.dout(n944),.clk(gclk));
	jnot g0873(.din(n944),.dout(n945),.clk(gclk));
	jand g0874(.dina(w_n690_0[1]),.dinb(w_G97_2[1]),.dout(n946),.clk(gclk));
	jand g0875(.dina(w_n684_0[0]),.dinb(w_n137_0[0]),.dout(n947),.clk(gclk));
	jor g0876(.dina(w_dff_B_AwPZqyvy3_0),.dinb(w_n802_0[0]),.dout(n948),.clk(gclk));
	jor g0877(.dina(n948),.dinb(w_dff_B_LY7bYntw8_1),.dout(n949),.clk(gclk));
	jand g0878(.dina(w_n653_4[2]),.dinb(w_G50_2[2]),.dout(n950),.clk(gclk));
	jand g0879(.dina(w_n638_4[2]),.dinb(w_G58_2[0]),.dout(n951),.clk(gclk));
	jor g0880(.dina(n951),.dinb(n950),.dout(n952),.clk(gclk));
	jand g0881(.dina(w_n646_4[2]),.dinb(w_G159_2[0]),.dout(n953),.clk(gclk));
	jand g0882(.dina(w_n633_3[2]),.dinb(w_G68_1[2]),.dout(n954),.clk(gclk));
	jor g0883(.dina(n954),.dinb(n953),.dout(n955),.clk(gclk));
	jand g0884(.dina(w_n651_4[2]),.dinb(w_G150_2[0]),.dout(n956),.clk(gclk));
	jor g0885(.dina(n956),.dinb(w_n733_0[0]),.dout(n957),.clk(gclk));
	jand g0886(.dina(w_n640_4[2]),.dinb(w_G143_1[2]),.dout(n958),.clk(gclk));
	jand g0887(.dina(w_n629_3[0]),.dinb(w_G77_1[1]),.dout(n959),.clk(gclk));
	jor g0888(.dina(w_n959_0[1]),.dinb(n958),.dout(n960),.clk(gclk));
	jor g0889(.dina(n960),.dinb(w_dff_B_3538W6Se4_1),.dout(n961),.clk(gclk));
	jor g0890(.dina(n961),.dinb(w_dff_B_yRAbqoPj3_1),.dout(n962),.clk(gclk));
	jor g0891(.dina(n962),.dinb(w_dff_B_2fzj4tTD7_1),.dout(n963),.clk(gclk));
	jand g0892(.dina(n963),.dinb(w_n153_3[1]),.dout(n964),.clk(gclk));
	jand g0893(.dina(w_n638_4[1]),.dinb(w_G294_1[2]),.dout(n965),.clk(gclk));
	jand g0894(.dina(w_n640_4[1]),.dinb(w_G322_0[0]),.dout(n966),.clk(gclk));
	jor g0895(.dina(n966),.dinb(w_dff_B_QGb6dHNc8_1),.dout(n967),.clk(gclk));
	jand g0896(.dina(w_n646_4[1]),.dinb(w_G311_0[1]),.dout(n968),.clk(gclk));
	jand g0897(.dina(w_n651_4[1]),.dinb(w_G317_0[1]),.dout(n969),.clk(gclk));
	jor g0898(.dina(n969),.dinb(n968),.dout(n970),.clk(gclk));
	jand g0899(.dina(w_n653_4[1]),.dinb(w_G303_1[0]),.dout(n971),.clk(gclk));
	jor g0900(.dina(n971),.dinb(w_n649_0[0]),.dout(n972),.clk(gclk));
	jor g0901(.dina(n972),.dinb(n970),.dout(n973),.clk(gclk));
	jand g0902(.dina(w_n633_3[1]),.dinb(w_G283_2[0]),.dout(n974),.clk(gclk));
	jand g0903(.dina(w_n629_2[2]),.dinb(w_G116_2[2]),.dout(n975),.clk(gclk));
	jor g0904(.dina(n975),.dinb(w_dff_B_Y3pctb3y9_1),.dout(n976),.clk(gclk));
	jor g0905(.dina(n976),.dinb(n973),.dout(n977),.clk(gclk));
	jor g0906(.dina(n977),.dinb(w_dff_B_7whsfyG25_1),.dout(n978),.clk(gclk));
	jand g0907(.dina(n978),.dinb(w_G33_5[1]),.dout(n979),.clk(gclk));
	jor g0908(.dina(n979),.dinb(w_n680_2[1]),.dout(n980),.clk(gclk));
	jor g0909(.dina(n980),.dinb(n964),.dout(n981),.clk(gclk));
	jand g0910(.dina(n981),.dinb(w_n614_3[0]),.dout(n982),.clk(gclk));
	jand g0911(.dina(n982),.dinb(w_dff_B_7g4tZBYO7_1),.dout(n983),.clk(gclk));
	jand g0912(.dina(w_dff_B_Og2VNfOO6_0),.dinb(n945),.dout(n984),.clk(gclk));
	jnot g0913(.din(n984),.dout(n985),.clk(gclk));
	jand g0914(.dina(w_dff_B_JC0CyPB34_0),.dinb(n943),.dout(n986),.clk(gclk));
	jand g0915(.dina(n986),.dinb(w_dff_B_76G1R80I7_1),.dout(n987),.clk(gclk));
	jnot g0916(.din(w_n987_0[2]),.dout(w_dff_A_4z7A7QZb0_1),.clk(gclk));
	jand g0917(.dina(w_n766_0[0]),.dinb(w_n618_1[1]),.dout(n989),.clk(gclk));
	jnot g0918(.din(n989),.dout(n990),.clk(gclk));
	jand g0919(.dina(w_n651_4[0]),.dinb(w_G128_0[2]),.dout(n991),.clk(gclk));
	jand g0920(.dina(w_n640_4[0]),.dinb(w_G125_0[1]),.dout(n992),.clk(gclk));
	jor g0921(.dina(n992),.dinb(w_dff_B_MemRcEoA6_1),.dout(n993),.clk(gclk));
	jand g0922(.dina(w_n648_2[0]),.dinb(w_G50_2[1]),.dout(n994),.clk(gclk));
	jand g0923(.dina(w_n653_4[0]),.dinb(w_G137_1[0]),.dout(n995),.clk(gclk));
	jor g0924(.dina(n995),.dinb(n994),.dout(n996),.clk(gclk));
	jor g0925(.dina(n996),.dinb(w_G33_5[0]),.dout(n997),.clk(gclk));
	jor g0926(.dina(n997),.dinb(n993),.dout(n998),.clk(gclk));
	jand g0927(.dina(w_n638_4[0]),.dinb(w_G143_1[1]),.dout(n999),.clk(gclk));
	jand g0928(.dina(w_n633_3[0]),.dinb(w_G150_1[2]),.dout(n1000),.clk(gclk));
	jand g0929(.dina(w_n629_2[1]),.dinb(w_G159_1[2]),.dout(n1001),.clk(gclk));
	jand g0930(.dina(w_n646_4[0]),.dinb(w_G132_1[0]),.dout(n1002),.clk(gclk));
	jor g0931(.dina(w_dff_B_qpyT6lIT2_0),.dinb(n1001),.dout(n1003),.clk(gclk));
	jor g0932(.dina(n1003),.dinb(w_dff_B_mpEZYCdW1_1),.dout(n1004),.clk(gclk));
	jor g0933(.dina(n1004),.dinb(w_dff_B_8UkSvFVL7_1),.dout(n1005),.clk(gclk));
	jor g0934(.dina(n1005),.dinb(w_dff_B_CkUcccqP4_1),.dout(n1006),.clk(gclk));
	jand g0935(.dina(w_n651_3[2]),.dinb(w_G283_1[2]),.dout(n1007),.clk(gclk));
	jand g0936(.dina(w_n638_3[2]),.dinb(w_G97_2[0]),.dout(n1008),.clk(gclk));
	jor g0937(.dina(n1008),.dinb(w_n153_3[0]),.dout(n1009),.clk(gclk));
	jor g0938(.dina(n1009),.dinb(w_dff_B_CLm81odN6_1),.dout(n1010),.clk(gclk));
	jand g0939(.dina(w_n646_3[2]),.dinb(w_G116_2[1]),.dout(n1011),.clk(gclk));
	jand g0940(.dina(w_n640_3[2]),.dinb(w_G294_1[1]),.dout(n1012),.clk(gclk));
	jor g0941(.dina(n1012),.dinb(w_dff_B_Jp6T2fN52_1),.dout(n1013),.clk(gclk));
	jand g0942(.dina(w_n653_3[2]),.dinb(w_G107_2[0]),.dout(n1014),.clk(gclk));
	jor g0943(.dina(n1014),.dinb(w_n634_0[0]),.dout(n1015),.clk(gclk));
	jor g0944(.dina(w_dff_B_AaXitViX9_0),.dinb(n1013),.dout(n1016),.clk(gclk));
	jor g0945(.dina(n1016),.dinb(w_dff_B_8gPGC0Fu6_1),.dout(n1017),.clk(gclk));
	jor g0946(.dina(n1017),.dinb(w_n959_0[0]),.dout(n1018),.clk(gclk));
	jor g0947(.dina(n1018),.dinb(w_n718_0[0]),.dout(n1019),.clk(gclk));
	jand g0948(.dina(n1019),.dinb(w_dff_B_m88xIWPw1_1),.dout(n1020),.clk(gclk));
	jor g0949(.dina(n1020),.dinb(w_n680_2[0]),.dout(n1021),.clk(gclk));
	jand g0950(.dina(w_n741_1[0]),.dinb(w_n74_0[2]),.dout(n1022),.clk(gclk));
	jnot g0951(.din(n1022),.dout(n1023),.clk(gclk));
	jand g0952(.dina(w_dff_B_QKTeOl1e3_0),.dinb(n1021),.dout(n1024),.clk(gclk));
	jand g0953(.dina(n1024),.dinb(w_n614_2[2]),.dout(n1025),.clk(gclk));
	jand g0954(.dina(w_dff_B_B2gUorcj5_0),.dinb(n990),.dout(n1026),.clk(gclk));
	jnot g0955(.din(n1026),.dout(n1027),.clk(gclk));
	jor g0956(.dina(w_n600_0[2]),.dinb(w_n514_0[1]),.dout(n1028),.clk(gclk));
	jand g0957(.dina(w_dff_B_zOWbBvLs7_0),.dinb(w_n782_0[0]),.dout(n1029),.clk(gclk));
	jnot g0958(.din(w_n387_0[0]),.dout(n1030),.clk(gclk));
	jand g0959(.dina(w_n571_0[2]),.dinb(n1030),.dout(n1031),.clk(gclk));
	jnot g0960(.din(n1031),.dout(n1032),.clk(gclk));
	jand g0961(.dina(w_dff_B_Uz0lf2br0_0),.dinb(w_n748_0[0]),.dout(n1033),.clk(gclk));
	jor g0962(.dina(w_n567_1[2]),.dinb(w_n351_0[0]),.dout(n1034),.clk(gclk));
	jand g0963(.dina(w_n598_0[0]),.dinb(n1034),.dout(n1035),.clk(gclk));
	jand g0964(.dina(w_n703_0[1]),.dinb(n1035),.dout(n1036),.clk(gclk));
	jxor g0965(.dina(w_n1036_0[1]),.dinb(w_n771_1[0]),.dout(n1037),.clk(gclk));
	jxor g0966(.dina(n1037),.dinb(w_n1033_0[1]),.dout(n1038),.clk(gclk));
	jand g0967(.dina(n1038),.dinb(w_n1029_0[2]),.dout(n1039),.clk(gclk));
	jor g0968(.dina(w_n1039_0[1]),.dinb(w_n604_1[0]),.dout(n1040),.clk(gclk));
	jand g0969(.dina(w_n1040_0[1]),.dinb(w_n613_0[2]),.dout(n1041),.clk(gclk));
	jor g0970(.dina(w_n704_0[0]),.dinb(w_n600_0[1]),.dout(n1042),.clk(gclk));
	jor g0971(.dina(n1042),.dinb(w_n771_0[2]),.dout(n1043),.clk(gclk));
	jxor g0972(.dina(w_n775_0[0]),.dinb(w_n767_0[2]),.dout(n1044),.clk(gclk));
	jxor g0973(.dina(w_n1044_0[1]),.dinb(w_n1043_0[1]),.dout(n1045),.clk(gclk));
	jor g0974(.dina(w_n1045_0[1]),.dinb(w_n1041_0[1]),.dout(n1046),.clk(gclk));
	jnot g0975(.din(w_n1039_0[0]),.dout(n1047),.clk(gclk));
	jnot g0976(.din(w_n1043_0[0]),.dout(n1048),.clk(gclk));
	jxor g0977(.dina(w_n1044_0[0]),.dinb(w_n1048_0[1]),.dout(n1049),.clk(gclk));
	jor g0978(.dina(n1049),.dinb(w_n604_0[2]),.dout(n1050),.clk(gclk));
	jor g0979(.dina(n1050),.dinb(n1047),.dout(n1051),.clk(gclk));
	jand g0980(.dina(w_dff_B_1N7T31AP7_0),.dinb(n1046),.dout(n1052),.clk(gclk));
	jand g0981(.dina(n1052),.dinb(w_dff_B_4uF57oCj4_1),.dout(n1053),.clk(gclk));
	jnot g0982(.din(w_n1053_0[2]),.dout(w_dff_A_lKt9RnS31_1),.clk(gclk));
	jxor g0983(.dina(w_n1036_0[0]),.dinb(w_n772_0[0]),.dout(n1055),.clk(gclk));
	jxor g0984(.dina(n1055),.dinb(w_n1033_0[0]),.dout(n1056),.clk(gclk));
	jor g0985(.dina(w_n1045_0[0]),.dinb(w_n1056_0[1]),.dout(n1057),.clk(gclk));
	jand g0986(.dina(w_n1029_0[1]),.dinb(w_n613_0[1]),.dout(n1058),.clk(gclk));
	jand g0987(.dina(w_dff_B_XZ06BLZb3_0),.dinb(n1057),.dout(n1059),.clk(gclk));
	jand g0988(.dina(w_n1048_0[0]),.dinb(w_n767_0[1]),.dout(n1060),.clk(gclk));
	jand g0989(.dina(w_n566_0[1]),.dinb(w_n457_0[0]),.dout(n1061),.clk(gclk));
	jxor g0990(.dina(w_dff_B_QnLRwrnw8_0),.dinb(w_n473_0[0]),.dout(n1062),.clk(gclk));
	jxor g0991(.dina(w_n1062_0[1]),.dinb(w_n777_0[0]),.dout(n1063),.clk(gclk));
	jxor g0992(.dina(n1063),.dinb(w_dff_B_jIOqZmB33_1),.dout(n1064),.clk(gclk));
	jor g0993(.dina(n1064),.dinb(n1059),.dout(n1065),.clk(gclk));
	jor g0994(.dina(n1065),.dinb(w_n614_2[1]),.dout(n1066),.clk(gclk));
	jand g0995(.dina(w_n1062_0[0]),.dinb(w_n618_1[0]),.dout(n1067),.clk(gclk));
	jnot g0996(.din(n1067),.dout(n1068),.clk(gclk));
	jand g0997(.dina(w_G50_2[0]),.dinb(w_G41_0[0]),.dout(n1069),.clk(gclk));
	jor g0998(.dina(w_dff_B_dIaU5zlH8_0),.dinb(w_n680_1[2]),.dout(n1070),.clk(gclk));
	jand g0999(.dina(w_n638_3[1]),.dinb(w_G137_0[2]),.dout(n1071),.clk(gclk));
	jand g1000(.dina(w_n633_2[2]),.dinb(w_G143_1[0]),.dout(n1072),.clk(gclk));
	jand g1001(.dina(w_n651_3[1]),.dinb(w_G125_0[0]),.dout(n1073),.clk(gclk));
	jor g1002(.dina(n1073),.dinb(n1072),.dout(n1074),.clk(gclk));
	jor g1003(.dina(n1074),.dinb(w_dff_B_dfAUOGxt2_1),.dout(n1075),.clk(gclk));
	jand g1004(.dina(w_n640_3[1]),.dinb(w_dff_B_C7SLVvkC7_1),.dout(n1076),.clk(gclk));
	jand g1005(.dina(w_n629_2[0]),.dinb(w_G150_1[1]),.dout(n1077),.clk(gclk));
	jand g1006(.dina(w_n646_3[1]),.dinb(w_G128_0[1]),.dout(n1078),.clk(gclk));
	jor g1007(.dina(w_dff_B_TdsIXP264_0),.dinb(n1077),.dout(n1079),.clk(gclk));
	jor g1008(.dina(n1079),.dinb(w_dff_B_q2JofDlD2_1),.dout(n1080),.clk(gclk));
	jand g1009(.dina(w_n648_1[2]),.dinb(w_G159_1[1]),.dout(n1081),.clk(gclk));
	jand g1010(.dina(w_n653_3[1]),.dinb(w_G132_0[2]),.dout(n1082),.clk(gclk));
	jor g1011(.dina(n1082),.dinb(n1081),.dout(n1083),.clk(gclk));
	jor g1012(.dina(n1083),.dinb(w_G33_4[2]),.dout(n1084),.clk(gclk));
	jor g1013(.dina(w_dff_B_SRmOgYXh7_0),.dinb(n1080),.dout(n1085),.clk(gclk));
	jor g1014(.dina(n1085),.dinb(w_dff_B_seMa3UNg8_1),.dout(n1086),.clk(gclk));
	jand g1015(.dina(w_n653_3[0]),.dinb(w_G97_1[2]),.dout(n1087),.clk(gclk));
	jand g1016(.dina(w_n646_3[0]),.dinb(w_G107_1[2]),.dout(n1088),.clk(gclk));
	jor g1017(.dina(n1088),.dinb(n1087),.dout(n1089),.clk(gclk));
	jnot g1018(.din(n1089),.dout(n1090),.clk(gclk));
	jand g1019(.dina(w_n648_1[1]),.dinb(w_G58_1[2]),.dout(n1091),.clk(gclk));
	jnot g1020(.din(w_n1091_0[1]),.dout(n1092),.clk(gclk));
	jand g1021(.dina(n1092),.dinb(w_n887_0[0]),.dout(n1093),.clk(gclk));
	jand g1022(.dina(n1093),.dinb(n1090),.dout(n1094),.clk(gclk));
	jand g1023(.dina(w_n640_3[0]),.dinb(w_G283_1[1]),.dout(n1095),.clk(gclk));
	jor g1024(.dina(n1095),.dinb(w_n830_0[0]),.dout(n1096),.clk(gclk));
	jand g1025(.dina(w_n651_3[0]),.dinb(w_G116_2[0]),.dout(n1097),.clk(gclk));
	jand g1026(.dina(w_n638_3[0]),.dinb(w_G87_1[0]),.dout(n1098),.clk(gclk));
	jor g1027(.dina(n1098),.dinb(n1097),.dout(n1099),.clk(gclk));
	jor g1028(.dina(w_dff_B_vIG23IUk8_0),.dinb(n1096),.dout(n1100),.clk(gclk));
	jnot g1029(.din(n1100),.dout(n1101),.clk(gclk));
	jand g1030(.dina(n1101),.dinb(w_dff_B_6p2TD6t02_1),.dout(n1102),.clk(gclk));
	jand g1031(.dina(n1102),.dinb(w_G33_4[1]),.dout(n1103),.clk(gclk));
	jnot g1032(.din(n1103),.dout(n1104),.clk(gclk));
	jand g1033(.dina(n1104),.dinb(w_dff_B_UcePQ7nO9_1),.dout(n1105),.clk(gclk));
	jand g1034(.dina(n1105),.dinb(w_n163_0[1]),.dout(n1106),.clk(gclk));
	jor g1035(.dina(n1106),.dinb(w_dff_B_jY1lzMXy0_1),.dout(n1107),.clk(gclk));
	jand g1036(.dina(w_n741_0[2]),.dinb(w_n73_0[2]),.dout(n1108),.clk(gclk));
	jnot g1037(.din(n1108),.dout(n1109),.clk(gclk));
	jand g1038(.dina(w_dff_B_LpNv12ZK0_0),.dinb(n1107),.dout(n1110),.clk(gclk));
	jand g1039(.dina(n1110),.dinb(n1068),.dout(n1111),.clk(gclk));
	jand g1040(.dina(n1111),.dinb(w_n614_2[0]),.dout(n1112),.clk(gclk));
	jnot g1041(.din(n1112),.dout(n1113),.clk(gclk));
	jand g1042(.dina(w_dff_B_yX29Iaal8_0),.dinb(n1066),.dout(n1114),.clk(gclk));
	jnot g1043(.din(w_n1114_0[2]),.dout(w_dff_A_1rpzyvbw3_1),.clk(gclk));
	jand g1044(.dina(w_n771_0[1]),.dinb(w_n618_0[2]),.dout(n1116),.clk(gclk));
	jnot g1045(.din(n1116),.dout(n1117),.clk(gclk));
	jand g1046(.dina(w_n646_2[2]),.dinb(w_G283_1[0]),.dout(n1118),.clk(gclk));
	jand g1047(.dina(w_n633_2[1]),.dinb(w_G97_1[1]),.dout(n1119),.clk(gclk));
	jand g1048(.dina(w_n653_2[2]),.dinb(w_G116_1[2]),.dout(n1120),.clk(gclk));
	jor g1049(.dina(n1120),.dinb(n1119),.dout(n1121),.clk(gclk));
	jand g1050(.dina(w_n640_2[2]),.dinb(w_G303_0[2]),.dout(n1122),.clk(gclk));
	jor g1051(.dina(n1122),.dinb(n1121),.dout(n1123),.clk(gclk));
	jor g1052(.dina(n1123),.dinb(w_dff_B_JxhsXLS99_1),.dout(n1124),.clk(gclk));
	jor g1053(.dina(w_n884_0[0]),.dinb(w_n833_0[0]),.dout(n1125),.clk(gclk));
	jand g1054(.dina(w_n651_2[2]),.dinb(w_G294_1[0]),.dout(n1126),.clk(gclk));
	jand g1055(.dina(w_n638_2[2]),.dinb(w_G107_1[1]),.dout(n1127),.clk(gclk));
	jor g1056(.dina(n1127),.dinb(n1126),.dout(n1128),.clk(gclk));
	jor g1057(.dina(n1128),.dinb(w_n153_2[2]),.dout(n1129),.clk(gclk));
	jor g1058(.dina(n1129),.dinb(n1125),.dout(n1130),.clk(gclk));
	jor g1059(.dina(n1130),.dinb(n1124),.dout(n1131),.clk(gclk));
	jand g1060(.dina(w_n646_2[1]),.dinb(w_G137_0[1]),.dout(n1132),.clk(gclk));
	jand g1061(.dina(w_n633_2[0]),.dinb(w_G159_1[0]),.dout(n1133),.clk(gclk));
	jand g1062(.dina(w_n638_2[1]),.dinb(w_G150_1[0]),.dout(n1134),.clk(gclk));
	jor g1063(.dina(n1134),.dinb(n1133),.dout(n1135),.clk(gclk));
	jand g1064(.dina(w_n651_2[1]),.dinb(w_G132_0[1]),.dout(n1136),.clk(gclk));
	jand g1065(.dina(w_n629_1[2]),.dinb(w_G50_1[2]),.dout(n1137),.clk(gclk));
	jor g1066(.dina(n1137),.dinb(w_n1091_0[0]),.dout(n1138),.clk(gclk));
	jor g1067(.dina(n1138),.dinb(w_dff_B_JeNg2Ljz2_1),.dout(n1139),.clk(gclk));
	jand g1068(.dina(w_n653_2[1]),.dinb(w_G143_0[2]),.dout(n1140),.clk(gclk));
	jand g1069(.dina(w_n640_2[1]),.dinb(w_G128_0[0]),.dout(n1141),.clk(gclk));
	jor g1070(.dina(n1141),.dinb(w_dff_B_KZ9JUhvf0_1),.dout(n1142),.clk(gclk));
	jor g1071(.dina(n1142),.dinb(w_G33_4[0]),.dout(n1143),.clk(gclk));
	jor g1072(.dina(n1143),.dinb(n1139),.dout(n1144),.clk(gclk));
	jor g1073(.dina(n1144),.dinb(w_dff_B_PXEpW0aS6_1),.dout(n1145),.clk(gclk));
	jor g1074(.dina(n1145),.dinb(w_dff_B_OckltRcT2_1),.dout(n1146),.clk(gclk));
	jand g1075(.dina(n1146),.dinb(w_dff_B_UeGz7vFO4_1),.dout(n1147),.clk(gclk));
	jor g1076(.dina(n1147),.dinb(w_n680_1[1]),.dout(n1148),.clk(gclk));
	jand g1077(.dina(w_n741_0[1]),.dinb(w_n75_0[2]),.dout(n1149),.clk(gclk));
	jnot g1078(.din(n1149),.dout(n1150),.clk(gclk));
	jand g1079(.dina(w_dff_B_Alqur92y5_0),.dinb(n1148),.dout(n1151),.clk(gclk));
	jand g1080(.dina(w_dff_B_pgnI3aQB0_0),.dinb(n1117),.dout(n1152),.clk(gclk));
	jand g1081(.dina(n1152),.dinb(w_n614_1[2]),.dout(n1153),.clk(gclk));
	jnot g1082(.din(n1153),.dout(n1154),.clk(gclk));
	jor g1083(.dina(w_n1041_0[0]),.dinb(w_n1056_0[0]),.dout(n1155),.clk(gclk));
	jnot g1084(.din(w_n1029_0[0]),.dout(n1156),.clk(gclk));
	jor g1085(.dina(w_n1040_0[0]),.dinb(w_dff_B_wko8F1q72_1),.dout(n1157),.clk(gclk));
	jand g1086(.dina(w_dff_B_DuplOqxG0_0),.dinb(n1155),.dout(n1158),.clk(gclk));
	jand g1087(.dina(n1158),.dinb(w_dff_B_aPConhyT7_1),.dout(n1159),.clk(gclk));
	jnot g1088(.din(w_n1159_0[2]),.dout(w_dff_A_ZFDj4KzA8_1),.clk(gclk));
	jand g1089(.dina(w_n1114_0[1]),.dinb(w_n1053_0[1]),.dout(n1161),.clk(gclk));
	jand g1090(.dina(w_n1159_0[1]),.dinb(w_n759_0[0]),.dout(n1162),.clk(gclk));
	jand g1091(.dina(w_n987_0[1]),.dinb(w_n869_0[1]),.dout(n1163),.clk(gclk));
	jnot g1092(.din(w_G396_0),.dout(n1164),.clk(gclk));
	jand g1093(.dina(w_n937_0[1]),.dinb(w_n1164_0[1]),.dout(n1165),.clk(gclk));
	jand g1094(.dina(w_dff_B_HSI4VBVl1_0),.dinb(n1163),.dout(n1166),.clk(gclk));
	jand g1095(.dina(w_dff_B_NZyNgzld3_0),.dinb(n1162),.dout(n1167),.clk(gclk));
	jand g1096(.dina(n1167),.dinb(w_n1161_0[1]),.dout(n1168),.clk(gclk));
	jnot g1097(.din(w_n1168_0[1]),.dout(w_dff_A_U9Dhhxdh2_1),.clk(gclk));
	jnot g1098(.din(w_G343_0[0]),.dout(n1170),.clk(gclk));
	jand g1099(.dina(w_n1161_0[0]),.dinb(w_n1170_0[1]),.dout(n1171),.clk(gclk));
	jnot g1100(.din(w_G213_0[1]),.dout(n1172),.clk(gclk));
	jor g1101(.dina(w_n1168_0[0]),.dinb(w_dff_B_jy3F7UiK7_1),.dout(n1173),.clk(gclk));
	jor g1102(.dina(n1173),.dinb(w_dff_B_pLHv3hyp7_1),.dout(G409),.clk(gclk));
	jxor g1103(.dina(w_n937_0[0]),.dinb(w_n1164_0[0]),.dout(n1175),.clk(gclk));
	jxor g1104(.dina(w_n987_0[0]),.dinb(w_n869_0[0]),.dout(n1176),.clk(gclk));
	jxor g1105(.dina(n1176),.dinb(w_dff_B_cRQ7BKJr4_1),.dout(n1177),.clk(gclk));
	jand g1106(.dina(w_n1170_0[0]),.dinb(w_G213_0[0]),.dout(n1178),.clk(gclk));
	jxor g1107(.dina(w_n1159_0[0]),.dinb(w_G384_0),.dout(n1179),.clk(gclk));
	jxor g1108(.dina(w_n1179_0[1]),.dinb(w_dff_B_PsF3JsDJ6_1),.dout(n1180),.clk(gclk));
	jand g1109(.dina(n1180),.dinb(w_n1178_0[1]),.dout(n1181),.clk(gclk));
	jnot g1110(.din(w_n1178_0[0]),.dout(n1182),.clk(gclk));
	jxor g1111(.dina(w_n1114_0[0]),.dinb(w_n1053_0[0]),.dout(n1183),.clk(gclk));
	jxor g1112(.dina(n1183),.dinb(w_n1179_0[0]),.dout(n1184),.clk(gclk));
	jand g1113(.dina(w_n1184_0[1]),.dinb(w_dff_B_ep09lUf91_1),.dout(n1185),.clk(gclk));
	jor g1114(.dina(n1185),.dinb(n1181),.dout(n1186),.clk(gclk));
	jxor g1115(.dina(n1186),.dinb(w_n1177_0[1]),.dout(G405),.clk(gclk));
	jxor g1116(.dina(w_n1184_0[0]),.dinb(w_n1177_0[0]),.dout(w_dff_A_nMRnQXEZ3_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_dff_A_Z3J2hJSb1_2),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_dff_A_N5jP9i6U3_0),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_dff_A_aAR6pYCz9_1),.din(w_G1_0[1]));
	jspl3 jspl3_w_G13_0(.douta(w_G13_0[0]),.doutb(w_G13_0[1]),.doutc(w_G13_0[2]),.din(G13));
	jspl3 jspl3_w_G13_1(.douta(w_dff_A_a2pL4i4R6_0),.doutb(w_dff_A_DU8SRIU89_1),.doutc(w_G13_1[2]),.din(w_G13_0[0]));
	jspl jspl_w_G13_2(.douta(w_dff_A_e3s8cSwM6_0),.doutb(w_G13_2[1]),.din(w_G13_0[1]));
	jspl3 jspl3_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.doutc(w_dff_A_4X5ktXLG6_2),.din(G20));
	jspl3 jspl3_w_G20_1(.douta(w_dff_A_umfdCvHV8_0),.doutb(w_G20_1[1]),.doutc(w_G20_1[2]),.din(w_G20_0[0]));
	jspl3 jspl3_w_G20_2(.douta(w_G20_2[0]),.doutb(w_G20_2[1]),.doutc(w_dff_A_Za5J4EeW1_2),.din(w_G20_0[1]));
	jspl3 jspl3_w_G20_3(.douta(w_G20_3[0]),.doutb(w_G20_3[1]),.doutc(w_dff_A_CJmQAE0W4_2),.din(w_G20_0[2]));
	jspl3 jspl3_w_G20_4(.douta(w_G20_4[0]),.doutb(w_dff_A_Mk9d0q7l7_1),.doutc(w_dff_A_bzBoME3G6_2),.din(w_G20_1[0]));
	jspl3 jspl3_w_G20_5(.douta(w_dff_A_S8Ex2UsS9_0),.doutb(w_G20_5[1]),.doutc(w_G20_5[2]),.din(w_G20_1[1]));
	jspl3 jspl3_w_G20_6(.douta(w_dff_A_4naE8Tex9_0),.doutb(w_G20_6[1]),.doutc(w_dff_A_WDaLdjET0_2),.din(w_G20_1[2]));
	jspl3 jspl3_w_G33_0(.douta(w_dff_A_Fe2KaN991_0),.doutb(w_G33_0[1]),.doutc(w_G33_0[2]),.din(G33));
	jspl3 jspl3_w_G33_1(.douta(w_dff_A_2SGy3vXE7_0),.doutb(w_dff_A_iCkZqIXJ7_1),.doutc(w_G33_1[2]),.din(w_G33_0[0]));
	jspl3 jspl3_w_G33_2(.douta(w_G33_2[0]),.doutb(w_G33_2[1]),.doutc(w_G33_2[2]),.din(w_G33_0[1]));
	jspl3 jspl3_w_G33_3(.douta(w_G33_3[0]),.doutb(w_G33_3[1]),.doutc(w_G33_3[2]),.din(w_G33_0[2]));
	jspl3 jspl3_w_G33_4(.douta(w_dff_A_5O647Yik4_0),.doutb(w_dff_A_90HwEfKC6_1),.doutc(w_G33_4[2]),.din(w_G33_1[0]));
	jspl3 jspl3_w_G33_5(.douta(w_G33_5[0]),.doutb(w_dff_A_yuAZQRgU4_1),.doutc(w_G33_5[2]),.din(w_G33_1[1]));
	jspl3 jspl3_w_G33_6(.douta(w_dff_A_tvZyrkCr1_0),.doutb(w_dff_A_4ED3xgM51_1),.doutc(w_G33_6[2]),.din(w_G33_1[2]));
	jspl3 jspl3_w_G33_7(.douta(w_dff_A_KAokJYo86_0),.doutb(w_dff_A_awdv05eE1_1),.doutc(w_G33_7[2]),.din(w_G33_2[0]));
	jspl3 jspl3_w_G33_8(.douta(w_G33_8[0]),.doutb(w_dff_A_ugfSWE8Z0_1),.doutc(w_G33_8[2]),.din(w_G33_2[1]));
	jspl3 jspl3_w_G33_9(.douta(w_dff_A_LFqTsjbc6_0),.doutb(w_dff_A_YBop4ogN4_1),.doutc(w_G33_9[2]),.din(w_G33_2[2]));
	jspl3 jspl3_w_G33_10(.douta(w_G33_10[0]),.doutb(w_G33_10[1]),.doutc(w_G33_10[2]),.din(w_G33_3[0]));
	jspl3 jspl3_w_G33_11(.douta(w_G33_11[0]),.doutb(w_G33_11[1]),.doutc(w_G33_11[2]),.din(w_G33_3[1]));
	jspl3 jspl3_w_G33_12(.douta(w_G33_12[0]),.doutb(w_dff_A_4G19A59n2_1),.doutc(w_dff_A_6UMkh2iw9_2),.din(w_G33_3[2]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_G41_0[1]),.doutc(w_G41_0[2]),.din(G41));
	jspl3 jspl3_w_G45_0(.douta(w_G45_0[0]),.doutb(w_dff_A_aZAttY8G0_1),.doutc(w_G45_0[2]),.din(G45));
	jspl jspl_w_G45_1(.douta(w_G45_1[0]),.doutb(w_dff_A_gIp1idMr6_1),.din(w_G45_0[0]));
	jspl3 jspl3_w_G50_0(.douta(w_G50_0[0]),.doutb(w_G50_0[1]),.doutc(w_G50_0[2]),.din(G50));
	jspl3 jspl3_w_G50_1(.douta(w_dff_A_uRXQAEmO4_0),.doutb(w_G50_1[1]),.doutc(w_dff_A_TfYO4oLX8_2),.din(w_G50_0[0]));
	jspl3 jspl3_w_G50_2(.douta(w_G50_2[0]),.doutb(w_dff_A_N4Y2Mr3N2_1),.doutc(w_dff_A_nLJPHWsy8_2),.din(w_G50_0[1]));
	jspl3 jspl3_w_G50_3(.douta(w_dff_A_Yq1g9EbF9_0),.doutb(w_dff_A_W5vhrWtU2_1),.doutc(w_G50_3[2]),.din(w_G50_0[2]));
	jspl3 jspl3_w_G50_4(.douta(w_dff_A_myzgEm6o4_0),.doutb(w_dff_A_IatAuJ4D8_1),.doutc(w_G50_4[2]),.din(w_G50_1[0]));
	jspl3 jspl3_w_G50_5(.douta(w_G50_5[0]),.doutb(w_dff_A_5FfXtKws4_1),.doutc(w_G50_5[2]),.din(w_G50_1[1]));
	jspl3 jspl3_w_G58_0(.douta(w_G58_0[0]),.doutb(w_dff_A_ID44LOwM4_1),.doutc(w_G58_0[2]),.din(G58));
	jspl3 jspl3_w_G58_1(.douta(w_G58_1[0]),.doutb(w_G58_1[1]),.doutc(w_dff_A_oDEU0Bbw2_2),.din(w_G58_0[0]));
	jspl3 jspl3_w_G58_2(.douta(w_dff_A_tuXdhDwY1_0),.doutb(w_G58_2[1]),.doutc(w_dff_A_bAIyhmRv0_2),.din(w_G58_0[1]));
	jspl3 jspl3_w_G58_3(.douta(w_dff_A_QDZZMnUA1_0),.doutb(w_G58_3[1]),.doutc(w_dff_A_ziTFnVBC9_2),.din(w_G58_0[2]));
	jspl3 jspl3_w_G58_4(.douta(w_dff_A_JDcLtCSU8_0),.doutb(w_G58_4[1]),.doutc(w_dff_A_ga0eICyE4_2),.din(w_G58_1[0]));
	jspl3 jspl3_w_G58_5(.douta(w_dff_A_4T2OBKU75_0),.doutb(w_G58_5[1]),.doutc(w_G58_5[2]),.din(w_G58_1[1]));
	jspl3 jspl3_w_G68_0(.douta(w_G68_0[0]),.doutb(w_G68_0[1]),.doutc(w_dff_A_hIy1Evbj3_2),.din(G68));
	jspl3 jspl3_w_G68_1(.douta(w_G68_1[0]),.doutb(w_G68_1[1]),.doutc(w_dff_A_atCkOc2f6_2),.din(w_G68_0[0]));
	jspl3 jspl3_w_G68_2(.douta(w_G68_2[0]),.doutb(w_dff_A_xOXKEPir9_1),.doutc(w_dff_A_V27RGjLX5_2),.din(w_G68_0[1]));
	jspl3 jspl3_w_G68_3(.douta(w_G68_3[0]),.doutb(w_dff_A_gkhyvNus0_1),.doutc(w_dff_A_YbKn54312_2),.din(w_G68_0[2]));
	jspl3 jspl3_w_G68_4(.douta(w_dff_A_vb2mpHcf6_0),.doutb(w_G68_4[1]),.doutc(w_dff_A_OE7sgIuQ1_2),.din(w_G68_1[0]));
	jspl3 jspl3_w_G68_5(.douta(w_dff_A_GYNZU5xm9_0),.doutb(w_G68_5[1]),.doutc(w_G68_5[2]),.din(w_G68_1[1]));
	jspl3 jspl3_w_G77_0(.douta(w_G77_0[0]),.doutb(w_dff_A_TlHlMIDS6_1),.doutc(w_G77_0[2]),.din(G77));
	jspl3 jspl3_w_G77_1(.douta(w_G77_1[0]),.doutb(w_dff_A_t101vT8I6_1),.doutc(w_G77_1[2]),.din(w_G77_0[0]));
	jspl3 jspl3_w_G77_2(.douta(w_dff_A_PcNxiZVX6_0),.doutb(w_dff_A_IIsPcozW7_1),.doutc(w_G77_2[2]),.din(w_G77_0[1]));
	jspl3 jspl3_w_G77_3(.douta(w_dff_A_RnLehcsx9_0),.doutb(w_G77_3[1]),.doutc(w_dff_A_6R5e6Vpw8_2),.din(w_G77_0[2]));
	jspl3 jspl3_w_G77_4(.douta(w_dff_A_66Lb5xL71_0),.doutb(w_G77_4[1]),.doutc(w_G77_4[2]),.din(w_G77_1[0]));
	jspl3 jspl3_w_G87_0(.douta(w_dff_A_tP0ttjuI6_0),.doutb(w_G87_0[1]),.doutc(w_G87_0[2]),.din(G87));
	jspl3 jspl3_w_G87_1(.douta(w_G87_1[0]),.doutb(w_dff_A_O0UPS0rg6_1),.doutc(w_dff_A_u3LkBAgE3_2),.din(w_G87_0[0]));
	jspl3 jspl3_w_G87_2(.douta(w_dff_A_lb8DHTMQ0_0),.doutb(w_dff_A_sCFfnYDW2_1),.doutc(w_G87_2[2]),.din(w_G87_0[1]));
	jspl3 jspl3_w_G87_3(.douta(w_dff_A_FMuI1CcA8_0),.doutb(w_G87_3[1]),.doutc(w_G87_3[2]),.din(w_G87_0[2]));
	jspl3 jspl3_w_G97_0(.douta(w_G97_0[0]),.doutb(w_dff_A_ytpqUgnf0_1),.doutc(w_G97_0[2]),.din(G97));
	jspl3 jspl3_w_G97_1(.douta(w_G97_1[0]),.doutb(w_dff_A_l8TPzBcC4_1),.doutc(w_dff_A_6yYBYou13_2),.din(w_G97_0[0]));
	jspl3 jspl3_w_G97_2(.douta(w_G97_2[0]),.doutb(w_dff_A_YnKQKoVh5_1),.doutc(w_G97_2[2]),.din(w_G97_0[1]));
	jspl3 jspl3_w_G97_3(.douta(w_dff_A_P9BlaCSh4_0),.doutb(w_G97_3[1]),.doutc(w_G97_3[2]),.din(w_G97_0[2]));
	jspl3 jspl3_w_G97_4(.douta(w_dff_A_sDaQeqU74_0),.doutb(w_G97_4[1]),.doutc(w_G97_4[2]),.din(w_G97_1[0]));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_dff_A_JOflgydm7_1),.doutc(w_G107_0[2]),.din(G107));
	jspl3 jspl3_w_G107_1(.douta(w_G107_1[0]),.doutb(w_dff_A_6ineyHI54_1),.doutc(w_dff_A_AfTxsI4D4_2),.din(w_G107_0[0]));
	jspl3 jspl3_w_G107_2(.douta(w_G107_2[0]),.doutb(w_dff_A_GugwOcEI1_1),.doutc(w_G107_2[2]),.din(w_G107_0[1]));
	jspl3 jspl3_w_G107_3(.douta(w_dff_A_1053Xzse9_0),.doutb(w_G107_3[1]),.doutc(w_G107_3[2]),.din(w_G107_0[2]));
	jspl jspl_w_G107_4(.douta(w_dff_A_ieJJYPRg7_0),.doutb(w_G107_4[1]),.din(w_G107_1[0]));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_dff_A_6Jnib6tG3_1),.doutc(w_dff_A_7SiU0GIE8_2),.din(G116));
	jspl3 jspl3_w_G116_1(.douta(w_G116_1[0]),.doutb(w_G116_1[1]),.doutc(w_dff_A_7FnPaeON8_2),.din(w_G116_0[0]));
	jspl3 jspl3_w_G116_2(.douta(w_G116_2[0]),.doutb(w_G116_2[1]),.doutc(w_dff_A_cUW9NY2e1_2),.din(w_G116_0[1]));
	jspl3 jspl3_w_G116_3(.douta(w_G116_3[0]),.doutb(w_G116_3[1]),.doutc(w_G116_3[2]),.din(w_G116_0[2]));
	jspl3 jspl3_w_G116_4(.douta(w_dff_A_aCfmhJLD5_0),.doutb(w_G116_4[1]),.doutc(w_G116_4[2]),.din(w_G116_1[0]));
	jspl3 jspl3_w_G116_5(.douta(w_dff_A_cIXMQj1C0_0),.doutb(w_dff_A_VKaiihHm3_1),.doutc(w_G116_5[2]),.din(w_G116_1[1]));
	jspl jspl_w_G125_0(.douta(w_G125_0[0]),.doutb(w_dff_A_6fwpVXDc5_1),.din(w_dff_B_osGoo7l30_2));
	jspl3 jspl3_w_G128_0(.douta(w_dff_A_YWRtBQ7V5_0),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(w_dff_B_aXjaDQ4M0_3));
	jspl3 jspl3_w_G132_0(.douta(w_G132_0[0]),.doutb(w_G132_0[1]),.doutc(w_G132_0[2]),.din(w_dff_B_EDPlRGQZ8_3));
	jspl jspl_w_G132_1(.douta(w_G132_1[0]),.doutb(w_dff_A_97lxGxD29_1),.din(w_G132_0[0]));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(w_dff_B_24faEiGY7_3));
	jspl3 jspl3_w_G137_1(.douta(w_G137_1[0]),.doutb(w_dff_A_8cGpDfv52_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(w_dff_B_2fQBAMhR4_3));
	jspl3 jspl3_w_G143_1(.douta(w_G143_1[0]),.doutb(w_G143_1[1]),.doutc(w_dff_A_0FXdgbTT2_2),.din(w_G143_0[0]));
	jspl jspl_w_G143_2(.douta(w_G143_2[0]),.doutb(w_G143_2[1]),.din(w_G143_0[1]));
	jspl3 jspl3_w_G150_0(.douta(w_dff_A_xY4JYrGU6_0),.doutb(w_dff_A_fhwY2GGF7_1),.doutc(w_G150_0[2]),.din(w_dff_B_rVxBzmCT4_3));
	jspl3 jspl3_w_G150_1(.douta(w_G150_1[0]),.doutb(w_dff_A_JIa7x4XB8_1),.doutc(w_G150_1[2]),.din(w_G150_0[0]));
	jspl3 jspl3_w_G150_2(.douta(w_G150_2[0]),.doutb(w_dff_A_sDiaw4jP0_1),.doutc(w_G150_2[2]),.din(w_G150_0[1]));
	jspl jspl_w_G150_3(.douta(w_dff_A_nbkZK3gz7_0),.doutb(w_G150_3[1]),.din(w_G150_0[2]));
	jspl3 jspl3_w_G159_0(.douta(w_dff_A_gTmJHqmw8_0),.doutb(w_dff_A_02gL5xdu7_1),.doutc(w_G159_0[2]),.din(G159));
	jspl3 jspl3_w_G159_1(.douta(w_G159_1[0]),.doutb(w_G159_1[1]),.doutc(w_dff_A_oAPZEv3J5_2),.din(w_G159_0[0]));
	jspl3 jspl3_w_G159_2(.douta(w_G159_2[0]),.doutb(w_G159_2[1]),.doutc(w_G159_2[2]),.din(w_G159_0[1]));
	jspl3 jspl3_w_G159_3(.douta(w_dff_A_uCHVmEAR2_0),.doutb(w_dff_A_OjRpaYTH3_1),.doutc(w_G159_3[2]),.din(w_G159_0[2]));
	jspl3 jspl3_w_G169_0(.douta(w_dff_A_GBIGJCYs5_0),.doutb(w_dff_A_Gi5qJDve0_1),.doutc(w_G169_0[2]),.din(G169));
	jspl3 jspl3_w_G169_1(.douta(w_G169_1[0]),.doutb(w_dff_A_Zq0Bc14H4_1),.doutc(w_dff_A_n08iQj1A2_2),.din(w_G169_0[0]));
	jspl3 jspl3_w_G169_2(.douta(w_dff_A_gaaqrNnu9_0),.doutb(w_dff_A_CZyKlEfI8_1),.doutc(w_G169_2[2]),.din(w_G169_0[1]));
	jspl jspl_w_G169_3(.douta(w_G169_3[0]),.doutb(w_dff_A_53LigxUI3_1),.din(w_G169_0[2]));
	jspl3 jspl3_w_G179_0(.douta(w_dff_A_kBLVlvFw4_0),.doutb(w_G179_0[1]),.doutc(w_G179_0[2]),.din(G179));
	jspl3 jspl3_w_G179_1(.douta(w_G179_1[0]),.doutb(w_G179_1[1]),.doutc(w_G179_1[2]),.din(w_G179_0[0]));
	jspl3 jspl3_w_G179_2(.douta(w_dff_A_adNHm5Ts5_0),.doutb(w_dff_A_C1uqPPe31_1),.doutc(w_G179_2[2]),.din(w_G179_0[1]));
	jspl3 jspl3_w_G190_0(.douta(w_dff_A_AOAazSbn8_0),.doutb(w_G190_0[1]),.doutc(w_dff_A_TufCRslF2_2),.din(G190));
	jspl3 jspl3_w_G190_1(.douta(w_dff_A_e7aAggJJ6_0),.doutb(w_G190_1[1]),.doutc(w_G190_1[2]),.din(w_G190_0[0]));
	jspl3 jspl3_w_G190_2(.douta(w_dff_A_mj3y81XF0_0),.doutb(w_G190_2[1]),.doutc(w_dff_A_exnGLAXE9_2),.din(w_G190_0[1]));
	jspl3 jspl3_w_G190_3(.douta(w_dff_A_pI5UWDYu8_0),.doutb(w_dff_A_rkfMiR059_1),.doutc(w_G190_3[2]),.din(w_G190_0[2]));
	jspl3 jspl3_w_G190_4(.douta(w_G190_4[0]),.doutb(w_dff_A_3jLZoVp15_1),.doutc(w_dff_A_hxtQ4qkq4_2),.din(w_G190_1[0]));
	jspl3 jspl3_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.doutc(w_dff_A_7TIFVRkI6_2),.din(G200));
	jspl3 jspl3_w_G200_1(.douta(w_dff_A_WuJdh9tN4_0),.doutb(w_G200_1[1]),.doutc(w_dff_A_qJJ0psJq6_2),.din(w_G200_0[0]));
	jspl3 jspl3_w_G200_2(.douta(w_G200_2[0]),.doutb(w_dff_A_JVEiqZj74_1),.doutc(w_dff_A_RuwTxlmp4_2),.din(w_G200_0[1]));
	jspl jspl_w_G200_3(.douta(w_G200_3[0]),.doutb(w_G200_3[1]),.din(w_G200_0[2]));
	jspl3 jspl3_w_G213_0(.douta(w_dff_A_lJ5nagS34_0),.doutb(w_G213_0[1]),.doutc(w_dff_A_raF79JIE4_2),.din(G213));
	jspl jspl_w_G223_0(.douta(w_G223_0[0]),.doutb(w_G223_0[1]),.din(w_dff_B_zdMtXarI8_2));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_dff_A_8DaOgCE19_1),.doutc(w_dff_A_cOKP08oN6_2),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_dff_A_wBv5RdHQ9_0),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G232_0(.douta(w_G232_0[0]),.doutb(w_dff_A_5mpRZrMx0_1),.doutc(w_dff_A_rGcJMBIj6_2),.din(G232));
	jspl3 jspl3_w_G232_1(.douta(w_dff_A_40PAzvkt0_0),.doutb(w_G232_1[1]),.doutc(w_G232_1[2]),.din(w_G232_0[0]));
	jspl3 jspl3_w_G238_0(.douta(w_dff_A_WGcIau8i4_0),.doutb(w_dff_A_vm0PmMfd2_1),.doutc(w_G238_0[2]),.din(G238));
	jspl3 jspl3_w_G244_0(.douta(w_G244_0[0]),.doutb(w_dff_A_xBgHXuCO4_1),.doutc(w_dff_A_a4qbyPcr0_2),.din(G244));
	jspl jspl_w_G244_1(.douta(w_dff_A_DBtIjgyf7_0),.doutb(w_G244_1[1]),.din(w_G244_0[0]));
	jspl3 jspl3_w_G250_0(.douta(w_dff_A_UifMbqcT0_0),.doutb(w_G250_0[1]),.doutc(w_G250_0[2]),.din(G250));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_dff_A_LseBYIOK8_1),.doutc(w_dff_A_TGsmLIqQ6_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_XjVZ48HX4_0),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G264_0(.douta(w_dff_A_B212phLv9_0),.doutb(w_dff_A_ahXSG8UL4_1),.doutc(w_G264_0[2]),.din(G264));
	jspl3 jspl3_w_G270_0(.douta(w_dff_A_D30XsiAm4_0),.doutb(w_dff_A_AYEVyLfQ3_1),.doutc(w_G270_0[2]),.din(G270));
	jspl3 jspl3_w_G274_0(.douta(w_dff_A_u6jQZWCN8_0),.doutb(w_G274_0[1]),.doutc(w_dff_A_GSO5PdCL6_2),.din(G274));
	jspl3 jspl3_w_G283_0(.douta(w_dff_A_G7tY3cCa7_0),.doutb(w_dff_A_IrXp32UJ4_1),.doutc(w_G283_0[2]),.din(G283));
	jspl3 jspl3_w_G283_1(.douta(w_G283_1[0]),.doutb(w_dff_A_bvHEwYPn0_1),.doutc(w_G283_1[2]),.din(w_G283_0[0]));
	jspl3 jspl3_w_G283_2(.douta(w_G283_2[0]),.doutb(w_dff_A_XgHMaMKJ0_1),.doutc(w_G283_2[2]),.din(w_G283_0[1]));
	jspl3 jspl3_w_G283_3(.douta(w_dff_A_UMyuYaC41_0),.doutb(w_dff_A_OcKfnYpe3_1),.doutc(w_G283_3[2]),.din(w_G283_0[2]));
	jspl3 jspl3_w_G294_0(.douta(w_dff_A_M8PDc24u2_0),.doutb(w_dff_A_UGB6UDPz6_1),.doutc(w_G294_0[2]),.din(G294));
	jspl3 jspl3_w_G294_1(.douta(w_G294_1[0]),.doutb(w_dff_A_p726uaCi3_1),.doutc(w_G294_1[2]),.din(w_G294_0[0]));
	jspl3 jspl3_w_G294_2(.douta(w_G294_2[0]),.doutb(w_G294_2[1]),.doutc(w_G294_2[2]),.din(w_G294_0[1]));
	jspl jspl_w_G294_3(.douta(w_dff_A_7KXAvexG1_0),.doutb(w_G294_3[1]),.din(w_G294_0[2]));
	jspl3 jspl3_w_G303_0(.douta(w_dff_A_5em3aR5A7_0),.doutb(w_G303_0[1]),.doutc(w_dff_A_qt1GiljN0_2),.din(G303));
	jspl3 jspl3_w_G303_1(.douta(w_G303_1[0]),.doutb(w_G303_1[1]),.doutc(w_G303_1[2]),.din(w_G303_0[0]));
	jspl3 jspl3_w_G303_2(.douta(w_dff_A_hMpawB0o6_0),.doutb(w_dff_A_Z1eKN7YO8_1),.doutc(w_G303_2[2]),.din(w_G303_0[1]));
	jspl3 jspl3_w_G311_0(.douta(w_G311_0[0]),.doutb(w_G311_0[1]),.doutc(w_G311_0[2]),.din(w_dff_B_DleL7hkB5_3));
	jspl3 jspl3_w_G311_1(.douta(w_G311_1[0]),.doutb(w_dff_A_FduAQ6k65_1),.doutc(w_G311_1[2]),.din(w_G311_0[0]));
	jspl3 jspl3_w_G317_0(.douta(w_G317_0[0]),.doutb(w_G317_0[1]),.doutc(w_G317_0[2]),.din(w_dff_B_aZT4eAIR2_3));
	jspl jspl_w_G317_1(.douta(w_dff_A_wFVyREYN6_0),.doutb(w_G317_1[1]),.din(w_G317_0[0]));
	jspl3 jspl3_w_G322_0(.douta(w_dff_A_IgwH6UHi3_0),.doutb(w_G322_0[1]),.doutc(w_G322_0[2]),.din(w_dff_B_76RyYuVJ5_3));
	jspl jspl_w_G326_0(.douta(w_dff_A_UAHBuC8a9_0),.doutb(w_G326_0[1]),.din(w_dff_B_3IYLQbVv5_2));
	jspl3 jspl3_w_G330_0(.douta(w_dff_A_92WyQHFf7_0),.doutb(w_G330_0[1]),.doutc(w_dff_A_2LB4S6lL1_2),.din(w_dff_B_LllyakdK2_3));
	jspl jspl_w_G343_0(.douta(w_G343_0[0]),.doutb(w_dff_A_aA2Efb6n2_1),.din(G343));
	jspl3 jspl3_w_G1698_0(.douta(w_G1698_0[0]),.doutb(w_G1698_0[1]),.doutc(w_dff_A_rzrEgui05_2),.din(G1698));
	jspl jspl_w_G355_0(.douta(w_dff_A_2tQIXM091_0),.doutb(w_dff_A_heHbqSsj6_1),.din(G355_fa_));
	jspl jspl_w_G396_0(.douta(w_G396_0),.doutb(w_dff_A_0XfjDTOX8_1),.din(G396_fa_));
	jspl jspl_w_G384_0(.douta(w_dff_A_UDsUAlsV2_0),.doutb(w_dff_A_w0ospIK34_1),.din(G384_fa_));
	jspl3 jspl3_w_n72_0(.douta(w_n72_0[0]),.doutb(w_dff_A_UjcH846S9_1),.doutc(w_dff_A_AOrGp42Y8_2),.din(n72));
	jspl3 jspl3_w_n72_1(.douta(w_n72_1[0]),.doutb(w_n72_1[1]),.doutc(w_dff_A_ZVkHsFxW5_2),.din(w_n72_0[0]));
	jspl3 jspl3_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.doutc(w_dff_A_8fctjVtq2_2),.din(n73));
	jspl3 jspl3_w_n73_1(.douta(w_n73_1[0]),.doutb(w_dff_A_YyiYAuhi0_1),.doutc(w_dff_A_FadPCto76_2),.din(w_n73_0[0]));
	jspl3 jspl3_w_n73_2(.douta(w_dff_A_0l8nIW9H9_0),.doutb(w_n73_2[1]),.doutc(w_dff_A_o7WcTBV71_2),.din(w_n73_0[1]));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_dff_A_Q82G0qZs0_2),.din(n74));
	jspl3 jspl3_w_n74_1(.douta(w_n74_1[0]),.doutb(w_dff_A_JEG8Zf214_1),.doutc(w_dff_A_jI0YuI4j5_2),.din(w_n74_0[0]));
	jspl jspl_w_n74_2(.douta(w_n74_2[0]),.doutb(w_n74_2[1]),.din(w_n74_0[1]));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.doutc(w_dff_A_Evudwhde2_2),.din(n75));
	jspl3 jspl3_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.doutc(w_n75_1[2]),.din(w_n75_0[0]));
	jspl jspl_w_n75_2(.douta(w_n75_2[0]),.doutb(w_n75_2[1]),.din(w_n75_0[1]));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.din(n76));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl3 jspl3_w_n79_0(.douta(w_n79_0[0]),.doutb(w_dff_A_N68nDtWQ1_1),.doutc(w_n79_0[2]),.din(n79));
	jspl3 jspl3_w_n79_1(.douta(w_dff_A_OFeyg3eT2_0),.doutb(w_n79_1[1]),.doutc(w_dff_A_PRuOSv1q6_2),.din(w_n79_0[0]));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_dff_A_sukh36C02_1),.doutc(w_dff_A_pK4nazjv8_2),.din(n80));
	jspl3 jspl3_w_n80_1(.douta(w_n80_1[0]),.doutb(w_n80_1[1]),.doutc(w_n80_1[2]),.din(w_n80_0[0]));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_dff_A_NKXy33Zt9_2),.din(n81));
	jspl3 jspl3_w_n81_1(.douta(w_dff_A_wpDTwxvd2_0),.doutb(w_n81_1[1]),.doutc(w_n81_1[2]),.din(w_n81_0[0]));
	jspl jspl_w_n81_2(.douta(w_n81_2[0]),.doutb(w_n81_2[1]),.din(w_n81_0[1]));
	jspl3 jspl3_w_n84_0(.douta(w_n84_0[0]),.doutb(w_dff_A_4Z7QsvPG7_1),.doutc(w_dff_A_9Zcfe4AD1_2),.din(n84));
	jspl3 jspl3_w_n84_1(.douta(w_n84_1[0]),.doutb(w_n84_1[1]),.doutc(w_dff_A_JqIje15q7_2),.din(w_n84_0[0]));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl3 jspl3_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.doutc(w_n86_0[2]),.din(n86));
	jspl jspl_w_n89_0(.douta(w_n89_0[0]),.doutb(w_n89_0[1]),.din(n89));
	jspl3 jspl3_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.doutc(w_n91_0[2]),.din(n91));
	jspl3 jspl3_w_n91_1(.douta(w_n91_1[0]),.doutb(w_n91_1[1]),.doutc(w_n91_1[2]),.din(w_n91_0[0]));
	jspl3 jspl3_w_n94_0(.douta(w_dff_A_2fVsdO4y2_0),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.doutc(w_n96_0[2]),.din(n96));
	jspl3 jspl3_w_n105_0(.douta(w_n105_0[0]),.doutb(w_dff_A_TB5hfQ0o8_1),.doutc(w_dff_A_p1Lv5tZs8_2),.din(n105));
	jspl jspl_w_n105_1(.douta(w_dff_A_qgWVCfvQ1_0),.doutb(w_n105_1[1]),.din(w_n105_0[0]));
	jspl3 jspl3_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.doutc(w_n111_0[2]),.din(n111));
	jspl jspl_w_n112_0(.douta(w_dff_A_VV0G5Xfi3_0),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_dff_A_fqJ0YkIr5_1),.din(n120));
	jspl jspl_w_n126_0(.douta(w_dff_A_oZ09gIbv8_0),.doutb(w_n126_0[1]),.din(n126));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_dff_A_K5y6vMox0_1),.din(n130));
	jspl jspl_w_n134_0(.douta(w_n134_0[0]),.doutb(w_dff_A_IfmgPiJs5_1),.din(n134));
	jspl jspl_w_n137_0(.douta(w_dff_A_NxLNoeNl9_0),.doutb(w_n137_0[1]),.din(n137));
	jspl3 jspl3_w_n139_0(.douta(w_n139_0[0]),.doutb(w_n139_0[1]),.doutc(w_n139_0[2]),.din(n139));
	jspl3 jspl3_w_n139_1(.douta(w_dff_A_4m3fVzqZ7_0),.doutb(w_n139_1[1]),.doutc(w_dff_A_Xf56kWhH1_2),.din(w_n139_0[0]));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.doutc(w_n141_0[2]),.din(n141));
	jspl3 jspl3_w_n141_1(.douta(w_n141_1[0]),.doutb(w_dff_A_uBod4A164_1),.doutc(w_dff_A_6qfkpFnA6_2),.din(w_n141_0[0]));
	jspl3 jspl3_w_n141_2(.douta(w_dff_A_y5iOTmpa2_0),.doutb(w_n141_2[1]),.doutc(w_n141_2[2]),.din(w_n141_0[1]));
	jspl jspl_w_n141_3(.douta(w_dff_A_H7EoIeNt4_0),.doutb(w_n141_3[1]),.din(w_n141_0[2]));
	jspl3 jspl3_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.doutc(w_dff_A_VsLbwrtO3_2),.din(n142));
	jspl3 jspl3_w_n142_1(.douta(w_dff_A_RfddQYn10_0),.doutb(w_n142_1[1]),.doutc(w_n142_1[2]),.din(w_n142_0[0]));
	jspl jspl_w_n142_2(.douta(w_n142_2[0]),.doutb(w_n142_2[1]),.din(w_n142_0[1]));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n144_1(.douta(w_n144_1[0]),.doutb(w_n144_1[1]),.doutc(w_n144_1[2]),.din(w_n144_0[0]));
	jspl jspl_w_n144_2(.douta(w_n144_2[0]),.doutb(w_n144_2[1]),.din(w_n144_0[1]));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl jspl_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.din(n148));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_dff_A_QoYS69xf0_1),.doutc(w_dff_A_J6xfLXCV2_2),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_dff_A_6jCIhLww4_0),.doutb(w_n151_2[1]),.doutc(w_dff_A_0bioxm1z1_2),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_n151_3[0]),.doutb(w_n151_3[1]),.doutc(w_dff_A_PzhApn8n0_2),.din(w_n151_0[2]));
	jspl3 jspl3_w_n151_4(.douta(w_n151_4[0]),.doutb(w_dff_A_4MwNiXOn4_1),.doutc(w_n151_4[2]),.din(w_n151_1[0]));
	jspl3 jspl3_w_n151_5(.douta(w_dff_A_WruRIkvC8_0),.doutb(w_n151_5[1]),.doutc(w_n151_5[2]),.din(w_n151_1[1]));
	jspl jspl_w_n151_6(.douta(w_dff_A_lypYdccR6_0),.doutb(w_n151_6[1]),.din(w_n151_1[2]));
	jspl3 jspl3_w_n152_0(.douta(w_dff_A_oJeBx24G4_0),.doutb(w_n152_0[1]),.doutc(w_dff_A_UWfbyl1h1_2),.din(n152));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_dff_A_y8uCNX1z9_2),.din(n153));
	jspl3 jspl3_w_n153_1(.douta(w_dff_A_RNoxb2dK4_0),.doutb(w_n153_1[1]),.doutc(w_n153_1[2]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n153_2(.douta(w_n153_2[0]),.doutb(w_n153_2[1]),.doutc(w_dff_A_dZAaiECU3_2),.din(w_n153_0[1]));
	jspl3 jspl3_w_n153_3(.douta(w_n153_3[0]),.doutb(w_dff_A_tsGL62uo6_1),.doutc(w_dff_A_x9FcaIIF3_2),.din(w_n153_0[2]));
	jspl3 jspl3_w_n153_4(.douta(w_dff_A_3RdTVT158_0),.doutb(w_dff_A_zIyt1ZDW7_1),.doutc(w_n153_4[2]),.din(w_n153_1[0]));
	jspl3 jspl3_w_n153_5(.douta(w_dff_A_uk6JKueg4_0),.doutb(w_n153_5[1]),.doutc(w_n153_5[2]),.din(w_n153_1[1]));
	jspl3 jspl3_w_n153_6(.douta(w_n153_6[0]),.doutb(w_n153_6[1]),.doutc(w_n153_6[2]),.din(w_n153_1[2]));
	jspl3 jspl3_w_n153_7(.douta(w_n153_7[0]),.doutb(w_n153_7[1]),.doutc(w_n153_7[2]),.din(w_n153_2[0]));
	jspl jspl_w_n153_8(.douta(w_n153_8[0]),.doutb(w_n153_8[1]),.din(w_n153_2[1]));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_dff_A_agZidya10_1),.doutc(w_n161_0[2]),.din(n161));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_dff_A_Ug09h26b1_1),.doutc(w_dff_A_jIXxqQBl5_2),.din(n163));
	jspl jspl_w_n163_1(.douta(w_n163_1[0]),.doutb(w_dff_A_Ehupaxh00_1),.din(w_n163_0[0]));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_n164_0[2]),.din(n164));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_kNaDVNSq3_1),.din(n165));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_dff_A_XTFGpIVr3_1),.din(n167));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl3 jspl3_w_n168_1(.douta(w_n168_1[0]),.doutb(w_n168_1[1]),.doutc(w_n168_1[2]),.din(w_n168_0[0]));
	jspl3 jspl3_w_n168_2(.douta(w_dff_A_9QBz8RYs5_0),.doutb(w_n168_2[1]),.doutc(w_n168_2[2]),.din(w_n168_0[1]));
	jspl3 jspl3_w_n168_3(.douta(w_dff_A_0C1uqOXc6_0),.doutb(w_n168_3[1]),.doutc(w_dff_A_aIBsKakw8_2),.din(w_n168_0[2]));
	jspl3 jspl3_w_n168_4(.douta(w_dff_A_ezplO8FG1_0),.doutb(w_dff_A_UT5E5WLW6_1),.doutc(w_n168_4[2]),.din(w_n168_1[0]));
	jspl jspl_w_n168_5(.douta(w_n168_5[0]),.doutb(w_n168_5[1]),.din(w_n168_1[1]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_dff_A_YJlh3oE04_2),.din(w_dff_B_j1gpmBTM4_3));
	jspl3 jspl3_w_n172_0(.douta(w_n172_0[0]),.doutb(w_dff_A_a7OroNKR0_1),.doutc(w_dff_A_rPcvYyJw0_2),.din(n172));
	jspl3 jspl3_w_n172_1(.douta(w_n172_1[0]),.doutb(w_dff_A_NwQFKoZl5_1),.doutc(w_dff_A_dZmAmqcr4_2),.din(w_n172_0[0]));
	jspl3 jspl3_w_n172_2(.douta(w_n172_2[0]),.doutb(w_n172_2[1]),.doutc(w_n172_2[2]),.din(w_n172_0[1]));
	jspl3 jspl3_w_n172_3(.douta(w_n172_3[0]),.doutb(w_n172_3[1]),.doutc(w_n172_3[2]),.din(w_n172_0[2]));
	jspl3 jspl3_w_n172_4(.douta(w_n172_4[0]),.doutb(w_dff_A_re8iwzaB9_1),.doutc(w_dff_A_qhl06zxv1_2),.din(w_n172_1[0]));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl3 jspl3_w_n173_1(.douta(w_n173_1[0]),.doutb(w_n173_1[1]),.doutc(w_n173_1[2]),.din(w_n173_0[0]));
	jspl3 jspl3_w_n173_2(.douta(w_n173_2[0]),.doutb(w_n173_2[1]),.doutc(w_n173_2[2]),.din(w_n173_0[1]));
	jspl jspl_w_n173_3(.douta(w_n173_3[0]),.doutb(w_n173_3[1]),.din(w_n173_0[2]));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.doutc(w_n177_0[2]),.din(n177));
	jspl3 jspl3_w_n177_1(.douta(w_n177_1[0]),.doutb(w_n177_1[1]),.doutc(w_n177_1[2]),.din(w_n177_0[0]));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl jspl_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n186_0(.douta(w_n186_0[0]),.doutb(w_dff_A_SyzkO7SL4_1),.doutc(w_n186_0[2]),.din(n186));
	jspl3 jspl3_w_n186_1(.douta(w_n186_1[0]),.doutb(w_n186_1[1]),.doutc(w_n186_1[2]),.din(w_n186_0[0]));
	jspl3 jspl3_w_n189_0(.douta(w_dff_A_oKT7Ez0f7_0),.doutb(w_dff_A_FPx0BJSn6_1),.doutc(w_n189_0[2]),.din(n189));
	jspl3 jspl3_w_n189_1(.douta(w_n189_1[0]),.doutb(w_dff_A_CwkCNF3L1_1),.doutc(w_n189_1[2]),.din(w_n189_0[0]));
	jspl3 jspl3_w_n189_2(.douta(w_n189_2[0]),.doutb(w_dff_A_maUN2Flg6_1),.doutc(w_dff_A_gb7dweU23_2),.din(w_n189_0[1]));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_dff_A_Uw9rA5Q79_1),.din(n190));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_dff_A_oAfHk9in3_1),.doutc(w_n192_0[2]),.din(n192));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_dff_A_PyGxFW0l7_2),.din(n198));
	jspl3 jspl3_w_n199_0(.douta(w_dff_A_kq9R0Hx92_0),.doutb(w_n199_0[1]),.doutc(w_dff_A_d9JyWCYQ8_2),.din(w_dff_B_ffUfftvl6_3));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_dff_A_smOwfoRH9_1),.din(n201));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_dff_A_eQ84Agja2_1),.din(n202));
	jspl3 jspl3_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.doutc(w_n205_0[2]),.din(n205));
	jspl jspl_w_n205_1(.douta(w_n205_1[0]),.doutb(w_n205_1[1]),.din(w_n205_0[0]));
	jspl jspl_w_n207_0(.douta(w_dff_A_bViPQEmR9_0),.doutb(w_n207_0[1]),.din(n207));
	jspl3 jspl3_w_n212_0(.douta(w_n212_0[0]),.doutb(w_dff_A_BlTCyyYc9_1),.doutc(w_n212_0[2]),.din(n212));
	jspl jspl_w_n212_1(.douta(w_n212_1[0]),.doutb(w_n212_1[1]),.din(w_n212_0[0]));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_dff_A_hlo8UFjr6_1),.din(n213));
	jspl jspl_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.din(n215));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_dff_A_jTypQ46G6_1),.din(n218));
	jspl3 jspl3_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.doutc(w_dff_A_t9qhoLV72_2),.din(n224));
	jspl jspl_w_n224_1(.douta(w_dff_A_m0U3yfr82_0),.doutb(w_n224_1[1]),.din(w_n224_0[0]));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(n225));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_dff_A_ehyGtSRL7_1),.din(n229));
	jspl3 jspl3_w_n234_0(.douta(w_n234_0[0]),.doutb(w_dff_A_Bc6Smvon8_1),.doutc(w_n234_0[2]),.din(n234));
	jspl jspl_w_n234_1(.douta(w_n234_1[0]),.doutb(w_n234_1[1]),.din(w_n234_0[0]));
	jspl3 jspl3_w_n237_0(.douta(w_n237_0[0]),.doutb(w_dff_A_1H4g7aOH3_1),.doutc(w_n237_0[2]),.din(n237));
	jspl jspl_w_n238_0(.douta(w_n238_0[0]),.doutb(w_dff_A_pbCCveUn4_1),.din(n238));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_dff_A_MeHRTeA34_1),.doutc(w_dff_A_tCXveOjQ6_2),.din(n242));
	jspl jspl_w_n243_0(.douta(w_dff_A_lUeRqMzZ6_0),.doutb(w_n243_0[1]),.din(n243));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_dff_A_jJRwyNRU9_1),.din(n247));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_dff_A_5pvZ8Iej6_1),.din(n250));
	jspl jspl_w_n251_0(.douta(w_dff_A_LKGd0RP57_0),.doutb(w_n251_0[1]),.din(n251));
	jspl3 jspl3_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.doutc(w_n255_0[2]),.din(n255));
	jspl jspl_w_n255_1(.douta(w_n255_1[0]),.doutb(w_n255_1[1]),.din(w_n255_0[0]));
	jspl jspl_w_n256_0(.douta(w_n256_0[0]),.doutb(w_dff_A_y6QJ2NYk0_1),.din(n256));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_dff_A_Q2RwdHnB6_1),.din(n257));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_dff_A_d4Ac9V5o7_1),.din(n260));
	jspl3 jspl3_w_n261_0(.douta(w_n261_0[0]),.doutb(w_dff_A_7UT1Tdcn2_1),.doutc(w_dff_A_FZAOHU4A3_2),.din(n261));
	jspl3 jspl3_w_n261_1(.douta(w_n261_1[0]),.doutb(w_n261_1[1]),.doutc(w_n261_1[2]),.din(w_n261_0[0]));
	jspl3 jspl3_w_n262_0(.douta(w_dff_A_HmUdrO5U0_0),.doutb(w_dff_A_jIEF3LPd4_1),.doutc(w_n262_0[2]),.din(n262));
	jspl jspl_w_n269_0(.douta(w_dff_A_ZNRnTKv70_0),.doutb(w_n269_0[1]),.din(n269));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl3 jspl3_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.doutc(w_n279_0[2]),.din(n279));
	jspl jspl_w_n279_1(.douta(w_n279_1[0]),.doutb(w_n279_1[1]),.din(w_n279_0[0]));
	jspl jspl_w_n282_0(.douta(w_dff_A_IvJ5Yk489_0),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_dff_A_HKxjezPj9_1),.din(n283));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl jspl_w_n298_0(.douta(w_dff_A_09glOBoH0_0),.doutb(w_n298_0[1]),.din(n298));
	jspl3 jspl3_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.doutc(w_n308_0[2]),.din(n308));
	jspl3 jspl3_w_n308_1(.douta(w_n308_1[0]),.doutb(w_n308_1[1]),.doutc(w_n308_1[2]),.din(w_n308_0[0]));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_dff_A_lCjPuVzC0_1),.din(n309));
	jspl jspl_w_n310_0(.douta(w_dff_A_r52exDBL5_0),.doutb(w_n310_0[1]),.din(n310));
	jspl jspl_w_n312_0(.douta(w_dff_A_4f98VY5J0_0),.doutb(w_n312_0[1]),.din(n312));
	jspl jspl_w_n313_0(.douta(w_dff_A_PoKWS1oL5_0),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n315_0(.douta(w_dff_A_4u1g0nRA4_0),.doutb(w_n315_0[1]),.doutc(w_dff_A_sABhtlWN3_2),.din(n315));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_dff_A_v6Kexx641_1),.din(n321));
	jspl3 jspl3_w_n323_0(.douta(w_n323_0[0]),.doutb(w_dff_A_8l4yuvmS0_1),.doutc(w_dff_A_BhmWJ5Xk8_2),.din(n323));
	jspl3 jspl3_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.doutc(w_n330_0[2]),.din(n330));
	jspl jspl_w_n333_0(.douta(w_dff_A_JS0Y1SzS9_0),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n334_0(.douta(w_dff_A_iYvogae46_0),.doutb(w_n334_0[1]),.din(n334));
	jspl jspl_w_n344_0(.douta(w_n344_0[0]),.doutb(w_n344_0[1]),.din(n344));
	jspl jspl_w_n347_0(.douta(w_n347_0[0]),.doutb(w_dff_A_I6SmfvYh6_1),.din(n347));
	jspl jspl_w_n348_0(.douta(w_dff_A_CrFou7NL0_0),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n351_0(.douta(w_n351_0[0]),.doutb(w_dff_A_UUzuMJy37_1),.din(n351));
	jspl3 jspl3_w_n352_0(.douta(w_n352_0[0]),.doutb(w_dff_A_l5QVFNa52_1),.doutc(w_dff_A_OVOzVEbJ0_2),.din(n352));
	jspl jspl_w_n352_1(.douta(w_dff_A_Ur4fGXuz7_0),.doutb(w_n352_1[1]),.din(w_n352_0[0]));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_dff_A_NDct26XZ8_1),.doutc(w_dff_A_zzA9gOhC2_2),.din(n354));
	jspl jspl_w_n354_1(.douta(w_dff_A_uEuoVxFA7_0),.doutb(w_n354_1[1]),.din(w_n354_0[0]));
	jspl jspl_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.din(n355));
	jspl3 jspl3_w_n356_0(.douta(w_n356_0[0]),.doutb(w_dff_A_LB2BJLy78_1),.doutc(w_dff_A_CwoR9y7N7_2),.din(n356));
	jspl jspl_w_n356_1(.douta(w_dff_A_Mi458JfJ5_0),.doutb(w_n356_1[1]),.din(w_n356_0[0]));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_dff_A_u0zShoW77_1),.din(n357));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl jspl_w_n367_1(.douta(w_n367_1[0]),.doutb(w_n367_1[1]),.din(w_n367_0[0]));
	jspl jspl_w_n370_0(.douta(w_dff_A_34WEawZK6_0),.doutb(w_n370_0[1]),.din(w_dff_B_gHQTSLrz0_2));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl jspl_w_n378_0(.douta(w_dff_A_pgfK9uma1_0),.doutb(w_n378_0[1]),.din(n378));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_dff_A_PSySrwr68_1),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl3 jspl3_w_n388_0(.douta(w_dff_A_hvqDGvPG2_0),.doutb(w_dff_A_5ZUteJJl5_1),.doutc(w_n388_0[2]),.din(n388));
	jspl3 jspl3_w_n388_1(.douta(w_n388_1[0]),.doutb(w_dff_A_ONNWueaN8_1),.doutc(w_dff_A_JoHpLu1U0_2),.din(w_n388_0[0]));
	jspl jspl_w_n388_2(.douta(w_n388_2[0]),.doutb(w_dff_A_LR5W7OFQ5_1),.din(w_n388_0[1]));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n395_0(.douta(w_dff_A_YTi8Dgu26_0),.doutb(w_n395_0[1]),.din(n395));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_dff_A_xc49V2yN9_1),.din(n407));
	jspl3 jspl3_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.doutc(w_n414_0[2]),.din(n414));
	jspl3 jspl3_w_n417_0(.douta(w_n417_0[0]),.doutb(w_dff_A_Oh91G41R4_1),.doutc(w_dff_A_SKxkA4gY1_2),.din(n417));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_dff_A_FcdkyXoc5_1),.din(n420));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl jspl_w_n428_0(.douta(w_dff_A_UbfmXpYv9_0),.doutb(w_n428_0[1]),.din(n428));
	jspl jspl_w_n430_0(.douta(w_dff_A_Cqut5Hol2_0),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_dff_A_Zh3LZqwt0_1),.din(n435));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.doutc(w_n439_0[2]),.din(n439));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n450_0(.douta(w_dff_A_NLrLty692_0),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_dff_A_n48ZFbuf3_1),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl jspl_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.din(n473));
	jspl3 jspl3_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.doutc(w_n482_0[2]),.din(n482));
	jspl jspl_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n494_0(.douta(w_dff_A_uPxZXOvn9_0),.doutb(w_n494_0[1]),.din(n494));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_dff_A_I33LFH801_1),.din(n499));
	jspl jspl_w_n500_0(.douta(w_n500_0[0]),.doutb(w_n500_0[1]),.din(n500));
	jspl3 jspl3_w_n503_0(.douta(w_n503_0[0]),.doutb(w_dff_A_W5Ogq3VP7_1),.doutc(w_n503_0[2]),.din(n503));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_dff_A_qdkzIen67_1),.doutc(w_dff_A_kt9eReKY6_2),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_dff_A_EdOHaFaB2_0),.doutb(w_dff_A_HegGS2qX4_1),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl jspl_w_n507_2(.douta(w_n507_2[0]),.doutb(w_dff_A_V6jSsjcw7_1),.din(w_n507_0[1]));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl jspl_w_n512_0(.douta(w_dff_A_vSDsysS30_0),.doutb(w_n512_0[1]),.din(n512));
	jspl3 jspl3_w_n514_0(.douta(w_n514_0[0]),.doutb(w_dff_A_YS7cNnUb6_1),.doutc(w_dff_A_6ypzyubQ1_2),.din(n514));
	jspl jspl_w_n514_1(.douta(w_dff_A_obDpq9Wc4_0),.doutb(w_n514_1[1]),.din(w_n514_0[0]));
	jspl jspl_w_n520_0(.douta(w_dff_A_SqJOrxYE3_0),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_dff_A_Gm4CyLtF8_1),.din(n534));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_dff_A_fFhQYuH08_1),.din(n548));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_n559_0[1]),.din(n559));
	jspl jspl_w_n562_0(.douta(w_dff_A_Vep6fdi22_0),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_dff_A_az5jMjMD1_1),.doutc(w_dff_A_00kALzpj4_2),.din(n566));
	jspl jspl_w_n566_1(.douta(w_n566_1[0]),.doutb(w_n566_1[1]),.din(w_n566_0[0]));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_dff_A_AaWsLxke0_1),.doutc(w_dff_A_MzwhkeoN1_2),.din(n567));
	jspl3 jspl3_w_n567_1(.douta(w_dff_A_H10i0gnZ4_0),.doutb(w_n567_1[1]),.doutc(w_dff_A_hqzJ7BUz0_2),.din(w_n567_0[0]));
	jspl3 jspl3_w_n567_2(.douta(w_n567_2[0]),.doutb(w_n567_2[1]),.doutc(w_dff_A_RsAMSWpq3_2),.din(w_n567_0[1]));
	jspl3 jspl3_w_n567_3(.douta(w_dff_A_sdMQGsvz6_0),.doutb(w_dff_A_dTjGelrD5_1),.doutc(w_n567_3[2]),.din(w_n567_0[2]));
	jspl3 jspl3_w_n567_4(.douta(w_dff_A_6TImLwIf6_0),.doutb(w_n567_4[1]),.doutc(w_n567_4[2]),.din(w_n567_1[0]));
	jspl jspl_w_n567_5(.douta(w_n567_5[0]),.doutb(w_dff_A_fRorsgP65_1),.din(w_n567_1[1]));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_dff_A_WfzRtcFC0_1),.din(n569));
	jspl jspl_w_n570_0(.douta(w_dff_A_b8cO9g9e4_0),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_dff_A_0YNUmbHB5_1),.doutc(w_dff_A_tA6eYaIu4_2),.din(w_dff_B_fj0fuCCv9_3));
	jspl3 jspl3_w_n571_1(.douta(w_n571_1[0]),.doutb(w_dff_A_UDYrwmQr2_1),.doutc(w_n571_1[2]),.din(w_n571_0[0]));
	jspl jspl_w_n571_2(.douta(w_dff_A_ubAFFJDR1_0),.doutb(w_n571_2[1]),.din(w_n571_0[1]));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl jspl_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.din(n573));
	jspl jspl_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.din(n574));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n577_0(.douta(w_dff_A_f3ju7Xvn3_0),.doutb(w_n577_0[1]),.din(n577));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.doutc(w_dff_A_4EkeUj953_2),.din(n579));
	jspl jspl_w_n579_1(.douta(w_n579_1[0]),.doutb(w_dff_A_nBTj7VM28_1),.din(w_n579_0[0]));
	jspl3 jspl3_w_n580_0(.douta(w_n580_0[0]),.doutb(w_n580_0[1]),.doutc(w_n580_0[2]),.din(n580));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl jspl_w_n598_0(.douta(w_dff_A_mGCpcx5X1_0),.doutb(w_n598_0[1]),.din(n598));
	jspl3 jspl3_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.doutc(w_n600_0[2]),.din(n600));
	jspl3 jspl3_w_n600_1(.douta(w_dff_A_rV0vbByL7_0),.doutb(w_dff_A_wN72twRj6_1),.doutc(w_n600_1[2]),.din(w_n600_0[0]));
	jspl3 jspl3_w_n601_0(.douta(w_n601_0[0]),.doutb(w_dff_A_GsUCtSeh1_1),.doutc(w_n601_0[2]),.din(n601));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n604_0(.douta(w_dff_A_0NHp2NW70_0),.doutb(w_n604_0[1]),.doutc(w_dff_A_guTVlD6N5_2),.din(n604));
	jspl3 jspl3_w_n604_1(.douta(w_dff_A_q04uKjDl0_0),.doutb(w_dff_A_VK0Jemwn8_1),.doutc(w_n604_1[2]),.din(w_n604_0[0]));
	jspl3 jspl3_w_n604_2(.douta(w_dff_A_InXusHiD4_0),.doutb(w_n604_2[1]),.doutc(w_n604_2[2]),.din(w_n604_0[1]));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_dff_A_e63nU98t4_1),.doutc(w_dff_A_qEGBsBzK4_2),.din(w_dff_B_ZKL3QDgj6_3));
	jspl3 jspl3_w_n613_1(.douta(w_dff_A_WPwKHGLe3_0),.doutb(w_dff_A_zKqqXszk4_1),.doutc(w_n613_1[2]),.din(w_n613_0[0]));
	jspl3 jspl3_w_n614_0(.douta(w_n614_0[0]),.doutb(w_dff_A_TQSST8xv0_1),.doutc(w_dff_A_pMifdcYw3_2),.din(n614));
	jspl3 jspl3_w_n614_1(.douta(w_dff_A_ax2aeJKe0_0),.doutb(w_n614_1[1]),.doutc(w_dff_A_OF6GhCY34_2),.din(w_n614_0[0]));
	jspl3 jspl3_w_n614_2(.douta(w_dff_A_peMkkoOB8_0),.doutb(w_dff_A_gps9NreM1_1),.doutc(w_n614_2[2]),.din(w_n614_0[1]));
	jspl3 jspl3_w_n614_3(.douta(w_n614_3[0]),.doutb(w_dff_A_uhmDajlO9_1),.doutc(w_dff_A_XOHknlG88_2),.din(w_n614_0[2]));
	jspl3 jspl3_w_n614_4(.douta(w_n614_4[0]),.doutb(w_dff_A_aBqoN1gC4_1),.doutc(w_dff_A_VZajrdVB7_2),.din(w_n614_1[0]));
	jspl jspl_w_n614_5(.douta(w_dff_A_uHCxWV2a9_0),.doutb(w_n614_5[1]),.din(w_n614_1[1]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_dff_A_V5rlJOz46_2),.din(n618));
	jspl3 jspl3_w_n618_1(.douta(w_dff_A_vp9rvH7c9_0),.doutb(w_dff_A_om1uan588_1),.doutc(w_n618_1[2]),.din(w_n618_0[0]));
	jspl jspl_w_n618_2(.douta(w_dff_A_8kOfjuPP0_0),.doutb(w_n618_2[1]),.din(w_n618_0[1]));
	jspl3 jspl3_w_n619_0(.douta(w_dff_A_gUS2zuK58_0),.doutb(w_dff_A_pRUa8Ttq1_1),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n620_0(.douta(w_dff_A_cLTLoYju5_0),.doutb(w_n620_0[1]),.doutc(w_dff_A_M3oKymkX0_2),.din(n620));
	jspl jspl_w_n622_0(.douta(w_dff_A_LNnhatrx2_0),.doutb(w_n622_0[1]),.din(n622));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl3 jspl3_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.doutc(w_n626_0[2]),.din(n626));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(n628));
	jspl3 jspl3_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.doutc(w_n629_0[2]),.din(n629));
	jspl3 jspl3_w_n629_1(.douta(w_n629_1[0]),.doutb(w_n629_1[1]),.doutc(w_n629_1[2]),.din(w_n629_0[0]));
	jspl3 jspl3_w_n629_2(.douta(w_n629_2[0]),.doutb(w_n629_2[1]),.doutc(w_n629_2[2]),.din(w_n629_0[1]));
	jspl3 jspl3_w_n629_3(.douta(w_n629_3[0]),.doutb(w_n629_3[1]),.doutc(w_n629_3[2]),.din(w_n629_0[2]));
	jspl3 jspl3_w_n629_4(.douta(w_n629_4[0]),.doutb(w_n629_4[1]),.doutc(w_n629_4[2]),.din(w_n629_1[0]));
	jspl jspl_w_n629_5(.douta(w_n629_5[0]),.doutb(w_n629_5[1]),.din(w_n629_1[1]));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl3 jspl3_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.doutc(w_n633_0[2]),.din(n633));
	jspl3 jspl3_w_n633_1(.douta(w_n633_1[0]),.doutb(w_n633_1[1]),.doutc(w_n633_1[2]),.din(w_n633_0[0]));
	jspl3 jspl3_w_n633_2(.douta(w_n633_2[0]),.doutb(w_n633_2[1]),.doutc(w_n633_2[2]),.din(w_n633_0[1]));
	jspl3 jspl3_w_n633_3(.douta(w_n633_3[0]),.doutb(w_n633_3[1]),.doutc(w_n633_3[2]),.din(w_n633_0[2]));
	jspl3 jspl3_w_n633_4(.douta(w_n633_4[0]),.doutb(w_n633_4[1]),.doutc(w_n633_4[2]),.din(w_n633_1[0]));
	jspl3 jspl3_w_n633_5(.douta(w_n633_5[0]),.doutb(w_n633_5[1]),.doutc(w_n633_5[2]),.din(w_n633_1[1]));
	jspl jspl_w_n633_6(.douta(w_n633_6[0]),.doutb(w_n633_6[1]),.din(w_n633_1[2]));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(n637));
	jspl3 jspl3_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.doutc(w_n638_0[2]),.din(n638));
	jspl3 jspl3_w_n638_1(.douta(w_n638_1[0]),.doutb(w_n638_1[1]),.doutc(w_n638_1[2]),.din(w_n638_0[0]));
	jspl3 jspl3_w_n638_2(.douta(w_n638_2[0]),.doutb(w_n638_2[1]),.doutc(w_n638_2[2]),.din(w_n638_0[1]));
	jspl3 jspl3_w_n638_3(.douta(w_n638_3[0]),.doutb(w_n638_3[1]),.doutc(w_n638_3[2]),.din(w_n638_0[2]));
	jspl3 jspl3_w_n638_4(.douta(w_n638_4[0]),.doutb(w_n638_4[1]),.doutc(w_n638_4[2]),.din(w_n638_1[0]));
	jspl3 jspl3_w_n638_5(.douta(w_n638_5[0]),.doutb(w_n638_5[1]),.doutc(w_n638_5[2]),.din(w_n638_1[1]));
	jspl3 jspl3_w_n638_6(.douta(w_n638_6[0]),.doutb(w_n638_6[1]),.doutc(w_n638_6[2]),.din(w_n638_1[2]));
	jspl jspl_w_n638_7(.douta(w_n638_7[0]),.doutb(w_n638_7[1]),.din(w_n638_2[0]));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl3 jspl3_w_n640_2(.douta(w_n640_2[0]),.doutb(w_n640_2[1]),.doutc(w_n640_2[2]),.din(w_n640_0[1]));
	jspl3 jspl3_w_n640_3(.douta(w_n640_3[0]),.doutb(w_n640_3[1]),.doutc(w_n640_3[2]),.din(w_n640_0[2]));
	jspl3 jspl3_w_n640_4(.douta(w_n640_4[0]),.doutb(w_n640_4[1]),.doutc(w_n640_4[2]),.din(w_n640_1[0]));
	jspl3 jspl3_w_n640_5(.douta(w_n640_5[0]),.doutb(w_n640_5[1]),.doutc(w_n640_5[2]),.din(w_n640_1[1]));
	jspl3 jspl3_w_n640_6(.douta(w_n640_6[0]),.doutb(w_n640_6[1]),.doutc(w_n640_6[2]),.din(w_n640_1[2]));
	jspl jspl_w_n640_7(.douta(w_n640_7[0]),.doutb(w_n640_7[1]),.din(w_n640_2[0]));
	jspl3 jspl3_w_n646_0(.douta(w_n646_0[0]),.doutb(w_n646_0[1]),.doutc(w_n646_0[2]),.din(n646));
	jspl3 jspl3_w_n646_1(.douta(w_n646_1[0]),.doutb(w_n646_1[1]),.doutc(w_n646_1[2]),.din(w_n646_0[0]));
	jspl3 jspl3_w_n646_2(.douta(w_n646_2[0]),.doutb(w_n646_2[1]),.doutc(w_n646_2[2]),.din(w_n646_0[1]));
	jspl3 jspl3_w_n646_3(.douta(w_n646_3[0]),.doutb(w_n646_3[1]),.doutc(w_n646_3[2]),.din(w_n646_0[2]));
	jspl3 jspl3_w_n646_4(.douta(w_n646_4[0]),.doutb(w_n646_4[1]),.doutc(w_n646_4[2]),.din(w_n646_1[0]));
	jspl3 jspl3_w_n646_5(.douta(w_n646_5[0]),.doutb(w_n646_5[1]),.doutc(w_n646_5[2]),.din(w_n646_1[1]));
	jspl3 jspl3_w_n646_6(.douta(w_n646_6[0]),.doutb(w_n646_6[1]),.doutc(w_n646_6[2]),.din(w_n646_1[2]));
	jspl jspl_w_n646_7(.douta(w_n646_7[0]),.doutb(w_n646_7[1]),.din(w_n646_2[0]));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.doutc(w_n648_0[2]),.din(n648));
	jspl3 jspl3_w_n648_1(.douta(w_n648_1[0]),.doutb(w_n648_1[1]),.doutc(w_n648_1[2]),.din(w_n648_0[0]));
	jspl3 jspl3_w_n648_2(.douta(w_n648_2[0]),.doutb(w_n648_2[1]),.doutc(w_n648_2[2]),.din(w_n648_0[1]));
	jspl3 jspl3_w_n648_3(.douta(w_n648_3[0]),.doutb(w_n648_3[1]),.doutc(w_n648_3[2]),.din(w_n648_0[2]));
	jspl jspl_w_n648_4(.douta(w_n648_4[0]),.doutb(w_n648_4[1]),.din(w_n648_1[0]));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_dff_A_BaM0tXbx0_1),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.doutc(w_n651_0[2]),.din(n651));
	jspl3 jspl3_w_n651_1(.douta(w_n651_1[0]),.doutb(w_n651_1[1]),.doutc(w_n651_1[2]),.din(w_n651_0[0]));
	jspl3 jspl3_w_n651_2(.douta(w_n651_2[0]),.doutb(w_n651_2[1]),.doutc(w_n651_2[2]),.din(w_n651_0[1]));
	jspl3 jspl3_w_n651_3(.douta(w_n651_3[0]),.doutb(w_n651_3[1]),.doutc(w_n651_3[2]),.din(w_n651_0[2]));
	jspl3 jspl3_w_n651_4(.douta(w_n651_4[0]),.doutb(w_n651_4[1]),.doutc(w_n651_4[2]),.din(w_n651_1[0]));
	jspl3 jspl3_w_n651_5(.douta(w_n651_5[0]),.doutb(w_n651_5[1]),.doutc(w_n651_5[2]),.din(w_n651_1[1]));
	jspl3 jspl3_w_n651_6(.douta(w_n651_6[0]),.doutb(w_n651_6[1]),.doutc(w_n651_6[2]),.din(w_n651_1[2]));
	jspl jspl_w_n651_7(.douta(w_n651_7[0]),.doutb(w_n651_7[1]),.din(w_n651_2[0]));
	jspl3 jspl3_w_n653_0(.douta(w_n653_0[0]),.doutb(w_n653_0[1]),.doutc(w_n653_0[2]),.din(n653));
	jspl3 jspl3_w_n653_1(.douta(w_n653_1[0]),.doutb(w_n653_1[1]),.doutc(w_n653_1[2]),.din(w_n653_0[0]));
	jspl3 jspl3_w_n653_2(.douta(w_n653_2[0]),.doutb(w_n653_2[1]),.doutc(w_n653_2[2]),.din(w_n653_0[1]));
	jspl3 jspl3_w_n653_3(.douta(w_n653_3[0]),.doutb(w_n653_3[1]),.doutc(w_n653_3[2]),.din(w_n653_0[2]));
	jspl3 jspl3_w_n653_4(.douta(w_n653_4[0]),.doutb(w_n653_4[1]),.doutc(w_n653_4[2]),.din(w_n653_1[0]));
	jspl3 jspl3_w_n653_5(.douta(w_n653_5[0]),.doutb(w_n653_5[1]),.doutc(w_n653_5[2]),.din(w_n653_1[1]));
	jspl3 jspl3_w_n653_6(.douta(w_n653_6[0]),.doutb(w_n653_6[1]),.doutc(w_n653_6[2]),.din(w_n653_1[2]));
	jspl jspl_w_n653_7(.douta(w_n653_7[0]),.doutb(w_n653_7[1]),.din(w_n653_2[0]));
	jspl3 jspl3_w_n680_0(.douta(w_n680_0[0]),.doutb(w_dff_A_sQCRFlbg1_1),.doutc(w_n680_0[2]),.din(n680));
	jspl3 jspl3_w_n680_1(.douta(w_n680_1[0]),.doutb(w_dff_A_AieAZqdi9_1),.doutc(w_n680_1[2]),.din(w_n680_0[0]));
	jspl3 jspl3_w_n680_2(.douta(w_dff_A_U5NGfB3C5_0),.doutb(w_n680_2[1]),.doutc(w_dff_A_mQ5PH6K54_2),.din(w_n680_0[1]));
	jspl3 jspl3_w_n680_3(.douta(w_dff_A_GbYdWwlj5_0),.doutb(w_n680_3[1]),.doutc(w_dff_A_JmyOfB7B1_2),.din(w_n680_0[2]));
	jspl jspl_w_n680_4(.douta(w_n680_4[0]),.doutb(w_dff_A_wVzkdJBF7_1),.din(w_n680_1[0]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_dff_A_sHAus9Hg6_1),.din(n682));
	jspl3 jspl3_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.doutc(w_n684_0[2]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl3 jspl3_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.doutc(w_n690_0[2]),.din(n690));
	jspl jspl_w_n690_1(.douta(w_n690_1[0]),.doutb(w_n690_1[1]),.din(w_n690_0[0]));
	jspl jspl_w_n692_0(.douta(w_dff_A_Icil9oyk6_0),.doutb(w_n692_0[1]),.din(n692));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_dff_A_ByPGuawY7_1),.doutc(w_dff_A_qHvtVqkT7_2),.din(n703));
	jspl jspl_w_n703_1(.douta(w_dff_A_iOdcPdRN2_0),.doutb(w_n703_1[1]),.din(w_n703_0[0]));
	jspl jspl_w_n704_0(.douta(w_dff_A_JH3Amltv7_0),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n718_0(.douta(w_dff_A_tpD3wjjN6_0),.doutb(w_n718_0[1]),.din(w_dff_B_5UdxwxRG3_2));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n741_1(.douta(w_n741_1[0]),.doutb(w_n741_1[1]),.din(w_n741_0[0]));
	jspl jspl_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.din(n748));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl jspl_w_n759_0(.douta(w_dff_A_akZQpuOp2_0),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n766_0(.douta(w_n766_0[0]),.doutb(w_n766_0[1]),.din(n766));
	jspl3 jspl3_w_n767_0(.douta(w_n767_0[0]),.doutb(w_dff_A_Ney4EExm3_1),.doutc(w_dff_A_z0M12BCP9_2),.din(w_dff_B_p5X6eS3F5_3));
	jspl jspl_w_n767_1(.douta(w_n767_1[0]),.doutb(w_dff_A_JEo4JplL4_1),.din(w_n767_0[0]));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_dff_A_TJwIehfe4_2),.din(n771));
	jspl jspl_w_n771_1(.douta(w_dff_A_EPTeD56R1_0),.doutb(w_n771_1[1]),.din(w_n771_0[0]));
	jspl jspl_w_n772_0(.douta(w_dff_A_Z55c4btw4_0),.doutb(w_n772_0[1]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_dff_A_vvtvW8iE0_1),.din(n773));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n798_0(.douta(w_dff_A_NWjxawI12_0),.doutb(w_n798_0[1]),.din(n798));
	jspl3 jspl3_w_n802_0(.douta(w_n802_0[0]),.doutb(w_dff_A_eiDE24Oq2_1),.doutc(w_n802_0[2]),.din(n802));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_dff_A_jZ8bFWoo9_1),.din(n817));
	jspl jspl_w_n830_0(.douta(w_n830_0[0]),.doutb(w_n830_0[1]),.din(n830));
	jspl jspl_w_n833_0(.douta(w_dff_A_1gSwhNQf5_0),.doutb(w_n833_0[1]),.din(n833));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_dff_A_OG8upKwM1_1),.doutc(w_n845_0[2]),.din(n845));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl jspl_w_n861_0(.douta(w_dff_A_lk2PBJq41_0),.doutb(w_n861_0[1]),.din(n861));
	jspl3 jspl3_w_n863_0(.douta(w_dff_A_lbuSIHpA8_0),.doutb(w_n863_0[1]),.doutc(w_dff_A_gfTtQOA63_2),.din(n863));
	jspl3 jspl3_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.doutc(w_n869_0[2]),.din(n869));
	jspl jspl_w_n873_0(.douta(w_n873_0[0]),.doutb(w_n873_0[1]),.din(n873));
	jspl jspl_w_n875_0(.douta(w_n875_0[0]),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_dff_A_xR7b1os08_1),.din(n887));
	jspl3 jspl3_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.doutc(w_n937_0[2]),.din(n937));
	jspl jspl_w_n959_0(.douta(w_dff_A_AvSlXyCe7_0),.doutb(w_n959_0[1]),.din(n959));
	jspl3 jspl3_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.doutc(w_n987_0[2]),.din(n987));
	jspl3 jspl3_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.doutc(w_n1029_0[2]),.din(n1029));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1036_0(.douta(w_n1036_0[0]),.doutb(w_n1036_0[1]),.din(n1036));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.din(n1039));
	jspl jspl_w_n1040_0(.douta(w_n1040_0[0]),.doutb(w_n1040_0[1]),.din(n1040));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_dff_A_pXjCxg399_1),.din(n1043));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(n1044));
	jspl jspl_w_n1045_0(.douta(w_n1045_0[0]),.doutb(w_dff_A_qSzqW1xY9_1),.din(n1045));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(n1048));
	jspl3 jspl3_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.doutc(w_n1053_0[2]),.din(n1053));
	jspl jspl_w_n1056_0(.douta(w_dff_A_VvKWeSn83_0),.doutb(w_n1056_0[1]),.din(w_dff_B_IF4NufHq0_2));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_dff_A_NvbC047F9_1),.din(n1062));
	jspl jspl_w_n1091_0(.douta(w_dff_A_0yyXrzMH2_0),.doutb(w_n1091_0[1]),.din(n1091));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl3 jspl3_w_n1159_0(.douta(w_n1159_0[0]),.doutb(w_n1159_0[1]),.doutc(w_n1159_0[2]),.din(n1159));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_dff_A_NlX6DN6V3_1),.din(n1161));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(w_dff_B_W7UKalJt1_2));
	jspl jspl_w_n1168_0(.douta(w_n1168_0[0]),.doutb(w_n1168_0[1]),.din(n1168));
	jspl jspl_w_n1170_0(.douta(w_n1170_0[0]),.doutb(w_dff_A_WWo1OGan9_1),.din(n1170));
	jspl jspl_w_n1177_0(.douta(w_n1177_0[0]),.doutb(w_dff_A_Lz3Y5PGp7_1),.din(w_dff_B_Dq2Xk9Zs5_2));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_dff_A_cebzNpmp2_1),.din(n1178));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.din(n1184));
	jdff dff_B_ynZ5YnHd1_1(.din(n92),.dout(w_dff_B_ynZ5YnHd1_1),.clk(gclk));
	jdff dff_B_xrbgYCPy3_1(.din(w_dff_B_ynZ5YnHd1_1),.dout(w_dff_B_xrbgYCPy3_1),.clk(gclk));
	jdff dff_B_Pb9h1aHH6_1(.din(w_dff_B_xrbgYCPy3_1),.dout(w_dff_B_Pb9h1aHH6_1),.clk(gclk));
	jdff dff_B_q71j2OGx8_0(.din(n114),.dout(w_dff_B_q71j2OGx8_0),.clk(gclk));
	jdff dff_B_udMr7RwF5_0(.din(n109),.dout(w_dff_B_udMr7RwF5_0),.clk(gclk));
	jdff dff_B_9z3KwyPI0_1(.din(n93),.dout(w_dff_B_9z3KwyPI0_1),.clk(gclk));
	jdff dff_B_hbZGDMrg3_1(.din(w_dff_B_9z3KwyPI0_1),.dout(w_dff_B_hbZGDMrg3_1),.clk(gclk));
	jdff dff_B_zCONiVVC8_0(.din(n100),.dout(w_dff_B_zCONiVVC8_0),.clk(gclk));
	jdff dff_B_WG4S1uzv0_1(.din(n583),.dout(w_dff_B_WG4S1uzv0_1),.clk(gclk));
	jdff dff_B_e4hfOEbK7_1(.din(w_dff_B_WG4S1uzv0_1),.dout(w_dff_B_e4hfOEbK7_1),.clk(gclk));
	jdff dff_B_ZbTG51FI0_1(.din(w_dff_B_e4hfOEbK7_1),.dout(w_dff_B_ZbTG51FI0_1),.clk(gclk));
	jdff dff_B_t6YLDsJf6_1(.din(w_dff_B_ZbTG51FI0_1),.dout(w_dff_B_t6YLDsJf6_1),.clk(gclk));
	jdff dff_B_JHWAjE433_1(.din(w_dff_B_t6YLDsJf6_1),.dout(w_dff_B_JHWAjE433_1),.clk(gclk));
	jdff dff_B_Ws5GYjEw0_1(.din(w_dff_B_JHWAjE433_1),.dout(w_dff_B_Ws5GYjEw0_1),.clk(gclk));
	jdff dff_B_xB1RSBq43_1(.din(w_dff_B_Ws5GYjEw0_1),.dout(w_dff_B_xB1RSBq43_1),.clk(gclk));
	jdff dff_B_rpt2txpk2_1(.din(w_dff_B_xB1RSBq43_1),.dout(w_dff_B_rpt2txpk2_1),.clk(gclk));
	jdff dff_B_CXcfAsYh9_1(.din(w_dff_B_rpt2txpk2_1),.dout(w_dff_B_CXcfAsYh9_1),.clk(gclk));
	jdff dff_B_8FKXV26O9_1(.din(w_dff_B_CXcfAsYh9_1),.dout(w_dff_B_8FKXV26O9_1),.clk(gclk));
	jdff dff_B_N9BGqFE76_1(.din(w_dff_B_8FKXV26O9_1),.dout(w_dff_B_N9BGqFE76_1),.clk(gclk));
	jdff dff_B_VtB1sIV48_1(.din(w_dff_B_N9BGqFE76_1),.dout(w_dff_B_VtB1sIV48_1),.clk(gclk));
	jdff dff_B_mL75RmLX6_1(.din(w_dff_B_VtB1sIV48_1),.dout(w_dff_B_mL75RmLX6_1),.clk(gclk));
	jdff dff_B_N6Lw2OXO1_1(.din(w_dff_B_mL75RmLX6_1),.dout(w_dff_B_N6Lw2OXO1_1),.clk(gclk));
	jdff dff_B_S51GjHWv7_1(.din(w_dff_B_N6Lw2OXO1_1),.dout(w_dff_B_S51GjHWv7_1),.clk(gclk));
	jdff dff_B_prADZb7W6_1(.din(w_dff_B_S51GjHWv7_1),.dout(w_dff_B_prADZb7W6_1),.clk(gclk));
	jdff dff_B_fHOwcBxf0_0(.din(n607),.dout(w_dff_B_fHOwcBxf0_0),.clk(gclk));
	jdff dff_B_Jvtvvq538_0(.din(w_dff_B_fHOwcBxf0_0),.dout(w_dff_B_Jvtvvq538_0),.clk(gclk));
	jdff dff_B_3M27IcLs1_0(.din(w_dff_B_Jvtvvq538_0),.dout(w_dff_B_3M27IcLs1_0),.clk(gclk));
	jdff dff_B_I7gb4k2j7_0(.din(w_dff_B_3M27IcLs1_0),.dout(w_dff_B_I7gb4k2j7_0),.clk(gclk));
	jdff dff_B_Q0OU1C3u7_0(.din(w_dff_B_I7gb4k2j7_0),.dout(w_dff_B_Q0OU1C3u7_0),.clk(gclk));
	jdff dff_B_cFVEODNb8_0(.din(w_dff_B_Q0OU1C3u7_0),.dout(w_dff_B_cFVEODNb8_0),.clk(gclk));
	jdff dff_B_jOwdAJi95_0(.din(w_dff_B_cFVEODNb8_0),.dout(w_dff_B_jOwdAJi95_0),.clk(gclk));
	jdff dff_B_1m3mqAGi7_0(.din(w_dff_B_jOwdAJi95_0),.dout(w_dff_B_1m3mqAGi7_0),.clk(gclk));
	jdff dff_B_jnU9okez8_0(.din(w_dff_B_1m3mqAGi7_0),.dout(w_dff_B_jnU9okez8_0),.clk(gclk));
	jdff dff_B_oyimtRpZ0_0(.din(w_dff_B_jnU9okez8_0),.dout(w_dff_B_oyimtRpZ0_0),.clk(gclk));
	jdff dff_B_EAroxufK9_0(.din(w_dff_B_oyimtRpZ0_0),.dout(w_dff_B_EAroxufK9_0),.clk(gclk));
	jdff dff_B_0OMFfL6U4_0(.din(w_dff_B_EAroxufK9_0),.dout(w_dff_B_0OMFfL6U4_0),.clk(gclk));
	jdff dff_B_kUcR5PsM8_0(.din(w_dff_B_0OMFfL6U4_0),.dout(w_dff_B_kUcR5PsM8_0),.clk(gclk));
	jdff dff_B_mOPif1fF3_0(.din(w_dff_B_kUcR5PsM8_0),.dout(w_dff_B_mOPif1fF3_0),.clk(gclk));
	jdff dff_B_bLAKcHKe6_0(.din(n795),.dout(w_dff_B_bLAKcHKe6_0),.clk(gclk));
	jdff dff_B_SPiR5Gfq0_0(.din(w_dff_B_bLAKcHKe6_0),.dout(w_dff_B_SPiR5Gfq0_0),.clk(gclk));
	jdff dff_B_40lhxiL72_0(.din(w_dff_B_SPiR5Gfq0_0),.dout(w_dff_B_40lhxiL72_0),.clk(gclk));
	jdff dff_B_U7NvSjUt8_0(.din(w_dff_B_40lhxiL72_0),.dout(w_dff_B_U7NvSjUt8_0),.clk(gclk));
	jdff dff_B_c7m59G2O8_0(.din(w_dff_B_U7NvSjUt8_0),.dout(w_dff_B_c7m59G2O8_0),.clk(gclk));
	jdff dff_B_lUWwwYmu7_0(.din(w_dff_B_c7m59G2O8_0),.dout(w_dff_B_lUWwwYmu7_0),.clk(gclk));
	jdff dff_B_H9wIZlfo4_0(.din(w_dff_B_lUWwwYmu7_0),.dout(w_dff_B_H9wIZlfo4_0),.clk(gclk));
	jdff dff_B_1EC4mkL36_0(.din(w_dff_B_H9wIZlfo4_0),.dout(w_dff_B_1EC4mkL36_0),.clk(gclk));
	jdff dff_B_sNMgBzfb4_0(.din(w_dff_B_1EC4mkL36_0),.dout(w_dff_B_sNMgBzfb4_0),.clk(gclk));
	jdff dff_B_dYU2wWJk4_0(.din(w_dff_B_sNMgBzfb4_0),.dout(w_dff_B_dYU2wWJk4_0),.clk(gclk));
	jdff dff_B_KCoETwj26_0(.din(w_dff_B_dYU2wWJk4_0),.dout(w_dff_B_KCoETwj26_0),.clk(gclk));
	jdff dff_B_347UTkUS3_0(.din(w_dff_B_KCoETwj26_0),.dout(w_dff_B_347UTkUS3_0),.clk(gclk));
	jdff dff_B_6RgXlCOo7_0(.din(w_dff_B_347UTkUS3_0),.dout(w_dff_B_6RgXlCOo7_0),.clk(gclk));
	jdff dff_B_huhjNFeY1_0(.din(w_dff_B_6RgXlCOo7_0),.dout(w_dff_B_huhjNFeY1_0),.clk(gclk));
	jdff dff_B_1TU4w3Jl0_0(.din(w_dff_B_huhjNFeY1_0),.dout(w_dff_B_1TU4w3Jl0_0),.clk(gclk));
	jdff dff_B_fHVw0UMH6_0(.din(w_dff_B_1TU4w3Jl0_0),.dout(w_dff_B_fHVw0UMH6_0),.clk(gclk));
	jdff dff_B_eyzArHIQ3_0(.din(w_dff_B_fHVw0UMH6_0),.dout(w_dff_B_eyzArHIQ3_0),.clk(gclk));
	jdff dff_B_sq671Pcx0_0(.din(n794),.dout(w_dff_B_sq671Pcx0_0),.clk(gclk));
	jdff dff_A_rwvnvfyK3_1(.dout(w_n120_0[1]),.din(w_dff_A_rwvnvfyK3_1),.clk(gclk));
	jdff dff_A_Gv04fcjb4_1(.dout(w_dff_A_rwvnvfyK3_1),.din(w_dff_A_Gv04fcjb4_1),.clk(gclk));
	jdff dff_A_fqJ0YkIr5_1(.dout(w_dff_A_Gv04fcjb4_1),.din(w_dff_A_fqJ0YkIr5_1),.clk(gclk));
	jdff dff_B_AVjPnWhX9_0(.din(n791),.dout(w_dff_B_AVjPnWhX9_0),.clk(gclk));
	jdff dff_B_KpnIjPAZ5_1(.din(n762),.dout(w_dff_B_KpnIjPAZ5_1),.clk(gclk));
	jdff dff_B_TwPIIMOM4_1(.din(w_dff_B_KpnIjPAZ5_1),.dout(w_dff_B_TwPIIMOM4_1),.clk(gclk));
	jdff dff_B_cYnRrgGN4_1(.din(w_dff_B_TwPIIMOM4_1),.dout(w_dff_B_cYnRrgGN4_1),.clk(gclk));
	jdff dff_B_QsOWg22Z7_1(.din(w_dff_B_cYnRrgGN4_1),.dout(w_dff_B_QsOWg22Z7_1),.clk(gclk));
	jdff dff_B_9puWg91t9_1(.din(w_dff_B_QsOWg22Z7_1),.dout(w_dff_B_9puWg91t9_1),.clk(gclk));
	jdff dff_B_pdUogo6x0_1(.din(w_dff_B_9puWg91t9_1),.dout(w_dff_B_pdUogo6x0_1),.clk(gclk));
	jdff dff_B_7P58rKmj8_1(.din(w_dff_B_pdUogo6x0_1),.dout(w_dff_B_7P58rKmj8_1),.clk(gclk));
	jdff dff_B_k6DQEmqy0_1(.din(w_dff_B_7P58rKmj8_1),.dout(w_dff_B_k6DQEmqy0_1),.clk(gclk));
	jdff dff_B_KAQ6kGp86_1(.din(w_dff_B_k6DQEmqy0_1),.dout(w_dff_B_KAQ6kGp86_1),.clk(gclk));
	jdff dff_B_mfgfwltP7_1(.din(w_dff_B_KAQ6kGp86_1),.dout(w_dff_B_mfgfwltP7_1),.clk(gclk));
	jdff dff_B_IiyhBUHa3_1(.din(w_dff_B_mfgfwltP7_1),.dout(w_dff_B_IiyhBUHa3_1),.clk(gclk));
	jdff dff_B_xGeWlfHP1_1(.din(w_dff_B_IiyhBUHa3_1),.dout(w_dff_B_xGeWlfHP1_1),.clk(gclk));
	jdff dff_B_F7txf4wl7_1(.din(w_dff_B_xGeWlfHP1_1),.dout(w_dff_B_F7txf4wl7_1),.clk(gclk));
	jdff dff_B_FMWNkpb43_1(.din(w_dff_B_F7txf4wl7_1),.dout(w_dff_B_FMWNkpb43_1),.clk(gclk));
	jdff dff_B_rDYpXZLK3_1(.din(w_dff_B_FMWNkpb43_1),.dout(w_dff_B_rDYpXZLK3_1),.clk(gclk));
	jdff dff_B_F6XMW7zK9_1(.din(w_dff_B_rDYpXZLK3_1),.dout(w_dff_B_F6XMW7zK9_1),.clk(gclk));
	jdff dff_B_mCBbpt9J8_1(.din(w_dff_B_F6XMW7zK9_1),.dout(w_dff_B_mCBbpt9J8_1),.clk(gclk));
	jdff dff_B_mirvIYcZ8_1(.din(w_dff_B_mCBbpt9J8_1),.dout(w_dff_B_mirvIYcZ8_1),.clk(gclk));
	jdff dff_B_NNpb1PAP1_0(.din(n783),.dout(w_dff_B_NNpb1PAP1_0),.clk(gclk));
	jdff dff_A_VV0G5Xfi3_0(.dout(w_n112_0[0]),.din(w_dff_A_VV0G5Xfi3_0),.clk(gclk));
	jdff dff_B_MOGcl5UV4_1(.din(n1171),.dout(w_dff_B_MOGcl5UV4_1),.clk(gclk));
	jdff dff_B_pLHv3hyp7_1(.din(w_dff_B_MOGcl5UV4_1),.dout(w_dff_B_pLHv3hyp7_1),.clk(gclk));
	jdff dff_B_HfCFKUce9_1(.din(n1172),.dout(w_dff_B_HfCFKUce9_1),.clk(gclk));
	jdff dff_B_oUye4lm36_1(.din(w_dff_B_HfCFKUce9_1),.dout(w_dff_B_oUye4lm36_1),.clk(gclk));
	jdff dff_B_ccCmc88O3_1(.din(w_dff_B_oUye4lm36_1),.dout(w_dff_B_ccCmc88O3_1),.clk(gclk));
	jdff dff_B_Oyyhcu7R7_1(.din(w_dff_B_ccCmc88O3_1),.dout(w_dff_B_Oyyhcu7R7_1),.clk(gclk));
	jdff dff_B_3yH9xtxp0_1(.din(w_dff_B_Oyyhcu7R7_1),.dout(w_dff_B_3yH9xtxp0_1),.clk(gclk));
	jdff dff_B_fVa69rRd2_1(.din(w_dff_B_3yH9xtxp0_1),.dout(w_dff_B_fVa69rRd2_1),.clk(gclk));
	jdff dff_B_ISIuAwLU4_1(.din(w_dff_B_fVa69rRd2_1),.dout(w_dff_B_ISIuAwLU4_1),.clk(gclk));
	jdff dff_B_MiPcuc7d1_1(.din(w_dff_B_ISIuAwLU4_1),.dout(w_dff_B_MiPcuc7d1_1),.clk(gclk));
	jdff dff_B_i56ZNTFD4_1(.din(w_dff_B_MiPcuc7d1_1),.dout(w_dff_B_i56ZNTFD4_1),.clk(gclk));
	jdff dff_B_Yg9QwWVa5_1(.din(w_dff_B_i56ZNTFD4_1),.dout(w_dff_B_Yg9QwWVa5_1),.clk(gclk));
	jdff dff_B_uh65DdRn2_1(.din(w_dff_B_Yg9QwWVa5_1),.dout(w_dff_B_uh65DdRn2_1),.clk(gclk));
	jdff dff_B_lkpLCRPL1_1(.din(w_dff_B_uh65DdRn2_1),.dout(w_dff_B_lkpLCRPL1_1),.clk(gclk));
	jdff dff_B_OHSAB6HG1_1(.din(w_dff_B_lkpLCRPL1_1),.dout(w_dff_B_OHSAB6HG1_1),.clk(gclk));
	jdff dff_B_j1VOoZqi5_1(.din(w_dff_B_OHSAB6HG1_1),.dout(w_dff_B_j1VOoZqi5_1),.clk(gclk));
	jdff dff_B_LFokzkIg5_1(.din(w_dff_B_j1VOoZqi5_1),.dout(w_dff_B_LFokzkIg5_1),.clk(gclk));
	jdff dff_B_GcFzOQHz3_1(.din(w_dff_B_LFokzkIg5_1),.dout(w_dff_B_GcFzOQHz3_1),.clk(gclk));
	jdff dff_B_CP8Qiqn29_1(.din(w_dff_B_GcFzOQHz3_1),.dout(w_dff_B_CP8Qiqn29_1),.clk(gclk));
	jdff dff_B_ZhLnKxlj9_1(.din(w_dff_B_CP8Qiqn29_1),.dout(w_dff_B_ZhLnKxlj9_1),.clk(gclk));
	jdff dff_B_CE4hUIpS1_1(.din(w_dff_B_ZhLnKxlj9_1),.dout(w_dff_B_CE4hUIpS1_1),.clk(gclk));
	jdff dff_B_yqcq7O9G2_1(.din(w_dff_B_CE4hUIpS1_1),.dout(w_dff_B_yqcq7O9G2_1),.clk(gclk));
	jdff dff_B_FoniNyag2_1(.din(w_dff_B_yqcq7O9G2_1),.dout(w_dff_B_FoniNyag2_1),.clk(gclk));
	jdff dff_B_1tFGnpYG7_1(.din(w_dff_B_FoniNyag2_1),.dout(w_dff_B_1tFGnpYG7_1),.clk(gclk));
	jdff dff_B_iQ6wkzeT9_1(.din(w_dff_B_1tFGnpYG7_1),.dout(w_dff_B_iQ6wkzeT9_1),.clk(gclk));
	jdff dff_B_bFmJ5DuS4_1(.din(w_dff_B_iQ6wkzeT9_1),.dout(w_dff_B_bFmJ5DuS4_1),.clk(gclk));
	jdff dff_B_HkKtItOb4_1(.din(w_dff_B_bFmJ5DuS4_1),.dout(w_dff_B_HkKtItOb4_1),.clk(gclk));
	jdff dff_B_LvvcfnQ51_1(.din(w_dff_B_HkKtItOb4_1),.dout(w_dff_B_LvvcfnQ51_1),.clk(gclk));
	jdff dff_B_9RlCuJE84_1(.din(w_dff_B_LvvcfnQ51_1),.dout(w_dff_B_9RlCuJE84_1),.clk(gclk));
	jdff dff_B_jy3F7UiK7_1(.din(w_dff_B_9RlCuJE84_1),.dout(w_dff_B_jy3F7UiK7_1),.clk(gclk));
	jdff dff_B_NZyNgzld3_0(.din(n1166),.dout(w_dff_B_NZyNgzld3_0),.clk(gclk));
	jdff dff_B_HSI4VBVl1_0(.din(n1165),.dout(w_dff_B_HSI4VBVl1_0),.clk(gclk));
	jdff dff_A_NlX6DN6V3_1(.dout(w_n1161_0[1]),.din(w_dff_A_NlX6DN6V3_1),.clk(gclk));
	jdff dff_B_4Jva4wWJ7_1(.din(n1182),.dout(w_dff_B_4Jva4wWJ7_1),.clk(gclk));
	jdff dff_B_Yp126YZE0_1(.din(w_dff_B_4Jva4wWJ7_1),.dout(w_dff_B_Yp126YZE0_1),.clk(gclk));
	jdff dff_B_WjTJ54NR6_1(.din(w_dff_B_Yp126YZE0_1),.dout(w_dff_B_WjTJ54NR6_1),.clk(gclk));
	jdff dff_B_KxS9j7Ct8_1(.din(w_dff_B_WjTJ54NR6_1),.dout(w_dff_B_KxS9j7Ct8_1),.clk(gclk));
	jdff dff_B_ooJVhPtl4_1(.din(w_dff_B_KxS9j7Ct8_1),.dout(w_dff_B_ooJVhPtl4_1),.clk(gclk));
	jdff dff_B_Swa2GdbL7_1(.din(w_dff_B_ooJVhPtl4_1),.dout(w_dff_B_Swa2GdbL7_1),.clk(gclk));
	jdff dff_B_Gp7nP9S90_1(.din(w_dff_B_Swa2GdbL7_1),.dout(w_dff_B_Gp7nP9S90_1),.clk(gclk));
	jdff dff_B_XY1pnQ3s1_1(.din(w_dff_B_Gp7nP9S90_1),.dout(w_dff_B_XY1pnQ3s1_1),.clk(gclk));
	jdff dff_B_JRXFOd4X2_1(.din(w_dff_B_XY1pnQ3s1_1),.dout(w_dff_B_JRXFOd4X2_1),.clk(gclk));
	jdff dff_B_VWEfQuec5_1(.din(w_dff_B_JRXFOd4X2_1),.dout(w_dff_B_VWEfQuec5_1),.clk(gclk));
	jdff dff_B_hkHyVgjx6_1(.din(w_dff_B_VWEfQuec5_1),.dout(w_dff_B_hkHyVgjx6_1),.clk(gclk));
	jdff dff_B_ElenyalL8_1(.din(w_dff_B_hkHyVgjx6_1),.dout(w_dff_B_ElenyalL8_1),.clk(gclk));
	jdff dff_B_LL1UC17n5_1(.din(w_dff_B_ElenyalL8_1),.dout(w_dff_B_LL1UC17n5_1),.clk(gclk));
	jdff dff_B_onvbfAJl0_1(.din(w_dff_B_LL1UC17n5_1),.dout(w_dff_B_onvbfAJl0_1),.clk(gclk));
	jdff dff_B_7GqXLUBk4_1(.din(w_dff_B_onvbfAJl0_1),.dout(w_dff_B_7GqXLUBk4_1),.clk(gclk));
	jdff dff_B_TJrrlA0t2_1(.din(w_dff_B_7GqXLUBk4_1),.dout(w_dff_B_TJrrlA0t2_1),.clk(gclk));
	jdff dff_B_QJSsaXGL6_1(.din(w_dff_B_TJrrlA0t2_1),.dout(w_dff_B_QJSsaXGL6_1),.clk(gclk));
	jdff dff_B_AvtvG76D6_1(.din(w_dff_B_QJSsaXGL6_1),.dout(w_dff_B_AvtvG76D6_1),.clk(gclk));
	jdff dff_B_4YD8iW2l7_1(.din(w_dff_B_AvtvG76D6_1),.dout(w_dff_B_4YD8iW2l7_1),.clk(gclk));
	jdff dff_B_EZATfHu78_1(.din(w_dff_B_4YD8iW2l7_1),.dout(w_dff_B_EZATfHu78_1),.clk(gclk));
	jdff dff_B_rPPpTlqc4_1(.din(w_dff_B_EZATfHu78_1),.dout(w_dff_B_rPPpTlqc4_1),.clk(gclk));
	jdff dff_B_YTkb88oz0_1(.din(w_dff_B_rPPpTlqc4_1),.dout(w_dff_B_YTkb88oz0_1),.clk(gclk));
	jdff dff_B_hRMMJKQr8_1(.din(w_dff_B_YTkb88oz0_1),.dout(w_dff_B_hRMMJKQr8_1),.clk(gclk));
	jdff dff_B_0ug2eyZl8_1(.din(w_dff_B_hRMMJKQr8_1),.dout(w_dff_B_0ug2eyZl8_1),.clk(gclk));
	jdff dff_B_ep09lUf91_1(.din(w_dff_B_0ug2eyZl8_1),.dout(w_dff_B_ep09lUf91_1),.clk(gclk));
	jdff dff_B_tCTyTYsZ1_1(.din(G2897),.dout(w_dff_B_tCTyTYsZ1_1),.clk(gclk));
	jdff dff_B_nNZ0GruW3_1(.din(w_dff_B_tCTyTYsZ1_1),.dout(w_dff_B_nNZ0GruW3_1),.clk(gclk));
	jdff dff_B_Sb1jYBl36_1(.din(w_dff_B_nNZ0GruW3_1),.dout(w_dff_B_Sb1jYBl36_1),.clk(gclk));
	jdff dff_B_FoKlvykA8_1(.din(w_dff_B_Sb1jYBl36_1),.dout(w_dff_B_FoKlvykA8_1),.clk(gclk));
	jdff dff_B_92NfxHvE5_1(.din(w_dff_B_FoKlvykA8_1),.dout(w_dff_B_92NfxHvE5_1),.clk(gclk));
	jdff dff_B_akcrgVn10_1(.din(w_dff_B_92NfxHvE5_1),.dout(w_dff_B_akcrgVn10_1),.clk(gclk));
	jdff dff_B_LkkgUbfh9_1(.din(w_dff_B_akcrgVn10_1),.dout(w_dff_B_LkkgUbfh9_1),.clk(gclk));
	jdff dff_B_DdU91plB6_1(.din(w_dff_B_LkkgUbfh9_1),.dout(w_dff_B_DdU91plB6_1),.clk(gclk));
	jdff dff_B_NkrRuS4v6_1(.din(w_dff_B_DdU91plB6_1),.dout(w_dff_B_NkrRuS4v6_1),.clk(gclk));
	jdff dff_B_kGzofVkP0_1(.din(w_dff_B_NkrRuS4v6_1),.dout(w_dff_B_kGzofVkP0_1),.clk(gclk));
	jdff dff_B_FkDjUroM5_1(.din(w_dff_B_kGzofVkP0_1),.dout(w_dff_B_FkDjUroM5_1),.clk(gclk));
	jdff dff_B_a5qsdpPl0_1(.din(w_dff_B_FkDjUroM5_1),.dout(w_dff_B_a5qsdpPl0_1),.clk(gclk));
	jdff dff_B_geszqRin9_1(.din(w_dff_B_a5qsdpPl0_1),.dout(w_dff_B_geszqRin9_1),.clk(gclk));
	jdff dff_B_XPPkmska3_1(.din(w_dff_B_geszqRin9_1),.dout(w_dff_B_XPPkmska3_1),.clk(gclk));
	jdff dff_B_q6xrlLHy0_1(.din(w_dff_B_XPPkmska3_1),.dout(w_dff_B_q6xrlLHy0_1),.clk(gclk));
	jdff dff_B_u4YvyHno2_1(.din(w_dff_B_q6xrlLHy0_1),.dout(w_dff_B_u4YvyHno2_1),.clk(gclk));
	jdff dff_B_oiUAum5a2_1(.din(w_dff_B_u4YvyHno2_1),.dout(w_dff_B_oiUAum5a2_1),.clk(gclk));
	jdff dff_B_Dj4EA9br3_1(.din(w_dff_B_oiUAum5a2_1),.dout(w_dff_B_Dj4EA9br3_1),.clk(gclk));
	jdff dff_B_AVlSSToM7_1(.din(w_dff_B_Dj4EA9br3_1),.dout(w_dff_B_AVlSSToM7_1),.clk(gclk));
	jdff dff_B_2wh4DxzF3_1(.din(w_dff_B_AVlSSToM7_1),.dout(w_dff_B_2wh4DxzF3_1),.clk(gclk));
	jdff dff_B_kqcm35Et6_1(.din(w_dff_B_2wh4DxzF3_1),.dout(w_dff_B_kqcm35Et6_1),.clk(gclk));
	jdff dff_B_9Lneeevi3_1(.din(w_dff_B_kqcm35Et6_1),.dout(w_dff_B_9Lneeevi3_1),.clk(gclk));
	jdff dff_B_SccqQPVF0_1(.din(w_dff_B_9Lneeevi3_1),.dout(w_dff_B_SccqQPVF0_1),.clk(gclk));
	jdff dff_B_DpKEq05N3_1(.din(w_dff_B_SccqQPVF0_1),.dout(w_dff_B_DpKEq05N3_1),.clk(gclk));
	jdff dff_B_CkLQh78X3_1(.din(w_dff_B_DpKEq05N3_1),.dout(w_dff_B_CkLQh78X3_1),.clk(gclk));
	jdff dff_B_UM0Lkz9K1_1(.din(w_dff_B_CkLQh78X3_1),.dout(w_dff_B_UM0Lkz9K1_1),.clk(gclk));
	jdff dff_B_PsF3JsDJ6_1(.din(w_dff_B_UM0Lkz9K1_1),.dout(w_dff_B_PsF3JsDJ6_1),.clk(gclk));
	jdff dff_A_ILeDfsuw7_1(.dout(w_n1178_0[1]),.din(w_dff_A_ILeDfsuw7_1),.clk(gclk));
	jdff dff_A_pxawqQ3a3_1(.dout(w_dff_A_ILeDfsuw7_1),.din(w_dff_A_pxawqQ3a3_1),.clk(gclk));
	jdff dff_A_D2wsoZKF9_1(.dout(w_dff_A_pxawqQ3a3_1),.din(w_dff_A_D2wsoZKF9_1),.clk(gclk));
	jdff dff_A_Inn18rz07_1(.dout(w_dff_A_D2wsoZKF9_1),.din(w_dff_A_Inn18rz07_1),.clk(gclk));
	jdff dff_A_FXi9Q7wi5_1(.dout(w_dff_A_Inn18rz07_1),.din(w_dff_A_FXi9Q7wi5_1),.clk(gclk));
	jdff dff_A_AIxfc44U1_1(.dout(w_dff_A_FXi9Q7wi5_1),.din(w_dff_A_AIxfc44U1_1),.clk(gclk));
	jdff dff_A_iS0tUClF8_1(.dout(w_dff_A_AIxfc44U1_1),.din(w_dff_A_iS0tUClF8_1),.clk(gclk));
	jdff dff_A_OXTVixPV4_1(.dout(w_dff_A_iS0tUClF8_1),.din(w_dff_A_OXTVixPV4_1),.clk(gclk));
	jdff dff_A_kx9jF2yE1_1(.dout(w_dff_A_OXTVixPV4_1),.din(w_dff_A_kx9jF2yE1_1),.clk(gclk));
	jdff dff_A_f5EBb4x37_1(.dout(w_dff_A_kx9jF2yE1_1),.din(w_dff_A_f5EBb4x37_1),.clk(gclk));
	jdff dff_A_KaqR2Yu58_1(.dout(w_dff_A_f5EBb4x37_1),.din(w_dff_A_KaqR2Yu58_1),.clk(gclk));
	jdff dff_A_pEQqklk58_1(.dout(w_dff_A_KaqR2Yu58_1),.din(w_dff_A_pEQqklk58_1),.clk(gclk));
	jdff dff_A_PLmr5Ubr7_1(.dout(w_dff_A_pEQqklk58_1),.din(w_dff_A_PLmr5Ubr7_1),.clk(gclk));
	jdff dff_A_fApyZn363_1(.dout(w_dff_A_PLmr5Ubr7_1),.din(w_dff_A_fApyZn363_1),.clk(gclk));
	jdff dff_A_sTXFaWHj3_1(.dout(w_dff_A_fApyZn363_1),.din(w_dff_A_sTXFaWHj3_1),.clk(gclk));
	jdff dff_A_OmsWeqas0_1(.dout(w_dff_A_sTXFaWHj3_1),.din(w_dff_A_OmsWeqas0_1),.clk(gclk));
	jdff dff_A_KKksWgzY0_1(.dout(w_dff_A_OmsWeqas0_1),.din(w_dff_A_KKksWgzY0_1),.clk(gclk));
	jdff dff_A_hFSP9obF9_1(.dout(w_dff_A_KKksWgzY0_1),.din(w_dff_A_hFSP9obF9_1),.clk(gclk));
	jdff dff_A_YzSysODz5_1(.dout(w_dff_A_hFSP9obF9_1),.din(w_dff_A_YzSysODz5_1),.clk(gclk));
	jdff dff_A_YGXs8kLG2_1(.dout(w_dff_A_YzSysODz5_1),.din(w_dff_A_YGXs8kLG2_1),.clk(gclk));
	jdff dff_A_Q9MBdEoW4_1(.dout(w_dff_A_YGXs8kLG2_1),.din(w_dff_A_Q9MBdEoW4_1),.clk(gclk));
	jdff dff_A_oiDLfZe90_1(.dout(w_dff_A_Q9MBdEoW4_1),.din(w_dff_A_oiDLfZe90_1),.clk(gclk));
	jdff dff_A_FqziWXfs7_1(.dout(w_dff_A_oiDLfZe90_1),.din(w_dff_A_FqziWXfs7_1),.clk(gclk));
	jdff dff_A_ZZi18SpG5_1(.dout(w_dff_A_FqziWXfs7_1),.din(w_dff_A_ZZi18SpG5_1),.clk(gclk));
	jdff dff_A_HODbHNBK8_1(.dout(w_dff_A_ZZi18SpG5_1),.din(w_dff_A_HODbHNBK8_1),.clk(gclk));
	jdff dff_A_cebzNpmp2_1(.dout(w_dff_A_HODbHNBK8_1),.din(w_dff_A_cebzNpmp2_1),.clk(gclk));
	jdff dff_A_5IgX0xir6_1(.dout(w_n1170_0[1]),.din(w_dff_A_5IgX0xir6_1),.clk(gclk));
	jdff dff_A_vyPi09V38_1(.dout(w_dff_A_5IgX0xir6_1),.din(w_dff_A_vyPi09V38_1),.clk(gclk));
	jdff dff_A_9BDr473e2_1(.dout(w_dff_A_vyPi09V38_1),.din(w_dff_A_9BDr473e2_1),.clk(gclk));
	jdff dff_A_5ynAQ5FP8_1(.dout(w_dff_A_9BDr473e2_1),.din(w_dff_A_5ynAQ5FP8_1),.clk(gclk));
	jdff dff_A_3QWOje9G8_1(.dout(w_dff_A_5ynAQ5FP8_1),.din(w_dff_A_3QWOje9G8_1),.clk(gclk));
	jdff dff_A_Dw1jRvsm7_1(.dout(w_dff_A_3QWOje9G8_1),.din(w_dff_A_Dw1jRvsm7_1),.clk(gclk));
	jdff dff_A_rYyvzy0h3_1(.dout(w_dff_A_Dw1jRvsm7_1),.din(w_dff_A_rYyvzy0h3_1),.clk(gclk));
	jdff dff_A_CK34gOZr6_1(.dout(w_dff_A_rYyvzy0h3_1),.din(w_dff_A_CK34gOZr6_1),.clk(gclk));
	jdff dff_A_JoU1LoiZ6_1(.dout(w_dff_A_CK34gOZr6_1),.din(w_dff_A_JoU1LoiZ6_1),.clk(gclk));
	jdff dff_A_348Mxk9U0_1(.dout(w_dff_A_JoU1LoiZ6_1),.din(w_dff_A_348Mxk9U0_1),.clk(gclk));
	jdff dff_A_WvnTDaGw9_1(.dout(w_dff_A_348Mxk9U0_1),.din(w_dff_A_WvnTDaGw9_1),.clk(gclk));
	jdff dff_A_Y29Mh8P43_1(.dout(w_dff_A_WvnTDaGw9_1),.din(w_dff_A_Y29Mh8P43_1),.clk(gclk));
	jdff dff_A_34Hh8ZaC5_1(.dout(w_dff_A_Y29Mh8P43_1),.din(w_dff_A_34Hh8ZaC5_1),.clk(gclk));
	jdff dff_A_6j09Spgg0_1(.dout(w_dff_A_34Hh8ZaC5_1),.din(w_dff_A_6j09Spgg0_1),.clk(gclk));
	jdff dff_A_ksMFUMwP3_1(.dout(w_dff_A_6j09Spgg0_1),.din(w_dff_A_ksMFUMwP3_1),.clk(gclk));
	jdff dff_A_MagO818t6_1(.dout(w_dff_A_ksMFUMwP3_1),.din(w_dff_A_MagO818t6_1),.clk(gclk));
	jdff dff_A_VdYA3Qjv1_1(.dout(w_dff_A_MagO818t6_1),.din(w_dff_A_VdYA3Qjv1_1),.clk(gclk));
	jdff dff_A_mRX1fxRK9_1(.dout(w_dff_A_VdYA3Qjv1_1),.din(w_dff_A_mRX1fxRK9_1),.clk(gclk));
	jdff dff_A_Zm5e9g7P5_1(.dout(w_dff_A_mRX1fxRK9_1),.din(w_dff_A_Zm5e9g7P5_1),.clk(gclk));
	jdff dff_A_O5r1H6216_1(.dout(w_dff_A_Zm5e9g7P5_1),.din(w_dff_A_O5r1H6216_1),.clk(gclk));
	jdff dff_A_1gOiWsKn6_1(.dout(w_dff_A_O5r1H6216_1),.din(w_dff_A_1gOiWsKn6_1),.clk(gclk));
	jdff dff_A_3dzdKn6K9_1(.dout(w_dff_A_1gOiWsKn6_1),.din(w_dff_A_3dzdKn6K9_1),.clk(gclk));
	jdff dff_A_agWKvC6d4_1(.dout(w_dff_A_3dzdKn6K9_1),.din(w_dff_A_agWKvC6d4_1),.clk(gclk));
	jdff dff_A_6kZ25O5i0_1(.dout(w_dff_A_agWKvC6d4_1),.din(w_dff_A_6kZ25O5i0_1),.clk(gclk));
	jdff dff_A_pKK2AQ8o9_1(.dout(w_dff_A_6kZ25O5i0_1),.din(w_dff_A_pKK2AQ8o9_1),.clk(gclk));
	jdff dff_A_WWo1OGan9_1(.dout(w_dff_A_pKK2AQ8o9_1),.din(w_dff_A_WWo1OGan9_1),.clk(gclk));
	jdff dff_B_9IOKiBPx3_0(.din(n1113),.dout(w_dff_B_9IOKiBPx3_0),.clk(gclk));
	jdff dff_B_AmBrGIhR0_0(.din(w_dff_B_9IOKiBPx3_0),.dout(w_dff_B_AmBrGIhR0_0),.clk(gclk));
	jdff dff_B_M6ZwTmD70_0(.din(w_dff_B_AmBrGIhR0_0),.dout(w_dff_B_M6ZwTmD70_0),.clk(gclk));
	jdff dff_B_8kcLwFOF0_0(.din(w_dff_B_M6ZwTmD70_0),.dout(w_dff_B_8kcLwFOF0_0),.clk(gclk));
	jdff dff_B_FXcr77hx2_0(.din(w_dff_B_8kcLwFOF0_0),.dout(w_dff_B_FXcr77hx2_0),.clk(gclk));
	jdff dff_B_yGoT3d7y9_0(.din(w_dff_B_FXcr77hx2_0),.dout(w_dff_B_yGoT3d7y9_0),.clk(gclk));
	jdff dff_B_yX29Iaal8_0(.din(w_dff_B_yGoT3d7y9_0),.dout(w_dff_B_yX29Iaal8_0),.clk(gclk));
	jdff dff_B_2PGtm2bd1_0(.din(n1109),.dout(w_dff_B_2PGtm2bd1_0),.clk(gclk));
	jdff dff_B_b2c5cbPb0_0(.din(w_dff_B_2PGtm2bd1_0),.dout(w_dff_B_b2c5cbPb0_0),.clk(gclk));
	jdff dff_B_etvtQCR71_0(.din(w_dff_B_b2c5cbPb0_0),.dout(w_dff_B_etvtQCR71_0),.clk(gclk));
	jdff dff_B_xIkmAwaF3_0(.din(w_dff_B_etvtQCR71_0),.dout(w_dff_B_xIkmAwaF3_0),.clk(gclk));
	jdff dff_B_14GPHnhZ5_0(.din(w_dff_B_xIkmAwaF3_0),.dout(w_dff_B_14GPHnhZ5_0),.clk(gclk));
	jdff dff_B_1bzYNzPb2_0(.din(w_dff_B_14GPHnhZ5_0),.dout(w_dff_B_1bzYNzPb2_0),.clk(gclk));
	jdff dff_B_LpNv12ZK0_0(.din(w_dff_B_1bzYNzPb2_0),.dout(w_dff_B_LpNv12ZK0_0),.clk(gclk));
	jdff dff_B_2YJIO6bP1_1(.din(n1070),.dout(w_dff_B_2YJIO6bP1_1),.clk(gclk));
	jdff dff_B_TVj34eH45_1(.din(w_dff_B_2YJIO6bP1_1),.dout(w_dff_B_TVj34eH45_1),.clk(gclk));
	jdff dff_B_a2suvZFA7_1(.din(w_dff_B_TVj34eH45_1),.dout(w_dff_B_a2suvZFA7_1),.clk(gclk));
	jdff dff_B_vCoqdJZO5_1(.din(w_dff_B_a2suvZFA7_1),.dout(w_dff_B_vCoqdJZO5_1),.clk(gclk));
	jdff dff_B_qwclzErK5_1(.din(w_dff_B_vCoqdJZO5_1),.dout(w_dff_B_qwclzErK5_1),.clk(gclk));
	jdff dff_B_fmH78Oyd7_1(.din(w_dff_B_qwclzErK5_1),.dout(w_dff_B_fmH78Oyd7_1),.clk(gclk));
	jdff dff_B_WQ2yBKPr1_1(.din(w_dff_B_fmH78Oyd7_1),.dout(w_dff_B_WQ2yBKPr1_1),.clk(gclk));
	jdff dff_B_jY1lzMXy0_1(.din(w_dff_B_WQ2yBKPr1_1),.dout(w_dff_B_jY1lzMXy0_1),.clk(gclk));
	jdff dff_B_AgLcT7f60_1(.din(n1086),.dout(w_dff_B_AgLcT7f60_1),.clk(gclk));
	jdff dff_B_UcePQ7nO9_1(.din(w_dff_B_AgLcT7f60_1),.dout(w_dff_B_UcePQ7nO9_1),.clk(gclk));
	jdff dff_B_6p2TD6t02_1(.din(n1094),.dout(w_dff_B_6p2TD6t02_1),.clk(gclk));
	jdff dff_B_vIG23IUk8_0(.din(n1099),.dout(w_dff_B_vIG23IUk8_0),.clk(gclk));
	jdff dff_B_PAQIdhXW3_1(.din(n1075),.dout(w_dff_B_PAQIdhXW3_1),.clk(gclk));
	jdff dff_B_seMa3UNg8_1(.din(w_dff_B_PAQIdhXW3_1),.dout(w_dff_B_seMa3UNg8_1),.clk(gclk));
	jdff dff_B_SRmOgYXh7_0(.din(n1084),.dout(w_dff_B_SRmOgYXh7_0),.clk(gclk));
	jdff dff_B_q2JofDlD2_1(.din(n1076),.dout(w_dff_B_q2JofDlD2_1),.clk(gclk));
	jdff dff_B_TdsIXP264_0(.din(n1078),.dout(w_dff_B_TdsIXP264_0),.clk(gclk));
	jdff dff_B_7SvklPTh7_1(.din(G124),.dout(w_dff_B_7SvklPTh7_1),.clk(gclk));
	jdff dff_B_eqVYmkLb8_1(.din(w_dff_B_7SvklPTh7_1),.dout(w_dff_B_eqVYmkLb8_1),.clk(gclk));
	jdff dff_B_sDZ488Y14_1(.din(w_dff_B_eqVYmkLb8_1),.dout(w_dff_B_sDZ488Y14_1),.clk(gclk));
	jdff dff_B_C7SLVvkC7_1(.din(w_dff_B_sDZ488Y14_1),.dout(w_dff_B_C7SLVvkC7_1),.clk(gclk));
	jdff dff_B_dfAUOGxt2_1(.din(n1071),.dout(w_dff_B_dfAUOGxt2_1),.clk(gclk));
	jdff dff_B_Vn3lvBwj6_0(.din(n1069),.dout(w_dff_B_Vn3lvBwj6_0),.clk(gclk));
	jdff dff_B_f72n7whF8_0(.din(w_dff_B_Vn3lvBwj6_0),.dout(w_dff_B_f72n7whF8_0),.clk(gclk));
	jdff dff_B_dIaU5zlH8_0(.din(w_dff_B_f72n7whF8_0),.dout(w_dff_B_dIaU5zlH8_0),.clk(gclk));
	jdff dff_B_jIOqZmB33_1(.din(n1060),.dout(w_dff_B_jIOqZmB33_1),.clk(gclk));
	jdff dff_A_AQjdfNJy3_1(.dout(w_n1062_0[1]),.din(w_dff_A_AQjdfNJy3_1),.clk(gclk));
	jdff dff_A_RYql7SpD6_1(.dout(w_dff_A_AQjdfNJy3_1),.din(w_dff_A_RYql7SpD6_1),.clk(gclk));
	jdff dff_A_M7cIU7oP7_1(.dout(w_dff_A_RYql7SpD6_1),.din(w_dff_A_M7cIU7oP7_1),.clk(gclk));
	jdff dff_A_g66tHovf5_1(.dout(w_dff_A_M7cIU7oP7_1),.din(w_dff_A_g66tHovf5_1),.clk(gclk));
	jdff dff_A_OD4kqRMI8_1(.dout(w_dff_A_g66tHovf5_1),.din(w_dff_A_OD4kqRMI8_1),.clk(gclk));
	jdff dff_A_gBPuj7GC2_1(.dout(w_dff_A_OD4kqRMI8_1),.din(w_dff_A_gBPuj7GC2_1),.clk(gclk));
	jdff dff_A_4E3ZfTzQ6_1(.dout(w_dff_A_gBPuj7GC2_1),.din(w_dff_A_4E3ZfTzQ6_1),.clk(gclk));
	jdff dff_A_NvbC047F9_1(.dout(w_dff_A_4E3ZfTzQ6_1),.din(w_dff_A_NvbC047F9_1),.clk(gclk));
	jdff dff_B_t3YZ9YNv1_0(.din(n1061),.dout(w_dff_B_t3YZ9YNv1_0),.clk(gclk));
	jdff dff_B_QnLRwrnw8_0(.din(w_dff_B_t3YZ9YNv1_0),.dout(w_dff_B_QnLRwrnw8_0),.clk(gclk));
	jdff dff_B_nCJnhmBj5_1(.din(n764),.dout(w_dff_B_nCJnhmBj5_1),.clk(gclk));
	jdff dff_B_6uSLkFyL4_1(.din(w_dff_B_nCJnhmBj5_1),.dout(w_dff_B_6uSLkFyL4_1),.clk(gclk));
	jdff dff_B_vXSWPy6C5_1(.din(w_dff_B_6uSLkFyL4_1),.dout(w_dff_B_vXSWPy6C5_1),.clk(gclk));
	jdff dff_B_SfkCUuyu4_1(.din(w_dff_B_vXSWPy6C5_1),.dout(w_dff_B_SfkCUuyu4_1),.clk(gclk));
	jdff dff_B_E6LEHatv5_1(.din(w_dff_B_SfkCUuyu4_1),.dout(w_dff_B_E6LEHatv5_1),.clk(gclk));
	jdff dff_B_9mUJs9TO4_1(.din(w_dff_B_E6LEHatv5_1),.dout(w_dff_B_9mUJs9TO4_1),.clk(gclk));
	jdff dff_B_uCU5BhTa0_1(.din(w_dff_B_9mUJs9TO4_1),.dout(w_dff_B_uCU5BhTa0_1),.clk(gclk));
	jdff dff_B_4HRWX6FB9_1(.din(w_dff_B_uCU5BhTa0_1),.dout(w_dff_B_4HRWX6FB9_1),.clk(gclk));
	jdff dff_A_Iys6T4A83_1(.dout(w_n767_1[1]),.din(w_dff_A_Iys6T4A83_1),.clk(gclk));
	jdff dff_A_i2Gbulu39_1(.dout(w_dff_A_Iys6T4A83_1),.din(w_dff_A_i2Gbulu39_1),.clk(gclk));
	jdff dff_A_JEo4JplL4_1(.dout(w_dff_A_i2Gbulu39_1),.din(w_dff_A_JEo4JplL4_1),.clk(gclk));
	jdff dff_B_MzbukCNK4_0(.din(n763),.dout(w_dff_B_MzbukCNK4_0),.clk(gclk));
	jdff dff_B_s8dXbXUQ9_0(.din(w_dff_B_MzbukCNK4_0),.dout(w_dff_B_s8dXbXUQ9_0),.clk(gclk));
	jdff dff_B_qQRl7ORa8_0(.din(w_dff_B_s8dXbXUQ9_0),.dout(w_dff_B_qQRl7ORa8_0),.clk(gclk));
	jdff dff_B_6xmW4B3f8_0(.din(w_dff_B_qQRl7ORa8_0),.dout(w_dff_B_6xmW4B3f8_0),.clk(gclk));
	jdff dff_B_mDHgUgxZ7_0(.din(w_dff_B_6xmW4B3f8_0),.dout(w_dff_B_mDHgUgxZ7_0),.clk(gclk));
	jdff dff_B_uxtRcIsy7_0(.din(w_dff_B_mDHgUgxZ7_0),.dout(w_dff_B_uxtRcIsy7_0),.clk(gclk));
	jdff dff_B_XZ06BLZb3_0(.din(n1058),.dout(w_dff_B_XZ06BLZb3_0),.clk(gclk));
	jdff dff_B_soZKWZSH9_1(.din(n1027),.dout(w_dff_B_soZKWZSH9_1),.clk(gclk));
	jdff dff_B_DVJbvddl0_1(.din(w_dff_B_soZKWZSH9_1),.dout(w_dff_B_DVJbvddl0_1),.clk(gclk));
	jdff dff_B_t14mZ7Wt6_1(.din(w_dff_B_DVJbvddl0_1),.dout(w_dff_B_t14mZ7Wt6_1),.clk(gclk));
	jdff dff_B_TKIzkszB4_1(.din(w_dff_B_t14mZ7Wt6_1),.dout(w_dff_B_TKIzkszB4_1),.clk(gclk));
	jdff dff_B_YmC8U9uy1_1(.din(w_dff_B_TKIzkszB4_1),.dout(w_dff_B_YmC8U9uy1_1),.clk(gclk));
	jdff dff_B_NEDV5Qq39_1(.din(w_dff_B_YmC8U9uy1_1),.dout(w_dff_B_NEDV5Qq39_1),.clk(gclk));
	jdff dff_B_O181L9ZS5_1(.din(w_dff_B_NEDV5Qq39_1),.dout(w_dff_B_O181L9ZS5_1),.clk(gclk));
	jdff dff_B_4uF57oCj4_1(.din(w_dff_B_O181L9ZS5_1),.dout(w_dff_B_4uF57oCj4_1),.clk(gclk));
	jdff dff_B_1N7T31AP7_0(.din(n1051),.dout(w_dff_B_1N7T31AP7_0),.clk(gclk));
	jdff dff_A_L99Ypaxn3_1(.dout(w_n1045_0[1]),.din(w_dff_A_L99Ypaxn3_1),.clk(gclk));
	jdff dff_A_qSzqW1xY9_1(.dout(w_dff_A_L99Ypaxn3_1),.din(w_dff_A_qSzqW1xY9_1),.clk(gclk));
	jdff dff_B_Go0Z7t8Q7_1(.din(n769),.dout(w_dff_B_Go0Z7t8Q7_1),.clk(gclk));
	jdff dff_B_ED5gFEA37_1(.din(w_dff_B_Go0Z7t8Q7_1),.dout(w_dff_B_ED5gFEA37_1),.clk(gclk));
	jdff dff_A_vvtvW8iE0_1(.dout(w_n773_0[1]),.din(w_dff_A_vvtvW8iE0_1),.clk(gclk));
	jdff dff_A_XTyFZhMw1_1(.dout(w_n767_0[1]),.din(w_dff_A_XTyFZhMw1_1),.clk(gclk));
	jdff dff_A_PocpNMT54_1(.dout(w_dff_A_XTyFZhMw1_1),.din(w_dff_A_PocpNMT54_1),.clk(gclk));
	jdff dff_A_Mo2Sva0V8_1(.dout(w_dff_A_PocpNMT54_1),.din(w_dff_A_Mo2Sva0V8_1),.clk(gclk));
	jdff dff_A_Ney4EExm3_1(.dout(w_dff_A_Mo2Sva0V8_1),.din(w_dff_A_Ney4EExm3_1),.clk(gclk));
	jdff dff_A_ggCuepbO8_2(.dout(w_n767_0[2]),.din(w_dff_A_ggCuepbO8_2),.clk(gclk));
	jdff dff_A_mAfW15vs4_2(.dout(w_dff_A_ggCuepbO8_2),.din(w_dff_A_mAfW15vs4_2),.clk(gclk));
	jdff dff_A_z0M12BCP9_2(.dout(w_dff_A_mAfW15vs4_2),.din(w_dff_A_z0M12BCP9_2),.clk(gclk));
	jdff dff_B_nasyWk486_3(.din(n767),.dout(w_dff_B_nasyWk486_3),.clk(gclk));
	jdff dff_B_p5X6eS3F5_3(.din(w_dff_B_nasyWk486_3),.dout(w_dff_B_p5X6eS3F5_3),.clk(gclk));
	jdff dff_A_pXjCxg399_1(.dout(w_n1043_0[1]),.din(w_dff_A_pXjCxg399_1),.clk(gclk));
	jdff dff_B_B2gUorcj5_0(.din(n1025),.dout(w_dff_B_B2gUorcj5_0),.clk(gclk));
	jdff dff_B_6UKKzey64_0(.din(n1023),.dout(w_dff_B_6UKKzey64_0),.clk(gclk));
	jdff dff_B_8GJiAsB33_0(.din(w_dff_B_6UKKzey64_0),.dout(w_dff_B_8GJiAsB33_0),.clk(gclk));
	jdff dff_B_ELkhX7KN4_0(.din(w_dff_B_8GJiAsB33_0),.dout(w_dff_B_ELkhX7KN4_0),.clk(gclk));
	jdff dff_B_t3fUfV9F2_0(.din(w_dff_B_ELkhX7KN4_0),.dout(w_dff_B_t3fUfV9F2_0),.clk(gclk));
	jdff dff_B_QKTeOl1e3_0(.din(w_dff_B_t3fUfV9F2_0),.dout(w_dff_B_QKTeOl1e3_0),.clk(gclk));
	jdff dff_B_m88xIWPw1_1(.din(n1006),.dout(w_dff_B_m88xIWPw1_1),.clk(gclk));
	jdff dff_B_8gPGC0Fu6_1(.din(n1010),.dout(w_dff_B_8gPGC0Fu6_1),.clk(gclk));
	jdff dff_B_AaXitViX9_0(.din(n1015),.dout(w_dff_B_AaXitViX9_0),.clk(gclk));
	jdff dff_B_Jp6T2fN52_1(.din(n1011),.dout(w_dff_B_Jp6T2fN52_1),.clk(gclk));
	jdff dff_B_CLm81odN6_1(.din(n1007),.dout(w_dff_B_CLm81odN6_1),.clk(gclk));
	jdff dff_B_CkUcccqP4_1(.din(n998),.dout(w_dff_B_CkUcccqP4_1),.clk(gclk));
	jdff dff_B_eEs0hkWs3_1(.din(n999),.dout(w_dff_B_eEs0hkWs3_1),.clk(gclk));
	jdff dff_B_4qBjV5F97_1(.din(w_dff_B_eEs0hkWs3_1),.dout(w_dff_B_4qBjV5F97_1),.clk(gclk));
	jdff dff_B_8UkSvFVL7_1(.din(w_dff_B_4qBjV5F97_1),.dout(w_dff_B_8UkSvFVL7_1),.clk(gclk));
	jdff dff_B_0ccWCGf52_1(.din(n1000),.dout(w_dff_B_0ccWCGf52_1),.clk(gclk));
	jdff dff_B_mpEZYCdW1_1(.din(w_dff_B_0ccWCGf52_1),.dout(w_dff_B_mpEZYCdW1_1),.clk(gclk));
	jdff dff_B_qpyT6lIT2_0(.din(n1002),.dout(w_dff_B_qpyT6lIT2_0),.clk(gclk));
	jdff dff_B_MemRcEoA6_1(.din(n991),.dout(w_dff_B_MemRcEoA6_1),.clk(gclk));
	jdff dff_A_6fwpVXDc5_1(.dout(w_G125_0[1]),.din(w_dff_A_6fwpVXDc5_1),.clk(gclk));
	jdff dff_B_kYAY9cCE3_2(.din(G125),.dout(w_dff_B_kYAY9cCE3_2),.clk(gclk));
	jdff dff_B_DvAMv9hV5_2(.din(w_dff_B_kYAY9cCE3_2),.dout(w_dff_B_DvAMv9hV5_2),.clk(gclk));
	jdff dff_B_osGoo7l30_2(.din(w_dff_B_DvAMv9hV5_2),.dout(w_dff_B_osGoo7l30_2),.clk(gclk));
	jdff dff_A_ctnulHmK7_0(.dout(w_n614_2[0]),.din(w_dff_A_ctnulHmK7_0),.clk(gclk));
	jdff dff_A_wsO9wAL21_0(.dout(w_dff_A_ctnulHmK7_0),.din(w_dff_A_wsO9wAL21_0),.clk(gclk));
	jdff dff_A_peMkkoOB8_0(.dout(w_dff_A_wsO9wAL21_0),.din(w_dff_A_peMkkoOB8_0),.clk(gclk));
	jdff dff_A_lBHOKvxP8_1(.dout(w_n614_2[1]),.din(w_dff_A_lBHOKvxP8_1),.clk(gclk));
	jdff dff_A_lN4oWSO32_1(.dout(w_dff_A_lBHOKvxP8_1),.din(w_dff_A_lN4oWSO32_1),.clk(gclk));
	jdff dff_A_zJXLAHkh2_1(.dout(w_dff_A_lN4oWSO32_1),.din(w_dff_A_zJXLAHkh2_1),.clk(gclk));
	jdff dff_A_6XkRdgC42_1(.dout(w_dff_A_zJXLAHkh2_1),.din(w_dff_A_6XkRdgC42_1),.clk(gclk));
	jdff dff_A_UPHyR0D85_1(.dout(w_dff_A_6XkRdgC42_1),.din(w_dff_A_UPHyR0D85_1),.clk(gclk));
	jdff dff_A_IId9JDG40_1(.dout(w_dff_A_UPHyR0D85_1),.din(w_dff_A_IId9JDG40_1),.clk(gclk));
	jdff dff_A_8vlSL97B9_1(.dout(w_dff_A_IId9JDG40_1),.din(w_dff_A_8vlSL97B9_1),.clk(gclk));
	jdff dff_A_TkQ626Ep1_1(.dout(w_dff_A_8vlSL97B9_1),.din(w_dff_A_TkQ626Ep1_1),.clk(gclk));
	jdff dff_A_Eq3uJins8_1(.dout(w_dff_A_TkQ626Ep1_1),.din(w_dff_A_Eq3uJins8_1),.clk(gclk));
	jdff dff_A_e0sy6Ty21_1(.dout(w_dff_A_Eq3uJins8_1),.din(w_dff_A_e0sy6Ty21_1),.clk(gclk));
	jdff dff_A_gps9NreM1_1(.dout(w_dff_A_e0sy6Ty21_1),.din(w_dff_A_gps9NreM1_1),.clk(gclk));
	jdff dff_B_kwjGrP3X0_0(.din(n765),.dout(w_dff_B_kwjGrP3X0_0),.clk(gclk));
	jdff dff_B_pgpnDPot6_0(.din(w_dff_B_kwjGrP3X0_0),.dout(w_dff_B_pgpnDPot6_0),.clk(gclk));
	jdff dff_B_bbDuC9hg5_1(.din(n1154),.dout(w_dff_B_bbDuC9hg5_1),.clk(gclk));
	jdff dff_B_tofmwiV27_1(.din(w_dff_B_bbDuC9hg5_1),.dout(w_dff_B_tofmwiV27_1),.clk(gclk));
	jdff dff_B_O2CbvBPK1_1(.din(w_dff_B_tofmwiV27_1),.dout(w_dff_B_O2CbvBPK1_1),.clk(gclk));
	jdff dff_B_Q26YwzAT5_1(.din(w_dff_B_O2CbvBPK1_1),.dout(w_dff_B_Q26YwzAT5_1),.clk(gclk));
	jdff dff_B_zb8rwFO40_1(.din(w_dff_B_Q26YwzAT5_1),.dout(w_dff_B_zb8rwFO40_1),.clk(gclk));
	jdff dff_B_aPConhyT7_1(.din(w_dff_B_zb8rwFO40_1),.dout(w_dff_B_aPConhyT7_1),.clk(gclk));
	jdff dff_B_DuplOqxG0_0(.din(n1157),.dout(w_dff_B_DuplOqxG0_0),.clk(gclk));
	jdff dff_B_wko8F1q72_1(.din(n1156),.dout(w_dff_B_wko8F1q72_1),.clk(gclk));
	jdff dff_B_zOWbBvLs7_0(.din(n1028),.dout(w_dff_B_zOWbBvLs7_0),.clk(gclk));
	jdff dff_A_obDpq9Wc4_0(.dout(w_n514_1[0]),.din(w_dff_A_obDpq9Wc4_0),.clk(gclk));
	jdff dff_A_KtaDcr6o2_1(.dout(w_n514_0[1]),.din(w_dff_A_KtaDcr6o2_1),.clk(gclk));
	jdff dff_A_YS7cNnUb6_1(.dout(w_dff_A_KtaDcr6o2_1),.din(w_dff_A_YS7cNnUb6_1),.clk(gclk));
	jdff dff_A_76GUKfTK9_2(.dout(w_n514_0[2]),.din(w_dff_A_76GUKfTK9_2),.clk(gclk));
	jdff dff_A_6ypzyubQ1_2(.dout(w_dff_A_76GUKfTK9_2),.din(w_dff_A_6ypzyubQ1_2),.clk(gclk));
	jdff dff_A_Vep6fdi22_0(.dout(w_n562_0[0]),.din(w_dff_A_Vep6fdi22_0),.clk(gclk));
	jdff dff_B_codiG89P1_1(.din(n555),.dout(w_dff_B_codiG89P1_1),.clk(gclk));
	jdff dff_B_a6D3DV1K1_1(.din(w_dff_B_codiG89P1_1),.dout(w_dff_B_a6D3DV1K1_1),.clk(gclk));
	jdff dff_B_Xsm9xh5N4_1(.din(n556),.dout(w_dff_B_Xsm9xh5N4_1),.clk(gclk));
	jdff dff_B_3wtckWVD5_1(.din(w_dff_B_Xsm9xh5N4_1),.dout(w_dff_B_3wtckWVD5_1),.clk(gclk));
	jdff dff_B_K3A7R6M86_1(.din(w_dff_B_3wtckWVD5_1),.dout(w_dff_B_K3A7R6M86_1),.clk(gclk));
	jdff dff_B_GHDibozC2_1(.din(n557),.dout(w_dff_B_GHDibozC2_1),.clk(gclk));
	jdff dff_A_vSDsysS30_0(.dout(w_n512_0[0]),.din(w_dff_A_vSDsysS30_0),.clk(gclk));
	jdff dff_B_gWM7VLxp7_1(.din(n440),.dout(w_dff_B_gWM7VLxp7_1),.clk(gclk));
	jdff dff_A_W5Ogq3VP7_1(.dout(w_n503_0[1]),.din(w_dff_A_W5Ogq3VP7_1),.clk(gclk));
	jdff dff_A_I33LFH801_1(.dout(w_n499_0[1]),.din(w_dff_A_I33LFH801_1),.clk(gclk));
	jdff dff_A_JrOA0bvg9_1(.dout(w_n74_1[1]),.din(w_dff_A_JrOA0bvg9_1),.clk(gclk));
	jdff dff_A_jLEg05hM1_1(.dout(w_dff_A_JrOA0bvg9_1),.din(w_dff_A_jLEg05hM1_1),.clk(gclk));
	jdff dff_A_0KyCEXJH5_1(.dout(w_dff_A_jLEg05hM1_1),.din(w_dff_A_0KyCEXJH5_1),.clk(gclk));
	jdff dff_A_JEG8Zf214_1(.dout(w_dff_A_0KyCEXJH5_1),.din(w_dff_A_JEG8Zf214_1),.clk(gclk));
	jdff dff_A_196A7o9u3_2(.dout(w_n74_1[2]),.din(w_dff_A_196A7o9u3_2),.clk(gclk));
	jdff dff_A_XwUXAtVT4_2(.dout(w_dff_A_196A7o9u3_2),.din(w_dff_A_XwUXAtVT4_2),.clk(gclk));
	jdff dff_A_jI0YuI4j5_2(.dout(w_dff_A_XwUXAtVT4_2),.din(w_dff_A_jI0YuI4j5_2),.clk(gclk));
	jdff dff_A_uPxZXOvn9_0(.dout(w_n494_0[0]),.din(w_dff_A_uPxZXOvn9_0),.clk(gclk));
	jdff dff_B_eapyrZRK4_1(.din(n487),.dout(w_dff_B_eapyrZRK4_1),.clk(gclk));
	jdff dff_B_s7xqtnNw8_1(.din(n489),.dout(w_dff_B_s7xqtnNw8_1),.clk(gclk));
	jdff dff_B_fPSynR9i2_1(.din(w_dff_B_s7xqtnNw8_1),.dout(w_dff_B_fPSynR9i2_1),.clk(gclk));
	jdff dff_B_mDqj1ljP3_1(.din(n485),.dout(w_dff_B_mDqj1ljP3_1),.clk(gclk));
	jdff dff_B_IOgjobww9_1(.din(w_dff_B_mDqj1ljP3_1),.dout(w_dff_B_IOgjobww9_1),.clk(gclk));
	jdff dff_B_GY5YBRnb7_1(.din(n475),.dout(w_dff_B_GY5YBRnb7_1),.clk(gclk));
	jdff dff_B_uAVr2jzw7_1(.din(w_dff_B_GY5YBRnb7_1),.dout(w_dff_B_uAVr2jzw7_1),.clk(gclk));
	jdff dff_B_G3EgqqmC4_1(.din(n476),.dout(w_dff_B_G3EgqqmC4_1),.clk(gclk));
	jdff dff_A_n48ZFbuf3_1(.dout(w_n456_0[1]),.din(w_dff_A_n48ZFbuf3_1),.clk(gclk));
	jdff dff_A_NLrLty692_0(.dout(w_n450_0[0]),.din(w_dff_A_NLrLty692_0),.clk(gclk));
	jdff dff_B_OKK6X1Xx9_1(.din(n443),.dout(w_dff_B_OKK6X1Xx9_1),.clk(gclk));
	jdff dff_A_ETyHwJZZ6_0(.dout(w_n73_2[0]),.din(w_dff_A_ETyHwJZZ6_0),.clk(gclk));
	jdff dff_A_5GUiSh0H6_0(.dout(w_dff_A_ETyHwJZZ6_0),.din(w_dff_A_5GUiSh0H6_0),.clk(gclk));
	jdff dff_A_0l8nIW9H9_0(.dout(w_dff_A_5GUiSh0H6_0),.din(w_dff_A_0l8nIW9H9_0),.clk(gclk));
	jdff dff_A_o7WcTBV71_2(.dout(w_n73_2[2]),.din(w_dff_A_o7WcTBV71_2),.clk(gclk));
	jdff dff_A_kLHkaF9J4_2(.dout(w_n151_3[2]),.din(w_dff_A_kLHkaF9J4_2),.clk(gclk));
	jdff dff_A_PzhApn8n0_2(.dout(w_dff_A_kLHkaF9J4_2),.din(w_dff_A_PzhApn8n0_2),.clk(gclk));
	jdff dff_B_HPDhHTvl3_1(.din(n429),.dout(w_dff_B_HPDhHTvl3_1),.clk(gclk));
	jdff dff_A_Zh3LZqwt0_1(.dout(w_n435_0[1]),.din(w_dff_A_Zh3LZqwt0_1),.clk(gclk));
	jdff dff_A_Cqut5Hol2_0(.dout(w_n430_0[0]),.din(w_dff_A_Cqut5Hol2_0),.clk(gclk));
	jdff dff_B_QuYqfTew0_2(.din(G223),.dout(w_dff_B_QuYqfTew0_2),.clk(gclk));
	jdff dff_B_zdMtXarI8_2(.din(w_dff_B_QuYqfTew0_2),.dout(w_dff_B_zdMtXarI8_2),.clk(gclk));
	jdff dff_A_nzPHUKnK0_0(.dout(w_n428_0[0]),.din(w_dff_A_nzPHUKnK0_0),.clk(gclk));
	jdff dff_A_UbfmXpYv9_0(.dout(w_dff_A_nzPHUKnK0_0),.din(w_dff_A_UbfmXpYv9_0),.clk(gclk));
	jdff dff_A_MpttRNvE6_0(.dout(w_n1056_0[0]),.din(w_dff_A_MpttRNvE6_0),.clk(gclk));
	jdff dff_A_VvKWeSn83_0(.dout(w_dff_A_MpttRNvE6_0),.din(w_dff_A_VvKWeSn83_0),.clk(gclk));
	jdff dff_B_IF4NufHq0_2(.din(n1056),.dout(w_dff_B_IF4NufHq0_2),.clk(gclk));
	jdff dff_A_UUzuMJy37_1(.dout(w_n351_0[1]),.din(w_dff_A_UUzuMJy37_1),.clk(gclk));
	jdff dff_A_FtBHihML4_0(.dout(w_n772_0[0]),.din(w_dff_A_FtBHihML4_0),.clk(gclk));
	jdff dff_A_D96Dk9uZ6_0(.dout(w_dff_A_FtBHihML4_0),.din(w_dff_A_D96Dk9uZ6_0),.clk(gclk));
	jdff dff_A_Z55c4btw4_0(.dout(w_dff_A_D96Dk9uZ6_0),.din(w_dff_A_Z55c4btw4_0),.clk(gclk));
	jdff dff_A_aZSTRNcR3_0(.dout(w_n771_1[0]),.din(w_dff_A_aZSTRNcR3_0),.clk(gclk));
	jdff dff_A_Fv85uBtG6_0(.dout(w_dff_A_aZSTRNcR3_0),.din(w_dff_A_Fv85uBtG6_0),.clk(gclk));
	jdff dff_A_M6D2HWEZ2_0(.dout(w_dff_A_Fv85uBtG6_0),.din(w_dff_A_M6D2HWEZ2_0),.clk(gclk));
	jdff dff_A_EPTeD56R1_0(.dout(w_dff_A_M6D2HWEZ2_0),.din(w_dff_A_EPTeD56R1_0),.clk(gclk));
	jdff dff_B_wMi9uOsJ9_0(.din(n1032),.dout(w_dff_B_wMi9uOsJ9_0),.clk(gclk));
	jdff dff_B_4ZkfhsuZ8_0(.din(w_dff_B_wMi9uOsJ9_0),.dout(w_dff_B_4ZkfhsuZ8_0),.clk(gclk));
	jdff dff_B_Uz0lf2br0_0(.din(w_dff_B_4ZkfhsuZ8_0),.dout(w_dff_B_Uz0lf2br0_0),.clk(gclk));
	jdff dff_B_CrutxyLd1_0(.din(n1151),.dout(w_dff_B_CrutxyLd1_0),.clk(gclk));
	jdff dff_B_kSpOWxbn2_0(.din(w_dff_B_CrutxyLd1_0),.dout(w_dff_B_kSpOWxbn2_0),.clk(gclk));
	jdff dff_B_pgnI3aQB0_0(.din(w_dff_B_kSpOWxbn2_0),.dout(w_dff_B_pgnI3aQB0_0),.clk(gclk));
	jdff dff_B_PQ6gA8B69_0(.din(n1150),.dout(w_dff_B_PQ6gA8B69_0),.clk(gclk));
	jdff dff_B_EGXmiC7J3_0(.din(w_dff_B_PQ6gA8B69_0),.dout(w_dff_B_EGXmiC7J3_0),.clk(gclk));
	jdff dff_B_kfpXk8sW5_0(.din(w_dff_B_EGXmiC7J3_0),.dout(w_dff_B_kfpXk8sW5_0),.clk(gclk));
	jdff dff_B_hFunX7DE5_0(.din(w_dff_B_kfpXk8sW5_0),.dout(w_dff_B_hFunX7DE5_0),.clk(gclk));
	jdff dff_B_Alqur92y5_0(.din(w_dff_B_hFunX7DE5_0),.dout(w_dff_B_Alqur92y5_0),.clk(gclk));
	jdff dff_B_mz2u4UQD9_1(.din(n1131),.dout(w_dff_B_mz2u4UQD9_1),.clk(gclk));
	jdff dff_B_UeGz7vFO4_1(.din(w_dff_B_mz2u4UQD9_1),.dout(w_dff_B_UeGz7vFO4_1),.clk(gclk));
	jdff dff_B_VI8urFpX0_1(.din(n1132),.dout(w_dff_B_VI8urFpX0_1),.clk(gclk));
	jdff dff_B_qI34WO6Q9_1(.din(w_dff_B_VI8urFpX0_1),.dout(w_dff_B_qI34WO6Q9_1),.clk(gclk));
	jdff dff_B_WtBCHLNl5_1(.din(w_dff_B_qI34WO6Q9_1),.dout(w_dff_B_WtBCHLNl5_1),.clk(gclk));
	jdff dff_B_I96gKeLI7_1(.din(w_dff_B_WtBCHLNl5_1),.dout(w_dff_B_I96gKeLI7_1),.clk(gclk));
	jdff dff_B_OckltRcT2_1(.din(w_dff_B_I96gKeLI7_1),.dout(w_dff_B_OckltRcT2_1),.clk(gclk));
	jdff dff_B_cBcHvVMM1_1(.din(n1135),.dout(w_dff_B_cBcHvVMM1_1),.clk(gclk));
	jdff dff_B_c4620I9v0_1(.din(w_dff_B_cBcHvVMM1_1),.dout(w_dff_B_c4620I9v0_1),.clk(gclk));
	jdff dff_B_PXEpW0aS6_1(.din(w_dff_B_c4620I9v0_1),.dout(w_dff_B_PXEpW0aS6_1),.clk(gclk));
	jdff dff_B_KZ9JUhvf0_1(.din(n1140),.dout(w_dff_B_KZ9JUhvf0_1),.clk(gclk));
	jdff dff_A_YWRtBQ7V5_0(.dout(w_G128_0[0]),.din(w_dff_A_YWRtBQ7V5_0),.clk(gclk));
	jdff dff_B_W3iuT2RV1_3(.din(G128),.dout(w_dff_B_W3iuT2RV1_3),.clk(gclk));
	jdff dff_B_8O9yucme6_3(.din(w_dff_B_W3iuT2RV1_3),.dout(w_dff_B_8O9yucme6_3),.clk(gclk));
	jdff dff_B_aXjaDQ4M0_3(.din(w_dff_B_8O9yucme6_3),.dout(w_dff_B_aXjaDQ4M0_3),.clk(gclk));
	jdff dff_A_5O647Yik4_0(.dout(w_G33_4[0]),.din(w_dff_A_5O647Yik4_0),.clk(gclk));
	jdff dff_A_2F2Oudh08_1(.dout(w_G33_4[1]),.din(w_dff_A_2F2Oudh08_1),.clk(gclk));
	jdff dff_A_XtQxDIXw9_1(.dout(w_dff_A_2F2Oudh08_1),.din(w_dff_A_XtQxDIXw9_1),.clk(gclk));
	jdff dff_A_LOuZt1hJ2_1(.dout(w_dff_A_XtQxDIXw9_1),.din(w_dff_A_LOuZt1hJ2_1),.clk(gclk));
	jdff dff_A_90HwEfKC6_1(.dout(w_dff_A_LOuZt1hJ2_1),.din(w_dff_A_90HwEfKC6_1),.clk(gclk));
	jdff dff_B_FptpMnwi7_1(.din(n1136),.dout(w_dff_B_FptpMnwi7_1),.clk(gclk));
	jdff dff_B_JeNg2Ljz2_1(.din(w_dff_B_FptpMnwi7_1),.dout(w_dff_B_JeNg2Ljz2_1),.clk(gclk));
	jdff dff_A_0yyXrzMH2_0(.dout(w_n1091_0[0]),.din(w_dff_A_0yyXrzMH2_0),.clk(gclk));
	jdff dff_A_JIa7x4XB8_1(.dout(w_G150_1[1]),.din(w_dff_A_JIa7x4XB8_1),.clk(gclk));
	jdff dff_A_oAPZEv3J5_2(.dout(w_G159_1[2]),.din(w_dff_A_oAPZEv3J5_2),.clk(gclk));
	jdff dff_B_YPROuvuL0_1(.din(n1118),.dout(w_dff_B_YPROuvuL0_1),.clk(gclk));
	jdff dff_B_JxhsXLS99_1(.din(w_dff_B_YPROuvuL0_1),.dout(w_dff_B_JxhsXLS99_1),.clk(gclk));
	jdff dff_A_bvHEwYPn0_1(.dout(w_G283_1[1]),.din(w_dff_A_bvHEwYPn0_1),.clk(gclk));
	jdff dff_A_NcO9Sjbo1_2(.dout(w_n771_0[2]),.din(w_dff_A_NcO9Sjbo1_2),.clk(gclk));
	jdff dff_A_6eiINvJZ3_2(.dout(w_dff_A_NcO9Sjbo1_2),.din(w_dff_A_6eiINvJZ3_2),.clk(gclk));
	jdff dff_A_mdZgBqlb2_2(.dout(w_dff_A_6eiINvJZ3_2),.din(w_dff_A_mdZgBqlb2_2),.clk(gclk));
	jdff dff_A_TJwIehfe4_2(.dout(w_dff_A_mdZgBqlb2_2),.din(w_dff_A_TJwIehfe4_2),.clk(gclk));
	jdff dff_B_5c9wZdRa0_0(.din(n770),.dout(w_dff_B_5c9wZdRa0_0),.clk(gclk));
	jdff dff_B_IWopkhLh1_0(.din(w_dff_B_5c9wZdRa0_0),.dout(w_dff_B_IWopkhLh1_0),.clk(gclk));
	jdff dff_B_ZNbHQtQH4_0(.din(w_dff_B_IWopkhLh1_0),.dout(w_dff_B_ZNbHQtQH4_0),.clk(gclk));
	jdff dff_B_hQIfFVma4_0(.din(w_dff_B_ZNbHQtQH4_0),.dout(w_dff_B_hQIfFVma4_0),.clk(gclk));
	jdff dff_A_FcdkyXoc5_1(.dout(w_n420_0[1]),.din(w_dff_A_FcdkyXoc5_1),.clk(gclk));
	jdff dff_A_Oh91G41R4_1(.dout(w_n417_0[1]),.din(w_dff_A_Oh91G41R4_1),.clk(gclk));
	jdff dff_A_SKxkA4gY1_2(.dout(w_n417_0[2]),.din(w_dff_A_SKxkA4gY1_2),.clk(gclk));
	jdff dff_B_9sgztSk90_1(.din(n411),.dout(w_dff_B_9sgztSk90_1),.clk(gclk));
	jdff dff_B_bH0fzxpY2_1(.din(w_dff_B_9sgztSk90_1),.dout(w_dff_B_bH0fzxpY2_1),.clk(gclk));
	jdff dff_B_mqMdDvCO3_1(.din(n413),.dout(w_dff_B_mqMdDvCO3_1),.clk(gclk));
	jdff dff_B_BhPBEMs71_1(.din(w_dff_B_mqMdDvCO3_1),.dout(w_dff_B_BhPBEMs71_1),.clk(gclk));
	jdff dff_A_MchgcMM65_0(.dout(w_G68_4[0]),.din(w_dff_A_MchgcMM65_0),.clk(gclk));
	jdff dff_A_vb2mpHcf6_0(.dout(w_dff_A_MchgcMM65_0),.din(w_dff_A_vb2mpHcf6_0),.clk(gclk));
	jdff dff_A_SfnC8UI12_2(.dout(w_G68_4[2]),.din(w_dff_A_SfnC8UI12_2),.clk(gclk));
	jdff dff_A_0msoXEw23_2(.dout(w_dff_A_SfnC8UI12_2),.din(w_dff_A_0msoXEw23_2),.clk(gclk));
	jdff dff_A_IMx4AmGF3_2(.dout(w_dff_A_0msoXEw23_2),.din(w_dff_A_IMx4AmGF3_2),.clk(gclk));
	jdff dff_A_gwvRXqe98_2(.dout(w_dff_A_IMx4AmGF3_2),.din(w_dff_A_gwvRXqe98_2),.clk(gclk));
	jdff dff_A_OE7sgIuQ1_2(.dout(w_dff_A_gwvRXqe98_2),.din(w_dff_A_OE7sgIuQ1_2),.clk(gclk));
	jdff dff_B_lrgl6soP5_0(.din(n412),.dout(w_dff_B_lrgl6soP5_0),.clk(gclk));
	jdff dff_A_xc49V2yN9_1(.dout(w_n407_0[1]),.din(w_dff_A_xc49V2yN9_1),.clk(gclk));
	jdff dff_B_Vz7Z6xjQ8_1(.din(n397),.dout(w_dff_B_Vz7Z6xjQ8_1),.clk(gclk));
	jdff dff_B_947c0t5M6_1(.din(w_dff_B_Vz7Z6xjQ8_1),.dout(w_dff_B_947c0t5M6_1),.clk(gclk));
	jdff dff_B_EwVOvqLO1_1(.din(n398),.dout(w_dff_B_EwVOvqLO1_1),.clk(gclk));
	jdff dff_A_ZrygzSyX5_0(.dout(w_n168_2[0]),.din(w_dff_A_ZrygzSyX5_0),.clk(gclk));
	jdff dff_A_9QBz8RYs5_0(.dout(w_dff_A_ZrygzSyX5_0),.din(w_dff_A_9QBz8RYs5_0),.clk(gclk));
	jdff dff_A_e5E483ow0_0(.dout(w_G384_0),.din(w_dff_A_e5E483ow0_0),.clk(gclk));
	jdff dff_A_Q2U1rWYC3_0(.dout(w_dff_A_e5E483ow0_0),.din(w_dff_A_Q2U1rWYC3_0),.clk(gclk));
	jdff dff_A_UDsUAlsV2_0(.dout(w_dff_A_Q2U1rWYC3_0),.din(w_dff_A_UDsUAlsV2_0),.clk(gclk));
	jdff dff_A_g5xzbAJs4_0(.dout(w_n759_0[0]),.din(w_dff_A_g5xzbAJs4_0),.clk(gclk));
	jdff dff_A_vgLnRoeq5_0(.dout(w_dff_A_g5xzbAJs4_0),.din(w_dff_A_vgLnRoeq5_0),.clk(gclk));
	jdff dff_A_UydSEI1R7_0(.dout(w_dff_A_vgLnRoeq5_0),.din(w_dff_A_UydSEI1R7_0),.clk(gclk));
	jdff dff_A_akZQpuOp2_0(.dout(w_dff_A_UydSEI1R7_0),.din(w_dff_A_akZQpuOp2_0),.clk(gclk));
	jdff dff_B_rh4QLE558_1(.din(n747),.dout(w_dff_B_rh4QLE558_1),.clk(gclk));
	jdff dff_B_WE9fOSRN4_1(.din(w_dff_B_rh4QLE558_1),.dout(w_dff_B_WE9fOSRN4_1),.clk(gclk));
	jdff dff_B_UcjOiyLY9_0(.din(n751),.dout(w_dff_B_UcjOiyLY9_0),.clk(gclk));
	jdff dff_B_7B0RoYiB7_1(.din(n296),.dout(w_dff_B_7B0RoYiB7_1),.clk(gclk));
	jdff dff_A_EmMFb6Ux0_0(.dout(w_n395_0[0]),.din(w_dff_A_EmMFb6Ux0_0),.clk(gclk));
	jdff dff_A_zDloW7fa1_0(.dout(w_dff_A_EmMFb6Ux0_0),.din(w_dff_A_zDloW7fa1_0),.clk(gclk));
	jdff dff_A_YTi8Dgu26_0(.dout(w_dff_A_zDloW7fa1_0),.din(w_dff_A_YTi8Dgu26_0),.clk(gclk));
	jdff dff_B_hVfg89iI1_0(.din(n745),.dout(w_dff_B_hVfg89iI1_0),.clk(gclk));
	jdff dff_B_yiifLGK53_0(.din(w_dff_B_hVfg89iI1_0),.dout(w_dff_B_yiifLGK53_0),.clk(gclk));
	jdff dff_B_vhBtoQwU7_0(.din(w_dff_B_yiifLGK53_0),.dout(w_dff_B_vhBtoQwU7_0),.clk(gclk));
	jdff dff_B_iNYb9PqW3_0(.din(w_dff_B_vhBtoQwU7_0),.dout(w_dff_B_iNYb9PqW3_0),.clk(gclk));
	jdff dff_B_6axqDvYD6_0(.din(n743),.dout(w_dff_B_6axqDvYD6_0),.clk(gclk));
	jdff dff_B_a4VQMPiO2_0(.din(w_dff_B_6axqDvYD6_0),.dout(w_dff_B_a4VQMPiO2_0),.clk(gclk));
	jdff dff_B_yOlpVy2k4_0(.din(w_dff_B_a4VQMPiO2_0),.dout(w_dff_B_yOlpVy2k4_0),.clk(gclk));
	jdff dff_B_vaDBoLY89_0(.din(w_dff_B_yOlpVy2k4_0),.dout(w_dff_B_vaDBoLY89_0),.clk(gclk));
	jdff dff_B_QeiMDT8I5_1(.din(n740),.dout(w_dff_B_QeiMDT8I5_1),.clk(gclk));
	jdff dff_A_czxibepF3_0(.dout(w_n618_1[0]),.din(w_dff_A_czxibepF3_0),.clk(gclk));
	jdff dff_A_YimUmIaL6_0(.dout(w_dff_A_czxibepF3_0),.din(w_dff_A_YimUmIaL6_0),.clk(gclk));
	jdff dff_A_40nzIkoe9_0(.dout(w_dff_A_YimUmIaL6_0),.din(w_dff_A_40nzIkoe9_0),.clk(gclk));
	jdff dff_A_yXd4Uuu18_0(.dout(w_dff_A_40nzIkoe9_0),.din(w_dff_A_yXd4Uuu18_0),.clk(gclk));
	jdff dff_A_YXZheSm79_0(.dout(w_dff_A_yXd4Uuu18_0),.din(w_dff_A_YXZheSm79_0),.clk(gclk));
	jdff dff_A_D0lwcCld0_0(.dout(w_dff_A_YXZheSm79_0),.din(w_dff_A_D0lwcCld0_0),.clk(gclk));
	jdff dff_A_QGPlReu91_0(.dout(w_dff_A_D0lwcCld0_0),.din(w_dff_A_QGPlReu91_0),.clk(gclk));
	jdff dff_A_82kfVSlJ5_0(.dout(w_dff_A_QGPlReu91_0),.din(w_dff_A_82kfVSlJ5_0),.clk(gclk));
	jdff dff_A_vqqHyQld4_0(.dout(w_dff_A_82kfVSlJ5_0),.din(w_dff_A_vqqHyQld4_0),.clk(gclk));
	jdff dff_A_SCvhVDYY6_0(.dout(w_dff_A_vqqHyQld4_0),.din(w_dff_A_SCvhVDYY6_0),.clk(gclk));
	jdff dff_A_vp9rvH7c9_0(.dout(w_dff_A_SCvhVDYY6_0),.din(w_dff_A_vp9rvH7c9_0),.clk(gclk));
	jdff dff_A_xgxKAMrc7_1(.dout(w_n618_1[1]),.din(w_dff_A_xgxKAMrc7_1),.clk(gclk));
	jdff dff_A_W6tDfEn78_1(.dout(w_dff_A_xgxKAMrc7_1),.din(w_dff_A_W6tDfEn78_1),.clk(gclk));
	jdff dff_A_sWjbEFMw4_1(.dout(w_dff_A_W6tDfEn78_1),.din(w_dff_A_sWjbEFMw4_1),.clk(gclk));
	jdff dff_A_3WDz4osr6_1(.dout(w_dff_A_sWjbEFMw4_1),.din(w_dff_A_3WDz4osr6_1),.clk(gclk));
	jdff dff_A_xlixRGKu3_1(.dout(w_dff_A_3WDz4osr6_1),.din(w_dff_A_xlixRGKu3_1),.clk(gclk));
	jdff dff_A_VM8dThXw0_1(.dout(w_dff_A_xlixRGKu3_1),.din(w_dff_A_VM8dThXw0_1),.clk(gclk));
	jdff dff_A_pOrw0prw5_1(.dout(w_dff_A_VM8dThXw0_1),.din(w_dff_A_pOrw0prw5_1),.clk(gclk));
	jdff dff_A_eWucBi366_1(.dout(w_dff_A_pOrw0prw5_1),.din(w_dff_A_eWucBi366_1),.clk(gclk));
	jdff dff_A_u5hNhmDB3_1(.dout(w_dff_A_eWucBi366_1),.din(w_dff_A_u5hNhmDB3_1),.clk(gclk));
	jdff dff_A_Dz7BMP8p7_1(.dout(w_dff_A_u5hNhmDB3_1),.din(w_dff_A_Dz7BMP8p7_1),.clk(gclk));
	jdff dff_A_om1uan588_1(.dout(w_dff_A_Dz7BMP8p7_1),.din(w_dff_A_om1uan588_1),.clk(gclk));
	jdff dff_B_OhgEfmRx3_0(.din(n735),.dout(w_dff_B_OhgEfmRx3_0),.clk(gclk));
	jdff dff_B_c4JQbR9H5_0(.din(n726),.dout(w_dff_B_c4JQbR9H5_0),.clk(gclk));
	jdff dff_B_Qgk1zIAq1_1(.din(n723),.dout(w_dff_B_Qgk1zIAq1_1),.clk(gclk));
	jdff dff_B_oCrH7Lgx0_1(.din(n713),.dout(w_dff_B_oCrH7Lgx0_1),.clk(gclk));
	jdff dff_B_LPi0uogA1_1(.din(n716),.dout(w_dff_B_LPi0uogA1_1),.clk(gclk));
	jdff dff_A_n5GY4sdo6_0(.dout(w_n718_0[0]),.din(w_dff_A_n5GY4sdo6_0),.clk(gclk));
	jdff dff_A_9ipMDwCo7_0(.dout(w_dff_A_n5GY4sdo6_0),.din(w_dff_A_9ipMDwCo7_0),.clk(gclk));
	jdff dff_A_1uyzNcr30_0(.dout(w_dff_A_9ipMDwCo7_0),.din(w_dff_A_1uyzNcr30_0),.clk(gclk));
	jdff dff_A_tpD3wjjN6_0(.dout(w_dff_A_1uyzNcr30_0),.din(w_dff_A_tpD3wjjN6_0),.clk(gclk));
	jdff dff_B_5UdxwxRG3_2(.din(n718),.dout(w_dff_B_5UdxwxRG3_2),.clk(gclk));
	jdff dff_B_l3j8OZvY8_1(.din(n714),.dout(w_dff_B_l3j8OZvY8_1),.clk(gclk));
	jdff dff_A_97lxGxD29_1(.dout(w_G132_1[1]),.din(w_dff_A_97lxGxD29_1),.clk(gclk));
	jdff dff_B_WfF5hDW57_3(.din(G132),.dout(w_dff_B_WfF5hDW57_3),.clk(gclk));
	jdff dff_B_wPFcyzwI9_3(.din(w_dff_B_WfF5hDW57_3),.dout(w_dff_B_wPFcyzwI9_3),.clk(gclk));
	jdff dff_B_EDPlRGQZ8_3(.din(w_dff_B_wPFcyzwI9_3),.dout(w_dff_B_EDPlRGQZ8_3),.clk(gclk));
	jdff dff_B_yO4odglo3_1(.din(n707),.dout(w_dff_B_yO4odglo3_1),.clk(gclk));
	jdff dff_B_CsOHDHJM3_1(.din(w_dff_B_yO4odglo3_1),.dout(w_dff_B_CsOHDHJM3_1),.clk(gclk));
	jdff dff_B_0YsiHeIC6_0(.din(n711),.dout(w_dff_B_0YsiHeIC6_0),.clk(gclk));
	jdff dff_A_nbkZK3gz7_0(.dout(w_G150_3[0]),.din(w_dff_A_nbkZK3gz7_0),.clk(gclk));
	jdff dff_A_226JHW4E9_0(.dout(w_n704_0[0]),.din(w_dff_A_226JHW4E9_0),.clk(gclk));
	jdff dff_A_JH3Amltv7_0(.dout(w_dff_A_226JHW4E9_0),.din(w_dff_A_JH3Amltv7_0),.clk(gclk));
	jdff dff_A_TXIsUPNy8_0(.dout(w_n703_1[0]),.din(w_dff_A_TXIsUPNy8_0),.clk(gclk));
	jdff dff_A_39XrxDvY6_0(.dout(w_dff_A_TXIsUPNy8_0),.din(w_dff_A_39XrxDvY6_0),.clk(gclk));
	jdff dff_A_iOdcPdRN2_0(.dout(w_dff_A_39XrxDvY6_0),.din(w_dff_A_iOdcPdRN2_0),.clk(gclk));
	jdff dff_A_mjcIPlYI2_1(.dout(w_n703_0[1]),.din(w_dff_A_mjcIPlYI2_1),.clk(gclk));
	jdff dff_A_W95K5KKG3_1(.dout(w_dff_A_mjcIPlYI2_1),.din(w_dff_A_W95K5KKG3_1),.clk(gclk));
	jdff dff_A_ByPGuawY7_1(.dout(w_dff_A_W95K5KKG3_1),.din(w_dff_A_ByPGuawY7_1),.clk(gclk));
	jdff dff_A_qHvtVqkT7_2(.dout(w_n703_0[2]),.din(w_dff_A_qHvtVqkT7_2),.clk(gclk));
	jdff dff_B_vI1890VH2_0(.din(n702),.dout(w_dff_B_vI1890VH2_0),.clk(gclk));
	jdff dff_B_gmxxOQzu0_0(.din(w_dff_B_vI1890VH2_0),.dout(w_dff_B_gmxxOQzu0_0),.clk(gclk));
	jdff dff_B_tIvO4YzW4_0(.din(w_dff_B_gmxxOQzu0_0),.dout(w_dff_B_tIvO4YzW4_0),.clk(gclk));
	jdff dff_B_oEGQHARh0_0(.din(w_dff_B_tIvO4YzW4_0),.dout(w_dff_B_oEGQHARh0_0),.clk(gclk));
	jdff dff_B_LzxIiMpc8_0(.din(w_dff_B_oEGQHARh0_0),.dout(w_dff_B_LzxIiMpc8_0),.clk(gclk));
	jdff dff_A_sdMQGsvz6_0(.dout(w_n567_3[0]),.din(w_dff_A_sdMQGsvz6_0),.clk(gclk));
	jdff dff_A_ruwX4sgZ3_1(.dout(w_n567_3[1]),.din(w_dff_A_ruwX4sgZ3_1),.clk(gclk));
	jdff dff_A_wWlgZZ4S2_1(.dout(w_dff_A_ruwX4sgZ3_1),.din(w_dff_A_wWlgZZ4S2_1),.clk(gclk));
	jdff dff_A_RLsYC9xP9_1(.dout(w_dff_A_wWlgZZ4S2_1),.din(w_dff_A_RLsYC9xP9_1),.clk(gclk));
	jdff dff_A_t9pnQjqb7_1(.dout(w_dff_A_RLsYC9xP9_1),.din(w_dff_A_t9pnQjqb7_1),.clk(gclk));
	jdff dff_A_1cZgT8FT3_1(.dout(w_dff_A_t9pnQjqb7_1),.din(w_dff_A_1cZgT8FT3_1),.clk(gclk));
	jdff dff_A_aYTPkeyl4_1(.dout(w_dff_A_1cZgT8FT3_1),.din(w_dff_A_aYTPkeyl4_1),.clk(gclk));
	jdff dff_A_dTjGelrD5_1(.dout(w_dff_A_aYTPkeyl4_1),.din(w_dff_A_dTjGelrD5_1),.clk(gclk));
	jdff dff_A_LR5W7OFQ5_1(.dout(w_n388_2[1]),.din(w_dff_A_LR5W7OFQ5_1),.clk(gclk));
	jdff dff_B_qhibm7nF7_1(.din(n384),.dout(w_dff_B_qhibm7nF7_1),.clk(gclk));
	jdff dff_B_IAH45NQo8_1(.din(w_dff_B_qhibm7nF7_1),.dout(w_dff_B_IAH45NQo8_1),.clk(gclk));
	jdff dff_A_UZ27vMAF8_1(.dout(w_n383_0[1]),.din(w_dff_A_UZ27vMAF8_1),.clk(gclk));
	jdff dff_A_GdC3iBAj1_1(.dout(w_dff_A_UZ27vMAF8_1),.din(w_dff_A_GdC3iBAj1_1),.clk(gclk));
	jdff dff_A_PSySrwr68_1(.dout(w_dff_A_GdC3iBAj1_1),.din(w_dff_A_PSySrwr68_1),.clk(gclk));
	jdff dff_B_2DwCmg7O1_1(.din(n374),.dout(w_dff_B_2DwCmg7O1_1),.clk(gclk));
	jdff dff_B_2c83vRPV0_0(.din(n381),.dout(w_dff_B_2c83vRPV0_0),.clk(gclk));
	jdff dff_B_aEtb0mcV1_1(.din(n376),.dout(w_dff_B_aEtb0mcV1_1),.clk(gclk));
	jdff dff_A_pgfK9uma1_0(.dout(w_n378_0[0]),.din(w_dff_A_pgfK9uma1_0),.clk(gclk));
	jdff dff_A_34WEawZK6_0(.dout(w_n370_0[0]),.din(w_dff_A_34WEawZK6_0),.clk(gclk));
	jdff dff_B_gHQTSLrz0_2(.din(n370),.dout(w_dff_B_gHQTSLrz0_2),.clk(gclk));
	jdff dff_B_jLV0ghFw1_0(.din(n365),.dout(w_dff_B_jLV0ghFw1_0),.clk(gclk));
	jdff dff_B_pGicBI5G6_1(.din(n358),.dout(w_dff_B_pGicBI5G6_1),.clk(gclk));
	jdff dff_A_jxVQlUsh1_1(.dout(w_n357_0[1]),.din(w_dff_A_jxVQlUsh1_1),.clk(gclk));
	jdff dff_A_u0zShoW77_1(.dout(w_dff_A_jxVQlUsh1_1),.din(w_dff_A_u0zShoW77_1),.clk(gclk));
	jdff dff_A_Mi458JfJ5_0(.dout(w_n356_1[0]),.din(w_dff_A_Mi458JfJ5_0),.clk(gclk));
	jdff dff_A_LB2BJLy78_1(.dout(w_n356_0[1]),.din(w_dff_A_LB2BJLy78_1),.clk(gclk));
	jdff dff_A_CwoR9y7N7_2(.dout(w_n356_0[2]),.din(w_dff_A_CwoR9y7N7_2),.clk(gclk));
	jdff dff_A_uEuoVxFA7_0(.dout(w_n354_1[0]),.din(w_dff_A_uEuoVxFA7_0),.clk(gclk));
	jdff dff_A_NDct26XZ8_1(.dout(w_n354_0[1]),.din(w_dff_A_NDct26XZ8_1),.clk(gclk));
	jdff dff_A_zzA9gOhC2_2(.dout(w_n354_0[2]),.din(w_dff_A_zzA9gOhC2_2),.clk(gclk));
	jdff dff_A_7H2DEj1c7_1(.dout(w_n1177_0[1]),.din(w_dff_A_7H2DEj1c7_1),.clk(gclk));
	jdff dff_A_Lz3Y5PGp7_1(.dout(w_dff_A_7H2DEj1c7_1),.din(w_dff_A_Lz3Y5PGp7_1),.clk(gclk));
	jdff dff_B_hpwzkZhz7_2(.din(n1177),.dout(w_dff_B_hpwzkZhz7_2),.clk(gclk));
	jdff dff_B_Dq2Xk9Zs5_2(.din(w_dff_B_hpwzkZhz7_2),.dout(w_dff_B_Dq2Xk9Zs5_2),.clk(gclk));
	jdff dff_B_cRQ7BKJr4_1(.din(n1175),.dout(w_dff_B_cRQ7BKJr4_1),.clk(gclk));
	jdff dff_B_76G1R80I7_1(.din(n942),.dout(w_dff_B_76G1R80I7_1),.clk(gclk));
	jdff dff_B_MW8Bjtcc4_0(.din(n985),.dout(w_dff_B_MW8Bjtcc4_0),.clk(gclk));
	jdff dff_B_EEa8Na864_0(.din(w_dff_B_MW8Bjtcc4_0),.dout(w_dff_B_EEa8Na864_0),.clk(gclk));
	jdff dff_B_lnQ8HUb74_0(.din(w_dff_B_EEa8Na864_0),.dout(w_dff_B_lnQ8HUb74_0),.clk(gclk));
	jdff dff_B_L79gYsFG0_0(.din(w_dff_B_lnQ8HUb74_0),.dout(w_dff_B_L79gYsFG0_0),.clk(gclk));
	jdff dff_B_JC0CyPB34_0(.din(w_dff_B_L79gYsFG0_0),.dout(w_dff_B_JC0CyPB34_0),.clk(gclk));
	jdff dff_B_gNQYeVZj1_0(.din(n983),.dout(w_dff_B_gNQYeVZj1_0),.clk(gclk));
	jdff dff_B_Og2VNfOO6_0(.din(w_dff_B_gNQYeVZj1_0),.dout(w_dff_B_Og2VNfOO6_0),.clk(gclk));
	jdff dff_B_Q6ihH8472_1(.din(n949),.dout(w_dff_B_Q6ihH8472_1),.clk(gclk));
	jdff dff_B_p0uyDgDK6_1(.din(w_dff_B_Q6ihH8472_1),.dout(w_dff_B_p0uyDgDK6_1),.clk(gclk));
	jdff dff_B_LpW2euEs6_1(.din(w_dff_B_p0uyDgDK6_1),.dout(w_dff_B_LpW2euEs6_1),.clk(gclk));
	jdff dff_B_7g4tZBYO7_1(.din(w_dff_B_LpW2euEs6_1),.dout(w_dff_B_7g4tZBYO7_1),.clk(gclk));
	jdff dff_B_7whsfyG25_1(.din(n967),.dout(w_dff_B_7whsfyG25_1),.clk(gclk));
	jdff dff_B_Y3pctb3y9_1(.din(n974),.dout(w_dff_B_Y3pctb3y9_1),.clk(gclk));
	jdff dff_A_cUW9NY2e1_2(.dout(w_G116_2[2]),.din(w_dff_A_cUW9NY2e1_2),.clk(gclk));
	jdff dff_B_QGb6dHNc8_1(.din(n965),.dout(w_dff_B_QGb6dHNc8_1),.clk(gclk));
	jdff dff_A_p726uaCi3_1(.dout(w_G294_1[1]),.din(w_dff_A_p726uaCi3_1),.clk(gclk));
	jdff dff_B_oesYkrT41_1(.din(n952),.dout(w_dff_B_oesYkrT41_1),.clk(gclk));
	jdff dff_B_1o1k8E266_1(.din(w_dff_B_oesYkrT41_1),.dout(w_dff_B_1o1k8E266_1),.clk(gclk));
	jdff dff_B_2fzj4tTD7_1(.din(w_dff_B_1o1k8E266_1),.dout(w_dff_B_2fzj4tTD7_1),.clk(gclk));
	jdff dff_B_00tOmlcV1_1(.din(n955),.dout(w_dff_B_00tOmlcV1_1),.clk(gclk));
	jdff dff_B_yRAbqoPj3_1(.din(w_dff_B_00tOmlcV1_1),.dout(w_dff_B_yRAbqoPj3_1),.clk(gclk));
	jdff dff_B_3538W6Se4_1(.din(n957),.dout(w_dff_B_3538W6Se4_1),.clk(gclk));
	jdff dff_A_n1qPfFTw9_0(.dout(w_n959_0[0]),.din(w_dff_A_n1qPfFTw9_0),.clk(gclk));
	jdff dff_A_ceXLqub56_0(.dout(w_dff_A_n1qPfFTw9_0),.din(w_dff_A_ceXLqub56_0),.clk(gclk));
	jdff dff_A_AvSlXyCe7_0(.dout(w_dff_A_ceXLqub56_0),.din(w_dff_A_AvSlXyCe7_0),.clk(gclk));
	jdff dff_A_0FXdgbTT2_2(.dout(w_G143_1[2]),.din(w_dff_A_0FXdgbTT2_2),.clk(gclk));
	jdff dff_A_Fweb03Sm6_1(.dout(w_G50_2[1]),.din(w_dff_A_Fweb03Sm6_1),.clk(gclk));
	jdff dff_A_zkS5FPqg8_1(.dout(w_dff_A_Fweb03Sm6_1),.din(w_dff_A_zkS5FPqg8_1),.clk(gclk));
	jdff dff_A_N4Y2Mr3N2_1(.dout(w_dff_A_zkS5FPqg8_1),.din(w_dff_A_N4Y2Mr3N2_1),.clk(gclk));
	jdff dff_A_0JtXnC2e8_2(.dout(w_G50_2[2]),.din(w_dff_A_0JtXnC2e8_2),.clk(gclk));
	jdff dff_A_q93wIPSs7_2(.dout(w_dff_A_0JtXnC2e8_2),.din(w_dff_A_q93wIPSs7_2),.clk(gclk));
	jdff dff_A_nLJPHWsy8_2(.dout(w_dff_A_q93wIPSs7_2),.din(w_dff_A_nLJPHWsy8_2),.clk(gclk));
	jdff dff_B_lm0hFwU34_1(.din(n946),.dout(w_dff_B_lm0hFwU34_1),.clk(gclk));
	jdff dff_B_LY7bYntw8_1(.din(w_dff_B_lm0hFwU34_1),.dout(w_dff_B_LY7bYntw8_1),.clk(gclk));
	jdff dff_B_AwPZqyvy3_0(.din(n947),.dout(w_dff_B_AwPZqyvy3_0),.clk(gclk));
	jdff dff_A_NxLNoeNl9_0(.dout(w_n137_0[0]),.din(w_dff_A_NxLNoeNl9_0),.clk(gclk));
	jdff dff_B_DZJ2aS4s0_0(.din(n136),.dout(w_dff_B_DZJ2aS4s0_0),.clk(gclk));
	jdff dff_B_bmkZyDxZ1_1(.din(n939),.dout(w_dff_B_bmkZyDxZ1_1),.clk(gclk));
	jdff dff_B_JvjjaOGR2_1(.din(n843),.dout(w_dff_B_JvjjaOGR2_1),.clk(gclk));
	jdff dff_B_P5QO7Brl0_1(.din(w_dff_B_JvjjaOGR2_1),.dout(w_dff_B_P5QO7Brl0_1),.clk(gclk));
	jdff dff_B_wnA5m0lB7_1(.din(w_dff_B_P5QO7Brl0_1),.dout(w_dff_B_wnA5m0lB7_1),.clk(gclk));
	jdff dff_B_vujsMn4w8_1(.din(w_dff_B_wnA5m0lB7_1),.dout(w_dff_B_vujsMn4w8_1),.clk(gclk));
	jdff dff_B_pMhcoQm33_1(.din(w_dff_B_vujsMn4w8_1),.dout(w_dff_B_pMhcoQm33_1),.clk(gclk));
	jdff dff_B_u5krdrV44_1(.din(w_dff_B_pMhcoQm33_1),.dout(w_dff_B_u5krdrV44_1),.clk(gclk));
	jdff dff_B_vSBWEpvC8_1(.din(w_dff_B_u5krdrV44_1),.dout(w_dff_B_vSBWEpvC8_1),.clk(gclk));
	jdff dff_B_DrZ5NFFL2_1(.din(n856),.dout(w_dff_B_DrZ5NFFL2_1),.clk(gclk));
	jdff dff_B_EYZKU5ko9_1(.din(w_dff_B_DrZ5NFFL2_1),.dout(w_dff_B_EYZKU5ko9_1),.clk(gclk));
	jdff dff_B_2qZ3BbhQ9_0(.din(n866),.dout(w_dff_B_2qZ3BbhQ9_0),.clk(gclk));
	jdff dff_A_ufV6lJRQ8_0(.dout(w_n863_0[0]),.din(w_dff_A_ufV6lJRQ8_0),.clk(gclk));
	jdff dff_A_oowgKUsw6_0(.dout(w_dff_A_ufV6lJRQ8_0),.din(w_dff_A_oowgKUsw6_0),.clk(gclk));
	jdff dff_A_lbuSIHpA8_0(.dout(w_dff_A_oowgKUsw6_0),.din(w_dff_A_lbuSIHpA8_0),.clk(gclk));
	jdff dff_A_gfTtQOA63_2(.dout(w_n863_0[2]),.din(w_dff_A_gfTtQOA63_2),.clk(gclk));
	jdff dff_B_YAk8KxDc6_1(.din(n847),.dout(w_dff_B_YAk8KxDc6_1),.clk(gclk));
	jdff dff_B_FRUsGpKl3_1(.din(n848),.dout(w_dff_B_FRUsGpKl3_1),.clk(gclk));
	jdff dff_B_500HLwzz0_1(.din(w_dff_B_FRUsGpKl3_1),.dout(w_dff_B_500HLwzz0_1),.clk(gclk));
	jdff dff_B_8phYCkmE0_1(.din(w_dff_B_500HLwzz0_1),.dout(w_dff_B_8phYCkmE0_1),.clk(gclk));
	jdff dff_B_ZAfep1yA9_1(.din(w_dff_B_8phYCkmE0_1),.dout(w_dff_B_ZAfep1yA9_1),.clk(gclk));
	jdff dff_B_drb9tgyI3_0(.din(n851),.dout(w_dff_B_drb9tgyI3_0),.clk(gclk));
	jdff dff_A_6SXdzCnI2_1(.dout(w_n569_0[1]),.din(w_dff_A_6SXdzCnI2_1),.clk(gclk));
	jdff dff_A_WfzRtcFC0_1(.dout(w_dff_A_6SXdzCnI2_1),.din(w_dff_A_WfzRtcFC0_1),.clk(gclk));
	jdff dff_A_CrFou7NL0_0(.dout(w_n348_0[0]),.din(w_dff_A_CrFou7NL0_0),.clk(gclk));
	jdff dff_A_AcbZ4Tay0_0(.dout(w_n333_0[0]),.din(w_dff_A_AcbZ4Tay0_0),.clk(gclk));
	jdff dff_A_JS0Y1SzS9_0(.dout(w_dff_A_AcbZ4Tay0_0),.din(w_dff_A_JS0Y1SzS9_0),.clk(gclk));
	jdff dff_B_tascgUPq3_0(.din(n846),.dout(w_dff_B_tascgUPq3_0),.clk(gclk));
	jdff dff_B_olPxfAgE5_0(.din(w_dff_B_tascgUPq3_0),.dout(w_dff_B_olPxfAgE5_0),.clk(gclk));
	jdff dff_A_zBDMi8J16_1(.dout(w_n845_0[1]),.din(w_dff_A_zBDMi8J16_1),.clk(gclk));
	jdff dff_A_41v9qUwg2_1(.dout(w_dff_A_zBDMi8J16_1),.din(w_dff_A_41v9qUwg2_1),.clk(gclk));
	jdff dff_A_jsVmobp23_1(.dout(w_dff_A_41v9qUwg2_1),.din(w_dff_A_jsVmobp23_1),.clk(gclk));
	jdff dff_A_OG8upKwM1_1(.dout(w_dff_A_jsVmobp23_1),.din(w_dff_A_OG8upKwM1_1),.clk(gclk));
	jdff dff_B_tDkrTTgd8_0(.din(n844),.dout(w_dff_B_tDkrTTgd8_0),.clk(gclk));
	jdff dff_B_XrN8ujoq0_0(.din(w_dff_B_tDkrTTgd8_0),.dout(w_dff_B_XrN8ujoq0_0),.clk(gclk));
	jdff dff_B_JiavlIFh1_0(.din(w_dff_B_XrN8ujoq0_0),.dout(w_dff_B_JiavlIFh1_0),.clk(gclk));
	jdff dff_A_yxo8XTQb4_1(.dout(w_n579_1[1]),.din(w_dff_A_yxo8XTQb4_1),.clk(gclk));
	jdff dff_A_nBTj7VM28_1(.dout(w_dff_A_yxo8XTQb4_1),.din(w_dff_A_nBTj7VM28_1),.clk(gclk));
	jdff dff_B_reR9chzK7_0(.din(n841),.dout(w_dff_B_reR9chzK7_0),.clk(gclk));
	jdff dff_B_lryXG1jZ6_1(.din(n806),.dout(w_dff_B_lryXG1jZ6_1),.clk(gclk));
	jdff dff_B_dnmNCXeR4_1(.din(w_dff_B_lryXG1jZ6_1),.dout(w_dff_B_dnmNCXeR4_1),.clk(gclk));
	jdff dff_B_tbPUkQaw0_1(.din(w_dff_B_dnmNCXeR4_1),.dout(w_dff_B_tbPUkQaw0_1),.clk(gclk));
	jdff dff_B_3oQ96Ro83_1(.din(n825),.dout(w_dff_B_3oQ96Ro83_1),.clk(gclk));
	jdff dff_B_PwACYx4m9_1(.din(w_dff_B_3oQ96Ro83_1),.dout(w_dff_B_PwACYx4m9_1),.clk(gclk));
	jdff dff_B_wcfSg0N25_1(.din(n828),.dout(w_dff_B_wcfSg0N25_1),.clk(gclk));
	jdff dff_B_RxJFYEeT9_1(.din(w_dff_B_wcfSg0N25_1),.dout(w_dff_B_RxJFYEeT9_1),.clk(gclk));
	jdff dff_B_evK5ALlS6_0(.din(n834),.dout(w_dff_B_evK5ALlS6_0),.clk(gclk));
	jdff dff_A_1gSwhNQf5_0(.dout(w_n833_0[0]),.din(w_dff_A_1gSwhNQf5_0),.clk(gclk));
	jdff dff_B_xumulVta2_1(.din(n829),.dout(w_dff_B_xumulVta2_1),.clk(gclk));
	jdff dff_A_RooK4Q3D0_0(.dout(w_G58_3[0]),.din(w_dff_A_RooK4Q3D0_0),.clk(gclk));
	jdff dff_A_bG2djZ6W8_0(.dout(w_dff_A_RooK4Q3D0_0),.din(w_dff_A_bG2djZ6W8_0),.clk(gclk));
	jdff dff_A_QDZZMnUA1_0(.dout(w_dff_A_bG2djZ6W8_0),.din(w_dff_A_QDZZMnUA1_0),.clk(gclk));
	jdff dff_A_YJiz5Z9H3_2(.dout(w_G58_3[2]),.din(w_dff_A_YJiz5Z9H3_2),.clk(gclk));
	jdff dff_A_3ZEmc1Qq4_2(.dout(w_dff_A_YJiz5Z9H3_2),.din(w_dff_A_3ZEmc1Qq4_2),.clk(gclk));
	jdff dff_A_GR0woiLp9_2(.dout(w_dff_A_3ZEmc1Qq4_2),.din(w_dff_A_GR0woiLp9_2),.clk(gclk));
	jdff dff_A_ziTFnVBC9_2(.dout(w_dff_A_GR0woiLp9_2),.din(w_dff_A_ziTFnVBC9_2),.clk(gclk));
	jdff dff_B_OSTqnc9o9_3(.din(G143),.dout(w_dff_B_OSTqnc9o9_3),.clk(gclk));
	jdff dff_B_yZBK22iS5_3(.din(w_dff_B_OSTqnc9o9_3),.dout(w_dff_B_yZBK22iS5_3),.clk(gclk));
	jdff dff_B_2fQBAMhR4_3(.din(w_dff_B_yZBK22iS5_3),.dout(w_dff_B_2fQBAMhR4_3),.clk(gclk));
	jdff dff_B_J4G9mpnt1_1(.din(n823),.dout(w_dff_B_J4G9mpnt1_1),.clk(gclk));
	jdff dff_A_8cGpDfv52_1(.dout(w_G137_1[1]),.din(w_dff_A_8cGpDfv52_1),.clk(gclk));
	jdff dff_B_3A6t9QDM7_3(.din(G137),.dout(w_dff_B_3A6t9QDM7_3),.clk(gclk));
	jdff dff_B_Ux9afbeq9_3(.din(w_dff_B_3A6t9QDM7_3),.dout(w_dff_B_Ux9afbeq9_3),.clk(gclk));
	jdff dff_B_24faEiGY7_3(.din(w_dff_B_Ux9afbeq9_3),.dout(w_dff_B_24faEiGY7_3),.clk(gclk));
	jdff dff_B_Pa7mNo931_1(.din(n809),.dout(w_dff_B_Pa7mNo931_1),.clk(gclk));
	jdff dff_B_E0lqSfHI1_1(.din(w_dff_B_Pa7mNo931_1),.dout(w_dff_B_E0lqSfHI1_1),.clk(gclk));
	jdff dff_B_ITBo9cRh8_1(.din(w_dff_B_E0lqSfHI1_1),.dout(w_dff_B_ITBo9cRh8_1),.clk(gclk));
	jdff dff_B_tBpgZeHR6_1(.din(n812),.dout(w_dff_B_tBpgZeHR6_1),.clk(gclk));
	jdff dff_B_IcFqzFcb4_1(.din(w_dff_B_tBpgZeHR6_1),.dout(w_dff_B_IcFqzFcb4_1),.clk(gclk));
	jdff dff_A_GugwOcEI1_1(.dout(w_G107_2[1]),.din(w_dff_A_GugwOcEI1_1),.clk(gclk));
	jdff dff_B_ORF3evCs4_1(.din(n813),.dout(w_dff_B_ORF3evCs4_1),.clk(gclk));
	jdff dff_A_s7wx6l3t2_0(.dout(w_n680_3[0]),.din(w_dff_A_s7wx6l3t2_0),.clk(gclk));
	jdff dff_A_Hn3xa1Rf4_0(.dout(w_dff_A_s7wx6l3t2_0),.din(w_dff_A_Hn3xa1Rf4_0),.clk(gclk));
	jdff dff_A_HKxft28O8_0(.dout(w_dff_A_Hn3xa1Rf4_0),.din(w_dff_A_HKxft28O8_0),.clk(gclk));
	jdff dff_A_TQ8QPLsV9_0(.dout(w_dff_A_HKxft28O8_0),.din(w_dff_A_TQ8QPLsV9_0),.clk(gclk));
	jdff dff_A_oyhoAt5v5_0(.dout(w_dff_A_TQ8QPLsV9_0),.din(w_dff_A_oyhoAt5v5_0),.clk(gclk));
	jdff dff_A_XaaQSeDR1_0(.dout(w_dff_A_oyhoAt5v5_0),.din(w_dff_A_XaaQSeDR1_0),.clk(gclk));
	jdff dff_A_GbYdWwlj5_0(.dout(w_dff_A_XaaQSeDR1_0),.din(w_dff_A_GbYdWwlj5_0),.clk(gclk));
	jdff dff_A_UNfPpoSj7_2(.dout(w_n680_3[2]),.din(w_dff_A_UNfPpoSj7_2),.clk(gclk));
	jdff dff_A_xDs9WJzV1_2(.dout(w_dff_A_UNfPpoSj7_2),.din(w_dff_A_xDs9WJzV1_2),.clk(gclk));
	jdff dff_A_JMSQkLdp9_2(.dout(w_dff_A_xDs9WJzV1_2),.din(w_dff_A_JMSQkLdp9_2),.clk(gclk));
	jdff dff_A_1xwARsnp4_2(.dout(w_dff_A_JMSQkLdp9_2),.din(w_dff_A_1xwARsnp4_2),.clk(gclk));
	jdff dff_A_n8K1NTCA0_2(.dout(w_dff_A_1xwARsnp4_2),.din(w_dff_A_n8K1NTCA0_2),.clk(gclk));
	jdff dff_A_JmyOfB7B1_2(.dout(w_dff_A_n8K1NTCA0_2),.din(w_dff_A_JmyOfB7B1_2),.clk(gclk));
	jdff dff_B_3EdAInlv4_1(.din(n801),.dout(w_dff_B_3EdAInlv4_1),.clk(gclk));
	jdff dff_B_9kC6cd7E5_1(.din(w_dff_B_3EdAInlv4_1),.dout(w_dff_B_9kC6cd7E5_1),.clk(gclk));
	jdff dff_B_jHdHPdUh9_0(.din(n803),.dout(w_dff_B_jHdHPdUh9_0),.clk(gclk));
	jdff dff_A_oZ09gIbv8_0(.dout(w_n126_0[0]),.din(w_dff_A_oZ09gIbv8_0),.clk(gclk));
	jdff dff_B_PHRg72GV4_0(.din(n125),.dout(w_dff_B_PHRg72GV4_0),.clk(gclk));
	jdff dff_A_f2O2TfQE2_1(.dout(w_n614_4[1]),.din(w_dff_A_f2O2TfQE2_1),.clk(gclk));
	jdff dff_A_ROk1wMdd7_1(.dout(w_dff_A_f2O2TfQE2_1),.din(w_dff_A_ROk1wMdd7_1),.clk(gclk));
	jdff dff_A_O1iMba9j5_1(.dout(w_dff_A_ROk1wMdd7_1),.din(w_dff_A_O1iMba9j5_1),.clk(gclk));
	jdff dff_A_N5L1lzpW5_1(.dout(w_dff_A_O1iMba9j5_1),.din(w_dff_A_N5L1lzpW5_1),.clk(gclk));
	jdff dff_A_QjXIX3JX3_1(.dout(w_dff_A_N5L1lzpW5_1),.din(w_dff_A_QjXIX3JX3_1),.clk(gclk));
	jdff dff_A_q4424rMo6_1(.dout(w_dff_A_QjXIX3JX3_1),.din(w_dff_A_q4424rMo6_1),.clk(gclk));
	jdff dff_A_qQHdypN76_1(.dout(w_dff_A_q4424rMo6_1),.din(w_dff_A_qQHdypN76_1),.clk(gclk));
	jdff dff_A_p8ELpzs83_1(.dout(w_dff_A_qQHdypN76_1),.din(w_dff_A_p8ELpzs83_1),.clk(gclk));
	jdff dff_A_NPPMvooM8_1(.dout(w_dff_A_p8ELpzs83_1),.din(w_dff_A_NPPMvooM8_1),.clk(gclk));
	jdff dff_A_zsDmacJB5_1(.dout(w_dff_A_NPPMvooM8_1),.din(w_dff_A_zsDmacJB5_1),.clk(gclk));
	jdff dff_A_7SMRNitG2_1(.dout(w_dff_A_zsDmacJB5_1),.din(w_dff_A_7SMRNitG2_1),.clk(gclk));
	jdff dff_A_aBqoN1gC4_1(.dout(w_dff_A_7SMRNitG2_1),.din(w_dff_A_aBqoN1gC4_1),.clk(gclk));
	jdff dff_A_rhnNNtjf9_2(.dout(w_n614_4[2]),.din(w_dff_A_rhnNNtjf9_2),.clk(gclk));
	jdff dff_A_TuA7yQBL6_2(.dout(w_dff_A_rhnNNtjf9_2),.din(w_dff_A_TuA7yQBL6_2),.clk(gclk));
	jdff dff_A_U4G2hbYB4_2(.dout(w_dff_A_TuA7yQBL6_2),.din(w_dff_A_U4G2hbYB4_2),.clk(gclk));
	jdff dff_A_VZajrdVB7_2(.dout(w_dff_A_U4G2hbYB4_2),.din(w_dff_A_VZajrdVB7_2),.clk(gclk));
	jdff dff_A_FNF8GtI49_0(.dout(w_n798_0[0]),.din(w_dff_A_FNF8GtI49_0),.clk(gclk));
	jdff dff_A_cda3Ibtk0_0(.dout(w_dff_A_FNF8GtI49_0),.din(w_dff_A_cda3Ibtk0_0),.clk(gclk));
	jdff dff_A_ZoqZzlTJ5_0(.dout(w_dff_A_cda3Ibtk0_0),.din(w_dff_A_ZoqZzlTJ5_0),.clk(gclk));
	jdff dff_A_PY053j2E3_0(.dout(w_dff_A_ZoqZzlTJ5_0),.din(w_dff_A_PY053j2E3_0),.clk(gclk));
	jdff dff_A_NWjxawI12_0(.dout(w_dff_A_PY053j2E3_0),.din(w_dff_A_NWjxawI12_0),.clk(gclk));
	jdff dff_B_aw7lozyC2_0(.din(n797),.dout(w_dff_B_aw7lozyC2_0),.clk(gclk));
	jdff dff_B_n68jINf37_0(.din(w_dff_B_aw7lozyC2_0),.dout(w_dff_B_n68jINf37_0),.clk(gclk));
	jdff dff_A_CsKIKhNk8_2(.dout(w_n567_2[2]),.din(w_dff_A_CsKIKhNk8_2),.clk(gclk));
	jdff dff_A_6ClywbqX8_2(.dout(w_dff_A_CsKIKhNk8_2),.din(w_dff_A_6ClywbqX8_2),.clk(gclk));
	jdff dff_A_yv9RxOo11_2(.dout(w_dff_A_6ClywbqX8_2),.din(w_dff_A_yv9RxOo11_2),.clk(gclk));
	jdff dff_A_oCgTu8PU1_2(.dout(w_dff_A_yv9RxOo11_2),.din(w_dff_A_oCgTu8PU1_2),.clk(gclk));
	jdff dff_A_om3QB3IG7_2(.dout(w_dff_A_oCgTu8PU1_2),.din(w_dff_A_om3QB3IG7_2),.clk(gclk));
	jdff dff_A_kIFH2Ysa1_2(.dout(w_dff_A_om3QB3IG7_2),.din(w_dff_A_kIFH2Ysa1_2),.clk(gclk));
	jdff dff_A_b1lHgAcI0_2(.dout(w_dff_A_kIFH2Ysa1_2),.din(w_dff_A_b1lHgAcI0_2),.clk(gclk));
	jdff dff_A_OKjBty4r9_2(.dout(w_dff_A_b1lHgAcI0_2),.din(w_dff_A_OKjBty4r9_2),.clk(gclk));
	jdff dff_A_RsAMSWpq3_2(.dout(w_dff_A_OKjBty4r9_2),.din(w_dff_A_RsAMSWpq3_2),.clk(gclk));
	jdff dff_B_mBIfwTu57_0(.din(n936),.dout(w_dff_B_mBIfwTu57_0),.clk(gclk));
	jdff dff_B_HxCQNKHB7_0(.din(w_dff_B_mBIfwTu57_0),.dout(w_dff_B_HxCQNKHB7_0),.clk(gclk));
	jdff dff_B_Qes4Prln1_0(.din(w_dff_B_HxCQNKHB7_0),.dout(w_dff_B_Qes4Prln1_0),.clk(gclk));
	jdff dff_B_9gG2pNCA3_0(.din(w_dff_B_Qes4Prln1_0),.dout(w_dff_B_9gG2pNCA3_0),.clk(gclk));
	jdff dff_B_jlxAK9nM9_0(.din(w_dff_B_9gG2pNCA3_0),.dout(w_dff_B_jlxAK9nM9_0),.clk(gclk));
	jdff dff_B_9cMgXHwX2_0(.din(n932),.dout(w_dff_B_9cMgXHwX2_0),.clk(gclk));
	jdff dff_B_t2YV5ulg4_0(.din(w_dff_B_9cMgXHwX2_0),.dout(w_dff_B_t2YV5ulg4_0),.clk(gclk));
	jdff dff_B_RF4hpguR9_1(.din(n917),.dout(w_dff_B_RF4hpguR9_1),.clk(gclk));
	jdff dff_B_A3jLiNuo4_1(.din(w_dff_B_RF4hpguR9_1),.dout(w_dff_B_A3jLiNuo4_1),.clk(gclk));
	jdff dff_B_BNt8wNsu8_1(.din(w_dff_B_A3jLiNuo4_1),.dout(w_dff_B_BNt8wNsu8_1),.clk(gclk));
	jdff dff_B_tyQKaLlA7_0(.din(n929),.dout(w_dff_B_tyQKaLlA7_0),.clk(gclk));
	jdff dff_B_KdZ70WhS7_0(.din(w_dff_B_tyQKaLlA7_0),.dout(w_dff_B_KdZ70WhS7_0),.clk(gclk));
	jdff dff_B_7ESZrZng0_0(.din(n927),.dout(w_dff_B_7ESZrZng0_0),.clk(gclk));
	jdff dff_A_8psWY8rS6_1(.dout(w_n73_1[1]),.din(w_dff_A_8psWY8rS6_1),.clk(gclk));
	jdff dff_A_YyiYAuhi0_1(.dout(w_dff_A_8psWY8rS6_1),.din(w_dff_A_YyiYAuhi0_1),.clk(gclk));
	jdff dff_A_XMNBXna95_2(.dout(w_n73_1[2]),.din(w_dff_A_XMNBXna95_2),.clk(gclk));
	jdff dff_A_6uaoxXlx0_2(.dout(w_dff_A_XMNBXna95_2),.din(w_dff_A_6uaoxXlx0_2),.clk(gclk));
	jdff dff_A_DSLseczh2_2(.dout(w_dff_A_6uaoxXlx0_2),.din(w_dff_A_DSLseczh2_2),.clk(gclk));
	jdff dff_A_FadPCto76_2(.dout(w_dff_A_DSLseczh2_2),.din(w_dff_A_FadPCto76_2),.clk(gclk));
	jdff dff_A_4iOF6mXk2_2(.dout(w_n73_0[2]),.din(w_dff_A_4iOF6mXk2_2),.clk(gclk));
	jdff dff_A_Sd7ZNSfY2_2(.dout(w_dff_A_4iOF6mXk2_2),.din(w_dff_A_Sd7ZNSfY2_2),.clk(gclk));
	jdff dff_A_CVp4pTp89_2(.dout(w_dff_A_Sd7ZNSfY2_2),.din(w_dff_A_CVp4pTp89_2),.clk(gclk));
	jdff dff_A_8fctjVtq2_2(.dout(w_dff_A_CVp4pTp89_2),.din(w_dff_A_8fctjVtq2_2),.clk(gclk));
	jdff dff_B_6MfxNJ1F1_0(.din(n922),.dout(w_dff_B_6MfxNJ1F1_0),.clk(gclk));
	jdff dff_B_Q4nvGl6c1_0(.din(n921),.dout(w_dff_B_Q4nvGl6c1_0),.clk(gclk));
	jdff dff_A_K5y6vMox0_1(.dout(w_n130_0[1]),.din(w_dff_A_K5y6vMox0_1),.clk(gclk));
	jdff dff_B_3f5k93LL3_0(.din(n129),.dout(w_dff_B_3f5k93LL3_0),.clk(gclk));
	jdff dff_A_iXiu8ig33_0(.dout(w_G232_1[0]),.din(w_dff_A_iXiu8ig33_0),.clk(gclk));
	jdff dff_A_40PAzvkt0_0(.dout(w_dff_A_iXiu8ig33_0),.din(w_dff_A_40PAzvkt0_0),.clk(gclk));
	jdff dff_A_rNztm4fG1_1(.dout(w_G232_0[1]),.din(w_dff_A_rNztm4fG1_1),.clk(gclk));
	jdff dff_A_De6k9eKv4_1(.dout(w_dff_A_rNztm4fG1_1),.din(w_dff_A_De6k9eKv4_1),.clk(gclk));
	jdff dff_A_5mpRZrMx0_1(.dout(w_dff_A_De6k9eKv4_1),.din(w_dff_A_5mpRZrMx0_1),.clk(gclk));
	jdff dff_A_PfoVU7vB4_2(.dout(w_G232_0[2]),.din(w_dff_A_PfoVU7vB4_2),.clk(gclk));
	jdff dff_A_rGcJMBIj6_2(.dout(w_dff_A_PfoVU7vB4_2),.din(w_dff_A_rGcJMBIj6_2),.clk(gclk));
	jdff dff_A_WPNxCxhU7_0(.dout(w_G226_1[0]),.din(w_dff_A_WPNxCxhU7_0),.clk(gclk));
	jdff dff_A_wBv5RdHQ9_0(.dout(w_dff_A_WPNxCxhU7_0),.din(w_dff_A_wBv5RdHQ9_0),.clk(gclk));
	jdff dff_A_OHByhVgl2_1(.dout(w_G226_0[1]),.din(w_dff_A_OHByhVgl2_1),.clk(gclk));
	jdff dff_A_8DaOgCE19_1(.dout(w_dff_A_OHByhVgl2_1),.din(w_dff_A_8DaOgCE19_1),.clk(gclk));
	jdff dff_A_Sn8UzVX90_2(.dout(w_G226_0[2]),.din(w_dff_A_Sn8UzVX90_2),.clk(gclk));
	jdff dff_A_AEw2G3VR6_2(.dout(w_dff_A_Sn8UzVX90_2),.din(w_dff_A_AEw2G3VR6_2),.clk(gclk));
	jdff dff_A_cOKP08oN6_2(.dout(w_dff_A_AEw2G3VR6_2),.din(w_dff_A_cOKP08oN6_2),.clk(gclk));
	jdff dff_A_e6d3Dqpr7_1(.dout(w_n802_0[1]),.din(w_dff_A_e6d3Dqpr7_1),.clk(gclk));
	jdff dff_A_fJHbRvmw7_1(.dout(w_dff_A_e6d3Dqpr7_1),.din(w_dff_A_fJHbRvmw7_1),.clk(gclk));
	jdff dff_A_gH7AkekS8_1(.dout(w_dff_A_fJHbRvmw7_1),.din(w_dff_A_gH7AkekS8_1),.clk(gclk));
	jdff dff_A_eiDE24Oq2_1(.dout(w_dff_A_gH7AkekS8_1),.din(w_dff_A_eiDE24Oq2_1),.clk(gclk));
	jdff dff_B_LDgdsH4j0_0(.din(n913),.dout(w_dff_B_LDgdsH4j0_0),.clk(gclk));
	jdff dff_B_mJyPI1ZB7_0(.din(w_dff_B_LDgdsH4j0_0),.dout(w_dff_B_mJyPI1ZB7_0),.clk(gclk));
	jdff dff_B_K0aRBr5x9_1(.din(n898),.dout(w_dff_B_K0aRBr5x9_1),.clk(gclk));
	jdff dff_B_TGNX02BM7_1(.din(w_dff_B_K0aRBr5x9_1),.dout(w_dff_B_TGNX02BM7_1),.clk(gclk));
	jdff dff_B_XsJZ1J8F9_1(.din(w_dff_B_TGNX02BM7_1),.dout(w_dff_B_XsJZ1J8F9_1),.clk(gclk));
	jdff dff_B_gNEDBGez0_1(.din(w_dff_B_XsJZ1J8F9_1),.dout(w_dff_B_gNEDBGez0_1),.clk(gclk));
	jdff dff_B_USA1XYU61_0(.din(n909),.dout(w_dff_B_USA1XYU61_0),.clk(gclk));
	jdff dff_A_JHKb9dFG7_1(.dout(w_n153_3[1]),.din(w_dff_A_JHKb9dFG7_1),.clk(gclk));
	jdff dff_A_aPMWqlyr2_1(.dout(w_dff_A_JHKb9dFG7_1),.din(w_dff_A_aPMWqlyr2_1),.clk(gclk));
	jdff dff_A_AszVSaBX6_1(.dout(w_dff_A_aPMWqlyr2_1),.din(w_dff_A_AszVSaBX6_1),.clk(gclk));
	jdff dff_A_qFW8mvb81_1(.dout(w_dff_A_AszVSaBX6_1),.din(w_dff_A_qFW8mvb81_1),.clk(gclk));
	jdff dff_A_tsGL62uo6_1(.dout(w_dff_A_qFW8mvb81_1),.din(w_dff_A_tsGL62uo6_1),.clk(gclk));
	jdff dff_A_yoJMUpJN0_2(.dout(w_n153_3[2]),.din(w_dff_A_yoJMUpJN0_2),.clk(gclk));
	jdff dff_A_x9FcaIIF3_2(.dout(w_dff_A_yoJMUpJN0_2),.din(w_dff_A_x9FcaIIF3_2),.clk(gclk));
	jdff dff_B_ITkbkyJf1_1(.din(n902),.dout(w_dff_B_ITkbkyJf1_1),.clk(gclk));
	jdff dff_B_uJOhXaQ34_1(.din(n899),.dout(w_dff_B_uJOhXaQ34_1),.clk(gclk));
	jdff dff_A_XgHMaMKJ0_1(.dout(w_G283_2[1]),.din(w_dff_A_XgHMaMKJ0_1),.clk(gclk));
	jdff dff_B_PERCOOkK4_1(.din(n883),.dout(w_dff_B_PERCOOkK4_1),.clk(gclk));
	jdff dff_B_h4qqhYoZ3_1(.din(n888),.dout(w_dff_B_h4qqhYoZ3_1),.clk(gclk));
	jdff dff_B_O3Odp1da0_0(.din(n892),.dout(w_dff_B_O3Odp1da0_0),.clk(gclk));
	jdff dff_B_v9iNmF707_0(.din(w_dff_B_O3Odp1da0_0),.dout(w_dff_B_v9iNmF707_0),.clk(gclk));
	jdff dff_B_RwoL5VWu8_1(.din(n889),.dout(w_dff_B_RwoL5VWu8_1),.clk(gclk));
	jdff dff_A_sDiaw4jP0_1(.dout(w_G150_2[1]),.din(w_dff_A_sDiaw4jP0_1),.clk(gclk));
	jdff dff_A_xY4JYrGU6_0(.dout(w_G150_0[0]),.din(w_dff_A_xY4JYrGU6_0),.clk(gclk));
	jdff dff_A_fhwY2GGF7_1(.dout(w_G150_0[1]),.din(w_dff_A_fhwY2GGF7_1),.clk(gclk));
	jdff dff_B_lOVN20O51_3(.din(G150),.dout(w_dff_B_lOVN20O51_3),.clk(gclk));
	jdff dff_B_rVxBzmCT4_3(.din(w_dff_B_lOVN20O51_3),.dout(w_dff_B_rVxBzmCT4_3),.clk(gclk));
	jdff dff_A_CxId2X4p1_0(.dout(w_G50_3[0]),.din(w_dff_A_CxId2X4p1_0),.clk(gclk));
	jdff dff_A_YeNUUbk43_0(.dout(w_dff_A_CxId2X4p1_0),.din(w_dff_A_YeNUUbk43_0),.clk(gclk));
	jdff dff_A_Yq1g9EbF9_0(.dout(w_dff_A_YeNUUbk43_0),.din(w_dff_A_Yq1g9EbF9_0),.clk(gclk));
	jdff dff_A_QovUWjK44_1(.dout(w_G50_3[1]),.din(w_dff_A_QovUWjK44_1),.clk(gclk));
	jdff dff_A_PCgw152I9_1(.dout(w_dff_A_QovUWjK44_1),.din(w_dff_A_PCgw152I9_1),.clk(gclk));
	jdff dff_A_W5vhrWtU2_1(.dout(w_dff_A_PCgw152I9_1),.din(w_dff_A_W5vhrWtU2_1),.clk(gclk));
	jdff dff_A_xR7b1os08_1(.dout(w_n887_0[1]),.din(w_dff_A_xR7b1os08_1),.clk(gclk));
	jdff dff_A_PcNxiZVX6_0(.dout(w_G77_2[0]),.din(w_dff_A_PcNxiZVX6_0),.clk(gclk));
	jdff dff_A_IIsPcozW7_1(.dout(w_G77_2[1]),.din(w_dff_A_IIsPcozW7_1),.clk(gclk));
	jdff dff_A_O0UPS0rg6_1(.dout(w_G87_1[1]),.din(w_dff_A_O0UPS0rg6_1),.clk(gclk));
	jdff dff_A_u3LkBAgE3_2(.dout(w_G87_1[2]),.din(w_dff_A_u3LkBAgE3_2),.clk(gclk));
	jdff dff_B_UF5t5H872_1(.din(n878),.dout(w_dff_B_UF5t5H872_1),.clk(gclk));
	jdff dff_B_8Vywqy5C4_1(.din(w_dff_B_UF5t5H872_1),.dout(w_dff_B_8Vywqy5C4_1),.clk(gclk));
	jdff dff_A_C1qcDK9h2_1(.dout(w_G68_2[1]),.din(w_dff_A_C1qcDK9h2_1),.clk(gclk));
	jdff dff_A_vSeCGvWH5_1(.dout(w_dff_A_C1qcDK9h2_1),.din(w_dff_A_vSeCGvWH5_1),.clk(gclk));
	jdff dff_A_xOXKEPir9_1(.dout(w_dff_A_vSeCGvWH5_1),.din(w_dff_A_xOXKEPir9_1),.clk(gclk));
	jdff dff_A_A5yn995E5_2(.dout(w_G68_2[2]),.din(w_dff_A_A5yn995E5_2),.clk(gclk));
	jdff dff_A_5zADzc499_2(.dout(w_dff_A_A5yn995E5_2),.din(w_dff_A_5zADzc499_2),.clk(gclk));
	jdff dff_A_8LkxneID7_2(.dout(w_dff_A_5zADzc499_2),.din(w_dff_A_8LkxneID7_2),.clk(gclk));
	jdff dff_A_V27RGjLX5_2(.dout(w_dff_A_8LkxneID7_2),.din(w_dff_A_V27RGjLX5_2),.clk(gclk));
	jdff dff_A_jZ8bFWoo9_1(.dout(w_n817_0[1]),.din(w_dff_A_jZ8bFWoo9_1),.clk(gclk));
	jdff dff_A_YnKQKoVh5_1(.dout(w_G97_2[1]),.din(w_dff_A_YnKQKoVh5_1),.clk(gclk));
	jdff dff_A_MzxxoxCA9_1(.dout(w_G33_5[1]),.din(w_dff_A_MzxxoxCA9_1),.clk(gclk));
	jdff dff_A_DVdKI9wv2_1(.dout(w_dff_A_MzxxoxCA9_1),.din(w_dff_A_DVdKI9wv2_1),.clk(gclk));
	jdff dff_A_yuAZQRgU4_1(.dout(w_dff_A_DVdKI9wv2_1),.din(w_dff_A_yuAZQRgU4_1),.clk(gclk));
	jdff dff_A_ef7BMETH9_0(.dout(w_G58_2[0]),.din(w_dff_A_ef7BMETH9_0),.clk(gclk));
	jdff dff_A_tuXdhDwY1_0(.dout(w_dff_A_ef7BMETH9_0),.din(w_dff_A_tuXdhDwY1_0),.clk(gclk));
	jdff dff_A_Ipm7vSBl0_2(.dout(w_G58_2[2]),.din(w_dff_A_Ipm7vSBl0_2),.clk(gclk));
	jdff dff_A_bAIyhmRv0_2(.dout(w_dff_A_Ipm7vSBl0_2),.din(w_dff_A_bAIyhmRv0_2),.clk(gclk));
	jdff dff_A_JvW1s6wj8_0(.dout(w_n680_2[0]),.din(w_dff_A_JvW1s6wj8_0),.clk(gclk));
	jdff dff_A_U5NGfB3C5_0(.dout(w_dff_A_JvW1s6wj8_0),.din(w_dff_A_U5NGfB3C5_0),.clk(gclk));
	jdff dff_A_4jPOWda36_2(.dout(w_n680_2[2]),.din(w_dff_A_4jPOWda36_2),.clk(gclk));
	jdff dff_A_VXiDgnTl0_2(.dout(w_dff_A_4jPOWda36_2),.din(w_dff_A_VXiDgnTl0_2),.clk(gclk));
	jdff dff_A_mQ5PH6K54_2(.dout(w_dff_A_VXiDgnTl0_2),.din(w_dff_A_mQ5PH6K54_2),.clk(gclk));
	jdff dff_A_BZKHOI4D0_1(.dout(w_n614_3[1]),.din(w_dff_A_BZKHOI4D0_1),.clk(gclk));
	jdff dff_A_w0RmUAOp6_1(.dout(w_dff_A_BZKHOI4D0_1),.din(w_dff_A_w0RmUAOp6_1),.clk(gclk));
	jdff dff_A_qcIAzvu09_1(.dout(w_dff_A_w0RmUAOp6_1),.din(w_dff_A_qcIAzvu09_1),.clk(gclk));
	jdff dff_A_uhmDajlO9_1(.dout(w_dff_A_qcIAzvu09_1),.din(w_dff_A_uhmDajlO9_1),.clk(gclk));
	jdff dff_A_dHVanQTw5_2(.dout(w_n614_3[2]),.din(w_dff_A_dHVanQTw5_2),.clk(gclk));
	jdff dff_A_Nyew7vER2_2(.dout(w_dff_A_dHVanQTw5_2),.din(w_dff_A_Nyew7vER2_2),.clk(gclk));
	jdff dff_A_wqkhJfN54_2(.dout(w_dff_A_Nyew7vER2_2),.din(w_dff_A_wqkhJfN54_2),.clk(gclk));
	jdff dff_A_Zi7TV5ts4_2(.dout(w_dff_A_wqkhJfN54_2),.din(w_dff_A_Zi7TV5ts4_2),.clk(gclk));
	jdff dff_A_hwu55APx7_2(.dout(w_dff_A_Zi7TV5ts4_2),.din(w_dff_A_hwu55APx7_2),.clk(gclk));
	jdff dff_A_K1yCmZ129_2(.dout(w_dff_A_hwu55APx7_2),.din(w_dff_A_K1yCmZ129_2),.clk(gclk));
	jdff dff_A_FmQ1WqRS3_2(.dout(w_dff_A_K1yCmZ129_2),.din(w_dff_A_FmQ1WqRS3_2),.clk(gclk));
	jdff dff_A_nkb3mWIg6_2(.dout(w_dff_A_FmQ1WqRS3_2),.din(w_dff_A_nkb3mWIg6_2),.clk(gclk));
	jdff dff_A_XOHknlG88_2(.dout(w_dff_A_nkb3mWIg6_2),.din(w_dff_A_XOHknlG88_2),.clk(gclk));
	jdff dff_A_Lq4xPcLF3_1(.dout(w_n601_0[1]),.din(w_dff_A_Lq4xPcLF3_1),.clk(gclk));
	jdff dff_A_GsUCtSeh1_1(.dout(w_dff_A_Lq4xPcLF3_1),.din(w_dff_A_GsUCtSeh1_1),.clk(gclk));
	jdff dff_A_rV0vbByL7_0(.dout(w_n600_1[0]),.din(w_dff_A_rV0vbByL7_0),.clk(gclk));
	jdff dff_A_mUoU2YLO5_1(.dout(w_n600_1[1]),.din(w_dff_A_mUoU2YLO5_1),.clk(gclk));
	jdff dff_A_wN72twRj6_1(.dout(w_dff_A_mUoU2YLO5_1),.din(w_dff_A_wN72twRj6_1),.clk(gclk));
	jdff dff_B_STIrPms96_0(.din(n599),.dout(w_dff_B_STIrPms96_0),.clk(gclk));
	jdff dff_A_psZ4pvPn6_0(.dout(w_n598_0[0]),.din(w_dff_A_psZ4pvPn6_0),.clk(gclk));
	jdff dff_A_mGCpcx5X1_0(.dout(w_dff_A_psZ4pvPn6_0),.din(w_dff_A_mGCpcx5X1_0),.clk(gclk));
	jdff dff_A_xy45DvJ30_1(.dout(w_n571_1[1]),.din(w_dff_A_xy45DvJ30_1),.clk(gclk));
	jdff dff_A_D6gbvKTe2_1(.dout(w_dff_A_xy45DvJ30_1),.din(w_dff_A_D6gbvKTe2_1),.clk(gclk));
	jdff dff_A_dcoKiQBF6_1(.dout(w_dff_A_D6gbvKTe2_1),.din(w_dff_A_dcoKiQBF6_1),.clk(gclk));
	jdff dff_A_BlOSIGtz5_1(.dout(w_dff_A_dcoKiQBF6_1),.din(w_dff_A_BlOSIGtz5_1),.clk(gclk));
	jdff dff_A_UDYrwmQr2_1(.dout(w_dff_A_BlOSIGtz5_1),.din(w_dff_A_UDYrwmQr2_1),.clk(gclk));
	jdff dff_B_vcISusnL7_0(.din(n589),.dout(w_dff_B_vcISusnL7_0),.clk(gclk));
	jdff dff_B_rBoAC2sS8_0(.din(w_dff_B_vcISusnL7_0),.dout(w_dff_B_rBoAC2sS8_0),.clk(gclk));
	jdff dff_A_WW3mbcMB1_1(.dout(w_n548_0[1]),.din(w_dff_A_WW3mbcMB1_1),.clk(gclk));
	jdff dff_A_fFhQYuH08_1(.dout(w_dff_A_WW3mbcMB1_1),.din(w_dff_A_fFhQYuH08_1),.clk(gclk));
	jdff dff_A_I6SmfvYh6_1(.dout(w_n347_0[1]),.din(w_dff_A_I6SmfvYh6_1),.clk(gclk));
	jdff dff_A_I6R4qOpr9_1(.dout(w_n189_1[1]),.din(w_dff_A_I6R4qOpr9_1),.clk(gclk));
	jdff dff_A_CwkCNF3L1_1(.dout(w_dff_A_I6R4qOpr9_1),.din(w_dff_A_CwkCNF3L1_1),.clk(gclk));
	jdff dff_A_IvJ5Yk489_0(.dout(w_n282_0[0]),.din(w_dff_A_IvJ5Yk489_0),.clk(gclk));
	jdff dff_B_OrLSHVmi8_1(.din(n525),.dout(w_dff_B_OrLSHVmi8_1),.clk(gclk));
	jdff dff_B_azq4YLDP6_1(.din(n538),.dout(w_dff_B_azq4YLDP6_1),.clk(gclk));
	jdff dff_B_acPEU2UT6_1(.din(n324),.dout(w_dff_B_acPEU2UT6_1),.clk(gclk));
	jdff dff_A_8l4yuvmS0_1(.dout(w_n323_0[1]),.din(w_dff_A_8l4yuvmS0_1),.clk(gclk));
	jdff dff_A_BhmWJ5Xk8_2(.dout(w_n323_0[2]),.din(w_dff_A_BhmWJ5Xk8_2),.clk(gclk));
	jdff dff_B_L6k4xnL21_1(.din(n314),.dout(w_dff_B_L6k4xnL21_1),.clk(gclk));
	jdff dff_B_RxrF3lmL5_1(.din(w_dff_B_L6k4xnL21_1),.dout(w_dff_B_RxrF3lmL5_1),.clk(gclk));
	jdff dff_A_CJmQAE0W4_2(.dout(w_G20_3[2]),.din(w_dff_A_CJmQAE0W4_2),.clk(gclk));
	jdff dff_A_uBod4A164_1(.dout(w_n141_1[1]),.din(w_dff_A_uBod4A164_1),.clk(gclk));
	jdff dff_A_6qfkpFnA6_2(.dout(w_n141_1[2]),.din(w_dff_A_6qfkpFnA6_2),.clk(gclk));
	jdff dff_A_VOUHRpC53_0(.dout(w_n334_0[0]),.din(w_dff_A_VOUHRpC53_0),.clk(gclk));
	jdff dff_A_iYvogae46_0(.dout(w_dff_A_VOUHRpC53_0),.din(w_dff_A_iYvogae46_0),.clk(gclk));
	jdff dff_A_gaaqrNnu9_0(.dout(w_G169_2[0]),.din(w_dff_A_gaaqrNnu9_0),.clk(gclk));
	jdff dff_A_myzdZv9H0_1(.dout(w_G169_2[1]),.din(w_dff_A_myzdZv9H0_1),.clk(gclk));
	jdff dff_A_CZyKlEfI8_1(.dout(w_dff_A_myzdZv9H0_1),.din(w_dff_A_CZyKlEfI8_1),.clk(gclk));
	jdff dff_B_vGb3QaKr3_0(.din(n342),.dout(w_dff_B_vGb3QaKr3_0),.clk(gclk));
	jdff dff_A_UH2mw9IG9_1(.dout(w_n321_0[1]),.din(w_dff_A_UH2mw9IG9_1),.clk(gclk));
	jdff dff_A_v6Kexx641_1(.dout(w_dff_A_UH2mw9IG9_1),.din(w_dff_A_v6Kexx641_1),.clk(gclk));
	jdff dff_B_aDt2lZxg4_1(.din(n336),.dout(w_dff_B_aDt2lZxg4_1),.clk(gclk));
	jdff dff_A_lGjIW0tb1_2(.dout(w_n72_1[2]),.din(w_dff_A_lGjIW0tb1_2),.clk(gclk));
	jdff dff_A_ZVkHsFxW5_2(.dout(w_dff_A_lGjIW0tb1_2),.din(w_dff_A_ZVkHsFxW5_2),.clk(gclk));
	jdff dff_A_Wn6G64x50_1(.dout(w_n72_0[1]),.din(w_dff_A_Wn6G64x50_1),.clk(gclk));
	jdff dff_A_P5CCnnsY7_1(.dout(w_dff_A_Wn6G64x50_1),.din(w_dff_A_P5CCnnsY7_1),.clk(gclk));
	jdff dff_A_vIN32VZI0_1(.dout(w_dff_A_P5CCnnsY7_1),.din(w_dff_A_vIN32VZI0_1),.clk(gclk));
	jdff dff_A_UjcH846S9_1(.dout(w_dff_A_vIN32VZI0_1),.din(w_dff_A_UjcH846S9_1),.clk(gclk));
	jdff dff_A_ugurzdDE3_2(.dout(w_n72_0[2]),.din(w_dff_A_ugurzdDE3_2),.clk(gclk));
	jdff dff_A_AOrGp42Y8_2(.dout(w_dff_A_ugurzdDE3_2),.din(w_dff_A_AOrGp42Y8_2),.clk(gclk));
	jdff dff_A_4IRxXou16_0(.dout(w_n315_0[0]),.din(w_dff_A_4IRxXou16_0),.clk(gclk));
	jdff dff_A_4u1g0nRA4_0(.dout(w_dff_A_4IRxXou16_0),.din(w_dff_A_4u1g0nRA4_0),.clk(gclk));
	jdff dff_A_c0kaHqI69_2(.dout(w_n315_0[2]),.din(w_dff_A_c0kaHqI69_2),.clk(gclk));
	jdff dff_A_sABhtlWN3_2(.dout(w_dff_A_c0kaHqI69_2),.din(w_dff_A_sABhtlWN3_2),.clk(gclk));
	jdff dff_A_ugfSWE8Z0_1(.dout(w_G33_8[1]),.din(w_dff_A_ugfSWE8Z0_1),.clk(gclk));
	jdff dff_A_S3P8vT1S3_0(.dout(w_n313_0[0]),.din(w_dff_A_S3P8vT1S3_0),.clk(gclk));
	jdff dff_A_hyYF8zgZ9_0(.dout(w_dff_A_S3P8vT1S3_0),.din(w_dff_A_hyYF8zgZ9_0),.clk(gclk));
	jdff dff_A_PoKWS1oL5_0(.dout(w_dff_A_hyYF8zgZ9_0),.din(w_dff_A_PoKWS1oL5_0),.clk(gclk));
	jdff dff_A_4f98VY5J0_0(.dout(w_n312_0[0]),.din(w_dff_A_4f98VY5J0_0),.clk(gclk));
	jdff dff_A_r52exDBL5_0(.dout(w_n310_0[0]),.din(w_dff_A_r52exDBL5_0),.clk(gclk));
	jdff dff_A_UL17uMyz6_1(.dout(w_n309_0[1]),.din(w_dff_A_UL17uMyz6_1),.clk(gclk));
	jdff dff_A_lCjPuVzC0_1(.dout(w_dff_A_UL17uMyz6_1),.din(w_dff_A_lCjPuVzC0_1),.clk(gclk));
	jdff dff_A_zQqKriJB3_0(.dout(w_n94_0[0]),.din(w_dff_A_zQqKriJB3_0),.clk(gclk));
	jdff dff_A_KOZBvQqa7_0(.dout(w_dff_A_zQqKriJB3_0),.din(w_dff_A_KOZBvQqa7_0),.clk(gclk));
	jdff dff_A_2fVsdO4y2_0(.dout(w_dff_A_KOZBvQqa7_0),.din(w_dff_A_2fVsdO4y2_0),.clk(gclk));
	jdff dff_A_DBtIjgyf7_0(.dout(w_G244_1[0]),.din(w_dff_A_DBtIjgyf7_0),.clk(gclk));
	jdff dff_A_T04A5Jm83_0(.dout(w_n298_0[0]),.din(w_dff_A_T04A5Jm83_0),.clk(gclk));
	jdff dff_A_09glOBoH0_0(.dout(w_dff_A_T04A5Jm83_0),.din(w_dff_A_09glOBoH0_0),.clk(gclk));
	jdff dff_A_EW6FVQyj1_0(.dout(w_G190_3[0]),.din(w_dff_A_EW6FVQyj1_0),.clk(gclk));
	jdff dff_A_pI5UWDYu8_0(.dout(w_dff_A_EW6FVQyj1_0),.din(w_dff_A_pI5UWDYu8_0),.clk(gclk));
	jdff dff_A_K3q8J32N3_1(.dout(w_G190_3[1]),.din(w_dff_A_K3q8J32N3_1),.clk(gclk));
	jdff dff_A_rkfMiR059_1(.dout(w_dff_A_K3q8J32N3_1),.din(w_dff_A_rkfMiR059_1),.clk(gclk));
	jdff dff_A_Gm4CyLtF8_1(.dout(w_n534_0[1]),.din(w_dff_A_Gm4CyLtF8_1),.clk(gclk));
	jdff dff_A_V6jSsjcw7_1(.dout(w_n507_2[1]),.din(w_dff_A_V6jSsjcw7_1),.clk(gclk));
	jdff dff_B_zLrZuBmg2_0(.din(n270),.dout(w_dff_B_zLrZuBmg2_0),.clk(gclk));
	jdff dff_B_0yChTZMT8_1(.din(n263),.dout(w_dff_B_0yChTZMT8_1),.clk(gclk));
	jdff dff_A_WruRIkvC8_0(.dout(w_n151_5[0]),.din(w_dff_A_WruRIkvC8_0),.clk(gclk));
	jdff dff_A_Maqp9vwT3_1(.dout(w_n261_0[1]),.din(w_dff_A_Maqp9vwT3_1),.clk(gclk));
	jdff dff_A_7UT1Tdcn2_1(.dout(w_dff_A_Maqp9vwT3_1),.din(w_dff_A_7UT1Tdcn2_1),.clk(gclk));
	jdff dff_A_IAiOz3ZI6_2(.dout(w_n261_0[2]),.din(w_dff_A_IAiOz3ZI6_2),.clk(gclk));
	jdff dff_A_FZAOHU4A3_2(.dout(w_dff_A_IAiOz3ZI6_2),.din(w_dff_A_FZAOHU4A3_2),.clk(gclk));
	jdff dff_A_HKxjezPj9_1(.dout(w_n283_0[1]),.din(w_dff_A_HKxjezPj9_1),.clk(gclk));
	jdff dff_A_0C1uqOXc6_0(.dout(w_n168_3[0]),.din(w_dff_A_0C1uqOXc6_0),.clk(gclk));
	jdff dff_A_ojfbe8eC4_2(.dout(w_n168_3[2]),.din(w_dff_A_ojfbe8eC4_2),.clk(gclk));
	jdff dff_A_aIBsKakw8_2(.dout(w_dff_A_ojfbe8eC4_2),.din(w_dff_A_aIBsKakw8_2),.clk(gclk));
	jdff dff_A_Q4Evzbr60_0(.dout(w_n269_0[0]),.din(w_dff_A_Q4Evzbr60_0),.clk(gclk));
	jdff dff_A_ZNRnTKv70_0(.dout(w_dff_A_Q4Evzbr60_0),.din(w_dff_A_ZNRnTKv70_0),.clk(gclk));
	jdff dff_A_s9hBFqu00_0(.dout(w_n262_0[0]),.din(w_dff_A_s9hBFqu00_0),.clk(gclk));
	jdff dff_A_HmUdrO5U0_0(.dout(w_dff_A_s9hBFqu00_0),.din(w_dff_A_HmUdrO5U0_0),.clk(gclk));
	jdff dff_A_cu6nqP592_1(.dout(w_n262_0[1]),.din(w_dff_A_cu6nqP592_1),.clk(gclk));
	jdff dff_A_jIEF3LPd4_1(.dout(w_dff_A_cu6nqP592_1),.din(w_dff_A_jIEF3LPd4_1),.clk(gclk));
	jdff dff_A_LFqTsjbc6_0(.dout(w_G33_9[0]),.din(w_dff_A_LFqTsjbc6_0),.clk(gclk));
	jdff dff_A_YBop4ogN4_1(.dout(w_G33_9[1]),.din(w_dff_A_YBop4ogN4_1),.clk(gclk));
	jdff dff_A_d4Ac9V5o7_1(.dout(w_n260_0[1]),.din(w_dff_A_d4Ac9V5o7_1),.clk(gclk));
	jdff dff_A_Mk9d0q7l7_1(.dout(w_G20_4[1]),.din(w_dff_A_Mk9d0q7l7_1),.clk(gclk));
	jdff dff_A_ptBuZUVv8_2(.dout(w_G20_4[2]),.din(w_dff_A_ptBuZUVv8_2),.clk(gclk));
	jdff dff_A_bzBoME3G6_2(.dout(w_dff_A_ptBuZUVv8_2),.din(w_dff_A_bzBoME3G6_2),.clk(gclk));
	jdff dff_A_Q2RwdHnB6_1(.dout(w_n257_0[1]),.din(w_dff_A_Q2RwdHnB6_1),.clk(gclk));
	jdff dff_A_y6QJ2NYk0_1(.dout(w_n256_0[1]),.din(w_dff_A_y6QJ2NYk0_1),.clk(gclk));
	jdff dff_A_LKGd0RP57_0(.dout(w_n251_0[0]),.din(w_dff_A_LKGd0RP57_0),.clk(gclk));
	jdff dff_A_5pvZ8Iej6_1(.dout(w_n250_0[1]),.din(w_dff_A_5pvZ8Iej6_1),.clk(gclk));
	jdff dff_A_jJRwyNRU9_1(.dout(w_n247_0[1]),.din(w_dff_A_jJRwyNRU9_1),.clk(gclk));
	jdff dff_A_VMpsqkN26_0(.dout(w_G238_0[0]),.din(w_dff_A_VMpsqkN26_0),.clk(gclk));
	jdff dff_A_MgaHJqQP3_0(.dout(w_dff_A_VMpsqkN26_0),.din(w_dff_A_MgaHJqQP3_0),.clk(gclk));
	jdff dff_A_WGcIau8i4_0(.dout(w_dff_A_MgaHJqQP3_0),.din(w_dff_A_WGcIau8i4_0),.clk(gclk));
	jdff dff_A_kslexxj42_1(.dout(w_G238_0[1]),.din(w_dff_A_kslexxj42_1),.clk(gclk));
	jdff dff_A_vm0PmMfd2_1(.dout(w_dff_A_kslexxj42_1),.din(w_dff_A_vm0PmMfd2_1),.clk(gclk));
	jdff dff_A_lUeRqMzZ6_0(.dout(w_n243_0[0]),.din(w_dff_A_lUeRqMzZ6_0),.clk(gclk));
	jdff dff_A_Lyne1nuA5_1(.dout(w_G244_0[1]),.din(w_dff_A_Lyne1nuA5_1),.clk(gclk));
	jdff dff_A_xBgHXuCO4_1(.dout(w_dff_A_Lyne1nuA5_1),.din(w_dff_A_xBgHXuCO4_1),.clk(gclk));
	jdff dff_A_Yh9u04z25_2(.dout(w_G244_0[2]),.din(w_dff_A_Yh9u04z25_2),.clk(gclk));
	jdff dff_A_a4qbyPcr0_2(.dout(w_dff_A_Yh9u04z25_2),.din(w_dff_A_a4qbyPcr0_2),.clk(gclk));
	jdff dff_A_ONNWueaN8_1(.dout(w_n388_1[1]),.din(w_dff_A_ONNWueaN8_1),.clk(gclk));
	jdff dff_A_JHn4h5fV4_2(.dout(w_n388_1[2]),.din(w_dff_A_JHn4h5fV4_2),.clk(gclk));
	jdff dff_A_JoHpLu1U0_2(.dout(w_dff_A_JHn4h5fV4_2),.din(w_dff_A_JoHpLu1U0_2),.clk(gclk));
	jdff dff_A_xbHy7meL8_0(.dout(w_n520_0[0]),.din(w_dff_A_xbHy7meL8_0),.clk(gclk));
	jdff dff_A_SqJOrxYE3_0(.dout(w_dff_A_xbHy7meL8_0),.din(w_dff_A_SqJOrxYE3_0),.clk(gclk));
	jdff dff_A_h97w8Uuz8_0(.dout(w_n604_1[0]),.din(w_dff_A_h97w8Uuz8_0),.clk(gclk));
	jdff dff_A_q04uKjDl0_0(.dout(w_dff_A_h97w8Uuz8_0),.din(w_dff_A_q04uKjDl0_0),.clk(gclk));
	jdff dff_A_XbByAM9Z5_1(.dout(w_n604_1[1]),.din(w_dff_A_XbByAM9Z5_1),.clk(gclk));
	jdff dff_A_VK0Jemwn8_1(.dout(w_dff_A_XbByAM9Z5_1),.din(w_dff_A_VK0Jemwn8_1),.clk(gclk));
	jdff dff_A_lk2PBJq41_0(.dout(w_n861_0[0]),.din(w_dff_A_lk2PBJq41_0),.clk(gclk));
	jdff dff_B_Fsh1G4pF3_0(.din(n858),.dout(w_dff_B_Fsh1G4pF3_0),.clk(gclk));
	jdff dff_A_4EkeUj953_2(.dout(w_n579_0[2]),.din(w_dff_A_4EkeUj953_2),.clk(gclk));
	jdff dff_B_7izUGPf87_0(.din(n578),.dout(w_dff_B_7izUGPf87_0),.clk(gclk));
	jdff dff_B_7kdH1aLg2_0(.din(w_dff_B_7izUGPf87_0),.dout(w_dff_B_7kdH1aLg2_0),.clk(gclk));
	jdff dff_B_YHsPo9ub3_0(.din(w_dff_B_7kdH1aLg2_0),.dout(w_dff_B_YHsPo9ub3_0),.clk(gclk));
	jdff dff_A_pyvMT0dW7_0(.dout(w_n571_2[0]),.din(w_dff_A_pyvMT0dW7_0),.clk(gclk));
	jdff dff_A_ubAFFJDR1_0(.dout(w_dff_A_pyvMT0dW7_0),.din(w_dff_A_ubAFFJDR1_0),.clk(gclk));
	jdff dff_A_eNjzWxfS2_1(.dout(w_n571_0[1]),.din(w_dff_A_eNjzWxfS2_1),.clk(gclk));
	jdff dff_A_0YNUmbHB5_1(.dout(w_dff_A_eNjzWxfS2_1),.din(w_dff_A_0YNUmbHB5_1),.clk(gclk));
	jdff dff_A_BeM6e52w4_2(.dout(w_n571_0[2]),.din(w_dff_A_BeM6e52w4_2),.clk(gclk));
	jdff dff_A_tA6eYaIu4_2(.dout(w_dff_A_BeM6e52w4_2),.din(w_dff_A_tA6eYaIu4_2),.clk(gclk));
	jdff dff_B_FCYgFZDb8_3(.din(n571),.dout(w_dff_B_FCYgFZDb8_3),.clk(gclk));
	jdff dff_B_Dgf2wMUK4_3(.din(w_dff_B_FCYgFZDb8_3),.dout(w_dff_B_Dgf2wMUK4_3),.clk(gclk));
	jdff dff_B_0mSZYAmZ8_3(.din(w_dff_B_Dgf2wMUK4_3),.dout(w_dff_B_0mSZYAmZ8_3),.clk(gclk));
	jdff dff_B_leZnMZJz3_3(.din(w_dff_B_0mSZYAmZ8_3),.dout(w_dff_B_leZnMZJz3_3),.clk(gclk));
	jdff dff_B_fj0fuCCv9_3(.din(w_dff_B_leZnMZJz3_3),.dout(w_dff_B_fj0fuCCv9_3),.clk(gclk));
	jdff dff_A_C6mqboJQ1_1(.dout(w_n567_5[1]),.din(w_dff_A_C6mqboJQ1_1),.clk(gclk));
	jdff dff_A_yg7TGh7s4_1(.dout(w_dff_A_C6mqboJQ1_1),.din(w_dff_A_yg7TGh7s4_1),.clk(gclk));
	jdff dff_A_dMFM4oPT9_1(.dout(w_dff_A_yg7TGh7s4_1),.din(w_dff_A_dMFM4oPT9_1),.clk(gclk));
	jdff dff_A_0v9d9oYZ3_1(.dout(w_dff_A_dMFM4oPT9_1),.din(w_dff_A_0v9d9oYZ3_1),.clk(gclk));
	jdff dff_A_Nbk5Aqs47_1(.dout(w_dff_A_0v9d9oYZ3_1),.din(w_dff_A_Nbk5Aqs47_1),.clk(gclk));
	jdff dff_A_fRorsgP65_1(.dout(w_dff_A_Nbk5Aqs47_1),.din(w_dff_A_fRorsgP65_1),.clk(gclk));
	jdff dff_A_b8cO9g9e4_0(.dout(w_n570_0[0]),.din(w_dff_A_b8cO9g9e4_0),.clk(gclk));
	jdff dff_A_Gva2bMP27_1(.dout(w_n242_0[1]),.din(w_dff_A_Gva2bMP27_1),.clk(gclk));
	jdff dff_A_MeHRTeA34_1(.dout(w_dff_A_Gva2bMP27_1),.din(w_dff_A_MeHRTeA34_1),.clk(gclk));
	jdff dff_A_tCXveOjQ6_2(.dout(w_n242_0[2]),.din(w_dff_A_tCXveOjQ6_2),.clk(gclk));
	jdff dff_A_pbCCveUn4_1(.dout(w_n238_0[1]),.din(w_dff_A_pbCCveUn4_1),.clk(gclk));
	jdff dff_A_UM007gqd4_1(.dout(w_n237_0[1]),.din(w_dff_A_UM007gqd4_1),.clk(gclk));
	jdff dff_A_1H4g7aOH3_1(.dout(w_dff_A_UM007gqd4_1),.din(w_dff_A_1H4g7aOH3_1),.clk(gclk));
	jdff dff_A_sSWuGHby9_1(.dout(w_n234_0[1]),.din(w_dff_A_sSWuGHby9_1),.clk(gclk));
	jdff dff_A_KXepKQry7_1(.dout(w_dff_A_sSWuGHby9_1),.din(w_dff_A_KXepKQry7_1),.clk(gclk));
	jdff dff_A_Bc6Smvon8_1(.dout(w_dff_A_KXepKQry7_1),.din(w_dff_A_Bc6Smvon8_1),.clk(gclk));
	jdff dff_B_H5DWbEEY9_1(.din(n226),.dout(w_dff_B_H5DWbEEY9_1),.clk(gclk));
	jdff dff_A_ehyGtSRL7_1(.dout(w_n229_0[1]),.din(w_dff_A_ehyGtSRL7_1),.clk(gclk));
	jdff dff_B_l6ynPKtQ1_1(.din(n227),.dout(w_dff_B_l6ynPKtQ1_1),.clk(gclk));
	jdff dff_B_vjIuho306_1(.din(w_dff_B_l6ynPKtQ1_1),.dout(w_dff_B_vjIuho306_1),.clk(gclk));
	jdff dff_A_m0U3yfr82_0(.dout(w_n224_1[0]),.din(w_dff_A_m0U3yfr82_0),.clk(gclk));
	jdff dff_A_t9qhoLV72_2(.dout(w_n224_0[2]),.din(w_dff_A_t9qhoLV72_2),.clk(gclk));
	jdff dff_B_3956jpsI0_0(.din(n223),.dout(w_dff_B_3956jpsI0_0),.clk(gclk));
	jdff dff_B_v4umk7t39_1(.din(n217),.dout(w_dff_B_v4umk7t39_1),.clk(gclk));
	jdff dff_A_jTypQ46G6_1(.dout(w_n218_0[1]),.din(w_dff_A_jTypQ46G6_1),.clk(gclk));
	jdff dff_A_y5iOTmpa2_0(.dout(w_n141_2[0]),.din(w_dff_A_y5iOTmpa2_0),.clk(gclk));
	jdff dff_B_b6QY8yMK0_0(.din(n216),.dout(w_dff_B_b6QY8yMK0_0),.clk(gclk));
	jdff dff_A_wpDTwxvd2_0(.dout(w_n81_1[0]),.din(w_dff_A_wpDTwxvd2_0),.clk(gclk));
	jdff dff_A_hlo8UFjr6_1(.dout(w_n213_0[1]),.din(w_dff_A_hlo8UFjr6_1),.clk(gclk));
	jdff dff_A_E0X6eWJ73_1(.dout(w_n212_0[1]),.din(w_dff_A_E0X6eWJ73_1),.clk(gclk));
	jdff dff_A_BlTCyyYc9_1(.dout(w_dff_A_E0X6eWJ73_1),.din(w_dff_A_BlTCyyYc9_1),.clk(gclk));
	jdff dff_A_bViPQEmR9_0(.dout(w_n207_0[0]),.din(w_dff_A_bViPQEmR9_0),.clk(gclk));
	jdff dff_A_JqIje15q7_2(.dout(w_n84_1[2]),.din(w_dff_A_JqIje15q7_2),.clk(gclk));
	jdff dff_A_4Z7QsvPG7_1(.dout(w_n84_0[1]),.din(w_dff_A_4Z7QsvPG7_1),.clk(gclk));
	jdff dff_A_9Zcfe4AD1_2(.dout(w_n84_0[2]),.din(w_dff_A_9Zcfe4AD1_2),.clk(gclk));
	jdff dff_A_XtgaX3F38_0(.dout(w_G250_0[0]),.din(w_dff_A_XtgaX3F38_0),.clk(gclk));
	jdff dff_A_UifMbqcT0_0(.dout(w_dff_A_XtgaX3F38_0),.din(w_dff_A_UifMbqcT0_0),.clk(gclk));
	jdff dff_A_eQ84Agja2_1(.dout(w_n202_0[1]),.din(w_dff_A_eQ84Agja2_1),.clk(gclk));
	jdff dff_A_GS59ELfG3_1(.dout(w_n201_0[1]),.din(w_dff_A_GS59ELfG3_1),.clk(gclk));
	jdff dff_A_smOwfoRH9_1(.dout(w_dff_A_GS59ELfG3_1),.din(w_dff_A_smOwfoRH9_1),.clk(gclk));
	jdff dff_A_dZlq84rC4_0(.dout(w_n168_4[0]),.din(w_dff_A_dZlq84rC4_0),.clk(gclk));
	jdff dff_A_ezplO8FG1_0(.dout(w_dff_A_dZlq84rC4_0),.din(w_dff_A_ezplO8FG1_0),.clk(gclk));
	jdff dff_A_9GkQ8nxk7_1(.dout(w_n168_4[1]),.din(w_dff_A_9GkQ8nxk7_1),.clk(gclk));
	jdff dff_A_UT5E5WLW6_1(.dout(w_dff_A_9GkQ8nxk7_1),.din(w_dff_A_UT5E5WLW6_1),.clk(gclk));
	jdff dff_A_zwpxlafl6_0(.dout(w_n199_0[0]),.din(w_dff_A_zwpxlafl6_0),.clk(gclk));
	jdff dff_A_mCUAmSWn7_0(.dout(w_dff_A_zwpxlafl6_0),.din(w_dff_A_mCUAmSWn7_0),.clk(gclk));
	jdff dff_A_kq9R0Hx92_0(.dout(w_dff_A_mCUAmSWn7_0),.din(w_dff_A_kq9R0Hx92_0),.clk(gclk));
	jdff dff_A_d9JyWCYQ8_2(.dout(w_n199_0[2]),.din(w_dff_A_d9JyWCYQ8_2),.clk(gclk));
	jdff dff_B_1o0b1wRq7_3(.din(n199),.dout(w_dff_B_1o0b1wRq7_3),.clk(gclk));
	jdff dff_B_2fIvKTzI6_3(.din(w_dff_B_1o0b1wRq7_3),.dout(w_dff_B_2fIvKTzI6_3),.clk(gclk));
	jdff dff_B_n66BveGg3_3(.din(w_dff_B_2fIvKTzI6_3),.dout(w_dff_B_n66BveGg3_3),.clk(gclk));
	jdff dff_B_dQmmLHRO0_3(.din(w_dff_B_n66BveGg3_3),.dout(w_dff_B_dQmmLHRO0_3),.clk(gclk));
	jdff dff_B_kMTbtHbg6_3(.din(w_dff_B_dQmmLHRO0_3),.dout(w_dff_B_kMTbtHbg6_3),.clk(gclk));
	jdff dff_B_ffUfftvl6_3(.din(w_dff_B_kMTbtHbg6_3),.dout(w_dff_B_ffUfftvl6_3),.clk(gclk));
	jdff dff_A_2TRl5kqn1_0(.dout(w_n577_0[0]),.din(w_dff_A_2TRl5kqn1_0),.clk(gclk));
	jdff dff_A_f3ju7Xvn3_0(.dout(w_dff_A_2TRl5kqn1_0),.din(w_dff_A_f3ju7Xvn3_0),.clk(gclk));
	jdff dff_B_iXyxHpsb3_2(.din(n1164),.dout(w_dff_B_iXyxHpsb3_2),.clk(gclk));
	jdff dff_B_mXIarFpT2_2(.din(w_dff_B_iXyxHpsb3_2),.dout(w_dff_B_mXIarFpT2_2),.clk(gclk));
	jdff dff_B_CnME2FJ40_2(.din(w_dff_B_mXIarFpT2_2),.dout(w_dff_B_CnME2FJ40_2),.clk(gclk));
	jdff dff_B_W7UKalJt1_2(.din(w_dff_B_CnME2FJ40_2),.dout(w_dff_B_W7UKalJt1_2),.clk(gclk));
	jdff dff_B_7dexFQRr4_1(.din(n617),.dout(w_dff_B_7dexFQRr4_1),.clk(gclk));
	jdff dff_B_3KsAx5iO0_0(.din(n698),.dout(w_dff_B_3KsAx5iO0_0),.clk(gclk));
	jdff dff_B_hoiOK8je7_0(.din(n697),.dout(w_dff_B_hoiOK8je7_0),.clk(gclk));
	jdff dff_B_eIU6FKJH2_0(.din(w_dff_B_hoiOK8je7_0),.dout(w_dff_B_eIU6FKJH2_0),.clk(gclk));
	jdff dff_B_H2ok2CHD2_0(.din(n694),.dout(w_dff_B_H2ok2CHD2_0),.clk(gclk));
	jdff dff_B_2uiw1TE68_0(.din(w_dff_B_H2ok2CHD2_0),.dout(w_dff_B_2uiw1TE68_0),.clk(gclk));
	jdff dff_A_Icil9oyk6_0(.dout(w_n692_0[0]),.din(w_dff_A_Icil9oyk6_0),.clk(gclk));
	jdff dff_A_HV5MqwNv4_0(.dout(w_n153_4[0]),.din(w_dff_A_HV5MqwNv4_0),.clk(gclk));
	jdff dff_A_wCY4BIU75_0(.dout(w_dff_A_HV5MqwNv4_0),.din(w_dff_A_wCY4BIU75_0),.clk(gclk));
	jdff dff_A_FJXwIsoD3_0(.dout(w_dff_A_wCY4BIU75_0),.din(w_dff_A_FJXwIsoD3_0),.clk(gclk));
	jdff dff_A_B099aipu7_0(.dout(w_dff_A_FJXwIsoD3_0),.din(w_dff_A_B099aipu7_0),.clk(gclk));
	jdff dff_A_I9OoPHr58_0(.dout(w_dff_A_B099aipu7_0),.din(w_dff_A_I9OoPHr58_0),.clk(gclk));
	jdff dff_A_3RdTVT158_0(.dout(w_dff_A_I9OoPHr58_0),.din(w_dff_A_3RdTVT158_0),.clk(gclk));
	jdff dff_A_0mHxmi5c9_1(.dout(w_n153_4[1]),.din(w_dff_A_0mHxmi5c9_1),.clk(gclk));
	jdff dff_A_prntjCou7_1(.dout(w_dff_A_0mHxmi5c9_1),.din(w_dff_A_prntjCou7_1),.clk(gclk));
	jdff dff_A_YJ7N1I1O6_1(.dout(w_dff_A_prntjCou7_1),.din(w_dff_A_YJ7N1I1O6_1),.clk(gclk));
	jdff dff_A_u93sXQNP5_1(.dout(w_dff_A_YJ7N1I1O6_1),.din(w_dff_A_u93sXQNP5_1),.clk(gclk));
	jdff dff_A_zIyt1ZDW7_1(.dout(w_dff_A_u93sXQNP5_1),.din(w_dff_A_zIyt1ZDW7_1),.clk(gclk));
	jdff dff_A_2tQIXM091_0(.dout(w_G355_0),.din(w_dff_A_2tQIXM091_0),.clk(gclk));
	jdff dff_A_BXp19r1I9_2(.dout(w_n81_0[2]),.din(w_dff_A_BXp19r1I9_2),.clk(gclk));
	jdff dff_A_Gtl4BAO57_2(.dout(w_dff_A_BXp19r1I9_2),.din(w_dff_A_Gtl4BAO57_2),.clk(gclk));
	jdff dff_A_NKXy33Zt9_2(.dout(w_dff_A_Gtl4BAO57_2),.din(w_dff_A_NKXy33Zt9_2),.clk(gclk));
	jdff dff_A_FSrO6w4K0_0(.dout(w_G107_4[0]),.din(w_dff_A_FSrO6w4K0_0),.clk(gclk));
	jdff dff_A_bZCkoJDo6_0(.dout(w_dff_A_FSrO6w4K0_0),.din(w_dff_A_bZCkoJDo6_0),.clk(gclk));
	jdff dff_A_6VTTiOdz4_0(.dout(w_dff_A_bZCkoJDo6_0),.din(w_dff_A_6VTTiOdz4_0),.clk(gclk));
	jdff dff_A_Y0dcH6Gw9_0(.dout(w_dff_A_6VTTiOdz4_0),.din(w_dff_A_Y0dcH6Gw9_0),.clk(gclk));
	jdff dff_A_DcO9EYeb0_0(.dout(w_dff_A_Y0dcH6Gw9_0),.din(w_dff_A_DcO9EYeb0_0),.clk(gclk));
	jdff dff_A_ieJJYPRg7_0(.dout(w_dff_A_DcO9EYeb0_0),.din(w_dff_A_ieJJYPRg7_0),.clk(gclk));
	jdff dff_A_VBAT3ybe9_1(.dout(w_G107_1[1]),.din(w_dff_A_VBAT3ybe9_1),.clk(gclk));
	jdff dff_A_2Ub4ESG99_1(.dout(w_dff_A_VBAT3ybe9_1),.din(w_dff_A_2Ub4ESG99_1),.clk(gclk));
	jdff dff_A_6ineyHI54_1(.dout(w_dff_A_2Ub4ESG99_1),.din(w_dff_A_6ineyHI54_1),.clk(gclk));
	jdff dff_A_zThGJpvx2_2(.dout(w_G107_1[2]),.din(w_dff_A_zThGJpvx2_2),.clk(gclk));
	jdff dff_A_diHCYZvR4_2(.dout(w_dff_A_zThGJpvx2_2),.din(w_dff_A_diHCYZvR4_2),.clk(gclk));
	jdff dff_A_AfTxsI4D4_2(.dout(w_dff_A_diHCYZvR4_2),.din(w_dff_A_AfTxsI4D4_2),.clk(gclk));
	jdff dff_A_ZqrpNP8R5_1(.dout(w_n80_0[1]),.din(w_dff_A_ZqrpNP8R5_1),.clk(gclk));
	jdff dff_A_sukh36C02_1(.dout(w_dff_A_ZqrpNP8R5_1),.din(w_dff_A_sukh36C02_1),.clk(gclk));
	jdff dff_A_uCHG4j7O2_2(.dout(w_n80_0[2]),.din(w_dff_A_uCHG4j7O2_2),.clk(gclk));
	jdff dff_A_hrCraXZX3_2(.dout(w_dff_A_uCHG4j7O2_2),.din(w_dff_A_hrCraXZX3_2),.clk(gclk));
	jdff dff_A_D9v8rz468_2(.dout(w_dff_A_hrCraXZX3_2),.din(w_dff_A_D9v8rz468_2),.clk(gclk));
	jdff dff_A_pK4nazjv8_2(.dout(w_dff_A_D9v8rz468_2),.din(w_dff_A_pK4nazjv8_2),.clk(gclk));
	jdff dff_A_AUfBtQ1c5_0(.dout(w_n79_1[0]),.din(w_dff_A_AUfBtQ1c5_0),.clk(gclk));
	jdff dff_A_PPGohfHm8_0(.dout(w_dff_A_AUfBtQ1c5_0),.din(w_dff_A_PPGohfHm8_0),.clk(gclk));
	jdff dff_A_Ib35Ox4U7_0(.dout(w_dff_A_PPGohfHm8_0),.din(w_dff_A_Ib35Ox4U7_0),.clk(gclk));
	jdff dff_A_OFeyg3eT2_0(.dout(w_dff_A_Ib35Ox4U7_0),.din(w_dff_A_OFeyg3eT2_0),.clk(gclk));
	jdff dff_A_PRuOSv1q6_2(.dout(w_n79_1[2]),.din(w_dff_A_PRuOSv1q6_2),.clk(gclk));
	jdff dff_A_pJD95jjG5_1(.dout(w_n79_0[1]),.din(w_dff_A_pJD95jjG5_1),.clk(gclk));
	jdff dff_A_N68nDtWQ1_1(.dout(w_dff_A_pJD95jjG5_1),.din(w_dff_A_N68nDtWQ1_1),.clk(gclk));
	jdff dff_A_FMuI1CcA8_0(.dout(w_G87_3[0]),.din(w_dff_A_FMuI1CcA8_0),.clk(gclk));
	jdff dff_B_g2BUHUmX1_1(.din(n683),.dout(w_dff_B_g2BUHUmX1_1),.clk(gclk));
	jdff dff_B_AroFzrwl4_1(.din(w_dff_B_g2BUHUmX1_1),.dout(w_dff_B_AroFzrwl4_1),.clk(gclk));
	jdff dff_B_EOO2UkWM2_1(.din(w_dff_B_AroFzrwl4_1),.dout(w_dff_B_EOO2UkWM2_1),.clk(gclk));
	jdff dff_B_zs0to0HM6_1(.din(w_dff_B_EOO2UkWM2_1),.dout(w_dff_B_zs0to0HM6_1),.clk(gclk));
	jdff dff_A_JrF3vsGJ7_2(.dout(w_n75_0[2]),.din(w_dff_A_JrF3vsGJ7_2),.clk(gclk));
	jdff dff_A_Gul787wf1_2(.dout(w_dff_A_JrF3vsGJ7_2),.din(w_dff_A_Gul787wf1_2),.clk(gclk));
	jdff dff_A_N1DAoVzM8_2(.dout(w_dff_A_Gul787wf1_2),.din(w_dff_A_N1DAoVzM8_2),.clk(gclk));
	jdff dff_A_Evudwhde2_2(.dout(w_dff_A_N1DAoVzM8_2),.din(w_dff_A_Evudwhde2_2),.clk(gclk));
	jdff dff_A_KpwcKUwN2_2(.dout(w_n74_0[2]),.din(w_dff_A_KpwcKUwN2_2),.clk(gclk));
	jdff dff_A_gusQRcRR1_2(.dout(w_dff_A_KpwcKUwN2_2),.din(w_dff_A_gusQRcRR1_2),.clk(gclk));
	jdff dff_A_Pgt8R5mk2_2(.dout(w_dff_A_gusQRcRR1_2),.din(w_dff_A_Pgt8R5mk2_2),.clk(gclk));
	jdff dff_A_Q82G0qZs0_2(.dout(w_dff_A_Pgt8R5mk2_2),.din(w_dff_A_Q82G0qZs0_2),.clk(gclk));
	jdff dff_A_xSsMCRBr7_0(.dout(w_G33_6[0]),.din(w_dff_A_xSsMCRBr7_0),.clk(gclk));
	jdff dff_A_lW4jTWas2_0(.dout(w_dff_A_xSsMCRBr7_0),.din(w_dff_A_lW4jTWas2_0),.clk(gclk));
	jdff dff_A_3elhcIgK5_0(.dout(w_dff_A_lW4jTWas2_0),.din(w_dff_A_3elhcIgK5_0),.clk(gclk));
	jdff dff_A_Qz9JojIl6_0(.dout(w_dff_A_3elhcIgK5_0),.din(w_dff_A_Qz9JojIl6_0),.clk(gclk));
	jdff dff_A_FvVptbhJ6_0(.dout(w_dff_A_Qz9JojIl6_0),.din(w_dff_A_FvVptbhJ6_0),.clk(gclk));
	jdff dff_A_tvZyrkCr1_0(.dout(w_dff_A_FvVptbhJ6_0),.din(w_dff_A_tvZyrkCr1_0),.clk(gclk));
	jdff dff_A_SprqBrJ81_1(.dout(w_G33_6[1]),.din(w_dff_A_SprqBrJ81_1),.clk(gclk));
	jdff dff_A_jlWWod3j4_1(.dout(w_dff_A_SprqBrJ81_1),.din(w_dff_A_jlWWod3j4_1),.clk(gclk));
	jdff dff_A_4ED3xgM51_1(.dout(w_dff_A_jlWWod3j4_1),.din(w_dff_A_4ED3xgM51_1),.clk(gclk));
	jdff dff_A_iVZsRrpd7_0(.dout(w_G33_1[0]),.din(w_dff_A_iVZsRrpd7_0),.clk(gclk));
	jdff dff_A_2SGy3vXE7_0(.dout(w_dff_A_iVZsRrpd7_0),.din(w_dff_A_2SGy3vXE7_0),.clk(gclk));
	jdff dff_A_UfpkqPRw4_1(.dout(w_G33_1[1]),.din(w_dff_A_UfpkqPRw4_1),.clk(gclk));
	jdff dff_A_iCkZqIXJ7_1(.dout(w_dff_A_UfpkqPRw4_1),.din(w_dff_A_iCkZqIXJ7_1),.clk(gclk));
	jdff dff_A_IfmgPiJs5_1(.dout(w_n134_0[1]),.din(w_dff_A_IfmgPiJs5_1),.clk(gclk));
	jdff dff_A_66Lb5xL71_0(.dout(w_G77_4[0]),.din(w_dff_A_66Lb5xL71_0),.clk(gclk));
	jdff dff_A_kk3grUL39_1(.dout(w_G77_1[1]),.din(w_dff_A_kk3grUL39_1),.clk(gclk));
	jdff dff_A_DLOvlq2Y9_1(.dout(w_dff_A_kk3grUL39_1),.din(w_dff_A_DLOvlq2Y9_1),.clk(gclk));
	jdff dff_A_U3yMFeo12_1(.dout(w_dff_A_DLOvlq2Y9_1),.din(w_dff_A_U3yMFeo12_1),.clk(gclk));
	jdff dff_A_t101vT8I6_1(.dout(w_dff_A_U3yMFeo12_1),.din(w_dff_A_t101vT8I6_1),.clk(gclk));
	jdff dff_A_GYNZU5xm9_0(.dout(w_G68_5[0]),.din(w_dff_A_GYNZU5xm9_0),.clk(gclk));
	jdff dff_A_Z5goGDQd7_2(.dout(w_G68_1[2]),.din(w_dff_A_Z5goGDQd7_2),.clk(gclk));
	jdff dff_A_ywlBQ1Eu4_2(.dout(w_dff_A_Z5goGDQd7_2),.din(w_dff_A_ywlBQ1Eu4_2),.clk(gclk));
	jdff dff_A_atCkOc2f6_2(.dout(w_dff_A_ywlBQ1Eu4_2),.din(w_dff_A_atCkOc2f6_2),.clk(gclk));
	jdff dff_A_4T2OBKU75_0(.dout(w_G58_5[0]),.din(w_dff_A_4T2OBKU75_0),.clk(gclk));
	jdff dff_A_uevzUhaB9_1(.dout(w_G50_5[1]),.din(w_dff_A_uevzUhaB9_1),.clk(gclk));
	jdff dff_A_YHrPatvI4_1(.dout(w_dff_A_uevzUhaB9_1),.din(w_dff_A_YHrPatvI4_1),.clk(gclk));
	jdff dff_A_5FfXtKws4_1(.dout(w_dff_A_YHrPatvI4_1),.din(w_dff_A_5FfXtKws4_1),.clk(gclk));
	jdff dff_A_Ur4fGXuz7_0(.dout(w_n352_1[0]),.din(w_dff_A_Ur4fGXuz7_0),.clk(gclk));
	jdff dff_A_tvIXBdGs1_1(.dout(w_n352_0[1]),.din(w_dff_A_tvIXBdGs1_1),.clk(gclk));
	jdff dff_A_Om6iWjaW9_1(.dout(w_dff_A_tvIXBdGs1_1),.din(w_dff_A_Om6iWjaW9_1),.clk(gclk));
	jdff dff_A_skZTG5Uq4_1(.dout(w_dff_A_Om6iWjaW9_1),.din(w_dff_A_skZTG5Uq4_1),.clk(gclk));
	jdff dff_A_l5QVFNa52_1(.dout(w_dff_A_skZTG5Uq4_1),.din(w_dff_A_l5QVFNa52_1),.clk(gclk));
	jdff dff_A_3kGape6e9_2(.dout(w_n352_0[2]),.din(w_dff_A_3kGape6e9_2),.clk(gclk));
	jdff dff_A_Igq2p78F1_2(.dout(w_dff_A_3kGape6e9_2),.din(w_dff_A_Igq2p78F1_2),.clk(gclk));
	jdff dff_A_OVOzVEbJ0_2(.dout(w_dff_A_Igq2p78F1_2),.din(w_dff_A_OVOzVEbJ0_2),.clk(gclk));
	jdff dff_A_HR4uFf1G5_1(.dout(w_n682_0[1]),.din(w_dff_A_HR4uFf1G5_1),.clk(gclk));
	jdff dff_A_jvgRanVX8_1(.dout(w_dff_A_HR4uFf1G5_1),.din(w_dff_A_jvgRanVX8_1),.clk(gclk));
	jdff dff_A_W5TRT1jw1_1(.dout(w_dff_A_jvgRanVX8_1),.din(w_dff_A_W5TRT1jw1_1),.clk(gclk));
	jdff dff_A_sHAus9Hg6_1(.dout(w_dff_A_W5TRT1jw1_1),.din(w_dff_A_sHAus9Hg6_1),.clk(gclk));
	jdff dff_A_6lkBff8a2_1(.dout(w_n680_4[1]),.din(w_dff_A_6lkBff8a2_1),.clk(gclk));
	jdff dff_A_r3xTgCrX5_1(.dout(w_dff_A_6lkBff8a2_1),.din(w_dff_A_r3xTgCrX5_1),.clk(gclk));
	jdff dff_A_cHLg8j5i1_1(.dout(w_dff_A_r3xTgCrX5_1),.din(w_dff_A_cHLg8j5i1_1),.clk(gclk));
	jdff dff_A_KxzTbend0_1(.dout(w_dff_A_cHLg8j5i1_1),.din(w_dff_A_KxzTbend0_1),.clk(gclk));
	jdff dff_A_L1OUvBOX5_1(.dout(w_dff_A_KxzTbend0_1),.din(w_dff_A_L1OUvBOX5_1),.clk(gclk));
	jdff dff_A_gLdsm9MT0_1(.dout(w_dff_A_L1OUvBOX5_1),.din(w_dff_A_gLdsm9MT0_1),.clk(gclk));
	jdff dff_A_vOdaRpIR9_1(.dout(w_dff_A_gLdsm9MT0_1),.din(w_dff_A_vOdaRpIR9_1),.clk(gclk));
	jdff dff_A_wVzkdJBF7_1(.dout(w_dff_A_vOdaRpIR9_1),.din(w_dff_A_wVzkdJBF7_1),.clk(gclk));
	jdff dff_A_WB1iM4RD7_1(.dout(w_n680_1[1]),.din(w_dff_A_WB1iM4RD7_1),.clk(gclk));
	jdff dff_A_HlhaDl444_1(.dout(w_dff_A_WB1iM4RD7_1),.din(w_dff_A_HlhaDl444_1),.clk(gclk));
	jdff dff_A_bUjDrnwq9_1(.dout(w_dff_A_HlhaDl444_1),.din(w_dff_A_bUjDrnwq9_1),.clk(gclk));
	jdff dff_A_Uld5ZWv42_1(.dout(w_dff_A_bUjDrnwq9_1),.din(w_dff_A_Uld5ZWv42_1),.clk(gclk));
	jdff dff_A_pB17JVLV8_1(.dout(w_dff_A_Uld5ZWv42_1),.din(w_dff_A_pB17JVLV8_1),.clk(gclk));
	jdff dff_A_RYyAyxtK4_1(.dout(w_dff_A_pB17JVLV8_1),.din(w_dff_A_RYyAyxtK4_1),.clk(gclk));
	jdff dff_A_AieAZqdi9_1(.dout(w_dff_A_RYyAyxtK4_1),.din(w_dff_A_AieAZqdi9_1),.clk(gclk));
	jdff dff_A_3UeoD8xh0_1(.dout(w_n680_0[1]),.din(w_dff_A_3UeoD8xh0_1),.clk(gclk));
	jdff dff_A_mJel1wGl0_1(.dout(w_dff_A_3UeoD8xh0_1),.din(w_dff_A_mJel1wGl0_1),.clk(gclk));
	jdff dff_A_iTbNsJcu3_1(.dout(w_dff_A_mJel1wGl0_1),.din(w_dff_A_iTbNsJcu3_1),.clk(gclk));
	jdff dff_A_VLgwlKXU5_1(.dout(w_dff_A_iTbNsJcu3_1),.din(w_dff_A_VLgwlKXU5_1),.clk(gclk));
	jdff dff_A_sQCRFlbg1_1(.dout(w_dff_A_VLgwlKXU5_1),.din(w_dff_A_sQCRFlbg1_1),.clk(gclk));
	jdff dff_A_pilupIAD1_1(.dout(w_G169_1[1]),.din(w_dff_A_pilupIAD1_1),.clk(gclk));
	jdff dff_A_LlXQbDvJ1_1(.dout(w_dff_A_pilupIAD1_1),.din(w_dff_A_LlXQbDvJ1_1),.clk(gclk));
	jdff dff_A_3QuVspq13_1(.dout(w_dff_A_LlXQbDvJ1_1),.din(w_dff_A_3QuVspq13_1),.clk(gclk));
	jdff dff_A_qabvBadO0_1(.dout(w_dff_A_3QuVspq13_1),.din(w_dff_A_qabvBadO0_1),.clk(gclk));
	jdff dff_A_vBIy6OKn2_1(.dout(w_dff_A_qabvBadO0_1),.din(w_dff_A_vBIy6OKn2_1),.clk(gclk));
	jdff dff_A_Zq0Bc14H4_1(.dout(w_dff_A_vBIy6OKn2_1),.din(w_dff_A_Zq0Bc14H4_1),.clk(gclk));
	jdff dff_A_S1Gy7Grj3_2(.dout(w_G169_1[2]),.din(w_dff_A_S1Gy7Grj3_2),.clk(gclk));
	jdff dff_A_oXYJQoHw7_2(.dout(w_dff_A_S1Gy7Grj3_2),.din(w_dff_A_oXYJQoHw7_2),.clk(gclk));
	jdff dff_A_PVds1BQh4_2(.dout(w_dff_A_oXYJQoHw7_2),.din(w_dff_A_PVds1BQh4_2),.clk(gclk));
	jdff dff_A_VG8jbie57_2(.dout(w_dff_A_PVds1BQh4_2),.din(w_dff_A_VG8jbie57_2),.clk(gclk));
	jdff dff_A_Eibqprn34_2(.dout(w_dff_A_VG8jbie57_2),.din(w_dff_A_Eibqprn34_2),.clk(gclk));
	jdff dff_A_abaKJPaS9_2(.dout(w_dff_A_Eibqprn34_2),.din(w_dff_A_abaKJPaS9_2),.clk(gclk));
	jdff dff_A_huDPOu0W6_2(.dout(w_dff_A_abaKJPaS9_2),.din(w_dff_A_huDPOu0W6_2),.clk(gclk));
	jdff dff_A_n08iQj1A2_2(.dout(w_dff_A_huDPOu0W6_2),.din(w_dff_A_n08iQj1A2_2),.clk(gclk));
	jdff dff_A_NOo5No7a1_1(.dout(w_n151_4[1]),.din(w_dff_A_NOo5No7a1_1),.clk(gclk));
	jdff dff_A_ja4D9moc2_1(.dout(w_dff_A_NOo5No7a1_1),.din(w_dff_A_ja4D9moc2_1),.clk(gclk));
	jdff dff_A_4MwNiXOn4_1(.dout(w_dff_A_ja4D9moc2_1),.din(w_dff_A_4MwNiXOn4_1),.clk(gclk));
	jdff dff_B_epnIwufb4_0(.din(n676),.dout(w_dff_B_epnIwufb4_0),.clk(gclk));
	jdff dff_B_IPXw9dON6_0(.din(w_dff_B_epnIwufb4_0),.dout(w_dff_B_IPXw9dON6_0),.clk(gclk));
	jdff dff_B_zQEgkBVr2_1(.din(n661),.dout(w_dff_B_zQEgkBVr2_1),.clk(gclk));
	jdff dff_B_SI3vpvEF0_1(.din(w_dff_B_zQEgkBVr2_1),.dout(w_dff_B_SI3vpvEF0_1),.clk(gclk));
	jdff dff_B_duIrmeBB7_1(.din(w_dff_B_SI3vpvEF0_1),.dout(w_dff_B_duIrmeBB7_1),.clk(gclk));
	jdff dff_B_2WX1sdRp1_1(.din(w_dff_B_duIrmeBB7_1),.dout(w_dff_B_2WX1sdRp1_1),.clk(gclk));
	jdff dff_B_PGB7mGTc7_0(.din(n672),.dout(w_dff_B_PGB7mGTc7_0),.clk(gclk));
	jdff dff_A_wFVyREYN6_0(.dout(w_G317_1[0]),.din(w_dff_A_wFVyREYN6_0),.clk(gclk));
	jdff dff_B_15zbGLLk8_3(.din(G317),.dout(w_dff_B_15zbGLLk8_3),.clk(gclk));
	jdff dff_B_PFBmPIhI2_3(.din(w_dff_B_15zbGLLk8_3),.dout(w_dff_B_PFBmPIhI2_3),.clk(gclk));
	jdff dff_B_aZT4eAIR2_3(.din(w_dff_B_PFBmPIhI2_3),.dout(w_dff_B_aZT4eAIR2_3),.clk(gclk));
	jdff dff_A_FduAQ6k65_1(.dout(w_G311_1[1]),.din(w_dff_A_FduAQ6k65_1),.clk(gclk));
	jdff dff_B_YFWQiIGl2_3(.din(G311),.dout(w_dff_B_YFWQiIGl2_3),.clk(gclk));
	jdff dff_B_b8tum4Cb1_3(.din(w_dff_B_YFWQiIGl2_3),.dout(w_dff_B_b8tum4Cb1_3),.clk(gclk));
	jdff dff_B_DleL7hkB5_3(.din(w_dff_B_b8tum4Cb1_3),.dout(w_dff_B_DleL7hkB5_3),.clk(gclk));
	jdff dff_B_Qoi6h4hS8_1(.din(G329),.dout(w_dff_B_Qoi6h4hS8_1),.clk(gclk));
	jdff dff_B_MkNT7zZD7_1(.din(w_dff_B_Qoi6h4hS8_1),.dout(w_dff_B_MkNT7zZD7_1),.clk(gclk));
	jdff dff_B_hpPNEX8y4_1(.din(w_dff_B_MkNT7zZD7_1),.dout(w_dff_B_hpPNEX8y4_1),.clk(gclk));
	jdff dff_B_U5SKTSDO0_1(.din(w_dff_B_hpPNEX8y4_1),.dout(w_dff_B_U5SKTSDO0_1),.clk(gclk));
	jdff dff_B_s0siIhop1_0(.din(n665),.dout(w_dff_B_s0siIhop1_0),.clk(gclk));
	jdff dff_B_Xa6NuVoZ9_0(.din(w_dff_B_s0siIhop1_0),.dout(w_dff_B_Xa6NuVoZ9_0),.clk(gclk));
	jdff dff_A_UAHBuC8a9_0(.dout(w_G326_0[0]),.din(w_dff_A_UAHBuC8a9_0),.clk(gclk));
	jdff dff_B_ctEQa78R7_2(.din(G326),.dout(w_dff_B_ctEQa78R7_2),.clk(gclk));
	jdff dff_B_uWuWFUxP0_2(.din(w_dff_B_ctEQa78R7_2),.dout(w_dff_B_uWuWFUxP0_2),.clk(gclk));
	jdff dff_B_3IYLQbVv5_2(.din(w_dff_B_uWuWFUxP0_2),.dout(w_dff_B_3IYLQbVv5_2),.clk(gclk));
	jdff dff_B_MdHqP3XU9_1(.din(n662),.dout(w_dff_B_MdHqP3XU9_1),.clk(gclk));
	jdff dff_A_RvwD4hSX8_0(.dout(w_G294_3[0]),.din(w_dff_A_RvwD4hSX8_0),.clk(gclk));
	jdff dff_A_HFE3nYvt1_0(.dout(w_dff_A_RvwD4hSX8_0),.din(w_dff_A_HFE3nYvt1_0),.clk(gclk));
	jdff dff_A_InUxnsUw6_0(.dout(w_dff_A_HFE3nYvt1_0),.din(w_dff_A_InUxnsUw6_0),.clk(gclk));
	jdff dff_A_7KXAvexG1_0(.dout(w_dff_A_InUxnsUw6_0),.din(w_dff_A_7KXAvexG1_0),.clk(gclk));
	jdff dff_A_nCtp9fmY5_0(.dout(w_G294_0[0]),.din(w_dff_A_nCtp9fmY5_0),.clk(gclk));
	jdff dff_A_imFC1NFv1_0(.dout(w_dff_A_nCtp9fmY5_0),.din(w_dff_A_imFC1NFv1_0),.clk(gclk));
	jdff dff_A_M8PDc24u2_0(.dout(w_dff_A_imFC1NFv1_0),.din(w_dff_A_M8PDc24u2_0),.clk(gclk));
	jdff dff_A_dfPF7vOD9_1(.dout(w_G294_0[1]),.din(w_dff_A_dfPF7vOD9_1),.clk(gclk));
	jdff dff_A_XA49QrCj3_1(.dout(w_dff_A_dfPF7vOD9_1),.din(w_dff_A_XA49QrCj3_1),.clk(gclk));
	jdff dff_A_UGB6UDPz6_1(.dout(w_dff_A_XA49QrCj3_1),.din(w_dff_A_UGB6UDPz6_1),.clk(gclk));
	jdff dff_A_IgwH6UHi3_0(.dout(w_G322_0[0]),.din(w_dff_A_IgwH6UHi3_0),.clk(gclk));
	jdff dff_B_nT9B3m7w1_3(.din(G322),.dout(w_dff_B_nT9B3m7w1_3),.clk(gclk));
	jdff dff_B_DuNi19WN8_3(.din(w_dff_B_nT9B3m7w1_3),.dout(w_dff_B_DuNi19WN8_3),.clk(gclk));
	jdff dff_B_76RyYuVJ5_3(.din(w_dff_B_DuNi19WN8_3),.dout(w_dff_B_76RyYuVJ5_3),.clk(gclk));
	jdff dff_B_XZYEa8my8_0(.din(n658),.dout(w_dff_B_XZYEa8my8_0),.clk(gclk));
	jdff dff_B_ZpGwgD9l5_1(.din(n647),.dout(w_dff_B_ZpGwgD9l5_1),.clk(gclk));
	jdff dff_B_WwaOHHlo8_1(.din(w_dff_B_ZpGwgD9l5_1),.dout(w_dff_B_WwaOHHlo8_1),.clk(gclk));
	jdff dff_A_Rpv7GXwZ4_1(.dout(w_G68_3[1]),.din(w_dff_A_Rpv7GXwZ4_1),.clk(gclk));
	jdff dff_A_gkhyvNus0_1(.dout(w_dff_A_Rpv7GXwZ4_1),.din(w_dff_A_gkhyvNus0_1),.clk(gclk));
	jdff dff_A_99bYBXMd5_2(.dout(w_G68_3[2]),.din(w_dff_A_99bYBXMd5_2),.clk(gclk));
	jdff dff_A_YbKn54312_2(.dout(w_dff_A_99bYBXMd5_2),.din(w_dff_A_YbKn54312_2),.clk(gclk));
	jdff dff_A_hIy1Evbj3_2(.dout(w_G68_0[2]),.din(w_dff_A_hIy1Evbj3_2),.clk(gclk));
	jdff dff_A_Lvr95I756_0(.dout(w_G50_4[0]),.din(w_dff_A_Lvr95I756_0),.clk(gclk));
	jdff dff_A_myzgEm6o4_0(.dout(w_dff_A_Lvr95I756_0),.din(w_dff_A_myzgEm6o4_0),.clk(gclk));
	jdff dff_A_bPu9byLN0_1(.dout(w_G50_4[1]),.din(w_dff_A_bPu9byLN0_1),.clk(gclk));
	jdff dff_A_IatAuJ4D8_1(.dout(w_dff_A_bPu9byLN0_1),.din(w_dff_A_IatAuJ4D8_1),.clk(gclk));
	jdff dff_A_uRXQAEmO4_0(.dout(w_G50_1[0]),.din(w_dff_A_uRXQAEmO4_0),.clk(gclk));
	jdff dff_A_TYmLuvgm0_2(.dout(w_G50_1[2]),.din(w_dff_A_TYmLuvgm0_2),.clk(gclk));
	jdff dff_A_iPQOF0Vq4_2(.dout(w_dff_A_TYmLuvgm0_2),.din(w_dff_A_iPQOF0Vq4_2),.clk(gclk));
	jdff dff_A_PLpIwZTf2_2(.dout(w_dff_A_iPQOF0Vq4_2),.din(w_dff_A_PLpIwZTf2_2),.clk(gclk));
	jdff dff_A_TfYO4oLX8_2(.dout(w_dff_A_PLpIwZTf2_2),.din(w_dff_A_TfYO4oLX8_2),.clk(gclk));
	jdff dff_A_BaM0tXbx0_1(.dout(w_n649_0[1]),.din(w_dff_A_BaM0tXbx0_1),.clk(gclk));
	jdff dff_A_rwpDjkM27_0(.dout(w_G107_3[0]),.din(w_dff_A_rwpDjkM27_0),.clk(gclk));
	jdff dff_A_u7tOXK7N1_0(.dout(w_dff_A_rwpDjkM27_0),.din(w_dff_A_u7tOXK7N1_0),.clk(gclk));
	jdff dff_A_1053Xzse9_0(.dout(w_dff_A_u7tOXK7N1_0),.din(w_dff_A_1053Xzse9_0),.clk(gclk));
	jdff dff_A_PSu8SQtN0_1(.dout(w_G107_0[1]),.din(w_dff_A_PSu8SQtN0_1),.clk(gclk));
	jdff dff_A_mLeTIMsk2_1(.dout(w_dff_A_PSu8SQtN0_1),.din(w_dff_A_mLeTIMsk2_1),.clk(gclk));
	jdff dff_A_JOflgydm7_1(.dout(w_dff_A_mLeTIMsk2_1),.din(w_dff_A_JOflgydm7_1),.clk(gclk));
	jdff dff_A_lbRvUuZh2_0(.dout(w_G58_4[0]),.din(w_dff_A_lbRvUuZh2_0),.clk(gclk));
	jdff dff_A_GjeJFaG75_0(.dout(w_dff_A_lbRvUuZh2_0),.din(w_dff_A_GjeJFaG75_0),.clk(gclk));
	jdff dff_A_JDcLtCSU8_0(.dout(w_dff_A_GjeJFaG75_0),.din(w_dff_A_JDcLtCSU8_0),.clk(gclk));
	jdff dff_A_jcmTerpl0_2(.dout(w_G58_4[2]),.din(w_dff_A_jcmTerpl0_2),.clk(gclk));
	jdff dff_A_ga0eICyE4_2(.dout(w_dff_A_jcmTerpl0_2),.din(w_dff_A_ga0eICyE4_2),.clk(gclk));
	jdff dff_A_S2EvNYYq9_2(.dout(w_G58_1[2]),.din(w_dff_A_S2EvNYYq9_2),.clk(gclk));
	jdff dff_A_a8oYTciW2_2(.dout(w_dff_A_S2EvNYYq9_2),.din(w_dff_A_a8oYTciW2_2),.clk(gclk));
	jdff dff_A_oDEU0Bbw2_2(.dout(w_dff_A_a8oYTciW2_2),.din(w_dff_A_oDEU0Bbw2_2),.clk(gclk));
	jdff dff_A_ID44LOwM4_1(.dout(w_G58_0[1]),.din(w_dff_A_ID44LOwM4_1),.clk(gclk));
	jdff dff_B_cx0kmtJb8_1(.din(n636),.dout(w_dff_B_cx0kmtJb8_1),.clk(gclk));
	jdff dff_B_cTi4cvda5_1(.din(n639),.dout(w_dff_B_cTi4cvda5_1),.clk(gclk));
	jdff dff_A_Ud0i2WQE0_0(.dout(w_G159_3[0]),.din(w_dff_A_Ud0i2WQE0_0),.clk(gclk));
	jdff dff_A_LySYsfzo0_0(.dout(w_dff_A_Ud0i2WQE0_0),.din(w_dff_A_LySYsfzo0_0),.clk(gclk));
	jdff dff_A_uCHVmEAR2_0(.dout(w_dff_A_LySYsfzo0_0),.din(w_dff_A_uCHVmEAR2_0),.clk(gclk));
	jdff dff_A_RRvMJjBr1_1(.dout(w_G159_3[1]),.din(w_dff_A_RRvMJjBr1_1),.clk(gclk));
	jdff dff_A_easMpTaD7_1(.dout(w_dff_A_RRvMJjBr1_1),.din(w_dff_A_easMpTaD7_1),.clk(gclk));
	jdff dff_A_wBMgzwlS3_1(.dout(w_dff_A_easMpTaD7_1),.din(w_dff_A_wBMgzwlS3_1),.clk(gclk));
	jdff dff_A_OjRpaYTH3_1(.dout(w_dff_A_wBMgzwlS3_1),.din(w_dff_A_OjRpaYTH3_1),.clk(gclk));
	jdff dff_A_jPZB0Uh39_0(.dout(w_G159_0[0]),.din(w_dff_A_jPZB0Uh39_0),.clk(gclk));
	jdff dff_A_fgpOljVt1_0(.dout(w_dff_A_jPZB0Uh39_0),.din(w_dff_A_fgpOljVt1_0),.clk(gclk));
	jdff dff_A_gTmJHqmw8_0(.dout(w_dff_A_fgpOljVt1_0),.din(w_dff_A_gTmJHqmw8_0),.clk(gclk));
	jdff dff_A_BoUr2vNR5_1(.dout(w_G159_0[1]),.din(w_dff_A_BoUr2vNR5_1),.clk(gclk));
	jdff dff_A_7aLUCqxE7_1(.dout(w_dff_A_BoUr2vNR5_1),.din(w_dff_A_7aLUCqxE7_1),.clk(gclk));
	jdff dff_A_02gL5xdu7_1(.dout(w_dff_A_7aLUCqxE7_1),.din(w_dff_A_02gL5xdu7_1),.clk(gclk));
	jdff dff_A_FNTuUT801_0(.dout(w_n388_0[0]),.din(w_dff_A_FNTuUT801_0),.clk(gclk));
	jdff dff_A_HTBDeNDf9_0(.dout(w_dff_A_FNTuUT801_0),.din(w_dff_A_HTBDeNDf9_0),.clk(gclk));
	jdff dff_A_VJu7bfcK9_0(.dout(w_dff_A_HTBDeNDf9_0),.din(w_dff_A_VJu7bfcK9_0),.clk(gclk));
	jdff dff_A_rJbWsbZI0_0(.dout(w_dff_A_VJu7bfcK9_0),.din(w_dff_A_rJbWsbZI0_0),.clk(gclk));
	jdff dff_A_dhPSkfWg5_0(.dout(w_dff_A_rJbWsbZI0_0),.din(w_dff_A_dhPSkfWg5_0),.clk(gclk));
	jdff dff_A_hvqDGvPG2_0(.dout(w_dff_A_dhPSkfWg5_0),.din(w_dff_A_hvqDGvPG2_0),.clk(gclk));
	jdff dff_A_0DNBLfcy6_1(.dout(w_n388_0[1]),.din(w_dff_A_0DNBLfcy6_1),.clk(gclk));
	jdff dff_A_roSSWwob9_1(.dout(w_dff_A_0DNBLfcy6_1),.din(w_dff_A_roSSWwob9_1),.clk(gclk));
	jdff dff_A_Gn1Ngk807_1(.dout(w_dff_A_roSSWwob9_1),.din(w_dff_A_Gn1Ngk807_1),.clk(gclk));
	jdff dff_A_wRJmGnUW9_1(.dout(w_dff_A_Gn1Ngk807_1),.din(w_dff_A_wRJmGnUW9_1),.clk(gclk));
	jdff dff_A_nEejx1Yk7_1(.dout(w_dff_A_wRJmGnUW9_1),.din(w_dff_A_nEejx1Yk7_1),.clk(gclk));
	jdff dff_A_eFTL9DI97_1(.dout(w_dff_A_nEejx1Yk7_1),.din(w_dff_A_eFTL9DI97_1),.clk(gclk));
	jdff dff_A_5ZUteJJl5_1(.dout(w_dff_A_eFTL9DI97_1),.din(w_dff_A_5ZUteJJl5_1),.clk(gclk));
	jdff dff_A_OVgrBv1T6_1(.dout(w_G200_2[1]),.din(w_dff_A_OVgrBv1T6_1),.clk(gclk));
	jdff dff_A_CtOhJ50s6_1(.dout(w_dff_A_OVgrBv1T6_1),.din(w_dff_A_CtOhJ50s6_1),.clk(gclk));
	jdff dff_A_NnTjfPfF4_1(.dout(w_dff_A_CtOhJ50s6_1),.din(w_dff_A_NnTjfPfF4_1),.clk(gclk));
	jdff dff_A_Z8NYjraw5_1(.dout(w_dff_A_NnTjfPfF4_1),.din(w_dff_A_Z8NYjraw5_1),.clk(gclk));
	jdff dff_A_VaIGOAew9_1(.dout(w_dff_A_Z8NYjraw5_1),.din(w_dff_A_VaIGOAew9_1),.clk(gclk));
	jdff dff_A_cNXzxi6f5_1(.dout(w_dff_A_VaIGOAew9_1),.din(w_dff_A_cNXzxi6f5_1),.clk(gclk));
	jdff dff_A_9LhzQicR2_1(.dout(w_dff_A_cNXzxi6f5_1),.din(w_dff_A_9LhzQicR2_1),.clk(gclk));
	jdff dff_A_JVEiqZj74_1(.dout(w_dff_A_9LhzQicR2_1),.din(w_dff_A_JVEiqZj74_1),.clk(gclk));
	jdff dff_A_juqI9PiX2_2(.dout(w_G200_2[2]),.din(w_dff_A_juqI9PiX2_2),.clk(gclk));
	jdff dff_A_dv0y0SBw3_2(.dout(w_dff_A_juqI9PiX2_2),.din(w_dff_A_dv0y0SBw3_2),.clk(gclk));
	jdff dff_A_uf482u1O4_2(.dout(w_dff_A_dv0y0SBw3_2),.din(w_dff_A_uf482u1O4_2),.clk(gclk));
	jdff dff_A_ZGUTahiJ3_2(.dout(w_dff_A_uf482u1O4_2),.din(w_dff_A_ZGUTahiJ3_2),.clk(gclk));
	jdff dff_A_9gTQKhFJ3_2(.dout(w_dff_A_ZGUTahiJ3_2),.din(w_dff_A_9gTQKhFJ3_2),.clk(gclk));
	jdff dff_A_ddD7f9Uq0_2(.dout(w_dff_A_9gTQKhFJ3_2),.din(w_dff_A_ddD7f9Uq0_2),.clk(gclk));
	jdff dff_A_RuwTxlmp4_2(.dout(w_dff_A_ddD7f9Uq0_2),.din(w_dff_A_RuwTxlmp4_2),.clk(gclk));
	jdff dff_A_7bb0sUTJ1_0(.dout(w_G77_3[0]),.din(w_dff_A_7bb0sUTJ1_0),.clk(gclk));
	jdff dff_A_50Fg1vgp4_0(.dout(w_dff_A_7bb0sUTJ1_0),.din(w_dff_A_50Fg1vgp4_0),.clk(gclk));
	jdff dff_A_RnLehcsx9_0(.dout(w_dff_A_50Fg1vgp4_0),.din(w_dff_A_RnLehcsx9_0),.clk(gclk));
	jdff dff_A_i9CGDgPG3_2(.dout(w_G77_3[2]),.din(w_dff_A_i9CGDgPG3_2),.clk(gclk));
	jdff dff_A_MlJChBlm4_2(.dout(w_dff_A_i9CGDgPG3_2),.din(w_dff_A_MlJChBlm4_2),.clk(gclk));
	jdff dff_A_6R5e6Vpw8_2(.dout(w_dff_A_MlJChBlm4_2),.din(w_dff_A_6R5e6Vpw8_2),.clk(gclk));
	jdff dff_A_H00ab9SS9_1(.dout(w_G77_0[1]),.din(w_dff_A_H00ab9SS9_1),.clk(gclk));
	jdff dff_A_TlHlMIDS6_1(.dout(w_dff_A_H00ab9SS9_1),.din(w_dff_A_TlHlMIDS6_1),.clk(gclk));
	jdff dff_A_WHNRDtKO3_0(.dout(w_G33_7[0]),.din(w_dff_A_WHNRDtKO3_0),.clk(gclk));
	jdff dff_A_QzjSqOyr6_0(.dout(w_dff_A_WHNRDtKO3_0),.din(w_dff_A_QzjSqOyr6_0),.clk(gclk));
	jdff dff_A_iZdiPAK29_0(.dout(w_dff_A_QzjSqOyr6_0),.din(w_dff_A_iZdiPAK29_0),.clk(gclk));
	jdff dff_A_i9Y28Gpo5_0(.dout(w_dff_A_iZdiPAK29_0),.din(w_dff_A_i9Y28Gpo5_0),.clk(gclk));
	jdff dff_A_eH5pr1Dt4_0(.dout(w_dff_A_i9Y28Gpo5_0),.din(w_dff_A_eH5pr1Dt4_0),.clk(gclk));
	jdff dff_A_KAokJYo86_0(.dout(w_dff_A_eH5pr1Dt4_0),.din(w_dff_A_KAokJYo86_0),.clk(gclk));
	jdff dff_A_awdv05eE1_1(.dout(w_G33_7[1]),.din(w_dff_A_awdv05eE1_1),.clk(gclk));
	jdff dff_B_HSexzlMl6_0(.din(n635),.dout(w_dff_B_HSexzlMl6_0),.clk(gclk));
	jdff dff_A_f6htjZ0h2_0(.dout(w_G87_2[0]),.din(w_dff_A_f6htjZ0h2_0),.clk(gclk));
	jdff dff_A_ctYTbV0I7_0(.dout(w_dff_A_f6htjZ0h2_0),.din(w_dff_A_ctYTbV0I7_0),.clk(gclk));
	jdff dff_A_lb8DHTMQ0_0(.dout(w_dff_A_ctYTbV0I7_0),.din(w_dff_A_lb8DHTMQ0_0),.clk(gclk));
	jdff dff_A_2w6f3LV65_1(.dout(w_G87_2[1]),.din(w_dff_A_2w6f3LV65_1),.clk(gclk));
	jdff dff_A_8vQCB9x34_1(.dout(w_dff_A_2w6f3LV65_1),.din(w_dff_A_8vQCB9x34_1),.clk(gclk));
	jdff dff_A_sCFfnYDW2_1(.dout(w_dff_A_8vQCB9x34_1),.din(w_dff_A_sCFfnYDW2_1),.clk(gclk));
	jdff dff_A_1cN0h2PT2_0(.dout(w_G87_0[0]),.din(w_dff_A_1cN0h2PT2_0),.clk(gclk));
	jdff dff_A_gV5tDO9v0_0(.dout(w_dff_A_1cN0h2PT2_0),.din(w_dff_A_gV5tDO9v0_0),.clk(gclk));
	jdff dff_A_tP0ttjuI6_0(.dout(w_dff_A_gV5tDO9v0_0),.din(w_dff_A_tP0ttjuI6_0),.clk(gclk));
	jdff dff_A_WuJdh9tN4_0(.dout(w_G200_1[0]),.din(w_dff_A_WuJdh9tN4_0),.clk(gclk));
	jdff dff_A_2SLOiQmU2_2(.dout(w_G200_1[2]),.din(w_dff_A_2SLOiQmU2_2),.clk(gclk));
	jdff dff_A_JTPDVDkf9_2(.dout(w_dff_A_2SLOiQmU2_2),.din(w_dff_A_JTPDVDkf9_2),.clk(gclk));
	jdff dff_A_5qPkdKiB1_2(.dout(w_dff_A_JTPDVDkf9_2),.din(w_dff_A_5qPkdKiB1_2),.clk(gclk));
	jdff dff_A_oMVEQn4J3_2(.dout(w_dff_A_5qPkdKiB1_2),.din(w_dff_A_oMVEQn4J3_2),.clk(gclk));
	jdff dff_A_naVGPcSL9_2(.dout(w_dff_A_oMVEQn4J3_2),.din(w_dff_A_naVGPcSL9_2),.clk(gclk));
	jdff dff_A_jcyD8gAL9_2(.dout(w_dff_A_naVGPcSL9_2),.din(w_dff_A_jcyD8gAL9_2),.clk(gclk));
	jdff dff_A_tyIazhTB1_2(.dout(w_dff_A_jcyD8gAL9_2),.din(w_dff_A_tyIazhTB1_2),.clk(gclk));
	jdff dff_A_qJJ0psJq6_2(.dout(w_dff_A_tyIazhTB1_2),.din(w_dff_A_qJJ0psJq6_2),.clk(gclk));
	jdff dff_A_LNnhatrx2_0(.dout(w_n622_0[0]),.din(w_dff_A_LNnhatrx2_0),.clk(gclk));
	jdff dff_A_EdOHaFaB2_0(.dout(w_n507_1[0]),.din(w_dff_A_EdOHaFaB2_0),.clk(gclk));
	jdff dff_A_HegGS2qX4_1(.dout(w_n507_1[1]),.din(w_dff_A_HegGS2qX4_1),.clk(gclk));
	jdff dff_A_aJvojiDY3_1(.dout(w_n507_0[1]),.din(w_dff_A_aJvojiDY3_1),.clk(gclk));
	jdff dff_A_NSxwuF543_1(.dout(w_dff_A_aJvojiDY3_1),.din(w_dff_A_NSxwuF543_1),.clk(gclk));
	jdff dff_A_EgUzCAux4_1(.dout(w_dff_A_NSxwuF543_1),.din(w_dff_A_EgUzCAux4_1),.clk(gclk));
	jdff dff_A_UZiJZi3v3_1(.dout(w_dff_A_EgUzCAux4_1),.din(w_dff_A_UZiJZi3v3_1),.clk(gclk));
	jdff dff_A_yLXqfWQo9_1(.dout(w_dff_A_UZiJZi3v3_1),.din(w_dff_A_yLXqfWQo9_1),.clk(gclk));
	jdff dff_A_qdkzIen67_1(.dout(w_dff_A_yLXqfWQo9_1),.din(w_dff_A_qdkzIen67_1),.clk(gclk));
	jdff dff_A_kt9eReKY6_2(.dout(w_n507_0[2]),.din(w_dff_A_kt9eReKY6_2),.clk(gclk));
	jdff dff_A_U5zeaEBP4_0(.dout(w_G190_2[0]),.din(w_dff_A_U5zeaEBP4_0),.clk(gclk));
	jdff dff_A_mj3y81XF0_0(.dout(w_dff_A_U5zeaEBP4_0),.din(w_dff_A_mj3y81XF0_0),.clk(gclk));
	jdff dff_A_CirbFGOI2_2(.dout(w_G190_2[2]),.din(w_dff_A_CirbFGOI2_2),.clk(gclk));
	jdff dff_A_G1XrAQAe4_2(.dout(w_dff_A_CirbFGOI2_2),.din(w_dff_A_G1XrAQAe4_2),.clk(gclk));
	jdff dff_A_kwMSiL5q6_2(.dout(w_dff_A_G1XrAQAe4_2),.din(w_dff_A_kwMSiL5q6_2),.clk(gclk));
	jdff dff_A_VbPXRntC0_2(.dout(w_dff_A_kwMSiL5q6_2),.din(w_dff_A_VbPXRntC0_2),.clk(gclk));
	jdff dff_A_QiMpmbzV4_2(.dout(w_dff_A_VbPXRntC0_2),.din(w_dff_A_QiMpmbzV4_2),.clk(gclk));
	jdff dff_A_ggKQXFRs6_2(.dout(w_dff_A_QiMpmbzV4_2),.din(w_dff_A_ggKQXFRs6_2),.clk(gclk));
	jdff dff_A_wOdYPzuO0_2(.dout(w_dff_A_ggKQXFRs6_2),.din(w_dff_A_wOdYPzuO0_2),.clk(gclk));
	jdff dff_A_exnGLAXE9_2(.dout(w_dff_A_wOdYPzuO0_2),.din(w_dff_A_exnGLAXE9_2),.clk(gclk));
	jdff dff_A_Za5J4EeW1_2(.dout(w_G20_2[2]),.din(w_dff_A_Za5J4EeW1_2),.clk(gclk));
	jdff dff_A_uAnlLjrn6_0(.dout(w_G97_3[0]),.din(w_dff_A_uAnlLjrn6_0),.clk(gclk));
	jdff dff_A_uhWG3V3B0_0(.dout(w_dff_A_uAnlLjrn6_0),.din(w_dff_A_uhWG3V3B0_0),.clk(gclk));
	jdff dff_A_bKjz2g4f0_0(.dout(w_dff_A_uhWG3V3B0_0),.din(w_dff_A_bKjz2g4f0_0),.clk(gclk));
	jdff dff_A_P9BlaCSh4_0(.dout(w_dff_A_bKjz2g4f0_0),.din(w_dff_A_P9BlaCSh4_0),.clk(gclk));
	jdff dff_A_SdTEQVUl4_0(.dout(w_n620_0[0]),.din(w_dff_A_SdTEQVUl4_0),.clk(gclk));
	jdff dff_A_EuxU2Int0_0(.dout(w_dff_A_SdTEQVUl4_0),.din(w_dff_A_EuxU2Int0_0),.clk(gclk));
	jdff dff_A_tmBL4v1l1_0(.dout(w_dff_A_EuxU2Int0_0),.din(w_dff_A_tmBL4v1l1_0),.clk(gclk));
	jdff dff_A_SZgxCPfN6_0(.dout(w_dff_A_tmBL4v1l1_0),.din(w_dff_A_SZgxCPfN6_0),.clk(gclk));
	jdff dff_A_2QJJym2f7_0(.dout(w_dff_A_SZgxCPfN6_0),.din(w_dff_A_2QJJym2f7_0),.clk(gclk));
	jdff dff_A_AiEo29PQ1_0(.dout(w_dff_A_2QJJym2f7_0),.din(w_dff_A_AiEo29PQ1_0),.clk(gclk));
	jdff dff_A_Gqltzonz4_0(.dout(w_dff_A_AiEo29PQ1_0),.din(w_dff_A_Gqltzonz4_0),.clk(gclk));
	jdff dff_A_6RJezA6N7_0(.dout(w_dff_A_Gqltzonz4_0),.din(w_dff_A_6RJezA6N7_0),.clk(gclk));
	jdff dff_A_cLTLoYju5_0(.dout(w_dff_A_6RJezA6N7_0),.din(w_dff_A_cLTLoYju5_0),.clk(gclk));
	jdff dff_A_xbB1niDx1_2(.dout(w_n620_0[2]),.din(w_dff_A_xbB1niDx1_2),.clk(gclk));
	jdff dff_A_HzjUXLGv1_2(.dout(w_dff_A_xbB1niDx1_2),.din(w_dff_A_HzjUXLGv1_2),.clk(gclk));
	jdff dff_A_uX9FTeu49_2(.dout(w_dff_A_HzjUXLGv1_2),.din(w_dff_A_uX9FTeu49_2),.clk(gclk));
	jdff dff_A_xm2zcuXS4_2(.dout(w_dff_A_uX9FTeu49_2),.din(w_dff_A_xm2zcuXS4_2),.clk(gclk));
	jdff dff_A_z9eqSGSK2_2(.dout(w_dff_A_xm2zcuXS4_2),.din(w_dff_A_z9eqSGSK2_2),.clk(gclk));
	jdff dff_A_6U9VqsfF3_2(.dout(w_dff_A_z9eqSGSK2_2),.din(w_dff_A_6U9VqsfF3_2),.clk(gclk));
	jdff dff_A_sH8FbVQ41_2(.dout(w_dff_A_6U9VqsfF3_2),.din(w_dff_A_sH8FbVQ41_2),.clk(gclk));
	jdff dff_A_ejUtGVit9_2(.dout(w_dff_A_sH8FbVQ41_2),.din(w_dff_A_ejUtGVit9_2),.clk(gclk));
	jdff dff_A_hh3UPOJj3_2(.dout(w_dff_A_ejUtGVit9_2),.din(w_dff_A_hh3UPOJj3_2),.clk(gclk));
	jdff dff_A_M3oKymkX0_2(.dout(w_dff_A_hh3UPOJj3_2),.din(w_dff_A_M3oKymkX0_2),.clk(gclk));
	jdff dff_A_pAH16aaE0_0(.dout(w_n619_0[0]),.din(w_dff_A_pAH16aaE0_0),.clk(gclk));
	jdff dff_A_EhRKcNdn1_0(.dout(w_dff_A_pAH16aaE0_0),.din(w_dff_A_EhRKcNdn1_0),.clk(gclk));
	jdff dff_A_kbRTm1KI5_0(.dout(w_dff_A_EhRKcNdn1_0),.din(w_dff_A_kbRTm1KI5_0),.clk(gclk));
	jdff dff_A_3F6v94TU0_0(.dout(w_dff_A_kbRTm1KI5_0),.din(w_dff_A_3F6v94TU0_0),.clk(gclk));
	jdff dff_A_jiZw6dXz8_0(.dout(w_dff_A_3F6v94TU0_0),.din(w_dff_A_jiZw6dXz8_0),.clk(gclk));
	jdff dff_A_gyGu27sC8_0(.dout(w_dff_A_jiZw6dXz8_0),.din(w_dff_A_gyGu27sC8_0),.clk(gclk));
	jdff dff_A_HzuVDqZY0_0(.dout(w_dff_A_gyGu27sC8_0),.din(w_dff_A_HzuVDqZY0_0),.clk(gclk));
	jdff dff_A_5ahwCGFI4_0(.dout(w_dff_A_HzuVDqZY0_0),.din(w_dff_A_5ahwCGFI4_0),.clk(gclk));
	jdff dff_A_pNIealtt9_0(.dout(w_dff_A_5ahwCGFI4_0),.din(w_dff_A_pNIealtt9_0),.clk(gclk));
	jdff dff_A_gUS2zuK58_0(.dout(w_dff_A_pNIealtt9_0),.din(w_dff_A_gUS2zuK58_0),.clk(gclk));
	jdff dff_A_FigNKfxo7_1(.dout(w_n619_0[1]),.din(w_dff_A_FigNKfxo7_1),.clk(gclk));
	jdff dff_A_260bEBTC6_1(.dout(w_dff_A_FigNKfxo7_1),.din(w_dff_A_260bEBTC6_1),.clk(gclk));
	jdff dff_A_VEn8q4z92_1(.dout(w_dff_A_260bEBTC6_1),.din(w_dff_A_VEn8q4z92_1),.clk(gclk));
	jdff dff_A_msprWaCP2_1(.dout(w_dff_A_VEn8q4z92_1),.din(w_dff_A_msprWaCP2_1),.clk(gclk));
	jdff dff_A_zdJ6DOrn3_1(.dout(w_dff_A_msprWaCP2_1),.din(w_dff_A_zdJ6DOrn3_1),.clk(gclk));
	jdff dff_A_2mkDxWwO8_1(.dout(w_dff_A_zdJ6DOrn3_1),.din(w_dff_A_2mkDxWwO8_1),.clk(gclk));
	jdff dff_A_XVHiTYCN8_1(.dout(w_dff_A_2mkDxWwO8_1),.din(w_dff_A_XVHiTYCN8_1),.clk(gclk));
	jdff dff_A_Gr4gVzGG9_1(.dout(w_dff_A_XVHiTYCN8_1),.din(w_dff_A_Gr4gVzGG9_1),.clk(gclk));
	jdff dff_A_pRUa8Ttq1_1(.dout(w_dff_A_Gr4gVzGG9_1),.din(w_dff_A_pRUa8Ttq1_1),.clk(gclk));
	jdff dff_A_zJ3ZWgMV1_0(.dout(w_n618_2[0]),.din(w_dff_A_zJ3ZWgMV1_0),.clk(gclk));
	jdff dff_A_4yptJBWd6_0(.dout(w_dff_A_zJ3ZWgMV1_0),.din(w_dff_A_4yptJBWd6_0),.clk(gclk));
	jdff dff_A_yjrrCu7o5_0(.dout(w_dff_A_4yptJBWd6_0),.din(w_dff_A_yjrrCu7o5_0),.clk(gclk));
	jdff dff_A_ibZVVIeY2_0(.dout(w_dff_A_yjrrCu7o5_0),.din(w_dff_A_ibZVVIeY2_0),.clk(gclk));
	jdff dff_A_DuypDAPN2_0(.dout(w_dff_A_ibZVVIeY2_0),.din(w_dff_A_DuypDAPN2_0),.clk(gclk));
	jdff dff_A_2kPYGMWC2_0(.dout(w_dff_A_DuypDAPN2_0),.din(w_dff_A_2kPYGMWC2_0),.clk(gclk));
	jdff dff_A_35poXltV8_0(.dout(w_dff_A_2kPYGMWC2_0),.din(w_dff_A_35poXltV8_0),.clk(gclk));
	jdff dff_A_TwCJsRjF2_0(.dout(w_dff_A_35poXltV8_0),.din(w_dff_A_TwCJsRjF2_0),.clk(gclk));
	jdff dff_A_SgxLCfYC5_0(.dout(w_dff_A_TwCJsRjF2_0),.din(w_dff_A_SgxLCfYC5_0),.clk(gclk));
	jdff dff_A_tFbVVaAs8_0(.dout(w_dff_A_SgxLCfYC5_0),.din(w_dff_A_tFbVVaAs8_0),.clk(gclk));
	jdff dff_A_oUZrYATW0_0(.dout(w_dff_A_tFbVVaAs8_0),.din(w_dff_A_oUZrYATW0_0),.clk(gclk));
	jdff dff_A_QFvgbUU20_0(.dout(w_dff_A_oUZrYATW0_0),.din(w_dff_A_QFvgbUU20_0),.clk(gclk));
	jdff dff_A_8kOfjuPP0_0(.dout(w_dff_A_QFvgbUU20_0),.din(w_dff_A_8kOfjuPP0_0),.clk(gclk));
	jdff dff_A_k7wsKiL36_2(.dout(w_n618_0[2]),.din(w_dff_A_k7wsKiL36_2),.clk(gclk));
	jdff dff_A_xf7JuvVR3_2(.dout(w_dff_A_k7wsKiL36_2),.din(w_dff_A_xf7JuvVR3_2),.clk(gclk));
	jdff dff_A_qemMsgKK9_2(.dout(w_dff_A_xf7JuvVR3_2),.din(w_dff_A_qemMsgKK9_2),.clk(gclk));
	jdff dff_A_HYhoACAY5_2(.dout(w_dff_A_qemMsgKK9_2),.din(w_dff_A_HYhoACAY5_2),.clk(gclk));
	jdff dff_A_w3mQjxe81_2(.dout(w_dff_A_HYhoACAY5_2),.din(w_dff_A_w3mQjxe81_2),.clk(gclk));
	jdff dff_A_zCGulpcr7_2(.dout(w_dff_A_w3mQjxe81_2),.din(w_dff_A_zCGulpcr7_2),.clk(gclk));
	jdff dff_A_0NDY6e3v0_2(.dout(w_dff_A_zCGulpcr7_2),.din(w_dff_A_0NDY6e3v0_2),.clk(gclk));
	jdff dff_A_W0WBHR8e2_2(.dout(w_dff_A_0NDY6e3v0_2),.din(w_dff_A_W0WBHR8e2_2),.clk(gclk));
	jdff dff_A_K0Pad6Ns8_2(.dout(w_dff_A_W0WBHR8e2_2),.din(w_dff_A_K0Pad6Ns8_2),.clk(gclk));
	jdff dff_A_4kzqbnWJ8_2(.dout(w_dff_A_K0Pad6Ns8_2),.din(w_dff_A_4kzqbnWJ8_2),.clk(gclk));
	jdff dff_A_yjipZPyy5_2(.dout(w_dff_A_4kzqbnWJ8_2),.din(w_dff_A_yjipZPyy5_2),.clk(gclk));
	jdff dff_A_V5rlJOz46_2(.dout(w_dff_A_yjipZPyy5_2),.din(w_dff_A_V5rlJOz46_2),.clk(gclk));
	jdff dff_A_I9dstlAO9_0(.dout(w_n153_5[0]),.din(w_dff_A_I9dstlAO9_0),.clk(gclk));
	jdff dff_A_JEtBTcVc0_0(.dout(w_dff_A_I9dstlAO9_0),.din(w_dff_A_JEtBTcVc0_0),.clk(gclk));
	jdff dff_A_xWn1uct69_0(.dout(w_dff_A_JEtBTcVc0_0),.din(w_dff_A_xWn1uct69_0),.clk(gclk));
	jdff dff_A_uk6JKueg4_0(.dout(w_dff_A_xWn1uct69_0),.din(w_dff_A_uk6JKueg4_0),.clk(gclk));
	jdff dff_A_cj41HD791_0(.dout(w_n153_1[0]),.din(w_dff_A_cj41HD791_0),.clk(gclk));
	jdff dff_A_RNoxb2dK4_0(.dout(w_dff_A_cj41HD791_0),.din(w_dff_A_RNoxb2dK4_0),.clk(gclk));
	jdff dff_B_w3v2F4oM6_1(.din(n615),.dout(w_dff_B_w3v2F4oM6_1),.clk(gclk));
	jdff dff_B_HIhbgpsC2_1(.din(w_dff_B_w3v2F4oM6_1),.dout(w_dff_B_HIhbgpsC2_1),.clk(gclk));
	jdff dff_B_mV0nW1Tm9_1(.din(w_dff_B_HIhbgpsC2_1),.dout(w_dff_B_mV0nW1Tm9_1),.clk(gclk));
	jdff dff_B_60ChBBxI3_1(.din(w_dff_B_mV0nW1Tm9_1),.dout(w_dff_B_60ChBBxI3_1),.clk(gclk));
	jdff dff_B_FKThuiyb9_1(.din(w_dff_B_60ChBBxI3_1),.dout(w_dff_B_FKThuiyb9_1),.clk(gclk));
	jdff dff_B_Od5Gk1gw0_1(.din(w_dff_B_FKThuiyb9_1),.dout(w_dff_B_Od5Gk1gw0_1),.clk(gclk));
	jdff dff_B_B3u4cSBY8_1(.din(w_dff_B_Od5Gk1gw0_1),.dout(w_dff_B_B3u4cSBY8_1),.clk(gclk));
	jdff dff_B_q8k9MOuf7_1(.din(w_dff_B_B3u4cSBY8_1),.dout(w_dff_B_q8k9MOuf7_1),.clk(gclk));
	jdff dff_B_KvJ7e3XT4_0(.din(n575),.dout(w_dff_B_KvJ7e3XT4_0),.clk(gclk));
	jdff dff_B_0Vssa9tt8_0(.din(w_dff_B_KvJ7e3XT4_0),.dout(w_dff_B_0Vssa9tt8_0),.clk(gclk));
	jdff dff_B_7xDTL5ru8_0(.din(w_dff_B_0Vssa9tt8_0),.dout(w_dff_B_7xDTL5ru8_0),.clk(gclk));
	jdff dff_B_jvbrpiFg4_0(.din(w_dff_B_7xDTL5ru8_0),.dout(w_dff_B_jvbrpiFg4_0),.clk(gclk));
	jdff dff_A_m7ctGy0p4_0(.dout(w_n567_4[0]),.din(w_dff_A_m7ctGy0p4_0),.clk(gclk));
	jdff dff_A_QGRxRHqV0_0(.dout(w_dff_A_m7ctGy0p4_0),.din(w_dff_A_QGRxRHqV0_0),.clk(gclk));
	jdff dff_A_NClwg5zS3_0(.dout(w_dff_A_QGRxRHqV0_0),.din(w_dff_A_NClwg5zS3_0),.clk(gclk));
	jdff dff_A_28EEJ0Sn8_0(.dout(w_dff_A_NClwg5zS3_0),.din(w_dff_A_28EEJ0Sn8_0),.clk(gclk));
	jdff dff_A_3rZZEYLc6_0(.dout(w_dff_A_28EEJ0Sn8_0),.din(w_dff_A_3rZZEYLc6_0),.clk(gclk));
	jdff dff_A_MEGH1NvO4_0(.dout(w_dff_A_3rZZEYLc6_0),.din(w_dff_A_MEGH1NvO4_0),.clk(gclk));
	jdff dff_A_uCmTs7TH7_0(.dout(w_dff_A_MEGH1NvO4_0),.din(w_dff_A_uCmTs7TH7_0),.clk(gclk));
	jdff dff_A_6TImLwIf6_0(.dout(w_dff_A_uCmTs7TH7_0),.din(w_dff_A_6TImLwIf6_0),.clk(gclk));
	jdff dff_A_kYHBqgOM8_0(.dout(w_n567_1[0]),.din(w_dff_A_kYHBqgOM8_0),.clk(gclk));
	jdff dff_A_VWP2JInt9_0(.dout(w_dff_A_kYHBqgOM8_0),.din(w_dff_A_VWP2JInt9_0),.clk(gclk));
	jdff dff_A_H10i0gnZ4_0(.dout(w_dff_A_VWP2JInt9_0),.din(w_dff_A_H10i0gnZ4_0),.clk(gclk));
	jdff dff_A_UdIxKefW1_2(.dout(w_n567_1[2]),.din(w_dff_A_UdIxKefW1_2),.clk(gclk));
	jdff dff_A_RFYth3pu9_2(.dout(w_dff_A_UdIxKefW1_2),.din(w_dff_A_RFYth3pu9_2),.clk(gclk));
	jdff dff_A_O7ydR7cm8_2(.dout(w_dff_A_RFYth3pu9_2),.din(w_dff_A_O7ydR7cm8_2),.clk(gclk));
	jdff dff_A_OV09zMKu6_2(.dout(w_dff_A_O7ydR7cm8_2),.din(w_dff_A_OV09zMKu6_2),.clk(gclk));
	jdff dff_A_0HMKhCxd2_2(.dout(w_dff_A_OV09zMKu6_2),.din(w_dff_A_0HMKhCxd2_2),.clk(gclk));
	jdff dff_A_393srodo3_2(.dout(w_dff_A_0HMKhCxd2_2),.din(w_dff_A_393srodo3_2),.clk(gclk));
	jdff dff_A_LTo0MXWQ5_2(.dout(w_dff_A_393srodo3_2),.din(w_dff_A_LTo0MXWQ5_2),.clk(gclk));
	jdff dff_A_BovatdL55_2(.dout(w_dff_A_LTo0MXWQ5_2),.din(w_dff_A_BovatdL55_2),.clk(gclk));
	jdff dff_A_icapLlXC4_2(.dout(w_dff_A_BovatdL55_2),.din(w_dff_A_icapLlXC4_2),.clk(gclk));
	jdff dff_A_hqzJ7BUz0_2(.dout(w_dff_A_icapLlXC4_2),.din(w_dff_A_hqzJ7BUz0_2),.clk(gclk));
	jdff dff_A_zyQLVVjd6_1(.dout(w_n567_0[1]),.din(w_dff_A_zyQLVVjd6_1),.clk(gclk));
	jdff dff_A_Oye7c9t85_1(.dout(w_dff_A_zyQLVVjd6_1),.din(w_dff_A_Oye7c9t85_1),.clk(gclk));
	jdff dff_A_AaWsLxke0_1(.dout(w_dff_A_Oye7c9t85_1),.din(w_dff_A_AaWsLxke0_1),.clk(gclk));
	jdff dff_A_cByZCHFb3_2(.dout(w_n567_0[2]),.din(w_dff_A_cByZCHFb3_2),.clk(gclk));
	jdff dff_A_MzwhkeoN1_2(.dout(w_dff_A_cByZCHFb3_2),.din(w_dff_A_MzwhkeoN1_2),.clk(gclk));
	jdff dff_A_VwmtA1gA7_1(.dout(w_n566_0[1]),.din(w_dff_A_VwmtA1gA7_1),.clk(gclk));
	jdff dff_A_Z2XBsqBC9_1(.dout(w_dff_A_VwmtA1gA7_1),.din(w_dff_A_Z2XBsqBC9_1),.clk(gclk));
	jdff dff_A_AfCrQjjM0_1(.dout(w_dff_A_Z2XBsqBC9_1),.din(w_dff_A_AfCrQjjM0_1),.clk(gclk));
	jdff dff_A_PuTXQgIf1_1(.dout(w_dff_A_AfCrQjjM0_1),.din(w_dff_A_PuTXQgIf1_1),.clk(gclk));
	jdff dff_A_az5jMjMD1_1(.dout(w_dff_A_PuTXQgIf1_1),.din(w_dff_A_az5jMjMD1_1),.clk(gclk));
	jdff dff_A_q0CypoSz6_2(.dout(w_n566_0[2]),.din(w_dff_A_q0CypoSz6_2),.clk(gclk));
	jdff dff_A_QXZO0qHl4_2(.dout(w_dff_A_q0CypoSz6_2),.din(w_dff_A_QXZO0qHl4_2),.clk(gclk));
	jdff dff_A_IHj1ibR70_2(.dout(w_dff_A_QXZO0qHl4_2),.din(w_dff_A_IHj1ibR70_2),.clk(gclk));
	jdff dff_A_JJmQXtTo5_2(.dout(w_dff_A_IHj1ibR70_2),.din(w_dff_A_JJmQXtTo5_2),.clk(gclk));
	jdff dff_A_00kALzpj4_2(.dout(w_dff_A_JJmQXtTo5_2),.din(w_dff_A_00kALzpj4_2),.clk(gclk));
	jdff dff_A_lJ5nagS34_0(.dout(w_G213_0[0]),.din(w_dff_A_lJ5nagS34_0),.clk(gclk));
	jdff dff_A_fFX9Wa6W5_2(.dout(w_G213_0[2]),.din(w_dff_A_fFX9Wa6W5_2),.clk(gclk));
	jdff dff_A_raF79JIE4_2(.dout(w_dff_A_fFX9Wa6W5_2),.din(w_dff_A_raF79JIE4_2),.clk(gclk));
	jdff dff_A_5xFSuWWJ2_1(.dout(w_G343_0[1]),.din(w_dff_A_5xFSuWWJ2_1),.clk(gclk));
	jdff dff_A_VH4fbc1h7_1(.dout(w_dff_A_5xFSuWWJ2_1),.din(w_dff_A_VH4fbc1h7_1),.clk(gclk));
	jdff dff_A_mLMEhh1X3_1(.dout(w_dff_A_VH4fbc1h7_1),.din(w_dff_A_mLMEhh1X3_1),.clk(gclk));
	jdff dff_A_aA2Efb6n2_1(.dout(w_dff_A_mLMEhh1X3_1),.din(w_dff_A_aA2Efb6n2_1),.clk(gclk));
	jdff dff_A_PyGxFW0l7_2(.dout(w_n198_0[2]),.din(w_dff_A_PyGxFW0l7_2),.clk(gclk));
	jdff dff_B_GES3CfPU6_1(.din(n193),.dout(w_dff_B_GES3CfPU6_1),.clk(gclk));
	jdff dff_B_tISGEVh33_1(.din(w_dff_B_GES3CfPU6_1),.dout(w_dff_B_tISGEVh33_1),.clk(gclk));
	jdff dff_A_3jLZoVp15_1(.dout(w_G190_4[1]),.din(w_dff_A_3jLZoVp15_1),.clk(gclk));
	jdff dff_A_ZmYTtGjP7_2(.dout(w_G190_4[2]),.din(w_dff_A_ZmYTtGjP7_2),.clk(gclk));
	jdff dff_A_hxtQ4qkq4_2(.dout(w_dff_A_ZmYTtGjP7_2),.din(w_dff_A_hxtQ4qkq4_2),.clk(gclk));
	jdff dff_A_eXXOSfVr4_0(.dout(w_G190_1[0]),.din(w_dff_A_eXXOSfVr4_0),.clk(gclk));
	jdff dff_A_pg2YfUI82_0(.dout(w_dff_A_eXXOSfVr4_0),.din(w_dff_A_pg2YfUI82_0),.clk(gclk));
	jdff dff_A_gKdiZiIb8_0(.dout(w_dff_A_pg2YfUI82_0),.din(w_dff_A_gKdiZiIb8_0),.clk(gclk));
	jdff dff_A_25PEjoF99_0(.dout(w_dff_A_gKdiZiIb8_0),.din(w_dff_A_25PEjoF99_0),.clk(gclk));
	jdff dff_A_e7aAggJJ6_0(.dout(w_dff_A_25PEjoF99_0),.din(w_dff_A_e7aAggJJ6_0),.clk(gclk));
	jdff dff_A_oUdYKSkV9_0(.dout(w_G190_0[0]),.din(w_dff_A_oUdYKSkV9_0),.clk(gclk));
	jdff dff_A_AOAazSbn8_0(.dout(w_dff_A_oUdYKSkV9_0),.din(w_dff_A_AOAazSbn8_0),.clk(gclk));
	jdff dff_A_268u0N709_2(.dout(w_G190_0[2]),.din(w_dff_A_268u0N709_2),.clk(gclk));
	jdff dff_A_KUBNllBB7_2(.dout(w_dff_A_268u0N709_2),.din(w_dff_A_KUBNllBB7_2),.clk(gclk));
	jdff dff_A_ZC8WDYmo0_2(.dout(w_dff_A_KUBNllBB7_2),.din(w_dff_A_ZC8WDYmo0_2),.clk(gclk));
	jdff dff_A_mrfJpwXB4_2(.dout(w_dff_A_ZC8WDYmo0_2),.din(w_dff_A_mrfJpwXB4_2),.clk(gclk));
	jdff dff_A_WrRtgUhA4_2(.dout(w_dff_A_mrfJpwXB4_2),.din(w_dff_A_WrRtgUhA4_2),.clk(gclk));
	jdff dff_A_Xcuel7Tg7_2(.dout(w_dff_A_WrRtgUhA4_2),.din(w_dff_A_Xcuel7Tg7_2),.clk(gclk));
	jdff dff_A_TufCRslF2_2(.dout(w_dff_A_Xcuel7Tg7_2),.din(w_dff_A_TufCRslF2_2),.clk(gclk));
	jdff dff_A_iPX7Z4Cu9_2(.dout(w_G200_0[2]),.din(w_dff_A_iPX7Z4Cu9_2),.clk(gclk));
	jdff dff_A_VefTAxdH1_2(.dout(w_dff_A_iPX7Z4Cu9_2),.din(w_dff_A_VefTAxdH1_2),.clk(gclk));
	jdff dff_A_cXO4wwz39_2(.dout(w_dff_A_VefTAxdH1_2),.din(w_dff_A_cXO4wwz39_2),.clk(gclk));
	jdff dff_A_Ldn2NI1j8_2(.dout(w_dff_A_cXO4wwz39_2),.din(w_dff_A_Ldn2NI1j8_2),.clk(gclk));
	jdff dff_A_ttA7cKY37_2(.dout(w_dff_A_Ldn2NI1j8_2),.din(w_dff_A_ttA7cKY37_2),.clk(gclk));
	jdff dff_A_jOAji8bc1_2(.dout(w_dff_A_ttA7cKY37_2),.din(w_dff_A_jOAji8bc1_2),.clk(gclk));
	jdff dff_A_8rxErzIf8_2(.dout(w_dff_A_jOAji8bc1_2),.din(w_dff_A_8rxErzIf8_2),.clk(gclk));
	jdff dff_A_7TIFVRkI6_2(.dout(w_dff_A_8rxErzIf8_2),.din(w_dff_A_7TIFVRkI6_2),.clk(gclk));
	jdff dff_A_NUfNMVn58_1(.dout(w_n192_0[1]),.din(w_dff_A_NUfNMVn58_1),.clk(gclk));
	jdff dff_A_oAfHk9in3_1(.dout(w_dff_A_NUfNMVn58_1),.din(w_dff_A_oAfHk9in3_1),.clk(gclk));
	jdff dff_B_2RLYosgE9_1(.din(n162),.dout(w_dff_B_2RLYosgE9_1),.clk(gclk));
	jdff dff_B_4iA5VZ472_1(.din(w_dff_B_2RLYosgE9_1),.dout(w_dff_B_4iA5VZ472_1),.clk(gclk));
	jdff dff_A_Uw9rA5Q79_1(.dout(w_n190_0[1]),.din(w_dff_A_Uw9rA5Q79_1),.clk(gclk));
	jdff dff_A_maUN2Flg6_1(.dout(w_n189_2[1]),.din(w_dff_A_maUN2Flg6_1),.clk(gclk));
	jdff dff_A_gb7dweU23_2(.dout(w_n189_2[2]),.din(w_dff_A_gb7dweU23_2),.clk(gclk));
	jdff dff_A_PeA8ptfg2_0(.dout(w_n189_0[0]),.din(w_dff_A_PeA8ptfg2_0),.clk(gclk));
	jdff dff_A_VNirrpwN2_0(.dout(w_dff_A_PeA8ptfg2_0),.din(w_dff_A_VNirrpwN2_0),.clk(gclk));
	jdff dff_A_50kHApfg2_0(.dout(w_dff_A_VNirrpwN2_0),.din(w_dff_A_50kHApfg2_0),.clk(gclk));
	jdff dff_A_o4b01Lh21_0(.dout(w_dff_A_50kHApfg2_0),.din(w_dff_A_o4b01Lh21_0),.clk(gclk));
	jdff dff_A_Ji9HKJb18_0(.dout(w_dff_A_o4b01Lh21_0),.din(w_dff_A_Ji9HKJb18_0),.clk(gclk));
	jdff dff_A_oKT7Ez0f7_0(.dout(w_dff_A_Ji9HKJb18_0),.din(w_dff_A_oKT7Ez0f7_0),.clk(gclk));
	jdff dff_A_xpS69ZrS3_1(.dout(w_n189_0[1]),.din(w_dff_A_xpS69ZrS3_1),.clk(gclk));
	jdff dff_A_yJts9i7G6_1(.dout(w_dff_A_xpS69ZrS3_1),.din(w_dff_A_yJts9i7G6_1),.clk(gclk));
	jdff dff_A_2yzE9Y8S6_1(.dout(w_dff_A_yJts9i7G6_1),.din(w_dff_A_2yzE9Y8S6_1),.clk(gclk));
	jdff dff_A_eM4pA4l30_1(.dout(w_dff_A_2yzE9Y8S6_1),.din(w_dff_A_eM4pA4l30_1),.clk(gclk));
	jdff dff_A_vn0SLuPI6_1(.dout(w_dff_A_eM4pA4l30_1),.din(w_dff_A_vn0SLuPI6_1),.clk(gclk));
	jdff dff_A_FPx0BJSn6_1(.dout(w_dff_A_vn0SLuPI6_1),.din(w_dff_A_FPx0BJSn6_1),.clk(gclk));
	jdff dff_A_UFx35RBF0_0(.dout(w_G179_2[0]),.din(w_dff_A_UFx35RBF0_0),.clk(gclk));
	jdff dff_A_uVC9z8PY3_0(.dout(w_dff_A_UFx35RBF0_0),.din(w_dff_A_uVC9z8PY3_0),.clk(gclk));
	jdff dff_A_HS9Rn81n8_0(.dout(w_dff_A_uVC9z8PY3_0),.din(w_dff_A_HS9Rn81n8_0),.clk(gclk));
	jdff dff_A_bSnjeapd9_0(.dout(w_dff_A_HS9Rn81n8_0),.din(w_dff_A_bSnjeapd9_0),.clk(gclk));
	jdff dff_A_Gbdxrt8p0_0(.dout(w_dff_A_bSnjeapd9_0),.din(w_dff_A_Gbdxrt8p0_0),.clk(gclk));
	jdff dff_A_jzvCaJzW7_0(.dout(w_dff_A_Gbdxrt8p0_0),.din(w_dff_A_jzvCaJzW7_0),.clk(gclk));
	jdff dff_A_W5jceAN66_0(.dout(w_dff_A_jzvCaJzW7_0),.din(w_dff_A_W5jceAN66_0),.clk(gclk));
	jdff dff_A_adNHm5Ts5_0(.dout(w_dff_A_W5jceAN66_0),.din(w_dff_A_adNHm5Ts5_0),.clk(gclk));
	jdff dff_A_VNW6KaN29_1(.dout(w_G179_2[1]),.din(w_dff_A_VNW6KaN29_1),.clk(gclk));
	jdff dff_A_Pncs4or61_1(.dout(w_dff_A_VNW6KaN29_1),.din(w_dff_A_Pncs4or61_1),.clk(gclk));
	jdff dff_A_cQgTutSB9_1(.dout(w_dff_A_Pncs4or61_1),.din(w_dff_A_cQgTutSB9_1),.clk(gclk));
	jdff dff_A_n8LNq6bN8_1(.dout(w_dff_A_cQgTutSB9_1),.din(w_dff_A_n8LNq6bN8_1),.clk(gclk));
	jdff dff_A_JGeeLpHH8_1(.dout(w_dff_A_n8LNq6bN8_1),.din(w_dff_A_JGeeLpHH8_1),.clk(gclk));
	jdff dff_A_6CZSu0Gw2_1(.dout(w_dff_A_JGeeLpHH8_1),.din(w_dff_A_6CZSu0Gw2_1),.clk(gclk));
	jdff dff_A_zdPn62Q54_1(.dout(w_dff_A_6CZSu0Gw2_1),.din(w_dff_A_zdPn62Q54_1),.clk(gclk));
	jdff dff_A_C1uqPPe31_1(.dout(w_dff_A_zdPn62Q54_1),.din(w_dff_A_C1uqPPe31_1),.clk(gclk));
	jdff dff_A_9CGFR2918_0(.dout(w_G179_0[0]),.din(w_dff_A_9CGFR2918_0),.clk(gclk));
	jdff dff_A_cB6r0kEd9_0(.dout(w_dff_A_9CGFR2918_0),.din(w_dff_A_cB6r0kEd9_0),.clk(gclk));
	jdff dff_A_PJ0ANXx23_0(.dout(w_dff_A_cB6r0kEd9_0),.din(w_dff_A_PJ0ANXx23_0),.clk(gclk));
	jdff dff_A_d28yZRUN3_0(.dout(w_dff_A_PJ0ANXx23_0),.din(w_dff_A_d28yZRUN3_0),.clk(gclk));
	jdff dff_A_8qmwtbr90_0(.dout(w_dff_A_d28yZRUN3_0),.din(w_dff_A_8qmwtbr90_0),.clk(gclk));
	jdff dff_A_dJhGqiUZ6_0(.dout(w_dff_A_8qmwtbr90_0),.din(w_dff_A_dJhGqiUZ6_0),.clk(gclk));
	jdff dff_A_RyIK6iYs2_0(.dout(w_dff_A_dJhGqiUZ6_0),.din(w_dff_A_RyIK6iYs2_0),.clk(gclk));
	jdff dff_A_kBLVlvFw4_0(.dout(w_dff_A_RyIK6iYs2_0),.din(w_dff_A_kBLVlvFw4_0),.clk(gclk));
	jdff dff_A_SyzkO7SL4_1(.dout(w_n186_0[1]),.din(w_dff_A_SyzkO7SL4_1),.clk(gclk));
	jdff dff_B_GcnqWhjj5_0(.din(n184),.dout(w_dff_B_GcnqWhjj5_0),.clk(gclk));
	jdff dff_A_21LTCwyy0_0(.dout(w_G270_0[0]),.din(w_dff_A_21LTCwyy0_0),.clk(gclk));
	jdff dff_A_5Os4Co0L7_0(.dout(w_dff_A_21LTCwyy0_0),.din(w_dff_A_5Os4Co0L7_0),.clk(gclk));
	jdff dff_A_D30XsiAm4_0(.dout(w_dff_A_5Os4Co0L7_0),.din(w_dff_A_D30XsiAm4_0),.clk(gclk));
	jdff dff_A_AYEVyLfQ3_1(.dout(w_G270_0[1]),.din(w_dff_A_AYEVyLfQ3_1),.clk(gclk));
	jdff dff_B_dI5peQw07_1(.din(n174),.dout(w_dff_B_dI5peQw07_1),.clk(gclk));
	jdff dff_B_SJl0iTHM2_1(.din(n175),.dout(w_dff_B_SJl0iTHM2_1),.clk(gclk));
	jdff dff_B_BgZDjfnJ5_1(.din(w_dff_B_SJl0iTHM2_1),.dout(w_dff_B_BgZDjfnJ5_1),.clk(gclk));
	jdff dff_A_Yay1H0sT4_0(.dout(w_G257_1[0]),.din(w_dff_A_Yay1H0sT4_0),.clk(gclk));
	jdff dff_A_XjVZ48HX4_0(.dout(w_dff_A_Yay1H0sT4_0),.din(w_dff_A_XjVZ48HX4_0),.clk(gclk));
	jdff dff_A_8O7tS3tU4_1(.dout(w_G257_0[1]),.din(w_dff_A_8O7tS3tU4_1),.clk(gclk));
	jdff dff_A_axQXsGFK3_1(.dout(w_dff_A_8O7tS3tU4_1),.din(w_dff_A_axQXsGFK3_1),.clk(gclk));
	jdff dff_A_LseBYIOK8_1(.dout(w_dff_A_axQXsGFK3_1),.din(w_dff_A_LseBYIOK8_1),.clk(gclk));
	jdff dff_A_DwDyRc4z4_2(.dout(w_G257_0[2]),.din(w_dff_A_DwDyRc4z4_2),.clk(gclk));
	jdff dff_A_TGsmLIqQ6_2(.dout(w_dff_A_DwDyRc4z4_2),.din(w_dff_A_TGsmLIqQ6_2),.clk(gclk));
	jdff dff_A_sAjQKnIV0_0(.dout(w_G303_2[0]),.din(w_dff_A_sAjQKnIV0_0),.clk(gclk));
	jdff dff_A_25Ixg5Bz5_0(.dout(w_dff_A_sAjQKnIV0_0),.din(w_dff_A_25Ixg5Bz5_0),.clk(gclk));
	jdff dff_A_hMpawB0o6_0(.dout(w_dff_A_25Ixg5Bz5_0),.din(w_dff_A_hMpawB0o6_0),.clk(gclk));
	jdff dff_A_J7DcwswV9_1(.dout(w_G303_2[1]),.din(w_dff_A_J7DcwswV9_1),.clk(gclk));
	jdff dff_A_VvwDY8HE4_1(.dout(w_dff_A_J7DcwswV9_1),.din(w_dff_A_VvwDY8HE4_1),.clk(gclk));
	jdff dff_A_Z1eKN7YO8_1(.dout(w_dff_A_VvwDY8HE4_1),.din(w_dff_A_Z1eKN7YO8_1),.clk(gclk));
	jdff dff_A_tA4WwVps9_0(.dout(w_G303_0[0]),.din(w_dff_A_tA4WwVps9_0),.clk(gclk));
	jdff dff_A_MY4gmzcB6_0(.dout(w_dff_A_tA4WwVps9_0),.din(w_dff_A_MY4gmzcB6_0),.clk(gclk));
	jdff dff_A_5em3aR5A7_0(.dout(w_dff_A_MY4gmzcB6_0),.din(w_dff_A_5em3aR5A7_0),.clk(gclk));
	jdff dff_A_Yu7uDWyd5_2(.dout(w_G303_0[2]),.din(w_dff_A_Yu7uDWyd5_2),.clk(gclk));
	jdff dff_A_jhzE4bo43_2(.dout(w_dff_A_Yu7uDWyd5_2),.din(w_dff_A_jhzE4bo43_2),.clk(gclk));
	jdff dff_A_K6oeFYj22_2(.dout(w_dff_A_jhzE4bo43_2),.din(w_dff_A_K6oeFYj22_2),.clk(gclk));
	jdff dff_A_qt1GiljN0_2(.dout(w_dff_A_K6oeFYj22_2),.din(w_dff_A_qt1GiljN0_2),.clk(gclk));
	jdff dff_A_rzrEgui05_2(.dout(w_G1698_0[2]),.din(w_dff_A_rzrEgui05_2),.clk(gclk));
	jdff dff_A_m34ss2Ex2_0(.dout(w_G264_0[0]),.din(w_dff_A_m34ss2Ex2_0),.clk(gclk));
	jdff dff_A_2kBUp0gP7_0(.dout(w_dff_A_m34ss2Ex2_0),.din(w_dff_A_2kBUp0gP7_0),.clk(gclk));
	jdff dff_A_B212phLv9_0(.dout(w_dff_A_2kBUp0gP7_0),.din(w_dff_A_B212phLv9_0),.clk(gclk));
	jdff dff_A_iK7dFzir4_1(.dout(w_G264_0[1]),.din(w_dff_A_iK7dFzir4_1),.clk(gclk));
	jdff dff_A_ahXSG8UL4_1(.dout(w_dff_A_iK7dFzir4_1),.din(w_dff_A_ahXSG8UL4_1),.clk(gclk));
	jdff dff_A_ceBD7C2p2_1(.dout(w_n172_4[1]),.din(w_dff_A_ceBD7C2p2_1),.clk(gclk));
	jdff dff_A_re8iwzaB9_1(.dout(w_dff_A_ceBD7C2p2_1),.din(w_dff_A_re8iwzaB9_1),.clk(gclk));
	jdff dff_A_GVkq5jlA9_2(.dout(w_n172_4[2]),.din(w_dff_A_GVkq5jlA9_2),.clk(gclk));
	jdff dff_A_qhl06zxv1_2(.dout(w_dff_A_GVkq5jlA9_2),.din(w_dff_A_qhl06zxv1_2),.clk(gclk));
	jdff dff_A_XKjLqvyA4_1(.dout(w_n172_1[1]),.din(w_dff_A_XKjLqvyA4_1),.clk(gclk));
	jdff dff_A_NwQFKoZl5_1(.dout(w_dff_A_XKjLqvyA4_1),.din(w_dff_A_NwQFKoZl5_1),.clk(gclk));
	jdff dff_A_bW7EyHf57_2(.dout(w_n172_1[2]),.din(w_dff_A_bW7EyHf57_2),.clk(gclk));
	jdff dff_A_dZmAmqcr4_2(.dout(w_dff_A_bW7EyHf57_2),.din(w_dff_A_dZmAmqcr4_2),.clk(gclk));
	jdff dff_A_MW926Uyt6_1(.dout(w_n172_0[1]),.din(w_dff_A_MW926Uyt6_1),.clk(gclk));
	jdff dff_A_a7OroNKR0_1(.dout(w_dff_A_MW926Uyt6_1),.din(w_dff_A_a7OroNKR0_1),.clk(gclk));
	jdff dff_A_4NqUh69t6_2(.dout(w_n172_0[2]),.din(w_dff_A_4NqUh69t6_2),.clk(gclk));
	jdff dff_A_rPcvYyJw0_2(.dout(w_dff_A_4NqUh69t6_2),.din(w_dff_A_rPcvYyJw0_2),.clk(gclk));
	jdff dff_A_YJlh3oE04_2(.dout(w_n170_0[2]),.din(w_dff_A_YJlh3oE04_2),.clk(gclk));
	jdff dff_B_j1gpmBTM4_3(.din(n170),.dout(w_dff_B_j1gpmBTM4_3),.clk(gclk));
	jdff dff_A_XTFGpIVr3_1(.dout(w_n167_0[1]),.din(w_dff_A_XTFGpIVr3_1),.clk(gclk));
	jdff dff_A_yD4Oi5hU0_0(.dout(w_G274_0[0]),.din(w_dff_A_yD4Oi5hU0_0),.clk(gclk));
	jdff dff_A_u6jQZWCN8_0(.dout(w_dff_A_yD4Oi5hU0_0),.din(w_dff_A_u6jQZWCN8_0),.clk(gclk));
	jdff dff_A_NSZ2h9dl9_2(.dout(w_G274_0[2]),.din(w_dff_A_NSZ2h9dl9_2),.clk(gclk));
	jdff dff_A_03ahk3n16_2(.dout(w_dff_A_NSZ2h9dl9_2),.din(w_dff_A_03ahk3n16_2),.clk(gclk));
	jdff dff_A_GSO5PdCL6_2(.dout(w_dff_A_03ahk3n16_2),.din(w_dff_A_GSO5PdCL6_2),.clk(gclk));
	jdff dff_A_kNaDVNSq3_1(.dout(w_n165_0[1]),.din(w_dff_A_kNaDVNSq3_1),.clk(gclk));
	jdff dff_A_gIp1idMr6_1(.dout(w_G45_1[1]),.din(w_dff_A_gIp1idMr6_1),.clk(gclk));
	jdff dff_A_jjyOFsE86_0(.dout(w_n142_1[0]),.din(w_dff_A_jjyOFsE86_0),.clk(gclk));
	jdff dff_A_NeFbVxgv6_0(.dout(w_dff_A_jjyOFsE86_0),.din(w_dff_A_NeFbVxgv6_0),.clk(gclk));
	jdff dff_A_MncSweYv9_0(.dout(w_dff_A_NeFbVxgv6_0),.din(w_dff_A_MncSweYv9_0),.clk(gclk));
	jdff dff_A_gw5ysKeH9_0(.dout(w_dff_A_MncSweYv9_0),.din(w_dff_A_gw5ysKeH9_0),.clk(gclk));
	jdff dff_A_pLAuYhxD6_0(.dout(w_dff_A_gw5ysKeH9_0),.din(w_dff_A_pLAuYhxD6_0),.clk(gclk));
	jdff dff_A_xCWnU4zI3_0(.dout(w_dff_A_pLAuYhxD6_0),.din(w_dff_A_xCWnU4zI3_0),.clk(gclk));
	jdff dff_A_duVIurAX0_0(.dout(w_dff_A_xCWnU4zI3_0),.din(w_dff_A_duVIurAX0_0),.clk(gclk));
	jdff dff_A_H7Vs399g6_0(.dout(w_dff_A_duVIurAX0_0),.din(w_dff_A_H7Vs399g6_0),.clk(gclk));
	jdff dff_A_8yMCUGnd6_0(.dout(w_dff_A_H7Vs399g6_0),.din(w_dff_A_8yMCUGnd6_0),.clk(gclk));
	jdff dff_A_ei1SxWmQ4_0(.dout(w_dff_A_8yMCUGnd6_0),.din(w_dff_A_ei1SxWmQ4_0),.clk(gclk));
	jdff dff_A_XdMqc9jc1_0(.dout(w_dff_A_ei1SxWmQ4_0),.din(w_dff_A_XdMqc9jc1_0),.clk(gclk));
	jdff dff_A_fqjEorEV0_0(.dout(w_dff_A_XdMqc9jc1_0),.din(w_dff_A_fqjEorEV0_0),.clk(gclk));
	jdff dff_A_4moNnSnd2_0(.dout(w_dff_A_fqjEorEV0_0),.din(w_dff_A_4moNnSnd2_0),.clk(gclk));
	jdff dff_A_p9d7fzAb5_0(.dout(w_dff_A_4moNnSnd2_0),.din(w_dff_A_p9d7fzAb5_0),.clk(gclk));
	jdff dff_A_DdA5je7k2_0(.dout(w_dff_A_p9d7fzAb5_0),.din(w_dff_A_DdA5je7k2_0),.clk(gclk));
	jdff dff_A_LwCLSk4Q9_0(.dout(w_dff_A_DdA5je7k2_0),.din(w_dff_A_LwCLSk4Q9_0),.clk(gclk));
	jdff dff_A_F2uvRqSV5_0(.dout(w_dff_A_LwCLSk4Q9_0),.din(w_dff_A_F2uvRqSV5_0),.clk(gclk));
	jdff dff_A_RfddQYn10_0(.dout(w_dff_A_F2uvRqSV5_0),.din(w_dff_A_RfddQYn10_0),.clk(gclk));
	jdff dff_A_Ehupaxh00_1(.dout(w_n163_1[1]),.din(w_dff_A_Ehupaxh00_1),.clk(gclk));
	jdff dff_A_XM8BCtkG6_1(.dout(w_G169_3[1]),.din(w_dff_A_XM8BCtkG6_1),.clk(gclk));
	jdff dff_A_BVNBrHJ22_1(.dout(w_dff_A_XM8BCtkG6_1),.din(w_dff_A_BVNBrHJ22_1),.clk(gclk));
	jdff dff_A_SFIRQzNx1_1(.dout(w_dff_A_BVNBrHJ22_1),.din(w_dff_A_SFIRQzNx1_1),.clk(gclk));
	jdff dff_A_wP7iAD9G9_1(.dout(w_dff_A_SFIRQzNx1_1),.din(w_dff_A_wP7iAD9G9_1),.clk(gclk));
	jdff dff_A_9MtHASw25_1(.dout(w_dff_A_wP7iAD9G9_1),.din(w_dff_A_9MtHASw25_1),.clk(gclk));
	jdff dff_A_OEB2aHrV7_1(.dout(w_dff_A_9MtHASw25_1),.din(w_dff_A_OEB2aHrV7_1),.clk(gclk));
	jdff dff_A_WrA9bOyU1_1(.dout(w_dff_A_OEB2aHrV7_1),.din(w_dff_A_WrA9bOyU1_1),.clk(gclk));
	jdff dff_A_53LigxUI3_1(.dout(w_dff_A_WrA9bOyU1_1),.din(w_dff_A_53LigxUI3_1),.clk(gclk));
	jdff dff_A_GBIGJCYs5_0(.dout(w_G169_0[0]),.din(w_dff_A_GBIGJCYs5_0),.clk(gclk));
	jdff dff_A_QgG4Hyin7_1(.dout(w_G169_0[1]),.din(w_dff_A_QgG4Hyin7_1),.clk(gclk));
	jdff dff_A_lQQRhe7H8_1(.dout(w_dff_A_QgG4Hyin7_1),.din(w_dff_A_lQQRhe7H8_1),.clk(gclk));
	jdff dff_A_yt34euw66_1(.dout(w_dff_A_lQQRhe7H8_1),.din(w_dff_A_yt34euw66_1),.clk(gclk));
	jdff dff_A_ON8lIAsy5_1(.dout(w_dff_A_yt34euw66_1),.din(w_dff_A_ON8lIAsy5_1),.clk(gclk));
	jdff dff_A_iyrgdOn12_1(.dout(w_dff_A_ON8lIAsy5_1),.din(w_dff_A_iyrgdOn12_1),.clk(gclk));
	jdff dff_A_Zd6KN2l20_1(.dout(w_dff_A_iyrgdOn12_1),.din(w_dff_A_Zd6KN2l20_1),.clk(gclk));
	jdff dff_A_Gi5qJDve0_1(.dout(w_dff_A_Zd6KN2l20_1),.din(w_dff_A_Gi5qJDve0_1),.clk(gclk));
	jdff dff_A_N0M2Dwtu1_1(.dout(w_n161_0[1]),.din(w_dff_A_N0M2Dwtu1_1),.clk(gclk));
	jdff dff_A_agZidya10_1(.dout(w_dff_A_N0M2Dwtu1_1),.din(w_dff_A_agZidya10_1),.clk(gclk));
	jdff dff_B_izbAE8qO7_0(.din(n159),.dout(w_dff_B_izbAE8qO7_0),.clk(gclk));
	jdff dff_B_M2hcu2Iu9_0(.din(w_dff_B_izbAE8qO7_0),.dout(w_dff_B_M2hcu2Iu9_0),.clk(gclk));
	jdff dff_A_wyilZyJB0_0(.dout(w_n105_1[0]),.din(w_dff_A_wyilZyJB0_0),.clk(gclk));
	jdff dff_A_qgWVCfvQ1_0(.dout(w_dff_A_wyilZyJB0_0),.din(w_dff_A_qgWVCfvQ1_0),.clk(gclk));
	jdff dff_A_awxo882Y8_1(.dout(w_n105_0[1]),.din(w_dff_A_awxo882Y8_1),.clk(gclk));
	jdff dff_A_AzWh0D143_1(.dout(w_dff_A_awxo882Y8_1),.din(w_dff_A_AzWh0D143_1),.clk(gclk));
	jdff dff_A_TB5hfQ0o8_1(.dout(w_dff_A_AzWh0D143_1),.din(w_dff_A_TB5hfQ0o8_1),.clk(gclk));
	jdff dff_A_6gcDyPwH1_2(.dout(w_n105_0[2]),.din(w_dff_A_6gcDyPwH1_2),.clk(gclk));
	jdff dff_A_p1Lv5tZs8_2(.dout(w_dff_A_6gcDyPwH1_2),.din(w_dff_A_p1Lv5tZs8_2),.clk(gclk));
	jdff dff_B_ZZIFyYAI8_1(.din(n150),.dout(w_dff_B_ZZIFyYAI8_1),.clk(gclk));
	jdff dff_B_FzHTR9pu7_1(.din(w_dff_B_ZZIFyYAI8_1),.dout(w_dff_B_FzHTR9pu7_1),.clk(gclk));
	jdff dff_B_QKp3wjYK2_1(.din(w_dff_B_FzHTR9pu7_1),.dout(w_dff_B_QKp3wjYK2_1),.clk(gclk));
	jdff dff_A_sDaQeqU74_0(.dout(w_G97_4[0]),.din(w_dff_A_sDaQeqU74_0),.clk(gclk));
	jdff dff_A_WKeEDn6S5_1(.dout(w_G97_1[1]),.din(w_dff_A_WKeEDn6S5_1),.clk(gclk));
	jdff dff_A_CueYVveM3_1(.dout(w_dff_A_WKeEDn6S5_1),.din(w_dff_A_CueYVveM3_1),.clk(gclk));
	jdff dff_A_l8TPzBcC4_1(.dout(w_dff_A_CueYVveM3_1),.din(w_dff_A_l8TPzBcC4_1),.clk(gclk));
	jdff dff_A_Yg7is76d4_2(.dout(w_G97_1[2]),.din(w_dff_A_Yg7is76d4_2),.clk(gclk));
	jdff dff_A_xewqMdmD6_2(.dout(w_dff_A_Yg7is76d4_2),.din(w_dff_A_xewqMdmD6_2),.clk(gclk));
	jdff dff_A_6yYBYou13_2(.dout(w_dff_A_xewqMdmD6_2),.din(w_dff_A_6yYBYou13_2),.clk(gclk));
	jdff dff_A_jbusTZln6_1(.dout(w_G97_0[1]),.din(w_dff_A_jbusTZln6_1),.clk(gclk));
	jdff dff_A_0EFK6krm0_1(.dout(w_dff_A_jbusTZln6_1),.din(w_dff_A_0EFK6krm0_1),.clk(gclk));
	jdff dff_A_ytpqUgnf0_1(.dout(w_dff_A_0EFK6krm0_1),.din(w_dff_A_ytpqUgnf0_1),.clk(gclk));
	jdff dff_A_p63nj3rN5_2(.dout(w_n153_2[2]),.din(w_dff_A_p63nj3rN5_2),.clk(gclk));
	jdff dff_A_wGwwfJCx9_2(.dout(w_dff_A_p63nj3rN5_2),.din(w_dff_A_wGwwfJCx9_2),.clk(gclk));
	jdff dff_A_hPOLBwJu3_2(.dout(w_dff_A_wGwwfJCx9_2),.din(w_dff_A_hPOLBwJu3_2),.clk(gclk));
	jdff dff_A_dZAaiECU3_2(.dout(w_dff_A_hPOLBwJu3_2),.din(w_dff_A_dZAaiECU3_2),.clk(gclk));
	jdff dff_A_Xo8Car738_2(.dout(w_n153_0[2]),.din(w_dff_A_Xo8Car738_2),.clk(gclk));
	jdff dff_A_tJ7Qxpoe3_2(.dout(w_dff_A_Xo8Car738_2),.din(w_dff_A_tJ7Qxpoe3_2),.clk(gclk));
	jdff dff_A_y8uCNX1z9_2(.dout(w_dff_A_tJ7Qxpoe3_2),.din(w_dff_A_y8uCNX1z9_2),.clk(gclk));
	jdff dff_A_9ngiHv6q8_0(.dout(w_n152_0[0]),.din(w_dff_A_9ngiHv6q8_0),.clk(gclk));
	jdff dff_A_oJeBx24G4_0(.dout(w_dff_A_9ngiHv6q8_0),.din(w_dff_A_oJeBx24G4_0),.clk(gclk));
	jdff dff_A_UWfbyl1h1_2(.dout(w_n152_0[2]),.din(w_dff_A_UWfbyl1h1_2),.clk(gclk));
	jdff dff_A_bxpFVpxw1_0(.dout(w_G283_3[0]),.din(w_dff_A_bxpFVpxw1_0),.clk(gclk));
	jdff dff_A_DcWhLFiX8_0(.dout(w_dff_A_bxpFVpxw1_0),.din(w_dff_A_DcWhLFiX8_0),.clk(gclk));
	jdff dff_A_UMyuYaC41_0(.dout(w_dff_A_DcWhLFiX8_0),.din(w_dff_A_UMyuYaC41_0),.clk(gclk));
	jdff dff_A_VPcXu3Td2_1(.dout(w_G283_3[1]),.din(w_dff_A_VPcXu3Td2_1),.clk(gclk));
	jdff dff_A_0daeuNOR1_1(.dout(w_dff_A_VPcXu3Td2_1),.din(w_dff_A_0daeuNOR1_1),.clk(gclk));
	jdff dff_A_OcKfnYpe3_1(.dout(w_dff_A_0daeuNOR1_1),.din(w_dff_A_OcKfnYpe3_1),.clk(gclk));
	jdff dff_A_NqqpT5bS4_0(.dout(w_G283_0[0]),.din(w_dff_A_NqqpT5bS4_0),.clk(gclk));
	jdff dff_A_DXX6RVdY6_0(.dout(w_dff_A_NqqpT5bS4_0),.din(w_dff_A_DXX6RVdY6_0),.clk(gclk));
	jdff dff_A_G7tY3cCa7_0(.dout(w_dff_A_DXX6RVdY6_0),.din(w_dff_A_G7tY3cCa7_0),.clk(gclk));
	jdff dff_A_raukKi4E5_1(.dout(w_G283_0[1]),.din(w_dff_A_raukKi4E5_1),.clk(gclk));
	jdff dff_A_W7JmUWlk9_1(.dout(w_dff_A_raukKi4E5_1),.din(w_dff_A_W7JmUWlk9_1),.clk(gclk));
	jdff dff_A_IrXp32UJ4_1(.dout(w_dff_A_W7JmUWlk9_1),.din(w_dff_A_IrXp32UJ4_1),.clk(gclk));
	jdff dff_A_lypYdccR6_0(.dout(w_n151_6[0]),.din(w_dff_A_lypYdccR6_0),.clk(gclk));
	jdff dff_A_QoYS69xf0_1(.dout(w_n151_1[1]),.din(w_dff_A_QoYS69xf0_1),.clk(gclk));
	jdff dff_A_rMTa615l0_2(.dout(w_n151_1[2]),.din(w_dff_A_rMTa615l0_2),.clk(gclk));
	jdff dff_A_J6xfLXCV2_2(.dout(w_dff_A_rMTa615l0_2),.din(w_dff_A_J6xfLXCV2_2),.clk(gclk));
	jdff dff_A_rB8oE75a0_0(.dout(w_G116_4[0]),.din(w_dff_A_rB8oE75a0_0),.clk(gclk));
	jdff dff_A_rrN7MSkv5_0(.dout(w_dff_A_rB8oE75a0_0),.din(w_dff_A_rrN7MSkv5_0),.clk(gclk));
	jdff dff_A_aCfmhJLD5_0(.dout(w_dff_A_rrN7MSkv5_0),.din(w_dff_A_aCfmhJLD5_0),.clk(gclk));
	jdff dff_B_myevPPDS9_0(.din(n146),.dout(w_dff_B_myevPPDS9_0),.clk(gclk));
	jdff dff_B_TWpw5Lkn9_0(.din(w_dff_B_myevPPDS9_0),.dout(w_dff_B_TWpw5Lkn9_0),.clk(gclk));
	jdff dff_A_1QcmdyLC6_0(.dout(w_n141_3[0]),.din(w_dff_A_1QcmdyLC6_0),.clk(gclk));
	jdff dff_A_H7EoIeNt4_0(.dout(w_dff_A_1QcmdyLC6_0),.din(w_dff_A_H7EoIeNt4_0),.clk(gclk));
	jdff dff_A_4G19A59n2_1(.dout(w_G33_12[1]),.din(w_dff_A_4G19A59n2_1),.clk(gclk));
	jdff dff_A_6UMkh2iw9_2(.dout(w_G33_12[2]),.din(w_dff_A_6UMkh2iw9_2),.clk(gclk));
	jdff dff_A_JUyi6zAp5_0(.dout(w_G33_0[0]),.din(w_dff_A_JUyi6zAp5_0),.clk(gclk));
	jdff dff_A_7hmPxE388_0(.dout(w_dff_A_JUyi6zAp5_0),.din(w_dff_A_7hmPxE388_0),.clk(gclk));
	jdff dff_A_Fe2KaN991_0(.dout(w_dff_A_7hmPxE388_0),.din(w_dff_A_Fe2KaN991_0),.clk(gclk));
	jdff dff_A_4m3fVzqZ7_0(.dout(w_n139_1[0]),.din(w_dff_A_4m3fVzqZ7_0),.clk(gclk));
	jdff dff_A_Xf56kWhH1_2(.dout(w_n139_1[2]),.din(w_dff_A_Xf56kWhH1_2),.clk(gclk));
	jdff dff_A_TYwDA2GO3_0(.dout(w_G13_1[0]),.din(w_dff_A_TYwDA2GO3_0),.clk(gclk));
	jdff dff_A_a2pL4i4R6_0(.dout(w_dff_A_TYwDA2GO3_0),.din(w_dff_A_a2pL4i4R6_0),.clk(gclk));
	jdff dff_A_DU8SRIU89_1(.dout(w_G13_1[1]),.din(w_dff_A_DU8SRIU89_1),.clk(gclk));
	jdff dff_A_XtbjMlao6_0(.dout(w_G116_5[0]),.din(w_dff_A_XtbjMlao6_0),.clk(gclk));
	jdff dff_A_fBrIb4Yj7_0(.dout(w_dff_A_XtbjMlao6_0),.din(w_dff_A_fBrIb4Yj7_0),.clk(gclk));
	jdff dff_A_t1IPvC8r1_0(.dout(w_dff_A_fBrIb4Yj7_0),.din(w_dff_A_t1IPvC8r1_0),.clk(gclk));
	jdff dff_A_ksJxD0uI3_0(.dout(w_dff_A_t1IPvC8r1_0),.din(w_dff_A_ksJxD0uI3_0),.clk(gclk));
	jdff dff_A_Y9rTJxB16_0(.dout(w_dff_A_ksJxD0uI3_0),.din(w_dff_A_Y9rTJxB16_0),.clk(gclk));
	jdff dff_A_cIXMQj1C0_0(.dout(w_dff_A_Y9rTJxB16_0),.din(w_dff_A_cIXMQj1C0_0),.clk(gclk));
	jdff dff_A_VKaiihHm3_1(.dout(w_G116_5[1]),.din(w_dff_A_VKaiihHm3_1),.clk(gclk));
	jdff dff_A_AhkhnfD37_2(.dout(w_G116_1[2]),.din(w_dff_A_AhkhnfD37_2),.clk(gclk));
	jdff dff_A_FPq6sE740_2(.dout(w_dff_A_AhkhnfD37_2),.din(w_dff_A_FPq6sE740_2),.clk(gclk));
	jdff dff_A_7FnPaeON8_2(.dout(w_dff_A_FPq6sE740_2),.din(w_dff_A_7FnPaeON8_2),.clk(gclk));
	jdff dff_A_1mvVggJS4_1(.dout(w_G116_0[1]),.din(w_dff_A_1mvVggJS4_1),.clk(gclk));
	jdff dff_A_wYohYmHl8_1(.dout(w_dff_A_1mvVggJS4_1),.din(w_dff_A_wYohYmHl8_1),.clk(gclk));
	jdff dff_A_6Jnib6tG3_1(.dout(w_dff_A_wYohYmHl8_1),.din(w_dff_A_6Jnib6tG3_1),.clk(gclk));
	jdff dff_A_v6Tm0TTV7_2(.dout(w_G116_0[2]),.din(w_dff_A_v6Tm0TTV7_2),.clk(gclk));
	jdff dff_A_OWUQhYUJ5_2(.dout(w_dff_A_v6Tm0TTV7_2),.din(w_dff_A_OWUQhYUJ5_2),.clk(gclk));
	jdff dff_A_7SiU0GIE8_2(.dout(w_dff_A_OWUQhYUJ5_2),.din(w_dff_A_7SiU0GIE8_2),.clk(gclk));
	jdff dff_A_92WyQHFf7_0(.dout(w_G330_0[0]),.din(w_dff_A_92WyQHFf7_0),.clk(gclk));
	jdff dff_A_2LB4S6lL1_2(.dout(w_G330_0[2]),.din(w_dff_A_2LB4S6lL1_2),.clk(gclk));
	jdff dff_B_KJmYe58O5_3(.din(G330),.dout(w_dff_B_KJmYe58O5_3),.clk(gclk));
	jdff dff_B_ni0jTr7x7_3(.din(w_dff_B_KJmYe58O5_3),.dout(w_dff_B_ni0jTr7x7_3),.clk(gclk));
	jdff dff_B_6bk3x7n79_3(.din(w_dff_B_ni0jTr7x7_3),.dout(w_dff_B_6bk3x7n79_3),.clk(gclk));
	jdff dff_B_rHPmGMoo8_3(.din(w_dff_B_6bk3x7n79_3),.dout(w_dff_B_rHPmGMoo8_3),.clk(gclk));
	jdff dff_B_90HfVKk17_3(.din(w_dff_B_rHPmGMoo8_3),.dout(w_dff_B_90HfVKk17_3),.clk(gclk));
	jdff dff_B_5gC5FILO3_3(.din(w_dff_B_90HfVKk17_3),.dout(w_dff_B_5gC5FILO3_3),.clk(gclk));
	jdff dff_B_qbxsD1Wv8_3(.din(w_dff_B_5gC5FILO3_3),.dout(w_dff_B_qbxsD1Wv8_3),.clk(gclk));
	jdff dff_B_MahJQJth5_3(.din(w_dff_B_qbxsD1Wv8_3),.dout(w_dff_B_MahJQJth5_3),.clk(gclk));
	jdff dff_B_3lrWq1ZZ2_3(.din(w_dff_B_MahJQJth5_3),.dout(w_dff_B_3lrWq1ZZ2_3),.clk(gclk));
	jdff dff_B_9VXUoVH00_3(.din(w_dff_B_3lrWq1ZZ2_3),.dout(w_dff_B_9VXUoVH00_3),.clk(gclk));
	jdff dff_B_D5Bx6L4k1_3(.din(w_dff_B_9VXUoVH00_3),.dout(w_dff_B_D5Bx6L4k1_3),.clk(gclk));
	jdff dff_B_XISZZfl35_3(.din(w_dff_B_D5Bx6L4k1_3),.dout(w_dff_B_XISZZfl35_3),.clk(gclk));
	jdff dff_B_LllyakdK2_3(.din(w_dff_B_XISZZfl35_3),.dout(w_dff_B_LllyakdK2_3),.clk(gclk));
	jdff dff_A_EIouoLnc5_0(.dout(w_n614_5[0]),.din(w_dff_A_EIouoLnc5_0),.clk(gclk));
	jdff dff_A_QGN3FYtA1_0(.dout(w_dff_A_EIouoLnc5_0),.din(w_dff_A_QGN3FYtA1_0),.clk(gclk));
	jdff dff_A_VPZDvZ3B7_0(.dout(w_dff_A_QGN3FYtA1_0),.din(w_dff_A_VPZDvZ3B7_0),.clk(gclk));
	jdff dff_A_tOSKmY9K7_0(.dout(w_dff_A_VPZDvZ3B7_0),.din(w_dff_A_tOSKmY9K7_0),.clk(gclk));
	jdff dff_A_tYyIqU8I4_0(.dout(w_dff_A_tOSKmY9K7_0),.din(w_dff_A_tYyIqU8I4_0),.clk(gclk));
	jdff dff_A_PednxCB11_0(.dout(w_dff_A_tYyIqU8I4_0),.din(w_dff_A_PednxCB11_0),.clk(gclk));
	jdff dff_A_yc5yqWwW4_0(.dout(w_dff_A_PednxCB11_0),.din(w_dff_A_yc5yqWwW4_0),.clk(gclk));
	jdff dff_A_nMsuSsbP8_0(.dout(w_dff_A_yc5yqWwW4_0),.din(w_dff_A_nMsuSsbP8_0),.clk(gclk));
	jdff dff_A_Rnhv3WZw1_0(.dout(w_dff_A_nMsuSsbP8_0),.din(w_dff_A_Rnhv3WZw1_0),.clk(gclk));
	jdff dff_A_uHCxWV2a9_0(.dout(w_dff_A_Rnhv3WZw1_0),.din(w_dff_A_uHCxWV2a9_0),.clk(gclk));
	jdff dff_A_pe4VyM901_0(.dout(w_n614_1[0]),.din(w_dff_A_pe4VyM901_0),.clk(gclk));
	jdff dff_A_ax2aeJKe0_0(.dout(w_dff_A_pe4VyM901_0),.din(w_dff_A_ax2aeJKe0_0),.clk(gclk));
	jdff dff_A_riJUsCaV4_2(.dout(w_n614_1[2]),.din(w_dff_A_riJUsCaV4_2),.clk(gclk));
	jdff dff_A_NtHf2mZN3_2(.dout(w_dff_A_riJUsCaV4_2),.din(w_dff_A_NtHf2mZN3_2),.clk(gclk));
	jdff dff_A_8c6wB8ym4_2(.dout(w_dff_A_NtHf2mZN3_2),.din(w_dff_A_8c6wB8ym4_2),.clk(gclk));
	jdff dff_A_fOXKGzIH2_2(.dout(w_dff_A_8c6wB8ym4_2),.din(w_dff_A_fOXKGzIH2_2),.clk(gclk));
	jdff dff_A_ZWk61n8A7_2(.dout(w_dff_A_fOXKGzIH2_2),.din(w_dff_A_ZWk61n8A7_2),.clk(gclk));
	jdff dff_A_NgFE8Z6K9_2(.dout(w_dff_A_ZWk61n8A7_2),.din(w_dff_A_NgFE8Z6K9_2),.clk(gclk));
	jdff dff_A_lWijELjg8_2(.dout(w_dff_A_NgFE8Z6K9_2),.din(w_dff_A_lWijELjg8_2),.clk(gclk));
	jdff dff_A_sucSOSwM4_2(.dout(w_dff_A_lWijELjg8_2),.din(w_dff_A_sucSOSwM4_2),.clk(gclk));
	jdff dff_A_gidrEGX38_2(.dout(w_dff_A_sucSOSwM4_2),.din(w_dff_A_gidrEGX38_2),.clk(gclk));
	jdff dff_A_2eUFjgy66_2(.dout(w_dff_A_gidrEGX38_2),.din(w_dff_A_2eUFjgy66_2),.clk(gclk));
	jdff dff_A_OF6GhCY34_2(.dout(w_dff_A_2eUFjgy66_2),.din(w_dff_A_OF6GhCY34_2),.clk(gclk));
	jdff dff_A_LJbc8UgO7_1(.dout(w_n614_0[1]),.din(w_dff_A_LJbc8UgO7_1),.clk(gclk));
	jdff dff_A_1ETxCsuV3_1(.dout(w_dff_A_LJbc8UgO7_1),.din(w_dff_A_1ETxCsuV3_1),.clk(gclk));
	jdff dff_A_L1rxmO587_1(.dout(w_dff_A_1ETxCsuV3_1),.din(w_dff_A_L1rxmO587_1),.clk(gclk));
	jdff dff_A_dRxpiVZy0_1(.dout(w_dff_A_L1rxmO587_1),.din(w_dff_A_dRxpiVZy0_1),.clk(gclk));
	jdff dff_A_X7aHFhnq1_1(.dout(w_dff_A_dRxpiVZy0_1),.din(w_dff_A_X7aHFhnq1_1),.clk(gclk));
	jdff dff_A_8v5wyk799_1(.dout(w_dff_A_X7aHFhnq1_1),.din(w_dff_A_8v5wyk799_1),.clk(gclk));
	jdff dff_A_TQSST8xv0_1(.dout(w_dff_A_8v5wyk799_1),.din(w_dff_A_TQSST8xv0_1),.clk(gclk));
	jdff dff_A_fp8UZbm02_2(.dout(w_n614_0[2]),.din(w_dff_A_fp8UZbm02_2),.clk(gclk));
	jdff dff_A_qshZv7hQ7_2(.dout(w_dff_A_fp8UZbm02_2),.din(w_dff_A_qshZv7hQ7_2),.clk(gclk));
	jdff dff_A_FcQcbM5U6_2(.dout(w_dff_A_qshZv7hQ7_2),.din(w_dff_A_FcQcbM5U6_2),.clk(gclk));
	jdff dff_A_fOMhSwhw7_2(.dout(w_dff_A_FcQcbM5U6_2),.din(w_dff_A_fOMhSwhw7_2),.clk(gclk));
	jdff dff_A_pMifdcYw3_2(.dout(w_dff_A_fOMhSwhw7_2),.din(w_dff_A_pMifdcYw3_2),.clk(gclk));
	jdff dff_A_9O5Nxu9W0_0(.dout(w_n613_1[0]),.din(w_dff_A_9O5Nxu9W0_0),.clk(gclk));
	jdff dff_A_eOOd4Wzs3_0(.dout(w_dff_A_9O5Nxu9W0_0),.din(w_dff_A_eOOd4Wzs3_0),.clk(gclk));
	jdff dff_A_sfT8hdn89_0(.dout(w_dff_A_eOOd4Wzs3_0),.din(w_dff_A_sfT8hdn89_0),.clk(gclk));
	jdff dff_A_AelXYhZ19_0(.dout(w_dff_A_sfT8hdn89_0),.din(w_dff_A_AelXYhZ19_0),.clk(gclk));
	jdff dff_A_s2AiT7Rh9_0(.dout(w_dff_A_AelXYhZ19_0),.din(w_dff_A_s2AiT7Rh9_0),.clk(gclk));
	jdff dff_A_8AQttcRs1_0(.dout(w_dff_A_s2AiT7Rh9_0),.din(w_dff_A_8AQttcRs1_0),.clk(gclk));
	jdff dff_A_NnUSno4B3_0(.dout(w_dff_A_8AQttcRs1_0),.din(w_dff_A_NnUSno4B3_0),.clk(gclk));
	jdff dff_A_n64U0nQk4_0(.dout(w_dff_A_NnUSno4B3_0),.din(w_dff_A_n64U0nQk4_0),.clk(gclk));
	jdff dff_A_OkecXknK2_0(.dout(w_dff_A_n64U0nQk4_0),.din(w_dff_A_OkecXknK2_0),.clk(gclk));
	jdff dff_A_TpMP28h14_0(.dout(w_dff_A_OkecXknK2_0),.din(w_dff_A_TpMP28h14_0),.clk(gclk));
	jdff dff_A_MyorrT4o6_0(.dout(w_dff_A_TpMP28h14_0),.din(w_dff_A_MyorrT4o6_0),.clk(gclk));
	jdff dff_A_6cth4LiG5_0(.dout(w_dff_A_MyorrT4o6_0),.din(w_dff_A_6cth4LiG5_0),.clk(gclk));
	jdff dff_A_5zyMBQ4e6_0(.dout(w_dff_A_6cth4LiG5_0),.din(w_dff_A_5zyMBQ4e6_0),.clk(gclk));
	jdff dff_A_WPwKHGLe3_0(.dout(w_dff_A_5zyMBQ4e6_0),.din(w_dff_A_WPwKHGLe3_0),.clk(gclk));
	jdff dff_A_aSvgI4nP6_1(.dout(w_n613_1[1]),.din(w_dff_A_aSvgI4nP6_1),.clk(gclk));
	jdff dff_A_tFYi5S421_1(.dout(w_dff_A_aSvgI4nP6_1),.din(w_dff_A_tFYi5S421_1),.clk(gclk));
	jdff dff_A_C23dacP67_1(.dout(w_dff_A_tFYi5S421_1),.din(w_dff_A_C23dacP67_1),.clk(gclk));
	jdff dff_A_x3oAx41T3_1(.dout(w_dff_A_C23dacP67_1),.din(w_dff_A_x3oAx41T3_1),.clk(gclk));
	jdff dff_A_DlW4a4Wk7_1(.dout(w_dff_A_x3oAx41T3_1),.din(w_dff_A_DlW4a4Wk7_1),.clk(gclk));
	jdff dff_A_r1h7pgr00_1(.dout(w_dff_A_DlW4a4Wk7_1),.din(w_dff_A_r1h7pgr00_1),.clk(gclk));
	jdff dff_A_eUW2J06r9_1(.dout(w_dff_A_r1h7pgr00_1),.din(w_dff_A_eUW2J06r9_1),.clk(gclk));
	jdff dff_A_9Coo9IHi9_1(.dout(w_dff_A_eUW2J06r9_1),.din(w_dff_A_9Coo9IHi9_1),.clk(gclk));
	jdff dff_A_GY1MIUoT5_1(.dout(w_dff_A_9Coo9IHi9_1),.din(w_dff_A_GY1MIUoT5_1),.clk(gclk));
	jdff dff_A_VaePAUu87_1(.dout(w_dff_A_GY1MIUoT5_1),.din(w_dff_A_VaePAUu87_1),.clk(gclk));
	jdff dff_A_iVqHq4Hr1_1(.dout(w_dff_A_VaePAUu87_1),.din(w_dff_A_iVqHq4Hr1_1),.clk(gclk));
	jdff dff_A_QF5aFoH61_1(.dout(w_dff_A_iVqHq4Hr1_1),.din(w_dff_A_QF5aFoH61_1),.clk(gclk));
	jdff dff_A_9VP9IOha1_1(.dout(w_dff_A_QF5aFoH61_1),.din(w_dff_A_9VP9IOha1_1),.clk(gclk));
	jdff dff_A_zKqqXszk4_1(.dout(w_dff_A_9VP9IOha1_1),.din(w_dff_A_zKqqXszk4_1),.clk(gclk));
	jdff dff_A_wuQD9Hzj0_1(.dout(w_n613_0[1]),.din(w_dff_A_wuQD9Hzj0_1),.clk(gclk));
	jdff dff_A_VIhe6DUA7_1(.dout(w_dff_A_wuQD9Hzj0_1),.din(w_dff_A_VIhe6DUA7_1),.clk(gclk));
	jdff dff_A_WbCy81H91_1(.dout(w_dff_A_VIhe6DUA7_1),.din(w_dff_A_WbCy81H91_1),.clk(gclk));
	jdff dff_A_V4OFxZ083_1(.dout(w_dff_A_WbCy81H91_1),.din(w_dff_A_V4OFxZ083_1),.clk(gclk));
	jdff dff_A_tkGJ9t5y6_1(.dout(w_dff_A_V4OFxZ083_1),.din(w_dff_A_tkGJ9t5y6_1),.clk(gclk));
	jdff dff_A_DQGtUc2l6_1(.dout(w_dff_A_tkGJ9t5y6_1),.din(w_dff_A_DQGtUc2l6_1),.clk(gclk));
	jdff dff_A_vfWf3gR25_1(.dout(w_dff_A_DQGtUc2l6_1),.din(w_dff_A_vfWf3gR25_1),.clk(gclk));
	jdff dff_A_nqPUHYk00_1(.dout(w_dff_A_vfWf3gR25_1),.din(w_dff_A_nqPUHYk00_1),.clk(gclk));
	jdff dff_A_x1s2U30T8_1(.dout(w_dff_A_nqPUHYk00_1),.din(w_dff_A_x1s2U30T8_1),.clk(gclk));
	jdff dff_A_CtcEoa8n2_1(.dout(w_dff_A_x1s2U30T8_1),.din(w_dff_A_CtcEoa8n2_1),.clk(gclk));
	jdff dff_A_v9xiFeg96_1(.dout(w_dff_A_CtcEoa8n2_1),.din(w_dff_A_v9xiFeg96_1),.clk(gclk));
	jdff dff_A_5C1hva4C5_1(.dout(w_dff_A_v9xiFeg96_1),.din(w_dff_A_5C1hva4C5_1),.clk(gclk));
	jdff dff_A_2x6djRsS9_1(.dout(w_dff_A_5C1hva4C5_1),.din(w_dff_A_2x6djRsS9_1),.clk(gclk));
	jdff dff_A_KoqiKnEX4_1(.dout(w_dff_A_2x6djRsS9_1),.din(w_dff_A_KoqiKnEX4_1),.clk(gclk));
	jdff dff_A_e63nU98t4_1(.dout(w_dff_A_KoqiKnEX4_1),.din(w_dff_A_e63nU98t4_1),.clk(gclk));
	jdff dff_A_kFe3LRGZ8_2(.dout(w_n613_0[2]),.din(w_dff_A_kFe3LRGZ8_2),.clk(gclk));
	jdff dff_A_wA86aAFS4_2(.dout(w_dff_A_kFe3LRGZ8_2),.din(w_dff_A_wA86aAFS4_2),.clk(gclk));
	jdff dff_A_d4rvyG4T9_2(.dout(w_dff_A_wA86aAFS4_2),.din(w_dff_A_d4rvyG4T9_2),.clk(gclk));
	jdff dff_A_0wVrAMwP3_2(.dout(w_dff_A_d4rvyG4T9_2),.din(w_dff_A_0wVrAMwP3_2),.clk(gclk));
	jdff dff_A_496hTPo42_2(.dout(w_dff_A_0wVrAMwP3_2),.din(w_dff_A_496hTPo42_2),.clk(gclk));
	jdff dff_A_fOGu7ZWA5_2(.dout(w_dff_A_496hTPo42_2),.din(w_dff_A_fOGu7ZWA5_2),.clk(gclk));
	jdff dff_A_0CweugFC8_2(.dout(w_dff_A_fOGu7ZWA5_2),.din(w_dff_A_0CweugFC8_2),.clk(gclk));
	jdff dff_A_4DpscUuV9_2(.dout(w_dff_A_0CweugFC8_2),.din(w_dff_A_4DpscUuV9_2),.clk(gclk));
	jdff dff_A_GsdaWvN54_2(.dout(w_dff_A_4DpscUuV9_2),.din(w_dff_A_GsdaWvN54_2),.clk(gclk));
	jdff dff_A_IHTSHDyC1_2(.dout(w_dff_A_GsdaWvN54_2),.din(w_dff_A_IHTSHDyC1_2),.clk(gclk));
	jdff dff_A_M8HdTe4Q8_2(.dout(w_dff_A_IHTSHDyC1_2),.din(w_dff_A_M8HdTe4Q8_2),.clk(gclk));
	jdff dff_A_VrYoCOTw7_2(.dout(w_dff_A_M8HdTe4Q8_2),.din(w_dff_A_VrYoCOTw7_2),.clk(gclk));
	jdff dff_A_AJeI4UoQ8_2(.dout(w_dff_A_VrYoCOTw7_2),.din(w_dff_A_AJeI4UoQ8_2),.clk(gclk));
	jdff dff_A_4G8okOjd0_2(.dout(w_dff_A_AJeI4UoQ8_2),.din(w_dff_A_4G8okOjd0_2),.clk(gclk));
	jdff dff_A_JXIXWcGo8_2(.dout(w_dff_A_4G8okOjd0_2),.din(w_dff_A_JXIXWcGo8_2),.clk(gclk));
	jdff dff_A_Rj63iQgT8_2(.dout(w_dff_A_JXIXWcGo8_2),.din(w_dff_A_Rj63iQgT8_2),.clk(gclk));
	jdff dff_A_qEGBsBzK4_2(.dout(w_dff_A_Rj63iQgT8_2),.din(w_dff_A_qEGBsBzK4_2),.clk(gclk));
	jdff dff_B_ZKL3QDgj6_3(.din(n613),.dout(w_dff_B_ZKL3QDgj6_3),.clk(gclk));
	jdff dff_A_egaZa6cr5_1(.dout(w_G45_0[1]),.din(w_dff_A_egaZa6cr5_1),.clk(gclk));
	jdff dff_A_JMvy7szU2_1(.dout(w_dff_A_egaZa6cr5_1),.din(w_dff_A_JMvy7szU2_1),.clk(gclk));
	jdff dff_A_aZAttY8G0_1(.dout(w_dff_A_JMvy7szU2_1),.din(w_dff_A_aZAttY8G0_1),.clk(gclk));
	jdff dff_A_6jCIhLww4_0(.dout(w_n151_2[0]),.din(w_dff_A_6jCIhLww4_0),.clk(gclk));
	jdff dff_A_XHe6xMWF4_2(.dout(w_n151_2[2]),.din(w_dff_A_XHe6xMWF4_2),.clk(gclk));
	jdff dff_A_0bioxm1z1_2(.dout(w_dff_A_XHe6xMWF4_2),.din(w_dff_A_0bioxm1z1_2),.clk(gclk));
	jdff dff_A_S8Ex2UsS9_0(.dout(w_G20_5[0]),.din(w_dff_A_S8Ex2UsS9_0),.clk(gclk));
	jdff dff_A_VsLbwrtO3_2(.dout(w_n142_0[2]),.din(w_dff_A_VsLbwrtO3_2),.clk(gclk));
	jdff dff_A_yAMMVBFC6_0(.dout(w_G1_1[0]),.din(w_dff_A_yAMMVBFC6_0),.clk(gclk));
	jdff dff_A_N5jP9i6U3_0(.dout(w_dff_A_yAMMVBFC6_0),.din(w_dff_A_N5jP9i6U3_0),.clk(gclk));
	jdff dff_A_qSKEbZh49_0(.dout(w_n604_2[0]),.din(w_dff_A_qSKEbZh49_0),.clk(gclk));
	jdff dff_A_H35nGzRP5_0(.dout(w_dff_A_qSKEbZh49_0),.din(w_dff_A_H35nGzRP5_0),.clk(gclk));
	jdff dff_A_aI1RUtP61_0(.dout(w_dff_A_H35nGzRP5_0),.din(w_dff_A_aI1RUtP61_0),.clk(gclk));
	jdff dff_A_F7ERN3hQ1_0(.dout(w_dff_A_aI1RUtP61_0),.din(w_dff_A_F7ERN3hQ1_0),.clk(gclk));
	jdff dff_A_iVRRV7Sw1_0(.dout(w_dff_A_F7ERN3hQ1_0),.din(w_dff_A_iVRRV7Sw1_0),.clk(gclk));
	jdff dff_A_cWYLC7ju0_0(.dout(w_dff_A_iVRRV7Sw1_0),.din(w_dff_A_cWYLC7ju0_0),.clk(gclk));
	jdff dff_A_ywYiSN8k3_0(.dout(w_dff_A_cWYLC7ju0_0),.din(w_dff_A_ywYiSN8k3_0),.clk(gclk));
	jdff dff_A_YTEdMcQC8_0(.dout(w_dff_A_ywYiSN8k3_0),.din(w_dff_A_YTEdMcQC8_0),.clk(gclk));
	jdff dff_A_wEp1EegM7_0(.dout(w_dff_A_YTEdMcQC8_0),.din(w_dff_A_wEp1EegM7_0),.clk(gclk));
	jdff dff_A_AX1G0bb44_0(.dout(w_dff_A_wEp1EegM7_0),.din(w_dff_A_AX1G0bb44_0),.clk(gclk));
	jdff dff_A_1qPTpA1q6_0(.dout(w_dff_A_AX1G0bb44_0),.din(w_dff_A_1qPTpA1q6_0),.clk(gclk));
	jdff dff_A_79mn2xNf3_0(.dout(w_dff_A_1qPTpA1q6_0),.din(w_dff_A_79mn2xNf3_0),.clk(gclk));
	jdff dff_A_HDp4Rv4b7_0(.dout(w_dff_A_79mn2xNf3_0),.din(w_dff_A_HDp4Rv4b7_0),.clk(gclk));
	jdff dff_A_InXusHiD4_0(.dout(w_dff_A_HDp4Rv4b7_0),.din(w_dff_A_InXusHiD4_0),.clk(gclk));
	jdff dff_A_2J4xUV9f5_0(.dout(w_n604_0[0]),.din(w_dff_A_2J4xUV9f5_0),.clk(gclk));
	jdff dff_A_wmUZLzCh4_0(.dout(w_dff_A_2J4xUV9f5_0),.din(w_dff_A_wmUZLzCh4_0),.clk(gclk));
	jdff dff_A_p3nTqZD10_0(.dout(w_dff_A_wmUZLzCh4_0),.din(w_dff_A_p3nTqZD10_0),.clk(gclk));
	jdff dff_A_wQHYfsYp4_0(.dout(w_dff_A_p3nTqZD10_0),.din(w_dff_A_wQHYfsYp4_0),.clk(gclk));
	jdff dff_A_RHuUdByJ7_0(.dout(w_dff_A_wQHYfsYp4_0),.din(w_dff_A_RHuUdByJ7_0),.clk(gclk));
	jdff dff_A_Abwx3fK25_0(.dout(w_dff_A_RHuUdByJ7_0),.din(w_dff_A_Abwx3fK25_0),.clk(gclk));
	jdff dff_A_taupPDeH9_0(.dout(w_dff_A_Abwx3fK25_0),.din(w_dff_A_taupPDeH9_0),.clk(gclk));
	jdff dff_A_Tszw1cSD1_0(.dout(w_dff_A_taupPDeH9_0),.din(w_dff_A_Tszw1cSD1_0),.clk(gclk));
	jdff dff_A_96EuYVYl3_0(.dout(w_dff_A_Tszw1cSD1_0),.din(w_dff_A_96EuYVYl3_0),.clk(gclk));
	jdff dff_A_WDZpszBJ8_0(.dout(w_dff_A_96EuYVYl3_0),.din(w_dff_A_WDZpszBJ8_0),.clk(gclk));
	jdff dff_A_1aQXot4l1_0(.dout(w_dff_A_WDZpszBJ8_0),.din(w_dff_A_1aQXot4l1_0),.clk(gclk));
	jdff dff_A_61jEzgoa0_0(.dout(w_dff_A_1aQXot4l1_0),.din(w_dff_A_61jEzgoa0_0),.clk(gclk));
	jdff dff_A_PUd3i7Rp2_0(.dout(w_dff_A_61jEzgoa0_0),.din(w_dff_A_PUd3i7Rp2_0),.clk(gclk));
	jdff dff_A_0NHp2NW70_0(.dout(w_dff_A_PUd3i7Rp2_0),.din(w_dff_A_0NHp2NW70_0),.clk(gclk));
	jdff dff_A_3cnhfRbG6_2(.dout(w_n604_0[2]),.din(w_dff_A_3cnhfRbG6_2),.clk(gclk));
	jdff dff_A_2noCDfoW2_2(.dout(w_dff_A_3cnhfRbG6_2),.din(w_dff_A_2noCDfoW2_2),.clk(gclk));
	jdff dff_A_NQJiFtDC4_2(.dout(w_dff_A_2noCDfoW2_2),.din(w_dff_A_NQJiFtDC4_2),.clk(gclk));
	jdff dff_A_j50Xlt662_2(.dout(w_dff_A_NQJiFtDC4_2),.din(w_dff_A_j50Xlt662_2),.clk(gclk));
	jdff dff_A_hTCvXI2g6_2(.dout(w_dff_A_j50Xlt662_2),.din(w_dff_A_hTCvXI2g6_2),.clk(gclk));
	jdff dff_A_N1HLg4Qb8_2(.dout(w_dff_A_hTCvXI2g6_2),.din(w_dff_A_N1HLg4Qb8_2),.clk(gclk));
	jdff dff_A_isP7eMnG7_2(.dout(w_dff_A_N1HLg4Qb8_2),.din(w_dff_A_isP7eMnG7_2),.clk(gclk));
	jdff dff_A_G9GbJgRh8_2(.dout(w_dff_A_isP7eMnG7_2),.din(w_dff_A_G9GbJgRh8_2),.clk(gclk));
	jdff dff_A_obwNyN3M3_2(.dout(w_dff_A_G9GbJgRh8_2),.din(w_dff_A_obwNyN3M3_2),.clk(gclk));
	jdff dff_A_dUxOj9k29_2(.dout(w_dff_A_obwNyN3M3_2),.din(w_dff_A_dUxOj9k29_2),.clk(gclk));
	jdff dff_A_dyi1Gi8L2_2(.dout(w_dff_A_dUxOj9k29_2),.din(w_dff_A_dyi1Gi8L2_2),.clk(gclk));
	jdff dff_A_ezUndS1G2_2(.dout(w_dff_A_dyi1Gi8L2_2),.din(w_dff_A_ezUndS1G2_2),.clk(gclk));
	jdff dff_A_XeLfyT332_2(.dout(w_dff_A_ezUndS1G2_2),.din(w_dff_A_XeLfyT332_2),.clk(gclk));
	jdff dff_A_4RapG7jq9_2(.dout(w_dff_A_XeLfyT332_2),.din(w_dff_A_4RapG7jq9_2),.clk(gclk));
	jdff dff_A_wDowTD480_2(.dout(w_dff_A_4RapG7jq9_2),.din(w_dff_A_wDowTD480_2),.clk(gclk));
	jdff dff_A_guTVlD6N5_2(.dout(w_dff_A_wDowTD480_2),.din(w_dff_A_guTVlD6N5_2),.clk(gclk));
	jdff dff_A_e3s8cSwM6_0(.dout(w_G13_2[0]),.din(w_dff_A_e3s8cSwM6_0),.clk(gclk));
	jdff dff_A_aAR6pYCz9_1(.dout(w_G1_2[1]),.din(w_dff_A_aAR6pYCz9_1),.clk(gclk));
	jdff dff_A_NOPU9yVk7_2(.dout(w_G1_0[2]),.din(w_dff_A_NOPU9yVk7_2),.clk(gclk));
	jdff dff_A_5tQGUpOt2_2(.dout(w_dff_A_NOPU9yVk7_2),.din(w_dff_A_5tQGUpOt2_2),.clk(gclk));
	jdff dff_A_rq0kkRTd8_2(.dout(w_dff_A_5tQGUpOt2_2),.din(w_dff_A_rq0kkRTd8_2),.clk(gclk));
	jdff dff_A_Z3J2hJSb1_2(.dout(w_dff_A_rq0kkRTd8_2),.din(w_dff_A_Z3J2hJSb1_2),.clk(gclk));
	jdff dff_A_8ZETPY5M4_0(.dout(w_G20_6[0]),.din(w_dff_A_8ZETPY5M4_0),.clk(gclk));
	jdff dff_A_4naE8Tex9_0(.dout(w_dff_A_8ZETPY5M4_0),.din(w_dff_A_4naE8Tex9_0),.clk(gclk));
	jdff dff_A_K1JJceJN9_2(.dout(w_G20_6[2]),.din(w_dff_A_K1JJceJN9_2),.clk(gclk));
	jdff dff_A_WDaLdjET0_2(.dout(w_dff_A_K1JJceJN9_2),.din(w_dff_A_WDaLdjET0_2),.clk(gclk));
	jdff dff_A_umfdCvHV8_0(.dout(w_G20_1[0]),.din(w_dff_A_umfdCvHV8_0),.clk(gclk));
	jdff dff_A_4X5ktXLG6_2(.dout(w_G20_0[2]),.din(w_dff_A_4X5ktXLG6_2),.clk(gclk));
	jdff dff_A_kTSf2yCF4_1(.dout(w_n163_0[1]),.din(w_dff_A_kTSf2yCF4_1),.clk(gclk));
	jdff dff_A_qD6GtDDf0_1(.dout(w_dff_A_kTSf2yCF4_1),.din(w_dff_A_qD6GtDDf0_1),.clk(gclk));
	jdff dff_A_skFdznOb0_1(.dout(w_dff_A_qD6GtDDf0_1),.din(w_dff_A_skFdznOb0_1),.clk(gclk));
	jdff dff_A_xir4isHr5_1(.dout(w_dff_A_skFdznOb0_1),.din(w_dff_A_xir4isHr5_1),.clk(gclk));
	jdff dff_A_jkhOXIw50_1(.dout(w_dff_A_xir4isHr5_1),.din(w_dff_A_jkhOXIw50_1),.clk(gclk));
	jdff dff_A_4vkk07dQ3_1(.dout(w_dff_A_jkhOXIw50_1),.din(w_dff_A_4vkk07dQ3_1),.clk(gclk));
	jdff dff_A_T1y13SqN0_1(.dout(w_dff_A_4vkk07dQ3_1),.din(w_dff_A_T1y13SqN0_1),.clk(gclk));
	jdff dff_A_DGZgzgEp6_1(.dout(w_dff_A_T1y13SqN0_1),.din(w_dff_A_DGZgzgEp6_1),.clk(gclk));
	jdff dff_A_cY9hvLqp3_1(.dout(w_dff_A_DGZgzgEp6_1),.din(w_dff_A_cY9hvLqp3_1),.clk(gclk));
	jdff dff_A_RBGcIbgw2_1(.dout(w_dff_A_cY9hvLqp3_1),.din(w_dff_A_RBGcIbgw2_1),.clk(gclk));
	jdff dff_A_Ug09h26b1_1(.dout(w_dff_A_RBGcIbgw2_1),.din(w_dff_A_Ug09h26b1_1),.clk(gclk));
	jdff dff_A_nTFcBRwC5_2(.dout(w_n163_0[2]),.din(w_dff_A_nTFcBRwC5_2),.clk(gclk));
	jdff dff_A_jIXxqQBl5_2(.dout(w_dff_A_nTFcBRwC5_2),.din(w_dff_A_jIXxqQBl5_2),.clk(gclk));
	jdff dff_A_Ai93AJFG8_2(.dout(w_dff_A_8wK8UJoV2_0),.din(w_dff_A_Ai93AJFG8_2),.clk(gclk));
	jdff dff_A_8wK8UJoV2_0(.dout(w_dff_A_6BjZhAeX9_0),.din(w_dff_A_8wK8UJoV2_0),.clk(gclk));
	jdff dff_A_6BjZhAeX9_0(.dout(w_dff_A_S5KM9Trm0_0),.din(w_dff_A_6BjZhAeX9_0),.clk(gclk));
	jdff dff_A_S5KM9Trm0_0(.dout(w_dff_A_c8gsiFJd5_0),.din(w_dff_A_S5KM9Trm0_0),.clk(gclk));
	jdff dff_A_c8gsiFJd5_0(.dout(w_dff_A_SOvO5oUh8_0),.din(w_dff_A_c8gsiFJd5_0),.clk(gclk));
	jdff dff_A_SOvO5oUh8_0(.dout(w_dff_A_tz7QtjWd6_0),.din(w_dff_A_SOvO5oUh8_0),.clk(gclk));
	jdff dff_A_tz7QtjWd6_0(.dout(w_dff_A_AVbjljYj0_0),.din(w_dff_A_tz7QtjWd6_0),.clk(gclk));
	jdff dff_A_AVbjljYj0_0(.dout(w_dff_A_bzLOMo5p2_0),.din(w_dff_A_AVbjljYj0_0),.clk(gclk));
	jdff dff_A_bzLOMo5p2_0(.dout(w_dff_A_EuImGtAL1_0),.din(w_dff_A_bzLOMo5p2_0),.clk(gclk));
	jdff dff_A_EuImGtAL1_0(.dout(w_dff_A_il6Dvlg90_0),.din(w_dff_A_EuImGtAL1_0),.clk(gclk));
	jdff dff_A_il6Dvlg90_0(.dout(w_dff_A_ICHD9OEJ4_0),.din(w_dff_A_il6Dvlg90_0),.clk(gclk));
	jdff dff_A_ICHD9OEJ4_0(.dout(w_dff_A_ugjitDbz9_0),.din(w_dff_A_ICHD9OEJ4_0),.clk(gclk));
	jdff dff_A_ugjitDbz9_0(.dout(w_dff_A_Vpq56JlK0_0),.din(w_dff_A_ugjitDbz9_0),.clk(gclk));
	jdff dff_A_Vpq56JlK0_0(.dout(w_dff_A_MFrcOJQK7_0),.din(w_dff_A_Vpq56JlK0_0),.clk(gclk));
	jdff dff_A_MFrcOJQK7_0(.dout(w_dff_A_jn2ogL1S9_0),.din(w_dff_A_MFrcOJQK7_0),.clk(gclk));
	jdff dff_A_jn2ogL1S9_0(.dout(w_dff_A_bC1ONhvq0_0),.din(w_dff_A_jn2ogL1S9_0),.clk(gclk));
	jdff dff_A_bC1ONhvq0_0(.dout(w_dff_A_USFsF0Q75_0),.din(w_dff_A_bC1ONhvq0_0),.clk(gclk));
	jdff dff_A_USFsF0Q75_0(.dout(w_dff_A_eOJ13Mva0_0),.din(w_dff_A_USFsF0Q75_0),.clk(gclk));
	jdff dff_A_eOJ13Mva0_0(.dout(w_dff_A_Q01RmBgn9_0),.din(w_dff_A_eOJ13Mva0_0),.clk(gclk));
	jdff dff_A_Q01RmBgn9_0(.dout(w_dff_A_QyRcSd7n2_0),.din(w_dff_A_Q01RmBgn9_0),.clk(gclk));
	jdff dff_A_QyRcSd7n2_0(.dout(w_dff_A_jOVPISwb2_0),.din(w_dff_A_QyRcSd7n2_0),.clk(gclk));
	jdff dff_A_jOVPISwb2_0(.dout(w_dff_A_IRyFOeZM1_0),.din(w_dff_A_jOVPISwb2_0),.clk(gclk));
	jdff dff_A_IRyFOeZM1_0(.dout(w_dff_A_xiulzJwB2_0),.din(w_dff_A_IRyFOeZM1_0),.clk(gclk));
	jdff dff_A_xiulzJwB2_0(.dout(w_dff_A_3NHEjUHK0_0),.din(w_dff_A_xiulzJwB2_0),.clk(gclk));
	jdff dff_A_3NHEjUHK0_0(.dout(w_dff_A_E6yqJQNg3_0),.din(w_dff_A_3NHEjUHK0_0),.clk(gclk));
	jdff dff_A_E6yqJQNg3_0(.dout(w_dff_A_kWSj6xz52_0),.din(w_dff_A_E6yqJQNg3_0),.clk(gclk));
	jdff dff_A_kWSj6xz52_0(.dout(G353),.din(w_dff_A_kWSj6xz52_0),.clk(gclk));
	jdff dff_A_heHbqSsj6_1(.dout(w_dff_A_6FpreaDL9_0),.din(w_dff_A_heHbqSsj6_1),.clk(gclk));
	jdff dff_A_6FpreaDL9_0(.dout(w_dff_A_oBlulQxO4_0),.din(w_dff_A_6FpreaDL9_0),.clk(gclk));
	jdff dff_A_oBlulQxO4_0(.dout(w_dff_A_zSHMdOlg5_0),.din(w_dff_A_oBlulQxO4_0),.clk(gclk));
	jdff dff_A_zSHMdOlg5_0(.dout(w_dff_A_3ouQPzKh8_0),.din(w_dff_A_zSHMdOlg5_0),.clk(gclk));
	jdff dff_A_3ouQPzKh8_0(.dout(w_dff_A_4Z0zJ60r3_0),.din(w_dff_A_3ouQPzKh8_0),.clk(gclk));
	jdff dff_A_4Z0zJ60r3_0(.dout(w_dff_A_BM61Geu76_0),.din(w_dff_A_4Z0zJ60r3_0),.clk(gclk));
	jdff dff_A_BM61Geu76_0(.dout(w_dff_A_P98P93Vo1_0),.din(w_dff_A_BM61Geu76_0),.clk(gclk));
	jdff dff_A_P98P93Vo1_0(.dout(w_dff_A_1bFkcBog0_0),.din(w_dff_A_P98P93Vo1_0),.clk(gclk));
	jdff dff_A_1bFkcBog0_0(.dout(w_dff_A_C5vjGe879_0),.din(w_dff_A_1bFkcBog0_0),.clk(gclk));
	jdff dff_A_C5vjGe879_0(.dout(w_dff_A_fxx806kt2_0),.din(w_dff_A_C5vjGe879_0),.clk(gclk));
	jdff dff_A_fxx806kt2_0(.dout(w_dff_A_nRxvoZy43_0),.din(w_dff_A_fxx806kt2_0),.clk(gclk));
	jdff dff_A_nRxvoZy43_0(.dout(w_dff_A_T1Ru8qFm5_0),.din(w_dff_A_nRxvoZy43_0),.clk(gclk));
	jdff dff_A_T1Ru8qFm5_0(.dout(w_dff_A_ZTSJahtc0_0),.din(w_dff_A_T1Ru8qFm5_0),.clk(gclk));
	jdff dff_A_ZTSJahtc0_0(.dout(w_dff_A_CqozIHur5_0),.din(w_dff_A_ZTSJahtc0_0),.clk(gclk));
	jdff dff_A_CqozIHur5_0(.dout(w_dff_A_VQDCUjM34_0),.din(w_dff_A_CqozIHur5_0),.clk(gclk));
	jdff dff_A_VQDCUjM34_0(.dout(w_dff_A_O3bEJz710_0),.din(w_dff_A_VQDCUjM34_0),.clk(gclk));
	jdff dff_A_O3bEJz710_0(.dout(w_dff_A_1GVJ6AsH9_0),.din(w_dff_A_O3bEJz710_0),.clk(gclk));
	jdff dff_A_1GVJ6AsH9_0(.dout(w_dff_A_N0on1wpE3_0),.din(w_dff_A_1GVJ6AsH9_0),.clk(gclk));
	jdff dff_A_N0on1wpE3_0(.dout(w_dff_A_mknWWI8a5_0),.din(w_dff_A_N0on1wpE3_0),.clk(gclk));
	jdff dff_A_mknWWI8a5_0(.dout(w_dff_A_7zuE67D02_0),.din(w_dff_A_mknWWI8a5_0),.clk(gclk));
	jdff dff_A_7zuE67D02_0(.dout(w_dff_A_rmUqLk1b0_0),.din(w_dff_A_7zuE67D02_0),.clk(gclk));
	jdff dff_A_rmUqLk1b0_0(.dout(w_dff_A_p1L3MV9H0_0),.din(w_dff_A_rmUqLk1b0_0),.clk(gclk));
	jdff dff_A_p1L3MV9H0_0(.dout(w_dff_A_WhhtPLAe0_0),.din(w_dff_A_p1L3MV9H0_0),.clk(gclk));
	jdff dff_A_WhhtPLAe0_0(.dout(w_dff_A_8mTF0rtj6_0),.din(w_dff_A_WhhtPLAe0_0),.clk(gclk));
	jdff dff_A_8mTF0rtj6_0(.dout(w_dff_A_mE5NcZom7_0),.din(w_dff_A_8mTF0rtj6_0),.clk(gclk));
	jdff dff_A_mE5NcZom7_0(.dout(w_dff_A_09oKH6DA8_0),.din(w_dff_A_mE5NcZom7_0),.clk(gclk));
	jdff dff_A_09oKH6DA8_0(.dout(w_dff_A_MhNMV9bW1_0),.din(w_dff_A_09oKH6DA8_0),.clk(gclk));
	jdff dff_A_MhNMV9bW1_0(.dout(G355),.din(w_dff_A_MhNMV9bW1_0),.clk(gclk));
	jdff dff_A_dcDQDPxH8_2(.dout(w_dff_A_2JWF9wm07_0),.din(w_dff_A_dcDQDPxH8_2),.clk(gclk));
	jdff dff_A_2JWF9wm07_0(.dout(w_dff_A_eOMG95CX1_0),.din(w_dff_A_2JWF9wm07_0),.clk(gclk));
	jdff dff_A_eOMG95CX1_0(.dout(w_dff_A_2tAQ40B94_0),.din(w_dff_A_eOMG95CX1_0),.clk(gclk));
	jdff dff_A_2tAQ40B94_0(.dout(w_dff_A_k3cg0RrP9_0),.din(w_dff_A_2tAQ40B94_0),.clk(gclk));
	jdff dff_A_k3cg0RrP9_0(.dout(w_dff_A_OKX3pUMK6_0),.din(w_dff_A_k3cg0RrP9_0),.clk(gclk));
	jdff dff_A_OKX3pUMK6_0(.dout(w_dff_A_8qzrIc9S6_0),.din(w_dff_A_OKX3pUMK6_0),.clk(gclk));
	jdff dff_A_8qzrIc9S6_0(.dout(w_dff_A_zWpc0EmV8_0),.din(w_dff_A_8qzrIc9S6_0),.clk(gclk));
	jdff dff_A_zWpc0EmV8_0(.dout(w_dff_A_xeiXKon84_0),.din(w_dff_A_zWpc0EmV8_0),.clk(gclk));
	jdff dff_A_xeiXKon84_0(.dout(w_dff_A_WMmrDgGo0_0),.din(w_dff_A_xeiXKon84_0),.clk(gclk));
	jdff dff_A_WMmrDgGo0_0(.dout(w_dff_A_fXDVISIz7_0),.din(w_dff_A_WMmrDgGo0_0),.clk(gclk));
	jdff dff_A_fXDVISIz7_0(.dout(w_dff_A_5KRr7hOJ1_0),.din(w_dff_A_fXDVISIz7_0),.clk(gclk));
	jdff dff_A_5KRr7hOJ1_0(.dout(w_dff_A_wNyduM9r0_0),.din(w_dff_A_5KRr7hOJ1_0),.clk(gclk));
	jdff dff_A_wNyduM9r0_0(.dout(w_dff_A_TWoDI0xq5_0),.din(w_dff_A_wNyduM9r0_0),.clk(gclk));
	jdff dff_A_TWoDI0xq5_0(.dout(w_dff_A_mVa35RVi0_0),.din(w_dff_A_TWoDI0xq5_0),.clk(gclk));
	jdff dff_A_mVa35RVi0_0(.dout(w_dff_A_5iZI7iGb1_0),.din(w_dff_A_mVa35RVi0_0),.clk(gclk));
	jdff dff_A_5iZI7iGb1_0(.dout(w_dff_A_MLO4bTuK9_0),.din(w_dff_A_5iZI7iGb1_0),.clk(gclk));
	jdff dff_A_MLO4bTuK9_0(.dout(w_dff_A_eylU7JFY2_0),.din(w_dff_A_MLO4bTuK9_0),.clk(gclk));
	jdff dff_A_eylU7JFY2_0(.dout(w_dff_A_SJifkAxx4_0),.din(w_dff_A_eylU7JFY2_0),.clk(gclk));
	jdff dff_A_SJifkAxx4_0(.dout(w_dff_A_ADLAh3eJ8_0),.din(w_dff_A_SJifkAxx4_0),.clk(gclk));
	jdff dff_A_ADLAh3eJ8_0(.dout(w_dff_A_MiEXD3jG9_0),.din(w_dff_A_ADLAh3eJ8_0),.clk(gclk));
	jdff dff_A_MiEXD3jG9_0(.dout(w_dff_A_S8FkLZxb3_0),.din(w_dff_A_MiEXD3jG9_0),.clk(gclk));
	jdff dff_A_S8FkLZxb3_0(.dout(w_dff_A_1F2vq7cY6_0),.din(w_dff_A_S8FkLZxb3_0),.clk(gclk));
	jdff dff_A_1F2vq7cY6_0(.dout(G361),.din(w_dff_A_1F2vq7cY6_0),.clk(gclk));
	jdff dff_A_LguSs9EC9_2(.dout(w_dff_A_CFNiCZF28_0),.din(w_dff_A_LguSs9EC9_2),.clk(gclk));
	jdff dff_A_CFNiCZF28_0(.dout(w_dff_A_SxW2B5cl0_0),.din(w_dff_A_CFNiCZF28_0),.clk(gclk));
	jdff dff_A_SxW2B5cl0_0(.dout(w_dff_A_viKuLYhm9_0),.din(w_dff_A_SxW2B5cl0_0),.clk(gclk));
	jdff dff_A_viKuLYhm9_0(.dout(w_dff_A_cK1OG4ZC5_0),.din(w_dff_A_viKuLYhm9_0),.clk(gclk));
	jdff dff_A_cK1OG4ZC5_0(.dout(w_dff_A_mRQio0LQ0_0),.din(w_dff_A_cK1OG4ZC5_0),.clk(gclk));
	jdff dff_A_mRQio0LQ0_0(.dout(w_dff_A_6xS7V23c1_0),.din(w_dff_A_mRQio0LQ0_0),.clk(gclk));
	jdff dff_A_6xS7V23c1_0(.dout(w_dff_A_dHku9i8q2_0),.din(w_dff_A_6xS7V23c1_0),.clk(gclk));
	jdff dff_A_dHku9i8q2_0(.dout(w_dff_A_qUW0RoQM1_0),.din(w_dff_A_dHku9i8q2_0),.clk(gclk));
	jdff dff_A_qUW0RoQM1_0(.dout(w_dff_A_Nihax5y29_0),.din(w_dff_A_qUW0RoQM1_0),.clk(gclk));
	jdff dff_A_Nihax5y29_0(.dout(w_dff_A_UAe7Fu759_0),.din(w_dff_A_Nihax5y29_0),.clk(gclk));
	jdff dff_A_UAe7Fu759_0(.dout(w_dff_A_vqd355fq0_0),.din(w_dff_A_UAe7Fu759_0),.clk(gclk));
	jdff dff_A_vqd355fq0_0(.dout(w_dff_A_fhGLWfSZ6_0),.din(w_dff_A_vqd355fq0_0),.clk(gclk));
	jdff dff_A_fhGLWfSZ6_0(.dout(w_dff_A_AGd7AVLH3_0),.din(w_dff_A_fhGLWfSZ6_0),.clk(gclk));
	jdff dff_A_AGd7AVLH3_0(.dout(w_dff_A_uzyAGsou2_0),.din(w_dff_A_AGd7AVLH3_0),.clk(gclk));
	jdff dff_A_uzyAGsou2_0(.dout(w_dff_A_VyaPxz1f2_0),.din(w_dff_A_uzyAGsou2_0),.clk(gclk));
	jdff dff_A_VyaPxz1f2_0(.dout(w_dff_A_8RHrabNL8_0),.din(w_dff_A_VyaPxz1f2_0),.clk(gclk));
	jdff dff_A_8RHrabNL8_0(.dout(w_dff_A_UFIMXzq03_0),.din(w_dff_A_8RHrabNL8_0),.clk(gclk));
	jdff dff_A_UFIMXzq03_0(.dout(w_dff_A_RToiNRdE6_0),.din(w_dff_A_UFIMXzq03_0),.clk(gclk));
	jdff dff_A_RToiNRdE6_0(.dout(w_dff_A_mvxanOFS4_0),.din(w_dff_A_RToiNRdE6_0),.clk(gclk));
	jdff dff_A_mvxanOFS4_0(.dout(w_dff_A_Y3Md220M2_0),.din(w_dff_A_mvxanOFS4_0),.clk(gclk));
	jdff dff_A_Y3Md220M2_0(.dout(w_dff_A_K9ynOQIK4_0),.din(w_dff_A_Y3Md220M2_0),.clk(gclk));
	jdff dff_A_K9ynOQIK4_0(.dout(w_dff_A_qRv3Kthb3_0),.din(w_dff_A_K9ynOQIK4_0),.clk(gclk));
	jdff dff_A_qRv3Kthb3_0(.dout(w_dff_A_QrDGQSQd8_0),.din(w_dff_A_qRv3Kthb3_0),.clk(gclk));
	jdff dff_A_QrDGQSQd8_0(.dout(w_dff_A_qiXxe7Fc9_0),.din(w_dff_A_QrDGQSQd8_0),.clk(gclk));
	jdff dff_A_qiXxe7Fc9_0(.dout(w_dff_A_q1pa0OsA6_0),.din(w_dff_A_qiXxe7Fc9_0),.clk(gclk));
	jdff dff_A_q1pa0OsA6_0(.dout(G358),.din(w_dff_A_q1pa0OsA6_0),.clk(gclk));
	jdff dff_A_jxO7Gb1E1_2(.dout(w_dff_A_2lCTvU9h2_0),.din(w_dff_A_jxO7Gb1E1_2),.clk(gclk));
	jdff dff_A_2lCTvU9h2_0(.dout(w_dff_A_sMhKaenh0_0),.din(w_dff_A_2lCTvU9h2_0),.clk(gclk));
	jdff dff_A_sMhKaenh0_0(.dout(w_dff_A_tJd3NBRk9_0),.din(w_dff_A_sMhKaenh0_0),.clk(gclk));
	jdff dff_A_tJd3NBRk9_0(.dout(w_dff_A_k5TFpQE33_0),.din(w_dff_A_tJd3NBRk9_0),.clk(gclk));
	jdff dff_A_k5TFpQE33_0(.dout(w_dff_A_qjN0MhyM1_0),.din(w_dff_A_k5TFpQE33_0),.clk(gclk));
	jdff dff_A_qjN0MhyM1_0(.dout(w_dff_A_8mzykBEF3_0),.din(w_dff_A_qjN0MhyM1_0),.clk(gclk));
	jdff dff_A_8mzykBEF3_0(.dout(w_dff_A_O5cozlGr7_0),.din(w_dff_A_8mzykBEF3_0),.clk(gclk));
	jdff dff_A_O5cozlGr7_0(.dout(w_dff_A_kMvDyWg85_0),.din(w_dff_A_O5cozlGr7_0),.clk(gclk));
	jdff dff_A_kMvDyWg85_0(.dout(w_dff_A_xGH5Ivs95_0),.din(w_dff_A_kMvDyWg85_0),.clk(gclk));
	jdff dff_A_xGH5Ivs95_0(.dout(w_dff_A_ueyEnQai1_0),.din(w_dff_A_xGH5Ivs95_0),.clk(gclk));
	jdff dff_A_ueyEnQai1_0(.dout(w_dff_A_1csAG2rb0_0),.din(w_dff_A_ueyEnQai1_0),.clk(gclk));
	jdff dff_A_1csAG2rb0_0(.dout(w_dff_A_YmqN1DgV8_0),.din(w_dff_A_1csAG2rb0_0),.clk(gclk));
	jdff dff_A_YmqN1DgV8_0(.dout(w_dff_A_Ojk52XmW4_0),.din(w_dff_A_YmqN1DgV8_0),.clk(gclk));
	jdff dff_A_Ojk52XmW4_0(.dout(w_dff_A_j1ky04Bg4_0),.din(w_dff_A_Ojk52XmW4_0),.clk(gclk));
	jdff dff_A_j1ky04Bg4_0(.dout(w_dff_A_AJaRT1qj2_0),.din(w_dff_A_j1ky04Bg4_0),.clk(gclk));
	jdff dff_A_AJaRT1qj2_0(.dout(w_dff_A_QmxGzTpy0_0),.din(w_dff_A_AJaRT1qj2_0),.clk(gclk));
	jdff dff_A_QmxGzTpy0_0(.dout(w_dff_A_HdJhXA425_0),.din(w_dff_A_QmxGzTpy0_0),.clk(gclk));
	jdff dff_A_HdJhXA425_0(.dout(w_dff_A_MoOazLC59_0),.din(w_dff_A_HdJhXA425_0),.clk(gclk));
	jdff dff_A_MoOazLC59_0(.dout(w_dff_A_946hA4991_0),.din(w_dff_A_MoOazLC59_0),.clk(gclk));
	jdff dff_A_946hA4991_0(.dout(w_dff_A_9FAkzqTC5_0),.din(w_dff_A_946hA4991_0),.clk(gclk));
	jdff dff_A_9FAkzqTC5_0(.dout(w_dff_A_qP85N9KR9_0),.din(w_dff_A_9FAkzqTC5_0),.clk(gclk));
	jdff dff_A_qP85N9KR9_0(.dout(w_dff_A_Cq8yWShR4_0),.din(w_dff_A_qP85N9KR9_0),.clk(gclk));
	jdff dff_A_Cq8yWShR4_0(.dout(w_dff_A_meWnGMiq9_0),.din(w_dff_A_Cq8yWShR4_0),.clk(gclk));
	jdff dff_A_meWnGMiq9_0(.dout(w_dff_A_cmSYvPGX9_0),.din(w_dff_A_meWnGMiq9_0),.clk(gclk));
	jdff dff_A_cmSYvPGX9_0(.dout(w_dff_A_HbUE7IYu9_0),.din(w_dff_A_cmSYvPGX9_0),.clk(gclk));
	jdff dff_A_HbUE7IYu9_0(.dout(w_dff_A_HJpBciPx2_0),.din(w_dff_A_HbUE7IYu9_0),.clk(gclk));
	jdff dff_A_HJpBciPx2_0(.dout(G351),.din(w_dff_A_HJpBciPx2_0),.clk(gclk));
	jdff dff_A_JAByGg7B5_2(.dout(w_dff_A_EoICxVBu2_0),.din(w_dff_A_JAByGg7B5_2),.clk(gclk));
	jdff dff_A_EoICxVBu2_0(.dout(w_dff_A_gjrpNmAA2_0),.din(w_dff_A_EoICxVBu2_0),.clk(gclk));
	jdff dff_A_gjrpNmAA2_0(.dout(w_dff_A_FAjOD6Oi6_0),.din(w_dff_A_gjrpNmAA2_0),.clk(gclk));
	jdff dff_A_FAjOD6Oi6_0(.dout(w_dff_A_d6sMEsnZ6_0),.din(w_dff_A_FAjOD6Oi6_0),.clk(gclk));
	jdff dff_A_d6sMEsnZ6_0(.dout(w_dff_A_85CUouSP3_0),.din(w_dff_A_d6sMEsnZ6_0),.clk(gclk));
	jdff dff_A_85CUouSP3_0(.dout(w_dff_A_lFczkg4K6_0),.din(w_dff_A_85CUouSP3_0),.clk(gclk));
	jdff dff_A_lFczkg4K6_0(.dout(w_dff_A_VmKEePlN2_0),.din(w_dff_A_lFczkg4K6_0),.clk(gclk));
	jdff dff_A_VmKEePlN2_0(.dout(w_dff_A_XzLmBfRQ1_0),.din(w_dff_A_VmKEePlN2_0),.clk(gclk));
	jdff dff_A_XzLmBfRQ1_0(.dout(w_dff_A_urGzhT8P2_0),.din(w_dff_A_XzLmBfRQ1_0),.clk(gclk));
	jdff dff_A_urGzhT8P2_0(.dout(w_dff_A_4gVZ4j902_0),.din(w_dff_A_urGzhT8P2_0),.clk(gclk));
	jdff dff_A_4gVZ4j902_0(.dout(w_dff_A_C4EbJt2q8_0),.din(w_dff_A_4gVZ4j902_0),.clk(gclk));
	jdff dff_A_C4EbJt2q8_0(.dout(w_dff_A_iCJ2GGev6_0),.din(w_dff_A_C4EbJt2q8_0),.clk(gclk));
	jdff dff_A_iCJ2GGev6_0(.dout(w_dff_A_S4Ge7OwR4_0),.din(w_dff_A_iCJ2GGev6_0),.clk(gclk));
	jdff dff_A_S4Ge7OwR4_0(.dout(G372),.din(w_dff_A_S4Ge7OwR4_0),.clk(gclk));
	jdff dff_A_qRdAfI1F8_2(.dout(w_dff_A_OyvXMKs59_0),.din(w_dff_A_qRdAfI1F8_2),.clk(gclk));
	jdff dff_A_OyvXMKs59_0(.dout(w_dff_A_c0es5wGK8_0),.din(w_dff_A_OyvXMKs59_0),.clk(gclk));
	jdff dff_A_c0es5wGK8_0(.dout(w_dff_A_7Zfn1xMY5_0),.din(w_dff_A_c0es5wGK8_0),.clk(gclk));
	jdff dff_A_7Zfn1xMY5_0(.dout(w_dff_A_fknHQfj16_0),.din(w_dff_A_7Zfn1xMY5_0),.clk(gclk));
	jdff dff_A_fknHQfj16_0(.dout(w_dff_A_85QK85lL7_0),.din(w_dff_A_fknHQfj16_0),.clk(gclk));
	jdff dff_A_85QK85lL7_0(.dout(w_dff_A_5GmK2co63_0),.din(w_dff_A_85QK85lL7_0),.clk(gclk));
	jdff dff_A_5GmK2co63_0(.dout(w_dff_A_oEKfbMSB8_0),.din(w_dff_A_5GmK2co63_0),.clk(gclk));
	jdff dff_A_oEKfbMSB8_0(.dout(w_dff_A_a4QoQGjb7_0),.din(w_dff_A_oEKfbMSB8_0),.clk(gclk));
	jdff dff_A_a4QoQGjb7_0(.dout(w_dff_A_FFSEMvOO7_0),.din(w_dff_A_a4QoQGjb7_0),.clk(gclk));
	jdff dff_A_FFSEMvOO7_0(.dout(w_dff_A_o8MDBcjX5_0),.din(w_dff_A_FFSEMvOO7_0),.clk(gclk));
	jdff dff_A_o8MDBcjX5_0(.dout(w_dff_A_4m1UV7fw5_0),.din(w_dff_A_o8MDBcjX5_0),.clk(gclk));
	jdff dff_A_4m1UV7fw5_0(.dout(G369),.din(w_dff_A_4m1UV7fw5_0),.clk(gclk));
	jdff dff_A_UHzT0RaE1_2(.dout(w_dff_A_KjTc5jEp4_0),.din(w_dff_A_UHzT0RaE1_2),.clk(gclk));
	jdff dff_A_KjTc5jEp4_0(.dout(w_dff_A_BN5PaiSn9_0),.din(w_dff_A_KjTc5jEp4_0),.clk(gclk));
	jdff dff_A_BN5PaiSn9_0(.dout(w_dff_A_ZLF4pp3d5_0),.din(w_dff_A_BN5PaiSn9_0),.clk(gclk));
	jdff dff_A_ZLF4pp3d5_0(.dout(w_dff_A_lgoO7Orz8_0),.din(w_dff_A_ZLF4pp3d5_0),.clk(gclk));
	jdff dff_A_lgoO7Orz8_0(.dout(w_dff_A_ZVNovf346_0),.din(w_dff_A_lgoO7Orz8_0),.clk(gclk));
	jdff dff_A_ZVNovf346_0(.dout(w_dff_A_m3L8a7Bg5_0),.din(w_dff_A_ZVNovf346_0),.clk(gclk));
	jdff dff_A_m3L8a7Bg5_0(.dout(w_dff_A_6yVs5rtw8_0),.din(w_dff_A_m3L8a7Bg5_0),.clk(gclk));
	jdff dff_A_6yVs5rtw8_0(.dout(w_dff_A_hok2NpAF2_0),.din(w_dff_A_6yVs5rtw8_0),.clk(gclk));
	jdff dff_A_hok2NpAF2_0(.dout(w_dff_A_EdHWmoz13_0),.din(w_dff_A_hok2NpAF2_0),.clk(gclk));
	jdff dff_A_EdHWmoz13_0(.dout(w_dff_A_s7KFIQBH1_0),.din(w_dff_A_EdHWmoz13_0),.clk(gclk));
	jdff dff_A_s7KFIQBH1_0(.dout(w_dff_A_e250Ta4u5_0),.din(w_dff_A_s7KFIQBH1_0),.clk(gclk));
	jdff dff_A_e250Ta4u5_0(.dout(w_dff_A_cDq0uFlu5_0),.din(w_dff_A_e250Ta4u5_0),.clk(gclk));
	jdff dff_A_cDq0uFlu5_0(.dout(w_dff_A_Q2ojPoe65_0),.din(w_dff_A_cDq0uFlu5_0),.clk(gclk));
	jdff dff_A_Q2ojPoe65_0(.dout(G399),.din(w_dff_A_Q2ojPoe65_0),.clk(gclk));
	jdff dff_A_PHITdRC31_2(.dout(w_dff_A_Mib1ZxWW6_0),.din(w_dff_A_PHITdRC31_2),.clk(gclk));
	jdff dff_A_Mib1ZxWW6_0(.dout(w_dff_A_GkwRoEH73_0),.din(w_dff_A_Mib1ZxWW6_0),.clk(gclk));
	jdff dff_A_GkwRoEH73_0(.dout(w_dff_A_GDYQeMP93_0),.din(w_dff_A_GkwRoEH73_0),.clk(gclk));
	jdff dff_A_GDYQeMP93_0(.dout(w_dff_A_KRnIQjkJ0_0),.din(w_dff_A_GDYQeMP93_0),.clk(gclk));
	jdff dff_A_KRnIQjkJ0_0(.dout(w_dff_A_s9buAJxf5_0),.din(w_dff_A_KRnIQjkJ0_0),.clk(gclk));
	jdff dff_A_s9buAJxf5_0(.dout(w_dff_A_izzAIYDC1_0),.din(w_dff_A_s9buAJxf5_0),.clk(gclk));
	jdff dff_A_izzAIYDC1_0(.dout(w_dff_A_aDbrixL86_0),.din(w_dff_A_izzAIYDC1_0),.clk(gclk));
	jdff dff_A_aDbrixL86_0(.dout(w_dff_A_qFi8lNVn2_0),.din(w_dff_A_aDbrixL86_0),.clk(gclk));
	jdff dff_A_qFi8lNVn2_0(.dout(G364),.din(w_dff_A_qFi8lNVn2_0),.clk(gclk));
	jdff dff_A_0XfjDTOX8_1(.dout(w_dff_A_OFpUOMpJ2_0),.din(w_dff_A_0XfjDTOX8_1),.clk(gclk));
	jdff dff_A_OFpUOMpJ2_0(.dout(w_dff_A_gpCErC2J7_0),.din(w_dff_A_OFpUOMpJ2_0),.clk(gclk));
	jdff dff_A_gpCErC2J7_0(.dout(w_dff_A_1XaNwXtd4_0),.din(w_dff_A_gpCErC2J7_0),.clk(gclk));
	jdff dff_A_1XaNwXtd4_0(.dout(w_dff_A_zaFEr2Qo4_0),.din(w_dff_A_1XaNwXtd4_0),.clk(gclk));
	jdff dff_A_zaFEr2Qo4_0(.dout(w_dff_A_fjYciVHo3_0),.din(w_dff_A_zaFEr2Qo4_0),.clk(gclk));
	jdff dff_A_fjYciVHo3_0(.dout(w_dff_A_2mzac4AP3_0),.din(w_dff_A_fjYciVHo3_0),.clk(gclk));
	jdff dff_A_2mzac4AP3_0(.dout(w_dff_A_xToQ7eE15_0),.din(w_dff_A_2mzac4AP3_0),.clk(gclk));
	jdff dff_A_xToQ7eE15_0(.dout(w_dff_A_C3fHhtX00_0),.din(w_dff_A_xToQ7eE15_0),.clk(gclk));
	jdff dff_A_C3fHhtX00_0(.dout(w_dff_A_B1rZOdhm8_0),.din(w_dff_A_C3fHhtX00_0),.clk(gclk));
	jdff dff_A_B1rZOdhm8_0(.dout(w_dff_A_RWQgGR7b9_0),.din(w_dff_A_B1rZOdhm8_0),.clk(gclk));
	jdff dff_A_RWQgGR7b9_0(.dout(w_dff_A_TJTCX4ic6_0),.din(w_dff_A_RWQgGR7b9_0),.clk(gclk));
	jdff dff_A_TJTCX4ic6_0(.dout(w_dff_A_pYpDbVvt6_0),.din(w_dff_A_TJTCX4ic6_0),.clk(gclk));
	jdff dff_A_pYpDbVvt6_0(.dout(G396),.din(w_dff_A_pYpDbVvt6_0),.clk(gclk));
	jdff dff_A_w0ospIK34_1(.dout(w_dff_A_s3gw2Kpf0_0),.din(w_dff_A_w0ospIK34_1),.clk(gclk));
	jdff dff_A_s3gw2Kpf0_0(.dout(w_dff_A_OsULOYGU0_0),.din(w_dff_A_s3gw2Kpf0_0),.clk(gclk));
	jdff dff_A_OsULOYGU0_0(.dout(w_dff_A_Hs7YH4XS1_0),.din(w_dff_A_OsULOYGU0_0),.clk(gclk));
	jdff dff_A_Hs7YH4XS1_0(.dout(w_dff_A_kxVVvueZ2_0),.din(w_dff_A_Hs7YH4XS1_0),.clk(gclk));
	jdff dff_A_kxVVvueZ2_0(.dout(w_dff_A_zwwGGmF66_0),.din(w_dff_A_kxVVvueZ2_0),.clk(gclk));
	jdff dff_A_zwwGGmF66_0(.dout(w_dff_A_Qw83aOJF4_0),.din(w_dff_A_zwwGGmF66_0),.clk(gclk));
	jdff dff_A_Qw83aOJF4_0(.dout(w_dff_A_iP8xR4Dp5_0),.din(w_dff_A_Qw83aOJF4_0),.clk(gclk));
	jdff dff_A_iP8xR4Dp5_0(.dout(G384),.din(w_dff_A_iP8xR4Dp5_0),.clk(gclk));
	jdff dff_A_s1BWpEPJ7_2(.dout(w_dff_A_xIPw46ed7_0),.din(w_dff_A_s1BWpEPJ7_2),.clk(gclk));
	jdff dff_A_xIPw46ed7_0(.dout(w_dff_A_Za09WhNt1_0),.din(w_dff_A_xIPw46ed7_0),.clk(gclk));
	jdff dff_A_Za09WhNt1_0(.dout(w_dff_A_KKwkaz148_0),.din(w_dff_A_Za09WhNt1_0),.clk(gclk));
	jdff dff_A_KKwkaz148_0(.dout(w_dff_A_Egy2GMK16_0),.din(w_dff_A_KKwkaz148_0),.clk(gclk));
	jdff dff_A_Egy2GMK16_0(.dout(w_dff_A_hKoYBXx60_0),.din(w_dff_A_Egy2GMK16_0),.clk(gclk));
	jdff dff_A_hKoYBXx60_0(.dout(w_dff_A_L68NbBTi7_0),.din(w_dff_A_hKoYBXx60_0),.clk(gclk));
	jdff dff_A_L68NbBTi7_0(.dout(G367),.din(w_dff_A_L68NbBTi7_0),.clk(gclk));
	jdff dff_A_9T1uPaDL7_1(.dout(w_dff_A_Bt9wVzTt8_0),.din(w_dff_A_9T1uPaDL7_1),.clk(gclk));
	jdff dff_A_Bt9wVzTt8_0(.dout(w_dff_A_XsprfBTq5_0),.din(w_dff_A_Bt9wVzTt8_0),.clk(gclk));
	jdff dff_A_XsprfBTq5_0(.dout(w_dff_A_BPJNqi4P9_0),.din(w_dff_A_XsprfBTq5_0),.clk(gclk));
	jdff dff_A_BPJNqi4P9_0(.dout(w_dff_A_2VS1HYFM1_0),.din(w_dff_A_BPJNqi4P9_0),.clk(gclk));
	jdff dff_A_2VS1HYFM1_0(.dout(w_dff_A_ebIqPRx40_0),.din(w_dff_A_2VS1HYFM1_0),.clk(gclk));
	jdff dff_A_ebIqPRx40_0(.dout(G387),.din(w_dff_A_ebIqPRx40_0),.clk(gclk));
	jdff dff_A_AxGVX6TL1_1(.dout(w_dff_A_P9xmPpsY4_0),.din(w_dff_A_AxGVX6TL1_1),.clk(gclk));
	jdff dff_A_P9xmPpsY4_0(.dout(w_dff_A_bEHImB6t9_0),.din(w_dff_A_P9xmPpsY4_0),.clk(gclk));
	jdff dff_A_bEHImB6t9_0(.dout(w_dff_A_cdgl24GK6_0),.din(w_dff_A_bEHImB6t9_0),.clk(gclk));
	jdff dff_A_cdgl24GK6_0(.dout(w_dff_A_P1VdzwAK9_0),.din(w_dff_A_cdgl24GK6_0),.clk(gclk));
	jdff dff_A_P1VdzwAK9_0(.dout(w_dff_A_21LJ38qi8_0),.din(w_dff_A_P1VdzwAK9_0),.clk(gclk));
	jdff dff_A_21LJ38qi8_0(.dout(w_dff_A_Jq6zQMHU6_0),.din(w_dff_A_21LJ38qi8_0),.clk(gclk));
	jdff dff_A_Jq6zQMHU6_0(.dout(G393),.din(w_dff_A_Jq6zQMHU6_0),.clk(gclk));
	jdff dff_A_4z7A7QZb0_1(.dout(w_dff_A_70oyHGSA9_0),.din(w_dff_A_4z7A7QZb0_1),.clk(gclk));
	jdff dff_A_70oyHGSA9_0(.dout(w_dff_A_K8cjy4tB5_0),.din(w_dff_A_70oyHGSA9_0),.clk(gclk));
	jdff dff_A_K8cjy4tB5_0(.dout(w_dff_A_wsfjiJc34_0),.din(w_dff_A_K8cjy4tB5_0),.clk(gclk));
	jdff dff_A_wsfjiJc34_0(.dout(w_dff_A_DlL4fp6E6_0),.din(w_dff_A_wsfjiJc34_0),.clk(gclk));
	jdff dff_A_DlL4fp6E6_0(.dout(w_dff_A_C38MetWn2_0),.din(w_dff_A_DlL4fp6E6_0),.clk(gclk));
	jdff dff_A_C38MetWn2_0(.dout(G390),.din(w_dff_A_C38MetWn2_0),.clk(gclk));
	jdff dff_A_lKt9RnS31_1(.dout(w_dff_A_eOvyUM789_0),.din(w_dff_A_lKt9RnS31_1),.clk(gclk));
	jdff dff_A_eOvyUM789_0(.dout(w_dff_A_zrE6ZEQR2_0),.din(w_dff_A_eOvyUM789_0),.clk(gclk));
	jdff dff_A_zrE6ZEQR2_0(.dout(w_dff_A_Tyi4ypDL0_0),.din(w_dff_A_zrE6ZEQR2_0),.clk(gclk));
	jdff dff_A_Tyi4ypDL0_0(.dout(G378),.din(w_dff_A_Tyi4ypDL0_0),.clk(gclk));
	jdff dff_A_1rpzyvbw3_1(.dout(w_dff_A_0f7I85Sz6_0),.din(w_dff_A_1rpzyvbw3_1),.clk(gclk));
	jdff dff_A_0f7I85Sz6_0(.dout(w_dff_A_ZtU3tyDA1_0),.din(w_dff_A_0f7I85Sz6_0),.clk(gclk));
	jdff dff_A_ZtU3tyDA1_0(.dout(w_dff_A_OFjJ8rbw8_0),.din(w_dff_A_ZtU3tyDA1_0),.clk(gclk));
	jdff dff_A_OFjJ8rbw8_0(.dout(G375),.din(w_dff_A_OFjJ8rbw8_0),.clk(gclk));
	jdff dff_A_ZFDj4KzA8_1(.dout(w_dff_A_GLrwuIti6_0),.din(w_dff_A_ZFDj4KzA8_1),.clk(gclk));
	jdff dff_A_GLrwuIti6_0(.dout(w_dff_A_ntiPQ6aK5_0),.din(w_dff_A_GLrwuIti6_0),.clk(gclk));
	jdff dff_A_ntiPQ6aK5_0(.dout(w_dff_A_Pr5W43mi1_0),.din(w_dff_A_ntiPQ6aK5_0),.clk(gclk));
	jdff dff_A_Pr5W43mi1_0(.dout(G381),.din(w_dff_A_Pr5W43mi1_0),.clk(gclk));
	jdff dff_A_U9Dhhxdh2_1(.dout(G407),.din(w_dff_A_U9Dhhxdh2_1),.clk(gclk));
	jdff dff_A_nMRnQXEZ3_2(.dout(w_dff_A_c0IRpd548_0),.din(w_dff_A_nMRnQXEZ3_2),.clk(gclk));
	jdff dff_A_c0IRpd548_0(.dout(G402),.din(w_dff_A_c0IRpd548_0),.clk(gclk));
endmodule

