/*

c432:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jdff: 1153
	jand: 111
	jor: 110

Summary:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jdff: 1153
	jand: 111
	jor: 110
*/

module c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n43;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n150;
	wire n151;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n217;
	wire n218;
	wire n219;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n235;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n244;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n262;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G4gat_0;
	wire[2:0] w_G8gat_0;
	wire[2:0] w_G11gat_0;
	wire[2:0] w_G14gat_0;
	wire[2:0] w_G17gat_0;
	wire[2:0] w_G21gat_0;
	wire[1:0] w_G21gat_1;
	wire[1:0] w_G24gat_0;
	wire[1:0] w_G27gat_0;
	wire[1:0] w_G30gat_0;
	wire[2:0] w_G34gat_0;
	wire[2:0] w_G37gat_0;
	wire[1:0] w_G40gat_0;
	wire[2:0] w_G43gat_0;
	wire[1:0] w_G43gat_1;
	wire[1:0] w_G47gat_0;
	wire[2:0] w_G50gat_0;
	wire[1:0] w_G53gat_0;
	wire[2:0] w_G56gat_0;
	wire[2:0] w_G60gat_0;
	wire[2:0] w_G63gat_0;
	wire[1:0] w_G66gat_0;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G73gat_0;
	wire[1:0] w_G76gat_0;
	wire[1:0] w_G79gat_0;
	wire[2:0] w_G82gat_0;
	wire[2:0] w_G86gat_0;
	wire[1:0] w_G86gat_1;
	wire[2:0] w_G89gat_0;
	wire[2:0] w_G92gat_0;
	wire[2:0] w_G95gat_0;
	wire[2:0] w_G99gat_0;
	wire[2:0] w_G102gat_0;
	wire[1:0] w_G105gat_0;
	wire[2:0] w_G108gat_0;
	wire[2:0] w_G112gat_0;
	wire[1:0] w_G115gat_0;
	wire[2:0] w_G223gat_0;
	wire[2:0] w_G223gat_1;
	wire[2:0] w_G223gat_2;
	wire[1:0] w_G223gat_3;
	wire G223gat_fa_;
	wire[2:0] w_G329gat_0;
	wire[2:0] w_G329gat_1;
	wire[2:0] w_G329gat_2;
	wire[2:0] w_G329gat_3;
	wire[2:0] w_G329gat_4;
	wire[2:0] w_G329gat_5;
	wire w_G329gat_6;
	wire G329gat_fa_;
	wire[2:0] w_G370gat_0;
	wire[2:0] w_G370gat_1;
	wire w_G370gat_2;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire[1:0] w_n43_0;
	wire[1:0] w_n44_0;
	wire[1:0] w_n47_0;
	wire[1:0] w_n52_0;
	wire[1:0] w_n53_0;
	wire[1:0] w_n56_0;
	wire[1:0] w_n58_0;
	wire[1:0] w_n61_0;
	wire[1:0] w_n63_0;
	wire[1:0] w_n69_0;
	wire[1:0] w_n71_0;
	wire[1:0] w_n72_0;
	wire[1:0] w_n73_0;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[1:0] w_n79_0;
	wire[1:0] w_n82_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n87_0;
	wire[1:0] w_n89_0;
	wire[2:0] w_n94_0;
	wire[2:0] w_n94_1;
	wire[2:0] w_n94_2;
	wire[2:0] w_n94_3;
	wire[1:0] w_n94_4;
	wire[1:0] w_n96_0;
	wire[1:0] w_n98_0;
	wire[1:0] w_n100_0;
	wire[1:0] w_n107_0;
	wire[1:0] w_n109_0;
	wire[2:0] w_n114_0;
	wire[1:0] w_n115_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n121_0;
	wire[1:0] w_n123_0;
	wire[2:0] w_n126_0;
	wire[1:0] w_n128_0;
	wire[2:0] w_n130_0;
	wire[1:0] w_n132_0;
	wire[1:0] w_n139_0;
	wire[1:0] w_n141_0;
	wire[1:0] w_n142_0;
	wire[1:0] w_n145_0;
	wire[1:0] w_n146_0;
	wire[1:0] w_n147_0;
	wire[1:0] w_n150_0;
	wire[1:0] w_n151_0;
	wire[1:0] w_n154_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n159_0;
	wire[1:0] w_n164_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n174_0;
	wire[1:0] w_n177_0;
	wire[2:0] w_n182_0;
	wire[2:0] w_n182_1;
	wire[2:0] w_n182_2;
	wire[1:0] w_n182_3;
	wire[1:0] w_n184_0;
	wire[1:0] w_n188_0;
	wire[1:0] w_n191_0;
	wire[1:0] w_n193_0;
	wire[1:0] w_n197_0;
	wire[1:0] w_n198_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n205_0;
	wire[1:0] w_n217_0;
	wire[1:0] w_n219_0;
	wire[1:0] w_n222_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n231_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n260_0;
	wire[2:0] w_n271_0;
	wire[2:0] w_n271_1;
	wire[2:0] w_n271_2;
	wire[1:0] w_n271_3;
	wire[1:0] w_n274_0;
	wire[1:0] w_n281_0;
	wire[1:0] w_n283_0;
	wire[1:0] w_n286_0;
	wire[1:0] w_n290_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n296_0;
	wire[1:0] w_n303_0;
	wire[1:0] w_n305_0;
	wire[1:0] w_n313_0;
	wire[1:0] w_n314_0;
	wire[2:0] w_n317_0;
	wire[1:0] w_n319_0;
	wire w_dff_B_E84WjtqU9_1;
	wire w_dff_B_b9HyKMji5_1;
	wire w_dff_B_qeEHfVCL7_1;
	wire w_dff_B_brIiDbPX4_0;
	wire w_dff_B_PyLHbrk94_0;
	wire w_dff_B_PqG1ajbQ5_0;
	wire w_dff_B_jNwrjMXK6_0;
	wire w_dff_B_uBsrld240_0;
	wire w_dff_B_ssGiefmH9_1;
	wire w_dff_A_63oNAdLK8_0;
	wire w_dff_B_OQVJCjD14_0;
	wire w_dff_B_yJb4L9dF8_0;
	wire w_dff_B_GRe8qVV25_0;
	wire w_dff_B_immWqEAs3_0;
	wire w_dff_B_5cwfiVA75_0;
	wire w_dff_A_LMnmGZJm4_0;
	wire w_dff_B_FhGW1nOI6_1;
	wire w_dff_B_lX9AQn0i9_0;
	wire w_dff_B_jefqsd6x1_0;
	wire w_dff_B_8qO7u2pw1_0;
	wire w_dff_B_qrSNogx69_0;
	wire w_dff_B_6ReuljeS7_0;
	wire w_dff_A_bhanmIps5_0;
	wire w_dff_A_we74WJ5x3_0;
	wire w_dff_A_HiEgvwr16_0;
	wire w_dff_A_LhdOrUZ06_0;
	wire w_dff_A_UWlYa7UW3_0;
	wire w_dff_A_Wxwv153g2_0;
	wire w_dff_A_mRCu6KOv1_0;
	wire w_dff_B_Pt70dW2M2_1;
	wire w_dff_B_RGMPKndI4_1;
	wire w_dff_B_7cuj51sA5_1;
	wire w_dff_B_v7onULsi4_1;
	wire w_dff_B_9HZyP6Zc0_1;
	wire w_dff_B_osD97IsC4_1;
	wire w_dff_B_BXLEhURq1_1;
	wire w_dff_B_1B5oGgdT8_1;
	wire w_dff_B_6GpfLvS53_1;
	wire w_dff_B_Do7VOgU68_1;
	wire w_dff_B_D2q8IV318_1;
	wire w_dff_B_On0SCoFm1_1;
	wire w_dff_B_A8tYvMnT1_1;
	wire w_dff_B_GXgKwjET1_1;
	wire w_dff_B_f1PbK5JV1_1;
	wire w_dff_B_JchGTsiz1_1;
	wire w_dff_B_QYQQMzsr4_1;
	wire w_dff_B_5h4ow6XR1_1;
	wire w_dff_B_KJ6kQ9ow5_1;
	wire w_dff_B_bTfpLFxD2_1;
	wire w_dff_B_TaFCL5fq0_1;
	wire w_dff_B_bYlbaeYM8_1;
	wire w_dff_B_gpnxk3wg2_1;
	wire w_dff_B_B7uisLfx7_1;
	wire w_dff_B_2wFSzp307_1;
	wire w_dff_B_K1thgq319_1;
	wire w_dff_B_uTuShrve9_1;
	wire w_dff_B_0v3JXI7t8_0;
	wire w_dff_B_zcZgJHWH2_0;
	wire w_dff_B_wR8dz6dx4_0;
	wire w_dff_A_xKJdmaWY3_1;
	wire w_dff_A_JxDwUKru5_1;
	wire w_dff_A_rH4XgQez6_1;
	wire w_dff_A_FX0Locty1_1;
	wire w_dff_A_G9mKx2417_1;
	wire w_dff_A_7RxalIYA6_1;
	wire w_dff_B_y8DmVsDm4_1;
	wire w_dff_B_3s5pqZGe8_0;
	wire w_dff_B_qJUcp0DF8_0;
	wire w_dff_B_De8g2oe11_0;
	wire w_dff_B_knX7jJXR9_0;
	wire w_dff_B_biS7DsnS2_0;
	wire w_dff_B_AxRQ3LvL6_1;
	wire w_dff_B_ogrRlWLn5_0;
	wire w_dff_B_6wxqCpKy4_0;
	wire w_dff_B_BzcxujOr8_0;
	wire w_dff_B_ct5lXz6H6_0;
	wire w_dff_A_cFHfMqxb5_0;
	wire w_dff_A_sOeOPPvk6_0;
	wire w_dff_A_ILdHlcoY5_0;
	wire w_dff_A_rPIuqBvc7_0;
	wire w_dff_A_HsczOm9L7_0;
	wire w_dff_A_t8PbktgK8_0;
	wire w_dff_A_35Waeda05_0;
	wire w_dff_A_f8rAJGZn9_0;
	wire w_dff_A_VopBQ54b6_0;
	wire w_dff_A_CpLrv76n4_0;
	wire w_dff_A_6IO6HRAS4_0;
	wire w_dff_A_MfOkD83t9_0;
	wire w_dff_A_exauHlsj2_0;
	wire w_dff_A_BGslSIQO3_0;
	wire w_dff_A_34zFNiej2_0;
	wire w_dff_A_EdUu0n264_0;
	wire w_dff_A_brlJoA973_0;
	wire w_dff_A_v9VcLd3g7_0;
	wire w_dff_B_QrmimWgB9_0;
	wire w_dff_B_nAh1Dqaq0_0;
	wire w_dff_B_qFZ28XBB5_0;
	wire w_dff_B_J09rXRIQ9_0;
	wire w_dff_B_hFem99714_0;
	wire w_dff_B_Nl3mb62H5_0;
	wire w_dff_B_2TnlZEFq4_1;
	wire w_dff_B_A6RWogJ76_1;
	wire w_dff_B_Lmvqt5U65_1;
	wire w_dff_A_Gxyn36e49_0;
	wire w_dff_A_BPcPin6M4_0;
	wire w_dff_A_vl4FimtG9_0;
	wire w_dff_A_ReyVoHjd7_0;
	wire w_dff_A_qyrcAqG02_0;
	wire w_dff_A_uWXJDqR56_0;
	wire w_dff_A_YiRU4dyJ8_0;
	wire w_dff_A_URdEWoJq1_0;
	wire w_dff_A_GcCtW2Bk8_0;
	wire w_dff_A_ILCPC6pi0_0;
	wire w_dff_A_yc8ikB592_0;
	wire w_dff_B_BXQdMy1D2_2;
	wire w_dff_B_YvDbImdz1_2;
	wire w_dff_B_J54WOYsi1_2;
	wire w_dff_B_5wjd3s9X3_2;
	wire w_dff_B_X0bT0CAM4_2;
	wire w_dff_B_Pf9E87fF5_2;
	wire w_dff_B_EeTdyLnm5_2;
	wire w_dff_B_GKHCdxW71_2;
	wire w_dff_B_Ai9M8hI28_2;
	wire w_dff_B_Ej7AXUqa7_2;
	wire w_dff_B_GewKCm6z4_2;
	wire w_dff_B_iI5YOLjt6_2;
	wire w_dff_B_bPCAM6l94_2;
	wire w_dff_B_Xc4m6MZ12_2;
	wire w_dff_A_utroPy4g4_0;
	wire w_dff_A_c5IvWWXm1_0;
	wire w_dff_A_JsiZLXWc6_0;
	wire w_dff_A_0l8e7Srp5_0;
	wire w_dff_A_BeTwbTta5_0;
	wire w_dff_A_qXG8zpi81_0;
	wire w_dff_A_aquxKKMG8_0;
	wire w_dff_A_vzFMzJ0s6_0;
	wire w_dff_A_8MUZIVM40_0;
	wire w_dff_A_8F4L9rEQ2_0;
	wire w_dff_A_C0gpur6a9_0;
	wire w_dff_A_fLHyWBkp6_0;
	wire w_dff_A_SVCRgDDz1_0;
	wire w_dff_A_NSGXEAav9_0;
	wire w_dff_A_pTPvviVi8_0;
	wire w_dff_A_8FZZKRYL6_1;
	wire w_dff_A_Md7vrpUJ3_1;
	wire w_dff_A_iVHeoyJr4_1;
	wire w_dff_A_d54mL2Om9_1;
	wire w_dff_A_K09wiWK30_0;
	wire w_dff_A_Buj8wYlS7_0;
	wire w_dff_A_KYC09Ls34_0;
	wire w_dff_A_7fQt6V3F4_0;
	wire w_dff_A_lTgL6P0O2_0;
	wire w_dff_A_1lx8uWHB5_0;
	wire w_dff_A_8CavIptA0_0;
	wire w_dff_A_aHV4aXfV4_0;
	wire w_dff_A_NEDzp6qH5_0;
	wire w_dff_A_0nqLD8yi9_0;
	wire w_dff_A_oe4tlPCg9_0;
	wire w_dff_B_2YcemIQ92_2;
	wire w_dff_B_tiulCnbL2_2;
	wire w_dff_B_QmYJJC3n9_2;
	wire w_dff_B_1u29ajOh1_2;
	wire w_dff_B_MywoQ7js6_2;
	wire w_dff_B_s9cZoVTR0_2;
	wire w_dff_B_FK9puWpO4_2;
	wire w_dff_B_FVREnZD71_2;
	wire w_dff_A_cQwLVOFm7_0;
	wire w_dff_A_m7jWDz0S8_0;
	wire w_dff_A_DW59HpH40_0;
	wire w_dff_A_0KVgAVg85_0;
	wire w_dff_A_J9e7HbqY0_0;
	wire w_dff_A_vKW4BJrW4_0;
	wire w_dff_A_EiWeU5AG8_0;
	wire w_dff_A_DysaCDw63_0;
	wire w_dff_A_nUqJJRf63_0;
	wire w_dff_A_MZWkJju34_0;
	wire w_dff_A_YHUwgax27_0;
	wire w_dff_A_92M2Zl8z8_0;
	wire w_dff_A_JQajJs659_0;
	wire w_dff_A_C34rz9Fg0_0;
	wire w_dff_A_FMGlxFBl8_0;
	wire w_dff_A_3UWegJy00_0;
	wire w_dff_A_oqTTcQyO7_0;
	wire w_dff_A_prfLRcRV9_0;
	wire w_dff_A_LB8w7xGO3_0;
	wire w_dff_A_cF2UM3na6_0;
	wire w_dff_B_JAtH6QYN6_1;
	wire w_dff_B_hknoBpDP2_1;
	wire w_dff_B_DlPlRZMf2_1;
	wire w_dff_B_Oi1GTYA27_1;
	wire w_dff_B_S0fUgJk15_1;
	wire w_dff_B_OTZRNQks9_1;
	wire w_dff_B_14PyE8ru3_1;
	wire w_dff_B_5iSKiwbu5_1;
	wire w_dff_B_lmSBl0DE6_1;
	wire w_dff_B_QaaHamPu0_1;
	wire w_dff_B_sg2gjBky1_1;
	wire w_dff_B_9ISUfuz87_1;
	wire w_dff_B_ip6L2EgA2_1;
	wire w_dff_B_9un0dYnS5_1;
	wire w_dff_B_pHw88pEo3_1;
	wire w_dff_B_BkoH1c7b4_1;
	wire w_dff_B_17QKc4032_1;
	wire w_dff_B_lY72b7Xi2_1;
	wire w_dff_B_uI2FUQZx0_1;
	wire w_dff_B_mdbxgMUr0_1;
	wire w_dff_B_SxTdgAXJ1_1;
	wire w_dff_B_3132phCB1_1;
	wire w_dff_B_oeRnJ07C6_1;
	wire w_dff_B_iun8o7aA0_1;
	wire w_dff_B_HCkoYt0G3_1;
	wire w_dff_B_uTCzO6Hi1_1;
	wire w_dff_A_EGoBSwq17_0;
	wire w_dff_A_2xI4MMCA4_0;
	wire w_dff_A_nKU2a0Vu7_0;
	wire w_dff_A_yyqq8xVU6_0;
	wire w_dff_A_AXZdTIEi1_0;
	wire w_dff_A_FVHJF5re9_0;
	wire w_dff_A_1h2Dwb9x6_0;
	wire w_dff_A_WcHWZvVs0_0;
	wire w_dff_A_3SBLw8T22_0;
	wire w_dff_A_05ial6b11_0;
	wire w_dff_A_xDYdVTql6_0;
	wire w_dff_A_fqOMxiy43_0;
	wire w_dff_A_CSfFWcDW9_0;
	wire w_dff_A_vupmUNby3_0;
	wire w_dff_A_ZHfG6End6_0;
	wire w_dff_A_4B1Y14dG6_1;
	wire w_dff_A_fY67RCm50_1;
	wire w_dff_A_5aq5BgUk0_1;
	wire w_dff_A_5WXQxHvf4_1;
	wire w_dff_A_N7RMsra07_1;
	wire w_dff_A_ttO0wQNS8_1;
	wire w_dff_A_hvodjvo19_1;
	wire w_dff_A_9Tt24nFE8_1;
	wire w_dff_A_qG53VjYE0_1;
	wire w_dff_A_MCyEELYN1_1;
	wire w_dff_A_CXtccuCO5_1;
	wire w_dff_A_OXbuJOhc8_1;
	wire w_dff_A_Pg9Yihf36_1;
	wire w_dff_A_2txbwMG71_1;
	wire w_dff_A_MaAgopZo4_1;
	wire w_dff_A_bKmBPZRg6_1;
	wire w_dff_A_OxR6szJ24_1;
	wire w_dff_A_ZVkNtnPK5_1;
	wire w_dff_A_jU2YAEAb7_1;
	wire w_dff_A_SRPEcVSu0_1;
	wire w_dff_A_GIavFXJY4_0;
	wire w_dff_A_h5nScqoq6_0;
	wire w_dff_A_bmkzxTd32_0;
	wire w_dff_A_t6BzmpDP7_0;
	wire w_dff_A_bSlRV5rd6_0;
	wire w_dff_A_EaVkdNfv5_0;
	wire w_dff_B_OFiT3GSp7_2;
	wire w_dff_B_RVlDbZ9m5_2;
	wire w_dff_B_cC7ubkQR1_2;
	wire w_dff_B_mQCHZgxH2_2;
	wire w_dff_B_2HGfSuSX4_2;
	wire w_dff_B_tbPTYDfA0_2;
	wire w_dff_B_wyfG7C8O2_2;
	wire w_dff_B_gGq2oYPE6_2;
	wire w_dff_B_KiPOa9Mz8_2;
	wire w_dff_B_qkYuge6v6_2;
	wire w_dff_B_y1rL8AYV0_2;
	wire w_dff_B_A10GNPnt2_2;
	wire w_dff_B_FbCWni4c0_2;
	wire w_dff_A_iu1WqPGS5_0;
	wire w_dff_A_QB91sCtJ1_0;
	wire w_dff_A_sMMDcdY31_0;
	wire w_dff_A_ayzV43KE6_0;
	wire w_dff_A_wcIEbD2x8_0;
	wire w_dff_A_HqxwDOul0_0;
	wire w_dff_A_VDAhH8S32_0;
	wire w_dff_A_UHZ0AsGE3_0;
	wire w_dff_A_4DJfSLme3_0;
	wire w_dff_A_Lwyjt1Bi4_0;
	wire w_dff_A_TJWqEGNl2_0;
	wire w_dff_A_9mjOUV812_0;
	wire w_dff_A_VwzK9wRe3_0;
	wire w_dff_A_1VuSXTht4_0;
	wire w_dff_A_16Mc6rX52_0;
	wire w_dff_A_ixNMUFVr3_0;
	wire w_dff_A_x7kcPeyr0_0;
	wire w_dff_A_PtVh3klS2_0;
	wire w_dff_A_tnePtMzo9_0;
	wire w_dff_A_6AlgyhNC8_0;
	wire w_dff_A_As8JnspT9_1;
	wire w_dff_A_MqMPAM8g8_1;
	wire w_dff_A_ZatDco8P9_1;
	wire w_dff_A_86c3BzAz2_1;
	wire w_dff_A_KQaawdCQ0_1;
	wire w_dff_A_xrOA8BGO2_1;
	wire w_dff_A_dZYOYQUF7_1;
	wire w_dff_A_fVk5TWhd6_1;
	wire w_dff_A_nZQQ6A4D3_1;
	wire w_dff_A_G9tl59HE2_1;
	wire w_dff_A_Y957lquf4_1;
	wire w_dff_A_VB0sQ4Hs6_1;
	wire w_dff_A_C7BTkScG1_1;
	wire w_dff_A_pVnNe7Ql2_1;
	wire w_dff_A_k4Y51fI90_0;
	wire w_dff_A_ZEYuEmjA2_0;
	wire w_dff_A_1kLqxltu3_0;
	wire w_dff_A_femnjQoD9_0;
	wire w_dff_A_iN4N0kGU2_0;
	wire w_dff_A_fS7LI9u52_0;
	wire w_dff_A_PXdOYgUc3_0;
	wire w_dff_A_9EHkEeAd8_0;
	wire w_dff_A_Kkzt62QM3_0;
	wire w_dff_A_WeIUFYL15_0;
	wire w_dff_A_x4Avr8QU9_0;
	wire w_dff_A_5vpnn1Hd2_0;
	wire w_dff_B_aM77vvQf2_2;
	wire w_dff_B_4yFEp7qB2_2;
	wire w_dff_B_Gwg8VPr55_2;
	wire w_dff_B_s9r5tMvl0_2;
	wire w_dff_B_8Xzm0hvr0_2;
	wire w_dff_B_lY5v2AR60_2;
	wire w_dff_B_HoljFIyH1_2;
	wire w_dff_B_7w6Ty0cH2_2;
	wire w_dff_B_KJLzsaIP2_2;
	wire w_dff_B_2neI1Evm1_2;
	wire w_dff_B_iHgdOBnX0_2;
	wire w_dff_B_gKPkkoLp1_2;
	wire w_dff_B_DTbtNB9T8_2;
	wire w_dff_A_RBEnPNtx5_0;
	wire w_dff_A_UxsZlsHM9_0;
	wire w_dff_A_CVFKzrvw5_0;
	wire w_dff_A_Ffcnbr041_0;
	wire w_dff_A_FVdGMKIu8_0;
	wire w_dff_A_KxsXErZn8_0;
	wire w_dff_A_G03M6b2O4_0;
	wire w_dff_A_RMwHhFwb4_0;
	wire w_dff_A_1iaXrsKi2_0;
	wire w_dff_A_PQW8m0Zz5_0;
	wire w_dff_A_HhqMSUCE3_0;
	wire w_dff_A_QAFcLRcE5_0;
	wire w_dff_A_PM6y6Rac5_0;
	wire w_dff_A_fuz1QEUW2_0;
	wire w_dff_A_QVMlWibB4_0;
	wire w_dff_A_TsTr8HVb4_0;
	wire w_dff_A_FBjetoBE9_0;
	wire w_dff_A_EdBUKRpG0_0;
	wire w_dff_A_nT7qtMo65_0;
	wire w_dff_A_D4Qlff1r3_0;
	wire w_dff_A_RPite0FH3_1;
	wire w_dff_A_EkWQoan84_1;
	wire w_dff_A_YD5yqhga5_1;
	wire w_dff_A_MDTRry8g2_1;
	wire w_dff_A_xqOc8yYE8_1;
	wire w_dff_A_AnpFQgZC3_1;
	wire w_dff_A_7K0OEzMt0_1;
	wire w_dff_B_PEalnbEV7_0;
	wire w_dff_B_ziLYTqk45_0;
	wire w_dff_B_mjnAvtN12_0;
	wire w_dff_B_EJ7mrd9b3_0;
	wire w_dff_B_6ncqurZe4_0;
	wire w_dff_A_ND367Ak01_0;
	wire w_dff_A_z15boVMH8_0;
	wire w_dff_A_FVMnuiyI7_0;
	wire w_dff_A_OKMn6FoW1_0;
	wire w_dff_A_TpvHyZ6w5_0;
	wire w_dff_A_hujdfCwR5_0;
	wire w_dff_A_3vP2MEBK1_0;
	wire w_dff_A_ZZbiFHxe9_0;
	wire w_dff_A_20UkTApF4_0;
	wire w_dff_A_QkA2Cbpy2_0;
	wire w_dff_A_M9pP9sKD7_0;
	wire w_dff_A_fNheglJ38_0;
	wire w_dff_A_1MLnXUWn3_0;
	wire w_dff_A_FtZ0zyZN3_0;
	wire w_dff_A_5dlSNhTG7_0;
	wire w_dff_A_S0eMVCQg5_0;
	wire w_dff_A_kPIoaThd5_0;
	wire w_dff_A_E4SvCZKX6_0;
	wire w_dff_A_IL5ZPbh26_0;
	wire w_dff_A_55F6uHpY0_0;
	wire w_dff_A_mmTeX8682_0;
	wire w_dff_A_5yGrNJrr8_0;
	wire w_dff_A_Yaq6pThX1_0;
	wire w_dff_A_j0pUy80B5_0;
	wire w_dff_A_yaHGqrTN8_0;
	wire w_dff_A_tsRvy61C7_0;
	wire w_dff_A_xGJQImtM9_0;
	wire w_dff_A_sNgvTVzH1_0;
	wire w_dff_A_mw0Elirt8_0;
	wire w_dff_A_3NOVNtP00_0;
	wire w_dff_A_hxBmxHZL4_0;
	wire w_dff_A_XeTWTHoh5_0;
	wire w_dff_A_yaRqaiCT1_0;
	wire w_dff_A_JoSfo5vs7_0;
	wire w_dff_A_EAw1ZGuB9_0;
	wire w_dff_A_tJmv72Z84_0;
	wire w_dff_A_8EFlvp4J9_0;
	wire w_dff_A_RSoaLTfG0_0;
	wire w_dff_A_i8Zztezs4_0;
	wire w_dff_A_Nb4pAod21_0;
	wire w_dff_A_Myvlt2t65_0;
	wire w_dff_A_Vi320bna1_0;
	wire w_dff_A_zwrhq5XR9_0;
	wire w_dff_A_ghXPkxnc5_0;
	wire w_dff_A_SI3AbHif1_0;
	wire w_dff_B_YUN2JMjJ6_1;
	wire w_dff_A_BJHSwyQx8_0;
	wire w_dff_A_tzT4W7pv5_0;
	wire w_dff_A_KpLEh9Nu4_0;
	wire w_dff_A_g2C6mCoA6_0;
	wire w_dff_A_K6YDEDBB2_0;
	wire w_dff_A_CLTiIAIk1_0;
	wire w_dff_A_FZjuf3g77_0;
	wire w_dff_A_2vwPjiJL8_0;
	wire w_dff_A_0vRLJBEb8_0;
	wire w_dff_A_AleaHKx53_0;
	wire w_dff_A_owB79coh6_0;
	wire w_dff_A_KrOIrhnz6_0;
	wire w_dff_B_PhXamBYL5_1;
	wire w_dff_B_pTSn0IBv6_1;
	wire w_dff_B_ALspOavY2_1;
	wire w_dff_B_3m7qSE6r0_1;
	wire w_dff_B_cCWLRHyF8_1;
	wire w_dff_B_U5uq0R0n0_1;
	wire w_dff_A_4ZHIWnzA2_0;
	wire w_dff_A_9EIJR6911_0;
	wire w_dff_A_3NZ7AJHN7_0;
	wire w_dff_A_f8IuNFel1_0;
	wire w_dff_B_AkYWyoNi7_2;
	wire w_dff_B_N2hdPM6Q1_0;
	wire w_dff_B_k0oKSxZz6_0;
	wire w_dff_B_6Ya57KKM4_0;
	wire w_dff_B_J5sydVXs4_0;
	wire w_dff_A_dXqkiOAU8_0;
	wire w_dff_A_pAt8pkO59_0;
	wire w_dff_A_hdoSAK8G1_0;
	wire w_dff_A_VRgXca2F3_0;
	wire w_dff_A_xYBILegS7_0;
	wire w_dff_A_BB2erPz25_0;
	wire w_dff_A_9aOj0izt2_0;
	wire w_dff_A_SKkCYDpZ5_0;
	wire w_dff_A_cvorLVXz3_0;
	wire w_dff_A_tpRIXYBS3_0;
	wire w_dff_A_NCLTK07C8_0;
	wire w_dff_A_1LY0ds4S1_0;
	wire w_dff_A_BbvkIzyJ6_0;
	wire w_dff_A_Thzz6PHF7_0;
	wire w_dff_A_znumnVVH6_0;
	wire w_dff_A_hgmNFIf31_0;
	wire w_dff_A_77ukaDLg7_0;
	wire w_dff_A_femGqmDM7_0;
	wire w_dff_A_U3sk8za80_0;
	wire w_dff_A_DAbPBAop5_0;
	wire w_dff_A_gDMg3dVH5_0;
	wire w_dff_A_bHqQwJqX2_0;
	wire w_dff_A_Rx2Dkhn52_0;
	wire w_dff_B_pdLOxC067_2;
	wire w_dff_B_hWWK1P840_2;
	wire w_dff_B_0s5a6xyR5_2;
	wire w_dff_B_kGkSn32F0_2;
	wire w_dff_B_C1fnISYO9_2;
	wire w_dff_B_OyKpGCGx9_2;
	wire w_dff_B_IDlmOMsx9_2;
	wire w_dff_B_UJP0Ddyk4_2;
	wire w_dff_B_y3wFeHkE4_2;
	wire w_dff_B_kX6bMGpm6_2;
	wire w_dff_B_dBcBY3pX1_2;
	wire w_dff_B_tD1JO75M7_2;
	wire w_dff_B_R0nRX52Z0_2;
	wire w_dff_B_ptDOWvoi1_2;
	wire w_dff_A_lHI0qlei8_0;
	wire w_dff_A_u8LNLsDM7_0;
	wire w_dff_A_TrDj6usd7_0;
	wire w_dff_A_o3heIQwe7_0;
	wire w_dff_A_1DiCN2SE6_0;
	wire w_dff_A_IZWfG0Lt4_0;
	wire w_dff_A_GMWXHIOT4_0;
	wire w_dff_A_JG7gYZDR4_0;
	wire w_dff_A_KBsHaoqG0_0;
	wire w_dff_A_O6t7W3kg8_0;
	wire w_dff_A_YDw0EU7O7_0;
	wire w_dff_A_lcXDKDi94_0;
	wire w_dff_A_WmywqqHu6_0;
	wire w_dff_A_pbkj0S0E2_0;
	wire w_dff_A_qE4HPvK16_0;
	wire w_dff_A_pzLyM3gx7_1;
	wire w_dff_A_zBABjna93_1;
	wire w_dff_A_MsasnzLU9_1;
	wire w_dff_A_cP8VsnHO1_1;
	wire w_dff_A_JeaOdzIB6_1;
	wire w_dff_A_JNGfH7qg4_1;
	wire w_dff_A_BrRnh4N75_0;
	wire w_dff_A_nOrIbI2l9_0;
	wire w_dff_A_AdX6YHTy3_0;
	wire w_dff_A_RSASyS4r5_0;
	wire w_dff_A_miWn5h5e1_0;
	wire w_dff_A_8ZQC5ilP0_0;
	wire w_dff_A_xtnGSsQG6_0;
	wire w_dff_A_FysE8gZR8_0;
	wire w_dff_A_MOoBy9eR6_0;
	wire w_dff_A_HCy3xjCo5_0;
	wire w_dff_A_Zy3wGKlo0_0;
	wire w_dff_A_vBJ43En75_0;
	wire w_dff_B_e3BDnmtq8_2;
	wire w_dff_B_d2JeyH4E2_2;
	wire w_dff_B_UbCuBvmm9_2;
	wire w_dff_B_hQwbeBWj0_2;
	wire w_dff_B_5hU28amv6_2;
	wire w_dff_B_5VaHrKr32_2;
	wire w_dff_B_GAX9VgP40_2;
	wire w_dff_A_bBUItHpo9_0;
	wire w_dff_A_N49Y5pdL3_0;
	wire w_dff_A_WKna2wMk9_0;
	wire w_dff_A_qgkIiCyx0_0;
	wire w_dff_A_TFxqJ3Iw1_0;
	wire w_dff_A_N4fYCRD64_0;
	wire w_dff_A_8RG6u1X27_0;
	wire w_dff_A_wa1cESpL0_0;
	wire w_dff_A_bNP1P9KA6_0;
	wire w_dff_A_phYwgwFP5_0;
	wire w_dff_A_WPuFpHnU9_0;
	wire w_dff_A_Uz8owtnF2_0;
	wire w_dff_A_8hZSAhgg7_0;
	wire w_dff_A_7NOKzKGz5_0;
	wire w_dff_A_aNRS81IT1_0;
	wire w_dff_A_bvacKOWW7_0;
	wire w_dff_A_Xf476TJt8_0;
	wire w_dff_A_3lvclMmW7_0;
	wire w_dff_A_nKJbfG0F3_0;
	wire w_dff_A_2DolGJBw8_0;
	wire w_dff_A_slBXbMmL5_1;
	wire w_dff_A_JDwlrsJB1_1;
	wire w_dff_A_vPCPcutH4_1;
	wire w_dff_A_B6fkMwmI7_1;
	wire w_dff_A_0NKTxPqa0_0;
	wire w_dff_A_aDoKFDYl3_0;
	wire w_dff_A_S9rIC2Lj5_0;
	wire w_dff_A_l6mBzRnm6_0;
	wire w_dff_A_DcnG9xyW5_0;
	wire w_dff_A_bgm1NLjI3_0;
	wire w_dff_A_EPfnWR8I7_0;
	wire w_dff_B_FO7OnCup9_1;
	wire w_dff_B_W4NMkniy8_1;
	wire w_dff_A_4kiezU4t7_0;
	wire w_dff_A_JjNGq4TP7_0;
	wire w_dff_A_Y0ChjMwC4_0;
	wire w_dff_A_rsos5Fm00_0;
	wire w_dff_A_zrmGGB885_0;
	wire w_dff_A_L7UkzfMe6_0;
	wire w_dff_A_qOfXCRrd5_0;
	wire w_dff_A_tAC1vEVq3_0;
	wire w_dff_A_Q7enk1ph6_0;
	wire w_dff_A_ORMBbBKv0_0;
	wire w_dff_A_JeYl2SgM1_0;
	wire w_dff_A_Yds801NX3_1;
	wire w_dff_A_wC0HanK92_1;
	wire w_dff_A_7o98vxHV9_1;
	wire w_dff_A_XMDxYmPO5_1;
	wire w_dff_A_tO3P15gs0_1;
	wire w_dff_B_etPOqWoX6_3;
	wire w_dff_B_zcnCxPAJ4_3;
	wire w_dff_B_nzUlwps71_3;
	wire w_dff_B_a4rYuHcC1_3;
	wire w_dff_B_7l1AWG7J3_3;
	wire w_dff_B_aKs3vIiu9_3;
	wire w_dff_B_EzKS0AVu8_3;
	wire w_dff_A_mcgw9Ud00_0;
	wire w_dff_A_VIkFKt1a2_0;
	wire w_dff_A_8NeDOyXR5_0;
	wire w_dff_A_xetB8bEd4_0;
	wire w_dff_A_SpFOPOTi6_0;
	wire w_dff_A_2WIHBanQ2_0;
	wire w_dff_A_cwD07wTi9_0;
	wire w_dff_A_oiRTHhbG8_0;
	wire w_dff_A_UZM8Wk3A5_1;
	wire w_dff_A_1vWXWuOn0_1;
	wire w_dff_A_2fjhSJ0N7_1;
	wire w_dff_A_oRrvzPiG2_1;
	wire w_dff_A_HCmVVddG2_1;
	wire w_dff_A_Qc06GbXM9_1;
	wire w_dff_A_kKhWHCdr7_1;
	wire w_dff_A_y96emqx31_1;
	wire w_dff_A_AW856LJC9_1;
	wire w_dff_A_kWw48Eko2_1;
	wire w_dff_A_DTf9QwgS4_1;
	wire w_dff_A_B894nJWu0_1;
	wire w_dff_A_PtjufDcc3_1;
	wire w_dff_A_ATVsHW0w7_2;
	wire w_dff_A_hypxtFVw3_2;
	wire w_dff_A_2ySw7LK83_2;
	wire w_dff_A_Jkl7f8Sw0_2;
	wire w_dff_A_E1G6jHtS0_2;
	wire w_dff_A_AYZHWwhS7_2;
	wire w_dff_A_qx90NEen5_2;
	wire w_dff_A_I2ZQzOpn0_2;
	wire w_dff_A_zExR2g2s7_2;
	wire w_dff_A_ooD55aNS0_2;
	wire w_dff_A_m9XC5wV75_2;
	wire w_dff_A_AtWLHQnD3_2;
	wire w_dff_A_WshjxAfQ5_2;
	wire w_dff_A_r3iUyr916_0;
	wire w_dff_A_jbdTcvks0_0;
	wire w_dff_A_xoEPukCl6_0;
	wire w_dff_A_spmvP23Z7_0;
	wire w_dff_A_o2LkBOIf7_0;
	wire w_dff_A_ZIsEgJ3T1_0;
	wire w_dff_A_pP8qmPLt9_0;
	wire w_dff_A_haE2X7L63_0;
	wire w_dff_A_vm1ylt3D2_0;
	wire w_dff_A_68hyfJC96_0;
	wire w_dff_A_3b6KP1Xr0_0;
	wire w_dff_A_N6wzs6ac4_1;
	wire w_dff_A_pXKmNmg82_1;
	wire w_dff_A_BCsn4f764_1;
	wire w_dff_A_gC6VUEAN1_1;
	wire w_dff_A_lHnmXJzK4_1;
	wire w_dff_B_s7j9ayXP8_3;
	wire w_dff_B_uEIqphoG9_3;
	wire w_dff_B_CRyaFUlM7_3;
	wire w_dff_B_CneCEBHj1_3;
	wire w_dff_B_RXJVo6698_3;
	wire w_dff_B_RMj0V95O8_3;
	wire w_dff_B_YeLHtNcC6_3;
	wire w_dff_A_dpeMo0y88_0;
	wire w_dff_A_ijkCNXde3_0;
	wire w_dff_A_7NuyewkD5_0;
	wire w_dff_A_ZZbdYIde3_0;
	wire w_dff_A_kj0XBpzp1_0;
	wire w_dff_A_Zn33bEhK9_0;
	wire w_dff_A_GsVNaxDu9_0;
	wire w_dff_A_yjVedfVQ4_0;
	wire w_dff_A_cUR0wbUU5_1;
	wire w_dff_A_wgigKsqo3_1;
	wire w_dff_A_25UuoGTf8_1;
	wire w_dff_A_70nrB0SL1_1;
	wire w_dff_A_s3CgOHqm4_1;
	wire w_dff_A_Xb2ovPJj1_1;
	wire w_dff_A_AU1BrwiZ6_1;
	wire w_dff_A_fczzsLAC1_1;
	wire w_dff_A_gnbRYeN84_1;
	wire w_dff_A_gKc0JG244_1;
	wire w_dff_A_SXTi0Hnn7_1;
	wire w_dff_A_pfcs9OfN8_1;
	wire w_dff_A_ypIElH5r9_1;
	wire w_dff_A_DhsNUEGQ8_2;
	wire w_dff_A_Q8iZl7Tt0_2;
	wire w_dff_A_FVuehxU57_2;
	wire w_dff_A_ur0vCEWL3_2;
	wire w_dff_A_eZRR2YPH3_2;
	wire w_dff_A_1x0zOaXT2_2;
	wire w_dff_A_iiorh9oP7_2;
	wire w_dff_A_BFrMIyUE7_2;
	wire w_dff_A_oeRkc5fA4_2;
	wire w_dff_A_b5aC0idQ3_2;
	wire w_dff_A_HU0MXQbV5_2;
	wire w_dff_A_BQt1wvsX2_2;
	wire w_dff_A_UJJOc4yD7_2;
	wire w_dff_B_5k3CBSX92_0;
	wire w_dff_A_4GlHeu0d9_1;
	wire w_dff_A_FZdUlzIc4_1;
	wire w_dff_A_8eFUU7KG9_1;
	wire w_dff_A_rOoHaY983_1;
	wire w_dff_A_pH0zxLsr9_1;
	wire w_dff_A_csgzIfQc0_0;
	wire w_dff_A_ozmYMCsi8_0;
	wire w_dff_A_YkHsRswo6_0;
	wire w_dff_A_bwUtO71m0_0;
	wire w_dff_A_3RpX77g78_0;
	wire w_dff_A_IRC0wbBQ1_0;
	wire w_dff_A_LZUBIv3c0_0;
	wire w_dff_A_gbEoHlYD1_0;
	wire w_dff_A_Zav5IAPQ4_0;
	wire w_dff_A_EuiKlArQ6_0;
	wire w_dff_A_ukI5AOSk4_0;
	wire w_dff_A_8d6iiiZY5_0;
	wire w_dff_A_8CCDWlrJ8_0;
	wire w_dff_B_4Zhg5uju9_1;
	wire w_dff_B_5bSR4sar3_1;
	wire w_dff_B_aE9ibtFv9_1;
	wire w_dff_B_LXkBdS2c5_1;
	wire w_dff_B_TzKsz0210_1;
	wire w_dff_B_9OUGm1OT6_1;
	wire w_dff_B_ffqh8P5m4_1;
	wire w_dff_A_u2o2vyNT8_0;
	wire w_dff_A_oFDmHfkx9_0;
	wire w_dff_A_Czeu6EaD2_0;
	wire w_dff_A_WGJgCACE1_0;
	wire w_dff_A_wtGrbgPE3_0;
	wire w_dff_A_1VKlLrV49_0;
	wire w_dff_A_fWOGl1ss9_0;
	wire w_dff_A_DrY94SJ54_0;
	wire w_dff_A_4UGFVwQa4_0;
	wire w_dff_A_uHjulb3A4_0;
	wire w_dff_A_ufPezCq83_0;
	wire w_dff_A_HYuZOdDo6_0;
	wire w_dff_A_o998TikY5_0;
	wire w_dff_A_zmSJXJog7_1;
	wire w_dff_A_3ic0lOvY4_1;
	wire w_dff_A_HDFCE9Ra2_1;
	wire w_dff_A_b3rBmTOY6_1;
	wire w_dff_A_aE22zqi41_1;
	wire w_dff_A_SPppKltk8_1;
	wire w_dff_A_Gosjnvc37_1;
	wire w_dff_A_8tObnMCA4_1;
	wire w_dff_A_v6NCN8Ps2_0;
	wire w_dff_A_jRWMkcb75_0;
	wire w_dff_A_OUGX0bC37_0;
	wire w_dff_A_PynhZ6tm3_0;
	wire w_dff_A_3Viobn0g9_0;
	wire w_dff_A_5YzlYxxv2_0;
	wire w_dff_A_srRqU8ZK1_0;
	wire w_dff_A_vzpAS6T33_0;
	wire w_dff_A_RJhHZLGL4_0;
	wire w_dff_A_2TzZKNIi4_0;
	wire w_dff_A_6Eh1bGgI3_0;
	wire w_dff_A_rw37N18g7_0;
	wire w_dff_A_Z82C6c1h0_0;
	wire w_dff_A_g9BeVl5L8_0;
	wire w_dff_A_oMLDARsX4_0;
	wire w_dff_A_Tlez3jKg0_0;
	wire w_dff_A_wkJiHxiJ2_0;
	wire w_dff_A_nN3psxv05_0;
	wire w_dff_A_ZjkH1l7G1_0;
	wire w_dff_A_LuWWhUkT2_0;
	wire w_dff_A_45KJcNxX6_0;
	wire w_dff_A_NtwJQERd5_2;
	wire w_dff_A_9Xpsc3pP8_2;
	wire w_dff_A_TH3MORgO4_2;
	wire w_dff_A_cEHnoUO15_2;
	wire w_dff_A_o2iQjXpM8_2;
	wire w_dff_A_pBNECicw9_2;
	wire w_dff_A_MeAqEvjp5_2;
	wire w_dff_A_m4Ae2IwH6_2;
	wire w_dff_A_Z1NYtCaj8_0;
	wire w_dff_A_xPS0zrTu1_0;
	wire w_dff_A_CSPzgjIt2_0;
	wire w_dff_A_iUMSITCT7_0;
	wire w_dff_A_IkwzG5A59_0;
	wire w_dff_A_9PWh6pjL1_0;
	wire w_dff_A_vFMq1rc39_0;
	wire w_dff_A_eeQFhTtw6_0;
	wire w_dff_A_CzzW6dEP2_0;
	wire w_dff_A_Jbgo1zMS7_0;
	wire w_dff_A_uuYeohou6_0;
	wire w_dff_B_D4Uj3POd5_2;
	wire w_dff_B_jBOghPDW2_2;
	wire w_dff_B_EnVZQBKX5_2;
	wire w_dff_B_wIHAtp7e7_2;
	wire w_dff_B_ay4QpemX4_2;
	wire w_dff_B_rJT8FTI67_2;
	wire w_dff_B_KjPWA0K59_2;
	wire w_dff_A_mpdH62qh1_0;
	wire w_dff_A_LWPdWuu84_0;
	wire w_dff_A_ZgUd1Aqt4_0;
	wire w_dff_A_eHl7k7d01_0;
	wire w_dff_A_Y8Z93HIb2_0;
	wire w_dff_A_q6CIHo5f9_0;
	wire w_dff_A_6smhHEjT0_0;
	wire w_dff_A_KV79Bzcm5_0;
	wire w_dff_A_dTKI1MBX9_0;
	wire w_dff_A_LAsYhJGn5_0;
	wire w_dff_A_SWVyRYqy8_0;
	wire w_dff_A_cnDCD1Ii8_0;
	wire w_dff_A_y9vALicB7_0;
	wire w_dff_A_a3vxG4wM6_1;
	wire w_dff_A_O3xE5l1p0_1;
	wire w_dff_A_5qN9hEe05_1;
	wire w_dff_A_4ppkeQfq3_1;
	wire w_dff_A_axWTm94x0_1;
	wire w_dff_A_tAjaqahn7_1;
	wire w_dff_A_u4zUTZK49_1;
	wire w_dff_A_jPiuEvLn5_1;
	wire w_dff_B_3q3uJTXK0_1;
	wire w_dff_B_Webltddt5_1;
	wire w_dff_B_OMjQFVzL0_1;
	wire w_dff_B_rDK8Seyi0_1;
	wire w_dff_B_yOtpg76R4_1;
	wire w_dff_B_rXtq5zsS2_1;
	wire w_dff_B_qdZUrO3T3_1;
	wire w_dff_A_JQEkHYdL3_0;
	wire w_dff_A_GWKBBymA1_0;
	wire w_dff_A_cmp2ENYx3_0;
	wire w_dff_A_xUSZTpTH2_0;
	wire w_dff_A_IWEqc1R23_0;
	wire w_dff_A_TbvIWBjq9_0;
	wire w_dff_A_1DRn7nos2_0;
	wire w_dff_A_rNQHft9w8_0;
	wire w_dff_A_GtNESeLD1_1;
	wire w_dff_A_aQ06KyK50_1;
	wire w_dff_A_ddpr6iII0_1;
	wire w_dff_A_T2CNLzLk1_1;
	wire w_dff_A_YAoRYpXC9_1;
	wire w_dff_A_5Fwu2crh3_1;
	wire w_dff_A_VrpypLOt1_1;
	wire w_dff_A_Bhr7B5352_1;
	wire w_dff_A_Q2IWkCYc1_1;
	wire w_dff_A_nouaKRpp6_1;
	wire w_dff_A_R4Oqs7rj8_1;
	wire w_dff_A_h0YrqkuB4_1;
	wire w_dff_A_pePc5qPA2_1;
	wire w_dff_A_rcvFle4e1_0;
	wire w_dff_A_cEkoftK35_0;
	wire w_dff_A_eHAKwe5L3_0;
	wire w_dff_A_FDVUoyVr7_0;
	wire w_dff_A_Ge5QTCjz0_0;
	wire w_dff_A_adLR2nLQ3_0;
	wire w_dff_A_R7AqDXEe5_0;
	wire w_dff_A_86vIatVO8_0;
	wire w_dff_A_UBAAwaDD8_0;
	wire w_dff_A_bVLVR48x8_0;
	wire w_dff_A_9ffzE9Xe7_0;
	wire w_dff_B_PzTm6c3O2_2;
	wire w_dff_B_i36PFyDq2_2;
	wire w_dff_B_9ptiehQW1_2;
	wire w_dff_B_XuIelDCn7_2;
	wire w_dff_B_bpY9c6ax3_2;
	wire w_dff_B_afBjiZUz2_2;
	wire w_dff_B_QCuW35tF1_2;
	wire w_dff_A_SZC6wqwR3_0;
	wire w_dff_A_M1ayiIXN7_0;
	wire w_dff_A_wo1WZE3S5_0;
	wire w_dff_A_wk4O4tJM6_0;
	wire w_dff_A_ILSV9DuX4_0;
	wire w_dff_A_aZLPuYJc0_0;
	wire w_dff_A_9aJeOWYx5_0;
	wire w_dff_A_EXY3HEom4_0;
	wire w_dff_A_MCDfcXLz8_0;
	wire w_dff_A_MNCvkhyj0_0;
	wire w_dff_A_14vY5lFt3_0;
	wire w_dff_A_pIJhu4c47_0;
	wire w_dff_A_J7Ni8DGh5_0;
	wire w_dff_A_utQirwwC3_1;
	wire w_dff_A_AxrFN8I25_1;
	wire w_dff_A_GFC64FIF3_1;
	wire w_dff_A_ZBIECQ5C5_1;
	wire w_dff_A_NEOCZtZ75_1;
	wire w_dff_A_DA87H3Es4_1;
	wire w_dff_A_ElfvlMue3_1;
	wire w_dff_A_Y58ckHoR2_1;
	wire w_dff_A_ekFSqqlX4_0;
	wire w_dff_A_tjMdoZay6_0;
	wire w_dff_A_cY4WZPW24_0;
	wire w_dff_A_YDql6qcL0_0;
	wire w_dff_A_IbwO6GSw7_0;
	wire w_dff_A_llwuIglX9_0;
	wire w_dff_B_yXaZP9Tk3_1;
	wire w_dff_B_GeUr3TFo8_1;
	wire w_dff_A_Q2lTggFU9_0;
	wire w_dff_A_AzQ8sAxq0_0;
	wire w_dff_A_1MF7ElMj4_0;
	wire w_dff_A_UNXucoXh5_0;
	wire w_dff_A_9wFwPlxX5_0;
	wire w_dff_A_LSQjTqpw4_0;
	wire w_dff_A_ZraDmxQ62_0;
	wire w_dff_A_Mio5T8Af3_0;
	wire w_dff_A_iYztd4Bf1_0;
	wire w_dff_A_lAR0vVB73_0;
	wire w_dff_A_iipd2KGQ2_0;
	wire w_dff_A_dhXW7ami4_0;
	wire w_dff_A_SWdrrLUX9_0;
	wire w_dff_A_Gqm0Tpox9_0;
	wire w_dff_A_rFfxckqV0_0;
	wire w_dff_A_JFhLedmD3_0;
	wire w_dff_A_4JRnfKCw4_0;
	wire w_dff_A_ZhhdXqXN7_0;
	wire w_dff_A_n3iobooB0_0;
	wire w_dff_A_H0FUpJj18_0;
	wire w_dff_A_9Wf5qaaL2_0;
	wire w_dff_A_oJCepPFk1_0;
	wire w_dff_A_xqO1nsWH4_0;
	wire w_dff_A_oDIYdEqg1_0;
	wire w_dff_A_ukL3jJRl9_0;
	wire w_dff_A_30SHR6zx5_0;
	wire w_dff_A_uWAAZltc2_0;
	wire w_dff_A_MPNdGI4x0_0;
	wire w_dff_A_D6BiZbl03_0;
	wire w_dff_A_jEQzpy3Y2_0;
	wire w_dff_A_ZYDcdArH4_0;
	wire w_dff_A_UMv943f01_0;
	wire w_dff_A_oQNsq2z73_0;
	wire w_dff_A_8dZ7FzZd5_0;
	wire w_dff_A_gVLds06A3_0;
	wire w_dff_A_HHCjlAO74_0;
	wire w_dff_A_bVddjTpq9_0;
	wire w_dff_A_IKCO1RKT1_0;
	wire w_dff_A_em9DAxQv6_0;
	wire w_dff_A_W85tryrl8_0;
	wire w_dff_A_XdMtB1fP9_0;
	wire w_dff_A_9G8u8If34_0;
	wire w_dff_A_5fIA5fmE1_0;
	wire w_dff_A_dQi7a2mO7_0;
	wire w_dff_A_LNNNHOMc6_0;
	wire w_dff_A_i3wfzIfI6_0;
	wire w_dff_A_qpbGa8nT5_0;
	wire w_dff_A_IMUSR4iz5_0;
	wire w_dff_A_wrwXWCbl9_0;
	wire w_dff_A_kqsSluya0_0;
	wire w_dff_A_nB5OHnJe9_0;
	wire w_dff_A_t5V3gYZH1_0;
	wire w_dff_A_DJwjTZyo0_0;
	wire w_dff_A_yBuIrjD62_0;
	wire w_dff_A_idV8RLow4_0;
	wire w_dff_B_eLiWCHHm6_2;
	wire w_dff_B_dh1QZYeF1_2;
	wire w_dff_B_CjY5rhLe9_2;
	wire w_dff_B_wj4h2j8T3_2;
	wire w_dff_B_vZoE3AT62_2;
	wire w_dff_B_9RWjf2qb1_2;
	wire w_dff_B_YvfeFDYf2_2;
	wire w_dff_A_i6bLeDAc4_0;
	wire w_dff_A_vC4L3q7D1_0;
	wire w_dff_A_KawixPpr7_0;
	wire w_dff_A_wqbPpEsF5_0;
	wire w_dff_A_Co7XTYEZ5_0;
	wire w_dff_A_gSWVosat9_0;
	wire w_dff_A_kRHPQ6DL8_0;
	wire w_dff_A_wSdM53il8_0;
	wire w_dff_A_ejcjulET7_0;
	wire w_dff_A_EW5RCved3_0;
	wire w_dff_A_vh36FAp74_0;
	wire w_dff_A_TRI6dzrh9_0;
	wire w_dff_A_2vpsb4yq7_0;
	wire w_dff_A_crKarmKn2_1;
	wire w_dff_A_3zKzzX0o9_1;
	wire w_dff_A_XloKwHC65_1;
	wire w_dff_A_6R0rSIKA8_1;
	wire w_dff_A_wwSvJ7zs2_1;
	wire w_dff_A_21dRWtTN0_1;
	wire w_dff_A_ke5TfXVn5_1;
	wire w_dff_A_JXS19OY08_1;
	wire w_dff_A_4vVSVNWb9_1;
	wire w_dff_A_pF42VPeW3_1;
	wire w_dff_A_wXbEfXpi6_1;
	wire w_dff_A_81SzDoTd9_1;
	wire w_dff_A_8Q4eDf5T1_1;
	wire w_dff_A_fT9wljA27_1;
	wire w_dff_B_MZVBPHjq7_1;
	wire w_dff_B_kYIEF2aV8_1;
	wire w_dff_A_1vJ2ygwZ1_0;
	wire w_dff_A_6RBbb3pF8_0;
	wire w_dff_A_QL0JVbtg7_0;
	wire w_dff_A_zN7L9Xib5_0;
	wire w_dff_A_P4LtSjGT5_0;
	wire w_dff_A_qsw5L1xA1_0;
	wire w_dff_A_FJepJW0D0_0;
	wire w_dff_A_tllPJFyQ9_2;
	wire w_dff_A_aFNVmE5J3_0;
	wire w_dff_A_q9UiaNJr3_0;
	wire w_dff_A_GWRWYNmk2_0;
	wire w_dff_A_W7duW0aV2_0;
	wire w_dff_A_yDrnNUkO3_0;
	wire w_dff_A_F3BcyRrH7_0;
	wire w_dff_A_ANIxLGii8_0;
	wire w_dff_A_mKfXLHxv0_0;
	wire w_dff_A_iBwruxZa9_0;
	wire w_dff_A_KWdeIHcj1_0;
	wire w_dff_A_uyyDderI0_0;
	wire w_dff_A_hOBi2wgc9_1;
	wire w_dff_A_GSIA5rLJ5_0;
	wire w_dff_A_723ZUFy59_0;
	wire w_dff_A_q5Fur47B7_0;
	wire w_dff_A_LbHL6NVU9_0;
	wire w_dff_A_bTB9zVMv4_0;
	wire w_dff_A_xEJAJHoi6_0;
	wire w_dff_A_GL4kS4WD9_0;
	wire w_dff_A_J6MpdPul1_0;
	wire w_dff_A_4pCo5JOC1_0;
	wire w_dff_A_lq3ZaFkm9_0;
	wire w_dff_A_vkNPP3Cd8_0;
	wire w_dff_A_h9q6CtEl3_1;
	wire w_dff_A_eYpRitAm5_0;
	wire w_dff_A_19lApDpL0_0;
	wire w_dff_A_CI2VMVur5_0;
	wire w_dff_A_4Lsd1Qer8_0;
	wire w_dff_A_56joeSDb3_0;
	wire w_dff_A_L7JyQjFO9_0;
	wire w_dff_A_Qc6vKUw11_0;
	wire w_dff_A_8P84km3w1_2;
	wire w_dff_A_r6nconcD2_0;
	wire w_dff_A_qmWZ6wVP1_0;
	wire w_dff_A_mlZFzwlZ2_0;
	wire w_dff_A_heu4L1Ns7_0;
	wire w_dff_A_gGvRmQIr2_0;
	wire w_dff_A_16be6FTn1_0;
	wire w_dff_A_z53fshU91_0;
	wire w_dff_A_eiLlJu3o9_0;
	wire w_dff_A_nwM5npPn8_0;
	wire w_dff_A_D9EtDKU45_0;
	wire w_dff_A_5wj2Tdsz1_0;
	wire w_dff_A_XzzsQ4iL7_1;
	wire w_dff_A_7kEGWqiZ8_0;
	wire w_dff_A_gROs3v982_0;
	wire w_dff_A_D2f2dGQv1_0;
	wire w_dff_A_iN9Vgaa21_0;
	wire w_dff_A_xgzCq0VH2_0;
	wire w_dff_A_R4XptZOV1_0;
	wire w_dff_A_VPLfegx98_0;
	wire w_dff_A_qB1wV2iS1_2;
	wire w_dff_A_Q9A4t4oZ2_0;
	wire w_dff_A_ijNO9qvH3_0;
	wire w_dff_A_6qP1UmU47_0;
	wire w_dff_A_ebFzpK3i2_0;
	wire w_dff_A_bpBTlwkC8_0;
	wire w_dff_A_U1eOvkav8_0;
	wire w_dff_A_mi5VXx440_0;
	wire w_dff_A_wz2EMHLE2_0;
	wire w_dff_A_WshWNZHf5_0;
	wire w_dff_A_HHmNheJy3_0;
	wire w_dff_A_AQOtljhc9_0;
	wire w_dff_A_MKhlq43s3_1;
	wire w_dff_A_6bT09feS3_0;
	wire w_dff_A_TLeHMkFY5_0;
	wire w_dff_A_o8nSjWMa0_0;
	wire w_dff_A_nTkSz7U96_0;
	wire w_dff_A_yA2vNyT90_0;
	wire w_dff_A_snST9etI2_0;
	wire w_dff_A_x6jLjakQ4_0;
	wire w_dff_A_H1t0GsEX5_2;
	wire w_dff_A_8WrG7YFw8_0;
	wire w_dff_A_LdgkSa4K8_0;
	wire w_dff_A_TDApIbAT0_0;
	wire w_dff_A_cutebYfY3_0;
	wire w_dff_A_ivBejZGA4_0;
	wire w_dff_A_ywGF07Yt5_0;
	wire w_dff_A_Mh2jNOs57_0;
	wire w_dff_A_AJfO7qUL3_0;
	wire w_dff_A_wajLPQZG6_0;
	wire w_dff_A_R19Yk38P5_0;
	wire w_dff_A_N0thLyMm9_0;
	wire w_dff_A_XJYSseO16_1;
	wire w_dff_A_gFEi0ILJ0_0;
	wire w_dff_A_L5ZhjltH9_0;
	wire w_dff_A_btfbrcGR5_0;
	wire w_dff_A_AD4OIk8E3_0;
	wire w_dff_A_9MNA8pJX2_1;
	wire w_dff_A_p2oaRg9A0_1;
	wire w_dff_A_XkeiPx5T6_2;
	wire w_dff_A_YLBqApx23_0;
	wire w_dff_A_5Clu7xMq9_0;
	wire w_dff_A_3BxagBXD6_0;
	wire w_dff_A_P8dVwl946_0;
	wire w_dff_A_LZjoW5Q68_0;
	wire w_dff_A_ZmRpUAqN5_0;
	wire w_dff_A_Il4LI20s8_1;
	wire w_dff_A_673eak7Z5_0;
	wire w_dff_A_JPTUn46c8_0;
	wire w_dff_A_xtCuV8GB0_0;
	wire w_dff_A_ptLf8Aei8_0;
	wire w_dff_A_DY5M21Eq8_0;
	wire w_dff_A_lE9BPisZ9_0;
	wire w_dff_A_bC3ynXnv7_0;
	wire w_dff_A_9GN6vBZw5_2;
	wire w_dff_A_6cZUH2EU9_0;
	wire w_dff_A_wISLR8sa1_0;
	wire w_dff_A_G0wiSCUW8_0;
	wire w_dff_A_3FZBqs5V4_0;
	wire w_dff_A_4sFDhFEl2_0;
	wire w_dff_A_NwJ9YEFb4_0;
	wire w_dff_A_PYGxBhqM6_0;
	wire w_dff_A_35RAxjnE0_0;
	wire w_dff_A_r117srsO3_0;
	wire w_dff_A_oCqD4GS20_0;
	wire w_dff_A_HkqsB3iX6_0;
	wire w_dff_A_FoogvTwZ9_1;
	wire w_dff_A_r7zmGIrz2_1;
	wire w_dff_A_jsqxPSei4_0;
	wire w_dff_A_hLMVnkT17_1;
	wire w_dff_A_owbfHAUL9_1;
	wire w_dff_A_GaW1e9fz9_1;
	wire w_dff_A_dSE75Enq1_1;
	wire w_dff_A_4hZwDtfK5_1;
	wire w_dff_A_gEgxyzuw3_1;
	wire w_dff_A_OMt7C9BY0_1;
	wire w_dff_A_Oq19nnOW7_1;
	wire w_dff_A_0LFFT8AU3_2;
	wire w_dff_A_cLHpH9ki5_0;
	wire w_dff_A_tzaD2OSm9_0;
	wire w_dff_A_zRYPA6M31_0;
	wire w_dff_A_NXNV4o3y8_0;
	wire w_dff_A_60Isjg0p8_0;
	wire w_dff_A_WYlnxJGX6_0;
	wire w_dff_A_LnK4VPRl1_0;
	wire w_dff_A_BHxn3vWE5_0;
	wire w_dff_A_QoauDusf9_0;
	wire w_dff_A_lMTmNFar2_0;
	wire w_dff_A_IwzqA2iF0_0;
	wire w_dff_A_nFiQWkQe2_0;
	wire w_dff_A_02sEIOQc0_0;
	wire w_dff_A_CQV93wuJ5_0;
	wire w_dff_A_2Rh298mt6_0;
	wire w_dff_A_8LxJD7Ka4_0;
	wire w_dff_A_98SxYP9q9_0;
	wire w_dff_A_R7wHTQLs5_0;
	wire w_dff_A_8Lbhp4gN7_0;
	wire w_dff_A_grhwHU0Q5_0;
	wire w_dff_A_GBMHBtLC7_0;
	wire w_dff_A_Ef0k35ne1_0;
	wire w_dff_A_u40iQJzv7_0;
	wire w_dff_A_6YUz5bTd3_0;
	wire w_dff_A_ArKlI0YR1_2;
	wire w_dff_A_yDeajRKO1_1;
	wire w_dff_A_q5Bwaxhn3_1;
	wire w_dff_A_yCPbTmvH4_1;
	wire w_dff_A_FnpqAHZ88_1;
	wire w_dff_A_qrGkmUSR3_1;
	wire w_dff_A_DpwkpF1e4_1;
	wire w_dff_A_uih7FaRx8_1;
	wire w_dff_A_cKzUmcT47_1;
	wire w_dff_A_KEF28kuZ3_1;
	wire w_dff_A_VlnhQV3B0_1;
	wire w_dff_A_4g6tQ1Jv2_1;
	wire w_dff_A_UkQF1isM7_1;
	wire w_dff_A_CoyOhJqe6_1;
	wire w_dff_A_Wp6m8flR3_1;
	wire w_dff_A_vzdET3bI2_1;
	wire w_dff_A_UpkpSmaE9_2;
	wire w_dff_A_FU6nqaMn8_0;
	wire w_dff_A_ZURtT3z48_0;
	wire w_dff_A_yWwXl4Ia8_0;
	wire w_dff_A_5KR7nyzA4_0;
	wire w_dff_A_TrpIRjTs6_0;
	wire w_dff_A_IH2i5YbZ3_0;
	wire w_dff_A_ojReUlWs0_0;
	wire w_dff_A_36M7VTwQ0_0;
	wire w_dff_A_6GJIz99K7_0;
	wire w_dff_A_g0bsMIUw6_0;
	wire w_dff_A_NBxdbV2b0_0;
	wire w_dff_A_LJAVZiyt7_0;
	wire w_dff_A_mCfbOrl39_0;
	wire w_dff_A_LnD9suQ63_0;
	wire w_dff_A_Pp9RYpVK6_0;
	wire w_dff_A_cpRx40lW9_0;
	wire w_dff_A_BYjuNU6O1_0;
	wire w_dff_A_HiA6zjCe3_0;
	wire w_dff_A_jHFVsp219_0;
	wire w_dff_A_Bu8Xx7qr6_1;
	wire w_dff_A_z0cbYEHf0_0;
	wire w_dff_A_icsYvCzl6_0;
	wire w_dff_A_SbCTtuPm8_0;
	wire w_dff_A_TCDSmcrq1_0;
	wire w_dff_A_2SlUWncV3_0;
	wire w_dff_A_7bG7OGGA5_0;
	wire w_dff_A_wy2ulCCa7_0;
	wire w_dff_A_G5HuG4MA3_0;
	wire w_dff_A_BD5BVYR26_0;
	wire w_dff_A_a1lcWSP85_0;
	wire w_dff_A_cJDUwa1p0_0;
	wire w_dff_A_Ogb9wPl73_0;
	wire w_dff_A_LssHnvSR5_1;
	wire w_dff_A_PgaZ1PXA1_0;
	wire w_dff_A_817POFMo8_0;
	wire w_dff_A_R5xiUOs84_0;
	wire w_dff_A_ZuERHQ0J4_0;
	wire w_dff_A_pOZByUTb2_0;
	wire w_dff_A_vdAnjuUY2_1;
	wire w_dff_A_OmxKvbDF0_0;
	jnot g000(.din(w_G76gat_0[1]),.dout(n43),.clk(gclk));
	jand g001(.dina(w_G82gat_0[2]),.dinb(w_n43_0[1]),.dout(n44),.clk(gclk));
	jnot g002(.din(w_G24gat_0[1]),.dout(n45),.clk(gclk));
	jand g003(.dina(w_G30gat_0[1]),.dinb(n45),.dout(n46),.clk(gclk));
	jnot g004(.din(w_G11gat_0[2]),.dout(n47),.clk(gclk));
	jand g005(.dina(w_G17gat_0[2]),.dinb(w_n47_0[1]),.dout(n48),.clk(gclk));
	jor g006(.dina(n48),.dinb(n46),.dout(n49),.clk(gclk));
	jor g007(.dina(n49),.dinb(w_n44_0[1]),.dout(n50),.clk(gclk));
	jnot g008(.din(w_G37gat_0[2]),.dout(n51),.clk(gclk));
	jand g009(.dina(w_G43gat_1[1]),.dinb(n51),.dout(n52),.clk(gclk));
	jnot g010(.din(w_G63gat_0[2]),.dout(n53),.clk(gclk));
	jand g011(.dina(w_G69gat_0[2]),.dinb(w_n53_0[1]),.dout(n54),.clk(gclk));
	jor g012(.dina(n54),.dinb(w_n52_0[1]),.dout(n55),.clk(gclk));
	jnot g013(.din(w_G102gat_0[2]),.dout(n56),.clk(gclk));
	jand g014(.dina(w_G108gat_0[2]),.dinb(w_n56_0[1]),.dout(n57),.clk(gclk));
	jnot g015(.din(w_G50gat_0[2]),.dout(n58),.clk(gclk));
	jand g016(.dina(w_G56gat_0[2]),.dinb(w_n58_0[1]),.dout(n59),.clk(gclk));
	jor g017(.dina(n59),.dinb(n57),.dout(n60),.clk(gclk));
	jnot g018(.din(w_G89gat_0[2]),.dout(n61),.clk(gclk));
	jand g019(.dina(w_G95gat_0[2]),.dinb(w_n61_0[1]),.dout(n62),.clk(gclk));
	jnot g020(.din(w_G1gat_0[2]),.dout(n63),.clk(gclk));
	jand g021(.dina(w_G4gat_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jor g022(.dina(n64),.dinb(n62),.dout(n65),.clk(gclk));
	jor g023(.dina(n65),.dinb(n60),.dout(n66),.clk(gclk));
	jor g024(.dina(n66),.dinb(w_dff_B_kYIEF2aV8_1),.dout(n67),.clk(gclk));
	jor g025(.dina(n67),.dinb(w_dff_B_MZVBPHjq7_1),.dout(G223gat_fa_),.clk(gclk));
	jnot g026(.din(w_G112gat_0[2]),.dout(n69),.clk(gclk));
	jnot g027(.din(w_n44_0[0]),.dout(n70),.clk(gclk));
	jnot g028(.din(w_G30gat_0[0]),.dout(n71),.clk(gclk));
	jor g029(.dina(w_n71_0[1]),.dinb(w_G24gat_0[0]),.dout(n72),.clk(gclk));
	jnot g030(.din(w_G17gat_0[1]),.dout(n73),.clk(gclk));
	jor g031(.dina(w_n73_0[1]),.dinb(w_G11gat_0[1]),.dout(n74),.clk(gclk));
	jand g032(.dina(n74),.dinb(w_n72_0[1]),.dout(n75),.clk(gclk));
	jand g033(.dina(n75),.dinb(n70),.dout(n76),.clk(gclk));
	jnot g034(.din(w_G43gat_1[0]),.dout(n77),.clk(gclk));
	jor g035(.dina(w_n77_0[1]),.dinb(w_G37gat_0[1]),.dout(n78),.clk(gclk));
	jnot g036(.din(w_G69gat_0[1]),.dout(n79),.clk(gclk));
	jor g037(.dina(w_n79_0[1]),.dinb(w_G63gat_0[1]),.dout(n80),.clk(gclk));
	jand g038(.dina(n80),.dinb(w_n78_0[1]),.dout(n81),.clk(gclk));
	jnot g039(.din(w_G108gat_0[1]),.dout(n82),.clk(gclk));
	jor g040(.dina(w_n82_0[1]),.dinb(w_G102gat_0[1]),.dout(n83),.clk(gclk));
	jnot g041(.din(w_G56gat_0[1]),.dout(n84),.clk(gclk));
	jor g042(.dina(w_n84_0[1]),.dinb(w_G50gat_0[1]),.dout(n85),.clk(gclk));
	jand g043(.dina(n85),.dinb(n83),.dout(n86),.clk(gclk));
	jnot g044(.din(w_G95gat_0[1]),.dout(n87),.clk(gclk));
	jor g045(.dina(w_n87_0[1]),.dinb(w_G89gat_0[1]),.dout(n88),.clk(gclk));
	jnot g046(.din(w_G4gat_0[1]),.dout(n89),.clk(gclk));
	jor g047(.dina(w_n89_0[1]),.dinb(w_G1gat_0[1]),.dout(n90),.clk(gclk));
	jand g048(.dina(n90),.dinb(n88),.dout(n91),.clk(gclk));
	jand g049(.dina(n91),.dinb(n86),.dout(n92),.clk(gclk));
	jand g050(.dina(n92),.dinb(w_dff_B_GeUr3TFo8_1),.dout(n93),.clk(gclk));
	jand g051(.dina(n93),.dinb(w_dff_B_yXaZP9Tk3_1),.dout(n94),.clk(gclk));
	jor g052(.dina(w_n94_4[1]),.dinb(w_n56_0[0]),.dout(n95),.clk(gclk));
	jand g053(.dina(n95),.dinb(w_G108gat_0[0]),.dout(n96),.clk(gclk));
	jand g054(.dina(w_n96_0[1]),.dinb(w_n69_0[1]),.dout(n97),.clk(gclk));
	jnot g055(.din(w_G8gat_0[2]),.dout(n98),.clk(gclk));
	jor g056(.dina(w_n94_4[0]),.dinb(w_n63_0[0]),.dout(n99),.clk(gclk));
	jand g057(.dina(n99),.dinb(w_G4gat_0[0]),.dout(n100),.clk(gclk));
	jand g058(.dina(w_n100_0[1]),.dinb(w_n98_0[1]),.dout(n101),.clk(gclk));
	jor g059(.dina(n101),.dinb(n97),.dout(n102),.clk(gclk));
	jnot g060(.din(w_G99gat_0[2]),.dout(n103),.clk(gclk));
	jor g061(.dina(w_n94_3[2]),.dinb(w_n61_0[0]),.dout(n104),.clk(gclk));
	jand g062(.dina(n104),.dinb(w_G95gat_0[0]),.dout(n105),.clk(gclk));
	jand g063(.dina(n105),.dinb(w_dff_B_qdZUrO3T3_1),.dout(n106),.clk(gclk));
	jnot g064(.din(w_G73gat_0[2]),.dout(n107),.clk(gclk));
	jor g065(.dina(w_n94_3[1]),.dinb(w_n53_0[0]),.dout(n108),.clk(gclk));
	jand g066(.dina(n108),.dinb(w_G69gat_0[0]),.dout(n109),.clk(gclk));
	jand g067(.dina(w_n109_0[1]),.dinb(w_n107_0[1]),.dout(n110),.clk(gclk));
	jor g068(.dina(n110),.dinb(n106),.dout(n111),.clk(gclk));
	jor g069(.dina(n111),.dinb(n102),.dout(n112),.clk(gclk));
	jxor g070(.dina(w_n94_3[0]),.dinb(w_n72_0[0]),.dout(n113),.clk(gclk));
	jor g071(.dina(n113),.dinb(w_n71_0[0]),.dout(n114),.clk(gclk));
	jor g072(.dina(w_n114_0[2]),.dinb(w_G34gat_0[2]),.dout(n115),.clk(gclk));
	jnot g073(.din(w_n115_0[1]),.dout(n116),.clk(gclk));
	jnot g074(.din(w_G60gat_0[2]),.dout(n117),.clk(gclk));
	jor g075(.dina(w_n94_2[2]),.dinb(w_n58_0[0]),.dout(n118),.clk(gclk));
	jand g076(.dina(n118),.dinb(w_G56gat_0[0]),.dout(n119),.clk(gclk));
	jand g077(.dina(w_n119_0[1]),.dinb(w_dff_B_ffqh8P5m4_1),.dout(n120),.clk(gclk));
	jxor g078(.dina(w_n94_2[1]),.dinb(w_n52_0[0]),.dout(n121),.clk(gclk));
	jnot g079(.din(w_G47gat_0[1]),.dout(n122),.clk(gclk));
	jand g080(.dina(n122),.dinb(w_G43gat_0[2]),.dout(n123),.clk(gclk));
	jand g081(.dina(w_n123_0[1]),.dinb(w_n121_0[1]),.dout(n124),.clk(gclk));
	jor g082(.dina(w_dff_B_5k3CBSX92_0),.dinb(n120),.dout(n125),.clk(gclk));
	jnot g083(.din(w_G86gat_1[1]),.dout(n126),.clk(gclk));
	jor g084(.dina(w_n94_2[0]),.dinb(w_n43_0[0]),.dout(n127),.clk(gclk));
	jand g085(.dina(n127),.dinb(w_G82gat_0[1]),.dout(n128),.clk(gclk));
	jand g086(.dina(w_n128_0[1]),.dinb(w_n126_0[2]),.dout(n129),.clk(gclk));
	jnot g087(.din(w_G21gat_1[1]),.dout(n130),.clk(gclk));
	jor g088(.dina(w_n94_1[2]),.dinb(w_n47_0[0]),.dout(n131),.clk(gclk));
	jand g089(.dina(n131),.dinb(w_G17gat_0[0]),.dout(n132),.clk(gclk));
	jand g090(.dina(w_n132_0[1]),.dinb(w_n130_0[2]),.dout(n133),.clk(gclk));
	jor g091(.dina(n133),.dinb(n129),.dout(n134),.clk(gclk));
	jor g092(.dina(n134),.dinb(n125),.dout(n135),.clk(gclk));
	jor g093(.dina(n135),.dinb(w_dff_B_W4NMkniy8_1),.dout(n136),.clk(gclk));
	jor g094(.dina(n136),.dinb(w_dff_B_FO7OnCup9_1),.dout(G329gat_fa_),.clk(gclk));
	jand g095(.dina(w_G223gat_3[1]),.dinb(w_G89gat_0[0]),.dout(n138),.clk(gclk));
	jor g096(.dina(n138),.dinb(w_n87_0[0]),.dout(n139),.clk(gclk));
	jand g097(.dina(w_G329gat_6),.dinb(w_G99gat_0[1]),.dout(n140),.clk(gclk));
	jor g098(.dina(n140),.dinb(w_n139_0[1]),.dout(n141),.clk(gclk));
	jor g099(.dina(w_n141_0[1]),.dinb(w_G105gat_0[1]),.dout(n142),.clk(gclk));
	jnot g100(.din(w_n142_0[1]),.dout(n143),.clk(gclk));
	jand g101(.dina(w_G223gat_3[0]),.dinb(w_G50gat_0[0]),.dout(n144),.clk(gclk));
	jor g102(.dina(n144),.dinb(w_n84_0[0]),.dout(n145),.clk(gclk));
	jor g103(.dina(w_n145_0[1]),.dinb(w_G60gat_0[1]),.dout(n146),.clk(gclk));
	jand g104(.dina(w_G329gat_5[2]),.dinb(w_n146_0[1]),.dout(n147),.clk(gclk));
	jnot g105(.din(w_n147_0[1]),.dout(n148),.clk(gclk));
	jnot g106(.din(w_G66gat_0[1]),.dout(n150),.clk(gclk));
	jand g107(.dina(w_n119_0[0]),.dinb(w_n150_0[1]),.dout(n151),.clk(gclk));
	jand g108(.dina(w_n151_0[1]),.dinb(n148),.dout(n153),.clk(gclk));
	jnot g109(.din(w_G79gat_0[1]),.dout(n154),.clk(gclk));
	jand g110(.dina(w_G223gat_2[2]),.dinb(w_G102gat_0[0]),.dout(n155),.clk(gclk));
	jor g111(.dina(n155),.dinb(w_n82_0[0]),.dout(n156),.clk(gclk));
	jor g112(.dina(w_n156_0[1]),.dinb(w_G112gat_0[1]),.dout(n157),.clk(gclk));
	jand g113(.dina(w_G223gat_2[1]),.dinb(w_G1gat_0[0]),.dout(n158),.clk(gclk));
	jor g114(.dina(n158),.dinb(w_n89_0[0]),.dout(n159),.clk(gclk));
	jor g115(.dina(w_n159_0[1]),.dinb(w_G8gat_0[1]),.dout(n160),.clk(gclk));
	jand g116(.dina(n160),.dinb(n157),.dout(n161),.clk(gclk));
	jor g117(.dina(w_n139_0[0]),.dinb(w_G99gat_0[0]),.dout(n162),.clk(gclk));
	jand g118(.dina(w_G223gat_2[0]),.dinb(w_G63gat_0[0]),.dout(n163),.clk(gclk));
	jor g119(.dina(n163),.dinb(w_n79_0[0]),.dout(n164),.clk(gclk));
	jor g120(.dina(w_n164_0[1]),.dinb(w_G73gat_0[1]),.dout(n165),.clk(gclk));
	jand g121(.dina(n165),.dinb(n162),.dout(n166),.clk(gclk));
	jand g122(.dina(n166),.dinb(n161),.dout(n167),.clk(gclk));
	jxor g123(.dina(w_n94_1[1]),.dinb(w_n78_0[0]),.dout(n168),.clk(gclk));
	jnot g124(.din(w_n123_0[0]),.dout(n169),.clk(gclk));
	jor g125(.dina(w_dff_B_J5sydVXs4_0),.dinb(n168),.dout(n170),.clk(gclk));
	jand g126(.dina(w_n170_0[1]),.dinb(w_n146_0[0]),.dout(n171),.clk(gclk));
	jnot g127(.din(w_G82gat_0[0]),.dout(n172),.clk(gclk));
	jand g128(.dina(w_G223gat_1[2]),.dinb(w_G76gat_0[0]),.dout(n173),.clk(gclk));
	jor g129(.dina(n173),.dinb(w_dff_B_U5uq0R0n0_1),.dout(n174),.clk(gclk));
	jor g130(.dina(w_n174_0[1]),.dinb(w_G86gat_1[0]),.dout(n175),.clk(gclk));
	jand g131(.dina(w_G223gat_1[1]),.dinb(w_G11gat_0[0]),.dout(n176),.clk(gclk));
	jor g132(.dina(n176),.dinb(w_n73_0[0]),.dout(n177),.clk(gclk));
	jor g133(.dina(w_n177_0[1]),.dinb(w_G21gat_1[0]),.dout(n178),.clk(gclk));
	jand g134(.dina(n178),.dinb(n175),.dout(n179),.clk(gclk));
	jand g135(.dina(n179),.dinb(n171),.dout(n180),.clk(gclk));
	jand g136(.dina(n180),.dinb(w_n115_0[0]),.dout(n181),.clk(gclk));
	jand g137(.dina(n181),.dinb(w_dff_B_YUN2JMjJ6_1),.dout(n182),.clk(gclk));
	jor g138(.dina(w_n182_3[1]),.dinb(w_n107_0[0]),.dout(n183),.clk(gclk));
	jand g139(.dina(n183),.dinb(w_n109_0[0]),.dout(n184),.clk(gclk));
	jand g140(.dina(w_n184_0[1]),.dinb(w_n154_0[1]),.dout(n185),.clk(gclk));
	jor g141(.dina(n185),.dinb(n153),.dout(n186),.clk(gclk));
	jor g142(.dina(n186),.dinb(n143),.dout(n187),.clk(gclk));
	jand g143(.dina(w_G329gat_5[1]),.dinb(w_n170_0[0]),.dout(n188),.clk(gclk));
	jnot g144(.din(w_n188_0[1]),.dout(n189),.clk(gclk));
	jnot g145(.din(w_G53gat_0[1]),.dout(n191),.clk(gclk));
	jand g146(.dina(w_n191_0[1]),.dinb(w_G43gat_0[1]),.dout(n192),.clk(gclk));
	jand g147(.dina(w_dff_B_6ncqurZe4_0),.dinb(w_n121_0[0]),.dout(n193),.clk(gclk));
	jand g148(.dina(w_n193_0[1]),.dinb(n189),.dout(n195),.clk(gclk));
	jor g149(.dina(w_n182_3[0]),.dinb(w_n130_0[1]),.dout(n196),.clk(gclk));
	jand g150(.dina(n196),.dinb(w_n132_0[0]),.dout(n197),.clk(gclk));
	jnot g151(.din(w_G27gat_0[1]),.dout(n198),.clk(gclk));
	jor g152(.dina(w_G329gat_5[0]),.dinb(w_G21gat_0[2]),.dout(n199),.clk(gclk));
	jand g153(.dina(n199),.dinb(w_n198_0[1]),.dout(n200),.clk(gclk));
	jand g154(.dina(n200),.dinb(w_n197_0[1]),.dout(n201),.clk(gclk));
	jor g155(.dina(n201),.dinb(n195),.dout(n202),.clk(gclk));
	jor g156(.dina(w_n182_2[2]),.dinb(w_n126_0[1]),.dout(n203),.clk(gclk));
	jand g157(.dina(n203),.dinb(w_n128_0[0]),.dout(n204),.clk(gclk));
	jnot g158(.din(w_G92gat_0[2]),.dout(n205),.clk(gclk));
	jor g159(.dina(w_G329gat_4[2]),.dinb(w_G86gat_0[2]),.dout(n206),.clk(gclk));
	jand g160(.dina(n206),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jand g161(.dina(n207),.dinb(w_n204_0[1]),.dout(n208),.clk(gclk));
	jnot g162(.din(w_G14gat_0[2]),.dout(n209),.clk(gclk));
	jor g163(.dina(w_n182_2[1]),.dinb(w_n98_0[0]),.dout(n210),.clk(gclk));
	jand g164(.dina(n210),.dinb(w_n100_0[0]),.dout(n211),.clk(gclk));
	jand g165(.dina(n211),.dinb(w_dff_B_uTCzO6Hi1_1),.dout(n212),.clk(gclk));
	jor g166(.dina(n212),.dinb(n208),.dout(n213),.clk(gclk));
	jnot g167(.din(w_G34gat_0[1]),.dout(n214),.clk(gclk));
	jor g168(.dina(w_n182_2[0]),.dinb(w_dff_B_9ISUfuz87_1),.dout(n215),.clk(gclk));
	jnot g169(.din(w_G40gat_0[1]),.dout(n217),.clk(gclk));
	jnot g170(.din(w_n114_0[1]),.dout(n218),.clk(gclk));
	jand g171(.dina(n218),.dinb(w_n217_0[1]),.dout(n219),.clk(gclk));
	jand g172(.dina(w_n219_0[1]),.dinb(n215),.dout(n221),.clk(gclk));
	jnot g173(.din(w_G115gat_0[1]),.dout(n222),.clk(gclk));
	jor g174(.dina(w_n182_1[2]),.dinb(w_n69_0[0]),.dout(n223),.clk(gclk));
	jand g175(.dina(n223),.dinb(w_n96_0[0]),.dout(n224),.clk(gclk));
	jand g176(.dina(w_n224_0[1]),.dinb(w_n222_0[1]),.dout(n225),.clk(gclk));
	jor g177(.dina(n225),.dinb(w_dff_B_Lmvqt5U65_1),.dout(n226),.clk(gclk));
	jor g178(.dina(n226),.dinb(n213),.dout(n227),.clk(gclk));
	jor g179(.dina(n227),.dinb(w_dff_B_A6RWogJ76_1),.dout(n228),.clk(gclk));
	jor g180(.dina(n228),.dinb(w_dff_B_2TnlZEFq4_1),.dout(G370gat_fa_),.clk(gclk));
	jand g181(.dina(w_G329gat_4[1]),.dinb(w_G8gat_0[0]),.dout(n230),.clk(gclk));
	jor g182(.dina(n230),.dinb(w_n159_0[0]),.dout(n231),.clk(gclk));
	jand g183(.dina(w_G370gat_2),.dinb(w_G14gat_0[1]),.dout(n232),.clk(gclk));
	jor g184(.dina(n232),.dinb(w_n231_0[1]),.dout(n233),.clk(gclk));
	jnot g185(.din(w_n151_0[0]),.dout(n235),.clk(gclk));
	jor g186(.dina(w_dff_B_ct5lXz6H6_0),.dinb(w_n147_0[0]),.dout(n237),.clk(gclk));
	jand g187(.dina(w_G329gat_4[0]),.dinb(w_G73gat_0[0]),.dout(n238),.clk(gclk));
	jor g188(.dina(n238),.dinb(w_n164_0[0]),.dout(n239),.clk(gclk));
	jor g189(.dina(n239),.dinb(w_G79gat_0[0]),.dout(n240),.clk(gclk));
	jand g190(.dina(n240),.dinb(w_dff_B_AxRQ3LvL6_1),.dout(n241),.clk(gclk));
	jand g191(.dina(n241),.dinb(w_n142_0[0]),.dout(n242),.clk(gclk));
	jnot g192(.din(w_n193_0[0]),.dout(n244),.clk(gclk));
	jor g193(.dina(w_dff_B_biS7DsnS2_0),.dinb(w_n188_0[0]),.dout(n246),.clk(gclk));
	jand g194(.dina(w_G329gat_3[2]),.dinb(w_G21gat_0[1]),.dout(n247),.clk(gclk));
	jor g195(.dina(n247),.dinb(w_n177_0[0]),.dout(n248),.clk(gclk));
	jand g196(.dina(w_n182_1[1]),.dinb(w_n130_0[0]),.dout(n249),.clk(gclk));
	jor g197(.dina(n249),.dinb(w_G27gat_0[0]),.dout(n250),.clk(gclk));
	jor g198(.dina(n250),.dinb(n248),.dout(n251),.clk(gclk));
	jand g199(.dina(n251),.dinb(w_dff_B_y8DmVsDm4_1),.dout(n252),.clk(gclk));
	jand g200(.dina(w_G329gat_3[1]),.dinb(w_G86gat_0[1]),.dout(n253),.clk(gclk));
	jor g201(.dina(n253),.dinb(w_n174_0[0]),.dout(n254),.clk(gclk));
	jand g202(.dina(w_n182_1[0]),.dinb(w_n126_0[0]),.dout(n255),.clk(gclk));
	jor g203(.dina(n255),.dinb(w_G92gat_0[1]),.dout(n256),.clk(gclk));
	jor g204(.dina(n256),.dinb(w_n254_0[1]),.dout(n257),.clk(gclk));
	jor g205(.dina(w_n231_0[0]),.dinb(w_G14gat_0[0]),.dout(n258),.clk(gclk));
	jand g206(.dina(n258),.dinb(n257),.dout(n259),.clk(gclk));
	jand g207(.dina(w_G329gat_3[0]),.dinb(w_G34gat_0[0]),.dout(n260),.clk(gclk));
	jnot g208(.din(w_n219_0[0]),.dout(n262),.clk(gclk));
	jor g209(.dina(w_dff_B_wR8dz6dx4_0),.dinb(w_n260_0[1]),.dout(n264),.clk(gclk));
	jand g210(.dina(w_G329gat_2[2]),.dinb(w_G112gat_0[0]),.dout(n265),.clk(gclk));
	jor g211(.dina(n265),.dinb(w_n156_0[0]),.dout(n266),.clk(gclk));
	jor g212(.dina(n266),.dinb(w_G115gat_0[0]),.dout(n267),.clk(gclk));
	jand g213(.dina(n267),.dinb(w_dff_B_uTuShrve9_1),.dout(n268),.clk(gclk));
	jand g214(.dina(n268),.dinb(n259),.dout(n269),.clk(gclk));
	jand g215(.dina(n269),.dinb(w_dff_B_K1thgq319_1),.dout(n270),.clk(gclk));
	jand g216(.dina(n270),.dinb(w_dff_B_2wFSzp307_1),.dout(n271),.clk(gclk));
	jor g217(.dina(w_n271_3[1]),.dinb(w_n150_0[0]),.dout(n272),.clk(gclk));
	jand g218(.dina(w_G329gat_2[1]),.dinb(w_G60gat_0[0]),.dout(n273),.clk(gclk));
	jor g219(.dina(n273),.dinb(w_n145_0[0]),.dout(n274),.clk(gclk));
	jnot g220(.din(w_n274_0[1]),.dout(n275),.clk(gclk));
	jand g221(.dina(w_dff_B_uBsrld240_0),.dinb(n272),.dout(n276),.clk(gclk));
	jor g222(.dina(w_n271_3[0]),.dinb(w_n191_0[0]),.dout(n277),.clk(gclk));
	jand g223(.dina(w_G329gat_2[0]),.dinb(w_G47gat_0[0]),.dout(n278),.clk(gclk));
	jand g224(.dina(w_G223gat_1[0]),.dinb(w_G37gat_0[0]),.dout(n279),.clk(gclk));
	jor g225(.dina(n279),.dinb(w_n77_0[0]),.dout(n280),.clk(gclk));
	jor g226(.dina(w_dff_B_Nl3mb62H5_0),.dinb(n278),.dout(n281),.clk(gclk));
	jnot g227(.din(w_n281_0[1]),.dout(n282),.clk(gclk));
	jand g228(.dina(w_dff_B_6ReuljeS7_0),.dinb(n277),.dout(n283),.clk(gclk));
	jor g229(.dina(w_n283_0[1]),.dinb(n276),.dout(n284),.clk(gclk));
	jor g230(.dina(w_n271_2[2]),.dinb(w_n198_0[0]),.dout(n285),.clk(gclk));
	jand g231(.dina(n285),.dinb(w_n197_0[0]),.dout(n286),.clk(gclk));
	jor g232(.dina(w_n271_2[1]),.dinb(w_n217_0[0]),.dout(n287),.clk(gclk));
	jor g233(.dina(w_n114_0[0]),.dinb(w_n260_0[0]),.dout(n290),.clk(gclk));
	jnot g234(.din(w_n290_0[1]),.dout(n291),.clk(gclk));
	jand g235(.dina(w_dff_B_5cwfiVA75_0),.dinb(n287),.dout(n292),.clk(gclk));
	jor g236(.dina(n292),.dinb(w_n286_0[1]),.dout(n293),.clk(gclk));
	jor g237(.dina(w_n293_0[1]),.dinb(n284),.dout(G430gat_fa_),.clk(gclk));
	jor g238(.dina(w_n271_2[0]),.dinb(w_n205_0[0]),.dout(n295),.clk(gclk));
	jand g239(.dina(n295),.dinb(w_n204_0[0]),.dout(n296),.clk(gclk));
	jor g240(.dina(w_n271_1[2]),.dinb(w_n222_0[0]),.dout(n297),.clk(gclk));
	jand g241(.dina(n297),.dinb(w_n224_0[0]),.dout(n298),.clk(gclk));
	jor g242(.dina(n298),.dinb(w_n296_0[1]),.dout(n299),.clk(gclk));
	jnot g243(.din(w_n141_0[0]),.dout(n300),.clk(gclk));
	jnot g244(.din(w_G105gat_0[0]),.dout(n301),.clk(gclk));
	jor g245(.dina(w_n271_1[1]),.dinb(w_dff_B_B7uisLfx7_1),.dout(n302),.clk(gclk));
	jand g246(.dina(n302),.dinb(w_dff_B_9HZyP6Zc0_1),.dout(n303),.clk(gclk));
	jor g247(.dina(w_n271_1[0]),.dinb(w_n154_0[0]),.dout(n304),.clk(gclk));
	jand g248(.dina(n304),.dinb(w_n184_0[0]),.dout(n305),.clk(gclk));
	jor g249(.dina(w_n305_0[1]),.dinb(w_n303_0[1]),.dout(n306),.clk(gclk));
	jor g250(.dina(n306),.dinb(n299),.dout(n307),.clk(gclk));
	jor g251(.dina(n307),.dinb(w_G430gat_0),.dout(n308),.clk(gclk));
	jand g252(.dina(n308),.dinb(w_dff_B_qeEHfVCL7_1),.dout(G421gat),.clk(gclk));
	jand g253(.dina(w_G370gat_1[2]),.dinb(w_G66gat_0[0]),.dout(n310),.clk(gclk));
	jor g254(.dina(w_n274_0[0]),.dinb(n310),.dout(n311),.clk(gclk));
	jand g255(.dina(w_G370gat_1[1]),.dinb(w_G53gat_0[0]),.dout(n312),.clk(gclk));
	jor g256(.dina(w_n281_0[0]),.dinb(n312),.dout(n313),.clk(gclk));
	jand g257(.dina(w_n313_0[1]),.dinb(n311),.dout(n314),.clk(gclk));
	jand g258(.dina(w_n296_0[0]),.dinb(w_n314_0[1]),.dout(n315),.clk(gclk));
	jand g259(.dina(w_G370gat_1[0]),.dinb(w_G40gat_0[0]),.dout(n316),.clk(gclk));
	jor g260(.dina(w_n290_0[0]),.dinb(n316),.dout(n317),.clk(gclk));
	jand g261(.dina(w_n305_0[0]),.dinb(w_n317_0[2]),.dout(n318),.clk(gclk));
	jand g262(.dina(n318),.dinb(w_n314_0[0]),.dout(n319),.clk(gclk));
	jor g263(.dina(w_n319_0[1]),.dinb(w_n293_0[0]),.dout(n320),.clk(gclk));
	jor g264(.dina(n320),.dinb(w_dff_B_ssGiefmH9_1),.dout(G431gat),.clk(gclk));
	jand g265(.dina(w_G370gat_0[2]),.dinb(w_G92gat_0[0]),.dout(n322),.clk(gclk));
	jor g266(.dina(n322),.dinb(w_n254_0[0]),.dout(n323),.clk(gclk));
	jand g267(.dina(n323),.dinb(w_n313_0[0]),.dout(n324),.clk(gclk));
	jand g268(.dina(w_n303_0[0]),.dinb(w_n317_0[1]),.dout(n325),.clk(gclk));
	jand g269(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jand g270(.dina(w_n317_0[0]),.dinb(w_n283_0[0]),.dout(n327),.clk(gclk));
	jor g271(.dina(n327),.dinb(w_n286_0[0]),.dout(n328),.clk(gclk));
	jor g272(.dina(n328),.dinb(w_n319_0[0]),.dout(n329),.clk(gclk));
	jor g273(.dina(n329),.dinb(w_dff_B_FhGW1nOI6_1),.dout(G432gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_uyyDderI0_0),.doutb(w_dff_A_hOBi2wgc9_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_dff_A_FJepJW0D0_0),.doutb(w_G4gat_0[1]),.doutc(w_dff_A_tllPJFyQ9_2),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_J7Ni8DGh5_0),.doutb(w_dff_A_Y58ckHoR2_1),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G11gat_0(.douta(w_dff_A_HkqsB3iX6_0),.doutb(w_dff_A_FoogvTwZ9_1),.doutc(w_G11gat_0[2]),.din(G11gat));
	jspl3 jspl3_w_G14gat_0(.douta(w_dff_A_ZHfG6End6_0),.doutb(w_dff_A_SRPEcVSu0_1),.doutc(w_G14gat_0[2]),.din(G14gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_dff_A_bC3ynXnv7_0),.doutb(w_G17gat_0[1]),.doutc(w_dff_A_9GN6vBZw5_2),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_G21gat_0[0]),.doutb(w_dff_A_PtjufDcc3_1),.doutc(w_dff_A_WshjxAfQ5_2),.din(G21gat));
	jspl jspl_w_G21gat_1(.douta(w_dff_A_oiRTHhbG8_0),.doutb(w_G21gat_1[1]),.din(w_G21gat_0[0]));
	jspl jspl_w_G24gat_0(.douta(w_dff_A_jsqxPSei4_0),.doutb(w_G24gat_0[1]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_dff_A_fuz1QEUW2_0),.doutb(w_G27gat_0[1]),.din(G27gat));
	jspl jspl_w_G30gat_0(.douta(w_G30gat_0[0]),.doutb(w_dff_A_r7zmGIrz2_1),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_dff_A_45KJcNxX6_0),.doutb(w_G34gat_0[1]),.doutc(w_dff_A_m4Ae2IwH6_2),.din(G34gat));
	jspl3 jspl3_w_G37gat_0(.douta(w_dff_A_ZmRpUAqN5_0),.doutb(w_dff_A_Il4LI20s8_1),.doutc(w_G37gat_0[2]),.din(G37gat));
	jspl jspl_w_G40gat_0(.douta(w_dff_A_cF2UM3na6_0),.doutb(w_G40gat_0[1]),.din(G40gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_G43gat_0[0]),.doutb(w_dff_A_p2oaRg9A0_1),.doutc(w_dff_A_XkeiPx5T6_2),.din(G43gat));
	jspl jspl_w_G43gat_1(.douta(w_G43gat_1[0]),.doutb(w_dff_A_9MNA8pJX2_1),.din(w_G43gat_0[0]));
	jspl jspl_w_G47gat_0(.douta(w_dff_A_8CCDWlrJ8_0),.doutb(w_G47gat_0[1]),.din(G47gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_dff_A_5wj2Tdsz1_0),.doutb(w_dff_A_XzzsQ4iL7_1),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_dff_A_i8Zztezs4_0),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_dff_A_Qc6vKUw11_0),.doutb(w_G56gat_0[1]),.doutc(w_dff_A_8P84km3w1_2),.din(G56gat));
	jspl3 jspl3_w_G60gat_0(.douta(w_dff_A_o998TikY5_0),.doutb(w_dff_A_8tObnMCA4_1),.doutc(w_G60gat_0[2]),.din(G60gat));
	jspl3 jspl3_w_G63gat_0(.douta(w_dff_A_N0thLyMm9_0),.doutb(w_dff_A_XJYSseO16_1),.doutc(w_G63gat_0[2]),.din(G63gat));
	jspl jspl_w_G66gat_0(.douta(w_dff_A_2DolGJBw8_0),.doutb(w_G66gat_0[1]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_dff_A_x6jLjakQ4_0),.doutb(w_G69gat_0[1]),.doutc(w_dff_A_H1t0GsEX5_2),.din(G69gat));
	jspl3 jspl3_w_G73gat_0(.douta(w_dff_A_y9vALicB7_0),.doutb(w_dff_A_jPiuEvLn5_1),.doutc(w_G73gat_0[2]),.din(G73gat));
	jspl jspl_w_G76gat_0(.douta(w_dff_A_IwzqA2iF0_0),.doutb(w_G76gat_0[1]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_dff_A_qE4HPvK16_0),.doutb(w_G79gat_0[1]),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_G82gat_0[0]),.doutb(w_dff_A_Oq19nnOW7_1),.doutc(w_dff_A_0LFFT8AU3_2),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_dff_A_ypIElH5r9_1),.doutc(w_dff_A_UJJOc4yD7_2),.din(G86gat));
	jspl jspl_w_G86gat_1(.douta(w_dff_A_yjVedfVQ4_0),.doutb(w_G86gat_1[1]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G89gat_0(.douta(w_dff_A_vkNPP3Cd8_0),.doutb(w_dff_A_h9q6CtEl3_1),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_6AlgyhNC8_0),.doutb(w_dff_A_pVnNe7Ql2_1),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_dff_A_6YUz5bTd3_0),.doutb(w_G95gat_0[1]),.doutc(w_dff_A_ArKlI0YR1_2),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_rNQHft9w8_0),.doutb(w_dff_A_pePc5qPA2_1),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl3 jspl3_w_G102gat_0(.douta(w_dff_A_AQOtljhc9_0),.doutb(w_dff_A_MKhlq43s3_1),.doutc(w_G102gat_0[2]),.din(G102gat));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_dff_A_vzdET3bI2_1),.din(G105gat));
	jspl3 jspl3_w_G108gat_0(.douta(w_dff_A_VPLfegx98_0),.doutb(w_G108gat_0[1]),.doutc(w_dff_A_qB1wV2iS1_2),.din(G108gat));
	jspl3 jspl3_w_G112gat_0(.douta(w_dff_A_2vpsb4yq7_0),.doutb(w_dff_A_JXS19OY08_1),.doutc(w_G112gat_0[2]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_dff_A_pTPvviVi8_0),.doutb(w_G115gat_0[1]),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(w_dff_A_UpkpSmaE9_2),.din(w_G223gat_0[2]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl3 jspl3_w_G329gat_4(.douta(w_G329gat_4[0]),.doutb(w_G329gat_4[1]),.doutc(w_G329gat_4[2]),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G329gat_5(.douta(w_G329gat_5[0]),.doutb(w_G329gat_5[1]),.doutc(w_G329gat_5[2]),.din(w_G329gat_1[1]));
	jspl jspl_w_G329gat_6(.douta(w_G329gat_6),.doutb(w_dff_A_Bu8Xx7qr6_1),.din(w_G329gat_1[2]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_G370gat_1[2]),.din(w_G370gat_0[0]));
	jspl jspl_w_G370gat_2(.douta(w_G370gat_2),.doutb(w_dff_A_LssHnvSR5_1),.din(w_G370gat_0[1]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(w_dff_A_vdAnjuUY2_1),.din(G430gat_fa_));
	jspl jspl_w_n43_0(.douta(w_dff_A_60Isjg0p8_0),.doutb(w_n43_0[1]),.din(n43));
	jspl jspl_w_n44_0(.douta(w_n44_0[0]),.doutb(w_dff_A_hLMVnkT17_1),.din(n44));
	jspl jspl_w_n47_0(.douta(w_dff_A_4sFDhFEl2_0),.doutb(w_n47_0[1]),.din(n47));
	jspl jspl_w_n52_0(.douta(w_dff_A_AD4OIk8E3_0),.doutb(w_n52_0[1]),.din(n52));
	jspl jspl_w_n53_0(.douta(w_dff_A_ivBejZGA4_0),.doutb(w_n53_0[1]),.din(n53));
	jspl jspl_w_n56_0(.douta(w_dff_A_bpBTlwkC8_0),.doutb(w_n56_0[1]),.din(n56));
	jspl jspl_w_n58_0(.douta(w_dff_A_gGvRmQIr2_0),.doutb(w_n58_0[1]),.din(n58));
	jspl jspl_w_n61_0(.douta(w_dff_A_bTB9zVMv4_0),.doutb(w_n61_0[1]),.din(n61));
	jspl jspl_w_n63_0(.douta(w_dff_A_yDrnNUkO3_0),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n69_0(.douta(w_dff_A_idV8RLow4_0),.doutb(w_n69_0[1]),.din(w_dff_B_YvfeFDYf2_2));
	jspl jspl_w_n71_0(.douta(w_dff_A_kqsSluya0_0),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n72_0(.douta(w_dff_A_dQi7a2mO7_0),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n73_0(.douta(w_dff_A_W85tryrl8_0),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n77_0(.douta(w_dff_A_8dZ7FzZd5_0),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_dff_A_MPNdGI4x0_0),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n79_0(.douta(w_dff_A_oDIYdEqg1_0),.doutb(w_n79_0[1]),.din(n79));
	jspl jspl_w_n82_0(.douta(w_dff_A_ZhhdXqXN7_0),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_dff_A_dhXW7ami4_0),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n87_0(.douta(w_dff_A_98SxYP9q9_0),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_dff_A_LSQjTqpw4_0),.doutb(w_n89_0[1]),.din(n89));
	jspl3 jspl3_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl3 jspl3_w_n94_1(.douta(w_n94_1[0]),.doutb(w_n94_1[1]),.doutc(w_n94_1[2]),.din(w_n94_0[0]));
	jspl3 jspl3_w_n94_2(.douta(w_n94_2[0]),.doutb(w_n94_2[1]),.doutc(w_n94_2[2]),.din(w_n94_0[1]));
	jspl3 jspl3_w_n94_3(.douta(w_n94_3[0]),.doutb(w_n94_3[1]),.doutc(w_n94_3[2]),.din(w_n94_0[2]));
	jspl jspl_w_n94_4(.douta(w_n94_4[0]),.doutb(w_n94_4[1]),.din(w_n94_1[0]));
	jspl jspl_w_n96_0(.douta(w_dff_A_llwuIglX9_0),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_dff_A_9ffzE9Xe7_0),.doutb(w_n98_0[1]),.din(w_dff_B_QCuW35tF1_2));
	jspl jspl_w_n100_0(.douta(w_dff_A_adLR2nLQ3_0),.doutb(w_n100_0[1]),.din(n100));
	jspl jspl_w_n107_0(.douta(w_dff_A_uuYeohou6_0),.doutb(w_n107_0[1]),.din(w_dff_B_KjPWA0K59_2));
	jspl jspl_w_n109_0(.douta(w_dff_A_9PWh6pjL1_0),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n114_0(.douta(w_dff_A_vzpAS6T33_0),.doutb(w_n114_0[1]),.doutc(w_n114_0[2]),.din(n114));
	jspl jspl_w_n115_0(.douta(w_dff_A_jRWMkcb75_0),.doutb(w_n115_0[1]),.din(n115));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n123_0(.douta(w_n123_0[0]),.doutb(w_dff_A_pH0zxLsr9_1),.din(n123));
	jspl3 jspl3_w_n126_0(.douta(w_dff_A_3b6KP1Xr0_0),.doutb(w_dff_A_lHnmXJzK4_1),.doutc(w_n126_0[2]),.din(w_dff_B_YeLHtNcC6_3));
	jspl jspl_w_n128_0(.douta(w_dff_A_ZIsEgJ3T1_0),.doutb(w_n128_0[1]),.din(n128));
	jspl3 jspl3_w_n130_0(.douta(w_dff_A_JeYl2SgM1_0),.doutb(w_dff_A_tO3P15gs0_1),.doutc(w_n130_0[2]),.din(w_dff_B_EzKS0AVu8_3));
	jspl jspl_w_n132_0(.douta(w_dff_A_L7UkzfMe6_0),.doutb(w_n132_0[1]),.din(n132));
	jspl jspl_w_n139_0(.douta(w_n139_0[0]),.doutb(w_dff_A_fT9wljA27_1),.din(n139));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_dff_A_EPfnWR8I7_0),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n145_0(.douta(w_dff_A_bgm1NLjI3_0),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_B6fkMwmI7_1),.din(n146));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl jspl_w_n150_0(.douta(w_dff_A_vBJ43En75_0),.doutb(w_n150_0[1]),.din(w_dff_B_GAX9VgP40_2));
	jspl jspl_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_JNGfH7qg4_1),.din(n151));
	jspl jspl_w_n154_0(.douta(w_dff_A_Rx2Dkhn52_0),.doutb(w_n154_0[1]),.din(w_dff_B_ptDOWvoi1_2));
	jspl jspl_w_n156_0(.douta(w_dff_A_femGqmDM7_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n159_0(.douta(w_dff_A_1LY0ds4S1_0),.doutb(w_n159_0[1]),.din(n159));
	jspl jspl_w_n164_0(.douta(w_dff_A_BB2erPz25_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n170_0(.douta(w_dff_A_f8IuNFel1_0),.doutb(w_n170_0[1]),.din(w_dff_B_AkYWyoNi7_2));
	jspl jspl_w_n174_0(.douta(w_dff_A_KrOIrhnz6_0),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n177_0(.douta(w_dff_A_CLTiIAIk1_0),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n182_2(.douta(w_n182_2[0]),.doutb(w_n182_2[1]),.doutc(w_n182_2[2]),.din(w_n182_0[1]));
	jspl jspl_w_n182_3(.douta(w_n182_3[0]),.doutb(w_n182_3[1]),.din(w_n182_0[2]));
	jspl jspl_w_n184_0(.douta(w_dff_A_SI3AbHif1_0),.doutb(w_n184_0[1]),.din(n184));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n191_0(.douta(w_dff_A_IL5ZPbh26_0),.doutb(w_n191_0[1]),.din(n191));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_dff_A_7K0OEzMt0_1),.din(n193));
	jspl jspl_w_n197_0(.douta(w_dff_A_D4Qlff1r3_0),.doutb(w_n197_0[1]),.din(n197));
	jspl jspl_w_n198_0(.douta(w_dff_A_5vpnn1Hd2_0),.doutb(w_n198_0[1]),.din(w_dff_B_DTbtNB9T8_2));
	jspl jspl_w_n204_0(.douta(w_dff_A_fS7LI9u52_0),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n205_0(.douta(w_dff_A_EaVkdNfv5_0),.doutb(w_n205_0[1]),.din(w_dff_B_FbCWni4c0_2));
	jspl jspl_w_n217_0(.douta(w_dff_A_oe4tlPCg9_0),.doutb(w_n217_0[1]),.din(w_dff_B_FVREnZD71_2));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_dff_A_d54mL2Om9_1),.din(n219));
	jspl jspl_w_n222_0(.douta(w_dff_A_yc8ikB592_0),.doutb(w_n222_0[1]),.din(w_dff_B_Xc4m6MZ12_2));
	jspl jspl_w_n224_0(.douta(w_dff_A_uWXJDqR56_0),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_dff_A_7RxalIYA6_1),.din(n231));
	jspl jspl_w_n254_0(.douta(w_dff_A_MfOkD83t9_0),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_n271_1[0]),.doutb(w_n271_1[1]),.doutc(w_n271_1[2]),.din(w_n271_0[0]));
	jspl3 jspl3_w_n271_2(.douta(w_n271_2[0]),.doutb(w_n271_2[1]),.doutc(w_n271_2[2]),.din(w_n271_0[1]));
	jspl jspl_w_n271_3(.douta(w_n271_3[0]),.doutb(w_n271_3[1]),.din(w_n271_0[2]));
	jspl jspl_w_n274_0(.douta(w_dff_A_mRCu6KOv1_0),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n281_0(.douta(w_dff_A_v9VcLd3g7_0),.doutb(w_n281_0[1]),.din(n281));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.din(n283));
	jspl jspl_w_n286_0(.douta(w_dff_A_bhanmIps5_0),.doutb(w_n286_0[1]),.din(n286));
	jspl jspl_w_n290_0(.douta(w_dff_A_t8PbktgK8_0),.doutb(w_n290_0[1]),.din(n290));
	jspl jspl_w_n293_0(.douta(w_dff_A_63oNAdLK8_0),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n296_0(.douta(w_dff_A_LMnmGZJm4_0),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(n305));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.din(n314));
	jspl3 jspl3_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.doutc(w_n317_0[2]),.din(n317));
	jspl jspl_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.din(n319));
	jdff dff_B_E84WjtqU9_1(.din(n233),.dout(w_dff_B_E84WjtqU9_1),.clk(gclk));
	jdff dff_B_b9HyKMji5_1(.din(w_dff_B_E84WjtqU9_1),.dout(w_dff_B_b9HyKMji5_1),.clk(gclk));
	jdff dff_B_qeEHfVCL7_1(.din(w_dff_B_b9HyKMji5_1),.dout(w_dff_B_qeEHfVCL7_1),.clk(gclk));
	jdff dff_B_brIiDbPX4_0(.din(n275),.dout(w_dff_B_brIiDbPX4_0),.clk(gclk));
	jdff dff_B_PyLHbrk94_0(.din(w_dff_B_brIiDbPX4_0),.dout(w_dff_B_PyLHbrk94_0),.clk(gclk));
	jdff dff_B_PqG1ajbQ5_0(.din(w_dff_B_PyLHbrk94_0),.dout(w_dff_B_PqG1ajbQ5_0),.clk(gclk));
	jdff dff_B_jNwrjMXK6_0(.din(w_dff_B_PqG1ajbQ5_0),.dout(w_dff_B_jNwrjMXK6_0),.clk(gclk));
	jdff dff_B_uBsrld240_0(.din(w_dff_B_jNwrjMXK6_0),.dout(w_dff_B_uBsrld240_0),.clk(gclk));
	jdff dff_B_ssGiefmH9_1(.din(n315),.dout(w_dff_B_ssGiefmH9_1),.clk(gclk));
	jdff dff_A_63oNAdLK8_0(.dout(w_n293_0[0]),.din(w_dff_A_63oNAdLK8_0),.clk(gclk));
	jdff dff_B_OQVJCjD14_0(.din(n291),.dout(w_dff_B_OQVJCjD14_0),.clk(gclk));
	jdff dff_B_yJb4L9dF8_0(.din(w_dff_B_OQVJCjD14_0),.dout(w_dff_B_yJb4L9dF8_0),.clk(gclk));
	jdff dff_B_GRe8qVV25_0(.din(w_dff_B_yJb4L9dF8_0),.dout(w_dff_B_GRe8qVV25_0),.clk(gclk));
	jdff dff_B_immWqEAs3_0(.din(w_dff_B_GRe8qVV25_0),.dout(w_dff_B_immWqEAs3_0),.clk(gclk));
	jdff dff_B_5cwfiVA75_0(.din(w_dff_B_immWqEAs3_0),.dout(w_dff_B_5cwfiVA75_0),.clk(gclk));
	jdff dff_A_LMnmGZJm4_0(.dout(w_n296_0[0]),.din(w_dff_A_LMnmGZJm4_0),.clk(gclk));
	jdff dff_B_FhGW1nOI6_1(.din(n326),.dout(w_dff_B_FhGW1nOI6_1),.clk(gclk));
	jdff dff_B_lX9AQn0i9_0(.din(n282),.dout(w_dff_B_lX9AQn0i9_0),.clk(gclk));
	jdff dff_B_jefqsd6x1_0(.din(w_dff_B_lX9AQn0i9_0),.dout(w_dff_B_jefqsd6x1_0),.clk(gclk));
	jdff dff_B_8qO7u2pw1_0(.din(w_dff_B_jefqsd6x1_0),.dout(w_dff_B_8qO7u2pw1_0),.clk(gclk));
	jdff dff_B_qrSNogx69_0(.din(w_dff_B_8qO7u2pw1_0),.dout(w_dff_B_qrSNogx69_0),.clk(gclk));
	jdff dff_B_6ReuljeS7_0(.din(w_dff_B_qrSNogx69_0),.dout(w_dff_B_6ReuljeS7_0),.clk(gclk));
	jdff dff_A_bhanmIps5_0(.dout(w_n286_0[0]),.din(w_dff_A_bhanmIps5_0),.clk(gclk));
	jdff dff_A_we74WJ5x3_0(.dout(w_n274_0[0]),.din(w_dff_A_we74WJ5x3_0),.clk(gclk));
	jdff dff_A_HiEgvwr16_0(.dout(w_dff_A_we74WJ5x3_0),.din(w_dff_A_HiEgvwr16_0),.clk(gclk));
	jdff dff_A_LhdOrUZ06_0(.dout(w_dff_A_HiEgvwr16_0),.din(w_dff_A_LhdOrUZ06_0),.clk(gclk));
	jdff dff_A_UWlYa7UW3_0(.dout(w_dff_A_LhdOrUZ06_0),.din(w_dff_A_UWlYa7UW3_0),.clk(gclk));
	jdff dff_A_Wxwv153g2_0(.dout(w_dff_A_UWlYa7UW3_0),.din(w_dff_A_Wxwv153g2_0),.clk(gclk));
	jdff dff_A_mRCu6KOv1_0(.dout(w_dff_A_Wxwv153g2_0),.din(w_dff_A_mRCu6KOv1_0),.clk(gclk));
	jdff dff_B_Pt70dW2M2_1(.din(n300),.dout(w_dff_B_Pt70dW2M2_1),.clk(gclk));
	jdff dff_B_RGMPKndI4_1(.din(w_dff_B_Pt70dW2M2_1),.dout(w_dff_B_RGMPKndI4_1),.clk(gclk));
	jdff dff_B_7cuj51sA5_1(.din(w_dff_B_RGMPKndI4_1),.dout(w_dff_B_7cuj51sA5_1),.clk(gclk));
	jdff dff_B_v7onULsi4_1(.din(w_dff_B_7cuj51sA5_1),.dout(w_dff_B_v7onULsi4_1),.clk(gclk));
	jdff dff_B_9HZyP6Zc0_1(.din(w_dff_B_v7onULsi4_1),.dout(w_dff_B_9HZyP6Zc0_1),.clk(gclk));
	jdff dff_B_osD97IsC4_1(.din(n301),.dout(w_dff_B_osD97IsC4_1),.clk(gclk));
	jdff dff_B_BXLEhURq1_1(.din(w_dff_B_osD97IsC4_1),.dout(w_dff_B_BXLEhURq1_1),.clk(gclk));
	jdff dff_B_1B5oGgdT8_1(.din(w_dff_B_BXLEhURq1_1),.dout(w_dff_B_1B5oGgdT8_1),.clk(gclk));
	jdff dff_B_6GpfLvS53_1(.din(w_dff_B_1B5oGgdT8_1),.dout(w_dff_B_6GpfLvS53_1),.clk(gclk));
	jdff dff_B_Do7VOgU68_1(.din(w_dff_B_6GpfLvS53_1),.dout(w_dff_B_Do7VOgU68_1),.clk(gclk));
	jdff dff_B_D2q8IV318_1(.din(w_dff_B_Do7VOgU68_1),.dout(w_dff_B_D2q8IV318_1),.clk(gclk));
	jdff dff_B_On0SCoFm1_1(.din(w_dff_B_D2q8IV318_1),.dout(w_dff_B_On0SCoFm1_1),.clk(gclk));
	jdff dff_B_A8tYvMnT1_1(.din(w_dff_B_On0SCoFm1_1),.dout(w_dff_B_A8tYvMnT1_1),.clk(gclk));
	jdff dff_B_GXgKwjET1_1(.din(w_dff_B_A8tYvMnT1_1),.dout(w_dff_B_GXgKwjET1_1),.clk(gclk));
	jdff dff_B_f1PbK5JV1_1(.din(w_dff_B_GXgKwjET1_1),.dout(w_dff_B_f1PbK5JV1_1),.clk(gclk));
	jdff dff_B_JchGTsiz1_1(.din(w_dff_B_f1PbK5JV1_1),.dout(w_dff_B_JchGTsiz1_1),.clk(gclk));
	jdff dff_B_QYQQMzsr4_1(.din(w_dff_B_JchGTsiz1_1),.dout(w_dff_B_QYQQMzsr4_1),.clk(gclk));
	jdff dff_B_5h4ow6XR1_1(.din(w_dff_B_QYQQMzsr4_1),.dout(w_dff_B_5h4ow6XR1_1),.clk(gclk));
	jdff dff_B_KJ6kQ9ow5_1(.din(w_dff_B_5h4ow6XR1_1),.dout(w_dff_B_KJ6kQ9ow5_1),.clk(gclk));
	jdff dff_B_bTfpLFxD2_1(.din(w_dff_B_KJ6kQ9ow5_1),.dout(w_dff_B_bTfpLFxD2_1),.clk(gclk));
	jdff dff_B_TaFCL5fq0_1(.din(w_dff_B_bTfpLFxD2_1),.dout(w_dff_B_TaFCL5fq0_1),.clk(gclk));
	jdff dff_B_bYlbaeYM8_1(.din(w_dff_B_TaFCL5fq0_1),.dout(w_dff_B_bYlbaeYM8_1),.clk(gclk));
	jdff dff_B_gpnxk3wg2_1(.din(w_dff_B_bYlbaeYM8_1),.dout(w_dff_B_gpnxk3wg2_1),.clk(gclk));
	jdff dff_B_B7uisLfx7_1(.din(w_dff_B_gpnxk3wg2_1),.dout(w_dff_B_B7uisLfx7_1),.clk(gclk));
	jdff dff_B_2wFSzp307_1(.din(n242),.dout(w_dff_B_2wFSzp307_1),.clk(gclk));
	jdff dff_B_K1thgq319_1(.din(n252),.dout(w_dff_B_K1thgq319_1),.clk(gclk));
	jdff dff_B_uTuShrve9_1(.din(n264),.dout(w_dff_B_uTuShrve9_1),.clk(gclk));
	jdff dff_B_0v3JXI7t8_0(.din(n262),.dout(w_dff_B_0v3JXI7t8_0),.clk(gclk));
	jdff dff_B_zcZgJHWH2_0(.din(w_dff_B_0v3JXI7t8_0),.dout(w_dff_B_zcZgJHWH2_0),.clk(gclk));
	jdff dff_B_wR8dz6dx4_0(.din(w_dff_B_zcZgJHWH2_0),.dout(w_dff_B_wR8dz6dx4_0),.clk(gclk));
	jdff dff_A_xKJdmaWY3_1(.dout(w_n231_0[1]),.din(w_dff_A_xKJdmaWY3_1),.clk(gclk));
	jdff dff_A_JxDwUKru5_1(.dout(w_dff_A_xKJdmaWY3_1),.din(w_dff_A_JxDwUKru5_1),.clk(gclk));
	jdff dff_A_rH4XgQez6_1(.dout(w_dff_A_JxDwUKru5_1),.din(w_dff_A_rH4XgQez6_1),.clk(gclk));
	jdff dff_A_FX0Locty1_1(.dout(w_dff_A_rH4XgQez6_1),.din(w_dff_A_FX0Locty1_1),.clk(gclk));
	jdff dff_A_G9mKx2417_1(.dout(w_dff_A_FX0Locty1_1),.din(w_dff_A_G9mKx2417_1),.clk(gclk));
	jdff dff_A_7RxalIYA6_1(.dout(w_dff_A_G9mKx2417_1),.din(w_dff_A_7RxalIYA6_1),.clk(gclk));
	jdff dff_B_y8DmVsDm4_1(.din(n246),.dout(w_dff_B_y8DmVsDm4_1),.clk(gclk));
	jdff dff_B_3s5pqZGe8_0(.din(n244),.dout(w_dff_B_3s5pqZGe8_0),.clk(gclk));
	jdff dff_B_qJUcp0DF8_0(.din(w_dff_B_3s5pqZGe8_0),.dout(w_dff_B_qJUcp0DF8_0),.clk(gclk));
	jdff dff_B_De8g2oe11_0(.din(w_dff_B_qJUcp0DF8_0),.dout(w_dff_B_De8g2oe11_0),.clk(gclk));
	jdff dff_B_knX7jJXR9_0(.din(w_dff_B_De8g2oe11_0),.dout(w_dff_B_knX7jJXR9_0),.clk(gclk));
	jdff dff_B_biS7DsnS2_0(.din(w_dff_B_knX7jJXR9_0),.dout(w_dff_B_biS7DsnS2_0),.clk(gclk));
	jdff dff_B_AxRQ3LvL6_1(.din(n237),.dout(w_dff_B_AxRQ3LvL6_1),.clk(gclk));
	jdff dff_B_ogrRlWLn5_0(.din(n235),.dout(w_dff_B_ogrRlWLn5_0),.clk(gclk));
	jdff dff_B_6wxqCpKy4_0(.din(w_dff_B_ogrRlWLn5_0),.dout(w_dff_B_6wxqCpKy4_0),.clk(gclk));
	jdff dff_B_BzcxujOr8_0(.din(w_dff_B_6wxqCpKy4_0),.dout(w_dff_B_BzcxujOr8_0),.clk(gclk));
	jdff dff_B_ct5lXz6H6_0(.din(w_dff_B_BzcxujOr8_0),.dout(w_dff_B_ct5lXz6H6_0),.clk(gclk));
	jdff dff_A_cFHfMqxb5_0(.dout(w_n290_0[0]),.din(w_dff_A_cFHfMqxb5_0),.clk(gclk));
	jdff dff_A_sOeOPPvk6_0(.dout(w_dff_A_cFHfMqxb5_0),.din(w_dff_A_sOeOPPvk6_0),.clk(gclk));
	jdff dff_A_ILdHlcoY5_0(.dout(w_dff_A_sOeOPPvk6_0),.din(w_dff_A_ILdHlcoY5_0),.clk(gclk));
	jdff dff_A_rPIuqBvc7_0(.dout(w_dff_A_ILdHlcoY5_0),.din(w_dff_A_rPIuqBvc7_0),.clk(gclk));
	jdff dff_A_HsczOm9L7_0(.dout(w_dff_A_rPIuqBvc7_0),.din(w_dff_A_HsczOm9L7_0),.clk(gclk));
	jdff dff_A_t8PbktgK8_0(.dout(w_dff_A_HsczOm9L7_0),.din(w_dff_A_t8PbktgK8_0),.clk(gclk));
	jdff dff_A_35Waeda05_0(.dout(w_n254_0[0]),.din(w_dff_A_35Waeda05_0),.clk(gclk));
	jdff dff_A_f8rAJGZn9_0(.dout(w_dff_A_35Waeda05_0),.din(w_dff_A_f8rAJGZn9_0),.clk(gclk));
	jdff dff_A_VopBQ54b6_0(.dout(w_dff_A_f8rAJGZn9_0),.din(w_dff_A_VopBQ54b6_0),.clk(gclk));
	jdff dff_A_CpLrv76n4_0(.dout(w_dff_A_VopBQ54b6_0),.din(w_dff_A_CpLrv76n4_0),.clk(gclk));
	jdff dff_A_6IO6HRAS4_0(.dout(w_dff_A_CpLrv76n4_0),.din(w_dff_A_6IO6HRAS4_0),.clk(gclk));
	jdff dff_A_MfOkD83t9_0(.dout(w_dff_A_6IO6HRAS4_0),.din(w_dff_A_MfOkD83t9_0),.clk(gclk));
	jdff dff_A_exauHlsj2_0(.dout(w_n281_0[0]),.din(w_dff_A_exauHlsj2_0),.clk(gclk));
	jdff dff_A_BGslSIQO3_0(.dout(w_dff_A_exauHlsj2_0),.din(w_dff_A_BGslSIQO3_0),.clk(gclk));
	jdff dff_A_34zFNiej2_0(.dout(w_dff_A_BGslSIQO3_0),.din(w_dff_A_34zFNiej2_0),.clk(gclk));
	jdff dff_A_EdUu0n264_0(.dout(w_dff_A_34zFNiej2_0),.din(w_dff_A_EdUu0n264_0),.clk(gclk));
	jdff dff_A_brlJoA973_0(.dout(w_dff_A_EdUu0n264_0),.din(w_dff_A_brlJoA973_0),.clk(gclk));
	jdff dff_A_v9VcLd3g7_0(.dout(w_dff_A_brlJoA973_0),.din(w_dff_A_v9VcLd3g7_0),.clk(gclk));
	jdff dff_B_QrmimWgB9_0(.din(n280),.dout(w_dff_B_QrmimWgB9_0),.clk(gclk));
	jdff dff_B_nAh1Dqaq0_0(.din(w_dff_B_QrmimWgB9_0),.dout(w_dff_B_nAh1Dqaq0_0),.clk(gclk));
	jdff dff_B_qFZ28XBB5_0(.din(w_dff_B_nAh1Dqaq0_0),.dout(w_dff_B_qFZ28XBB5_0),.clk(gclk));
	jdff dff_B_J09rXRIQ9_0(.din(w_dff_B_qFZ28XBB5_0),.dout(w_dff_B_J09rXRIQ9_0),.clk(gclk));
	jdff dff_B_hFem99714_0(.din(w_dff_B_J09rXRIQ9_0),.dout(w_dff_B_hFem99714_0),.clk(gclk));
	jdff dff_B_Nl3mb62H5_0(.din(w_dff_B_hFem99714_0),.dout(w_dff_B_Nl3mb62H5_0),.clk(gclk));
	jdff dff_B_2TnlZEFq4_1(.din(n187),.dout(w_dff_B_2TnlZEFq4_1),.clk(gclk));
	jdff dff_B_A6RWogJ76_1(.din(n202),.dout(w_dff_B_A6RWogJ76_1),.clk(gclk));
	jdff dff_B_Lmvqt5U65_1(.din(n221),.dout(w_dff_B_Lmvqt5U65_1),.clk(gclk));
	jdff dff_A_Gxyn36e49_0(.dout(w_n224_0[0]),.din(w_dff_A_Gxyn36e49_0),.clk(gclk));
	jdff dff_A_BPcPin6M4_0(.dout(w_dff_A_Gxyn36e49_0),.din(w_dff_A_BPcPin6M4_0),.clk(gclk));
	jdff dff_A_vl4FimtG9_0(.dout(w_dff_A_BPcPin6M4_0),.din(w_dff_A_vl4FimtG9_0),.clk(gclk));
	jdff dff_A_ReyVoHjd7_0(.dout(w_dff_A_vl4FimtG9_0),.din(w_dff_A_ReyVoHjd7_0),.clk(gclk));
	jdff dff_A_qyrcAqG02_0(.dout(w_dff_A_ReyVoHjd7_0),.din(w_dff_A_qyrcAqG02_0),.clk(gclk));
	jdff dff_A_uWXJDqR56_0(.dout(w_dff_A_qyrcAqG02_0),.din(w_dff_A_uWXJDqR56_0),.clk(gclk));
	jdff dff_A_YiRU4dyJ8_0(.dout(w_n222_0[0]),.din(w_dff_A_YiRU4dyJ8_0),.clk(gclk));
	jdff dff_A_URdEWoJq1_0(.dout(w_dff_A_YiRU4dyJ8_0),.din(w_dff_A_URdEWoJq1_0),.clk(gclk));
	jdff dff_A_GcCtW2Bk8_0(.dout(w_dff_A_URdEWoJq1_0),.din(w_dff_A_GcCtW2Bk8_0),.clk(gclk));
	jdff dff_A_ILCPC6pi0_0(.dout(w_dff_A_GcCtW2Bk8_0),.din(w_dff_A_ILCPC6pi0_0),.clk(gclk));
	jdff dff_A_yc8ikB592_0(.dout(w_dff_A_ILCPC6pi0_0),.din(w_dff_A_yc8ikB592_0),.clk(gclk));
	jdff dff_B_BXQdMy1D2_2(.din(n222),.dout(w_dff_B_BXQdMy1D2_2),.clk(gclk));
	jdff dff_B_YvDbImdz1_2(.din(w_dff_B_BXQdMy1D2_2),.dout(w_dff_B_YvDbImdz1_2),.clk(gclk));
	jdff dff_B_J54WOYsi1_2(.din(w_dff_B_YvDbImdz1_2),.dout(w_dff_B_J54WOYsi1_2),.clk(gclk));
	jdff dff_B_5wjd3s9X3_2(.din(w_dff_B_J54WOYsi1_2),.dout(w_dff_B_5wjd3s9X3_2),.clk(gclk));
	jdff dff_B_X0bT0CAM4_2(.din(w_dff_B_5wjd3s9X3_2),.dout(w_dff_B_X0bT0CAM4_2),.clk(gclk));
	jdff dff_B_Pf9E87fF5_2(.din(w_dff_B_X0bT0CAM4_2),.dout(w_dff_B_Pf9E87fF5_2),.clk(gclk));
	jdff dff_B_EeTdyLnm5_2(.din(w_dff_B_Pf9E87fF5_2),.dout(w_dff_B_EeTdyLnm5_2),.clk(gclk));
	jdff dff_B_GKHCdxW71_2(.din(w_dff_B_EeTdyLnm5_2),.dout(w_dff_B_GKHCdxW71_2),.clk(gclk));
	jdff dff_B_Ai9M8hI28_2(.din(w_dff_B_GKHCdxW71_2),.dout(w_dff_B_Ai9M8hI28_2),.clk(gclk));
	jdff dff_B_Ej7AXUqa7_2(.din(w_dff_B_Ai9M8hI28_2),.dout(w_dff_B_Ej7AXUqa7_2),.clk(gclk));
	jdff dff_B_GewKCm6z4_2(.din(w_dff_B_Ej7AXUqa7_2),.dout(w_dff_B_GewKCm6z4_2),.clk(gclk));
	jdff dff_B_iI5YOLjt6_2(.din(w_dff_B_GewKCm6z4_2),.dout(w_dff_B_iI5YOLjt6_2),.clk(gclk));
	jdff dff_B_bPCAM6l94_2(.din(w_dff_B_iI5YOLjt6_2),.dout(w_dff_B_bPCAM6l94_2),.clk(gclk));
	jdff dff_B_Xc4m6MZ12_2(.din(w_dff_B_bPCAM6l94_2),.dout(w_dff_B_Xc4m6MZ12_2),.clk(gclk));
	jdff dff_A_utroPy4g4_0(.dout(w_G115gat_0[0]),.din(w_dff_A_utroPy4g4_0),.clk(gclk));
	jdff dff_A_c5IvWWXm1_0(.dout(w_dff_A_utroPy4g4_0),.din(w_dff_A_c5IvWWXm1_0),.clk(gclk));
	jdff dff_A_JsiZLXWc6_0(.dout(w_dff_A_c5IvWWXm1_0),.din(w_dff_A_JsiZLXWc6_0),.clk(gclk));
	jdff dff_A_0l8e7Srp5_0(.dout(w_dff_A_JsiZLXWc6_0),.din(w_dff_A_0l8e7Srp5_0),.clk(gclk));
	jdff dff_A_BeTwbTta5_0(.dout(w_dff_A_0l8e7Srp5_0),.din(w_dff_A_BeTwbTta5_0),.clk(gclk));
	jdff dff_A_qXG8zpi81_0(.dout(w_dff_A_BeTwbTta5_0),.din(w_dff_A_qXG8zpi81_0),.clk(gclk));
	jdff dff_A_aquxKKMG8_0(.dout(w_dff_A_qXG8zpi81_0),.din(w_dff_A_aquxKKMG8_0),.clk(gclk));
	jdff dff_A_vzFMzJ0s6_0(.dout(w_dff_A_aquxKKMG8_0),.din(w_dff_A_vzFMzJ0s6_0),.clk(gclk));
	jdff dff_A_8MUZIVM40_0(.dout(w_dff_A_vzFMzJ0s6_0),.din(w_dff_A_8MUZIVM40_0),.clk(gclk));
	jdff dff_A_8F4L9rEQ2_0(.dout(w_dff_A_8MUZIVM40_0),.din(w_dff_A_8F4L9rEQ2_0),.clk(gclk));
	jdff dff_A_C0gpur6a9_0(.dout(w_dff_A_8F4L9rEQ2_0),.din(w_dff_A_C0gpur6a9_0),.clk(gclk));
	jdff dff_A_fLHyWBkp6_0(.dout(w_dff_A_C0gpur6a9_0),.din(w_dff_A_fLHyWBkp6_0),.clk(gclk));
	jdff dff_A_SVCRgDDz1_0(.dout(w_dff_A_fLHyWBkp6_0),.din(w_dff_A_SVCRgDDz1_0),.clk(gclk));
	jdff dff_A_NSGXEAav9_0(.dout(w_dff_A_SVCRgDDz1_0),.din(w_dff_A_NSGXEAav9_0),.clk(gclk));
	jdff dff_A_pTPvviVi8_0(.dout(w_dff_A_NSGXEAav9_0),.din(w_dff_A_pTPvviVi8_0),.clk(gclk));
	jdff dff_A_8FZZKRYL6_1(.dout(w_n219_0[1]),.din(w_dff_A_8FZZKRYL6_1),.clk(gclk));
	jdff dff_A_Md7vrpUJ3_1(.dout(w_dff_A_8FZZKRYL6_1),.din(w_dff_A_Md7vrpUJ3_1),.clk(gclk));
	jdff dff_A_iVHeoyJr4_1(.dout(w_dff_A_Md7vrpUJ3_1),.din(w_dff_A_iVHeoyJr4_1),.clk(gclk));
	jdff dff_A_d54mL2Om9_1(.dout(w_dff_A_iVHeoyJr4_1),.din(w_dff_A_d54mL2Om9_1),.clk(gclk));
	jdff dff_A_K09wiWK30_0(.dout(w_n217_0[0]),.din(w_dff_A_K09wiWK30_0),.clk(gclk));
	jdff dff_A_Buj8wYlS7_0(.dout(w_dff_A_K09wiWK30_0),.din(w_dff_A_Buj8wYlS7_0),.clk(gclk));
	jdff dff_A_KYC09Ls34_0(.dout(w_dff_A_Buj8wYlS7_0),.din(w_dff_A_KYC09Ls34_0),.clk(gclk));
	jdff dff_A_7fQt6V3F4_0(.dout(w_dff_A_KYC09Ls34_0),.din(w_dff_A_7fQt6V3F4_0),.clk(gclk));
	jdff dff_A_lTgL6P0O2_0(.dout(w_dff_A_7fQt6V3F4_0),.din(w_dff_A_lTgL6P0O2_0),.clk(gclk));
	jdff dff_A_1lx8uWHB5_0(.dout(w_dff_A_lTgL6P0O2_0),.din(w_dff_A_1lx8uWHB5_0),.clk(gclk));
	jdff dff_A_8CavIptA0_0(.dout(w_dff_A_1lx8uWHB5_0),.din(w_dff_A_8CavIptA0_0),.clk(gclk));
	jdff dff_A_aHV4aXfV4_0(.dout(w_dff_A_8CavIptA0_0),.din(w_dff_A_aHV4aXfV4_0),.clk(gclk));
	jdff dff_A_NEDzp6qH5_0(.dout(w_dff_A_aHV4aXfV4_0),.din(w_dff_A_NEDzp6qH5_0),.clk(gclk));
	jdff dff_A_0nqLD8yi9_0(.dout(w_dff_A_NEDzp6qH5_0),.din(w_dff_A_0nqLD8yi9_0),.clk(gclk));
	jdff dff_A_oe4tlPCg9_0(.dout(w_dff_A_0nqLD8yi9_0),.din(w_dff_A_oe4tlPCg9_0),.clk(gclk));
	jdff dff_B_2YcemIQ92_2(.din(n217),.dout(w_dff_B_2YcemIQ92_2),.clk(gclk));
	jdff dff_B_tiulCnbL2_2(.din(w_dff_B_2YcemIQ92_2),.dout(w_dff_B_tiulCnbL2_2),.clk(gclk));
	jdff dff_B_QmYJJC3n9_2(.din(w_dff_B_tiulCnbL2_2),.dout(w_dff_B_QmYJJC3n9_2),.clk(gclk));
	jdff dff_B_1u29ajOh1_2(.din(w_dff_B_QmYJJC3n9_2),.dout(w_dff_B_1u29ajOh1_2),.clk(gclk));
	jdff dff_B_MywoQ7js6_2(.din(w_dff_B_1u29ajOh1_2),.dout(w_dff_B_MywoQ7js6_2),.clk(gclk));
	jdff dff_B_s9cZoVTR0_2(.din(w_dff_B_MywoQ7js6_2),.dout(w_dff_B_s9cZoVTR0_2),.clk(gclk));
	jdff dff_B_FK9puWpO4_2(.din(w_dff_B_s9cZoVTR0_2),.dout(w_dff_B_FK9puWpO4_2),.clk(gclk));
	jdff dff_B_FVREnZD71_2(.din(w_dff_B_FK9puWpO4_2),.dout(w_dff_B_FVREnZD71_2),.clk(gclk));
	jdff dff_A_cQwLVOFm7_0(.dout(w_G40gat_0[0]),.din(w_dff_A_cQwLVOFm7_0),.clk(gclk));
	jdff dff_A_m7jWDz0S8_0(.dout(w_dff_A_cQwLVOFm7_0),.din(w_dff_A_m7jWDz0S8_0),.clk(gclk));
	jdff dff_A_DW59HpH40_0(.dout(w_dff_A_m7jWDz0S8_0),.din(w_dff_A_DW59HpH40_0),.clk(gclk));
	jdff dff_A_0KVgAVg85_0(.dout(w_dff_A_DW59HpH40_0),.din(w_dff_A_0KVgAVg85_0),.clk(gclk));
	jdff dff_A_J9e7HbqY0_0(.dout(w_dff_A_0KVgAVg85_0),.din(w_dff_A_J9e7HbqY0_0),.clk(gclk));
	jdff dff_A_vKW4BJrW4_0(.dout(w_dff_A_J9e7HbqY0_0),.din(w_dff_A_vKW4BJrW4_0),.clk(gclk));
	jdff dff_A_EiWeU5AG8_0(.dout(w_dff_A_vKW4BJrW4_0),.din(w_dff_A_EiWeU5AG8_0),.clk(gclk));
	jdff dff_A_DysaCDw63_0(.dout(w_dff_A_EiWeU5AG8_0),.din(w_dff_A_DysaCDw63_0),.clk(gclk));
	jdff dff_A_nUqJJRf63_0(.dout(w_dff_A_DysaCDw63_0),.din(w_dff_A_nUqJJRf63_0),.clk(gclk));
	jdff dff_A_MZWkJju34_0(.dout(w_dff_A_nUqJJRf63_0),.din(w_dff_A_MZWkJju34_0),.clk(gclk));
	jdff dff_A_YHUwgax27_0(.dout(w_dff_A_MZWkJju34_0),.din(w_dff_A_YHUwgax27_0),.clk(gclk));
	jdff dff_A_92M2Zl8z8_0(.dout(w_dff_A_YHUwgax27_0),.din(w_dff_A_92M2Zl8z8_0),.clk(gclk));
	jdff dff_A_JQajJs659_0(.dout(w_dff_A_92M2Zl8z8_0),.din(w_dff_A_JQajJs659_0),.clk(gclk));
	jdff dff_A_C34rz9Fg0_0(.dout(w_dff_A_JQajJs659_0),.din(w_dff_A_C34rz9Fg0_0),.clk(gclk));
	jdff dff_A_FMGlxFBl8_0(.dout(w_dff_A_C34rz9Fg0_0),.din(w_dff_A_FMGlxFBl8_0),.clk(gclk));
	jdff dff_A_3UWegJy00_0(.dout(w_dff_A_FMGlxFBl8_0),.din(w_dff_A_3UWegJy00_0),.clk(gclk));
	jdff dff_A_oqTTcQyO7_0(.dout(w_dff_A_3UWegJy00_0),.din(w_dff_A_oqTTcQyO7_0),.clk(gclk));
	jdff dff_A_prfLRcRV9_0(.dout(w_dff_A_oqTTcQyO7_0),.din(w_dff_A_prfLRcRV9_0),.clk(gclk));
	jdff dff_A_LB8w7xGO3_0(.dout(w_dff_A_prfLRcRV9_0),.din(w_dff_A_LB8w7xGO3_0),.clk(gclk));
	jdff dff_A_cF2UM3na6_0(.dout(w_dff_A_LB8w7xGO3_0),.din(w_dff_A_cF2UM3na6_0),.clk(gclk));
	jdff dff_B_JAtH6QYN6_1(.din(n214),.dout(w_dff_B_JAtH6QYN6_1),.clk(gclk));
	jdff dff_B_hknoBpDP2_1(.din(w_dff_B_JAtH6QYN6_1),.dout(w_dff_B_hknoBpDP2_1),.clk(gclk));
	jdff dff_B_DlPlRZMf2_1(.din(w_dff_B_hknoBpDP2_1),.dout(w_dff_B_DlPlRZMf2_1),.clk(gclk));
	jdff dff_B_Oi1GTYA27_1(.din(w_dff_B_DlPlRZMf2_1),.dout(w_dff_B_Oi1GTYA27_1),.clk(gclk));
	jdff dff_B_S0fUgJk15_1(.din(w_dff_B_Oi1GTYA27_1),.dout(w_dff_B_S0fUgJk15_1),.clk(gclk));
	jdff dff_B_OTZRNQks9_1(.din(w_dff_B_S0fUgJk15_1),.dout(w_dff_B_OTZRNQks9_1),.clk(gclk));
	jdff dff_B_14PyE8ru3_1(.din(w_dff_B_OTZRNQks9_1),.dout(w_dff_B_14PyE8ru3_1),.clk(gclk));
	jdff dff_B_5iSKiwbu5_1(.din(w_dff_B_14PyE8ru3_1),.dout(w_dff_B_5iSKiwbu5_1),.clk(gclk));
	jdff dff_B_lmSBl0DE6_1(.din(w_dff_B_5iSKiwbu5_1),.dout(w_dff_B_lmSBl0DE6_1),.clk(gclk));
	jdff dff_B_QaaHamPu0_1(.din(w_dff_B_lmSBl0DE6_1),.dout(w_dff_B_QaaHamPu0_1),.clk(gclk));
	jdff dff_B_sg2gjBky1_1(.din(w_dff_B_QaaHamPu0_1),.dout(w_dff_B_sg2gjBky1_1),.clk(gclk));
	jdff dff_B_9ISUfuz87_1(.din(w_dff_B_sg2gjBky1_1),.dout(w_dff_B_9ISUfuz87_1),.clk(gclk));
	jdff dff_B_ip6L2EgA2_1(.din(n209),.dout(w_dff_B_ip6L2EgA2_1),.clk(gclk));
	jdff dff_B_9un0dYnS5_1(.din(w_dff_B_ip6L2EgA2_1),.dout(w_dff_B_9un0dYnS5_1),.clk(gclk));
	jdff dff_B_pHw88pEo3_1(.din(w_dff_B_9un0dYnS5_1),.dout(w_dff_B_pHw88pEo3_1),.clk(gclk));
	jdff dff_B_BkoH1c7b4_1(.din(w_dff_B_pHw88pEo3_1),.dout(w_dff_B_BkoH1c7b4_1),.clk(gclk));
	jdff dff_B_17QKc4032_1(.din(w_dff_B_BkoH1c7b4_1),.dout(w_dff_B_17QKc4032_1),.clk(gclk));
	jdff dff_B_lY72b7Xi2_1(.din(w_dff_B_17QKc4032_1),.dout(w_dff_B_lY72b7Xi2_1),.clk(gclk));
	jdff dff_B_uI2FUQZx0_1(.din(w_dff_B_lY72b7Xi2_1),.dout(w_dff_B_uI2FUQZx0_1),.clk(gclk));
	jdff dff_B_mdbxgMUr0_1(.din(w_dff_B_uI2FUQZx0_1),.dout(w_dff_B_mdbxgMUr0_1),.clk(gclk));
	jdff dff_B_SxTdgAXJ1_1(.din(w_dff_B_mdbxgMUr0_1),.dout(w_dff_B_SxTdgAXJ1_1),.clk(gclk));
	jdff dff_B_3132phCB1_1(.din(w_dff_B_SxTdgAXJ1_1),.dout(w_dff_B_3132phCB1_1),.clk(gclk));
	jdff dff_B_oeRnJ07C6_1(.din(w_dff_B_3132phCB1_1),.dout(w_dff_B_oeRnJ07C6_1),.clk(gclk));
	jdff dff_B_iun8o7aA0_1(.din(w_dff_B_oeRnJ07C6_1),.dout(w_dff_B_iun8o7aA0_1),.clk(gclk));
	jdff dff_B_HCkoYt0G3_1(.din(w_dff_B_iun8o7aA0_1),.dout(w_dff_B_HCkoYt0G3_1),.clk(gclk));
	jdff dff_B_uTCzO6Hi1_1(.din(w_dff_B_HCkoYt0G3_1),.dout(w_dff_B_uTCzO6Hi1_1),.clk(gclk));
	jdff dff_A_EGoBSwq17_0(.dout(w_G14gat_0[0]),.din(w_dff_A_EGoBSwq17_0),.clk(gclk));
	jdff dff_A_2xI4MMCA4_0(.dout(w_dff_A_EGoBSwq17_0),.din(w_dff_A_2xI4MMCA4_0),.clk(gclk));
	jdff dff_A_nKU2a0Vu7_0(.dout(w_dff_A_2xI4MMCA4_0),.din(w_dff_A_nKU2a0Vu7_0),.clk(gclk));
	jdff dff_A_yyqq8xVU6_0(.dout(w_dff_A_nKU2a0Vu7_0),.din(w_dff_A_yyqq8xVU6_0),.clk(gclk));
	jdff dff_A_AXZdTIEi1_0(.dout(w_dff_A_yyqq8xVU6_0),.din(w_dff_A_AXZdTIEi1_0),.clk(gclk));
	jdff dff_A_FVHJF5re9_0(.dout(w_dff_A_AXZdTIEi1_0),.din(w_dff_A_FVHJF5re9_0),.clk(gclk));
	jdff dff_A_1h2Dwb9x6_0(.dout(w_dff_A_FVHJF5re9_0),.din(w_dff_A_1h2Dwb9x6_0),.clk(gclk));
	jdff dff_A_WcHWZvVs0_0(.dout(w_dff_A_1h2Dwb9x6_0),.din(w_dff_A_WcHWZvVs0_0),.clk(gclk));
	jdff dff_A_3SBLw8T22_0(.dout(w_dff_A_WcHWZvVs0_0),.din(w_dff_A_3SBLw8T22_0),.clk(gclk));
	jdff dff_A_05ial6b11_0(.dout(w_dff_A_3SBLw8T22_0),.din(w_dff_A_05ial6b11_0),.clk(gclk));
	jdff dff_A_xDYdVTql6_0(.dout(w_dff_A_05ial6b11_0),.din(w_dff_A_xDYdVTql6_0),.clk(gclk));
	jdff dff_A_fqOMxiy43_0(.dout(w_dff_A_xDYdVTql6_0),.din(w_dff_A_fqOMxiy43_0),.clk(gclk));
	jdff dff_A_CSfFWcDW9_0(.dout(w_dff_A_fqOMxiy43_0),.din(w_dff_A_CSfFWcDW9_0),.clk(gclk));
	jdff dff_A_vupmUNby3_0(.dout(w_dff_A_CSfFWcDW9_0),.din(w_dff_A_vupmUNby3_0),.clk(gclk));
	jdff dff_A_ZHfG6End6_0(.dout(w_dff_A_vupmUNby3_0),.din(w_dff_A_ZHfG6End6_0),.clk(gclk));
	jdff dff_A_4B1Y14dG6_1(.dout(w_G14gat_0[1]),.din(w_dff_A_4B1Y14dG6_1),.clk(gclk));
	jdff dff_A_fY67RCm50_1(.dout(w_dff_A_4B1Y14dG6_1),.din(w_dff_A_fY67RCm50_1),.clk(gclk));
	jdff dff_A_5aq5BgUk0_1(.dout(w_dff_A_fY67RCm50_1),.din(w_dff_A_5aq5BgUk0_1),.clk(gclk));
	jdff dff_A_5WXQxHvf4_1(.dout(w_dff_A_5aq5BgUk0_1),.din(w_dff_A_5WXQxHvf4_1),.clk(gclk));
	jdff dff_A_N7RMsra07_1(.dout(w_dff_A_5WXQxHvf4_1),.din(w_dff_A_N7RMsra07_1),.clk(gclk));
	jdff dff_A_ttO0wQNS8_1(.dout(w_dff_A_N7RMsra07_1),.din(w_dff_A_ttO0wQNS8_1),.clk(gclk));
	jdff dff_A_hvodjvo19_1(.dout(w_dff_A_ttO0wQNS8_1),.din(w_dff_A_hvodjvo19_1),.clk(gclk));
	jdff dff_A_9Tt24nFE8_1(.dout(w_dff_A_hvodjvo19_1),.din(w_dff_A_9Tt24nFE8_1),.clk(gclk));
	jdff dff_A_qG53VjYE0_1(.dout(w_dff_A_9Tt24nFE8_1),.din(w_dff_A_qG53VjYE0_1),.clk(gclk));
	jdff dff_A_MCyEELYN1_1(.dout(w_dff_A_qG53VjYE0_1),.din(w_dff_A_MCyEELYN1_1),.clk(gclk));
	jdff dff_A_CXtccuCO5_1(.dout(w_dff_A_MCyEELYN1_1),.din(w_dff_A_CXtccuCO5_1),.clk(gclk));
	jdff dff_A_OXbuJOhc8_1(.dout(w_dff_A_CXtccuCO5_1),.din(w_dff_A_OXbuJOhc8_1),.clk(gclk));
	jdff dff_A_Pg9Yihf36_1(.dout(w_dff_A_OXbuJOhc8_1),.din(w_dff_A_Pg9Yihf36_1),.clk(gclk));
	jdff dff_A_2txbwMG71_1(.dout(w_dff_A_Pg9Yihf36_1),.din(w_dff_A_2txbwMG71_1),.clk(gclk));
	jdff dff_A_MaAgopZo4_1(.dout(w_dff_A_2txbwMG71_1),.din(w_dff_A_MaAgopZo4_1),.clk(gclk));
	jdff dff_A_bKmBPZRg6_1(.dout(w_dff_A_MaAgopZo4_1),.din(w_dff_A_bKmBPZRg6_1),.clk(gclk));
	jdff dff_A_OxR6szJ24_1(.dout(w_dff_A_bKmBPZRg6_1),.din(w_dff_A_OxR6szJ24_1),.clk(gclk));
	jdff dff_A_ZVkNtnPK5_1(.dout(w_dff_A_OxR6szJ24_1),.din(w_dff_A_ZVkNtnPK5_1),.clk(gclk));
	jdff dff_A_jU2YAEAb7_1(.dout(w_dff_A_ZVkNtnPK5_1),.din(w_dff_A_jU2YAEAb7_1),.clk(gclk));
	jdff dff_A_SRPEcVSu0_1(.dout(w_dff_A_jU2YAEAb7_1),.din(w_dff_A_SRPEcVSu0_1),.clk(gclk));
	jdff dff_A_GIavFXJY4_0(.dout(w_n205_0[0]),.din(w_dff_A_GIavFXJY4_0),.clk(gclk));
	jdff dff_A_h5nScqoq6_0(.dout(w_dff_A_GIavFXJY4_0),.din(w_dff_A_h5nScqoq6_0),.clk(gclk));
	jdff dff_A_bmkzxTd32_0(.dout(w_dff_A_h5nScqoq6_0),.din(w_dff_A_bmkzxTd32_0),.clk(gclk));
	jdff dff_A_t6BzmpDP7_0(.dout(w_dff_A_bmkzxTd32_0),.din(w_dff_A_t6BzmpDP7_0),.clk(gclk));
	jdff dff_A_bSlRV5rd6_0(.dout(w_dff_A_t6BzmpDP7_0),.din(w_dff_A_bSlRV5rd6_0),.clk(gclk));
	jdff dff_A_EaVkdNfv5_0(.dout(w_dff_A_bSlRV5rd6_0),.din(w_dff_A_EaVkdNfv5_0),.clk(gclk));
	jdff dff_B_OFiT3GSp7_2(.din(n205),.dout(w_dff_B_OFiT3GSp7_2),.clk(gclk));
	jdff dff_B_RVlDbZ9m5_2(.din(w_dff_B_OFiT3GSp7_2),.dout(w_dff_B_RVlDbZ9m5_2),.clk(gclk));
	jdff dff_B_cC7ubkQR1_2(.din(w_dff_B_RVlDbZ9m5_2),.dout(w_dff_B_cC7ubkQR1_2),.clk(gclk));
	jdff dff_B_mQCHZgxH2_2(.din(w_dff_B_cC7ubkQR1_2),.dout(w_dff_B_mQCHZgxH2_2),.clk(gclk));
	jdff dff_B_2HGfSuSX4_2(.din(w_dff_B_mQCHZgxH2_2),.dout(w_dff_B_2HGfSuSX4_2),.clk(gclk));
	jdff dff_B_tbPTYDfA0_2(.din(w_dff_B_2HGfSuSX4_2),.dout(w_dff_B_tbPTYDfA0_2),.clk(gclk));
	jdff dff_B_wyfG7C8O2_2(.din(w_dff_B_tbPTYDfA0_2),.dout(w_dff_B_wyfG7C8O2_2),.clk(gclk));
	jdff dff_B_gGq2oYPE6_2(.din(w_dff_B_wyfG7C8O2_2),.dout(w_dff_B_gGq2oYPE6_2),.clk(gclk));
	jdff dff_B_KiPOa9Mz8_2(.din(w_dff_B_gGq2oYPE6_2),.dout(w_dff_B_KiPOa9Mz8_2),.clk(gclk));
	jdff dff_B_qkYuge6v6_2(.din(w_dff_B_KiPOa9Mz8_2),.dout(w_dff_B_qkYuge6v6_2),.clk(gclk));
	jdff dff_B_y1rL8AYV0_2(.din(w_dff_B_qkYuge6v6_2),.dout(w_dff_B_y1rL8AYV0_2),.clk(gclk));
	jdff dff_B_A10GNPnt2_2(.din(w_dff_B_y1rL8AYV0_2),.dout(w_dff_B_A10GNPnt2_2),.clk(gclk));
	jdff dff_B_FbCWni4c0_2(.din(w_dff_B_A10GNPnt2_2),.dout(w_dff_B_FbCWni4c0_2),.clk(gclk));
	jdff dff_A_iu1WqPGS5_0(.dout(w_G92gat_0[0]),.din(w_dff_A_iu1WqPGS5_0),.clk(gclk));
	jdff dff_A_QB91sCtJ1_0(.dout(w_dff_A_iu1WqPGS5_0),.din(w_dff_A_QB91sCtJ1_0),.clk(gclk));
	jdff dff_A_sMMDcdY31_0(.dout(w_dff_A_QB91sCtJ1_0),.din(w_dff_A_sMMDcdY31_0),.clk(gclk));
	jdff dff_A_ayzV43KE6_0(.dout(w_dff_A_sMMDcdY31_0),.din(w_dff_A_ayzV43KE6_0),.clk(gclk));
	jdff dff_A_wcIEbD2x8_0(.dout(w_dff_A_ayzV43KE6_0),.din(w_dff_A_wcIEbD2x8_0),.clk(gclk));
	jdff dff_A_HqxwDOul0_0(.dout(w_dff_A_wcIEbD2x8_0),.din(w_dff_A_HqxwDOul0_0),.clk(gclk));
	jdff dff_A_VDAhH8S32_0(.dout(w_dff_A_HqxwDOul0_0),.din(w_dff_A_VDAhH8S32_0),.clk(gclk));
	jdff dff_A_UHZ0AsGE3_0(.dout(w_dff_A_VDAhH8S32_0),.din(w_dff_A_UHZ0AsGE3_0),.clk(gclk));
	jdff dff_A_4DJfSLme3_0(.dout(w_dff_A_UHZ0AsGE3_0),.din(w_dff_A_4DJfSLme3_0),.clk(gclk));
	jdff dff_A_Lwyjt1Bi4_0(.dout(w_dff_A_4DJfSLme3_0),.din(w_dff_A_Lwyjt1Bi4_0),.clk(gclk));
	jdff dff_A_TJWqEGNl2_0(.dout(w_dff_A_Lwyjt1Bi4_0),.din(w_dff_A_TJWqEGNl2_0),.clk(gclk));
	jdff dff_A_9mjOUV812_0(.dout(w_dff_A_TJWqEGNl2_0),.din(w_dff_A_9mjOUV812_0),.clk(gclk));
	jdff dff_A_VwzK9wRe3_0(.dout(w_dff_A_9mjOUV812_0),.din(w_dff_A_VwzK9wRe3_0),.clk(gclk));
	jdff dff_A_1VuSXTht4_0(.dout(w_dff_A_VwzK9wRe3_0),.din(w_dff_A_1VuSXTht4_0),.clk(gclk));
	jdff dff_A_16Mc6rX52_0(.dout(w_dff_A_1VuSXTht4_0),.din(w_dff_A_16Mc6rX52_0),.clk(gclk));
	jdff dff_A_ixNMUFVr3_0(.dout(w_dff_A_16Mc6rX52_0),.din(w_dff_A_ixNMUFVr3_0),.clk(gclk));
	jdff dff_A_x7kcPeyr0_0(.dout(w_dff_A_ixNMUFVr3_0),.din(w_dff_A_x7kcPeyr0_0),.clk(gclk));
	jdff dff_A_PtVh3klS2_0(.dout(w_dff_A_x7kcPeyr0_0),.din(w_dff_A_PtVh3klS2_0),.clk(gclk));
	jdff dff_A_tnePtMzo9_0(.dout(w_dff_A_PtVh3klS2_0),.din(w_dff_A_tnePtMzo9_0),.clk(gclk));
	jdff dff_A_6AlgyhNC8_0(.dout(w_dff_A_tnePtMzo9_0),.din(w_dff_A_6AlgyhNC8_0),.clk(gclk));
	jdff dff_A_As8JnspT9_1(.dout(w_G92gat_0[1]),.din(w_dff_A_As8JnspT9_1),.clk(gclk));
	jdff dff_A_MqMPAM8g8_1(.dout(w_dff_A_As8JnspT9_1),.din(w_dff_A_MqMPAM8g8_1),.clk(gclk));
	jdff dff_A_ZatDco8P9_1(.dout(w_dff_A_MqMPAM8g8_1),.din(w_dff_A_ZatDco8P9_1),.clk(gclk));
	jdff dff_A_86c3BzAz2_1(.dout(w_dff_A_ZatDco8P9_1),.din(w_dff_A_86c3BzAz2_1),.clk(gclk));
	jdff dff_A_KQaawdCQ0_1(.dout(w_dff_A_86c3BzAz2_1),.din(w_dff_A_KQaawdCQ0_1),.clk(gclk));
	jdff dff_A_xrOA8BGO2_1(.dout(w_dff_A_KQaawdCQ0_1),.din(w_dff_A_xrOA8BGO2_1),.clk(gclk));
	jdff dff_A_dZYOYQUF7_1(.dout(w_dff_A_xrOA8BGO2_1),.din(w_dff_A_dZYOYQUF7_1),.clk(gclk));
	jdff dff_A_fVk5TWhd6_1(.dout(w_dff_A_dZYOYQUF7_1),.din(w_dff_A_fVk5TWhd6_1),.clk(gclk));
	jdff dff_A_nZQQ6A4D3_1(.dout(w_dff_A_fVk5TWhd6_1),.din(w_dff_A_nZQQ6A4D3_1),.clk(gclk));
	jdff dff_A_G9tl59HE2_1(.dout(w_dff_A_nZQQ6A4D3_1),.din(w_dff_A_G9tl59HE2_1),.clk(gclk));
	jdff dff_A_Y957lquf4_1(.dout(w_dff_A_G9tl59HE2_1),.din(w_dff_A_Y957lquf4_1),.clk(gclk));
	jdff dff_A_VB0sQ4Hs6_1(.dout(w_dff_A_Y957lquf4_1),.din(w_dff_A_VB0sQ4Hs6_1),.clk(gclk));
	jdff dff_A_C7BTkScG1_1(.dout(w_dff_A_VB0sQ4Hs6_1),.din(w_dff_A_C7BTkScG1_1),.clk(gclk));
	jdff dff_A_pVnNe7Ql2_1(.dout(w_dff_A_C7BTkScG1_1),.din(w_dff_A_pVnNe7Ql2_1),.clk(gclk));
	jdff dff_A_k4Y51fI90_0(.dout(w_n204_0[0]),.din(w_dff_A_k4Y51fI90_0),.clk(gclk));
	jdff dff_A_ZEYuEmjA2_0(.dout(w_dff_A_k4Y51fI90_0),.din(w_dff_A_ZEYuEmjA2_0),.clk(gclk));
	jdff dff_A_1kLqxltu3_0(.dout(w_dff_A_ZEYuEmjA2_0),.din(w_dff_A_1kLqxltu3_0),.clk(gclk));
	jdff dff_A_femnjQoD9_0(.dout(w_dff_A_1kLqxltu3_0),.din(w_dff_A_femnjQoD9_0),.clk(gclk));
	jdff dff_A_iN4N0kGU2_0(.dout(w_dff_A_femnjQoD9_0),.din(w_dff_A_iN4N0kGU2_0),.clk(gclk));
	jdff dff_A_fS7LI9u52_0(.dout(w_dff_A_iN4N0kGU2_0),.din(w_dff_A_fS7LI9u52_0),.clk(gclk));
	jdff dff_A_PXdOYgUc3_0(.dout(w_n198_0[0]),.din(w_dff_A_PXdOYgUc3_0),.clk(gclk));
	jdff dff_A_9EHkEeAd8_0(.dout(w_dff_A_PXdOYgUc3_0),.din(w_dff_A_9EHkEeAd8_0),.clk(gclk));
	jdff dff_A_Kkzt62QM3_0(.dout(w_dff_A_9EHkEeAd8_0),.din(w_dff_A_Kkzt62QM3_0),.clk(gclk));
	jdff dff_A_WeIUFYL15_0(.dout(w_dff_A_Kkzt62QM3_0),.din(w_dff_A_WeIUFYL15_0),.clk(gclk));
	jdff dff_A_x4Avr8QU9_0(.dout(w_dff_A_WeIUFYL15_0),.din(w_dff_A_x4Avr8QU9_0),.clk(gclk));
	jdff dff_A_5vpnn1Hd2_0(.dout(w_dff_A_x4Avr8QU9_0),.din(w_dff_A_5vpnn1Hd2_0),.clk(gclk));
	jdff dff_B_aM77vvQf2_2(.din(n198),.dout(w_dff_B_aM77vvQf2_2),.clk(gclk));
	jdff dff_B_4yFEp7qB2_2(.din(w_dff_B_aM77vvQf2_2),.dout(w_dff_B_4yFEp7qB2_2),.clk(gclk));
	jdff dff_B_Gwg8VPr55_2(.din(w_dff_B_4yFEp7qB2_2),.dout(w_dff_B_Gwg8VPr55_2),.clk(gclk));
	jdff dff_B_s9r5tMvl0_2(.din(w_dff_B_Gwg8VPr55_2),.dout(w_dff_B_s9r5tMvl0_2),.clk(gclk));
	jdff dff_B_8Xzm0hvr0_2(.din(w_dff_B_s9r5tMvl0_2),.dout(w_dff_B_8Xzm0hvr0_2),.clk(gclk));
	jdff dff_B_lY5v2AR60_2(.din(w_dff_B_8Xzm0hvr0_2),.dout(w_dff_B_lY5v2AR60_2),.clk(gclk));
	jdff dff_B_HoljFIyH1_2(.din(w_dff_B_lY5v2AR60_2),.dout(w_dff_B_HoljFIyH1_2),.clk(gclk));
	jdff dff_B_7w6Ty0cH2_2(.din(w_dff_B_HoljFIyH1_2),.dout(w_dff_B_7w6Ty0cH2_2),.clk(gclk));
	jdff dff_B_KJLzsaIP2_2(.din(w_dff_B_7w6Ty0cH2_2),.dout(w_dff_B_KJLzsaIP2_2),.clk(gclk));
	jdff dff_B_2neI1Evm1_2(.din(w_dff_B_KJLzsaIP2_2),.dout(w_dff_B_2neI1Evm1_2),.clk(gclk));
	jdff dff_B_iHgdOBnX0_2(.din(w_dff_B_2neI1Evm1_2),.dout(w_dff_B_iHgdOBnX0_2),.clk(gclk));
	jdff dff_B_gKPkkoLp1_2(.din(w_dff_B_iHgdOBnX0_2),.dout(w_dff_B_gKPkkoLp1_2),.clk(gclk));
	jdff dff_B_DTbtNB9T8_2(.din(w_dff_B_gKPkkoLp1_2),.dout(w_dff_B_DTbtNB9T8_2),.clk(gclk));
	jdff dff_A_RBEnPNtx5_0(.dout(w_G27gat_0[0]),.din(w_dff_A_RBEnPNtx5_0),.clk(gclk));
	jdff dff_A_UxsZlsHM9_0(.dout(w_dff_A_RBEnPNtx5_0),.din(w_dff_A_UxsZlsHM9_0),.clk(gclk));
	jdff dff_A_CVFKzrvw5_0(.dout(w_dff_A_UxsZlsHM9_0),.din(w_dff_A_CVFKzrvw5_0),.clk(gclk));
	jdff dff_A_Ffcnbr041_0(.dout(w_dff_A_CVFKzrvw5_0),.din(w_dff_A_Ffcnbr041_0),.clk(gclk));
	jdff dff_A_FVdGMKIu8_0(.dout(w_dff_A_Ffcnbr041_0),.din(w_dff_A_FVdGMKIu8_0),.clk(gclk));
	jdff dff_A_KxsXErZn8_0(.dout(w_dff_A_FVdGMKIu8_0),.din(w_dff_A_KxsXErZn8_0),.clk(gclk));
	jdff dff_A_G03M6b2O4_0(.dout(w_dff_A_KxsXErZn8_0),.din(w_dff_A_G03M6b2O4_0),.clk(gclk));
	jdff dff_A_RMwHhFwb4_0(.dout(w_dff_A_G03M6b2O4_0),.din(w_dff_A_RMwHhFwb4_0),.clk(gclk));
	jdff dff_A_1iaXrsKi2_0(.dout(w_dff_A_RMwHhFwb4_0),.din(w_dff_A_1iaXrsKi2_0),.clk(gclk));
	jdff dff_A_PQW8m0Zz5_0(.dout(w_dff_A_1iaXrsKi2_0),.din(w_dff_A_PQW8m0Zz5_0),.clk(gclk));
	jdff dff_A_HhqMSUCE3_0(.dout(w_dff_A_PQW8m0Zz5_0),.din(w_dff_A_HhqMSUCE3_0),.clk(gclk));
	jdff dff_A_QAFcLRcE5_0(.dout(w_dff_A_HhqMSUCE3_0),.din(w_dff_A_QAFcLRcE5_0),.clk(gclk));
	jdff dff_A_PM6y6Rac5_0(.dout(w_dff_A_QAFcLRcE5_0),.din(w_dff_A_PM6y6Rac5_0),.clk(gclk));
	jdff dff_A_fuz1QEUW2_0(.dout(w_dff_A_PM6y6Rac5_0),.din(w_dff_A_fuz1QEUW2_0),.clk(gclk));
	jdff dff_A_QVMlWibB4_0(.dout(w_n197_0[0]),.din(w_dff_A_QVMlWibB4_0),.clk(gclk));
	jdff dff_A_TsTr8HVb4_0(.dout(w_dff_A_QVMlWibB4_0),.din(w_dff_A_TsTr8HVb4_0),.clk(gclk));
	jdff dff_A_FBjetoBE9_0(.dout(w_dff_A_TsTr8HVb4_0),.din(w_dff_A_FBjetoBE9_0),.clk(gclk));
	jdff dff_A_EdBUKRpG0_0(.dout(w_dff_A_FBjetoBE9_0),.din(w_dff_A_EdBUKRpG0_0),.clk(gclk));
	jdff dff_A_nT7qtMo65_0(.dout(w_dff_A_EdBUKRpG0_0),.din(w_dff_A_nT7qtMo65_0),.clk(gclk));
	jdff dff_A_D4Qlff1r3_0(.dout(w_dff_A_nT7qtMo65_0),.din(w_dff_A_D4Qlff1r3_0),.clk(gclk));
	jdff dff_A_RPite0FH3_1(.dout(w_n193_0[1]),.din(w_dff_A_RPite0FH3_1),.clk(gclk));
	jdff dff_A_EkWQoan84_1(.dout(w_dff_A_RPite0FH3_1),.din(w_dff_A_EkWQoan84_1),.clk(gclk));
	jdff dff_A_YD5yqhga5_1(.dout(w_dff_A_EkWQoan84_1),.din(w_dff_A_YD5yqhga5_1),.clk(gclk));
	jdff dff_A_MDTRry8g2_1(.dout(w_dff_A_YD5yqhga5_1),.din(w_dff_A_MDTRry8g2_1),.clk(gclk));
	jdff dff_A_xqOc8yYE8_1(.dout(w_dff_A_MDTRry8g2_1),.din(w_dff_A_xqOc8yYE8_1),.clk(gclk));
	jdff dff_A_AnpFQgZC3_1(.dout(w_dff_A_xqOc8yYE8_1),.din(w_dff_A_AnpFQgZC3_1),.clk(gclk));
	jdff dff_A_7K0OEzMt0_1(.dout(w_dff_A_AnpFQgZC3_1),.din(w_dff_A_7K0OEzMt0_1),.clk(gclk));
	jdff dff_B_PEalnbEV7_0(.din(n192),.dout(w_dff_B_PEalnbEV7_0),.clk(gclk));
	jdff dff_B_ziLYTqk45_0(.din(w_dff_B_PEalnbEV7_0),.dout(w_dff_B_ziLYTqk45_0),.clk(gclk));
	jdff dff_B_mjnAvtN12_0(.din(w_dff_B_ziLYTqk45_0),.dout(w_dff_B_mjnAvtN12_0),.clk(gclk));
	jdff dff_B_EJ7mrd9b3_0(.din(w_dff_B_mjnAvtN12_0),.dout(w_dff_B_EJ7mrd9b3_0),.clk(gclk));
	jdff dff_B_6ncqurZe4_0(.din(w_dff_B_EJ7mrd9b3_0),.dout(w_dff_B_6ncqurZe4_0),.clk(gclk));
	jdff dff_A_ND367Ak01_0(.dout(w_n191_0[0]),.din(w_dff_A_ND367Ak01_0),.clk(gclk));
	jdff dff_A_z15boVMH8_0(.dout(w_dff_A_ND367Ak01_0),.din(w_dff_A_z15boVMH8_0),.clk(gclk));
	jdff dff_A_FVMnuiyI7_0(.dout(w_dff_A_z15boVMH8_0),.din(w_dff_A_FVMnuiyI7_0),.clk(gclk));
	jdff dff_A_OKMn6FoW1_0(.dout(w_dff_A_FVMnuiyI7_0),.din(w_dff_A_OKMn6FoW1_0),.clk(gclk));
	jdff dff_A_TpvHyZ6w5_0(.dout(w_dff_A_OKMn6FoW1_0),.din(w_dff_A_TpvHyZ6w5_0),.clk(gclk));
	jdff dff_A_hujdfCwR5_0(.dout(w_dff_A_TpvHyZ6w5_0),.din(w_dff_A_hujdfCwR5_0),.clk(gclk));
	jdff dff_A_3vP2MEBK1_0(.dout(w_dff_A_hujdfCwR5_0),.din(w_dff_A_3vP2MEBK1_0),.clk(gclk));
	jdff dff_A_ZZbiFHxe9_0(.dout(w_dff_A_3vP2MEBK1_0),.din(w_dff_A_ZZbiFHxe9_0),.clk(gclk));
	jdff dff_A_20UkTApF4_0(.dout(w_dff_A_ZZbiFHxe9_0),.din(w_dff_A_20UkTApF4_0),.clk(gclk));
	jdff dff_A_QkA2Cbpy2_0(.dout(w_dff_A_20UkTApF4_0),.din(w_dff_A_QkA2Cbpy2_0),.clk(gclk));
	jdff dff_A_M9pP9sKD7_0(.dout(w_dff_A_QkA2Cbpy2_0),.din(w_dff_A_M9pP9sKD7_0),.clk(gclk));
	jdff dff_A_fNheglJ38_0(.dout(w_dff_A_M9pP9sKD7_0),.din(w_dff_A_fNheglJ38_0),.clk(gclk));
	jdff dff_A_1MLnXUWn3_0(.dout(w_dff_A_fNheglJ38_0),.din(w_dff_A_1MLnXUWn3_0),.clk(gclk));
	jdff dff_A_FtZ0zyZN3_0(.dout(w_dff_A_1MLnXUWn3_0),.din(w_dff_A_FtZ0zyZN3_0),.clk(gclk));
	jdff dff_A_5dlSNhTG7_0(.dout(w_dff_A_FtZ0zyZN3_0),.din(w_dff_A_5dlSNhTG7_0),.clk(gclk));
	jdff dff_A_S0eMVCQg5_0(.dout(w_dff_A_5dlSNhTG7_0),.din(w_dff_A_S0eMVCQg5_0),.clk(gclk));
	jdff dff_A_kPIoaThd5_0(.dout(w_dff_A_S0eMVCQg5_0),.din(w_dff_A_kPIoaThd5_0),.clk(gclk));
	jdff dff_A_E4SvCZKX6_0(.dout(w_dff_A_kPIoaThd5_0),.din(w_dff_A_E4SvCZKX6_0),.clk(gclk));
	jdff dff_A_IL5ZPbh26_0(.dout(w_dff_A_E4SvCZKX6_0),.din(w_dff_A_IL5ZPbh26_0),.clk(gclk));
	jdff dff_A_55F6uHpY0_0(.dout(w_G53gat_0[0]),.din(w_dff_A_55F6uHpY0_0),.clk(gclk));
	jdff dff_A_mmTeX8682_0(.dout(w_dff_A_55F6uHpY0_0),.din(w_dff_A_mmTeX8682_0),.clk(gclk));
	jdff dff_A_5yGrNJrr8_0(.dout(w_dff_A_mmTeX8682_0),.din(w_dff_A_5yGrNJrr8_0),.clk(gclk));
	jdff dff_A_Yaq6pThX1_0(.dout(w_dff_A_5yGrNJrr8_0),.din(w_dff_A_Yaq6pThX1_0),.clk(gclk));
	jdff dff_A_j0pUy80B5_0(.dout(w_dff_A_Yaq6pThX1_0),.din(w_dff_A_j0pUy80B5_0),.clk(gclk));
	jdff dff_A_yaHGqrTN8_0(.dout(w_dff_A_j0pUy80B5_0),.din(w_dff_A_yaHGqrTN8_0),.clk(gclk));
	jdff dff_A_tsRvy61C7_0(.dout(w_dff_A_yaHGqrTN8_0),.din(w_dff_A_tsRvy61C7_0),.clk(gclk));
	jdff dff_A_xGJQImtM9_0(.dout(w_dff_A_tsRvy61C7_0),.din(w_dff_A_xGJQImtM9_0),.clk(gclk));
	jdff dff_A_sNgvTVzH1_0(.dout(w_dff_A_xGJQImtM9_0),.din(w_dff_A_sNgvTVzH1_0),.clk(gclk));
	jdff dff_A_mw0Elirt8_0(.dout(w_dff_A_sNgvTVzH1_0),.din(w_dff_A_mw0Elirt8_0),.clk(gclk));
	jdff dff_A_3NOVNtP00_0(.dout(w_dff_A_mw0Elirt8_0),.din(w_dff_A_3NOVNtP00_0),.clk(gclk));
	jdff dff_A_hxBmxHZL4_0(.dout(w_dff_A_3NOVNtP00_0),.din(w_dff_A_hxBmxHZL4_0),.clk(gclk));
	jdff dff_A_XeTWTHoh5_0(.dout(w_dff_A_hxBmxHZL4_0),.din(w_dff_A_XeTWTHoh5_0),.clk(gclk));
	jdff dff_A_yaRqaiCT1_0(.dout(w_dff_A_XeTWTHoh5_0),.din(w_dff_A_yaRqaiCT1_0),.clk(gclk));
	jdff dff_A_JoSfo5vs7_0(.dout(w_dff_A_yaRqaiCT1_0),.din(w_dff_A_JoSfo5vs7_0),.clk(gclk));
	jdff dff_A_EAw1ZGuB9_0(.dout(w_dff_A_JoSfo5vs7_0),.din(w_dff_A_EAw1ZGuB9_0),.clk(gclk));
	jdff dff_A_tJmv72Z84_0(.dout(w_dff_A_EAw1ZGuB9_0),.din(w_dff_A_tJmv72Z84_0),.clk(gclk));
	jdff dff_A_8EFlvp4J9_0(.dout(w_dff_A_tJmv72Z84_0),.din(w_dff_A_8EFlvp4J9_0),.clk(gclk));
	jdff dff_A_RSoaLTfG0_0(.dout(w_dff_A_8EFlvp4J9_0),.din(w_dff_A_RSoaLTfG0_0),.clk(gclk));
	jdff dff_A_i8Zztezs4_0(.dout(w_dff_A_RSoaLTfG0_0),.din(w_dff_A_i8Zztezs4_0),.clk(gclk));
	jdff dff_A_Nb4pAod21_0(.dout(w_n184_0[0]),.din(w_dff_A_Nb4pAod21_0),.clk(gclk));
	jdff dff_A_Myvlt2t65_0(.dout(w_dff_A_Nb4pAod21_0),.din(w_dff_A_Myvlt2t65_0),.clk(gclk));
	jdff dff_A_Vi320bna1_0(.dout(w_dff_A_Myvlt2t65_0),.din(w_dff_A_Vi320bna1_0),.clk(gclk));
	jdff dff_A_zwrhq5XR9_0(.dout(w_dff_A_Vi320bna1_0),.din(w_dff_A_zwrhq5XR9_0),.clk(gclk));
	jdff dff_A_ghXPkxnc5_0(.dout(w_dff_A_zwrhq5XR9_0),.din(w_dff_A_ghXPkxnc5_0),.clk(gclk));
	jdff dff_A_SI3AbHif1_0(.dout(w_dff_A_ghXPkxnc5_0),.din(w_dff_A_SI3AbHif1_0),.clk(gclk));
	jdff dff_B_YUN2JMjJ6_1(.din(n167),.dout(w_dff_B_YUN2JMjJ6_1),.clk(gclk));
	jdff dff_A_BJHSwyQx8_0(.dout(w_n177_0[0]),.din(w_dff_A_BJHSwyQx8_0),.clk(gclk));
	jdff dff_A_tzT4W7pv5_0(.dout(w_dff_A_BJHSwyQx8_0),.din(w_dff_A_tzT4W7pv5_0),.clk(gclk));
	jdff dff_A_KpLEh9Nu4_0(.dout(w_dff_A_tzT4W7pv5_0),.din(w_dff_A_KpLEh9Nu4_0),.clk(gclk));
	jdff dff_A_g2C6mCoA6_0(.dout(w_dff_A_KpLEh9Nu4_0),.din(w_dff_A_g2C6mCoA6_0),.clk(gclk));
	jdff dff_A_K6YDEDBB2_0(.dout(w_dff_A_g2C6mCoA6_0),.din(w_dff_A_K6YDEDBB2_0),.clk(gclk));
	jdff dff_A_CLTiIAIk1_0(.dout(w_dff_A_K6YDEDBB2_0),.din(w_dff_A_CLTiIAIk1_0),.clk(gclk));
	jdff dff_A_FZjuf3g77_0(.dout(w_n174_0[0]),.din(w_dff_A_FZjuf3g77_0),.clk(gclk));
	jdff dff_A_2vwPjiJL8_0(.dout(w_dff_A_FZjuf3g77_0),.din(w_dff_A_2vwPjiJL8_0),.clk(gclk));
	jdff dff_A_0vRLJBEb8_0(.dout(w_dff_A_2vwPjiJL8_0),.din(w_dff_A_0vRLJBEb8_0),.clk(gclk));
	jdff dff_A_AleaHKx53_0(.dout(w_dff_A_0vRLJBEb8_0),.din(w_dff_A_AleaHKx53_0),.clk(gclk));
	jdff dff_A_owB79coh6_0(.dout(w_dff_A_AleaHKx53_0),.din(w_dff_A_owB79coh6_0),.clk(gclk));
	jdff dff_A_KrOIrhnz6_0(.dout(w_dff_A_owB79coh6_0),.din(w_dff_A_KrOIrhnz6_0),.clk(gclk));
	jdff dff_B_PhXamBYL5_1(.din(n172),.dout(w_dff_B_PhXamBYL5_1),.clk(gclk));
	jdff dff_B_pTSn0IBv6_1(.din(w_dff_B_PhXamBYL5_1),.dout(w_dff_B_pTSn0IBv6_1),.clk(gclk));
	jdff dff_B_ALspOavY2_1(.din(w_dff_B_pTSn0IBv6_1),.dout(w_dff_B_ALspOavY2_1),.clk(gclk));
	jdff dff_B_3m7qSE6r0_1(.din(w_dff_B_ALspOavY2_1),.dout(w_dff_B_3m7qSE6r0_1),.clk(gclk));
	jdff dff_B_cCWLRHyF8_1(.din(w_dff_B_3m7qSE6r0_1),.dout(w_dff_B_cCWLRHyF8_1),.clk(gclk));
	jdff dff_B_U5uq0R0n0_1(.din(w_dff_B_cCWLRHyF8_1),.dout(w_dff_B_U5uq0R0n0_1),.clk(gclk));
	jdff dff_A_4ZHIWnzA2_0(.dout(w_n170_0[0]),.din(w_dff_A_4ZHIWnzA2_0),.clk(gclk));
	jdff dff_A_9EIJR6911_0(.dout(w_dff_A_4ZHIWnzA2_0),.din(w_dff_A_9EIJR6911_0),.clk(gclk));
	jdff dff_A_3NZ7AJHN7_0(.dout(w_dff_A_9EIJR6911_0),.din(w_dff_A_3NZ7AJHN7_0),.clk(gclk));
	jdff dff_A_f8IuNFel1_0(.dout(w_dff_A_3NZ7AJHN7_0),.din(w_dff_A_f8IuNFel1_0),.clk(gclk));
	jdff dff_B_AkYWyoNi7_2(.din(n170),.dout(w_dff_B_AkYWyoNi7_2),.clk(gclk));
	jdff dff_B_N2hdPM6Q1_0(.din(n169),.dout(w_dff_B_N2hdPM6Q1_0),.clk(gclk));
	jdff dff_B_k0oKSxZz6_0(.din(w_dff_B_N2hdPM6Q1_0),.dout(w_dff_B_k0oKSxZz6_0),.clk(gclk));
	jdff dff_B_6Ya57KKM4_0(.din(w_dff_B_k0oKSxZz6_0),.dout(w_dff_B_6Ya57KKM4_0),.clk(gclk));
	jdff dff_B_J5sydVXs4_0(.din(w_dff_B_6Ya57KKM4_0),.dout(w_dff_B_J5sydVXs4_0),.clk(gclk));
	jdff dff_A_dXqkiOAU8_0(.dout(w_n164_0[0]),.din(w_dff_A_dXqkiOAU8_0),.clk(gclk));
	jdff dff_A_pAt8pkO59_0(.dout(w_dff_A_dXqkiOAU8_0),.din(w_dff_A_pAt8pkO59_0),.clk(gclk));
	jdff dff_A_hdoSAK8G1_0(.dout(w_dff_A_pAt8pkO59_0),.din(w_dff_A_hdoSAK8G1_0),.clk(gclk));
	jdff dff_A_VRgXca2F3_0(.dout(w_dff_A_hdoSAK8G1_0),.din(w_dff_A_VRgXca2F3_0),.clk(gclk));
	jdff dff_A_xYBILegS7_0(.dout(w_dff_A_VRgXca2F3_0),.din(w_dff_A_xYBILegS7_0),.clk(gclk));
	jdff dff_A_BB2erPz25_0(.dout(w_dff_A_xYBILegS7_0),.din(w_dff_A_BB2erPz25_0),.clk(gclk));
	jdff dff_A_9aOj0izt2_0(.dout(w_n159_0[0]),.din(w_dff_A_9aOj0izt2_0),.clk(gclk));
	jdff dff_A_SKkCYDpZ5_0(.dout(w_dff_A_9aOj0izt2_0),.din(w_dff_A_SKkCYDpZ5_0),.clk(gclk));
	jdff dff_A_cvorLVXz3_0(.dout(w_dff_A_SKkCYDpZ5_0),.din(w_dff_A_cvorLVXz3_0),.clk(gclk));
	jdff dff_A_tpRIXYBS3_0(.dout(w_dff_A_cvorLVXz3_0),.din(w_dff_A_tpRIXYBS3_0),.clk(gclk));
	jdff dff_A_NCLTK07C8_0(.dout(w_dff_A_tpRIXYBS3_0),.din(w_dff_A_NCLTK07C8_0),.clk(gclk));
	jdff dff_A_1LY0ds4S1_0(.dout(w_dff_A_NCLTK07C8_0),.din(w_dff_A_1LY0ds4S1_0),.clk(gclk));
	jdff dff_A_BbvkIzyJ6_0(.dout(w_n156_0[0]),.din(w_dff_A_BbvkIzyJ6_0),.clk(gclk));
	jdff dff_A_Thzz6PHF7_0(.dout(w_dff_A_BbvkIzyJ6_0),.din(w_dff_A_Thzz6PHF7_0),.clk(gclk));
	jdff dff_A_znumnVVH6_0(.dout(w_dff_A_Thzz6PHF7_0),.din(w_dff_A_znumnVVH6_0),.clk(gclk));
	jdff dff_A_hgmNFIf31_0(.dout(w_dff_A_znumnVVH6_0),.din(w_dff_A_hgmNFIf31_0),.clk(gclk));
	jdff dff_A_77ukaDLg7_0(.dout(w_dff_A_hgmNFIf31_0),.din(w_dff_A_77ukaDLg7_0),.clk(gclk));
	jdff dff_A_femGqmDM7_0(.dout(w_dff_A_77ukaDLg7_0),.din(w_dff_A_femGqmDM7_0),.clk(gclk));
	jdff dff_A_U3sk8za80_0(.dout(w_n154_0[0]),.din(w_dff_A_U3sk8za80_0),.clk(gclk));
	jdff dff_A_DAbPBAop5_0(.dout(w_dff_A_U3sk8za80_0),.din(w_dff_A_DAbPBAop5_0),.clk(gclk));
	jdff dff_A_gDMg3dVH5_0(.dout(w_dff_A_DAbPBAop5_0),.din(w_dff_A_gDMg3dVH5_0),.clk(gclk));
	jdff dff_A_bHqQwJqX2_0(.dout(w_dff_A_gDMg3dVH5_0),.din(w_dff_A_bHqQwJqX2_0),.clk(gclk));
	jdff dff_A_Rx2Dkhn52_0(.dout(w_dff_A_bHqQwJqX2_0),.din(w_dff_A_Rx2Dkhn52_0),.clk(gclk));
	jdff dff_B_pdLOxC067_2(.din(n154),.dout(w_dff_B_pdLOxC067_2),.clk(gclk));
	jdff dff_B_hWWK1P840_2(.din(w_dff_B_pdLOxC067_2),.dout(w_dff_B_hWWK1P840_2),.clk(gclk));
	jdff dff_B_0s5a6xyR5_2(.din(w_dff_B_hWWK1P840_2),.dout(w_dff_B_0s5a6xyR5_2),.clk(gclk));
	jdff dff_B_kGkSn32F0_2(.din(w_dff_B_0s5a6xyR5_2),.dout(w_dff_B_kGkSn32F0_2),.clk(gclk));
	jdff dff_B_C1fnISYO9_2(.din(w_dff_B_kGkSn32F0_2),.dout(w_dff_B_C1fnISYO9_2),.clk(gclk));
	jdff dff_B_OyKpGCGx9_2(.din(w_dff_B_C1fnISYO9_2),.dout(w_dff_B_OyKpGCGx9_2),.clk(gclk));
	jdff dff_B_IDlmOMsx9_2(.din(w_dff_B_OyKpGCGx9_2),.dout(w_dff_B_IDlmOMsx9_2),.clk(gclk));
	jdff dff_B_UJP0Ddyk4_2(.din(w_dff_B_IDlmOMsx9_2),.dout(w_dff_B_UJP0Ddyk4_2),.clk(gclk));
	jdff dff_B_y3wFeHkE4_2(.din(w_dff_B_UJP0Ddyk4_2),.dout(w_dff_B_y3wFeHkE4_2),.clk(gclk));
	jdff dff_B_kX6bMGpm6_2(.din(w_dff_B_y3wFeHkE4_2),.dout(w_dff_B_kX6bMGpm6_2),.clk(gclk));
	jdff dff_B_dBcBY3pX1_2(.din(w_dff_B_kX6bMGpm6_2),.dout(w_dff_B_dBcBY3pX1_2),.clk(gclk));
	jdff dff_B_tD1JO75M7_2(.din(w_dff_B_dBcBY3pX1_2),.dout(w_dff_B_tD1JO75M7_2),.clk(gclk));
	jdff dff_B_R0nRX52Z0_2(.din(w_dff_B_tD1JO75M7_2),.dout(w_dff_B_R0nRX52Z0_2),.clk(gclk));
	jdff dff_B_ptDOWvoi1_2(.din(w_dff_B_R0nRX52Z0_2),.dout(w_dff_B_ptDOWvoi1_2),.clk(gclk));
	jdff dff_A_lHI0qlei8_0(.dout(w_G79gat_0[0]),.din(w_dff_A_lHI0qlei8_0),.clk(gclk));
	jdff dff_A_u8LNLsDM7_0(.dout(w_dff_A_lHI0qlei8_0),.din(w_dff_A_u8LNLsDM7_0),.clk(gclk));
	jdff dff_A_TrDj6usd7_0(.dout(w_dff_A_u8LNLsDM7_0),.din(w_dff_A_TrDj6usd7_0),.clk(gclk));
	jdff dff_A_o3heIQwe7_0(.dout(w_dff_A_TrDj6usd7_0),.din(w_dff_A_o3heIQwe7_0),.clk(gclk));
	jdff dff_A_1DiCN2SE6_0(.dout(w_dff_A_o3heIQwe7_0),.din(w_dff_A_1DiCN2SE6_0),.clk(gclk));
	jdff dff_A_IZWfG0Lt4_0(.dout(w_dff_A_1DiCN2SE6_0),.din(w_dff_A_IZWfG0Lt4_0),.clk(gclk));
	jdff dff_A_GMWXHIOT4_0(.dout(w_dff_A_IZWfG0Lt4_0),.din(w_dff_A_GMWXHIOT4_0),.clk(gclk));
	jdff dff_A_JG7gYZDR4_0(.dout(w_dff_A_GMWXHIOT4_0),.din(w_dff_A_JG7gYZDR4_0),.clk(gclk));
	jdff dff_A_KBsHaoqG0_0(.dout(w_dff_A_JG7gYZDR4_0),.din(w_dff_A_KBsHaoqG0_0),.clk(gclk));
	jdff dff_A_O6t7W3kg8_0(.dout(w_dff_A_KBsHaoqG0_0),.din(w_dff_A_O6t7W3kg8_0),.clk(gclk));
	jdff dff_A_YDw0EU7O7_0(.dout(w_dff_A_O6t7W3kg8_0),.din(w_dff_A_YDw0EU7O7_0),.clk(gclk));
	jdff dff_A_lcXDKDi94_0(.dout(w_dff_A_YDw0EU7O7_0),.din(w_dff_A_lcXDKDi94_0),.clk(gclk));
	jdff dff_A_WmywqqHu6_0(.dout(w_dff_A_lcXDKDi94_0),.din(w_dff_A_WmywqqHu6_0),.clk(gclk));
	jdff dff_A_pbkj0S0E2_0(.dout(w_dff_A_WmywqqHu6_0),.din(w_dff_A_pbkj0S0E2_0),.clk(gclk));
	jdff dff_A_qE4HPvK16_0(.dout(w_dff_A_pbkj0S0E2_0),.din(w_dff_A_qE4HPvK16_0),.clk(gclk));
	jdff dff_A_pzLyM3gx7_1(.dout(w_n151_0[1]),.din(w_dff_A_pzLyM3gx7_1),.clk(gclk));
	jdff dff_A_zBABjna93_1(.dout(w_dff_A_pzLyM3gx7_1),.din(w_dff_A_zBABjna93_1),.clk(gclk));
	jdff dff_A_MsasnzLU9_1(.dout(w_dff_A_zBABjna93_1),.din(w_dff_A_MsasnzLU9_1),.clk(gclk));
	jdff dff_A_cP8VsnHO1_1(.dout(w_dff_A_MsasnzLU9_1),.din(w_dff_A_cP8VsnHO1_1),.clk(gclk));
	jdff dff_A_JeaOdzIB6_1(.dout(w_dff_A_cP8VsnHO1_1),.din(w_dff_A_JeaOdzIB6_1),.clk(gclk));
	jdff dff_A_JNGfH7qg4_1(.dout(w_dff_A_JeaOdzIB6_1),.din(w_dff_A_JNGfH7qg4_1),.clk(gclk));
	jdff dff_A_BrRnh4N75_0(.dout(w_n150_0[0]),.din(w_dff_A_BrRnh4N75_0),.clk(gclk));
	jdff dff_A_nOrIbI2l9_0(.dout(w_dff_A_BrRnh4N75_0),.din(w_dff_A_nOrIbI2l9_0),.clk(gclk));
	jdff dff_A_AdX6YHTy3_0(.dout(w_dff_A_nOrIbI2l9_0),.din(w_dff_A_AdX6YHTy3_0),.clk(gclk));
	jdff dff_A_RSASyS4r5_0(.dout(w_dff_A_AdX6YHTy3_0),.din(w_dff_A_RSASyS4r5_0),.clk(gclk));
	jdff dff_A_miWn5h5e1_0(.dout(w_dff_A_RSASyS4r5_0),.din(w_dff_A_miWn5h5e1_0),.clk(gclk));
	jdff dff_A_8ZQC5ilP0_0(.dout(w_dff_A_miWn5h5e1_0),.din(w_dff_A_8ZQC5ilP0_0),.clk(gclk));
	jdff dff_A_xtnGSsQG6_0(.dout(w_dff_A_8ZQC5ilP0_0),.din(w_dff_A_xtnGSsQG6_0),.clk(gclk));
	jdff dff_A_FysE8gZR8_0(.dout(w_dff_A_xtnGSsQG6_0),.din(w_dff_A_FysE8gZR8_0),.clk(gclk));
	jdff dff_A_MOoBy9eR6_0(.dout(w_dff_A_FysE8gZR8_0),.din(w_dff_A_MOoBy9eR6_0),.clk(gclk));
	jdff dff_A_HCy3xjCo5_0(.dout(w_dff_A_MOoBy9eR6_0),.din(w_dff_A_HCy3xjCo5_0),.clk(gclk));
	jdff dff_A_Zy3wGKlo0_0(.dout(w_dff_A_HCy3xjCo5_0),.din(w_dff_A_Zy3wGKlo0_0),.clk(gclk));
	jdff dff_A_vBJ43En75_0(.dout(w_dff_A_Zy3wGKlo0_0),.din(w_dff_A_vBJ43En75_0),.clk(gclk));
	jdff dff_B_e3BDnmtq8_2(.din(n150),.dout(w_dff_B_e3BDnmtq8_2),.clk(gclk));
	jdff dff_B_d2JeyH4E2_2(.din(w_dff_B_e3BDnmtq8_2),.dout(w_dff_B_d2JeyH4E2_2),.clk(gclk));
	jdff dff_B_UbCuBvmm9_2(.din(w_dff_B_d2JeyH4E2_2),.dout(w_dff_B_UbCuBvmm9_2),.clk(gclk));
	jdff dff_B_hQwbeBWj0_2(.din(w_dff_B_UbCuBvmm9_2),.dout(w_dff_B_hQwbeBWj0_2),.clk(gclk));
	jdff dff_B_5hU28amv6_2(.din(w_dff_B_hQwbeBWj0_2),.dout(w_dff_B_5hU28amv6_2),.clk(gclk));
	jdff dff_B_5VaHrKr32_2(.din(w_dff_B_5hU28amv6_2),.dout(w_dff_B_5VaHrKr32_2),.clk(gclk));
	jdff dff_B_GAX9VgP40_2(.din(w_dff_B_5VaHrKr32_2),.dout(w_dff_B_GAX9VgP40_2),.clk(gclk));
	jdff dff_A_bBUItHpo9_0(.dout(w_G66gat_0[0]),.din(w_dff_A_bBUItHpo9_0),.clk(gclk));
	jdff dff_A_N49Y5pdL3_0(.dout(w_dff_A_bBUItHpo9_0),.din(w_dff_A_N49Y5pdL3_0),.clk(gclk));
	jdff dff_A_WKna2wMk9_0(.dout(w_dff_A_N49Y5pdL3_0),.din(w_dff_A_WKna2wMk9_0),.clk(gclk));
	jdff dff_A_qgkIiCyx0_0(.dout(w_dff_A_WKna2wMk9_0),.din(w_dff_A_qgkIiCyx0_0),.clk(gclk));
	jdff dff_A_TFxqJ3Iw1_0(.dout(w_dff_A_qgkIiCyx0_0),.din(w_dff_A_TFxqJ3Iw1_0),.clk(gclk));
	jdff dff_A_N4fYCRD64_0(.dout(w_dff_A_TFxqJ3Iw1_0),.din(w_dff_A_N4fYCRD64_0),.clk(gclk));
	jdff dff_A_8RG6u1X27_0(.dout(w_dff_A_N4fYCRD64_0),.din(w_dff_A_8RG6u1X27_0),.clk(gclk));
	jdff dff_A_wa1cESpL0_0(.dout(w_dff_A_8RG6u1X27_0),.din(w_dff_A_wa1cESpL0_0),.clk(gclk));
	jdff dff_A_bNP1P9KA6_0(.dout(w_dff_A_wa1cESpL0_0),.din(w_dff_A_bNP1P9KA6_0),.clk(gclk));
	jdff dff_A_phYwgwFP5_0(.dout(w_dff_A_bNP1P9KA6_0),.din(w_dff_A_phYwgwFP5_0),.clk(gclk));
	jdff dff_A_WPuFpHnU9_0(.dout(w_dff_A_phYwgwFP5_0),.din(w_dff_A_WPuFpHnU9_0),.clk(gclk));
	jdff dff_A_Uz8owtnF2_0(.dout(w_dff_A_WPuFpHnU9_0),.din(w_dff_A_Uz8owtnF2_0),.clk(gclk));
	jdff dff_A_8hZSAhgg7_0(.dout(w_dff_A_Uz8owtnF2_0),.din(w_dff_A_8hZSAhgg7_0),.clk(gclk));
	jdff dff_A_7NOKzKGz5_0(.dout(w_dff_A_8hZSAhgg7_0),.din(w_dff_A_7NOKzKGz5_0),.clk(gclk));
	jdff dff_A_aNRS81IT1_0(.dout(w_dff_A_7NOKzKGz5_0),.din(w_dff_A_aNRS81IT1_0),.clk(gclk));
	jdff dff_A_bvacKOWW7_0(.dout(w_dff_A_aNRS81IT1_0),.din(w_dff_A_bvacKOWW7_0),.clk(gclk));
	jdff dff_A_Xf476TJt8_0(.dout(w_dff_A_bvacKOWW7_0),.din(w_dff_A_Xf476TJt8_0),.clk(gclk));
	jdff dff_A_3lvclMmW7_0(.dout(w_dff_A_Xf476TJt8_0),.din(w_dff_A_3lvclMmW7_0),.clk(gclk));
	jdff dff_A_nKJbfG0F3_0(.dout(w_dff_A_3lvclMmW7_0),.din(w_dff_A_nKJbfG0F3_0),.clk(gclk));
	jdff dff_A_2DolGJBw8_0(.dout(w_dff_A_nKJbfG0F3_0),.din(w_dff_A_2DolGJBw8_0),.clk(gclk));
	jdff dff_A_slBXbMmL5_1(.dout(w_n146_0[1]),.din(w_dff_A_slBXbMmL5_1),.clk(gclk));
	jdff dff_A_JDwlrsJB1_1(.dout(w_dff_A_slBXbMmL5_1),.din(w_dff_A_JDwlrsJB1_1),.clk(gclk));
	jdff dff_A_vPCPcutH4_1(.dout(w_dff_A_JDwlrsJB1_1),.din(w_dff_A_vPCPcutH4_1),.clk(gclk));
	jdff dff_A_B6fkMwmI7_1(.dout(w_dff_A_vPCPcutH4_1),.din(w_dff_A_B6fkMwmI7_1),.clk(gclk));
	jdff dff_A_0NKTxPqa0_0(.dout(w_n145_0[0]),.din(w_dff_A_0NKTxPqa0_0),.clk(gclk));
	jdff dff_A_aDoKFDYl3_0(.dout(w_dff_A_0NKTxPqa0_0),.din(w_dff_A_aDoKFDYl3_0),.clk(gclk));
	jdff dff_A_S9rIC2Lj5_0(.dout(w_dff_A_aDoKFDYl3_0),.din(w_dff_A_S9rIC2Lj5_0),.clk(gclk));
	jdff dff_A_l6mBzRnm6_0(.dout(w_dff_A_S9rIC2Lj5_0),.din(w_dff_A_l6mBzRnm6_0),.clk(gclk));
	jdff dff_A_DcnG9xyW5_0(.dout(w_dff_A_l6mBzRnm6_0),.din(w_dff_A_DcnG9xyW5_0),.clk(gclk));
	jdff dff_A_bgm1NLjI3_0(.dout(w_dff_A_DcnG9xyW5_0),.din(w_dff_A_bgm1NLjI3_0),.clk(gclk));
	jdff dff_A_EPfnWR8I7_0(.dout(w_n142_0[0]),.din(w_dff_A_EPfnWR8I7_0),.clk(gclk));
	jdff dff_B_FO7OnCup9_1(.din(n112),.dout(w_dff_B_FO7OnCup9_1),.clk(gclk));
	jdff dff_B_W4NMkniy8_1(.din(n116),.dout(w_dff_B_W4NMkniy8_1),.clk(gclk));
	jdff dff_A_4kiezU4t7_0(.dout(w_n132_0[0]),.din(w_dff_A_4kiezU4t7_0),.clk(gclk));
	jdff dff_A_JjNGq4TP7_0(.dout(w_dff_A_4kiezU4t7_0),.din(w_dff_A_JjNGq4TP7_0),.clk(gclk));
	jdff dff_A_Y0ChjMwC4_0(.dout(w_dff_A_JjNGq4TP7_0),.din(w_dff_A_Y0ChjMwC4_0),.clk(gclk));
	jdff dff_A_rsos5Fm00_0(.dout(w_dff_A_Y0ChjMwC4_0),.din(w_dff_A_rsos5Fm00_0),.clk(gclk));
	jdff dff_A_zrmGGB885_0(.dout(w_dff_A_rsos5Fm00_0),.din(w_dff_A_zrmGGB885_0),.clk(gclk));
	jdff dff_A_L7UkzfMe6_0(.dout(w_dff_A_zrmGGB885_0),.din(w_dff_A_L7UkzfMe6_0),.clk(gclk));
	jdff dff_A_qOfXCRrd5_0(.dout(w_n130_0[0]),.din(w_dff_A_qOfXCRrd5_0),.clk(gclk));
	jdff dff_A_tAC1vEVq3_0(.dout(w_dff_A_qOfXCRrd5_0),.din(w_dff_A_tAC1vEVq3_0),.clk(gclk));
	jdff dff_A_Q7enk1ph6_0(.dout(w_dff_A_tAC1vEVq3_0),.din(w_dff_A_Q7enk1ph6_0),.clk(gclk));
	jdff dff_A_ORMBbBKv0_0(.dout(w_dff_A_Q7enk1ph6_0),.din(w_dff_A_ORMBbBKv0_0),.clk(gclk));
	jdff dff_A_JeYl2SgM1_0(.dout(w_dff_A_ORMBbBKv0_0),.din(w_dff_A_JeYl2SgM1_0),.clk(gclk));
	jdff dff_A_Yds801NX3_1(.dout(w_n130_0[1]),.din(w_dff_A_Yds801NX3_1),.clk(gclk));
	jdff dff_A_wC0HanK92_1(.dout(w_dff_A_Yds801NX3_1),.din(w_dff_A_wC0HanK92_1),.clk(gclk));
	jdff dff_A_7o98vxHV9_1(.dout(w_dff_A_wC0HanK92_1),.din(w_dff_A_7o98vxHV9_1),.clk(gclk));
	jdff dff_A_XMDxYmPO5_1(.dout(w_dff_A_7o98vxHV9_1),.din(w_dff_A_XMDxYmPO5_1),.clk(gclk));
	jdff dff_A_tO3P15gs0_1(.dout(w_dff_A_XMDxYmPO5_1),.din(w_dff_A_tO3P15gs0_1),.clk(gclk));
	jdff dff_B_etPOqWoX6_3(.din(n130),.dout(w_dff_B_etPOqWoX6_3),.clk(gclk));
	jdff dff_B_zcnCxPAJ4_3(.din(w_dff_B_etPOqWoX6_3),.dout(w_dff_B_zcnCxPAJ4_3),.clk(gclk));
	jdff dff_B_nzUlwps71_3(.din(w_dff_B_zcnCxPAJ4_3),.dout(w_dff_B_nzUlwps71_3),.clk(gclk));
	jdff dff_B_a4rYuHcC1_3(.din(w_dff_B_nzUlwps71_3),.dout(w_dff_B_a4rYuHcC1_3),.clk(gclk));
	jdff dff_B_7l1AWG7J3_3(.din(w_dff_B_a4rYuHcC1_3),.dout(w_dff_B_7l1AWG7J3_3),.clk(gclk));
	jdff dff_B_aKs3vIiu9_3(.din(w_dff_B_7l1AWG7J3_3),.dout(w_dff_B_aKs3vIiu9_3),.clk(gclk));
	jdff dff_B_EzKS0AVu8_3(.din(w_dff_B_aKs3vIiu9_3),.dout(w_dff_B_EzKS0AVu8_3),.clk(gclk));
	jdff dff_A_mcgw9Ud00_0(.dout(w_G21gat_1[0]),.din(w_dff_A_mcgw9Ud00_0),.clk(gclk));
	jdff dff_A_VIkFKt1a2_0(.dout(w_dff_A_mcgw9Ud00_0),.din(w_dff_A_VIkFKt1a2_0),.clk(gclk));
	jdff dff_A_8NeDOyXR5_0(.dout(w_dff_A_VIkFKt1a2_0),.din(w_dff_A_8NeDOyXR5_0),.clk(gclk));
	jdff dff_A_xetB8bEd4_0(.dout(w_dff_A_8NeDOyXR5_0),.din(w_dff_A_xetB8bEd4_0),.clk(gclk));
	jdff dff_A_SpFOPOTi6_0(.dout(w_dff_A_xetB8bEd4_0),.din(w_dff_A_SpFOPOTi6_0),.clk(gclk));
	jdff dff_A_2WIHBanQ2_0(.dout(w_dff_A_SpFOPOTi6_0),.din(w_dff_A_2WIHBanQ2_0),.clk(gclk));
	jdff dff_A_cwD07wTi9_0(.dout(w_dff_A_2WIHBanQ2_0),.din(w_dff_A_cwD07wTi9_0),.clk(gclk));
	jdff dff_A_oiRTHhbG8_0(.dout(w_dff_A_cwD07wTi9_0),.din(w_dff_A_oiRTHhbG8_0),.clk(gclk));
	jdff dff_A_UZM8Wk3A5_1(.dout(w_G21gat_0[1]),.din(w_dff_A_UZM8Wk3A5_1),.clk(gclk));
	jdff dff_A_1vWXWuOn0_1(.dout(w_dff_A_UZM8Wk3A5_1),.din(w_dff_A_1vWXWuOn0_1),.clk(gclk));
	jdff dff_A_2fjhSJ0N7_1(.dout(w_dff_A_1vWXWuOn0_1),.din(w_dff_A_2fjhSJ0N7_1),.clk(gclk));
	jdff dff_A_oRrvzPiG2_1(.dout(w_dff_A_2fjhSJ0N7_1),.din(w_dff_A_oRrvzPiG2_1),.clk(gclk));
	jdff dff_A_HCmVVddG2_1(.dout(w_dff_A_oRrvzPiG2_1),.din(w_dff_A_HCmVVddG2_1),.clk(gclk));
	jdff dff_A_Qc06GbXM9_1(.dout(w_dff_A_HCmVVddG2_1),.din(w_dff_A_Qc06GbXM9_1),.clk(gclk));
	jdff dff_A_kKhWHCdr7_1(.dout(w_dff_A_Qc06GbXM9_1),.din(w_dff_A_kKhWHCdr7_1),.clk(gclk));
	jdff dff_A_y96emqx31_1(.dout(w_dff_A_kKhWHCdr7_1),.din(w_dff_A_y96emqx31_1),.clk(gclk));
	jdff dff_A_AW856LJC9_1(.dout(w_dff_A_y96emqx31_1),.din(w_dff_A_AW856LJC9_1),.clk(gclk));
	jdff dff_A_kWw48Eko2_1(.dout(w_dff_A_AW856LJC9_1),.din(w_dff_A_kWw48Eko2_1),.clk(gclk));
	jdff dff_A_DTf9QwgS4_1(.dout(w_dff_A_kWw48Eko2_1),.din(w_dff_A_DTf9QwgS4_1),.clk(gclk));
	jdff dff_A_B894nJWu0_1(.dout(w_dff_A_DTf9QwgS4_1),.din(w_dff_A_B894nJWu0_1),.clk(gclk));
	jdff dff_A_PtjufDcc3_1(.dout(w_dff_A_B894nJWu0_1),.din(w_dff_A_PtjufDcc3_1),.clk(gclk));
	jdff dff_A_ATVsHW0w7_2(.dout(w_G21gat_0[2]),.din(w_dff_A_ATVsHW0w7_2),.clk(gclk));
	jdff dff_A_hypxtFVw3_2(.dout(w_dff_A_ATVsHW0w7_2),.din(w_dff_A_hypxtFVw3_2),.clk(gclk));
	jdff dff_A_2ySw7LK83_2(.dout(w_dff_A_hypxtFVw3_2),.din(w_dff_A_2ySw7LK83_2),.clk(gclk));
	jdff dff_A_Jkl7f8Sw0_2(.dout(w_dff_A_2ySw7LK83_2),.din(w_dff_A_Jkl7f8Sw0_2),.clk(gclk));
	jdff dff_A_E1G6jHtS0_2(.dout(w_dff_A_Jkl7f8Sw0_2),.din(w_dff_A_E1G6jHtS0_2),.clk(gclk));
	jdff dff_A_AYZHWwhS7_2(.dout(w_dff_A_E1G6jHtS0_2),.din(w_dff_A_AYZHWwhS7_2),.clk(gclk));
	jdff dff_A_qx90NEen5_2(.dout(w_dff_A_AYZHWwhS7_2),.din(w_dff_A_qx90NEen5_2),.clk(gclk));
	jdff dff_A_I2ZQzOpn0_2(.dout(w_dff_A_qx90NEen5_2),.din(w_dff_A_I2ZQzOpn0_2),.clk(gclk));
	jdff dff_A_zExR2g2s7_2(.dout(w_dff_A_I2ZQzOpn0_2),.din(w_dff_A_zExR2g2s7_2),.clk(gclk));
	jdff dff_A_ooD55aNS0_2(.dout(w_dff_A_zExR2g2s7_2),.din(w_dff_A_ooD55aNS0_2),.clk(gclk));
	jdff dff_A_m9XC5wV75_2(.dout(w_dff_A_ooD55aNS0_2),.din(w_dff_A_m9XC5wV75_2),.clk(gclk));
	jdff dff_A_AtWLHQnD3_2(.dout(w_dff_A_m9XC5wV75_2),.din(w_dff_A_AtWLHQnD3_2),.clk(gclk));
	jdff dff_A_WshjxAfQ5_2(.dout(w_dff_A_AtWLHQnD3_2),.din(w_dff_A_WshjxAfQ5_2),.clk(gclk));
	jdff dff_A_r3iUyr916_0(.dout(w_n128_0[0]),.din(w_dff_A_r3iUyr916_0),.clk(gclk));
	jdff dff_A_jbdTcvks0_0(.dout(w_dff_A_r3iUyr916_0),.din(w_dff_A_jbdTcvks0_0),.clk(gclk));
	jdff dff_A_xoEPukCl6_0(.dout(w_dff_A_jbdTcvks0_0),.din(w_dff_A_xoEPukCl6_0),.clk(gclk));
	jdff dff_A_spmvP23Z7_0(.dout(w_dff_A_xoEPukCl6_0),.din(w_dff_A_spmvP23Z7_0),.clk(gclk));
	jdff dff_A_o2LkBOIf7_0(.dout(w_dff_A_spmvP23Z7_0),.din(w_dff_A_o2LkBOIf7_0),.clk(gclk));
	jdff dff_A_ZIsEgJ3T1_0(.dout(w_dff_A_o2LkBOIf7_0),.din(w_dff_A_ZIsEgJ3T1_0),.clk(gclk));
	jdff dff_A_pP8qmPLt9_0(.dout(w_n126_0[0]),.din(w_dff_A_pP8qmPLt9_0),.clk(gclk));
	jdff dff_A_haE2X7L63_0(.dout(w_dff_A_pP8qmPLt9_0),.din(w_dff_A_haE2X7L63_0),.clk(gclk));
	jdff dff_A_vm1ylt3D2_0(.dout(w_dff_A_haE2X7L63_0),.din(w_dff_A_vm1ylt3D2_0),.clk(gclk));
	jdff dff_A_68hyfJC96_0(.dout(w_dff_A_vm1ylt3D2_0),.din(w_dff_A_68hyfJC96_0),.clk(gclk));
	jdff dff_A_3b6KP1Xr0_0(.dout(w_dff_A_68hyfJC96_0),.din(w_dff_A_3b6KP1Xr0_0),.clk(gclk));
	jdff dff_A_N6wzs6ac4_1(.dout(w_n126_0[1]),.din(w_dff_A_N6wzs6ac4_1),.clk(gclk));
	jdff dff_A_pXKmNmg82_1(.dout(w_dff_A_N6wzs6ac4_1),.din(w_dff_A_pXKmNmg82_1),.clk(gclk));
	jdff dff_A_BCsn4f764_1(.dout(w_dff_A_pXKmNmg82_1),.din(w_dff_A_BCsn4f764_1),.clk(gclk));
	jdff dff_A_gC6VUEAN1_1(.dout(w_dff_A_BCsn4f764_1),.din(w_dff_A_gC6VUEAN1_1),.clk(gclk));
	jdff dff_A_lHnmXJzK4_1(.dout(w_dff_A_gC6VUEAN1_1),.din(w_dff_A_lHnmXJzK4_1),.clk(gclk));
	jdff dff_B_s7j9ayXP8_3(.din(n126),.dout(w_dff_B_s7j9ayXP8_3),.clk(gclk));
	jdff dff_B_uEIqphoG9_3(.din(w_dff_B_s7j9ayXP8_3),.dout(w_dff_B_uEIqphoG9_3),.clk(gclk));
	jdff dff_B_CRyaFUlM7_3(.din(w_dff_B_uEIqphoG9_3),.dout(w_dff_B_CRyaFUlM7_3),.clk(gclk));
	jdff dff_B_CneCEBHj1_3(.din(w_dff_B_CRyaFUlM7_3),.dout(w_dff_B_CneCEBHj1_3),.clk(gclk));
	jdff dff_B_RXJVo6698_3(.din(w_dff_B_CneCEBHj1_3),.dout(w_dff_B_RXJVo6698_3),.clk(gclk));
	jdff dff_B_RMj0V95O8_3(.din(w_dff_B_RXJVo6698_3),.dout(w_dff_B_RMj0V95O8_3),.clk(gclk));
	jdff dff_B_YeLHtNcC6_3(.din(w_dff_B_RMj0V95O8_3),.dout(w_dff_B_YeLHtNcC6_3),.clk(gclk));
	jdff dff_A_dpeMo0y88_0(.dout(w_G86gat_1[0]),.din(w_dff_A_dpeMo0y88_0),.clk(gclk));
	jdff dff_A_ijkCNXde3_0(.dout(w_dff_A_dpeMo0y88_0),.din(w_dff_A_ijkCNXde3_0),.clk(gclk));
	jdff dff_A_7NuyewkD5_0(.dout(w_dff_A_ijkCNXde3_0),.din(w_dff_A_7NuyewkD5_0),.clk(gclk));
	jdff dff_A_ZZbdYIde3_0(.dout(w_dff_A_7NuyewkD5_0),.din(w_dff_A_ZZbdYIde3_0),.clk(gclk));
	jdff dff_A_kj0XBpzp1_0(.dout(w_dff_A_ZZbdYIde3_0),.din(w_dff_A_kj0XBpzp1_0),.clk(gclk));
	jdff dff_A_Zn33bEhK9_0(.dout(w_dff_A_kj0XBpzp1_0),.din(w_dff_A_Zn33bEhK9_0),.clk(gclk));
	jdff dff_A_GsVNaxDu9_0(.dout(w_dff_A_Zn33bEhK9_0),.din(w_dff_A_GsVNaxDu9_0),.clk(gclk));
	jdff dff_A_yjVedfVQ4_0(.dout(w_dff_A_GsVNaxDu9_0),.din(w_dff_A_yjVedfVQ4_0),.clk(gclk));
	jdff dff_A_cUR0wbUU5_1(.dout(w_G86gat_0[1]),.din(w_dff_A_cUR0wbUU5_1),.clk(gclk));
	jdff dff_A_wgigKsqo3_1(.dout(w_dff_A_cUR0wbUU5_1),.din(w_dff_A_wgigKsqo3_1),.clk(gclk));
	jdff dff_A_25UuoGTf8_1(.dout(w_dff_A_wgigKsqo3_1),.din(w_dff_A_25UuoGTf8_1),.clk(gclk));
	jdff dff_A_70nrB0SL1_1(.dout(w_dff_A_25UuoGTf8_1),.din(w_dff_A_70nrB0SL1_1),.clk(gclk));
	jdff dff_A_s3CgOHqm4_1(.dout(w_dff_A_70nrB0SL1_1),.din(w_dff_A_s3CgOHqm4_1),.clk(gclk));
	jdff dff_A_Xb2ovPJj1_1(.dout(w_dff_A_s3CgOHqm4_1),.din(w_dff_A_Xb2ovPJj1_1),.clk(gclk));
	jdff dff_A_AU1BrwiZ6_1(.dout(w_dff_A_Xb2ovPJj1_1),.din(w_dff_A_AU1BrwiZ6_1),.clk(gclk));
	jdff dff_A_fczzsLAC1_1(.dout(w_dff_A_AU1BrwiZ6_1),.din(w_dff_A_fczzsLAC1_1),.clk(gclk));
	jdff dff_A_gnbRYeN84_1(.dout(w_dff_A_fczzsLAC1_1),.din(w_dff_A_gnbRYeN84_1),.clk(gclk));
	jdff dff_A_gKc0JG244_1(.dout(w_dff_A_gnbRYeN84_1),.din(w_dff_A_gKc0JG244_1),.clk(gclk));
	jdff dff_A_SXTi0Hnn7_1(.dout(w_dff_A_gKc0JG244_1),.din(w_dff_A_SXTi0Hnn7_1),.clk(gclk));
	jdff dff_A_pfcs9OfN8_1(.dout(w_dff_A_SXTi0Hnn7_1),.din(w_dff_A_pfcs9OfN8_1),.clk(gclk));
	jdff dff_A_ypIElH5r9_1(.dout(w_dff_A_pfcs9OfN8_1),.din(w_dff_A_ypIElH5r9_1),.clk(gclk));
	jdff dff_A_DhsNUEGQ8_2(.dout(w_G86gat_0[2]),.din(w_dff_A_DhsNUEGQ8_2),.clk(gclk));
	jdff dff_A_Q8iZl7Tt0_2(.dout(w_dff_A_DhsNUEGQ8_2),.din(w_dff_A_Q8iZl7Tt0_2),.clk(gclk));
	jdff dff_A_FVuehxU57_2(.dout(w_dff_A_Q8iZl7Tt0_2),.din(w_dff_A_FVuehxU57_2),.clk(gclk));
	jdff dff_A_ur0vCEWL3_2(.dout(w_dff_A_FVuehxU57_2),.din(w_dff_A_ur0vCEWL3_2),.clk(gclk));
	jdff dff_A_eZRR2YPH3_2(.dout(w_dff_A_ur0vCEWL3_2),.din(w_dff_A_eZRR2YPH3_2),.clk(gclk));
	jdff dff_A_1x0zOaXT2_2(.dout(w_dff_A_eZRR2YPH3_2),.din(w_dff_A_1x0zOaXT2_2),.clk(gclk));
	jdff dff_A_iiorh9oP7_2(.dout(w_dff_A_1x0zOaXT2_2),.din(w_dff_A_iiorh9oP7_2),.clk(gclk));
	jdff dff_A_BFrMIyUE7_2(.dout(w_dff_A_iiorh9oP7_2),.din(w_dff_A_BFrMIyUE7_2),.clk(gclk));
	jdff dff_A_oeRkc5fA4_2(.dout(w_dff_A_BFrMIyUE7_2),.din(w_dff_A_oeRkc5fA4_2),.clk(gclk));
	jdff dff_A_b5aC0idQ3_2(.dout(w_dff_A_oeRkc5fA4_2),.din(w_dff_A_b5aC0idQ3_2),.clk(gclk));
	jdff dff_A_HU0MXQbV5_2(.dout(w_dff_A_b5aC0idQ3_2),.din(w_dff_A_HU0MXQbV5_2),.clk(gclk));
	jdff dff_A_BQt1wvsX2_2(.dout(w_dff_A_HU0MXQbV5_2),.din(w_dff_A_BQt1wvsX2_2),.clk(gclk));
	jdff dff_A_UJJOc4yD7_2(.dout(w_dff_A_BQt1wvsX2_2),.din(w_dff_A_UJJOc4yD7_2),.clk(gclk));
	jdff dff_B_5k3CBSX92_0(.din(n124),.dout(w_dff_B_5k3CBSX92_0),.clk(gclk));
	jdff dff_A_4GlHeu0d9_1(.dout(w_n123_0[1]),.din(w_dff_A_4GlHeu0d9_1),.clk(gclk));
	jdff dff_A_FZdUlzIc4_1(.dout(w_dff_A_4GlHeu0d9_1),.din(w_dff_A_FZdUlzIc4_1),.clk(gclk));
	jdff dff_A_8eFUU7KG9_1(.dout(w_dff_A_FZdUlzIc4_1),.din(w_dff_A_8eFUU7KG9_1),.clk(gclk));
	jdff dff_A_rOoHaY983_1(.dout(w_dff_A_8eFUU7KG9_1),.din(w_dff_A_rOoHaY983_1),.clk(gclk));
	jdff dff_A_pH0zxLsr9_1(.dout(w_dff_A_rOoHaY983_1),.din(w_dff_A_pH0zxLsr9_1),.clk(gclk));
	jdff dff_A_csgzIfQc0_0(.dout(w_G47gat_0[0]),.din(w_dff_A_csgzIfQc0_0),.clk(gclk));
	jdff dff_A_ozmYMCsi8_0(.dout(w_dff_A_csgzIfQc0_0),.din(w_dff_A_ozmYMCsi8_0),.clk(gclk));
	jdff dff_A_YkHsRswo6_0(.dout(w_dff_A_ozmYMCsi8_0),.din(w_dff_A_YkHsRswo6_0),.clk(gclk));
	jdff dff_A_bwUtO71m0_0(.dout(w_dff_A_YkHsRswo6_0),.din(w_dff_A_bwUtO71m0_0),.clk(gclk));
	jdff dff_A_3RpX77g78_0(.dout(w_dff_A_bwUtO71m0_0),.din(w_dff_A_3RpX77g78_0),.clk(gclk));
	jdff dff_A_IRC0wbBQ1_0(.dout(w_dff_A_3RpX77g78_0),.din(w_dff_A_IRC0wbBQ1_0),.clk(gclk));
	jdff dff_A_LZUBIv3c0_0(.dout(w_dff_A_IRC0wbBQ1_0),.din(w_dff_A_LZUBIv3c0_0),.clk(gclk));
	jdff dff_A_gbEoHlYD1_0(.dout(w_dff_A_LZUBIv3c0_0),.din(w_dff_A_gbEoHlYD1_0),.clk(gclk));
	jdff dff_A_Zav5IAPQ4_0(.dout(w_dff_A_gbEoHlYD1_0),.din(w_dff_A_Zav5IAPQ4_0),.clk(gclk));
	jdff dff_A_EuiKlArQ6_0(.dout(w_dff_A_Zav5IAPQ4_0),.din(w_dff_A_EuiKlArQ6_0),.clk(gclk));
	jdff dff_A_ukI5AOSk4_0(.dout(w_dff_A_EuiKlArQ6_0),.din(w_dff_A_ukI5AOSk4_0),.clk(gclk));
	jdff dff_A_8d6iiiZY5_0(.dout(w_dff_A_ukI5AOSk4_0),.din(w_dff_A_8d6iiiZY5_0),.clk(gclk));
	jdff dff_A_8CCDWlrJ8_0(.dout(w_dff_A_8d6iiiZY5_0),.din(w_dff_A_8CCDWlrJ8_0),.clk(gclk));
	jdff dff_B_4Zhg5uju9_1(.din(n117),.dout(w_dff_B_4Zhg5uju9_1),.clk(gclk));
	jdff dff_B_5bSR4sar3_1(.din(w_dff_B_4Zhg5uju9_1),.dout(w_dff_B_5bSR4sar3_1),.clk(gclk));
	jdff dff_B_aE9ibtFv9_1(.din(w_dff_B_5bSR4sar3_1),.dout(w_dff_B_aE9ibtFv9_1),.clk(gclk));
	jdff dff_B_LXkBdS2c5_1(.din(w_dff_B_aE9ibtFv9_1),.dout(w_dff_B_LXkBdS2c5_1),.clk(gclk));
	jdff dff_B_TzKsz0210_1(.din(w_dff_B_LXkBdS2c5_1),.dout(w_dff_B_TzKsz0210_1),.clk(gclk));
	jdff dff_B_9OUGm1OT6_1(.din(w_dff_B_TzKsz0210_1),.dout(w_dff_B_9OUGm1OT6_1),.clk(gclk));
	jdff dff_B_ffqh8P5m4_1(.din(w_dff_B_9OUGm1OT6_1),.dout(w_dff_B_ffqh8P5m4_1),.clk(gclk));
	jdff dff_A_u2o2vyNT8_0(.dout(w_G60gat_0[0]),.din(w_dff_A_u2o2vyNT8_0),.clk(gclk));
	jdff dff_A_oFDmHfkx9_0(.dout(w_dff_A_u2o2vyNT8_0),.din(w_dff_A_oFDmHfkx9_0),.clk(gclk));
	jdff dff_A_Czeu6EaD2_0(.dout(w_dff_A_oFDmHfkx9_0),.din(w_dff_A_Czeu6EaD2_0),.clk(gclk));
	jdff dff_A_WGJgCACE1_0(.dout(w_dff_A_Czeu6EaD2_0),.din(w_dff_A_WGJgCACE1_0),.clk(gclk));
	jdff dff_A_wtGrbgPE3_0(.dout(w_dff_A_WGJgCACE1_0),.din(w_dff_A_wtGrbgPE3_0),.clk(gclk));
	jdff dff_A_1VKlLrV49_0(.dout(w_dff_A_wtGrbgPE3_0),.din(w_dff_A_1VKlLrV49_0),.clk(gclk));
	jdff dff_A_fWOGl1ss9_0(.dout(w_dff_A_1VKlLrV49_0),.din(w_dff_A_fWOGl1ss9_0),.clk(gclk));
	jdff dff_A_DrY94SJ54_0(.dout(w_dff_A_fWOGl1ss9_0),.din(w_dff_A_DrY94SJ54_0),.clk(gclk));
	jdff dff_A_4UGFVwQa4_0(.dout(w_dff_A_DrY94SJ54_0),.din(w_dff_A_4UGFVwQa4_0),.clk(gclk));
	jdff dff_A_uHjulb3A4_0(.dout(w_dff_A_4UGFVwQa4_0),.din(w_dff_A_uHjulb3A4_0),.clk(gclk));
	jdff dff_A_ufPezCq83_0(.dout(w_dff_A_uHjulb3A4_0),.din(w_dff_A_ufPezCq83_0),.clk(gclk));
	jdff dff_A_HYuZOdDo6_0(.dout(w_dff_A_ufPezCq83_0),.din(w_dff_A_HYuZOdDo6_0),.clk(gclk));
	jdff dff_A_o998TikY5_0(.dout(w_dff_A_HYuZOdDo6_0),.din(w_dff_A_o998TikY5_0),.clk(gclk));
	jdff dff_A_zmSJXJog7_1(.dout(w_G60gat_0[1]),.din(w_dff_A_zmSJXJog7_1),.clk(gclk));
	jdff dff_A_3ic0lOvY4_1(.dout(w_dff_A_zmSJXJog7_1),.din(w_dff_A_3ic0lOvY4_1),.clk(gclk));
	jdff dff_A_HDFCE9Ra2_1(.dout(w_dff_A_3ic0lOvY4_1),.din(w_dff_A_HDFCE9Ra2_1),.clk(gclk));
	jdff dff_A_b3rBmTOY6_1(.dout(w_dff_A_HDFCE9Ra2_1),.din(w_dff_A_b3rBmTOY6_1),.clk(gclk));
	jdff dff_A_aE22zqi41_1(.dout(w_dff_A_b3rBmTOY6_1),.din(w_dff_A_aE22zqi41_1),.clk(gclk));
	jdff dff_A_SPppKltk8_1(.dout(w_dff_A_aE22zqi41_1),.din(w_dff_A_SPppKltk8_1),.clk(gclk));
	jdff dff_A_Gosjnvc37_1(.dout(w_dff_A_SPppKltk8_1),.din(w_dff_A_Gosjnvc37_1),.clk(gclk));
	jdff dff_A_8tObnMCA4_1(.dout(w_dff_A_Gosjnvc37_1),.din(w_dff_A_8tObnMCA4_1),.clk(gclk));
	jdff dff_A_v6NCN8Ps2_0(.dout(w_n115_0[0]),.din(w_dff_A_v6NCN8Ps2_0),.clk(gclk));
	jdff dff_A_jRWMkcb75_0(.dout(w_dff_A_v6NCN8Ps2_0),.din(w_dff_A_jRWMkcb75_0),.clk(gclk));
	jdff dff_A_OUGX0bC37_0(.dout(w_n114_0[0]),.din(w_dff_A_OUGX0bC37_0),.clk(gclk));
	jdff dff_A_PynhZ6tm3_0(.dout(w_dff_A_OUGX0bC37_0),.din(w_dff_A_PynhZ6tm3_0),.clk(gclk));
	jdff dff_A_3Viobn0g9_0(.dout(w_dff_A_PynhZ6tm3_0),.din(w_dff_A_3Viobn0g9_0),.clk(gclk));
	jdff dff_A_5YzlYxxv2_0(.dout(w_dff_A_3Viobn0g9_0),.din(w_dff_A_5YzlYxxv2_0),.clk(gclk));
	jdff dff_A_srRqU8ZK1_0(.dout(w_dff_A_5YzlYxxv2_0),.din(w_dff_A_srRqU8ZK1_0),.clk(gclk));
	jdff dff_A_vzpAS6T33_0(.dout(w_dff_A_srRqU8ZK1_0),.din(w_dff_A_vzpAS6T33_0),.clk(gclk));
	jdff dff_A_RJhHZLGL4_0(.dout(w_G34gat_0[0]),.din(w_dff_A_RJhHZLGL4_0),.clk(gclk));
	jdff dff_A_2TzZKNIi4_0(.dout(w_dff_A_RJhHZLGL4_0),.din(w_dff_A_2TzZKNIi4_0),.clk(gclk));
	jdff dff_A_6Eh1bGgI3_0(.dout(w_dff_A_2TzZKNIi4_0),.din(w_dff_A_6Eh1bGgI3_0),.clk(gclk));
	jdff dff_A_rw37N18g7_0(.dout(w_dff_A_6Eh1bGgI3_0),.din(w_dff_A_rw37N18g7_0),.clk(gclk));
	jdff dff_A_Z82C6c1h0_0(.dout(w_dff_A_rw37N18g7_0),.din(w_dff_A_Z82C6c1h0_0),.clk(gclk));
	jdff dff_A_g9BeVl5L8_0(.dout(w_dff_A_Z82C6c1h0_0),.din(w_dff_A_g9BeVl5L8_0),.clk(gclk));
	jdff dff_A_oMLDARsX4_0(.dout(w_dff_A_g9BeVl5L8_0),.din(w_dff_A_oMLDARsX4_0),.clk(gclk));
	jdff dff_A_Tlez3jKg0_0(.dout(w_dff_A_oMLDARsX4_0),.din(w_dff_A_Tlez3jKg0_0),.clk(gclk));
	jdff dff_A_wkJiHxiJ2_0(.dout(w_dff_A_Tlez3jKg0_0),.din(w_dff_A_wkJiHxiJ2_0),.clk(gclk));
	jdff dff_A_nN3psxv05_0(.dout(w_dff_A_wkJiHxiJ2_0),.din(w_dff_A_nN3psxv05_0),.clk(gclk));
	jdff dff_A_ZjkH1l7G1_0(.dout(w_dff_A_nN3psxv05_0),.din(w_dff_A_ZjkH1l7G1_0),.clk(gclk));
	jdff dff_A_LuWWhUkT2_0(.dout(w_dff_A_ZjkH1l7G1_0),.din(w_dff_A_LuWWhUkT2_0),.clk(gclk));
	jdff dff_A_45KJcNxX6_0(.dout(w_dff_A_LuWWhUkT2_0),.din(w_dff_A_45KJcNxX6_0),.clk(gclk));
	jdff dff_A_NtwJQERd5_2(.dout(w_G34gat_0[2]),.din(w_dff_A_NtwJQERd5_2),.clk(gclk));
	jdff dff_A_9Xpsc3pP8_2(.dout(w_dff_A_NtwJQERd5_2),.din(w_dff_A_9Xpsc3pP8_2),.clk(gclk));
	jdff dff_A_TH3MORgO4_2(.dout(w_dff_A_9Xpsc3pP8_2),.din(w_dff_A_TH3MORgO4_2),.clk(gclk));
	jdff dff_A_cEHnoUO15_2(.dout(w_dff_A_TH3MORgO4_2),.din(w_dff_A_cEHnoUO15_2),.clk(gclk));
	jdff dff_A_o2iQjXpM8_2(.dout(w_dff_A_cEHnoUO15_2),.din(w_dff_A_o2iQjXpM8_2),.clk(gclk));
	jdff dff_A_pBNECicw9_2(.dout(w_dff_A_o2iQjXpM8_2),.din(w_dff_A_pBNECicw9_2),.clk(gclk));
	jdff dff_A_MeAqEvjp5_2(.dout(w_dff_A_pBNECicw9_2),.din(w_dff_A_MeAqEvjp5_2),.clk(gclk));
	jdff dff_A_m4Ae2IwH6_2(.dout(w_dff_A_MeAqEvjp5_2),.din(w_dff_A_m4Ae2IwH6_2),.clk(gclk));
	jdff dff_A_Z1NYtCaj8_0(.dout(w_n109_0[0]),.din(w_dff_A_Z1NYtCaj8_0),.clk(gclk));
	jdff dff_A_xPS0zrTu1_0(.dout(w_dff_A_Z1NYtCaj8_0),.din(w_dff_A_xPS0zrTu1_0),.clk(gclk));
	jdff dff_A_CSPzgjIt2_0(.dout(w_dff_A_xPS0zrTu1_0),.din(w_dff_A_CSPzgjIt2_0),.clk(gclk));
	jdff dff_A_iUMSITCT7_0(.dout(w_dff_A_CSPzgjIt2_0),.din(w_dff_A_iUMSITCT7_0),.clk(gclk));
	jdff dff_A_IkwzG5A59_0(.dout(w_dff_A_iUMSITCT7_0),.din(w_dff_A_IkwzG5A59_0),.clk(gclk));
	jdff dff_A_9PWh6pjL1_0(.dout(w_dff_A_IkwzG5A59_0),.din(w_dff_A_9PWh6pjL1_0),.clk(gclk));
	jdff dff_A_vFMq1rc39_0(.dout(w_n107_0[0]),.din(w_dff_A_vFMq1rc39_0),.clk(gclk));
	jdff dff_A_eeQFhTtw6_0(.dout(w_dff_A_vFMq1rc39_0),.din(w_dff_A_eeQFhTtw6_0),.clk(gclk));
	jdff dff_A_CzzW6dEP2_0(.dout(w_dff_A_eeQFhTtw6_0),.din(w_dff_A_CzzW6dEP2_0),.clk(gclk));
	jdff dff_A_Jbgo1zMS7_0(.dout(w_dff_A_CzzW6dEP2_0),.din(w_dff_A_Jbgo1zMS7_0),.clk(gclk));
	jdff dff_A_uuYeohou6_0(.dout(w_dff_A_Jbgo1zMS7_0),.din(w_dff_A_uuYeohou6_0),.clk(gclk));
	jdff dff_B_D4Uj3POd5_2(.din(n107),.dout(w_dff_B_D4Uj3POd5_2),.clk(gclk));
	jdff dff_B_jBOghPDW2_2(.din(w_dff_B_D4Uj3POd5_2),.dout(w_dff_B_jBOghPDW2_2),.clk(gclk));
	jdff dff_B_EnVZQBKX5_2(.din(w_dff_B_jBOghPDW2_2),.dout(w_dff_B_EnVZQBKX5_2),.clk(gclk));
	jdff dff_B_wIHAtp7e7_2(.din(w_dff_B_EnVZQBKX5_2),.dout(w_dff_B_wIHAtp7e7_2),.clk(gclk));
	jdff dff_B_ay4QpemX4_2(.din(w_dff_B_wIHAtp7e7_2),.dout(w_dff_B_ay4QpemX4_2),.clk(gclk));
	jdff dff_B_rJT8FTI67_2(.din(w_dff_B_ay4QpemX4_2),.dout(w_dff_B_rJT8FTI67_2),.clk(gclk));
	jdff dff_B_KjPWA0K59_2(.din(w_dff_B_rJT8FTI67_2),.dout(w_dff_B_KjPWA0K59_2),.clk(gclk));
	jdff dff_A_mpdH62qh1_0(.dout(w_G73gat_0[0]),.din(w_dff_A_mpdH62qh1_0),.clk(gclk));
	jdff dff_A_LWPdWuu84_0(.dout(w_dff_A_mpdH62qh1_0),.din(w_dff_A_LWPdWuu84_0),.clk(gclk));
	jdff dff_A_ZgUd1Aqt4_0(.dout(w_dff_A_LWPdWuu84_0),.din(w_dff_A_ZgUd1Aqt4_0),.clk(gclk));
	jdff dff_A_eHl7k7d01_0(.dout(w_dff_A_ZgUd1Aqt4_0),.din(w_dff_A_eHl7k7d01_0),.clk(gclk));
	jdff dff_A_Y8Z93HIb2_0(.dout(w_dff_A_eHl7k7d01_0),.din(w_dff_A_Y8Z93HIb2_0),.clk(gclk));
	jdff dff_A_q6CIHo5f9_0(.dout(w_dff_A_Y8Z93HIb2_0),.din(w_dff_A_q6CIHo5f9_0),.clk(gclk));
	jdff dff_A_6smhHEjT0_0(.dout(w_dff_A_q6CIHo5f9_0),.din(w_dff_A_6smhHEjT0_0),.clk(gclk));
	jdff dff_A_KV79Bzcm5_0(.dout(w_dff_A_6smhHEjT0_0),.din(w_dff_A_KV79Bzcm5_0),.clk(gclk));
	jdff dff_A_dTKI1MBX9_0(.dout(w_dff_A_KV79Bzcm5_0),.din(w_dff_A_dTKI1MBX9_0),.clk(gclk));
	jdff dff_A_LAsYhJGn5_0(.dout(w_dff_A_dTKI1MBX9_0),.din(w_dff_A_LAsYhJGn5_0),.clk(gclk));
	jdff dff_A_SWVyRYqy8_0(.dout(w_dff_A_LAsYhJGn5_0),.din(w_dff_A_SWVyRYqy8_0),.clk(gclk));
	jdff dff_A_cnDCD1Ii8_0(.dout(w_dff_A_SWVyRYqy8_0),.din(w_dff_A_cnDCD1Ii8_0),.clk(gclk));
	jdff dff_A_y9vALicB7_0(.dout(w_dff_A_cnDCD1Ii8_0),.din(w_dff_A_y9vALicB7_0),.clk(gclk));
	jdff dff_A_a3vxG4wM6_1(.dout(w_G73gat_0[1]),.din(w_dff_A_a3vxG4wM6_1),.clk(gclk));
	jdff dff_A_O3xE5l1p0_1(.dout(w_dff_A_a3vxG4wM6_1),.din(w_dff_A_O3xE5l1p0_1),.clk(gclk));
	jdff dff_A_5qN9hEe05_1(.dout(w_dff_A_O3xE5l1p0_1),.din(w_dff_A_5qN9hEe05_1),.clk(gclk));
	jdff dff_A_4ppkeQfq3_1(.dout(w_dff_A_5qN9hEe05_1),.din(w_dff_A_4ppkeQfq3_1),.clk(gclk));
	jdff dff_A_axWTm94x0_1(.dout(w_dff_A_4ppkeQfq3_1),.din(w_dff_A_axWTm94x0_1),.clk(gclk));
	jdff dff_A_tAjaqahn7_1(.dout(w_dff_A_axWTm94x0_1),.din(w_dff_A_tAjaqahn7_1),.clk(gclk));
	jdff dff_A_u4zUTZK49_1(.dout(w_dff_A_tAjaqahn7_1),.din(w_dff_A_u4zUTZK49_1),.clk(gclk));
	jdff dff_A_jPiuEvLn5_1(.dout(w_dff_A_u4zUTZK49_1),.din(w_dff_A_jPiuEvLn5_1),.clk(gclk));
	jdff dff_B_3q3uJTXK0_1(.din(n103),.dout(w_dff_B_3q3uJTXK0_1),.clk(gclk));
	jdff dff_B_Webltddt5_1(.din(w_dff_B_3q3uJTXK0_1),.dout(w_dff_B_Webltddt5_1),.clk(gclk));
	jdff dff_B_OMjQFVzL0_1(.din(w_dff_B_Webltddt5_1),.dout(w_dff_B_OMjQFVzL0_1),.clk(gclk));
	jdff dff_B_rDK8Seyi0_1(.din(w_dff_B_OMjQFVzL0_1),.dout(w_dff_B_rDK8Seyi0_1),.clk(gclk));
	jdff dff_B_yOtpg76R4_1(.din(w_dff_B_rDK8Seyi0_1),.dout(w_dff_B_yOtpg76R4_1),.clk(gclk));
	jdff dff_B_rXtq5zsS2_1(.din(w_dff_B_yOtpg76R4_1),.dout(w_dff_B_rXtq5zsS2_1),.clk(gclk));
	jdff dff_B_qdZUrO3T3_1(.din(w_dff_B_rXtq5zsS2_1),.dout(w_dff_B_qdZUrO3T3_1),.clk(gclk));
	jdff dff_A_JQEkHYdL3_0(.dout(w_G99gat_0[0]),.din(w_dff_A_JQEkHYdL3_0),.clk(gclk));
	jdff dff_A_GWKBBymA1_0(.dout(w_dff_A_JQEkHYdL3_0),.din(w_dff_A_GWKBBymA1_0),.clk(gclk));
	jdff dff_A_cmp2ENYx3_0(.dout(w_dff_A_GWKBBymA1_0),.din(w_dff_A_cmp2ENYx3_0),.clk(gclk));
	jdff dff_A_xUSZTpTH2_0(.dout(w_dff_A_cmp2ENYx3_0),.din(w_dff_A_xUSZTpTH2_0),.clk(gclk));
	jdff dff_A_IWEqc1R23_0(.dout(w_dff_A_xUSZTpTH2_0),.din(w_dff_A_IWEqc1R23_0),.clk(gclk));
	jdff dff_A_TbvIWBjq9_0(.dout(w_dff_A_IWEqc1R23_0),.din(w_dff_A_TbvIWBjq9_0),.clk(gclk));
	jdff dff_A_1DRn7nos2_0(.dout(w_dff_A_TbvIWBjq9_0),.din(w_dff_A_1DRn7nos2_0),.clk(gclk));
	jdff dff_A_rNQHft9w8_0(.dout(w_dff_A_1DRn7nos2_0),.din(w_dff_A_rNQHft9w8_0),.clk(gclk));
	jdff dff_A_GtNESeLD1_1(.dout(w_G99gat_0[1]),.din(w_dff_A_GtNESeLD1_1),.clk(gclk));
	jdff dff_A_aQ06KyK50_1(.dout(w_dff_A_GtNESeLD1_1),.din(w_dff_A_aQ06KyK50_1),.clk(gclk));
	jdff dff_A_ddpr6iII0_1(.dout(w_dff_A_aQ06KyK50_1),.din(w_dff_A_ddpr6iII0_1),.clk(gclk));
	jdff dff_A_T2CNLzLk1_1(.dout(w_dff_A_ddpr6iII0_1),.din(w_dff_A_T2CNLzLk1_1),.clk(gclk));
	jdff dff_A_YAoRYpXC9_1(.dout(w_dff_A_T2CNLzLk1_1),.din(w_dff_A_YAoRYpXC9_1),.clk(gclk));
	jdff dff_A_5Fwu2crh3_1(.dout(w_dff_A_YAoRYpXC9_1),.din(w_dff_A_5Fwu2crh3_1),.clk(gclk));
	jdff dff_A_VrpypLOt1_1(.dout(w_dff_A_5Fwu2crh3_1),.din(w_dff_A_VrpypLOt1_1),.clk(gclk));
	jdff dff_A_Bhr7B5352_1(.dout(w_dff_A_VrpypLOt1_1),.din(w_dff_A_Bhr7B5352_1),.clk(gclk));
	jdff dff_A_Q2IWkCYc1_1(.dout(w_dff_A_Bhr7B5352_1),.din(w_dff_A_Q2IWkCYc1_1),.clk(gclk));
	jdff dff_A_nouaKRpp6_1(.dout(w_dff_A_Q2IWkCYc1_1),.din(w_dff_A_nouaKRpp6_1),.clk(gclk));
	jdff dff_A_R4Oqs7rj8_1(.dout(w_dff_A_nouaKRpp6_1),.din(w_dff_A_R4Oqs7rj8_1),.clk(gclk));
	jdff dff_A_h0YrqkuB4_1(.dout(w_dff_A_R4Oqs7rj8_1),.din(w_dff_A_h0YrqkuB4_1),.clk(gclk));
	jdff dff_A_pePc5qPA2_1(.dout(w_dff_A_h0YrqkuB4_1),.din(w_dff_A_pePc5qPA2_1),.clk(gclk));
	jdff dff_A_rcvFle4e1_0(.dout(w_n100_0[0]),.din(w_dff_A_rcvFle4e1_0),.clk(gclk));
	jdff dff_A_cEkoftK35_0(.dout(w_dff_A_rcvFle4e1_0),.din(w_dff_A_cEkoftK35_0),.clk(gclk));
	jdff dff_A_eHAKwe5L3_0(.dout(w_dff_A_cEkoftK35_0),.din(w_dff_A_eHAKwe5L3_0),.clk(gclk));
	jdff dff_A_FDVUoyVr7_0(.dout(w_dff_A_eHAKwe5L3_0),.din(w_dff_A_FDVUoyVr7_0),.clk(gclk));
	jdff dff_A_Ge5QTCjz0_0(.dout(w_dff_A_FDVUoyVr7_0),.din(w_dff_A_Ge5QTCjz0_0),.clk(gclk));
	jdff dff_A_adLR2nLQ3_0(.dout(w_dff_A_Ge5QTCjz0_0),.din(w_dff_A_adLR2nLQ3_0),.clk(gclk));
	jdff dff_A_R7AqDXEe5_0(.dout(w_n98_0[0]),.din(w_dff_A_R7AqDXEe5_0),.clk(gclk));
	jdff dff_A_86vIatVO8_0(.dout(w_dff_A_R7AqDXEe5_0),.din(w_dff_A_86vIatVO8_0),.clk(gclk));
	jdff dff_A_UBAAwaDD8_0(.dout(w_dff_A_86vIatVO8_0),.din(w_dff_A_UBAAwaDD8_0),.clk(gclk));
	jdff dff_A_bVLVR48x8_0(.dout(w_dff_A_UBAAwaDD8_0),.din(w_dff_A_bVLVR48x8_0),.clk(gclk));
	jdff dff_A_9ffzE9Xe7_0(.dout(w_dff_A_bVLVR48x8_0),.din(w_dff_A_9ffzE9Xe7_0),.clk(gclk));
	jdff dff_B_PzTm6c3O2_2(.din(n98),.dout(w_dff_B_PzTm6c3O2_2),.clk(gclk));
	jdff dff_B_i36PFyDq2_2(.din(w_dff_B_PzTm6c3O2_2),.dout(w_dff_B_i36PFyDq2_2),.clk(gclk));
	jdff dff_B_9ptiehQW1_2(.din(w_dff_B_i36PFyDq2_2),.dout(w_dff_B_9ptiehQW1_2),.clk(gclk));
	jdff dff_B_XuIelDCn7_2(.din(w_dff_B_9ptiehQW1_2),.dout(w_dff_B_XuIelDCn7_2),.clk(gclk));
	jdff dff_B_bpY9c6ax3_2(.din(w_dff_B_XuIelDCn7_2),.dout(w_dff_B_bpY9c6ax3_2),.clk(gclk));
	jdff dff_B_afBjiZUz2_2(.din(w_dff_B_bpY9c6ax3_2),.dout(w_dff_B_afBjiZUz2_2),.clk(gclk));
	jdff dff_B_QCuW35tF1_2(.din(w_dff_B_afBjiZUz2_2),.dout(w_dff_B_QCuW35tF1_2),.clk(gclk));
	jdff dff_A_SZC6wqwR3_0(.dout(w_G8gat_0[0]),.din(w_dff_A_SZC6wqwR3_0),.clk(gclk));
	jdff dff_A_M1ayiIXN7_0(.dout(w_dff_A_SZC6wqwR3_0),.din(w_dff_A_M1ayiIXN7_0),.clk(gclk));
	jdff dff_A_wo1WZE3S5_0(.dout(w_dff_A_M1ayiIXN7_0),.din(w_dff_A_wo1WZE3S5_0),.clk(gclk));
	jdff dff_A_wk4O4tJM6_0(.dout(w_dff_A_wo1WZE3S5_0),.din(w_dff_A_wk4O4tJM6_0),.clk(gclk));
	jdff dff_A_ILSV9DuX4_0(.dout(w_dff_A_wk4O4tJM6_0),.din(w_dff_A_ILSV9DuX4_0),.clk(gclk));
	jdff dff_A_aZLPuYJc0_0(.dout(w_dff_A_ILSV9DuX4_0),.din(w_dff_A_aZLPuYJc0_0),.clk(gclk));
	jdff dff_A_9aJeOWYx5_0(.dout(w_dff_A_aZLPuYJc0_0),.din(w_dff_A_9aJeOWYx5_0),.clk(gclk));
	jdff dff_A_EXY3HEom4_0(.dout(w_dff_A_9aJeOWYx5_0),.din(w_dff_A_EXY3HEom4_0),.clk(gclk));
	jdff dff_A_MCDfcXLz8_0(.dout(w_dff_A_EXY3HEom4_0),.din(w_dff_A_MCDfcXLz8_0),.clk(gclk));
	jdff dff_A_MNCvkhyj0_0(.dout(w_dff_A_MCDfcXLz8_0),.din(w_dff_A_MNCvkhyj0_0),.clk(gclk));
	jdff dff_A_14vY5lFt3_0(.dout(w_dff_A_MNCvkhyj0_0),.din(w_dff_A_14vY5lFt3_0),.clk(gclk));
	jdff dff_A_pIJhu4c47_0(.dout(w_dff_A_14vY5lFt3_0),.din(w_dff_A_pIJhu4c47_0),.clk(gclk));
	jdff dff_A_J7Ni8DGh5_0(.dout(w_dff_A_pIJhu4c47_0),.din(w_dff_A_J7Ni8DGh5_0),.clk(gclk));
	jdff dff_A_utQirwwC3_1(.dout(w_G8gat_0[1]),.din(w_dff_A_utQirwwC3_1),.clk(gclk));
	jdff dff_A_AxrFN8I25_1(.dout(w_dff_A_utQirwwC3_1),.din(w_dff_A_AxrFN8I25_1),.clk(gclk));
	jdff dff_A_GFC64FIF3_1(.dout(w_dff_A_AxrFN8I25_1),.din(w_dff_A_GFC64FIF3_1),.clk(gclk));
	jdff dff_A_ZBIECQ5C5_1(.dout(w_dff_A_GFC64FIF3_1),.din(w_dff_A_ZBIECQ5C5_1),.clk(gclk));
	jdff dff_A_NEOCZtZ75_1(.dout(w_dff_A_ZBIECQ5C5_1),.din(w_dff_A_NEOCZtZ75_1),.clk(gclk));
	jdff dff_A_DA87H3Es4_1(.dout(w_dff_A_NEOCZtZ75_1),.din(w_dff_A_DA87H3Es4_1),.clk(gclk));
	jdff dff_A_ElfvlMue3_1(.dout(w_dff_A_DA87H3Es4_1),.din(w_dff_A_ElfvlMue3_1),.clk(gclk));
	jdff dff_A_Y58ckHoR2_1(.dout(w_dff_A_ElfvlMue3_1),.din(w_dff_A_Y58ckHoR2_1),.clk(gclk));
	jdff dff_A_ekFSqqlX4_0(.dout(w_n96_0[0]),.din(w_dff_A_ekFSqqlX4_0),.clk(gclk));
	jdff dff_A_tjMdoZay6_0(.dout(w_dff_A_ekFSqqlX4_0),.din(w_dff_A_tjMdoZay6_0),.clk(gclk));
	jdff dff_A_cY4WZPW24_0(.dout(w_dff_A_tjMdoZay6_0),.din(w_dff_A_cY4WZPW24_0),.clk(gclk));
	jdff dff_A_YDql6qcL0_0(.dout(w_dff_A_cY4WZPW24_0),.din(w_dff_A_YDql6qcL0_0),.clk(gclk));
	jdff dff_A_IbwO6GSw7_0(.dout(w_dff_A_YDql6qcL0_0),.din(w_dff_A_IbwO6GSw7_0),.clk(gclk));
	jdff dff_A_llwuIglX9_0(.dout(w_dff_A_IbwO6GSw7_0),.din(w_dff_A_llwuIglX9_0),.clk(gclk));
	jdff dff_B_yXaZP9Tk3_1(.din(n76),.dout(w_dff_B_yXaZP9Tk3_1),.clk(gclk));
	jdff dff_B_GeUr3TFo8_1(.din(n81),.dout(w_dff_B_GeUr3TFo8_1),.clk(gclk));
	jdff dff_A_Q2lTggFU9_0(.dout(w_n89_0[0]),.din(w_dff_A_Q2lTggFU9_0),.clk(gclk));
	jdff dff_A_AzQ8sAxq0_0(.dout(w_dff_A_Q2lTggFU9_0),.din(w_dff_A_AzQ8sAxq0_0),.clk(gclk));
	jdff dff_A_1MF7ElMj4_0(.dout(w_dff_A_AzQ8sAxq0_0),.din(w_dff_A_1MF7ElMj4_0),.clk(gclk));
	jdff dff_A_UNXucoXh5_0(.dout(w_dff_A_1MF7ElMj4_0),.din(w_dff_A_UNXucoXh5_0),.clk(gclk));
	jdff dff_A_9wFwPlxX5_0(.dout(w_dff_A_UNXucoXh5_0),.din(w_dff_A_9wFwPlxX5_0),.clk(gclk));
	jdff dff_A_LSQjTqpw4_0(.dout(w_dff_A_9wFwPlxX5_0),.din(w_dff_A_LSQjTqpw4_0),.clk(gclk));
	jdff dff_A_ZraDmxQ62_0(.dout(w_n84_0[0]),.din(w_dff_A_ZraDmxQ62_0),.clk(gclk));
	jdff dff_A_Mio5T8Af3_0(.dout(w_dff_A_ZraDmxQ62_0),.din(w_dff_A_Mio5T8Af3_0),.clk(gclk));
	jdff dff_A_iYztd4Bf1_0(.dout(w_dff_A_Mio5T8Af3_0),.din(w_dff_A_iYztd4Bf1_0),.clk(gclk));
	jdff dff_A_lAR0vVB73_0(.dout(w_dff_A_iYztd4Bf1_0),.din(w_dff_A_lAR0vVB73_0),.clk(gclk));
	jdff dff_A_iipd2KGQ2_0(.dout(w_dff_A_lAR0vVB73_0),.din(w_dff_A_iipd2KGQ2_0),.clk(gclk));
	jdff dff_A_dhXW7ami4_0(.dout(w_dff_A_iipd2KGQ2_0),.din(w_dff_A_dhXW7ami4_0),.clk(gclk));
	jdff dff_A_SWdrrLUX9_0(.dout(w_n82_0[0]),.din(w_dff_A_SWdrrLUX9_0),.clk(gclk));
	jdff dff_A_Gqm0Tpox9_0(.dout(w_dff_A_SWdrrLUX9_0),.din(w_dff_A_Gqm0Tpox9_0),.clk(gclk));
	jdff dff_A_rFfxckqV0_0(.dout(w_dff_A_Gqm0Tpox9_0),.din(w_dff_A_rFfxckqV0_0),.clk(gclk));
	jdff dff_A_JFhLedmD3_0(.dout(w_dff_A_rFfxckqV0_0),.din(w_dff_A_JFhLedmD3_0),.clk(gclk));
	jdff dff_A_4JRnfKCw4_0(.dout(w_dff_A_JFhLedmD3_0),.din(w_dff_A_4JRnfKCw4_0),.clk(gclk));
	jdff dff_A_ZhhdXqXN7_0(.dout(w_dff_A_4JRnfKCw4_0),.din(w_dff_A_ZhhdXqXN7_0),.clk(gclk));
	jdff dff_A_n3iobooB0_0(.dout(w_n79_0[0]),.din(w_dff_A_n3iobooB0_0),.clk(gclk));
	jdff dff_A_H0FUpJj18_0(.dout(w_dff_A_n3iobooB0_0),.din(w_dff_A_H0FUpJj18_0),.clk(gclk));
	jdff dff_A_9Wf5qaaL2_0(.dout(w_dff_A_H0FUpJj18_0),.din(w_dff_A_9Wf5qaaL2_0),.clk(gclk));
	jdff dff_A_oJCepPFk1_0(.dout(w_dff_A_9Wf5qaaL2_0),.din(w_dff_A_oJCepPFk1_0),.clk(gclk));
	jdff dff_A_xqO1nsWH4_0(.dout(w_dff_A_oJCepPFk1_0),.din(w_dff_A_xqO1nsWH4_0),.clk(gclk));
	jdff dff_A_oDIYdEqg1_0(.dout(w_dff_A_xqO1nsWH4_0),.din(w_dff_A_oDIYdEqg1_0),.clk(gclk));
	jdff dff_A_ukL3jJRl9_0(.dout(w_n78_0[0]),.din(w_dff_A_ukL3jJRl9_0),.clk(gclk));
	jdff dff_A_30SHR6zx5_0(.dout(w_dff_A_ukL3jJRl9_0),.din(w_dff_A_30SHR6zx5_0),.clk(gclk));
	jdff dff_A_uWAAZltc2_0(.dout(w_dff_A_30SHR6zx5_0),.din(w_dff_A_uWAAZltc2_0),.clk(gclk));
	jdff dff_A_MPNdGI4x0_0(.dout(w_dff_A_uWAAZltc2_0),.din(w_dff_A_MPNdGI4x0_0),.clk(gclk));
	jdff dff_A_D6BiZbl03_0(.dout(w_n77_0[0]),.din(w_dff_A_D6BiZbl03_0),.clk(gclk));
	jdff dff_A_jEQzpy3Y2_0(.dout(w_dff_A_D6BiZbl03_0),.din(w_dff_A_jEQzpy3Y2_0),.clk(gclk));
	jdff dff_A_ZYDcdArH4_0(.dout(w_dff_A_jEQzpy3Y2_0),.din(w_dff_A_ZYDcdArH4_0),.clk(gclk));
	jdff dff_A_UMv943f01_0(.dout(w_dff_A_ZYDcdArH4_0),.din(w_dff_A_UMv943f01_0),.clk(gclk));
	jdff dff_A_oQNsq2z73_0(.dout(w_dff_A_UMv943f01_0),.din(w_dff_A_oQNsq2z73_0),.clk(gclk));
	jdff dff_A_8dZ7FzZd5_0(.dout(w_dff_A_oQNsq2z73_0),.din(w_dff_A_8dZ7FzZd5_0),.clk(gclk));
	jdff dff_A_gVLds06A3_0(.dout(w_n73_0[0]),.din(w_dff_A_gVLds06A3_0),.clk(gclk));
	jdff dff_A_HHCjlAO74_0(.dout(w_dff_A_gVLds06A3_0),.din(w_dff_A_HHCjlAO74_0),.clk(gclk));
	jdff dff_A_bVddjTpq9_0(.dout(w_dff_A_HHCjlAO74_0),.din(w_dff_A_bVddjTpq9_0),.clk(gclk));
	jdff dff_A_IKCO1RKT1_0(.dout(w_dff_A_bVddjTpq9_0),.din(w_dff_A_IKCO1RKT1_0),.clk(gclk));
	jdff dff_A_em9DAxQv6_0(.dout(w_dff_A_IKCO1RKT1_0),.din(w_dff_A_em9DAxQv6_0),.clk(gclk));
	jdff dff_A_W85tryrl8_0(.dout(w_dff_A_em9DAxQv6_0),.din(w_dff_A_W85tryrl8_0),.clk(gclk));
	jdff dff_A_XdMtB1fP9_0(.dout(w_n72_0[0]),.din(w_dff_A_XdMtB1fP9_0),.clk(gclk));
	jdff dff_A_9G8u8If34_0(.dout(w_dff_A_XdMtB1fP9_0),.din(w_dff_A_9G8u8If34_0),.clk(gclk));
	jdff dff_A_5fIA5fmE1_0(.dout(w_dff_A_9G8u8If34_0),.din(w_dff_A_5fIA5fmE1_0),.clk(gclk));
	jdff dff_A_dQi7a2mO7_0(.dout(w_dff_A_5fIA5fmE1_0),.din(w_dff_A_dQi7a2mO7_0),.clk(gclk));
	jdff dff_A_LNNNHOMc6_0(.dout(w_n71_0[0]),.din(w_dff_A_LNNNHOMc6_0),.clk(gclk));
	jdff dff_A_i3wfzIfI6_0(.dout(w_dff_A_LNNNHOMc6_0),.din(w_dff_A_i3wfzIfI6_0),.clk(gclk));
	jdff dff_A_qpbGa8nT5_0(.dout(w_dff_A_i3wfzIfI6_0),.din(w_dff_A_qpbGa8nT5_0),.clk(gclk));
	jdff dff_A_IMUSR4iz5_0(.dout(w_dff_A_qpbGa8nT5_0),.din(w_dff_A_IMUSR4iz5_0),.clk(gclk));
	jdff dff_A_wrwXWCbl9_0(.dout(w_dff_A_IMUSR4iz5_0),.din(w_dff_A_wrwXWCbl9_0),.clk(gclk));
	jdff dff_A_kqsSluya0_0(.dout(w_dff_A_wrwXWCbl9_0),.din(w_dff_A_kqsSluya0_0),.clk(gclk));
	jdff dff_A_nB5OHnJe9_0(.dout(w_n69_0[0]),.din(w_dff_A_nB5OHnJe9_0),.clk(gclk));
	jdff dff_A_t5V3gYZH1_0(.dout(w_dff_A_nB5OHnJe9_0),.din(w_dff_A_t5V3gYZH1_0),.clk(gclk));
	jdff dff_A_DJwjTZyo0_0(.dout(w_dff_A_t5V3gYZH1_0),.din(w_dff_A_DJwjTZyo0_0),.clk(gclk));
	jdff dff_A_yBuIrjD62_0(.dout(w_dff_A_DJwjTZyo0_0),.din(w_dff_A_yBuIrjD62_0),.clk(gclk));
	jdff dff_A_idV8RLow4_0(.dout(w_dff_A_yBuIrjD62_0),.din(w_dff_A_idV8RLow4_0),.clk(gclk));
	jdff dff_B_eLiWCHHm6_2(.din(n69),.dout(w_dff_B_eLiWCHHm6_2),.clk(gclk));
	jdff dff_B_dh1QZYeF1_2(.din(w_dff_B_eLiWCHHm6_2),.dout(w_dff_B_dh1QZYeF1_2),.clk(gclk));
	jdff dff_B_CjY5rhLe9_2(.din(w_dff_B_dh1QZYeF1_2),.dout(w_dff_B_CjY5rhLe9_2),.clk(gclk));
	jdff dff_B_wj4h2j8T3_2(.din(w_dff_B_CjY5rhLe9_2),.dout(w_dff_B_wj4h2j8T3_2),.clk(gclk));
	jdff dff_B_vZoE3AT62_2(.din(w_dff_B_wj4h2j8T3_2),.dout(w_dff_B_vZoE3AT62_2),.clk(gclk));
	jdff dff_B_9RWjf2qb1_2(.din(w_dff_B_vZoE3AT62_2),.dout(w_dff_B_9RWjf2qb1_2),.clk(gclk));
	jdff dff_B_YvfeFDYf2_2(.din(w_dff_B_9RWjf2qb1_2),.dout(w_dff_B_YvfeFDYf2_2),.clk(gclk));
	jdff dff_A_i6bLeDAc4_0(.dout(w_G112gat_0[0]),.din(w_dff_A_i6bLeDAc4_0),.clk(gclk));
	jdff dff_A_vC4L3q7D1_0(.dout(w_dff_A_i6bLeDAc4_0),.din(w_dff_A_vC4L3q7D1_0),.clk(gclk));
	jdff dff_A_KawixPpr7_0(.dout(w_dff_A_vC4L3q7D1_0),.din(w_dff_A_KawixPpr7_0),.clk(gclk));
	jdff dff_A_wqbPpEsF5_0(.dout(w_dff_A_KawixPpr7_0),.din(w_dff_A_wqbPpEsF5_0),.clk(gclk));
	jdff dff_A_Co7XTYEZ5_0(.dout(w_dff_A_wqbPpEsF5_0),.din(w_dff_A_Co7XTYEZ5_0),.clk(gclk));
	jdff dff_A_gSWVosat9_0(.dout(w_dff_A_Co7XTYEZ5_0),.din(w_dff_A_gSWVosat9_0),.clk(gclk));
	jdff dff_A_kRHPQ6DL8_0(.dout(w_dff_A_gSWVosat9_0),.din(w_dff_A_kRHPQ6DL8_0),.clk(gclk));
	jdff dff_A_wSdM53il8_0(.dout(w_dff_A_kRHPQ6DL8_0),.din(w_dff_A_wSdM53il8_0),.clk(gclk));
	jdff dff_A_ejcjulET7_0(.dout(w_dff_A_wSdM53il8_0),.din(w_dff_A_ejcjulET7_0),.clk(gclk));
	jdff dff_A_EW5RCved3_0(.dout(w_dff_A_ejcjulET7_0),.din(w_dff_A_EW5RCved3_0),.clk(gclk));
	jdff dff_A_vh36FAp74_0(.dout(w_dff_A_EW5RCved3_0),.din(w_dff_A_vh36FAp74_0),.clk(gclk));
	jdff dff_A_TRI6dzrh9_0(.dout(w_dff_A_vh36FAp74_0),.din(w_dff_A_TRI6dzrh9_0),.clk(gclk));
	jdff dff_A_2vpsb4yq7_0(.dout(w_dff_A_TRI6dzrh9_0),.din(w_dff_A_2vpsb4yq7_0),.clk(gclk));
	jdff dff_A_crKarmKn2_1(.dout(w_G112gat_0[1]),.din(w_dff_A_crKarmKn2_1),.clk(gclk));
	jdff dff_A_3zKzzX0o9_1(.dout(w_dff_A_crKarmKn2_1),.din(w_dff_A_3zKzzX0o9_1),.clk(gclk));
	jdff dff_A_XloKwHC65_1(.dout(w_dff_A_3zKzzX0o9_1),.din(w_dff_A_XloKwHC65_1),.clk(gclk));
	jdff dff_A_6R0rSIKA8_1(.dout(w_dff_A_XloKwHC65_1),.din(w_dff_A_6R0rSIKA8_1),.clk(gclk));
	jdff dff_A_wwSvJ7zs2_1(.dout(w_dff_A_6R0rSIKA8_1),.din(w_dff_A_wwSvJ7zs2_1),.clk(gclk));
	jdff dff_A_21dRWtTN0_1(.dout(w_dff_A_wwSvJ7zs2_1),.din(w_dff_A_21dRWtTN0_1),.clk(gclk));
	jdff dff_A_ke5TfXVn5_1(.dout(w_dff_A_21dRWtTN0_1),.din(w_dff_A_ke5TfXVn5_1),.clk(gclk));
	jdff dff_A_JXS19OY08_1(.dout(w_dff_A_ke5TfXVn5_1),.din(w_dff_A_JXS19OY08_1),.clk(gclk));
	jdff dff_A_4vVSVNWb9_1(.dout(w_n139_0[1]),.din(w_dff_A_4vVSVNWb9_1),.clk(gclk));
	jdff dff_A_pF42VPeW3_1(.dout(w_dff_A_4vVSVNWb9_1),.din(w_dff_A_pF42VPeW3_1),.clk(gclk));
	jdff dff_A_wXbEfXpi6_1(.dout(w_dff_A_pF42VPeW3_1),.din(w_dff_A_wXbEfXpi6_1),.clk(gclk));
	jdff dff_A_81SzDoTd9_1(.dout(w_dff_A_wXbEfXpi6_1),.din(w_dff_A_81SzDoTd9_1),.clk(gclk));
	jdff dff_A_8Q4eDf5T1_1(.dout(w_dff_A_81SzDoTd9_1),.din(w_dff_A_8Q4eDf5T1_1),.clk(gclk));
	jdff dff_A_fT9wljA27_1(.dout(w_dff_A_8Q4eDf5T1_1),.din(w_dff_A_fT9wljA27_1),.clk(gclk));
	jdff dff_B_MZVBPHjq7_1(.din(n50),.dout(w_dff_B_MZVBPHjq7_1),.clk(gclk));
	jdff dff_B_kYIEF2aV8_1(.din(n55),.dout(w_dff_B_kYIEF2aV8_1),.clk(gclk));
	jdff dff_A_1vJ2ygwZ1_0(.dout(w_G4gat_0[0]),.din(w_dff_A_1vJ2ygwZ1_0),.clk(gclk));
	jdff dff_A_6RBbb3pF8_0(.dout(w_dff_A_1vJ2ygwZ1_0),.din(w_dff_A_6RBbb3pF8_0),.clk(gclk));
	jdff dff_A_QL0JVbtg7_0(.dout(w_dff_A_6RBbb3pF8_0),.din(w_dff_A_QL0JVbtg7_0),.clk(gclk));
	jdff dff_A_zN7L9Xib5_0(.dout(w_dff_A_QL0JVbtg7_0),.din(w_dff_A_zN7L9Xib5_0),.clk(gclk));
	jdff dff_A_P4LtSjGT5_0(.dout(w_dff_A_zN7L9Xib5_0),.din(w_dff_A_P4LtSjGT5_0),.clk(gclk));
	jdff dff_A_qsw5L1xA1_0(.dout(w_dff_A_P4LtSjGT5_0),.din(w_dff_A_qsw5L1xA1_0),.clk(gclk));
	jdff dff_A_FJepJW0D0_0(.dout(w_dff_A_qsw5L1xA1_0),.din(w_dff_A_FJepJW0D0_0),.clk(gclk));
	jdff dff_A_tllPJFyQ9_2(.dout(w_G4gat_0[2]),.din(w_dff_A_tllPJFyQ9_2),.clk(gclk));
	jdff dff_A_aFNVmE5J3_0(.dout(w_n63_0[0]),.din(w_dff_A_aFNVmE5J3_0),.clk(gclk));
	jdff dff_A_q9UiaNJr3_0(.dout(w_dff_A_aFNVmE5J3_0),.din(w_dff_A_q9UiaNJr3_0),.clk(gclk));
	jdff dff_A_GWRWYNmk2_0(.dout(w_dff_A_q9UiaNJr3_0),.din(w_dff_A_GWRWYNmk2_0),.clk(gclk));
	jdff dff_A_W7duW0aV2_0(.dout(w_dff_A_GWRWYNmk2_0),.din(w_dff_A_W7duW0aV2_0),.clk(gclk));
	jdff dff_A_yDrnNUkO3_0(.dout(w_dff_A_W7duW0aV2_0),.din(w_dff_A_yDrnNUkO3_0),.clk(gclk));
	jdff dff_A_F3BcyRrH7_0(.dout(w_G1gat_0[0]),.din(w_dff_A_F3BcyRrH7_0),.clk(gclk));
	jdff dff_A_ANIxLGii8_0(.dout(w_dff_A_F3BcyRrH7_0),.din(w_dff_A_ANIxLGii8_0),.clk(gclk));
	jdff dff_A_mKfXLHxv0_0(.dout(w_dff_A_ANIxLGii8_0),.din(w_dff_A_mKfXLHxv0_0),.clk(gclk));
	jdff dff_A_iBwruxZa9_0(.dout(w_dff_A_mKfXLHxv0_0),.din(w_dff_A_iBwruxZa9_0),.clk(gclk));
	jdff dff_A_KWdeIHcj1_0(.dout(w_dff_A_iBwruxZa9_0),.din(w_dff_A_KWdeIHcj1_0),.clk(gclk));
	jdff dff_A_uyyDderI0_0(.dout(w_dff_A_KWdeIHcj1_0),.din(w_dff_A_uyyDderI0_0),.clk(gclk));
	jdff dff_A_hOBi2wgc9_1(.dout(w_G1gat_0[1]),.din(w_dff_A_hOBi2wgc9_1),.clk(gclk));
	jdff dff_A_GSIA5rLJ5_0(.dout(w_n61_0[0]),.din(w_dff_A_GSIA5rLJ5_0),.clk(gclk));
	jdff dff_A_723ZUFy59_0(.dout(w_dff_A_GSIA5rLJ5_0),.din(w_dff_A_723ZUFy59_0),.clk(gclk));
	jdff dff_A_q5Fur47B7_0(.dout(w_dff_A_723ZUFy59_0),.din(w_dff_A_q5Fur47B7_0),.clk(gclk));
	jdff dff_A_LbHL6NVU9_0(.dout(w_dff_A_q5Fur47B7_0),.din(w_dff_A_LbHL6NVU9_0),.clk(gclk));
	jdff dff_A_bTB9zVMv4_0(.dout(w_dff_A_LbHL6NVU9_0),.din(w_dff_A_bTB9zVMv4_0),.clk(gclk));
	jdff dff_A_xEJAJHoi6_0(.dout(w_G89gat_0[0]),.din(w_dff_A_xEJAJHoi6_0),.clk(gclk));
	jdff dff_A_GL4kS4WD9_0(.dout(w_dff_A_xEJAJHoi6_0),.din(w_dff_A_GL4kS4WD9_0),.clk(gclk));
	jdff dff_A_J6MpdPul1_0(.dout(w_dff_A_GL4kS4WD9_0),.din(w_dff_A_J6MpdPul1_0),.clk(gclk));
	jdff dff_A_4pCo5JOC1_0(.dout(w_dff_A_J6MpdPul1_0),.din(w_dff_A_4pCo5JOC1_0),.clk(gclk));
	jdff dff_A_lq3ZaFkm9_0(.dout(w_dff_A_4pCo5JOC1_0),.din(w_dff_A_lq3ZaFkm9_0),.clk(gclk));
	jdff dff_A_vkNPP3Cd8_0(.dout(w_dff_A_lq3ZaFkm9_0),.din(w_dff_A_vkNPP3Cd8_0),.clk(gclk));
	jdff dff_A_h9q6CtEl3_1(.dout(w_G89gat_0[1]),.din(w_dff_A_h9q6CtEl3_1),.clk(gclk));
	jdff dff_A_eYpRitAm5_0(.dout(w_G56gat_0[0]),.din(w_dff_A_eYpRitAm5_0),.clk(gclk));
	jdff dff_A_19lApDpL0_0(.dout(w_dff_A_eYpRitAm5_0),.din(w_dff_A_19lApDpL0_0),.clk(gclk));
	jdff dff_A_CI2VMVur5_0(.dout(w_dff_A_19lApDpL0_0),.din(w_dff_A_CI2VMVur5_0),.clk(gclk));
	jdff dff_A_4Lsd1Qer8_0(.dout(w_dff_A_CI2VMVur5_0),.din(w_dff_A_4Lsd1Qer8_0),.clk(gclk));
	jdff dff_A_56joeSDb3_0(.dout(w_dff_A_4Lsd1Qer8_0),.din(w_dff_A_56joeSDb3_0),.clk(gclk));
	jdff dff_A_L7JyQjFO9_0(.dout(w_dff_A_56joeSDb3_0),.din(w_dff_A_L7JyQjFO9_0),.clk(gclk));
	jdff dff_A_Qc6vKUw11_0(.dout(w_dff_A_L7JyQjFO9_0),.din(w_dff_A_Qc6vKUw11_0),.clk(gclk));
	jdff dff_A_8P84km3w1_2(.dout(w_G56gat_0[2]),.din(w_dff_A_8P84km3w1_2),.clk(gclk));
	jdff dff_A_r6nconcD2_0(.dout(w_n58_0[0]),.din(w_dff_A_r6nconcD2_0),.clk(gclk));
	jdff dff_A_qmWZ6wVP1_0(.dout(w_dff_A_r6nconcD2_0),.din(w_dff_A_qmWZ6wVP1_0),.clk(gclk));
	jdff dff_A_mlZFzwlZ2_0(.dout(w_dff_A_qmWZ6wVP1_0),.din(w_dff_A_mlZFzwlZ2_0),.clk(gclk));
	jdff dff_A_heu4L1Ns7_0(.dout(w_dff_A_mlZFzwlZ2_0),.din(w_dff_A_heu4L1Ns7_0),.clk(gclk));
	jdff dff_A_gGvRmQIr2_0(.dout(w_dff_A_heu4L1Ns7_0),.din(w_dff_A_gGvRmQIr2_0),.clk(gclk));
	jdff dff_A_16be6FTn1_0(.dout(w_G50gat_0[0]),.din(w_dff_A_16be6FTn1_0),.clk(gclk));
	jdff dff_A_z53fshU91_0(.dout(w_dff_A_16be6FTn1_0),.din(w_dff_A_z53fshU91_0),.clk(gclk));
	jdff dff_A_eiLlJu3o9_0(.dout(w_dff_A_z53fshU91_0),.din(w_dff_A_eiLlJu3o9_0),.clk(gclk));
	jdff dff_A_nwM5npPn8_0(.dout(w_dff_A_eiLlJu3o9_0),.din(w_dff_A_nwM5npPn8_0),.clk(gclk));
	jdff dff_A_D9EtDKU45_0(.dout(w_dff_A_nwM5npPn8_0),.din(w_dff_A_D9EtDKU45_0),.clk(gclk));
	jdff dff_A_5wj2Tdsz1_0(.dout(w_dff_A_D9EtDKU45_0),.din(w_dff_A_5wj2Tdsz1_0),.clk(gclk));
	jdff dff_A_XzzsQ4iL7_1(.dout(w_G50gat_0[1]),.din(w_dff_A_XzzsQ4iL7_1),.clk(gclk));
	jdff dff_A_7kEGWqiZ8_0(.dout(w_G108gat_0[0]),.din(w_dff_A_7kEGWqiZ8_0),.clk(gclk));
	jdff dff_A_gROs3v982_0(.dout(w_dff_A_7kEGWqiZ8_0),.din(w_dff_A_gROs3v982_0),.clk(gclk));
	jdff dff_A_D2f2dGQv1_0(.dout(w_dff_A_gROs3v982_0),.din(w_dff_A_D2f2dGQv1_0),.clk(gclk));
	jdff dff_A_iN9Vgaa21_0(.dout(w_dff_A_D2f2dGQv1_0),.din(w_dff_A_iN9Vgaa21_0),.clk(gclk));
	jdff dff_A_xgzCq0VH2_0(.dout(w_dff_A_iN9Vgaa21_0),.din(w_dff_A_xgzCq0VH2_0),.clk(gclk));
	jdff dff_A_R4XptZOV1_0(.dout(w_dff_A_xgzCq0VH2_0),.din(w_dff_A_R4XptZOV1_0),.clk(gclk));
	jdff dff_A_VPLfegx98_0(.dout(w_dff_A_R4XptZOV1_0),.din(w_dff_A_VPLfegx98_0),.clk(gclk));
	jdff dff_A_qB1wV2iS1_2(.dout(w_G108gat_0[2]),.din(w_dff_A_qB1wV2iS1_2),.clk(gclk));
	jdff dff_A_Q9A4t4oZ2_0(.dout(w_n56_0[0]),.din(w_dff_A_Q9A4t4oZ2_0),.clk(gclk));
	jdff dff_A_ijNO9qvH3_0(.dout(w_dff_A_Q9A4t4oZ2_0),.din(w_dff_A_ijNO9qvH3_0),.clk(gclk));
	jdff dff_A_6qP1UmU47_0(.dout(w_dff_A_ijNO9qvH3_0),.din(w_dff_A_6qP1UmU47_0),.clk(gclk));
	jdff dff_A_ebFzpK3i2_0(.dout(w_dff_A_6qP1UmU47_0),.din(w_dff_A_ebFzpK3i2_0),.clk(gclk));
	jdff dff_A_bpBTlwkC8_0(.dout(w_dff_A_ebFzpK3i2_0),.din(w_dff_A_bpBTlwkC8_0),.clk(gclk));
	jdff dff_A_U1eOvkav8_0(.dout(w_G102gat_0[0]),.din(w_dff_A_U1eOvkav8_0),.clk(gclk));
	jdff dff_A_mi5VXx440_0(.dout(w_dff_A_U1eOvkav8_0),.din(w_dff_A_mi5VXx440_0),.clk(gclk));
	jdff dff_A_wz2EMHLE2_0(.dout(w_dff_A_mi5VXx440_0),.din(w_dff_A_wz2EMHLE2_0),.clk(gclk));
	jdff dff_A_WshWNZHf5_0(.dout(w_dff_A_wz2EMHLE2_0),.din(w_dff_A_WshWNZHf5_0),.clk(gclk));
	jdff dff_A_HHmNheJy3_0(.dout(w_dff_A_WshWNZHf5_0),.din(w_dff_A_HHmNheJy3_0),.clk(gclk));
	jdff dff_A_AQOtljhc9_0(.dout(w_dff_A_HHmNheJy3_0),.din(w_dff_A_AQOtljhc9_0),.clk(gclk));
	jdff dff_A_MKhlq43s3_1(.dout(w_G102gat_0[1]),.din(w_dff_A_MKhlq43s3_1),.clk(gclk));
	jdff dff_A_6bT09feS3_0(.dout(w_G69gat_0[0]),.din(w_dff_A_6bT09feS3_0),.clk(gclk));
	jdff dff_A_TLeHMkFY5_0(.dout(w_dff_A_6bT09feS3_0),.din(w_dff_A_TLeHMkFY5_0),.clk(gclk));
	jdff dff_A_o8nSjWMa0_0(.dout(w_dff_A_TLeHMkFY5_0),.din(w_dff_A_o8nSjWMa0_0),.clk(gclk));
	jdff dff_A_nTkSz7U96_0(.dout(w_dff_A_o8nSjWMa0_0),.din(w_dff_A_nTkSz7U96_0),.clk(gclk));
	jdff dff_A_yA2vNyT90_0(.dout(w_dff_A_nTkSz7U96_0),.din(w_dff_A_yA2vNyT90_0),.clk(gclk));
	jdff dff_A_snST9etI2_0(.dout(w_dff_A_yA2vNyT90_0),.din(w_dff_A_snST9etI2_0),.clk(gclk));
	jdff dff_A_x6jLjakQ4_0(.dout(w_dff_A_snST9etI2_0),.din(w_dff_A_x6jLjakQ4_0),.clk(gclk));
	jdff dff_A_H1t0GsEX5_2(.dout(w_G69gat_0[2]),.din(w_dff_A_H1t0GsEX5_2),.clk(gclk));
	jdff dff_A_8WrG7YFw8_0(.dout(w_n53_0[0]),.din(w_dff_A_8WrG7YFw8_0),.clk(gclk));
	jdff dff_A_LdgkSa4K8_0(.dout(w_dff_A_8WrG7YFw8_0),.din(w_dff_A_LdgkSa4K8_0),.clk(gclk));
	jdff dff_A_TDApIbAT0_0(.dout(w_dff_A_LdgkSa4K8_0),.din(w_dff_A_TDApIbAT0_0),.clk(gclk));
	jdff dff_A_cutebYfY3_0(.dout(w_dff_A_TDApIbAT0_0),.din(w_dff_A_cutebYfY3_0),.clk(gclk));
	jdff dff_A_ivBejZGA4_0(.dout(w_dff_A_cutebYfY3_0),.din(w_dff_A_ivBejZGA4_0),.clk(gclk));
	jdff dff_A_ywGF07Yt5_0(.dout(w_G63gat_0[0]),.din(w_dff_A_ywGF07Yt5_0),.clk(gclk));
	jdff dff_A_Mh2jNOs57_0(.dout(w_dff_A_ywGF07Yt5_0),.din(w_dff_A_Mh2jNOs57_0),.clk(gclk));
	jdff dff_A_AJfO7qUL3_0(.dout(w_dff_A_Mh2jNOs57_0),.din(w_dff_A_AJfO7qUL3_0),.clk(gclk));
	jdff dff_A_wajLPQZG6_0(.dout(w_dff_A_AJfO7qUL3_0),.din(w_dff_A_wajLPQZG6_0),.clk(gclk));
	jdff dff_A_R19Yk38P5_0(.dout(w_dff_A_wajLPQZG6_0),.din(w_dff_A_R19Yk38P5_0),.clk(gclk));
	jdff dff_A_N0thLyMm9_0(.dout(w_dff_A_R19Yk38P5_0),.din(w_dff_A_N0thLyMm9_0),.clk(gclk));
	jdff dff_A_XJYSseO16_1(.dout(w_G63gat_0[1]),.din(w_dff_A_XJYSseO16_1),.clk(gclk));
	jdff dff_A_gFEi0ILJ0_0(.dout(w_n52_0[0]),.din(w_dff_A_gFEi0ILJ0_0),.clk(gclk));
	jdff dff_A_L5ZhjltH9_0(.dout(w_dff_A_gFEi0ILJ0_0),.din(w_dff_A_L5ZhjltH9_0),.clk(gclk));
	jdff dff_A_btfbrcGR5_0(.dout(w_dff_A_L5ZhjltH9_0),.din(w_dff_A_btfbrcGR5_0),.clk(gclk));
	jdff dff_A_AD4OIk8E3_0(.dout(w_dff_A_btfbrcGR5_0),.din(w_dff_A_AD4OIk8E3_0),.clk(gclk));
	jdff dff_A_9MNA8pJX2_1(.dout(w_G43gat_1[1]),.din(w_dff_A_9MNA8pJX2_1),.clk(gclk));
	jdff dff_A_p2oaRg9A0_1(.dout(w_G43gat_0[1]),.din(w_dff_A_p2oaRg9A0_1),.clk(gclk));
	jdff dff_A_XkeiPx5T6_2(.dout(w_G43gat_0[2]),.din(w_dff_A_XkeiPx5T6_2),.clk(gclk));
	jdff dff_A_YLBqApx23_0(.dout(w_G37gat_0[0]),.din(w_dff_A_YLBqApx23_0),.clk(gclk));
	jdff dff_A_5Clu7xMq9_0(.dout(w_dff_A_YLBqApx23_0),.din(w_dff_A_5Clu7xMq9_0),.clk(gclk));
	jdff dff_A_3BxagBXD6_0(.dout(w_dff_A_5Clu7xMq9_0),.din(w_dff_A_3BxagBXD6_0),.clk(gclk));
	jdff dff_A_P8dVwl946_0(.dout(w_dff_A_3BxagBXD6_0),.din(w_dff_A_P8dVwl946_0),.clk(gclk));
	jdff dff_A_LZjoW5Q68_0(.dout(w_dff_A_P8dVwl946_0),.din(w_dff_A_LZjoW5Q68_0),.clk(gclk));
	jdff dff_A_ZmRpUAqN5_0(.dout(w_dff_A_LZjoW5Q68_0),.din(w_dff_A_ZmRpUAqN5_0),.clk(gclk));
	jdff dff_A_Il4LI20s8_1(.dout(w_G37gat_0[1]),.din(w_dff_A_Il4LI20s8_1),.clk(gclk));
	jdff dff_A_673eak7Z5_0(.dout(w_G17gat_0[0]),.din(w_dff_A_673eak7Z5_0),.clk(gclk));
	jdff dff_A_JPTUn46c8_0(.dout(w_dff_A_673eak7Z5_0),.din(w_dff_A_JPTUn46c8_0),.clk(gclk));
	jdff dff_A_xtCuV8GB0_0(.dout(w_dff_A_JPTUn46c8_0),.din(w_dff_A_xtCuV8GB0_0),.clk(gclk));
	jdff dff_A_ptLf8Aei8_0(.dout(w_dff_A_xtCuV8GB0_0),.din(w_dff_A_ptLf8Aei8_0),.clk(gclk));
	jdff dff_A_DY5M21Eq8_0(.dout(w_dff_A_ptLf8Aei8_0),.din(w_dff_A_DY5M21Eq8_0),.clk(gclk));
	jdff dff_A_lE9BPisZ9_0(.dout(w_dff_A_DY5M21Eq8_0),.din(w_dff_A_lE9BPisZ9_0),.clk(gclk));
	jdff dff_A_bC3ynXnv7_0(.dout(w_dff_A_lE9BPisZ9_0),.din(w_dff_A_bC3ynXnv7_0),.clk(gclk));
	jdff dff_A_9GN6vBZw5_2(.dout(w_G17gat_0[2]),.din(w_dff_A_9GN6vBZw5_2),.clk(gclk));
	jdff dff_A_6cZUH2EU9_0(.dout(w_n47_0[0]),.din(w_dff_A_6cZUH2EU9_0),.clk(gclk));
	jdff dff_A_wISLR8sa1_0(.dout(w_dff_A_6cZUH2EU9_0),.din(w_dff_A_wISLR8sa1_0),.clk(gclk));
	jdff dff_A_G0wiSCUW8_0(.dout(w_dff_A_wISLR8sa1_0),.din(w_dff_A_G0wiSCUW8_0),.clk(gclk));
	jdff dff_A_3FZBqs5V4_0(.dout(w_dff_A_G0wiSCUW8_0),.din(w_dff_A_3FZBqs5V4_0),.clk(gclk));
	jdff dff_A_4sFDhFEl2_0(.dout(w_dff_A_3FZBqs5V4_0),.din(w_dff_A_4sFDhFEl2_0),.clk(gclk));
	jdff dff_A_NwJ9YEFb4_0(.dout(w_G11gat_0[0]),.din(w_dff_A_NwJ9YEFb4_0),.clk(gclk));
	jdff dff_A_PYGxBhqM6_0(.dout(w_dff_A_NwJ9YEFb4_0),.din(w_dff_A_PYGxBhqM6_0),.clk(gclk));
	jdff dff_A_35RAxjnE0_0(.dout(w_dff_A_PYGxBhqM6_0),.din(w_dff_A_35RAxjnE0_0),.clk(gclk));
	jdff dff_A_r117srsO3_0(.dout(w_dff_A_35RAxjnE0_0),.din(w_dff_A_r117srsO3_0),.clk(gclk));
	jdff dff_A_oCqD4GS20_0(.dout(w_dff_A_r117srsO3_0),.din(w_dff_A_oCqD4GS20_0),.clk(gclk));
	jdff dff_A_HkqsB3iX6_0(.dout(w_dff_A_oCqD4GS20_0),.din(w_dff_A_HkqsB3iX6_0),.clk(gclk));
	jdff dff_A_FoogvTwZ9_1(.dout(w_G11gat_0[1]),.din(w_dff_A_FoogvTwZ9_1),.clk(gclk));
	jdff dff_A_r7zmGIrz2_1(.dout(w_G30gat_0[1]),.din(w_dff_A_r7zmGIrz2_1),.clk(gclk));
	jdff dff_A_jsqxPSei4_0(.dout(w_G24gat_0[0]),.din(w_dff_A_jsqxPSei4_0),.clk(gclk));
	jdff dff_A_hLMVnkT17_1(.dout(w_n44_0[1]),.din(w_dff_A_hLMVnkT17_1),.clk(gclk));
	jdff dff_A_owbfHAUL9_1(.dout(w_G82gat_0[1]),.din(w_dff_A_owbfHAUL9_1),.clk(gclk));
	jdff dff_A_GaW1e9fz9_1(.dout(w_dff_A_owbfHAUL9_1),.din(w_dff_A_GaW1e9fz9_1),.clk(gclk));
	jdff dff_A_dSE75Enq1_1(.dout(w_dff_A_GaW1e9fz9_1),.din(w_dff_A_dSE75Enq1_1),.clk(gclk));
	jdff dff_A_4hZwDtfK5_1(.dout(w_dff_A_dSE75Enq1_1),.din(w_dff_A_4hZwDtfK5_1),.clk(gclk));
	jdff dff_A_gEgxyzuw3_1(.dout(w_dff_A_4hZwDtfK5_1),.din(w_dff_A_gEgxyzuw3_1),.clk(gclk));
	jdff dff_A_OMt7C9BY0_1(.dout(w_dff_A_gEgxyzuw3_1),.din(w_dff_A_OMt7C9BY0_1),.clk(gclk));
	jdff dff_A_Oq19nnOW7_1(.dout(w_dff_A_OMt7C9BY0_1),.din(w_dff_A_Oq19nnOW7_1),.clk(gclk));
	jdff dff_A_0LFFT8AU3_2(.dout(w_G82gat_0[2]),.din(w_dff_A_0LFFT8AU3_2),.clk(gclk));
	jdff dff_A_cLHpH9ki5_0(.dout(w_n43_0[0]),.din(w_dff_A_cLHpH9ki5_0),.clk(gclk));
	jdff dff_A_tzaD2OSm9_0(.dout(w_dff_A_cLHpH9ki5_0),.din(w_dff_A_tzaD2OSm9_0),.clk(gclk));
	jdff dff_A_zRYPA6M31_0(.dout(w_dff_A_tzaD2OSm9_0),.din(w_dff_A_zRYPA6M31_0),.clk(gclk));
	jdff dff_A_NXNV4o3y8_0(.dout(w_dff_A_zRYPA6M31_0),.din(w_dff_A_NXNV4o3y8_0),.clk(gclk));
	jdff dff_A_60Isjg0p8_0(.dout(w_dff_A_NXNV4o3y8_0),.din(w_dff_A_60Isjg0p8_0),.clk(gclk));
	jdff dff_A_WYlnxJGX6_0(.dout(w_G76gat_0[0]),.din(w_dff_A_WYlnxJGX6_0),.clk(gclk));
	jdff dff_A_LnK4VPRl1_0(.dout(w_dff_A_WYlnxJGX6_0),.din(w_dff_A_LnK4VPRl1_0),.clk(gclk));
	jdff dff_A_BHxn3vWE5_0(.dout(w_dff_A_LnK4VPRl1_0),.din(w_dff_A_BHxn3vWE5_0),.clk(gclk));
	jdff dff_A_QoauDusf9_0(.dout(w_dff_A_BHxn3vWE5_0),.din(w_dff_A_QoauDusf9_0),.clk(gclk));
	jdff dff_A_lMTmNFar2_0(.dout(w_dff_A_QoauDusf9_0),.din(w_dff_A_lMTmNFar2_0),.clk(gclk));
	jdff dff_A_IwzqA2iF0_0(.dout(w_dff_A_lMTmNFar2_0),.din(w_dff_A_IwzqA2iF0_0),.clk(gclk));
	jdff dff_A_nFiQWkQe2_0(.dout(w_n87_0[0]),.din(w_dff_A_nFiQWkQe2_0),.clk(gclk));
	jdff dff_A_02sEIOQc0_0(.dout(w_dff_A_nFiQWkQe2_0),.din(w_dff_A_02sEIOQc0_0),.clk(gclk));
	jdff dff_A_CQV93wuJ5_0(.dout(w_dff_A_02sEIOQc0_0),.din(w_dff_A_CQV93wuJ5_0),.clk(gclk));
	jdff dff_A_2Rh298mt6_0(.dout(w_dff_A_CQV93wuJ5_0),.din(w_dff_A_2Rh298mt6_0),.clk(gclk));
	jdff dff_A_8LxJD7Ka4_0(.dout(w_dff_A_2Rh298mt6_0),.din(w_dff_A_8LxJD7Ka4_0),.clk(gclk));
	jdff dff_A_98SxYP9q9_0(.dout(w_dff_A_8LxJD7Ka4_0),.din(w_dff_A_98SxYP9q9_0),.clk(gclk));
	jdff dff_A_R7wHTQLs5_0(.dout(w_G95gat_0[0]),.din(w_dff_A_R7wHTQLs5_0),.clk(gclk));
	jdff dff_A_8Lbhp4gN7_0(.dout(w_dff_A_R7wHTQLs5_0),.din(w_dff_A_8Lbhp4gN7_0),.clk(gclk));
	jdff dff_A_grhwHU0Q5_0(.dout(w_dff_A_8Lbhp4gN7_0),.din(w_dff_A_grhwHU0Q5_0),.clk(gclk));
	jdff dff_A_GBMHBtLC7_0(.dout(w_dff_A_grhwHU0Q5_0),.din(w_dff_A_GBMHBtLC7_0),.clk(gclk));
	jdff dff_A_Ef0k35ne1_0(.dout(w_dff_A_GBMHBtLC7_0),.din(w_dff_A_Ef0k35ne1_0),.clk(gclk));
	jdff dff_A_u40iQJzv7_0(.dout(w_dff_A_Ef0k35ne1_0),.din(w_dff_A_u40iQJzv7_0),.clk(gclk));
	jdff dff_A_6YUz5bTd3_0(.dout(w_dff_A_u40iQJzv7_0),.din(w_dff_A_6YUz5bTd3_0),.clk(gclk));
	jdff dff_A_ArKlI0YR1_2(.dout(w_G95gat_0[2]),.din(w_dff_A_ArKlI0YR1_2),.clk(gclk));
	jdff dff_A_yDeajRKO1_1(.dout(w_G105gat_0[1]),.din(w_dff_A_yDeajRKO1_1),.clk(gclk));
	jdff dff_A_q5Bwaxhn3_1(.dout(w_dff_A_yDeajRKO1_1),.din(w_dff_A_q5Bwaxhn3_1),.clk(gclk));
	jdff dff_A_yCPbTmvH4_1(.dout(w_dff_A_q5Bwaxhn3_1),.din(w_dff_A_yCPbTmvH4_1),.clk(gclk));
	jdff dff_A_FnpqAHZ88_1(.dout(w_dff_A_yCPbTmvH4_1),.din(w_dff_A_FnpqAHZ88_1),.clk(gclk));
	jdff dff_A_qrGkmUSR3_1(.dout(w_dff_A_FnpqAHZ88_1),.din(w_dff_A_qrGkmUSR3_1),.clk(gclk));
	jdff dff_A_DpwkpF1e4_1(.dout(w_dff_A_qrGkmUSR3_1),.din(w_dff_A_DpwkpF1e4_1),.clk(gclk));
	jdff dff_A_uih7FaRx8_1(.dout(w_dff_A_DpwkpF1e4_1),.din(w_dff_A_uih7FaRx8_1),.clk(gclk));
	jdff dff_A_cKzUmcT47_1(.dout(w_dff_A_uih7FaRx8_1),.din(w_dff_A_cKzUmcT47_1),.clk(gclk));
	jdff dff_A_KEF28kuZ3_1(.dout(w_dff_A_cKzUmcT47_1),.din(w_dff_A_KEF28kuZ3_1),.clk(gclk));
	jdff dff_A_VlnhQV3B0_1(.dout(w_dff_A_KEF28kuZ3_1),.din(w_dff_A_VlnhQV3B0_1),.clk(gclk));
	jdff dff_A_4g6tQ1Jv2_1(.dout(w_dff_A_VlnhQV3B0_1),.din(w_dff_A_4g6tQ1Jv2_1),.clk(gclk));
	jdff dff_A_UkQF1isM7_1(.dout(w_dff_A_4g6tQ1Jv2_1),.din(w_dff_A_UkQF1isM7_1),.clk(gclk));
	jdff dff_A_CoyOhJqe6_1(.dout(w_dff_A_UkQF1isM7_1),.din(w_dff_A_CoyOhJqe6_1),.clk(gclk));
	jdff dff_A_Wp6m8flR3_1(.dout(w_dff_A_CoyOhJqe6_1),.din(w_dff_A_Wp6m8flR3_1),.clk(gclk));
	jdff dff_A_vzdET3bI2_1(.dout(w_dff_A_Wp6m8flR3_1),.din(w_dff_A_vzdET3bI2_1),.clk(gclk));
	jdff dff_A_UpkpSmaE9_2(.dout(w_dff_A_FU6nqaMn8_0),.din(w_dff_A_UpkpSmaE9_2),.clk(gclk));
	jdff dff_A_FU6nqaMn8_0(.dout(w_dff_A_ZURtT3z48_0),.din(w_dff_A_FU6nqaMn8_0),.clk(gclk));
	jdff dff_A_ZURtT3z48_0(.dout(w_dff_A_yWwXl4Ia8_0),.din(w_dff_A_ZURtT3z48_0),.clk(gclk));
	jdff dff_A_yWwXl4Ia8_0(.dout(w_dff_A_5KR7nyzA4_0),.din(w_dff_A_yWwXl4Ia8_0),.clk(gclk));
	jdff dff_A_5KR7nyzA4_0(.dout(w_dff_A_TrpIRjTs6_0),.din(w_dff_A_5KR7nyzA4_0),.clk(gclk));
	jdff dff_A_TrpIRjTs6_0(.dout(w_dff_A_IH2i5YbZ3_0),.din(w_dff_A_TrpIRjTs6_0),.clk(gclk));
	jdff dff_A_IH2i5YbZ3_0(.dout(w_dff_A_ojReUlWs0_0),.din(w_dff_A_IH2i5YbZ3_0),.clk(gclk));
	jdff dff_A_ojReUlWs0_0(.dout(w_dff_A_36M7VTwQ0_0),.din(w_dff_A_ojReUlWs0_0),.clk(gclk));
	jdff dff_A_36M7VTwQ0_0(.dout(w_dff_A_6GJIz99K7_0),.din(w_dff_A_36M7VTwQ0_0),.clk(gclk));
	jdff dff_A_6GJIz99K7_0(.dout(w_dff_A_g0bsMIUw6_0),.din(w_dff_A_6GJIz99K7_0),.clk(gclk));
	jdff dff_A_g0bsMIUw6_0(.dout(w_dff_A_NBxdbV2b0_0),.din(w_dff_A_g0bsMIUw6_0),.clk(gclk));
	jdff dff_A_NBxdbV2b0_0(.dout(w_dff_A_LJAVZiyt7_0),.din(w_dff_A_NBxdbV2b0_0),.clk(gclk));
	jdff dff_A_LJAVZiyt7_0(.dout(w_dff_A_mCfbOrl39_0),.din(w_dff_A_LJAVZiyt7_0),.clk(gclk));
	jdff dff_A_mCfbOrl39_0(.dout(w_dff_A_LnD9suQ63_0),.din(w_dff_A_mCfbOrl39_0),.clk(gclk));
	jdff dff_A_LnD9suQ63_0(.dout(w_dff_A_Pp9RYpVK6_0),.din(w_dff_A_LnD9suQ63_0),.clk(gclk));
	jdff dff_A_Pp9RYpVK6_0(.dout(w_dff_A_cpRx40lW9_0),.din(w_dff_A_Pp9RYpVK6_0),.clk(gclk));
	jdff dff_A_cpRx40lW9_0(.dout(w_dff_A_BYjuNU6O1_0),.din(w_dff_A_cpRx40lW9_0),.clk(gclk));
	jdff dff_A_BYjuNU6O1_0(.dout(w_dff_A_HiA6zjCe3_0),.din(w_dff_A_BYjuNU6O1_0),.clk(gclk));
	jdff dff_A_HiA6zjCe3_0(.dout(w_dff_A_jHFVsp219_0),.din(w_dff_A_HiA6zjCe3_0),.clk(gclk));
	jdff dff_A_jHFVsp219_0(.dout(G223gat),.din(w_dff_A_jHFVsp219_0),.clk(gclk));
	jdff dff_A_Bu8Xx7qr6_1(.dout(w_dff_A_z0cbYEHf0_0),.din(w_dff_A_Bu8Xx7qr6_1),.clk(gclk));
	jdff dff_A_z0cbYEHf0_0(.dout(w_dff_A_icsYvCzl6_0),.din(w_dff_A_z0cbYEHf0_0),.clk(gclk));
	jdff dff_A_icsYvCzl6_0(.dout(w_dff_A_SbCTtuPm8_0),.din(w_dff_A_icsYvCzl6_0),.clk(gclk));
	jdff dff_A_SbCTtuPm8_0(.dout(w_dff_A_TCDSmcrq1_0),.din(w_dff_A_SbCTtuPm8_0),.clk(gclk));
	jdff dff_A_TCDSmcrq1_0(.dout(w_dff_A_2SlUWncV3_0),.din(w_dff_A_TCDSmcrq1_0),.clk(gclk));
	jdff dff_A_2SlUWncV3_0(.dout(w_dff_A_7bG7OGGA5_0),.din(w_dff_A_2SlUWncV3_0),.clk(gclk));
	jdff dff_A_7bG7OGGA5_0(.dout(w_dff_A_wy2ulCCa7_0),.din(w_dff_A_7bG7OGGA5_0),.clk(gclk));
	jdff dff_A_wy2ulCCa7_0(.dout(w_dff_A_G5HuG4MA3_0),.din(w_dff_A_wy2ulCCa7_0),.clk(gclk));
	jdff dff_A_G5HuG4MA3_0(.dout(w_dff_A_BD5BVYR26_0),.din(w_dff_A_G5HuG4MA3_0),.clk(gclk));
	jdff dff_A_BD5BVYR26_0(.dout(w_dff_A_a1lcWSP85_0),.din(w_dff_A_BD5BVYR26_0),.clk(gclk));
	jdff dff_A_a1lcWSP85_0(.dout(w_dff_A_cJDUwa1p0_0),.din(w_dff_A_a1lcWSP85_0),.clk(gclk));
	jdff dff_A_cJDUwa1p0_0(.dout(w_dff_A_Ogb9wPl73_0),.din(w_dff_A_cJDUwa1p0_0),.clk(gclk));
	jdff dff_A_Ogb9wPl73_0(.dout(G329gat),.din(w_dff_A_Ogb9wPl73_0),.clk(gclk));
	jdff dff_A_LssHnvSR5_1(.dout(w_dff_A_PgaZ1PXA1_0),.din(w_dff_A_LssHnvSR5_1),.clk(gclk));
	jdff dff_A_PgaZ1PXA1_0(.dout(w_dff_A_817POFMo8_0),.din(w_dff_A_PgaZ1PXA1_0),.clk(gclk));
	jdff dff_A_817POFMo8_0(.dout(w_dff_A_R5xiUOs84_0),.din(w_dff_A_817POFMo8_0),.clk(gclk));
	jdff dff_A_R5xiUOs84_0(.dout(w_dff_A_ZuERHQ0J4_0),.din(w_dff_A_R5xiUOs84_0),.clk(gclk));
	jdff dff_A_ZuERHQ0J4_0(.dout(w_dff_A_pOZByUTb2_0),.din(w_dff_A_ZuERHQ0J4_0),.clk(gclk));
	jdff dff_A_pOZByUTb2_0(.dout(G370gat),.din(w_dff_A_pOZByUTb2_0),.clk(gclk));
	jdff dff_A_vdAnjuUY2_1(.dout(w_dff_A_OmxKvbDF0_0),.din(w_dff_A_vdAnjuUY2_1),.clk(gclk));
	jdff dff_A_OmxKvbDF0_0(.dout(G430gat),.din(w_dff_A_OmxKvbDF0_0),.clk(gclk));
endmodule

