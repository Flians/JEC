/*

c5315:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jdff: 4692
	jand: 605
	jor: 419

Summary:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jdff: 4692
	jand: 605
	jor: 419
*/

module c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1157;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [1:0] w_G1_2;
	wire [2:0] w_G4_0;
	wire [1:0] w_G4_1;
	wire [1:0] w_G11_0;
	wire [1:0] w_G14_0;
	wire [1:0] w_G17_0;
	wire [1:0] w_G20_0;
	wire [1:0] w_G37_0;
	wire [1:0] w_G40_0;
	wire [1:0] w_G43_0;
	wire [1:0] w_G46_0;
	wire [1:0] w_G49_0;
	wire [1:0] w_G54_0;
	wire [1:0] w_G61_0;
	wire [1:0] w_G64_0;
	wire [1:0] w_G67_0;
	wire [1:0] w_G70_0;
	wire [1:0] w_G73_0;
	wire [1:0] w_G76_0;
	wire [1:0] w_G91_0;
	wire [1:0] w_G100_0;
	wire [1:0] w_G103_0;
	wire [1:0] w_G106_0;
	wire [1:0] w_G109_0;
	wire [1:0] w_G123_0;
	wire [1:0] w_G132_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G137_2;
	wire [2:0] w_G137_3;
	wire [2:0] w_G137_4;
	wire [2:0] w_G137_5;
	wire [2:0] w_G137_6;
	wire [2:0] w_G137_7;
	wire [2:0] w_G137_8;
	wire [1:0] w_G137_9;
	wire [2:0] w_G141_0;
	wire [2:0] w_G141_1;
	wire [2:0] w_G141_2;
	wire [1:0] w_G146_0;
	wire [1:0] w_G149_0;
	wire [1:0] w_G152_0;
	wire [1:0] w_G155_0;
	wire [1:0] w_G158_0;
	wire [1:0] w_G161_0;
	wire [1:0] w_G164_0;
	wire [1:0] w_G167_0;
	wire [1:0] w_G170_0;
	wire [1:0] w_G173_0;
	wire [1:0] w_G182_0;
	wire [1:0] w_G185_0;
	wire [1:0] w_G188_0;
	wire [1:0] w_G191_0;
	wire [1:0] w_G194_0;
	wire [1:0] w_G197_0;
	wire [1:0] w_G200_0;
	wire [1:0] w_G203_0;
	wire [2:0] w_G206_0;
	wire [2:0] w_G210_0;
	wire [2:0] w_G210_1;
	wire [2:0] w_G210_2;
	wire [2:0] w_G218_0;
	wire [2:0] w_G218_1;
	wire [2:0] w_G218_2;
	wire [2:0] w_G226_0;
	wire [2:0] w_G226_1;
	wire [2:0] w_G226_2;
	wire [2:0] w_G234_0;
	wire [2:0] w_G234_1;
	wire [1:0] w_G234_2;
	wire [2:0] w_G242_0;
	wire [2:0] w_G242_1;
	wire [1:0] w_G245_0;
	wire [2:0] w_G248_0;
	wire [2:0] w_G248_1;
	wire [2:0] w_G248_2;
	wire [2:0] w_G248_3;
	wire [2:0] w_G248_4;
	wire [1:0] w_G248_5;
	wire [2:0] w_G251_0;
	wire [2:0] w_G251_1;
	wire [2:0] w_G251_2;
	wire [2:0] w_G251_3;
	wire [2:0] w_G251_4;
	wire [2:0] w_G254_0;
	wire [2:0] w_G254_1;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [2:0] w_G257_2;
	wire [2:0] w_G265_0;
	wire [2:0] w_G265_1;
	wire [1:0] w_G265_2;
	wire [2:0] w_G273_0;
	wire [2:0] w_G273_1;
	wire [2:0] w_G273_2;
	wire [1:0] w_G280_0;
	wire [2:0] w_G281_0;
	wire [2:0] w_G281_1;
	wire [1:0] w_G281_2;
	wire [1:0] w_G289_0;
	wire [2:0] w_G293_0;
	wire [2:0] w_G299_0;
	wire [2:0] w_G302_0;
	wire [2:0] w_G308_0;
	wire [2:0] w_G308_1;
	wire [2:0] w_G316_0;
	wire [2:0] w_G316_1;
	wire [2:0] w_G324_0;
	wire [2:0] w_G324_1;
	wire [1:0] w_G331_0;
	wire [2:0] w_G332_0;
	wire [2:0] w_G332_1;
	wire [2:0] w_G332_2;
	wire [2:0] w_G332_3;
	wire [2:0] w_G332_4;
	wire [2:0] w_G335_0;
	wire [2:0] w_G335_1;
	wire [2:0] w_G335_2;
	wire [2:0] w_G335_3;
	wire [1:0] w_G335_4;
	wire [2:0] w_G341_0;
	wire [2:0] w_G341_1;
	wire [2:0] w_G341_2;
	wire [1:0] w_G348_0;
	wire [2:0] w_G351_0;
	wire [2:0] w_G351_1;
	wire [2:0] w_G351_2;
	wire [1:0] w_G358_0;
	wire [2:0] w_G361_0;
	wire [1:0] w_G369_0;
	wire [2:0] w_G374_0;
	wire [2:0] w_G389_0;
	wire [2:0] w_G400_0;
	wire [1:0] w_G400_1;
	wire [2:0] w_G411_0;
	wire [2:0] w_G422_0;
	wire [2:0] w_G422_1;
	wire [1:0] w_G422_2;
	wire [2:0] w_G435_0;
	wire [2:0] w_G435_1;
	wire [2:0] w_G446_0;
	wire [2:0] w_G446_1;
	wire [2:0] w_G457_0;
	wire [2:0] w_G457_1;
	wire [1:0] w_G457_2;
	wire [2:0] w_G468_0;
	wire [2:0] w_G468_1;
	wire [2:0] w_G479_0;
	wire [1:0] w_G479_1;
	wire [2:0] w_G490_0;
	wire [2:0] w_G490_1;
	wire [2:0] w_G503_0;
	wire [2:0] w_G503_1;
	wire [2:0] w_G514_0;
	wire [1:0] w_G514_1;
	wire [2:0] w_G523_0;
	wire [1:0] w_G523_1;
	wire [2:0] w_G534_0;
	wire [2:0] w_G534_1;
	wire [2:0] w_G545_0;
	wire [2:0] w_G549_0;
	wire [1:0] w_G552_0;
	wire [1:0] w_G559_0;
	wire [1:0] w_G562_0;
	wire [2:0] w_G1497_0;
	wire [2:0] w_G1689_0;
	wire [2:0] w_G1690_0;
	wire [2:0] w_G1691_0;
	wire [2:0] w_G1694_0;
	wire [2:0] w_G2174_0;
	wire [2:0] w_G2358_0;
	wire [2:0] w_G2358_1;
	wire [2:0] w_G2358_2;
	wire [1:0] w_G3173_0;
	wire [2:0] w_G3546_0;
	wire [2:0] w_G3546_1;
	wire [2:0] w_G3546_2;
	wire [2:0] w_G3546_3;
	wire [2:0] w_G3546_4;
	wire [1:0] w_G3546_5;
	wire [2:0] w_G3548_0;
	wire [2:0] w_G3548_1;
	wire [2:0] w_G3548_2;
	wire [2:0] w_G3548_3;
	wire [2:0] w_G3548_4;
	wire [1:0] w_G3552_0;
	wire [1:0] w_G3717_0;
	wire [2:0] w_G3724_0;
	wire [2:0] w_G4087_0;
	wire [2:0] w_G4088_0;
	wire [2:0] w_G4089_0;
	wire [2:0] w_G4090_0;
	wire [2:0] w_G4091_0;
	wire [2:0] w_G4091_1;
	wire [2:0] w_G4091_2;
	wire [2:0] w_G4092_0;
	wire [2:0] w_G4092_1;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G600_0;
	wire G600_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G611_0;
	wire G611_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire [2:0] w_G809_0;
	wire [2:0] w_G809_1;
	wire [2:0] w_G809_2;
	wire [1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G1000_0;
	wire G1000_fa_;
	wire w_G826_0;
	wire G826_fa_;
	wire w_G828_0;
	wire G828_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G867_0;
	wire G867_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire [1:0] w_n316_0;
	wire [1:0] w_n318_0;
	wire [2:0] w_n326_0;
	wire [2:0] w_n326_1;
	wire [1:0] w_n326_2;
	wire [1:0] w_n333_0;
	wire [1:0] w_n336_0;
	wire [1:0] w_n360_0;
	wire [1:0] w_n362_0;
	wire [2:0] w_n366_0;
	wire [2:0] w_n366_1;
	wire [2:0] w_n366_2;
	wire [2:0] w_n366_3;
	wire [2:0] w_n366_4;
	wire [2:0] w_n368_0;
	wire [2:0] w_n368_1;
	wire [2:0] w_n368_2;
	wire [2:0] w_n368_3;
	wire [2:0] w_n368_4;
	wire [1:0] w_n368_5;
	wire [2:0] w_n372_0;
	wire [1:0] w_n373_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n385_0;
	wire [2:0] w_n385_1;
	wire [2:0] w_n386_0;
	wire [2:0] w_n386_1;
	wire [2:0] w_n386_2;
	wire [2:0] w_n386_3;
	wire [2:0] w_n386_4;
	wire [2:0] w_n388_0;
	wire [2:0] w_n388_1;
	wire [2:0] w_n389_0;
	wire [2:0] w_n389_1;
	wire [2:0] w_n389_2;
	wire [2:0] w_n389_3;
	wire [2:0] w_n389_4;
	wire [1:0] w_n397_0;
	wire [2:0] w_n398_0;
	wire [2:0] w_n401_0;
	wire [2:0] w_n402_0;
	wire [2:0] w_n402_1;
	wire [1:0] w_n402_2;
	wire [1:0] w_n403_0;
	wire [2:0] w_n405_0;
	wire [2:0] w_n405_1;
	wire [1:0] w_n405_2;
	wire [1:0] w_n407_0;
	wire [1:0] w_n408_0;
	wire [2:0] w_n410_0;
	wire [1:0] w_n410_1;
	wire [1:0] w_n414_0;
	wire [1:0] w_n416_0;
	wire [2:0] w_n419_0;
	wire [2:0] w_n424_0;
	wire [2:0] w_n424_1;
	wire [1:0] w_n424_2;
	wire [1:0] w_n426_0;
	wire [1:0] w_n434_0;
	wire [2:0] w_n435_0;
	wire [2:0] w_n435_1;
	wire [2:0] w_n437_0;
	wire [2:0] w_n437_1;
	wire [1:0] w_n445_0;
	wire [2:0] w_n449_0;
	wire [2:0] w_n449_1;
	wire [2:0] w_n451_0;
	wire [1:0] w_n451_1;
	wire [1:0] w_n459_0;
	wire [2:0] w_n460_0;
	wire [2:0] w_n460_1;
	wire [2:0] w_n462_0;
	wire [1:0] w_n470_0;
	wire [2:0] w_n471_0;
	wire [1:0] w_n471_1;
	wire [2:0] w_n473_0;
	wire [2:0] w_n473_1;
	wire [1:0] w_n481_0;
	wire [2:0] w_n484_0;
	wire [1:0] w_n484_1;
	wire [2:0] w_n486_0;
	wire [1:0] w_n486_1;
	wire [1:0] w_n494_0;
	wire [2:0] w_n495_0;
	wire [2:0] w_n495_1;
	wire [2:0] w_n497_0;
	wire [1:0] w_n497_1;
	wire [1:0] w_n505_0;
	wire [2:0] w_n507_0;
	wire [1:0] w_n507_1;
	wire [1:0] w_n509_0;
	wire [1:0] w_n517_0;
	wire [2:0] w_n518_0;
	wire [1:0] w_n518_1;
	wire [2:0] w_n528_0;
	wire [2:0] w_n530_0;
	wire [1:0] w_n530_1;
	wire [1:0] w_n532_0;
	wire [1:0] w_n540_0;
	wire [2:0] w_n541_0;
	wire [1:0] w_n541_1;
	wire [1:0] w_n543_0;
	wire [1:0] w_n551_0;
	wire [2:0] w_n556_0;
	wire [2:0] w_n556_1;
	wire [2:0] w_n556_2;
	wire [2:0] w_n556_3;
	wire [2:0] w_n556_4;
	wire [1:0] w_n556_5;
	wire [2:0] w_n560_0;
	wire [1:0] w_n560_1;
	wire [2:0] w_n561_0;
	wire [1:0] w_n562_0;
	wire [2:0] w_n566_0;
	wire [2:0] w_n567_0;
	wire [1:0] w_n567_1;
	wire [1:0] w_n569_0;
	wire [1:0] w_n570_0;
	wire [2:0] w_n571_0;
	wire [1:0] w_n571_1;
	wire [2:0] w_n572_0;
	wire [2:0] w_n574_0;
	wire [2:0] w_n577_0;
	wire [2:0] w_n578_0;
	wire [2:0] w_n582_0;
	wire [1:0] w_n582_1;
	wire [2:0] w_n583_0;
	wire [1:0] w_n583_1;
	wire [1:0] w_n585_0;
	wire [2:0] w_n587_0;
	wire [1:0] w_n587_1;
	wire [2:0] w_n590_0;
	wire [1:0] w_n590_1;
	wire [1:0] w_n591_0;
	wire [2:0] w_n595_0;
	wire [1:0] w_n595_1;
	wire [2:0] w_n596_0;
	wire [2:0] w_n600_0;
	wire [1:0] w_n600_1;
	wire [1:0] w_n601_0;
	wire [2:0] w_n604_0;
	wire [2:0] w_n605_0;
	wire [2:0] w_n605_1;
	wire [2:0] w_n605_2;
	wire [2:0] w_n607_0;
	wire [2:0] w_n609_0;
	wire [2:0] w_n609_1;
	wire [2:0] w_n609_2;
	wire [2:0] w_n609_3;
	wire [2:0] w_n609_4;
	wire [2:0] w_n609_5;
	wire [2:0] w_n613_0;
	wire [2:0] w_n614_0;
	wire [2:0] w_n614_1;
	wire [1:0] w_n614_2;
	wire [2:0] w_n617_0;
	wire [1:0] w_n617_1;
	wire [2:0] w_n618_0;
	wire [1:0] w_n618_1;
	wire [2:0] w_n621_0;
	wire [2:0] w_n621_1;
	wire [1:0] w_n621_2;
	wire [2:0] w_n622_0;
	wire [1:0] w_n622_1;
	wire [1:0] w_n623_0;
	wire [2:0] w_n624_0;
	wire [2:0] w_n624_1;
	wire [2:0] w_n625_0;
	wire [2:0] w_n628_0;
	wire [2:0] w_n629_0;
	wire [1:0] w_n631_0;
	wire [2:0] w_n633_0;
	wire [1:0] w_n633_1;
	wire [2:0] w_n636_0;
	wire [1:0] w_n636_1;
	wire [2:0] w_n640_0;
	wire [2:0] w_n640_1;
	wire [1:0] w_n641_0;
	wire [1:0] w_n642_0;
	wire [2:0] w_n645_0;
	wire [2:0] w_n646_0;
	wire [2:0] w_n649_0;
	wire [1:0] w_n649_1;
	wire [1:0] w_n650_0;
	wire [2:0] w_n651_0;
	wire [1:0] w_n651_1;
	wire [1:0] w_n652_0;
	wire [1:0] w_n661_0;
	wire [1:0] w_n671_0;
	wire [1:0] w_n677_0;
	wire [1:0] w_n678_0;
	wire [1:0] w_n679_0;
	wire [1:0] w_n680_0;
	wire [2:0] w_n681_0;
	wire [2:0] w_n681_1;
	wire [1:0] w_n681_2;
	wire [1:0] w_n682_0;
	wire [2:0] w_n687_0;
	wire [1:0] w_n689_0;
	wire [2:0] w_n691_0;
	wire [2:0] w_n693_0;
	wire [2:0] w_n696_0;
	wire [1:0] w_n697_0;
	wire [1:0] w_n700_0;
	wire [1:0] w_n702_0;
	wire [2:0] w_n703_0;
	wire [1:0] w_n705_0;
	wire [1:0] w_n706_0;
	wire [2:0] w_n707_0;
	wire [1:0] w_n709_0;
	wire [1:0] w_n716_0;
	wire [2:0] w_n717_0;
	wire [1:0] w_n720_0;
	wire [2:0] w_n721_0;
	wire [1:0] w_n723_0;
	wire [1:0] w_n726_0;
	wire [2:0] w_n727_0;
	wire [2:0] w_n729_0;
	wire [1:0] w_n729_1;
	wire [2:0] w_n732_0;
	wire [1:0] w_n733_0;
	wire [1:0] w_n735_0;
	wire [1:0] w_n736_0;
	wire [2:0] w_n739_0;
	wire [1:0] w_n739_1;
	wire [1:0] w_n740_0;
	wire [1:0] w_n741_0;
	wire [1:0] w_n742_0;
	wire [2:0] w_n744_0;
	wire [2:0] w_n744_1;
	wire [2:0] w_n746_0;
	wire [2:0] w_n746_1;
	wire [2:0] w_n747_0;
	wire [2:0] w_n747_1;
	wire [2:0] w_n747_2;
	wire [2:0] w_n747_3;
	wire [2:0] w_n748_0;
	wire [2:0] w_n748_1;
	wire [2:0] w_n748_2;
	wire [2:0] w_n748_3;
	wire [1:0] w_n748_4;
	wire [2:0] w_n750_0;
	wire [1:0] w_n750_1;
	wire [2:0] w_n751_0;
	wire [2:0] w_n751_1;
	wire [1:0] w_n751_2;
	wire [2:0] w_n753_0;
	wire [2:0] w_n753_1;
	wire [2:0] w_n753_2;
	wire [2:0] w_n753_3;
	wire [2:0] w_n753_4;
	wire [2:0] w_n753_5;
	wire [2:0] w_n753_6;
	wire [2:0] w_n753_7;
	wire [1:0] w_n753_8;
	wire [1:0] w_n759_0;
	wire [1:0] w_n760_0;
	wire [1:0] w_n761_0;
	wire [2:0] w_n765_0;
	wire [2:0] w_n765_1;
	wire [2:0] w_n765_2;
	wire [2:0] w_n765_3;
	wire [2:0] w_n765_4;
	wire [2:0] w_n765_5;
	wire [1:0] w_n771_0;
	wire [1:0] w_n779_0;
	wire [2:0] w_n781_0;
	wire [2:0] w_n783_0;
	wire [1:0] w_n783_1;
	wire [1:0] w_n786_0;
	wire [1:0] w_n787_0;
	wire [2:0] w_n789_0;
	wire [2:0] w_n791_0;
	wire [1:0] w_n791_1;
	wire [1:0] w_n792_0;
	wire [2:0] w_n793_0;
	wire [2:0] w_n793_1;
	wire [2:0] w_n793_2;
	wire [2:0] w_n793_3;
	wire [1:0] w_n793_4;
	wire [2:0] w_n795_0;
	wire [1:0] w_n795_1;
	wire [1:0] w_n796_0;
	wire [2:0] w_n797_0;
	wire [2:0] w_n797_1;
	wire [2:0] w_n797_2;
	wire [2:0] w_n797_3;
	wire [1:0] w_n797_4;
	wire [2:0] w_n799_0;
	wire [2:0] w_n799_1;
	wire [2:0] w_n799_2;
	wire [2:0] w_n799_3;
	wire [1:0] w_n799_4;
	wire [2:0] w_n801_0;
	wire [2:0] w_n801_1;
	wire [2:0] w_n801_2;
	wire [2:0] w_n801_3;
	wire [1:0] w_n801_4;
	wire [2:0] w_n806_0;
	wire [1:0] w_n809_0;
	wire [1:0] w_n819_0;
	wire [1:0] w_n821_0;
	wire [2:0] w_n828_0;
	wire [1:0] w_n829_0;
	wire [1:0] w_n832_0;
	wire [1:0] w_n839_0;
	wire [2:0] w_n840_0;
	wire [2:0] w_n840_1;
	wire [2:0] w_n840_2;
	wire [2:0] w_n840_3;
	wire [1:0] w_n840_4;
	wire [1:0] w_n842_0;
	wire [2:0] w_n843_0;
	wire [2:0] w_n843_1;
	wire [2:0] w_n843_2;
	wire [2:0] w_n843_3;
	wire [1:0] w_n843_4;
	wire [2:0] w_n845_0;
	wire [2:0] w_n845_1;
	wire [2:0] w_n845_2;
	wire [2:0] w_n845_3;
	wire [1:0] w_n845_4;
	wire [2:0] w_n847_0;
	wire [2:0] w_n847_1;
	wire [2:0] w_n847_2;
	wire [2:0] w_n847_3;
	wire [1:0] w_n847_4;
	wire [1:0] w_n853_0;
	wire [1:0] w_n855_0;
	wire [1:0] w_n856_0;
	wire [1:0] w_n857_0;
	wire [1:0] w_n859_0;
	wire [1:0] w_n862_0;
	wire [1:0] w_n869_0;
	wire [1:0] w_n877_0;
	wire [1:0] w_n879_0;
	wire [1:0] w_n881_0;
	wire [1:0] w_n892_0;
	wire [1:0] w_n914_0;
	wire [1:0] w_n928_0;
	wire [2:0] w_n930_0;
	wire [1:0] w_n932_0;
	wire [2:0] w_n936_0;
	wire [1:0] w_n938_0;
	wire [1:0] w_n941_0;
	wire [1:0] w_n943_0;
	wire [1:0] w_n944_0;
	wire [1:0] w_n946_0;
	wire [2:0] w_n948_0;
	wire [1:0] w_n953_0;
	wire [1:0] w_n954_0;
	wire [1:0] w_n968_0;
	wire [1:0] w_n971_0;
	wire [1:0] w_n972_0;
	wire [1:0] w_n973_0;
	wire [1:0] w_n984_0;
	wire [2:0] w_n985_0;
	wire [2:0] w_n985_1;
	wire [2:0] w_n985_2;
	wire [2:0] w_n985_3;
	wire [1:0] w_n985_4;
	wire [1:0] w_n987_0;
	wire [2:0] w_n988_0;
	wire [2:0] w_n988_1;
	wire [2:0] w_n988_2;
	wire [2:0] w_n988_3;
	wire [1:0] w_n988_4;
	wire [2:0] w_n990_0;
	wire [2:0] w_n990_1;
	wire [2:0] w_n990_2;
	wire [2:0] w_n990_3;
	wire [1:0] w_n990_4;
	wire [2:0] w_n992_0;
	wire [2:0] w_n992_1;
	wire [2:0] w_n992_2;
	wire [2:0] w_n992_3;
	wire [1:0] w_n992_4;
	wire [1:0] w_n998_0;
	wire [2:0] w_n999_0;
	wire [2:0] w_n999_1;
	wire [2:0] w_n999_2;
	wire [2:0] w_n999_3;
	wire [1:0] w_n999_4;
	wire [1:0] w_n1001_0;
	wire [2:0] w_n1002_0;
	wire [2:0] w_n1002_1;
	wire [2:0] w_n1002_2;
	wire [2:0] w_n1002_3;
	wire [1:0] w_n1002_4;
	wire [2:0] w_n1004_0;
	wire [2:0] w_n1004_1;
	wire [2:0] w_n1004_2;
	wire [2:0] w_n1004_3;
	wire [1:0] w_n1004_4;
	wire [2:0] w_n1006_0;
	wire [2:0] w_n1006_1;
	wire [2:0] w_n1006_2;
	wire [2:0] w_n1006_3;
	wire [1:0] w_n1006_4;
	wire [2:0] w_n1012_0;
	wire [1:0] w_n1012_1;
	wire [2:0] w_n1014_0;
	wire [1:0] w_n1014_1;
	wire [2:0] w_n1021_0;
	wire [1:0] w_n1021_1;
	wire [2:0] w_n1023_0;
	wire [1:0] w_n1023_1;
	wire [2:0] w_n1030_0;
	wire [1:0] w_n1030_1;
	wire [2:0] w_n1032_0;
	wire [1:0] w_n1032_1;
	wire [2:0] w_n1039_0;
	wire [1:0] w_n1039_1;
	wire [2:0] w_n1041_0;
	wire [1:0] w_n1041_1;
	wire [1:0] w_n1142_0;
	wire [1:0] w_n1151_0;
	wire [2:0] w_n1163_0;
	wire [2:0] w_n1163_1;
	wire [2:0] w_n1197_0;
	wire [2:0] w_n1197_1;
	wire [2:0] w_n1205_0;
	wire [2:0] w_n1205_1;
	wire [2:0] w_n1235_0;
	wire [1:0] w_n1235_1;
	wire [2:0] w_n1242_0;
	wire [1:0] w_n1242_1;
	wire [2:0] w_n1244_0;
	wire [1:0] w_n1244_1;
	wire [2:0] w_n1251_0;
	wire [1:0] w_n1251_1;
	wire [2:0] w_n1253_0;
	wire [1:0] w_n1253_1;
	wire [1:0] w_n1358_0;
	wire [1:0] w_n1383_0;
	wire [1:0] w_n1391_0;
	wire [1:0] w_n1394_0;
	wire [1:0] w_n1398_0;
	wire [1:0] w_n1399_0;
	wire [1:0] w_n1409_0;
	wire [1:0] w_n1410_0;
	wire [1:0] w_n1411_0;
	wire [1:0] w_n1421_0;
	wire [1:0] w_n1425_0;
	wire [1:0] w_n1434_0;
	wire [1:0] w_n1438_0;
	wire [1:0] w_n1445_0;
	wire [1:0] w_n1446_0;
	wire [1:0] w_n1447_0;
	wire [1:0] w_n1452_0;
	wire [1:0] w_n1494_0;
	wire [1:0] w_n1533_0;
	wire [1:0] w_n1543_0;
	wire [1:0] w_n1545_0;
	wire [1:0] w_n1553_0;
	wire [1:0] w_n1555_0;
	wire [1:0] w_n1560_0;
	wire [1:0] w_n1568_0;
	wire [1:0] w_n1591_0;
	wire [1:0] w_n1597_0;
	wire [2:0] w_n1601_0;
	wire [1:0] w_n1602_0;
	wire [1:0] w_n1609_0;
	wire [1:0] w_n1610_0;
	wire [1:0] w_n1624_0;
	wire [1:0] w_n1629_0;
	wire [1:0] w_n1631_0;
	wire [1:0] w_n1634_0;
	wire w_dff_B_Id93cNMm3_1;
	wire w_dff_B_DSqho5bM5_0;
	wire w_dff_B_k7loCNst5_1;
	wire w_dff_B_gitFSkvp1_1;
	wire w_dff_B_iIiqK0wI0_2;
	wire w_dff_B_lCHdGDBG8_1;
	wire w_dff_B_3iwXC5Ze8_1;
	wire w_dff_B_WfzLEPFN3_0;
	wire w_dff_B_s29xw4Br7_1;
	wire w_dff_B_P9Y9rX433_1;
	wire w_dff_B_qQYrjorV2_0;
	wire w_dff_B_hA9gudFc2_1;
	wire w_dff_A_CPtyhCgc0_0;
	wire w_dff_A_dpaXL5n99_0;
	wire w_dff_A_77AqNmRZ4_0;
	wire w_dff_A_4jl8JVpv6_0;
	wire w_dff_A_WXVNPlky6_1;
	wire w_dff_A_muhFrUle4_1;
	wire w_dff_A_rRtH7eSm2_1;
	wire w_dff_A_7QRzfq9F4_1;
	wire w_dff_B_heedTL9O1_1;
	wire w_dff_B_inkwp1BG9_0;
	wire w_dff_B_dQvTcDHr1_1;
	wire w_dff_B_ovleiaxu5_1;
	wire w_dff_B_g5ylZoCc8_0;
	wire w_dff_B_dQxeAXvO7_1;
	wire w_dff_A_1ORJ7GLS6_0;
	wire w_dff_A_CMurshcQ6_1;
	wire w_dff_A_utxcD91K9_1;
	wire w_dff_A_12zpmsxd2_1;
	wire w_dff_A_eeMr8Due7_1;
	wire w_dff_A_Z5MG9Uvi3_1;
	wire w_dff_A_3DeliFwL5_2;
	wire w_dff_A_6n70IdMj6_2;
	wire w_dff_A_zLBQMaug5_2;
	wire w_dff_A_Ot0zYzPB2_2;
	wire w_dff_B_dk8GTSgy6_1;
	wire w_dff_B_FuxDKOSc6_1;
	wire w_dff_B_83XCQ04X6_0;
	wire w_dff_B_rTBel3Ui5_1;
	wire w_dff_B_fBBsNrfa9_1;
	wire w_dff_B_mEUW4q3f7_2;
	wire w_dff_B_EOZkHyo79_2;
	wire w_dff_B_wjOfmtcp1_2;
	wire w_dff_B_kq54St0X9_2;
	wire w_dff_B_e662TtVw6_1;
	wire w_dff_B_JbxfBhzd3_1;
	wire w_dff_B_acuTyYa16_1;
	wire w_dff_B_YYYGQkai2_1;
	wire w_dff_B_EkNSJ5Jv2_1;
	wire w_dff_B_p9mcHn1a3_1;
	wire w_dff_B_sQ1LnrdP9_1;
	wire w_dff_A_hmHkoDSJ2_1;
	wire w_dff_A_snnl1FyO3_1;
	wire w_dff_B_SDma8nWa1_3;
	wire w_dff_B_r4ed7AqC9_3;
	wire w_dff_B_7zdIdKpx6_3;
	wire w_dff_B_dI9q9fvR7_0;
	wire w_dff_B_XmCasODw0_2;
	wire w_dff_B_k4Ni3v0k9_2;
	wire w_dff_B_B2RShfql6_2;
	wire w_dff_B_AuYskGEF5_2;
	wire w_dff_B_3Mdt917A2_2;
	wire w_dff_A_584demJC4_0;
	wire w_dff_A_SO9kKnGd8_0;
	wire w_dff_A_3S8ZaUvv8_0;
	wire w_dff_A_F0FyPtwW1_0;
	wire w_dff_A_3qb3qbxk7_0;
	wire w_dff_A_bvaE7bz80_0;
	wire w_dff_B_6eEd5HAd3_0;
	wire w_dff_B_nPNkbsto3_0;
	wire w_dff_B_JJF1od7i7_0;
	wire w_dff_B_xGjOvOtH0_0;
	wire w_dff_B_mmIR7lIl0_0;
	wire w_dff_B_hOLlBpdr3_0;
	wire w_dff_B_hkTuO8SI5_0;
	wire w_dff_B_are00Gb59_0;
	wire w_dff_B_vBR5umxJ2_0;
	wire w_dff_B_PiEWqbwA4_0;
	wire w_dff_B_xNysK2R40_0;
	wire w_dff_B_tx0jMe6i2_0;
	wire w_dff_B_4HhBeV5W9_2;
	wire w_dff_B_nG3bsuQb7_2;
	wire w_dff_B_TTi3HKcw0_2;
	wire w_dff_B_bkgjFZb24_0;
	wire w_dff_B_5yVzVK379_0;
	wire w_dff_B_TcczeA249_0;
	wire w_dff_B_ndD6yr1S9_1;
	wire w_dff_B_y5H00sBe8_1;
	wire w_dff_B_SIf5AlHq5_1;
	wire w_dff_B_0C521gtF5_1;
	wire w_dff_B_raMBVX0g9_0;
	wire w_dff_B_tWjqZr2a1_0;
	wire w_dff_B_vcqIHBmT2_0;
	wire w_dff_B_ksLsfQMS2_0;
	wire w_dff_B_0G1dH7Rk3_0;
	wire w_dff_B_i6oJGg1L9_0;
	wire w_dff_B_eoOl4jo23_0;
	wire w_dff_B_xwx7QPtN4_0;
	wire w_dff_B_xinGAnSF1_0;
	wire w_dff_B_4099YKTg7_0;
	wire w_dff_B_Dp2fIXZN1_0;
	wire w_dff_B_THwIgXnc9_0;
	wire w_dff_B_KMwqRnSO9_0;
	wire w_dff_B_0YjR6u0w9_0;
	wire w_dff_B_W6kyvGYR7_0;
	wire w_dff_B_lkX286T74_0;
	wire w_dff_B_zQrjFDnb9_0;
	wire w_dff_B_UPcddqAS5_0;
	wire w_dff_B_TYlxeCwP3_2;
	wire w_dff_B_ycce6Lx65_2;
	wire w_dff_B_3lqw6BQP3_2;
	wire w_dff_B_chrVOFeU6_1;
	wire w_dff_B_9ZXX0n5X8_0;
	wire w_dff_B_81gYVq2G4_1;
	wire w_dff_B_EU7b06o62_1;
	wire w_dff_B_JgKebfju2_0;
	wire w_dff_B_9X5TAAfm0_0;
	wire w_dff_B_0Fmg88T65_1;
	wire w_dff_B_ippiVCQk1_1;
	wire w_dff_B_mvkwBMxs2_0;
	wire w_dff_B_ZwRsMymD1_1;
	wire w_dff_B_TJ0WxKdf1_0;
	wire w_dff_B_BEryW3mD9_0;
	wire w_dff_B_8kp36Tmz3_0;
	wire w_dff_B_cTT6ZgmG9_0;
	wire w_dff_B_fsMSFOzP9_0;
	wire w_dff_B_iLvON5Y48_0;
	wire w_dff_B_nEHltJjm0_0;
	wire w_dff_B_StdsBtGU2_0;
	wire w_dff_B_1nls4XEo9_0;
	wire w_dff_B_uSB73dQf4_0;
	wire w_dff_B_YJA3jG9g3_0;
	wire w_dff_B_lIOsDLVB3_0;
	wire w_dff_B_7oDXgmsj2_0;
	wire w_dff_B_tQiCExJB3_0;
	wire w_dff_A_siIh9YTQ4_0;
	wire w_dff_A_T9K8nkUe0_0;
	wire w_dff_A_NmzcGEOh0_0;
	wire w_dff_A_ZeZBAic30_0;
	wire w_dff_A_UffZVtVy7_0;
	wire w_dff_A_CtV7OBkU5_0;
	wire w_dff_A_4KOxYKIx5_0;
	wire w_dff_A_5pih1i2L9_0;
	wire w_dff_A_cM2ntAS04_0;
	wire w_dff_A_MPc2zuvu5_0;
	wire w_dff_A_lGXMKMcj6_0;
	wire w_dff_A_Nnrat7908_0;
	wire w_dff_A_n4Icl5t36_0;
	wire w_dff_A_XKe6QUf15_0;
	wire w_dff_A_DkCylNHW6_0;
	wire w_dff_B_S0KAFPTt1_0;
	wire w_dff_B_3noJ5F8U9_0;
	wire w_dff_B_DBiEtEMf6_0;
	wire w_dff_B_HdwOqerz1_0;
	wire w_dff_B_QcspVjQZ9_0;
	wire w_dff_B_XOJ1yKqR0_0;
	wire w_dff_B_fQ4IqU7U0_0;
	wire w_dff_B_lh8rfYao5_0;
	wire w_dff_B_SAB6UfdD7_0;
	wire w_dff_B_yOmprw5H3_0;
	wire w_dff_B_B2O0Sk7l4_0;
	wire w_dff_B_znZy9qvU2_0;
	wire w_dff_B_Qq9JiHcL5_0;
	wire w_dff_B_ffsg39Db4_0;
	wire w_dff_B_lcybjzNR4_0;
	wire w_dff_B_AAxLVVr25_0;
	wire w_dff_B_s8cdFx8V7_0;
	wire w_dff_B_yvaNLqw83_0;
	wire w_dff_B_SKYji9zI2_0;
	wire w_dff_B_jEQzjslZ4_0;
	wire w_dff_B_ALIeBAhq3_0;
	wire w_dff_B_UXPXI8BI6_0;
	wire w_dff_B_lcWxHoXi5_0;
	wire w_dff_B_WflnvAnp0_0;
	wire w_dff_B_NBbBKMGY2_0;
	wire w_dff_B_eQZuP0F98_0;
	wire w_dff_B_1dT86M9P1_0;
	wire w_dff_B_DrPeBPZ73_0;
	wire w_dff_B_CxP69g5l7_0;
	wire w_dff_B_ubqjtHnA6_0;
	wire w_dff_B_k5AHAt704_0;
	wire w_dff_B_DtlcdPho4_0;
	wire w_dff_B_6hnVM6k33_0;
	wire w_dff_A_b9DxND8P5_1;
	wire w_dff_A_GAy0RsyZ9_1;
	wire w_dff_A_i8BZwpIx3_2;
	wire w_dff_A_EzAR2vfD0_2;
	wire w_dff_A_gxRIdmRO6_2;
	wire w_dff_A_1vjksKh00_2;
	wire w_dff_A_3hxACZ724_1;
	wire w_dff_A_nA9xCYfF2_2;
	wire w_dff_A_Lfpu8aaD6_2;
	wire w_dff_B_VK4V7vCg1_0;
	wire w_dff_B_X84IcinJ8_0;
	wire w_dff_B_F0kYbrOg6_0;
	wire w_dff_B_2JmCzuXy8_0;
	wire w_dff_B_T7yu0DrN0_0;
	wire w_dff_B_megj8YUu7_0;
	wire w_dff_B_TwlMCvBa1_0;
	wire w_dff_B_Txm6iwGw9_0;
	wire w_dff_B_YCyunKXF5_0;
	wire w_dff_B_3EuztHLJ7_0;
	wire w_dff_B_SJhukanT5_0;
	wire w_dff_B_mZq6ymBp8_0;
	wire w_dff_B_KvchqE8I4_0;
	wire w_dff_B_YLKUDv2t1_0;
	wire w_dff_B_0QNOVFad6_2;
	wire w_dff_B_RaUeAJfS3_2;
	wire w_dff_B_lWeXAT4l1_2;
	wire w_dff_A_iEuz810I1_0;
	wire w_dff_A_j2DrEfx60_0;
	wire w_dff_A_xCZoYyqu2_0;
	wire w_dff_A_zoOfQhIk5_0;
	wire w_dff_A_GRzwZhCM5_0;
	wire w_dff_A_76G6ei0f1_0;
	wire w_dff_A_myzuL8GK8_0;
	wire w_dff_A_15d2twUx4_0;
	wire w_dff_A_r86EQqaE6_0;
	wire w_dff_A_RaPU5EZW3_0;
	wire w_dff_A_TpZCxc8j7_0;
	wire w_dff_A_dWmleysb5_0;
	wire w_dff_A_Rrfn7o2r5_0;
	wire w_dff_A_MRSr68jt7_0;
	wire w_dff_A_XDZ3xYaL9_0;
	wire w_dff_B_rOb8Gu7a6_0;
	wire w_dff_B_qsVRSY6K4_0;
	wire w_dff_B_c5OiLB299_0;
	wire w_dff_B_8uWItg6y1_0;
	wire w_dff_B_FFGeZrdd1_0;
	wire w_dff_B_qVawKd586_0;
	wire w_dff_B_0Uv407OR2_0;
	wire w_dff_B_nt38ReTw0_0;
	wire w_dff_B_ZvjbCkJz7_0;
	wire w_dff_B_skoIA8Hf5_0;
	wire w_dff_B_PBsKfb6g3_0;
	wire w_dff_B_QPJoRHpB9_0;
	wire w_dff_B_ZKONFJX52_2;
	wire w_dff_B_xKyJIKjB0_2;
	wire w_dff_B_mBRbiigd7_2;
	wire w_dff_B_PZl9L0Ym4_0;
	wire w_dff_B_KKLryKvr9_0;
	wire w_dff_B_zOylP07W0_0;
	wire w_dff_B_YrZPXZQH8_0;
	wire w_dff_B_gfrepL034_0;
	wire w_dff_B_PmFodKp56_0;
	wire w_dff_B_AnIR8f402_0;
	wire w_dff_B_U3vGkCaz8_0;
	wire w_dff_B_h6DRTrBX2_0;
	wire w_dff_B_eRBL8ZRO4_0;
	wire w_dff_B_rpkLrdoL7_0;
	wire w_dff_B_K4uE6dlT7_2;
	wire w_dff_B_S9df5jjs1_2;
	wire w_dff_B_xqM8Xbir9_2;
	wire w_dff_B_thv62NCx2_0;
	wire w_dff_B_ccpSNxHr2_0;
	wire w_dff_B_j39BeYFI8_0;
	wire w_dff_B_r3Vu4Yqw8_0;
	wire w_dff_B_9teD8Blt0_0;
	wire w_dff_B_uW1cntiw5_0;
	wire w_dff_B_fozBxNCC0_0;
	wire w_dff_B_tjLrggWN8_0;
	wire w_dff_B_NIVGXwuL9_0;
	wire w_dff_B_VVfb37309_0;
	wire w_dff_B_P4yay9r89_2;
	wire w_dff_B_w22BrIXB0_2;
	wire w_dff_B_IHXTYMqa1_2;
	wire w_dff_A_gmM4reVL0_1;
	wire w_dff_A_5mewilor6_1;
	wire w_dff_A_ste0IyhO2_2;
	wire w_dff_A_nx0IpDTI1_2;
	wire w_dff_A_DGHH2M3d7_2;
	wire w_dff_A_n7jGp1G37_2;
	wire w_dff_A_GYLz104K6_1;
	wire w_dff_A_rO3qYPbo2_2;
	wire w_dff_A_4wKiggY12_2;
	wire w_dff_B_Y2Zix5Sa1_0;
	wire w_dff_B_eHm6QLCe2_0;
	wire w_dff_B_KFhwNKMZ7_0;
	wire w_dff_B_XoJ6Wcqg3_0;
	wire w_dff_B_iIJeOkQ01_0;
	wire w_dff_B_ctWpjLVU2_0;
	wire w_dff_B_gg1U3cVV0_0;
	wire w_dff_B_Y7siAdOu4_0;
	wire w_dff_B_e7Cx7APb6_0;
	wire w_dff_B_8z9ikzWw8_0;
	wire w_dff_B_8N4MIl7e1_0;
	wire w_dff_B_Tdso8v7U5_0;
	wire w_dff_B_1Kt4iVGy4_0;
	wire w_dff_B_b2lq2Q2n7_0;
	wire w_dff_A_MyM5dgl37_0;
	wire w_dff_A_2tgNnHRA6_0;
	wire w_dff_A_LaueRLuW3_0;
	wire w_dff_A_wQu7aPfe9_0;
	wire w_dff_A_XjvKCxDn1_0;
	wire w_dff_A_F9YEEKZ20_0;
	wire w_dff_A_ZStwA7746_0;
	wire w_dff_A_7SgxEgOr4_0;
	wire w_dff_A_fo69tmbG0_0;
	wire w_dff_A_HbNzWxqy1_0;
	wire w_dff_A_0IuUq3qP9_0;
	wire w_dff_A_ykvi5NXc2_0;
	wire w_dff_A_ZrlNobvH1_0;
	wire w_dff_A_1EuSltka2_0;
	wire w_dff_A_XSyHe9qJ0_0;
	wire w_dff_B_dsAkIOls6_0;
	wire w_dff_B_iqL5QVgb3_0;
	wire w_dff_B_zYIkRZYU7_0;
	wire w_dff_B_pTcSqvVJ1_0;
	wire w_dff_B_ezoTYRWu4_0;
	wire w_dff_B_qwqwy70j8_0;
	wire w_dff_B_cD8QjL1l0_0;
	wire w_dff_B_5OMJYOqj2_0;
	wire w_dff_B_CWftwgeY8_0;
	wire w_dff_B_6OrtFTWs5_0;
	wire w_dff_B_d9CdKHzw7_0;
	wire w_dff_B_rfDhlykd3_0;
	wire w_dff_B_VtFPLDbu5_0;
	wire w_dff_B_ABtbWRYA3_0;
	wire w_dff_B_xpOAJV1S0_0;
	wire w_dff_B_oQue21gJ4_0;
	wire w_dff_B_gFJjeSU29_0;
	wire w_dff_B_fKMxE8QX4_0;
	wire w_dff_B_kwlxKjSu6_0;
	wire w_dff_B_YWU8t7go8_0;
	wire w_dff_B_76PEudjL8_0;
	wire w_dff_A_bwDk8wJS5_0;
	wire w_dff_A_y3mly7fF6_2;
	wire w_dff_A_CZH8B3ZO4_2;
	wire w_dff_A_dNH1hRh55_2;
	wire w_dff_A_c68Gy7OQ3_2;
	wire w_dff_B_oG0s388d4_0;
	wire w_dff_B_Re9gNGJE1_0;
	wire w_dff_B_fCmeMEMs2_0;
	wire w_dff_B_OtdQ3vFp6_0;
	wire w_dff_B_tadGsxag7_0;
	wire w_dff_B_gyA4NbWb8_0;
	wire w_dff_B_btZ3YHCc7_0;
	wire w_dff_B_vmAenznW3_0;
	wire w_dff_B_8GhYDpnR5_0;
	wire w_dff_B_2RcTZXdf2_0;
	wire w_dff_B_WAGQYCw72_0;
	wire w_dff_B_BrlY33gH4_0;
	wire w_dff_A_Edw0dPLH8_0;
	wire w_dff_A_1IpCWF9U5_0;
	wire w_dff_A_Dd6FveJz5_0;
	wire w_dff_A_ot3W3H814_0;
	wire w_dff_A_O4WcigL54_1;
	wire w_dff_A_FMUAtALP2_1;
	wire w_dff_A_GW5WSIsz3_0;
	wire w_dff_A_xRrmz9IE4_0;
	wire w_dff_A_f3xGREPE5_1;
	wire w_dff_B_SKrf3Cde8_0;
	wire w_dff_B_ST4Ndu5y9_0;
	wire w_dff_B_dP2IDRP77_0;
	wire w_dff_B_YkMBiu1n6_0;
	wire w_dff_B_U6Z4UY655_0;
	wire w_dff_B_rP59kVNh0_0;
	wire w_dff_B_gGfDCL4d3_0;
	wire w_dff_B_fyntxCTa5_0;
	wire w_dff_B_nDbgzLkI0_0;
	wire w_dff_B_9rKyvyJg0_0;
	wire w_dff_B_Vw92Ic3y1_0;
	wire w_dff_B_g7Khh2t65_0;
	wire w_dff_B_yTMNljsp9_0;
	wire w_dff_B_Q5CYsc8T9_0;
	wire w_dff_B_qpVakveK0_2;
	wire w_dff_B_3GXYxsTl9_2;
	wire w_dff_B_6uRl87Y29_2;
	wire w_dff_A_txp6AFKK4_0;
	wire w_dff_A_kPENjzXH4_0;
	wire w_dff_A_KCCsBxhm7_0;
	wire w_dff_A_TjNvWTAN0_0;
	wire w_dff_A_UYkLgkoW6_0;
	wire w_dff_A_7gxD2dLE5_0;
	wire w_dff_A_9f3ZTmi57_0;
	wire w_dff_B_p4yQhdvH5_0;
	wire w_dff_B_5bWTsV5t1_0;
	wire w_dff_B_y2nyBVQl7_0;
	wire w_dff_B_2MlRsDzR6_0;
	wire w_dff_B_zUbZh2AH1_0;
	wire w_dff_B_TAKE6U3t4_0;
	wire w_dff_B_ZgiS9Y6b0_0;
	wire w_dff_B_r8g0D6iJ3_0;
	wire w_dff_B_l5yiDbV36_1;
	wire w_dff_B_QJjsEbXt0_1;
	wire w_dff_B_6sGFwgL41_0;
	wire w_dff_B_fVsMa68i5_1;
	wire w_dff_A_fOleiBdk2_0;
	wire w_dff_A_y4LCp2Pi2_0;
	wire w_dff_A_FR3YClXm7_0;
	wire w_dff_A_dqmXt2a92_0;
	wire w_dff_A_QghXK8sy0_0;
	wire w_dff_A_PLgkUd441_0;
	wire w_dff_A_A8eDiGPQ8_0;
	wire w_dff_A_rhsUaOPN5_0;
	wire w_dff_B_CE2Vl1ea9_0;
	wire w_dff_B_DCAfXW7K4_0;
	wire w_dff_B_KHwbTEck1_0;
	wire w_dff_B_GGyalsZg4_0;
	wire w_dff_B_ogisMkkQ0_0;
	wire w_dff_B_g6X9K9FW6_0;
	wire w_dff_B_oZMF7rnb0_0;
	wire w_dff_B_MjeizViB9_0;
	wire w_dff_B_vxOFMEb27_0;
	wire w_dff_B_eQYXXswa6_0;
	wire w_dff_B_4mkfWb3v3_1;
	wire w_dff_B_25LjbvG77_1;
	wire w_dff_B_2SWRVRtF9_0;
	wire w_dff_B_RqnE4Ckq4_1;
	wire w_dff_B_4kYylFYj6_1;
	wire w_dff_B_AVJtX9VD2_1;
	wire w_dff_B_jlHZhAgo0_1;
	wire w_dff_B_0Aud0Oz35_1;
	wire w_dff_B_rhrXIeUF6_1;
	wire w_dff_B_EHwVUm3b2_1;
	wire w_dff_B_6MMxw6cE9_0;
	wire w_dff_B_JLQ03swz8_0;
	wire w_dff_B_naGe759P5_0;
	wire w_dff_B_TrWoTZwY8_0;
	wire w_dff_B_T0gOR15x1_0;
	wire w_dff_B_NvtaKItF0_0;
	wire w_dff_B_vXHoK1Bw5_0;
	wire w_dff_B_Q6aPBvyk1_0;
	wire w_dff_B_1waQ82K29_0;
	wire w_dff_B_0PbamN0N3_0;
	wire w_dff_B_Zkwko78p2_2;
	wire w_dff_B_2KqurAVh2_2;
	wire w_dff_B_9HPAWxIL1_2;
	wire w_dff_B_EQ4dCWyB1_0;
	wire w_dff_B_RNq2kfq04_0;
	wire w_dff_B_lXotI9so3_1;
	wire w_dff_B_H453Fxi78_1;
	wire w_dff_A_dmVkfCCc4_1;
	wire w_dff_B_uOWGZG217_0;
	wire w_dff_B_sMPIbE0P2_1;
	wire w_dff_A_TCaFfdVO2_0;
	wire w_dff_B_SCdRIpJo7_0;
	wire w_dff_B_6TiR4Avn9_0;
	wire w_dff_B_sglZAwff9_0;
	wire w_dff_B_sEKMPOcX8_0;
	wire w_dff_B_OJw71AoT6_0;
	wire w_dff_B_p60ZL6903_0;
	wire w_dff_B_0c9AXwHx1_1;
	wire w_dff_B_Dq5WLR2J7_1;
	wire w_dff_B_zpjQOf2U6_0;
	wire w_dff_B_cYahSXIn8_1;
	wire w_dff_B_FMmGyVGz9_0;
	wire w_dff_A_GltqHRr33_1;
	wire w_dff_A_cKMotMgo0_1;
	wire w_dff_A_lrYtObOH9_1;
	wire w_dff_A_D0fzhUMk0_1;
	wire w_dff_A_f4pgnVYu9_2;
	wire w_dff_A_QB56rGgY4_2;
	wire w_dff_A_kN0rlN7D8_0;
	wire w_dff_A_SQBn9wUY9_0;
	wire w_dff_A_vFivVuNl4_0;
	wire w_dff_A_inyEzEyT3_0;
	wire w_dff_A_UIGabkCu4_1;
	wire w_dff_A_QPr2FzPM5_1;
	wire w_dff_A_X1uiAiGC0_1;
	wire w_dff_A_e7EX4hop8_1;
	wire w_dff_B_s4pokhNX4_0;
	wire w_dff_B_IL8mvxNn9_0;
	wire w_dff_B_rUZ8gtx07_0;
	wire w_dff_B_rePXtQT82_0;
	wire w_dff_B_AbKNlnNx9_0;
	wire w_dff_B_v13gxwy20_0;
	wire w_dff_B_Z51mgOLi5_0;
	wire w_dff_B_Dpg5Z6Ou4_0;
	wire w_dff_B_0vdDPXmz7_0;
	wire w_dff_B_57rtjik33_0;
	wire w_dff_B_VTNitF7w1_0;
	wire w_dff_B_dOJaaTYT1_2;
	wire w_dff_B_uYTyBNBM2_2;
	wire w_dff_B_dOY9Sgmb6_2;
	wire w_dff_B_boAqdgSE9_0;
	wire w_dff_B_9lmp3lFb5_0;
	wire w_dff_B_2WmBJGSp0_0;
	wire w_dff_B_hQgBgHlP8_0;
	wire w_dff_B_ER99DSjI7_1;
	wire w_dff_B_iojmpH570_1;
	wire w_dff_B_XsQtfZjz4_0;
	wire w_dff_B_R1DgXB5Q0_1;
	wire w_dff_A_dQT0gd6k0_0;
	wire w_dff_A_HeInYmKg5_0;
	wire w_dff_A_TTCvWlQS7_0;
	wire w_dff_A_cWQZQc5t8_0;
	wire w_dff_A_7CWru7tZ0_0;
	wire w_dff_A_3JDVhz4W3_0;
	wire w_dff_B_k8hvkzF79_0;
	wire w_dff_B_hcmCq3ie7_0;
	wire w_dff_B_rRXoBqXY0_0;
	wire w_dff_B_mKbhzueB4_0;
	wire w_dff_B_U4YzXz4t6_0;
	wire w_dff_B_aXiWRMoZ0_0;
	wire w_dff_B_RSx2wWa70_0;
	wire w_dff_B_1WqIVF1L6_1;
	wire w_dff_B_AIEF4ijs8_1;
	wire w_dff_A_yEEkNlvz4_1;
	wire w_dff_B_Bojb8ccS4_0;
	wire w_dff_B_WBWgcu617_1;
	wire w_dff_B_03vhMbix5_0;
	wire w_dff_B_TVKhZIYw8_0;
	wire w_dff_B_sbx59ryn8_0;
	wire w_dff_B_Qd0dIKM25_0;
	wire w_dff_B_tMM8nhMj3_0;
	wire w_dff_B_IXxX6c2f0_0;
	wire w_dff_B_vuMNY9N62_0;
	wire w_dff_B_TFp41Crg5_0;
	wire w_dff_B_zMBaP8KC5_0;
	wire w_dff_B_YWk44sUP0_0;
	wire w_dff_B_hy53SsrT2_0;
	wire w_dff_B_vO706glE4_0;
	wire w_dff_B_6WCAemJ45_2;
	wire w_dff_B_kFVK53eQ7_2;
	wire w_dff_B_fm02c33D4_2;
	wire w_dff_A_iOZv9bvu4_0;
	wire w_dff_A_EhnspAGJ7_0;
	wire w_dff_A_dVVDTJGg2_0;
	wire w_dff_A_AO2Fb7lv2_0;
	wire w_dff_A_e7w3YjiL4_1;
	wire w_dff_A_GC7RmWww4_1;
	wire w_dff_B_OScALuvX8_0;
	wire w_dff_B_UwLl5j245_0;
	wire w_dff_B_M5SxCwSC1_0;
	wire w_dff_B_hiBEXKR64_0;
	wire w_dff_B_q7sIJVml5_0;
	wire w_dff_B_pWZ8gdsS9_0;
	wire w_dff_B_d6FpOrY91_1;
	wire w_dff_B_lNEbkQDY3_1;
	wire w_dff_B_qYhCDAB74_0;
	wire w_dff_B_I18ZZ34v1_1;
	wire w_dff_B_nfgQw7ht0_1;
	wire w_dff_B_9iog8XGt2_1;
	wire w_dff_B_YBI2nvkz0_1;
	wire w_dff_B_FMUbEqxb4_1;
	wire w_dff_A_hCMC9BxT9_2;
	wire w_dff_A_DcsFIBhn6_2;
	wire w_dff_A_adbeEL128_2;
	wire w_dff_A_XnJVWyVQ2_2;
	wire w_dff_B_XXhSP2CH3_3;
	wire w_dff_B_792OCErl1_3;
	wire w_dff_A_M0Pbx1Wj7_1;
	wire w_dff_A_tiltUMDh0_1;
	wire w_dff_A_4eAR3fuh0_2;
	wire w_dff_A_cLOTdFOI4_2;
	wire w_dff_A_i977vbLG0_2;
	wire w_dff_A_QBdu86M61_2;
	wire w_dff_A_MMJKujt49_0;
	wire w_dff_A_wxO2kF688_0;
	wire w_dff_A_fSFRTojg7_1;
	wire w_dff_B_q1g17QxW8_0;
	wire w_dff_B_6AJoBFaD1_0;
	wire w_dff_B_bIj9QglQ2_0;
	wire w_dff_B_NAjFVZ4G1_0;
	wire w_dff_B_LufNUIUy5_0;
	wire w_dff_B_zG0fkk6t3_0;
	wire w_dff_B_2nBctRa23_0;
	wire w_dff_B_7ZmmlJlu8_0;
	wire w_dff_B_IJoOo9HB6_1;
	wire w_dff_B_AiJ3oHxw6_1;
	wire w_dff_B_uuCq0Loz4_0;
	wire w_dff_B_hGD3gZm12_1;
	wire w_dff_B_utGnKuzG6_0;
	wire w_dff_A_1rR4Eh0M4_0;
	wire w_dff_A_6cgboUh24_0;
	wire w_dff_A_AALy9F1S9_0;
	wire w_dff_A_o1Ltpy1M8_0;
	wire w_dff_B_96mmDUl54_0;
	wire w_dff_B_UiKpCWv47_0;
	wire w_dff_B_jeIueljz0_0;
	wire w_dff_B_ipwJyREU9_0;
	wire w_dff_B_9QZPzyQ07_0;
	wire w_dff_B_eITe9ef42_0;
	wire w_dff_B_RoSOetZ70_0;
	wire w_dff_B_kY4Uz8h28_0;
	wire w_dff_B_NCuvBPCh0_0;
	wire w_dff_B_kPBmYc3V6_0;
	wire w_dff_B_U1ILsJjk4_0;
	wire w_dff_B_fONYaYHu7_0;
	wire w_dff_B_m3VQBE5F4_1;
	wire w_dff_B_4vJkQoic3_1;
	wire w_dff_B_fl9l574l5_1;
	wire w_dff_B_sEsIOO6B9_1;
	wire w_dff_B_VlWsDQyY4_1;
	wire w_dff_B_cAWCQ3GB5_1;
	wire w_dff_B_hnDtYCOQ2_0;
	wire w_dff_B_AYvu6gyr4_0;
	wire w_dff_B_kjfEXsjk7_0;
	wire w_dff_B_nMqtZAGB4_0;
	wire w_dff_B_ngeONwlG3_0;
	wire w_dff_B_TGmimn3W9_0;
	wire w_dff_B_dECqJNsv0_0;
	wire w_dff_B_Sg9wyukl9_0;
	wire w_dff_B_YamLtak89_0;
	wire w_dff_B_M3UGxdqe8_0;
	wire w_dff_B_3x5tHgxT4_0;
	wire w_dff_B_glttbpPm3_0;
	wire w_dff_B_LyayteW29_0;
	wire w_dff_B_Rye43WkJ3_0;
	wire w_dff_B_yC9Oqny89_0;
	wire w_dff_B_THKPYsQ40_0;
	wire w_dff_B_Fdj4RatZ1_1;
	wire w_dff_A_hKQYqhOv9_0;
	wire w_dff_A_ka9emVfG9_0;
	wire w_dff_A_uMQUu5Mt4_0;
	wire w_dff_A_zbAMO4ra6_0;
	wire w_dff_A_bBiesTm84_0;
	wire w_dff_A_7L3dMzNT2_0;
	wire w_dff_A_WcozmRnR8_0;
	wire w_dff_A_AcuIn80b5_0;
	wire w_dff_A_EpG7ZzI35_0;
	wire w_dff_A_uVAMcr3U1_0;
	wire w_dff_A_V5wPRyCH1_0;
	wire w_dff_A_EXwBExOx4_0;
	wire w_dff_A_8LXC2oEA5_2;
	wire w_dff_A_A5UoKsYg7_2;
	wire w_dff_A_wh9OqUnZ6_2;
	wire w_dff_A_WoXRAIiC4_2;
	wire w_dff_A_BN5s0OWO0_2;
	wire w_dff_A_QK6lzWmX6_2;
	wire w_dff_A_JbgB6ykI3_2;
	wire w_dff_A_OdBlXJcV2_2;
	wire w_dff_A_bJfjpC4g4_2;
	wire w_dff_A_fzJxdAU93_2;
	wire w_dff_A_k37QSIze9_2;
	wire w_dff_A_T2fBfKaU8_2;
	wire w_dff_A_RxAdn4vu3_2;
	wire w_dff_A_26IouIAS2_2;
	wire w_dff_A_0ilMfPlr6_2;
	wire w_dff_A_x8fElbcd4_2;
	wire w_dff_A_8jHWSEfk2_2;
	wire w_dff_A_4fATliDZ0_2;
	wire w_dff_A_y4bycuRs2_0;
	wire w_dff_A_Gal35TrV5_0;
	wire w_dff_A_EzOLEFkn2_0;
	wire w_dff_A_TFpmRgVb2_0;
	wire w_dff_A_hvaU3ANT8_0;
	wire w_dff_A_Bu5SEptC9_0;
	wire w_dff_A_jybOjyyD6_0;
	wire w_dff_A_KmaIF2qp6_0;
	wire w_dff_A_FRUcta711_0;
	wire w_dff_A_kvGKwaR46_0;
	wire w_dff_A_rE3kG1Y35_0;
	wire w_dff_A_kbfB5rmE9_0;
	wire w_dff_A_KPZKUBKl8_0;
	wire w_dff_B_8BN9JgJr4_2;
	wire w_dff_B_G0tIU59Z0_2;
	wire w_dff_B_nD7b9jDc3_2;
	wire w_dff_B_kEvZGrFN3_1;
	wire w_dff_B_vVo6NpYO0_0;
	wire w_dff_B_NIssC7zS7_0;
	wire w_dff_B_ZPdVBZ620_0;
	wire w_dff_A_hKPwJCt40_0;
	wire w_dff_B_omv28N7A3_1;
	wire w_dff_A_eGI5ioL92_0;
	wire w_dff_B_8xlMiN679_1;
	wire w_dff_B_UImnMwAf3_1;
	wire w_dff_B_53V4VH5V2_1;
	wire w_dff_B_Wzx6zhX68_1;
	wire w_dff_B_0kxmv4TN6_0;
	wire w_dff_B_zdUxXCoH5_1;
	wire w_dff_B_bNOwwZgX8_0;
	wire w_dff_A_OkzrOEWX9_0;
	wire w_dff_A_7UBBPQTy7_0;
	wire w_dff_A_Af7aqnpx1_0;
	wire w_dff_A_ZcjTCanV9_0;
	wire w_dff_B_Njv8LDIf3_0;
	wire w_dff_A_4T8SEnOh4_0;
	wire w_dff_B_5hsqcOvn3_0;
	wire w_dff_B_gnQGsW5I5_0;
	wire w_dff_B_khqqblDa1_0;
	wire w_dff_B_ciRoZKue4_0;
	wire w_dff_B_2xmnb8An4_0;
	wire w_dff_B_Z4vWh6kn7_0;
	wire w_dff_B_4PxaYOTQ7_0;
	wire w_dff_B_fptPdpyV5_0;
	wire w_dff_B_2UbHNWf24_0;
	wire w_dff_B_um3yBCOh7_0;
	wire w_dff_B_NSlHX2uf2_0;
	wire w_dff_B_cIQsVOIZ9_0;
	wire w_dff_B_Mu3dFL2x7_0;
	wire w_dff_B_s8tlO6rJ5_0;
	wire w_dff_B_oZvyQe5e2_0;
	wire w_dff_B_oq6JPoJK9_0;
	wire w_dff_B_fE20assw7_0;
	wire w_dff_B_QXWGfaW84_0;
	wire w_dff_B_F8m6nLQa7_0;
	wire w_dff_B_GQ0PLVdF9_0;
	wire w_dff_B_ntpr1OrJ8_0;
	wire w_dff_B_rrzqkxJX2_0;
	wire w_dff_B_UsKTbJOH2_0;
	wire w_dff_B_U57Tn4OJ6_0;
	wire w_dff_B_ygJarYfs0_0;
	wire w_dff_B_7UBwKGAW8_0;
	wire w_dff_B_nScdvI9E7_0;
	wire w_dff_B_zjTkoiaA0_0;
	wire w_dff_B_OcSfrWjB7_0;
	wire w_dff_B_k6dFFJ5d9_0;
	wire w_dff_B_eE9BHOiQ4_0;
	wire w_dff_B_Dperetc79_0;
	wire w_dff_B_qxKUMI2s8_0;
	wire w_dff_B_Z2kCsBUf6_0;
	wire w_dff_B_eUoyMdux2_0;
	wire w_dff_B_lrLLoZaM8_0;
	wire w_dff_B_UeAhgxOY3_2;
	wire w_dff_B_4zTjIPSx3_2;
	wire w_dff_B_KBen70oB1_2;
	wire w_dff_B_IJbKMdYW1_0;
	wire w_dff_B_LMt06rRg9_0;
	wire w_dff_B_UP1AnLUt5_0;
	wire w_dff_B_ELToS6ad7_0;
	wire w_dff_B_bZk81CwM9_0;
	wire w_dff_B_ofGUW5RS3_0;
	wire w_dff_B_1e2K5l962_0;
	wire w_dff_B_49xixjr13_0;
	wire w_dff_B_2Jrakhrj6_0;
	wire w_dff_B_p02BTYxB6_0;
	wire w_dff_B_YPMqT73X3_0;
	wire w_dff_B_7jP2SkIc2_0;
	wire w_dff_B_hvtHPjWP6_0;
	wire w_dff_B_0kRqpW4z8_0;
	wire w_dff_B_pa2Z2kjW5_0;
	wire w_dff_B_0JrtqFgk8_0;
	wire w_dff_B_Foucat1g1_0;
	wire w_dff_B_tyhcO2867_0;
	wire w_dff_B_oceMWlqv0_0;
	wire w_dff_B_xDaQlDmY9_0;
	wire w_dff_B_YihmyH3A4_0;
	wire w_dff_B_UmWlof7l5_0;
	wire w_dff_B_oqUcqDfa8_0;
	wire w_dff_B_3t7SR3Ek3_0;
	wire w_dff_B_neTNoa0G6_0;
	wire w_dff_B_qn2hLOcN9_0;
	wire w_dff_B_2okZtWdb2_0;
	wire w_dff_B_EgSggrT63_0;
	wire w_dff_B_jwmbYkEd7_0;
	wire w_dff_B_HXv8tPOX6_0;
	wire w_dff_B_fPpETqz82_0;
	wire w_dff_B_HaCTnfuG9_0;
	wire w_dff_B_qiaSDrf53_0;
	wire w_dff_B_3LcSg0uW3_0;
	wire w_dff_A_4KE5DLLY1_2;
	wire w_dff_A_DvvXWMSC4_2;
	wire w_dff_B_WvUzs1Ts3_0;
	wire w_dff_B_f2ZpQjlX1_0;
	wire w_dff_B_WejA4FLu8_0;
	wire w_dff_B_6YRv9iKj6_0;
	wire w_dff_B_wbheDars5_0;
	wire w_dff_B_oERyJoSr0_0;
	wire w_dff_B_BdTLhuto8_0;
	wire w_dff_B_7j6kMCPl8_0;
	wire w_dff_B_4I4tqIYh2_0;
	wire w_dff_B_VPFnzmRM6_0;
	wire w_dff_B_NMHZGI2e2_0;
	wire w_dff_B_SHPW11385_0;
	wire w_dff_B_x0tl3HEi2_0;
	wire w_dff_B_v0zLj5Od4_0;
	wire w_dff_B_1xKtCMCP1_0;
	wire w_dff_B_K4fKwws38_0;
	wire w_dff_B_LaUmfTSg0_0;
	wire w_dff_B_OWl8EKew6_0;
	wire w_dff_B_mOU4ExbL6_0;
	wire w_dff_B_zsL91hBh6_0;
	wire w_dff_B_WxKpJivV8_0;
	wire w_dff_B_8XrXzZY87_0;
	wire w_dff_B_AZqvnguG5_0;
	wire w_dff_B_eBZ5pvxp1_0;
	wire w_dff_B_ttVhzxHJ5_0;
	wire w_dff_B_QauO95Rq0_0;
	wire w_dff_B_qXkdGEae9_0;
	wire w_dff_B_efeCm2R40_0;
	wire w_dff_B_leDKtqH27_0;
	wire w_dff_B_h0OPKYgB1_0;
	wire w_dff_B_szqEZaur3_0;
	wire w_dff_B_HfR9NiRb5_0;
	wire w_dff_B_8DjwxO8J4_0;
	wire w_dff_B_LY7NLxU77_2;
	wire w_dff_B_7lNTWjgU2_2;
	wire w_dff_B_agihHWfT0_2;
	wire w_dff_B_Dsi6kEVv0_0;
	wire w_dff_B_caSoMYmE9_0;
	wire w_dff_B_6picSZTO7_0;
	wire w_dff_B_1WIk8esE8_0;
	wire w_dff_B_H6Ku1xD71_0;
	wire w_dff_B_KYqGTzkz7_0;
	wire w_dff_B_89eBLgjP3_0;
	wire w_dff_B_2YMC2gyN5_0;
	wire w_dff_B_CKx8PJfx1_0;
	wire w_dff_B_ZFAo4mrR0_0;
	wire w_dff_B_JvpU8GmB3_0;
	wire w_dff_B_GUVV8PFt9_0;
	wire w_dff_B_RZIRIXk37_0;
	wire w_dff_B_GZVaPspF7_0;
	wire w_dff_B_ILMNY9yM7_0;
	wire w_dff_B_jgcc0Xlp3_0;
	wire w_dff_B_p0dtSfDh5_0;
	wire w_dff_B_fJylF7gT3_2;
	wire w_dff_B_xZvxPhuO3_2;
	wire w_dff_B_o5pLiG8c7_2;
	wire w_dff_A_HPZV4S169_2;
	wire w_dff_A_JkQzaEnP2_2;
	wire w_dff_B_TlPbYDHg5_0;
	wire w_dff_B_VynV79Ea6_0;
	wire w_dff_B_SSIgrztB6_0;
	wire w_dff_B_UvqLAqdy1_0;
	wire w_dff_B_ssxuIrBs2_0;
	wire w_dff_B_U7oIt5kt7_0;
	wire w_dff_B_lfh1lHlH3_0;
	wire w_dff_B_ts0cGKd99_0;
	wire w_dff_B_J7em22F56_0;
	wire w_dff_B_fRMhin913_0;
	wire w_dff_B_paT4gHN20_0;
	wire w_dff_B_P1oVGmOm4_0;
	wire w_dff_B_mqNFGYbA8_0;
	wire w_dff_B_QWeznXfG3_0;
	wire w_dff_B_4ZPfSibY8_0;
	wire w_dff_B_2V4gCxYY5_0;
	wire w_dff_B_9XFcTKAY6_2;
	wire w_dff_B_d6P1H7FR3_2;
	wire w_dff_B_daimAzmN6_2;
	wire w_dff_B_bW8KinqO0_0;
	wire w_dff_B_iktnIL0L6_0;
	wire w_dff_B_M5BWNTpH4_0;
	wire w_dff_B_uYjMGAgs6_0;
	wire w_dff_B_QfF1cgp14_0;
	wire w_dff_B_j4yw23zc2_0;
	wire w_dff_B_HCPl31yi7_0;
	wire w_dff_B_YtYQyY3I9_0;
	wire w_dff_B_rHCZqgn79_0;
	wire w_dff_B_3SShvQfM7_0;
	wire w_dff_B_IU2UfoME2_0;
	wire w_dff_B_I9D5SnTh6_0;
	wire w_dff_B_PDGODrkG7_0;
	wire w_dff_B_jHhMLNMw5_0;
	wire w_dff_B_kCrwhqOF3_0;
	wire w_dff_B_CLS7VxaR5_0;
	wire w_dff_A_8LjImTsb6_0;
	wire w_dff_A_Le83ZYs52_0;
	wire w_dff_A_S2HGctti1_0;
	wire w_dff_A_oXqaLl9T1_0;
	wire w_dff_A_PNqV6Qcx1_0;
	wire w_dff_A_pQ3EGlQh9_1;
	wire w_dff_B_7sZ77vpw0_0;
	wire w_dff_B_gQVib5Ky2_0;
	wire w_dff_B_zDvvXsdD3_0;
	wire w_dff_B_3uUhCogx3_0;
	wire w_dff_B_6sKEyhKr3_0;
	wire w_dff_B_3XfNGyaC8_0;
	wire w_dff_B_m9Xf2G8T3_0;
	wire w_dff_B_TiFcmO2D4_0;
	wire w_dff_B_m0jBdFO43_0;
	wire w_dff_B_KL5axc5D2_0;
	wire w_dff_B_wdoOD40p2_0;
	wire w_dff_B_6H7XOcCL7_0;
	wire w_dff_B_LzblFryV0_0;
	wire w_dff_B_mi3BNH5X1_0;
	wire w_dff_B_QpuCc7aU9_0;
	wire w_dff_B_xkI0oTdo9_0;
	wire w_dff_B_wHs13Xsv8_0;
	wire w_dff_B_pqqzMUZl8_0;
	wire w_dff_B_eDGJMUsh1_0;
	wire w_dff_B_zDEWOE8r4_0;
	wire w_dff_B_ROW32n2Y7_0;
	wire w_dff_B_q9BTNHhf8_0;
	wire w_dff_B_kaE8LV7h8_0;
	wire w_dff_B_SzuDFWmC0_0;
	wire w_dff_B_kWLqNuTG3_0;
	wire w_dff_B_khNQBvbu6_0;
	wire w_dff_B_QnhusBw42_0;
	wire w_dff_B_6Og4tF8l2_0;
	wire w_dff_B_oyFq5PQM6_0;
	wire w_dff_B_f7rGyw7A4_0;
	wire w_dff_B_Qqyg0ppa1_0;
	wire w_dff_B_OQjliZDL7_0;
	wire w_dff_B_Gkx80q075_0;
	wire w_dff_B_2lnt7ZZc6_0;
	wire w_dff_A_jkwCsyvQ2_0;
	wire w_dff_A_ssvHqDnK6_1;
	wire w_dff_A_KOcAUxzg9_0;
	wire w_dff_A_VeVRreo87_1;
	wire w_dff_B_psgHtD3X4_0;
	wire w_dff_B_gxhjelfQ0_0;
	wire w_dff_B_4OjYtLMW3_0;
	wire w_dff_B_uF8pXqRS1_0;
	wire w_dff_B_lJKaaXEs2_0;
	wire w_dff_B_0kzx022p2_0;
	wire w_dff_B_KBWcRlxM8_0;
	wire w_dff_B_5HETUlqq4_0;
	wire w_dff_B_FqzyediK8_0;
	wire w_dff_B_DtjazNvV6_0;
	wire w_dff_B_IDd31ii58_0;
	wire w_dff_B_lhTzgnLZ5_0;
	wire w_dff_B_JafwXmKH7_0;
	wire w_dff_B_nC5DE3KI8_0;
	wire w_dff_B_KSjAw9yk3_0;
	wire w_dff_B_oE1JZ1uG7_0;
	wire w_dff_B_lClUUBK73_0;
	wire w_dff_B_oir3KOd09_0;
	wire w_dff_A_Q5iQULE34_0;
	wire w_dff_B_ACG9gMAr7_0;
	wire w_dff_B_qqXpbwvH5_0;
	wire w_dff_B_UBz4wztc2_0;
	wire w_dff_B_zqy8829E1_0;
	wire w_dff_B_yqPhX9sK0_0;
	wire w_dff_B_wNcDOGWv5_0;
	wire w_dff_B_88WzFsQN7_0;
	wire w_dff_B_6ERaSkNq8_0;
	wire w_dff_B_CegQKCXD2_0;
	wire w_dff_B_1G6AH4SC0_0;
	wire w_dff_B_WXtURZR96_0;
	wire w_dff_B_jJ2ZF4MG4_0;
	wire w_dff_B_QH3IzzPX0_0;
	wire w_dff_B_XoHIIzfZ5_0;
	wire w_dff_B_qNDrs8HS5_0;
	wire w_dff_B_hu36JLKP8_0;
	wire w_dff_B_Y9eZYFbZ9_2;
	wire w_dff_B_7JJA35wq4_2;
	wire w_dff_B_hUr9Tjjk0_2;
	wire w_dff_B_z4ZusqbI3_0;
	wire w_dff_B_SERaMATc5_0;
	wire w_dff_B_qQWxfnOR6_0;
	wire w_dff_B_6JgCC1x72_0;
	wire w_dff_B_SXznF4MS1_0;
	wire w_dff_B_y1AOhIBq7_0;
	wire w_dff_B_WYbBZJjj3_0;
	wire w_dff_B_FqOQgcdX0_0;
	wire w_dff_B_iJl25Ho34_0;
	wire w_dff_B_rjYRKcj64_0;
	wire w_dff_B_L7sOoYjC0_0;
	wire w_dff_B_vhl4Infz5_1;
	wire w_dff_B_X0uLgB6d7_1;
	wire w_dff_B_PwIGwvRL3_0;
	wire w_dff_B_1q36Kfhi6_0;
	wire w_dff_B_UNlSYR6n1_0;
	wire w_dff_B_DOuR6GSJ2_0;
	wire w_dff_B_LeaNdVMJ4_0;
	wire w_dff_B_GiLV8bMY9_0;
	wire w_dff_B_hUklCis55_0;
	wire w_dff_B_ox7P9IJy7_0;
	wire w_dff_B_x2KNZ6iI1_0;
	wire w_dff_B_IUk8gXyh9_0;
	wire w_dff_B_Jior3hBQ9_0;
	wire w_dff_B_7kBC6HHg6_0;
	wire w_dff_B_p4kYf6YZ4_1;
	wire w_dff_B_glA5B8U56_1;
	wire w_dff_B_bXdLyk5W1_0;
	wire w_dff_B_dYPgXtsD0_1;
	wire w_dff_B_IC0ps1fo6_0;
	wire w_dff_B_jq4fNhWr2_0;
	wire w_dff_B_cUqcTNe14_0;
	wire w_dff_B_PPDilmP60_0;
	wire w_dff_B_1StuuxkN7_0;
	wire w_dff_B_KIgBZSuJ3_0;
	wire w_dff_B_vbhBoZhC2_0;
	wire w_dff_B_U5vzV9CO5_0;
	wire w_dff_B_7ZOJJbIN4_0;
	wire w_dff_B_0gNvbhUZ2_0;
	wire w_dff_B_MQDLUuzm1_0;
	wire w_dff_B_iE3s2WX19_0;
	wire w_dff_B_36pvyGsG2_0;
	wire w_dff_B_IaAH95SD2_0;
	wire w_dff_B_jEhbxsjl3_0;
	wire w_dff_B_gjb4Oi0q0_0;
	wire w_dff_B_PVzDrUI07_0;
	wire w_dff_B_EOzGzui27_2;
	wire w_dff_B_i8SxsqYX0_2;
	wire w_dff_B_SKbHMiPW2_2;
	wire w_dff_B_PzwauFEn5_0;
	wire w_dff_B_T1WLndiE7_0;
	wire w_dff_B_wk2mTHoO6_0;
	wire w_dff_B_uftwXITn5_0;
	wire w_dff_B_Pprlg6Pk7_0;
	wire w_dff_B_z1rch9tb1_0;
	wire w_dff_B_iZHAJWmI6_0;
	wire w_dff_B_tFk35qCd0_0;
	wire w_dff_B_3Qy6W5L95_0;
	wire w_dff_B_hkmYepsr1_0;
	wire w_dff_B_IgMqFLy09_0;
	wire w_dff_B_ua2pDzep4_0;
	wire w_dff_B_JQ3weE2T6_1;
	wire w_dff_B_XSMluYwI5_1;
	wire w_dff_A_NuJTEUlq2_1;
	wire w_dff_B_RLn8NmTO6_1;
	wire w_dff_B_ko7vEbz17_1;
	wire w_dff_B_rTNjjYZQ2_1;
	wire w_dff_B_I6u7Xvyt7_1;
	wire w_dff_B_9awdeCEy5_1;
	wire w_dff_B_10FZb3Xe6_1;
	wire w_dff_B_1QTbg1t01_1;
	wire w_dff_B_DTEZEmzc3_1;
	wire w_dff_B_UsBq3o8C3_1;
	wire w_dff_B_gZZxHR9A9_1;
	wire w_dff_B_x4ipNBLy2_0;
	wire w_dff_B_G6R5a1ku6_0;
	wire w_dff_B_ydD3jYtZ2_0;
	wire w_dff_B_pcCgPbGV9_0;
	wire w_dff_B_d76h6jha4_0;
	wire w_dff_B_gjxnMQvY5_0;
	wire w_dff_B_XrZYz4ad6_0;
	wire w_dff_B_Tbt7paOx5_0;
	wire w_dff_B_rGvjwjYQ3_0;
	wire w_dff_B_XOIjbCTo2_0;
	wire w_dff_B_lC30vCYl0_0;
	wire w_dff_B_c3t1imLH3_0;
	wire w_dff_B_CFEHNOeE2_0;
	wire w_dff_B_APznchf67_1;
	wire w_dff_B_ZA4O3y686_1;
	wire w_dff_B_tG9adEFH1_0;
	wire w_dff_B_RjlglxQt3_1;
	wire w_dff_B_9hMU6lcc0_1;
	wire w_dff_B_AUupmtsm7_1;
	wire w_dff_B_HtxUaVVx9_1;
	wire w_dff_B_1C0tSIMy4_1;
	wire w_dff_B_HLW7vWet5_1;
	wire w_dff_B_XQIOUIOp3_1;
	wire w_dff_B_fv1ZyOmz0_1;
	wire w_dff_B_RfESNhlC1_1;
	wire w_dff_B_0hsauJ6R8_1;
	wire w_dff_B_gn54M3Ww9_1;
	wire w_dff_B_qPVtVFvi2_1;
	wire w_dff_B_IJW9hVqL8_1;
	wire w_dff_B_CC39pABg7_1;
	wire w_dff_B_MkVrTEoD9_1;
	wire w_dff_B_0H2DIDvE4_1;
	wire w_dff_B_lKxuVDm25_1;
	wire w_dff_B_S1QX8Zvs1_1;
	wire w_dff_B_ofUBp4UG4_1;
	wire w_dff_B_rRMNoTYZ7_1;
	wire w_dff_A_nWLaiN3j3_1;
	wire w_dff_A_RJa4Gq8s8_1;
	wire w_dff_A_MBuGZqLz6_1;
	wire w_dff_A_dhUJ9rvE6_1;
	wire w_dff_A_FilrnN435_1;
	wire w_dff_A_nahFt7xa8_1;
	wire w_dff_A_CqfnTfWi7_1;
	wire w_dff_A_anLfhxRS1_1;
	wire w_dff_A_Ogz8PFMW1_1;
	wire w_dff_A_HZjtsSJL1_1;
	wire w_dff_A_UhTU1Eae9_1;
	wire w_dff_A_PJayM3t63_1;
	wire w_dff_A_LgHOED8V7_1;
	wire w_dff_A_KXRjMjqW9_2;
	wire w_dff_A_dwuX4k8i2_2;
	wire w_dff_A_LTgyNi8J7_2;
	wire w_dff_A_JkOpa6Sh7_2;
	wire w_dff_A_eIOE29rS2_2;
	wire w_dff_A_fDzeVmLY4_2;
	wire w_dff_A_KudOem1w6_2;
	wire w_dff_A_TdZh7eaG9_2;
	wire w_dff_A_GBoCOpiM3_2;
	wire w_dff_A_MYgwYiWG7_2;
	wire w_dff_A_Fz0Ytbk11_2;
	wire w_dff_A_A5Gq2DXr3_2;
	wire w_dff_B_nkCdGZ7y3_0;
	wire w_dff_B_yCMt4mVz6_0;
	wire w_dff_B_QxcVWerE2_0;
	wire w_dff_B_YDjt6HPO6_0;
	wire w_dff_B_s29JAerm7_0;
	wire w_dff_B_kAboX37W9_0;
	wire w_dff_B_C8cMFetO5_0;
	wire w_dff_B_Lltmh7hF3_0;
	wire w_dff_B_JoVEzuEX1_0;
	wire w_dff_B_TGEMRHmX9_0;
	wire w_dff_B_ru1xUOcn8_0;
	wire w_dff_B_BNYDaigi9_0;
	wire w_dff_B_7jJuMPSE4_0;
	wire w_dff_B_pZZobhUw4_0;
	wire w_dff_B_tpSFld6Y9_0;
	wire w_dff_B_aAqwkRiN8_0;
	wire w_dff_B_E09Mezaa2_0;
	wire w_dff_B_CxepozI67_2;
	wire w_dff_B_klaNNE4T8_2;
	wire w_dff_B_lvXXY4k86_2;
	wire w_dff_B_Zj9p7RCB0_0;
	wire w_dff_B_Lnfhs4QJ8_0;
	wire w_dff_B_9wzovW1K1_0;
	wire w_dff_B_AYQXw4ah0_0;
	wire w_dff_B_EKrRSiUS5_0;
	wire w_dff_B_fCIcrYzg0_0;
	wire w_dff_B_vXM1eHmw1_0;
	wire w_dff_B_UaeLKGLt7_0;
	wire w_dff_B_lpELGz3b9_0;
	wire w_dff_B_EjCPy7S41_0;
	wire w_dff_B_x44aRKhf9_0;
	wire w_dff_B_V7eyhQDU8_0;
	wire w_dff_B_ODsq8MGz9_1;
	wire w_dff_B_5BhY4KmB4_1;
	wire w_dff_A_fVD0VTxf3_0;
	wire w_dff_A_j5OiPsNP5_0;
	wire w_dff_A_gWYGPnUF3_0;
	wire w_dff_A_tN7pN9zS4_0;
	wire w_dff_A_J8FNQi6d4_2;
	wire w_dff_A_LBlA3ipn0_2;
	wire w_dff_A_5jVlxlEd8_1;
	wire w_dff_A_IHZUTaxN7_1;
	wire w_dff_A_L8w0sTR85_1;
	wire w_dff_A_P39oH47z7_1;
	wire w_dff_A_8t14FyZA1_1;
	wire w_dff_A_pY7FLW693_1;
	wire w_dff_A_LPC2Hmgb2_1;
	wire w_dff_A_zUHE6OJp7_1;
	wire w_dff_A_8kFX6j9B3_2;
	wire w_dff_A_uLgdoARU2_2;
	wire w_dff_A_FT2KWkZO9_2;
	wire w_dff_A_zkyVJEDD9_2;
	wire w_dff_B_b3QgmtF84_3;
	wire w_dff_A_NxO5wa0G9_0;
	wire w_dff_A_v2tOVFxg8_0;
	wire w_dff_A_S9KUT1RQ5_0;
	wire w_dff_A_jS25Wu2N0_0;
	wire w_dff_A_0qt0LoFx1_0;
	wire w_dff_A_RlqxV35g6_0;
	wire w_dff_A_UG4xlEf71_0;
	wire w_dff_A_ZUTBvrie0_0;
	wire w_dff_A_rOaXI9Y85_1;
	wire w_dff_A_usYtItjc0_1;
	wire w_dff_A_osacSdo95_1;
	wire w_dff_A_QVXdpFrt1_0;
	wire w_dff_A_PddqTTdc0_1;
	wire w_dff_B_d3sjWix71_0;
	wire w_dff_B_A9hyVSUf9_0;
	wire w_dff_B_NUK6N2kP4_0;
	wire w_dff_B_3ZpBAuHt9_0;
	wire w_dff_B_dDNTTR8P3_0;
	wire w_dff_B_fxXG1myj6_0;
	wire w_dff_B_YXLkdU1c7_0;
	wire w_dff_B_fFUvJFBQ3_0;
	wire w_dff_B_5DHQsWWb3_0;
	wire w_dff_B_g2gwllFI2_0;
	wire w_dff_B_Nq2ZTkki8_0;
	wire w_dff_B_DpIp5SnS1_0;
	wire w_dff_B_7NIGw5Oa9_0;
	wire w_dff_B_CT8997VH1_1;
	wire w_dff_B_LjNP1xe75_1;
	wire w_dff_B_Cb6NJFBH6_3;
	wire w_dff_B_f8EmpGFW4_3;
	wire w_dff_A_JkGZyrSp0_1;
	wire w_dff_B_zfgiQdEd9_0;
	wire w_dff_B_4Q09WIFX4_3;
	wire w_dff_B_XX2WTl2R5_1;
	wire w_dff_A_EFjtmaS02_0;
	wire w_dff_A_b2cAoQXM2_1;
	wire w_dff_A_FvGkOaCi3_0;
	wire w_dff_A_SL2CkCQG0_1;
	wire w_dff_A_Rb2uXiFi0_0;
	wire w_dff_A_W6ugICTc9_0;
	wire w_dff_A_ntctoOUO0_0;
	wire w_dff_A_bnJMv21n0_0;
	wire w_dff_A_vkKShGM35_0;
	wire w_dff_A_0PYOUKfD7_1;
	wire w_dff_A_63Qn5KIc5_1;
	wire w_dff_A_5JtNalT21_1;
	wire w_dff_A_4FmLSURR9_1;
	wire w_dff_A_uTGBBX7c2_1;
	wire w_dff_A_pomlwqel7_1;
	wire w_dff_B_DTKs4Je02_0;
	wire w_dff_B_wDPyu4xs2_0;
	wire w_dff_B_I4ifPtmg6_0;
	wire w_dff_B_ZiaTwSdv9_0;
	wire w_dff_B_rlthOJX65_0;
	wire w_dff_B_hqaKMx2x5_0;
	wire w_dff_B_HWXO9WmH8_0;
	wire w_dff_B_huJjbbAv2_0;
	wire w_dff_B_ewH1lAGq8_0;
	wire w_dff_B_J6Yoh2Hq6_0;
	wire w_dff_B_ZWU5zdNs8_0;
	wire w_dff_B_SvYarsVD2_0;
	wire w_dff_B_VYJB5g7M7_0;
	wire w_dff_B_RntGXBae2_0;
	wire w_dff_B_azOiCFjl0_0;
	wire w_dff_B_ks6belN15_0;
	wire w_dff_B_nfMwAaDh9_0;
	wire w_dff_B_CDnC17cx4_0;
	wire w_dff_B_xSQVsPoZ2_2;
	wire w_dff_B_PEnNw0c31_2;
	wire w_dff_B_58usAc7i4_2;
	wire w_dff_B_eJUZaB8a5_0;
	wire w_dff_B_PzBOjRNh7_0;
	wire w_dff_B_d63iWvuT2_0;
	wire w_dff_B_DJpVwbnP6_0;
	wire w_dff_B_I2jWeDpn4_0;
	wire w_dff_B_Oj6apF427_0;
	wire w_dff_B_EvuBXMid2_0;
	wire w_dff_B_ckMwtmqC4_0;
	wire w_dff_B_CBRfLtzW5_0;
	wire w_dff_B_loyjdCvL4_0;
	wire w_dff_B_edH823860_0;
	wire w_dff_B_yNJqNkWF5_0;
	wire w_dff_B_J5ifSxXj6_0;
	wire w_dff_B_4yZCFnr61_1;
	wire w_dff_B_kWE29rax3_1;
	wire w_dff_A_Oy42UHnV4_1;
	wire w_dff_A_hzg3IKyz0_0;
	wire w_dff_B_HPz1yzyw0_2;
	wire w_dff_B_9gUly01L6_0;
	wire w_dff_B_XBueP9mY3_0;
	wire w_dff_B_2aJGrS2I8_0;
	wire w_dff_B_5Ubx6wng4_0;
	wire w_dff_A_YoUpGZEF4_0;
	wire w_dff_A_rPl93rKj3_0;
	wire w_dff_A_mrLIkdhc0_0;
	wire w_dff_A_HX7RCHHO4_0;
	wire w_dff_A_32h8KHfo0_0;
	wire w_dff_A_VTwCLqoy3_0;
	wire w_dff_A_TrW88K8S7_0;
	wire w_dff_A_TBOZGujq2_0;
	wire w_dff_A_MmPMhp1X7_0;
	wire w_dff_A_M3lqmndX0_0;
	wire w_dff_A_CHgitgri5_0;
	wire w_dff_A_uYvlz1NO4_0;
	wire w_dff_A_HeLRgrdp3_0;
	wire w_dff_A_9miJU0V01_0;
	wire w_dff_A_1huJGL037_0;
	wire w_dff_A_HwQ6OJs31_0;
	wire w_dff_A_TXqFKuK68_0;
	wire w_dff_A_q1y4R3CG4_0;
	wire w_dff_A_X0si2R2Z8_0;
	wire w_dff_A_69179VsI2_0;
	wire w_dff_A_wyGNDgss6_1;
	wire w_dff_A_4vjFKfps3_1;
	wire w_dff_A_z46HEOva8_1;
	wire w_dff_A_3FY1pyvB8_1;
	wire w_dff_A_v7267uGc8_1;
	wire w_dff_A_DiLJ8cCA6_1;
	wire w_dff_A_2Llhfgir8_1;
	wire w_dff_A_vLqVZ47g5_1;
	wire w_dff_A_Kd60217a3_1;
	wire w_dff_B_ftj9PPAC3_0;
	wire w_dff_B_dGKwyCEr2_0;
	wire w_dff_B_WepTQcQ25_0;
	wire w_dff_B_varN7BWI9_0;
	wire w_dff_B_X8KuPgAP6_0;
	wire w_dff_B_XZkzsrjA4_0;
	wire w_dff_B_vA3MOdfZ5_0;
	wire w_dff_B_TaAtuTab9_0;
	wire w_dff_B_Ign8YJUD7_0;
	wire w_dff_B_RqHIxS1O1_0;
	wire w_dff_B_P1vGgqKr0_0;
	wire w_dff_B_jKj3SKn22_0;
	wire w_dff_B_mdPyiKmd0_0;
	wire w_dff_B_eVuEP4Ca2_0;
	wire w_dff_B_PwIuOo4U9_0;
	wire w_dff_B_QVpp9gnE7_0;
	wire w_dff_B_S4Fe6U2p7_1;
	wire w_dff_B_iunU92P06_1;
	wire w_dff_A_IVzXe4al7_0;
	wire w_dff_A_haZpLyY01_2;
	wire w_dff_A_gn3eJPS54_2;
	wire w_dff_A_8JIFM9F91_2;
	wire w_dff_A_8Wcm2ddZ5_2;
	wire w_dff_B_yyeTZfAc2_1;
	wire w_dff_B_mN6QhgZ65_1;
	wire w_dff_B_TOeqyTOR4_1;
	wire w_dff_B_0Gox7zAp4_1;
	wire w_dff_B_j0TWinXw0_1;
	wire w_dff_B_hzkoANlZ1_1;
	wire w_dff_B_NWCCJe449_1;
	wire w_dff_B_SaJAM3N00_1;
	wire w_dff_B_TVmDremS7_1;
	wire w_dff_B_Qs7JBXrM6_1;
	wire w_dff_B_6fy14eq14_1;
	wire w_dff_B_kYixEY4a3_1;
	wire w_dff_B_HinJg8jy0_1;
	wire w_dff_B_PjRshg3R5_1;
	wire w_dff_B_Zkjoqe727_1;
	wire w_dff_B_SfmGU9ge5_1;
	wire w_dff_B_2Sr2ebjQ1_1;
	wire w_dff_B_6DbqdCFJ1_1;
	wire w_dff_B_bdh2mSot5_0;
	wire w_dff_A_WyfAoSHm2_1;
	wire w_dff_A_XyHvh8tW7_1;
	wire w_dff_A_9i4LzyXu3_1;
	wire w_dff_A_UMt1k7Kl5_1;
	wire w_dff_A_2hMQhhdO6_1;
	wire w_dff_A_R0DOJt8p2_1;
	wire w_dff_B_J2gxHcmX2_3;
	wire w_dff_B_Veimd5dm5_3;
	wire w_dff_B_FSgLnOcW1_3;
	wire w_dff_B_gvIUJVje8_3;
	wire w_dff_B_x5wLkZTT7_2;
	wire w_dff_B_sRnUQIOa6_2;
	wire w_dff_B_VevBZNSP7_2;
	wire w_dff_B_yQdwIGbX9_2;
	wire w_dff_B_MWUfwYei7_2;
	wire w_dff_B_jMgDRVhY1_2;
	wire w_dff_B_t5t3bqkt4_2;
	wire w_dff_B_888HJOmE2_2;
	wire w_dff_B_XYG7lamz1_2;
	wire w_dff_A_hWd10c6p4_1;
	wire w_dff_A_AiVdoE9f6_1;
	wire w_dff_A_kc7C7W6D4_1;
	wire w_dff_A_ByfD1gwT6_2;
	wire w_dff_A_cQoM0L162_2;
	wire w_dff_A_nNpSSEUv5_2;
	wire w_dff_A_S4pNyZOJ2_2;
	wire w_dff_A_P6KUHL7z1_0;
	wire w_dff_A_UhCBGmq06_0;
	wire w_dff_A_11kaPSjM9_0;
	wire w_dff_A_qrUWHeLz4_0;
	wire w_dff_A_uxhWYyQZ6_0;
	wire w_dff_A_1qWIZ3Oq3_0;
	wire w_dff_A_7jLEpLmB7_0;
	wire w_dff_A_RX6X5bl79_0;
	wire w_dff_A_FxjLs9uE6_0;
	wire w_dff_A_vlgcW8f95_0;
	wire w_dff_A_51RSWDjd1_0;
	wire w_dff_A_9SD8CUQk2_0;
	wire w_dff_A_abiRJ84q1_0;
	wire w_dff_A_iBdvOCbi2_1;
	wire w_dff_A_iDHxzIDQ1_1;
	wire w_dff_A_6kX2OLqW3_1;
	wire w_dff_A_cbqwSQcX3_1;
	wire w_dff_A_UcFqDnAN4_1;
	wire w_dff_A_NxSXq9pw3_1;
	wire w_dff_A_xVwWe8BZ7_1;
	wire w_dff_B_PSSVQYrh3_1;
	wire w_dff_B_GWrBT2oc0_1;
	wire w_dff_B_BPn9TLUF8_1;
	wire w_dff_B_V3j6wOGE2_1;
	wire w_dff_B_lgN5BTih8_1;
	wire w_dff_B_8BjmnNm32_1;
	wire w_dff_B_WVpGlc070_1;
	wire w_dff_B_1antOYHT0_1;
	wire w_dff_B_qYgqs6c76_1;
	wire w_dff_B_lmcnPDen9_1;
	wire w_dff_B_0NpLdZnA4_1;
	wire w_dff_B_Mkz1S36q9_1;
	wire w_dff_B_mOrDmNbH4_1;
	wire w_dff_B_pfK1Bm0p9_1;
	wire w_dff_B_uIKEDw5W5_1;
	wire w_dff_B_YsNcVzEP7_1;
	wire w_dff_B_KfYjRf515_1;
	wire w_dff_B_Ebp6XgBG9_1;
	wire w_dff_B_tlTNiJrb5_1;
	wire w_dff_B_MWXMhdj96_1;
	wire w_dff_B_8Uz3ufRE5_1;
	wire w_dff_B_ltAbWIpY0_1;
	wire w_dff_B_XSI6BZJ17_1;
	wire w_dff_B_I4krucv43_1;
	wire w_dff_B_HeM22eFF6_1;
	wire w_dff_B_T1L9PIeW3_1;
	wire w_dff_B_JABImF1M5_1;
	wire w_dff_B_ryMj8vOZ6_1;
	wire w_dff_B_LukVAR2m2_1;
	wire w_dff_B_rmeqPkzb6_1;
	wire w_dff_B_PYfzAJdU4_1;
	wire w_dff_B_dgJ8ImcE7_1;
	wire w_dff_B_B9eDp4U79_1;
	wire w_dff_B_g6TnYnbD2_1;
	wire w_dff_B_kVpeL4lv1_1;
	wire w_dff_B_OwUHNzMz9_1;
	wire w_dff_B_vuf4YPWQ8_1;
	wire w_dff_B_IIdqX6mj8_1;
	wire w_dff_B_MEO3d8q96_0;
	wire w_dff_B_VHEjOWlr0_0;
	wire w_dff_B_gb6Z3Xyr5_0;
	wire w_dff_B_7YHFJ8k35_0;
	wire w_dff_B_GmCHsWyE2_0;
	wire w_dff_B_Ak80ZyMS2_0;
	wire w_dff_B_wvvFKVFb1_0;
	wire w_dff_B_70wj62FA1_0;
	wire w_dff_B_OvL07NLV3_0;
	wire w_dff_B_3drzL6rn1_0;
	wire w_dff_B_oZixLIUj2_0;
	wire w_dff_B_FGwDbZqe6_0;
	wire w_dff_B_Zti4Bcwo5_0;
	wire w_dff_B_MqvdPi8I7_0;
	wire w_dff_B_VNS2lQhf0_0;
	wire w_dff_B_1rTQDNlf5_0;
	wire w_dff_B_F5zOduc43_0;
	wire w_dff_B_4cT38ERN0_0;
	wire w_dff_B_FstWOxMJ7_0;
	wire w_dff_B_kA3QnmlP5_0;
	wire w_dff_A_2BHRjPXu5_1;
	wire w_dff_A_LJVlJdj69_1;
	wire w_dff_A_4YpHF1Qd3_1;
	wire w_dff_A_Y5YYbz3i8_1;
	wire w_dff_A_4vHBkBSS9_1;
	wire w_dff_A_GV2pKAxt7_1;
	wire w_dff_A_4WxEcWCe0_1;
	wire w_dff_A_FE8svY6X9_1;
	wire w_dff_A_cYQJnmg89_1;
	wire w_dff_A_6WpXnb3N2_1;
	wire w_dff_A_GjMKJfzx8_1;
	wire w_dff_A_o4ULUWFk4_1;
	wire w_dff_A_pPqHdtgv5_1;
	wire w_dff_A_qovNcWLc4_1;
	wire w_dff_A_NVQNgztX5_2;
	wire w_dff_A_IkFHensy2_2;
	wire w_dff_A_Hgmw9N1F1_2;
	wire w_dff_A_4CWqr7sf6_2;
	wire w_dff_A_DOBDqk9r7_2;
	wire w_dff_A_Lojwy1gj1_2;
	wire w_dff_A_ZbrkCbDh2_2;
	wire w_dff_A_xDbl4HMC9_2;
	wire w_dff_A_U8B4g5eB9_2;
	wire w_dff_A_Ae5SNb7y0_2;
	wire w_dff_A_uQaMhm7w3_1;
	wire w_dff_A_HTvE6bvC6_1;
	wire w_dff_A_ORetPWpf6_1;
	wire w_dff_A_yu2u2imy1_1;
	wire w_dff_A_hCJ9zakk6_1;
	wire w_dff_A_9JP1G19y9_1;
	wire w_dff_A_0HOBUu6H1_1;
	wire w_dff_A_ANaYa1m63_1;
	wire w_dff_A_hmQ0hxrp3_1;
	wire w_dff_A_sVUU8jRG6_1;
	wire w_dff_A_la6I0zsv1_1;
	wire w_dff_A_8c8YIv9Z3_2;
	wire w_dff_B_zVdn96Cx9_3;
	wire w_dff_B_TMWmsUoR4_3;
	wire w_dff_B_40VEXi2C3_3;
	wire w_dff_B_KkIoLw2R3_3;
	wire w_dff_B_2EgDjwaa5_3;
	wire w_dff_B_fkxGB2wk5_3;
	wire w_dff_A_SynBGV085_1;
	wire w_dff_A_wKGgSIdq1_1;
	wire w_dff_A_xOqzB6Bb7_1;
	wire w_dff_A_ozvAaHc46_1;
	wire w_dff_A_Y4Q8Nrql6_1;
	wire w_dff_A_JCmx0ffA6_1;
	wire w_dff_A_OXO3dpd57_1;
	wire w_dff_A_GR1KqTtM4_1;
	wire w_dff_A_OFDBwyRn8_1;
	wire w_dff_A_hjzhQks09_1;
	wire w_dff_A_cWBI7L8L6_1;
	wire w_dff_A_ZAAGuerl8_1;
	wire w_dff_A_mHwsDrOt3_1;
	wire w_dff_A_awGli8B57_1;
	wire w_dff_A_zef5JSYo2_2;
	wire w_dff_A_1Lql7xGW3_2;
	wire w_dff_A_0DNp4rkF4_2;
	wire w_dff_A_zBUdklzJ2_2;
	wire w_dff_A_GVTjFlIY3_2;
	wire w_dff_A_jTp48KP56_2;
	wire w_dff_A_XKPibHSf7_2;
	wire w_dff_A_BncmWU7u7_2;
	wire w_dff_A_Pp0eBHjk0_2;
	wire w_dff_A_lGSOXHj04_2;
	wire w_dff_A_VWPGiUH60_1;
	wire w_dff_A_JUlOSG6o2_1;
	wire w_dff_A_RwwjwGFi3_1;
	wire w_dff_A_QVtGEvtA2_1;
	wire w_dff_A_sJ25soSa6_1;
	wire w_dff_A_yEwyVCMS4_1;
	wire w_dff_A_6G3CynG85_1;
	wire w_dff_A_I1FjocQF5_1;
	wire w_dff_A_FBNhkPIT1_1;
	wire w_dff_A_b4WFldKb4_1;
	wire w_dff_A_Uck6BVVc7_1;
	wire w_dff_A_gUyPHObs8_2;
	wire w_dff_A_b8It70LO1_2;
	wire w_dff_A_1qjmRQCl2_2;
	wire w_dff_A_uxzSyXNv7_2;
	wire w_dff_B_K9AGMGuF9_3;
	wire w_dff_B_ls42C8lp4_3;
	wire w_dff_B_iZ4BEQyX0_3;
	wire w_dff_B_t3wNn53i8_3;
	wire w_dff_B_BoAcDQIB4_3;
	wire w_dff_B_5nmvW88k8_3;
	wire w_dff_B_IRk8CjcP4_3;
	wire w_dff_A_6ma5F38f2_2;
	wire w_dff_A_FTuHRH8f2_1;
	wire w_dff_B_mx8n3Ai93_0;
	wire w_dff_B_pYp3CDu43_0;
	wire w_dff_B_TtueYOmb7_0;
	wire w_dff_B_mYjxnGuU6_0;
	wire w_dff_B_CMWquzL43_0;
	wire w_dff_B_WfZNkflh7_0;
	wire w_dff_B_qoGGw7bJ8_0;
	wire w_dff_B_vBExeG9j5_0;
	wire w_dff_B_70K05SSy7_0;
	wire w_dff_B_IEckeMl75_0;
	wire w_dff_B_bksrw7pz2_0;
	wire w_dff_B_LIty7jJU6_0;
	wire w_dff_B_E7Cpwizy1_0;
	wire w_dff_B_vGKvDKpH7_0;
	wire w_dff_B_fqtQOO3N8_0;
	wire w_dff_B_E9XrPimD5_0;
	wire w_dff_B_c4uEurZK0_0;
	wire w_dff_B_bvS3vdT85_0;
	wire w_dff_B_UYe82NPj3_0;
	wire w_dff_B_1tJj2pw78_0;
	wire w_dff_B_CPdioXsj6_2;
	wire w_dff_B_qMQsQAo42_2;
	wire w_dff_B_DbS2HEhc5_2;
	wire w_dff_A_VeM1GuY34_1;
	wire w_dff_A_6a1bTLaC6_1;
	wire w_dff_A_t720y4za9_1;
	wire w_dff_A_nKAuaDZ02_1;
	wire w_dff_A_wUwsDg1W0_1;
	wire w_dff_A_cVplHmUC6_1;
	wire w_dff_A_xUHOb8jG3_1;
	wire w_dff_A_JX3J5xJw3_1;
	wire w_dff_A_cWkChUra6_1;
	wire w_dff_A_7AHSfJsd7_1;
	wire w_dff_A_uyzX1rmX9_1;
	wire w_dff_A_eee57DFl7_1;
	wire w_dff_A_645HeLnO7_1;
	wire w_dff_A_0HiOG1SP1_1;
	wire w_dff_A_fK4K6jJQ3_2;
	wire w_dff_A_sEiEdIec8_2;
	wire w_dff_A_MwHMJvDL0_2;
	wire w_dff_A_kJ2H4MXc8_2;
	wire w_dff_A_1feiUy8v1_2;
	wire w_dff_A_7meb2ZSk9_2;
	wire w_dff_A_uc3PKkxM1_2;
	wire w_dff_A_cJgrrRaW3_2;
	wire w_dff_A_8xG2O6Ia9_2;
	wire w_dff_A_vuhtRYQD6_2;
	wire w_dff_A_rX4X66Vn6_1;
	wire w_dff_A_jDPgrLWs8_1;
	wire w_dff_A_GF5krNfO1_1;
	wire w_dff_A_yw0hccLG8_1;
	wire w_dff_A_acblp5LJ1_1;
	wire w_dff_A_r9fnHnR71_1;
	wire w_dff_A_nfyVuQPC0_1;
	wire w_dff_A_o0CrjVkS6_1;
	wire w_dff_A_zhWSMOFn1_1;
	wire w_dff_A_swpKsueu3_1;
	wire w_dff_A_mwCoMitu7_1;
	wire w_dff_A_b3PzTxgP3_2;
	wire w_dff_B_NFYmXjap0_3;
	wire w_dff_B_3R7hbTLo8_3;
	wire w_dff_B_AfquKikj8_3;
	wire w_dff_B_lDHjV6Yj7_3;
	wire w_dff_B_DKrBzNRP3_3;
	wire w_dff_B_NoFcKoJw2_3;
	wire w_dff_A_nkBkbhDA8_1;
	wire w_dff_A_scfkKZjy8_1;
	wire w_dff_A_5Owzi61p1_1;
	wire w_dff_A_JbVPKepv2_1;
	wire w_dff_A_73sVhA7w9_1;
	wire w_dff_A_nIwBCpXi4_1;
	wire w_dff_A_Il49YHsk4_1;
	wire w_dff_A_wKmW8qMj5_1;
	wire w_dff_A_TZaCrk1i3_1;
	wire w_dff_A_3oDxbYye3_1;
	wire w_dff_A_DIG9kD0N3_1;
	wire w_dff_A_cMMATo8X4_1;
	wire w_dff_A_RWlZCJbu3_1;
	wire w_dff_A_oPFxAwah3_1;
	wire w_dff_A_a7UFN0Uh7_2;
	wire w_dff_A_sRSC3A8A5_2;
	wire w_dff_A_Ta3DWYTB1_2;
	wire w_dff_A_w0BZivgt0_2;
	wire w_dff_A_5kjiY2cf5_2;
	wire w_dff_A_1I1ajFIP4_2;
	wire w_dff_A_FVbyTzEw9_2;
	wire w_dff_A_vXMhNBiR8_2;
	wire w_dff_A_kVbLXsRG9_2;
	wire w_dff_A_Jy2uufCu7_2;
	wire w_dff_A_e6TerabC0_1;
	wire w_dff_A_UGLdQg8w9_1;
	wire w_dff_A_HWTMfyzp4_1;
	wire w_dff_A_6ICfHWwi1_1;
	wire w_dff_A_iPYLaqK78_1;
	wire w_dff_A_yaxkx7d88_1;
	wire w_dff_A_UuH9XUSa5_1;
	wire w_dff_A_aaa9mnAP7_1;
	wire w_dff_A_FOV1LhKx1_1;
	wire w_dff_A_XTjON36r5_1;
	wire w_dff_A_I5c4OnJa6_1;
	wire w_dff_A_MxddZJHs5_2;
	wire w_dff_A_XZbvFUvd6_2;
	wire w_dff_A_UmX0EuCz9_2;
	wire w_dff_A_6bUW0NZ23_2;
	wire w_dff_B_Qtn3h0Tm6_3;
	wire w_dff_B_ELWWf9620_3;
	wire w_dff_B_r1lnAy1I3_3;
	wire w_dff_B_WA2DV3Vf0_3;
	wire w_dff_B_8R7J4r6g0_3;
	wire w_dff_B_03qcQDFT5_3;
	wire w_dff_B_Ua5DCBO99_3;
	wire w_dff_A_BadhDM3A4_1;
	wire w_dff_A_uFn2pNSI7_2;
	wire w_dff_B_xA0vYSin2_1;
	wire w_dff_B_n078xPUD8_0;
	wire w_dff_B_pt6MItKr0_0;
	wire w_dff_B_rosl3jPX7_0;
	wire w_dff_B_Rgbv2Gtx3_0;
	wire w_dff_B_BhTC6eJE4_0;
	wire w_dff_B_MoC5iSjJ4_0;
	wire w_dff_B_k3ACB6772_0;
	wire w_dff_B_o8CZ3GWW8_0;
	wire w_dff_B_8hTS6JfU3_0;
	wire w_dff_B_Ji3yWvM96_0;
	wire w_dff_B_h2uuehdI9_0;
	wire w_dff_B_CTQRxkAh3_0;
	wire w_dff_B_CHKDEOLe6_0;
	wire w_dff_B_37hP9ygD1_0;
	wire w_dff_B_Tlcay7sT3_0;
	wire w_dff_B_4silvIz19_0;
	wire w_dff_B_2h1HXx4o1_0;
	wire w_dff_B_NEceM8xN0_0;
	wire w_dff_B_QBM2HGO14_1;
	wire w_dff_B_WjCopaOU8_1;
	wire w_dff_B_N8wIuoDw7_1;
	wire w_dff_B_mJ4NKWRl2_1;
	wire w_dff_B_UwRxg3MX7_1;
	wire w_dff_B_lqs2ydvD0_1;
	wire w_dff_B_LARZFADt4_1;
	wire w_dff_B_ujqEeYer1_1;
	wire w_dff_B_hHxvGh243_1;
	wire w_dff_B_w8EFnRTn7_1;
	wire w_dff_B_qvajMSfs0_1;
	wire w_dff_B_wy5GZvL64_1;
	wire w_dff_B_BGnLcEqz5_1;
	wire w_dff_B_Ons9LCHV0_1;
	wire w_dff_B_fqiDJapU6_1;
	wire w_dff_B_tZ2zDv4U8_1;
	wire w_dff_B_8mQQFoVP2_1;
	wire w_dff_B_0knoR80E4_1;
	wire w_dff_B_mPyZHcJA0_1;
	wire w_dff_B_q3Yf7HM58_1;
	wire w_dff_A_zANiK10X9_0;
	wire w_dff_A_2PnpBSVi1_0;
	wire w_dff_A_DFUg5kjj4_0;
	wire w_dff_A_wvnkraax7_0;
	wire w_dff_A_bvbp1zIY8_0;
	wire w_dff_A_gpHh6toS5_0;
	wire w_dff_A_D8IjNm4D3_2;
	wire w_dff_A_n13TQpRP8_2;
	wire w_dff_A_V9gmVsjw0_2;
	wire w_dff_A_PnQXDKMq4_2;
	wire w_dff_A_lZzUJE1h5_2;
	wire w_dff_A_DxTfdG1h9_2;
	wire w_dff_A_nXm9wK0P5_2;
	wire w_dff_A_4Ql8qXpc2_2;
	wire w_dff_A_zk4VSNBZ8_2;
	wire w_dff_A_DHmrZ5j96_2;
	wire w_dff_A_8VvYjaXq2_2;
	wire w_dff_A_WQ6uCOAq7_2;
	wire w_dff_A_YJEoqH5y8_2;
	wire w_dff_A_rXImKdHt6_2;
	wire w_dff_A_pZ2PQGNC5_2;
	wire w_dff_A_LDgOPlyo7_2;
	wire w_dff_A_o2NXtWKY2_2;
	wire w_dff_A_Z7o0FbIx1_2;
	wire w_dff_A_cvvYCVZ33_1;
	wire w_dff_A_ZjkvOD6o5_1;
	wire w_dff_A_UfWuBhFF1_1;
	wire w_dff_A_TkueEScT3_1;
	wire w_dff_A_Y8I6zfIG7_1;
	wire w_dff_A_pdRsSaV75_1;
	wire w_dff_A_4yuWQuL74_1;
	wire w_dff_A_ECEsCU3W5_1;
	wire w_dff_A_8oUDouHL9_1;
	wire w_dff_A_gkGDwd6X0_1;
	wire w_dff_A_KD6QhGAK3_1;
	wire w_dff_A_JZ1ywGXq7_1;
	wire w_dff_A_jBBKyDco1_1;
	wire w_dff_A_yGWARj6r5_1;
	wire w_dff_A_K9wO8y109_1;
	wire w_dff_A_B9uKgh0B8_1;
	wire w_dff_A_yR3LGZKu2_2;
	wire w_dff_A_CRiNvvDn3_2;
	wire w_dff_A_lrUAb7493_2;
	wire w_dff_A_jWMlgr7T7_2;
	wire w_dff_A_HuxvSMAX5_2;
	wire w_dff_A_SUgE56ZD8_2;
	wire w_dff_A_P2IcOBYT4_2;
	wire w_dff_B_doFl3vwD2_1;
	wire w_dff_B_SUI2ZvpX9_1;
	wire w_dff_B_dXfk9olI7_1;
	wire w_dff_B_EPtCOdgg2_1;
	wire w_dff_B_x6QRsMbM7_1;
	wire w_dff_B_f1n1Y4Mm8_1;
	wire w_dff_B_OvCy6SmH8_1;
	wire w_dff_B_LZouneJq7_1;
	wire w_dff_B_KSKsdCZ91_1;
	wire w_dff_B_ugv3GUcQ4_1;
	wire w_dff_B_F34WJs6U2_1;
	wire w_dff_B_qYY2eNcY6_1;
	wire w_dff_B_WhrdeZgS6_1;
	wire w_dff_B_dqS2YwLH8_1;
	wire w_dff_B_DwhQ158Q2_1;
	wire w_dff_B_28FqjB0d4_1;
	wire w_dff_B_LP409KKA4_1;
	wire w_dff_B_XL4HHL9f7_1;
	wire w_dff_B_uSrom04Y5_1;
	wire w_dff_A_OHWGpSNV7_0;
	wire w_dff_A_h2N8nIye8_0;
	wire w_dff_A_8eXgH3K64_0;
	wire w_dff_A_xP8nRnYM1_0;
	wire w_dff_A_WhF8GNAk2_0;
	wire w_dff_A_EtEfJ8W07_0;
	wire w_dff_A_T9vIVRvM5_0;
	wire w_dff_A_YO0mP3XC1_2;
	wire w_dff_A_YoNUvkDx4_2;
	wire w_dff_A_iBAILy4o7_2;
	wire w_dff_A_feSVqn7k0_2;
	wire w_dff_A_ChpdGrbB6_2;
	wire w_dff_A_dABCwaV04_2;
	wire w_dff_A_InRfc20D5_2;
	wire w_dff_A_0luYfXCa4_2;
	wire w_dff_A_i3zcEiMj3_2;
	wire w_dff_A_4QLG6wQk6_2;
	wire w_dff_A_gtJvAjE86_2;
	wire w_dff_A_amNgEKYR2_2;
	wire w_dff_A_WXrBAOZO8_2;
	wire w_dff_A_FhYieZXV1_2;
	wire w_dff_A_6eZMbTnv8_2;
	wire w_dff_A_VDJHXKIq1_2;
	wire w_dff_A_zRfb5UVR3_2;
	wire w_dff_A_dyh85Ttw8_2;
	wire w_dff_A_MLToMRuZ9_2;
	wire w_dff_A_aeKAGSCg7_1;
	wire w_dff_A_pfKC3rsj5_1;
	wire w_dff_A_Jnk0oSli6_1;
	wire w_dff_A_9CdXQzzd2_1;
	wire w_dff_A_B34x5AsY1_1;
	wire w_dff_A_OswyhW3j2_1;
	wire w_dff_A_rAQPOaZk1_1;
	wire w_dff_A_snh6lWUk2_1;
	wire w_dff_A_odiIjmux2_1;
	wire w_dff_A_nvgoEXNm3_1;
	wire w_dff_A_aT01ZwOF8_1;
	wire w_dff_A_R2L2rZlr7_1;
	wire w_dff_A_4iqUQ62V3_1;
	wire w_dff_A_rKHVtsEn3_1;
	wire w_dff_A_Y0q6fX3z8_1;
	wire w_dff_A_kNhOidYe1_1;
	wire w_dff_A_iYxEkZyg0_1;
	wire w_dff_A_PqB0lklw9_2;
	wire w_dff_A_vWwPitHK1_2;
	wire w_dff_A_hpj13S168_2;
	wire w_dff_A_vqPZKqIW7_2;
	wire w_dff_A_HMpgyEEf3_2;
	wire w_dff_A_w8nAFFtp9_2;
	wire w_dff_A_XPh3pkSs5_2;
	wire w_dff_A_YVBetRxS7_2;
	wire w_dff_A_uSe7Axul1_2;
	wire w_dff_A_p0emwRUY2_2;
	wire w_dff_A_ICJEW9YY6_2;
	wire w_dff_A_TzPdTV922_1;
	wire w_dff_A_jZQpmhwB0_2;
	wire w_dff_B_BsnuMHo72_1;
	wire w_dff_B_0OQA9ptp4_0;
	wire w_dff_B_ZyxEP5N92_0;
	wire w_dff_B_OyDk8pw65_0;
	wire w_dff_B_hQKoiH9Y0_0;
	wire w_dff_B_r7cCnYQ74_0;
	wire w_dff_B_wS7Pabpk7_0;
	wire w_dff_B_eRCu8QB44_0;
	wire w_dff_B_NCtyN3dR2_0;
	wire w_dff_B_PpsFzXUk3_0;
	wire w_dff_B_v9lsnwlz1_0;
	wire w_dff_B_S72YKBWS7_0;
	wire w_dff_B_twFnlQqg3_0;
	wire w_dff_B_JtyBBIX31_0;
	wire w_dff_B_moRuQVvE6_0;
	wire w_dff_B_Ohgyme1S1_0;
	wire w_dff_B_6RFN7g056_0;
	wire w_dff_B_H6W0Emv19_0;
	wire w_dff_B_CGcUBzOR8_0;
	wire w_dff_B_bVOuko2y1_1;
	wire w_dff_B_U24SoQQf7_2;
	wire w_dff_B_oUZfakXc6_2;
	wire w_dff_B_JuqoCnrz3_2;
	wire w_dff_B_OKfdq3cA1_1;
	wire w_dff_B_8PX1GDoU5_1;
	wire w_dff_B_2r2ydSlc4_1;
	wire w_dff_B_hJTvTNBh9_1;
	wire w_dff_B_gdyVWrjk2_1;
	wire w_dff_B_TaKh9HbN9_1;
	wire w_dff_B_AZcMHsa48_1;
	wire w_dff_B_6lxmEqr84_1;
	wire w_dff_B_NtIZYNf47_1;
	wire w_dff_B_B0icVx8h9_1;
	wire w_dff_B_kIFZwWzd7_1;
	wire w_dff_B_2KSacEBF3_1;
	wire w_dff_B_sLSg93yN4_1;
	wire w_dff_B_ZANhEngS8_1;
	wire w_dff_B_uYxTnCUy7_1;
	wire w_dff_B_8uTCp8Hn8_1;
	wire w_dff_B_NRIVh24E0_1;
	wire w_dff_B_1I29x71r3_1;
	wire w_dff_B_dX64z8cV0_1;
	wire w_dff_B_iNw3Vakc1_0;
	wire w_dff_B_F6YrgLL71_0;
	wire w_dff_B_Rc4dgdeP1_0;
	wire w_dff_B_DlpLbvfb8_0;
	wire w_dff_B_rGm3yYio7_0;
	wire w_dff_B_93RtKOiA9_0;
	wire w_dff_B_cSGC9RYB8_0;
	wire w_dff_B_OMrgHnLd1_0;
	wire w_dff_B_qJzYmhjs5_0;
	wire w_dff_B_Stv8tSr94_0;
	wire w_dff_B_rP4eNdoI2_0;
	wire w_dff_B_1QiusGXx5_0;
	wire w_dff_B_mUy9AMw66_0;
	wire w_dff_B_ZFPbteDe2_0;
	wire w_dff_B_cvJSCxbs5_0;
	wire w_dff_B_Tya8Tj9E5_0;
	wire w_dff_B_2tVAfDUS6_0;
	wire w_dff_B_Shy0yNC95_0;
	wire w_dff_B_MRWuuE6D0_0;
	wire w_dff_A_FHG5wHSW6_1;
	wire w_dff_A_LU26bgDI7_1;
	wire w_dff_A_sYZxVC6p4_1;
	wire w_dff_A_26HXs43r8_1;
	wire w_dff_A_lZ7eUrRG4_1;
	wire w_dff_A_FUVFASAc3_1;
	wire w_dff_A_m2doOAnp6_1;
	wire w_dff_A_SL8JSuej4_1;
	wire w_dff_A_OPVl9SYl6_1;
	wire w_dff_A_9pWn6sQk9_1;
	wire w_dff_A_kAkLYPmA7_1;
	wire w_dff_A_bzrmhNfn7_1;
	wire w_dff_A_xoxhGbk60_1;
	wire w_dff_A_UTf2MXfn7_1;
	wire w_dff_A_ecD7gx984_1;
	wire w_dff_A_22JSAGlj9_1;
	wire w_dff_A_6MWHxteX0_1;
	wire w_dff_A_CCd8nReW7_1;
	wire w_dff_A_bzIOoVfs3_1;
	wire w_dff_A_8ibn2ThK1_1;
	wire w_dff_B_lUZDsqeU1_1;
	wire w_dff_B_z42zrVKM5_1;
	wire w_dff_B_QSnSHTIl6_1;
	wire w_dff_B_EFsU1XA45_1;
	wire w_dff_B_cKc2TOh76_1;
	wire w_dff_B_CQpW27lF9_1;
	wire w_dff_A_fgrJABZv7_1;
	wire w_dff_B_YlSAaHFt4_1;
	wire w_dff_B_F4g3du833_1;
	wire w_dff_B_LBs5Rtdw0_1;
	wire w_dff_B_REGeQgUa0_1;
	wire w_dff_B_ZPyW40H24_1;
	wire w_dff_B_rfRIYaNb9_1;
	wire w_dff_B_2aMxh9bk1_1;
	wire w_dff_B_0B84Cl4m5_1;
	wire w_dff_B_wBbD3bNt9_1;
	wire w_dff_B_d8pD8Ezv4_1;
	wire w_dff_B_ANg88wro8_0;
	wire w_dff_B_9GLwzPEr8_0;
	wire w_dff_A_QtvilpXc4_1;
	wire w_dff_A_uPM6mDAw0_1;
	wire w_dff_A_KzB0g1Nb1_1;
	wire w_dff_B_y9QNuL3z4_0;
	wire w_dff_B_dFCMmpUR1_1;
	wire w_dff_B_uHKiqOJY7_1;
	wire w_dff_B_cUJPDF5T8_1;
	wire w_dff_B_76hbirnt5_1;
	wire w_dff_B_R5ODUbWW7_1;
	wire w_dff_B_JVbrCqGZ3_1;
	wire w_dff_B_URvx2Jvn2_1;
	wire w_dff_B_SIU56iQI0_1;
	wire w_dff_B_BbDFpwmB6_1;
	wire w_dff_B_7U2Armpn8_1;
	wire w_dff_B_SQFxn9UY4_1;
	wire w_dff_B_7J4yUeo43_1;
	wire w_dff_B_CNapvRPK9_1;
	wire w_dff_B_9NzEBlA36_1;
	wire w_dff_B_ZqSJntMl5_1;
	wire w_dff_B_vj4uRcAr3_1;
	wire w_dff_B_jPIh30mM3_1;
	wire w_dff_B_fXge62pK6_0;
	wire w_dff_A_ChlsoDwO8_0;
	wire w_dff_A_0ay4vSmU3_0;
	wire w_dff_A_JXVu36Ka7_0;
	wire w_dff_B_AHQpbTXO6_1;
	wire w_dff_A_C6FdzPPt8_1;
	wire w_dff_A_w48cUdHX2_0;
	wire w_dff_A_EaANQjNV7_0;
	wire w_dff_A_aRyKXAax3_0;
	wire w_dff_A_TfB8AK0q8_0;
	wire w_dff_A_pBW3DPRX8_0;
	wire w_dff_A_rxs2INgK8_2;
	wire w_dff_A_UQB2RqFo7_2;
	wire w_dff_A_Tx2A3lWa6_2;
	wire w_dff_A_J04wO39a1_2;
	wire w_dff_A_H3wNa1iM6_2;
	wire w_dff_A_LOEMaROP6_2;
	wire w_dff_A_QOi2xMeJ2_1;
	wire w_dff_A_cwgcIkMW2_1;
	wire w_dff_A_EpDPndjc0_1;
	wire w_dff_A_gO8VDvG40_1;
	wire w_dff_A_JP3Ip3nE2_1;
	wire w_dff_A_VnwMUdos2_1;
	wire w_dff_A_rwbuN3lF2_2;
	wire w_dff_A_WutHriiW2_2;
	wire w_dff_B_xQFBRjFr0_2;
	wire w_dff_B_K3fr7C5p8_2;
	wire w_dff_B_NttktZYI2_2;
	wire w_dff_B_P4fo1Pmd8_2;
	wire w_dff_B_BaqOPZ646_2;
	wire w_dff_B_S7yHHKqo3_2;
	wire w_dff_B_HfrBjEFp6_2;
	wire w_dff_B_PJsAM0Am4_2;
	wire w_dff_B_tswFWHNN0_2;
	wire w_dff_A_pdGcakNm7_1;
	wire w_dff_A_ffwLEjuB8_1;
	wire w_dff_A_d3odaars2_1;
	wire w_dff_A_esJnoely4_1;
	wire w_dff_A_HlIqDWum0_1;
	wire w_dff_A_hho9pabx0_1;
	wire w_dff_A_wjyPR4Q55_1;
	wire w_dff_A_F0SmUnOV6_1;
	wire w_dff_A_Gghfwt0C2_1;
	wire w_dff_A_GfciHy3B3_1;
	wire w_dff_A_LefhVn3Z6_1;
	wire w_dff_A_WZyU70B86_1;
	wire w_dff_A_ySfB1G0n0_1;
	wire w_dff_A_ADSSagpo0_1;
	wire w_dff_A_K6f1eYEf2_2;
	wire w_dff_A_BRclw7Kc3_0;
	wire w_dff_A_kiNFkwt71_0;
	wire w_dff_A_jnlbi7kZ4_0;
	wire w_dff_A_Ru1gRn2Z3_0;
	wire w_dff_A_jSszOj0K5_0;
	wire w_dff_A_1HrCzaq51_0;
	wire w_dff_A_Kbxrl8Z16_0;
	wire w_dff_A_urhDNzTr3_0;
	wire w_dff_A_MMdQ1c6m6_0;
	wire w_dff_A_hIqyZcc48_0;
	wire w_dff_A_jIOBzIQ13_0;
	wire w_dff_A_xyxMXKFh7_0;
	wire w_dff_B_AOf3PMd74_1;
	wire w_dff_B_RSBxnL4w9_0;
	wire w_dff_B_fvTJbHeF9_0;
	wire w_dff_B_FcFEgFew3_0;
	wire w_dff_B_9ODYf6pV6_0;
	wire w_dff_A_aQ7HXJvB2_1;
	wire w_dff_A_MRlr7ald7_1;
	wire w_dff_A_J0qI5n7m6_1;
	wire w_dff_A_ALpZQIjD5_1;
	wire w_dff_A_JjHPO06u2_1;
	wire w_dff_B_6rqXqpJ01_2;
	wire w_dff_B_mwnP0hxW8_2;
	wire w_dff_B_KRKihJsA9_2;
	wire w_dff_B_fGNxAou53_2;
	wire w_dff_B_r2WXSA2G3_2;
	wire w_dff_B_x8jcFjAS6_0;
	wire w_dff_B_fdXgcZAc6_0;
	wire w_dff_B_63HPZrNT6_1;
	wire w_dff_B_Qwk5WDrA8_1;
	wire w_dff_B_eM51dZqn7_1;
	wire w_dff_A_CmsnOfjB2_1;
	wire w_dff_A_GOHXnMpZ8_1;
	wire w_dff_A_QrUn5Y1q2_1;
	wire w_dff_A_CoR02alG1_2;
	wire w_dff_A_oG4v0NJT1_2;
	wire w_dff_A_DF5FSiJD0_2;
	wire w_dff_A_rJR5CfaT1_2;
	wire w_dff_A_yikJDtD03_2;
	wire w_dff_A_Xkr6dqbD7_2;
	wire w_dff_A_SSqurgJA3_2;
	wire w_dff_B_5tBr8GmK5_3;
	wire w_dff_A_466xwsJd9_0;
	wire w_dff_A_3SyX6WOy6_0;
	wire w_dff_A_9ecManOQ7_0;
	wire w_dff_A_L64PkMmi3_0;
	wire w_dff_A_9VMwjoTv1_0;
	wire w_dff_A_eKYXsKcW3_0;
	wire w_dff_A_pDDuEHYq6_0;
	wire w_dff_A_38imH19D1_0;
	wire w_dff_A_g83TBW6C0_0;
	wire w_dff_B_GtX4MKB26_1;
	wire w_dff_A_IA24yFJu7_1;
	wire w_dff_A_BkPpqbEr6_0;
	wire w_dff_A_MQUS6LhM8_0;
	wire w_dff_A_OsDmPOrR7_0;
	wire w_dff_A_bqXPRDbF7_0;
	wire w_dff_A_AhheJNR09_0;
	wire w_dff_A_O7xdiAw80_0;
	wire w_dff_A_ROPVd4b70_0;
	wire w_dff_A_NABcI0GJ6_0;
	wire w_dff_A_mpgmD9Kb4_0;
	wire w_dff_A_dkW0DJwa4_2;
	wire w_dff_A_mkBWdZtU7_2;
	wire w_dff_A_zLgKIio29_2;
	wire w_dff_A_rIWb77up4_2;
	wire w_dff_A_edJapZXS5_2;
	wire w_dff_A_4o8dWzod0_2;
	wire w_dff_B_HkACRLua4_0;
	wire w_dff_B_EbanuIL94_1;
	wire w_dff_A_gIfxbOeB2_0;
	wire w_dff_A_W8bNgbnM3_0;
	wire w_dff_A_KMn58kOm9_0;
	wire w_dff_A_j9Cq96bD8_0;
	wire w_dff_A_lXQfBWHf5_0;
	wire w_dff_A_Mrsvtuqe3_0;
	wire w_dff_A_adanFM526_0;
	wire w_dff_A_o3SGJcYE7_0;
	wire w_dff_A_3gixdF4m1_0;
	wire w_dff_A_2UKq2RSX8_0;
	wire w_dff_A_4qExMfTp2_0;
	wire w_dff_A_5SPZsnnS9_0;
	wire w_dff_A_XMc8XPuB1_0;
	wire w_dff_B_aa12GdHb2_0;
	wire w_dff_B_lFMH0nP49_1;
	wire w_dff_A_wCzkzTI42_1;
	wire w_dff_A_kMCd1Vpa5_2;
	wire w_dff_A_sXGtEOkU8_2;
	wire w_dff_A_K8bEREo46_2;
	wire w_dff_A_OjVjRNuA3_2;
	wire w_dff_A_zlIap0zn3_2;
	wire w_dff_A_FEP2jJOW5_2;
	wire w_dff_A_3BiEFrMv1_2;
	wire w_dff_A_Uet3vZWn5_2;
	wire w_dff_A_8dmrSXMb2_2;
	wire w_dff_A_j7FfwYML2_2;
	wire w_dff_A_SZza9EIx1_2;
	wire w_dff_B_8Vk4FzSE9_1;
	wire w_dff_B_BVkNQ79x1_1;
	wire w_dff_B_1uHcbsMd7_0;
	wire w_dff_B_TNEGyBiS4_0;
	wire w_dff_B_l1uAx0AP2_0;
	wire w_dff_A_TVYzYBxD9_0;
	wire w_dff_A_MRAMZT0G8_0;
	wire w_dff_A_SNSIvQLJ8_0;
	wire w_dff_A_71H4QDix5_1;
	wire w_dff_A_A1l2JSGf8_1;
	wire w_dff_A_bAIxOVC57_1;
	wire w_dff_A_ieu9LqiI2_1;
	wire w_dff_B_sRRrq9fT4_0;
	wire w_dff_A_h4DbwCpQ5_0;
	wire w_dff_A_TV5Z6BNA5_2;
	wire w_dff_A_P6llDIia8_0;
	wire w_dff_B_ow5BU3l15_0;
	wire w_dff_A_rN5QuUBu0_0;
	wire w_dff_A_xnDHd5k14_0;
	wire w_dff_A_U47ZbNnc1_0;
	wire w_dff_A_VY8skPAt1_0;
	wire w_dff_A_0yb5aQ5q4_0;
	wire w_dff_A_B9B5aRkE4_0;
	wire w_dff_A_5wChciOM6_0;
	wire w_dff_A_ej0PMbLP8_0;
	wire w_dff_A_AYdZ9OPD3_0;
	wire w_dff_A_DoYuYt3o0_0;
	wire w_dff_A_FzmSQcjZ8_0;
	wire w_dff_A_YFG3IsSo3_2;
	wire w_dff_A_eUw2U2AD1_2;
	wire w_dff_A_DNcLtVZT6_2;
	wire w_dff_A_DrSCtFhK1_2;
	wire w_dff_A_A3LqPYKu4_2;
	wire w_dff_A_3DUO5WVG8_2;
	wire w_dff_A_cChJUGIa0_2;
	wire w_dff_A_TBhpKZhG1_2;
	wire w_dff_B_Utw847178_1;
	wire w_dff_B_fIkYYlr24_1;
	wire w_dff_B_q9lg12EA5_1;
	wire w_dff_B_gV0ujE1p6_1;
	wire w_dff_B_3ZUXkE3q4_1;
	wire w_dff_B_qOGmSgWp9_1;
	wire w_dff_B_cNPK8Tiq9_1;
	wire w_dff_B_0R7JY9iW9_1;
	wire w_dff_B_efuL0FT03_1;
	wire w_dff_B_dt5rETtL5_1;
	wire w_dff_B_B3RK3ujN2_1;
	wire w_dff_B_mNPRY81a1_1;
	wire w_dff_B_xkh3ej2l3_1;
	wire w_dff_B_354K2EW42_1;
	wire w_dff_B_xTDbuQrc6_1;
	wire w_dff_A_fMv0x7dt0_0;
	wire w_dff_A_KGO1f1I56_0;
	wire w_dff_A_s9lrbxa57_1;
	wire w_dff_A_rNSxHSxU8_1;
	wire w_dff_A_p56n7AdR3_1;
	wire w_dff_A_bbNVnxrp4_1;
	wire w_dff_A_enNF7sed7_1;
	wire w_dff_A_IYre53nc7_1;
	wire w_dff_A_FYFbEOeg7_0;
	wire w_dff_A_AT1Avun83_0;
	wire w_dff_A_umPSBfAm7_1;
	wire w_dff_A_eUL5RS502_1;
	wire w_dff_A_S2LToxqY5_1;
	wire w_dff_A_d3P4bKgJ3_1;
	wire w_dff_A_VbcRc7wU1_2;
	wire w_dff_A_YVKjARmo8_2;
	wire w_dff_A_5N4U0R7P9_0;
	wire w_dff_A_22LW2eOR1_0;
	wire w_dff_A_YUvWpXW59_0;
	wire w_dff_A_zQPB9WuL5_1;
	wire w_dff_A_jbpgR47I0_0;
	wire w_dff_A_6hgNxPZ11_2;
	wire w_dff_A_15kIWfyz3_0;
	wire w_dff_A_CyVrelK90_0;
	wire w_dff_A_PexqyRIy5_0;
	wire w_dff_A_pyxSFSNG2_0;
	wire w_dff_A_HwhzBRUb9_1;
	wire w_dff_A_uWtMHdEi7_1;
	wire w_dff_A_dFHUU87T3_2;
	wire w_dff_A_oIBi9uCt9_2;
	wire w_dff_A_OpERxBMY3_2;
	wire w_dff_A_dv9qDyKm0_2;
	wire w_dff_B_2GSH3u6a3_1;
	wire w_dff_A_wdTD53Z07_0;
	wire w_dff_A_iJNkOBcs6_2;
	wire w_dff_A_Q2Ystg7B1_1;
	wire w_dff_A_9zo8w2nC0_0;
	wire w_dff_A_2OpYfxyO8_0;
	wire w_dff_A_grOdrvAe0_0;
	wire w_dff_A_gseW7AfT9_0;
	wire w_dff_A_PsI6B1CX7_0;
	wire w_dff_A_gJrDnbTx0_0;
	wire w_dff_A_HBen2u2L4_0;
	wire w_dff_B_JemMZoOb4_1;
	wire w_dff_B_l1aSVjxa3_1;
	wire w_dff_A_229310Pj4_1;
	wire w_dff_A_nEKMBtUX7_1;
	wire w_dff_A_7pO45wdU2_1;
	wire w_dff_A_fEPYXVYS3_1;
	wire w_dff_A_XeoILYub2_1;
	wire w_dff_A_wDvfa1v54_1;
	wire w_dff_A_Ps483HaZ6_1;
	wire w_dff_A_viYBww8f6_1;
	wire w_dff_A_LuXkb1gQ3_1;
	wire w_dff_A_c55wTJCO0_1;
	wire w_dff_A_lxZmYScW6_1;
	wire w_dff_A_H20UwY2C7_1;
	wire w_dff_A_v533jOmM9_1;
	wire w_dff_A_W9shQgB82_1;
	wire w_dff_A_j6tD9JNz9_1;
	wire w_dff_A_YoCgkczG0_1;
	wire w_dff_A_p4dN46MK3_1;
	wire w_dff_A_GBdJ8qxM0_1;
	wire w_dff_A_eI23THGf9_2;
	wire w_dff_A_gVNAxhYM2_2;
	wire w_dff_A_XYLxVUDh7_2;
	wire w_dff_A_drA0dc717_2;
	wire w_dff_A_2GxEKn7v5_2;
	wire w_dff_A_tlY3woxf6_2;
	wire w_dff_A_zOM3h7rE3_2;
	wire w_dff_A_KMxa9F4G3_2;
	wire w_dff_A_8ld0AhPF6_2;
	wire w_dff_A_U2nEUDmM9_2;
	wire w_dff_A_hcffjs9U1_0;
	wire w_dff_A_ZDq3w5ma4_0;
	wire w_dff_B_7Zrzttfu0_1;
	wire w_dff_B_hfwAfqic5_1;
	wire w_dff_B_aN7DnGVD7_1;
	wire w_dff_B_MNXlIaF17_1;
	wire w_dff_A_Fn8Bdpbb4_1;
	wire w_dff_A_k31sob227_0;
	wire w_dff_A_JKwks8bX3_0;
	wire w_dff_A_86MfvnTh9_0;
	wire w_dff_A_Zlou7Hha4_0;
	wire w_dff_A_0SmFqPbu6_1;
	wire w_dff_A_wBrNA6kY6_1;
	wire w_dff_A_vgOyOihe1_1;
	wire w_dff_A_lS6kLNkC3_2;
	wire w_dff_A_ABaQaqS04_2;
	wire w_dff_A_F5NgWOo37_2;
	wire w_dff_A_pwLbgITt6_2;
	wire w_dff_A_Pix1T5Ii7_1;
	wire w_dff_A_2Z0K9zBT8_1;
	wire w_dff_B_5ZvWoKPI1_1;
	wire w_dff_B_a6IBdNjb5_1;
	wire w_dff_A_oRe2HLmT5_2;
	wire w_dff_B_l9V0R11f7_3;
	wire w_dff_A_tiWIMtFl5_0;
	wire w_dff_A_SyTGvP4b2_0;
	wire w_dff_A_YqbMMSiH2_0;
	wire w_dff_A_JNMCiPQM9_1;
	wire w_dff_B_5j4gjsAx5_1;
	wire w_dff_A_UjBQH0Zl5_1;
	wire w_dff_A_B8ChI9y29_1;
	wire w_dff_A_mVrS8o4v7_1;
	wire w_dff_A_VeZtSxbX9_2;
	wire w_dff_A_D7QHmD778_2;
	wire w_dff_A_Lm3Wb03d5_2;
	wire w_dff_A_fMakeybT3_0;
	wire w_dff_A_PQWTlDM18_2;
	wire w_dff_A_qVwVWVcQ5_1;
	wire w_dff_A_co0w1ynH1_2;
	wire w_dff_A_XxixcFjb6_2;
	wire w_dff_A_RkoxuewP3_1;
	wire w_dff_B_CKFMWMZG7_1;
	wire w_dff_B_vc2CbMzP1_1;
	wire w_dff_B_B0WxHOIX3_1;
	wire w_dff_B_nUiidziz7_1;
	wire w_dff_B_kgP3d0345_1;
	wire w_dff_A_ttX26wiQ4_0;
	wire w_dff_A_4sasHgEi3_0;
	wire w_dff_A_IGH3UTH66_0;
	wire w_dff_A_t3kZlWYQ2_1;
	wire w_dff_A_B9NRc5n21_1;
	wire w_dff_A_aEpA6uPn7_1;
	wire w_dff_A_scUGrfox5_1;
	wire w_dff_A_fwBz1ci64_1;
	wire w_dff_A_PYBRhA2j5_2;
	wire w_dff_A_LvCUOXXt4_2;
	wire w_dff_A_SDo89qRs2_2;
	wire w_dff_A_uICwoGZT6_0;
	wire w_dff_B_zavP2zuO7_1;
	wire w_dff_B_niiqv8J41_1;
	wire w_dff_A_ISTEQ5Zl6_0;
	wire w_dff_A_08cq8yE56_0;
	wire w_dff_A_xQReP0PA4_0;
	wire w_dff_A_lOm9er0S6_0;
	wire w_dff_A_vcbZ96Yk7_0;
	wire w_dff_A_KXyZwOVb4_1;
	wire w_dff_A_nQy1rt4A1_1;
	wire w_dff_A_Pxom4RSw4_1;
	wire w_dff_A_oa0EixC20_2;
	wire w_dff_A_9PnPWOgg8_2;
	wire w_dff_A_DFmdfCgD2_2;
	wire w_dff_A_dltZK1Z17_0;
	wire w_dff_A_W0RigKhz8_0;
	wire w_dff_A_CapWvRY64_1;
	wire w_dff_A_r1l9bUN20_0;
	wire w_dff_A_fPmmE3xD9_2;
	wire w_dff_A_e4wCn9PN4_1;
	wire w_dff_B_PWP6gSHG7_1;
	wire w_dff_B_Ycv7c5LF4_1;
	wire w_dff_A_yvXDm0ym2_0;
	wire w_dff_A_swV2kJDX7_2;
	wire w_dff_A_mrHgL0da5_2;
	wire w_dff_A_w0Ny0zwc1_0;
	wire w_dff_A_wIkX4I6r0_1;
	wire w_dff_A_37sMpk473_1;
	wire w_dff_A_rfAUD5jN9_1;
	wire w_dff_A_pg6AqhMU6_2;
	wire w_dff_A_8rATMYQt0_2;
	wire w_dff_A_kjapD70J7_1;
	wire w_dff_A_LHr0g24r7_2;
	wire w_dff_A_eIiTMP0c2_2;
	wire w_dff_A_QYCTBoZC8_2;
	wire w_dff_A_af19hOMD6_2;
	wire w_dff_A_BZOLwxXs5_2;
	wire w_dff_A_3cWjdMqw2_2;
	wire w_dff_A_wfSd7gzC5_2;
	wire w_dff_A_OuQiUOlc6_2;
	wire w_dff_A_xkSxuZlZ0_2;
	wire w_dff_A_7I1tCCSc0_2;
	wire w_dff_A_ZBsC8Br30_2;
	wire w_dff_A_Hlfz5tLw4_2;
	wire w_dff_A_64vyYzxK4_0;
	wire w_dff_A_sEBCiPbv9_0;
	wire w_dff_A_vVt0nama4_0;
	wire w_dff_A_nITTOkrd7_0;
	wire w_dff_A_OPJm0w7Y9_0;
	wire w_dff_A_ayovNCNM2_0;
	wire w_dff_A_PTUN5wli3_2;
	wire w_dff_A_r2h4RkPj9_2;
	wire w_dff_A_RFaQ96J16_2;
	wire w_dff_A_YOzNbAII1_2;
	wire w_dff_A_AY38Xu2F2_2;
	wire w_dff_A_U7VDY1450_2;
	wire w_dff_A_pGhWEDCn9_2;
	wire w_dff_A_uB5ORrbZ4_2;
	wire w_dff_A_CZaORwpN2_2;
	wire w_dff_A_pC2Mo1fT7_2;
	wire w_dff_A_khWV93EV6_2;
	wire w_dff_A_b2z9rtlA0_2;
	wire w_dff_A_W6o0McAd1_2;
	wire w_dff_A_8JDSD9gO1_2;
	wire w_dff_A_TUGSEb6r3_2;
	wire w_dff_A_CdOctyaS7_2;
	wire w_dff_A_KEAJMF1s8_2;
	wire w_dff_A_IMnGiKEn7_2;
	wire w_dff_A_dk9yo68N9_1;
	wire w_dff_A_04zl8Bxc6_1;
	wire w_dff_A_gbA2SURq8_1;
	wire w_dff_A_TVlTtE6r7_1;
	wire w_dff_A_4ym3sVNQ8_1;
	wire w_dff_A_Ag4lhDMZ7_1;
	wire w_dff_A_kIlvUKcO3_1;
	wire w_dff_A_mtxJGkWf4_1;
	wire w_dff_A_3F0yJgCq5_1;
	wire w_dff_A_1yFmmmqE0_1;
	wire w_dff_A_51HlVrDt5_1;
	wire w_dff_A_kNEKMNe02_1;
	wire w_dff_A_zI6r6zWP1_1;
	wire w_dff_A_bIKN2Bid9_1;
	wire w_dff_A_f2ED1Poh3_1;
	wire w_dff_A_q4v7VrV62_1;
	wire w_dff_A_HZx7zHi24_2;
	wire w_dff_A_QtZZ1elG6_2;
	wire w_dff_A_2P6TUELz8_2;
	wire w_dff_A_vLjItTvK2_2;
	wire w_dff_A_ROOgjzFz8_2;
	wire w_dff_A_5YMBjLyY9_2;
	wire w_dff_A_Amqs3Bit9_2;
	wire w_dff_B_6OeN7K636_1;
	wire w_dff_B_1L6o6Cko8_1;
	wire w_dff_B_ImqgfV7J8_1;
	wire w_dff_B_EtkgiWtu9_1;
	wire w_dff_B_cGk6N2sD5_1;
	wire w_dff_B_S3mB3zSa6_1;
	wire w_dff_B_CJd9RD5S0_1;
	wire w_dff_B_uVr5f8oh2_1;
	wire w_dff_B_2wz2D0Pr1_1;
	wire w_dff_B_8hrJ0wYW1_1;
	wire w_dff_B_R5F530526_1;
	wire w_dff_B_souuacIB0_1;
	wire w_dff_B_JRWM6lha9_1;
	wire w_dff_B_lyvI4CwF3_1;
	wire w_dff_B_4GmtljTw5_1;
	wire w_dff_B_76yLKDrR8_1;
	wire w_dff_B_Yx8Y5mBm5_1;
	wire w_dff_B_jNzKA38i4_1;
	wire w_dff_B_n3cs1FfX4_1;
	wire w_dff_B_EhJkZzbA4_0;
	wire w_dff_B_HS69KahT6_0;
	wire w_dff_B_ThUFz0mE9_0;
	wire w_dff_B_HnE2ciiS9_0;
	wire w_dff_B_93OsQDIC7_0;
	wire w_dff_B_H20Gu3l83_0;
	wire w_dff_B_A7CSZ7zs0_0;
	wire w_dff_B_hj6k4AW68_0;
	wire w_dff_B_LtaItCx80_0;
	wire w_dff_B_mBGTLlPb7_0;
	wire w_dff_B_hjTfYdzz3_0;
	wire w_dff_B_hmLUvkg22_0;
	wire w_dff_B_CIp1uF8m0_0;
	wire w_dff_B_tGGze2J71_0;
	wire w_dff_B_yCJCVwuc5_0;
	wire w_dff_B_2khqw2AR0_0;
	wire w_dff_B_gQ3HQZ7w5_0;
	wire w_dff_B_AsoKSNIU2_0;
	wire w_dff_B_88vVCwdc4_0;
	wire w_dff_B_Qf1PQoZZ5_1;
	wire w_dff_B_GncxnPhC1_1;
	wire w_dff_B_c4GH5yc22_1;
	wire w_dff_B_6zxqdXAJ4_1;
	wire w_dff_B_mcGzYXIk5_1;
	wire w_dff_B_L99eLpKe4_1;
	wire w_dff_B_Jrysdmbr7_1;
	wire w_dff_B_KSw97FQY9_1;
	wire w_dff_B_pKrQqRjP2_0;
	wire w_dff_B_5sQTU8zG9_0;
	wire w_dff_B_nhICFsvk8_1;
	wire w_dff_B_EtgMCAiT2_0;
	wire w_dff_B_WVLqhli38_0;
	wire w_dff_B_0qPXDqtW9_0;
	wire w_dff_B_I3DZOT0N9_0;
	wire w_dff_B_EVlwy7Ax0_1;
	wire w_dff_B_2MbpbnbB1_1;
	wire w_dff_B_J2KV0Fnw6_1;
	wire w_dff_B_0aGJ5bAa9_1;
	wire w_dff_B_1qJTC31r1_1;
	wire w_dff_B_2yjrLfHS5_1;
	wire w_dff_B_YeW9ImRd9_1;
	wire w_dff_B_3KhERs6R8_1;
	wire w_dff_B_1CoSnAiy8_1;
	wire w_dff_B_XdrxUKX55_1;
	wire w_dff_B_O9rHUWWP6_1;
	wire w_dff_B_ybm314OY6_1;
	wire w_dff_B_wBB2siGO4_1;
	wire w_dff_B_Pwv1sH3P1_1;
	wire w_dff_B_Y8zfDsM18_1;
	wire w_dff_B_sMf275Oj5_1;
	wire w_dff_B_CdlBZLKv8_1;
	wire w_dff_B_TB6HaPrd4_1;
	wire w_dff_B_6Th0vuFA4_1;
	wire w_dff_B_U2djDFY16_1;
	wire w_dff_B_2XTWqIPU0_1;
	wire w_dff_B_K30Kxw1G5_1;
	wire w_dff_B_To8vsBxy8_1;
	wire w_dff_A_VeQVEag42_0;
	wire w_dff_A_zx1Zjokm5_1;
	wire w_dff_B_5bPD11Zu0_2;
	wire w_dff_B_8f7Rwor92_2;
	wire w_dff_B_b8zsgBWp5_2;
	wire w_dff_B_Ro7kTiWC3_2;
	wire w_dff_A_xCxv6HKT2_0;
	wire w_dff_A_HUQ0FT1o3_0;
	wire w_dff_A_2Z8mXk8k5_0;
	wire w_dff_A_Z01nOi0E2_0;
	wire w_dff_A_xySRvejU7_1;
	wire w_dff_A_cq8EeuVL6_1;
	wire w_dff_B_Aqgco1yP8_1;
	wire w_dff_B_R3AsyGgd0_0;
	wire w_dff_B_2c3jPkB65_1;
	wire w_dff_A_kbnB72tY6_0;
	wire w_dff_A_jvBsZeVC2_0;
	wire w_dff_B_JwbTmWEP5_2;
	wire w_dff_B_bV4ITsi30_2;
	wire w_dff_B_PMsOGxPU2_2;
	wire w_dff_B_o6QtMK7q2_2;
	wire w_dff_B_XU6W4ozn0_2;
	wire w_dff_B_Dy6tX2Yq7_2;
	wire w_dff_B_zwWypTr77_0;
	wire w_dff_B_Owq66JFL6_0;
	wire w_dff_B_ulmeB7oI0_0;
	wire w_dff_B_yWXPpkU14_0;
	wire w_dff_B_Cxu0AvQP9_0;
	wire w_dff_B_SqxMVJQv9_0;
	wire w_dff_B_SWU0Og0K2_0;
	wire w_dff_B_F6fTFBFL8_0;
	wire w_dff_A_3ja49RM29_2;
	wire w_dff_A_wWqxvnFh5_2;
	wire w_dff_A_Gtb5rL9D6_2;
	wire w_dff_A_RHBgMXWQ6_2;
	wire w_dff_A_aj8ithYg8_2;
	wire w_dff_A_S6JWOdGf1_2;
	wire w_dff_A_WrZMAIQo0_2;
	wire w_dff_A_tc2FYKIM4_2;
	wire w_dff_A_OciTwPi61_2;
	wire w_dff_A_fHwo9xj71_2;
	wire w_dff_A_jmPxkNvb8_2;
	wire w_dff_A_YNBRqcRa7_2;
	wire w_dff_A_nHigQEHp3_1;
	wire w_dff_A_VEZ2Lyt87_1;
	wire w_dff_A_WC2N9Msk0_1;
	wire w_dff_A_YAC9j1oB7_1;
	wire w_dff_A_Dl0Ry4UP1_1;
	wire w_dff_A_0MglTAon8_1;
	wire w_dff_A_y2HKCHyV4_1;
	wire w_dff_A_0EKC9WTT4_1;
	wire w_dff_A_IhjvjxkU8_1;
	wire w_dff_A_tpeqpbPU1_2;
	wire w_dff_A_VbBdf96I2_2;
	wire w_dff_A_swWSomix1_2;
	wire w_dff_A_4WZEEWt28_2;
	wire w_dff_A_ic1Sd5dt8_2;
	wire w_dff_A_cisqXhkJ5_2;
	wire w_dff_A_Ad3UL6lH1_2;
	wire w_dff_A_QjPZEWqj8_2;
	wire w_dff_A_PFBHx6OY6_2;
	wire w_dff_B_blt8YHHv2_3;
	wire w_dff_B_ue2FJvjL9_3;
	wire w_dff_A_mWZi5Wvh4_1;
	wire w_dff_A_rt1CipLT7_1;
	wire w_dff_A_IMU7GyEl9_1;
	wire w_dff_A_Bi2zBv3k9_0;
	wire w_dff_B_xyvvpyID3_1;
	wire w_dff_B_QoISKYFR2_1;
	wire w_dff_B_Gw3mBlYD2_0;
	wire w_dff_B_RdkYRMhY3_1;
	wire w_dff_B_8MNPYt2H8_2;
	wire w_dff_A_MVAVHnvF7_0;
	wire w_dff_B_lJJhKMIC2_0;
	wire w_dff_B_OGZ3SmVF3_1;
	wire w_dff_A_4PZcCC7F9_1;
	wire w_dff_A_rU9nK9bv2_1;
	wire w_dff_A_N3VTAcw44_1;
	wire w_dff_A_PcBj3BQH4_1;
	wire w_dff_A_XcUoOKCH7_1;
	wire w_dff_A_X4NFrEQU5_1;
	wire w_dff_A_9kFtfxdw7_1;
	wire w_dff_A_Dt7atwku0_1;
	wire w_dff_A_vb0eqkuN8_1;
	wire w_dff_B_QCKE4Vj84_2;
	wire w_dff_B_njDmDYvj6_2;
	wire w_dff_B_rI3rDfQO6_2;
	wire w_dff_A_RcQxCNTJ4_0;
	wire w_dff_A_lJFZsVQE5_0;
	wire w_dff_A_PEsInGMZ2_0;
	wire w_dff_A_qojEt2kH7_0;
	wire w_dff_A_F0ZZ8ljA9_0;
	wire w_dff_B_EBnxoP7t6_1;
	wire w_dff_B_eO5eMZRj6_1;
	wire w_dff_B_LWCDxLKe9_0;
	wire w_dff_A_pEJMJpr07_0;
	wire w_dff_B_MniNMeSj0_0;
	wire w_dff_B_zyEKpJaB5_0;
	wire w_dff_A_1F8jFF1c1_0;
	wire w_dff_A_qfSiuZc81_0;
	wire w_dff_A_rBYzm1ut3_0;
	wire w_dff_A_PDsN4Y8C0_0;
	wire w_dff_A_HNJiObHX0_0;
	wire w_dff_A_RbbxnHEB6_0;
	wire w_dff_A_s3a2UhOY3_0;
	wire w_dff_A_rNtdnGCB4_1;
	wire w_dff_A_Pi97kgwG7_1;
	wire w_dff_A_bZmkYIdN2_1;
	wire w_dff_A_F5A5MZ505_1;
	wire w_dff_A_ixbpSxxm4_0;
	wire w_dff_A_Zn2BH9Cy0_0;
	wire w_dff_A_M3mLHJYX1_0;
	wire w_dff_A_CtxohyMF6_0;
	wire w_dff_A_PA9ynngi7_0;
	wire w_dff_A_0pE0wOE56_0;
	wire w_dff_B_TQvuXTWR4_2;
	wire w_dff_B_Vhp7DYjM5_2;
	wire w_dff_A_Rzp9MT8F9_0;
	wire w_dff_A_VyHLCHxB8_1;
	wire w_dff_A_giEofqP28_1;
	wire w_dff_A_9OAdvTyj2_1;
	wire w_dff_A_yfszB5K62_0;
	wire w_dff_A_a9ABx1MJ6_0;
	wire w_dff_A_nXjwNtcd7_0;
	wire w_dff_A_vaZlhGfN7_0;
	wire w_dff_A_G8o9lxgE4_0;
	wire w_dff_A_g5x9RPCW1_0;
	wire w_dff_A_cBTUSIlK9_0;
	wire w_dff_A_Kq47wWt17_0;
	wire w_dff_A_cgE24JCS8_0;
	wire w_dff_A_IJB7r4Tb8_0;
	wire w_dff_A_3LWJ42QH3_0;
	wire w_dff_A_QIPZdZ9U2_0;
	wire w_dff_A_0YIluyBg5_2;
	wire w_dff_A_x5RSzLg95_2;
	wire w_dff_A_KlZqlUxc6_2;
	wire w_dff_A_tjtZVJ2u2_2;
	wire w_dff_A_1N9g9ILt1_2;
	wire w_dff_A_UwO2FDe47_2;
	wire w_dff_A_0kENtmZp5_2;
	wire w_dff_A_017YlmjG8_2;
	wire w_dff_A_GzSCvmyJ9_2;
	wire w_dff_A_gmdSfpsv8_2;
	wire w_dff_B_FboPHIRO5_1;
	wire w_dff_B_RUghDjnJ6_1;
	wire w_dff_B_hrQg93Qp0_1;
	wire w_dff_B_15CS6bYn4_1;
	wire w_dff_B_T1NSR8jE9_1;
	wire w_dff_B_iF0KyPtM9_1;
	wire w_dff_B_tgCupd6O2_1;
	wire w_dff_B_2VIl7vl08_1;
	wire w_dff_B_Uc3tdeoM0_1;
	wire w_dff_A_YAqQIAnL3_1;
	wire w_dff_A_evSASmTu6_0;
	wire w_dff_A_kGXM6RqT9_0;
	wire w_dff_A_yuFEVChI9_1;
	wire w_dff_A_7pXUF9fR4_1;
	wire w_dff_A_Plj7rlTI0_1;
	wire w_dff_A_qDDp2ip11_1;
	wire w_dff_A_5IIaAJoR1_2;
	wire w_dff_A_SRrG980J0_2;
	wire w_dff_A_gTlyjfpT1_2;
	wire w_dff_A_z8mKH3gn7_1;
	wire w_dff_A_m1AaSk9P7_1;
	wire w_dff_A_OkQ4V4ul0_0;
	wire w_dff_A_nMug4MFz8_0;
	wire w_dff_A_aNeRiGDk3_0;
	wire w_dff_A_Q8688C4e3_1;
	wire w_dff_B_n06xFyHa9_2;
	wire w_dff_A_quGm9qOq7_0;
	wire w_dff_A_R7x0xSWu1_1;
	wire w_dff_A_y24sHRf73_1;
	wire w_dff_A_vDwub33C8_1;
	wire w_dff_A_mMhdil6U0_1;
	wire w_dff_A_AHYVuzOx6_1;
	wire w_dff_B_sgRjECoX8_1;
	wire w_dff_B_XMxOAZNd4_1;
	wire w_dff_B_udTWXWny9_2;
	wire w_dff_B_UtgxsUNu9_2;
	wire w_dff_B_JPFUb9cB6_2;
	wire w_dff_B_tFhesDRj6_2;
	wire w_dff_B_L9ZMFgnB6_2;
	wire w_dff_B_1pShMc1D2_2;
	wire w_dff_B_Dkqd5guL7_2;
	wire w_dff_B_WknH7xHK3_2;
	wire w_dff_B_Fg5lBWpv4_2;
	wire w_dff_B_kuwmshAL9_2;
	wire w_dff_A_Ysk3cZVl4_2;
	wire w_dff_A_dm6gyHFT9_2;
	wire w_dff_A_TDrrSPXo7_2;
	wire w_dff_A_FskTuqoE1_2;
	wire w_dff_A_legCigtL3_2;
	wire w_dff_A_gyPtAf1f2_1;
	wire w_dff_A_Ssov5t7J6_1;
	wire w_dff_A_JScAPa3A8_1;
	wire w_dff_A_HJZTXVlc5_1;
	wire w_dff_A_5fld2Bhh1_1;
	wire w_dff_A_dkZK43yW7_1;
	wire w_dff_A_H8aPmCPQ7_1;
	wire w_dff_B_SyGdP9t01_0;
	wire w_dff_A_MVqbkzH00_0;
	wire w_dff_B_zXsy4sDE9_1;
	wire w_dff_A_E2vqs1Gz9_0;
	wire w_dff_A_Rx7my7XR1_0;
	wire w_dff_A_F72lr6t99_1;
	wire w_dff_A_OYI0EwiM0_1;
	wire w_dff_A_SVbnN9s24_1;
	wire w_dff_A_TlknoW6D7_1;
	wire w_dff_A_EmzmYA7F1_1;
	wire w_dff_A_IsFo5hR41_1;
	wire w_dff_A_FS1dtY4e7_1;
	wire w_dff_A_bKObz1oh2_1;
	wire w_dff_A_qdG8UMs30_1;
	wire w_dff_A_tTROXtQE4_1;
	wire w_dff_A_VaI15jXt6_1;
	wire w_dff_A_irDksPBB8_1;
	wire w_dff_A_QjppZzxw4_1;
	wire w_dff_A_2NXqZb9L5_1;
	wire w_dff_A_0Rqlm6JO6_1;
	wire w_dff_A_BIFyI2Ba4_1;
	wire w_dff_B_jK6rhq0e3_0;
	wire w_dff_B_gwnaqesO9_1;
	wire w_dff_A_f7lUCiew2_0;
	wire w_dff_A_giWd21D36_2;
	wire w_dff_A_8oKXciT03_1;
	wire w_dff_A_T5WUaTeX7_1;
	wire w_dff_A_rqE1AeFv5_1;
	wire w_dff_A_J7TlupEE3_1;
	wire w_dff_A_vyzf7wGv7_1;
	wire w_dff_A_aW4fAWQe5_1;
	wire w_dff_A_8AIJ25oZ5_1;
	wire w_dff_A_5Q8c7W6x3_1;
	wire w_dff_A_PWdd2DEy6_1;
	wire w_dff_A_8PrYpk353_1;
	wire w_dff_A_S5lETVX55_1;
	wire w_dff_A_fiYCsWVX3_1;
	wire w_dff_A_s7dU7DEJ4_1;
	wire w_dff_A_hQMLIAPg0_1;
	wire w_dff_A_Xrkgt8Uq2_1;
	wire w_dff_A_QzXpiAQL1_1;
	wire w_dff_A_UfmvrRkC4_1;
	wire w_dff_A_hzxSu0t47_2;
	wire w_dff_A_PlNFSRZF0_2;
	wire w_dff_A_WB2Uv4N09_2;
	wire w_dff_A_QuvMuqkL5_2;
	wire w_dff_A_pEF531yR7_2;
	wire w_dff_A_2Iy5PONt3_2;
	wire w_dff_A_v0uVrX126_2;
	wire w_dff_A_JuSmpmgD2_2;
	wire w_dff_A_HsNOgYfh5_2;
	wire w_dff_A_xthy18NE9_2;
	wire w_dff_A_t40zNYXZ9_2;
	wire w_dff_A_nQRxAP3K2_2;
	wire w_dff_A_K5oSnFpI3_2;
	wire w_dff_A_zpJyU6uJ7_2;
	wire w_dff_A_GZprBdzv7_2;
	wire w_dff_A_EfOBnjDB0_2;
	wire w_dff_A_Zs4y31Dq2_2;
	wire w_dff_A_zg1pibig3_2;
	wire w_dff_A_3geM0Cms6_2;
	wire w_dff_A_txTqEs2L8_2;
	wire w_dff_A_HGT1TjPl5_2;
	wire w_dff_A_1RahILR75_2;
	wire w_dff_A_yg7oj4gc8_2;
	wire w_dff_A_7NfPz0Xh7_2;
	wire w_dff_A_DaipWDjI3_2;
	wire w_dff_A_2isySGdC3_2;
	wire w_dff_A_4XKB28U33_2;
	wire w_dff_B_tFWjCfY76_2;
	wire w_dff_B_ypoCYK9M4_1;
	wire w_dff_B_9VCie3KC0_1;
	wire w_dff_A_W71XNuJJ0_0;
	wire w_dff_A_RIOyuKSd2_2;
	wire w_dff_A_AYrARYnc4_2;
	wire w_dff_A_tpZMpNCi1_0;
	wire w_dff_A_IBV2KcPm6_0;
	wire w_dff_A_KdrmsbCd1_1;
	wire w_dff_A_k47UJfMu3_1;
	wire w_dff_A_LzTv22fS0_2;
	wire w_dff_B_3IdeH9Np3_1;
	wire w_dff_B_acLe9BB14_1;
	wire w_dff_A_BuHAXN7I3_2;
	wire w_dff_A_cR87xW9l6_2;
	wire w_dff_B_9tSn0Y3k1_3;
	wire w_dff_B_hmWGLqJC7_1;
	wire w_dff_A_AHWfAdJj2_1;
	wire w_dff_A_EXVkxyFG1_0;
	wire w_dff_A_8QLBYNJY8_0;
	wire w_dff_A_emFgZITx2_1;
	wire w_dff_A_WQTppcFP4_0;
	wire w_dff_B_FBmqfDmr8_1;
	wire w_dff_B_MuDZpq9d7_1;
	wire w_dff_A_XBsqqt4V8_0;
	wire w_dff_A_g7GwuWCI6_2;
	wire w_dff_A_KKnWbrl30_2;
	wire w_dff_A_epP7q5ez9_0;
	wire w_dff_A_GiVZV48h2_1;
	wire w_dff_A_3gDDM7YM7_1;
	wire w_dff_A_2BKmGxKs5_2;
	wire w_dff_A_tgC1v8gX3_2;
	wire w_dff_A_6TXoc7rK1_2;
	wire w_dff_A_Nvzu5XCg3_0;
	wire w_dff_A_VmEvoykn8_2;
	wire w_dff_B_TnDCwe8l9_1;
	wire w_dff_B_0XVfhXz86_1;
	wire w_dff_A_hcaBnGNJ4_0;
	wire w_dff_A_dkRzf9Fo3_2;
	wire w_dff_A_aL3GOddb6_2;
	wire w_dff_A_6NnZ85746_0;
	wire w_dff_A_uzHU8Ycj9_0;
	wire w_dff_A_zxoV718G2_1;
	wire w_dff_A_5f3YffZc9_0;
	wire w_dff_A_i4yijk0O8_2;
	wire w_dff_B_1P3BHLgR7_1;
	wire w_dff_B_RzIglBOu5_1;
	wire w_dff_B_9WJTBuJM3_1;
	wire w_dff_B_Dbht9dBE8_1;
	wire w_dff_A_EizV1JxL4_1;
	wire w_dff_A_cjga727m6_1;
	wire w_dff_A_DSYuGwNq6_0;
	wire w_dff_A_utIED0WE2_0;
	wire w_dff_A_yQ2rIpMw1_0;
	wire w_dff_A_sWDiBuh02_0;
	wire w_dff_A_JUV4H6lN0_2;
	wire w_dff_A_siA6kNFd3_2;
	wire w_dff_A_TRyHePPu3_1;
	wire w_dff_A_UBKQ6Prb5_2;
	wire w_dff_B_VwSpmpmP0_1;
	wire w_dff_B_ft2Gh3C70_1;
	wire w_dff_B_nQshTVjR8_2;
	wire w_dff_A_Rg98vPlY4_0;
	wire w_dff_A_vZnYrOku2_0;
	wire w_dff_A_zPwGSvjv5_0;
	wire w_dff_A_ePZeCHJY0_1;
	wire w_dff_B_nEin9Box4_1;
	wire w_dff_A_5rnoyF4a9_1;
	wire w_dff_A_BKcFDSnW7_1;
	wire w_dff_A_gU7880GW8_1;
	wire w_dff_A_3ddKH4RU8_2;
	wire w_dff_A_EqCpre9Y7_2;
	wire w_dff_A_F12oIkZY4_2;
	wire w_dff_A_7sPGyeUk4_0;
	wire w_dff_B_XAClLi7a5_1;
	wire w_dff_B_ObJKJAL65_1;
	wire w_dff_B_VElSIzjE4_2;
	wire w_dff_A_3BiR3btB8_0;
	wire w_dff_B_bhkwObJ23_1;
	wire w_dff_A_uazgisl77_1;
	wire w_dff_A_hmoDB3ZB7_0;
	wire w_dff_A_XJZbC1zp8_0;
	wire w_dff_A_u7SX3Bg06_0;
	wire w_dff_A_VwRRsoqh0_2;
	wire w_dff_A_3mpWkusM1_2;
	wire w_dff_A_FkEO5EKi9_1;
	wire w_dff_A_8ErAXYhy7_2;
	wire w_dff_A_oh0mZN6n0_1;
	wire w_dff_A_UvE4980e5_2;
	wire w_dff_A_UIM1XxVP6_0;
	wire w_dff_B_mmaQjxYO6_1;
	wire w_dff_B_Vte1rW7f8_1;
	wire w_dff_A_vBnwzuFg4_0;
	wire w_dff_A_gbBNtmKH0_0;
	wire w_dff_A_etOclqIw0_0;
	wire w_dff_A_YeycLRNs9_0;
	wire w_dff_A_sl8a1jJF6_1;
	wire w_dff_A_5acy51VL2_1;
	wire w_dff_A_SLdMtM8b8_1;
	wire w_dff_A_d3aCecw68_1;
	wire w_dff_A_YcZ4Jqcu3_1;
	wire w_dff_A_mw3Zve2w6_1;
	wire w_dff_A_Yi7meXIa0_2;
	wire w_dff_A_tol8jPOT1_2;
	wire w_dff_A_8xvh3C4x5_2;
	wire w_dff_A_fLq7odAN5_2;
	wire w_dff_A_Iri93B0L9_0;
	wire w_dff_B_cQGu051n7_1;
	wire w_dff_B_gleghccY1_1;
	wire w_dff_A_WP939Db63_0;
	wire w_dff_A_m8xX8rCk2_1;
	wire w_dff_A_cJfO8GK75_1;
	wire w_dff_A_hCUj84rT2_2;
	wire w_dff_A_DcYzTp8C6_2;
	wire w_dff_A_eoHESROo4_1;
	wire w_dff_A_yes0HgDd1_1;
	wire w_dff_A_kgki6oiX8_1;
	wire w_dff_A_3aaz8XkD0_1;
	wire w_dff_A_4vYs8wAb7_2;
	wire w_dff_A_1TuDV9NO0_0;
	wire w_dff_A_EgU4L2EN6_0;
	wire w_dff_A_ffFxNKV48_0;
	wire w_dff_A_Jgsa7gf44_0;
	wire w_dff_A_8PTPxEZU2_1;
	wire w_dff_A_eMy77nlV4_1;
	wire w_dff_A_KBCP7C4J6_1;
	wire w_dff_A_1UlOwWN55_2;
	wire w_dff_A_SAia8h8T3_2;
	wire w_dff_A_aieTzyUI2_2;
	wire w_dff_A_5srVuwcl4_2;
	wire w_dff_A_KEFDYI724_1;
	wire w_dff_A_UWfb0VmV7_2;
	wire w_dff_A_kc6Gp8Ba3_0;
	wire w_dff_A_xxiY3hzF4_2;
	wire w_dff_A_viGpsNUS2_0;
	wire w_dff_A_73wzFBMd0_0;
	wire w_dff_A_eusntHHy5_0;
	wire w_dff_A_ef7UMty77_0;
	wire w_dff_A_YSEkqc135_0;
	wire w_dff_A_BBXnGp3V1_0;
	wire w_dff_A_F0NkKZMh2_0;
	wire w_dff_A_xZchiVRd2_0;
	wire w_dff_A_f6xoYpup5_0;
	wire w_dff_A_MpgP6oaC4_0;
	wire w_dff_A_I4mWuMdI9_0;
	wire w_dff_A_X5iFbqWZ6_1;
	wire w_dff_A_paExvVgh1_0;
	wire w_dff_A_z9T9hpxY0_0;
	wire w_dff_A_UKZDXthg8_0;
	wire w_dff_A_xmJ00wV22_0;
	wire w_dff_A_yV3IXiGf0_0;
	wire w_dff_A_m54Pr7NK1_0;
	wire w_dff_A_WnuzEvYQ9_0;
	wire w_dff_A_uA2oguuJ4_2;
	wire w_dff_A_Z8XlFiam4_2;
	wire w_dff_A_V2vDih6Z4_2;
	wire w_dff_A_B3VACOQO5_2;
	wire w_dff_A_YdI9tNGe6_2;
	wire w_dff_A_25CNjiae8_2;
	wire w_dff_A_GA86mqIH2_2;
	wire w_dff_A_OXYgzVS37_2;
	wire w_dff_A_rSPrbVlt1_2;
	wire w_dff_A_P7dYRDUJ9_2;
	wire w_dff_A_yj4tkaQ32_2;
	wire w_dff_A_eqbKIpKc0_2;
	wire w_dff_A_NxKFlP6E5_2;
	wire w_dff_A_KpIEWaYu1_2;
	wire w_dff_A_cA8amEaP6_2;
	wire w_dff_A_0IEw0WLI3_2;
	wire w_dff_A_a9MBk0zK8_2;
	wire w_dff_A_jMDahzlB6_2;
	wire w_dff_A_EYUNAq5J7_2;
	wire w_dff_A_U9LGVDfH9_1;
	wire w_dff_A_pqBhYW279_1;
	wire w_dff_A_1tJYaH7l4_1;
	wire w_dff_A_0x5ZJo1h4_1;
	wire w_dff_A_8lB0GH520_1;
	wire w_dff_A_CFa9rKFI5_1;
	wire w_dff_A_bmZURhFr1_1;
	wire w_dff_A_Eri2EBMQ1_1;
	wire w_dff_A_ZCRpgCFQ0_1;
	wire w_dff_A_IljkbICw2_1;
	wire w_dff_A_eK0j9ZaM5_1;
	wire w_dff_A_UyraIZti2_1;
	wire w_dff_A_KcEHa6Yr4_1;
	wire w_dff_A_bH6cEhzw1_1;
	wire w_dff_A_mOFV86Bz2_1;
	wire w_dff_A_1Ox31FK61_1;
	wire w_dff_A_XUckKp2H8_1;
	wire w_dff_A_8Ep4cE458_2;
	wire w_dff_A_NBBAmwgZ2_2;
	wire w_dff_A_buy3CmPo8_2;
	wire w_dff_A_BFHhjxBJ5_2;
	wire w_dff_A_Dyiuatp05_2;
	wire w_dff_A_WAXdgUYi1_2;
	wire w_dff_A_LCgryU6H4_2;
	wire w_dff_A_mBeDuA271_2;
	wire w_dff_A_XWAPLWbL5_2;
	wire w_dff_A_ui7oAtrb7_2;
	wire w_dff_A_9XPHNBBU0_2;
	wire w_dff_A_sIWnwDEh7_1;
	wire w_dff_A_FgyHJt2a3_2;
	wire w_dff_B_I4fAPK9e7_2;
	wire w_dff_B_4H455TCA6_2;
	wire w_dff_B_ZZ47TlVM0_2;
	wire w_dff_B_dRf9BErv4_2;
	wire w_dff_B_STXNS9JG9_2;
	wire w_dff_B_XASqlK6q9_2;
	wire w_dff_B_BlCSfxRv7_2;
	wire w_dff_B_JUaKTUWs0_2;
	wire w_dff_B_82I58rjp0_2;
	wire w_dff_B_Mvh5p9V32_2;
	wire w_dff_B_D3YV7bYd5_2;
	wire w_dff_B_6zTa0c6n0_2;
	wire w_dff_B_F2GTTvIS0_2;
	wire w_dff_B_yjTMlEDO2_2;
	wire w_dff_B_xN6DHAUf0_2;
	wire w_dff_B_lzCdJ9k40_2;
	wire w_dff_B_nHxI0s1Y8_2;
	wire w_dff_B_E3zpKwOW7_2;
	wire w_dff_B_uOSiCRB66_2;
	wire w_dff_B_yrnmnuY47_2;
	wire w_dff_B_YYSXf3Cw1_2;
	wire w_dff_B_Y8KiCjfk3_2;
	wire w_dff_B_qJRpuyjt6_2;
	wire w_dff_B_SUr3R1MO3_2;
	wire w_dff_A_Er0lPOGE3_2;
	wire w_dff_A_JSk4D0w16_2;
	wire w_dff_A_0o1yUlot0_2;
	wire w_dff_A_eyin0HN03_2;
	wire w_dff_A_gZs5dwrj8_2;
	wire w_dff_A_9UTA3UMW8_2;
	wire w_dff_A_ixkDvfLk6_2;
	wire w_dff_A_X7PDkg0r9_2;
	wire w_dff_A_aYbBW02x0_2;
	wire w_dff_A_tTdMNgQg1_2;
	wire w_dff_A_HiGLvP440_2;
	wire w_dff_A_8v3DeU6y5_2;
	wire w_dff_A_Ohp9CgnO1_2;
	wire w_dff_A_eSsG7fWD5_2;
	wire w_dff_A_ZGCSzzn94_2;
	wire w_dff_A_KZHb8zjT1_2;
	wire w_dff_A_KTxw2vow3_2;
	wire w_dff_A_SRCD7BNj2_2;
	wire w_dff_A_pKCtvoOt9_2;
	wire w_dff_A_o9V2RABJ1_2;
	wire w_dff_A_KOoTQLek9_2;
	wire w_dff_A_IntbbyyG8_2;
	wire w_dff_A_vbqnXyDv5_2;
	wire w_dff_A_URHU4IuH9_0;
	wire w_dff_A_uu1NyUgA1_0;
	wire w_dff_A_aIBjR3T21_0;
	wire w_dff_A_H8jccFVF9_0;
	wire w_dff_A_fFriHcp03_0;
	wire w_dff_A_qiJpGME05_0;
	wire w_dff_A_tpzyB56f6_0;
	wire w_dff_A_Tj6fM6md4_0;
	wire w_dff_A_klsyIl0w4_0;
	wire w_dff_A_XpyP0Agr4_0;
	wire w_dff_A_EUchdzbn9_0;
	wire w_dff_A_Z0RAvOnB2_0;
	wire w_dff_A_A9U70sOV4_0;
	wire w_dff_A_tbZV8FCz1_0;
	wire w_dff_A_TqW5byGS9_0;
	wire w_dff_A_w46tlnWm0_0;
	wire w_dff_A_EZFj4lep1_1;
	wire w_dff_A_DzxPqTsI9_1;
	wire w_dff_A_EcQsoT9g3_1;
	wire w_dff_A_Nyiiwyuu1_1;
	wire w_dff_A_R2AOgfTK1_1;
	wire w_dff_A_CKvgTkiE3_1;
	wire w_dff_A_jvrLVt7O3_1;
	wire w_dff_A_gcqKeMoa8_1;
	wire w_dff_A_ggVqkWvU9_1;
	wire w_dff_A_i1Rasi4v5_1;
	wire w_dff_A_ZmlcfrZO8_1;
	wire w_dff_A_EBC8N9T79_1;
	wire w_dff_A_js2yMspE4_0;
	wire w_dff_A_ETMMXGaF0_0;
	wire w_dff_A_J4U27oSg2_0;
	wire w_dff_A_yw8o5U4R2_0;
	wire w_dff_A_tJc0cKRv9_0;
	wire w_dff_A_rZAseHNZ2_0;
	wire w_dff_A_VBTPSrG00_0;
	wire w_dff_A_9fyArUqG1_0;
	wire w_dff_A_uvRscf898_0;
	wire w_dff_A_przgP03g2_0;
	wire w_dff_A_swLddxws3_0;
	wire w_dff_A_nam4BOlK4_0;
	wire w_dff_A_ohgHWyp62_0;
	wire w_dff_A_Nx0DBZ8l6_0;
	wire w_dff_A_ovoHPIdI6_0;
	wire w_dff_A_vm0Sb9pr3_0;
	wire w_dff_A_wb4zkTA16_0;
	wire w_dff_A_GPiQ5TuP8_0;
	wire w_dff_A_3Jvt1A2P3_0;
	wire w_dff_A_a8ceP99Q8_0;
	wire w_dff_A_UIbrAWwd8_0;
	wire w_dff_A_fnZgtWOm9_0;
	wire w_dff_A_8VO7QJRY0_0;
	wire w_dff_A_8iXvTUpm7_0;
	wire w_dff_A_4dUJQMso6_0;
	wire w_dff_A_kk7cd6j65_1;
	wire w_dff_A_Afz9WXRJ5_0;
	wire w_dff_A_QTfMMhmG7_0;
	wire w_dff_A_UwQjHgiN5_0;
	wire w_dff_A_6fDo3UPn2_0;
	wire w_dff_A_2ci3SdFX7_0;
	wire w_dff_A_cll7EyyK5_0;
	wire w_dff_A_z3lprCox2_0;
	wire w_dff_A_IjdktLEQ4_0;
	wire w_dff_A_QkR49ma34_0;
	wire w_dff_A_6KvwVae57_0;
	wire w_dff_A_ZDRkilbs7_0;
	wire w_dff_A_9J2KbRkJ1_0;
	wire w_dff_A_erEWjDxi5_0;
	wire w_dff_A_WYboSFBI7_0;
	wire w_dff_A_51ysUhir2_0;
	wire w_dff_A_OwtHNWEa3_0;
	wire w_dff_A_potMbMC38_0;
	wire w_dff_A_gZb5bDv29_0;
	wire w_dff_A_8iW0Sl4i6_0;
	wire w_dff_A_dapypv925_0;
	wire w_dff_A_oRvrw7KV7_0;
	wire w_dff_A_kKNB3afA4_0;
	wire w_dff_A_A0f1L1Lt5_0;
	wire w_dff_A_afSXXLl07_0;
	wire w_dff_A_TK4XX8yx8_0;
	wire w_dff_A_a27FDOlD2_1;
	wire w_dff_A_7kA1e56U5_0;
	wire w_dff_A_dpgSKpl85_0;
	wire w_dff_A_DMyUoc0k3_0;
	wire w_dff_A_vXrsnBNS9_0;
	wire w_dff_A_FjUPWESn4_0;
	wire w_dff_A_JlvJ4awX3_0;
	wire w_dff_A_RfMBeTad3_0;
	wire w_dff_A_lyYrReaj8_0;
	wire w_dff_A_p6NWMAvP8_0;
	wire w_dff_A_ktLqLAGX5_0;
	wire w_dff_A_nsKCijmv8_0;
	wire w_dff_A_LHIomuu80_0;
	wire w_dff_A_6wFpFbRk4_0;
	wire w_dff_A_rcvUU5IZ6_0;
	wire w_dff_A_8qSdgszb4_0;
	wire w_dff_A_yFexwtY77_0;
	wire w_dff_A_xda3Vy0d6_0;
	wire w_dff_A_qzY6k9bV1_0;
	wire w_dff_A_LmZ0mUY13_0;
	wire w_dff_A_itLtmvNN7_0;
	wire w_dff_A_ljAecS813_0;
	wire w_dff_A_xXPOArSh9_0;
	wire w_dff_A_jendyGrO6_0;
	wire w_dff_A_f7A6Kc5N3_0;
	wire w_dff_A_ZmdUGqAM2_0;
	wire w_dff_A_x1fDTMpv4_1;
	wire w_dff_A_3eJkcZNv9_0;
	wire w_dff_A_X9tajY7k8_0;
	wire w_dff_A_xA0mRPKS0_0;
	wire w_dff_A_rLehVRFX3_0;
	wire w_dff_A_etlAf4X79_0;
	wire w_dff_A_64z72IBX9_0;
	wire w_dff_A_mh6W16JF8_0;
	wire w_dff_A_Fm2SPi825_0;
	wire w_dff_A_Qp7NrPNx3_0;
	wire w_dff_A_ZJ9sOzGb5_0;
	wire w_dff_A_oG8MZvNo1_0;
	wire w_dff_A_yguufseH2_0;
	wire w_dff_A_9yPlCXyn4_0;
	wire w_dff_A_Yo1dwklH7_0;
	wire w_dff_A_7BLirZBO5_0;
	wire w_dff_A_oqmu97qb3_0;
	wire w_dff_A_MDSAPr0g9_0;
	wire w_dff_A_e3wYAzRF4_0;
	wire w_dff_A_QoQM8ycS2_0;
	wire w_dff_A_FMf0Y2x02_0;
	wire w_dff_A_O69NHFZw0_0;
	wire w_dff_A_EfjyputL3_0;
	wire w_dff_A_RAJk3tgW3_0;
	wire w_dff_A_17NypG9V3_0;
	wire w_dff_A_Md6sOKZ80_1;
	wire w_dff_A_XvKxEYeb3_0;
	wire w_dff_A_i3XhF68D7_0;
	wire w_dff_A_8xqEaYYx2_0;
	wire w_dff_A_jtvLgiD99_0;
	wire w_dff_A_iXZdZlzp7_0;
	wire w_dff_A_XlzTt09d7_0;
	wire w_dff_A_HktJ1QZd2_0;
	wire w_dff_A_47HNa0811_0;
	wire w_dff_A_syDUelsQ0_0;
	wire w_dff_A_152ntPtq1_0;
	wire w_dff_A_IdCc1g4u1_0;
	wire w_dff_A_nMrDRXjR8_0;
	wire w_dff_A_1CQ8pp6U0_0;
	wire w_dff_A_b7PLKkUf2_0;
	wire w_dff_A_OPoYeikb9_0;
	wire w_dff_A_0lGNWpoZ8_0;
	wire w_dff_A_orosTVSG8_0;
	wire w_dff_A_Mb4puldy6_0;
	wire w_dff_A_LRDgmMRD0_0;
	wire w_dff_A_FJsbvNw90_0;
	wire w_dff_A_DQmwjfCt4_0;
	wire w_dff_A_HRGuZvis1_0;
	wire w_dff_A_DCOAnzVo8_0;
	wire w_dff_A_mybCOiNB9_0;
	wire w_dff_A_95yRjwe90_1;
	wire w_dff_A_NGnFQ2mj3_0;
	wire w_dff_A_Df8ddHxv7_0;
	wire w_dff_A_Q92jIBqk5_0;
	wire w_dff_A_NKYpk9oX1_0;
	wire w_dff_A_T0RH3nWO7_0;
	wire w_dff_A_zalk2Z9V1_0;
	wire w_dff_A_lpdgsik56_0;
	wire w_dff_A_YZTgR7Uj7_0;
	wire w_dff_A_ZDRfD1Ay2_0;
	wire w_dff_A_PNqNJOAs8_0;
	wire w_dff_A_kkFJ5V7M9_0;
	wire w_dff_A_rEzTzose3_0;
	wire w_dff_A_ONqr2cy19_0;
	wire w_dff_A_K1mUvgZK7_0;
	wire w_dff_A_hHnvlRYC9_0;
	wire w_dff_A_fKJnZX4L7_0;
	wire w_dff_A_DpPOdRXR4_0;
	wire w_dff_A_QpbcdHhU9_0;
	wire w_dff_A_0Jh4CTBc1_0;
	wire w_dff_A_stYB7YaL3_0;
	wire w_dff_A_AGBLizWo8_0;
	wire w_dff_A_pK6j8JNo6_0;
	wire w_dff_A_L1JQmsCW1_0;
	wire w_dff_A_xTZ1dCBt8_0;
	wire w_dff_A_AtXnEyBC7_1;
	wire w_dff_A_FouQWFaB4_0;
	wire w_dff_A_5ZHZUS7M6_0;
	wire w_dff_A_GmgpDGDR2_0;
	wire w_dff_A_PriqH0wm6_0;
	wire w_dff_A_sMmzXXj41_0;
	wire w_dff_A_Wl47g9D92_0;
	wire w_dff_A_pu988qNr8_0;
	wire w_dff_A_TiDgNwFx9_0;
	wire w_dff_A_qfXhWJqT3_0;
	wire w_dff_A_ucyWdUIR6_0;
	wire w_dff_A_e59Izlyj0_0;
	wire w_dff_A_NCxwK95s0_0;
	wire w_dff_A_EHU2iTZ85_0;
	wire w_dff_A_I3LmKJ0a0_0;
	wire w_dff_A_RGgYilYt3_0;
	wire w_dff_A_jYc7f8nn5_0;
	wire w_dff_A_Jo20Jtiw2_0;
	wire w_dff_A_uoq4Zv620_0;
	wire w_dff_A_dhqS9DYw0_0;
	wire w_dff_A_1EcuuRWd2_0;
	wire w_dff_A_tqaP1fcJ2_0;
	wire w_dff_A_T6cWsFWg9_0;
	wire w_dff_A_PFp8LOMS9_0;
	wire w_dff_A_eIIO9z1t3_0;
	wire w_dff_A_d5oFxJLf5_1;
	wire w_dff_A_quqgr5Ep4_0;
	wire w_dff_A_nDQWTRPm9_0;
	wire w_dff_A_IXPg4fPj5_0;
	wire w_dff_A_OT9aXnPz7_0;
	wire w_dff_A_bgBFMxfz9_0;
	wire w_dff_A_1CRCRvHU6_0;
	wire w_dff_A_4dYcBy0D5_0;
	wire w_dff_A_YZE2bGGd5_0;
	wire w_dff_A_Gf0si6rP2_0;
	wire w_dff_A_pu2G6fmg5_0;
	wire w_dff_A_y2EVG8CJ1_0;
	wire w_dff_A_1H3gRmuE6_0;
	wire w_dff_A_uLkpO3pV7_0;
	wire w_dff_A_rAJ53Wdx1_0;
	wire w_dff_A_0HpOOd7h2_0;
	wire w_dff_A_T8Kb0OIX8_0;
	wire w_dff_A_scDPLGRk8_0;
	wire w_dff_A_7RWBD3Em3_0;
	wire w_dff_A_AsPJgWuK7_0;
	wire w_dff_A_quc44TPB0_0;
	wire w_dff_A_YG3pGkx39_0;
	wire w_dff_A_Q0csuqQ08_0;
	wire w_dff_A_MEDAvAne0_0;
	wire w_dff_A_YbC1Kx7X5_0;
	wire w_dff_A_psklSFAO5_1;
	wire w_dff_A_syrspiJb8_0;
	wire w_dff_A_XSH3hame1_0;
	wire w_dff_A_K8z4jh8m4_0;
	wire w_dff_A_LLaQKBrF0_0;
	wire w_dff_A_eu9UKrS33_0;
	wire w_dff_A_N57dancA2_0;
	wire w_dff_A_Xb1Xrrqc1_0;
	wire w_dff_A_8byz53nP5_0;
	wire w_dff_A_ylQtX0ZS3_0;
	wire w_dff_A_YZHKLBLI0_0;
	wire w_dff_A_A0PZnddb2_0;
	wire w_dff_A_3MCGZOZF1_0;
	wire w_dff_A_9UjTvXEI2_0;
	wire w_dff_A_yx2royOW5_0;
	wire w_dff_A_5ommu2eA0_0;
	wire w_dff_A_IdFX6uti6_0;
	wire w_dff_A_KoxbzP5h4_0;
	wire w_dff_A_eOMRKb965_0;
	wire w_dff_A_UcSv1Yyw5_0;
	wire w_dff_A_HMmeEGFG3_0;
	wire w_dff_A_MX8T0eGB3_0;
	wire w_dff_A_cq4jRdSq2_0;
	wire w_dff_A_pvGf9Poj9_0;
	wire w_dff_A_1L88bpv31_0;
	wire w_dff_A_TwNsD2rL2_1;
	wire w_dff_A_zLtiV7Hl9_0;
	wire w_dff_A_duLohmMZ1_0;
	wire w_dff_A_hjWfbfeb6_0;
	wire w_dff_A_OSSPYYo76_0;
	wire w_dff_A_E6ZTtMGZ3_0;
	wire w_dff_A_0IPypipt7_0;
	wire w_dff_A_Z2xrnaVM5_0;
	wire w_dff_A_Hg0nen860_0;
	wire w_dff_A_XDf9c3wR6_0;
	wire w_dff_A_buoU9x751_0;
	wire w_dff_A_h7ZSJErN6_0;
	wire w_dff_A_g9BseHpq7_0;
	wire w_dff_A_7xrpUrne1_0;
	wire w_dff_A_DZ7eClga0_0;
	wire w_dff_A_gWzVaXk65_0;
	wire w_dff_A_KZcGxfVS7_0;
	wire w_dff_A_dv9B6CSK3_0;
	wire w_dff_A_LajfI1038_0;
	wire w_dff_A_QeLeoSHx3_0;
	wire w_dff_A_bPIA2cJk9_0;
	wire w_dff_A_CgEWVihV8_0;
	wire w_dff_A_KflzC4fR3_0;
	wire w_dff_A_n19JPVCU6_0;
	wire w_dff_A_Egpwz42Y4_0;
	wire w_dff_A_g9Y6z9mT9_1;
	wire w_dff_A_xoVR1WGa0_0;
	wire w_dff_A_GbRR1pC52_0;
	wire w_dff_A_SRYHYUhx9_0;
	wire w_dff_A_2Bze2Tpt1_0;
	wire w_dff_A_8qPQBUGx5_0;
	wire w_dff_A_Anzu2NlP5_0;
	wire w_dff_A_Og5HVl4t3_0;
	wire w_dff_A_RKVFx3rx9_0;
	wire w_dff_A_oKhytRBm2_0;
	wire w_dff_A_cj2SuduW6_0;
	wire w_dff_A_VAivyzf87_0;
	wire w_dff_A_uP6xiXyD9_0;
	wire w_dff_A_nEF9ZX820_0;
	wire w_dff_A_Y9Y79gPP0_0;
	wire w_dff_A_bA9IK4OQ6_0;
	wire w_dff_A_qR2bPC1j4_0;
	wire w_dff_A_j646Whri1_0;
	wire w_dff_A_9ekTT3Ee1_0;
	wire w_dff_A_CTxqaQiW0_0;
	wire w_dff_A_9eDpmNFz8_0;
	wire w_dff_A_ArXhC84a1_0;
	wire w_dff_A_FUPUOTjR9_0;
	wire w_dff_A_K8MWOyGH7_0;
	wire w_dff_A_zQTFQxmk5_0;
	wire w_dff_A_wMjzKV3T2_1;
	wire w_dff_A_gmVc3HeH7_0;
	wire w_dff_A_YPmVzXo50_0;
	wire w_dff_A_xqcHp5R21_0;
	wire w_dff_A_rVueodNB8_0;
	wire w_dff_A_eHzjibSc4_0;
	wire w_dff_A_5uZGPdgs1_0;
	wire w_dff_A_HRzcRnuI6_0;
	wire w_dff_A_rLCtRtjC3_0;
	wire w_dff_A_XwsGc7vW0_0;
	wire w_dff_A_K6oDWatf0_0;
	wire w_dff_A_Rshwbgwf2_0;
	wire w_dff_A_QR3LTFu02_0;
	wire w_dff_A_WBggRGbi8_0;
	wire w_dff_A_OeeRPS5c6_0;
	wire w_dff_A_ZONYte9y6_0;
	wire w_dff_A_V31Tc6V30_0;
	wire w_dff_A_H93WLYsM3_0;
	wire w_dff_A_xwm1JBI16_0;
	wire w_dff_A_Zx9bzyRT9_0;
	wire w_dff_A_zo4VTCwN4_0;
	wire w_dff_A_TwlQBUXs8_0;
	wire w_dff_A_5ZZaC6uo4_0;
	wire w_dff_A_ZcXqDxnv5_0;
	wire w_dff_A_uxhrSHau9_0;
	wire w_dff_A_ngmk1eik7_2;
	wire w_dff_A_rCDjaHpI3_0;
	wire w_dff_A_8Fp46olI2_0;
	wire w_dff_A_D00HEcCH4_0;
	wire w_dff_A_gH1Kf8c15_0;
	wire w_dff_A_8KpQHMKD2_0;
	wire w_dff_A_VLlphInN5_0;
	wire w_dff_A_sEYst0N12_0;
	wire w_dff_A_oDNmbRjH9_0;
	wire w_dff_A_ZnmBmKwa8_0;
	wire w_dff_A_dpsqOQpb0_0;
	wire w_dff_A_OjUtfoEE1_0;
	wire w_dff_A_9BfVnHtw1_0;
	wire w_dff_A_QQFFRuzS3_0;
	wire w_dff_A_px73EUeB5_0;
	wire w_dff_A_M5txvtd66_0;
	wire w_dff_A_haqALR7a5_0;
	wire w_dff_A_GMIVcFp51_0;
	wire w_dff_A_VthD3EiR5_0;
	wire w_dff_A_Qo5xvpQj6_0;
	wire w_dff_A_b2JQRBmH9_0;
	wire w_dff_A_ifWuJqJ83_0;
	wire w_dff_A_Zz5O4hms8_0;
	wire w_dff_A_3QCPLwDI3_0;
	wire w_dff_A_nNDblEMt0_0;
	wire w_dff_A_WaFIGnAa9_1;
	wire w_dff_A_93k3q9BE5_0;
	wire w_dff_A_9hnNWfb10_0;
	wire w_dff_A_2sykZE7m1_0;
	wire w_dff_A_rNgubPbI6_0;
	wire w_dff_A_iVnlT7Q32_0;
	wire w_dff_A_c9kx7tNO6_0;
	wire w_dff_A_SOLqzsQl7_0;
	wire w_dff_A_d7pt807o9_0;
	wire w_dff_A_ooIhtFkB7_0;
	wire w_dff_A_nZQSRnHI9_0;
	wire w_dff_A_QxlC37c31_0;
	wire w_dff_A_nJjLr0CU5_0;
	wire w_dff_A_tjkX94Uo2_0;
	wire w_dff_A_4ncXZcSP6_0;
	wire w_dff_A_ul7MAnSa8_0;
	wire w_dff_A_A9lO3CyH0_0;
	wire w_dff_A_tei56dez2_0;
	wire w_dff_A_dbgaP0Rd6_0;
	wire w_dff_A_zIE918rM8_0;
	wire w_dff_A_jHC6zbkX0_0;
	wire w_dff_A_yXCkIIaN8_0;
	wire w_dff_A_Kd84SJZL2_0;
	wire w_dff_A_XpduZ7gz3_0;
	wire w_dff_A_ZcQWVm3f9_0;
	wire w_dff_A_A8hVAlbl2_1;
	wire w_dff_A_KH2E4U4e4_0;
	wire w_dff_A_tkfU81ia3_0;
	wire w_dff_A_nCnTvZXH7_0;
	wire w_dff_A_92PqVcHB6_0;
	wire w_dff_A_tNAYM1pR1_0;
	wire w_dff_A_wVXn3hKW8_0;
	wire w_dff_A_rIPsPQuG7_0;
	wire w_dff_A_zgWqaAK52_0;
	wire w_dff_A_dtvCJSli3_0;
	wire w_dff_A_yJayNhdq3_0;
	wire w_dff_A_2GEzOe1q2_0;
	wire w_dff_A_L5oDVMKh8_0;
	wire w_dff_A_BowNEFNZ4_0;
	wire w_dff_A_VKRxySFe8_0;
	wire w_dff_A_WLAFVOWO8_0;
	wire w_dff_A_Bgsxl5rv3_0;
	wire w_dff_A_QgrlKjMZ9_0;
	wire w_dff_A_9CvrZqXc7_0;
	wire w_dff_A_cNkqUffv4_0;
	wire w_dff_A_ajt3F2WD9_0;
	wire w_dff_A_dqDyWFJM1_0;
	wire w_dff_A_UXRWSh954_0;
	wire w_dff_A_5VHLvVjS9_0;
	wire w_dff_A_yt3bbOY15_0;
	wire w_dff_A_6894XwHg4_1;
	wire w_dff_A_VUbwMfnm3_0;
	wire w_dff_A_zr9POrwW8_0;
	wire w_dff_A_sMbWaRLX6_0;
	wire w_dff_A_1XPA7sXR5_0;
	wire w_dff_A_kFXeJVb30_0;
	wire w_dff_A_y2PETxVf7_0;
	wire w_dff_A_x4CznEat7_0;
	wire w_dff_A_PRj8j7ey4_0;
	wire w_dff_A_FrficphV1_0;
	wire w_dff_A_s5TIPeLb3_0;
	wire w_dff_A_2kcw91Yq1_0;
	wire w_dff_A_8sfHadIK8_0;
	wire w_dff_A_OSf0b74V5_0;
	wire w_dff_A_dRVYuHOA4_0;
	wire w_dff_A_2M1msprE8_0;
	wire w_dff_A_gOzqewLt1_0;
	wire w_dff_A_a5EILIGX6_0;
	wire w_dff_A_582nY0w96_0;
	wire w_dff_A_QMTVzXzd3_0;
	wire w_dff_A_cIUchttw2_0;
	wire w_dff_A_C5aoSTNr3_0;
	wire w_dff_A_kIt2ysnS1_0;
	wire w_dff_A_5JgXSuOx1_0;
	wire w_dff_A_nKfqeR3a3_0;
	wire w_dff_A_HHWOph5b7_1;
	wire w_dff_A_ZAzv3gLz8_0;
	wire w_dff_A_Kels9HHA8_0;
	wire w_dff_A_LkcUbwPK6_0;
	wire w_dff_A_B9sJDTNd5_0;
	wire w_dff_A_1DfwWTjw2_0;
	wire w_dff_A_C13xRN3G3_0;
	wire w_dff_A_9h366wQY5_0;
	wire w_dff_A_aHEwNMML6_0;
	wire w_dff_A_rtXwMPxD3_0;
	wire w_dff_A_0qSHGKcc8_0;
	wire w_dff_A_eDZD0ueg6_0;
	wire w_dff_A_48n1I4sP6_0;
	wire w_dff_A_5VSxk5bT8_0;
	wire w_dff_A_tlqG2zrB3_0;
	wire w_dff_A_hntE2EzT4_0;
	wire w_dff_A_frLa6Gon1_0;
	wire w_dff_A_teqW8fCd1_0;
	wire w_dff_A_DrdRFazP4_0;
	wire w_dff_A_Wn06qBZI2_0;
	wire w_dff_A_QnuJmDG62_0;
	wire w_dff_A_6aFDZH2V1_0;
	wire w_dff_A_MivsMC8G0_0;
	wire w_dff_A_G6V5Phx14_0;
	wire w_dff_A_BBo1gajo5_0;
	wire w_dff_A_YkzxoQtB2_2;
	wire w_dff_A_mmoyTtaK6_0;
	wire w_dff_A_UYGS9ZSh3_0;
	wire w_dff_A_QmOblBJQ6_0;
	wire w_dff_A_eP4zlPHi9_0;
	wire w_dff_A_odDFbvq47_0;
	wire w_dff_A_GykK2TQp8_0;
	wire w_dff_A_kegSiuQZ0_0;
	wire w_dff_A_LsPpmI8K4_0;
	wire w_dff_A_P7vfS4vW8_0;
	wire w_dff_A_wYl99yhY5_0;
	wire w_dff_A_mdSwKMO74_0;
	wire w_dff_A_uZ27h9L10_0;
	wire w_dff_A_7dZeTwjs7_0;
	wire w_dff_A_xdFoL6JW4_0;
	wire w_dff_A_J9zpjoO99_0;
	wire w_dff_A_SpWTup9B5_0;
	wire w_dff_A_Iizw5isy6_0;
	wire w_dff_A_WW3mjIsK2_0;
	wire w_dff_A_Qax9Srjc9_0;
	wire w_dff_A_bVqY3Jc39_0;
	wire w_dff_A_hdUwCm208_0;
	wire w_dff_A_Uo588KnT3_0;
	wire w_dff_A_sMAmJ0391_0;
	wire w_dff_A_SYGTJskO0_0;
	wire w_dff_A_gMoTHiyF2_2;
	wire w_dff_A_VTjsgKuU1_0;
	wire w_dff_A_b2ZEFNbE4_0;
	wire w_dff_A_apAu1UK38_0;
	wire w_dff_A_1xrwjf0X2_0;
	wire w_dff_A_D61E1PyV9_0;
	wire w_dff_A_7QbUsl7H7_0;
	wire w_dff_A_mdLjyh2k4_0;
	wire w_dff_A_VROJQ4Gx0_0;
	wire w_dff_A_1sAMcDo47_0;
	wire w_dff_A_CijIXDxo4_0;
	wire w_dff_A_St6DHmPu7_0;
	wire w_dff_A_snPcbtFQ5_0;
	wire w_dff_A_qyj4bKDl1_0;
	wire w_dff_A_FZlwYflm1_0;
	wire w_dff_A_IcH8j55H2_0;
	wire w_dff_A_dGM0tJA56_0;
	wire w_dff_A_6CXnUImU7_0;
	wire w_dff_A_SHy3muHk4_0;
	wire w_dff_A_hwHC8ITx6_0;
	wire w_dff_A_zmw4w8hz5_0;
	wire w_dff_A_sYxNjcml1_0;
	wire w_dff_A_l5LsU9RF8_0;
	wire w_dff_A_t8HbDwEf1_0;
	wire w_dff_A_YXrgNVZe8_2;
	wire w_dff_A_XBiahQiV1_0;
	wire w_dff_A_VHUl1q965_0;
	wire w_dff_A_5kJR66x03_0;
	wire w_dff_A_k8G3Iiji4_0;
	wire w_dff_A_SBLV8qSQ0_0;
	wire w_dff_A_eu8hscUt3_0;
	wire w_dff_A_pD89C3Zv5_0;
	wire w_dff_A_VlRmVwy42_0;
	wire w_dff_A_YONZH3dx4_0;
	wire w_dff_A_DPkgoYry5_0;
	wire w_dff_A_dzQlXcd66_0;
	wire w_dff_A_Y0zh1ZFY3_0;
	wire w_dff_A_MqYoul0z3_0;
	wire w_dff_A_ClAPdzkd6_0;
	wire w_dff_A_dtA90Sy32_0;
	wire w_dff_A_VjPpPFTp6_0;
	wire w_dff_A_ApezIZL96_0;
	wire w_dff_A_QSzkMrGA6_0;
	wire w_dff_A_tx9EFmX79_0;
	wire w_dff_A_4onzlFIs1_0;
	wire w_dff_A_A8BHtBpx3_0;
	wire w_dff_A_pSIcjSir7_0;
	wire w_dff_A_ufMWgX2S9_0;
	wire w_dff_A_1vhZ3Duu7_1;
	wire w_dff_A_xaBEhCvg3_0;
	wire w_dff_A_pMzJ0rrY7_0;
	wire w_dff_A_fO54PrRc4_0;
	wire w_dff_A_eWGuX4Hb2_0;
	wire w_dff_A_NR5x9ZaJ0_0;
	wire w_dff_A_MWxkboMK8_0;
	wire w_dff_A_UKXlgs5R2_0;
	wire w_dff_A_uK8usMXv9_0;
	wire w_dff_A_7dLbHxSa0_0;
	wire w_dff_A_4aFYLfiw4_0;
	wire w_dff_A_OKojFEkQ4_0;
	wire w_dff_A_fbpJGHyl3_0;
	wire w_dff_A_FhDDhKGI1_0;
	wire w_dff_A_LHAumLIi6_0;
	wire w_dff_A_HsLX4xME8_0;
	wire w_dff_A_CfemMX3W6_0;
	wire w_dff_A_i1NQu6Jo8_0;
	wire w_dff_A_x9aHuxnc3_0;
	wire w_dff_A_RZLM3YlS2_0;
	wire w_dff_A_rRg7ndCF2_0;
	wire w_dff_A_2h9pkyBl4_0;
	wire w_dff_A_HCWGWcV32_0;
	wire w_dff_A_blhjv9jP2_0;
	wire w_dff_A_2BQXXCY79_1;
	wire w_dff_A_xRGig8377_0;
	wire w_dff_A_RIhUx2nw8_0;
	wire w_dff_A_aJAoDH2g5_0;
	wire w_dff_A_xyljvqlp7_0;
	wire w_dff_A_kYNBknzr6_0;
	wire w_dff_A_e4dVA2Wt2_0;
	wire w_dff_A_LAGxNsX03_0;
	wire w_dff_A_kgcAoagA8_0;
	wire w_dff_A_PBlo9OsH1_0;
	wire w_dff_A_JM4zImIa8_0;
	wire w_dff_A_iP1J6CzE5_0;
	wire w_dff_A_MhWhCN8g5_0;
	wire w_dff_A_TEZCAOzt6_0;
	wire w_dff_A_ujoQjHiV7_0;
	wire w_dff_A_rN5FmHAw0_0;
	wire w_dff_A_aF6gTfrh1_0;
	wire w_dff_A_7gd1M7G10_0;
	wire w_dff_A_jWpSByPW4_0;
	wire w_dff_A_0Xqw2c5Z1_0;
	wire w_dff_A_zoN5m0oc5_0;
	wire w_dff_A_2Gpg6zHf6_0;
	wire w_dff_A_xEoyoL3u4_0;
	wire w_dff_A_4EYDmp5c0_0;
	wire w_dff_A_6BNVEGbH7_0;
	wire w_dff_A_XHnryFNT6_0;
	wire w_dff_A_RJ7IrVGd3_1;
	wire w_dff_A_EQ37yykE3_0;
	wire w_dff_A_VLt9xiM65_0;
	wire w_dff_A_DSCdIuQx6_0;
	wire w_dff_A_iApKW7MT5_0;
	wire w_dff_A_CUKLLEQw9_0;
	wire w_dff_A_o0AZu8551_0;
	wire w_dff_A_qR4tpdR63_0;
	wire w_dff_A_Y78l4tbm7_0;
	wire w_dff_A_t0iMmbE84_0;
	wire w_dff_A_aprY7Hxz7_0;
	wire w_dff_A_T6rcURAQ7_0;
	wire w_dff_A_cSNB2yKf2_0;
	wire w_dff_A_IgglOpA07_0;
	wire w_dff_A_9kxFLE7j3_0;
	wire w_dff_A_l8NvcR8K1_0;
	wire w_dff_A_CSYG8x4H4_0;
	wire w_dff_A_pHJ7DrXq5_0;
	wire w_dff_A_rpGTnU5z4_0;
	wire w_dff_A_2Hrmf9zX9_0;
	wire w_dff_A_0yDnFnFU8_0;
	wire w_dff_A_ORSg5U0o0_0;
	wire w_dff_A_hxUxrhRC9_0;
	wire w_dff_A_Fl09Z4x47_0;
	wire w_dff_A_ReZpeQio9_0;
	wire w_dff_A_hwsWkcta6_0;
	wire w_dff_A_88VaWVqO6_1;
	wire w_dff_A_KafEuoPR1_0;
	wire w_dff_A_y8BZduW51_0;
	wire w_dff_A_0otdT7wu5_0;
	wire w_dff_A_wi4BtpDo2_0;
	wire w_dff_A_EOmIOPxI8_0;
	wire w_dff_A_rJwRTXNY3_0;
	wire w_dff_A_2pBZzS9a0_0;
	wire w_dff_A_OZjfciZ72_0;
	wire w_dff_A_SlnPlGr07_0;
	wire w_dff_A_k3fXH3ul1_0;
	wire w_dff_A_RiZrk0bw3_0;
	wire w_dff_A_DNyaSlRn9_0;
	wire w_dff_A_4Gw6z5kt8_0;
	wire w_dff_A_X9B1OuZc4_0;
	wire w_dff_A_2VIMb5Cm1_0;
	wire w_dff_A_cYzohbvw3_0;
	wire w_dff_A_FsVl5IM42_0;
	wire w_dff_A_INu8qnWm9_0;
	wire w_dff_A_8mtilUTZ5_0;
	wire w_dff_A_PqAGtkmO5_0;
	wire w_dff_A_anoYIH2a4_0;
	wire w_dff_A_mrfNQf350_0;
	wire w_dff_A_JQf7NqGh5_0;
	wire w_dff_A_FjF4b82V7_0;
	wire w_dff_A_jwap2BjM8_0;
	wire w_dff_A_QSbbVJ567_1;
	wire w_dff_A_QaZHnHBu1_0;
	wire w_dff_A_b0Q9CeWZ6_0;
	wire w_dff_A_q8qnf7pK3_0;
	wire w_dff_A_JlJcvdNA9_0;
	wire w_dff_A_TWurAjsC4_0;
	wire w_dff_A_Cc5q8fmD4_0;
	wire w_dff_A_a3SwUa8v9_0;
	wire w_dff_A_T8pQasFM0_0;
	wire w_dff_A_cenyqIl21_0;
	wire w_dff_A_MmF2BjKi5_0;
	wire w_dff_A_aCTppGsN4_0;
	wire w_dff_A_fEsJgHJk9_0;
	wire w_dff_A_TW6FMMtF0_0;
	wire w_dff_A_L5WsDwWb4_0;
	wire w_dff_A_kIj1TW136_0;
	wire w_dff_A_Es77KwOD5_0;
	wire w_dff_A_ZvSmXE3U3_0;
	wire w_dff_A_YhyW6Jog0_0;
	wire w_dff_A_j5E0o9H89_0;
	wire w_dff_A_cXT5Wqs20_0;
	wire w_dff_A_0VjhFhUN5_0;
	wire w_dff_A_qjYREwnY3_0;
	wire w_dff_A_DesNHXqO3_0;
	wire w_dff_A_oROOZXXm2_0;
	wire w_dff_A_vqllTW0F0_0;
	wire w_dff_A_QFHYc7Fj1_1;
	wire w_dff_A_PMZF4mUi7_0;
	wire w_dff_A_uMG66Qip9_0;
	wire w_dff_A_tBtDY7Dj9_0;
	wire w_dff_A_8tU4DtWU5_0;
	wire w_dff_A_czryexAs0_0;
	wire w_dff_A_NU64LTm80_0;
	wire w_dff_A_OZfb0iRl5_0;
	wire w_dff_A_jquXzVdc4_0;
	wire w_dff_A_IT3xMGJ89_0;
	wire w_dff_A_FyGmX1Lx0_0;
	wire w_dff_A_t4BVRV3q9_0;
	wire w_dff_A_KEWsQdWT0_0;
	wire w_dff_A_fBF1V4431_0;
	wire w_dff_A_02EqBpfb9_0;
	wire w_dff_A_yovzNn3U8_0;
	wire w_dff_A_9u5Ufmuo3_0;
	wire w_dff_A_pYnQYhqq5_0;
	wire w_dff_A_4fMweFG82_0;
	wire w_dff_A_ndtvTD3M6_0;
	wire w_dff_A_XH45lJcj2_0;
	wire w_dff_A_Rrs8FY0R6_0;
	wire w_dff_A_ShDWRVng2_0;
	wire w_dff_A_9UtbIp9q9_0;
	wire w_dff_A_MikKOYaC1_0;
	wire w_dff_A_aTsBRGqL6_0;
	wire w_dff_A_0OPq6GU27_1;
	wire w_dff_A_ISi2XYXx9_0;
	wire w_dff_A_XuQgYQ138_0;
	wire w_dff_A_UBTHxJvq6_0;
	wire w_dff_A_bhTwe7ii2_0;
	wire w_dff_A_0Drf1Qww0_0;
	wire w_dff_A_EbAhbqOP8_0;
	wire w_dff_A_sGW2EcJY2_0;
	wire w_dff_A_nH53o9AR5_0;
	wire w_dff_A_uOnF7NKK8_0;
	wire w_dff_A_PiVhECcY8_0;
	wire w_dff_A_fV546wwq1_0;
	wire w_dff_A_zUyqGHW02_0;
	wire w_dff_A_v0fWeeZW3_0;
	wire w_dff_A_7ujRWc1N2_0;
	wire w_dff_A_3GxMm94q8_0;
	wire w_dff_A_EDVHbBsq2_0;
	wire w_dff_A_BVvSRfeC8_0;
	wire w_dff_A_abvTzoZR6_0;
	wire w_dff_A_zymTnHTE3_0;
	wire w_dff_A_7p8fuMN78_0;
	wire w_dff_A_VDEYP1cj6_0;
	wire w_dff_A_gs9mOI0f8_0;
	wire w_dff_A_WmsrZvsf4_0;
	wire w_dff_A_QpbmHz4K1_0;
	wire w_dff_A_9LMyKtbq7_2;
	wire w_dff_A_LeX4LYJX0_0;
	wire w_dff_A_31sOqvSO5_0;
	wire w_dff_A_feVftU9h6_0;
	wire w_dff_A_xUGPZ3vK8_0;
	wire w_dff_A_Mu1m9N2G5_0;
	wire w_dff_A_QvVAdbMb9_0;
	wire w_dff_A_mz4tHFXy9_0;
	wire w_dff_A_ankZ8yng9_0;
	wire w_dff_A_tQw9pSRx5_0;
	wire w_dff_A_5D6J6niT6_0;
	wire w_dff_A_4hyGW6N78_0;
	wire w_dff_A_HSU2GkO85_0;
	wire w_dff_A_rmPzrKzX1_0;
	wire w_dff_A_8LjF2bIZ4_0;
	wire w_dff_A_Qq1VabVP3_0;
	wire w_dff_A_J8ETL6sl0_0;
	wire w_dff_A_pKy6pIv48_0;
	wire w_dff_A_gYQTGHsH9_0;
	wire w_dff_A_omIm2yxE2_0;
	wire w_dff_A_IAowf1US3_0;
	wire w_dff_A_JmMCQgqB9_0;
	wire w_dff_A_OotEsjpD2_0;
	wire w_dff_A_4FDeHSQK4_2;
	wire w_dff_A_53F08RXh9_0;
	wire w_dff_A_bwvFUUO72_0;
	wire w_dff_A_A5EdTfQo3_0;
	wire w_dff_A_ZFRSGBK33_0;
	wire w_dff_A_zWCgwJ4T9_0;
	wire w_dff_A_YfNqVm6O9_0;
	wire w_dff_A_5gVsKW0k9_0;
	wire w_dff_A_QrXXHDQH4_0;
	wire w_dff_A_xl3S76Rj6_0;
	wire w_dff_A_2RrXjq8U9_0;
	wire w_dff_A_gvcGSg713_0;
	wire w_dff_A_dOowzlRw3_0;
	wire w_dff_A_aWPlizYh8_0;
	wire w_dff_A_s0gU8yuk9_0;
	wire w_dff_A_aAet1x6W0_0;
	wire w_dff_A_YnBY93x42_0;
	wire w_dff_A_WmY2AXVv1_0;
	wire w_dff_A_4e7QblSY1_0;
	wire w_dff_A_GgJPlDrh0_0;
	wire w_dff_A_Q7wGKW2c0_0;
	wire w_dff_A_aXxieiC35_0;
	wire w_dff_A_4tE1sT3T7_0;
	wire w_dff_A_v0aZb5kz5_0;
	wire w_dff_A_uN1e9ym35_1;
	wire w_dff_A_DDE8BJzV5_0;
	wire w_dff_A_TSonxKRY3_0;
	wire w_dff_A_rCza6zCY6_0;
	wire w_dff_A_khmZ2pxx1_0;
	wire w_dff_A_XngQgKQy3_0;
	wire w_dff_A_7fnFMIBm4_0;
	wire w_dff_A_AIDI0fd23_0;
	wire w_dff_A_KgGs29KD8_0;
	wire w_dff_A_wEa3E1EL0_0;
	wire w_dff_A_LKZzLQPY9_0;
	wire w_dff_A_e0xTxuDQ8_0;
	wire w_dff_A_DqdAE0c33_0;
	wire w_dff_A_gbRStlEe3_0;
	wire w_dff_A_Zpg4qWUR8_0;
	wire w_dff_A_PDyuMfC12_0;
	wire w_dff_A_Zqu5CR5b2_0;
	wire w_dff_A_drXXU6Wl0_0;
	wire w_dff_A_r8wfL2rL3_0;
	wire w_dff_A_x6ak8e884_0;
	wire w_dff_A_Gp1Zj1qL1_0;
	wire w_dff_A_dBzxZnWH7_0;
	wire w_dff_A_OES7JWNi8_0;
	wire w_dff_A_6Vlmlz5H5_0;
	wire w_dff_A_9RerqaJa3_0;
	wire w_dff_A_EikSB4526_0;
	wire w_dff_A_NnNpN7LE0_1;
	wire w_dff_A_98i8w2QX4_0;
	wire w_dff_A_9dYQ0MBV4_0;
	wire w_dff_A_DhBOJ4mI0_0;
	wire w_dff_A_NOiHHKfc2_0;
	wire w_dff_A_VTOlczNQ1_0;
	wire w_dff_A_KhdQQ4Ov4_0;
	wire w_dff_A_ZiODlsO86_0;
	wire w_dff_A_jDwPP2oX9_0;
	wire w_dff_A_wGH08fmO7_0;
	wire w_dff_A_Ym82e2Zy0_0;
	wire w_dff_A_yseIjvsq8_0;
	wire w_dff_A_IlsbZwWv8_0;
	wire w_dff_A_BoRetuJU2_0;
	wire w_dff_A_DaNirjya4_0;
	wire w_dff_A_NxuwoN3R6_0;
	wire w_dff_A_Cm3wGoB99_0;
	wire w_dff_A_Qc4MAacK3_0;
	wire w_dff_A_sJAmPAgd3_0;
	wire w_dff_A_RXmgIt4l6_0;
	wire w_dff_A_T7iJOIGc1_0;
	wire w_dff_A_VHaoAV704_0;
	wire w_dff_A_SEL3KXPi7_0;
	wire w_dff_A_rMQA6tWD0_0;
	wire w_dff_A_75qgGpF97_0;
	wire w_dff_A_6pcevl1s5_0;
	wire w_dff_A_2LtSmUnw2_1;
	wire w_dff_A_DCEKpMZe3_0;
	wire w_dff_A_0RrCnvrw0_0;
	wire w_dff_A_ucFluxaL0_0;
	wire w_dff_A_JFZVaWzo0_0;
	wire w_dff_A_xGJ73V7C3_0;
	wire w_dff_A_hXk3t87U7_0;
	wire w_dff_A_lvOqVOJH5_0;
	wire w_dff_A_Dj34yWJ18_0;
	wire w_dff_A_KRYBHC5Y6_0;
	wire w_dff_A_4u9beA0C5_0;
	wire w_dff_A_w4d3SPld0_0;
	wire w_dff_A_ARXar45I3_0;
	wire w_dff_A_SkSXS6uy7_0;
	wire w_dff_A_jiEc8ZSq2_0;
	wire w_dff_A_XQ7Z9yFc3_0;
	wire w_dff_A_9dvFI3ha0_0;
	wire w_dff_A_4Wv4Koqv0_0;
	wire w_dff_A_XGyd3ihA6_0;
	wire w_dff_A_UhiWgx794_0;
	wire w_dff_A_94BZuozg1_0;
	wire w_dff_A_prXiWfPG5_0;
	wire w_dff_A_oW37fLM99_0;
	wire w_dff_A_PRPlMr0e0_0;
	wire w_dff_A_7XjXvFRw8_0;
	wire w_dff_A_0kCIwMLz2_0;
	wire w_dff_A_bhCkHx8o1_1;
	wire w_dff_A_zLAD9MAs6_0;
	wire w_dff_A_b6PyrG9D0_0;
	wire w_dff_A_lvAjtu2Q0_0;
	wire w_dff_A_T2xVdAGo9_0;
	wire w_dff_A_jixHMTo23_0;
	wire w_dff_A_mECcdmDu5_0;
	wire w_dff_A_FNhYLUNV5_0;
	wire w_dff_A_8OQW41Jt0_0;
	wire w_dff_A_7yVhsTkT7_0;
	wire w_dff_A_AY4Qnx3m1_0;
	wire w_dff_A_2KyOlAVx1_0;
	wire w_dff_A_cGMDKwWw0_0;
	wire w_dff_A_b697pHxQ3_0;
	wire w_dff_A_XwvzxxTH2_0;
	wire w_dff_A_QEI5p7Ym3_0;
	wire w_dff_A_i89gtJ4S1_0;
	wire w_dff_A_hkTJ0VYW7_0;
	wire w_dff_A_frv7p8y58_0;
	wire w_dff_A_pX3Q8Uax0_0;
	wire w_dff_A_X8Oysb7a4_0;
	wire w_dff_A_SJshBxdt8_0;
	wire w_dff_A_wgAF5rYA2_0;
	wire w_dff_A_nCKnPfb64_0;
	wire w_dff_A_CGUXvuJH3_0;
	wire w_dff_A_SZHdqKEr8_0;
	wire w_dff_A_RvDEgF9N8_1;
	wire w_dff_A_IznpfcOq9_0;
	wire w_dff_A_uC2juEjC4_0;
	wire w_dff_A_BEDOENFC3_0;
	wire w_dff_A_QjCXCqBQ4_0;
	wire w_dff_A_o8QopJDN1_0;
	wire w_dff_A_vKCqEmq32_0;
	wire w_dff_A_zqgyP5oj2_0;
	wire w_dff_A_Mm1v7Vpq4_0;
	wire w_dff_A_SEvXjhlY9_0;
	wire w_dff_A_aV8lqEBR2_0;
	wire w_dff_A_gtfNUY6z8_0;
	wire w_dff_A_WgVb8MiY2_0;
	wire w_dff_A_utU4WP8j4_0;
	wire w_dff_A_wYt4UxtS9_0;
	wire w_dff_A_LChqDAVs6_0;
	wire w_dff_A_WFQUi4jm7_0;
	wire w_dff_A_fh5MCp210_0;
	wire w_dff_A_3BRew9G51_0;
	wire w_dff_A_7voMf0we2_0;
	wire w_dff_A_aMG0QwnA1_0;
	wire w_dff_A_rhrrGLpy9_0;
	wire w_dff_A_6ajUOm4r9_0;
	wire w_dff_A_OCYlJY7m3_0;
	wire w_dff_A_uHcHn3hs4_0;
	wire w_dff_A_qZ1mA9zs2_0;
	wire w_dff_A_T8dVu50g8_1;
	wire w_dff_A_zCnTskqc8_0;
	wire w_dff_A_gHTbkyaV1_0;
	wire w_dff_A_olhd6I4n0_0;
	wire w_dff_A_wPRKyTpU9_0;
	wire w_dff_A_Hx7mchhX6_0;
	wire w_dff_A_FNdUpmAq0_0;
	wire w_dff_A_JpvWkjLX2_0;
	wire w_dff_A_6kbN3b4b6_0;
	wire w_dff_A_9TxPnvMs2_0;
	wire w_dff_A_jyClKqdg3_0;
	wire w_dff_A_C72m2Eqj5_0;
	wire w_dff_A_GUGD6aYS7_0;
	wire w_dff_A_tqigecYc7_0;
	wire w_dff_A_ECmDm9Ct1_0;
	wire w_dff_A_iCCmfY0J1_0;
	wire w_dff_A_eM0jEiUq3_0;
	wire w_dff_A_4wD3UChI2_0;
	wire w_dff_A_6cuahdtq3_0;
	wire w_dff_A_bARsrghJ2_0;
	wire w_dff_A_bYhM0UFD5_0;
	wire w_dff_A_2ntibkXR3_0;
	wire w_dff_A_cgYWLNPD1_0;
	wire w_dff_A_HVpuMc0R9_0;
	wire w_dff_A_ThLUgkNN4_0;
	wire w_dff_A_tjW8NLMX1_2;
	wire w_dff_A_H9TNAipS8_0;
	wire w_dff_A_sil2BaHk4_0;
	wire w_dff_A_VLwvdYqM6_0;
	wire w_dff_A_rX4nh5r81_0;
	wire w_dff_A_vch1eA7O4_0;
	wire w_dff_A_7Uklk3uY4_0;
	wire w_dff_A_hl8XfH9q8_0;
	wire w_dff_A_dY4JM8Ma9_0;
	wire w_dff_A_GZ03g1l60_0;
	wire w_dff_A_gWiapdnz4_0;
	wire w_dff_A_jDBS4Kto3_0;
	wire w_dff_A_P93ZEZVW4_0;
	wire w_dff_A_lg3M9YNX1_0;
	wire w_dff_A_qXoz65Xu8_0;
	wire w_dff_A_XUmZkIFP7_0;
	wire w_dff_A_AQvfuaaX8_0;
	wire w_dff_A_kg737fNl7_0;
	wire w_dff_A_SNaRIK6p4_0;
	wire w_dff_A_Wkobyo4c0_0;
	wire w_dff_A_6aUo4ehg0_0;
	wire w_dff_A_kxfuJvZt2_0;
	wire w_dff_A_uZFyizaT3_2;
	wire w_dff_A_Iup5Etr22_0;
	wire w_dff_A_zEyb8kbB2_0;
	wire w_dff_A_KMKmbzve9_0;
	wire w_dff_A_tCRS59BQ5_0;
	wire w_dff_A_3A0r1Zwr9_0;
	wire w_dff_A_ynd2r14n7_0;
	wire w_dff_A_9QrrjaJT4_0;
	wire w_dff_A_ozVDdAKz4_0;
	wire w_dff_A_3oAHYtvh7_0;
	wire w_dff_A_O0EBbhyD2_0;
	wire w_dff_A_SgG66Y1N3_0;
	wire w_dff_A_FR8mPSDU0_0;
	wire w_dff_A_EZgT09lv2_0;
	wire w_dff_A_mdVCiKD18_0;
	wire w_dff_A_pLRXoKy13_0;
	wire w_dff_A_ilRRf97M4_0;
	wire w_dff_A_A3p5oRWj4_0;
	wire w_dff_A_oHAqSUbo6_0;
	wire w_dff_A_xrM4FbYP1_0;
	wire w_dff_A_10oEFGMw0_0;
	wire w_dff_A_IDmsZhwS0_0;
	wire w_dff_A_aInYLOFA7_2;
	wire w_dff_A_ZzjTEjGE7_0;
	wire w_dff_A_hvGCZTZv2_0;
	wire w_dff_A_dk8TRHFN4_0;
	wire w_dff_A_3Ga9Nzbe8_0;
	wire w_dff_A_DBBTDaqh3_0;
	wire w_dff_A_ACcmO2X72_0;
	wire w_dff_A_ORXd5Uni3_0;
	wire w_dff_A_qkeM14Wh7_0;
	wire w_dff_A_HeTKmtDF6_0;
	wire w_dff_A_aWji6Cq39_0;
	wire w_dff_A_uuD7Po8Z1_0;
	wire w_dff_A_5GOF8sjO1_0;
	wire w_dff_A_4GQM5DdY2_0;
	wire w_dff_A_ry4Va7jZ7_0;
	wire w_dff_A_DIqvilCI7_0;
	wire w_dff_A_a4WbtcNh0_0;
	wire w_dff_A_TvK4fqcj2_0;
	wire w_dff_A_w9GpjKFG1_0;
	wire w_dff_A_g32NSzLX6_0;
	wire w_dff_A_IFl1JOmu2_0;
	wire w_dff_A_Hq8CUuOH4_0;
	wire w_dff_A_1RnTGjF92_2;
	wire w_dff_A_XpeFdbpX0_0;
	wire w_dff_A_qXnvJGO68_0;
	wire w_dff_A_hPdSzwCK3_0;
	wire w_dff_A_Aw2K0WOu6_0;
	wire w_dff_A_Lim1RbxU1_0;
	wire w_dff_A_gVqOoBCH6_0;
	wire w_dff_A_clBYr3K46_0;
	wire w_dff_A_k5oBvWcm8_0;
	wire w_dff_A_nV9mWPoL6_0;
	wire w_dff_A_vgpmPwJH4_0;
	wire w_dff_A_tagrcOs30_0;
	wire w_dff_A_IQ12Qa1e2_0;
	wire w_dff_A_UWdADaUp5_0;
	wire w_dff_A_Hk7d1xco6_0;
	wire w_dff_A_G54k42aC6_0;
	wire w_dff_A_heO1fFTY3_0;
	wire w_dff_A_zDmiktN89_0;
	wire w_dff_A_4u5QF0U34_0;
	wire w_dff_A_HVzwcJTv6_0;
	wire w_dff_A_WK95aYuy6_0;
	wire w_dff_A_dU76sXvb9_0;
	wire w_dff_A_jHzqXZsV3_0;
	wire w_dff_A_MTvHxVse2_2;
	wire w_dff_A_hBJW0UE92_0;
	wire w_dff_A_dy8GyFLw3_0;
	wire w_dff_A_iPZrgL0e7_0;
	wire w_dff_A_vYlvHLsT8_0;
	wire w_dff_A_GaaDZ0Cp9_0;
	wire w_dff_A_T47ab6ca4_0;
	wire w_dff_A_jYjs7tBs0_0;
	wire w_dff_A_8hUwGXOE5_0;
	wire w_dff_A_v7nK7nE98_0;
	wire w_dff_A_wrw7TbOF9_0;
	wire w_dff_A_wztYHFfo8_0;
	wire w_dff_A_UAx68KMz9_0;
	wire w_dff_A_Vl0CtV079_0;
	wire w_dff_A_2cPrXCWR7_0;
	wire w_dff_A_F84Qf7T07_0;
	wire w_dff_A_CyKOGwFh5_0;
	wire w_dff_A_IdE90A2W3_0;
	wire w_dff_A_AbukKjR94_0;
	wire w_dff_A_nRVSS5K52_0;
	wire w_dff_A_uxirQxCC7_0;
	wire w_dff_A_QgILRn1A0_2;
	wire w_dff_A_rJEdO5Bd8_0;
	wire w_dff_A_ONVyIf2B8_0;
	wire w_dff_A_Diyd9NdS1_0;
	wire w_dff_A_YFEfdFOq8_0;
	wire w_dff_A_nsDddu9i0_0;
	wire w_dff_A_WwWJaJPh2_0;
	wire w_dff_A_H7AXLq781_0;
	wire w_dff_A_GGInvWlw1_0;
	wire w_dff_A_mPbDdSW04_0;
	wire w_dff_A_mAjVKfb88_0;
	wire w_dff_A_JxsdCr5v8_0;
	wire w_dff_A_mG9LsSU07_0;
	wire w_dff_A_ceylxuyL0_0;
	wire w_dff_A_Qw3y8sc13_0;
	wire w_dff_A_H7WRDg3Q7_0;
	wire w_dff_A_Rfx2JrZF2_0;
	wire w_dff_A_0CYqhtmb9_0;
	wire w_dff_A_FsE5HE270_0;
	wire w_dff_A_M1KVHirV2_0;
	wire w_dff_A_aZo1DHpL7_0;
	wire w_dff_A_0GmzN7ei2_2;
	wire w_dff_A_duon9KZm0_0;
	wire w_dff_A_zAKwyIc84_0;
	wire w_dff_A_mBPgKd0S5_0;
	wire w_dff_A_SLtzBcl09_0;
	wire w_dff_A_ekZ0o5Kc1_0;
	wire w_dff_A_tjAcEdqW8_0;
	wire w_dff_A_R6i15A043_0;
	wire w_dff_A_UUGW9Jqa0_0;
	wire w_dff_A_VNKoP4VG1_0;
	wire w_dff_A_6kqBOXer0_0;
	wire w_dff_A_kH2wlUKi1_0;
	wire w_dff_A_LbLNEQLS3_0;
	wire w_dff_A_10js08Js5_0;
	wire w_dff_A_eeOB5FER8_0;
	wire w_dff_A_NyySJDko3_0;
	wire w_dff_A_6JavPM1P1_0;
	wire w_dff_A_A89uGD5j2_0;
	wire w_dff_A_TU3vFcyh3_0;
	wire w_dff_A_ck8ovaT59_0;
	wire w_dff_A_VTUk3OHL6_0;
	wire w_dff_A_0tDgTm6S3_2;
	wire w_dff_A_jzhstoLj0_0;
	wire w_dff_A_nUx6zhfL5_0;
	wire w_dff_A_XjufneCv9_0;
	wire w_dff_A_UvBoPF852_0;
	wire w_dff_A_hjuMrogZ7_0;
	wire w_dff_A_R8kemgtX8_0;
	wire w_dff_A_r3H9kFdA5_0;
	wire w_dff_A_6DdDNP5z0_0;
	wire w_dff_A_8vrG5R2g8_0;
	wire w_dff_A_gs3auYyT9_0;
	wire w_dff_A_GakBwCVH6_0;
	wire w_dff_A_qo3XzztQ9_0;
	wire w_dff_A_YLapVxBp0_0;
	wire w_dff_A_lSmte0YH2_0;
	wire w_dff_A_tQ2AxIQU9_0;
	wire w_dff_A_OP2lL9df7_0;
	wire w_dff_A_ZwzSGMdN1_0;
	wire w_dff_A_YZcJYF1H1_0;
	wire w_dff_A_q4ijwy397_0;
	wire w_dff_A_WmIreB3a9_0;
	wire w_dff_A_MDA1CyFJ0_2;
	wire w_dff_A_lOytSnZh2_0;
	wire w_dff_A_Vwr0DdND6_0;
	wire w_dff_A_EcwGGLiT4_0;
	wire w_dff_A_kEeA7pO89_0;
	wire w_dff_A_EjAI1DBK7_0;
	wire w_dff_A_080ubyZE2_0;
	wire w_dff_A_ZJmhIdV58_0;
	wire w_dff_A_rKaC1NUK0_0;
	wire w_dff_A_l4kRRui19_0;
	wire w_dff_A_KrnvwBLl7_0;
	wire w_dff_A_ag3fLpp56_0;
	wire w_dff_A_Ax5Uy56q6_0;
	wire w_dff_A_Hv0zqIUP4_0;
	wire w_dff_A_YOg9rkaN6_0;
	wire w_dff_A_nPJjfh300_0;
	wire w_dff_A_1XsTjUlC5_0;
	wire w_dff_A_JI54GYgt8_2;
	wire w_dff_A_w0BV9Hwn9_0;
	wire w_dff_A_JRxSQKDk0_0;
	wire w_dff_A_eh6D1e7U1_0;
	wire w_dff_A_BTHJQcXM5_0;
	wire w_dff_A_cDVLQgpE8_0;
	wire w_dff_A_sbTycoJG4_0;
	wire w_dff_A_jQYkZMLj8_0;
	wire w_dff_A_6FLfHyDC3_0;
	wire w_dff_A_1M0IZtja1_0;
	wire w_dff_A_XiVTC9CX2_0;
	wire w_dff_A_khFTa7cK8_0;
	wire w_dff_A_gfIZ3ys35_0;
	wire w_dff_A_5o39kAha7_0;
	wire w_dff_A_SM6zpNTd5_0;
	wire w_dff_A_8Uh82O9k9_0;
	wire w_dff_A_vhiEA8VD0_0;
	wire w_dff_A_QgbmpZht9_2;
	wire w_dff_A_GMILkGLM9_0;
	wire w_dff_A_VlpjscMX6_0;
	wire w_dff_A_yKboFWFA5_0;
	wire w_dff_A_KX9Tqpgr0_0;
	wire w_dff_A_NsyMePNK7_0;
	wire w_dff_A_VjAGNj3F7_0;
	wire w_dff_A_moX6JpjN0_0;
	wire w_dff_A_Lr7p19I87_0;
	wire w_dff_A_mL4SnxAD9_0;
	wire w_dff_A_wDWFw27g5_0;
	wire w_dff_A_HmxKfANZ3_0;
	wire w_dff_A_mz0dJCbt9_0;
	wire w_dff_A_GULorWJ72_0;
	wire w_dff_A_iQdzLS0R2_0;
	wire w_dff_A_0OgvtRqK7_2;
	wire w_dff_A_cSb0UA0b2_0;
	wire w_dff_A_XcHrV9VL9_0;
	wire w_dff_A_4jSMUs2g9_0;
	wire w_dff_A_oUSY9uU15_0;
	wire w_dff_A_Vaw4VKmV6_0;
	wire w_dff_A_juh1xyHG3_0;
	wire w_dff_A_Q0wTUQkw1_0;
	wire w_dff_A_kbJX1bYZ4_0;
	wire w_dff_A_H7nS2ORk9_0;
	wire w_dff_A_1zcunMHv4_0;
	wire w_dff_A_6EvOP3fu0_0;
	wire w_dff_A_wqiLaPqg7_0;
	wire w_dff_A_yzKXFTsU4_0;
	wire w_dff_A_OpiAFAgk7_0;
	wire w_dff_A_8yGStRn20_0;
	wire w_dff_A_RaNgJZ0x9_0;
	wire w_dff_A_WZtzsak76_2;
	wire w_dff_A_cT7U8lKk6_0;
	wire w_dff_A_suS6PqyK1_0;
	wire w_dff_A_PInrur1m3_0;
	wire w_dff_A_neArHU5K6_0;
	wire w_dff_A_50ZKOalW7_0;
	wire w_dff_A_27h0MhW31_0;
	wire w_dff_A_kMTM2Ou99_0;
	wire w_dff_A_bJc3GcsB8_0;
	wire w_dff_A_jm0biYLj5_0;
	wire w_dff_A_JytWYUNK9_0;
	wire w_dff_A_Z2F8HuOt0_0;
	wire w_dff_A_WNgr8LQn6_0;
	wire w_dff_A_os8tY1mZ1_0;
	wire w_dff_A_jZmj1A6T9_0;
	wire w_dff_A_x1YibhHq6_0;
	wire w_dff_A_eLgRMScw4_0;
	wire w_dff_A_aqgWgVCw7_2;
	wire w_dff_A_O1rFA57x9_0;
	wire w_dff_A_7PQ4g2Kp1_0;
	wire w_dff_A_9Qe5Fee53_0;
	wire w_dff_A_4ToV2gLw2_0;
	wire w_dff_A_VfvOAFy55_0;
	wire w_dff_A_XbPDiyvr6_0;
	wire w_dff_A_MC29mWjU4_0;
	wire w_dff_A_h5ic0Zw61_0;
	wire w_dff_A_Lav6XARH1_0;
	wire w_dff_A_YHyRqu6v2_0;
	wire w_dff_A_E98IyfpV3_0;
	wire w_dff_A_HzqF36XT4_0;
	wire w_dff_A_XZoiT8XU2_0;
	wire w_dff_A_Z16LTNoq6_0;
	wire w_dff_A_ExzIBIS38_1;
	wire w_dff_A_dtNI1rGH3_0;
	wire w_dff_A_FNDp067N1_0;
	wire w_dff_A_xV7j1vtZ2_0;
	wire w_dff_A_Mbdo1fJG4_0;
	wire w_dff_A_FwPVKu9g9_0;
	wire w_dff_A_vV9WBLU51_0;
	wire w_dff_A_7IbmsY3R9_0;
	wire w_dff_A_3TYXNsXY0_0;
	wire w_dff_A_1wyZqhUV3_0;
	wire w_dff_A_4w8sKzXo0_0;
	wire w_dff_A_NJ3Sotag4_0;
	wire w_dff_A_DbYTJV8b8_0;
	wire w_dff_A_hQ1JA2t21_0;
	wire w_dff_A_1ur4pzOk2_0;
	wire w_dff_A_R0NBYpVr0_0;
	wire w_dff_A_hmiUOb7Z4_0;
	wire w_dff_A_ow0Cb9UT8_0;
	wire w_dff_A_cvczcfHv9_0;
	wire w_dff_A_m0IDceCV9_0;
	wire w_dff_A_sinQH8b84_0;
	wire w_dff_A_eF25cZUD2_1;
	wire w_dff_A_NT17urFK9_0;
	wire w_dff_A_IxLx04z91_0;
	wire w_dff_A_5wUPmnbG6_0;
	wire w_dff_A_icRxBarg5_0;
	wire w_dff_A_Mam7M0j77_0;
	wire w_dff_A_qRNFJs2l4_0;
	wire w_dff_A_2UFy3Wgo0_0;
	wire w_dff_A_KpDxxA5a9_0;
	wire w_dff_A_RmcJZGW83_0;
	wire w_dff_A_l1OlhjxF7_0;
	wire w_dff_A_2zAfa6a85_0;
	wire w_dff_A_B4Pxk3qv3_0;
	wire w_dff_A_j1qw7Aax9_0;
	wire w_dff_A_ZL6gaiFr9_0;
	wire w_dff_A_zAWVk2s33_0;
	wire w_dff_A_Yw9bDhUO8_0;
	wire w_dff_A_Zi4ClYjW8_0;
	wire w_dff_A_aIZ3bLTn5_0;
	wire w_dff_A_tv8cw3Th2_0;
	wire w_dff_A_Tz0ymolQ7_0;
	wire w_dff_A_mfoVLXEC9_2;
	wire w_dff_A_agD0E8LR5_0;
	wire w_dff_A_eEYs9Fey2_0;
	wire w_dff_A_4gBT5zXA3_0;
	wire w_dff_A_EP4GlbTC9_0;
	wire w_dff_A_eBdOUDx58_0;
	wire w_dff_A_bgH74ekf0_0;
	wire w_dff_A_T5NmPRPy0_0;
	wire w_dff_A_oMBoHOQK8_0;
	wire w_dff_A_BzwpgGgq8_0;
	wire w_dff_A_PjLHKwBi4_0;
	wire w_dff_A_PXBX8FA26_0;
	wire w_dff_A_qJmjJP2c4_2;
	wire w_dff_A_qXRAtiND2_0;
	wire w_dff_A_Jbk10W3U2_0;
	wire w_dff_A_RHWDoGBm5_0;
	wire w_dff_A_2mJQbMZB9_0;
	wire w_dff_A_fyVjTgFU0_0;
	wire w_dff_A_kIpIJOjR6_0;
	wire w_dff_A_jyJCDh204_0;
	wire w_dff_A_aM6fNRj28_0;
	wire w_dff_A_v4gygKSV0_0;
	wire w_dff_A_KTkZyOXT9_0;
	wire w_dff_A_k4ucQ4pX3_0;
	wire w_dff_A_yfLRIfqS6_2;
	wire w_dff_A_1xgzYpP76_0;
	wire w_dff_A_zPAqavb28_0;
	wire w_dff_A_FNI2N5oB0_0;
	wire w_dff_A_qxSqAmE30_0;
	wire w_dff_A_5kmgiiRM4_0;
	wire w_dff_A_fZpHNZqr8_0;
	wire w_dff_A_1O928NQu3_0;
	wire w_dff_A_C6KvVvRw4_0;
	wire w_dff_A_NzqAHX8J0_0;
	wire w_dff_A_xhWMExsS6_0;
	wire w_dff_A_D0YIkcmq8_0;
	wire w_dff_A_pW3zWuB61_2;
	wire w_dff_A_iuhgNjMk9_0;
	wire w_dff_A_0btv8qbN4_0;
	wire w_dff_A_Fvk6Rn4J5_0;
	wire w_dff_A_ucJdm4dT2_0;
	wire w_dff_A_qkcwqVzg9_0;
	wire w_dff_A_dFplCsJf4_0;
	wire w_dff_A_8JPelck91_0;
	wire w_dff_A_PRTB8Ws46_0;
	wire w_dff_A_U2gk24EX5_0;
	wire w_dff_A_TDcCbFpz4_0;
	wire w_dff_A_jytQ3geU6_0;
	wire w_dff_A_St9eEOx71_1;
	wire w_dff_A_28mVbJ1Z5_0;
	wire w_dff_A_goPkPOBL5_0;
	wire w_dff_A_b7hYGBal6_0;
	wire w_dff_A_YlYZW9CP0_0;
	wire w_dff_A_54xN6qlU2_0;
	wire w_dff_A_1EkmCJbj1_0;
	wire w_dff_A_dhvbG9Hp7_0;
	wire w_dff_A_Toz8Cyf38_0;
	wire w_dff_A_9z8b24NF3_0;
	wire w_dff_A_Oi2rYkvS8_0;
	wire w_dff_A_TZIFYD3p2_0;
	wire w_dff_A_3B1wfRkm1_0;
	wire w_dff_A_zkPkpbQs3_0;
	wire w_dff_A_kQaVA9b58_0;
	wire w_dff_A_080eNj162_0;
	wire w_dff_A_gbqxKkWf3_0;
	wire w_dff_A_mWCct4wI7_0;
	wire w_dff_A_7peJnpA54_0;
	wire w_dff_A_YdqD4BPM6_1;
	wire w_dff_A_HTJ3dgCR4_0;
	wire w_dff_A_uZRmZeWc7_0;
	wire w_dff_A_5NiqtKD21_0;
	wire w_dff_A_ZbxeuFVB9_0;
	wire w_dff_A_v6c3OxBq7_0;
	wire w_dff_A_IaM5GIxE4_0;
	wire w_dff_A_mX0o1eqC2_0;
	wire w_dff_A_zqHrxjU17_0;
	wire w_dff_A_kq9v8JyC2_0;
	wire w_dff_A_JwpVFd7m3_0;
	wire w_dff_A_wEb8cgZo2_0;
	wire w_dff_A_mmNzRu3N0_0;
	wire w_dff_A_wwsAQM7y3_0;
	wire w_dff_A_WRqjnmJp9_0;
	wire w_dff_A_Y9r4UMe27_0;
	wire w_dff_A_RD1lG3ow5_0;
	wire w_dff_A_ltiR10Xa4_0;
	wire w_dff_A_CnsGiYrK3_1;
	wire w_dff_A_83EKGves6_0;
	wire w_dff_A_vJPsZl701_0;
	wire w_dff_A_y2Xoglld7_0;
	wire w_dff_A_8SvZ74Qm2_0;
	wire w_dff_A_pOp9XGEc4_0;
	wire w_dff_A_C6CLZAK44_0;
	wire w_dff_A_fq9BW8Aj6_0;
	wire w_dff_A_UlaYkN8l8_0;
	wire w_dff_A_DhcYCfRX8_0;
	wire w_dff_A_4llKW2k82_0;
	wire w_dff_A_Z9I3IhsS7_0;
	wire w_dff_A_uy0SWKff0_0;
	wire w_dff_A_eaUrWHnD8_0;
	wire w_dff_A_LbwBuooE3_0;
	wire w_dff_A_SwDsi6jB6_0;
	wire w_dff_A_NXQF4HCr1_0;
	wire w_dff_A_yjsLMZjX3_0;
	wire w_dff_A_k5yPLMrJ3_1;
	wire w_dff_A_fvq3IfaD1_0;
	wire w_dff_A_k6II2E9H3_0;
	wire w_dff_A_sa7mXR8O1_0;
	wire w_dff_A_aINk9Eez8_0;
	wire w_dff_A_JFc5wbhj1_0;
	wire w_dff_A_kwa8IYkA3_0;
	wire w_dff_A_GvPDbonV7_2;
	wire w_dff_A_nOSyCAkd3_0;
	wire w_dff_A_jU9lzuWV8_0;
	wire w_dff_A_PKIvM7vx3_0;
	wire w_dff_A_ZQ72ZoxQ3_0;
	wire w_dff_A_cviQh5KU4_0;
	wire w_dff_A_Ynk9Rojw0_0;
	wire w_dff_A_8BGQ4quh3_0;
	wire w_dff_A_WXGd0sNX2_0;
	wire w_dff_A_3Wg9Z3FU3_0;
	wire w_dff_A_Ic59kQtS7_0;
	wire w_dff_A_BWxXN7Q49_0;
	wire w_dff_A_599oNvDw3_0;
	wire w_dff_A_wDus7Xlx0_0;
	wire w_dff_A_zizyxwgW1_0;
	wire w_dff_A_ZffOHOwP8_1;
	wire w_dff_A_oW5c9Yys4_0;
	wire w_dff_A_aoX9PM4h8_0;
	wire w_dff_A_l1oc758E6_0;
	wire w_dff_A_5fYMrykJ1_0;
	wire w_dff_A_GINYGC9z5_0;
	wire w_dff_A_A6p88IdL0_0;
	wire w_dff_A_0QIqRIev7_0;
	wire w_dff_A_p4Ml6w9n1_0;
	wire w_dff_A_p2ELthUi3_0;
	wire w_dff_A_U0md0XSE7_0;
	wire w_dff_A_8CNkI0eU4_0;
	wire w_dff_A_msTcj59W3_1;
	wire w_dff_A_G5MbsiEP4_0;
	wire w_dff_A_bOsgKylV9_0;
	wire w_dff_A_30rWTXLk2_0;
	wire w_dff_A_6X6SDLcT4_0;
	wire w_dff_A_jUpFiyuG7_0;
	wire w_dff_A_ZTjhmtnF4_0;
	wire w_dff_A_kFPYv3nn6_0;
	wire w_dff_A_sNo9Dghe2_0;
	wire w_dff_A_HiM0Gdkd7_0;
	wire w_dff_A_oTtU9Rbv7_0;
	wire w_dff_A_SWTTSma93_0;
	wire w_dff_A_0XJcPhsN7_0;
	wire w_dff_A_tkE1fDqo8_0;
	wire w_dff_A_DncwKVdg0_1;
	wire w_dff_A_tnnEG8Ec3_0;
	wire w_dff_A_9RApjLTs8_0;
	wire w_dff_A_vGznwiUd3_0;
	wire w_dff_A_2ITdwgpn3_0;
	wire w_dff_A_NLL83CuD4_0;
	wire w_dff_A_ncehto3S7_0;
	wire w_dff_A_kas13WDr1_0;
	wire w_dff_A_XHruMOpB4_0;
	wire w_dff_A_r1SwHZWk8_0;
	wire w_dff_A_Sq7VWW7F2_0;
	wire w_dff_A_duDx3le64_0;
	wire w_dff_A_DL6aqxX38_0;
	wire w_dff_A_eFrnj7hA1_0;
	wire w_dff_A_NVcIuwAK2_0;
	wire w_dff_A_8Sppg9R88_0;
	wire w_dff_A_8TrmV4bo1_2;
	wire w_dff_A_fzwUM4R65_0;
	wire w_dff_A_0TgI2VJp1_0;
	wire w_dff_A_exINZv4C0_0;
	wire w_dff_A_FUM9BEya1_0;
	wire w_dff_A_TRWfubfV1_0;
	wire w_dff_A_XH9IXdoh1_0;
	wire w_dff_A_C4theoMg4_0;
	wire w_dff_A_lfP9KjOp0_0;
	wire w_dff_A_IGWmh2l21_0;
	wire w_dff_A_yOj7mIoi4_0;
	wire w_dff_A_oqpB9X5S2_0;
	wire w_dff_A_gdq1cazK1_0;
	wire w_dff_A_6MRdUHit8_0;
	wire w_dff_A_NrW5qRyb0_0;
	wire w_dff_A_IXVtm8zU8_1;
	wire w_dff_A_mB5v21pN5_0;
	wire w_dff_A_sTsNouiN8_0;
	wire w_dff_A_S4my90vB1_0;
	wire w_dff_A_cwFEfvcJ1_0;
	wire w_dff_A_EoNNZtM72_0;
	wire w_dff_A_rlLH4CzB7_0;
	wire w_dff_A_DXI2DKSU4_0;
	wire w_dff_A_8aLZA2Wn5_0;
	wire w_dff_A_hEMT2bfT0_0;
	wire w_dff_A_NIZhYMSx1_1;
	wire w_dff_A_jFbfgyKv5_0;
	wire w_dff_A_eh8TOSl19_0;
	wire w_dff_A_1bpmZKHO7_0;
	wire w_dff_A_8NmM8OaC8_0;
	wire w_dff_A_GfU1i5mF8_0;
	wire w_dff_A_vnlUsT7q5_0;
	wire w_dff_A_eqLJrOBc0_0;
	wire w_dff_A_gd9cEWXz6_0;
	wire w_dff_A_MXURVI2L3_0;
	wire w_dff_A_TSBzS8134_0;
	wire w_dff_A_o2n5yBar4_0;
	wire w_dff_A_wxyThvto1_1;
	wire w_dff_A_Oq0L4EC19_0;
	wire w_dff_A_fXrKLlaH6_0;
	wire w_dff_A_T4RqAqNP5_0;
	wire w_dff_A_DJcXeLtS2_0;
	wire w_dff_A_VNLv3DNN9_0;
	wire w_dff_A_4PTJZ3kK0_0;
	wire w_dff_A_TP6gSsnx5_0;
	wire w_dff_A_gbDFa50o7_0;
	wire w_dff_A_KRg67GBY7_0;
	wire w_dff_A_7ghoOdvN1_0;
	wire w_dff_A_ZL9nOHXE2_0;
	wire w_dff_A_ohaO0QbP3_0;
	wire w_dff_A_y2fvlRfV5_1;
	wire w_dff_A_LnYSCbXn9_0;
	wire w_dff_A_f6lpTfON3_0;
	wire w_dff_A_CciD38DR3_0;
	wire w_dff_A_LrwxJvo53_0;
	wire w_dff_A_eNXeGQas8_0;
	wire w_dff_A_o6GTmLG27_0;
	wire w_dff_A_PFpfjHWI0_0;
	wire w_dff_A_kuafdsuF8_0;
	wire w_dff_A_SHCZbjsl4_0;
	wire w_dff_A_miEUHJyN4_0;
	wire w_dff_A_I8dm8M1B8_0;
	wire w_dff_A_vvM4LYCS8_0;
	wire w_dff_A_N3gyNNC57_0;
	wire w_dff_A_hy3XRMt16_1;
	wire w_dff_A_nlJ6vhn78_0;
	wire w_dff_A_YgsIYrS27_0;
	wire w_dff_A_sVtdwruG0_0;
	wire w_dff_A_TvKM6GDk6_0;
	wire w_dff_A_By65h7ve9_0;
	wire w_dff_A_q2ep5t2e9_0;
	wire w_dff_A_6pvA1WnF9_0;
	wire w_dff_A_ZG5ktrdT5_0;
	wire w_dff_A_EKkAAozQ3_0;
	wire w_dff_A_LqGWjEKb4_0;
	wire w_dff_A_yyBRG0eW2_0;
	wire w_dff_A_3cu7Ywe51_0;
	wire w_dff_A_wBIAyGJL9_0;
	wire w_dff_A_ocAGjrj65_0;
	wire w_dff_A_lavgTu5v9_0;
	wire w_dff_A_z2no7W9H4_0;
	wire w_dff_A_yV3M3vWw4_1;
	wire w_dff_A_nxPx0cIa5_0;
	wire w_dff_A_5kYh2G7x1_0;
	wire w_dff_A_T8lqoWCL7_0;
	wire w_dff_A_Ypktngn25_0;
	wire w_dff_A_slSZQgGt1_0;
	wire w_dff_A_l5VXW8zM2_0;
	wire w_dff_A_4hkbVbUF9_0;
	wire w_dff_A_4Hk71Rpv7_0;
	wire w_dff_A_wcunGtT17_0;
	wire w_dff_A_njRTuOBR8_0;
	wire w_dff_A_slk0RpSk6_0;
	wire w_dff_A_pfBskIu99_0;
	wire w_dff_A_OhDAgSNI0_0;
	wire w_dff_A_PIs04hum8_0;
	wire w_dff_A_8LmpDHTm3_0;
	wire w_dff_A_A6MBRDD45_0;
	wire w_dff_A_DHHKKRtK9_0;
	wire w_dff_A_wcbljaey5_0;
	wire w_dff_A_rzj3Gxf21_2;
	wire w_dff_A_S48jCoEZ7_0;
	wire w_dff_A_436cEISi1_0;
	wire w_dff_A_MX9ZfvsT3_0;
	wire w_dff_A_KSpr5fVE0_0;
	wire w_dff_A_OurWUoh22_2;
	wire w_dff_A_a4YtDaw40_0;
	wire w_dff_A_6pYyqoxk1_0;
	wire w_dff_A_ThUQVMEj6_0;
	wire w_dff_A_SHcAE3dZ9_0;
	wire w_dff_A_GT0N0tKO8_0;
	wire w_dff_A_P9zOJhhd5_0;
	wire w_dff_A_M4wuqmaJ9_0;
	wire w_dff_A_CdLv686k3_2;
	wire w_dff_A_wVnRgiAg5_0;
	wire w_dff_A_Rv1xzE9Q1_0;
	wire w_dff_A_t8FSO4NZ3_0;
	wire w_dff_A_qvkchFAl0_0;
	wire w_dff_A_IBXzG8LL3_0;
	wire w_dff_A_Am64hqcN0_0;
	wire w_dff_A_XBItEODN1_0;
	wire w_dff_A_YY3Ejfev2_0;
	wire w_dff_A_xvs258ej6_0;
	wire w_dff_A_pAvuaBLZ7_0;
	wire w_dff_A_yYjyoZsI5_0;
	wire w_dff_A_W6VhlTt27_0;
	wire w_dff_A_wuqM8eDK6_0;
	wire w_dff_A_eISRmwvG1_2;
	wire w_dff_A_DuJnvwwJ7_0;
	wire w_dff_A_IhZ6kUNN7_0;
	wire w_dff_A_79epYESg6_0;
	wire w_dff_A_xNo22IQ48_0;
	wire w_dff_A_mbfguTpo1_0;
	wire w_dff_A_TyWnQ3Gf6_0;
	wire w_dff_A_qtOORKx37_0;
	wire w_dff_A_iIR2E4HM4_0;
	wire w_dff_A_vo6ZiUby3_0;
	wire w_dff_A_55iAiWu90_0;
	wire w_dff_A_3oMyx8CQ1_0;
	wire w_dff_A_z9amqPRY5_0;
	wire w_dff_A_GzH6xKpN8_0;
	wire w_dff_A_pbgvSBrL9_2;
	wire w_dff_A_yXroYVSS5_0;
	wire w_dff_A_GCfkkTRs0_0;
	wire w_dff_A_v7RLv10f3_0;
	wire w_dff_A_vMTtlUYk2_0;
	wire w_dff_A_wFZsi1fI6_0;
	wire w_dff_A_BhPHxHby8_0;
	wire w_dff_A_eFLyZN3r9_2;
	wire w_dff_A_qO2PfSKg0_0;
	wire w_dff_A_YYQfVngw2_0;
	wire w_dff_A_tFBjUQuU0_0;
	wire w_dff_A_iB1mXwn10_0;
	wire w_dff_A_Sxr1TNJc6_0;
	wire w_dff_A_aU2zvkL33_0;
	wire w_dff_A_MrPJLRpt8_0;
	wire w_dff_A_QTOLHuFS9_0;
	wire w_dff_A_SmweK2rc4_2;
	wire w_dff_A_kCf0gnem7_0;
	wire w_dff_A_mncjqRI36_0;
	wire w_dff_A_J6oIVXMM4_0;
	wire w_dff_A_wv7nFki81_0;
	wire w_dff_A_D4g7LYgi0_0;
	wire w_dff_A_XyJRopmA2_0;
	wire w_dff_A_7oUpz2pl4_0;
	wire w_dff_A_11VyRUfz4_0;
	wire w_dff_A_vNTKL5wL6_0;
	wire w_dff_A_19H5GxO39_2;
	wire w_dff_A_CkplTEF39_0;
	wire w_dff_A_VpQ895LF5_0;
	wire w_dff_A_LPzmIaxm7_0;
	wire w_dff_A_T98IUh9p5_0;
	wire w_dff_A_kEinjJWw5_0;
	wire w_dff_A_p35Tfkqo2_0;
	wire w_dff_A_CF4nTgrd4_0;
	wire w_dff_A_333Bxx204_0;
	wire w_dff_A_vIISzsln7_0;
	wire w_dff_A_vXSVgGy34_0;
	wire w_dff_A_pYaVT0Rd8_2;
	wire w_dff_A_Pf47elGq7_0;
	wire w_dff_A_Cq73wuwD4_0;
	wire w_dff_A_gJojppiQ8_0;
	wire w_dff_A_RbW9zctz4_0;
	wire w_dff_A_6l2Ydi907_0;
	wire w_dff_A_05xG1v6s4_0;
	wire w_dff_A_zWQ5oN7u7_2;
	wire w_dff_A_kZqLK9Oe2_0;
	wire w_dff_A_RrjdQ1Ie4_0;
	wire w_dff_A_f81B8eNJ3_0;
	wire w_dff_A_Xjvw3LUK6_0;
	wire w_dff_A_0DkL6X2v5_0;
	wire w_dff_A_UHprJJi11_0;
	wire w_dff_A_bZ7fGTv52_0;
	wire w_dff_A_cxwBHQIU5_0;
	wire w_dff_A_3Phyc5ei6_2;
	wire w_dff_A_fbbGPwTf2_0;
	wire w_dff_A_OSuH9g8x7_0;
	wire w_dff_A_Gv1QOu920_0;
	wire w_dff_A_ZTMCKfLC4_0;
	wire w_dff_A_N6lVp1zz8_0;
	wire w_dff_A_ezaOVLRV0_0;
	wire w_dff_A_bmrWEQNl7_0;
	wire w_dff_A_xHk89ZmV2_0;
	wire w_dff_A_i4XbFAfI4_0;
	wire w_dff_A_kR71S9B18_2;
	wire w_dff_A_aCA6XL235_0;
	wire w_dff_A_TakHbnji0_0;
	wire w_dff_A_QJtBWF2X1_0;
	wire w_dff_A_KW4ljHCu3_0;
	wire w_dff_A_Ru72osg75_0;
	wire w_dff_A_IenheodB6_0;
	wire w_dff_A_MCNNZQST9_0;
	wire w_dff_A_Lwtw3oUA6_0;
	wire w_dff_A_vBUBildu3_0;
	wire w_dff_A_T5KTvmcx1_0;
	wire w_dff_A_K4P7N6hP0_2;
	wire w_dff_A_EMuOqUc83_0;
	wire w_dff_A_I0icv16C9_0;
	wire w_dff_A_AqOhtOe31_0;
	wire w_dff_A_rRZTnKA65_0;
	wire w_dff_A_AkyEd3kP8_0;
	wire w_dff_A_ezoq8C9i9_2;
	wire w_dff_A_r7ofSOrF0_0;
	wire w_dff_A_JfKnqpVd0_0;
	wire w_dff_A_gkw2YFHw9_0;
	wire w_dff_A_HwHOl2M93_0;
	wire w_dff_A_8bQOTEfo0_0;
	wire w_dff_A_taEuKB0R6_0;
	wire w_dff_A_w2qqhGHj4_0;
	wire w_dff_A_8Xgfz7I19_0;
	wire w_dff_A_3St8Wg039_0;
	wire w_dff_A_gnv61TFV1_2;
	wire w_dff_A_mMfZiepW4_0;
	wire w_dff_A_CkU8mcFC0_0;
	wire w_dff_A_9SL0YjeN3_0;
	wire w_dff_A_lH1SOfWF7_0;
	wire w_dff_A_GkkDKFhC6_0;
	wire w_dff_A_ezHOAA2O4_0;
	wire w_dff_A_gC63kOGS8_0;
	wire w_dff_A_QTUfGkKg6_0;
	wire w_dff_A_rJmF9iXA4_2;
	wire w_dff_A_wuCNB4UR3_0;
	wire w_dff_A_CUGWhDlB8_0;
	wire w_dff_A_j4GLjSqq9_0;
	wire w_dff_A_eva3bVmB9_0;
	wire w_dff_A_jRtr63dN5_0;
	wire w_dff_A_IpUQfIyO6_0;
	wire w_dff_A_roGkLfMO2_0;
	wire w_dff_A_Ox1Xngjw7_2;
	wire w_dff_A_CI8vtukZ7_0;
	wire w_dff_A_fSKr5kwp3_0;
	wire w_dff_A_LVci0KQs4_0;
	wire w_dff_A_EFKPCJSO0_0;
	wire w_dff_A_8A0phuLi9_0;
	wire w_dff_A_McN35ANS3_2;
	wire w_dff_A_BosRwV852_0;
	wire w_dff_A_qlzsTmU16_0;
	wire w_dff_A_W79NsMZG5_0;
	wire w_dff_A_6txG9rdT9_0;
	wire w_dff_A_kzKdnUt37_0;
	wire w_dff_A_2NJkJHVQ0_0;
	wire w_dff_A_qWXZYGSi6_0;
	wire w_dff_A_o0iUeAoK2_0;
	wire w_dff_A_5qvAay5z2_0;
	wire w_dff_A_EEV2iFkR2_2;
	wire w_dff_A_t7TnUSKN7_0;
	wire w_dff_A_1fQoPR9M5_0;
	wire w_dff_A_fiJjTg9N5_0;
	wire w_dff_A_zW4POg2M2_0;
	wire w_dff_A_U8jJeBae8_0;
	wire w_dff_A_mC2kIqIz9_0;
	wire w_dff_A_k1mwG7fn4_0;
	wire w_dff_A_hP4eKqU42_0;
	wire w_dff_A_x965G86B7_2;
	wire w_dff_A_zXf9E0Og1_0;
	wire w_dff_A_70xlT3x62_0;
	wire w_dff_A_Lm8y4DcO9_0;
	wire w_dff_A_a06eyMM67_0;
	wire w_dff_A_eeeVtZlV6_0;
	wire w_dff_A_3r2jDFcY2_0;
	wire w_dff_A_w55egnzk1_0;
	wire w_dff_A_YIjMVBcl3_2;
	wire w_dff_A_YDP4YiCG6_0;
	wire w_dff_A_BX6lASSb2_0;
	wire w_dff_A_K6m8maJW8_0;
	wire w_dff_A_KrXez6WB0_0;
	wire w_dff_A_VUuDR6GP3_2;
	wire w_dff_A_2UUTflwp7_0;
	wire w_dff_A_AqNe3o8C0_0;
	wire w_dff_A_cJHUWzDP6_0;
	wire w_dff_A_ZQGg0kSb7_0;
	wire w_dff_A_UJdi8eDm4_0;
	wire w_dff_A_cRGRjQb90_0;
	wire w_dff_A_jx2THHHv0_0;
	wire w_dff_A_55bRIRtq1_0;
	wire w_dff_A_dRifuz8t7_1;
	wire w_dff_A_Lj2wljKi8_0;
	wire w_dff_A_n9v9kLba2_0;
	wire w_dff_A_L1aXTwpM2_0;
	wire w_dff_A_5hZJmb488_0;
	wire w_dff_A_8Pa9YStv0_1;
	wire w_dff_A_8FDlU7Z94_0;
	wire w_dff_A_YA723v3U1_0;
	wire w_dff_A_dKnmV6xp3_0;
	wire w_dff_A_4f4smzWv7_0;
	wire w_dff_A_r2WU4mxa7_0;
	wire w_dff_A_0eCZVfks5_0;
	wire w_dff_A_unZc6zDF5_0;
	wire w_dff_A_WWL5M9oO4_1;
	wire w_dff_A_MwQ62wHi0_0;
	wire w_dff_A_bXXqA2gj0_0;
	wire w_dff_A_vQzWbjcD8_0;
	wire w_dff_A_89pAjEOo2_0;
	wire w_dff_A_Z6Md5XyQ1_0;
	wire w_dff_A_V6uqVzyG3_0;
	wire w_dff_A_L7SR8ykS2_0;
	wire w_dff_A_mLyNlAgr2_1;
	wire w_dff_A_mraoG5du0_0;
	wire w_dff_A_YEawgPrx4_0;
	wire w_dff_A_B7gsoJio3_0;
	wire w_dff_A_uV8eFwMf2_0;
	wire w_dff_A_nGiSCrPh2_0;
	wire w_dff_A_8Ynurn2G0_0;
	wire w_dff_A_gxQ3cpsS0_0;
	wire w_dff_A_aljJRhok0_0;
	wire w_dff_A_dWiR3lKc9_2;
	wire w_dff_A_REBnqDrA5_0;
	wire w_dff_A_sKBWvyPh9_0;
	wire w_dff_A_5ToOHbWm8_0;
	wire w_dff_A_LoIhxFRI9_0;
	wire w_dff_A_2HMndqNF9_0;
	wire w_dff_A_WS56Qo9Z5_0;
	wire w_dff_A_6UAEFGew6_0;
	wire w_dff_A_SYj6CJqL4_0;
	wire w_dff_A_hV5cQzcV5_0;
	wire w_dff_A_eyz1tPcM8_0;
	wire w_dff_A_oe773Z964_0;
	wire w_dff_A_HBm8Pqso5_0;
	wire w_dff_A_WPtnuktD0_0;
	wire w_dff_A_3ikstzRv4_0;
	wire w_dff_A_5gC9Os1p4_0;
	wire w_dff_A_YbUu0rt76_1;
	wire w_dff_A_uMJxHwHR9_0;
	wire w_dff_A_ELEPugdY3_0;
	wire w_dff_A_Cn3iv0w64_0;
	wire w_dff_A_jFPW27Js2_1;
	wire w_dff_A_XD6j3chI0_0;
	wire w_dff_A_z6FqgfEj7_0;
	wire w_dff_A_LFRXAEMs0_0;
	wire w_dff_A_EMv9EHTg6_0;
	wire w_dff_A_yZxRu1CP2_1;
	wire w_dff_A_t0UT0z536_0;
	wire w_dff_A_wyGvadyG9_0;
	wire w_dff_A_8R4oR8H47_0;
	wire w_dff_A_JPMgzgEx2_0;
	wire w_dff_A_Q7zqQz1Q8_0;
	wire w_dff_A_CR2Xnq2k7_0;
	wire w_dff_A_3kPjIFex3_1;
	wire w_dff_A_asAFbCei9_0;
	wire w_dff_A_cCdNDXPH6_0;
	wire w_dff_A_XvoRUMQB7_0;
	wire w_dff_A_XErBjIMI5_0;
	wire w_dff_A_LUW5uCGe2_0;
	wire w_dff_A_c6BudVkf4_0;
	wire w_dff_A_c349SEMu3_0;
	wire w_dff_A_nWpQUXif7_2;
	wire w_dff_A_qnQCP2FW6_0;
	wire w_dff_A_w46jqcqI5_0;
	wire w_dff_A_wC6dLpOY8_2;
	wire w_dff_A_DJoEsS8a5_0;
	wire w_dff_A_ZDnS8Dex4_0;
	wire w_dff_A_aOg13yvN6_2;
	wire w_dff_A_BoKCrHaW0_0;
	wire w_dff_A_iJi8hbqm4_0;
	wire w_dff_A_jjn7m34c5_0;
	wire w_dff_A_Gz7SUmwg3_2;
	wire w_dff_A_vR67JDpJ5_0;
	wire w_dff_A_gKNKnbk48_0;
	wire w_dff_A_WOszV7J96_0;
	wire w_dff_A_Kj9RkwBZ2_2;
	wire w_dff_A_YAt4ZZqV2_0;
	wire w_dff_A_en51KzfX7_0;
	wire w_dff_A_5aBGWT594_0;
	wire w_dff_A_SC7UKnfq8_0;
	wire w_dff_A_r913b9Tx0_2;
	wire w_dff_A_MyLslFcV2_0;
	wire w_dff_A_KyIDrp7O3_0;
	wire w_dff_A_MUyDFMxZ5_0;
	wire w_dff_A_B7zzNCht4_2;
	wire w_dff_A_gzPPoZzQ1_0;
	wire w_dff_A_Pb2PdW7y6_0;
	wire w_dff_A_3L2PEZOQ6_0;
	wire w_dff_A_zAFhLVgo8_2;
	wire w_dff_A_PHqc0E8t0_0;
	wire w_dff_A_qPJeZuC07_0;
	wire w_dff_A_qmraD4Nd5_0;
	wire w_dff_A_btpGjl9F0_0;
	wire w_dff_A_IHkscreG0_2;
	wire w_dff_A_vvc2VZZb5_0;
	wire w_dff_A_AcozqTrH7_0;
	wire w_dff_A_Po0WJqnD9_0;
	wire w_dff_A_waPH8W0z0_2;
	wire w_dff_A_W3CeAKtQ5_0;
	wire w_dff_A_8F4EYnfM6_0;
	wire w_dff_A_Ma7drrNq3_2;
	wire w_dff_A_To0ayZgd9_0;
	wire w_dff_A_4p4Wrc8s2_0;
	wire w_dff_A_CSW3oR7E2_2;
	wire w_dff_A_ZApLNaRm5_0;
	wire w_dff_A_jCh5PqgI7_2;
	wire w_dff_A_LQ1RT4Xg3_0;
	wire w_dff_A_1TfznRbi4_0;
	wire w_dff_A_yIsjDxSq4_0;
	wire w_dff_A_QI9HYEpX5_2;
	wire w_dff_A_TD904Lgl4_0;
	wire w_dff_A_6eNES9vT4_0;
	wire w_dff_A_MbjnhRRh3_2;
	wire w_dff_A_qARrPKVs1_0;
	wire w_dff_A_seMwHF2r9_0;
	wire w_dff_A_j5GasjKW1_2;
	wire w_dff_A_rwYucOoo7_0;
	wire w_dff_A_JuKIKgog1_2;
	wire w_dff_A_xoyA0ozh6_0;
	wire w_dff_A_YZNLLjuP3_0;
	wire w_dff_A_novSlxr97_0;
	wire w_dff_A_fExTKHZC7_2;
	wire w_dff_A_udOtkEGA8_0;
	wire w_dff_A_lIrjR9Jj0_0;
	wire w_dff_A_0Qtxkv1O2_0;
	wire w_dff_A_1182Ow2c0_2;
	wire w_dff_A_GtGQe1WM9_2;
	jnot g0000(.din(w_G545_0[2]),.dout(w_dff_A_x1fDTMpv4_1),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(G366),.dout(G600_fa_),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(w_dff_A_d5oFxJLf5_1),.clk(gclk));
	jnot g0005(.din(G338),.dout(G611_fa_),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(w_dff_A_ngmk1eik7_2),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(w_dff_A_WaFIGnAa9_1),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(w_dff_A_A8hVAlbl2_1),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(w_dff_A_6894XwHg4_1),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(w_dff_A_HHWOph5b7_1),.clk(gclk));
	jand g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(w_dff_A_YkzxoQtB2_2),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_Id93cNMm3_1),.dout(w_dff_A_gMoTHiyF2_2),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jor g0016(.dina(w_dff_B_DSqho5bM5_0),.dinb(w_n316_0[1]),.dout(w_dff_A_YXrgNVZe8_2),.clk(gclk));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(w_dff_A_1vhZ3Duu7_1),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jor g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_),.clk(gclk));
	jor g0022(.dina(w_G809_3[1]),.dinb(w_dff_B_k7loCNst5_1),.dout(w_dff_A_9LMyKtbq7_2),.clk(gclk));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jor g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330),.clk(gclk));
	jor g0030(.dina(n330),.dinb(w_dff_B_gitFSkvp1_1),.dout(w_dff_A_tjW8NLMX1_2),.clk(gclk));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jor g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336),.clk(gclk));
	jor g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(w_dff_A_uZFyizaT3_2),.clk(gclk));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jor g0038(.dina(w_G809_2[1]),.dinb(w_dff_B_lCHdGDBG8_1),.dout(w_dff_A_1RnTGjF92_2),.clk(gclk));
	jand g0039(.dina(w_n326_1[2]),.dinb(w_dff_B_s29xw4Br7_1),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jor g0041(.dina(w_dff_B_WfzLEPFN3_0),.dinb(w_G809_2[0]),.dout(n342),.clk(gclk));
	jor g0042(.dina(n342),.dinb(w_dff_B_3iwXC5Ze8_1),.dout(n343),.clk(gclk));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(w_dff_A_MTvHxVse2_2),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(w_dff_B_hA9gudFc2_1),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jor g0046(.dina(w_dff_B_qQYrjorV2_0),.dinb(w_G809_1[2]),.dout(n347),.clk(gclk));
	jor g0047(.dina(n347),.dinb(w_dff_B_P9Y9rX433_1),.dout(n348),.clk(gclk));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(w_dff_A_QgILRn1A0_2),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(w_dff_B_dQvTcDHr1_1),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jor g0051(.dina(w_dff_B_inkwp1BG9_0),.dinb(w_G809_1[1]),.dout(n352),.clk(gclk));
	jor g0052(.dina(n352),.dinb(w_dff_B_heedTL9O1_1),.dout(n353),.clk(gclk));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(w_dff_A_0GmzN7ei2_2),.clk(gclk));
	jand g0054(.dina(w_n326_0[2]),.dinb(w_dff_B_dQxeAXvO7_1),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_G2358_0[2]),.dinb(G80),.dout(n356),.clk(gclk));
	jor g0056(.dina(w_dff_B_g5ylZoCc8_0),.dinb(w_G809_1[0]),.dout(n357),.clk(gclk));
	jor g0057(.dina(n357),.dinb(w_dff_B_ovleiaxu5_1),.dout(n358),.clk(gclk));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(w_dff_A_0tDgTm6S3_2),.clk(gclk));
	jnot g0059(.din(w_G308_1[2]),.dout(n360),.clk(gclk));
	jand g0060(.dina(w_n360_0[1]),.dinb(w_G251_4[2]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G479_1[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(w_G308_1[1]),.dinb(w_G248_5[1]),.dout(n363),.clk(gclk));
	jor g0063(.dina(n363),.dinb(w_n362_0[1]),.dout(n364),.clk(gclk));
	jor g0064(.dina(n364),.dinb(n361),.dout(n365),.clk(gclk));
	jnot g0065(.din(w_G254_1[2]),.dout(n366),.clk(gclk));
	jand g0066(.dina(w_n360_0[0]),.dinb(w_n366_4[2]),.dout(n367),.clk(gclk));
	jnot g0067(.din(w_G242_1[2]),.dout(n368),.clk(gclk));
	jand g0068(.dina(w_G308_1[0]),.dinb(w_n368_5[1]),.dout(n369),.clk(gclk));
	jor g0069(.dina(n369),.dinb(w_G479_1[0]),.dout(n370),.clk(gclk));
	jor g0070(.dina(n370),.dinb(w_dff_B_niiqv8J41_1),.dout(n371),.clk(gclk));
	jand g0071(.dina(n371),.dinb(w_dff_B_zavP2zuO7_1),.dout(n372),.clk(gclk));
	jnot g0072(.din(w_G316_1[2]),.dout(n373),.clk(gclk));
	jand g0073(.dina(w_n373_0[1]),.dinb(w_G251_4[1]),.dout(n374),.clk(gclk));
	jnot g0074(.din(w_G490_1[2]),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_G316_1[1]),.dinb(w_G248_5[0]),.dout(n376),.clk(gclk));
	jor g0076(.dina(n376),.dinb(n375),.dout(n377),.clk(gclk));
	jor g0077(.dina(n377),.dinb(n374),.dout(n378),.clk(gclk));
	jand g0078(.dina(w_n373_0[0]),.dinb(w_n366_4[1]),.dout(n379),.clk(gclk));
	jand g0079(.dina(w_G316_1[0]),.dinb(w_n368_5[0]),.dout(n380),.clk(gclk));
	jor g0080(.dina(n380),.dinb(w_G490_1[1]),.dout(n381),.clk(gclk));
	jor g0081(.dina(n381),.dinb(w_dff_B_kgP3d0345_1),.dout(n382),.clk(gclk));
	jand g0082(.dina(n382),.dinb(w_dff_B_nUiidziz7_1),.dout(n383),.clk(gclk));
	jand g0083(.dina(w_n383_0[2]),.dinb(w_n372_0[2]),.dout(n384),.clk(gclk));
	jnot g0084(.din(w_G351_2[2]),.dout(n385),.clk(gclk));
	jnot g0085(.din(G3550),.dout(n386),.clk(gclk));
	jand g0086(.dina(w_n386_4[2]),.dinb(w_n385_1[2]),.dout(n387),.clk(gclk));
	jnot g0087(.din(w_G534_1[2]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G3552_0[1]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n389_4[2]),.dinb(w_G351_2[1]),.dout(n390),.clk(gclk));
	jor g0090(.dina(n390),.dinb(w_n388_1[2]),.dout(n391),.clk(gclk));
	jor g0091(.dina(n391),.dinb(w_dff_B_sMPIbE0P2_1),.dout(n392),.clk(gclk));
	jand g0092(.dina(w_G3548_4[2]),.dinb(w_n385_1[1]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3546_5[1]),.dinb(w_G351_2[0]),.dout(n394),.clk(gclk));
	jor g0094(.dina(n394),.dinb(w_G534_1[1]),.dout(n395),.clk(gclk));
	jor g0095(.dina(n395),.dinb(n393),.dout(n396),.clk(gclk));
	jand g0096(.dina(w_dff_B_uOWGZG217_0),.dinb(n392),.dout(n397),.clk(gclk));
	jnot g0097(.din(w_G293_0[2]),.dout(n398),.clk(gclk));
	jand g0098(.dina(w_n398_0[2]),.dinb(w_n366_4[0]),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G293_0[1]),.dinb(w_n368_4[2]),.dout(n400),.clk(gclk));
	jor g0100(.dina(n400),.dinb(n399),.dout(n401),.clk(gclk));
	jnot g0101(.din(w_G251_4[0]),.dout(n402),.clk(gclk));
	jnot g0102(.din(w_G302_0[2]),.dout(n403),.clk(gclk));
	jand g0103(.dina(w_n403_0[1]),.dinb(w_n402_2[1]),.dout(n404),.clk(gclk));
	jnot g0104(.din(w_G248_4[2]),.dout(n405),.clk(gclk));
	jand g0105(.dina(w_G302_0[1]),.dinb(w_n405_2[1]),.dout(n406),.clk(gclk));
	jor g0106(.dina(n406),.dinb(n404),.dout(n407),.clk(gclk));
	jnot g0107(.din(w_n407_0[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_n408_0[1]),.dinb(w_n401_0[2]),.dout(n409),.clk(gclk));
	jnot g0109(.din(w_G514_1[1]),.dout(n410),.clk(gclk));
	jnot g0110(.din(w_G3546_5[0]),.dout(n411),.clk(gclk));
	jand g0111(.dina(n411),.dinb(w_n410_1[1]),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G3552_0[0]),.dinb(w_G514_1[0]),.dout(n413),.clk(gclk));
	jor g0113(.dina(w_dff_B_qYhCDAB74_0),.dinb(n412),.dout(n414),.clk(gclk));
	jnot g0114(.din(w_n414_0[1]),.dout(n415),.clk(gclk));
	jnot g0115(.din(w_G361_0[2]),.dout(n416),.clk(gclk));
	jand g0116(.dina(w_n416_0[1]),.dinb(w_n402_2[0]),.dout(n417),.clk(gclk));
	jand g0117(.dina(w_G361_0[1]),.dinb(w_n405_2[0]),.dout(n418),.clk(gclk));
	jor g0118(.dina(n418),.dinb(n417),.dout(n419),.clk(gclk));
	jnot g0119(.din(w_n419_0[2]),.dout(n420),.clk(gclk));
	jand g0120(.dina(n420),.dinb(n415),.dout(n421),.clk(gclk));
	jand g0121(.dina(n421),.dinb(n409),.dout(n422),.clk(gclk));
	jand g0122(.dina(n422),.dinb(w_n397_0[1]),.dout(n423),.clk(gclk));
	jnot g0123(.din(w_G324_1[2]),.dout(n424),.clk(gclk));
	jand g0124(.dina(w_n386_4[1]),.dinb(w_n424_2[1]),.dout(n425),.clk(gclk));
	jnot g0125(.din(w_G503_1[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_n389_4[1]),.dinb(w_G324_1[1]),.dout(n427),.clk(gclk));
	jor g0127(.dina(n427),.dinb(w_n426_0[1]),.dout(n428),.clk(gclk));
	jor g0128(.dina(n428),.dinb(w_dff_B_fVsMa68i5_1),.dout(n429),.clk(gclk));
	jand g0129(.dina(w_G3548_4[1]),.dinb(w_n424_2[0]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G3546_4[2]),.dinb(w_G324_1[0]),.dout(n431),.clk(gclk));
	jor g0131(.dina(n431),.dinb(w_G503_1[1]),.dout(n432),.clk(gclk));
	jor g0132(.dina(n432),.dinb(n430),.dout(n433),.clk(gclk));
	jand g0133(.dina(w_dff_B_6sGFwgL41_0),.dinb(n429),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G341_2[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n386_4[0]),.dinb(w_n435_1[2]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G523_1[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n389_4[0]),.dinb(w_G341_2[1]),.dout(n438),.clk(gclk));
	jor g0138(.dina(n438),.dinb(w_n437_1[2]),.dout(n439),.clk(gclk));
	jor g0139(.dina(n439),.dinb(w_dff_B_R1DgXB5Q0_1),.dout(n440),.clk(gclk));
	jand g0140(.dina(w_G3548_4[0]),.dinb(w_n435_1[1]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3546_4[1]),.dinb(w_G341_2[0]),.dout(n442),.clk(gclk));
	jor g0142(.dina(n442),.dinb(w_G523_1[0]),.dout(n443),.clk(gclk));
	jor g0143(.dina(n443),.dinb(n441),.dout(n444),.clk(gclk));
	jand g0144(.dina(w_dff_B_XsQtfZjz4_0),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(w_n434_0[1]),.dout(n446),.clk(gclk));
	jand g0146(.dina(w_dff_B_83XCQ04X6_0),.dinb(n423),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(w_dff_B_FuxDKOSc6_1),.dout(w_dff_A_MDA1CyFJ0_2),.clk(gclk));
	jnot g0148(.din(w_G265_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n386_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G400_1[1]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n389_3[2]),.dinb(w_G265_2[0]),.dout(n452),.clk(gclk));
	jor g0152(.dina(n452),.dinb(w_n451_1[1]),.dout(n453),.clk(gclk));
	jor g0153(.dina(n453),.dinb(w_dff_B_WBWgcu617_1),.dout(n454),.clk(gclk));
	jand g0154(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3546_4[0]),.dinb(w_G265_1[2]),.dout(n456),.clk(gclk));
	jor g0156(.dina(n456),.dinb(w_G400_1[0]),.dout(n457),.clk(gclk));
	jor g0157(.dina(n457),.dinb(n455),.dout(n458),.clk(gclk));
	jand g0158(.dina(w_dff_B_Bojb8ccS4_0),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n386_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n389_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jor g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464),.clk(gclk));
	jor g0164(.dina(n464),.dinb(w_dff_B_RqnE4Ckq4_1),.dout(n465),.clk(gclk));
	jand g0165(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n467),.clk(gclk));
	jor g0167(.dina(n467),.dinb(w_G435_1[1]),.dout(n468),.clk(gclk));
	jor g0168(.dina(n468),.dinb(n466),.dout(n469),.clk(gclk));
	jand g0169(.dina(w_dff_B_2SWRVRtF9_0),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G257_2[2]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n386_3[0]),.dinb(w_n471_1[1]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G389_0[2]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n389_3[0]),.dinb(w_G257_2[1]),.dout(n474),.clk(gclk));
	jor g0174(.dina(n474),.dinb(w_n473_1[2]),.dout(n475),.clk(gclk));
	jor g0175(.dina(n475),.dinb(w_dff_B_hGD3gZm12_1),.dout(n476),.clk(gclk));
	jand g0176(.dina(w_G3548_3[0]),.dinb(w_n471_1[0]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3546_3[1]),.dinb(w_G257_2[0]),.dout(n478),.clk(gclk));
	jor g0178(.dina(n478),.dinb(w_G389_0[1]),.dout(n479),.clk(gclk));
	jor g0179(.dina(n479),.dinb(n477),.dout(n480),.clk(gclk));
	jand g0180(.dina(w_dff_B_uuCq0Loz4_0),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jand g0182(.dina(n482),.dinb(w_n459_0[1]),.dout(n483),.clk(gclk));
	jnot g0183(.din(w_G273_2[2]),.dout(n484),.clk(gclk));
	jand g0184(.dina(w_n386_2[2]),.dinb(w_n484_1[1]),.dout(n485),.clk(gclk));
	jnot g0185(.din(w_G411_0[2]),.dout(n486),.clk(gclk));
	jand g0186(.dina(w_n389_2[2]),.dinb(w_G273_2[1]),.dout(n487),.clk(gclk));
	jor g0187(.dina(n487),.dinb(w_n486_1[1]),.dout(n488),.clk(gclk));
	jor g0188(.dina(n488),.dinb(w_dff_B_cYahSXIn8_1),.dout(n489),.clk(gclk));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n484_1[0]),.dout(n490),.clk(gclk));
	jand g0190(.dina(w_G3546_3[0]),.dinb(w_G273_2[0]),.dout(n491),.clk(gclk));
	jor g0191(.dina(n491),.dinb(w_G411_0[1]),.dout(n492),.clk(gclk));
	jor g0192(.dina(n492),.dinb(n490),.dout(n493),.clk(gclk));
	jand g0193(.dina(w_dff_B_zpjQOf2U6_0),.dinb(n489),.dout(n494),.clk(gclk));
	jnot g0194(.din(w_G281_2[1]),.dout(n495),.clk(gclk));
	jand g0195(.dina(w_n386_2[1]),.dinb(w_n495_1[2]),.dout(n496),.clk(gclk));
	jnot g0196(.din(w_G374_0[2]),.dout(n497),.clk(gclk));
	jand g0197(.dina(w_n389_2[1]),.dinb(w_G281_2[0]),.dout(n498),.clk(gclk));
	jor g0198(.dina(n498),.dinb(w_n497_1[1]),.dout(n499),.clk(gclk));
	jor g0199(.dina(n499),.dinb(w_dff_B_ZwRsMymD1_1),.dout(n500),.clk(gclk));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n495_1[1]),.dout(n501),.clk(gclk));
	jand g0201(.dina(w_G3546_2[2]),.dinb(w_G281_1[2]),.dout(n502),.clk(gclk));
	jor g0202(.dina(n502),.dinb(w_G374_0[1]),.dout(n503),.clk(gclk));
	jor g0203(.dina(n503),.dinb(n501),.dout(n504),.clk(gclk));
	jand g0204(.dina(w_dff_B_mvkwBMxs2_0),.dinb(n500),.dout(n505),.clk(gclk));
	jand g0205(.dina(w_n505_0[1]),.dinb(w_n494_0[1]),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[2]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n386_2[0]),.dinb(w_n507_1[1]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n389_2[0]),.dinb(w_G218_2[1]),.dout(n510),.clk(gclk));
	jor g0210(.dina(n510),.dinb(w_n509_0[1]),.dout(n511),.clk(gclk));
	jor g0211(.dina(n511),.dinb(w_dff_B_RjlglxQt3_1),.dout(n512),.clk(gclk));
	jand g0212(.dina(w_G3548_2[0]),.dinb(w_n507_1[0]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3546_2[1]),.dinb(w_G218_2[0]),.dout(n514),.clk(gclk));
	jor g0214(.dina(n514),.dinb(w_G468_1[1]),.dout(n515),.clk(gclk));
	jor g0215(.dina(n515),.dinb(n513),.dout(n516),.clk(gclk));
	jand g0216(.dina(w_dff_B_tG9adEFH1_0),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G206_0[2]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_G251_3[2]),.dinb(w_n518_1[1]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G446_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_G248_4[1]),.dinb(w_G206_0[1]),.dout(n521),.clk(gclk));
	jor g0221(.dina(n521),.dinb(n520),.dout(n522),.clk(gclk));
	jor g0222(.dina(n522),.dinb(n519),.dout(n523),.clk(gclk));
	jand g0223(.dina(w_n366_3[2]),.dinb(w_n518_1[0]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_n368_4[1]),.dinb(w_G206_0[0]),.dout(n525),.clk(gclk));
	jor g0225(.dina(n525),.dinb(w_G446_1[1]),.dout(n526),.clk(gclk));
	jor g0226(.dina(n526),.dinb(w_dff_B_Vte1rW7f8_1),.dout(n527),.clk(gclk));
	jand g0227(.dina(n527),.dinb(w_dff_B_mmaQjxYO6_1),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[2]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G226_2[2]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n386_1[2]),.dinb(w_n530_1[1]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G422_2[1]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n389_1[2]),.dinb(w_G226_2[1]),.dout(n533),.clk(gclk));
	jor g0233(.dina(n533),.dinb(w_n532_0[1]),.dout(n534),.clk(gclk));
	jor g0234(.dina(n534),.dinb(w_dff_B_dYPgXtsD0_1),.dout(n535),.clk(gclk));
	jand g0235(.dina(w_G3548_1[2]),.dinb(w_n530_1[0]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3546_2[0]),.dinb(w_G226_2[0]),.dout(n537),.clk(gclk));
	jor g0237(.dina(n537),.dinb(w_G422_2[0]),.dout(n538),.clk(gclk));
	jor g0238(.dina(n538),.dinb(n536),.dout(n539),.clk(gclk));
	jand g0239(.dina(w_dff_B_bXdLyk5W1_0),.dinb(n535),.dout(n540),.clk(gclk));
	jnot g0240(.din(w_G210_2[2]),.dout(n541),.clk(gclk));
	jand g0241(.dina(w_n386_1[1]),.dinb(w_n541_1[1]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G457_2[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_n389_1[1]),.dinb(w_G210_2[1]),.dout(n544),.clk(gclk));
	jor g0244(.dina(n544),.dinb(w_n543_0[1]),.dout(n545),.clk(gclk));
	jor g0245(.dina(n545),.dinb(w_dff_B_XX2WTl2R5_1),.dout(n546),.clk(gclk));
	jand g0246(.dina(w_G3548_1[1]),.dinb(w_n541_1[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_G3546_1[2]),.dinb(w_G210_2[0]),.dout(n548),.clk(gclk));
	jor g0248(.dina(n548),.dinb(w_G457_2[0]),.dout(n549),.clk(gclk));
	jor g0249(.dina(n549),.dinb(n547),.dout(n550),.clk(gclk));
	jand g0250(.dina(w_dff_B_zfgiQdEd9_0),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[1]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(w_dff_B_fBBsNrfa9_1),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_dff_B_rTBel3Ui5_1),.dout(w_dff_A_JI54GYgt8_2),.clk(gclk));
	jnot g0255(.din(w_G335_4[1]),.dout(n556),.clk(gclk));
	jor g0256(.dina(w_n556_5[1]),.dinb(w_dff_B_XMxOAZNd4_1),.dout(n557),.clk(gclk));
	jand g0257(.dina(w_n556_5[0]),.dinb(w_n460_1[0]),.dout(n558),.clk(gclk));
	jnot g0258(.din(n558),.dout(n559),.clk(gclk));
	jand g0259(.dina(n559),.dinb(w_dff_B_sgRjECoX8_1),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_1[1]),.dinb(w_G435_1[0]),.dout(n561),.clk(gclk));
	jnot g0261(.din(w_n561_0[2]),.dout(n562),.clk(gclk));
	jnot g0262(.din(G288),.dout(n563),.clk(gclk));
	jand g0263(.dina(w_G335_4[0]),.dinb(n563),.dout(n564),.clk(gclk));
	jand g0264(.dina(w_n556_4[2]),.dinb(w_n495_1[0]),.dout(n565),.clk(gclk));
	jor g0265(.dina(n565),.dinb(n564),.dout(n566),.clk(gclk));
	jxor g0266(.dina(w_n566_0[2]),.dinb(w_n497_1[0]),.dout(n567),.clk(gclk));
	jor g0267(.dina(w_n556_4[1]),.dinb(w_G280_0[1]),.dout(n568),.clk(gclk));
	jor g0268(.dina(w_G335_3[2]),.dinb(w_G273_1[2]),.dout(n569),.clk(gclk));
	jand g0269(.dina(w_n569_0[1]),.dinb(n568),.dout(n570),.clk(gclk));
	jxor g0270(.dina(w_n570_0[1]),.dinb(w_n486_1[0]),.dout(n571),.clk(gclk));
	jnot g0271(.din(w_n571_1[1]),.dout(n572),.clk(gclk));
	jand g0272(.dina(w_n572_0[2]),.dinb(w_n567_1[1]),.dout(n573),.clk(gclk));
	jnot g0273(.din(n573),.dout(n574),.clk(gclk));
	jor g0274(.dina(w_n556_4[0]),.dinb(w_dff_B_zXsy4sDE9_1),.dout(n575),.clk(gclk));
	jor g0275(.dina(w_G335_3[1]),.dinb(w_G257_1[2]),.dout(n576),.clk(gclk));
	jand g0276(.dina(w_dff_B_SyGdP9t01_0),.dinb(n575),.dout(n577),.clk(gclk));
	jxor g0277(.dina(w_n577_0[2]),.dinb(w_n473_1[1]),.dout(n578),.clk(gclk));
	jnot g0278(.din(G272),.dout(n579),.clk(gclk));
	jand g0279(.dina(w_G335_3[0]),.dinb(n579),.dout(n580),.clk(gclk));
	jand g0280(.dina(w_n556_3[2]),.dinb(w_n449_1[0]),.dout(n581),.clk(gclk));
	jor g0281(.dina(n581),.dinb(n580),.dout(n582),.clk(gclk));
	jxor g0282(.dina(w_n582_1[1]),.dinb(w_G400_0[2]),.dout(n583),.clk(gclk));
	jor g0283(.dina(w_n583_1[1]),.dinb(w_n578_0[2]),.dout(n584),.clk(gclk));
	jor g0284(.dina(w_dff_B_zyEKpJaB5_0),.dinb(w_n574_0[2]),.dout(n585),.clk(gclk));
	jor g0285(.dina(w_n585_0[1]),.dinb(w_n562_0[1]),.dout(n586),.clk(gclk));
	jnot g0286(.din(n586),.dout(n587),.clk(gclk));
	jor g0287(.dina(w_n556_3[1]),.dinb(w_dff_B_gwnaqesO9_1),.dout(n588),.clk(gclk));
	jor g0288(.dina(w_G335_2[2]),.dinb(w_G210_1[2]),.dout(n589),.clk(gclk));
	jand g0289(.dina(w_dff_B_jK6rhq0e3_0),.dinb(n588),.dout(n590),.clk(gclk));
	jxor g0290(.dina(w_n590_1[1]),.dinb(w_G457_1[2]),.dout(n591),.clk(gclk));
	jor g0291(.dina(w_n556_3[0]),.dinb(w_dff_B_eO5eMZRj6_1),.dout(n592),.clk(gclk));
	jand g0292(.dina(w_n556_2[2]),.dinb(w_n518_0[2]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jand g0294(.dina(n594),.dinb(w_dff_B_EBnxoP7t6_1),.dout(n595),.clk(gclk));
	jxor g0295(.dina(w_n595_1[1]),.dinb(w_G446_1[0]),.dout(n596),.clk(gclk));
	jand g0296(.dina(w_n596_0[2]),.dinb(w_n591_0[1]),.dout(n597),.clk(gclk));
	jor g0297(.dina(w_n556_2[1]),.dinb(w_dff_B_RdkYRMhY3_1),.dout(n598),.clk(gclk));
	jor g0298(.dina(w_G335_2[1]),.dinb(w_G226_1[2]),.dout(n599),.clk(gclk));
	jand g0299(.dina(w_dff_B_Gw3mBlYD2_0),.dinb(n598),.dout(n600),.clk(gclk));
	jxor g0300(.dina(w_n600_1[1]),.dinb(w_G422_1[2]),.dout(n601),.clk(gclk));
	jor g0301(.dina(w_n556_2[0]),.dinb(w_dff_B_OGZ3SmVF3_1),.dout(n602),.clk(gclk));
	jor g0302(.dina(w_G335_2[0]),.dinb(w_G218_1[2]),.dout(n603),.clk(gclk));
	jand g0303(.dina(w_dff_B_lJJhKMIC2_0),.dinb(n602),.dout(n604),.clk(gclk));
	jxor g0304(.dina(w_n604_0[2]),.dinb(w_G468_1[0]),.dout(n605),.clk(gclk));
	jand g0305(.dina(w_n605_2[2]),.dinb(w_n601_0[1]),.dout(n606),.clk(gclk));
	jand g0306(.dina(w_dff_B_dI9q9fvR7_0),.dinb(n597),.dout(n607),.clk(gclk));
	jand g0307(.dina(w_n607_0[2]),.dinb(w_n587_1[1]),.dout(w_dff_A_QgbmpZht9_2),.clk(gclk));
	jnot g0308(.din(w_G332_4[2]),.dout(n609),.clk(gclk));
	jor g0309(.dina(w_n609_5[2]),.dinb(w_G331_0[1]),.dout(n610),.clk(gclk));
	jand g0310(.dina(w_n609_5[1]),.dinb(w_n424_1[2]),.dout(n611),.clk(gclk));
	jnot g0311(.din(n611),.dout(n612),.clk(gclk));
	jand g0312(.dina(n612),.dinb(w_dff_B_2GSH3u6a3_1),.dout(n613),.clk(gclk));
	jxor g0313(.dina(w_n613_0[2]),.dinb(w_G503_1[0]),.dout(n614),.clk(gclk));
	jor g0314(.dina(w_G358_0[0]),.dinb(w_n609_5[0]),.dout(n615),.clk(gclk));
	jor g0315(.dina(w_G351_1[2]),.dinb(w_G332_4[1]),.dout(n616),.clk(gclk));
	jand g0316(.dina(w_dff_B_ow5BU3l15_0),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_n388_1[1]),.dout(n618),.clk(gclk));
	jand g0318(.dina(w_G600_0),.dinb(w_G332_4[0]),.dout(n619),.clk(gclk));
	jand g0319(.dina(w_n416_0[0]),.dinb(w_n609_4[2]),.dout(n620),.clk(gclk));
	jor g0320(.dina(n620),.dinb(n619),.dout(n621),.clk(gclk));
	jnot g0321(.din(w_n621_2[1]),.dout(n622),.clk(gclk));
	jor g0322(.dina(w_n622_1[1]),.dinb(w_n618_1[1]),.dout(n623),.clk(gclk));
	jand g0323(.dina(w_G611_0),.dinb(w_G332_3[2]),.dout(n624),.clk(gclk));
	jxor g0324(.dina(w_n624_1[2]),.dinb(w_G514_0[2]),.dout(n625),.clk(gclk));
	jor g0325(.dina(w_G348_0[0]),.dinb(w_n609_4[1]),.dout(n626),.clk(gclk));
	jor g0326(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n627),.clk(gclk));
	jand g0327(.dina(w_dff_B_sRRrq9fT4_0),.dinb(n626),.dout(n628),.clk(gclk));
	jxor g0328(.dina(w_n628_0[2]),.dinb(w_n437_1[1]),.dout(n629),.clk(gclk));
	jor g0329(.dina(w_n629_0[2]),.dinb(w_n625_0[2]),.dout(n630),.clk(gclk));
	jor g0330(.dina(n630),.dinb(w_n623_0[1]),.dout(n631),.clk(gclk));
	jnot g0331(.din(w_n631_0[1]),.dout(n632),.clk(gclk));
	jand g0332(.dina(n632),.dinb(w_n614_2[1]),.dout(n633),.clk(gclk));
	jand g0333(.dina(w_G332_3[0]),.dinb(w_G593_0),.dout(n634),.clk(gclk));
	jand g0334(.dina(w_n609_4[0]),.dinb(w_n398_0[1]),.dout(n635),.clk(gclk));
	jor g0335(.dina(n635),.dinb(n634),.dout(n636),.clk(gclk));
	jor g0336(.dina(w_n609_3[2]),.dinb(w_dff_B_BVkNQ79x1_1),.dout(n637),.clk(gclk));
	jand g0337(.dina(w_n609_3[1]),.dinb(w_n403_0[0]),.dout(n638),.clk(gclk));
	jnot g0338(.din(n638),.dout(n639),.clk(gclk));
	jand g0339(.dina(n639),.dinb(w_dff_B_8Vk4FzSE9_1),.dout(n640),.clk(gclk));
	jnot g0340(.din(w_n640_1[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n641_0[1]),.dinb(w_n636_1[1]),.dout(n642),.clk(gclk));
	jor g0342(.dina(w_n609_3[0]),.dinb(w_dff_B_lFMH0nP49_1),.dout(n643),.clk(gclk));
	jor g0343(.dina(w_G332_2[2]),.dinb(w_G308_0[2]),.dout(n644),.clk(gclk));
	jand g0344(.dina(w_dff_B_aa12GdHb2_0),.dinb(n643),.dout(n645),.clk(gclk));
	jxor g0345(.dina(w_n645_0[2]),.dinb(w_G479_0[2]),.dout(n646),.clk(gclk));
	jor g0346(.dina(w_n609_2[2]),.dinb(w_dff_B_EbanuIL94_1),.dout(n647),.clk(gclk));
	jor g0347(.dina(w_G332_2[1]),.dinb(w_G316_0[2]),.dout(n648),.clk(gclk));
	jand g0348(.dina(w_dff_B_HkACRLua4_0),.dinb(n647),.dout(n649),.clk(gclk));
	jxor g0349(.dina(w_n649_1[1]),.dinb(w_G490_1[0]),.dout(n650),.clk(gclk));
	jand g0350(.dina(w_n650_0[1]),.dinb(w_n646_0[2]),.dout(n651),.clk(gclk));
	jand g0351(.dina(w_n651_1[1]),.dinb(w_n642_0[1]),.dout(n652),.clk(gclk));
	jand g0352(.dina(w_n652_0[1]),.dinb(w_n633_1[1]),.dout(w_dff_A_0OgvtRqK7_2),.clk(gclk));
	jxor g0353(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n654),.clk(gclk));
	jxor g0354(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n655),.clk(gclk));
	jxor g0355(.dina(n655),.dinb(n654),.dout(n656),.clk(gclk));
	jxor g0356(.dina(w_G369_0[1]),.dinb(w_G361_0[0]),.dout(n657),.clk(gclk));
	jxor g0357(.dina(n657),.dinb(w_n424_1[1]),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_G302_0[0]),.dinb(w_n398_0[0]),.dout(n659),.clk(gclk));
	jxor g0359(.dina(n659),.dinb(n658),.dout(n660),.clk(gclk));
	jxor g0360(.dina(n660),.dinb(w_dff_B_omv28N7A3_1),.dout(n661),.clk(gclk));
	jnot g0361(.din(w_n661_0[1]),.dout(w_dff_A_ExzIBIS38_1),.clk(gclk));
	jxor g0362(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G273_1[1]),.dinb(w_G265_1[1]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(n663),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(n667),.dinb(n666),.dout(n668),.clk(gclk));
	jxor g0368(.dina(w_G210_1[1]),.dinb(w_n518_0[1]),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n668),.dout(n670),.clk(gclk));
	jxor g0370(.dina(n670),.dinb(w_dff_B_8xlMiN679_1),.dout(n671),.clk(gclk));
	jnot g0371(.din(w_n671_0[1]),.dout(w_dff_A_eF25cZUD2_1),.clk(gclk));
	jnot g0372(.din(w_n560_1[0]),.dout(n673),.clk(gclk));
	jand g0373(.dina(n673),.dinb(w_n462_0[1]),.dout(n674),.clk(gclk));
	jnot g0374(.din(n674),.dout(n675),.clk(gclk));
	jand g0375(.dina(w_n560_0[2]),.dinb(w_G435_0[2]),.dout(n676),.clk(gclk));
	jnot g0376(.din(w_n577_0[1]),.dout(n677),.clk(gclk));
	jand g0377(.dina(w_n677_0[1]),.dinb(w_n473_1[0]),.dout(n678),.clk(gclk));
	jor g0378(.dina(w_n677_0[0]),.dinb(w_n473_0[2]),.dout(n679),.clk(gclk));
	jand g0379(.dina(w_n582_1[0]),.dinb(w_n451_1[0]),.dout(n680),.clk(gclk));
	jor g0380(.dina(w_n566_0[1]),.dinb(w_n497_0[2]),.dout(n681),.clk(gclk));
	jor g0381(.dina(w_n571_1[0]),.dinb(w_n681_2[1]),.dout(n682),.clk(gclk));
	jnot g0382(.din(w_G280_0[0]),.dout(n683),.clk(gclk));
	jand g0383(.dina(w_G335_1[2]),.dinb(n683),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n569_0[0]),.dout(n685),.clk(gclk));
	jor g0385(.dina(n685),.dinb(n684),.dout(n686),.clk(gclk));
	jor g0386(.dina(n686),.dinb(w_n486_0[2]),.dout(n687),.clk(gclk));
	jor g0387(.dina(w_n582_0[2]),.dinb(w_n451_0[2]),.dout(n688),.clk(gclk));
	jand g0388(.dina(n688),.dinb(w_n687_0[2]),.dout(n689),.clk(gclk));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n682_0[1]),.dout(n690),.clk(gclk));
	jor g0390(.dina(n690),.dinb(w_n680_0[1]),.dout(n691),.clk(gclk));
	jand g0391(.dina(w_n691_0[2]),.dinb(w_n679_0[1]),.dout(n692),.clk(gclk));
	jor g0392(.dina(n692),.dinb(w_n678_0[1]),.dout(n693),.clk(gclk));
	jnot g0393(.din(w_n693_0[2]),.dout(n694),.clk(gclk));
	jor g0394(.dina(n694),.dinb(w_dff_B_Uc3tdeoM0_1),.dout(n695),.clk(gclk));
	jand g0395(.dina(n695),.dinb(w_dff_B_15CS6bYn4_1),.dout(n696),.clk(gclk));
	jand g0396(.dina(w_n696_0[2]),.dinb(w_n607_0[1]),.dout(n697),.clk(gclk));
	jand g0397(.dina(w_n595_1[0]),.dinb(w_G446_0[2]),.dout(n698),.clk(gclk));
	jor g0398(.dina(w_n595_0[2]),.dinb(w_G446_0[1]),.dout(n699),.clk(gclk));
	jor g0399(.dina(w_n590_1[0]),.dinb(w_G457_1[1]),.dout(n700),.clk(gclk));
	jand g0400(.dina(w_n590_0[2]),.dinb(w_G457_1[0]),.dout(n701),.clk(gclk));
	jand g0401(.dina(w_n604_0[1]),.dinb(w_G468_0[2]),.dout(n702),.clk(gclk));
	jand g0402(.dina(w_n600_1[0]),.dinb(w_G422_1[1]),.dout(n703),.clk(gclk));
	jand g0403(.dina(w_n605_2[1]),.dinb(w_n703_0[2]),.dout(n704),.clk(gclk));
	jor g0404(.dina(n704),.dinb(w_n702_0[1]),.dout(n705),.clk(gclk));
	jor g0405(.dina(w_n705_0[1]),.dinb(w_dff_B_QoISKYFR2_1),.dout(n706),.clk(gclk));
	jand g0406(.dina(w_n706_0[1]),.dinb(w_n700_0[1]),.dout(n707),.clk(gclk));
	jand g0407(.dina(w_n707_0[2]),.dinb(w_dff_B_sQ1LnrdP9_1),.dout(n708),.clk(gclk));
	jor g0408(.dina(n708),.dinb(w_dff_B_YYYGQkai2_1),.dout(n709),.clk(gclk));
	jor g0409(.dina(w_n709_0[1]),.dinb(w_n697_0[1]),.dout(w_dff_A_mfoVLXEC9_2),.clk(gclk));
	jand g0410(.dina(w_n613_0[1]),.dinb(w_G503_0[2]),.dout(n711),.clk(gclk));
	jor g0411(.dina(w_n624_1[1]),.dinb(w_n410_1[0]),.dout(n712),.clk(gclk));
	jand g0412(.dina(w_n624_1[0]),.dinb(w_n410_0[2]),.dout(n713),.clk(gclk));
	jand g0413(.dina(w_G599_0),.dinb(w_G332_2[0]),.dout(n714),.clk(gclk));
	jand g0414(.dina(w_n435_1[0]),.dinb(w_n609_2[1]),.dout(n715),.clk(gclk));
	jor g0415(.dina(n715),.dinb(n714),.dout(n716),.clk(gclk));
	jand g0416(.dina(w_n716_0[1]),.dinb(w_n437_1[0]),.dout(n717),.clk(gclk));
	jand g0417(.dina(w_G612_0),.dinb(w_G332_1[2]),.dout(n718),.clk(gclk));
	jand g0418(.dina(w_n385_1[0]),.dinb(w_n609_2[0]),.dout(n719),.clk(gclk));
	jor g0419(.dina(n719),.dinb(n718),.dout(n720),.clk(gclk));
	jand g0420(.dina(w_n720_0[1]),.dinb(w_n388_1[0]),.dout(n721),.clk(gclk));
	jor g0421(.dina(w_n621_2[0]),.dinb(w_n721_0[2]),.dout(n722),.clk(gclk));
	jor g0422(.dina(w_n720_0[0]),.dinb(w_n388_0[2]),.dout(n723),.clk(gclk));
	jor g0423(.dina(w_n716_0[0]),.dinb(w_n437_0[2]),.dout(n724),.clk(gclk));
	jand g0424(.dina(n724),.dinb(w_n723_0[1]),.dout(n725),.clk(gclk));
	jand g0425(.dina(n725),.dinb(n722),.dout(n726),.clk(gclk));
	jor g0426(.dina(w_n726_0[1]),.dinb(w_n717_0[2]),.dout(n727),.clk(gclk));
	jor g0427(.dina(w_n727_0[2]),.dinb(w_dff_B_xTDbuQrc6_1),.dout(n728),.clk(gclk));
	jand g0428(.dina(n728),.dinb(w_dff_B_B3RK3ujN2_1),.dout(n729),.clk(gclk));
	jnot g0429(.din(w_n729_1[1]),.dout(n730),.clk(gclk));
	jand g0430(.dina(n730),.dinb(w_n614_2[0]),.dout(n731),.clk(gclk));
	jor g0431(.dina(n731),.dinb(w_dff_B_qOGmSgWp9_1),.dout(n732),.clk(gclk));
	jand g0432(.dina(w_n732_0[2]),.dinb(w_n651_1[0]),.dout(n733),.clk(gclk));
	jnot g0433(.din(w_n642_0[0]),.dout(n734),.clk(gclk));
	jnot g0434(.din(w_n645_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[1]),.dinb(w_n362_0[0]),.dout(n736),.clk(gclk));
	jnot g0436(.din(w_n736_0[1]),.dout(n737),.clk(gclk));
	jand g0437(.dina(w_n645_0[0]),.dinb(w_G479_0[1]),.dout(n738),.clk(gclk));
	jand g0438(.dina(w_n649_1[0]),.dinb(w_G490_0[2]),.dout(n739),.clk(gclk));
	jor g0439(.dina(w_n739_1[1]),.dinb(n738),.dout(n740),.clk(gclk));
	jand g0440(.dina(w_n740_0[1]),.dinb(n737),.dout(n741),.clk(gclk));
	jor g0441(.dina(w_n741_0[1]),.dinb(n734),.dout(n742),.clk(gclk));
	jor g0442(.dina(w_n742_0[1]),.dinb(w_n733_0[1]),.dout(w_dff_A_qJmjJP2c4_2),.clk(gclk));
	jnot g0443(.din(w_G54_0[1]),.dout(n744),.clk(gclk));
	jxor g0444(.dina(w_n621_1[2]),.dinb(w_n744_1[2]),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_G4092_1[2]),.dout(n746),.clk(gclk));
	jand g0446(.dina(w_n746_1[2]),.dinb(w_G4091_2[2]),.dout(n747),.clk(gclk));
	jnot g0447(.din(w_n747_3[2]),.dout(n748),.clk(gclk));
	jor g0448(.dina(w_n748_4[1]),.dinb(n745),.dout(n749),.clk(gclk));
	jnot g0449(.din(w_G4091_2[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n746_1[1]),.dinb(w_n750_1[1]),.dout(n751),.clk(gclk));
	jand g0451(.dina(w_n751_2[1]),.dinb(w_n419_0[1]),.dout(n752),.clk(gclk));
	jand g0452(.dina(w_G4092_1[1]),.dinb(w_n750_1[0]),.dout(n753),.clk(gclk));
	jand g0453(.dina(w_n753_8[1]),.dinb(w_dff_B_EU7b06o62_1),.dout(n754),.clk(gclk));
	jor g0454(.dina(w_dff_B_9ZXX0n5X8_0),.dinb(n752),.dout(n755),.clk(gclk));
	jnot g0455(.din(n755),.dout(n756),.clk(gclk));
	jand g0456(.dina(n756),.dinb(w_dff_B_chrVOFeU6_1),.dout(G822_fa_),.clk(gclk));
	jnot g0457(.din(w_n618_1[0]),.dout(n758),.clk(gclk));
	jand g0458(.dina(w_n621_1[1]),.dinb(w_n744_1[1]),.dout(n759),.clk(gclk));
	jnot g0459(.din(w_n759_0[1]),.dout(n760),.clk(gclk));
	jand g0460(.dina(w_n760_0[1]),.dinb(n758),.dout(n761),.clk(gclk));
	jand g0461(.dina(w_n759_0[0]),.dinb(w_n618_0[2]),.dout(n762),.clk(gclk));
	jor g0462(.dina(n762),.dinb(w_n748_4[0]),.dout(n763),.clk(gclk));
	jor g0463(.dina(n763),.dinb(w_n761_0[1]),.dout(n764),.clk(gclk));
	jnot g0464(.din(w_n751_2[0]),.dout(n765),.clk(gclk));
	jor g0465(.dina(w_n765_5[2]),.dinb(w_n397_0[0]),.dout(n766),.clk(gclk));
	jand g0466(.dina(w_n753_8[0]),.dinb(w_dff_B_H453Fxi78_1),.dout(n767),.clk(gclk));
	jnot g0467(.din(n767),.dout(n768),.clk(gclk));
	jand g0468(.dina(w_dff_B_RNq2kfq04_0),.dinb(n766),.dout(n769),.clk(gclk));
	jand g0469(.dina(n769),.dinb(n764),.dout(G838_fa_),.clk(gclk));
	jxor g0470(.dina(w_n567_1[0]),.dinb(w_G4_1[1]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n771_0[1]),.dinb(w_n747_3[1]),.dout(n772),.clk(gclk));
	jnot g0472(.din(n772),.dout(n773),.clk(gclk));
	jor g0473(.dina(w_n765_5[1]),.dinb(w_n505_0[0]),.dout(n774),.clk(gclk));
	jand g0474(.dina(w_n753_7[2]),.dinb(w_dff_B_ippiVCQk1_1),.dout(n775),.clk(gclk));
	jnot g0475(.din(n775),.dout(n776),.clk(gclk));
	jand g0476(.dina(w_dff_B_9X5TAAfm0_0),.dinb(n774),.dout(n777),.clk(gclk));
	jand g0477(.dina(n777),.dinb(n773),.dout(G861_fa_),.clk(gclk));
	jnot g0478(.din(w_n636_1[0]),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n633_1[0]),.dinb(w_G54_0[0]),.dout(n780),.clk(gclk));
	jor g0480(.dina(w_dff_B_5Ubx6wng4_0),.dinb(w_n732_0[1]),.dout(n781),.clk(gclk));
	jand g0481(.dina(w_n781_0[2]),.dinb(w_n651_0[2]),.dout(n782),.clk(gclk));
	jor g0482(.dina(n782),.dinb(w_n741_0[0]),.dout(n783),.clk(gclk));
	jnot g0483(.din(w_n783_1[1]),.dout(n784),.clk(gclk));
	jor g0484(.dina(n784),.dinb(w_n779_0[1]),.dout(n785),.clk(gclk));
	jxor g0485(.dina(w_n640_1[1]),.dinb(w_n779_0[0]),.dout(n786),.clk(gclk));
	jnot g0486(.din(w_n786_0[1]),.dout(n787),.clk(gclk));
	jor g0487(.dina(w_n787_0[1]),.dinb(w_n783_1[0]),.dout(n788),.clk(gclk));
	jand g0488(.dina(w_dff_B_9gUly01L6_0),.dinb(n785),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n789_0[2]),.dout(w_dff_A_k5yPLMrJ3_1),.clk(gclk));
	jnot g0490(.din(w_G861_0),.dout(n791),.clk(gclk));
	jnot g0491(.din(w_G4087_0[2]),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_G4088_0[2]),.dinb(w_n792_0[1]),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n793_4[1]),.dinb(w_n791_1[1]),.dout(n794),.clk(gclk));
	jnot g0494(.din(w_G822_0),.dout(n795),.clk(gclk));
	jnot g0495(.din(w_G4088_0[1]),.dout(n796),.clk(gclk));
	jand g0496(.dina(w_n796_0[1]),.dinb(w_n792_0[0]),.dout(n797),.clk(gclk));
	jand g0497(.dina(w_n797_4[1]),.dinb(w_n795_1[1]),.dout(n798),.clk(gclk));
	jand g0498(.dina(w_n796_0[0]),.dinb(w_G4087_0[1]),.dout(n799),.clk(gclk));
	jand g0499(.dina(w_n799_4[1]),.dinb(w_G11_0[1]),.dout(n800),.clk(gclk));
	jand g0500(.dina(w_G4088_0[0]),.dinb(w_G4087_0[0]),.dout(n801),.clk(gclk));
	jand g0501(.dina(w_n801_4[1]),.dinb(w_G61_0[1]),.dout(n802),.clk(gclk));
	jor g0502(.dina(w_dff_B_hOLlBpdr3_0),.dinb(n800),.dout(n803),.clk(gclk));
	jor g0503(.dina(w_dff_B_mmIR7lIl0_0),.dinb(n798),.dout(n804),.clk(gclk));
	jor g0504(.dina(n804),.dinb(n794),.dout(w_dff_A_GvPDbonV7_2),.clk(gclk));
	jand g0505(.dina(w_n729_1[0]),.dinb(w_n631_0[0]),.dout(n806),.clk(gclk));
	jand g0506(.dina(w_n729_0[2]),.dinb(w_n744_1[0]),.dout(n807),.clk(gclk));
	jor g0507(.dina(n807),.dinb(w_n806_0[2]),.dout(n808),.clk(gclk));
	jxor g0508(.dina(n808),.dinb(w_n614_1[2]),.dout(n809),.clk(gclk));
	jor g0509(.dina(w_n809_0[1]),.dinb(w_n748_3[2]),.dout(n810),.clk(gclk));
	jor g0510(.dina(w_n765_5[0]),.dinb(w_n434_0[0]),.dout(n811),.clk(gclk));
	jand g0511(.dina(w_n753_7[1]),.dinb(w_dff_B_QJjsEbXt0_1),.dout(n812),.clk(gclk));
	jnot g0512(.din(n812),.dout(n813),.clk(gclk));
	jand g0513(.dina(w_dff_B_r8g0D6iJ3_0),.dinb(n811),.dout(n814),.clk(gclk));
	jand g0514(.dina(w_dff_B_TAKE6U3t4_0),.dinb(n810),.dout(G832_fa_),.clk(gclk));
	jnot g0515(.din(w_n625_0[1]),.dout(n816),.clk(gclk));
	jand g0516(.dina(w_n727_0[1]),.dinb(w_n744_0[2]),.dout(n817),.clk(gclk));
	jand g0517(.dina(w_n726_0[0]),.dinb(w_n623_0[0]),.dout(n818),.clk(gclk));
	jor g0518(.dina(n818),.dinb(w_n717_0[1]),.dout(n819),.clk(gclk));
	jor g0519(.dina(w_n819_0[1]),.dinb(n817),.dout(n820),.clk(gclk));
	jxor g0520(.dina(n820),.dinb(w_dff_B_FMUbEqxb4_1),.dout(n821),.clk(gclk));
	jor g0521(.dina(w_n821_0[1]),.dinb(w_n748_3[1]),.dout(n822),.clk(gclk));
	jand g0522(.dina(w_n751_1[2]),.dinb(w_n414_0[0]),.dout(n823),.clk(gclk));
	jand g0523(.dina(w_n753_7[0]),.dinb(w_dff_B_lNEbkQDY3_1),.dout(n824),.clk(gclk));
	jor g0524(.dina(w_dff_B_pWZ8gdsS9_0),.dinb(n823),.dout(n825),.clk(gclk));
	jnot g0525(.din(n825),.dout(n826),.clk(gclk));
	jand g0526(.dina(w_dff_B_q7sIJVml5_0),.dinb(n822),.dout(G834_fa_),.clk(gclk));
	jor g0527(.dina(w_n617_1[0]),.dinb(w_G534_1[0]),.dout(n828),.clk(gclk));
	jand g0528(.dina(w_n617_0[2]),.dinb(w_G534_0[2]),.dout(n829),.clk(gclk));
	jor g0529(.dina(w_n760_0[0]),.dinb(w_n829_0[1]),.dout(n830),.clk(gclk));
	jand g0530(.dina(n830),.dinb(w_n828_0[2]),.dout(n831),.clk(gclk));
	jxor g0531(.dina(n831),.dinb(w_n629_0[1]),.dout(n832),.clk(gclk));
	jor g0532(.dina(w_n832_0[1]),.dinb(w_n748_3[0]),.dout(n833),.clk(gclk));
	jor g0533(.dina(w_n765_4[2]),.dinb(w_n445_0[0]),.dout(n834),.clk(gclk));
	jand g0534(.dina(w_n753_6[2]),.dinb(w_dff_B_iojmpH570_1),.dout(n835),.clk(gclk));
	jnot g0535(.din(n835),.dout(n836),.clk(gclk));
	jand g0536(.dina(w_dff_B_hQgBgHlP8_0),.dinb(n834),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_dff_B_9lmp3lFb5_0),.dinb(n833),.dout(G836_fa_),.clk(gclk));
	jnot g0538(.din(w_G4090_0[2]),.dout(n839),.clk(gclk));
	jand g0539(.dina(w_n839_0[1]),.dinb(w_G4089_0[2]),.dout(n840),.clk(gclk));
	jand g0540(.dina(w_n840_4[1]),.dinb(w_n791_1[0]),.dout(n841),.clk(gclk));
	jnot g0541(.din(w_G4089_0[1]),.dout(n842),.clk(gclk));
	jand g0542(.dina(w_n839_0[0]),.dinb(w_n842_0[1]),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n843_4[1]),.dinb(w_n795_1[0]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_G4090_0[1]),.dinb(w_n842_0[0]),.dout(n845),.clk(gclk));
	jand g0545(.dina(w_n845_4[1]),.dinb(w_G11_0[0]),.dout(n846),.clk(gclk));
	jand g0546(.dina(w_G4090_0[0]),.dinb(w_G4089_0[0]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_4[1]),.dinb(w_G61_0[0]),.dout(n848),.clk(gclk));
	jor g0548(.dina(w_dff_B_tx0jMe6i2_0),.dinb(n846),.dout(n849),.clk(gclk));
	jor g0549(.dina(w_dff_B_xNysK2R40_0),.dinb(n844),.dout(n850),.clk(gclk));
	jor g0550(.dina(n850),.dinb(n841),.dout(w_dff_A_8TrmV4bo1_2),.clk(gclk));
	jnot g0551(.din(w_n678_0[0]),.dout(n852),.clk(gclk));
	jnot g0552(.din(w_n679_0[0]),.dout(n853),.clk(gclk));
	jor g0553(.dina(w_n583_1[0]),.dinb(w_n574_0[1]),.dout(n854),.clk(gclk));
	jand g0554(.dina(n854),.dinb(w_n691_0[1]),.dout(n855),.clk(gclk));
	jnot g0555(.din(w_n855_0[1]),.dout(n856),.clk(gclk));
	jnot g0556(.din(w_n691_0[0]),.dout(n857),.clk(gclk));
	jor g0557(.dina(w_n857_0[1]),.dinb(w_G4_1[0]),.dout(n858),.clk(gclk));
	jand g0558(.dina(w_dff_B_utGnKuzG6_0),.dinb(w_n856_0[1]),.dout(n859),.clk(gclk));
	jor g0559(.dina(w_n859_0[1]),.dinb(w_n853_0[1]),.dout(n860),.clk(gclk));
	jand g0560(.dina(n860),.dinb(w_dff_B_EHwVUm3b2_1),.dout(n861),.clk(gclk));
	jxor g0561(.dina(n861),.dinb(w_n562_0[0]),.dout(n862),.clk(gclk));
	jor g0562(.dina(w_n862_0[1]),.dinb(w_n748_2[2]),.dout(n863),.clk(gclk));
	jor g0563(.dina(w_n765_4[1]),.dinb(w_n470_0[0]),.dout(n864),.clk(gclk));
	jand g0564(.dina(w_n753_6[1]),.dinb(w_dff_B_25LjbvG77_1),.dout(n865),.clk(gclk));
	jnot g0565(.din(n865),.dout(n866),.clk(gclk));
	jand g0566(.dina(w_dff_B_eQYXXswa6_0),.dinb(n864),.dout(n867),.clk(gclk));
	jand g0567(.dina(w_dff_B_MjeizViB9_0),.dinb(n863),.dout(G871_fa_),.clk(gclk));
	jxor g0568(.dina(w_n859_0[0]),.dinb(w_n578_0[1]),.dout(n869),.clk(gclk));
	jor g0569(.dina(w_n869_0[1]),.dinb(w_n748_2[1]),.dout(n870),.clk(gclk));
	jor g0570(.dina(w_n765_4[0]),.dinb(w_n481_0[0]),.dout(n871),.clk(gclk));
	jand g0571(.dina(w_n753_6[0]),.dinb(w_dff_B_AiJ3oHxw6_1),.dout(n872),.clk(gclk));
	jnot g0572(.din(n872),.dout(n873),.clk(gclk));
	jand g0573(.dina(w_dff_B_7ZmmlJlu8_0),.dinb(n871),.dout(n874),.clk(gclk));
	jand g0574(.dina(w_dff_B_zG0fkk6t3_0),.dinb(n870),.dout(G873_fa_),.clk(gclk));
	jand g0575(.dina(w_n567_0[2]),.dinb(w_G4_0[2]),.dout(n876),.clk(gclk));
	jnot g0576(.din(n876),.dout(n877),.clk(gclk));
	jand g0577(.dina(w_n877_0[1]),.dinb(w_n681_2[0]),.dout(n878),.clk(gclk));
	jor g0578(.dina(n878),.dinb(w_n571_0[2]),.dout(n879),.clk(gclk));
	jand g0579(.dina(w_n879_0[1]),.dinb(w_n687_0[1]),.dout(n880),.clk(gclk));
	jxor g0580(.dina(n880),.dinb(w_n583_0[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n881_0[1]),.dinb(w_n747_3[0]),.dout(n882),.clk(gclk));
	jnot g0582(.din(n882),.dout(n883),.clk(gclk));
	jor g0583(.dina(w_n765_3[2]),.dinb(w_n459_0[0]),.dout(n884),.clk(gclk));
	jand g0584(.dina(w_n753_5[2]),.dinb(w_dff_B_AIEF4ijs8_1),.dout(n885),.clk(gclk));
	jnot g0585(.din(n885),.dout(n886),.clk(gclk));
	jand g0586(.dina(w_dff_B_RSx2wWa70_0),.dinb(n884),.dout(n887),.clk(gclk));
	jand g0587(.dina(w_dff_B_U4YzXz4t6_0),.dinb(n883),.dout(G875_fa_),.clk(gclk));
	jand g0588(.dina(w_n571_0[1]),.dinb(w_n681_1[2]),.dout(n889),.clk(gclk));
	jand g0589(.dina(w_dff_B_FMmGyVGz9_0),.dinb(w_n877_0[0]),.dout(n890),.clk(gclk));
	jnot g0590(.din(n890),.dout(n891),.clk(gclk));
	jand g0591(.dina(n891),.dinb(w_n879_0[0]),.dout(n892),.clk(gclk));
	jand g0592(.dina(w_n892_0[1]),.dinb(w_n747_2[2]),.dout(n893),.clk(gclk));
	jnot g0593(.din(n893),.dout(n894),.clk(gclk));
	jor g0594(.dina(w_n765_3[1]),.dinb(w_n494_0[0]),.dout(n895),.clk(gclk));
	jand g0595(.dina(w_n753_5[1]),.dinb(w_dff_B_Dq5WLR2J7_1),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jand g0597(.dina(w_dff_B_p60ZL6903_0),.dinb(n895),.dout(n898),.clk(gclk));
	jand g0598(.dina(w_dff_B_sEKMPOcX8_0),.dinb(n894),.dout(G877_fa_),.clk(gclk));
	jxor g0599(.dina(w_n649_0[2]),.dinb(w_n735_0[0]),.dout(n900),.clk(gclk));
	jxor g0600(.dina(n900),.dinb(w_n786_0[0]),.dout(n901),.clk(gclk));
	jxor g0601(.dina(n901),.dinb(w_n621_1[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_G369_0[0]),.dinb(w_n609_1[2]),.dout(n903),.clk(gclk));
	jand g0603(.dina(G372),.dinb(w_G332_1[1]),.dout(n904),.clk(gclk));
	jor g0604(.dina(w_dff_B_bNOwwZgX8_0),.dinb(n903),.dout(n905),.clk(gclk));
	jxor g0605(.dina(n905),.dinb(w_n617_0[1]),.dout(n906),.clk(gclk));
	jxor g0606(.dina(n906),.dinb(w_n628_0[1]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_G331_0[0]),.dout(n908),.clk(gclk));
	jand g0608(.dina(w_n624_0[2]),.dinb(w_dff_B_zdUxXCoH5_1),.dout(n909),.clk(gclk));
	jnot g0609(.din(w_n624_0[1]),.dout(n910),.clk(gclk));
	jand g0610(.dina(w_dff_B_0kxmv4TN6_0),.dinb(w_n613_0[0]),.dout(n911),.clk(gclk));
	jor g0611(.dina(n911),.dinb(w_dff_B_Wzx6zhX68_1),.dout(n912),.clk(gclk));
	jxor g0612(.dina(n912),.dinb(w_dff_B_UImnMwAf3_1),.dout(n913),.clk(gclk));
	jxor g0613(.dina(n913),.dinb(n902),.dout(n914),.clk(gclk));
	jnot g0614(.din(w_n914_0[1]),.dout(w_dff_A_hy3XRMt16_1),.clk(gclk));
	jxor g0615(.dina(w_n577_0[0]),.dinb(w_n566_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n582_0[1]),.dinb(w_n570_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(n917),.dinb(n916),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_n590_0[1]),.dout(n919),.clk(gclk));
	jand g0619(.dina(w_n556_1[2]),.dinb(w_G289_0[0]),.dout(n920),.clk(gclk));
	jand g0620(.dina(w_G335_1[1]),.dinb(G292),.dout(n921),.clk(gclk));
	jor g0621(.dina(w_dff_B_Njv8LDIf3_0),.dinb(n920),.dout(n922),.clk(gclk));
	jxor g0622(.dina(n922),.dinb(w_n600_0[2]),.dout(n923),.clk(gclk));
	jxor g0623(.dina(n923),.dinb(w_n560_0[1]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n604_0[0]),.dinb(w_n595_0[1]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jxor g0626(.dina(n926),.dinb(n919),.dout(G1000_fa_),.clk(gclk));
	jnot g0627(.din(w_n596_0[1]),.dout(n928),.clk(gclk));
	jnot g0628(.din(w_n707_0[1]),.dout(n929),.clk(gclk));
	jnot g0629(.din(w_n700_0[0]),.dout(n930),.clk(gclk));
	jnot g0630(.din(w_n605_2[0]),.dout(n931),.clk(gclk));
	jnot g0631(.din(w_n601_0[0]),.dout(n932),.clk(gclk));
	jnot g0632(.din(w_n696_0[1]),.dout(n933),.clk(gclk));
	jand g0633(.dina(w_n587_1[0]),.dinb(w_G4_0[1]),.dout(n934),.clk(gclk));
	jnot g0634(.din(n934),.dout(n935),.clk(gclk));
	jand g0635(.dina(w_dff_B_bdh2mSot5_0),.dinb(n933),.dout(n936),.clk(gclk));
	jor g0636(.dina(w_n936_0[2]),.dinb(w_n932_0[1]),.dout(n937),.clk(gclk));
	jor g0637(.dina(n937),.dinb(w_dff_B_6DbqdCFJ1_1),.dout(n938),.clk(gclk));
	jor g0638(.dina(w_n938_0[1]),.dinb(w_n930_0[2]),.dout(n939),.clk(gclk));
	jand g0639(.dina(n939),.dinb(w_dff_B_SaJAM3N00_1),.dout(n940),.clk(gclk));
	jxor g0640(.dina(n940),.dinb(w_n928_0[1]),.dout(n941),.clk(gclk));
	jnot g0641(.din(w_n941_0[1]),.dout(n942),.clk(gclk));
	jnot g0642(.din(w_n591_0[0]),.dout(n943),.clk(gclk));
	jnot g0643(.din(w_n705_0[0]),.dout(n944),.clk(gclk));
	jand g0644(.dina(w_n938_0[0]),.dinb(w_n944_0[1]),.dout(n945),.clk(gclk));
	jxor g0645(.dina(n945),.dinb(w_n943_0[1]),.dout(n946),.clk(gclk));
	jnot g0646(.din(w_n946_0[1]),.dout(n947),.clk(gclk));
	jor g0647(.dina(w_n600_0[1]),.dinb(w_G422_1[0]),.dout(n948),.clk(gclk));
	jnot g0648(.din(w_n948_0[2]),.dout(n949),.clk(gclk));
	jnot g0649(.din(w_n703_0[1]),.dout(n950),.clk(gclk));
	jand g0650(.dina(w_n936_0[1]),.dinb(w_dff_B_rRMNoTYZ7_1),.dout(n951),.clk(gclk));
	jor g0651(.dina(n951),.dinb(w_dff_B_gn54M3Ww9_1),.dout(n952),.clk(gclk));
	jxor g0652(.dina(n952),.dinb(w_n605_1[2]),.dout(n953),.clk(gclk));
	jxor g0653(.dina(w_n936_0[0]),.dinb(w_n932_0[0]),.dout(n954),.clk(gclk));
	jnot g0654(.din(w_n954_0[1]),.dout(n955),.clk(gclk));
	jnot g0655(.din(w_n881_0[0]),.dout(n956),.clk(gclk));
	jnot g0656(.din(w_n771_0[0]),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n892_0[0]),.dout(n958),.clk(gclk));
	jand g0658(.dina(n958),.dinb(w_dff_B_0C521gtF5_1),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(n956),.dout(n960),.clk(gclk));
	jand g0660(.dina(n960),.dinb(w_n869_0[0]),.dout(n961),.clk(gclk));
	jand g0661(.dina(w_dff_B_TcczeA249_0),.dinb(w_n862_0[0]),.dout(n962),.clk(gclk));
	jand g0662(.dina(w_dff_B_5yVzVK379_0),.dinb(n955),.dout(n963),.clk(gclk));
	jand g0663(.dina(n963),.dinb(w_n953_0[1]),.dout(n964),.clk(gclk));
	jand g0664(.dina(w_dff_B_bkgjFZb24_0),.dinb(n947),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(n942),.dout(w_dff_A_rzj3Gxf21_2),.clk(gclk));
	jnot g0666(.din(w_n646_0[1]),.dout(n967),.clk(gclk));
	jor g0667(.dina(w_n649_0[1]),.dinb(w_G490_0[1]),.dout(n968),.clk(gclk));
	jor g0668(.dina(w_n781_0[1]),.dinb(w_n739_1[0]),.dout(n969),.clk(gclk));
	jand g0669(.dina(n969),.dinb(w_n968_0[1]),.dout(n970),.clk(gclk));
	jxor g0670(.dina(n970),.dinb(w_dff_B_gZZxHR9A9_1),.dout(n971),.clk(gclk));
	jxor g0671(.dina(w_n783_0[2]),.dinb(w_n640_1[0]),.dout(n972),.clk(gclk));
	jxor g0672(.dina(w_n781_0[0]),.dinb(w_n650_0[0]),.dout(n973),.clk(gclk));
	jnot g0673(.din(w_n973_0[1]),.dout(n974),.clk(gclk));
	jor g0674(.dina(w_n621_0[2]),.dinb(w_n744_0[1]),.dout(n975),.clk(gclk));
	jand g0675(.dina(n975),.dinb(w_n636_0[2]),.dout(n976),.clk(gclk));
	jand g0676(.dina(w_dff_B_i6oJGg1L9_0),.dinb(w_n761_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(w_dff_B_0G1dH7Rk3_0),.dinb(w_n832_0[0]),.dout(n978),.clk(gclk));
	jand g0678(.dina(w_dff_B_ksLsfQMS2_0),.dinb(w_n821_0[0]),.dout(n979),.clk(gclk));
	jand g0679(.dina(w_dff_B_vcqIHBmT2_0),.dinb(w_n809_0[0]),.dout(n980),.clk(gclk));
	jand g0680(.dina(w_dff_B_tWjqZr2a1_0),.dinb(n974),.dout(n981),.clk(gclk));
	jand g0681(.dina(n981),.dinb(w_n972_0[1]),.dout(n982),.clk(gclk));
	jand g0682(.dina(n982),.dinb(w_n971_0[1]),.dout(w_dff_A_OurWUoh22_2),.clk(gclk));
	jnot g0683(.din(w_G1690_0[2]),.dout(n984),.clk(gclk));
	jand g0684(.dina(w_n984_0[1]),.dinb(w_G1689_0[2]),.dout(n985),.clk(gclk));
	jand g0685(.dina(w_n985_4[1]),.dinb(w_n791_0[2]),.dout(n986),.clk(gclk));
	jnot g0686(.din(w_G1689_0[1]),.dout(n987),.clk(gclk));
	jand g0687(.dina(w_n984_0[0]),.dinb(w_n987_0[1]),.dout(n988),.clk(gclk));
	jand g0688(.dina(w_n988_4[1]),.dinb(w_n795_0[2]),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_G1690_0[1]),.dinb(w_n987_0[0]),.dout(n990),.clk(gclk));
	jand g0690(.dina(w_n990_4[1]),.dinb(w_G182_0[1]),.dout(n991),.clk(gclk));
	jand g0691(.dina(w_G1690_0[0]),.dinb(w_G1689_0[0]),.dout(n992),.clk(gclk));
	jand g0692(.dina(w_n992_4[1]),.dinb(w_G185_0[1]),.dout(n993),.clk(gclk));
	jor g0693(.dina(w_dff_B_THwIgXnc9_0),.dinb(n991),.dout(n994),.clk(gclk));
	jor g0694(.dina(w_dff_B_Dp2fIXZN1_0),.dinb(n989),.dout(n995),.clk(gclk));
	jor g0695(.dina(n995),.dinb(n986),.dout(n996),.clk(gclk));
	jand g0696(.dina(n996),.dinb(w_G137_9[1]),.dout(w_dff_A_CdLv686k3_2),.clk(gclk));
	jnot g0697(.din(w_G1694_0[2]),.dout(n998),.clk(gclk));
	jand g0698(.dina(w_n998_0[1]),.dinb(w_G1691_0[2]),.dout(n999),.clk(gclk));
	jand g0699(.dina(w_n999_4[1]),.dinb(w_n791_0[1]),.dout(n1000),.clk(gclk));
	jnot g0700(.din(w_G1691_0[1]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_n998_0[0]),.dinb(w_n1001_0[1]),.dout(n1002),.clk(gclk));
	jand g0702(.dina(w_n1002_4[1]),.dinb(w_n795_0[1]),.dout(n1003),.clk(gclk));
	jand g0703(.dina(w_G1694_0[1]),.dinb(w_n1001_0[0]),.dout(n1004),.clk(gclk));
	jand g0704(.dina(w_n1004_4[1]),.dinb(w_G182_0[0]),.dout(n1005),.clk(gclk));
	jand g0705(.dina(w_G1694_0[0]),.dinb(w_G1691_0[0]),.dout(n1006),.clk(gclk));
	jand g0706(.dina(w_n1006_4[1]),.dinb(w_G185_0[0]),.dout(n1007),.clk(gclk));
	jor g0707(.dina(w_dff_B_UPcddqAS5_0),.dinb(n1005),.dout(n1008),.clk(gclk));
	jor g0708(.dina(w_dff_B_zQrjFDnb9_0),.dinb(n1003),.dout(n1009),.clk(gclk));
	jor g0709(.dina(n1009),.dinb(n1000),.dout(n1010),.clk(gclk));
	jand g0710(.dina(n1010),.dinb(w_G137_9[0]),.dout(w_dff_A_eISRmwvG1_2),.clk(gclk));
	jnot g0711(.din(w_G871_0),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_1[1]),.dinb(w_n793_4[0]),.dout(n1013),.clk(gclk));
	jnot g0713(.din(w_G832_0),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_1[1]),.dinb(w_n797_4[0]),.dout(n1015),.clk(gclk));
	jand g0715(.dina(w_n799_4[0]),.dinb(w_G43_0[1]),.dout(n1016),.clk(gclk));
	jand g0716(.dina(w_n801_4[0]),.dinb(w_G37_0[1]),.dout(n1017),.clk(gclk));
	jor g0717(.dina(w_dff_B_tQiCExJB3_0),.dinb(n1016),.dout(n1018),.clk(gclk));
	jor g0718(.dina(w_dff_B_7oDXgmsj2_0),.dinb(n1015),.dout(n1019),.clk(gclk));
	jor g0719(.dina(w_dff_B_TJ0WxKdf1_0),.dinb(n1013),.dout(w_dff_A_pbgvSBrL9_2),.clk(gclk));
	jnot g0720(.din(w_G873_0),.dout(n1021),.clk(gclk));
	jand g0721(.dina(w_n1021_1[1]),.dinb(w_n793_3[2]),.dout(n1022),.clk(gclk));
	jnot g0722(.din(w_G834_0),.dout(n1023),.clk(gclk));
	jand g0723(.dina(w_n1023_1[1]),.dinb(w_n797_3[2]),.dout(n1024),.clk(gclk));
	jand g0724(.dina(w_n799_3[2]),.dinb(w_G76_0[1]),.dout(n1025),.clk(gclk));
	jand g0725(.dina(w_n801_3[2]),.dinb(w_G20_0[1]),.dout(n1026),.clk(gclk));
	jor g0726(.dina(w_dff_B_znZy9qvU2_0),.dinb(n1025),.dout(n1027),.clk(gclk));
	jor g0727(.dina(w_dff_B_B2O0Sk7l4_0),.dinb(n1024),.dout(n1028),.clk(gclk));
	jor g0728(.dina(w_dff_B_S0KAFPTt1_0),.dinb(n1022),.dout(w_dff_A_eFLyZN3r9_2),.clk(gclk));
	jnot g0729(.din(w_G875_0),.dout(n1030),.clk(gclk));
	jand g0730(.dina(w_n1030_1[1]),.dinb(w_n793_3[1]),.dout(n1031),.clk(gclk));
	jnot g0731(.din(w_G836_0),.dout(n1032),.clk(gclk));
	jand g0732(.dina(w_n1032_1[1]),.dinb(w_n797_3[1]),.dout(n1033),.clk(gclk));
	jand g0733(.dina(w_n799_3[1]),.dinb(w_G73_0[1]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(w_n801_3[1]),.dinb(w_G17_0[1]),.dout(n1035),.clk(gclk));
	jor g0735(.dina(w_dff_B_lcWxHoXi5_0),.dinb(n1034),.dout(n1036),.clk(gclk));
	jor g0736(.dina(w_dff_B_UXPXI8BI6_0),.dinb(n1033),.dout(n1037),.clk(gclk));
	jor g0737(.dina(w_dff_B_ffsg39Db4_0),.dinb(n1031),.dout(w_dff_A_SmweK2rc4_2),.clk(gclk));
	jnot g0738(.din(w_G877_0),.dout(n1039),.clk(gclk));
	jand g0739(.dina(w_n1039_1[1]),.dinb(w_n793_3[0]),.dout(n1040),.clk(gclk));
	jnot g0740(.din(w_G838_0),.dout(n1041),.clk(gclk));
	jand g0741(.dina(w_n797_3[0]),.dinb(w_n1041_1[1]),.dout(n1042),.clk(gclk));
	jand g0742(.dina(w_n799_3[0]),.dinb(w_G67_0[1]),.dout(n1043),.clk(gclk));
	jand g0743(.dina(w_n801_3[0]),.dinb(w_G70_0[1]),.dout(n1044),.clk(gclk));
	jor g0744(.dina(w_dff_B_6hnVM6k33_0),.dinb(n1043),.dout(n1045),.clk(gclk));
	jor g0745(.dina(w_dff_B_DtlcdPho4_0),.dinb(n1042),.dout(n1046),.clk(gclk));
	jor g0746(.dina(w_dff_B_eQZuP0F98_0),.dinb(n1040),.dout(w_dff_A_19H5GxO39_2),.clk(gclk));
	jand g0747(.dina(w_n1012_1[0]),.dinb(w_n840_4[0]),.dout(n1048),.clk(gclk));
	jand g0748(.dina(w_n843_4[0]),.dinb(w_n1014_1[0]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(w_n845_4[0]),.dinb(w_G43_0[0]),.dout(n1050),.clk(gclk));
	jand g0750(.dina(w_n847_4[0]),.dinb(w_G37_0[0]),.dout(n1051),.clk(gclk));
	jor g0751(.dina(w_dff_B_YLKUDv2t1_0),.dinb(n1050),.dout(n1052),.clk(gclk));
	jor g0752(.dina(w_dff_B_KvchqE8I4_0),.dinb(n1049),.dout(n1053),.clk(gclk));
	jor g0753(.dina(w_dff_B_VK4V7vCg1_0),.dinb(n1048),.dout(w_dff_A_pYaVT0Rd8_2),.clk(gclk));
	jand g0754(.dina(w_n1021_1[0]),.dinb(w_n840_3[2]),.dout(n1055),.clk(gclk));
	jand g0755(.dina(w_n843_3[2]),.dinb(w_n1023_1[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(w_n845_3[2]),.dinb(w_G76_0[0]),.dout(n1057),.clk(gclk));
	jand g0757(.dina(w_n847_3[2]),.dinb(w_G20_0[0]),.dout(n1058),.clk(gclk));
	jor g0758(.dina(w_dff_B_QPJoRHpB9_0),.dinb(n1057),.dout(n1059),.clk(gclk));
	jor g0759(.dina(w_dff_B_PBsKfb6g3_0),.dinb(n1056),.dout(n1060),.clk(gclk));
	jor g0760(.dina(w_dff_B_rOb8Gu7a6_0),.dinb(n1055),.dout(w_dff_A_zWQ5oN7u7_2),.clk(gclk));
	jand g0761(.dina(w_n1030_1[0]),.dinb(w_n840_3[1]),.dout(n1062),.clk(gclk));
	jand g0762(.dina(w_n843_3[1]),.dinb(w_n1032_1[0]),.dout(n1063),.clk(gclk));
	jand g0763(.dina(w_n845_3[1]),.dinb(w_G73_0[0]),.dout(n1064),.clk(gclk));
	jand g0764(.dina(w_n847_3[1]),.dinb(w_G17_0[0]),.dout(n1065),.clk(gclk));
	jor g0765(.dina(w_dff_B_rpkLrdoL7_0),.dinb(n1064),.dout(n1066),.clk(gclk));
	jor g0766(.dina(w_dff_B_eRBL8ZRO4_0),.dinb(n1063),.dout(n1067),.clk(gclk));
	jor g0767(.dina(w_dff_B_KKLryKvr9_0),.dinb(n1062),.dout(w_dff_A_3Phyc5ei6_2),.clk(gclk));
	jand g0768(.dina(w_n1039_1[0]),.dinb(w_n840_3[0]),.dout(n1069),.clk(gclk));
	jand g0769(.dina(w_n843_3[0]),.dinb(w_n1041_1[0]),.dout(n1070),.clk(gclk));
	jand g0770(.dina(w_n845_3[0]),.dinb(w_G67_0[0]),.dout(n1071),.clk(gclk));
	jand g0771(.dina(w_n847_3[0]),.dinb(w_G70_0[0]),.dout(n1072),.clk(gclk));
	jor g0772(.dina(w_dff_B_VVfb37309_0),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0773(.dina(w_dff_B_NIVGXwuL9_0),.dinb(n1070),.dout(n1074),.clk(gclk));
	jor g0774(.dina(w_dff_B_j39BeYFI8_0),.dinb(n1069),.dout(w_dff_A_kR71S9B18_2),.clk(gclk));
	jand g0775(.dina(w_n985_4[0]),.dinb(w_n1012_0[2]),.dout(n1076),.clk(gclk));
	jand g0776(.dina(w_n988_4[0]),.dinb(w_n1014_0[2]),.dout(n1077),.clk(gclk));
	jand g0777(.dina(w_n990_4[0]),.dinb(w_G200_0[1]),.dout(n1078),.clk(gclk));
	jand g0778(.dina(w_n992_4[0]),.dinb(w_G170_0[1]),.dout(n1079),.clk(gclk));
	jor g0779(.dina(w_dff_B_b2lq2Q2n7_0),.dinb(n1078),.dout(n1080),.clk(gclk));
	jor g0780(.dina(w_dff_B_1Kt4iVGy4_0),.dinb(n1077),.dout(n1081),.clk(gclk));
	jor g0781(.dina(w_dff_B_Y2Zix5Sa1_0),.dinb(n1076),.dout(n1082),.clk(gclk));
	jand g0782(.dina(n1082),.dinb(w_G137_8[2]),.dout(w_dff_A_K4P7N6hP0_2),.clk(gclk));
	jand g0783(.dina(w_n985_3[2]),.dinb(w_n1039_0[2]),.dout(n1084),.clk(gclk));
	jand g0784(.dina(w_n988_3[2]),.dinb(w_n1041_0[2]),.dout(n1085),.clk(gclk));
	jand g0785(.dina(w_n990_3[2]),.dinb(w_G188_0[1]),.dout(n1086),.clk(gclk));
	jand g0786(.dina(w_n992_3[2]),.dinb(w_G158_0[1]),.dout(n1087),.clk(gclk));
	jor g0787(.dina(w_dff_B_6OrtFTWs5_0),.dinb(n1086),.dout(n1088),.clk(gclk));
	jor g0788(.dina(w_dff_B_CWftwgeY8_0),.dinb(n1085),.dout(n1089),.clk(gclk));
	jor g0789(.dina(w_dff_B_zYIkRZYU7_0),.dinb(n1084),.dout(n1090),.clk(gclk));
	jand g0790(.dina(n1090),.dinb(w_G137_8[1]),.dout(w_dff_A_ezoq8C9i9_2),.clk(gclk));
	jand g0791(.dina(w_n985_3[1]),.dinb(w_n1030_0[2]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(w_n988_3[1]),.dinb(w_n1032_0[2]),.dout(n1093),.clk(gclk));
	jand g0793(.dina(w_n990_3[1]),.dinb(w_G155_0[1]),.dout(n1094),.clk(gclk));
	jand g0794(.dina(w_n992_3[1]),.dinb(w_G152_0[1]),.dout(n1095),.clk(gclk));
	jor g0795(.dina(w_dff_B_76PEudjL8_0),.dinb(n1094),.dout(n1096),.clk(gclk));
	jor g0796(.dina(w_dff_B_YWU8t7go8_0),.dinb(n1093),.dout(n1097),.clk(gclk));
	jor g0797(.dina(w_dff_B_rfDhlykd3_0),.dinb(n1092),.dout(n1098),.clk(gclk));
	jand g0798(.dina(n1098),.dinb(w_G137_8[0]),.dout(w_dff_A_gnv61TFV1_2),.clk(gclk));
	jand g0799(.dina(w_n985_3[0]),.dinb(w_n1021_0[2]),.dout(n1100),.clk(gclk));
	jand g0800(.dina(w_n988_3[0]),.dinb(w_n1023_0[2]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(w_n990_3[0]),.dinb(w_G149_0[1]),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n992_3[0]),.dinb(w_G146_0[1]),.dout(n1103),.clk(gclk));
	jor g0803(.dina(w_dff_B_BrlY33gH4_0),.dinb(n1102),.dout(n1104),.clk(gclk));
	jor g0804(.dina(w_dff_B_WAGQYCw72_0),.dinb(n1101),.dout(n1105),.clk(gclk));
	jor g0805(.dina(w_dff_B_oG0s388d4_0),.dinb(n1100),.dout(n1106),.clk(gclk));
	jand g0806(.dina(n1106),.dinb(w_G137_7[2]),.dout(w_dff_A_rJmF9iXA4_2),.clk(gclk));
	jand g0807(.dina(w_n999_4[0]),.dinb(w_n1012_0[1]),.dout(n1108),.clk(gclk));
	jand g0808(.dina(w_n1002_4[0]),.dinb(w_n1014_0[1]),.dout(n1109),.clk(gclk));
	jand g0809(.dina(w_n1004_4[0]),.dinb(w_G200_0[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(w_n1006_4[0]),.dinb(w_G170_0[0]),.dout(n1111),.clk(gclk));
	jor g0811(.dina(w_dff_B_Q5CYsc8T9_0),.dinb(n1110),.dout(n1112),.clk(gclk));
	jor g0812(.dina(w_dff_B_yTMNljsp9_0),.dinb(n1109),.dout(n1113),.clk(gclk));
	jor g0813(.dina(w_dff_B_SKrf3Cde8_0),.dinb(n1108),.dout(n1114),.clk(gclk));
	jand g0814(.dina(n1114),.dinb(w_G137_7[1]),.dout(w_dff_A_Ox1Xngjw7_2),.clk(gclk));
	jand g0815(.dina(w_n999_3[2]),.dinb(w_n1039_0[1]),.dout(n1116),.clk(gclk));
	jand g0816(.dina(w_n1002_3[2]),.dinb(w_n1041_0[1]),.dout(n1117),.clk(gclk));
	jand g0817(.dina(w_n1004_3[2]),.dinb(w_G188_0[0]),.dout(n1118),.clk(gclk));
	jand g0818(.dina(w_n1006_3[2]),.dinb(w_G158_0[0]),.dout(n1119),.clk(gclk));
	jor g0819(.dina(w_dff_B_0PbamN0N3_0),.dinb(n1118),.dout(n1120),.clk(gclk));
	jor g0820(.dina(w_dff_B_1waQ82K29_0),.dinb(n1117),.dout(n1121),.clk(gclk));
	jor g0821(.dina(w_dff_B_naGe759P5_0),.dinb(n1116),.dout(n1122),.clk(gclk));
	jand g0822(.dina(n1122),.dinb(w_G137_7[0]),.dout(w_dff_A_McN35ANS3_2),.clk(gclk));
	jand g0823(.dina(w_n999_3[1]),.dinb(w_n1030_0[1]),.dout(n1124),.clk(gclk));
	jand g0824(.dina(w_n1002_3[1]),.dinb(w_n1032_0[1]),.dout(n1125),.clk(gclk));
	jand g0825(.dina(w_n1004_3[1]),.dinb(w_G155_0[0]),.dout(n1126),.clk(gclk));
	jand g0826(.dina(w_n1006_3[1]),.dinb(w_G152_0[0]),.dout(n1127),.clk(gclk));
	jor g0827(.dina(w_dff_B_VTNitF7w1_0),.dinb(n1126),.dout(n1128),.clk(gclk));
	jor g0828(.dina(w_dff_B_57rtjik33_0),.dinb(n1125),.dout(n1129),.clk(gclk));
	jor g0829(.dina(w_dff_B_IL8mvxNn9_0),.dinb(n1124),.dout(n1130),.clk(gclk));
	jand g0830(.dina(n1130),.dinb(w_G137_6[2]),.dout(w_dff_A_EEV2iFkR2_2),.clk(gclk));
	jand g0831(.dina(w_n999_3[0]),.dinb(w_n1021_0[1]),.dout(n1132),.clk(gclk));
	jand g0832(.dina(w_n1002_3[0]),.dinb(w_n1023_0[1]),.dout(n1133),.clk(gclk));
	jand g0833(.dina(w_n1004_3[0]),.dinb(w_G149_0[0]),.dout(n1134),.clk(gclk));
	jand g0834(.dina(w_n1006_3[0]),.dinb(w_G146_0[0]),.dout(n1135),.clk(gclk));
	jor g0835(.dina(w_dff_B_vO706glE4_0),.dinb(n1134),.dout(n1136),.clk(gclk));
	jor g0836(.dina(w_dff_B_hy53SsrT2_0),.dinb(n1133),.dout(n1137),.clk(gclk));
	jor g0837(.dina(w_dff_B_03vhMbix5_0),.dinb(n1132),.dout(n1138),.clk(gclk));
	jand g0838(.dina(n1138),.dinb(w_G137_6[1]),.dout(w_dff_A_x965G86B7_2),.clk(gclk));
	jand g0839(.dina(w_n789_0[1]),.dinb(w_G3724_0[2]),.dout(n1140),.clk(gclk));
	jnot g0840(.din(w_G3717_0[1]),.dout(n1141),.clk(gclk));
	jnot g0841(.din(w_G3724_0[1]),.dout(n1142),.clk(gclk));
	jand g0842(.dina(w_n1142_0[1]),.dinb(w_G123_0[1]),.dout(n1143),.clk(gclk));
	jor g0843(.dina(n1143),.dinb(w_dff_B_Fdj4RatZ1_1),.dout(n1144),.clk(gclk));
	jor g0844(.dina(w_dff_B_THKPYsQ40_0),.dinb(n1140),.dout(n1145),.clk(gclk));
	jnot g0845(.din(G135),.dout(n1146),.clk(gclk));
	jnot g0846(.din(G4115),.dout(n1147),.clk(gclk));
	jor g0847(.dina(n1147),.dinb(n1146),.dout(n1148),.clk(gclk));
	jxor g0848(.dina(w_n636_0[1]),.dinb(w_G132_0[1]),.dout(n1149),.clk(gclk));
	jand g0849(.dina(n1149),.dinb(w_G3724_0[0]),.dout(n1150),.clk(gclk));
	jnot g0850(.din(w_n401_0[1]),.dout(n1151),.clk(gclk));
	jand g0851(.dina(w_n1151_0[1]),.dinb(w_n1142_0[0]),.dout(n1152),.clk(gclk));
	jor g0852(.dina(n1152),.dinb(w_G3717_0[0]),.dout(n1153),.clk(gclk));
	jor g0853(.dina(n1153),.dinb(w_dff_B_cAWCQ3GB5_1),.dout(n1154),.clk(gclk));
	jand g0854(.dina(n1154),.dinb(w_dff_B_VlWsDQyY4_1),.dout(n1155),.clk(gclk));
	jand g0855(.dina(w_dff_B_fONYaYHu7_0),.dinb(n1145),.dout(w_dff_A_YIjMVBcl3_2),.clk(gclk));
	jor g0856(.dina(w_n783_0[1]),.dinb(w_n640_0[2]),.dout(n1157),.clk(gclk));
	jxor g0857(.dina(n1157),.dinb(w_G132_0[0]),.dout(w_dff_A_VUuDR6GP3_2),.clk(gclk));
	jand g0858(.dina(w_n789_0[0]),.dinb(w_n747_2[1]),.dout(n1159),.clk(gclk));
	jand g0859(.dina(w_n753_5[0]),.dinb(w_G123_0[0]),.dout(n1160),.clk(gclk));
	jand g0860(.dina(w_n751_1[1]),.dinb(w_n1151_0[0]),.dout(n1161),.clk(gclk));
	jor g0861(.dina(n1161),.dinb(w_dff_B_kWE29rax3_1),.dout(n1162),.clk(gclk));
	jor g0862(.dina(w_dff_B_J5ifSxXj6_0),.dinb(n1159),.dout(n1163),.clk(gclk));
	jnot g0863(.din(w_n1163_1[2]),.dout(w_dff_A_dRifuz8t7_1),.clk(gclk));
	jor g0864(.dina(w_n972_0[0]),.dinb(w_n748_2[0]),.dout(n1165),.clk(gclk));
	jand g0865(.dina(w_n751_1[0]),.dinb(w_n407_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n753_4[2]),.dinb(w_dff_B_5BhY4KmB4_1),.dout(n1167),.clk(gclk));
	jor g0867(.dina(w_dff_B_V7eyhQDU8_0),.dinb(n1166),.dout(n1168),.clk(gclk));
	jnot g0868(.din(n1168),.dout(n1169),.clk(gclk));
	jand g0869(.dina(w_dff_B_x44aRKhf9_0),.dinb(n1165),.dout(G826_fa_),.clk(gclk));
	jor g0870(.dina(w_n971_0[0]),.dinb(w_n748_1[2]),.dout(n1171),.clk(gclk));
	jor g0871(.dina(w_n765_3[0]),.dinb(w_n372_0[1]),.dout(n1172),.clk(gclk));
	jand g0872(.dina(w_n753_4[1]),.dinb(w_dff_B_XSMluYwI5_1),.dout(n1173),.clk(gclk));
	jnot g0873(.din(n1173),.dout(n1174),.clk(gclk));
	jand g0874(.dina(w_dff_B_ua2pDzep4_0),.dinb(n1172),.dout(n1175),.clk(gclk));
	jand g0875(.dina(w_dff_B_hkmYepsr1_0),.dinb(n1171),.dout(G828_fa_),.clk(gclk));
	jand g0876(.dina(w_n973_0[0]),.dinb(w_n747_2[0]),.dout(n1177),.clk(gclk));
	jnot g0877(.din(n1177),.dout(n1178),.clk(gclk));
	jor g0878(.dina(w_n765_2[2]),.dinb(w_n383_0[1]),.dout(n1179),.clk(gclk));
	jand g0879(.dina(w_n753_4[0]),.dinb(w_dff_B_X0uLgB6d7_1),.dout(n1180),.clk(gclk));
	jnot g0880(.din(n1180),.dout(n1181),.clk(gclk));
	jand g0881(.dina(w_dff_B_L7sOoYjC0_0),.dinb(n1179),.dout(n1182),.clk(gclk));
	jand g0882(.dina(w_dff_B_iJl25Ho34_0),.dinb(n1178),.dout(G830_fa_),.clk(gclk));
	jnot g0883(.din(w_G1000_0),.dout(n1184),.clk(gclk));
	jand g0884(.dina(w_G559_0[0]),.dinb(w_G245_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(n1185),.dinb(w_n318_0[0]),.dout(n1186),.clk(gclk));
	jand g0886(.dina(n1186),.dinb(w_G601_0),.dout(n1187),.clk(gclk));
	jand g0887(.dina(w_dff_B_ZPdVBZ620_0),.dinb(w_n661_0[0]),.dout(n1188),.clk(gclk));
	jand g0888(.dina(n1188),.dinb(w_n671_0[0]),.dout(n1189),.clk(gclk));
	jand g0889(.dina(w_dff_B_NIssC7zS7_0),.dinb(w_n914_0[0]),.dout(n1190),.clk(gclk));
	jand g0890(.dina(n1190),.dinb(w_dff_B_kEvZGrFN3_1),.dout(w_dff_A_dWiR3lKc9_2),.clk(gclk));
	jand g0891(.dina(w_n941_0[0]),.dinb(w_n747_1[2]),.dout(n1192),.clk(gclk));
	jnot g0892(.din(w_n528_0[1]),.dout(n1193),.clk(gclk));
	jand g0893(.dina(w_n751_0[2]),.dinb(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_n753_3[2]),.dinb(w_dff_B_iunU92P06_1),.dout(n1195),.clk(gclk));
	jor g0895(.dina(w_dff_B_QVpp9gnE7_0),.dinb(n1194),.dout(n1196),.clk(gclk));
	jor g0896(.dina(w_dff_B_jKj3SKn22_0),.dinb(n1192),.dout(n1197),.clk(gclk));
	jnot g0897(.din(w_n1197_1[2]),.dout(w_dff_A_YbUu0rt76_1),.clk(gclk));
	jand g0898(.dina(w_n946_0[0]),.dinb(w_n747_1[1]),.dout(n1199),.clk(gclk));
	jor g0899(.dina(w_n765_2[1]),.dinb(w_n551_0[0]),.dout(n1200),.clk(gclk));
	jand g0900(.dina(w_n753_3[1]),.dinb(w_dff_B_LjNP1xe75_1),.dout(n1201),.clk(gclk));
	jnot g0901(.din(n1201),.dout(n1202),.clk(gclk));
	jand g0902(.dina(w_dff_B_7NIGw5Oa9_0),.dinb(n1200),.dout(n1203),.clk(gclk));
	jnot g0903(.din(n1203),.dout(n1204),.clk(gclk));
	jor g0904(.dina(w_dff_B_Nq2ZTkki8_0),.dinb(n1199),.dout(n1205),.clk(gclk));
	jnot g0905(.din(w_n1205_1[2]),.dout(w_dff_A_jFPW27Js2_1),.clk(gclk));
	jor g0906(.dina(w_n953_0[0]),.dinb(w_n748_1[1]),.dout(n1207),.clk(gclk));
	jor g0907(.dina(w_n765_2[0]),.dinb(w_n517_0[0]),.dout(n1208),.clk(gclk));
	jand g0908(.dina(w_n753_3[0]),.dinb(w_dff_B_ZA4O3y686_1),.dout(n1209),.clk(gclk));
	jnot g0909(.din(n1209),.dout(n1210),.clk(gclk));
	jand g0910(.dina(w_dff_B_CFEHNOeE2_0),.dinb(n1208),.dout(n1211),.clk(gclk));
	jand g0911(.dina(w_dff_B_lC30vCYl0_0),.dinb(n1207),.dout(G867_fa_),.clk(gclk));
	jand g0912(.dina(w_n954_0[0]),.dinb(w_n747_1[0]),.dout(n1213),.clk(gclk));
	jnot g0913(.din(n1213),.dout(n1214),.clk(gclk));
	jor g0914(.dina(w_n765_1[2]),.dinb(w_n540_0[0]),.dout(n1215),.clk(gclk));
	jand g0915(.dina(w_n753_2[2]),.dinb(w_dff_B_glA5B8U56_1),.dout(n1216),.clk(gclk));
	jnot g0916(.din(n1216),.dout(n1217),.clk(gclk));
	jand g0917(.dina(w_dff_B_7kBC6HHg6_0),.dinb(n1215),.dout(n1218),.clk(gclk));
	jand g0918(.dina(w_dff_B_IUk8gXyh9_0),.dinb(n1214),.dout(G869_fa_),.clk(gclk));
	jand g0919(.dina(w_n1197_1[1]),.dinb(w_n840_2[2]),.dout(n1220),.clk(gclk));
	jand g0920(.dina(w_n1163_1[1]),.dinb(w_n843_2[2]),.dout(n1221),.clk(gclk));
	jand g0921(.dina(w_n845_2[2]),.dinb(w_G109_0[1]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(w_n847_2[2]),.dinb(w_G106_0[1]),.dout(n1223),.clk(gclk));
	jor g0923(.dina(w_dff_B_QXWGfaW84_0),.dinb(n1222),.dout(n1224),.clk(gclk));
	jor g0924(.dina(w_dff_B_fE20assw7_0),.dinb(n1221),.dout(n1225),.clk(gclk));
	jor g0925(.dina(n1225),.dinb(n1220),.dout(w_dff_A_nWpQUXif7_2),.clk(gclk));
	jand g0926(.dina(w_n1197_1[0]),.dinb(w_n793_2[2]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_n1163_1[0]),.dinb(w_n797_2[2]),.dout(n1228),.clk(gclk));
	jand g0928(.dina(w_n799_2[2]),.dinb(w_G109_0[0]),.dout(n1229),.clk(gclk));
	jand g0929(.dina(w_n801_2[2]),.dinb(w_G106_0[0]),.dout(n1230),.clk(gclk));
	jor g0930(.dina(w_dff_B_lrLLoZaM8_0),.dinb(n1229),.dout(n1231),.clk(gclk));
	jor g0931(.dina(w_dff_B_eUoyMdux2_0),.dinb(n1228),.dout(n1232),.clk(gclk));
	jor g0932(.dina(n1232),.dinb(n1227),.dout(w_dff_A_wC6dLpOY8_2),.clk(gclk));
	jand g0933(.dina(w_n1205_1[1]),.dinb(w_n793_2[1]),.dout(n1234),.clk(gclk));
	jnot g0934(.din(w_G826_0),.dout(n1235),.clk(gclk));
	jand g0935(.dina(w_n1235_1[1]),.dinb(w_n797_2[1]),.dout(n1236),.clk(gclk));
	jand g0936(.dina(w_n799_2[1]),.dinb(w_G46_0[1]),.dout(n1237),.clk(gclk));
	jand g0937(.dina(w_n801_2[1]),.dinb(w_G49_0[1]),.dout(n1238),.clk(gclk));
	jor g0938(.dina(w_dff_B_Foucat1g1_0),.dinb(n1237),.dout(n1239),.clk(gclk));
	jor g0939(.dina(w_dff_B_0JrtqFgk8_0),.dinb(n1236),.dout(n1240),.clk(gclk));
	jor g0940(.dina(n1240),.dinb(n1234),.dout(w_dff_A_aOg13yvN6_2),.clk(gclk));
	jnot g0941(.din(w_G867_0),.dout(n1242),.clk(gclk));
	jand g0942(.dina(w_n1242_1[1]),.dinb(w_n793_2[0]),.dout(n1243),.clk(gclk));
	jnot g0943(.din(w_G828_0),.dout(n1244),.clk(gclk));
	jand g0944(.dina(w_n1244_1[1]),.dinb(w_n797_2[0]),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n799_2[0]),.dinb(w_G100_0[1]),.dout(n1246),.clk(gclk));
	jand g0946(.dina(w_n801_2[0]),.dinb(w_G103_0[1]),.dout(n1247),.clk(gclk));
	jor g0947(.dina(w_dff_B_3LcSg0uW3_0),.dinb(n1246),.dout(n1248),.clk(gclk));
	jor g0948(.dina(w_dff_B_qiaSDrf53_0),.dinb(n1245),.dout(n1249),.clk(gclk));
	jor g0949(.dina(n1249),.dinb(n1243),.dout(w_dff_A_Gz7SUmwg3_2),.clk(gclk));
	jnot g0950(.din(w_G869_0),.dout(n1251),.clk(gclk));
	jand g0951(.dina(w_n1251_1[1]),.dinb(w_n793_1[2]),.dout(n1252),.clk(gclk));
	jnot g0952(.din(w_G830_0),.dout(n1253),.clk(gclk));
	jand g0953(.dina(w_n1253_1[1]),.dinb(w_n797_1[2]),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n799_1[2]),.dinb(w_G91_0[1]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n801_1[2]),.dinb(w_G40_0[1]),.dout(n1256),.clk(gclk));
	jor g0956(.dina(w_dff_B_K4fKwws38_0),.dinb(n1255),.dout(n1257),.clk(gclk));
	jor g0957(.dina(w_dff_B_1xKtCMCP1_0),.dinb(n1254),.dout(n1258),.clk(gclk));
	jor g0958(.dina(n1258),.dinb(n1252),.dout(w_dff_A_Kj9RkwBZ2_2),.clk(gclk));
	jand g0959(.dina(w_n1205_1[0]),.dinb(w_n840_2[1]),.dout(n1260),.clk(gclk));
	jand g0960(.dina(w_n1235_1[0]),.dinb(w_n843_2[1]),.dout(n1261),.clk(gclk));
	jand g0961(.dina(w_n845_2[1]),.dinb(w_G46_0[0]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(w_n847_2[1]),.dinb(w_G49_0[0]),.dout(n1263),.clk(gclk));
	jor g0963(.dina(w_dff_B_8DjwxO8J4_0),.dinb(n1262),.dout(n1264),.clk(gclk));
	jor g0964(.dina(w_dff_B_HfR9NiRb5_0),.dinb(n1261),.dout(n1265),.clk(gclk));
	jor g0965(.dina(n1265),.dinb(n1260),.dout(w_dff_A_r913b9Tx0_2),.clk(gclk));
	jand g0966(.dina(w_n1242_1[0]),.dinb(w_n840_2[0]),.dout(n1267),.clk(gclk));
	jand g0967(.dina(w_n1244_1[0]),.dinb(w_n843_2[0]),.dout(n1268),.clk(gclk));
	jand g0968(.dina(w_n845_2[0]),.dinb(w_G100_0[0]),.dout(n1269),.clk(gclk));
	jand g0969(.dina(w_n847_2[0]),.dinb(w_G103_0[0]),.dout(n1270),.clk(gclk));
	jor g0970(.dina(w_dff_B_p0dtSfDh5_0),.dinb(n1269),.dout(n1271),.clk(gclk));
	jor g0971(.dina(w_dff_B_jgcc0Xlp3_0),.dinb(n1268),.dout(n1272),.clk(gclk));
	jor g0972(.dina(n1272),.dinb(n1267),.dout(w_dff_A_B7zzNCht4_2),.clk(gclk));
	jand g0973(.dina(w_n1251_1[0]),.dinb(w_n840_1[2]),.dout(n1274),.clk(gclk));
	jand g0974(.dina(w_n1253_1[0]),.dinb(w_n843_1[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(w_n845_1[2]),.dinb(w_G91_0[0]),.dout(n1276),.clk(gclk));
	jand g0976(.dina(w_n847_1[2]),.dinb(w_G40_0[0]),.dout(n1277),.clk(gclk));
	jor g0977(.dina(w_dff_B_2V4gCxYY5_0),.dinb(n1276),.dout(n1278),.clk(gclk));
	jor g0978(.dina(w_dff_B_4ZPfSibY8_0),.dinb(n1275),.dout(n1279),.clk(gclk));
	jor g0979(.dina(n1279),.dinb(n1274),.dout(w_dff_A_zAFhLVgo8_2),.clk(gclk));
	jand g0980(.dina(w_n1251_0[2]),.dinb(w_n985_2[2]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(w_n1253_0[2]),.dinb(w_n988_2[2]),.dout(n1282),.clk(gclk));
	jand g0982(.dina(w_n990_2[2]),.dinb(w_G203_0[1]),.dout(n1283),.clk(gclk));
	jand g0983(.dina(w_n992_2[2]),.dinb(w_G173_0[1]),.dout(n1284),.clk(gclk));
	jor g0984(.dina(w_dff_B_CLS7VxaR5_0),.dinb(n1283),.dout(n1285),.clk(gclk));
	jor g0985(.dina(w_dff_B_kCrwhqOF3_0),.dinb(n1282),.dout(n1286),.clk(gclk));
	jor g0986(.dina(n1286),.dinb(n1281),.dout(n1287),.clk(gclk));
	jand g0987(.dina(n1287),.dinb(w_G137_6[0]),.dout(w_dff_A_IHkscreG0_2),.clk(gclk));
	jand g0988(.dina(w_n1242_0[2]),.dinb(w_n985_2[1]),.dout(n1289),.clk(gclk));
	jand g0989(.dina(w_n1244_0[2]),.dinb(w_n988_2[1]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(w_n990_2[1]),.dinb(w_G197_0[1]),.dout(n1291),.clk(gclk));
	jand g0991(.dina(w_n992_2[1]),.dinb(w_G167_0[1]),.dout(n1292),.clk(gclk));
	jor g0992(.dina(w_dff_B_wHs13Xsv8_0),.dinb(n1291),.dout(n1293),.clk(gclk));
	jor g0993(.dina(w_dff_B_xkI0oTdo9_0),.dinb(n1290),.dout(n1294),.clk(gclk));
	jor g0994(.dina(n1294),.dinb(n1289),.dout(n1295),.clk(gclk));
	jand g0995(.dina(n1295),.dinb(w_G137_5[2]),.dout(w_dff_A_waPH8W0z0_2),.clk(gclk));
	jand g0996(.dina(w_n1205_0[2]),.dinb(w_n985_2[0]),.dout(n1297),.clk(gclk));
	jand g0997(.dina(w_n1235_0[2]),.dinb(w_n988_2[0]),.dout(n1298),.clk(gclk));
	jand g0998(.dina(w_n990_2[0]),.dinb(w_G194_0[1]),.dout(n1299),.clk(gclk));
	jand g0999(.dina(w_n992_2[0]),.dinb(w_G164_0[1]),.dout(n1300),.clk(gclk));
	jor g1000(.dina(w_dff_B_2lnt7ZZc6_0),.dinb(n1299),.dout(n1301),.clk(gclk));
	jor g1001(.dina(w_dff_B_Gkx80q075_0),.dinb(n1298),.dout(n1302),.clk(gclk));
	jor g1002(.dina(n1302),.dinb(n1297),.dout(n1303),.clk(gclk));
	jand g1003(.dina(n1303),.dinb(w_G137_5[1]),.dout(w_dff_A_Ma7drrNq3_2),.clk(gclk));
	jand g1004(.dina(w_n1197_0[2]),.dinb(w_n985_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(w_n1163_0[2]),.dinb(w_n988_1[2]),.dout(n1306),.clk(gclk));
	jand g1006(.dina(w_n990_1[2]),.dinb(w_G191_0[1]),.dout(n1307),.clk(gclk));
	jand g1007(.dina(w_n992_1[2]),.dinb(w_G161_0[1]),.dout(n1308),.clk(gclk));
	jor g1008(.dina(w_dff_B_oir3KOd09_0),.dinb(n1307),.dout(n1309),.clk(gclk));
	jor g1009(.dina(w_dff_B_lClUUBK73_0),.dinb(n1306),.dout(n1310),.clk(gclk));
	jor g1010(.dina(n1310),.dinb(n1305),.dout(n1311),.clk(gclk));
	jand g1011(.dina(n1311),.dinb(w_G137_5[0]),.dout(w_dff_A_CSW3oR7E2_2),.clk(gclk));
	jand g1012(.dina(w_n1251_0[1]),.dinb(w_n999_2[2]),.dout(n1313),.clk(gclk));
	jand g1013(.dina(w_n1253_0[1]),.dinb(w_n1002_2[2]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(w_n1004_2[2]),.dinb(w_G203_0[0]),.dout(n1315),.clk(gclk));
	jand g1015(.dina(w_n1006_2[2]),.dinb(w_G173_0[0]),.dout(n1316),.clk(gclk));
	jor g1016(.dina(w_dff_B_hu36JLKP8_0),.dinb(n1315),.dout(n1317),.clk(gclk));
	jor g1017(.dina(w_dff_B_qNDrs8HS5_0),.dinb(n1314),.dout(n1318),.clk(gclk));
	jor g1018(.dina(n1318),.dinb(n1313),.dout(n1319),.clk(gclk));
	jand g1019(.dina(n1319),.dinb(w_G137_4[2]),.dout(w_dff_A_jCh5PqgI7_2),.clk(gclk));
	jand g1020(.dina(w_n1242_0[1]),.dinb(w_n999_2[1]),.dout(n1321),.clk(gclk));
	jand g1021(.dina(w_n1244_0[1]),.dinb(w_n1002_2[1]),.dout(n1322),.clk(gclk));
	jand g1022(.dina(w_n1004_2[1]),.dinb(w_G197_0[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(w_n1006_2[1]),.dinb(w_G167_0[0]),.dout(n1324),.clk(gclk));
	jor g1024(.dina(w_dff_B_PVzDrUI07_0),.dinb(n1323),.dout(n1325),.clk(gclk));
	jor g1025(.dina(w_dff_B_gjb4Oi0q0_0),.dinb(n1322),.dout(n1326),.clk(gclk));
	jor g1026(.dina(n1326),.dinb(n1321),.dout(n1327),.clk(gclk));
	jand g1027(.dina(n1327),.dinb(w_G137_4[1]),.dout(w_dff_A_QI9HYEpX5_2),.clk(gclk));
	jand g1028(.dina(w_n1205_0[1]),.dinb(w_n999_2[0]),.dout(n1329),.clk(gclk));
	jand g1029(.dina(w_n1235_0[1]),.dinb(w_n1002_2[0]),.dout(n1330),.clk(gclk));
	jand g1030(.dina(w_n1004_2[0]),.dinb(w_G194_0[0]),.dout(n1331),.clk(gclk));
	jand g1031(.dina(w_n1006_2[0]),.dinb(w_G164_0[0]),.dout(n1332),.clk(gclk));
	jor g1032(.dina(w_dff_B_E09Mezaa2_0),.dinb(n1331),.dout(n1333),.clk(gclk));
	jor g1033(.dina(w_dff_B_aAqwkRiN8_0),.dinb(n1330),.dout(n1334),.clk(gclk));
	jor g1034(.dina(n1334),.dinb(n1329),.dout(n1335),.clk(gclk));
	jand g1035(.dina(n1335),.dinb(w_G137_4[0]),.dout(w_dff_A_MbjnhRRh3_2),.clk(gclk));
	jand g1036(.dina(w_n1197_0[1]),.dinb(w_n999_1[2]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(w_n1163_0[1]),.dinb(w_n1002_1[2]),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n1004_1[2]),.dinb(w_G191_0[0]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n1006_1[2]),.dinb(w_G161_0[0]),.dout(n1340),.clk(gclk));
	jor g1040(.dina(w_dff_B_CDnC17cx4_0),.dinb(n1339),.dout(n1341),.clk(gclk));
	jor g1041(.dina(w_dff_B_nfMwAaDh9_0),.dinb(n1338),.dout(n1342),.clk(gclk));
	jor g1042(.dina(n1342),.dinb(n1337),.dout(n1343),.clk(gclk));
	jand g1043(.dina(n1343),.dinb(w_G137_3[2]),.dout(w_dff_A_j5GasjKW1_2),.clk(gclk));
	jor g1044(.dina(w_G4091_2[0]),.dinb(G120),.dout(n1345),.clk(gclk));
	jand g1045(.dina(w_n435_0[2]),.dinb(w_G251_3[1]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1347),.clk(gclk));
	jor g1047(.dina(n1347),.dinb(w_n437_0[1]),.dout(n1348),.clk(gclk));
	jor g1048(.dina(n1348),.dinb(n1346),.dout(n1349),.clk(gclk));
	jand g1049(.dina(w_n435_0[1]),.dinb(w_n366_3[1]),.dout(n1350),.clk(gclk));
	jand g1050(.dina(w_G341_0[2]),.dinb(w_n368_4[0]),.dout(n1351),.clk(gclk));
	jor g1051(.dina(n1351),.dinb(w_G523_0[2]),.dout(n1352),.clk(gclk));
	jor g1052(.dina(n1352),.dinb(w_dff_B_Ycv7c5LF4_1),.dout(n1353),.clk(gclk));
	jand g1053(.dina(n1353),.dinb(w_dff_B_PWP6gSHG7_1),.dout(n1354),.clk(gclk));
	jxor g1054(.dina(w_n408_0[0]),.dinb(w_n401_0[0]),.dout(n1355),.clk(gclk));
	jxor g1055(.dina(w_n383_0[0]),.dinb(w_n372_0[0]),.dout(n1356),.clk(gclk));
	jxor g1056(.dina(n1356),.dinb(w_dff_B_B0WxHOIX3_1),.dout(n1357),.clk(gclk));
	jxor g1057(.dina(n1357),.dinb(w_dff_B_vc2CbMzP1_1),.dout(n1358),.clk(gclk));
	jnot g1058(.din(w_n1358_0[1]),.dout(n1359),.clk(gclk));
	jor g1059(.dina(w_n410_0[1]),.dinb(w_G248_3[2]),.dout(n1360),.clk(gclk));
	jor g1060(.dina(w_G514_0[1]),.dinb(w_n368_3[2]),.dout(n1361),.clk(gclk));
	jand g1061(.dina(n1361),.dinb(n1360),.dout(n1362),.clk(gclk));
	jxor g1062(.dina(n1362),.dinb(w_n419_0[0]),.dout(n1363),.clk(gclk));
	jor g1063(.dina(w_G351_1[0]),.dinb(w_n402_1[2]),.dout(n1364),.clk(gclk));
	jor g1064(.dina(w_n385_0[2]),.dinb(w_n405_1[2]),.dout(n1365),.clk(gclk));
	jand g1065(.dina(n1365),.dinb(w_G534_0[1]),.dout(n1366),.clk(gclk));
	jand g1066(.dina(n1366),.dinb(w_dff_B_5j4gjsAx5_1),.dout(n1367),.clk(gclk));
	jor g1067(.dina(w_G351_0[2]),.dinb(w_G254_1[1]),.dout(n1368),.clk(gclk));
	jor g1068(.dina(w_n385_0[1]),.dinb(w_G242_1[1]),.dout(n1369),.clk(gclk));
	jand g1069(.dina(n1369),.dinb(w_n388_0[1]),.dout(n1370),.clk(gclk));
	jand g1070(.dina(n1370),.dinb(w_dff_B_a6IBdNjb5_1),.dout(n1371),.clk(gclk));
	jor g1071(.dina(n1371),.dinb(n1367),.dout(n1372),.clk(gclk));
	jand g1072(.dina(w_n424_1[0]),.dinb(w_G251_3[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(w_G324_0[2]),.dinb(w_G248_3[1]),.dout(n1374),.clk(gclk));
	jor g1074(.dina(n1374),.dinb(w_n426_0[0]),.dout(n1375),.clk(gclk));
	jor g1075(.dina(n1375),.dinb(n1373),.dout(n1376),.clk(gclk));
	jand g1076(.dina(w_n424_0[2]),.dinb(w_n366_3[0]),.dout(n1377),.clk(gclk));
	jand g1077(.dina(w_G324_0[1]),.dinb(w_n368_3[1]),.dout(n1378),.clk(gclk));
	jor g1078(.dina(n1378),.dinb(w_G503_0[1]),.dout(n1379),.clk(gclk));
	jor g1079(.dina(n1379),.dinb(w_dff_B_MNXlIaF17_1),.dout(n1380),.clk(gclk));
	jand g1080(.dina(n1380),.dinb(w_dff_B_aN7DnGVD7_1),.dout(n1381),.clk(gclk));
	jxor g1081(.dina(n1381),.dinb(n1372),.dout(n1382),.clk(gclk));
	jxor g1082(.dina(n1382),.dinb(w_dff_B_hfwAfqic5_1),.dout(n1383),.clk(gclk));
	jnot g1083(.din(w_n1383_0[1]),.dout(n1384),.clk(gclk));
	jand g1084(.dina(w_n1383_0[0]),.dinb(n1359),.dout(n1385),.clk(gclk));
	jor g1085(.dina(n1385),.dinb(w_G4091_1[2]),.dout(n1386),.clk(gclk));
	jor g1086(.dina(n1345),.dinb(w_n746_1[0]),.dout(n1388),.clk(gclk));
	jand g1087(.dina(n1384),.dinb(w_n1358_0[0]),.dout(n1389),.clk(gclk));
	jor g1088(.dina(n1386),.dinb(w_dff_B_l1aSVjxa3_1),.dout(n1390),.clk(gclk));
	jand g1089(.dina(n1390),.dinb(w_n746_0[2]),.dout(n1391),.clk(gclk));
	jnot g1090(.din(w_n1391_0[1]),.dout(n1392),.clk(gclk));
	jand g1091(.dina(w_n633_0[2]),.dinb(w_G2174_0[2]),.dout(n1393),.clk(gclk));
	jor g1092(.dina(w_dff_B_l1uAx0AP2_0),.dinb(w_n732_0[0]),.dout(n1394),.clk(gclk));
	jand g1093(.dina(w_n736_0[0]),.dinb(w_n640_0[1]),.dout(n1395),.clk(gclk));
	jor g1094(.dina(w_n740_0[0]),.dinb(w_n641_0[0]),.dout(n1396),.clk(gclk));
	jand g1095(.dina(n1396),.dinb(w_n646_0[0]),.dout(n1397),.clk(gclk));
	jor g1096(.dina(n1397),.dinb(w_dff_B_GtX4MKB26_1),.dout(n1398),.clk(gclk));
	jnot g1097(.din(w_n1398_0[1]),.dout(n1399),.clk(gclk));
	jand g1098(.dina(w_n1399_0[1]),.dinb(w_n739_0[2]),.dout(n1400),.clk(gclk));
	jnot g1099(.din(w_n739_0[1]),.dout(n1401),.clk(gclk));
	jand g1100(.dina(w_n1398_0[0]),.dinb(w_dff_B_eM51dZqn7_1),.dout(n1402),.clk(gclk));
	jor g1101(.dina(n1402),.dinb(w_n651_0[1]),.dout(n1403),.clk(gclk));
	jor g1102(.dina(n1403),.dinb(n1400),.dout(n1404),.clk(gclk));
	jand g1103(.dina(w_dff_B_fdXgcZAc6_0),.dinb(w_n1394_0[1]),.dout(n1405),.clk(gclk));
	jnot g1104(.din(w_n1394_0[0]),.dout(n1406),.clk(gclk));
	jxor g1105(.dina(w_n1399_0[0]),.dinb(w_n968_0[0]),.dout(n1407),.clk(gclk));
	jand g1106(.dina(w_dff_B_9ODYf6pV6_0),.dinb(n1406),.dout(n1408),.clk(gclk));
	jor g1107(.dina(n1408),.dinb(w_dff_B_AOf3PMd74_1),.dout(n1409),.clk(gclk));
	jnot g1108(.din(w_n1409_0[1]),.dout(n1410),.clk(gclk));
	jxor g1109(.dina(w_n629_0[0]),.dinb(w_n625_0[0]),.dout(n1411),.clk(gclk));
	jnot g1110(.din(w_n1411_0[1]),.dout(n1412),.clk(gclk));
	jxor g1111(.dina(w_n806_0[1]),.dinb(w_n828_0[1]),.dout(n1413),.clk(gclk));
	jnot g1112(.din(w_n614_1[1]),.dout(n1414),.clk(gclk));
	jnot g1113(.din(w_n717_0[0]),.dout(n1415),.clk(gclk));
	jand g1114(.dina(w_n622_1[0]),.dinb(w_n828_0[0]),.dout(n1416),.clk(gclk));
	jand g1115(.dina(w_n628_0[0]),.dinb(w_G523_0[1]),.dout(n1417),.clk(gclk));
	jor g1116(.dina(n1417),.dinb(w_n829_0[0]),.dout(n1418),.clk(gclk));
	jor g1117(.dina(n1418),.dinb(n1416),.dout(n1419),.clk(gclk));
	jand g1118(.dina(n1419),.dinb(w_dff_B_AHQpbTXO6_1),.dout(n1420),.clk(gclk));
	jxor g1119(.dina(w_n622_0[2]),.dinb(w_n618_0[1]),.dout(n1421),.clk(gclk));
	jnot g1120(.din(w_n1421_0[1]),.dout(n1422),.clk(gclk));
	jor g1121(.dina(w_dff_B_fXge62pK6_0),.dinb(n1420),.dout(n1423),.clk(gclk));
	jor g1122(.dina(w_n1421_0[0]),.dinb(w_n819_0[0]),.dout(n1424),.clk(gclk));
	jand g1123(.dina(n1424),.dinb(w_dff_B_jPIh30mM3_1),.dout(n1425),.clk(gclk));
	jxor g1124(.dina(w_n1425_0[1]),.dinb(w_dff_B_vj4uRcAr3_1),.dout(n1426),.clk(gclk));
	jand g1125(.dina(n1426),.dinb(n1413),.dout(n1427),.clk(gclk));
	jnot g1126(.din(w_G2174_0[1]),.dout(n1428),.clk(gclk));
	jxor g1127(.dina(w_n806_0[0]),.dinb(w_n721_0[1]),.dout(n1429),.clk(gclk));
	jxor g1128(.dina(w_n1425_0[0]),.dinb(w_n614_1[0]),.dout(n1430),.clk(gclk));
	jand g1129(.dina(n1430),.dinb(n1429),.dout(n1431),.clk(gclk));
	jor g1130(.dina(n1431),.dinb(w_dff_B_7J4yUeo43_1),.dout(n1432),.clk(gclk));
	jor g1131(.dina(n1432),.dinb(w_dff_B_dFCMmpUR1_1),.dout(n1433),.clk(gclk));
	jxor g1132(.dina(w_n729_0[1]),.dinb(w_n614_0[2]),.dout(n1434),.clk(gclk));
	jnot g1133(.din(w_n1434_0[1]),.dout(n1435),.clk(gclk));
	jor g1134(.dina(w_n622_0[1]),.dinb(w_n721_0[0]),.dout(n1436),.clk(gclk));
	jand g1135(.dina(n1436),.dinb(w_n723_0[0]),.dout(n1437),.clk(gclk));
	jxor g1136(.dina(w_dff_B_y9QNuL3z4_0),.dinb(w_n727_0[0]),.dout(n1438),.clk(gclk));
	jand g1137(.dina(w_n1438_0[1]),.dinb(n1435),.dout(n1439),.clk(gclk));
	jnot g1138(.din(w_n1438_0[0]),.dout(n1440),.clk(gclk));
	jand g1139(.dina(w_dff_B_9GLwzPEr8_0),.dinb(w_n1434_0[0]),.dout(n1441),.clk(gclk));
	jor g1140(.dina(n1441),.dinb(w_G2174_0[0]),.dout(n1442),.clk(gclk));
	jor g1141(.dina(n1442),.dinb(n1439),.dout(n1443),.clk(gclk));
	jand g1142(.dina(w_dff_B_ANg88wro8_0),.dinb(n1433),.dout(n1444),.clk(gclk));
	jxor g1143(.dina(n1444),.dinb(w_n787_0[0]),.dout(n1445),.clk(gclk));
	jxor g1144(.dina(w_n1445_0[1]),.dinb(w_dff_B_d8pD8Ezv4_1),.dout(n1446),.clk(gclk));
	jor g1145(.dina(w_n1446_0[1]),.dinb(w_n1410_0[1]),.dout(n1447),.clk(gclk));
	jxor g1146(.dina(w_n1445_0[0]),.dinb(w_n1411_0[0]),.dout(n1448),.clk(gclk));
	jor g1147(.dina(n1448),.dinb(w_n1409_0[0]),.dout(n1449),.clk(gclk));
	jand g1148(.dina(n1449),.dinb(w_G4091_1[1]),.dout(n1450),.clk(gclk));
	jand g1149(.dina(n1450),.dinb(w_n1447_0[1]),.dout(n1451),.clk(gclk));
	jor g1150(.dina(n1451),.dinb(w_dff_B_CQpW27lF9_1),.dout(n1452),.clk(gclk));
	jand g1151(.dina(w_n1452_0[1]),.dinb(w_dff_B_tlTNiJrb5_1),.dout(w_dff_A_JuKIKgog1_2),.clk(gclk));
	jor g1152(.dina(w_G4091_1[0]),.dinb(G118),.dout(n1454),.clk(gclk));
	jand g1153(.dina(w_G251_2[2]),.dinb(w_n460_0[2]),.dout(n1455),.clk(gclk));
	jand g1154(.dina(w_G248_3[0]),.dinb(w_G234_1[0]),.dout(n1456),.clk(gclk));
	jor g1155(.dina(n1456),.dinb(w_n462_0[0]),.dout(n1457),.clk(gclk));
	jor g1156(.dina(n1457),.dinb(n1455),.dout(n1458),.clk(gclk));
	jand g1157(.dina(w_n366_2[2]),.dinb(w_n460_0[1]),.dout(n1459),.clk(gclk));
	jand g1158(.dina(w_n368_3[0]),.dinb(w_G234_0[2]),.dout(n1460),.clk(gclk));
	jor g1159(.dina(n1460),.dinb(w_G435_0[1]),.dout(n1461),.clk(gclk));
	jor g1160(.dina(n1461),.dinb(w_dff_B_gleghccY1_1),.dout(n1462),.clk(gclk));
	jand g1161(.dina(n1462),.dinb(w_dff_B_cQGu051n7_1),.dout(n1463),.clk(gclk));
	jor g1162(.dina(w_n402_1[1]),.dinb(w_G226_1[0]),.dout(n1464),.clk(gclk));
	jor g1163(.dina(w_n405_1[1]),.dinb(w_n530_0[2]),.dout(n1465),.clk(gclk));
	jand g1164(.dina(n1465),.dinb(w_G422_0[2]),.dout(n1466),.clk(gclk));
	jand g1165(.dina(n1466),.dinb(w_dff_B_bhkwObJ23_1),.dout(n1467),.clk(gclk));
	jor g1166(.dina(w_G254_1[0]),.dinb(w_G226_0[2]),.dout(n1468),.clk(gclk));
	jor g1167(.dina(w_G242_1[0]),.dinb(w_n530_0[1]),.dout(n1469),.clk(gclk));
	jand g1168(.dina(n1469),.dinb(w_n532_0[0]),.dout(n1470),.clk(gclk));
	jand g1169(.dina(n1470),.dinb(w_dff_B_ObJKJAL65_1),.dout(n1471),.clk(gclk));
	jor g1170(.dina(n1471),.dinb(n1467),.dout(n1472),.clk(gclk));
	jxor g1171(.dina(n1472),.dinb(w_n528_0[0]),.dout(n1473),.clk(gclk));
	jor g1172(.dina(w_n402_1[0]),.dinb(w_G218_1[0]),.dout(n1474),.clk(gclk));
	jor g1173(.dina(w_n405_1[0]),.dinb(w_n507_0[2]),.dout(n1475),.clk(gclk));
	jand g1174(.dina(n1475),.dinb(w_G468_0[1]),.dout(n1476),.clk(gclk));
	jand g1175(.dina(n1476),.dinb(w_dff_B_nEin9Box4_1),.dout(n1477),.clk(gclk));
	jor g1176(.dina(w_G254_0[2]),.dinb(w_G218_0[2]),.dout(n1478),.clk(gclk));
	jor g1177(.dina(w_G242_0[2]),.dinb(w_n507_0[1]),.dout(n1479),.clk(gclk));
	jand g1178(.dina(n1479),.dinb(w_n509_0[0]),.dout(n1480),.clk(gclk));
	jand g1179(.dina(n1480),.dinb(w_dff_B_ft2Gh3C70_1),.dout(n1481),.clk(gclk));
	jor g1180(.dina(n1481),.dinb(n1477),.dout(n1482),.clk(gclk));
	jand g1181(.dina(w_G251_2[1]),.dinb(w_n541_0[2]),.dout(n1483),.clk(gclk));
	jand g1182(.dina(w_G248_2[2]),.dinb(w_G210_1[0]),.dout(n1484),.clk(gclk));
	jor g1183(.dina(n1484),.dinb(w_n543_0[0]),.dout(n1485),.clk(gclk));
	jor g1184(.dina(n1485),.dinb(n1483),.dout(n1486),.clk(gclk));
	jand g1185(.dina(w_n366_2[1]),.dinb(w_n541_0[1]),.dout(n1487),.clk(gclk));
	jand g1186(.dina(w_n368_2[2]),.dinb(w_G210_0[2]),.dout(n1488),.clk(gclk));
	jor g1187(.dina(n1488),.dinb(w_G457_0[2]),.dout(n1489),.clk(gclk));
	jor g1188(.dina(n1489),.dinb(w_dff_B_Dbht9dBE8_1),.dout(n1490),.clk(gclk));
	jand g1189(.dina(n1490),.dinb(w_dff_B_9WJTBuJM3_1),.dout(n1491),.clk(gclk));
	jxor g1190(.dina(n1491),.dinb(n1482),.dout(n1492),.clk(gclk));
	jxor g1191(.dina(n1492),.dinb(n1473),.dout(n1493),.clk(gclk));
	jxor g1192(.dina(n1493),.dinb(w_dff_B_RzIglBOu5_1),.dout(n1494),.clk(gclk));
	jand g1193(.dina(w_n495_0[2]),.dinb(w_G251_2[0]),.dout(n1495),.clk(gclk));
	jand g1194(.dina(w_G281_1[0]),.dinb(w_G248_2[1]),.dout(n1496),.clk(gclk));
	jor g1195(.dina(n1496),.dinb(w_n497_0[1]),.dout(n1497),.clk(gclk));
	jor g1196(.dina(n1497),.dinb(n1495),.dout(n1498),.clk(gclk));
	jand g1197(.dina(w_n495_0[1]),.dinb(w_n366_2[0]),.dout(n1499),.clk(gclk));
	jand g1198(.dina(w_G281_0[2]),.dinb(w_n368_2[1]),.dout(n1500),.clk(gclk));
	jor g1199(.dina(n1500),.dinb(w_G374_0[0]),.dout(n1501),.clk(gclk));
	jor g1200(.dina(n1501),.dinb(w_dff_B_0XVfhXz86_1),.dout(n1502),.clk(gclk));
	jand g1201(.dina(n1502),.dinb(w_dff_B_TnDCwe8l9_1),.dout(n1503),.clk(gclk));
	jand g1202(.dina(w_n449_0[2]),.dinb(w_G251_1[2]),.dout(n1504),.clk(gclk));
	jand g1203(.dina(w_G265_1[0]),.dinb(w_G248_2[0]),.dout(n1505),.clk(gclk));
	jor g1204(.dina(n1505),.dinb(w_n451_0[1]),.dout(n1506),.clk(gclk));
	jor g1205(.dina(n1506),.dinb(n1504),.dout(n1507),.clk(gclk));
	jand g1206(.dina(w_n449_0[1]),.dinb(w_n366_1[2]),.dout(n1508),.clk(gclk));
	jand g1207(.dina(w_G265_0[2]),.dinb(w_n368_2[0]),.dout(n1509),.clk(gclk));
	jor g1208(.dina(n1509),.dinb(w_G400_0[1]),.dout(n1510),.clk(gclk));
	jor g1209(.dina(n1510),.dinb(w_dff_B_MuDZpq9d7_1),.dout(n1511),.clk(gclk));
	jand g1210(.dina(n1511),.dinb(w_dff_B_FBmqfDmr8_1),.dout(n1512),.clk(gclk));
	jxor g1211(.dina(n1512),.dinb(n1503),.dout(n1513),.clk(gclk));
	jor g1212(.dina(w_G257_1[0]),.dinb(w_n402_0[2]),.dout(n1514),.clk(gclk));
	jor g1213(.dina(w_n471_0[2]),.dinb(w_n405_0[2]),.dout(n1515),.clk(gclk));
	jand g1214(.dina(n1515),.dinb(w_G389_0[0]),.dout(n1516),.clk(gclk));
	jand g1215(.dina(n1516),.dinb(w_dff_B_hmWGLqJC7_1),.dout(n1517),.clk(gclk));
	jor g1216(.dina(w_G257_0[2]),.dinb(w_G254_0[1]),.dout(n1518),.clk(gclk));
	jor g1217(.dina(w_n471_0[1]),.dinb(w_G242_0[1]),.dout(n1519),.clk(gclk));
	jand g1218(.dina(n1519),.dinb(w_n473_0[1]),.dout(n1520),.clk(gclk));
	jand g1219(.dina(n1520),.dinb(w_dff_B_acLe9BB14_1),.dout(n1521),.clk(gclk));
	jor g1220(.dina(n1521),.dinb(n1517),.dout(n1522),.clk(gclk));
	jand g1221(.dina(w_n484_0[2]),.dinb(w_G251_1[1]),.dout(n1523),.clk(gclk));
	jand g1222(.dina(w_G273_1[0]),.dinb(w_G248_1[2]),.dout(n1524),.clk(gclk));
	jor g1223(.dina(n1524),.dinb(w_n486_0[1]),.dout(n1525),.clk(gclk));
	jor g1224(.dina(n1525),.dinb(n1523),.dout(n1526),.clk(gclk));
	jand g1225(.dina(w_n484_0[1]),.dinb(w_n366_1[1]),.dout(n1527),.clk(gclk));
	jand g1226(.dina(w_G273_0[2]),.dinb(w_n368_1[2]),.dout(n1528),.clk(gclk));
	jor g1227(.dina(n1528),.dinb(w_G411_0[0]),.dout(n1529),.clk(gclk));
	jor g1228(.dina(n1529),.dinb(w_dff_B_9VCie3KC0_1),.dout(n1530),.clk(gclk));
	jand g1229(.dina(n1530),.dinb(w_dff_B_ypoCYK9M4_1),.dout(n1531),.clk(gclk));
	jxor g1230(.dina(n1531),.dinb(n1522),.dout(n1532),.clk(gclk));
	jxor g1231(.dina(n1532),.dinb(n1513),.dout(n1533),.clk(gclk));
	jand g1232(.dina(w_n1533_0[1]),.dinb(w_n1494_0[1]),.dout(n1534),.clk(gclk));
	jnot g1233(.din(n1534),.dout(n1535),.clk(gclk));
	jor g1234(.dina(w_n1533_0[0]),.dinb(w_n1494_0[0]),.dout(n1536),.clk(gclk));
	jand g1235(.dina(n1536),.dinb(w_n750_0[2]),.dout(n1537),.clk(gclk));
	jand g1236(.dina(n1537),.dinb(n1535),.dout(n1538),.clk(gclk));
	jor g1237(.dina(n1454),.dinb(w_n746_0[1]),.dout(n1539),.clk(gclk));
	jor g1238(.dina(n1538),.dinb(w_G4092_1[0]),.dout(n1540),.clk(gclk));
	jxor g1239(.dina(w_n583_0[1]),.dinb(w_n578_0[0]),.dout(n1541),.clk(gclk));
	jxor g1240(.dina(n1541),.dinb(w_n943_0[0]),.dout(n1542),.clk(gclk));
	jnot g1241(.din(n1542),.dout(n1543),.clk(gclk));
	jand g1242(.dina(w_n587_0[2]),.dinb(w_G1497_0[2]),.dout(n1544),.clk(gclk));
	jor g1243(.dina(w_dff_B_LWCDxLKe9_0),.dinb(w_n696_0[0]),.dout(n1545),.clk(gclk));
	jnot g1244(.din(w_n1545_0[1]),.dout(n1546),.clk(gclk));
	jor g1245(.dina(w_n944_0[0]),.dinb(w_n930_0[1]),.dout(n1547),.clk(gclk));
	jand g1246(.dina(n1547),.dinb(w_n706_0[0]),.dout(n1548),.clk(gclk));
	jxor g1247(.dina(n1548),.dinb(w_n928_0[0]),.dout(n1549),.clk(gclk));
	jxor g1248(.dina(w_n605_1[1]),.dinb(w_n948_0[1]),.dout(n1550),.clk(gclk));
	jxor g1249(.dina(w_dff_B_F6fTFBFL8_0),.dinb(n1549),.dout(n1551),.clk(gclk));
	jand g1250(.dina(w_dff_B_ulmeB7oI0_0),.dinb(n1546),.dout(n1552),.clk(gclk));
	jxor g1251(.dina(w_n605_1[0]),.dinb(w_n703_0[0]),.dout(n1553),.clk(gclk));
	jand g1252(.dina(w_n605_0[2]),.dinb(w_n948_0[0]),.dout(n1554),.clk(gclk));
	jor g1253(.dina(n1554),.dinb(w_n702_0[0]),.dout(n1555),.clk(gclk));
	jnot g1254(.din(w_n1555_0[1]),.dout(n1556),.clk(gclk));
	jor g1255(.dina(n1556),.dinb(w_n930_0[0]),.dout(n1557),.clk(gclk));
	jor g1256(.dina(w_n1555_0[0]),.dinb(w_n707_0[0]),.dout(n1558),.clk(gclk));
	jand g1257(.dina(n1558),.dinb(w_dff_B_2c3jPkB65_1),.dout(n1559),.clk(gclk));
	jxor g1258(.dina(n1559),.dinb(w_n596_0[0]),.dout(n1560),.clk(gclk));
	jand g1259(.dina(w_n1560_0[1]),.dinb(w_n1553_0[1]),.dout(n1561),.clk(gclk));
	jnot g1260(.din(n1561),.dout(n1562),.clk(gclk));
	jor g1261(.dina(w_n1560_0[0]),.dinb(w_n1553_0[0]),.dout(n1563),.clk(gclk));
	jand g1262(.dina(w_dff_B_R3AsyGgd0_0),.dinb(w_n1545_0[0]),.dout(n1564),.clk(gclk));
	jand g1263(.dina(n1564),.dinb(w_dff_B_Aqgco1yP8_1),.dout(n1565),.clk(gclk));
	jor g1264(.dina(n1565),.dinb(n1552),.dout(n1566),.clk(gclk));
	jnot g1265(.din(w_G1497_0[1]),.dout(n1567),.clk(gclk));
	jand g1266(.dina(w_n682_0[0]),.dinb(w_n687_0[0]),.dout(n1568),.clk(gclk));
	jand g1267(.dina(w_n1568_0[1]),.dinb(w_n574_0[0]),.dout(n1569),.clk(gclk));
	jxor g1268(.dina(n1569),.dinb(w_n561_0[1]),.dout(n1570),.clk(gclk));
	jxor g1269(.dina(w_n572_0[1]),.dinb(w_n681_1[1]),.dout(n1571),.clk(gclk));
	jor g1270(.dina(w_n856_0[0]),.dinb(w_n853_0[0]),.dout(n1572),.clk(gclk));
	jand g1271(.dina(w_n693_0[1]),.dinb(w_n585_0[0]),.dout(n1573),.clk(gclk));
	jor g1272(.dina(n1573),.dinb(w_n855_0[0]),.dout(n1574),.clk(gclk));
	jand g1273(.dina(n1574),.dinb(n1572),.dout(n1575),.clk(gclk));
	jxor g1274(.dina(n1575),.dinb(w_dff_B_To8vsBxy8_1),.dout(n1576),.clk(gclk));
	jxor g1275(.dina(n1576),.dinb(w_dff_B_CdlBZLKv8_1),.dout(n1577),.clk(gclk));
	jor g1276(.dina(n1577),.dinb(w_dff_B_wBB2siGO4_1),.dout(n1578),.clk(gclk));
	jxor g1277(.dina(w_n693_0[0]),.dinb(w_n572_0[0]),.dout(n1579),.clk(gclk));
	jor g1278(.dina(w_n857_0[0]),.dinb(w_n681_1[0]),.dout(n1580),.clk(gclk));
	jnot g1279(.din(w_n681_0[2]),.dout(n1581),.clk(gclk));
	jor g1280(.dina(w_n680_0[0]),.dinb(n1581),.dout(n1582),.clk(gclk));
	jor g1281(.dina(n1582),.dinb(w_n689_0[0]),.dout(n1583),.clk(gclk));
	jxor g1282(.dina(n1583),.dinb(w_n567_0[1]),.dout(n1584),.clk(gclk));
	jand g1283(.dina(w_dff_B_I3DZOT0N9_0),.dinb(n1580),.dout(n1585),.clk(gclk));
	jxor g1284(.dina(w_n1568_0[0]),.dinb(w_n561_0[0]),.dout(n1586),.clk(gclk));
	jxor g1285(.dina(w_dff_B_0qPXDqtW9_0),.dinb(n1585),.dout(n1587),.clk(gclk));
	jxor g1286(.dina(n1587),.dinb(w_dff_B_nhICFsvk8_1),.dout(n1588),.clk(gclk));
	jor g1287(.dina(n1588),.dinb(w_G1497_0[0]),.dout(n1589),.clk(gclk));
	jand g1288(.dina(w_dff_B_5sQTU8zG9_0),.dinb(n1578),.dout(n1590),.clk(gclk));
	jxor g1289(.dina(n1590),.dinb(n1566),.dout(n1591),.clk(gclk));
	jand g1290(.dina(w_n1591_0[1]),.dinb(w_n1543_0[1]),.dout(n1592),.clk(gclk));
	jnot g1291(.din(n1592),.dout(n1593),.clk(gclk));
	jor g1292(.dina(w_n1591_0[0]),.dinb(w_n1543_0[0]),.dout(n1594),.clk(gclk));
	jand g1293(.dina(n1594),.dinb(w_G4091_0[2]),.dout(n1595),.clk(gclk));
	jand g1294(.dina(n1595),.dinb(n1593),.dout(n1596),.clk(gclk));
	jor g1295(.dina(n1596),.dinb(w_dff_B_KSw97FQY9_1),.dout(n1597),.clk(gclk));
	jand g1296(.dina(w_n1597_0[1]),.dinb(w_dff_B_IIdqX6mj8_1),.dout(w_dff_A_fExTKHZC7_2),.clk(gclk));
	jand g1297(.dina(w_G4092_0[2]),.dinb(G97),.dout(n1599),.clk(gclk));
	jnot g1298(.din(n1599),.dout(n1600),.clk(gclk));
	jand g1299(.dina(w_dff_B_88vVCwdc4_0),.dinb(w_n1597_0[0]),.dout(n1601),.clk(gclk));
	jnot g1300(.din(w_n1601_0[2]),.dout(n1602),.clk(gclk));
	jand g1301(.dina(w_n1602_0[1]),.dinb(w_n793_1[1]),.dout(n1603),.clk(gclk));
	jnot g1302(.din(w_n1447_0[0]),.dout(n1604),.clk(gclk));
	jand g1303(.dina(w_n1446_0[0]),.dinb(w_n1410_0[0]),.dout(n1605),.clk(gclk));
	jor g1304(.dina(n1605),.dinb(w_n750_0[1]),.dout(n1606),.clk(gclk));
	jor g1305(.dina(n1606),.dinb(n1604),.dout(n1607),.clk(gclk));
	jand g1306(.dina(n1607),.dinb(w_n1391_0[0]),.dout(n1608),.clk(gclk));
	jand g1307(.dina(w_G4092_0[1]),.dinb(G94),.dout(n1609),.clk(gclk));
	jor g1308(.dina(w_n1609_0[1]),.dinb(n1608),.dout(n1610),.clk(gclk));
	jand g1309(.dina(w_n1610_0[1]),.dinb(w_n797_1[1]),.dout(n1611),.clk(gclk));
	jand g1310(.dina(w_n799_1[1]),.dinb(w_G14_0[1]),.dout(n1612),.clk(gclk));
	jand g1311(.dina(w_n801_1[1]),.dinb(w_G64_0[1]),.dout(n1613),.clk(gclk));
	jor g1312(.dina(w_dff_B_kA3QnmlP5_0),.dinb(n1612),.dout(n1614),.clk(gclk));
	jor g1313(.dina(w_dff_B_FstWOxMJ7_0),.dinb(n1611),.dout(n1615),.clk(gclk));
	jor g1314(.dina(n1615),.dinb(n1603),.dout(w_dff_A_1182Ow2c0_2),.clk(gclk));
	jand g1315(.dina(w_n1602_0[0]),.dinb(w_n840_1[1]),.dout(n1617),.clk(gclk));
	jand g1316(.dina(w_n1610_0[0]),.dinb(w_n843_1[1]),.dout(n1618),.clk(gclk));
	jand g1317(.dina(w_n845_1[1]),.dinb(w_G14_0[0]),.dout(n1619),.clk(gclk));
	jand g1318(.dina(w_n847_1[1]),.dinb(w_G64_0[0]),.dout(n1620),.clk(gclk));
	jor g1319(.dina(w_dff_B_1tJj2pw78_0),.dinb(n1619),.dout(n1621),.clk(gclk));
	jor g1320(.dina(w_dff_B_UYe82NPj3_0),.dinb(n1618),.dout(n1622),.clk(gclk));
	jor g1321(.dina(n1622),.dinb(n1617),.dout(w_dff_A_GtGQe1WM9_2),.clk(gclk));
	jnot g1322(.din(w_G137_3[1]),.dout(n1624),.clk(gclk));
	jnot g1323(.din(w_n985_1[1]),.dout(n1625),.clk(gclk));
	jor g1324(.dina(w_n1601_0[1]),.dinb(w_dff_B_uSrom04Y5_1),.dout(n1626),.clk(gclk));
	jnot g1325(.din(w_n988_1[1]),.dout(n1627),.clk(gclk));
	jnot g1326(.din(w_n1609_0[0]),.dout(n1628),.clk(gclk));
	jand g1327(.dina(w_dff_B_MRWuuE6D0_0),.dinb(w_n1452_0[0]),.dout(n1629),.clk(gclk));
	jor g1328(.dina(w_n1629_0[1]),.dinb(w_dff_B_q3Yf7HM58_1),.dout(n1630),.clk(gclk));
	jnot g1329(.din(G179),.dout(n1631),.clk(gclk));
	jnot g1330(.din(w_n992_1[1]),.dout(n1632),.clk(gclk));
	jor g1331(.dina(n1632),.dinb(w_n1631_0[1]),.dout(n1633),.clk(gclk));
	jnot g1332(.din(G176),.dout(n1634),.clk(gclk));
	jnot g1333(.din(w_n990_1[1]),.dout(n1635),.clk(gclk));
	jor g1334(.dina(n1635),.dinb(w_n1634_0[1]),.dout(n1636),.clk(gclk));
	jand g1335(.dina(n1636),.dinb(w_dff_B_QBM2HGO14_1),.dout(n1637),.clk(gclk));
	jand g1336(.dina(w_dff_B_NEceM8xN0_0),.dinb(n1630),.dout(n1638),.clk(gclk));
	jand g1337(.dina(n1638),.dinb(w_dff_B_xA0vYSin2_1),.dout(n1639),.clk(gclk));
	jor g1338(.dina(n1639),.dinb(w_n1624_0[1]),.dout(G658),.clk(gclk));
	jnot g1339(.din(w_n999_1[1]),.dout(n1641),.clk(gclk));
	jor g1340(.dina(w_n1601_0[0]),.dinb(w_dff_B_n3cs1FfX4_1),.dout(n1642),.clk(gclk));
	jnot g1341(.din(w_n1002_1[1]),.dout(n1643),.clk(gclk));
	jor g1342(.dina(w_n1629_0[0]),.dinb(w_dff_B_dX64z8cV0_1),.dout(n1644),.clk(gclk));
	jnot g1343(.din(w_n1006_1[1]),.dout(n1645),.clk(gclk));
	jor g1344(.dina(n1645),.dinb(w_n1631_0[0]),.dout(n1646),.clk(gclk));
	jnot g1345(.din(w_n1004_1[1]),.dout(n1647),.clk(gclk));
	jor g1346(.dina(n1647),.dinb(w_n1634_0[0]),.dout(n1648),.clk(gclk));
	jand g1347(.dina(n1648),.dinb(w_dff_B_bVOuko2y1_1),.dout(n1649),.clk(gclk));
	jand g1348(.dina(w_dff_B_CGcUBzOR8_0),.dinb(n1644),.dout(n1650),.clk(gclk));
	jand g1349(.dina(n1650),.dinb(w_dff_B_BsnuMHo72_1),.dout(n1651),.clk(gclk));
	jor g1350(.dina(n1651),.dinb(w_n1624_0[0]),.dout(G690),.clk(gclk));
	buf g1351(.din(w_G141_1[0]),.dout(w_dff_A_EBC8N9T79_1));
	buf g1352(.din(w_G293_0[0]),.dout(w_dff_A_kk7cd6j65_1));
	buf g1353(.din(w_G3173_0[0]),.dout(w_dff_A_a27FDOlD2_1));
	jnot g1354(.din(w_G545_0[1]),.dout(w_dff_A_psklSFAO5_1),.clk(gclk));
	jnot g1355(.din(w_G545_0[0]),.dout(w_dff_A_TwNsD2rL2_1),.clk(gclk));
	buf g1356(.din(w_G137_3[0]),.dout(w_dff_A_2BQXXCY79_1));
	buf g1357(.din(w_G141_0[2]),.dout(w_dff_A_RJ7IrVGd3_1));
	buf g1358(.din(w_G1_2[0]),.dout(w_dff_A_88VaWVqO6_1));
	buf g1359(.din(w_G549_0[1]),.dout(w_dff_A_QSbbVJ567_1));
	buf g1360(.din(w_G299_0[1]),.dout(w_dff_A_QFHYc7Fj1_1));
	jnot g1361(.din(w_G549_0[0]),.dout(w_dff_A_0OPq6GU27_1),.clk(gclk));
	buf g1362(.din(w_G1_1[2]),.dout(w_dff_A_uN1e9ym35_1));
	buf g1363(.din(w_G1_1[1]),.dout(w_dff_A_NnNpN7LE0_1));
	buf g1364(.din(w_G1_1[0]),.dout(w_dff_A_2LtSmUnw2_1));
	buf g1365(.din(w_G1_0[2]),.dout(w_dff_A_bhCkHx8o1_1));
	buf g1366(.din(w_G299_0[0]),.dout(w_dff_A_RvDEgF9N8_1));
	jor g1367(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(w_dff_A_aInYLOFA7_2),.clk(gclk));
	jand g1368(.dina(w_n652_0[0]),.dinb(w_n633_0[1]),.dout(w_dff_A_WZtzsak76_2),.clk(gclk));
	jand g1369(.dina(w_n607_0[0]),.dinb(w_n587_0[1]),.dout(w_dff_A_aqgWgVCw7_2),.clk(gclk));
	jor g1370(.dina(w_n709_0[0]),.dinb(w_n697_0[0]),.dout(w_dff_A_yfLRIfqS6_2),.clk(gclk));
	jor g1371(.dina(w_n742_0[0]),.dinb(w_n733_0[0]),.dout(w_dff_A_pW3zWuB61_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_dff_A_R0DOJt8p2_1),.doutc(w_G4_0[2]),.din(w_dff_B_gvIUJVje8_3));
	jspl jspl_w_G4_1(.douta(w_dff_A_o1Ltpy1M8_0),.doutb(w_G4_1[1]),.din(w_G4_0[0]));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(w_dff_B_TTi3HKcw0_2));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(w_dff_B_DbS2HEhc5_2));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(w_dff_B_K4uE6dlT7_2));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(w_dff_B_ZKONFJX52_2));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(w_dff_B_0QNOVFad6_2));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(w_dff_B_9XFcTKAY6_2));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(w_dff_B_lWeXAT4l1_2));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(w_dff_B_agihHWfT0_2));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(w_dff_B_LY7NLxU77_2));
	jspl jspl_w_G54_0(.douta(w_dff_A_TBOZGujq2_0),.doutb(w_G54_0[1]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(w_dff_B_4HhBeV5W9_2));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(w_dff_B_CPdioXsj6_2));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(w_dff_B_IHXTYMqa1_2));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(w_dff_B_P4yay9r89_2));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(w_dff_B_xqM8Xbir9_2));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(w_dff_B_mBRbiigd7_2));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(w_dff_B_daimAzmN6_2));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(w_dff_B_o5pLiG8c7_2));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(w_dff_B_fJylF7gT3_2));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(w_dff_B_UeAhgxOY3_2));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(w_dff_B_KBen70oB1_2));
	jspl jspl_w_G123_0(.douta(w_dff_A_hzg3IKyz0_0),.doutb(w_G123_0[1]),.din(w_dff_B_HPz1yzyw0_2));
	jspl jspl_w_G132_0(.douta(w_dff_A_KPZKUBKl8_0),.doutb(w_G132_0[1]),.din(w_dff_B_nD7b9jDc3_2));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_w46tlnWm0_0),.doutb(w_dff_A_ZmlcfrZO8_1),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_vkKShGM35_0),.doutb(w_dff_A_pomlwqel7_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_inyEzEyT3_0),.doutb(w_dff_A_e7EX4hop8_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_dff_A_vbqnXyDv5_2),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_dff_A_FvGkOaCi3_0),.doutb(w_dff_A_SL2CkCQG0_1),.doutc(w_G137_4[2]),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_dff_A_Q5iQULE34_0),.doutb(w_G137_5[1]),.doutc(w_G137_5[2]),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_PNqV6Qcx1_0),.doutb(w_dff_A_pQ3EGlQh9_1),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_D0fzhUMk0_1),.doutc(w_dff_A_QB56rGgY4_2),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_dff_A_bwDk8wJS5_0),.doutb(w_G137_8[1]),.doutc(w_dff_A_c68Gy7OQ3_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_G137_9[0]),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_Z5MG9Uvi3_1),.doutc(w_dff_A_Ot0zYzPB2_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_4jl8JVpv6_0),.doutb(w_dff_A_7QRzfq9F4_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(w_dff_B_6WCAemJ45_2));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(w_dff_B_fm02c33D4_2));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(w_dff_B_dOJaaTYT1_2));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(w_dff_B_dOY9Sgmb6_2));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(w_dff_B_Zkwko78p2_2));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(w_dff_B_xSQVsPoZ2_2));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(w_dff_B_CxepozI67_2));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(w_dff_B_EOzGzui27_2));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(w_dff_B_qpVakveK0_2));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(w_dff_B_Y9eZYFbZ9_2));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(w_dff_B_3lqw6BQP3_2));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(w_dff_B_TYlxeCwP3_2));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(w_dff_B_9HPAWxIL1_2));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(w_dff_B_58usAc7i4_2));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(w_dff_B_lvXXY4k86_2));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(w_dff_B_SKbHMiPW2_2));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(w_dff_B_6uRl87Y29_2));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(w_dff_B_hUr9Tjjk0_2));
	jspl3 jspl3_w_G206_0(.douta(w_dff_A_Iri93B0L9_0),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_dff_A_UBKQ6Prb5_2),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_dff_A_EizV1JxL4_1),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl3 jspl3_w_G210_2(.douta(w_G210_2[0]),.doutb(w_dff_A_TRyHePPu3_1),.doutc(w_G210_2[2]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_dff_A_7sPGyeUk4_0),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl3 jspl3_w_G218_2(.douta(w_G218_2[0]),.doutb(w_dff_A_5rnoyF4a9_1),.doutc(w_G218_2[2]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_G226_0[2]),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_dff_A_UIM1XxVP6_0),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G226_2(.douta(w_G226_2[0]),.doutb(w_dff_A_uazgisl77_1),.doutc(w_G226_2[2]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_dff_A_xxiY3hzF4_2),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_dff_A_kc6Gp8Ba3_0),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_dff_A_cJfO8GK75_1),.doutc(w_dff_A_hCUj84rT2_2),.din(G242));
	jspl3 jspl3_w_G242_1(.douta(w_dff_A_WP939Db63_0),.doutb(w_dff_A_m8xX8rCk2_1),.doutc(w_G242_1[2]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_G245_0[0]),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_dff_A_DcYzTp8C6_2),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl jspl_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_dff_A_KEFDYI724_1),.doutc(w_dff_A_UWfb0VmV7_2),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_G251_1[0]),.doutb(w_dff_A_oh0mZN6n0_1),.doutc(w_dff_A_UvE4980e5_2),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_dff_A_FkEO5EKi9_1),.doutc(w_dff_A_8ErAXYhy7_2),.din(w_G251_1[0]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl3 jspl3_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.doutc(w_G254_1[2]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_G257_0[2]),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_WQTppcFP4_0),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G257_2(.douta(w_G257_2[0]),.doutb(w_dff_A_AHWfAdJj2_1),.doutc(w_G257_2[2]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_dff_A_VmEvoykn8_2),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_G265_1[1]),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl jspl_w_G265_2(.douta(w_dff_A_Nvzu5XCg3_0),.doutb(w_G265_2[1]),.din(w_G265_0[1]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_dff_A_LzTv22fS0_2),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_G273_1[1]),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl3 jspl3_w_G273_2(.douta(w_G273_2[0]),.doutb(w_dff_A_k47UJfMu3_1),.doutc(w_G273_2[2]),.din(w_G273_0[1]));
	jspl jspl_w_G280_0(.douta(w_G280_0[0]),.doutb(w_dff_A_m1AaSk9P7_1),.din(G280));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_dff_A_i4yijk0O8_2),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_dff_A_5f3YffZc9_0),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_dff_A_4T8SEnOh4_0),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_dff_A_e4wCn9PN4_1),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_dff_A_W0RigKhz8_0),.doutb(w_dff_A_CapWvRY64_1),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_dff_A_dltZK1Z17_0),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_G316_0[2]),.din(G316));
	jspl3 jspl3_w_G316_1(.douta(w_dff_A_uICwoGZT6_0),.doutb(w_G316_1[1]),.doutc(w_G316_1[2]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_dff_A_2Z0K9zBT8_1),.doutc(w_G324_0[2]),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_dff_A_Pix1T5Ii7_1),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_dff_A_Q2Ystg7B1_1),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_G332_1[1]),.doutc(w_dff_A_iJNkOBcs6_2),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_dff_A_22LW2eOR1_0),.doutb(w_G332_2[1]),.doutc(w_G332_2[2]),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_dff_A_jbpgR47I0_0),.doutb(w_G332_3[1]),.doutc(w_dff_A_6hgNxPZ11_2),.din(w_G332_0[2]));
	jspl3 jspl3_w_G332_4(.douta(w_dff_A_wdTD53Z07_0),.doutb(w_G332_4[1]),.doutc(w_G332_4[2]),.din(w_G332_1[0]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl3 jspl3_w_G335_1(.douta(w_G335_1[0]),.doutb(w_G335_1[1]),.doutc(w_dff_A_giWd21D36_2),.din(w_G335_0[0]));
	jspl3 jspl3_w_G335_2(.douta(w_G335_2[0]),.doutb(w_G335_2[1]),.doutc(w_G335_2[2]),.din(w_G335_0[1]));
	jspl3 jspl3_w_G335_3(.douta(w_dff_A_MVqbkzH00_0),.doutb(w_G335_3[1]),.doutc(w_G335_3[2]),.din(w_G335_0[2]));
	jspl jspl_w_G335_4(.douta(w_dff_A_f7lUCiew2_0),.doutb(w_G335_4[1]),.din(w_G335_1[0]));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_dff_A_LHr0g24r7_2),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_dff_A_kjapD70J7_1),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_dff_A_5N4U0R7P9_0),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_G351_0[2]),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_dff_A_fMakeybT3_0),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_dff_A_UjBQH0Zl5_1),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_dff_A_FYFbEOeg7_0),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_dff_A_RkoxuewP3_1),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G369_0(.douta(w_dff_A_OkzrOEWX9_0),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_dff_A_uzHU8Ycj9_0),.doutb(w_dff_A_zxoV718G2_1),.doutc(w_G374_0[2]),.din(G374));
	jspl3 jspl3_w_G389_0(.douta(w_dff_A_8QLBYNJY8_0),.doutb(w_dff_A_emFgZITx2_1),.doutc(w_G389_0[2]),.din(G389));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_dff_A_3gDDM7YM7_1),.doutc(w_dff_A_6TXoc7rK1_2),.din(G400));
	jspl jspl_w_G400_1(.douta(w_dff_A_epP7q5ez9_0),.doutb(w_G400_1[1]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_dff_A_IBV2KcPm6_0),.doutb(w_dff_A_KdrmsbCd1_1),.doutc(w_G411_0[2]),.din(G411));
	jspl3 jspl3_w_G422_0(.douta(w_dff_A_u7SX3Bg06_0),.doutb(w_G422_0[1]),.doutc(w_dff_A_3mpWkusM1_2),.din(G422));
	jspl3 jspl3_w_G422_1(.douta(w_G422_1[0]),.doutb(w_G422_1[1]),.doutc(w_G422_1[2]),.din(w_G422_0[0]));
	jspl jspl_w_G422_2(.douta(w_dff_A_3BiR3btB8_0),.doutb(w_G422_2[1]),.din(w_G422_0[1]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_dff_A_KBCP7C4J6_1),.doutc(w_dff_A_5srVuwcl4_2),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_dff_A_Jgsa7gf44_0),.doutb(w_dff_A_8PTPxEZU2_1),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_dff_A_mw3Zve2w6_1),.doutc(w_dff_A_fLq7odAN5_2),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_dff_A_YeycLRNs9_0),.doutb(w_dff_A_5acy51VL2_1),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_dff_A_sWDiBuh02_0),.doutb(w_G457_0[1]),.doutc(w_dff_A_siA6kNFd3_2),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_G457_1[0]),.doutb(w_G457_1[1]),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl jspl_w_G457_2(.douta(w_dff_A_DSYuGwNq6_0),.doutb(w_G457_2[1]),.din(w_G457_0[1]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_dff_A_gU7880GW8_1),.doutc(w_dff_A_F12oIkZY4_2),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_dff_A_zPwGSvjv5_0),.doutb(w_dff_A_ePZeCHJY0_1),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_G479_0[0]),.doutb(w_dff_A_Pxom4RSw4_1),.doutc(w_dff_A_DFmdfCgD2_2),.din(G479));
	jspl jspl_w_G479_1(.douta(w_dff_A_vcbZ96Yk7_0),.doutb(w_G479_1[1]),.din(w_G479_0[0]));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_dff_A_fwBz1ci64_1),.doutc(w_dff_A_SDo89qRs2_2),.din(G490));
	jspl3 jspl3_w_G490_1(.douta(w_dff_A_IGH3UTH66_0),.doutb(w_dff_A_B9NRc5n21_1),.doutc(w_G490_1[2]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_G503_0[0]),.doutb(w_dff_A_vgOyOihe1_1),.doutc(w_dff_A_pwLbgITt6_2),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_dff_A_Zlou7Hha4_0),.doutb(w_dff_A_0SmFqPbu6_1),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl3 jspl3_w_G514_0(.douta(w_G514_0[0]),.doutb(w_dff_A_qVwVWVcQ5_1),.doutc(w_dff_A_XxixcFjb6_2),.din(G514));
	jspl jspl_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.din(w_G514_0[0]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_dff_A_rfAUD5jN9_1),.doutc(w_dff_A_8rATMYQt0_2),.din(G523));
	jspl jspl_w_G523_1(.douta(w_dff_A_w0Ny0zwc1_0),.doutb(w_G523_1[1]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_G534_0[0]),.doutb(w_dff_A_mVrS8o4v7_1),.doutc(w_dff_A_Lm3Wb03d5_2),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_dff_A_YqbMMSiH2_0),.doutb(w_dff_A_JNMCiPQM9_1),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_G559_0[0]),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_dff_A_QIPZdZ9U2_0),.doutb(w_G1497_0[1]),.doutc(w_dff_A_gmdSfpsv8_2),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_G1689_0[1]),.doutc(w_dff_A_jZQpmhwB0_2),.din(G1689));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_dff_A_TzPdTV922_1),.doutc(w_G1690_0[2]),.din(G1690));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_G1691_0[1]),.doutc(w_dff_A_FgyHJt2a3_2),.din(G1691));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_dff_A_sIWnwDEh7_1),.doutc(w_G1694_0[2]),.din(G1694));
	jspl3 jspl3_w_G2174_0(.douta(w_dff_A_FzmSQcjZ8_0),.doutb(w_G2174_0[1]),.doutc(w_dff_A_TBhpKZhG1_2),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_dff_A_1ORJ7GLS6_0),.doutb(w_dff_A_CMurshcQ6_1),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(w_dff_B_4Q09WIFX4_3));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_dff_A_AcuIn80b5_0),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_dff_A_EXwBExOx4_0),.doutb(w_G3724_0[1]),.doutc(w_dff_A_4fATliDZ0_2),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_dff_A_FTuHRH8f2_1),.doutc(w_G4087_0[2]),.din(G4087));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_dff_A_6ma5F38f2_2),.din(G4088));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_dff_A_uFn2pNSI7_2),.din(G4089));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_dff_A_BadhDM3A4_1),.doutc(w_G4090_0[2]),.din(G4090));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_G4091_0[1]),.doutc(w_dff_A_4XKB28U33_2),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_G4091_1[0]),.doutb(w_dff_A_GBdJ8qxM0_1),.doutc(w_dff_A_U2nEUDmM9_2),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_G4091_2[0]),.doutb(w_G4091_2[1]),.doutc(w_dff_A_HsNOgYfh5_2),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_G4092_0[1]),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_dff_A_I4mWuMdI9_0),.doutb(w_dff_A_X5iFbqWZ6_1),.doutc(w_G4092_1[2]),.din(w_G4092_0[0]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(w_dff_A_Md6sOKZ80_1),.din(G599_fa_));
	jspl jspl_w_G600_0(.douta(w_G600_0),.doutb(w_dff_A_95yRjwe90_1),.din(G600_fa_));
	jspl jspl_w_G601_0(.douta(w_dff_A_hKPwJCt40_0),.doutb(w_dff_A_AtXnEyBC7_1),.din(G601_fa_));
	jspl jspl_w_G611_0(.douta(w_G611_0),.doutb(w_dff_A_g9Y6z9mT9_1),.din(G611_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(w_dff_A_wMjzKV3T2_1),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_G809_1[0]),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_G809_2[2]),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_G809_3[0]),.doutb(w_G809_3[1]),.doutc(w_dff_A_4FDeHSQK4_2),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(w_dff_A_T8dVu50g8_1),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(w_dff_A_St9eEOx71_1),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(w_dff_A_YdqD4BPM6_1),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(w_dff_A_CnsGiYrK3_1),.din(G861_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(w_dff_A_ZffOHOwP8_1),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(w_dff_A_msTcj59W3_1),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(w_dff_A_DncwKVdg0_1),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(w_dff_A_IXVtm8zU8_1),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(w_dff_A_NIZhYMSx1_1),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(w_dff_A_wxyThvto1_1),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(w_dff_A_y2fvlRfV5_1),.din(G877_fa_));
	jspl jspl_w_G1000_0(.douta(w_G1000_0),.doutb(w_dff_A_yV3M3vWw4_1),.din(G1000_fa_));
	jspl jspl_w_G826_0(.douta(w_G826_0),.doutb(w_dff_A_8Pa9YStv0_1),.din(G826_fa_));
	jspl jspl_w_G828_0(.douta(w_G828_0),.doutb(w_dff_A_WWL5M9oO4_1),.din(G828_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(w_dff_A_mLyNlAgr2_1),.din(G830_fa_));
	jspl jspl_w_G867_0(.douta(w_G867_0),.doutb(w_dff_A_yZxRu1CP2_1),.din(G867_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(w_dff_A_3kPjIFex3_1),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(w_dff_B_iIiqK0wI0_2));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_dff_A_xQReP0PA4_0),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n366_2(.douta(w_n366_2[0]),.doutb(w_n366_2[1]),.doutc(w_n366_2[2]),.din(w_n366_0[1]));
	jspl3 jspl3_w_n366_3(.douta(w_n366_3[0]),.doutb(w_n366_3[1]),.doutc(w_n366_3[2]),.din(w_n366_0[2]));
	jspl3 jspl3_w_n366_4(.douta(w_n366_4[0]),.doutb(w_n366_4[1]),.doutc(w_n366_4[2]),.din(w_n366_1[0]));
	jspl3 jspl3_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.doutc(w_n368_0[2]),.din(n368));
	jspl3 jspl3_w_n368_1(.douta(w_n368_1[0]),.doutb(w_n368_1[1]),.doutc(w_n368_1[2]),.din(w_n368_0[0]));
	jspl3 jspl3_w_n368_2(.douta(w_n368_2[0]),.doutb(w_n368_2[1]),.doutc(w_n368_2[2]),.din(w_n368_0[1]));
	jspl3 jspl3_w_n368_3(.douta(w_n368_3[0]),.doutb(w_n368_3[1]),.doutc(w_n368_3[2]),.din(w_n368_0[2]));
	jspl3 jspl3_w_n368_4(.douta(w_n368_4[0]),.doutb(w_n368_4[1]),.doutc(w_n368_4[2]),.din(w_n368_1[0]));
	jspl jspl_w_n368_5(.douta(w_n368_5[0]),.doutb(w_n368_5[1]),.din(w_n368_1[1]));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.doutc(w_n372_0[2]),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl3 jspl3_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.doutc(w_n385_1[2]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n386_1(.douta(w_n386_1[0]),.doutb(w_n386_1[1]),.doutc(w_n386_1[2]),.din(w_n386_0[0]));
	jspl3 jspl3_w_n386_2(.douta(w_n386_2[0]),.doutb(w_n386_2[1]),.doutc(w_n386_2[2]),.din(w_n386_0[1]));
	jspl3 jspl3_w_n386_3(.douta(w_n386_3[0]),.doutb(w_n386_3[1]),.doutc(w_n386_3[2]),.din(w_n386_0[2]));
	jspl3 jspl3_w_n386_4(.douta(w_n386_4[0]),.doutb(w_n386_4[1]),.doutc(w_n386_4[2]),.din(w_n386_1[0]));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_dff_A_oRe2HLmT5_2),.din(w_dff_B_l9V0R11f7_3));
	jspl3 jspl3_w_n388_1(.douta(w_dff_A_AT1Avun83_0),.doutb(w_dff_A_umPSBfAm7_1),.doutc(w_n388_1[2]),.din(w_n388_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_n389_0[2]),.din(n389));
	jspl3 jspl3_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.doutc(w_n389_1[2]),.din(w_n389_0[0]));
	jspl3 jspl3_w_n389_2(.douta(w_n389_2[0]),.doutb(w_n389_2[1]),.doutc(w_n389_2[2]),.din(w_n389_0[1]));
	jspl3 jspl3_w_n389_3(.douta(w_n389_3[0]),.doutb(w_n389_3[1]),.doutc(w_n389_3[2]),.din(w_n389_0[2]));
	jspl3 jspl3_w_n389_4(.douta(w_n389_4[0]),.doutb(w_n389_4[1]),.doutc(w_n389_4[2]),.din(w_n389_1[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_dff_A_dmVkfCCc4_1),.din(n397));
	jspl3 jspl3_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.doutc(w_n398_0[2]),.din(n398));
	jspl3 jspl3_w_n401_0(.douta(w_dff_A_r1l9bUN20_0),.doutb(w_n401_0[1]),.doutc(w_dff_A_fPmmE3xD9_2),.din(n401));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n402_1(.douta(w_n402_1[0]),.doutb(w_n402_1[1]),.doutc(w_n402_1[2]),.din(w_n402_0[0]));
	jspl jspl_w_n402_2(.douta(w_n402_2[0]),.doutb(w_n402_2[1]),.din(w_n402_0[1]));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl3 jspl3_w_n405_1(.douta(w_n405_1[0]),.doutb(w_n405_1[1]),.doutc(w_n405_1[2]),.din(w_n405_0[0]));
	jspl jspl_w_n405_2(.douta(w_n405_2[0]),.doutb(w_n405_2[1]),.din(w_n405_0[1]));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_dff_A_PQWTlDM18_2),.din(n410));
	jspl jspl_w_n410_1(.douta(w_dff_A_15kIWfyz3_0),.doutb(w_n410_1[1]),.din(w_n410_0[0]));
	jspl jspl_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.din(n414));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(n416));
	jspl3 jspl3_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.doutc(w_n419_0[2]),.din(n419));
	jspl3 jspl3_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.doutc(w_n424_0[2]),.din(n424));
	jspl3 jspl3_w_n424_1(.douta(w_n424_1[0]),.doutb(w_n424_1[1]),.doutc(w_n424_1[2]),.din(w_n424_0[0]));
	jspl jspl_w_n424_2(.douta(w_n424_2[0]),.doutb(w_n424_2[1]),.din(w_n424_0[1]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_dff_A_Fn8Bdpbb4_1),.din(n426));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl3 jspl3_w_n437_0(.douta(w_dff_A_yvXDm0ym2_0),.doutb(w_n437_0[1]),.doutc(w_dff_A_mrHgL0da5_2),.din(n437));
	jspl3 jspl3_w_n437_1(.douta(w_dff_A_YUvWpXW59_0),.doutb(w_dff_A_zQPB9WuL5_1),.doutc(w_n437_1[2]),.din(w_n437_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_dff_A_XBsqqt4V8_0),.doutb(w_n451_0[1]),.doutc(w_dff_A_KKnWbrl30_2),.din(n451));
	jspl jspl_w_n451_1(.douta(w_dff_A_quGm9qOq7_0),.doutb(w_n451_1[1]),.din(w_n451_0[0]));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_dff_A_yEEkNlvz4_1),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_3aaz8XkD0_1),.doutc(w_dff_A_4vYs8wAb7_2),.din(n462));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl jspl_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.doutc(w_dff_A_cR87xW9l6_2),.din(w_dff_B_9tSn0Y3k1_3));
	jspl3 jspl3_w_n473_1(.douta(w_dff_A_Rx7my7XR1_0),.doutb(w_dff_A_F72lr6t99_1),.doutc(w_n473_1[2]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.doutc(w_n484_0[2]),.din(n484));
	jspl jspl_w_n484_1(.douta(w_n484_1[0]),.doutb(w_n484_1[1]),.din(w_n484_0[0]));
	jspl3 jspl3_w_n486_0(.douta(w_dff_A_W71XNuJJ0_0),.doutb(w_n486_0[1]),.doutc(w_dff_A_AYrARYnc4_2),.din(n486));
	jspl jspl_w_n486_1(.douta(w_dff_A_OkQ4V4ul0_0),.doutb(w_n486_1[1]),.din(w_n486_0[0]));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl3 jspl3_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.doutc(w_n495_0[2]),.din(n495));
	jspl3 jspl3_w_n495_1(.douta(w_n495_1[0]),.doutb(w_n495_1[1]),.doutc(w_n495_1[2]),.din(w_n495_0[0]));
	jspl3 jspl3_w_n497_0(.douta(w_dff_A_hcaBnGNJ4_0),.doutb(w_n497_0[1]),.doutc(w_dff_A_aL3GOddb6_2),.din(n497));
	jspl jspl_w_n497_1(.douta(w_dff_A_ixbpSxxm4_0),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl jspl_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.din(w_n507_0[0]));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_nQshTVjR8_2));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl jspl_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.doutc(w_n528_0[2]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl jspl_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.din(w_n530_0[0]));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(w_dff_B_VElSIzjE4_2));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl3 jspl3_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.doutc(w_n541_0[2]),.din(n541));
	jspl jspl_w_n541_1(.douta(w_n541_1[0]),.doutb(w_n541_1[1]),.din(w_n541_0[0]));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_dff_A_cjga727m6_1),.din(n543));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl jspl_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl jspl_w_n560_1(.douta(w_n560_1[0]),.doutb(w_n560_1[1]),.din(w_n560_0[0]));
	jspl3 jspl3_w_n561_0(.douta(w_dff_A_Rzp9MT8F9_0),.doutb(w_dff_A_9OAdvTyj2_1),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n562_0(.douta(w_dff_A_0pE0wOE56_0),.doutb(w_n562_0[1]),.din(w_dff_B_Vhp7DYjM5_2));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_dff_A_F5A5MZ505_1),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n567_1(.douta(w_n567_1[0]),.doutb(w_dff_A_rNtdnGCB4_1),.din(w_n567_0[0]));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_dff_A_z8mKH3gn7_1),.din(n569));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_dff_A_gTlyjfpT1_2),.din(n571));
	jspl jspl_w_n571_1(.douta(w_n571_1[0]),.doutb(w_n571_1[1]),.din(w_n571_0[0]));
	jspl3 jspl3_w_n572_0(.douta(w_dff_A_s3a2UhOY3_0),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.doutc(w_n577_0[2]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_dff_A_H8aPmCPQ7_1),.doutc(w_n578_0[2]),.din(n578));
	jspl3 jspl3_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.doutc(w_n582_0[2]),.din(n582));
	jspl jspl_w_n582_1(.douta(w_n582_1[0]),.doutb(w_n582_1[1]),.din(w_n582_0[0]));
	jspl3 jspl3_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.doutc(w_dff_A_legCigtL3_2),.din(n583));
	jspl jspl_w_n583_1(.douta(w_dff_A_rBYzm1ut3_0),.doutb(w_n583_1[1]),.din(w_n583_0[0]));
	jspl jspl_w_n585_0(.douta(w_dff_A_pEJMJpr07_0),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.doutc(w_n587_0[2]),.din(n587));
	jspl jspl_w_n587_1(.douta(w_n587_1[0]),.doutb(w_n587_1[1]),.din(w_n587_0[0]));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_dff_A_BIFyI2Ba4_1),.doutc(w_n590_0[2]),.din(n590));
	jspl jspl_w_n590_1(.douta(w_n590_1[0]),.doutb(w_n590_1[1]),.din(w_n590_0[0]));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_dff_A_2NXqZb9L5_1),.din(n591));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.doutc(w_n595_0[2]),.din(n595));
	jspl jspl_w_n595_1(.douta(w_n595_1[0]),.doutb(w_n595_1[1]),.din(w_n595_0[0]));
	jspl3 jspl3_w_n596_0(.douta(w_dff_A_F0ZZ8ljA9_0),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl3 jspl3_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.doutc(w_n600_0[2]),.din(n600));
	jspl jspl_w_n600_1(.douta(w_n600_1[0]),.doutb(w_n600_1[1]),.din(w_n600_0[0]));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl3 jspl3_w_n604_0(.douta(w_dff_A_MVAVHnvF7_0),.doutb(w_n604_0[1]),.doutc(w_n604_0[2]),.din(n604));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_dff_A_YNBRqcRa7_2),.din(w_n605_0[0]));
	jspl3 jspl3_w_n605_2(.douta(w_n605_2[0]),.doutb(w_n605_2[1]),.doutc(w_n605_2[2]),.din(w_n605_0[1]));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_dff_A_snnl1FyO3_1),.doutc(w_n607_0[2]),.din(w_dff_B_7zdIdKpx6_3));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n609_1(.douta(w_n609_1[0]),.doutb(w_n609_1[1]),.doutc(w_n609_1[2]),.din(w_n609_0[0]));
	jspl3 jspl3_w_n609_2(.douta(w_n609_2[0]),.doutb(w_n609_2[1]),.doutc(w_n609_2[2]),.din(w_n609_0[1]));
	jspl3 jspl3_w_n609_3(.douta(w_n609_3[0]),.doutb(w_n609_3[1]),.doutc(w_n609_3[2]),.din(w_n609_0[2]));
	jspl3 jspl3_w_n609_4(.douta(w_n609_4[0]),.doutb(w_n609_4[1]),.doutc(w_n609_4[2]),.din(w_n609_1[0]));
	jspl3 jspl3_w_n609_5(.douta(w_n609_5[0]),.doutb(w_n609_5[1]),.doutc(w_n609_5[2]),.din(w_n609_1[1]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n614_0(.douta(w_n614_0[0]),.doutb(w_dff_A_uWtMHdEi7_1),.doutc(w_dff_A_dv9qDyKm0_2),.din(n614));
	jspl3 jspl3_w_n614_1(.douta(w_dff_A_pBW3DPRX8_0),.doutb(w_n614_1[1]),.doutc(w_dff_A_LOEMaROP6_2),.din(w_n614_0[0]));
	jspl jspl_w_n614_2(.douta(w_dff_A_pyxSFSNG2_0),.doutb(w_n614_2[1]),.din(w_n614_0[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl jspl_w_n618_1(.douta(w_n618_1[0]),.doutb(w_n618_1[1]),.din(w_n618_0[0]));
	jspl3 jspl3_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.doutc(w_n621_0[2]),.din(n621));
	jspl3 jspl3_w_n621_1(.douta(w_dff_A_ZcjTCanV9_0),.doutb(w_n621_1[1]),.doutc(w_n621_1[2]),.din(w_n621_0[0]));
	jspl jspl_w_n621_2(.douta(w_dff_A_KGO1f1I56_0),.doutb(w_n621_2[1]),.din(w_n621_0[1]));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_n622_0[2]),.din(n622));
	jspl jspl_w_n622_1(.douta(w_n622_1[0]),.doutb(w_n622_1[1]),.din(w_n622_0[0]));
	jspl jspl_w_n623_0(.douta(w_dff_A_P6llDIia8_0),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.doutc(w_n624_0[2]),.din(n624));
	jspl3 jspl3_w_n624_1(.douta(w_n624_1[0]),.doutb(w_n624_1[1]),.doutc(w_n624_1[2]),.din(w_n624_0[0]));
	jspl3 jspl3_w_n625_0(.douta(w_dff_A_h4DbwCpQ5_0),.doutb(w_n625_0[1]),.doutc(w_dff_A_TV5Z6BNA5_2),.din(n625));
	jspl3 jspl3_w_n628_0(.douta(w_n628_0[0]),.doutb(w_dff_A_ieu9LqiI2_1),.doutc(w_n628_0[2]),.din(n628));
	jspl3 jspl3_w_n629_0(.douta(w_n629_0[0]),.doutb(w_dff_A_bAIxOVC57_1),.doutc(w_n629_0[2]),.din(n629));
	jspl jspl_w_n631_0(.douta(w_dff_A_SNSIvQLJ8_0),.doutb(w_n631_0[1]),.din(n631));
	jspl3 jspl3_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.doutc(w_n633_0[2]),.din(n633));
	jspl jspl_w_n633_1(.douta(w_n633_1[0]),.doutb(w_n633_1[1]),.din(w_n633_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_dff_A_K6f1eYEf2_2),.din(n636));
	jspl jspl_w_n636_1(.douta(w_n636_1[0]),.doutb(w_dff_A_ADSSagpo0_1),.din(w_n636_0[0]));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_dff_A_wCzkzTI42_1),.doutc(w_dff_A_SZza9EIx1_2),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_dff_A_4qExMfTp2_0),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.doutc(w_n645_0[2]),.din(n645));
	jspl3 jspl3_w_n646_0(.douta(w_dff_A_XMc8XPuB1_0),.doutb(w_n646_0[1]),.doutc(w_n646_0[2]),.din(n646));
	jspl3 jspl3_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.doutc(w_dff_A_4o8dWzod0_2),.din(n649));
	jspl jspl_w_n649_1(.douta(w_n649_1[0]),.doutb(w_n649_1[1]),.din(w_n649_0[0]));
	jspl jspl_w_n650_0(.douta(w_dff_A_g83TBW6C0_0),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n651_0(.douta(w_n651_0[0]),.doutb(w_dff_A_QrUn5Y1q2_1),.doutc(w_dff_A_SSqurgJA3_2),.din(w_dff_B_5tBr8GmK5_3));
	jspl jspl_w_n651_1(.douta(w_dff_A_bvaE7bz80_0),.doutb(w_n651_1[1]),.din(w_n651_0[0]));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(w_dff_B_mEUW4q3f7_2));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl jspl_w_n671_0(.douta(w_dff_A_eGI5ioL92_0),.doutb(w_n671_0[1]),.din(n671));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_dff_A_AHYVuzOx6_1),.din(n678));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_dff_A_y24sHRf73_1),.din(n679));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_dff_A_Q8688C4e3_1),.din(w_dff_B_n06xFyHa9_2));
	jspl3 jspl3_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.doutc(w_n681_0[2]),.din(n681));
	jspl3 jspl3_w_n681_1(.douta(w_dff_A_Z01nOi0E2_0),.doutb(w_dff_A_xySRvejU7_1),.doutc(w_n681_1[2]),.din(w_n681_0[0]));
	jspl jspl_w_n681_2(.douta(w_dff_A_aNeRiGDk3_0),.doutb(w_n681_2[1]),.din(w_n681_0[1]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl3 jspl3_w_n687_0(.douta(w_dff_A_kGXM6RqT9_0),.doutb(w_dff_A_qDDp2ip11_1),.doutc(w_n687_0[2]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_dff_A_evSASmTu6_0),.doutb(w_n689_0[1]),.din(n689));
	jspl3 jspl3_w_n691_0(.douta(w_n691_0[0]),.doutb(w_dff_A_YAqQIAnL3_1),.doutc(w_n691_0[2]),.din(n691));
	jspl3 jspl3_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.doutc(w_n693_0[2]),.din(n693));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.doutc(w_n696_0[2]),.din(n696));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_dff_A_IMU7GyEl9_1),.din(n700));
	jspl jspl_w_n702_0(.douta(w_n702_0[0]),.doutb(w_n702_0[1]),.din(w_dff_B_8MNPYt2H8_2));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl jspl_w_n706_0(.douta(w_dff_A_Bi2zBv3k9_0),.doutb(w_n706_0[1]),.din(n706));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.doutc(w_n707_0[2]),.din(n707));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(w_dff_B_kq54St0X9_2));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_dff_A_d3P4bKgJ3_1),.doutc(w_dff_A_YVKjARmo8_2),.din(n717));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl3 jspl3_w_n721_0(.douta(w_n721_0[0]),.doutb(w_dff_A_IYre53nc7_1),.doutc(w_n721_0[2]),.din(n721));
	jspl jspl_w_n723_0(.douta(w_dff_A_fMv0x7dt0_0),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl3 jspl3_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.doutc(w_n727_0[2]),.din(n727));
	jspl3 jspl3_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.doutc(w_n729_0[2]),.din(n729));
	jspl jspl_w_n729_1(.douta(w_n729_1[0]),.doutb(w_n729_1[1]),.din(w_n729_0[0]));
	jspl3 jspl3_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.doutc(w_n732_0[2]),.din(n732));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.din(n735));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl3 jspl3_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.doutc(w_dff_A_edJapZXS5_2),.din(n739));
	jspl jspl_w_n739_1(.douta(w_dff_A_mpgmD9Kb4_0),.doutb(w_n739_1[1]),.din(w_n739_0[0]));
	jspl jspl_w_n740_0(.douta(w_n740_0[0]),.doutb(w_dff_A_IA24yFJu7_1),.din(n740));
	jspl jspl_w_n741_0(.douta(w_dff_A_1huJGL037_0),.doutb(w_n741_0[1]),.din(n741));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(w_dff_B_3Mdt917A2_2));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_dff_A_XnJVWyVQ2_2),.din(w_dff_B_792OCErl1_3));
	jspl3 jspl3_w_n744_1(.douta(w_dff_A_3JDVhz4W3_0),.doutb(w_n744_1[1]),.doutc(w_n744_1[2]),.din(w_n744_0[0]));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.doutc(w_dff_A_Hlfz5tLw4_2),.din(n746));
	jspl3 jspl3_w_n746_1(.douta(w_n746_1[0]),.doutb(w_n746_1[1]),.doutc(w_n746_1[2]),.din(w_n746_0[0]));
	jspl3 jspl3_w_n747_0(.douta(w_dff_A_abiRJ84q1_0),.doutb(w_dff_A_xVwWe8BZ7_1),.doutc(w_n747_0[2]),.din(n747));
	jspl3 jspl3_w_n747_1(.douta(w_n747_1[0]),.doutb(w_dff_A_kc7C7W6D4_1),.doutc(w_dff_A_S4pNyZOJ2_2),.din(w_n747_0[0]));
	jspl3 jspl3_w_n747_2(.douta(w_dff_A_69179VsI2_0),.doutb(w_dff_A_Kd60217a3_1),.doutc(w_n747_2[2]),.din(w_n747_0[1]));
	jspl3 jspl3_w_n747_3(.douta(w_dff_A_ZUTBvrie0_0),.doutb(w_dff_A_osacSdo95_1),.doutc(w_n747_3[2]),.din(w_n747_0[2]));
	jspl3 jspl3_w_n748_0(.douta(w_n748_0[0]),.doutb(w_dff_A_zUHE6OJp7_1),.doutc(w_dff_A_zkyVJEDD9_2),.din(w_dff_B_b3QgmtF84_3));
	jspl3 jspl3_w_n748_1(.douta(w_n748_1[0]),.doutb(w_dff_A_LgHOED8V7_1),.doutc(w_dff_A_A5Gq2DXr3_2),.din(w_n748_0[0]));
	jspl3 jspl3_w_n748_2(.douta(w_dff_A_tN7pN9zS4_0),.doutb(w_n748_2[1]),.doutc(w_dff_A_LBlA3ipn0_2),.din(w_n748_0[1]));
	jspl3 jspl3_w_n748_3(.douta(w_n748_3[0]),.doutb(w_dff_A_tiltUMDh0_1),.doutc(w_dff_A_QBdu86M61_2),.din(w_n748_0[2]));
	jspl jspl_w_n748_4(.douta(w_dff_A_TCaFfdVO2_0),.doutb(w_n748_4[1]),.din(w_n748_1[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_dff_A_UfmvrRkC4_1),.doutc(w_dff_A_JuSmpmgD2_2),.din(n750));
	jspl jspl_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n751_0(.douta(w_dff_A_IVzXe4al7_0),.doutb(w_n751_0[1]),.doutc(w_dff_A_8Wcm2ddZ5_2),.din(n751));
	jspl3 jspl3_w_n751_1(.douta(w_n751_1[0]),.doutb(w_dff_A_Oy42UHnV4_1),.doutc(w_n751_1[2]),.din(w_n751_0[0]));
	jspl jspl_w_n751_2(.douta(w_n751_2[0]),.doutb(w_dff_A_JkGZyrSp0_1),.din(w_n751_0[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.doutc(w_n753_0[2]),.din(n753));
	jspl3 jspl3_w_n753_1(.douta(w_n753_1[0]),.doutb(w_n753_1[1]),.doutc(w_n753_1[2]),.din(w_n753_0[0]));
	jspl3 jspl3_w_n753_2(.douta(w_n753_2[0]),.doutb(w_n753_2[1]),.doutc(w_n753_2[2]),.din(w_n753_0[1]));
	jspl3 jspl3_w_n753_3(.douta(w_n753_3[0]),.doutb(w_n753_3[1]),.doutc(w_n753_3[2]),.din(w_n753_0[2]));
	jspl3 jspl3_w_n753_4(.douta(w_n753_4[0]),.doutb(w_n753_4[1]),.doutc(w_n753_4[2]),.din(w_n753_1[0]));
	jspl3 jspl3_w_n753_5(.douta(w_n753_5[0]),.doutb(w_n753_5[1]),.doutc(w_n753_5[2]),.din(w_n753_1[1]));
	jspl3 jspl3_w_n753_6(.douta(w_n753_6[0]),.doutb(w_n753_6[1]),.doutc(w_n753_6[2]),.din(w_n753_1[2]));
	jspl3 jspl3_w_n753_7(.douta(w_n753_7[0]),.doutb(w_n753_7[1]),.doutc(w_n753_7[2]),.din(w_n753_2[0]));
	jspl jspl_w_n753_8(.douta(w_n753_8[0]),.doutb(w_n753_8[1]),.din(w_n753_2[1]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.din(n761));
	jspl3 jspl3_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.doutc(w_n765_0[2]),.din(w_dff_B_f8EmpGFW4_3));
	jspl3 jspl3_w_n765_1(.douta(w_n765_1[0]),.doutb(w_n765_1[1]),.doutc(w_n765_1[2]),.din(w_n765_0[0]));
	jspl3 jspl3_w_n765_2(.douta(w_n765_2[0]),.doutb(w_n765_2[1]),.doutc(w_n765_2[2]),.din(w_n765_0[1]));
	jspl3 jspl3_w_n765_3(.douta(w_n765_3[0]),.doutb(w_n765_3[1]),.doutc(w_n765_3[2]),.din(w_n765_0[2]));
	jspl3 jspl3_w_n765_4(.douta(w_n765_4[0]),.doutb(w_n765_4[1]),.doutc(w_n765_4[2]),.din(w_n765_1[0]));
	jspl3 jspl3_w_n765_5(.douta(w_n765_5[0]),.doutb(w_n765_5[1]),.doutc(w_n765_5[2]),.din(w_n765_1[1]));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_dff_A_WZyU70B86_1),.din(n779));
	jspl3 jspl3_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.doutc(w_n781_0[2]),.din(n781));
	jspl3 jspl3_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.doutc(w_n783_0[2]),.din(n783));
	jspl jspl_w_n783_1(.douta(w_n783_1[0]),.doutb(w_n783_1[1]),.din(w_n783_0[0]));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_tswFWHNN0_2));
	jspl3 jspl3_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.doutc(w_n789_0[2]),.din(n789));
	jspl3 jspl3_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.doutc(w_n791_0[2]),.din(n791));
	jspl jspl_w_n791_1(.douta(w_n791_1[0]),.doutb(w_n791_1[1]),.din(w_n791_0[0]));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl3 jspl3_w_n793_0(.douta(w_n793_0[0]),.doutb(w_dff_A_Uck6BVVc7_1),.doutc(w_dff_A_uxzSyXNv7_2),.din(w_dff_B_IRk8CjcP4_3));
	jspl3 jspl3_w_n793_1(.douta(w_n793_1[0]),.doutb(w_dff_A_awGli8B57_1),.doutc(w_dff_A_lGSOXHj04_2),.din(w_n793_0[0]));
	jspl3 jspl3_w_n793_2(.douta(w_n793_2[0]),.doutb(w_n793_2[1]),.doutc(w_dff_A_DvvXWMSC4_2),.din(w_n793_0[1]));
	jspl3 jspl3_w_n793_3(.douta(w_n793_3[0]),.doutb(w_dff_A_3hxACZ724_1),.doutc(w_dff_A_Lfpu8aaD6_2),.din(w_n793_0[2]));
	jspl jspl_w_n793_4(.douta(w_dff_A_DkCylNHW6_0),.doutb(w_n793_4[1]),.din(w_n793_1[0]));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_dff_A_la6I0zsv1_1),.doutc(w_dff_A_8c8YIv9Z3_2),.din(w_dff_B_fkxGB2wk5_3));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_dff_A_qovNcWLc4_1),.doutc(w_dff_A_Ae5SNb7y0_2),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_dff_A_4KE5DLLY1_2),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_n797_3[0]),.doutb(w_dff_A_GAy0RsyZ9_1),.doutc(w_dff_A_1vjksKh00_2),.din(w_n797_0[2]));
	jspl jspl_w_n797_4(.douta(w_dff_A_4KOxYKIx5_0),.doutb(w_n797_4[1]),.din(w_n797_1[0]));
	jspl3 jspl3_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.doutc(w_n799_0[2]),.din(n799));
	jspl3 jspl3_w_n799_1(.douta(w_n799_1[0]),.doutb(w_n799_1[1]),.doutc(w_n799_1[2]),.din(w_n799_0[0]));
	jspl3 jspl3_w_n799_2(.douta(w_n799_2[0]),.doutb(w_n799_2[1]),.doutc(w_n799_2[2]),.din(w_n799_0[1]));
	jspl3 jspl3_w_n799_3(.douta(w_n799_3[0]),.doutb(w_n799_3[1]),.doutc(w_n799_3[2]),.din(w_n799_0[2]));
	jspl jspl_w_n799_4(.douta(w_n799_4[0]),.doutb(w_n799_4[1]),.din(w_n799_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl3 jspl3_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.doutc(w_n801_1[2]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n801_2(.douta(w_n801_2[0]),.doutb(w_n801_2[1]),.doutc(w_n801_2[2]),.din(w_n801_0[1]));
	jspl3 jspl3_w_n801_3(.douta(w_n801_3[0]),.doutb(w_n801_3[1]),.doutc(w_n801_3[2]),.din(w_n801_0[2]));
	jspl jspl_w_n801_4(.douta(w_n801_4[0]),.doutb(w_n801_4[1]),.din(w_n801_1[0]));
	jspl3 jspl3_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.doutc(w_n806_0[2]),.din(n806));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(n821));
	jspl3 jspl3_w_n828_0(.douta(w_n828_0[0]),.doutb(w_dff_A_VnwMUdos2_1),.doutc(w_dff_A_WutHriiW2_2),.din(n828));
	jspl jspl_w_n829_0(.douta(w_n829_0[0]),.doutb(w_dff_A_C6FdzPPt8_1),.din(n829));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl3 jspl3_w_n840_0(.douta(w_n840_0[0]),.doutb(w_dff_A_I5c4OnJa6_1),.doutc(w_dff_A_6bUW0NZ23_2),.din(w_dff_B_Ua5DCBO99_3));
	jspl3 jspl3_w_n840_1(.douta(w_n840_1[0]),.doutb(w_dff_A_oPFxAwah3_1),.doutc(w_dff_A_Jy2uufCu7_2),.din(w_n840_0[0]));
	jspl3 jspl3_w_n840_2(.douta(w_n840_2[0]),.doutb(w_n840_2[1]),.doutc(w_dff_A_JkQzaEnP2_2),.din(w_n840_0[1]));
	jspl3 jspl3_w_n840_3(.douta(w_n840_3[0]),.doutb(w_dff_A_GYLz104K6_1),.doutc(w_dff_A_4wKiggY12_2),.din(w_n840_0[2]));
	jspl jspl_w_n840_4(.douta(w_dff_A_XDZ3xYaL9_0),.doutb(w_n840_4[1]),.din(w_n840_1[0]));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(n842));
	jspl3 jspl3_w_n843_0(.douta(w_n843_0[0]),.doutb(w_dff_A_mwCoMitu7_1),.doutc(w_dff_A_b3PzTxgP3_2),.din(w_dff_B_NoFcKoJw2_3));
	jspl3 jspl3_w_n843_1(.douta(w_n843_1[0]),.doutb(w_dff_A_0HiOG1SP1_1),.doutc(w_dff_A_vuhtRYQD6_2),.din(w_n843_0[0]));
	jspl3 jspl3_w_n843_2(.douta(w_n843_2[0]),.doutb(w_n843_2[1]),.doutc(w_dff_A_HPZV4S169_2),.din(w_n843_0[1]));
	jspl3 jspl3_w_n843_3(.douta(w_n843_3[0]),.doutb(w_dff_A_5mewilor6_1),.doutc(w_dff_A_n7jGp1G37_2),.din(w_n843_0[2]));
	jspl jspl_w_n843_4(.douta(w_dff_A_myzuL8GK8_0),.doutb(w_n843_4[1]),.din(w_n843_1[0]));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.doutc(w_n845_0[2]),.din(n845));
	jspl3 jspl3_w_n845_1(.douta(w_n845_1[0]),.doutb(w_n845_1[1]),.doutc(w_n845_1[2]),.din(w_n845_0[0]));
	jspl3 jspl3_w_n845_2(.douta(w_n845_2[0]),.doutb(w_n845_2[1]),.doutc(w_n845_2[2]),.din(w_n845_0[1]));
	jspl3 jspl3_w_n845_3(.douta(w_n845_3[0]),.doutb(w_n845_3[1]),.doutc(w_n845_3[2]),.din(w_n845_0[2]));
	jspl jspl_w_n845_4(.douta(w_n845_4[0]),.doutb(w_n845_4[1]),.din(w_n845_1[0]));
	jspl3 jspl3_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.doutc(w_n847_0[2]),.din(n847));
	jspl3 jspl3_w_n847_1(.douta(w_n847_1[0]),.doutb(w_n847_1[1]),.doutc(w_n847_1[2]),.din(w_n847_0[0]));
	jspl3 jspl3_w_n847_2(.douta(w_n847_2[0]),.doutb(w_n847_2[1]),.doutc(w_n847_2[2]),.din(w_n847_0[1]));
	jspl3 jspl3_w_n847_3(.douta(w_n847_3[0]),.doutb(w_n847_3[1]),.doutc(w_n847_3[2]),.din(w_n847_0[2]));
	jspl jspl_w_n847_4(.douta(w_n847_4[0]),.doutb(w_n847_4[1]),.din(w_n847_1[0]));
	jspl jspl_w_n853_0(.douta(w_n853_0[0]),.doutb(w_dff_A_zx1Zjokm5_1),.din(w_dff_B_Ro7kTiWC3_2));
	jspl jspl_w_n855_0(.douta(w_dff_A_VeQVEag42_0),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(n857));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(n862));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.din(n877));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n928_0(.douta(w_n928_0[0]),.doutb(w_dff_A_vb0eqkuN8_1),.din(w_dff_B_rI3rDfQO6_2));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_dff_A_PFBHx6OY6_2),.din(w_dff_B_ue2FJvjL9_3));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(w_dff_B_XYG7lamz1_2));
	jspl3 jspl3_w_n936_0(.douta(w_n936_0[0]),.doutb(w_n936_0[1]),.doutc(w_n936_0[2]),.din(n936));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(n938));
	jspl jspl_w_n941_0(.douta(w_n941_0[0]),.doutb(w_n941_0[1]),.din(n941));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_dff_A_QjppZzxw4_1),.din(n943));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_dff_A_IhjvjxkU8_1),.din(n944));
	jspl jspl_w_n946_0(.douta(w_n946_0[0]),.doutb(w_n946_0[1]),.din(n946));
	jspl3 jspl3_w_n948_0(.douta(w_n948_0[0]),.doutb(w_n948_0[1]),.doutc(w_n948_0[2]),.din(n948));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n968_0(.douta(w_n968_0[0]),.doutb(w_dff_A_JjHPO06u2_1),.din(w_dff_B_r2WXSA2G3_2));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_dff_A_NuJTEUlq2_1),.din(n971));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.din(n973));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl3 jspl3_w_n985_0(.douta(w_n985_0[0]),.doutb(w_dff_A_iYxEkZyg0_1),.doutc(w_dff_A_ICJEW9YY6_2),.din(n985));
	jspl3 jspl3_w_n985_1(.douta(w_dff_A_T9vIVRvM5_0),.doutb(w_n985_1[1]),.doutc(w_dff_A_MLToMRuZ9_2),.din(w_n985_0[0]));
	jspl3 jspl3_w_n985_2(.douta(w_dff_A_KOcAUxzg9_0),.doutb(w_dff_A_VeVRreo87_1),.doutc(w_n985_2[2]),.din(w_n985_0[1]));
	jspl3 jspl3_w_n985_3(.douta(w_dff_A_xRrmz9IE4_0),.doutb(w_dff_A_f3xGREPE5_1),.doutc(w_n985_3[2]),.din(w_n985_0[2]));
	jspl jspl_w_n985_4(.douta(w_dff_A_XSyHe9qJ0_0),.doutb(w_n985_4[1]),.din(w_n985_1[0]));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_dff_A_B9uKgh0B8_1),.doutc(w_dff_A_P2IcOBYT4_2),.din(n988));
	jspl3 jspl3_w_n988_1(.douta(w_dff_A_gpHh6toS5_0),.doutb(w_n988_1[1]),.doutc(w_dff_A_Z7o0FbIx1_2),.din(w_n988_0[0]));
	jspl3 jspl3_w_n988_2(.douta(w_dff_A_jkwCsyvQ2_0),.doutb(w_dff_A_ssvHqDnK6_1),.doutc(w_n988_2[2]),.din(w_n988_0[1]));
	jspl3 jspl3_w_n988_3(.douta(w_dff_A_ot3W3H814_0),.doutb(w_dff_A_FMUAtALP2_1),.doutc(w_n988_3[2]),.din(w_n988_0[2]));
	jspl jspl_w_n988_4(.douta(w_dff_A_ZStwA7746_0),.doutb(w_n988_4[1]),.din(w_n988_1[0]));
	jspl3 jspl3_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.doutc(w_n990_0[2]),.din(n990));
	jspl3 jspl3_w_n990_1(.douta(w_n990_1[0]),.doutb(w_n990_1[1]),.doutc(w_n990_1[2]),.din(w_n990_0[0]));
	jspl3 jspl3_w_n990_2(.douta(w_n990_2[0]),.doutb(w_n990_2[1]),.doutc(w_n990_2[2]),.din(w_n990_0[1]));
	jspl3 jspl3_w_n990_3(.douta(w_n990_3[0]),.doutb(w_n990_3[1]),.doutc(w_n990_3[2]),.din(w_n990_0[2]));
	jspl jspl_w_n990_4(.douta(w_n990_4[0]),.doutb(w_n990_4[1]),.din(w_n990_1[0]));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl3 jspl3_w_n992_1(.douta(w_n992_1[0]),.doutb(w_n992_1[1]),.doutc(w_n992_1[2]),.din(w_n992_0[0]));
	jspl3 jspl3_w_n992_2(.douta(w_n992_2[0]),.doutb(w_n992_2[1]),.doutc(w_n992_2[2]),.din(w_n992_0[1]));
	jspl3 jspl3_w_n992_3(.douta(w_n992_3[0]),.doutb(w_n992_3[1]),.doutc(w_n992_3[2]),.din(w_n992_0[2]));
	jspl jspl_w_n992_4(.douta(w_n992_4[0]),.doutb(w_n992_4[1]),.din(w_n992_1[0]));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_dff_A_XUckKp2H8_1),.doutc(w_dff_A_9XPHNBBU0_2),.din(n999));
	jspl3 jspl3_w_n999_1(.douta(w_dff_A_WnuzEvYQ9_0),.doutb(w_n999_1[1]),.doutc(w_dff_A_EYUNAq5J7_2),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_dff_A_EFjtmaS02_0),.doutb(w_dff_A_b2cAoQXM2_1),.doutc(w_n999_2[2]),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_dff_A_wxO2kF688_0),.doutb(w_dff_A_fSFRTojg7_1),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl jspl_w_n999_4(.douta(w_dff_A_rhsUaOPN5_0),.doutb(w_n999_4[1]),.din(w_n999_1[0]));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_dff_A_q4v7VrV62_1),.doutc(w_dff_A_Amqs3Bit9_2),.din(n1002));
	jspl3 jspl3_w_n1002_1(.douta(w_dff_A_ayovNCNM2_0),.doutb(w_n1002_1[1]),.doutc(w_dff_A_IMnGiKEn7_2),.din(w_n1002_0[0]));
	jspl3 jspl3_w_n1002_2(.douta(w_dff_A_QVXdpFrt1_0),.doutb(w_dff_A_PddqTTdc0_1),.doutc(w_n1002_2[2]),.din(w_n1002_0[1]));
	jspl3 jspl3_w_n1002_3(.douta(w_dff_A_AO2Fb7lv2_0),.doutb(w_dff_A_GC7RmWww4_1),.doutc(w_n1002_3[2]),.din(w_n1002_0[2]));
	jspl jspl_w_n1002_4(.douta(w_dff_A_9f3ZTmi57_0),.doutb(w_n1002_4[1]),.din(w_n1002_1[0]));
	jspl3 jspl3_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.doutc(w_n1004_0[2]),.din(n1004));
	jspl3 jspl3_w_n1004_1(.douta(w_n1004_1[0]),.doutb(w_n1004_1[1]),.doutc(w_n1004_1[2]),.din(w_n1004_0[0]));
	jspl3 jspl3_w_n1004_2(.douta(w_n1004_2[0]),.doutb(w_n1004_2[1]),.doutc(w_n1004_2[2]),.din(w_n1004_0[1]));
	jspl3 jspl3_w_n1004_3(.douta(w_n1004_3[0]),.doutb(w_n1004_3[1]),.doutc(w_n1004_3[2]),.din(w_n1004_0[2]));
	jspl jspl_w_n1004_4(.douta(w_n1004_4[0]),.doutb(w_n1004_4[1]),.din(w_n1004_1[0]));
	jspl3 jspl3_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.doutc(w_n1006_0[2]),.din(n1006));
	jspl3 jspl3_w_n1006_1(.douta(w_n1006_1[0]),.doutb(w_n1006_1[1]),.doutc(w_n1006_1[2]),.din(w_n1006_0[0]));
	jspl3 jspl3_w_n1006_2(.douta(w_n1006_2[0]),.doutb(w_n1006_2[1]),.doutc(w_n1006_2[2]),.din(w_n1006_0[1]));
	jspl3 jspl3_w_n1006_3(.douta(w_n1006_3[0]),.doutb(w_n1006_3[1]),.doutc(w_n1006_3[2]),.din(w_n1006_0[2]));
	jspl jspl_w_n1006_4(.douta(w_n1006_4[0]),.doutb(w_n1006_4[1]),.din(w_n1006_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl jspl_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl jspl_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.doutc(w_n1023_0[2]),.din(n1023));
	jspl jspl_w_n1023_1(.douta(w_n1023_1[0]),.doutb(w_n1023_1[1]),.din(w_n1023_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.doutc(w_n1039_0[2]),.din(n1039));
	jspl jspl_w_n1039_1(.douta(w_n1039_1[0]),.doutb(w_n1039_1[1]),.din(w_n1039_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl jspl_w_n1142_0(.douta(w_dff_A_uMQUu5Mt4_0),.doutb(w_n1142_0[1]),.din(n1142));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(n1151));
	jspl3 jspl3_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.doutc(w_n1163_0[2]),.din(n1163));
	jspl3 jspl3_w_n1163_1(.douta(w_n1163_1[0]),.doutb(w_n1163_1[1]),.doutc(w_n1163_1[2]),.din(w_n1163_0[0]));
	jspl3 jspl3_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.doutc(w_n1197_0[2]),.din(n1197));
	jspl3 jspl3_w_n1197_1(.douta(w_n1197_1[0]),.doutb(w_n1197_1[1]),.doutc(w_n1197_1[2]),.din(w_n1197_0[0]));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.doutc(w_n1235_0[2]),.din(n1235));
	jspl jspl_w_n1235_1(.douta(w_n1235_1[0]),.doutb(w_n1235_1[1]),.din(w_n1235_0[0]));
	jspl3 jspl3_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.doutc(w_n1242_0[2]),.din(n1242));
	jspl jspl_w_n1242_1(.douta(w_n1242_1[0]),.doutb(w_n1242_1[1]),.din(w_n1242_0[0]));
	jspl3 jspl3_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.doutc(w_n1244_0[2]),.din(n1244));
	jspl jspl_w_n1244_1(.douta(w_n1244_1[0]),.doutb(w_n1244_1[1]),.din(w_n1244_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl jspl_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.doutc(w_n1253_0[2]),.din(n1253));
	jspl jspl_w_n1253_1(.douta(w_n1253_1[0]),.doutb(w_n1253_1[1]),.din(w_n1253_0[0]));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1383_0(.douta(w_dff_A_ZDq3w5ma4_0),.doutb(w_n1383_0[1]),.din(n1383));
	jspl jspl_w_n1391_0(.douta(w_dff_A_HBen2u2L4_0),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(n1399));
	jspl jspl_w_n1409_0(.douta(w_dff_A_xyxMXKFh7_0),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(n1410));
	jspl jspl_w_n1411_0(.douta(w_dff_A_jIOBzIQ13_0),.doutb(w_n1411_0[1]),.din(n1411));
	jspl jspl_w_n1421_0(.douta(w_dff_A_JXVu36Ka7_0),.doutb(w_n1421_0[1]),.din(n1421));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_dff_A_KzB0g1Nb1_1),.din(n1438));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_dff_A_fgrJABZv7_1),.din(n1447));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(n1494));
	jspl jspl_w_n1533_0(.douta(w_n1533_0[0]),.doutb(w_n1533_0[1]),.din(w_dff_B_tFWjCfY76_2));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(w_dff_B_kuwmshAL9_2));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(w_dff_B_Dy6tX2Yq7_2));
	jspl jspl_w_n1555_0(.douta(w_dff_A_jvBsZeVC2_0),.doutb(w_n1555_0[1]),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_dff_A_cq8EeuVL6_1),.din(n1568));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(n1597));
	jspl3 jspl3_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.doutc(w_n1601_0[2]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_dff_A_8ibn2ThK1_1),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.din(w_dff_B_SUr3R1MO3_2));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(w_dff_B_JuqoCnrz3_2));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(w_dff_B_oUZfakXc6_2));
	jdff dff_B_Id93cNMm3_1(.din(G136),.dout(w_dff_B_Id93cNMm3_1),.clk(gclk));
	jdff dff_B_DSqho5bM5_0(.din(G2824),.dout(w_dff_B_DSqho5bM5_0),.clk(gclk));
	jdff dff_B_k7loCNst5_1(.din(n320),.dout(w_dff_B_k7loCNst5_1),.clk(gclk));
	jdff dff_B_gitFSkvp1_1(.din(n327),.dout(w_dff_B_gitFSkvp1_1),.clk(gclk));
	jdff dff_B_iIiqK0wI0_2(.din(n333),.dout(w_dff_B_iIiqK0wI0_2),.clk(gclk));
	jdff dff_B_lCHdGDBG8_1(.din(n338),.dout(w_dff_B_lCHdGDBG8_1),.clk(gclk));
	jdff dff_B_3iwXC5Ze8_1(.din(n340),.dout(w_dff_B_3iwXC5Ze8_1),.clk(gclk));
	jdff dff_B_WfzLEPFN3_0(.din(n341),.dout(w_dff_B_WfzLEPFN3_0),.clk(gclk));
	jdff dff_B_s29xw4Br7_1(.din(G24),.dout(w_dff_B_s29xw4Br7_1),.clk(gclk));
	jdff dff_B_P9Y9rX433_1(.din(n345),.dout(w_dff_B_P9Y9rX433_1),.clk(gclk));
	jdff dff_B_qQYrjorV2_0(.din(n346),.dout(w_dff_B_qQYrjorV2_0),.clk(gclk));
	jdff dff_B_hA9gudFc2_1(.din(G26),.dout(w_dff_B_hA9gudFc2_1),.clk(gclk));
	jdff dff_A_CPtyhCgc0_0(.dout(w_G141_2[0]),.din(w_dff_A_CPtyhCgc0_0),.clk(gclk));
	jdff dff_A_dpaXL5n99_0(.dout(w_dff_A_CPtyhCgc0_0),.din(w_dff_A_dpaXL5n99_0),.clk(gclk));
	jdff dff_A_77AqNmRZ4_0(.dout(w_dff_A_dpaXL5n99_0),.din(w_dff_A_77AqNmRZ4_0),.clk(gclk));
	jdff dff_A_4jl8JVpv6_0(.dout(w_dff_A_77AqNmRZ4_0),.din(w_dff_A_4jl8JVpv6_0),.clk(gclk));
	jdff dff_A_WXVNPlky6_1(.dout(w_G141_2[1]),.din(w_dff_A_WXVNPlky6_1),.clk(gclk));
	jdff dff_A_muhFrUle4_1(.dout(w_dff_A_WXVNPlky6_1),.din(w_dff_A_muhFrUle4_1),.clk(gclk));
	jdff dff_A_rRtH7eSm2_1(.dout(w_dff_A_muhFrUle4_1),.din(w_dff_A_rRtH7eSm2_1),.clk(gclk));
	jdff dff_A_7QRzfq9F4_1(.dout(w_dff_A_rRtH7eSm2_1),.din(w_dff_A_7QRzfq9F4_1),.clk(gclk));
	jdff dff_B_heedTL9O1_1(.din(n350),.dout(w_dff_B_heedTL9O1_1),.clk(gclk));
	jdff dff_B_inkwp1BG9_0(.din(n351),.dout(w_dff_B_inkwp1BG9_0),.clk(gclk));
	jdff dff_B_dQvTcDHr1_1(.din(G79),.dout(w_dff_B_dQvTcDHr1_1),.clk(gclk));
	jdff dff_B_ovleiaxu5_1(.din(n355),.dout(w_dff_B_ovleiaxu5_1),.clk(gclk));
	jdff dff_B_g5ylZoCc8_0(.din(n356),.dout(w_dff_B_g5ylZoCc8_0),.clk(gclk));
	jdff dff_B_dQxeAXvO7_1(.din(G82),.dout(w_dff_B_dQxeAXvO7_1),.clk(gclk));
	jdff dff_A_1ORJ7GLS6_0(.dout(w_G2358_2[0]),.din(w_dff_A_1ORJ7GLS6_0),.clk(gclk));
	jdff dff_A_CMurshcQ6_1(.dout(w_G2358_2[1]),.din(w_dff_A_CMurshcQ6_1),.clk(gclk));
	jdff dff_A_utxcD91K9_1(.dout(w_G141_1[1]),.din(w_dff_A_utxcD91K9_1),.clk(gclk));
	jdff dff_A_12zpmsxd2_1(.dout(w_dff_A_utxcD91K9_1),.din(w_dff_A_12zpmsxd2_1),.clk(gclk));
	jdff dff_A_eeMr8Due7_1(.dout(w_dff_A_12zpmsxd2_1),.din(w_dff_A_eeMr8Due7_1),.clk(gclk));
	jdff dff_A_Z5MG9Uvi3_1(.dout(w_dff_A_eeMr8Due7_1),.din(w_dff_A_Z5MG9Uvi3_1),.clk(gclk));
	jdff dff_A_3DeliFwL5_2(.dout(w_G141_1[2]),.din(w_dff_A_3DeliFwL5_2),.clk(gclk));
	jdff dff_A_6n70IdMj6_2(.dout(w_dff_A_3DeliFwL5_2),.din(w_dff_A_6n70IdMj6_2),.clk(gclk));
	jdff dff_A_zLBQMaug5_2(.dout(w_dff_A_6n70IdMj6_2),.din(w_dff_A_zLBQMaug5_2),.clk(gclk));
	jdff dff_A_Ot0zYzPB2_2(.dout(w_dff_A_zLBQMaug5_2),.din(w_dff_A_Ot0zYzPB2_2),.clk(gclk));
	jdff dff_B_dk8GTSgy6_1(.din(n384),.dout(w_dff_B_dk8GTSgy6_1),.clk(gclk));
	jdff dff_B_FuxDKOSc6_1(.din(w_dff_B_dk8GTSgy6_1),.dout(w_dff_B_FuxDKOSc6_1),.clk(gclk));
	jdff dff_B_83XCQ04X6_0(.din(n446),.dout(w_dff_B_83XCQ04X6_0),.clk(gclk));
	jdff dff_B_rTBel3Ui5_1(.din(n483),.dout(w_dff_B_rTBel3Ui5_1),.clk(gclk));
	jdff dff_B_fBBsNrfa9_1(.din(n506),.dout(w_dff_B_fBBsNrfa9_1),.clk(gclk));
	jdff dff_B_mEUW4q3f7_2(.din(n652),.dout(w_dff_B_mEUW4q3f7_2),.clk(gclk));
	jdff dff_B_EOZkHyo79_2(.din(n709),.dout(w_dff_B_EOZkHyo79_2),.clk(gclk));
	jdff dff_B_wjOfmtcp1_2(.din(w_dff_B_EOZkHyo79_2),.dout(w_dff_B_wjOfmtcp1_2),.clk(gclk));
	jdff dff_B_kq54St0X9_2(.din(w_dff_B_wjOfmtcp1_2),.dout(w_dff_B_kq54St0X9_2),.clk(gclk));
	jdff dff_B_e662TtVw6_1(.din(n698),.dout(w_dff_B_e662TtVw6_1),.clk(gclk));
	jdff dff_B_JbxfBhzd3_1(.din(w_dff_B_e662TtVw6_1),.dout(w_dff_B_JbxfBhzd3_1),.clk(gclk));
	jdff dff_B_acuTyYa16_1(.din(w_dff_B_JbxfBhzd3_1),.dout(w_dff_B_acuTyYa16_1),.clk(gclk));
	jdff dff_B_YYYGQkai2_1(.din(w_dff_B_acuTyYa16_1),.dout(w_dff_B_YYYGQkai2_1),.clk(gclk));
	jdff dff_B_EkNSJ5Jv2_1(.din(n699),.dout(w_dff_B_EkNSJ5Jv2_1),.clk(gclk));
	jdff dff_B_p9mcHn1a3_1(.din(w_dff_B_EkNSJ5Jv2_1),.dout(w_dff_B_p9mcHn1a3_1),.clk(gclk));
	jdff dff_B_sQ1LnrdP9_1(.din(w_dff_B_p9mcHn1a3_1),.dout(w_dff_B_sQ1LnrdP9_1),.clk(gclk));
	jdff dff_A_hmHkoDSJ2_1(.dout(w_n607_0[1]),.din(w_dff_A_hmHkoDSJ2_1),.clk(gclk));
	jdff dff_A_snnl1FyO3_1(.dout(w_dff_A_hmHkoDSJ2_1),.din(w_dff_A_snnl1FyO3_1),.clk(gclk));
	jdff dff_B_SDma8nWa1_3(.din(n607),.dout(w_dff_B_SDma8nWa1_3),.clk(gclk));
	jdff dff_B_r4ed7AqC9_3(.din(w_dff_B_SDma8nWa1_3),.dout(w_dff_B_r4ed7AqC9_3),.clk(gclk));
	jdff dff_B_7zdIdKpx6_3(.din(w_dff_B_r4ed7AqC9_3),.dout(w_dff_B_7zdIdKpx6_3),.clk(gclk));
	jdff dff_B_dI9q9fvR7_0(.din(n606),.dout(w_dff_B_dI9q9fvR7_0),.clk(gclk));
	jdff dff_B_XmCasODw0_2(.din(n742),.dout(w_dff_B_XmCasODw0_2),.clk(gclk));
	jdff dff_B_k4Ni3v0k9_2(.din(w_dff_B_XmCasODw0_2),.dout(w_dff_B_k4Ni3v0k9_2),.clk(gclk));
	jdff dff_B_B2RShfql6_2(.din(w_dff_B_k4Ni3v0k9_2),.dout(w_dff_B_B2RShfql6_2),.clk(gclk));
	jdff dff_B_AuYskGEF5_2(.din(w_dff_B_B2RShfql6_2),.dout(w_dff_B_AuYskGEF5_2),.clk(gclk));
	jdff dff_B_3Mdt917A2_2(.din(w_dff_B_AuYskGEF5_2),.dout(w_dff_B_3Mdt917A2_2),.clk(gclk));
	jdff dff_A_584demJC4_0(.dout(w_n651_1[0]),.din(w_dff_A_584demJC4_0),.clk(gclk));
	jdff dff_A_SO9kKnGd8_0(.dout(w_dff_A_584demJC4_0),.din(w_dff_A_SO9kKnGd8_0),.clk(gclk));
	jdff dff_A_3S8ZaUvv8_0(.dout(w_dff_A_SO9kKnGd8_0),.din(w_dff_A_3S8ZaUvv8_0),.clk(gclk));
	jdff dff_A_F0FyPtwW1_0(.dout(w_dff_A_3S8ZaUvv8_0),.din(w_dff_A_F0FyPtwW1_0),.clk(gclk));
	jdff dff_A_3qb3qbxk7_0(.dout(w_dff_A_F0FyPtwW1_0),.din(w_dff_A_3qb3qbxk7_0),.clk(gclk));
	jdff dff_A_bvaE7bz80_0(.dout(w_dff_A_3qb3qbxk7_0),.din(w_dff_A_bvaE7bz80_0),.clk(gclk));
	jdff dff_B_6eEd5HAd3_0(.din(n803),.dout(w_dff_B_6eEd5HAd3_0),.clk(gclk));
	jdff dff_B_nPNkbsto3_0(.din(w_dff_B_6eEd5HAd3_0),.dout(w_dff_B_nPNkbsto3_0),.clk(gclk));
	jdff dff_B_JJF1od7i7_0(.din(w_dff_B_nPNkbsto3_0),.dout(w_dff_B_JJF1od7i7_0),.clk(gclk));
	jdff dff_B_xGjOvOtH0_0(.din(w_dff_B_JJF1od7i7_0),.dout(w_dff_B_xGjOvOtH0_0),.clk(gclk));
	jdff dff_B_mmIR7lIl0_0(.din(w_dff_B_xGjOvOtH0_0),.dout(w_dff_B_mmIR7lIl0_0),.clk(gclk));
	jdff dff_B_hOLlBpdr3_0(.din(n802),.dout(w_dff_B_hOLlBpdr3_0),.clk(gclk));
	jdff dff_B_hkTuO8SI5_0(.din(n849),.dout(w_dff_B_hkTuO8SI5_0),.clk(gclk));
	jdff dff_B_are00Gb59_0(.din(w_dff_B_hkTuO8SI5_0),.dout(w_dff_B_are00Gb59_0),.clk(gclk));
	jdff dff_B_vBR5umxJ2_0(.din(w_dff_B_are00Gb59_0),.dout(w_dff_B_vBR5umxJ2_0),.clk(gclk));
	jdff dff_B_PiEWqbwA4_0(.din(w_dff_B_vBR5umxJ2_0),.dout(w_dff_B_PiEWqbwA4_0),.clk(gclk));
	jdff dff_B_xNysK2R40_0(.din(w_dff_B_PiEWqbwA4_0),.dout(w_dff_B_xNysK2R40_0),.clk(gclk));
	jdff dff_B_tx0jMe6i2_0(.din(n848),.dout(w_dff_B_tx0jMe6i2_0),.clk(gclk));
	jdff dff_B_4HhBeV5W9_2(.din(G61),.dout(w_dff_B_4HhBeV5W9_2),.clk(gclk));
	jdff dff_B_nG3bsuQb7_2(.din(G11),.dout(w_dff_B_nG3bsuQb7_2),.clk(gclk));
	jdff dff_B_TTi3HKcw0_2(.din(w_dff_B_nG3bsuQb7_2),.dout(w_dff_B_TTi3HKcw0_2),.clk(gclk));
	jdff dff_B_bkgjFZb24_0(.din(n964),.dout(w_dff_B_bkgjFZb24_0),.clk(gclk));
	jdff dff_B_5yVzVK379_0(.din(n962),.dout(w_dff_B_5yVzVK379_0),.clk(gclk));
	jdff dff_B_TcczeA249_0(.din(n961),.dout(w_dff_B_TcczeA249_0),.clk(gclk));
	jdff dff_B_ndD6yr1S9_1(.din(n957),.dout(w_dff_B_ndD6yr1S9_1),.clk(gclk));
	jdff dff_B_y5H00sBe8_1(.din(w_dff_B_ndD6yr1S9_1),.dout(w_dff_B_y5H00sBe8_1),.clk(gclk));
	jdff dff_B_SIf5AlHq5_1(.din(w_dff_B_y5H00sBe8_1),.dout(w_dff_B_SIf5AlHq5_1),.clk(gclk));
	jdff dff_B_0C521gtF5_1(.din(w_dff_B_SIf5AlHq5_1),.dout(w_dff_B_0C521gtF5_1),.clk(gclk));
	jdff dff_B_raMBVX0g9_0(.din(n980),.dout(w_dff_B_raMBVX0g9_0),.clk(gclk));
	jdff dff_B_tWjqZr2a1_0(.din(w_dff_B_raMBVX0g9_0),.dout(w_dff_B_tWjqZr2a1_0),.clk(gclk));
	jdff dff_B_vcqIHBmT2_0(.din(n979),.dout(w_dff_B_vcqIHBmT2_0),.clk(gclk));
	jdff dff_B_ksLsfQMS2_0(.din(n978),.dout(w_dff_B_ksLsfQMS2_0),.clk(gclk));
	jdff dff_B_0G1dH7Rk3_0(.din(n977),.dout(w_dff_B_0G1dH7Rk3_0),.clk(gclk));
	jdff dff_B_i6oJGg1L9_0(.din(n976),.dout(w_dff_B_i6oJGg1L9_0),.clk(gclk));
	jdff dff_B_eoOl4jo23_0(.din(n994),.dout(w_dff_B_eoOl4jo23_0),.clk(gclk));
	jdff dff_B_xwx7QPtN4_0(.din(w_dff_B_eoOl4jo23_0),.dout(w_dff_B_xwx7QPtN4_0),.clk(gclk));
	jdff dff_B_xinGAnSF1_0(.din(w_dff_B_xwx7QPtN4_0),.dout(w_dff_B_xinGAnSF1_0),.clk(gclk));
	jdff dff_B_4099YKTg7_0(.din(w_dff_B_xinGAnSF1_0),.dout(w_dff_B_4099YKTg7_0),.clk(gclk));
	jdff dff_B_Dp2fIXZN1_0(.din(w_dff_B_4099YKTg7_0),.dout(w_dff_B_Dp2fIXZN1_0),.clk(gclk));
	jdff dff_B_THwIgXnc9_0(.din(n993),.dout(w_dff_B_THwIgXnc9_0),.clk(gclk));
	jdff dff_B_KMwqRnSO9_0(.din(n1008),.dout(w_dff_B_KMwqRnSO9_0),.clk(gclk));
	jdff dff_B_0YjR6u0w9_0(.din(w_dff_B_KMwqRnSO9_0),.dout(w_dff_B_0YjR6u0w9_0),.clk(gclk));
	jdff dff_B_W6kyvGYR7_0(.din(w_dff_B_0YjR6u0w9_0),.dout(w_dff_B_W6kyvGYR7_0),.clk(gclk));
	jdff dff_B_lkX286T74_0(.din(w_dff_B_W6kyvGYR7_0),.dout(w_dff_B_lkX286T74_0),.clk(gclk));
	jdff dff_B_zQrjFDnb9_0(.din(w_dff_B_lkX286T74_0),.dout(w_dff_B_zQrjFDnb9_0),.clk(gclk));
	jdff dff_B_UPcddqAS5_0(.din(n1007),.dout(w_dff_B_UPcddqAS5_0),.clk(gclk));
	jdff dff_B_TYlxeCwP3_2(.din(G185),.dout(w_dff_B_TYlxeCwP3_2),.clk(gclk));
	jdff dff_B_ycce6Lx65_2(.din(G182),.dout(w_dff_B_ycce6Lx65_2),.clk(gclk));
	jdff dff_B_3lqw6BQP3_2(.din(w_dff_B_ycce6Lx65_2),.dout(w_dff_B_3lqw6BQP3_2),.clk(gclk));
	jdff dff_B_chrVOFeU6_1(.din(n749),.dout(w_dff_B_chrVOFeU6_1),.clk(gclk));
	jdff dff_B_9ZXX0n5X8_0(.din(n754),.dout(w_dff_B_9ZXX0n5X8_0),.clk(gclk));
	jdff dff_B_81gYVq2G4_1(.din(G131),.dout(w_dff_B_81gYVq2G4_1),.clk(gclk));
	jdff dff_B_EU7b06o62_1(.din(w_dff_B_81gYVq2G4_1),.dout(w_dff_B_EU7b06o62_1),.clk(gclk));
	jdff dff_B_JgKebfju2_0(.din(n776),.dout(w_dff_B_JgKebfju2_0),.clk(gclk));
	jdff dff_B_9X5TAAfm0_0(.din(w_dff_B_JgKebfju2_0),.dout(w_dff_B_9X5TAAfm0_0),.clk(gclk));
	jdff dff_B_0Fmg88T65_1(.din(G117),.dout(w_dff_B_0Fmg88T65_1),.clk(gclk));
	jdff dff_B_ippiVCQk1_1(.din(w_dff_B_0Fmg88T65_1),.dout(w_dff_B_ippiVCQk1_1),.clk(gclk));
	jdff dff_B_mvkwBMxs2_0(.din(n504),.dout(w_dff_B_mvkwBMxs2_0),.clk(gclk));
	jdff dff_B_ZwRsMymD1_1(.din(n496),.dout(w_dff_B_ZwRsMymD1_1),.clk(gclk));
	jdff dff_B_TJ0WxKdf1_0(.din(n1019),.dout(w_dff_B_TJ0WxKdf1_0),.clk(gclk));
	jdff dff_B_BEryW3mD9_0(.din(n1018),.dout(w_dff_B_BEryW3mD9_0),.clk(gclk));
	jdff dff_B_8kp36Tmz3_0(.din(w_dff_B_BEryW3mD9_0),.dout(w_dff_B_8kp36Tmz3_0),.clk(gclk));
	jdff dff_B_cTT6ZgmG9_0(.din(w_dff_B_8kp36Tmz3_0),.dout(w_dff_B_cTT6ZgmG9_0),.clk(gclk));
	jdff dff_B_fsMSFOzP9_0(.din(w_dff_B_cTT6ZgmG9_0),.dout(w_dff_B_fsMSFOzP9_0),.clk(gclk));
	jdff dff_B_iLvON5Y48_0(.din(w_dff_B_fsMSFOzP9_0),.dout(w_dff_B_iLvON5Y48_0),.clk(gclk));
	jdff dff_B_nEHltJjm0_0(.din(w_dff_B_iLvON5Y48_0),.dout(w_dff_B_nEHltJjm0_0),.clk(gclk));
	jdff dff_B_StdsBtGU2_0(.din(w_dff_B_nEHltJjm0_0),.dout(w_dff_B_StdsBtGU2_0),.clk(gclk));
	jdff dff_B_1nls4XEo9_0(.din(w_dff_B_StdsBtGU2_0),.dout(w_dff_B_1nls4XEo9_0),.clk(gclk));
	jdff dff_B_uSB73dQf4_0(.din(w_dff_B_1nls4XEo9_0),.dout(w_dff_B_uSB73dQf4_0),.clk(gclk));
	jdff dff_B_YJA3jG9g3_0(.din(w_dff_B_uSB73dQf4_0),.dout(w_dff_B_YJA3jG9g3_0),.clk(gclk));
	jdff dff_B_lIOsDLVB3_0(.din(w_dff_B_YJA3jG9g3_0),.dout(w_dff_B_lIOsDLVB3_0),.clk(gclk));
	jdff dff_B_7oDXgmsj2_0(.din(w_dff_B_lIOsDLVB3_0),.dout(w_dff_B_7oDXgmsj2_0),.clk(gclk));
	jdff dff_B_tQiCExJB3_0(.din(n1017),.dout(w_dff_B_tQiCExJB3_0),.clk(gclk));
	jdff dff_A_siIh9YTQ4_0(.dout(w_n797_4[0]),.din(w_dff_A_siIh9YTQ4_0),.clk(gclk));
	jdff dff_A_T9K8nkUe0_0(.dout(w_dff_A_siIh9YTQ4_0),.din(w_dff_A_T9K8nkUe0_0),.clk(gclk));
	jdff dff_A_NmzcGEOh0_0(.dout(w_dff_A_T9K8nkUe0_0),.din(w_dff_A_NmzcGEOh0_0),.clk(gclk));
	jdff dff_A_ZeZBAic30_0(.dout(w_dff_A_NmzcGEOh0_0),.din(w_dff_A_ZeZBAic30_0),.clk(gclk));
	jdff dff_A_UffZVtVy7_0(.dout(w_dff_A_ZeZBAic30_0),.din(w_dff_A_UffZVtVy7_0),.clk(gclk));
	jdff dff_A_CtV7OBkU5_0(.dout(w_dff_A_UffZVtVy7_0),.din(w_dff_A_CtV7OBkU5_0),.clk(gclk));
	jdff dff_A_4KOxYKIx5_0(.dout(w_dff_A_CtV7OBkU5_0),.din(w_dff_A_4KOxYKIx5_0),.clk(gclk));
	jdff dff_A_5pih1i2L9_0(.dout(w_n793_4[0]),.din(w_dff_A_5pih1i2L9_0),.clk(gclk));
	jdff dff_A_cM2ntAS04_0(.dout(w_dff_A_5pih1i2L9_0),.din(w_dff_A_cM2ntAS04_0),.clk(gclk));
	jdff dff_A_MPc2zuvu5_0(.dout(w_dff_A_cM2ntAS04_0),.din(w_dff_A_MPc2zuvu5_0),.clk(gclk));
	jdff dff_A_lGXMKMcj6_0(.dout(w_dff_A_MPc2zuvu5_0),.din(w_dff_A_lGXMKMcj6_0),.clk(gclk));
	jdff dff_A_Nnrat7908_0(.dout(w_dff_A_lGXMKMcj6_0),.din(w_dff_A_Nnrat7908_0),.clk(gclk));
	jdff dff_A_n4Icl5t36_0(.dout(w_dff_A_Nnrat7908_0),.din(w_dff_A_n4Icl5t36_0),.clk(gclk));
	jdff dff_A_XKe6QUf15_0(.dout(w_dff_A_n4Icl5t36_0),.din(w_dff_A_XKe6QUf15_0),.clk(gclk));
	jdff dff_A_DkCylNHW6_0(.dout(w_dff_A_XKe6QUf15_0),.din(w_dff_A_DkCylNHW6_0),.clk(gclk));
	jdff dff_B_S0KAFPTt1_0(.din(n1028),.dout(w_dff_B_S0KAFPTt1_0),.clk(gclk));
	jdff dff_B_3noJ5F8U9_0(.din(n1027),.dout(w_dff_B_3noJ5F8U9_0),.clk(gclk));
	jdff dff_B_DBiEtEMf6_0(.din(w_dff_B_3noJ5F8U9_0),.dout(w_dff_B_DBiEtEMf6_0),.clk(gclk));
	jdff dff_B_HdwOqerz1_0(.din(w_dff_B_DBiEtEMf6_0),.dout(w_dff_B_HdwOqerz1_0),.clk(gclk));
	jdff dff_B_QcspVjQZ9_0(.din(w_dff_B_HdwOqerz1_0),.dout(w_dff_B_QcspVjQZ9_0),.clk(gclk));
	jdff dff_B_XOJ1yKqR0_0(.din(w_dff_B_QcspVjQZ9_0),.dout(w_dff_B_XOJ1yKqR0_0),.clk(gclk));
	jdff dff_B_fQ4IqU7U0_0(.din(w_dff_B_XOJ1yKqR0_0),.dout(w_dff_B_fQ4IqU7U0_0),.clk(gclk));
	jdff dff_B_lh8rfYao5_0(.din(w_dff_B_fQ4IqU7U0_0),.dout(w_dff_B_lh8rfYao5_0),.clk(gclk));
	jdff dff_B_SAB6UfdD7_0(.din(w_dff_B_lh8rfYao5_0),.dout(w_dff_B_SAB6UfdD7_0),.clk(gclk));
	jdff dff_B_yOmprw5H3_0(.din(w_dff_B_SAB6UfdD7_0),.dout(w_dff_B_yOmprw5H3_0),.clk(gclk));
	jdff dff_B_B2O0Sk7l4_0(.din(w_dff_B_yOmprw5H3_0),.dout(w_dff_B_B2O0Sk7l4_0),.clk(gclk));
	jdff dff_B_znZy9qvU2_0(.din(n1026),.dout(w_dff_B_znZy9qvU2_0),.clk(gclk));
	jdff dff_B_Qq9JiHcL5_0(.din(n1037),.dout(w_dff_B_Qq9JiHcL5_0),.clk(gclk));
	jdff dff_B_ffsg39Db4_0(.din(w_dff_B_Qq9JiHcL5_0),.dout(w_dff_B_ffsg39Db4_0),.clk(gclk));
	jdff dff_B_lcybjzNR4_0(.din(n1036),.dout(w_dff_B_lcybjzNR4_0),.clk(gclk));
	jdff dff_B_AAxLVVr25_0(.din(w_dff_B_lcybjzNR4_0),.dout(w_dff_B_AAxLVVr25_0),.clk(gclk));
	jdff dff_B_s8cdFx8V7_0(.din(w_dff_B_AAxLVVr25_0),.dout(w_dff_B_s8cdFx8V7_0),.clk(gclk));
	jdff dff_B_yvaNLqw83_0(.din(w_dff_B_s8cdFx8V7_0),.dout(w_dff_B_yvaNLqw83_0),.clk(gclk));
	jdff dff_B_SKYji9zI2_0(.din(w_dff_B_yvaNLqw83_0),.dout(w_dff_B_SKYji9zI2_0),.clk(gclk));
	jdff dff_B_jEQzjslZ4_0(.din(w_dff_B_SKYji9zI2_0),.dout(w_dff_B_jEQzjslZ4_0),.clk(gclk));
	jdff dff_B_ALIeBAhq3_0(.din(w_dff_B_jEQzjslZ4_0),.dout(w_dff_B_ALIeBAhq3_0),.clk(gclk));
	jdff dff_B_UXPXI8BI6_0(.din(w_dff_B_ALIeBAhq3_0),.dout(w_dff_B_UXPXI8BI6_0),.clk(gclk));
	jdff dff_B_lcWxHoXi5_0(.din(n1035),.dout(w_dff_B_lcWxHoXi5_0),.clk(gclk));
	jdff dff_B_WflnvAnp0_0(.din(n1046),.dout(w_dff_B_WflnvAnp0_0),.clk(gclk));
	jdff dff_B_NBbBKMGY2_0(.din(w_dff_B_WflnvAnp0_0),.dout(w_dff_B_NBbBKMGY2_0),.clk(gclk));
	jdff dff_B_eQZuP0F98_0(.din(w_dff_B_NBbBKMGY2_0),.dout(w_dff_B_eQZuP0F98_0),.clk(gclk));
	jdff dff_B_1dT86M9P1_0(.din(n1045),.dout(w_dff_B_1dT86M9P1_0),.clk(gclk));
	jdff dff_B_DrPeBPZ73_0(.din(w_dff_B_1dT86M9P1_0),.dout(w_dff_B_DrPeBPZ73_0),.clk(gclk));
	jdff dff_B_CxP69g5l7_0(.din(w_dff_B_DrPeBPZ73_0),.dout(w_dff_B_CxP69g5l7_0),.clk(gclk));
	jdff dff_B_ubqjtHnA6_0(.din(w_dff_B_CxP69g5l7_0),.dout(w_dff_B_ubqjtHnA6_0),.clk(gclk));
	jdff dff_B_k5AHAt704_0(.din(w_dff_B_ubqjtHnA6_0),.dout(w_dff_B_k5AHAt704_0),.clk(gclk));
	jdff dff_B_DtlcdPho4_0(.din(w_dff_B_k5AHAt704_0),.dout(w_dff_B_DtlcdPho4_0),.clk(gclk));
	jdff dff_B_6hnVM6k33_0(.din(n1044),.dout(w_dff_B_6hnVM6k33_0),.clk(gclk));
	jdff dff_A_b9DxND8P5_1(.dout(w_n797_3[1]),.din(w_dff_A_b9DxND8P5_1),.clk(gclk));
	jdff dff_A_GAy0RsyZ9_1(.dout(w_dff_A_b9DxND8P5_1),.din(w_dff_A_GAy0RsyZ9_1),.clk(gclk));
	jdff dff_A_i8BZwpIx3_2(.dout(w_n797_3[2]),.din(w_dff_A_i8BZwpIx3_2),.clk(gclk));
	jdff dff_A_EzAR2vfD0_2(.dout(w_dff_A_i8BZwpIx3_2),.din(w_dff_A_EzAR2vfD0_2),.clk(gclk));
	jdff dff_A_gxRIdmRO6_2(.dout(w_dff_A_EzAR2vfD0_2),.din(w_dff_A_gxRIdmRO6_2),.clk(gclk));
	jdff dff_A_1vjksKh00_2(.dout(w_dff_A_gxRIdmRO6_2),.din(w_dff_A_1vjksKh00_2),.clk(gclk));
	jdff dff_A_3hxACZ724_1(.dout(w_n793_3[1]),.din(w_dff_A_3hxACZ724_1),.clk(gclk));
	jdff dff_A_nA9xCYfF2_2(.dout(w_n793_3[2]),.din(w_dff_A_nA9xCYfF2_2),.clk(gclk));
	jdff dff_A_Lfpu8aaD6_2(.dout(w_dff_A_nA9xCYfF2_2),.din(w_dff_A_Lfpu8aaD6_2),.clk(gclk));
	jdff dff_B_VK4V7vCg1_0(.din(n1053),.dout(w_dff_B_VK4V7vCg1_0),.clk(gclk));
	jdff dff_B_X84IcinJ8_0(.din(n1052),.dout(w_dff_B_X84IcinJ8_0),.clk(gclk));
	jdff dff_B_F0kYbrOg6_0(.din(w_dff_B_X84IcinJ8_0),.dout(w_dff_B_F0kYbrOg6_0),.clk(gclk));
	jdff dff_B_2JmCzuXy8_0(.din(w_dff_B_F0kYbrOg6_0),.dout(w_dff_B_2JmCzuXy8_0),.clk(gclk));
	jdff dff_B_T7yu0DrN0_0(.din(w_dff_B_2JmCzuXy8_0),.dout(w_dff_B_T7yu0DrN0_0),.clk(gclk));
	jdff dff_B_megj8YUu7_0(.din(w_dff_B_T7yu0DrN0_0),.dout(w_dff_B_megj8YUu7_0),.clk(gclk));
	jdff dff_B_TwlMCvBa1_0(.din(w_dff_B_megj8YUu7_0),.dout(w_dff_B_TwlMCvBa1_0),.clk(gclk));
	jdff dff_B_Txm6iwGw9_0(.din(w_dff_B_TwlMCvBa1_0),.dout(w_dff_B_Txm6iwGw9_0),.clk(gclk));
	jdff dff_B_YCyunKXF5_0(.din(w_dff_B_Txm6iwGw9_0),.dout(w_dff_B_YCyunKXF5_0),.clk(gclk));
	jdff dff_B_3EuztHLJ7_0(.din(w_dff_B_YCyunKXF5_0),.dout(w_dff_B_3EuztHLJ7_0),.clk(gclk));
	jdff dff_B_SJhukanT5_0(.din(w_dff_B_3EuztHLJ7_0),.dout(w_dff_B_SJhukanT5_0),.clk(gclk));
	jdff dff_B_mZq6ymBp8_0(.din(w_dff_B_SJhukanT5_0),.dout(w_dff_B_mZq6ymBp8_0),.clk(gclk));
	jdff dff_B_KvchqE8I4_0(.din(w_dff_B_mZq6ymBp8_0),.dout(w_dff_B_KvchqE8I4_0),.clk(gclk));
	jdff dff_B_YLKUDv2t1_0(.din(n1051),.dout(w_dff_B_YLKUDv2t1_0),.clk(gclk));
	jdff dff_B_0QNOVFad6_2(.din(G37),.dout(w_dff_B_0QNOVFad6_2),.clk(gclk));
	jdff dff_B_RaUeAJfS3_2(.din(G43),.dout(w_dff_B_RaUeAJfS3_2),.clk(gclk));
	jdff dff_B_lWeXAT4l1_2(.din(w_dff_B_RaUeAJfS3_2),.dout(w_dff_B_lWeXAT4l1_2),.clk(gclk));
	jdff dff_A_iEuz810I1_0(.dout(w_n843_4[0]),.din(w_dff_A_iEuz810I1_0),.clk(gclk));
	jdff dff_A_j2DrEfx60_0(.dout(w_dff_A_iEuz810I1_0),.din(w_dff_A_j2DrEfx60_0),.clk(gclk));
	jdff dff_A_xCZoYyqu2_0(.dout(w_dff_A_j2DrEfx60_0),.din(w_dff_A_xCZoYyqu2_0),.clk(gclk));
	jdff dff_A_zoOfQhIk5_0(.dout(w_dff_A_xCZoYyqu2_0),.din(w_dff_A_zoOfQhIk5_0),.clk(gclk));
	jdff dff_A_GRzwZhCM5_0(.dout(w_dff_A_zoOfQhIk5_0),.din(w_dff_A_GRzwZhCM5_0),.clk(gclk));
	jdff dff_A_76G6ei0f1_0(.dout(w_dff_A_GRzwZhCM5_0),.din(w_dff_A_76G6ei0f1_0),.clk(gclk));
	jdff dff_A_myzuL8GK8_0(.dout(w_dff_A_76G6ei0f1_0),.din(w_dff_A_myzuL8GK8_0),.clk(gclk));
	jdff dff_A_15d2twUx4_0(.dout(w_n840_4[0]),.din(w_dff_A_15d2twUx4_0),.clk(gclk));
	jdff dff_A_r86EQqaE6_0(.dout(w_dff_A_15d2twUx4_0),.din(w_dff_A_r86EQqaE6_0),.clk(gclk));
	jdff dff_A_RaPU5EZW3_0(.dout(w_dff_A_r86EQqaE6_0),.din(w_dff_A_RaPU5EZW3_0),.clk(gclk));
	jdff dff_A_TpZCxc8j7_0(.dout(w_dff_A_RaPU5EZW3_0),.din(w_dff_A_TpZCxc8j7_0),.clk(gclk));
	jdff dff_A_dWmleysb5_0(.dout(w_dff_A_TpZCxc8j7_0),.din(w_dff_A_dWmleysb5_0),.clk(gclk));
	jdff dff_A_Rrfn7o2r5_0(.dout(w_dff_A_dWmleysb5_0),.din(w_dff_A_Rrfn7o2r5_0),.clk(gclk));
	jdff dff_A_MRSr68jt7_0(.dout(w_dff_A_Rrfn7o2r5_0),.din(w_dff_A_MRSr68jt7_0),.clk(gclk));
	jdff dff_A_XDZ3xYaL9_0(.dout(w_dff_A_MRSr68jt7_0),.din(w_dff_A_XDZ3xYaL9_0),.clk(gclk));
	jdff dff_B_rOb8Gu7a6_0(.din(n1060),.dout(w_dff_B_rOb8Gu7a6_0),.clk(gclk));
	jdff dff_B_qsVRSY6K4_0(.din(n1059),.dout(w_dff_B_qsVRSY6K4_0),.clk(gclk));
	jdff dff_B_c5OiLB299_0(.din(w_dff_B_qsVRSY6K4_0),.dout(w_dff_B_c5OiLB299_0),.clk(gclk));
	jdff dff_B_8uWItg6y1_0(.din(w_dff_B_c5OiLB299_0),.dout(w_dff_B_8uWItg6y1_0),.clk(gclk));
	jdff dff_B_FFGeZrdd1_0(.din(w_dff_B_8uWItg6y1_0),.dout(w_dff_B_FFGeZrdd1_0),.clk(gclk));
	jdff dff_B_qVawKd586_0(.din(w_dff_B_FFGeZrdd1_0),.dout(w_dff_B_qVawKd586_0),.clk(gclk));
	jdff dff_B_0Uv407OR2_0(.din(w_dff_B_qVawKd586_0),.dout(w_dff_B_0Uv407OR2_0),.clk(gclk));
	jdff dff_B_nt38ReTw0_0(.din(w_dff_B_0Uv407OR2_0),.dout(w_dff_B_nt38ReTw0_0),.clk(gclk));
	jdff dff_B_ZvjbCkJz7_0(.din(w_dff_B_nt38ReTw0_0),.dout(w_dff_B_ZvjbCkJz7_0),.clk(gclk));
	jdff dff_B_skoIA8Hf5_0(.din(w_dff_B_ZvjbCkJz7_0),.dout(w_dff_B_skoIA8Hf5_0),.clk(gclk));
	jdff dff_B_PBsKfb6g3_0(.din(w_dff_B_skoIA8Hf5_0),.dout(w_dff_B_PBsKfb6g3_0),.clk(gclk));
	jdff dff_B_QPJoRHpB9_0(.din(n1058),.dout(w_dff_B_QPJoRHpB9_0),.clk(gclk));
	jdff dff_B_ZKONFJX52_2(.din(G20),.dout(w_dff_B_ZKONFJX52_2),.clk(gclk));
	jdff dff_B_xKyJIKjB0_2(.din(G76),.dout(w_dff_B_xKyJIKjB0_2),.clk(gclk));
	jdff dff_B_mBRbiigd7_2(.din(w_dff_B_xKyJIKjB0_2),.dout(w_dff_B_mBRbiigd7_2),.clk(gclk));
	jdff dff_B_PZl9L0Ym4_0(.din(n1067),.dout(w_dff_B_PZl9L0Ym4_0),.clk(gclk));
	jdff dff_B_KKLryKvr9_0(.din(w_dff_B_PZl9L0Ym4_0),.dout(w_dff_B_KKLryKvr9_0),.clk(gclk));
	jdff dff_B_zOylP07W0_0(.din(n1066),.dout(w_dff_B_zOylP07W0_0),.clk(gclk));
	jdff dff_B_YrZPXZQH8_0(.din(w_dff_B_zOylP07W0_0),.dout(w_dff_B_YrZPXZQH8_0),.clk(gclk));
	jdff dff_B_gfrepL034_0(.din(w_dff_B_YrZPXZQH8_0),.dout(w_dff_B_gfrepL034_0),.clk(gclk));
	jdff dff_B_PmFodKp56_0(.din(w_dff_B_gfrepL034_0),.dout(w_dff_B_PmFodKp56_0),.clk(gclk));
	jdff dff_B_AnIR8f402_0(.din(w_dff_B_PmFodKp56_0),.dout(w_dff_B_AnIR8f402_0),.clk(gclk));
	jdff dff_B_U3vGkCaz8_0(.din(w_dff_B_AnIR8f402_0),.dout(w_dff_B_U3vGkCaz8_0),.clk(gclk));
	jdff dff_B_h6DRTrBX2_0(.din(w_dff_B_U3vGkCaz8_0),.dout(w_dff_B_h6DRTrBX2_0),.clk(gclk));
	jdff dff_B_eRBL8ZRO4_0(.din(w_dff_B_h6DRTrBX2_0),.dout(w_dff_B_eRBL8ZRO4_0),.clk(gclk));
	jdff dff_B_rpkLrdoL7_0(.din(n1065),.dout(w_dff_B_rpkLrdoL7_0),.clk(gclk));
	jdff dff_B_K4uE6dlT7_2(.din(G17),.dout(w_dff_B_K4uE6dlT7_2),.clk(gclk));
	jdff dff_B_S9df5jjs1_2(.din(G73),.dout(w_dff_B_S9df5jjs1_2),.clk(gclk));
	jdff dff_B_xqM8Xbir9_2(.din(w_dff_B_S9df5jjs1_2),.dout(w_dff_B_xqM8Xbir9_2),.clk(gclk));
	jdff dff_B_thv62NCx2_0(.din(n1074),.dout(w_dff_B_thv62NCx2_0),.clk(gclk));
	jdff dff_B_ccpSNxHr2_0(.din(w_dff_B_thv62NCx2_0),.dout(w_dff_B_ccpSNxHr2_0),.clk(gclk));
	jdff dff_B_j39BeYFI8_0(.din(w_dff_B_ccpSNxHr2_0),.dout(w_dff_B_j39BeYFI8_0),.clk(gclk));
	jdff dff_B_r3Vu4Yqw8_0(.din(n1073),.dout(w_dff_B_r3Vu4Yqw8_0),.clk(gclk));
	jdff dff_B_9teD8Blt0_0(.din(w_dff_B_r3Vu4Yqw8_0),.dout(w_dff_B_9teD8Blt0_0),.clk(gclk));
	jdff dff_B_uW1cntiw5_0(.din(w_dff_B_9teD8Blt0_0),.dout(w_dff_B_uW1cntiw5_0),.clk(gclk));
	jdff dff_B_fozBxNCC0_0(.din(w_dff_B_uW1cntiw5_0),.dout(w_dff_B_fozBxNCC0_0),.clk(gclk));
	jdff dff_B_tjLrggWN8_0(.din(w_dff_B_fozBxNCC0_0),.dout(w_dff_B_tjLrggWN8_0),.clk(gclk));
	jdff dff_B_NIVGXwuL9_0(.din(w_dff_B_tjLrggWN8_0),.dout(w_dff_B_NIVGXwuL9_0),.clk(gclk));
	jdff dff_B_VVfb37309_0(.din(n1072),.dout(w_dff_B_VVfb37309_0),.clk(gclk));
	jdff dff_B_P4yay9r89_2(.din(G70),.dout(w_dff_B_P4yay9r89_2),.clk(gclk));
	jdff dff_B_w22BrIXB0_2(.din(G67),.dout(w_dff_B_w22BrIXB0_2),.clk(gclk));
	jdff dff_B_IHXTYMqa1_2(.din(w_dff_B_w22BrIXB0_2),.dout(w_dff_B_IHXTYMqa1_2),.clk(gclk));
	jdff dff_A_gmM4reVL0_1(.dout(w_n843_3[1]),.din(w_dff_A_gmM4reVL0_1),.clk(gclk));
	jdff dff_A_5mewilor6_1(.dout(w_dff_A_gmM4reVL0_1),.din(w_dff_A_5mewilor6_1),.clk(gclk));
	jdff dff_A_ste0IyhO2_2(.dout(w_n843_3[2]),.din(w_dff_A_ste0IyhO2_2),.clk(gclk));
	jdff dff_A_nx0IpDTI1_2(.dout(w_dff_A_ste0IyhO2_2),.din(w_dff_A_nx0IpDTI1_2),.clk(gclk));
	jdff dff_A_DGHH2M3d7_2(.dout(w_dff_A_nx0IpDTI1_2),.din(w_dff_A_DGHH2M3d7_2),.clk(gclk));
	jdff dff_A_n7jGp1G37_2(.dout(w_dff_A_DGHH2M3d7_2),.din(w_dff_A_n7jGp1G37_2),.clk(gclk));
	jdff dff_A_GYLz104K6_1(.dout(w_n840_3[1]),.din(w_dff_A_GYLz104K6_1),.clk(gclk));
	jdff dff_A_rO3qYPbo2_2(.dout(w_n840_3[2]),.din(w_dff_A_rO3qYPbo2_2),.clk(gclk));
	jdff dff_A_4wKiggY12_2(.dout(w_dff_A_rO3qYPbo2_2),.din(w_dff_A_4wKiggY12_2),.clk(gclk));
	jdff dff_B_Y2Zix5Sa1_0(.din(n1081),.dout(w_dff_B_Y2Zix5Sa1_0),.clk(gclk));
	jdff dff_B_eHm6QLCe2_0(.din(n1080),.dout(w_dff_B_eHm6QLCe2_0),.clk(gclk));
	jdff dff_B_KFhwNKMZ7_0(.din(w_dff_B_eHm6QLCe2_0),.dout(w_dff_B_KFhwNKMZ7_0),.clk(gclk));
	jdff dff_B_XoJ6Wcqg3_0(.din(w_dff_B_KFhwNKMZ7_0),.dout(w_dff_B_XoJ6Wcqg3_0),.clk(gclk));
	jdff dff_B_iIJeOkQ01_0(.din(w_dff_B_XoJ6Wcqg3_0),.dout(w_dff_B_iIJeOkQ01_0),.clk(gclk));
	jdff dff_B_ctWpjLVU2_0(.din(w_dff_B_iIJeOkQ01_0),.dout(w_dff_B_ctWpjLVU2_0),.clk(gclk));
	jdff dff_B_gg1U3cVV0_0(.din(w_dff_B_ctWpjLVU2_0),.dout(w_dff_B_gg1U3cVV0_0),.clk(gclk));
	jdff dff_B_Y7siAdOu4_0(.din(w_dff_B_gg1U3cVV0_0),.dout(w_dff_B_Y7siAdOu4_0),.clk(gclk));
	jdff dff_B_e7Cx7APb6_0(.din(w_dff_B_Y7siAdOu4_0),.dout(w_dff_B_e7Cx7APb6_0),.clk(gclk));
	jdff dff_B_8z9ikzWw8_0(.din(w_dff_B_e7Cx7APb6_0),.dout(w_dff_B_8z9ikzWw8_0),.clk(gclk));
	jdff dff_B_8N4MIl7e1_0(.din(w_dff_B_8z9ikzWw8_0),.dout(w_dff_B_8N4MIl7e1_0),.clk(gclk));
	jdff dff_B_Tdso8v7U5_0(.din(w_dff_B_8N4MIl7e1_0),.dout(w_dff_B_Tdso8v7U5_0),.clk(gclk));
	jdff dff_B_1Kt4iVGy4_0(.din(w_dff_B_Tdso8v7U5_0),.dout(w_dff_B_1Kt4iVGy4_0),.clk(gclk));
	jdff dff_B_b2lq2Q2n7_0(.din(n1079),.dout(w_dff_B_b2lq2Q2n7_0),.clk(gclk));
	jdff dff_A_MyM5dgl37_0(.dout(w_n988_4[0]),.din(w_dff_A_MyM5dgl37_0),.clk(gclk));
	jdff dff_A_2tgNnHRA6_0(.dout(w_dff_A_MyM5dgl37_0),.din(w_dff_A_2tgNnHRA6_0),.clk(gclk));
	jdff dff_A_LaueRLuW3_0(.dout(w_dff_A_2tgNnHRA6_0),.din(w_dff_A_LaueRLuW3_0),.clk(gclk));
	jdff dff_A_wQu7aPfe9_0(.dout(w_dff_A_LaueRLuW3_0),.din(w_dff_A_wQu7aPfe9_0),.clk(gclk));
	jdff dff_A_XjvKCxDn1_0(.dout(w_dff_A_wQu7aPfe9_0),.din(w_dff_A_XjvKCxDn1_0),.clk(gclk));
	jdff dff_A_F9YEEKZ20_0(.dout(w_dff_A_XjvKCxDn1_0),.din(w_dff_A_F9YEEKZ20_0),.clk(gclk));
	jdff dff_A_ZStwA7746_0(.dout(w_dff_A_F9YEEKZ20_0),.din(w_dff_A_ZStwA7746_0),.clk(gclk));
	jdff dff_A_7SgxEgOr4_0(.dout(w_n985_4[0]),.din(w_dff_A_7SgxEgOr4_0),.clk(gclk));
	jdff dff_A_fo69tmbG0_0(.dout(w_dff_A_7SgxEgOr4_0),.din(w_dff_A_fo69tmbG0_0),.clk(gclk));
	jdff dff_A_HbNzWxqy1_0(.dout(w_dff_A_fo69tmbG0_0),.din(w_dff_A_HbNzWxqy1_0),.clk(gclk));
	jdff dff_A_0IuUq3qP9_0(.dout(w_dff_A_HbNzWxqy1_0),.din(w_dff_A_0IuUq3qP9_0),.clk(gclk));
	jdff dff_A_ykvi5NXc2_0(.dout(w_dff_A_0IuUq3qP9_0),.din(w_dff_A_ykvi5NXc2_0),.clk(gclk));
	jdff dff_A_ZrlNobvH1_0(.dout(w_dff_A_ykvi5NXc2_0),.din(w_dff_A_ZrlNobvH1_0),.clk(gclk));
	jdff dff_A_1EuSltka2_0(.dout(w_dff_A_ZrlNobvH1_0),.din(w_dff_A_1EuSltka2_0),.clk(gclk));
	jdff dff_A_XSyHe9qJ0_0(.dout(w_dff_A_1EuSltka2_0),.din(w_dff_A_XSyHe9qJ0_0),.clk(gclk));
	jdff dff_B_dsAkIOls6_0(.din(n1089),.dout(w_dff_B_dsAkIOls6_0),.clk(gclk));
	jdff dff_B_iqL5QVgb3_0(.din(w_dff_B_dsAkIOls6_0),.dout(w_dff_B_iqL5QVgb3_0),.clk(gclk));
	jdff dff_B_zYIkRZYU7_0(.din(w_dff_B_iqL5QVgb3_0),.dout(w_dff_B_zYIkRZYU7_0),.clk(gclk));
	jdff dff_B_pTcSqvVJ1_0(.din(n1088),.dout(w_dff_B_pTcSqvVJ1_0),.clk(gclk));
	jdff dff_B_ezoTYRWu4_0(.din(w_dff_B_pTcSqvVJ1_0),.dout(w_dff_B_ezoTYRWu4_0),.clk(gclk));
	jdff dff_B_qwqwy70j8_0(.din(w_dff_B_ezoTYRWu4_0),.dout(w_dff_B_qwqwy70j8_0),.clk(gclk));
	jdff dff_B_cD8QjL1l0_0(.din(w_dff_B_qwqwy70j8_0),.dout(w_dff_B_cD8QjL1l0_0),.clk(gclk));
	jdff dff_B_5OMJYOqj2_0(.din(w_dff_B_cD8QjL1l0_0),.dout(w_dff_B_5OMJYOqj2_0),.clk(gclk));
	jdff dff_B_CWftwgeY8_0(.din(w_dff_B_5OMJYOqj2_0),.dout(w_dff_B_CWftwgeY8_0),.clk(gclk));
	jdff dff_B_6OrtFTWs5_0(.din(n1087),.dout(w_dff_B_6OrtFTWs5_0),.clk(gclk));
	jdff dff_B_d9CdKHzw7_0(.din(n1097),.dout(w_dff_B_d9CdKHzw7_0),.clk(gclk));
	jdff dff_B_rfDhlykd3_0(.din(w_dff_B_d9CdKHzw7_0),.dout(w_dff_B_rfDhlykd3_0),.clk(gclk));
	jdff dff_B_VtFPLDbu5_0(.din(n1096),.dout(w_dff_B_VtFPLDbu5_0),.clk(gclk));
	jdff dff_B_ABtbWRYA3_0(.din(w_dff_B_VtFPLDbu5_0),.dout(w_dff_B_ABtbWRYA3_0),.clk(gclk));
	jdff dff_B_xpOAJV1S0_0(.din(w_dff_B_ABtbWRYA3_0),.dout(w_dff_B_xpOAJV1S0_0),.clk(gclk));
	jdff dff_B_oQue21gJ4_0(.din(w_dff_B_xpOAJV1S0_0),.dout(w_dff_B_oQue21gJ4_0),.clk(gclk));
	jdff dff_B_gFJjeSU29_0(.din(w_dff_B_oQue21gJ4_0),.dout(w_dff_B_gFJjeSU29_0),.clk(gclk));
	jdff dff_B_fKMxE8QX4_0(.din(w_dff_B_gFJjeSU29_0),.dout(w_dff_B_fKMxE8QX4_0),.clk(gclk));
	jdff dff_B_kwlxKjSu6_0(.din(w_dff_B_fKMxE8QX4_0),.dout(w_dff_B_kwlxKjSu6_0),.clk(gclk));
	jdff dff_B_YWU8t7go8_0(.din(w_dff_B_kwlxKjSu6_0),.dout(w_dff_B_YWU8t7go8_0),.clk(gclk));
	jdff dff_B_76PEudjL8_0(.din(n1095),.dout(w_dff_B_76PEudjL8_0),.clk(gclk));
	jdff dff_A_bwDk8wJS5_0(.dout(w_G137_8[0]),.din(w_dff_A_bwDk8wJS5_0),.clk(gclk));
	jdff dff_A_y3mly7fF6_2(.dout(w_G137_8[2]),.din(w_dff_A_y3mly7fF6_2),.clk(gclk));
	jdff dff_A_CZH8B3ZO4_2(.dout(w_dff_A_y3mly7fF6_2),.din(w_dff_A_CZH8B3ZO4_2),.clk(gclk));
	jdff dff_A_dNH1hRh55_2(.dout(w_dff_A_CZH8B3ZO4_2),.din(w_dff_A_dNH1hRh55_2),.clk(gclk));
	jdff dff_A_c68Gy7OQ3_2(.dout(w_dff_A_dNH1hRh55_2),.din(w_dff_A_c68Gy7OQ3_2),.clk(gclk));
	jdff dff_B_oG0s388d4_0(.din(n1105),.dout(w_dff_B_oG0s388d4_0),.clk(gclk));
	jdff dff_B_Re9gNGJE1_0(.din(n1104),.dout(w_dff_B_Re9gNGJE1_0),.clk(gclk));
	jdff dff_B_fCmeMEMs2_0(.din(w_dff_B_Re9gNGJE1_0),.dout(w_dff_B_fCmeMEMs2_0),.clk(gclk));
	jdff dff_B_OtdQ3vFp6_0(.din(w_dff_B_fCmeMEMs2_0),.dout(w_dff_B_OtdQ3vFp6_0),.clk(gclk));
	jdff dff_B_tadGsxag7_0(.din(w_dff_B_OtdQ3vFp6_0),.dout(w_dff_B_tadGsxag7_0),.clk(gclk));
	jdff dff_B_gyA4NbWb8_0(.din(w_dff_B_tadGsxag7_0),.dout(w_dff_B_gyA4NbWb8_0),.clk(gclk));
	jdff dff_B_btZ3YHCc7_0(.din(w_dff_B_gyA4NbWb8_0),.dout(w_dff_B_btZ3YHCc7_0),.clk(gclk));
	jdff dff_B_vmAenznW3_0(.din(w_dff_B_btZ3YHCc7_0),.dout(w_dff_B_vmAenznW3_0),.clk(gclk));
	jdff dff_B_8GhYDpnR5_0(.din(w_dff_B_vmAenznW3_0),.dout(w_dff_B_8GhYDpnR5_0),.clk(gclk));
	jdff dff_B_2RcTZXdf2_0(.din(w_dff_B_8GhYDpnR5_0),.dout(w_dff_B_2RcTZXdf2_0),.clk(gclk));
	jdff dff_B_WAGQYCw72_0(.din(w_dff_B_2RcTZXdf2_0),.dout(w_dff_B_WAGQYCw72_0),.clk(gclk));
	jdff dff_B_BrlY33gH4_0(.din(n1103),.dout(w_dff_B_BrlY33gH4_0),.clk(gclk));
	jdff dff_A_Edw0dPLH8_0(.dout(w_n988_3[0]),.din(w_dff_A_Edw0dPLH8_0),.clk(gclk));
	jdff dff_A_1IpCWF9U5_0(.dout(w_dff_A_Edw0dPLH8_0),.din(w_dff_A_1IpCWF9U5_0),.clk(gclk));
	jdff dff_A_Dd6FveJz5_0(.dout(w_dff_A_1IpCWF9U5_0),.din(w_dff_A_Dd6FveJz5_0),.clk(gclk));
	jdff dff_A_ot3W3H814_0(.dout(w_dff_A_Dd6FveJz5_0),.din(w_dff_A_ot3W3H814_0),.clk(gclk));
	jdff dff_A_O4WcigL54_1(.dout(w_n988_3[1]),.din(w_dff_A_O4WcigL54_1),.clk(gclk));
	jdff dff_A_FMUAtALP2_1(.dout(w_dff_A_O4WcigL54_1),.din(w_dff_A_FMUAtALP2_1),.clk(gclk));
	jdff dff_A_GW5WSIsz3_0(.dout(w_n985_3[0]),.din(w_dff_A_GW5WSIsz3_0),.clk(gclk));
	jdff dff_A_xRrmz9IE4_0(.dout(w_dff_A_GW5WSIsz3_0),.din(w_dff_A_xRrmz9IE4_0),.clk(gclk));
	jdff dff_A_f3xGREPE5_1(.dout(w_n985_3[1]),.din(w_dff_A_f3xGREPE5_1),.clk(gclk));
	jdff dff_B_SKrf3Cde8_0(.din(n1113),.dout(w_dff_B_SKrf3Cde8_0),.clk(gclk));
	jdff dff_B_ST4Ndu5y9_0(.din(n1112),.dout(w_dff_B_ST4Ndu5y9_0),.clk(gclk));
	jdff dff_B_dP2IDRP77_0(.din(w_dff_B_ST4Ndu5y9_0),.dout(w_dff_B_dP2IDRP77_0),.clk(gclk));
	jdff dff_B_YkMBiu1n6_0(.din(w_dff_B_dP2IDRP77_0),.dout(w_dff_B_YkMBiu1n6_0),.clk(gclk));
	jdff dff_B_U6Z4UY655_0(.din(w_dff_B_YkMBiu1n6_0),.dout(w_dff_B_U6Z4UY655_0),.clk(gclk));
	jdff dff_B_rP59kVNh0_0(.din(w_dff_B_U6Z4UY655_0),.dout(w_dff_B_rP59kVNh0_0),.clk(gclk));
	jdff dff_B_gGfDCL4d3_0(.din(w_dff_B_rP59kVNh0_0),.dout(w_dff_B_gGfDCL4d3_0),.clk(gclk));
	jdff dff_B_fyntxCTa5_0(.din(w_dff_B_gGfDCL4d3_0),.dout(w_dff_B_fyntxCTa5_0),.clk(gclk));
	jdff dff_B_nDbgzLkI0_0(.din(w_dff_B_fyntxCTa5_0),.dout(w_dff_B_nDbgzLkI0_0),.clk(gclk));
	jdff dff_B_9rKyvyJg0_0(.din(w_dff_B_nDbgzLkI0_0),.dout(w_dff_B_9rKyvyJg0_0),.clk(gclk));
	jdff dff_B_Vw92Ic3y1_0(.din(w_dff_B_9rKyvyJg0_0),.dout(w_dff_B_Vw92Ic3y1_0),.clk(gclk));
	jdff dff_B_g7Khh2t65_0(.din(w_dff_B_Vw92Ic3y1_0),.dout(w_dff_B_g7Khh2t65_0),.clk(gclk));
	jdff dff_B_yTMNljsp9_0(.din(w_dff_B_g7Khh2t65_0),.dout(w_dff_B_yTMNljsp9_0),.clk(gclk));
	jdff dff_B_Q5CYsc8T9_0(.din(n1111),.dout(w_dff_B_Q5CYsc8T9_0),.clk(gclk));
	jdff dff_B_qpVakveK0_2(.din(G170),.dout(w_dff_B_qpVakveK0_2),.clk(gclk));
	jdff dff_B_3GXYxsTl9_2(.din(G200),.dout(w_dff_B_3GXYxsTl9_2),.clk(gclk));
	jdff dff_B_6uRl87Y29_2(.din(w_dff_B_3GXYxsTl9_2),.dout(w_dff_B_6uRl87Y29_2),.clk(gclk));
	jdff dff_A_txp6AFKK4_0(.dout(w_n1002_4[0]),.din(w_dff_A_txp6AFKK4_0),.clk(gclk));
	jdff dff_A_kPENjzXH4_0(.dout(w_dff_A_txp6AFKK4_0),.din(w_dff_A_kPENjzXH4_0),.clk(gclk));
	jdff dff_A_KCCsBxhm7_0(.dout(w_dff_A_kPENjzXH4_0),.din(w_dff_A_KCCsBxhm7_0),.clk(gclk));
	jdff dff_A_TjNvWTAN0_0(.dout(w_dff_A_KCCsBxhm7_0),.din(w_dff_A_TjNvWTAN0_0),.clk(gclk));
	jdff dff_A_UYkLgkoW6_0(.dout(w_dff_A_TjNvWTAN0_0),.din(w_dff_A_UYkLgkoW6_0),.clk(gclk));
	jdff dff_A_7gxD2dLE5_0(.dout(w_dff_A_UYkLgkoW6_0),.din(w_dff_A_7gxD2dLE5_0),.clk(gclk));
	jdff dff_A_9f3ZTmi57_0(.dout(w_dff_A_7gxD2dLE5_0),.din(w_dff_A_9f3ZTmi57_0),.clk(gclk));
	jdff dff_B_p4yQhdvH5_0(.din(n814),.dout(w_dff_B_p4yQhdvH5_0),.clk(gclk));
	jdff dff_B_5bWTsV5t1_0(.din(w_dff_B_p4yQhdvH5_0),.dout(w_dff_B_5bWTsV5t1_0),.clk(gclk));
	jdff dff_B_y2nyBVQl7_0(.din(w_dff_B_5bWTsV5t1_0),.dout(w_dff_B_y2nyBVQl7_0),.clk(gclk));
	jdff dff_B_2MlRsDzR6_0(.din(w_dff_B_y2nyBVQl7_0),.dout(w_dff_B_2MlRsDzR6_0),.clk(gclk));
	jdff dff_B_zUbZh2AH1_0(.din(w_dff_B_2MlRsDzR6_0),.dout(w_dff_B_zUbZh2AH1_0),.clk(gclk));
	jdff dff_B_TAKE6U3t4_0(.din(w_dff_B_zUbZh2AH1_0),.dout(w_dff_B_TAKE6U3t4_0),.clk(gclk));
	jdff dff_B_ZgiS9Y6b0_0(.din(n813),.dout(w_dff_B_ZgiS9Y6b0_0),.clk(gclk));
	jdff dff_B_r8g0D6iJ3_0(.din(w_dff_B_ZgiS9Y6b0_0),.dout(w_dff_B_r8g0D6iJ3_0),.clk(gclk));
	jdff dff_B_l5yiDbV36_1(.din(G52),.dout(w_dff_B_l5yiDbV36_1),.clk(gclk));
	jdff dff_B_QJjsEbXt0_1(.din(w_dff_B_l5yiDbV36_1),.dout(w_dff_B_QJjsEbXt0_1),.clk(gclk));
	jdff dff_B_6sGFwgL41_0(.din(n433),.dout(w_dff_B_6sGFwgL41_0),.clk(gclk));
	jdff dff_B_fVsMa68i5_1(.din(n425),.dout(w_dff_B_fVsMa68i5_1),.clk(gclk));
	jdff dff_A_fOleiBdk2_0(.dout(w_n999_4[0]),.din(w_dff_A_fOleiBdk2_0),.clk(gclk));
	jdff dff_A_y4LCp2Pi2_0(.dout(w_dff_A_fOleiBdk2_0),.din(w_dff_A_y4LCp2Pi2_0),.clk(gclk));
	jdff dff_A_FR3YClXm7_0(.dout(w_dff_A_y4LCp2Pi2_0),.din(w_dff_A_FR3YClXm7_0),.clk(gclk));
	jdff dff_A_dqmXt2a92_0(.dout(w_dff_A_FR3YClXm7_0),.din(w_dff_A_dqmXt2a92_0),.clk(gclk));
	jdff dff_A_QghXK8sy0_0(.dout(w_dff_A_dqmXt2a92_0),.din(w_dff_A_QghXK8sy0_0),.clk(gclk));
	jdff dff_A_PLgkUd441_0(.dout(w_dff_A_QghXK8sy0_0),.din(w_dff_A_PLgkUd441_0),.clk(gclk));
	jdff dff_A_A8eDiGPQ8_0(.dout(w_dff_A_PLgkUd441_0),.din(w_dff_A_A8eDiGPQ8_0),.clk(gclk));
	jdff dff_A_rhsUaOPN5_0(.dout(w_dff_A_A8eDiGPQ8_0),.din(w_dff_A_rhsUaOPN5_0),.clk(gclk));
	jdff dff_B_CE2Vl1ea9_0(.din(n867),.dout(w_dff_B_CE2Vl1ea9_0),.clk(gclk));
	jdff dff_B_DCAfXW7K4_0(.din(w_dff_B_CE2Vl1ea9_0),.dout(w_dff_B_DCAfXW7K4_0),.clk(gclk));
	jdff dff_B_KHwbTEck1_0(.din(w_dff_B_DCAfXW7K4_0),.dout(w_dff_B_KHwbTEck1_0),.clk(gclk));
	jdff dff_B_GGyalsZg4_0(.din(w_dff_B_KHwbTEck1_0),.dout(w_dff_B_GGyalsZg4_0),.clk(gclk));
	jdff dff_B_ogisMkkQ0_0(.din(w_dff_B_GGyalsZg4_0),.dout(w_dff_B_ogisMkkQ0_0),.clk(gclk));
	jdff dff_B_g6X9K9FW6_0(.din(w_dff_B_ogisMkkQ0_0),.dout(w_dff_B_g6X9K9FW6_0),.clk(gclk));
	jdff dff_B_oZMF7rnb0_0(.din(w_dff_B_g6X9K9FW6_0),.dout(w_dff_B_oZMF7rnb0_0),.clk(gclk));
	jdff dff_B_MjeizViB9_0(.din(w_dff_B_oZMF7rnb0_0),.dout(w_dff_B_MjeizViB9_0),.clk(gclk));
	jdff dff_B_vxOFMEb27_0(.din(n866),.dout(w_dff_B_vxOFMEb27_0),.clk(gclk));
	jdff dff_B_eQYXXswa6_0(.din(w_dff_B_vxOFMEb27_0),.dout(w_dff_B_eQYXXswa6_0),.clk(gclk));
	jdff dff_B_4mkfWb3v3_1(.din(G122),.dout(w_dff_B_4mkfWb3v3_1),.clk(gclk));
	jdff dff_B_25LjbvG77_1(.din(w_dff_B_4mkfWb3v3_1),.dout(w_dff_B_25LjbvG77_1),.clk(gclk));
	jdff dff_B_2SWRVRtF9_0(.din(n469),.dout(w_dff_B_2SWRVRtF9_0),.clk(gclk));
	jdff dff_B_RqnE4Ckq4_1(.din(n461),.dout(w_dff_B_RqnE4Ckq4_1),.clk(gclk));
	jdff dff_B_4kYylFYj6_1(.din(n852),.dout(w_dff_B_4kYylFYj6_1),.clk(gclk));
	jdff dff_B_AVJtX9VD2_1(.din(w_dff_B_4kYylFYj6_1),.dout(w_dff_B_AVJtX9VD2_1),.clk(gclk));
	jdff dff_B_jlHZhAgo0_1(.din(w_dff_B_AVJtX9VD2_1),.dout(w_dff_B_jlHZhAgo0_1),.clk(gclk));
	jdff dff_B_0Aud0Oz35_1(.din(w_dff_B_jlHZhAgo0_1),.dout(w_dff_B_0Aud0Oz35_1),.clk(gclk));
	jdff dff_B_rhrXIeUF6_1(.din(w_dff_B_0Aud0Oz35_1),.dout(w_dff_B_rhrXIeUF6_1),.clk(gclk));
	jdff dff_B_EHwVUm3b2_1(.din(w_dff_B_rhrXIeUF6_1),.dout(w_dff_B_EHwVUm3b2_1),.clk(gclk));
	jdff dff_B_6MMxw6cE9_0(.din(n1121),.dout(w_dff_B_6MMxw6cE9_0),.clk(gclk));
	jdff dff_B_JLQ03swz8_0(.din(w_dff_B_6MMxw6cE9_0),.dout(w_dff_B_JLQ03swz8_0),.clk(gclk));
	jdff dff_B_naGe759P5_0(.din(w_dff_B_JLQ03swz8_0),.dout(w_dff_B_naGe759P5_0),.clk(gclk));
	jdff dff_B_TrWoTZwY8_0(.din(n1120),.dout(w_dff_B_TrWoTZwY8_0),.clk(gclk));
	jdff dff_B_T0gOR15x1_0(.din(w_dff_B_TrWoTZwY8_0),.dout(w_dff_B_T0gOR15x1_0),.clk(gclk));
	jdff dff_B_NvtaKItF0_0(.din(w_dff_B_T0gOR15x1_0),.dout(w_dff_B_NvtaKItF0_0),.clk(gclk));
	jdff dff_B_vXHoK1Bw5_0(.din(w_dff_B_NvtaKItF0_0),.dout(w_dff_B_vXHoK1Bw5_0),.clk(gclk));
	jdff dff_B_Q6aPBvyk1_0(.din(w_dff_B_vXHoK1Bw5_0),.dout(w_dff_B_Q6aPBvyk1_0),.clk(gclk));
	jdff dff_B_1waQ82K29_0(.din(w_dff_B_Q6aPBvyk1_0),.dout(w_dff_B_1waQ82K29_0),.clk(gclk));
	jdff dff_B_0PbamN0N3_0(.din(n1119),.dout(w_dff_B_0PbamN0N3_0),.clk(gclk));
	jdff dff_B_Zkwko78p2_2(.din(G158),.dout(w_dff_B_Zkwko78p2_2),.clk(gclk));
	jdff dff_B_2KqurAVh2_2(.din(G188),.dout(w_dff_B_2KqurAVh2_2),.clk(gclk));
	jdff dff_B_9HPAWxIL1_2(.din(w_dff_B_2KqurAVh2_2),.dout(w_dff_B_9HPAWxIL1_2),.clk(gclk));
	jdff dff_B_EQ4dCWyB1_0(.din(n768),.dout(w_dff_B_EQ4dCWyB1_0),.clk(gclk));
	jdff dff_B_RNq2kfq04_0(.din(w_dff_B_EQ4dCWyB1_0),.dout(w_dff_B_RNq2kfq04_0),.clk(gclk));
	jdff dff_B_lXotI9so3_1(.din(G129),.dout(w_dff_B_lXotI9so3_1),.clk(gclk));
	jdff dff_B_H453Fxi78_1(.din(w_dff_B_lXotI9so3_1),.dout(w_dff_B_H453Fxi78_1),.clk(gclk));
	jdff dff_A_dmVkfCCc4_1(.dout(w_n397_0[1]),.din(w_dff_A_dmVkfCCc4_1),.clk(gclk));
	jdff dff_B_uOWGZG217_0(.din(n396),.dout(w_dff_B_uOWGZG217_0),.clk(gclk));
	jdff dff_B_sMPIbE0P2_1(.din(n387),.dout(w_dff_B_sMPIbE0P2_1),.clk(gclk));
	jdff dff_A_TCaFfdVO2_0(.dout(w_n748_4[0]),.din(w_dff_A_TCaFfdVO2_0),.clk(gclk));
	jdff dff_B_SCdRIpJo7_0(.din(n898),.dout(w_dff_B_SCdRIpJo7_0),.clk(gclk));
	jdff dff_B_6TiR4Avn9_0(.din(w_dff_B_SCdRIpJo7_0),.dout(w_dff_B_6TiR4Avn9_0),.clk(gclk));
	jdff dff_B_sglZAwff9_0(.din(w_dff_B_6TiR4Avn9_0),.dout(w_dff_B_sglZAwff9_0),.clk(gclk));
	jdff dff_B_sEKMPOcX8_0(.din(w_dff_B_sglZAwff9_0),.dout(w_dff_B_sEKMPOcX8_0),.clk(gclk));
	jdff dff_B_OJw71AoT6_0(.din(n897),.dout(w_dff_B_OJw71AoT6_0),.clk(gclk));
	jdff dff_B_p60ZL6903_0(.din(w_dff_B_OJw71AoT6_0),.dout(w_dff_B_p60ZL6903_0),.clk(gclk));
	jdff dff_B_0c9AXwHx1_1(.din(G126),.dout(w_dff_B_0c9AXwHx1_1),.clk(gclk));
	jdff dff_B_Dq5WLR2J7_1(.din(w_dff_B_0c9AXwHx1_1),.dout(w_dff_B_Dq5WLR2J7_1),.clk(gclk));
	jdff dff_B_zpjQOf2U6_0(.din(n493),.dout(w_dff_B_zpjQOf2U6_0),.clk(gclk));
	jdff dff_B_cYahSXIn8_1(.din(n485),.dout(w_dff_B_cYahSXIn8_1),.clk(gclk));
	jdff dff_B_FMmGyVGz9_0(.din(n889),.dout(w_dff_B_FMmGyVGz9_0),.clk(gclk));
	jdff dff_A_GltqHRr33_1(.dout(w_G137_7[1]),.din(w_dff_A_GltqHRr33_1),.clk(gclk));
	jdff dff_A_cKMotMgo0_1(.dout(w_dff_A_GltqHRr33_1),.din(w_dff_A_cKMotMgo0_1),.clk(gclk));
	jdff dff_A_lrYtObOH9_1(.dout(w_dff_A_cKMotMgo0_1),.din(w_dff_A_lrYtObOH9_1),.clk(gclk));
	jdff dff_A_D0fzhUMk0_1(.dout(w_dff_A_lrYtObOH9_1),.din(w_dff_A_D0fzhUMk0_1),.clk(gclk));
	jdff dff_A_f4pgnVYu9_2(.dout(w_G137_7[2]),.din(w_dff_A_f4pgnVYu9_2),.clk(gclk));
	jdff dff_A_QB56rGgY4_2(.dout(w_dff_A_f4pgnVYu9_2),.din(w_dff_A_QB56rGgY4_2),.clk(gclk));
	jdff dff_A_kN0rlN7D8_0(.dout(w_G137_2[0]),.din(w_dff_A_kN0rlN7D8_0),.clk(gclk));
	jdff dff_A_SQBn9wUY9_0(.dout(w_dff_A_kN0rlN7D8_0),.din(w_dff_A_SQBn9wUY9_0),.clk(gclk));
	jdff dff_A_vFivVuNl4_0(.dout(w_dff_A_SQBn9wUY9_0),.din(w_dff_A_vFivVuNl4_0),.clk(gclk));
	jdff dff_A_inyEzEyT3_0(.dout(w_dff_A_vFivVuNl4_0),.din(w_dff_A_inyEzEyT3_0),.clk(gclk));
	jdff dff_A_UIGabkCu4_1(.dout(w_G137_2[1]),.din(w_dff_A_UIGabkCu4_1),.clk(gclk));
	jdff dff_A_QPr2FzPM5_1(.dout(w_dff_A_UIGabkCu4_1),.din(w_dff_A_QPr2FzPM5_1),.clk(gclk));
	jdff dff_A_X1uiAiGC0_1(.dout(w_dff_A_QPr2FzPM5_1),.din(w_dff_A_X1uiAiGC0_1),.clk(gclk));
	jdff dff_A_e7EX4hop8_1(.dout(w_dff_A_X1uiAiGC0_1),.din(w_dff_A_e7EX4hop8_1),.clk(gclk));
	jdff dff_B_s4pokhNX4_0(.din(n1129),.dout(w_dff_B_s4pokhNX4_0),.clk(gclk));
	jdff dff_B_IL8mvxNn9_0(.din(w_dff_B_s4pokhNX4_0),.dout(w_dff_B_IL8mvxNn9_0),.clk(gclk));
	jdff dff_B_rUZ8gtx07_0(.din(n1128),.dout(w_dff_B_rUZ8gtx07_0),.clk(gclk));
	jdff dff_B_rePXtQT82_0(.din(w_dff_B_rUZ8gtx07_0),.dout(w_dff_B_rePXtQT82_0),.clk(gclk));
	jdff dff_B_AbKNlnNx9_0(.din(w_dff_B_rePXtQT82_0),.dout(w_dff_B_AbKNlnNx9_0),.clk(gclk));
	jdff dff_B_v13gxwy20_0(.din(w_dff_B_AbKNlnNx9_0),.dout(w_dff_B_v13gxwy20_0),.clk(gclk));
	jdff dff_B_Z51mgOLi5_0(.din(w_dff_B_v13gxwy20_0),.dout(w_dff_B_Z51mgOLi5_0),.clk(gclk));
	jdff dff_B_Dpg5Z6Ou4_0(.din(w_dff_B_Z51mgOLi5_0),.dout(w_dff_B_Dpg5Z6Ou4_0),.clk(gclk));
	jdff dff_B_0vdDPXmz7_0(.din(w_dff_B_Dpg5Z6Ou4_0),.dout(w_dff_B_0vdDPXmz7_0),.clk(gclk));
	jdff dff_B_57rtjik33_0(.din(w_dff_B_0vdDPXmz7_0),.dout(w_dff_B_57rtjik33_0),.clk(gclk));
	jdff dff_B_VTNitF7w1_0(.din(n1127),.dout(w_dff_B_VTNitF7w1_0),.clk(gclk));
	jdff dff_B_dOJaaTYT1_2(.din(G152),.dout(w_dff_B_dOJaaTYT1_2),.clk(gclk));
	jdff dff_B_uYTyBNBM2_2(.din(G155),.dout(w_dff_B_uYTyBNBM2_2),.clk(gclk));
	jdff dff_B_dOY9Sgmb6_2(.din(w_dff_B_uYTyBNBM2_2),.dout(w_dff_B_dOY9Sgmb6_2),.clk(gclk));
	jdff dff_B_boAqdgSE9_0(.din(n837),.dout(w_dff_B_boAqdgSE9_0),.clk(gclk));
	jdff dff_B_9lmp3lFb5_0(.din(w_dff_B_boAqdgSE9_0),.dout(w_dff_B_9lmp3lFb5_0),.clk(gclk));
	jdff dff_B_2WmBJGSp0_0(.din(n836),.dout(w_dff_B_2WmBJGSp0_0),.clk(gclk));
	jdff dff_B_hQgBgHlP8_0(.din(w_dff_B_2WmBJGSp0_0),.dout(w_dff_B_hQgBgHlP8_0),.clk(gclk));
	jdff dff_B_ER99DSjI7_1(.din(G119),.dout(w_dff_B_ER99DSjI7_1),.clk(gclk));
	jdff dff_B_iojmpH570_1(.din(w_dff_B_ER99DSjI7_1),.dout(w_dff_B_iojmpH570_1),.clk(gclk));
	jdff dff_B_XsQtfZjz4_0(.din(n444),.dout(w_dff_B_XsQtfZjz4_0),.clk(gclk));
	jdff dff_B_R1DgXB5Q0_1(.din(n436),.dout(w_dff_B_R1DgXB5Q0_1),.clk(gclk));
	jdff dff_A_dQT0gd6k0_0(.dout(w_n744_1[0]),.din(w_dff_A_dQT0gd6k0_0),.clk(gclk));
	jdff dff_A_HeInYmKg5_0(.dout(w_dff_A_dQT0gd6k0_0),.din(w_dff_A_HeInYmKg5_0),.clk(gclk));
	jdff dff_A_TTCvWlQS7_0(.dout(w_dff_A_HeInYmKg5_0),.din(w_dff_A_TTCvWlQS7_0),.clk(gclk));
	jdff dff_A_cWQZQc5t8_0(.dout(w_dff_A_TTCvWlQS7_0),.din(w_dff_A_cWQZQc5t8_0),.clk(gclk));
	jdff dff_A_7CWru7tZ0_0(.dout(w_dff_A_cWQZQc5t8_0),.din(w_dff_A_7CWru7tZ0_0),.clk(gclk));
	jdff dff_A_3JDVhz4W3_0(.dout(w_dff_A_7CWru7tZ0_0),.din(w_dff_A_3JDVhz4W3_0),.clk(gclk));
	jdff dff_B_k8hvkzF79_0(.din(n887),.dout(w_dff_B_k8hvkzF79_0),.clk(gclk));
	jdff dff_B_hcmCq3ie7_0(.din(w_dff_B_k8hvkzF79_0),.dout(w_dff_B_hcmCq3ie7_0),.clk(gclk));
	jdff dff_B_rRXoBqXY0_0(.din(w_dff_B_hcmCq3ie7_0),.dout(w_dff_B_rRXoBqXY0_0),.clk(gclk));
	jdff dff_B_mKbhzueB4_0(.din(w_dff_B_rRXoBqXY0_0),.dout(w_dff_B_mKbhzueB4_0),.clk(gclk));
	jdff dff_B_U4YzXz4t6_0(.din(w_dff_B_mKbhzueB4_0),.dout(w_dff_B_U4YzXz4t6_0),.clk(gclk));
	jdff dff_B_aXiWRMoZ0_0(.din(n886),.dout(w_dff_B_aXiWRMoZ0_0),.clk(gclk));
	jdff dff_B_RSx2wWa70_0(.din(w_dff_B_aXiWRMoZ0_0),.dout(w_dff_B_RSx2wWa70_0),.clk(gclk));
	jdff dff_B_1WqIVF1L6_1(.din(G127),.dout(w_dff_B_1WqIVF1L6_1),.clk(gclk));
	jdff dff_B_AIEF4ijs8_1(.din(w_dff_B_1WqIVF1L6_1),.dout(w_dff_B_AIEF4ijs8_1),.clk(gclk));
	jdff dff_A_yEEkNlvz4_1(.dout(w_n459_0[1]),.din(w_dff_A_yEEkNlvz4_1),.clk(gclk));
	jdff dff_B_Bojb8ccS4_0(.din(n458),.dout(w_dff_B_Bojb8ccS4_0),.clk(gclk));
	jdff dff_B_WBWgcu617_1(.din(n450),.dout(w_dff_B_WBWgcu617_1),.clk(gclk));
	jdff dff_B_03vhMbix5_0(.din(n1137),.dout(w_dff_B_03vhMbix5_0),.clk(gclk));
	jdff dff_B_TVKhZIYw8_0(.din(n1136),.dout(w_dff_B_TVKhZIYw8_0),.clk(gclk));
	jdff dff_B_sbx59ryn8_0(.din(w_dff_B_TVKhZIYw8_0),.dout(w_dff_B_sbx59ryn8_0),.clk(gclk));
	jdff dff_B_Qd0dIKM25_0(.din(w_dff_B_sbx59ryn8_0),.dout(w_dff_B_Qd0dIKM25_0),.clk(gclk));
	jdff dff_B_tMM8nhMj3_0(.din(w_dff_B_Qd0dIKM25_0),.dout(w_dff_B_tMM8nhMj3_0),.clk(gclk));
	jdff dff_B_IXxX6c2f0_0(.din(w_dff_B_tMM8nhMj3_0),.dout(w_dff_B_IXxX6c2f0_0),.clk(gclk));
	jdff dff_B_vuMNY9N62_0(.din(w_dff_B_IXxX6c2f0_0),.dout(w_dff_B_vuMNY9N62_0),.clk(gclk));
	jdff dff_B_TFp41Crg5_0(.din(w_dff_B_vuMNY9N62_0),.dout(w_dff_B_TFp41Crg5_0),.clk(gclk));
	jdff dff_B_zMBaP8KC5_0(.din(w_dff_B_TFp41Crg5_0),.dout(w_dff_B_zMBaP8KC5_0),.clk(gclk));
	jdff dff_B_YWk44sUP0_0(.din(w_dff_B_zMBaP8KC5_0),.dout(w_dff_B_YWk44sUP0_0),.clk(gclk));
	jdff dff_B_hy53SsrT2_0(.din(w_dff_B_YWk44sUP0_0),.dout(w_dff_B_hy53SsrT2_0),.clk(gclk));
	jdff dff_B_vO706glE4_0(.din(n1135),.dout(w_dff_B_vO706glE4_0),.clk(gclk));
	jdff dff_B_6WCAemJ45_2(.din(G146),.dout(w_dff_B_6WCAemJ45_2),.clk(gclk));
	jdff dff_B_kFVK53eQ7_2(.din(G149),.dout(w_dff_B_kFVK53eQ7_2),.clk(gclk));
	jdff dff_B_fm02c33D4_2(.din(w_dff_B_kFVK53eQ7_2),.dout(w_dff_B_fm02c33D4_2),.clk(gclk));
	jdff dff_A_iOZv9bvu4_0(.dout(w_n1002_3[0]),.din(w_dff_A_iOZv9bvu4_0),.clk(gclk));
	jdff dff_A_EhnspAGJ7_0(.dout(w_dff_A_iOZv9bvu4_0),.din(w_dff_A_EhnspAGJ7_0),.clk(gclk));
	jdff dff_A_dVVDTJGg2_0(.dout(w_dff_A_EhnspAGJ7_0),.din(w_dff_A_dVVDTJGg2_0),.clk(gclk));
	jdff dff_A_AO2Fb7lv2_0(.dout(w_dff_A_dVVDTJGg2_0),.din(w_dff_A_AO2Fb7lv2_0),.clk(gclk));
	jdff dff_A_e7w3YjiL4_1(.dout(w_n1002_3[1]),.din(w_dff_A_e7w3YjiL4_1),.clk(gclk));
	jdff dff_A_GC7RmWww4_1(.dout(w_dff_A_e7w3YjiL4_1),.din(w_dff_A_GC7RmWww4_1),.clk(gclk));
	jdff dff_B_OScALuvX8_0(.din(n826),.dout(w_dff_B_OScALuvX8_0),.clk(gclk));
	jdff dff_B_UwLl5j245_0(.din(w_dff_B_OScALuvX8_0),.dout(w_dff_B_UwLl5j245_0),.clk(gclk));
	jdff dff_B_M5SxCwSC1_0(.din(w_dff_B_UwLl5j245_0),.dout(w_dff_B_M5SxCwSC1_0),.clk(gclk));
	jdff dff_B_hiBEXKR64_0(.din(w_dff_B_M5SxCwSC1_0),.dout(w_dff_B_hiBEXKR64_0),.clk(gclk));
	jdff dff_B_q7sIJVml5_0(.din(w_dff_B_hiBEXKR64_0),.dout(w_dff_B_q7sIJVml5_0),.clk(gclk));
	jdff dff_B_pWZ8gdsS9_0(.din(n824),.dout(w_dff_B_pWZ8gdsS9_0),.clk(gclk));
	jdff dff_B_d6FpOrY91_1(.din(G130),.dout(w_dff_B_d6FpOrY91_1),.clk(gclk));
	jdff dff_B_lNEbkQDY3_1(.din(w_dff_B_d6FpOrY91_1),.dout(w_dff_B_lNEbkQDY3_1),.clk(gclk));
	jdff dff_B_qYhCDAB74_0(.din(n413),.dout(w_dff_B_qYhCDAB74_0),.clk(gclk));
	jdff dff_B_I18ZZ34v1_1(.din(n816),.dout(w_dff_B_I18ZZ34v1_1),.clk(gclk));
	jdff dff_B_nfgQw7ht0_1(.din(w_dff_B_I18ZZ34v1_1),.dout(w_dff_B_nfgQw7ht0_1),.clk(gclk));
	jdff dff_B_9iog8XGt2_1(.din(w_dff_B_nfgQw7ht0_1),.dout(w_dff_B_9iog8XGt2_1),.clk(gclk));
	jdff dff_B_YBI2nvkz0_1(.din(w_dff_B_9iog8XGt2_1),.dout(w_dff_B_YBI2nvkz0_1),.clk(gclk));
	jdff dff_B_FMUbEqxb4_1(.din(w_dff_B_YBI2nvkz0_1),.dout(w_dff_B_FMUbEqxb4_1),.clk(gclk));
	jdff dff_A_hCMC9BxT9_2(.dout(w_n744_0[2]),.din(w_dff_A_hCMC9BxT9_2),.clk(gclk));
	jdff dff_A_DcsFIBhn6_2(.dout(w_dff_A_hCMC9BxT9_2),.din(w_dff_A_DcsFIBhn6_2),.clk(gclk));
	jdff dff_A_adbeEL128_2(.dout(w_dff_A_DcsFIBhn6_2),.din(w_dff_A_adbeEL128_2),.clk(gclk));
	jdff dff_A_XnJVWyVQ2_2(.dout(w_dff_A_adbeEL128_2),.din(w_dff_A_XnJVWyVQ2_2),.clk(gclk));
	jdff dff_B_XXhSP2CH3_3(.din(n744),.dout(w_dff_B_XXhSP2CH3_3),.clk(gclk));
	jdff dff_B_792OCErl1_3(.din(w_dff_B_XXhSP2CH3_3),.dout(w_dff_B_792OCErl1_3),.clk(gclk));
	jdff dff_A_M0Pbx1Wj7_1(.dout(w_n748_3[1]),.din(w_dff_A_M0Pbx1Wj7_1),.clk(gclk));
	jdff dff_A_tiltUMDh0_1(.dout(w_dff_A_M0Pbx1Wj7_1),.din(w_dff_A_tiltUMDh0_1),.clk(gclk));
	jdff dff_A_4eAR3fuh0_2(.dout(w_n748_3[2]),.din(w_dff_A_4eAR3fuh0_2),.clk(gclk));
	jdff dff_A_cLOTdFOI4_2(.dout(w_dff_A_4eAR3fuh0_2),.din(w_dff_A_cLOTdFOI4_2),.clk(gclk));
	jdff dff_A_i977vbLG0_2(.dout(w_dff_A_cLOTdFOI4_2),.din(w_dff_A_i977vbLG0_2),.clk(gclk));
	jdff dff_A_QBdu86M61_2(.dout(w_dff_A_i977vbLG0_2),.din(w_dff_A_QBdu86M61_2),.clk(gclk));
	jdff dff_A_MMJKujt49_0(.dout(w_n999_3[0]),.din(w_dff_A_MMJKujt49_0),.clk(gclk));
	jdff dff_A_wxO2kF688_0(.dout(w_dff_A_MMJKujt49_0),.din(w_dff_A_wxO2kF688_0),.clk(gclk));
	jdff dff_A_fSFRTojg7_1(.dout(w_n999_3[1]),.din(w_dff_A_fSFRTojg7_1),.clk(gclk));
	jdff dff_B_q1g17QxW8_0(.din(n874),.dout(w_dff_B_q1g17QxW8_0),.clk(gclk));
	jdff dff_B_6AJoBFaD1_0(.din(w_dff_B_q1g17QxW8_0),.dout(w_dff_B_6AJoBFaD1_0),.clk(gclk));
	jdff dff_B_bIj9QglQ2_0(.din(w_dff_B_6AJoBFaD1_0),.dout(w_dff_B_bIj9QglQ2_0),.clk(gclk));
	jdff dff_B_NAjFVZ4G1_0(.din(w_dff_B_bIj9QglQ2_0),.dout(w_dff_B_NAjFVZ4G1_0),.clk(gclk));
	jdff dff_B_LufNUIUy5_0(.din(w_dff_B_NAjFVZ4G1_0),.dout(w_dff_B_LufNUIUy5_0),.clk(gclk));
	jdff dff_B_zG0fkk6t3_0(.din(w_dff_B_LufNUIUy5_0),.dout(w_dff_B_zG0fkk6t3_0),.clk(gclk));
	jdff dff_B_2nBctRa23_0(.din(n873),.dout(w_dff_B_2nBctRa23_0),.clk(gclk));
	jdff dff_B_7ZmmlJlu8_0(.din(w_dff_B_2nBctRa23_0),.dout(w_dff_B_7ZmmlJlu8_0),.clk(gclk));
	jdff dff_B_IJoOo9HB6_1(.din(G128),.dout(w_dff_B_IJoOo9HB6_1),.clk(gclk));
	jdff dff_B_AiJ3oHxw6_1(.din(w_dff_B_IJoOo9HB6_1),.dout(w_dff_B_AiJ3oHxw6_1),.clk(gclk));
	jdff dff_B_uuCq0Loz4_0(.din(n480),.dout(w_dff_B_uuCq0Loz4_0),.clk(gclk));
	jdff dff_B_hGD3gZm12_1(.din(n472),.dout(w_dff_B_hGD3gZm12_1),.clk(gclk));
	jdff dff_B_utGnKuzG6_0(.din(n858),.dout(w_dff_B_utGnKuzG6_0),.clk(gclk));
	jdff dff_A_1rR4Eh0M4_0(.dout(w_G4_1[0]),.din(w_dff_A_1rR4Eh0M4_0),.clk(gclk));
	jdff dff_A_6cgboUh24_0(.dout(w_dff_A_1rR4Eh0M4_0),.din(w_dff_A_6cgboUh24_0),.clk(gclk));
	jdff dff_A_AALy9F1S9_0(.dout(w_dff_A_6cgboUh24_0),.din(w_dff_A_AALy9F1S9_0),.clk(gclk));
	jdff dff_A_o1Ltpy1M8_0(.dout(w_dff_A_AALy9F1S9_0),.din(w_dff_A_o1Ltpy1M8_0),.clk(gclk));
	jdff dff_B_96mmDUl54_0(.din(n1155),.dout(w_dff_B_96mmDUl54_0),.clk(gclk));
	jdff dff_B_UiKpCWv47_0(.din(w_dff_B_96mmDUl54_0),.dout(w_dff_B_UiKpCWv47_0),.clk(gclk));
	jdff dff_B_jeIueljz0_0(.din(w_dff_B_UiKpCWv47_0),.dout(w_dff_B_jeIueljz0_0),.clk(gclk));
	jdff dff_B_ipwJyREU9_0(.din(w_dff_B_jeIueljz0_0),.dout(w_dff_B_ipwJyREU9_0),.clk(gclk));
	jdff dff_B_9QZPzyQ07_0(.din(w_dff_B_ipwJyREU9_0),.dout(w_dff_B_9QZPzyQ07_0),.clk(gclk));
	jdff dff_B_eITe9ef42_0(.din(w_dff_B_9QZPzyQ07_0),.dout(w_dff_B_eITe9ef42_0),.clk(gclk));
	jdff dff_B_RoSOetZ70_0(.din(w_dff_B_eITe9ef42_0),.dout(w_dff_B_RoSOetZ70_0),.clk(gclk));
	jdff dff_B_kY4Uz8h28_0(.din(w_dff_B_RoSOetZ70_0),.dout(w_dff_B_kY4Uz8h28_0),.clk(gclk));
	jdff dff_B_NCuvBPCh0_0(.din(w_dff_B_kY4Uz8h28_0),.dout(w_dff_B_NCuvBPCh0_0),.clk(gclk));
	jdff dff_B_kPBmYc3V6_0(.din(w_dff_B_NCuvBPCh0_0),.dout(w_dff_B_kPBmYc3V6_0),.clk(gclk));
	jdff dff_B_U1ILsJjk4_0(.din(w_dff_B_kPBmYc3V6_0),.dout(w_dff_B_U1ILsJjk4_0),.clk(gclk));
	jdff dff_B_fONYaYHu7_0(.din(w_dff_B_U1ILsJjk4_0),.dout(w_dff_B_fONYaYHu7_0),.clk(gclk));
	jdff dff_B_m3VQBE5F4_1(.din(n1148),.dout(w_dff_B_m3VQBE5F4_1),.clk(gclk));
	jdff dff_B_4vJkQoic3_1(.din(w_dff_B_m3VQBE5F4_1),.dout(w_dff_B_4vJkQoic3_1),.clk(gclk));
	jdff dff_B_fl9l574l5_1(.din(w_dff_B_4vJkQoic3_1),.dout(w_dff_B_fl9l574l5_1),.clk(gclk));
	jdff dff_B_sEsIOO6B9_1(.din(w_dff_B_fl9l574l5_1),.dout(w_dff_B_sEsIOO6B9_1),.clk(gclk));
	jdff dff_B_VlWsDQyY4_1(.din(w_dff_B_sEsIOO6B9_1),.dout(w_dff_B_VlWsDQyY4_1),.clk(gclk));
	jdff dff_B_cAWCQ3GB5_1(.din(n1150),.dout(w_dff_B_cAWCQ3GB5_1),.clk(gclk));
	jdff dff_B_hnDtYCOQ2_0(.din(n1144),.dout(w_dff_B_hnDtYCOQ2_0),.clk(gclk));
	jdff dff_B_AYvu6gyr4_0(.din(w_dff_B_hnDtYCOQ2_0),.dout(w_dff_B_AYvu6gyr4_0),.clk(gclk));
	jdff dff_B_kjfEXsjk7_0(.din(w_dff_B_AYvu6gyr4_0),.dout(w_dff_B_kjfEXsjk7_0),.clk(gclk));
	jdff dff_B_nMqtZAGB4_0(.din(w_dff_B_kjfEXsjk7_0),.dout(w_dff_B_nMqtZAGB4_0),.clk(gclk));
	jdff dff_B_ngeONwlG3_0(.din(w_dff_B_nMqtZAGB4_0),.dout(w_dff_B_ngeONwlG3_0),.clk(gclk));
	jdff dff_B_TGmimn3W9_0(.din(w_dff_B_ngeONwlG3_0),.dout(w_dff_B_TGmimn3W9_0),.clk(gclk));
	jdff dff_B_dECqJNsv0_0(.din(w_dff_B_TGmimn3W9_0),.dout(w_dff_B_dECqJNsv0_0),.clk(gclk));
	jdff dff_B_Sg9wyukl9_0(.din(w_dff_B_dECqJNsv0_0),.dout(w_dff_B_Sg9wyukl9_0),.clk(gclk));
	jdff dff_B_YamLtak89_0(.din(w_dff_B_Sg9wyukl9_0),.dout(w_dff_B_YamLtak89_0),.clk(gclk));
	jdff dff_B_M3UGxdqe8_0(.din(w_dff_B_YamLtak89_0),.dout(w_dff_B_M3UGxdqe8_0),.clk(gclk));
	jdff dff_B_3x5tHgxT4_0(.din(w_dff_B_M3UGxdqe8_0),.dout(w_dff_B_3x5tHgxT4_0),.clk(gclk));
	jdff dff_B_glttbpPm3_0(.din(w_dff_B_3x5tHgxT4_0),.dout(w_dff_B_glttbpPm3_0),.clk(gclk));
	jdff dff_B_LyayteW29_0(.din(w_dff_B_glttbpPm3_0),.dout(w_dff_B_LyayteW29_0),.clk(gclk));
	jdff dff_B_Rye43WkJ3_0(.din(w_dff_B_LyayteW29_0),.dout(w_dff_B_Rye43WkJ3_0),.clk(gclk));
	jdff dff_B_yC9Oqny89_0(.din(w_dff_B_Rye43WkJ3_0),.dout(w_dff_B_yC9Oqny89_0),.clk(gclk));
	jdff dff_B_THKPYsQ40_0(.din(w_dff_B_yC9Oqny89_0),.dout(w_dff_B_THKPYsQ40_0),.clk(gclk));
	jdff dff_B_Fdj4RatZ1_1(.din(n1141),.dout(w_dff_B_Fdj4RatZ1_1),.clk(gclk));
	jdff dff_A_hKQYqhOv9_0(.dout(w_n1142_0[0]),.din(w_dff_A_hKQYqhOv9_0),.clk(gclk));
	jdff dff_A_ka9emVfG9_0(.dout(w_dff_A_hKQYqhOv9_0),.din(w_dff_A_ka9emVfG9_0),.clk(gclk));
	jdff dff_A_uMQUu5Mt4_0(.dout(w_dff_A_ka9emVfG9_0),.din(w_dff_A_uMQUu5Mt4_0),.clk(gclk));
	jdff dff_A_zbAMO4ra6_0(.dout(w_G3717_0[0]),.din(w_dff_A_zbAMO4ra6_0),.clk(gclk));
	jdff dff_A_bBiesTm84_0(.dout(w_dff_A_zbAMO4ra6_0),.din(w_dff_A_bBiesTm84_0),.clk(gclk));
	jdff dff_A_7L3dMzNT2_0(.dout(w_dff_A_bBiesTm84_0),.din(w_dff_A_7L3dMzNT2_0),.clk(gclk));
	jdff dff_A_WcozmRnR8_0(.dout(w_dff_A_7L3dMzNT2_0),.din(w_dff_A_WcozmRnR8_0),.clk(gclk));
	jdff dff_A_AcuIn80b5_0(.dout(w_dff_A_WcozmRnR8_0),.din(w_dff_A_AcuIn80b5_0),.clk(gclk));
	jdff dff_A_EpG7ZzI35_0(.dout(w_G3724_0[0]),.din(w_dff_A_EpG7ZzI35_0),.clk(gclk));
	jdff dff_A_uVAMcr3U1_0(.dout(w_dff_A_EpG7ZzI35_0),.din(w_dff_A_uVAMcr3U1_0),.clk(gclk));
	jdff dff_A_V5wPRyCH1_0(.dout(w_dff_A_uVAMcr3U1_0),.din(w_dff_A_V5wPRyCH1_0),.clk(gclk));
	jdff dff_A_EXwBExOx4_0(.dout(w_dff_A_V5wPRyCH1_0),.din(w_dff_A_EXwBExOx4_0),.clk(gclk));
	jdff dff_A_8LXC2oEA5_2(.dout(w_G3724_0[2]),.din(w_dff_A_8LXC2oEA5_2),.clk(gclk));
	jdff dff_A_A5UoKsYg7_2(.dout(w_dff_A_8LXC2oEA5_2),.din(w_dff_A_A5UoKsYg7_2),.clk(gclk));
	jdff dff_A_wh9OqUnZ6_2(.dout(w_dff_A_A5UoKsYg7_2),.din(w_dff_A_wh9OqUnZ6_2),.clk(gclk));
	jdff dff_A_WoXRAIiC4_2(.dout(w_dff_A_wh9OqUnZ6_2),.din(w_dff_A_WoXRAIiC4_2),.clk(gclk));
	jdff dff_A_BN5s0OWO0_2(.dout(w_dff_A_WoXRAIiC4_2),.din(w_dff_A_BN5s0OWO0_2),.clk(gclk));
	jdff dff_A_QK6lzWmX6_2(.dout(w_dff_A_BN5s0OWO0_2),.din(w_dff_A_QK6lzWmX6_2),.clk(gclk));
	jdff dff_A_JbgB6ykI3_2(.dout(w_dff_A_QK6lzWmX6_2),.din(w_dff_A_JbgB6ykI3_2),.clk(gclk));
	jdff dff_A_OdBlXJcV2_2(.dout(w_dff_A_JbgB6ykI3_2),.din(w_dff_A_OdBlXJcV2_2),.clk(gclk));
	jdff dff_A_bJfjpC4g4_2(.dout(w_dff_A_OdBlXJcV2_2),.din(w_dff_A_bJfjpC4g4_2),.clk(gclk));
	jdff dff_A_fzJxdAU93_2(.dout(w_dff_A_bJfjpC4g4_2),.din(w_dff_A_fzJxdAU93_2),.clk(gclk));
	jdff dff_A_k37QSIze9_2(.dout(w_dff_A_fzJxdAU93_2),.din(w_dff_A_k37QSIze9_2),.clk(gclk));
	jdff dff_A_T2fBfKaU8_2(.dout(w_dff_A_k37QSIze9_2),.din(w_dff_A_T2fBfKaU8_2),.clk(gclk));
	jdff dff_A_RxAdn4vu3_2(.dout(w_dff_A_T2fBfKaU8_2),.din(w_dff_A_RxAdn4vu3_2),.clk(gclk));
	jdff dff_A_26IouIAS2_2(.dout(w_dff_A_RxAdn4vu3_2),.din(w_dff_A_26IouIAS2_2),.clk(gclk));
	jdff dff_A_0ilMfPlr6_2(.dout(w_dff_A_26IouIAS2_2),.din(w_dff_A_0ilMfPlr6_2),.clk(gclk));
	jdff dff_A_x8fElbcd4_2(.dout(w_dff_A_0ilMfPlr6_2),.din(w_dff_A_x8fElbcd4_2),.clk(gclk));
	jdff dff_A_8jHWSEfk2_2(.dout(w_dff_A_x8fElbcd4_2),.din(w_dff_A_8jHWSEfk2_2),.clk(gclk));
	jdff dff_A_4fATliDZ0_2(.dout(w_dff_A_8jHWSEfk2_2),.din(w_dff_A_4fATliDZ0_2),.clk(gclk));
	jdff dff_A_y4bycuRs2_0(.dout(w_G132_0[0]),.din(w_dff_A_y4bycuRs2_0),.clk(gclk));
	jdff dff_A_Gal35TrV5_0(.dout(w_dff_A_y4bycuRs2_0),.din(w_dff_A_Gal35TrV5_0),.clk(gclk));
	jdff dff_A_EzOLEFkn2_0(.dout(w_dff_A_Gal35TrV5_0),.din(w_dff_A_EzOLEFkn2_0),.clk(gclk));
	jdff dff_A_TFpmRgVb2_0(.dout(w_dff_A_EzOLEFkn2_0),.din(w_dff_A_TFpmRgVb2_0),.clk(gclk));
	jdff dff_A_hvaU3ANT8_0(.dout(w_dff_A_TFpmRgVb2_0),.din(w_dff_A_hvaU3ANT8_0),.clk(gclk));
	jdff dff_A_Bu5SEptC9_0(.dout(w_dff_A_hvaU3ANT8_0),.din(w_dff_A_Bu5SEptC9_0),.clk(gclk));
	jdff dff_A_jybOjyyD6_0(.dout(w_dff_A_Bu5SEptC9_0),.din(w_dff_A_jybOjyyD6_0),.clk(gclk));
	jdff dff_A_KmaIF2qp6_0(.dout(w_dff_A_jybOjyyD6_0),.din(w_dff_A_KmaIF2qp6_0),.clk(gclk));
	jdff dff_A_FRUcta711_0(.dout(w_dff_A_KmaIF2qp6_0),.din(w_dff_A_FRUcta711_0),.clk(gclk));
	jdff dff_A_kvGKwaR46_0(.dout(w_dff_A_FRUcta711_0),.din(w_dff_A_kvGKwaR46_0),.clk(gclk));
	jdff dff_A_rE3kG1Y35_0(.dout(w_dff_A_kvGKwaR46_0),.din(w_dff_A_rE3kG1Y35_0),.clk(gclk));
	jdff dff_A_kbfB5rmE9_0(.dout(w_dff_A_rE3kG1Y35_0),.din(w_dff_A_kbfB5rmE9_0),.clk(gclk));
	jdff dff_A_KPZKUBKl8_0(.dout(w_dff_A_kbfB5rmE9_0),.din(w_dff_A_KPZKUBKl8_0),.clk(gclk));
	jdff dff_B_8BN9JgJr4_2(.din(G132),.dout(w_dff_B_8BN9JgJr4_2),.clk(gclk));
	jdff dff_B_G0tIU59Z0_2(.din(w_dff_B_8BN9JgJr4_2),.dout(w_dff_B_G0tIU59Z0_2),.clk(gclk));
	jdff dff_B_nD7b9jDc3_2(.din(w_dff_B_G0tIU59Z0_2),.dout(w_dff_B_nD7b9jDc3_2),.clk(gclk));
	jdff dff_B_kEvZGrFN3_1(.din(n1184),.dout(w_dff_B_kEvZGrFN3_1),.clk(gclk));
	jdff dff_B_vVo6NpYO0_0(.din(n1189),.dout(w_dff_B_vVo6NpYO0_0),.clk(gclk));
	jdff dff_B_NIssC7zS7_0(.din(w_dff_B_vVo6NpYO0_0),.dout(w_dff_B_NIssC7zS7_0),.clk(gclk));
	jdff dff_B_ZPdVBZ620_0(.din(n1187),.dout(w_dff_B_ZPdVBZ620_0),.clk(gclk));
	jdff dff_A_hKPwJCt40_0(.dout(w_G601_0),.din(w_dff_A_hKPwJCt40_0),.clk(gclk));
	jdff dff_B_omv28N7A3_1(.din(n656),.dout(w_dff_B_omv28N7A3_1),.clk(gclk));
	jdff dff_A_eGI5ioL92_0(.dout(w_n671_0[0]),.din(w_dff_A_eGI5ioL92_0),.clk(gclk));
	jdff dff_B_8xlMiN679_1(.din(n665),.dout(w_dff_B_8xlMiN679_1),.clk(gclk));
	jdff dff_B_UImnMwAf3_1(.din(n907),.dout(w_dff_B_UImnMwAf3_1),.clk(gclk));
	jdff dff_B_53V4VH5V2_1(.din(n909),.dout(w_dff_B_53V4VH5V2_1),.clk(gclk));
	jdff dff_B_Wzx6zhX68_1(.din(w_dff_B_53V4VH5V2_1),.dout(w_dff_B_Wzx6zhX68_1),.clk(gclk));
	jdff dff_B_0kxmv4TN6_0(.din(n910),.dout(w_dff_B_0kxmv4TN6_0),.clk(gclk));
	jdff dff_B_zdUxXCoH5_1(.din(n908),.dout(w_dff_B_zdUxXCoH5_1),.clk(gclk));
	jdff dff_B_bNOwwZgX8_0(.din(n904),.dout(w_dff_B_bNOwwZgX8_0),.clk(gclk));
	jdff dff_A_OkzrOEWX9_0(.dout(w_G369_0[0]),.din(w_dff_A_OkzrOEWX9_0),.clk(gclk));
	jdff dff_A_7UBBPQTy7_0(.dout(w_n621_1[0]),.din(w_dff_A_7UBBPQTy7_0),.clk(gclk));
	jdff dff_A_Af7aqnpx1_0(.dout(w_dff_A_7UBBPQTy7_0),.din(w_dff_A_Af7aqnpx1_0),.clk(gclk));
	jdff dff_A_ZcjTCanV9_0(.dout(w_dff_A_Af7aqnpx1_0),.din(w_dff_A_ZcjTCanV9_0),.clk(gclk));
	jdff dff_B_Njv8LDIf3_0(.din(n921),.dout(w_dff_B_Njv8LDIf3_0),.clk(gclk));
	jdff dff_A_4T8SEnOh4_0(.dout(w_G289_0[0]),.din(w_dff_A_4T8SEnOh4_0),.clk(gclk));
	jdff dff_B_5hsqcOvn3_0(.din(n1224),.dout(w_dff_B_5hsqcOvn3_0),.clk(gclk));
	jdff dff_B_gnQGsW5I5_0(.din(w_dff_B_5hsqcOvn3_0),.dout(w_dff_B_gnQGsW5I5_0),.clk(gclk));
	jdff dff_B_khqqblDa1_0(.din(w_dff_B_gnQGsW5I5_0),.dout(w_dff_B_khqqblDa1_0),.clk(gclk));
	jdff dff_B_ciRoZKue4_0(.din(w_dff_B_khqqblDa1_0),.dout(w_dff_B_ciRoZKue4_0),.clk(gclk));
	jdff dff_B_2xmnb8An4_0(.din(w_dff_B_ciRoZKue4_0),.dout(w_dff_B_2xmnb8An4_0),.clk(gclk));
	jdff dff_B_Z4vWh6kn7_0(.din(w_dff_B_2xmnb8An4_0),.dout(w_dff_B_Z4vWh6kn7_0),.clk(gclk));
	jdff dff_B_4PxaYOTQ7_0(.din(w_dff_B_Z4vWh6kn7_0),.dout(w_dff_B_4PxaYOTQ7_0),.clk(gclk));
	jdff dff_B_fptPdpyV5_0(.din(w_dff_B_4PxaYOTQ7_0),.dout(w_dff_B_fptPdpyV5_0),.clk(gclk));
	jdff dff_B_2UbHNWf24_0(.din(w_dff_B_fptPdpyV5_0),.dout(w_dff_B_2UbHNWf24_0),.clk(gclk));
	jdff dff_B_um3yBCOh7_0(.din(w_dff_B_2UbHNWf24_0),.dout(w_dff_B_um3yBCOh7_0),.clk(gclk));
	jdff dff_B_NSlHX2uf2_0(.din(w_dff_B_um3yBCOh7_0),.dout(w_dff_B_NSlHX2uf2_0),.clk(gclk));
	jdff dff_B_cIQsVOIZ9_0(.din(w_dff_B_NSlHX2uf2_0),.dout(w_dff_B_cIQsVOIZ9_0),.clk(gclk));
	jdff dff_B_Mu3dFL2x7_0(.din(w_dff_B_cIQsVOIZ9_0),.dout(w_dff_B_Mu3dFL2x7_0),.clk(gclk));
	jdff dff_B_s8tlO6rJ5_0(.din(w_dff_B_Mu3dFL2x7_0),.dout(w_dff_B_s8tlO6rJ5_0),.clk(gclk));
	jdff dff_B_oZvyQe5e2_0(.din(w_dff_B_s8tlO6rJ5_0),.dout(w_dff_B_oZvyQe5e2_0),.clk(gclk));
	jdff dff_B_oq6JPoJK9_0(.din(w_dff_B_oZvyQe5e2_0),.dout(w_dff_B_oq6JPoJK9_0),.clk(gclk));
	jdff dff_B_fE20assw7_0(.din(w_dff_B_oq6JPoJK9_0),.dout(w_dff_B_fE20assw7_0),.clk(gclk));
	jdff dff_B_QXWGfaW84_0(.din(n1223),.dout(w_dff_B_QXWGfaW84_0),.clk(gclk));
	jdff dff_B_F8m6nLQa7_0(.din(n1231),.dout(w_dff_B_F8m6nLQa7_0),.clk(gclk));
	jdff dff_B_GQ0PLVdF9_0(.din(w_dff_B_F8m6nLQa7_0),.dout(w_dff_B_GQ0PLVdF9_0),.clk(gclk));
	jdff dff_B_ntpr1OrJ8_0(.din(w_dff_B_GQ0PLVdF9_0),.dout(w_dff_B_ntpr1OrJ8_0),.clk(gclk));
	jdff dff_B_rrzqkxJX2_0(.din(w_dff_B_ntpr1OrJ8_0),.dout(w_dff_B_rrzqkxJX2_0),.clk(gclk));
	jdff dff_B_UsKTbJOH2_0(.din(w_dff_B_rrzqkxJX2_0),.dout(w_dff_B_UsKTbJOH2_0),.clk(gclk));
	jdff dff_B_U57Tn4OJ6_0(.din(w_dff_B_UsKTbJOH2_0),.dout(w_dff_B_U57Tn4OJ6_0),.clk(gclk));
	jdff dff_B_ygJarYfs0_0(.din(w_dff_B_U57Tn4OJ6_0),.dout(w_dff_B_ygJarYfs0_0),.clk(gclk));
	jdff dff_B_7UBwKGAW8_0(.din(w_dff_B_ygJarYfs0_0),.dout(w_dff_B_7UBwKGAW8_0),.clk(gclk));
	jdff dff_B_nScdvI9E7_0(.din(w_dff_B_7UBwKGAW8_0),.dout(w_dff_B_nScdvI9E7_0),.clk(gclk));
	jdff dff_B_zjTkoiaA0_0(.din(w_dff_B_nScdvI9E7_0),.dout(w_dff_B_zjTkoiaA0_0),.clk(gclk));
	jdff dff_B_OcSfrWjB7_0(.din(w_dff_B_zjTkoiaA0_0),.dout(w_dff_B_OcSfrWjB7_0),.clk(gclk));
	jdff dff_B_k6dFFJ5d9_0(.din(w_dff_B_OcSfrWjB7_0),.dout(w_dff_B_k6dFFJ5d9_0),.clk(gclk));
	jdff dff_B_eE9BHOiQ4_0(.din(w_dff_B_k6dFFJ5d9_0),.dout(w_dff_B_eE9BHOiQ4_0),.clk(gclk));
	jdff dff_B_Dperetc79_0(.din(w_dff_B_eE9BHOiQ4_0),.dout(w_dff_B_Dperetc79_0),.clk(gclk));
	jdff dff_B_qxKUMI2s8_0(.din(w_dff_B_Dperetc79_0),.dout(w_dff_B_qxKUMI2s8_0),.clk(gclk));
	jdff dff_B_Z2kCsBUf6_0(.din(w_dff_B_qxKUMI2s8_0),.dout(w_dff_B_Z2kCsBUf6_0),.clk(gclk));
	jdff dff_B_eUoyMdux2_0(.din(w_dff_B_Z2kCsBUf6_0),.dout(w_dff_B_eUoyMdux2_0),.clk(gclk));
	jdff dff_B_lrLLoZaM8_0(.din(n1230),.dout(w_dff_B_lrLLoZaM8_0),.clk(gclk));
	jdff dff_B_UeAhgxOY3_2(.din(G106),.dout(w_dff_B_UeAhgxOY3_2),.clk(gclk));
	jdff dff_B_4zTjIPSx3_2(.din(G109),.dout(w_dff_B_4zTjIPSx3_2),.clk(gclk));
	jdff dff_B_KBen70oB1_2(.din(w_dff_B_4zTjIPSx3_2),.dout(w_dff_B_KBen70oB1_2),.clk(gclk));
	jdff dff_B_IJbKMdYW1_0(.din(n1239),.dout(w_dff_B_IJbKMdYW1_0),.clk(gclk));
	jdff dff_B_LMt06rRg9_0(.din(w_dff_B_IJbKMdYW1_0),.dout(w_dff_B_LMt06rRg9_0),.clk(gclk));
	jdff dff_B_UP1AnLUt5_0(.din(w_dff_B_LMt06rRg9_0),.dout(w_dff_B_UP1AnLUt5_0),.clk(gclk));
	jdff dff_B_ELToS6ad7_0(.din(w_dff_B_UP1AnLUt5_0),.dout(w_dff_B_ELToS6ad7_0),.clk(gclk));
	jdff dff_B_bZk81CwM9_0(.din(w_dff_B_ELToS6ad7_0),.dout(w_dff_B_bZk81CwM9_0),.clk(gclk));
	jdff dff_B_ofGUW5RS3_0(.din(w_dff_B_bZk81CwM9_0),.dout(w_dff_B_ofGUW5RS3_0),.clk(gclk));
	jdff dff_B_1e2K5l962_0(.din(w_dff_B_ofGUW5RS3_0),.dout(w_dff_B_1e2K5l962_0),.clk(gclk));
	jdff dff_B_49xixjr13_0(.din(w_dff_B_1e2K5l962_0),.dout(w_dff_B_49xixjr13_0),.clk(gclk));
	jdff dff_B_2Jrakhrj6_0(.din(w_dff_B_49xixjr13_0),.dout(w_dff_B_2Jrakhrj6_0),.clk(gclk));
	jdff dff_B_p02BTYxB6_0(.din(w_dff_B_2Jrakhrj6_0),.dout(w_dff_B_p02BTYxB6_0),.clk(gclk));
	jdff dff_B_YPMqT73X3_0(.din(w_dff_B_p02BTYxB6_0),.dout(w_dff_B_YPMqT73X3_0),.clk(gclk));
	jdff dff_B_7jP2SkIc2_0(.din(w_dff_B_YPMqT73X3_0),.dout(w_dff_B_7jP2SkIc2_0),.clk(gclk));
	jdff dff_B_hvtHPjWP6_0(.din(w_dff_B_7jP2SkIc2_0),.dout(w_dff_B_hvtHPjWP6_0),.clk(gclk));
	jdff dff_B_0kRqpW4z8_0(.din(w_dff_B_hvtHPjWP6_0),.dout(w_dff_B_0kRqpW4z8_0),.clk(gclk));
	jdff dff_B_pa2Z2kjW5_0(.din(w_dff_B_0kRqpW4z8_0),.dout(w_dff_B_pa2Z2kjW5_0),.clk(gclk));
	jdff dff_B_0JrtqFgk8_0(.din(w_dff_B_pa2Z2kjW5_0),.dout(w_dff_B_0JrtqFgk8_0),.clk(gclk));
	jdff dff_B_Foucat1g1_0(.din(n1238),.dout(w_dff_B_Foucat1g1_0),.clk(gclk));
	jdff dff_B_tyhcO2867_0(.din(n1248),.dout(w_dff_B_tyhcO2867_0),.clk(gclk));
	jdff dff_B_oceMWlqv0_0(.din(w_dff_B_tyhcO2867_0),.dout(w_dff_B_oceMWlqv0_0),.clk(gclk));
	jdff dff_B_xDaQlDmY9_0(.din(w_dff_B_oceMWlqv0_0),.dout(w_dff_B_xDaQlDmY9_0),.clk(gclk));
	jdff dff_B_YihmyH3A4_0(.din(w_dff_B_xDaQlDmY9_0),.dout(w_dff_B_YihmyH3A4_0),.clk(gclk));
	jdff dff_B_UmWlof7l5_0(.din(w_dff_B_YihmyH3A4_0),.dout(w_dff_B_UmWlof7l5_0),.clk(gclk));
	jdff dff_B_oqUcqDfa8_0(.din(w_dff_B_UmWlof7l5_0),.dout(w_dff_B_oqUcqDfa8_0),.clk(gclk));
	jdff dff_B_3t7SR3Ek3_0(.din(w_dff_B_oqUcqDfa8_0),.dout(w_dff_B_3t7SR3Ek3_0),.clk(gclk));
	jdff dff_B_neTNoa0G6_0(.din(w_dff_B_3t7SR3Ek3_0),.dout(w_dff_B_neTNoa0G6_0),.clk(gclk));
	jdff dff_B_qn2hLOcN9_0(.din(w_dff_B_neTNoa0G6_0),.dout(w_dff_B_qn2hLOcN9_0),.clk(gclk));
	jdff dff_B_2okZtWdb2_0(.din(w_dff_B_qn2hLOcN9_0),.dout(w_dff_B_2okZtWdb2_0),.clk(gclk));
	jdff dff_B_EgSggrT63_0(.din(w_dff_B_2okZtWdb2_0),.dout(w_dff_B_EgSggrT63_0),.clk(gclk));
	jdff dff_B_jwmbYkEd7_0(.din(w_dff_B_EgSggrT63_0),.dout(w_dff_B_jwmbYkEd7_0),.clk(gclk));
	jdff dff_B_HXv8tPOX6_0(.din(w_dff_B_jwmbYkEd7_0),.dout(w_dff_B_HXv8tPOX6_0),.clk(gclk));
	jdff dff_B_fPpETqz82_0(.din(w_dff_B_HXv8tPOX6_0),.dout(w_dff_B_fPpETqz82_0),.clk(gclk));
	jdff dff_B_HaCTnfuG9_0(.din(w_dff_B_fPpETqz82_0),.dout(w_dff_B_HaCTnfuG9_0),.clk(gclk));
	jdff dff_B_qiaSDrf53_0(.din(w_dff_B_HaCTnfuG9_0),.dout(w_dff_B_qiaSDrf53_0),.clk(gclk));
	jdff dff_B_3LcSg0uW3_0(.din(n1247),.dout(w_dff_B_3LcSg0uW3_0),.clk(gclk));
	jdff dff_A_4KE5DLLY1_2(.dout(w_n797_2[2]),.din(w_dff_A_4KE5DLLY1_2),.clk(gclk));
	jdff dff_A_DvvXWMSC4_2(.dout(w_n793_2[2]),.din(w_dff_A_DvvXWMSC4_2),.clk(gclk));
	jdff dff_B_WvUzs1Ts3_0(.din(n1257),.dout(w_dff_B_WvUzs1Ts3_0),.clk(gclk));
	jdff dff_B_f2ZpQjlX1_0(.din(w_dff_B_WvUzs1Ts3_0),.dout(w_dff_B_f2ZpQjlX1_0),.clk(gclk));
	jdff dff_B_WejA4FLu8_0(.din(w_dff_B_f2ZpQjlX1_0),.dout(w_dff_B_WejA4FLu8_0),.clk(gclk));
	jdff dff_B_6YRv9iKj6_0(.din(w_dff_B_WejA4FLu8_0),.dout(w_dff_B_6YRv9iKj6_0),.clk(gclk));
	jdff dff_B_wbheDars5_0(.din(w_dff_B_6YRv9iKj6_0),.dout(w_dff_B_wbheDars5_0),.clk(gclk));
	jdff dff_B_oERyJoSr0_0(.din(w_dff_B_wbheDars5_0),.dout(w_dff_B_oERyJoSr0_0),.clk(gclk));
	jdff dff_B_BdTLhuto8_0(.din(w_dff_B_oERyJoSr0_0),.dout(w_dff_B_BdTLhuto8_0),.clk(gclk));
	jdff dff_B_7j6kMCPl8_0(.din(w_dff_B_BdTLhuto8_0),.dout(w_dff_B_7j6kMCPl8_0),.clk(gclk));
	jdff dff_B_4I4tqIYh2_0(.din(w_dff_B_7j6kMCPl8_0),.dout(w_dff_B_4I4tqIYh2_0),.clk(gclk));
	jdff dff_B_VPFnzmRM6_0(.din(w_dff_B_4I4tqIYh2_0),.dout(w_dff_B_VPFnzmRM6_0),.clk(gclk));
	jdff dff_B_NMHZGI2e2_0(.din(w_dff_B_VPFnzmRM6_0),.dout(w_dff_B_NMHZGI2e2_0),.clk(gclk));
	jdff dff_B_SHPW11385_0(.din(w_dff_B_NMHZGI2e2_0),.dout(w_dff_B_SHPW11385_0),.clk(gclk));
	jdff dff_B_x0tl3HEi2_0(.din(w_dff_B_SHPW11385_0),.dout(w_dff_B_x0tl3HEi2_0),.clk(gclk));
	jdff dff_B_v0zLj5Od4_0(.din(w_dff_B_x0tl3HEi2_0),.dout(w_dff_B_v0zLj5Od4_0),.clk(gclk));
	jdff dff_B_1xKtCMCP1_0(.din(w_dff_B_v0zLj5Od4_0),.dout(w_dff_B_1xKtCMCP1_0),.clk(gclk));
	jdff dff_B_K4fKwws38_0(.din(n1256),.dout(w_dff_B_K4fKwws38_0),.clk(gclk));
	jdff dff_B_LaUmfTSg0_0(.din(n1264),.dout(w_dff_B_LaUmfTSg0_0),.clk(gclk));
	jdff dff_B_OWl8EKew6_0(.din(w_dff_B_LaUmfTSg0_0),.dout(w_dff_B_OWl8EKew6_0),.clk(gclk));
	jdff dff_B_mOU4ExbL6_0(.din(w_dff_B_OWl8EKew6_0),.dout(w_dff_B_mOU4ExbL6_0),.clk(gclk));
	jdff dff_B_zsL91hBh6_0(.din(w_dff_B_mOU4ExbL6_0),.dout(w_dff_B_zsL91hBh6_0),.clk(gclk));
	jdff dff_B_WxKpJivV8_0(.din(w_dff_B_zsL91hBh6_0),.dout(w_dff_B_WxKpJivV8_0),.clk(gclk));
	jdff dff_B_8XrXzZY87_0(.din(w_dff_B_WxKpJivV8_0),.dout(w_dff_B_8XrXzZY87_0),.clk(gclk));
	jdff dff_B_AZqvnguG5_0(.din(w_dff_B_8XrXzZY87_0),.dout(w_dff_B_AZqvnguG5_0),.clk(gclk));
	jdff dff_B_eBZ5pvxp1_0(.din(w_dff_B_AZqvnguG5_0),.dout(w_dff_B_eBZ5pvxp1_0),.clk(gclk));
	jdff dff_B_ttVhzxHJ5_0(.din(w_dff_B_eBZ5pvxp1_0),.dout(w_dff_B_ttVhzxHJ5_0),.clk(gclk));
	jdff dff_B_QauO95Rq0_0(.din(w_dff_B_ttVhzxHJ5_0),.dout(w_dff_B_QauO95Rq0_0),.clk(gclk));
	jdff dff_B_qXkdGEae9_0(.din(w_dff_B_QauO95Rq0_0),.dout(w_dff_B_qXkdGEae9_0),.clk(gclk));
	jdff dff_B_efeCm2R40_0(.din(w_dff_B_qXkdGEae9_0),.dout(w_dff_B_efeCm2R40_0),.clk(gclk));
	jdff dff_B_leDKtqH27_0(.din(w_dff_B_efeCm2R40_0),.dout(w_dff_B_leDKtqH27_0),.clk(gclk));
	jdff dff_B_h0OPKYgB1_0(.din(w_dff_B_leDKtqH27_0),.dout(w_dff_B_h0OPKYgB1_0),.clk(gclk));
	jdff dff_B_szqEZaur3_0(.din(w_dff_B_h0OPKYgB1_0),.dout(w_dff_B_szqEZaur3_0),.clk(gclk));
	jdff dff_B_HfR9NiRb5_0(.din(w_dff_B_szqEZaur3_0),.dout(w_dff_B_HfR9NiRb5_0),.clk(gclk));
	jdff dff_B_8DjwxO8J4_0(.din(n1263),.dout(w_dff_B_8DjwxO8J4_0),.clk(gclk));
	jdff dff_B_LY7NLxU77_2(.din(G49),.dout(w_dff_B_LY7NLxU77_2),.clk(gclk));
	jdff dff_B_7lNTWjgU2_2(.din(G46),.dout(w_dff_B_7lNTWjgU2_2),.clk(gclk));
	jdff dff_B_agihHWfT0_2(.din(w_dff_B_7lNTWjgU2_2),.dout(w_dff_B_agihHWfT0_2),.clk(gclk));
	jdff dff_B_Dsi6kEVv0_0(.din(n1271),.dout(w_dff_B_Dsi6kEVv0_0),.clk(gclk));
	jdff dff_B_caSoMYmE9_0(.din(w_dff_B_Dsi6kEVv0_0),.dout(w_dff_B_caSoMYmE9_0),.clk(gclk));
	jdff dff_B_6picSZTO7_0(.din(w_dff_B_caSoMYmE9_0),.dout(w_dff_B_6picSZTO7_0),.clk(gclk));
	jdff dff_B_1WIk8esE8_0(.din(w_dff_B_6picSZTO7_0),.dout(w_dff_B_1WIk8esE8_0),.clk(gclk));
	jdff dff_B_H6Ku1xD71_0(.din(w_dff_B_1WIk8esE8_0),.dout(w_dff_B_H6Ku1xD71_0),.clk(gclk));
	jdff dff_B_KYqGTzkz7_0(.din(w_dff_B_H6Ku1xD71_0),.dout(w_dff_B_KYqGTzkz7_0),.clk(gclk));
	jdff dff_B_89eBLgjP3_0(.din(w_dff_B_KYqGTzkz7_0),.dout(w_dff_B_89eBLgjP3_0),.clk(gclk));
	jdff dff_B_2YMC2gyN5_0(.din(w_dff_B_89eBLgjP3_0),.dout(w_dff_B_2YMC2gyN5_0),.clk(gclk));
	jdff dff_B_CKx8PJfx1_0(.din(w_dff_B_2YMC2gyN5_0),.dout(w_dff_B_CKx8PJfx1_0),.clk(gclk));
	jdff dff_B_ZFAo4mrR0_0(.din(w_dff_B_CKx8PJfx1_0),.dout(w_dff_B_ZFAo4mrR0_0),.clk(gclk));
	jdff dff_B_JvpU8GmB3_0(.din(w_dff_B_ZFAo4mrR0_0),.dout(w_dff_B_JvpU8GmB3_0),.clk(gclk));
	jdff dff_B_GUVV8PFt9_0(.din(w_dff_B_JvpU8GmB3_0),.dout(w_dff_B_GUVV8PFt9_0),.clk(gclk));
	jdff dff_B_RZIRIXk37_0(.din(w_dff_B_GUVV8PFt9_0),.dout(w_dff_B_RZIRIXk37_0),.clk(gclk));
	jdff dff_B_GZVaPspF7_0(.din(w_dff_B_RZIRIXk37_0),.dout(w_dff_B_GZVaPspF7_0),.clk(gclk));
	jdff dff_B_ILMNY9yM7_0(.din(w_dff_B_GZVaPspF7_0),.dout(w_dff_B_ILMNY9yM7_0),.clk(gclk));
	jdff dff_B_jgcc0Xlp3_0(.din(w_dff_B_ILMNY9yM7_0),.dout(w_dff_B_jgcc0Xlp3_0),.clk(gclk));
	jdff dff_B_p0dtSfDh5_0(.din(n1270),.dout(w_dff_B_p0dtSfDh5_0),.clk(gclk));
	jdff dff_B_fJylF7gT3_2(.din(G103),.dout(w_dff_B_fJylF7gT3_2),.clk(gclk));
	jdff dff_B_xZvxPhuO3_2(.din(G100),.dout(w_dff_B_xZvxPhuO3_2),.clk(gclk));
	jdff dff_B_o5pLiG8c7_2(.din(w_dff_B_xZvxPhuO3_2),.dout(w_dff_B_o5pLiG8c7_2),.clk(gclk));
	jdff dff_A_HPZV4S169_2(.dout(w_n843_2[2]),.din(w_dff_A_HPZV4S169_2),.clk(gclk));
	jdff dff_A_JkQzaEnP2_2(.dout(w_n840_2[2]),.din(w_dff_A_JkQzaEnP2_2),.clk(gclk));
	jdff dff_B_TlPbYDHg5_0(.din(n1278),.dout(w_dff_B_TlPbYDHg5_0),.clk(gclk));
	jdff dff_B_VynV79Ea6_0(.din(w_dff_B_TlPbYDHg5_0),.dout(w_dff_B_VynV79Ea6_0),.clk(gclk));
	jdff dff_B_SSIgrztB6_0(.din(w_dff_B_VynV79Ea6_0),.dout(w_dff_B_SSIgrztB6_0),.clk(gclk));
	jdff dff_B_UvqLAqdy1_0(.din(w_dff_B_SSIgrztB6_0),.dout(w_dff_B_UvqLAqdy1_0),.clk(gclk));
	jdff dff_B_ssxuIrBs2_0(.din(w_dff_B_UvqLAqdy1_0),.dout(w_dff_B_ssxuIrBs2_0),.clk(gclk));
	jdff dff_B_U7oIt5kt7_0(.din(w_dff_B_ssxuIrBs2_0),.dout(w_dff_B_U7oIt5kt7_0),.clk(gclk));
	jdff dff_B_lfh1lHlH3_0(.din(w_dff_B_U7oIt5kt7_0),.dout(w_dff_B_lfh1lHlH3_0),.clk(gclk));
	jdff dff_B_ts0cGKd99_0(.din(w_dff_B_lfh1lHlH3_0),.dout(w_dff_B_ts0cGKd99_0),.clk(gclk));
	jdff dff_B_J7em22F56_0(.din(w_dff_B_ts0cGKd99_0),.dout(w_dff_B_J7em22F56_0),.clk(gclk));
	jdff dff_B_fRMhin913_0(.din(w_dff_B_J7em22F56_0),.dout(w_dff_B_fRMhin913_0),.clk(gclk));
	jdff dff_B_paT4gHN20_0(.din(w_dff_B_fRMhin913_0),.dout(w_dff_B_paT4gHN20_0),.clk(gclk));
	jdff dff_B_P1oVGmOm4_0(.din(w_dff_B_paT4gHN20_0),.dout(w_dff_B_P1oVGmOm4_0),.clk(gclk));
	jdff dff_B_mqNFGYbA8_0(.din(w_dff_B_P1oVGmOm4_0),.dout(w_dff_B_mqNFGYbA8_0),.clk(gclk));
	jdff dff_B_QWeznXfG3_0(.din(w_dff_B_mqNFGYbA8_0),.dout(w_dff_B_QWeznXfG3_0),.clk(gclk));
	jdff dff_B_4ZPfSibY8_0(.din(w_dff_B_QWeznXfG3_0),.dout(w_dff_B_4ZPfSibY8_0),.clk(gclk));
	jdff dff_B_2V4gCxYY5_0(.din(n1277),.dout(w_dff_B_2V4gCxYY5_0),.clk(gclk));
	jdff dff_B_9XFcTKAY6_2(.din(G40),.dout(w_dff_B_9XFcTKAY6_2),.clk(gclk));
	jdff dff_B_d6P1H7FR3_2(.din(G91),.dout(w_dff_B_d6P1H7FR3_2),.clk(gclk));
	jdff dff_B_daimAzmN6_2(.din(w_dff_B_d6P1H7FR3_2),.dout(w_dff_B_daimAzmN6_2),.clk(gclk));
	jdff dff_B_bW8KinqO0_0(.din(n1285),.dout(w_dff_B_bW8KinqO0_0),.clk(gclk));
	jdff dff_B_iktnIL0L6_0(.din(w_dff_B_bW8KinqO0_0),.dout(w_dff_B_iktnIL0L6_0),.clk(gclk));
	jdff dff_B_M5BWNTpH4_0(.din(w_dff_B_iktnIL0L6_0),.dout(w_dff_B_M5BWNTpH4_0),.clk(gclk));
	jdff dff_B_uYjMGAgs6_0(.din(w_dff_B_M5BWNTpH4_0),.dout(w_dff_B_uYjMGAgs6_0),.clk(gclk));
	jdff dff_B_QfF1cgp14_0(.din(w_dff_B_uYjMGAgs6_0),.dout(w_dff_B_QfF1cgp14_0),.clk(gclk));
	jdff dff_B_j4yw23zc2_0(.din(w_dff_B_QfF1cgp14_0),.dout(w_dff_B_j4yw23zc2_0),.clk(gclk));
	jdff dff_B_HCPl31yi7_0(.din(w_dff_B_j4yw23zc2_0),.dout(w_dff_B_HCPl31yi7_0),.clk(gclk));
	jdff dff_B_YtYQyY3I9_0(.din(w_dff_B_HCPl31yi7_0),.dout(w_dff_B_YtYQyY3I9_0),.clk(gclk));
	jdff dff_B_rHCZqgn79_0(.din(w_dff_B_YtYQyY3I9_0),.dout(w_dff_B_rHCZqgn79_0),.clk(gclk));
	jdff dff_B_3SShvQfM7_0(.din(w_dff_B_rHCZqgn79_0),.dout(w_dff_B_3SShvQfM7_0),.clk(gclk));
	jdff dff_B_IU2UfoME2_0(.din(w_dff_B_3SShvQfM7_0),.dout(w_dff_B_IU2UfoME2_0),.clk(gclk));
	jdff dff_B_I9D5SnTh6_0(.din(w_dff_B_IU2UfoME2_0),.dout(w_dff_B_I9D5SnTh6_0),.clk(gclk));
	jdff dff_B_PDGODrkG7_0(.din(w_dff_B_I9D5SnTh6_0),.dout(w_dff_B_PDGODrkG7_0),.clk(gclk));
	jdff dff_B_jHhMLNMw5_0(.din(w_dff_B_PDGODrkG7_0),.dout(w_dff_B_jHhMLNMw5_0),.clk(gclk));
	jdff dff_B_kCrwhqOF3_0(.din(w_dff_B_jHhMLNMw5_0),.dout(w_dff_B_kCrwhqOF3_0),.clk(gclk));
	jdff dff_B_CLS7VxaR5_0(.din(n1284),.dout(w_dff_B_CLS7VxaR5_0),.clk(gclk));
	jdff dff_A_8LjImTsb6_0(.dout(w_G137_6[0]),.din(w_dff_A_8LjImTsb6_0),.clk(gclk));
	jdff dff_A_Le83ZYs52_0(.dout(w_dff_A_8LjImTsb6_0),.din(w_dff_A_Le83ZYs52_0),.clk(gclk));
	jdff dff_A_S2HGctti1_0(.dout(w_dff_A_Le83ZYs52_0),.din(w_dff_A_S2HGctti1_0),.clk(gclk));
	jdff dff_A_oXqaLl9T1_0(.dout(w_dff_A_S2HGctti1_0),.din(w_dff_A_oXqaLl9T1_0),.clk(gclk));
	jdff dff_A_PNqV6Qcx1_0(.dout(w_dff_A_oXqaLl9T1_0),.din(w_dff_A_PNqV6Qcx1_0),.clk(gclk));
	jdff dff_A_pQ3EGlQh9_1(.dout(w_G137_6[1]),.din(w_dff_A_pQ3EGlQh9_1),.clk(gclk));
	jdff dff_B_7sZ77vpw0_0(.din(n1293),.dout(w_dff_B_7sZ77vpw0_0),.clk(gclk));
	jdff dff_B_gQVib5Ky2_0(.din(w_dff_B_7sZ77vpw0_0),.dout(w_dff_B_gQVib5Ky2_0),.clk(gclk));
	jdff dff_B_zDvvXsdD3_0(.din(w_dff_B_gQVib5Ky2_0),.dout(w_dff_B_zDvvXsdD3_0),.clk(gclk));
	jdff dff_B_3uUhCogx3_0(.din(w_dff_B_zDvvXsdD3_0),.dout(w_dff_B_3uUhCogx3_0),.clk(gclk));
	jdff dff_B_6sKEyhKr3_0(.din(w_dff_B_3uUhCogx3_0),.dout(w_dff_B_6sKEyhKr3_0),.clk(gclk));
	jdff dff_B_3XfNGyaC8_0(.din(w_dff_B_6sKEyhKr3_0),.dout(w_dff_B_3XfNGyaC8_0),.clk(gclk));
	jdff dff_B_m9Xf2G8T3_0(.din(w_dff_B_3XfNGyaC8_0),.dout(w_dff_B_m9Xf2G8T3_0),.clk(gclk));
	jdff dff_B_TiFcmO2D4_0(.din(w_dff_B_m9Xf2G8T3_0),.dout(w_dff_B_TiFcmO2D4_0),.clk(gclk));
	jdff dff_B_m0jBdFO43_0(.din(w_dff_B_TiFcmO2D4_0),.dout(w_dff_B_m0jBdFO43_0),.clk(gclk));
	jdff dff_B_KL5axc5D2_0(.din(w_dff_B_m0jBdFO43_0),.dout(w_dff_B_KL5axc5D2_0),.clk(gclk));
	jdff dff_B_wdoOD40p2_0(.din(w_dff_B_KL5axc5D2_0),.dout(w_dff_B_wdoOD40p2_0),.clk(gclk));
	jdff dff_B_6H7XOcCL7_0(.din(w_dff_B_wdoOD40p2_0),.dout(w_dff_B_6H7XOcCL7_0),.clk(gclk));
	jdff dff_B_LzblFryV0_0(.din(w_dff_B_6H7XOcCL7_0),.dout(w_dff_B_LzblFryV0_0),.clk(gclk));
	jdff dff_B_mi3BNH5X1_0(.din(w_dff_B_LzblFryV0_0),.dout(w_dff_B_mi3BNH5X1_0),.clk(gclk));
	jdff dff_B_QpuCc7aU9_0(.din(w_dff_B_mi3BNH5X1_0),.dout(w_dff_B_QpuCc7aU9_0),.clk(gclk));
	jdff dff_B_xkI0oTdo9_0(.din(w_dff_B_QpuCc7aU9_0),.dout(w_dff_B_xkI0oTdo9_0),.clk(gclk));
	jdff dff_B_wHs13Xsv8_0(.din(n1292),.dout(w_dff_B_wHs13Xsv8_0),.clk(gclk));
	jdff dff_B_pqqzMUZl8_0(.din(n1301),.dout(w_dff_B_pqqzMUZl8_0),.clk(gclk));
	jdff dff_B_eDGJMUsh1_0(.din(w_dff_B_pqqzMUZl8_0),.dout(w_dff_B_eDGJMUsh1_0),.clk(gclk));
	jdff dff_B_zDEWOE8r4_0(.din(w_dff_B_eDGJMUsh1_0),.dout(w_dff_B_zDEWOE8r4_0),.clk(gclk));
	jdff dff_B_ROW32n2Y7_0(.din(w_dff_B_zDEWOE8r4_0),.dout(w_dff_B_ROW32n2Y7_0),.clk(gclk));
	jdff dff_B_q9BTNHhf8_0(.din(w_dff_B_ROW32n2Y7_0),.dout(w_dff_B_q9BTNHhf8_0),.clk(gclk));
	jdff dff_B_kaE8LV7h8_0(.din(w_dff_B_q9BTNHhf8_0),.dout(w_dff_B_kaE8LV7h8_0),.clk(gclk));
	jdff dff_B_SzuDFWmC0_0(.din(w_dff_B_kaE8LV7h8_0),.dout(w_dff_B_SzuDFWmC0_0),.clk(gclk));
	jdff dff_B_kWLqNuTG3_0(.din(w_dff_B_SzuDFWmC0_0),.dout(w_dff_B_kWLqNuTG3_0),.clk(gclk));
	jdff dff_B_khNQBvbu6_0(.din(w_dff_B_kWLqNuTG3_0),.dout(w_dff_B_khNQBvbu6_0),.clk(gclk));
	jdff dff_B_QnhusBw42_0(.din(w_dff_B_khNQBvbu6_0),.dout(w_dff_B_QnhusBw42_0),.clk(gclk));
	jdff dff_B_6Og4tF8l2_0(.din(w_dff_B_QnhusBw42_0),.dout(w_dff_B_6Og4tF8l2_0),.clk(gclk));
	jdff dff_B_oyFq5PQM6_0(.din(w_dff_B_6Og4tF8l2_0),.dout(w_dff_B_oyFq5PQM6_0),.clk(gclk));
	jdff dff_B_f7rGyw7A4_0(.din(w_dff_B_oyFq5PQM6_0),.dout(w_dff_B_f7rGyw7A4_0),.clk(gclk));
	jdff dff_B_Qqyg0ppa1_0(.din(w_dff_B_f7rGyw7A4_0),.dout(w_dff_B_Qqyg0ppa1_0),.clk(gclk));
	jdff dff_B_OQjliZDL7_0(.din(w_dff_B_Qqyg0ppa1_0),.dout(w_dff_B_OQjliZDL7_0),.clk(gclk));
	jdff dff_B_Gkx80q075_0(.din(w_dff_B_OQjliZDL7_0),.dout(w_dff_B_Gkx80q075_0),.clk(gclk));
	jdff dff_B_2lnt7ZZc6_0(.din(n1300),.dout(w_dff_B_2lnt7ZZc6_0),.clk(gclk));
	jdff dff_A_jkwCsyvQ2_0(.dout(w_n988_2[0]),.din(w_dff_A_jkwCsyvQ2_0),.clk(gclk));
	jdff dff_A_ssvHqDnK6_1(.dout(w_n988_2[1]),.din(w_dff_A_ssvHqDnK6_1),.clk(gclk));
	jdff dff_A_KOcAUxzg9_0(.dout(w_n985_2[0]),.din(w_dff_A_KOcAUxzg9_0),.clk(gclk));
	jdff dff_A_VeVRreo87_1(.dout(w_n985_2[1]),.din(w_dff_A_VeVRreo87_1),.clk(gclk));
	jdff dff_B_psgHtD3X4_0(.din(n1309),.dout(w_dff_B_psgHtD3X4_0),.clk(gclk));
	jdff dff_B_gxhjelfQ0_0(.din(w_dff_B_psgHtD3X4_0),.dout(w_dff_B_gxhjelfQ0_0),.clk(gclk));
	jdff dff_B_4OjYtLMW3_0(.din(w_dff_B_gxhjelfQ0_0),.dout(w_dff_B_4OjYtLMW3_0),.clk(gclk));
	jdff dff_B_uF8pXqRS1_0(.din(w_dff_B_4OjYtLMW3_0),.dout(w_dff_B_uF8pXqRS1_0),.clk(gclk));
	jdff dff_B_lJKaaXEs2_0(.din(w_dff_B_uF8pXqRS1_0),.dout(w_dff_B_lJKaaXEs2_0),.clk(gclk));
	jdff dff_B_0kzx022p2_0(.din(w_dff_B_lJKaaXEs2_0),.dout(w_dff_B_0kzx022p2_0),.clk(gclk));
	jdff dff_B_KBWcRlxM8_0(.din(w_dff_B_0kzx022p2_0),.dout(w_dff_B_KBWcRlxM8_0),.clk(gclk));
	jdff dff_B_5HETUlqq4_0(.din(w_dff_B_KBWcRlxM8_0),.dout(w_dff_B_5HETUlqq4_0),.clk(gclk));
	jdff dff_B_FqzyediK8_0(.din(w_dff_B_5HETUlqq4_0),.dout(w_dff_B_FqzyediK8_0),.clk(gclk));
	jdff dff_B_DtjazNvV6_0(.din(w_dff_B_FqzyediK8_0),.dout(w_dff_B_DtjazNvV6_0),.clk(gclk));
	jdff dff_B_IDd31ii58_0(.din(w_dff_B_DtjazNvV6_0),.dout(w_dff_B_IDd31ii58_0),.clk(gclk));
	jdff dff_B_lhTzgnLZ5_0(.din(w_dff_B_IDd31ii58_0),.dout(w_dff_B_lhTzgnLZ5_0),.clk(gclk));
	jdff dff_B_JafwXmKH7_0(.din(w_dff_B_lhTzgnLZ5_0),.dout(w_dff_B_JafwXmKH7_0),.clk(gclk));
	jdff dff_B_nC5DE3KI8_0(.din(w_dff_B_JafwXmKH7_0),.dout(w_dff_B_nC5DE3KI8_0),.clk(gclk));
	jdff dff_B_KSjAw9yk3_0(.din(w_dff_B_nC5DE3KI8_0),.dout(w_dff_B_KSjAw9yk3_0),.clk(gclk));
	jdff dff_B_oE1JZ1uG7_0(.din(w_dff_B_KSjAw9yk3_0),.dout(w_dff_B_oE1JZ1uG7_0),.clk(gclk));
	jdff dff_B_lClUUBK73_0(.din(w_dff_B_oE1JZ1uG7_0),.dout(w_dff_B_lClUUBK73_0),.clk(gclk));
	jdff dff_B_oir3KOd09_0(.din(n1308),.dout(w_dff_B_oir3KOd09_0),.clk(gclk));
	jdff dff_A_Q5iQULE34_0(.dout(w_G137_5[0]),.din(w_dff_A_Q5iQULE34_0),.clk(gclk));
	jdff dff_B_ACG9gMAr7_0(.din(n1317),.dout(w_dff_B_ACG9gMAr7_0),.clk(gclk));
	jdff dff_B_qqXpbwvH5_0(.din(w_dff_B_ACG9gMAr7_0),.dout(w_dff_B_qqXpbwvH5_0),.clk(gclk));
	jdff dff_B_UBz4wztc2_0(.din(w_dff_B_qqXpbwvH5_0),.dout(w_dff_B_UBz4wztc2_0),.clk(gclk));
	jdff dff_B_zqy8829E1_0(.din(w_dff_B_UBz4wztc2_0),.dout(w_dff_B_zqy8829E1_0),.clk(gclk));
	jdff dff_B_yqPhX9sK0_0(.din(w_dff_B_zqy8829E1_0),.dout(w_dff_B_yqPhX9sK0_0),.clk(gclk));
	jdff dff_B_wNcDOGWv5_0(.din(w_dff_B_yqPhX9sK0_0),.dout(w_dff_B_wNcDOGWv5_0),.clk(gclk));
	jdff dff_B_88WzFsQN7_0(.din(w_dff_B_wNcDOGWv5_0),.dout(w_dff_B_88WzFsQN7_0),.clk(gclk));
	jdff dff_B_6ERaSkNq8_0(.din(w_dff_B_88WzFsQN7_0),.dout(w_dff_B_6ERaSkNq8_0),.clk(gclk));
	jdff dff_B_CegQKCXD2_0(.din(w_dff_B_6ERaSkNq8_0),.dout(w_dff_B_CegQKCXD2_0),.clk(gclk));
	jdff dff_B_1G6AH4SC0_0(.din(w_dff_B_CegQKCXD2_0),.dout(w_dff_B_1G6AH4SC0_0),.clk(gclk));
	jdff dff_B_WXtURZR96_0(.din(w_dff_B_1G6AH4SC0_0),.dout(w_dff_B_WXtURZR96_0),.clk(gclk));
	jdff dff_B_jJ2ZF4MG4_0(.din(w_dff_B_WXtURZR96_0),.dout(w_dff_B_jJ2ZF4MG4_0),.clk(gclk));
	jdff dff_B_QH3IzzPX0_0(.din(w_dff_B_jJ2ZF4MG4_0),.dout(w_dff_B_QH3IzzPX0_0),.clk(gclk));
	jdff dff_B_XoHIIzfZ5_0(.din(w_dff_B_QH3IzzPX0_0),.dout(w_dff_B_XoHIIzfZ5_0),.clk(gclk));
	jdff dff_B_qNDrs8HS5_0(.din(w_dff_B_XoHIIzfZ5_0),.dout(w_dff_B_qNDrs8HS5_0),.clk(gclk));
	jdff dff_B_hu36JLKP8_0(.din(n1316),.dout(w_dff_B_hu36JLKP8_0),.clk(gclk));
	jdff dff_B_Y9eZYFbZ9_2(.din(G173),.dout(w_dff_B_Y9eZYFbZ9_2),.clk(gclk));
	jdff dff_B_7JJA35wq4_2(.din(G203),.dout(w_dff_B_7JJA35wq4_2),.clk(gclk));
	jdff dff_B_hUr9Tjjk0_2(.din(w_dff_B_7JJA35wq4_2),.dout(w_dff_B_hUr9Tjjk0_2),.clk(gclk));
	jdff dff_B_z4ZusqbI3_0(.din(n1182),.dout(w_dff_B_z4ZusqbI3_0),.clk(gclk));
	jdff dff_B_SERaMATc5_0(.din(w_dff_B_z4ZusqbI3_0),.dout(w_dff_B_SERaMATc5_0),.clk(gclk));
	jdff dff_B_qQWxfnOR6_0(.din(w_dff_B_SERaMATc5_0),.dout(w_dff_B_qQWxfnOR6_0),.clk(gclk));
	jdff dff_B_6JgCC1x72_0(.din(w_dff_B_qQWxfnOR6_0),.dout(w_dff_B_6JgCC1x72_0),.clk(gclk));
	jdff dff_B_SXznF4MS1_0(.din(w_dff_B_6JgCC1x72_0),.dout(w_dff_B_SXznF4MS1_0),.clk(gclk));
	jdff dff_B_y1AOhIBq7_0(.din(w_dff_B_SXznF4MS1_0),.dout(w_dff_B_y1AOhIBq7_0),.clk(gclk));
	jdff dff_B_WYbBZJjj3_0(.din(w_dff_B_y1AOhIBq7_0),.dout(w_dff_B_WYbBZJjj3_0),.clk(gclk));
	jdff dff_B_FqOQgcdX0_0(.din(w_dff_B_WYbBZJjj3_0),.dout(w_dff_B_FqOQgcdX0_0),.clk(gclk));
	jdff dff_B_iJl25Ho34_0(.din(w_dff_B_FqOQgcdX0_0),.dout(w_dff_B_iJl25Ho34_0),.clk(gclk));
	jdff dff_B_rjYRKcj64_0(.din(n1181),.dout(w_dff_B_rjYRKcj64_0),.clk(gclk));
	jdff dff_B_L7sOoYjC0_0(.din(w_dff_B_rjYRKcj64_0),.dout(w_dff_B_L7sOoYjC0_0),.clk(gclk));
	jdff dff_B_vhl4Infz5_1(.din(G112),.dout(w_dff_B_vhl4Infz5_1),.clk(gclk));
	jdff dff_B_X0uLgB6d7_1(.din(w_dff_B_vhl4Infz5_1),.dout(w_dff_B_X0uLgB6d7_1),.clk(gclk));
	jdff dff_B_PwIGwvRL3_0(.din(n1218),.dout(w_dff_B_PwIGwvRL3_0),.clk(gclk));
	jdff dff_B_1q36Kfhi6_0(.din(w_dff_B_PwIGwvRL3_0),.dout(w_dff_B_1q36Kfhi6_0),.clk(gclk));
	jdff dff_B_UNlSYR6n1_0(.din(w_dff_B_1q36Kfhi6_0),.dout(w_dff_B_UNlSYR6n1_0),.clk(gclk));
	jdff dff_B_DOuR6GSJ2_0(.din(w_dff_B_UNlSYR6n1_0),.dout(w_dff_B_DOuR6GSJ2_0),.clk(gclk));
	jdff dff_B_LeaNdVMJ4_0(.din(w_dff_B_DOuR6GSJ2_0),.dout(w_dff_B_LeaNdVMJ4_0),.clk(gclk));
	jdff dff_B_GiLV8bMY9_0(.din(w_dff_B_LeaNdVMJ4_0),.dout(w_dff_B_GiLV8bMY9_0),.clk(gclk));
	jdff dff_B_hUklCis55_0(.din(w_dff_B_GiLV8bMY9_0),.dout(w_dff_B_hUklCis55_0),.clk(gclk));
	jdff dff_B_ox7P9IJy7_0(.din(w_dff_B_hUklCis55_0),.dout(w_dff_B_ox7P9IJy7_0),.clk(gclk));
	jdff dff_B_x2KNZ6iI1_0(.din(w_dff_B_ox7P9IJy7_0),.dout(w_dff_B_x2KNZ6iI1_0),.clk(gclk));
	jdff dff_B_IUk8gXyh9_0(.din(w_dff_B_x2KNZ6iI1_0),.dout(w_dff_B_IUk8gXyh9_0),.clk(gclk));
	jdff dff_B_Jior3hBQ9_0(.din(n1217),.dout(w_dff_B_Jior3hBQ9_0),.clk(gclk));
	jdff dff_B_7kBC6HHg6_0(.din(w_dff_B_Jior3hBQ9_0),.dout(w_dff_B_7kBC6HHg6_0),.clk(gclk));
	jdff dff_B_p4kYf6YZ4_1(.din(G113),.dout(w_dff_B_p4kYf6YZ4_1),.clk(gclk));
	jdff dff_B_glA5B8U56_1(.din(w_dff_B_p4kYf6YZ4_1),.dout(w_dff_B_glA5B8U56_1),.clk(gclk));
	jdff dff_B_bXdLyk5W1_0(.din(n539),.dout(w_dff_B_bXdLyk5W1_0),.clk(gclk));
	jdff dff_B_dYPgXtsD0_1(.din(n531),.dout(w_dff_B_dYPgXtsD0_1),.clk(gclk));
	jdff dff_B_IC0ps1fo6_0(.din(n1325),.dout(w_dff_B_IC0ps1fo6_0),.clk(gclk));
	jdff dff_B_jq4fNhWr2_0(.din(w_dff_B_IC0ps1fo6_0),.dout(w_dff_B_jq4fNhWr2_0),.clk(gclk));
	jdff dff_B_cUqcTNe14_0(.din(w_dff_B_jq4fNhWr2_0),.dout(w_dff_B_cUqcTNe14_0),.clk(gclk));
	jdff dff_B_PPDilmP60_0(.din(w_dff_B_cUqcTNe14_0),.dout(w_dff_B_PPDilmP60_0),.clk(gclk));
	jdff dff_B_1StuuxkN7_0(.din(w_dff_B_PPDilmP60_0),.dout(w_dff_B_1StuuxkN7_0),.clk(gclk));
	jdff dff_B_KIgBZSuJ3_0(.din(w_dff_B_1StuuxkN7_0),.dout(w_dff_B_KIgBZSuJ3_0),.clk(gclk));
	jdff dff_B_vbhBoZhC2_0(.din(w_dff_B_KIgBZSuJ3_0),.dout(w_dff_B_vbhBoZhC2_0),.clk(gclk));
	jdff dff_B_U5vzV9CO5_0(.din(w_dff_B_vbhBoZhC2_0),.dout(w_dff_B_U5vzV9CO5_0),.clk(gclk));
	jdff dff_B_7ZOJJbIN4_0(.din(w_dff_B_U5vzV9CO5_0),.dout(w_dff_B_7ZOJJbIN4_0),.clk(gclk));
	jdff dff_B_0gNvbhUZ2_0(.din(w_dff_B_7ZOJJbIN4_0),.dout(w_dff_B_0gNvbhUZ2_0),.clk(gclk));
	jdff dff_B_MQDLUuzm1_0(.din(w_dff_B_0gNvbhUZ2_0),.dout(w_dff_B_MQDLUuzm1_0),.clk(gclk));
	jdff dff_B_iE3s2WX19_0(.din(w_dff_B_MQDLUuzm1_0),.dout(w_dff_B_iE3s2WX19_0),.clk(gclk));
	jdff dff_B_36pvyGsG2_0(.din(w_dff_B_iE3s2WX19_0),.dout(w_dff_B_36pvyGsG2_0),.clk(gclk));
	jdff dff_B_IaAH95SD2_0(.din(w_dff_B_36pvyGsG2_0),.dout(w_dff_B_IaAH95SD2_0),.clk(gclk));
	jdff dff_B_jEhbxsjl3_0(.din(w_dff_B_IaAH95SD2_0),.dout(w_dff_B_jEhbxsjl3_0),.clk(gclk));
	jdff dff_B_gjb4Oi0q0_0(.din(w_dff_B_jEhbxsjl3_0),.dout(w_dff_B_gjb4Oi0q0_0),.clk(gclk));
	jdff dff_B_PVzDrUI07_0(.din(n1324),.dout(w_dff_B_PVzDrUI07_0),.clk(gclk));
	jdff dff_B_EOzGzui27_2(.din(G167),.dout(w_dff_B_EOzGzui27_2),.clk(gclk));
	jdff dff_B_i8SxsqYX0_2(.din(G197),.dout(w_dff_B_i8SxsqYX0_2),.clk(gclk));
	jdff dff_B_SKbHMiPW2_2(.din(w_dff_B_i8SxsqYX0_2),.dout(w_dff_B_SKbHMiPW2_2),.clk(gclk));
	jdff dff_B_PzwauFEn5_0(.din(n1175),.dout(w_dff_B_PzwauFEn5_0),.clk(gclk));
	jdff dff_B_T1WLndiE7_0(.din(w_dff_B_PzwauFEn5_0),.dout(w_dff_B_T1WLndiE7_0),.clk(gclk));
	jdff dff_B_wk2mTHoO6_0(.din(w_dff_B_T1WLndiE7_0),.dout(w_dff_B_wk2mTHoO6_0),.clk(gclk));
	jdff dff_B_uftwXITn5_0(.din(w_dff_B_wk2mTHoO6_0),.dout(w_dff_B_uftwXITn5_0),.clk(gclk));
	jdff dff_B_Pprlg6Pk7_0(.din(w_dff_B_uftwXITn5_0),.dout(w_dff_B_Pprlg6Pk7_0),.clk(gclk));
	jdff dff_B_z1rch9tb1_0(.din(w_dff_B_Pprlg6Pk7_0),.dout(w_dff_B_z1rch9tb1_0),.clk(gclk));
	jdff dff_B_iZHAJWmI6_0(.din(w_dff_B_z1rch9tb1_0),.dout(w_dff_B_iZHAJWmI6_0),.clk(gclk));
	jdff dff_B_tFk35qCd0_0(.din(w_dff_B_iZHAJWmI6_0),.dout(w_dff_B_tFk35qCd0_0),.clk(gclk));
	jdff dff_B_3Qy6W5L95_0(.din(w_dff_B_tFk35qCd0_0),.dout(w_dff_B_3Qy6W5L95_0),.clk(gclk));
	jdff dff_B_hkmYepsr1_0(.din(w_dff_B_3Qy6W5L95_0),.dout(w_dff_B_hkmYepsr1_0),.clk(gclk));
	jdff dff_B_IgMqFLy09_0(.din(n1174),.dout(w_dff_B_IgMqFLy09_0),.clk(gclk));
	jdff dff_B_ua2pDzep4_0(.din(w_dff_B_IgMqFLy09_0),.dout(w_dff_B_ua2pDzep4_0),.clk(gclk));
	jdff dff_B_JQ3weE2T6_1(.din(G116),.dout(w_dff_B_JQ3weE2T6_1),.clk(gclk));
	jdff dff_B_XSMluYwI5_1(.din(w_dff_B_JQ3weE2T6_1),.dout(w_dff_B_XSMluYwI5_1),.clk(gclk));
	jdff dff_A_NuJTEUlq2_1(.dout(w_n971_0[1]),.din(w_dff_A_NuJTEUlq2_1),.clk(gclk));
	jdff dff_B_RLn8NmTO6_1(.din(n967),.dout(w_dff_B_RLn8NmTO6_1),.clk(gclk));
	jdff dff_B_ko7vEbz17_1(.din(w_dff_B_RLn8NmTO6_1),.dout(w_dff_B_ko7vEbz17_1),.clk(gclk));
	jdff dff_B_rTNjjYZQ2_1(.din(w_dff_B_ko7vEbz17_1),.dout(w_dff_B_rTNjjYZQ2_1),.clk(gclk));
	jdff dff_B_I6u7Xvyt7_1(.din(w_dff_B_rTNjjYZQ2_1),.dout(w_dff_B_I6u7Xvyt7_1),.clk(gclk));
	jdff dff_B_9awdeCEy5_1(.din(w_dff_B_I6u7Xvyt7_1),.dout(w_dff_B_9awdeCEy5_1),.clk(gclk));
	jdff dff_B_10FZb3Xe6_1(.din(w_dff_B_9awdeCEy5_1),.dout(w_dff_B_10FZb3Xe6_1),.clk(gclk));
	jdff dff_B_1QTbg1t01_1(.din(w_dff_B_10FZb3Xe6_1),.dout(w_dff_B_1QTbg1t01_1),.clk(gclk));
	jdff dff_B_DTEZEmzc3_1(.din(w_dff_B_1QTbg1t01_1),.dout(w_dff_B_DTEZEmzc3_1),.clk(gclk));
	jdff dff_B_UsBq3o8C3_1(.din(w_dff_B_DTEZEmzc3_1),.dout(w_dff_B_UsBq3o8C3_1),.clk(gclk));
	jdff dff_B_gZZxHR9A9_1(.din(w_dff_B_UsBq3o8C3_1),.dout(w_dff_B_gZZxHR9A9_1),.clk(gclk));
	jdff dff_B_x4ipNBLy2_0(.din(n1211),.dout(w_dff_B_x4ipNBLy2_0),.clk(gclk));
	jdff dff_B_G6R5a1ku6_0(.din(w_dff_B_x4ipNBLy2_0),.dout(w_dff_B_G6R5a1ku6_0),.clk(gclk));
	jdff dff_B_ydD3jYtZ2_0(.din(w_dff_B_G6R5a1ku6_0),.dout(w_dff_B_ydD3jYtZ2_0),.clk(gclk));
	jdff dff_B_pcCgPbGV9_0(.din(w_dff_B_ydD3jYtZ2_0),.dout(w_dff_B_pcCgPbGV9_0),.clk(gclk));
	jdff dff_B_d76h6jha4_0(.din(w_dff_B_pcCgPbGV9_0),.dout(w_dff_B_d76h6jha4_0),.clk(gclk));
	jdff dff_B_gjxnMQvY5_0(.din(w_dff_B_d76h6jha4_0),.dout(w_dff_B_gjxnMQvY5_0),.clk(gclk));
	jdff dff_B_XrZYz4ad6_0(.din(w_dff_B_gjxnMQvY5_0),.dout(w_dff_B_XrZYz4ad6_0),.clk(gclk));
	jdff dff_B_Tbt7paOx5_0(.din(w_dff_B_XrZYz4ad6_0),.dout(w_dff_B_Tbt7paOx5_0),.clk(gclk));
	jdff dff_B_rGvjwjYQ3_0(.din(w_dff_B_Tbt7paOx5_0),.dout(w_dff_B_rGvjwjYQ3_0),.clk(gclk));
	jdff dff_B_XOIjbCTo2_0(.din(w_dff_B_rGvjwjYQ3_0),.dout(w_dff_B_XOIjbCTo2_0),.clk(gclk));
	jdff dff_B_lC30vCYl0_0(.din(w_dff_B_XOIjbCTo2_0),.dout(w_dff_B_lC30vCYl0_0),.clk(gclk));
	jdff dff_B_c3t1imLH3_0(.din(n1210),.dout(w_dff_B_c3t1imLH3_0),.clk(gclk));
	jdff dff_B_CFEHNOeE2_0(.din(w_dff_B_c3t1imLH3_0),.dout(w_dff_B_CFEHNOeE2_0),.clk(gclk));
	jdff dff_B_APznchf67_1(.din(G53),.dout(w_dff_B_APznchf67_1),.clk(gclk));
	jdff dff_B_ZA4O3y686_1(.din(w_dff_B_APznchf67_1),.dout(w_dff_B_ZA4O3y686_1),.clk(gclk));
	jdff dff_B_tG9adEFH1_0(.din(n516),.dout(w_dff_B_tG9adEFH1_0),.clk(gclk));
	jdff dff_B_RjlglxQt3_1(.din(n508),.dout(w_dff_B_RjlglxQt3_1),.clk(gclk));
	jdff dff_B_9hMU6lcc0_1(.din(n949),.dout(w_dff_B_9hMU6lcc0_1),.clk(gclk));
	jdff dff_B_AUupmtsm7_1(.din(w_dff_B_9hMU6lcc0_1),.dout(w_dff_B_AUupmtsm7_1),.clk(gclk));
	jdff dff_B_HtxUaVVx9_1(.din(w_dff_B_AUupmtsm7_1),.dout(w_dff_B_HtxUaVVx9_1),.clk(gclk));
	jdff dff_B_1C0tSIMy4_1(.din(w_dff_B_HtxUaVVx9_1),.dout(w_dff_B_1C0tSIMy4_1),.clk(gclk));
	jdff dff_B_HLW7vWet5_1(.din(w_dff_B_1C0tSIMy4_1),.dout(w_dff_B_HLW7vWet5_1),.clk(gclk));
	jdff dff_B_XQIOUIOp3_1(.din(w_dff_B_HLW7vWet5_1),.dout(w_dff_B_XQIOUIOp3_1),.clk(gclk));
	jdff dff_B_fv1ZyOmz0_1(.din(w_dff_B_XQIOUIOp3_1),.dout(w_dff_B_fv1ZyOmz0_1),.clk(gclk));
	jdff dff_B_RfESNhlC1_1(.din(w_dff_B_fv1ZyOmz0_1),.dout(w_dff_B_RfESNhlC1_1),.clk(gclk));
	jdff dff_B_0hsauJ6R8_1(.din(w_dff_B_RfESNhlC1_1),.dout(w_dff_B_0hsauJ6R8_1),.clk(gclk));
	jdff dff_B_gn54M3Ww9_1(.din(w_dff_B_0hsauJ6R8_1),.dout(w_dff_B_gn54M3Ww9_1),.clk(gclk));
	jdff dff_B_qPVtVFvi2_1(.din(n950),.dout(w_dff_B_qPVtVFvi2_1),.clk(gclk));
	jdff dff_B_IJW9hVqL8_1(.din(w_dff_B_qPVtVFvi2_1),.dout(w_dff_B_IJW9hVqL8_1),.clk(gclk));
	jdff dff_B_CC39pABg7_1(.din(w_dff_B_IJW9hVqL8_1),.dout(w_dff_B_CC39pABg7_1),.clk(gclk));
	jdff dff_B_MkVrTEoD9_1(.din(w_dff_B_CC39pABg7_1),.dout(w_dff_B_MkVrTEoD9_1),.clk(gclk));
	jdff dff_B_0H2DIDvE4_1(.din(w_dff_B_MkVrTEoD9_1),.dout(w_dff_B_0H2DIDvE4_1),.clk(gclk));
	jdff dff_B_lKxuVDm25_1(.din(w_dff_B_0H2DIDvE4_1),.dout(w_dff_B_lKxuVDm25_1),.clk(gclk));
	jdff dff_B_S1QX8Zvs1_1(.din(w_dff_B_lKxuVDm25_1),.dout(w_dff_B_S1QX8Zvs1_1),.clk(gclk));
	jdff dff_B_ofUBp4UG4_1(.din(w_dff_B_S1QX8Zvs1_1),.dout(w_dff_B_ofUBp4UG4_1),.clk(gclk));
	jdff dff_B_rRMNoTYZ7_1(.din(w_dff_B_ofUBp4UG4_1),.dout(w_dff_B_rRMNoTYZ7_1),.clk(gclk));
	jdff dff_A_nWLaiN3j3_1(.dout(w_n748_1[1]),.din(w_dff_A_nWLaiN3j3_1),.clk(gclk));
	jdff dff_A_RJa4Gq8s8_1(.dout(w_dff_A_nWLaiN3j3_1),.din(w_dff_A_RJa4Gq8s8_1),.clk(gclk));
	jdff dff_A_MBuGZqLz6_1(.dout(w_dff_A_RJa4Gq8s8_1),.din(w_dff_A_MBuGZqLz6_1),.clk(gclk));
	jdff dff_A_dhUJ9rvE6_1(.dout(w_dff_A_MBuGZqLz6_1),.din(w_dff_A_dhUJ9rvE6_1),.clk(gclk));
	jdff dff_A_FilrnN435_1(.dout(w_dff_A_dhUJ9rvE6_1),.din(w_dff_A_FilrnN435_1),.clk(gclk));
	jdff dff_A_nahFt7xa8_1(.dout(w_dff_A_FilrnN435_1),.din(w_dff_A_nahFt7xa8_1),.clk(gclk));
	jdff dff_A_CqfnTfWi7_1(.dout(w_dff_A_nahFt7xa8_1),.din(w_dff_A_CqfnTfWi7_1),.clk(gclk));
	jdff dff_A_anLfhxRS1_1(.dout(w_dff_A_CqfnTfWi7_1),.din(w_dff_A_anLfhxRS1_1),.clk(gclk));
	jdff dff_A_Ogz8PFMW1_1(.dout(w_dff_A_anLfhxRS1_1),.din(w_dff_A_Ogz8PFMW1_1),.clk(gclk));
	jdff dff_A_HZjtsSJL1_1(.dout(w_dff_A_Ogz8PFMW1_1),.din(w_dff_A_HZjtsSJL1_1),.clk(gclk));
	jdff dff_A_UhTU1Eae9_1(.dout(w_dff_A_HZjtsSJL1_1),.din(w_dff_A_UhTU1Eae9_1),.clk(gclk));
	jdff dff_A_PJayM3t63_1(.dout(w_dff_A_UhTU1Eae9_1),.din(w_dff_A_PJayM3t63_1),.clk(gclk));
	jdff dff_A_LgHOED8V7_1(.dout(w_dff_A_PJayM3t63_1),.din(w_dff_A_LgHOED8V7_1),.clk(gclk));
	jdff dff_A_KXRjMjqW9_2(.dout(w_n748_1[2]),.din(w_dff_A_KXRjMjqW9_2),.clk(gclk));
	jdff dff_A_dwuX4k8i2_2(.dout(w_dff_A_KXRjMjqW9_2),.din(w_dff_A_dwuX4k8i2_2),.clk(gclk));
	jdff dff_A_LTgyNi8J7_2(.dout(w_dff_A_dwuX4k8i2_2),.din(w_dff_A_LTgyNi8J7_2),.clk(gclk));
	jdff dff_A_JkOpa6Sh7_2(.dout(w_dff_A_LTgyNi8J7_2),.din(w_dff_A_JkOpa6Sh7_2),.clk(gclk));
	jdff dff_A_eIOE29rS2_2(.dout(w_dff_A_JkOpa6Sh7_2),.din(w_dff_A_eIOE29rS2_2),.clk(gclk));
	jdff dff_A_fDzeVmLY4_2(.dout(w_dff_A_eIOE29rS2_2),.din(w_dff_A_fDzeVmLY4_2),.clk(gclk));
	jdff dff_A_KudOem1w6_2(.dout(w_dff_A_fDzeVmLY4_2),.din(w_dff_A_KudOem1w6_2),.clk(gclk));
	jdff dff_A_TdZh7eaG9_2(.dout(w_dff_A_KudOem1w6_2),.din(w_dff_A_TdZh7eaG9_2),.clk(gclk));
	jdff dff_A_GBoCOpiM3_2(.dout(w_dff_A_TdZh7eaG9_2),.din(w_dff_A_GBoCOpiM3_2),.clk(gclk));
	jdff dff_A_MYgwYiWG7_2(.dout(w_dff_A_GBoCOpiM3_2),.din(w_dff_A_MYgwYiWG7_2),.clk(gclk));
	jdff dff_A_Fz0Ytbk11_2(.dout(w_dff_A_MYgwYiWG7_2),.din(w_dff_A_Fz0Ytbk11_2),.clk(gclk));
	jdff dff_A_A5Gq2DXr3_2(.dout(w_dff_A_Fz0Ytbk11_2),.din(w_dff_A_A5Gq2DXr3_2),.clk(gclk));
	jdff dff_B_nkCdGZ7y3_0(.din(n1333),.dout(w_dff_B_nkCdGZ7y3_0),.clk(gclk));
	jdff dff_B_yCMt4mVz6_0(.din(w_dff_B_nkCdGZ7y3_0),.dout(w_dff_B_yCMt4mVz6_0),.clk(gclk));
	jdff dff_B_QxcVWerE2_0(.din(w_dff_B_yCMt4mVz6_0),.dout(w_dff_B_QxcVWerE2_0),.clk(gclk));
	jdff dff_B_YDjt6HPO6_0(.din(w_dff_B_QxcVWerE2_0),.dout(w_dff_B_YDjt6HPO6_0),.clk(gclk));
	jdff dff_B_s29JAerm7_0(.din(w_dff_B_YDjt6HPO6_0),.dout(w_dff_B_s29JAerm7_0),.clk(gclk));
	jdff dff_B_kAboX37W9_0(.din(w_dff_B_s29JAerm7_0),.dout(w_dff_B_kAboX37W9_0),.clk(gclk));
	jdff dff_B_C8cMFetO5_0(.din(w_dff_B_kAboX37W9_0),.dout(w_dff_B_C8cMFetO5_0),.clk(gclk));
	jdff dff_B_Lltmh7hF3_0(.din(w_dff_B_C8cMFetO5_0),.dout(w_dff_B_Lltmh7hF3_0),.clk(gclk));
	jdff dff_B_JoVEzuEX1_0(.din(w_dff_B_Lltmh7hF3_0),.dout(w_dff_B_JoVEzuEX1_0),.clk(gclk));
	jdff dff_B_TGEMRHmX9_0(.din(w_dff_B_JoVEzuEX1_0),.dout(w_dff_B_TGEMRHmX9_0),.clk(gclk));
	jdff dff_B_ru1xUOcn8_0(.din(w_dff_B_TGEMRHmX9_0),.dout(w_dff_B_ru1xUOcn8_0),.clk(gclk));
	jdff dff_B_BNYDaigi9_0(.din(w_dff_B_ru1xUOcn8_0),.dout(w_dff_B_BNYDaigi9_0),.clk(gclk));
	jdff dff_B_7jJuMPSE4_0(.din(w_dff_B_BNYDaigi9_0),.dout(w_dff_B_7jJuMPSE4_0),.clk(gclk));
	jdff dff_B_pZZobhUw4_0(.din(w_dff_B_7jJuMPSE4_0),.dout(w_dff_B_pZZobhUw4_0),.clk(gclk));
	jdff dff_B_tpSFld6Y9_0(.din(w_dff_B_pZZobhUw4_0),.dout(w_dff_B_tpSFld6Y9_0),.clk(gclk));
	jdff dff_B_aAqwkRiN8_0(.din(w_dff_B_tpSFld6Y9_0),.dout(w_dff_B_aAqwkRiN8_0),.clk(gclk));
	jdff dff_B_E09Mezaa2_0(.din(n1332),.dout(w_dff_B_E09Mezaa2_0),.clk(gclk));
	jdff dff_B_CxepozI67_2(.din(G164),.dout(w_dff_B_CxepozI67_2),.clk(gclk));
	jdff dff_B_klaNNE4T8_2(.din(G194),.dout(w_dff_B_klaNNE4T8_2),.clk(gclk));
	jdff dff_B_lvXXY4k86_2(.din(w_dff_B_klaNNE4T8_2),.dout(w_dff_B_lvXXY4k86_2),.clk(gclk));
	jdff dff_B_Zj9p7RCB0_0(.din(n1169),.dout(w_dff_B_Zj9p7RCB0_0),.clk(gclk));
	jdff dff_B_Lnfhs4QJ8_0(.din(w_dff_B_Zj9p7RCB0_0),.dout(w_dff_B_Lnfhs4QJ8_0),.clk(gclk));
	jdff dff_B_9wzovW1K1_0(.din(w_dff_B_Lnfhs4QJ8_0),.dout(w_dff_B_9wzovW1K1_0),.clk(gclk));
	jdff dff_B_AYQXw4ah0_0(.din(w_dff_B_9wzovW1K1_0),.dout(w_dff_B_AYQXw4ah0_0),.clk(gclk));
	jdff dff_B_EKrRSiUS5_0(.din(w_dff_B_AYQXw4ah0_0),.dout(w_dff_B_EKrRSiUS5_0),.clk(gclk));
	jdff dff_B_fCIcrYzg0_0(.din(w_dff_B_EKrRSiUS5_0),.dout(w_dff_B_fCIcrYzg0_0),.clk(gclk));
	jdff dff_B_vXM1eHmw1_0(.din(w_dff_B_fCIcrYzg0_0),.dout(w_dff_B_vXM1eHmw1_0),.clk(gclk));
	jdff dff_B_UaeLKGLt7_0(.din(w_dff_B_vXM1eHmw1_0),.dout(w_dff_B_UaeLKGLt7_0),.clk(gclk));
	jdff dff_B_lpELGz3b9_0(.din(w_dff_B_UaeLKGLt7_0),.dout(w_dff_B_lpELGz3b9_0),.clk(gclk));
	jdff dff_B_EjCPy7S41_0(.din(w_dff_B_lpELGz3b9_0),.dout(w_dff_B_EjCPy7S41_0),.clk(gclk));
	jdff dff_B_x44aRKhf9_0(.din(w_dff_B_EjCPy7S41_0),.dout(w_dff_B_x44aRKhf9_0),.clk(gclk));
	jdff dff_B_V7eyhQDU8_0(.din(n1167),.dout(w_dff_B_V7eyhQDU8_0),.clk(gclk));
	jdff dff_B_ODsq8MGz9_1(.din(G121),.dout(w_dff_B_ODsq8MGz9_1),.clk(gclk));
	jdff dff_B_5BhY4KmB4_1(.din(w_dff_B_ODsq8MGz9_1),.dout(w_dff_B_5BhY4KmB4_1),.clk(gclk));
	jdff dff_A_fVD0VTxf3_0(.dout(w_n748_2[0]),.din(w_dff_A_fVD0VTxf3_0),.clk(gclk));
	jdff dff_A_j5OiPsNP5_0(.dout(w_dff_A_fVD0VTxf3_0),.din(w_dff_A_j5OiPsNP5_0),.clk(gclk));
	jdff dff_A_gWYGPnUF3_0(.dout(w_dff_A_j5OiPsNP5_0),.din(w_dff_A_gWYGPnUF3_0),.clk(gclk));
	jdff dff_A_tN7pN9zS4_0(.dout(w_dff_A_gWYGPnUF3_0),.din(w_dff_A_tN7pN9zS4_0),.clk(gclk));
	jdff dff_A_J8FNQi6d4_2(.dout(w_n748_2[2]),.din(w_dff_A_J8FNQi6d4_2),.clk(gclk));
	jdff dff_A_LBlA3ipn0_2(.dout(w_dff_A_J8FNQi6d4_2),.din(w_dff_A_LBlA3ipn0_2),.clk(gclk));
	jdff dff_A_5jVlxlEd8_1(.dout(w_n748_0[1]),.din(w_dff_A_5jVlxlEd8_1),.clk(gclk));
	jdff dff_A_IHZUTaxN7_1(.dout(w_dff_A_5jVlxlEd8_1),.din(w_dff_A_IHZUTaxN7_1),.clk(gclk));
	jdff dff_A_L8w0sTR85_1(.dout(w_dff_A_IHZUTaxN7_1),.din(w_dff_A_L8w0sTR85_1),.clk(gclk));
	jdff dff_A_P39oH47z7_1(.dout(w_dff_A_L8w0sTR85_1),.din(w_dff_A_P39oH47z7_1),.clk(gclk));
	jdff dff_A_8t14FyZA1_1(.dout(w_dff_A_P39oH47z7_1),.din(w_dff_A_8t14FyZA1_1),.clk(gclk));
	jdff dff_A_pY7FLW693_1(.dout(w_dff_A_8t14FyZA1_1),.din(w_dff_A_pY7FLW693_1),.clk(gclk));
	jdff dff_A_LPC2Hmgb2_1(.dout(w_dff_A_pY7FLW693_1),.din(w_dff_A_LPC2Hmgb2_1),.clk(gclk));
	jdff dff_A_zUHE6OJp7_1(.dout(w_dff_A_LPC2Hmgb2_1),.din(w_dff_A_zUHE6OJp7_1),.clk(gclk));
	jdff dff_A_8kFX6j9B3_2(.dout(w_n748_0[2]),.din(w_dff_A_8kFX6j9B3_2),.clk(gclk));
	jdff dff_A_uLgdoARU2_2(.dout(w_dff_A_8kFX6j9B3_2),.din(w_dff_A_uLgdoARU2_2),.clk(gclk));
	jdff dff_A_FT2KWkZO9_2(.dout(w_dff_A_uLgdoARU2_2),.din(w_dff_A_FT2KWkZO9_2),.clk(gclk));
	jdff dff_A_zkyVJEDD9_2(.dout(w_dff_A_FT2KWkZO9_2),.din(w_dff_A_zkyVJEDD9_2),.clk(gclk));
	jdff dff_B_b3QgmtF84_3(.din(n748),.dout(w_dff_B_b3QgmtF84_3),.clk(gclk));
	jdff dff_A_NxO5wa0G9_0(.dout(w_n747_3[0]),.din(w_dff_A_NxO5wa0G9_0),.clk(gclk));
	jdff dff_A_v2tOVFxg8_0(.dout(w_dff_A_NxO5wa0G9_0),.din(w_dff_A_v2tOVFxg8_0),.clk(gclk));
	jdff dff_A_S9KUT1RQ5_0(.dout(w_dff_A_v2tOVFxg8_0),.din(w_dff_A_S9KUT1RQ5_0),.clk(gclk));
	jdff dff_A_jS25Wu2N0_0(.dout(w_dff_A_S9KUT1RQ5_0),.din(w_dff_A_jS25Wu2N0_0),.clk(gclk));
	jdff dff_A_0qt0LoFx1_0(.dout(w_dff_A_jS25Wu2N0_0),.din(w_dff_A_0qt0LoFx1_0),.clk(gclk));
	jdff dff_A_RlqxV35g6_0(.dout(w_dff_A_0qt0LoFx1_0),.din(w_dff_A_RlqxV35g6_0),.clk(gclk));
	jdff dff_A_UG4xlEf71_0(.dout(w_dff_A_RlqxV35g6_0),.din(w_dff_A_UG4xlEf71_0),.clk(gclk));
	jdff dff_A_ZUTBvrie0_0(.dout(w_dff_A_UG4xlEf71_0),.din(w_dff_A_ZUTBvrie0_0),.clk(gclk));
	jdff dff_A_rOaXI9Y85_1(.dout(w_n747_3[1]),.din(w_dff_A_rOaXI9Y85_1),.clk(gclk));
	jdff dff_A_usYtItjc0_1(.dout(w_dff_A_rOaXI9Y85_1),.din(w_dff_A_usYtItjc0_1),.clk(gclk));
	jdff dff_A_osacSdo95_1(.dout(w_dff_A_usYtItjc0_1),.din(w_dff_A_osacSdo95_1),.clk(gclk));
	jdff dff_A_QVXdpFrt1_0(.dout(w_n1002_2[0]),.din(w_dff_A_QVXdpFrt1_0),.clk(gclk));
	jdff dff_A_PddqTTdc0_1(.dout(w_n1002_2[1]),.din(w_dff_A_PddqTTdc0_1),.clk(gclk));
	jdff dff_B_d3sjWix71_0(.din(n1204),.dout(w_dff_B_d3sjWix71_0),.clk(gclk));
	jdff dff_B_A9hyVSUf9_0(.din(w_dff_B_d3sjWix71_0),.dout(w_dff_B_A9hyVSUf9_0),.clk(gclk));
	jdff dff_B_NUK6N2kP4_0(.din(w_dff_B_A9hyVSUf9_0),.dout(w_dff_B_NUK6N2kP4_0),.clk(gclk));
	jdff dff_B_3ZpBAuHt9_0(.din(w_dff_B_NUK6N2kP4_0),.dout(w_dff_B_3ZpBAuHt9_0),.clk(gclk));
	jdff dff_B_dDNTTR8P3_0(.din(w_dff_B_3ZpBAuHt9_0),.dout(w_dff_B_dDNTTR8P3_0),.clk(gclk));
	jdff dff_B_fxXG1myj6_0(.din(w_dff_B_dDNTTR8P3_0),.dout(w_dff_B_fxXG1myj6_0),.clk(gclk));
	jdff dff_B_YXLkdU1c7_0(.din(w_dff_B_fxXG1myj6_0),.dout(w_dff_B_YXLkdU1c7_0),.clk(gclk));
	jdff dff_B_fFUvJFBQ3_0(.din(w_dff_B_YXLkdU1c7_0),.dout(w_dff_B_fFUvJFBQ3_0),.clk(gclk));
	jdff dff_B_5DHQsWWb3_0(.din(w_dff_B_fFUvJFBQ3_0),.dout(w_dff_B_5DHQsWWb3_0),.clk(gclk));
	jdff dff_B_g2gwllFI2_0(.din(w_dff_B_5DHQsWWb3_0),.dout(w_dff_B_g2gwllFI2_0),.clk(gclk));
	jdff dff_B_Nq2ZTkki8_0(.din(w_dff_B_g2gwllFI2_0),.dout(w_dff_B_Nq2ZTkki8_0),.clk(gclk));
	jdff dff_B_DpIp5SnS1_0(.din(n1202),.dout(w_dff_B_DpIp5SnS1_0),.clk(gclk));
	jdff dff_B_7NIGw5Oa9_0(.din(w_dff_B_DpIp5SnS1_0),.dout(w_dff_B_7NIGw5Oa9_0),.clk(gclk));
	jdff dff_B_CT8997VH1_1(.din(G114),.dout(w_dff_B_CT8997VH1_1),.clk(gclk));
	jdff dff_B_LjNP1xe75_1(.din(w_dff_B_CT8997VH1_1),.dout(w_dff_B_LjNP1xe75_1),.clk(gclk));
	jdff dff_B_Cb6NJFBH6_3(.din(n765),.dout(w_dff_B_Cb6NJFBH6_3),.clk(gclk));
	jdff dff_B_f8EmpGFW4_3(.din(w_dff_B_Cb6NJFBH6_3),.dout(w_dff_B_f8EmpGFW4_3),.clk(gclk));
	jdff dff_A_JkGZyrSp0_1(.dout(w_n751_2[1]),.din(w_dff_A_JkGZyrSp0_1),.clk(gclk));
	jdff dff_B_zfgiQdEd9_0(.din(n550),.dout(w_dff_B_zfgiQdEd9_0),.clk(gclk));
	jdff dff_B_4Q09WIFX4_3(.din(G3548),.dout(w_dff_B_4Q09WIFX4_3),.clk(gclk));
	jdff dff_B_XX2WTl2R5_1(.din(n542),.dout(w_dff_B_XX2WTl2R5_1),.clk(gclk));
	jdff dff_A_EFjtmaS02_0(.dout(w_n999_2[0]),.din(w_dff_A_EFjtmaS02_0),.clk(gclk));
	jdff dff_A_b2cAoQXM2_1(.dout(w_n999_2[1]),.din(w_dff_A_b2cAoQXM2_1),.clk(gclk));
	jdff dff_A_FvGkOaCi3_0(.dout(w_G137_4[0]),.din(w_dff_A_FvGkOaCi3_0),.clk(gclk));
	jdff dff_A_SL2CkCQG0_1(.dout(w_G137_4[1]),.din(w_dff_A_SL2CkCQG0_1),.clk(gclk));
	jdff dff_A_Rb2uXiFi0_0(.dout(w_G137_1[0]),.din(w_dff_A_Rb2uXiFi0_0),.clk(gclk));
	jdff dff_A_W6ugICTc9_0(.dout(w_dff_A_Rb2uXiFi0_0),.din(w_dff_A_W6ugICTc9_0),.clk(gclk));
	jdff dff_A_ntctoOUO0_0(.dout(w_dff_A_W6ugICTc9_0),.din(w_dff_A_ntctoOUO0_0),.clk(gclk));
	jdff dff_A_bnJMv21n0_0(.dout(w_dff_A_ntctoOUO0_0),.din(w_dff_A_bnJMv21n0_0),.clk(gclk));
	jdff dff_A_vkKShGM35_0(.dout(w_dff_A_bnJMv21n0_0),.din(w_dff_A_vkKShGM35_0),.clk(gclk));
	jdff dff_A_0PYOUKfD7_1(.dout(w_G137_1[1]),.din(w_dff_A_0PYOUKfD7_1),.clk(gclk));
	jdff dff_A_63Qn5KIc5_1(.dout(w_dff_A_0PYOUKfD7_1),.din(w_dff_A_63Qn5KIc5_1),.clk(gclk));
	jdff dff_A_5JtNalT21_1(.dout(w_dff_A_63Qn5KIc5_1),.din(w_dff_A_5JtNalT21_1),.clk(gclk));
	jdff dff_A_4FmLSURR9_1(.dout(w_dff_A_5JtNalT21_1),.din(w_dff_A_4FmLSURR9_1),.clk(gclk));
	jdff dff_A_uTGBBX7c2_1(.dout(w_dff_A_4FmLSURR9_1),.din(w_dff_A_uTGBBX7c2_1),.clk(gclk));
	jdff dff_A_pomlwqel7_1(.dout(w_dff_A_uTGBBX7c2_1),.din(w_dff_A_pomlwqel7_1),.clk(gclk));
	jdff dff_B_DTKs4Je02_0(.din(n1341),.dout(w_dff_B_DTKs4Je02_0),.clk(gclk));
	jdff dff_B_wDPyu4xs2_0(.din(w_dff_B_DTKs4Je02_0),.dout(w_dff_B_wDPyu4xs2_0),.clk(gclk));
	jdff dff_B_I4ifPtmg6_0(.din(w_dff_B_wDPyu4xs2_0),.dout(w_dff_B_I4ifPtmg6_0),.clk(gclk));
	jdff dff_B_ZiaTwSdv9_0(.din(w_dff_B_I4ifPtmg6_0),.dout(w_dff_B_ZiaTwSdv9_0),.clk(gclk));
	jdff dff_B_rlthOJX65_0(.din(w_dff_B_ZiaTwSdv9_0),.dout(w_dff_B_rlthOJX65_0),.clk(gclk));
	jdff dff_B_hqaKMx2x5_0(.din(w_dff_B_rlthOJX65_0),.dout(w_dff_B_hqaKMx2x5_0),.clk(gclk));
	jdff dff_B_HWXO9WmH8_0(.din(w_dff_B_hqaKMx2x5_0),.dout(w_dff_B_HWXO9WmH8_0),.clk(gclk));
	jdff dff_B_huJjbbAv2_0(.din(w_dff_B_HWXO9WmH8_0),.dout(w_dff_B_huJjbbAv2_0),.clk(gclk));
	jdff dff_B_ewH1lAGq8_0(.din(w_dff_B_huJjbbAv2_0),.dout(w_dff_B_ewH1lAGq8_0),.clk(gclk));
	jdff dff_B_J6Yoh2Hq6_0(.din(w_dff_B_ewH1lAGq8_0),.dout(w_dff_B_J6Yoh2Hq6_0),.clk(gclk));
	jdff dff_B_ZWU5zdNs8_0(.din(w_dff_B_J6Yoh2Hq6_0),.dout(w_dff_B_ZWU5zdNs8_0),.clk(gclk));
	jdff dff_B_SvYarsVD2_0(.din(w_dff_B_ZWU5zdNs8_0),.dout(w_dff_B_SvYarsVD2_0),.clk(gclk));
	jdff dff_B_VYJB5g7M7_0(.din(w_dff_B_SvYarsVD2_0),.dout(w_dff_B_VYJB5g7M7_0),.clk(gclk));
	jdff dff_B_RntGXBae2_0(.din(w_dff_B_VYJB5g7M7_0),.dout(w_dff_B_RntGXBae2_0),.clk(gclk));
	jdff dff_B_azOiCFjl0_0(.din(w_dff_B_RntGXBae2_0),.dout(w_dff_B_azOiCFjl0_0),.clk(gclk));
	jdff dff_B_ks6belN15_0(.din(w_dff_B_azOiCFjl0_0),.dout(w_dff_B_ks6belN15_0),.clk(gclk));
	jdff dff_B_nfMwAaDh9_0(.din(w_dff_B_ks6belN15_0),.dout(w_dff_B_nfMwAaDh9_0),.clk(gclk));
	jdff dff_B_CDnC17cx4_0(.din(n1340),.dout(w_dff_B_CDnC17cx4_0),.clk(gclk));
	jdff dff_B_xSQVsPoZ2_2(.din(G161),.dout(w_dff_B_xSQVsPoZ2_2),.clk(gclk));
	jdff dff_B_PEnNw0c31_2(.din(G191),.dout(w_dff_B_PEnNw0c31_2),.clk(gclk));
	jdff dff_B_58usAc7i4_2(.din(w_dff_B_PEnNw0c31_2),.dout(w_dff_B_58usAc7i4_2),.clk(gclk));
	jdff dff_B_eJUZaB8a5_0(.din(n1162),.dout(w_dff_B_eJUZaB8a5_0),.clk(gclk));
	jdff dff_B_PzBOjRNh7_0(.din(w_dff_B_eJUZaB8a5_0),.dout(w_dff_B_PzBOjRNh7_0),.clk(gclk));
	jdff dff_B_d63iWvuT2_0(.din(w_dff_B_PzBOjRNh7_0),.dout(w_dff_B_d63iWvuT2_0),.clk(gclk));
	jdff dff_B_DJpVwbnP6_0(.din(w_dff_B_d63iWvuT2_0),.dout(w_dff_B_DJpVwbnP6_0),.clk(gclk));
	jdff dff_B_I2jWeDpn4_0(.din(w_dff_B_DJpVwbnP6_0),.dout(w_dff_B_I2jWeDpn4_0),.clk(gclk));
	jdff dff_B_Oj6apF427_0(.din(w_dff_B_I2jWeDpn4_0),.dout(w_dff_B_Oj6apF427_0),.clk(gclk));
	jdff dff_B_EvuBXMid2_0(.din(w_dff_B_Oj6apF427_0),.dout(w_dff_B_EvuBXMid2_0),.clk(gclk));
	jdff dff_B_ckMwtmqC4_0(.din(w_dff_B_EvuBXMid2_0),.dout(w_dff_B_ckMwtmqC4_0),.clk(gclk));
	jdff dff_B_CBRfLtzW5_0(.din(w_dff_B_ckMwtmqC4_0),.dout(w_dff_B_CBRfLtzW5_0),.clk(gclk));
	jdff dff_B_loyjdCvL4_0(.din(w_dff_B_CBRfLtzW5_0),.dout(w_dff_B_loyjdCvL4_0),.clk(gclk));
	jdff dff_B_edH823860_0(.din(w_dff_B_loyjdCvL4_0),.dout(w_dff_B_edH823860_0),.clk(gclk));
	jdff dff_B_yNJqNkWF5_0(.din(w_dff_B_edH823860_0),.dout(w_dff_B_yNJqNkWF5_0),.clk(gclk));
	jdff dff_B_J5ifSxXj6_0(.din(w_dff_B_yNJqNkWF5_0),.dout(w_dff_B_J5ifSxXj6_0),.clk(gclk));
	jdff dff_B_4yZCFnr61_1(.din(n1160),.dout(w_dff_B_4yZCFnr61_1),.clk(gclk));
	jdff dff_B_kWE29rax3_1(.din(w_dff_B_4yZCFnr61_1),.dout(w_dff_B_kWE29rax3_1),.clk(gclk));
	jdff dff_A_Oy42UHnV4_1(.dout(w_n751_1[1]),.din(w_dff_A_Oy42UHnV4_1),.clk(gclk));
	jdff dff_A_hzg3IKyz0_0(.dout(w_G123_0[0]),.din(w_dff_A_hzg3IKyz0_0),.clk(gclk));
	jdff dff_B_HPz1yzyw0_2(.din(G123),.dout(w_dff_B_HPz1yzyw0_2),.clk(gclk));
	jdff dff_B_9gUly01L6_0(.din(n788),.dout(w_dff_B_9gUly01L6_0),.clk(gclk));
	jdff dff_B_XBueP9mY3_0(.din(n780),.dout(w_dff_B_XBueP9mY3_0),.clk(gclk));
	jdff dff_B_2aJGrS2I8_0(.din(w_dff_B_XBueP9mY3_0),.dout(w_dff_B_2aJGrS2I8_0),.clk(gclk));
	jdff dff_B_5Ubx6wng4_0(.din(w_dff_B_2aJGrS2I8_0),.dout(w_dff_B_5Ubx6wng4_0),.clk(gclk));
	jdff dff_A_YoUpGZEF4_0(.dout(w_G54_0[0]),.din(w_dff_A_YoUpGZEF4_0),.clk(gclk));
	jdff dff_A_rPl93rKj3_0(.dout(w_dff_A_YoUpGZEF4_0),.din(w_dff_A_rPl93rKj3_0),.clk(gclk));
	jdff dff_A_mrLIkdhc0_0(.dout(w_dff_A_rPl93rKj3_0),.din(w_dff_A_mrLIkdhc0_0),.clk(gclk));
	jdff dff_A_HX7RCHHO4_0(.dout(w_dff_A_mrLIkdhc0_0),.din(w_dff_A_HX7RCHHO4_0),.clk(gclk));
	jdff dff_A_32h8KHfo0_0(.dout(w_dff_A_HX7RCHHO4_0),.din(w_dff_A_32h8KHfo0_0),.clk(gclk));
	jdff dff_A_VTwCLqoy3_0(.dout(w_dff_A_32h8KHfo0_0),.din(w_dff_A_VTwCLqoy3_0),.clk(gclk));
	jdff dff_A_TrW88K8S7_0(.dout(w_dff_A_VTwCLqoy3_0),.din(w_dff_A_TrW88K8S7_0),.clk(gclk));
	jdff dff_A_TBOZGujq2_0(.dout(w_dff_A_TrW88K8S7_0),.din(w_dff_A_TBOZGujq2_0),.clk(gclk));
	jdff dff_A_MmPMhp1X7_0(.dout(w_n741_0[0]),.din(w_dff_A_MmPMhp1X7_0),.clk(gclk));
	jdff dff_A_M3lqmndX0_0(.dout(w_dff_A_MmPMhp1X7_0),.din(w_dff_A_M3lqmndX0_0),.clk(gclk));
	jdff dff_A_CHgitgri5_0(.dout(w_dff_A_M3lqmndX0_0),.din(w_dff_A_CHgitgri5_0),.clk(gclk));
	jdff dff_A_uYvlz1NO4_0(.dout(w_dff_A_CHgitgri5_0),.din(w_dff_A_uYvlz1NO4_0),.clk(gclk));
	jdff dff_A_HeLRgrdp3_0(.dout(w_dff_A_uYvlz1NO4_0),.din(w_dff_A_HeLRgrdp3_0),.clk(gclk));
	jdff dff_A_9miJU0V01_0(.dout(w_dff_A_HeLRgrdp3_0),.din(w_dff_A_9miJU0V01_0),.clk(gclk));
	jdff dff_A_1huJGL037_0(.dout(w_dff_A_9miJU0V01_0),.din(w_dff_A_1huJGL037_0),.clk(gclk));
	jdff dff_A_HwQ6OJs31_0(.dout(w_n747_2[0]),.din(w_dff_A_HwQ6OJs31_0),.clk(gclk));
	jdff dff_A_TXqFKuK68_0(.dout(w_dff_A_HwQ6OJs31_0),.din(w_dff_A_TXqFKuK68_0),.clk(gclk));
	jdff dff_A_q1y4R3CG4_0(.dout(w_dff_A_TXqFKuK68_0),.din(w_dff_A_q1y4R3CG4_0),.clk(gclk));
	jdff dff_A_X0si2R2Z8_0(.dout(w_dff_A_q1y4R3CG4_0),.din(w_dff_A_X0si2R2Z8_0),.clk(gclk));
	jdff dff_A_69179VsI2_0(.dout(w_dff_A_X0si2R2Z8_0),.din(w_dff_A_69179VsI2_0),.clk(gclk));
	jdff dff_A_wyGNDgss6_1(.dout(w_n747_2[1]),.din(w_dff_A_wyGNDgss6_1),.clk(gclk));
	jdff dff_A_4vjFKfps3_1(.dout(w_dff_A_wyGNDgss6_1),.din(w_dff_A_4vjFKfps3_1),.clk(gclk));
	jdff dff_A_z46HEOva8_1(.dout(w_dff_A_4vjFKfps3_1),.din(w_dff_A_z46HEOva8_1),.clk(gclk));
	jdff dff_A_3FY1pyvB8_1(.dout(w_dff_A_z46HEOva8_1),.din(w_dff_A_3FY1pyvB8_1),.clk(gclk));
	jdff dff_A_v7267uGc8_1(.dout(w_dff_A_3FY1pyvB8_1),.din(w_dff_A_v7267uGc8_1),.clk(gclk));
	jdff dff_A_DiLJ8cCA6_1(.dout(w_dff_A_v7267uGc8_1),.din(w_dff_A_DiLJ8cCA6_1),.clk(gclk));
	jdff dff_A_2Llhfgir8_1(.dout(w_dff_A_DiLJ8cCA6_1),.din(w_dff_A_2Llhfgir8_1),.clk(gclk));
	jdff dff_A_vLqVZ47g5_1(.dout(w_dff_A_2Llhfgir8_1),.din(w_dff_A_vLqVZ47g5_1),.clk(gclk));
	jdff dff_A_Kd60217a3_1(.dout(w_dff_A_vLqVZ47g5_1),.din(w_dff_A_Kd60217a3_1),.clk(gclk));
	jdff dff_B_ftj9PPAC3_0(.din(n1196),.dout(w_dff_B_ftj9PPAC3_0),.clk(gclk));
	jdff dff_B_dGKwyCEr2_0(.din(w_dff_B_ftj9PPAC3_0),.dout(w_dff_B_dGKwyCEr2_0),.clk(gclk));
	jdff dff_B_WepTQcQ25_0(.din(w_dff_B_dGKwyCEr2_0),.dout(w_dff_B_WepTQcQ25_0),.clk(gclk));
	jdff dff_B_varN7BWI9_0(.din(w_dff_B_WepTQcQ25_0),.dout(w_dff_B_varN7BWI9_0),.clk(gclk));
	jdff dff_B_X8KuPgAP6_0(.din(w_dff_B_varN7BWI9_0),.dout(w_dff_B_X8KuPgAP6_0),.clk(gclk));
	jdff dff_B_XZkzsrjA4_0(.din(w_dff_B_X8KuPgAP6_0),.dout(w_dff_B_XZkzsrjA4_0),.clk(gclk));
	jdff dff_B_vA3MOdfZ5_0(.din(w_dff_B_XZkzsrjA4_0),.dout(w_dff_B_vA3MOdfZ5_0),.clk(gclk));
	jdff dff_B_TaAtuTab9_0(.din(w_dff_B_vA3MOdfZ5_0),.dout(w_dff_B_TaAtuTab9_0),.clk(gclk));
	jdff dff_B_Ign8YJUD7_0(.din(w_dff_B_TaAtuTab9_0),.dout(w_dff_B_Ign8YJUD7_0),.clk(gclk));
	jdff dff_B_RqHIxS1O1_0(.din(w_dff_B_Ign8YJUD7_0),.dout(w_dff_B_RqHIxS1O1_0),.clk(gclk));
	jdff dff_B_P1vGgqKr0_0(.din(w_dff_B_RqHIxS1O1_0),.dout(w_dff_B_P1vGgqKr0_0),.clk(gclk));
	jdff dff_B_jKj3SKn22_0(.din(w_dff_B_P1vGgqKr0_0),.dout(w_dff_B_jKj3SKn22_0),.clk(gclk));
	jdff dff_B_mdPyiKmd0_0(.din(n1195),.dout(w_dff_B_mdPyiKmd0_0),.clk(gclk));
	jdff dff_B_eVuEP4Ca2_0(.din(w_dff_B_mdPyiKmd0_0),.dout(w_dff_B_eVuEP4Ca2_0),.clk(gclk));
	jdff dff_B_PwIuOo4U9_0(.din(w_dff_B_eVuEP4Ca2_0),.dout(w_dff_B_PwIuOo4U9_0),.clk(gclk));
	jdff dff_B_QVpp9gnE7_0(.din(w_dff_B_PwIuOo4U9_0),.dout(w_dff_B_QVpp9gnE7_0),.clk(gclk));
	jdff dff_B_S4Fe6U2p7_1(.din(G115),.dout(w_dff_B_S4Fe6U2p7_1),.clk(gclk));
	jdff dff_B_iunU92P06_1(.din(w_dff_B_S4Fe6U2p7_1),.dout(w_dff_B_iunU92P06_1),.clk(gclk));
	jdff dff_A_IVzXe4al7_0(.dout(w_n751_0[0]),.din(w_dff_A_IVzXe4al7_0),.clk(gclk));
	jdff dff_A_haZpLyY01_2(.dout(w_n751_0[2]),.din(w_dff_A_haZpLyY01_2),.clk(gclk));
	jdff dff_A_gn3eJPS54_2(.dout(w_dff_A_haZpLyY01_2),.din(w_dff_A_gn3eJPS54_2),.clk(gclk));
	jdff dff_A_8JIFM9F91_2(.dout(w_dff_A_gn3eJPS54_2),.din(w_dff_A_8JIFM9F91_2),.clk(gclk));
	jdff dff_A_8Wcm2ddZ5_2(.dout(w_dff_A_8JIFM9F91_2),.din(w_dff_A_8Wcm2ddZ5_2),.clk(gclk));
	jdff dff_B_yyeTZfAc2_1(.din(n929),.dout(w_dff_B_yyeTZfAc2_1),.clk(gclk));
	jdff dff_B_mN6QhgZ65_1(.din(w_dff_B_yyeTZfAc2_1),.dout(w_dff_B_mN6QhgZ65_1),.clk(gclk));
	jdff dff_B_TOeqyTOR4_1(.din(w_dff_B_mN6QhgZ65_1),.dout(w_dff_B_TOeqyTOR4_1),.clk(gclk));
	jdff dff_B_0Gox7zAp4_1(.din(w_dff_B_TOeqyTOR4_1),.dout(w_dff_B_0Gox7zAp4_1),.clk(gclk));
	jdff dff_B_j0TWinXw0_1(.din(w_dff_B_0Gox7zAp4_1),.dout(w_dff_B_j0TWinXw0_1),.clk(gclk));
	jdff dff_B_hzkoANlZ1_1(.din(w_dff_B_j0TWinXw0_1),.dout(w_dff_B_hzkoANlZ1_1),.clk(gclk));
	jdff dff_B_NWCCJe449_1(.din(w_dff_B_hzkoANlZ1_1),.dout(w_dff_B_NWCCJe449_1),.clk(gclk));
	jdff dff_B_SaJAM3N00_1(.din(w_dff_B_NWCCJe449_1),.dout(w_dff_B_SaJAM3N00_1),.clk(gclk));
	jdff dff_B_TVmDremS7_1(.din(n931),.dout(w_dff_B_TVmDremS7_1),.clk(gclk));
	jdff dff_B_Qs7JBXrM6_1(.din(w_dff_B_TVmDremS7_1),.dout(w_dff_B_Qs7JBXrM6_1),.clk(gclk));
	jdff dff_B_6fy14eq14_1(.din(w_dff_B_Qs7JBXrM6_1),.dout(w_dff_B_6fy14eq14_1),.clk(gclk));
	jdff dff_B_kYixEY4a3_1(.din(w_dff_B_6fy14eq14_1),.dout(w_dff_B_kYixEY4a3_1),.clk(gclk));
	jdff dff_B_HinJg8jy0_1(.din(w_dff_B_kYixEY4a3_1),.dout(w_dff_B_HinJg8jy0_1),.clk(gclk));
	jdff dff_B_PjRshg3R5_1(.din(w_dff_B_HinJg8jy0_1),.dout(w_dff_B_PjRshg3R5_1),.clk(gclk));
	jdff dff_B_Zkjoqe727_1(.din(w_dff_B_PjRshg3R5_1),.dout(w_dff_B_Zkjoqe727_1),.clk(gclk));
	jdff dff_B_SfmGU9ge5_1(.din(w_dff_B_Zkjoqe727_1),.dout(w_dff_B_SfmGU9ge5_1),.clk(gclk));
	jdff dff_B_2Sr2ebjQ1_1(.din(w_dff_B_SfmGU9ge5_1),.dout(w_dff_B_2Sr2ebjQ1_1),.clk(gclk));
	jdff dff_B_6DbqdCFJ1_1(.din(w_dff_B_2Sr2ebjQ1_1),.dout(w_dff_B_6DbqdCFJ1_1),.clk(gclk));
	jdff dff_B_bdh2mSot5_0(.din(n935),.dout(w_dff_B_bdh2mSot5_0),.clk(gclk));
	jdff dff_A_WyfAoSHm2_1(.dout(w_G4_0[1]),.din(w_dff_A_WyfAoSHm2_1),.clk(gclk));
	jdff dff_A_XyHvh8tW7_1(.dout(w_dff_A_WyfAoSHm2_1),.din(w_dff_A_XyHvh8tW7_1),.clk(gclk));
	jdff dff_A_9i4LzyXu3_1(.dout(w_dff_A_XyHvh8tW7_1),.din(w_dff_A_9i4LzyXu3_1),.clk(gclk));
	jdff dff_A_UMt1k7Kl5_1(.dout(w_dff_A_9i4LzyXu3_1),.din(w_dff_A_UMt1k7Kl5_1),.clk(gclk));
	jdff dff_A_2hMQhhdO6_1(.dout(w_dff_A_UMt1k7Kl5_1),.din(w_dff_A_2hMQhhdO6_1),.clk(gclk));
	jdff dff_A_R0DOJt8p2_1(.dout(w_dff_A_2hMQhhdO6_1),.din(w_dff_A_R0DOJt8p2_1),.clk(gclk));
	jdff dff_B_J2gxHcmX2_3(.din(G4),.dout(w_dff_B_J2gxHcmX2_3),.clk(gclk));
	jdff dff_B_Veimd5dm5_3(.din(w_dff_B_J2gxHcmX2_3),.dout(w_dff_B_Veimd5dm5_3),.clk(gclk));
	jdff dff_B_FSgLnOcW1_3(.din(w_dff_B_Veimd5dm5_3),.dout(w_dff_B_FSgLnOcW1_3),.clk(gclk));
	jdff dff_B_gvIUJVje8_3(.din(w_dff_B_FSgLnOcW1_3),.dout(w_dff_B_gvIUJVje8_3),.clk(gclk));
	jdff dff_B_x5wLkZTT7_2(.din(n932),.dout(w_dff_B_x5wLkZTT7_2),.clk(gclk));
	jdff dff_B_sRnUQIOa6_2(.din(w_dff_B_x5wLkZTT7_2),.dout(w_dff_B_sRnUQIOa6_2),.clk(gclk));
	jdff dff_B_VevBZNSP7_2(.din(w_dff_B_sRnUQIOa6_2),.dout(w_dff_B_VevBZNSP7_2),.clk(gclk));
	jdff dff_B_yQdwIGbX9_2(.din(w_dff_B_VevBZNSP7_2),.dout(w_dff_B_yQdwIGbX9_2),.clk(gclk));
	jdff dff_B_MWUfwYei7_2(.din(w_dff_B_yQdwIGbX9_2),.dout(w_dff_B_MWUfwYei7_2),.clk(gclk));
	jdff dff_B_jMgDRVhY1_2(.din(w_dff_B_MWUfwYei7_2),.dout(w_dff_B_jMgDRVhY1_2),.clk(gclk));
	jdff dff_B_t5t3bqkt4_2(.din(w_dff_B_jMgDRVhY1_2),.dout(w_dff_B_t5t3bqkt4_2),.clk(gclk));
	jdff dff_B_888HJOmE2_2(.din(w_dff_B_t5t3bqkt4_2),.dout(w_dff_B_888HJOmE2_2),.clk(gclk));
	jdff dff_B_XYG7lamz1_2(.din(w_dff_B_888HJOmE2_2),.dout(w_dff_B_XYG7lamz1_2),.clk(gclk));
	jdff dff_A_hWd10c6p4_1(.dout(w_n747_1[1]),.din(w_dff_A_hWd10c6p4_1),.clk(gclk));
	jdff dff_A_AiVdoE9f6_1(.dout(w_dff_A_hWd10c6p4_1),.din(w_dff_A_AiVdoE9f6_1),.clk(gclk));
	jdff dff_A_kc7C7W6D4_1(.dout(w_dff_A_AiVdoE9f6_1),.din(w_dff_A_kc7C7W6D4_1),.clk(gclk));
	jdff dff_A_ByfD1gwT6_2(.dout(w_n747_1[2]),.din(w_dff_A_ByfD1gwT6_2),.clk(gclk));
	jdff dff_A_cQoM0L162_2(.dout(w_dff_A_ByfD1gwT6_2),.din(w_dff_A_cQoM0L162_2),.clk(gclk));
	jdff dff_A_nNpSSEUv5_2(.dout(w_dff_A_cQoM0L162_2),.din(w_dff_A_nNpSSEUv5_2),.clk(gclk));
	jdff dff_A_S4pNyZOJ2_2(.dout(w_dff_A_nNpSSEUv5_2),.din(w_dff_A_S4pNyZOJ2_2),.clk(gclk));
	jdff dff_A_P6KUHL7z1_0(.dout(w_n747_0[0]),.din(w_dff_A_P6KUHL7z1_0),.clk(gclk));
	jdff dff_A_UhCBGmq06_0(.dout(w_dff_A_P6KUHL7z1_0),.din(w_dff_A_UhCBGmq06_0),.clk(gclk));
	jdff dff_A_11kaPSjM9_0(.dout(w_dff_A_UhCBGmq06_0),.din(w_dff_A_11kaPSjM9_0),.clk(gclk));
	jdff dff_A_qrUWHeLz4_0(.dout(w_dff_A_11kaPSjM9_0),.din(w_dff_A_qrUWHeLz4_0),.clk(gclk));
	jdff dff_A_uxhWYyQZ6_0(.dout(w_dff_A_qrUWHeLz4_0),.din(w_dff_A_uxhWYyQZ6_0),.clk(gclk));
	jdff dff_A_1qWIZ3Oq3_0(.dout(w_dff_A_uxhWYyQZ6_0),.din(w_dff_A_1qWIZ3Oq3_0),.clk(gclk));
	jdff dff_A_7jLEpLmB7_0(.dout(w_dff_A_1qWIZ3Oq3_0),.din(w_dff_A_7jLEpLmB7_0),.clk(gclk));
	jdff dff_A_RX6X5bl79_0(.dout(w_dff_A_7jLEpLmB7_0),.din(w_dff_A_RX6X5bl79_0),.clk(gclk));
	jdff dff_A_FxjLs9uE6_0(.dout(w_dff_A_RX6X5bl79_0),.din(w_dff_A_FxjLs9uE6_0),.clk(gclk));
	jdff dff_A_vlgcW8f95_0(.dout(w_dff_A_FxjLs9uE6_0),.din(w_dff_A_vlgcW8f95_0),.clk(gclk));
	jdff dff_A_51RSWDjd1_0(.dout(w_dff_A_vlgcW8f95_0),.din(w_dff_A_51RSWDjd1_0),.clk(gclk));
	jdff dff_A_9SD8CUQk2_0(.dout(w_dff_A_51RSWDjd1_0),.din(w_dff_A_9SD8CUQk2_0),.clk(gclk));
	jdff dff_A_abiRJ84q1_0(.dout(w_dff_A_9SD8CUQk2_0),.din(w_dff_A_abiRJ84q1_0),.clk(gclk));
	jdff dff_A_iBdvOCbi2_1(.dout(w_n747_0[1]),.din(w_dff_A_iBdvOCbi2_1),.clk(gclk));
	jdff dff_A_iDHxzIDQ1_1(.dout(w_dff_A_iBdvOCbi2_1),.din(w_dff_A_iDHxzIDQ1_1),.clk(gclk));
	jdff dff_A_6kX2OLqW3_1(.dout(w_dff_A_iDHxzIDQ1_1),.din(w_dff_A_6kX2OLqW3_1),.clk(gclk));
	jdff dff_A_cbqwSQcX3_1(.dout(w_dff_A_6kX2OLqW3_1),.din(w_dff_A_cbqwSQcX3_1),.clk(gclk));
	jdff dff_A_UcFqDnAN4_1(.dout(w_dff_A_cbqwSQcX3_1),.din(w_dff_A_UcFqDnAN4_1),.clk(gclk));
	jdff dff_A_NxSXq9pw3_1(.dout(w_dff_A_UcFqDnAN4_1),.din(w_dff_A_NxSXq9pw3_1),.clk(gclk));
	jdff dff_A_xVwWe8BZ7_1(.dout(w_dff_A_NxSXq9pw3_1),.din(w_dff_A_xVwWe8BZ7_1),.clk(gclk));
	jdff dff_B_PSSVQYrh3_1(.din(n1388),.dout(w_dff_B_PSSVQYrh3_1),.clk(gclk));
	jdff dff_B_GWrBT2oc0_1(.din(w_dff_B_PSSVQYrh3_1),.dout(w_dff_B_GWrBT2oc0_1),.clk(gclk));
	jdff dff_B_BPn9TLUF8_1(.din(w_dff_B_GWrBT2oc0_1),.dout(w_dff_B_BPn9TLUF8_1),.clk(gclk));
	jdff dff_B_V3j6wOGE2_1(.din(w_dff_B_BPn9TLUF8_1),.dout(w_dff_B_V3j6wOGE2_1),.clk(gclk));
	jdff dff_B_lgN5BTih8_1(.din(w_dff_B_V3j6wOGE2_1),.dout(w_dff_B_lgN5BTih8_1),.clk(gclk));
	jdff dff_B_8BjmnNm32_1(.din(w_dff_B_lgN5BTih8_1),.dout(w_dff_B_8BjmnNm32_1),.clk(gclk));
	jdff dff_B_WVpGlc070_1(.din(w_dff_B_8BjmnNm32_1),.dout(w_dff_B_WVpGlc070_1),.clk(gclk));
	jdff dff_B_1antOYHT0_1(.din(w_dff_B_WVpGlc070_1),.dout(w_dff_B_1antOYHT0_1),.clk(gclk));
	jdff dff_B_qYgqs6c76_1(.din(w_dff_B_1antOYHT0_1),.dout(w_dff_B_qYgqs6c76_1),.clk(gclk));
	jdff dff_B_lmcnPDen9_1(.din(w_dff_B_qYgqs6c76_1),.dout(w_dff_B_lmcnPDen9_1),.clk(gclk));
	jdff dff_B_0NpLdZnA4_1(.din(w_dff_B_lmcnPDen9_1),.dout(w_dff_B_0NpLdZnA4_1),.clk(gclk));
	jdff dff_B_Mkz1S36q9_1(.din(w_dff_B_0NpLdZnA4_1),.dout(w_dff_B_Mkz1S36q9_1),.clk(gclk));
	jdff dff_B_mOrDmNbH4_1(.din(w_dff_B_Mkz1S36q9_1),.dout(w_dff_B_mOrDmNbH4_1),.clk(gclk));
	jdff dff_B_pfK1Bm0p9_1(.din(w_dff_B_mOrDmNbH4_1),.dout(w_dff_B_pfK1Bm0p9_1),.clk(gclk));
	jdff dff_B_uIKEDw5W5_1(.din(w_dff_B_pfK1Bm0p9_1),.dout(w_dff_B_uIKEDw5W5_1),.clk(gclk));
	jdff dff_B_YsNcVzEP7_1(.din(w_dff_B_uIKEDw5W5_1),.dout(w_dff_B_YsNcVzEP7_1),.clk(gclk));
	jdff dff_B_KfYjRf515_1(.din(w_dff_B_YsNcVzEP7_1),.dout(w_dff_B_KfYjRf515_1),.clk(gclk));
	jdff dff_B_Ebp6XgBG9_1(.din(w_dff_B_KfYjRf515_1),.dout(w_dff_B_Ebp6XgBG9_1),.clk(gclk));
	jdff dff_B_tlTNiJrb5_1(.din(w_dff_B_Ebp6XgBG9_1),.dout(w_dff_B_tlTNiJrb5_1),.clk(gclk));
	jdff dff_B_MWXMhdj96_1(.din(n1539),.dout(w_dff_B_MWXMhdj96_1),.clk(gclk));
	jdff dff_B_8Uz3ufRE5_1(.din(w_dff_B_MWXMhdj96_1),.dout(w_dff_B_8Uz3ufRE5_1),.clk(gclk));
	jdff dff_B_ltAbWIpY0_1(.din(w_dff_B_8Uz3ufRE5_1),.dout(w_dff_B_ltAbWIpY0_1),.clk(gclk));
	jdff dff_B_XSI6BZJ17_1(.din(w_dff_B_ltAbWIpY0_1),.dout(w_dff_B_XSI6BZJ17_1),.clk(gclk));
	jdff dff_B_I4krucv43_1(.din(w_dff_B_XSI6BZJ17_1),.dout(w_dff_B_I4krucv43_1),.clk(gclk));
	jdff dff_B_HeM22eFF6_1(.din(w_dff_B_I4krucv43_1),.dout(w_dff_B_HeM22eFF6_1),.clk(gclk));
	jdff dff_B_T1L9PIeW3_1(.din(w_dff_B_HeM22eFF6_1),.dout(w_dff_B_T1L9PIeW3_1),.clk(gclk));
	jdff dff_B_JABImF1M5_1(.din(w_dff_B_T1L9PIeW3_1),.dout(w_dff_B_JABImF1M5_1),.clk(gclk));
	jdff dff_B_ryMj8vOZ6_1(.din(w_dff_B_JABImF1M5_1),.dout(w_dff_B_ryMj8vOZ6_1),.clk(gclk));
	jdff dff_B_LukVAR2m2_1(.din(w_dff_B_ryMj8vOZ6_1),.dout(w_dff_B_LukVAR2m2_1),.clk(gclk));
	jdff dff_B_rmeqPkzb6_1(.din(w_dff_B_LukVAR2m2_1),.dout(w_dff_B_rmeqPkzb6_1),.clk(gclk));
	jdff dff_B_PYfzAJdU4_1(.din(w_dff_B_rmeqPkzb6_1),.dout(w_dff_B_PYfzAJdU4_1),.clk(gclk));
	jdff dff_B_dgJ8ImcE7_1(.din(w_dff_B_PYfzAJdU4_1),.dout(w_dff_B_dgJ8ImcE7_1),.clk(gclk));
	jdff dff_B_B9eDp4U79_1(.din(w_dff_B_dgJ8ImcE7_1),.dout(w_dff_B_B9eDp4U79_1),.clk(gclk));
	jdff dff_B_g6TnYnbD2_1(.din(w_dff_B_B9eDp4U79_1),.dout(w_dff_B_g6TnYnbD2_1),.clk(gclk));
	jdff dff_B_kVpeL4lv1_1(.din(w_dff_B_g6TnYnbD2_1),.dout(w_dff_B_kVpeL4lv1_1),.clk(gclk));
	jdff dff_B_OwUHNzMz9_1(.din(w_dff_B_kVpeL4lv1_1),.dout(w_dff_B_OwUHNzMz9_1),.clk(gclk));
	jdff dff_B_vuf4YPWQ8_1(.din(w_dff_B_OwUHNzMz9_1),.dout(w_dff_B_vuf4YPWQ8_1),.clk(gclk));
	jdff dff_B_IIdqX6mj8_1(.din(w_dff_B_vuf4YPWQ8_1),.dout(w_dff_B_IIdqX6mj8_1),.clk(gclk));
	jdff dff_B_MEO3d8q96_0(.din(n1614),.dout(w_dff_B_MEO3d8q96_0),.clk(gclk));
	jdff dff_B_VHEjOWlr0_0(.din(w_dff_B_MEO3d8q96_0),.dout(w_dff_B_VHEjOWlr0_0),.clk(gclk));
	jdff dff_B_gb6Z3Xyr5_0(.din(w_dff_B_VHEjOWlr0_0),.dout(w_dff_B_gb6Z3Xyr5_0),.clk(gclk));
	jdff dff_B_7YHFJ8k35_0(.din(w_dff_B_gb6Z3Xyr5_0),.dout(w_dff_B_7YHFJ8k35_0),.clk(gclk));
	jdff dff_B_GmCHsWyE2_0(.din(w_dff_B_7YHFJ8k35_0),.dout(w_dff_B_GmCHsWyE2_0),.clk(gclk));
	jdff dff_B_Ak80ZyMS2_0(.din(w_dff_B_GmCHsWyE2_0),.dout(w_dff_B_Ak80ZyMS2_0),.clk(gclk));
	jdff dff_B_wvvFKVFb1_0(.din(w_dff_B_Ak80ZyMS2_0),.dout(w_dff_B_wvvFKVFb1_0),.clk(gclk));
	jdff dff_B_70wj62FA1_0(.din(w_dff_B_wvvFKVFb1_0),.dout(w_dff_B_70wj62FA1_0),.clk(gclk));
	jdff dff_B_OvL07NLV3_0(.din(w_dff_B_70wj62FA1_0),.dout(w_dff_B_OvL07NLV3_0),.clk(gclk));
	jdff dff_B_3drzL6rn1_0(.din(w_dff_B_OvL07NLV3_0),.dout(w_dff_B_3drzL6rn1_0),.clk(gclk));
	jdff dff_B_oZixLIUj2_0(.din(w_dff_B_3drzL6rn1_0),.dout(w_dff_B_oZixLIUj2_0),.clk(gclk));
	jdff dff_B_FGwDbZqe6_0(.din(w_dff_B_oZixLIUj2_0),.dout(w_dff_B_FGwDbZqe6_0),.clk(gclk));
	jdff dff_B_Zti4Bcwo5_0(.din(w_dff_B_FGwDbZqe6_0),.dout(w_dff_B_Zti4Bcwo5_0),.clk(gclk));
	jdff dff_B_MqvdPi8I7_0(.din(w_dff_B_Zti4Bcwo5_0),.dout(w_dff_B_MqvdPi8I7_0),.clk(gclk));
	jdff dff_B_VNS2lQhf0_0(.din(w_dff_B_MqvdPi8I7_0),.dout(w_dff_B_VNS2lQhf0_0),.clk(gclk));
	jdff dff_B_1rTQDNlf5_0(.din(w_dff_B_VNS2lQhf0_0),.dout(w_dff_B_1rTQDNlf5_0),.clk(gclk));
	jdff dff_B_F5zOduc43_0(.din(w_dff_B_1rTQDNlf5_0),.dout(w_dff_B_F5zOduc43_0),.clk(gclk));
	jdff dff_B_4cT38ERN0_0(.din(w_dff_B_F5zOduc43_0),.dout(w_dff_B_4cT38ERN0_0),.clk(gclk));
	jdff dff_B_FstWOxMJ7_0(.din(w_dff_B_4cT38ERN0_0),.dout(w_dff_B_FstWOxMJ7_0),.clk(gclk));
	jdff dff_B_kA3QnmlP5_0(.din(n1613),.dout(w_dff_B_kA3QnmlP5_0),.clk(gclk));
	jdff dff_A_2BHRjPXu5_1(.dout(w_n797_1[1]),.din(w_dff_A_2BHRjPXu5_1),.clk(gclk));
	jdff dff_A_LJVlJdj69_1(.dout(w_dff_A_2BHRjPXu5_1),.din(w_dff_A_LJVlJdj69_1),.clk(gclk));
	jdff dff_A_4YpHF1Qd3_1(.dout(w_dff_A_LJVlJdj69_1),.din(w_dff_A_4YpHF1Qd3_1),.clk(gclk));
	jdff dff_A_Y5YYbz3i8_1(.dout(w_dff_A_4YpHF1Qd3_1),.din(w_dff_A_Y5YYbz3i8_1),.clk(gclk));
	jdff dff_A_4vHBkBSS9_1(.dout(w_dff_A_Y5YYbz3i8_1),.din(w_dff_A_4vHBkBSS9_1),.clk(gclk));
	jdff dff_A_GV2pKAxt7_1(.dout(w_dff_A_4vHBkBSS9_1),.din(w_dff_A_GV2pKAxt7_1),.clk(gclk));
	jdff dff_A_4WxEcWCe0_1(.dout(w_dff_A_GV2pKAxt7_1),.din(w_dff_A_4WxEcWCe0_1),.clk(gclk));
	jdff dff_A_FE8svY6X9_1(.dout(w_dff_A_4WxEcWCe0_1),.din(w_dff_A_FE8svY6X9_1),.clk(gclk));
	jdff dff_A_cYQJnmg89_1(.dout(w_dff_A_FE8svY6X9_1),.din(w_dff_A_cYQJnmg89_1),.clk(gclk));
	jdff dff_A_6WpXnb3N2_1(.dout(w_dff_A_cYQJnmg89_1),.din(w_dff_A_6WpXnb3N2_1),.clk(gclk));
	jdff dff_A_GjMKJfzx8_1(.dout(w_dff_A_6WpXnb3N2_1),.din(w_dff_A_GjMKJfzx8_1),.clk(gclk));
	jdff dff_A_o4ULUWFk4_1(.dout(w_dff_A_GjMKJfzx8_1),.din(w_dff_A_o4ULUWFk4_1),.clk(gclk));
	jdff dff_A_pPqHdtgv5_1(.dout(w_dff_A_o4ULUWFk4_1),.din(w_dff_A_pPqHdtgv5_1),.clk(gclk));
	jdff dff_A_qovNcWLc4_1(.dout(w_dff_A_pPqHdtgv5_1),.din(w_dff_A_qovNcWLc4_1),.clk(gclk));
	jdff dff_A_NVQNgztX5_2(.dout(w_n797_1[2]),.din(w_dff_A_NVQNgztX5_2),.clk(gclk));
	jdff dff_A_IkFHensy2_2(.dout(w_dff_A_NVQNgztX5_2),.din(w_dff_A_IkFHensy2_2),.clk(gclk));
	jdff dff_A_Hgmw9N1F1_2(.dout(w_dff_A_IkFHensy2_2),.din(w_dff_A_Hgmw9N1F1_2),.clk(gclk));
	jdff dff_A_4CWqr7sf6_2(.dout(w_dff_A_Hgmw9N1F1_2),.din(w_dff_A_4CWqr7sf6_2),.clk(gclk));
	jdff dff_A_DOBDqk9r7_2(.dout(w_dff_A_4CWqr7sf6_2),.din(w_dff_A_DOBDqk9r7_2),.clk(gclk));
	jdff dff_A_Lojwy1gj1_2(.dout(w_dff_A_DOBDqk9r7_2),.din(w_dff_A_Lojwy1gj1_2),.clk(gclk));
	jdff dff_A_ZbrkCbDh2_2(.dout(w_dff_A_Lojwy1gj1_2),.din(w_dff_A_ZbrkCbDh2_2),.clk(gclk));
	jdff dff_A_xDbl4HMC9_2(.dout(w_dff_A_ZbrkCbDh2_2),.din(w_dff_A_xDbl4HMC9_2),.clk(gclk));
	jdff dff_A_U8B4g5eB9_2(.dout(w_dff_A_xDbl4HMC9_2),.din(w_dff_A_U8B4g5eB9_2),.clk(gclk));
	jdff dff_A_Ae5SNb7y0_2(.dout(w_dff_A_U8B4g5eB9_2),.din(w_dff_A_Ae5SNb7y0_2),.clk(gclk));
	jdff dff_A_uQaMhm7w3_1(.dout(w_n797_0[1]),.din(w_dff_A_uQaMhm7w3_1),.clk(gclk));
	jdff dff_A_HTvE6bvC6_1(.dout(w_dff_A_uQaMhm7w3_1),.din(w_dff_A_HTvE6bvC6_1),.clk(gclk));
	jdff dff_A_ORetPWpf6_1(.dout(w_dff_A_HTvE6bvC6_1),.din(w_dff_A_ORetPWpf6_1),.clk(gclk));
	jdff dff_A_yu2u2imy1_1(.dout(w_dff_A_ORetPWpf6_1),.din(w_dff_A_yu2u2imy1_1),.clk(gclk));
	jdff dff_A_hCJ9zakk6_1(.dout(w_dff_A_yu2u2imy1_1),.din(w_dff_A_hCJ9zakk6_1),.clk(gclk));
	jdff dff_A_9JP1G19y9_1(.dout(w_dff_A_hCJ9zakk6_1),.din(w_dff_A_9JP1G19y9_1),.clk(gclk));
	jdff dff_A_0HOBUu6H1_1(.dout(w_dff_A_9JP1G19y9_1),.din(w_dff_A_0HOBUu6H1_1),.clk(gclk));
	jdff dff_A_ANaYa1m63_1(.dout(w_dff_A_0HOBUu6H1_1),.din(w_dff_A_ANaYa1m63_1),.clk(gclk));
	jdff dff_A_hmQ0hxrp3_1(.dout(w_dff_A_ANaYa1m63_1),.din(w_dff_A_hmQ0hxrp3_1),.clk(gclk));
	jdff dff_A_sVUU8jRG6_1(.dout(w_dff_A_hmQ0hxrp3_1),.din(w_dff_A_sVUU8jRG6_1),.clk(gclk));
	jdff dff_A_la6I0zsv1_1(.dout(w_dff_A_sVUU8jRG6_1),.din(w_dff_A_la6I0zsv1_1),.clk(gclk));
	jdff dff_A_8c8YIv9Z3_2(.dout(w_n797_0[2]),.din(w_dff_A_8c8YIv9Z3_2),.clk(gclk));
	jdff dff_B_zVdn96Cx9_3(.din(n797),.dout(w_dff_B_zVdn96Cx9_3),.clk(gclk));
	jdff dff_B_TMWmsUoR4_3(.din(w_dff_B_zVdn96Cx9_3),.dout(w_dff_B_TMWmsUoR4_3),.clk(gclk));
	jdff dff_B_40VEXi2C3_3(.din(w_dff_B_TMWmsUoR4_3),.dout(w_dff_B_40VEXi2C3_3),.clk(gclk));
	jdff dff_B_KkIoLw2R3_3(.din(w_dff_B_40VEXi2C3_3),.dout(w_dff_B_KkIoLw2R3_3),.clk(gclk));
	jdff dff_B_2EgDjwaa5_3(.din(w_dff_B_KkIoLw2R3_3),.dout(w_dff_B_2EgDjwaa5_3),.clk(gclk));
	jdff dff_B_fkxGB2wk5_3(.din(w_dff_B_2EgDjwaa5_3),.dout(w_dff_B_fkxGB2wk5_3),.clk(gclk));
	jdff dff_A_SynBGV085_1(.dout(w_n793_1[1]),.din(w_dff_A_SynBGV085_1),.clk(gclk));
	jdff dff_A_wKGgSIdq1_1(.dout(w_dff_A_SynBGV085_1),.din(w_dff_A_wKGgSIdq1_1),.clk(gclk));
	jdff dff_A_xOqzB6Bb7_1(.dout(w_dff_A_wKGgSIdq1_1),.din(w_dff_A_xOqzB6Bb7_1),.clk(gclk));
	jdff dff_A_ozvAaHc46_1(.dout(w_dff_A_xOqzB6Bb7_1),.din(w_dff_A_ozvAaHc46_1),.clk(gclk));
	jdff dff_A_Y4Q8Nrql6_1(.dout(w_dff_A_ozvAaHc46_1),.din(w_dff_A_Y4Q8Nrql6_1),.clk(gclk));
	jdff dff_A_JCmx0ffA6_1(.dout(w_dff_A_Y4Q8Nrql6_1),.din(w_dff_A_JCmx0ffA6_1),.clk(gclk));
	jdff dff_A_OXO3dpd57_1(.dout(w_dff_A_JCmx0ffA6_1),.din(w_dff_A_OXO3dpd57_1),.clk(gclk));
	jdff dff_A_GR1KqTtM4_1(.dout(w_dff_A_OXO3dpd57_1),.din(w_dff_A_GR1KqTtM4_1),.clk(gclk));
	jdff dff_A_OFDBwyRn8_1(.dout(w_dff_A_GR1KqTtM4_1),.din(w_dff_A_OFDBwyRn8_1),.clk(gclk));
	jdff dff_A_hjzhQks09_1(.dout(w_dff_A_OFDBwyRn8_1),.din(w_dff_A_hjzhQks09_1),.clk(gclk));
	jdff dff_A_cWBI7L8L6_1(.dout(w_dff_A_hjzhQks09_1),.din(w_dff_A_cWBI7L8L6_1),.clk(gclk));
	jdff dff_A_ZAAGuerl8_1(.dout(w_dff_A_cWBI7L8L6_1),.din(w_dff_A_ZAAGuerl8_1),.clk(gclk));
	jdff dff_A_mHwsDrOt3_1(.dout(w_dff_A_ZAAGuerl8_1),.din(w_dff_A_mHwsDrOt3_1),.clk(gclk));
	jdff dff_A_awGli8B57_1(.dout(w_dff_A_mHwsDrOt3_1),.din(w_dff_A_awGli8B57_1),.clk(gclk));
	jdff dff_A_zef5JSYo2_2(.dout(w_n793_1[2]),.din(w_dff_A_zef5JSYo2_2),.clk(gclk));
	jdff dff_A_1Lql7xGW3_2(.dout(w_dff_A_zef5JSYo2_2),.din(w_dff_A_1Lql7xGW3_2),.clk(gclk));
	jdff dff_A_0DNp4rkF4_2(.dout(w_dff_A_1Lql7xGW3_2),.din(w_dff_A_0DNp4rkF4_2),.clk(gclk));
	jdff dff_A_zBUdklzJ2_2(.dout(w_dff_A_0DNp4rkF4_2),.din(w_dff_A_zBUdklzJ2_2),.clk(gclk));
	jdff dff_A_GVTjFlIY3_2(.dout(w_dff_A_zBUdklzJ2_2),.din(w_dff_A_GVTjFlIY3_2),.clk(gclk));
	jdff dff_A_jTp48KP56_2(.dout(w_dff_A_GVTjFlIY3_2),.din(w_dff_A_jTp48KP56_2),.clk(gclk));
	jdff dff_A_XKPibHSf7_2(.dout(w_dff_A_jTp48KP56_2),.din(w_dff_A_XKPibHSf7_2),.clk(gclk));
	jdff dff_A_BncmWU7u7_2(.dout(w_dff_A_XKPibHSf7_2),.din(w_dff_A_BncmWU7u7_2),.clk(gclk));
	jdff dff_A_Pp0eBHjk0_2(.dout(w_dff_A_BncmWU7u7_2),.din(w_dff_A_Pp0eBHjk0_2),.clk(gclk));
	jdff dff_A_lGSOXHj04_2(.dout(w_dff_A_Pp0eBHjk0_2),.din(w_dff_A_lGSOXHj04_2),.clk(gclk));
	jdff dff_A_VWPGiUH60_1(.dout(w_n793_0[1]),.din(w_dff_A_VWPGiUH60_1),.clk(gclk));
	jdff dff_A_JUlOSG6o2_1(.dout(w_dff_A_VWPGiUH60_1),.din(w_dff_A_JUlOSG6o2_1),.clk(gclk));
	jdff dff_A_RwwjwGFi3_1(.dout(w_dff_A_JUlOSG6o2_1),.din(w_dff_A_RwwjwGFi3_1),.clk(gclk));
	jdff dff_A_QVtGEvtA2_1(.dout(w_dff_A_RwwjwGFi3_1),.din(w_dff_A_QVtGEvtA2_1),.clk(gclk));
	jdff dff_A_sJ25soSa6_1(.dout(w_dff_A_QVtGEvtA2_1),.din(w_dff_A_sJ25soSa6_1),.clk(gclk));
	jdff dff_A_yEwyVCMS4_1(.dout(w_dff_A_sJ25soSa6_1),.din(w_dff_A_yEwyVCMS4_1),.clk(gclk));
	jdff dff_A_6G3CynG85_1(.dout(w_dff_A_yEwyVCMS4_1),.din(w_dff_A_6G3CynG85_1),.clk(gclk));
	jdff dff_A_I1FjocQF5_1(.dout(w_dff_A_6G3CynG85_1),.din(w_dff_A_I1FjocQF5_1),.clk(gclk));
	jdff dff_A_FBNhkPIT1_1(.dout(w_dff_A_I1FjocQF5_1),.din(w_dff_A_FBNhkPIT1_1),.clk(gclk));
	jdff dff_A_b4WFldKb4_1(.dout(w_dff_A_FBNhkPIT1_1),.din(w_dff_A_b4WFldKb4_1),.clk(gclk));
	jdff dff_A_Uck6BVVc7_1(.dout(w_dff_A_b4WFldKb4_1),.din(w_dff_A_Uck6BVVc7_1),.clk(gclk));
	jdff dff_A_gUyPHObs8_2(.dout(w_n793_0[2]),.din(w_dff_A_gUyPHObs8_2),.clk(gclk));
	jdff dff_A_b8It70LO1_2(.dout(w_dff_A_gUyPHObs8_2),.din(w_dff_A_b8It70LO1_2),.clk(gclk));
	jdff dff_A_1qjmRQCl2_2(.dout(w_dff_A_b8It70LO1_2),.din(w_dff_A_1qjmRQCl2_2),.clk(gclk));
	jdff dff_A_uxzSyXNv7_2(.dout(w_dff_A_1qjmRQCl2_2),.din(w_dff_A_uxzSyXNv7_2),.clk(gclk));
	jdff dff_B_K9AGMGuF9_3(.din(n793),.dout(w_dff_B_K9AGMGuF9_3),.clk(gclk));
	jdff dff_B_ls42C8lp4_3(.din(w_dff_B_K9AGMGuF9_3),.dout(w_dff_B_ls42C8lp4_3),.clk(gclk));
	jdff dff_B_iZ4BEQyX0_3(.din(w_dff_B_ls42C8lp4_3),.dout(w_dff_B_iZ4BEQyX0_3),.clk(gclk));
	jdff dff_B_t3wNn53i8_3(.din(w_dff_B_iZ4BEQyX0_3),.dout(w_dff_B_t3wNn53i8_3),.clk(gclk));
	jdff dff_B_BoAcDQIB4_3(.din(w_dff_B_t3wNn53i8_3),.dout(w_dff_B_BoAcDQIB4_3),.clk(gclk));
	jdff dff_B_5nmvW88k8_3(.din(w_dff_B_BoAcDQIB4_3),.dout(w_dff_B_5nmvW88k8_3),.clk(gclk));
	jdff dff_B_IRk8CjcP4_3(.din(w_dff_B_5nmvW88k8_3),.dout(w_dff_B_IRk8CjcP4_3),.clk(gclk));
	jdff dff_A_6ma5F38f2_2(.dout(w_G4088_0[2]),.din(w_dff_A_6ma5F38f2_2),.clk(gclk));
	jdff dff_A_FTuHRH8f2_1(.dout(w_G4087_0[1]),.din(w_dff_A_FTuHRH8f2_1),.clk(gclk));
	jdff dff_B_mx8n3Ai93_0(.din(n1621),.dout(w_dff_B_mx8n3Ai93_0),.clk(gclk));
	jdff dff_B_pYp3CDu43_0(.din(w_dff_B_mx8n3Ai93_0),.dout(w_dff_B_pYp3CDu43_0),.clk(gclk));
	jdff dff_B_TtueYOmb7_0(.din(w_dff_B_pYp3CDu43_0),.dout(w_dff_B_TtueYOmb7_0),.clk(gclk));
	jdff dff_B_mYjxnGuU6_0(.din(w_dff_B_TtueYOmb7_0),.dout(w_dff_B_mYjxnGuU6_0),.clk(gclk));
	jdff dff_B_CMWquzL43_0(.din(w_dff_B_mYjxnGuU6_0),.dout(w_dff_B_CMWquzL43_0),.clk(gclk));
	jdff dff_B_WfZNkflh7_0(.din(w_dff_B_CMWquzL43_0),.dout(w_dff_B_WfZNkflh7_0),.clk(gclk));
	jdff dff_B_qoGGw7bJ8_0(.din(w_dff_B_WfZNkflh7_0),.dout(w_dff_B_qoGGw7bJ8_0),.clk(gclk));
	jdff dff_B_vBExeG9j5_0(.din(w_dff_B_qoGGw7bJ8_0),.dout(w_dff_B_vBExeG9j5_0),.clk(gclk));
	jdff dff_B_70K05SSy7_0(.din(w_dff_B_vBExeG9j5_0),.dout(w_dff_B_70K05SSy7_0),.clk(gclk));
	jdff dff_B_IEckeMl75_0(.din(w_dff_B_70K05SSy7_0),.dout(w_dff_B_IEckeMl75_0),.clk(gclk));
	jdff dff_B_bksrw7pz2_0(.din(w_dff_B_IEckeMl75_0),.dout(w_dff_B_bksrw7pz2_0),.clk(gclk));
	jdff dff_B_LIty7jJU6_0(.din(w_dff_B_bksrw7pz2_0),.dout(w_dff_B_LIty7jJU6_0),.clk(gclk));
	jdff dff_B_E7Cpwizy1_0(.din(w_dff_B_LIty7jJU6_0),.dout(w_dff_B_E7Cpwizy1_0),.clk(gclk));
	jdff dff_B_vGKvDKpH7_0(.din(w_dff_B_E7Cpwizy1_0),.dout(w_dff_B_vGKvDKpH7_0),.clk(gclk));
	jdff dff_B_fqtQOO3N8_0(.din(w_dff_B_vGKvDKpH7_0),.dout(w_dff_B_fqtQOO3N8_0),.clk(gclk));
	jdff dff_B_E9XrPimD5_0(.din(w_dff_B_fqtQOO3N8_0),.dout(w_dff_B_E9XrPimD5_0),.clk(gclk));
	jdff dff_B_c4uEurZK0_0(.din(w_dff_B_E9XrPimD5_0),.dout(w_dff_B_c4uEurZK0_0),.clk(gclk));
	jdff dff_B_bvS3vdT85_0(.din(w_dff_B_c4uEurZK0_0),.dout(w_dff_B_bvS3vdT85_0),.clk(gclk));
	jdff dff_B_UYe82NPj3_0(.din(w_dff_B_bvS3vdT85_0),.dout(w_dff_B_UYe82NPj3_0),.clk(gclk));
	jdff dff_B_1tJj2pw78_0(.din(n1620),.dout(w_dff_B_1tJj2pw78_0),.clk(gclk));
	jdff dff_B_CPdioXsj6_2(.din(G64),.dout(w_dff_B_CPdioXsj6_2),.clk(gclk));
	jdff dff_B_qMQsQAo42_2(.din(G14),.dout(w_dff_B_qMQsQAo42_2),.clk(gclk));
	jdff dff_B_DbS2HEhc5_2(.din(w_dff_B_qMQsQAo42_2),.dout(w_dff_B_DbS2HEhc5_2),.clk(gclk));
	jdff dff_A_VeM1GuY34_1(.dout(w_n843_1[1]),.din(w_dff_A_VeM1GuY34_1),.clk(gclk));
	jdff dff_A_6a1bTLaC6_1(.dout(w_dff_A_VeM1GuY34_1),.din(w_dff_A_6a1bTLaC6_1),.clk(gclk));
	jdff dff_A_t720y4za9_1(.dout(w_dff_A_6a1bTLaC6_1),.din(w_dff_A_t720y4za9_1),.clk(gclk));
	jdff dff_A_nKAuaDZ02_1(.dout(w_dff_A_t720y4za9_1),.din(w_dff_A_nKAuaDZ02_1),.clk(gclk));
	jdff dff_A_wUwsDg1W0_1(.dout(w_dff_A_nKAuaDZ02_1),.din(w_dff_A_wUwsDg1W0_1),.clk(gclk));
	jdff dff_A_cVplHmUC6_1(.dout(w_dff_A_wUwsDg1W0_1),.din(w_dff_A_cVplHmUC6_1),.clk(gclk));
	jdff dff_A_xUHOb8jG3_1(.dout(w_dff_A_cVplHmUC6_1),.din(w_dff_A_xUHOb8jG3_1),.clk(gclk));
	jdff dff_A_JX3J5xJw3_1(.dout(w_dff_A_xUHOb8jG3_1),.din(w_dff_A_JX3J5xJw3_1),.clk(gclk));
	jdff dff_A_cWkChUra6_1(.dout(w_dff_A_JX3J5xJw3_1),.din(w_dff_A_cWkChUra6_1),.clk(gclk));
	jdff dff_A_7AHSfJsd7_1(.dout(w_dff_A_cWkChUra6_1),.din(w_dff_A_7AHSfJsd7_1),.clk(gclk));
	jdff dff_A_uyzX1rmX9_1(.dout(w_dff_A_7AHSfJsd7_1),.din(w_dff_A_uyzX1rmX9_1),.clk(gclk));
	jdff dff_A_eee57DFl7_1(.dout(w_dff_A_uyzX1rmX9_1),.din(w_dff_A_eee57DFl7_1),.clk(gclk));
	jdff dff_A_645HeLnO7_1(.dout(w_dff_A_eee57DFl7_1),.din(w_dff_A_645HeLnO7_1),.clk(gclk));
	jdff dff_A_0HiOG1SP1_1(.dout(w_dff_A_645HeLnO7_1),.din(w_dff_A_0HiOG1SP1_1),.clk(gclk));
	jdff dff_A_fK4K6jJQ3_2(.dout(w_n843_1[2]),.din(w_dff_A_fK4K6jJQ3_2),.clk(gclk));
	jdff dff_A_sEiEdIec8_2(.dout(w_dff_A_fK4K6jJQ3_2),.din(w_dff_A_sEiEdIec8_2),.clk(gclk));
	jdff dff_A_MwHMJvDL0_2(.dout(w_dff_A_sEiEdIec8_2),.din(w_dff_A_MwHMJvDL0_2),.clk(gclk));
	jdff dff_A_kJ2H4MXc8_2(.dout(w_dff_A_MwHMJvDL0_2),.din(w_dff_A_kJ2H4MXc8_2),.clk(gclk));
	jdff dff_A_1feiUy8v1_2(.dout(w_dff_A_kJ2H4MXc8_2),.din(w_dff_A_1feiUy8v1_2),.clk(gclk));
	jdff dff_A_7meb2ZSk9_2(.dout(w_dff_A_1feiUy8v1_2),.din(w_dff_A_7meb2ZSk9_2),.clk(gclk));
	jdff dff_A_uc3PKkxM1_2(.dout(w_dff_A_7meb2ZSk9_2),.din(w_dff_A_uc3PKkxM1_2),.clk(gclk));
	jdff dff_A_cJgrrRaW3_2(.dout(w_dff_A_uc3PKkxM1_2),.din(w_dff_A_cJgrrRaW3_2),.clk(gclk));
	jdff dff_A_8xG2O6Ia9_2(.dout(w_dff_A_cJgrrRaW3_2),.din(w_dff_A_8xG2O6Ia9_2),.clk(gclk));
	jdff dff_A_vuhtRYQD6_2(.dout(w_dff_A_8xG2O6Ia9_2),.din(w_dff_A_vuhtRYQD6_2),.clk(gclk));
	jdff dff_A_rX4X66Vn6_1(.dout(w_n843_0[1]),.din(w_dff_A_rX4X66Vn6_1),.clk(gclk));
	jdff dff_A_jDPgrLWs8_1(.dout(w_dff_A_rX4X66Vn6_1),.din(w_dff_A_jDPgrLWs8_1),.clk(gclk));
	jdff dff_A_GF5krNfO1_1(.dout(w_dff_A_jDPgrLWs8_1),.din(w_dff_A_GF5krNfO1_1),.clk(gclk));
	jdff dff_A_yw0hccLG8_1(.dout(w_dff_A_GF5krNfO1_1),.din(w_dff_A_yw0hccLG8_1),.clk(gclk));
	jdff dff_A_acblp5LJ1_1(.dout(w_dff_A_yw0hccLG8_1),.din(w_dff_A_acblp5LJ1_1),.clk(gclk));
	jdff dff_A_r9fnHnR71_1(.dout(w_dff_A_acblp5LJ1_1),.din(w_dff_A_r9fnHnR71_1),.clk(gclk));
	jdff dff_A_nfyVuQPC0_1(.dout(w_dff_A_r9fnHnR71_1),.din(w_dff_A_nfyVuQPC0_1),.clk(gclk));
	jdff dff_A_o0CrjVkS6_1(.dout(w_dff_A_nfyVuQPC0_1),.din(w_dff_A_o0CrjVkS6_1),.clk(gclk));
	jdff dff_A_zhWSMOFn1_1(.dout(w_dff_A_o0CrjVkS6_1),.din(w_dff_A_zhWSMOFn1_1),.clk(gclk));
	jdff dff_A_swpKsueu3_1(.dout(w_dff_A_zhWSMOFn1_1),.din(w_dff_A_swpKsueu3_1),.clk(gclk));
	jdff dff_A_mwCoMitu7_1(.dout(w_dff_A_swpKsueu3_1),.din(w_dff_A_mwCoMitu7_1),.clk(gclk));
	jdff dff_A_b3PzTxgP3_2(.dout(w_n843_0[2]),.din(w_dff_A_b3PzTxgP3_2),.clk(gclk));
	jdff dff_B_NFYmXjap0_3(.din(n843),.dout(w_dff_B_NFYmXjap0_3),.clk(gclk));
	jdff dff_B_3R7hbTLo8_3(.din(w_dff_B_NFYmXjap0_3),.dout(w_dff_B_3R7hbTLo8_3),.clk(gclk));
	jdff dff_B_AfquKikj8_3(.din(w_dff_B_3R7hbTLo8_3),.dout(w_dff_B_AfquKikj8_3),.clk(gclk));
	jdff dff_B_lDHjV6Yj7_3(.din(w_dff_B_AfquKikj8_3),.dout(w_dff_B_lDHjV6Yj7_3),.clk(gclk));
	jdff dff_B_DKrBzNRP3_3(.din(w_dff_B_lDHjV6Yj7_3),.dout(w_dff_B_DKrBzNRP3_3),.clk(gclk));
	jdff dff_B_NoFcKoJw2_3(.din(w_dff_B_DKrBzNRP3_3),.dout(w_dff_B_NoFcKoJw2_3),.clk(gclk));
	jdff dff_A_nkBkbhDA8_1(.dout(w_n840_1[1]),.din(w_dff_A_nkBkbhDA8_1),.clk(gclk));
	jdff dff_A_scfkKZjy8_1(.dout(w_dff_A_nkBkbhDA8_1),.din(w_dff_A_scfkKZjy8_1),.clk(gclk));
	jdff dff_A_5Owzi61p1_1(.dout(w_dff_A_scfkKZjy8_1),.din(w_dff_A_5Owzi61p1_1),.clk(gclk));
	jdff dff_A_JbVPKepv2_1(.dout(w_dff_A_5Owzi61p1_1),.din(w_dff_A_JbVPKepv2_1),.clk(gclk));
	jdff dff_A_73sVhA7w9_1(.dout(w_dff_A_JbVPKepv2_1),.din(w_dff_A_73sVhA7w9_1),.clk(gclk));
	jdff dff_A_nIwBCpXi4_1(.dout(w_dff_A_73sVhA7w9_1),.din(w_dff_A_nIwBCpXi4_1),.clk(gclk));
	jdff dff_A_Il49YHsk4_1(.dout(w_dff_A_nIwBCpXi4_1),.din(w_dff_A_Il49YHsk4_1),.clk(gclk));
	jdff dff_A_wKmW8qMj5_1(.dout(w_dff_A_Il49YHsk4_1),.din(w_dff_A_wKmW8qMj5_1),.clk(gclk));
	jdff dff_A_TZaCrk1i3_1(.dout(w_dff_A_wKmW8qMj5_1),.din(w_dff_A_TZaCrk1i3_1),.clk(gclk));
	jdff dff_A_3oDxbYye3_1(.dout(w_dff_A_TZaCrk1i3_1),.din(w_dff_A_3oDxbYye3_1),.clk(gclk));
	jdff dff_A_DIG9kD0N3_1(.dout(w_dff_A_3oDxbYye3_1),.din(w_dff_A_DIG9kD0N3_1),.clk(gclk));
	jdff dff_A_cMMATo8X4_1(.dout(w_dff_A_DIG9kD0N3_1),.din(w_dff_A_cMMATo8X4_1),.clk(gclk));
	jdff dff_A_RWlZCJbu3_1(.dout(w_dff_A_cMMATo8X4_1),.din(w_dff_A_RWlZCJbu3_1),.clk(gclk));
	jdff dff_A_oPFxAwah3_1(.dout(w_dff_A_RWlZCJbu3_1),.din(w_dff_A_oPFxAwah3_1),.clk(gclk));
	jdff dff_A_a7UFN0Uh7_2(.dout(w_n840_1[2]),.din(w_dff_A_a7UFN0Uh7_2),.clk(gclk));
	jdff dff_A_sRSC3A8A5_2(.dout(w_dff_A_a7UFN0Uh7_2),.din(w_dff_A_sRSC3A8A5_2),.clk(gclk));
	jdff dff_A_Ta3DWYTB1_2(.dout(w_dff_A_sRSC3A8A5_2),.din(w_dff_A_Ta3DWYTB1_2),.clk(gclk));
	jdff dff_A_w0BZivgt0_2(.dout(w_dff_A_Ta3DWYTB1_2),.din(w_dff_A_w0BZivgt0_2),.clk(gclk));
	jdff dff_A_5kjiY2cf5_2(.dout(w_dff_A_w0BZivgt0_2),.din(w_dff_A_5kjiY2cf5_2),.clk(gclk));
	jdff dff_A_1I1ajFIP4_2(.dout(w_dff_A_5kjiY2cf5_2),.din(w_dff_A_1I1ajFIP4_2),.clk(gclk));
	jdff dff_A_FVbyTzEw9_2(.dout(w_dff_A_1I1ajFIP4_2),.din(w_dff_A_FVbyTzEw9_2),.clk(gclk));
	jdff dff_A_vXMhNBiR8_2(.dout(w_dff_A_FVbyTzEw9_2),.din(w_dff_A_vXMhNBiR8_2),.clk(gclk));
	jdff dff_A_kVbLXsRG9_2(.dout(w_dff_A_vXMhNBiR8_2),.din(w_dff_A_kVbLXsRG9_2),.clk(gclk));
	jdff dff_A_Jy2uufCu7_2(.dout(w_dff_A_kVbLXsRG9_2),.din(w_dff_A_Jy2uufCu7_2),.clk(gclk));
	jdff dff_A_e6TerabC0_1(.dout(w_n840_0[1]),.din(w_dff_A_e6TerabC0_1),.clk(gclk));
	jdff dff_A_UGLdQg8w9_1(.dout(w_dff_A_e6TerabC0_1),.din(w_dff_A_UGLdQg8w9_1),.clk(gclk));
	jdff dff_A_HWTMfyzp4_1(.dout(w_dff_A_UGLdQg8w9_1),.din(w_dff_A_HWTMfyzp4_1),.clk(gclk));
	jdff dff_A_6ICfHWwi1_1(.dout(w_dff_A_HWTMfyzp4_1),.din(w_dff_A_6ICfHWwi1_1),.clk(gclk));
	jdff dff_A_iPYLaqK78_1(.dout(w_dff_A_6ICfHWwi1_1),.din(w_dff_A_iPYLaqK78_1),.clk(gclk));
	jdff dff_A_yaxkx7d88_1(.dout(w_dff_A_iPYLaqK78_1),.din(w_dff_A_yaxkx7d88_1),.clk(gclk));
	jdff dff_A_UuH9XUSa5_1(.dout(w_dff_A_yaxkx7d88_1),.din(w_dff_A_UuH9XUSa5_1),.clk(gclk));
	jdff dff_A_aaa9mnAP7_1(.dout(w_dff_A_UuH9XUSa5_1),.din(w_dff_A_aaa9mnAP7_1),.clk(gclk));
	jdff dff_A_FOV1LhKx1_1(.dout(w_dff_A_aaa9mnAP7_1),.din(w_dff_A_FOV1LhKx1_1),.clk(gclk));
	jdff dff_A_XTjON36r5_1(.dout(w_dff_A_FOV1LhKx1_1),.din(w_dff_A_XTjON36r5_1),.clk(gclk));
	jdff dff_A_I5c4OnJa6_1(.dout(w_dff_A_XTjON36r5_1),.din(w_dff_A_I5c4OnJa6_1),.clk(gclk));
	jdff dff_A_MxddZJHs5_2(.dout(w_n840_0[2]),.din(w_dff_A_MxddZJHs5_2),.clk(gclk));
	jdff dff_A_XZbvFUvd6_2(.dout(w_dff_A_MxddZJHs5_2),.din(w_dff_A_XZbvFUvd6_2),.clk(gclk));
	jdff dff_A_UmX0EuCz9_2(.dout(w_dff_A_XZbvFUvd6_2),.din(w_dff_A_UmX0EuCz9_2),.clk(gclk));
	jdff dff_A_6bUW0NZ23_2(.dout(w_dff_A_UmX0EuCz9_2),.din(w_dff_A_6bUW0NZ23_2),.clk(gclk));
	jdff dff_B_Qtn3h0Tm6_3(.din(n840),.dout(w_dff_B_Qtn3h0Tm6_3),.clk(gclk));
	jdff dff_B_ELWWf9620_3(.din(w_dff_B_Qtn3h0Tm6_3),.dout(w_dff_B_ELWWf9620_3),.clk(gclk));
	jdff dff_B_r1lnAy1I3_3(.din(w_dff_B_ELWWf9620_3),.dout(w_dff_B_r1lnAy1I3_3),.clk(gclk));
	jdff dff_B_WA2DV3Vf0_3(.din(w_dff_B_r1lnAy1I3_3),.dout(w_dff_B_WA2DV3Vf0_3),.clk(gclk));
	jdff dff_B_8R7J4r6g0_3(.din(w_dff_B_WA2DV3Vf0_3),.dout(w_dff_B_8R7J4r6g0_3),.clk(gclk));
	jdff dff_B_03qcQDFT5_3(.din(w_dff_B_8R7J4r6g0_3),.dout(w_dff_B_03qcQDFT5_3),.clk(gclk));
	jdff dff_B_Ua5DCBO99_3(.din(w_dff_B_03qcQDFT5_3),.dout(w_dff_B_Ua5DCBO99_3),.clk(gclk));
	jdff dff_A_BadhDM3A4_1(.dout(w_G4090_0[1]),.din(w_dff_A_BadhDM3A4_1),.clk(gclk));
	jdff dff_A_uFn2pNSI7_2(.dout(w_G4089_0[2]),.din(w_dff_A_uFn2pNSI7_2),.clk(gclk));
	jdff dff_B_xA0vYSin2_1(.din(n1626),.dout(w_dff_B_xA0vYSin2_1),.clk(gclk));
	jdff dff_B_n078xPUD8_0(.din(n1637),.dout(w_dff_B_n078xPUD8_0),.clk(gclk));
	jdff dff_B_pt6MItKr0_0(.din(w_dff_B_n078xPUD8_0),.dout(w_dff_B_pt6MItKr0_0),.clk(gclk));
	jdff dff_B_rosl3jPX7_0(.din(w_dff_B_pt6MItKr0_0),.dout(w_dff_B_rosl3jPX7_0),.clk(gclk));
	jdff dff_B_Rgbv2Gtx3_0(.din(w_dff_B_rosl3jPX7_0),.dout(w_dff_B_Rgbv2Gtx3_0),.clk(gclk));
	jdff dff_B_BhTC6eJE4_0(.din(w_dff_B_Rgbv2Gtx3_0),.dout(w_dff_B_BhTC6eJE4_0),.clk(gclk));
	jdff dff_B_MoC5iSjJ4_0(.din(w_dff_B_BhTC6eJE4_0),.dout(w_dff_B_MoC5iSjJ4_0),.clk(gclk));
	jdff dff_B_k3ACB6772_0(.din(w_dff_B_MoC5iSjJ4_0),.dout(w_dff_B_k3ACB6772_0),.clk(gclk));
	jdff dff_B_o8CZ3GWW8_0(.din(w_dff_B_k3ACB6772_0),.dout(w_dff_B_o8CZ3GWW8_0),.clk(gclk));
	jdff dff_B_8hTS6JfU3_0(.din(w_dff_B_o8CZ3GWW8_0),.dout(w_dff_B_8hTS6JfU3_0),.clk(gclk));
	jdff dff_B_Ji3yWvM96_0(.din(w_dff_B_8hTS6JfU3_0),.dout(w_dff_B_Ji3yWvM96_0),.clk(gclk));
	jdff dff_B_h2uuehdI9_0(.din(w_dff_B_Ji3yWvM96_0),.dout(w_dff_B_h2uuehdI9_0),.clk(gclk));
	jdff dff_B_CTQRxkAh3_0(.din(w_dff_B_h2uuehdI9_0),.dout(w_dff_B_CTQRxkAh3_0),.clk(gclk));
	jdff dff_B_CHKDEOLe6_0(.din(w_dff_B_CTQRxkAh3_0),.dout(w_dff_B_CHKDEOLe6_0),.clk(gclk));
	jdff dff_B_37hP9ygD1_0(.din(w_dff_B_CHKDEOLe6_0),.dout(w_dff_B_37hP9ygD1_0),.clk(gclk));
	jdff dff_B_Tlcay7sT3_0(.din(w_dff_B_37hP9ygD1_0),.dout(w_dff_B_Tlcay7sT3_0),.clk(gclk));
	jdff dff_B_4silvIz19_0(.din(w_dff_B_Tlcay7sT3_0),.dout(w_dff_B_4silvIz19_0),.clk(gclk));
	jdff dff_B_2h1HXx4o1_0(.din(w_dff_B_4silvIz19_0),.dout(w_dff_B_2h1HXx4o1_0),.clk(gclk));
	jdff dff_B_NEceM8xN0_0(.din(w_dff_B_2h1HXx4o1_0),.dout(w_dff_B_NEceM8xN0_0),.clk(gclk));
	jdff dff_B_QBM2HGO14_1(.din(n1633),.dout(w_dff_B_QBM2HGO14_1),.clk(gclk));
	jdff dff_B_WjCopaOU8_1(.din(n1627),.dout(w_dff_B_WjCopaOU8_1),.clk(gclk));
	jdff dff_B_N8wIuoDw7_1(.din(w_dff_B_WjCopaOU8_1),.dout(w_dff_B_N8wIuoDw7_1),.clk(gclk));
	jdff dff_B_mJ4NKWRl2_1(.din(w_dff_B_N8wIuoDw7_1),.dout(w_dff_B_mJ4NKWRl2_1),.clk(gclk));
	jdff dff_B_UwRxg3MX7_1(.din(w_dff_B_mJ4NKWRl2_1),.dout(w_dff_B_UwRxg3MX7_1),.clk(gclk));
	jdff dff_B_lqs2ydvD0_1(.din(w_dff_B_UwRxg3MX7_1),.dout(w_dff_B_lqs2ydvD0_1),.clk(gclk));
	jdff dff_B_LARZFADt4_1(.din(w_dff_B_lqs2ydvD0_1),.dout(w_dff_B_LARZFADt4_1),.clk(gclk));
	jdff dff_B_ujqEeYer1_1(.din(w_dff_B_LARZFADt4_1),.dout(w_dff_B_ujqEeYer1_1),.clk(gclk));
	jdff dff_B_hHxvGh243_1(.din(w_dff_B_ujqEeYer1_1),.dout(w_dff_B_hHxvGh243_1),.clk(gclk));
	jdff dff_B_w8EFnRTn7_1(.din(w_dff_B_hHxvGh243_1),.dout(w_dff_B_w8EFnRTn7_1),.clk(gclk));
	jdff dff_B_qvajMSfs0_1(.din(w_dff_B_w8EFnRTn7_1),.dout(w_dff_B_qvajMSfs0_1),.clk(gclk));
	jdff dff_B_wy5GZvL64_1(.din(w_dff_B_qvajMSfs0_1),.dout(w_dff_B_wy5GZvL64_1),.clk(gclk));
	jdff dff_B_BGnLcEqz5_1(.din(w_dff_B_wy5GZvL64_1),.dout(w_dff_B_BGnLcEqz5_1),.clk(gclk));
	jdff dff_B_Ons9LCHV0_1(.din(w_dff_B_BGnLcEqz5_1),.dout(w_dff_B_Ons9LCHV0_1),.clk(gclk));
	jdff dff_B_fqiDJapU6_1(.din(w_dff_B_Ons9LCHV0_1),.dout(w_dff_B_fqiDJapU6_1),.clk(gclk));
	jdff dff_B_tZ2zDv4U8_1(.din(w_dff_B_fqiDJapU6_1),.dout(w_dff_B_tZ2zDv4U8_1),.clk(gclk));
	jdff dff_B_8mQQFoVP2_1(.din(w_dff_B_tZ2zDv4U8_1),.dout(w_dff_B_8mQQFoVP2_1),.clk(gclk));
	jdff dff_B_0knoR80E4_1(.din(w_dff_B_8mQQFoVP2_1),.dout(w_dff_B_0knoR80E4_1),.clk(gclk));
	jdff dff_B_mPyZHcJA0_1(.din(w_dff_B_0knoR80E4_1),.dout(w_dff_B_mPyZHcJA0_1),.clk(gclk));
	jdff dff_B_q3Yf7HM58_1(.din(w_dff_B_mPyZHcJA0_1),.dout(w_dff_B_q3Yf7HM58_1),.clk(gclk));
	jdff dff_A_zANiK10X9_0(.dout(w_n988_1[0]),.din(w_dff_A_zANiK10X9_0),.clk(gclk));
	jdff dff_A_2PnpBSVi1_0(.dout(w_dff_A_zANiK10X9_0),.din(w_dff_A_2PnpBSVi1_0),.clk(gclk));
	jdff dff_A_DFUg5kjj4_0(.dout(w_dff_A_2PnpBSVi1_0),.din(w_dff_A_DFUg5kjj4_0),.clk(gclk));
	jdff dff_A_wvnkraax7_0(.dout(w_dff_A_DFUg5kjj4_0),.din(w_dff_A_wvnkraax7_0),.clk(gclk));
	jdff dff_A_bvbp1zIY8_0(.dout(w_dff_A_wvnkraax7_0),.din(w_dff_A_bvbp1zIY8_0),.clk(gclk));
	jdff dff_A_gpHh6toS5_0(.dout(w_dff_A_bvbp1zIY8_0),.din(w_dff_A_gpHh6toS5_0),.clk(gclk));
	jdff dff_A_D8IjNm4D3_2(.dout(w_n988_1[2]),.din(w_dff_A_D8IjNm4D3_2),.clk(gclk));
	jdff dff_A_n13TQpRP8_2(.dout(w_dff_A_D8IjNm4D3_2),.din(w_dff_A_n13TQpRP8_2),.clk(gclk));
	jdff dff_A_V9gmVsjw0_2(.dout(w_dff_A_n13TQpRP8_2),.din(w_dff_A_V9gmVsjw0_2),.clk(gclk));
	jdff dff_A_PnQXDKMq4_2(.dout(w_dff_A_V9gmVsjw0_2),.din(w_dff_A_PnQXDKMq4_2),.clk(gclk));
	jdff dff_A_lZzUJE1h5_2(.dout(w_dff_A_PnQXDKMq4_2),.din(w_dff_A_lZzUJE1h5_2),.clk(gclk));
	jdff dff_A_DxTfdG1h9_2(.dout(w_dff_A_lZzUJE1h5_2),.din(w_dff_A_DxTfdG1h9_2),.clk(gclk));
	jdff dff_A_nXm9wK0P5_2(.dout(w_dff_A_DxTfdG1h9_2),.din(w_dff_A_nXm9wK0P5_2),.clk(gclk));
	jdff dff_A_4Ql8qXpc2_2(.dout(w_dff_A_nXm9wK0P5_2),.din(w_dff_A_4Ql8qXpc2_2),.clk(gclk));
	jdff dff_A_zk4VSNBZ8_2(.dout(w_dff_A_4Ql8qXpc2_2),.din(w_dff_A_zk4VSNBZ8_2),.clk(gclk));
	jdff dff_A_DHmrZ5j96_2(.dout(w_dff_A_zk4VSNBZ8_2),.din(w_dff_A_DHmrZ5j96_2),.clk(gclk));
	jdff dff_A_8VvYjaXq2_2(.dout(w_dff_A_DHmrZ5j96_2),.din(w_dff_A_8VvYjaXq2_2),.clk(gclk));
	jdff dff_A_WQ6uCOAq7_2(.dout(w_dff_A_8VvYjaXq2_2),.din(w_dff_A_WQ6uCOAq7_2),.clk(gclk));
	jdff dff_A_YJEoqH5y8_2(.dout(w_dff_A_WQ6uCOAq7_2),.din(w_dff_A_YJEoqH5y8_2),.clk(gclk));
	jdff dff_A_rXImKdHt6_2(.dout(w_dff_A_YJEoqH5y8_2),.din(w_dff_A_rXImKdHt6_2),.clk(gclk));
	jdff dff_A_pZ2PQGNC5_2(.dout(w_dff_A_rXImKdHt6_2),.din(w_dff_A_pZ2PQGNC5_2),.clk(gclk));
	jdff dff_A_LDgOPlyo7_2(.dout(w_dff_A_pZ2PQGNC5_2),.din(w_dff_A_LDgOPlyo7_2),.clk(gclk));
	jdff dff_A_o2NXtWKY2_2(.dout(w_dff_A_LDgOPlyo7_2),.din(w_dff_A_o2NXtWKY2_2),.clk(gclk));
	jdff dff_A_Z7o0FbIx1_2(.dout(w_dff_A_o2NXtWKY2_2),.din(w_dff_A_Z7o0FbIx1_2),.clk(gclk));
	jdff dff_A_cvvYCVZ33_1(.dout(w_n988_0[1]),.din(w_dff_A_cvvYCVZ33_1),.clk(gclk));
	jdff dff_A_ZjkvOD6o5_1(.dout(w_dff_A_cvvYCVZ33_1),.din(w_dff_A_ZjkvOD6o5_1),.clk(gclk));
	jdff dff_A_UfWuBhFF1_1(.dout(w_dff_A_ZjkvOD6o5_1),.din(w_dff_A_UfWuBhFF1_1),.clk(gclk));
	jdff dff_A_TkueEScT3_1(.dout(w_dff_A_UfWuBhFF1_1),.din(w_dff_A_TkueEScT3_1),.clk(gclk));
	jdff dff_A_Y8I6zfIG7_1(.dout(w_dff_A_TkueEScT3_1),.din(w_dff_A_Y8I6zfIG7_1),.clk(gclk));
	jdff dff_A_pdRsSaV75_1(.dout(w_dff_A_Y8I6zfIG7_1),.din(w_dff_A_pdRsSaV75_1),.clk(gclk));
	jdff dff_A_4yuWQuL74_1(.dout(w_dff_A_pdRsSaV75_1),.din(w_dff_A_4yuWQuL74_1),.clk(gclk));
	jdff dff_A_ECEsCU3W5_1(.dout(w_dff_A_4yuWQuL74_1),.din(w_dff_A_ECEsCU3W5_1),.clk(gclk));
	jdff dff_A_8oUDouHL9_1(.dout(w_dff_A_ECEsCU3W5_1),.din(w_dff_A_8oUDouHL9_1),.clk(gclk));
	jdff dff_A_gkGDwd6X0_1(.dout(w_dff_A_8oUDouHL9_1),.din(w_dff_A_gkGDwd6X0_1),.clk(gclk));
	jdff dff_A_KD6QhGAK3_1(.dout(w_dff_A_gkGDwd6X0_1),.din(w_dff_A_KD6QhGAK3_1),.clk(gclk));
	jdff dff_A_JZ1ywGXq7_1(.dout(w_dff_A_KD6QhGAK3_1),.din(w_dff_A_JZ1ywGXq7_1),.clk(gclk));
	jdff dff_A_jBBKyDco1_1(.dout(w_dff_A_JZ1ywGXq7_1),.din(w_dff_A_jBBKyDco1_1),.clk(gclk));
	jdff dff_A_yGWARj6r5_1(.dout(w_dff_A_jBBKyDco1_1),.din(w_dff_A_yGWARj6r5_1),.clk(gclk));
	jdff dff_A_K9wO8y109_1(.dout(w_dff_A_yGWARj6r5_1),.din(w_dff_A_K9wO8y109_1),.clk(gclk));
	jdff dff_A_B9uKgh0B8_1(.dout(w_dff_A_K9wO8y109_1),.din(w_dff_A_B9uKgh0B8_1),.clk(gclk));
	jdff dff_A_yR3LGZKu2_2(.dout(w_n988_0[2]),.din(w_dff_A_yR3LGZKu2_2),.clk(gclk));
	jdff dff_A_CRiNvvDn3_2(.dout(w_dff_A_yR3LGZKu2_2),.din(w_dff_A_CRiNvvDn3_2),.clk(gclk));
	jdff dff_A_lrUAb7493_2(.dout(w_dff_A_CRiNvvDn3_2),.din(w_dff_A_lrUAb7493_2),.clk(gclk));
	jdff dff_A_jWMlgr7T7_2(.dout(w_dff_A_lrUAb7493_2),.din(w_dff_A_jWMlgr7T7_2),.clk(gclk));
	jdff dff_A_HuxvSMAX5_2(.dout(w_dff_A_jWMlgr7T7_2),.din(w_dff_A_HuxvSMAX5_2),.clk(gclk));
	jdff dff_A_SUgE56ZD8_2(.dout(w_dff_A_HuxvSMAX5_2),.din(w_dff_A_SUgE56ZD8_2),.clk(gclk));
	jdff dff_A_P2IcOBYT4_2(.dout(w_dff_A_SUgE56ZD8_2),.din(w_dff_A_P2IcOBYT4_2),.clk(gclk));
	jdff dff_B_doFl3vwD2_1(.din(n1625),.dout(w_dff_B_doFl3vwD2_1),.clk(gclk));
	jdff dff_B_SUI2ZvpX9_1(.din(w_dff_B_doFl3vwD2_1),.dout(w_dff_B_SUI2ZvpX9_1),.clk(gclk));
	jdff dff_B_dXfk9olI7_1(.din(w_dff_B_SUI2ZvpX9_1),.dout(w_dff_B_dXfk9olI7_1),.clk(gclk));
	jdff dff_B_EPtCOdgg2_1(.din(w_dff_B_dXfk9olI7_1),.dout(w_dff_B_EPtCOdgg2_1),.clk(gclk));
	jdff dff_B_x6QRsMbM7_1(.din(w_dff_B_EPtCOdgg2_1),.dout(w_dff_B_x6QRsMbM7_1),.clk(gclk));
	jdff dff_B_f1n1Y4Mm8_1(.din(w_dff_B_x6QRsMbM7_1),.dout(w_dff_B_f1n1Y4Mm8_1),.clk(gclk));
	jdff dff_B_OvCy6SmH8_1(.din(w_dff_B_f1n1Y4Mm8_1),.dout(w_dff_B_OvCy6SmH8_1),.clk(gclk));
	jdff dff_B_LZouneJq7_1(.din(w_dff_B_OvCy6SmH8_1),.dout(w_dff_B_LZouneJq7_1),.clk(gclk));
	jdff dff_B_KSKsdCZ91_1(.din(w_dff_B_LZouneJq7_1),.dout(w_dff_B_KSKsdCZ91_1),.clk(gclk));
	jdff dff_B_ugv3GUcQ4_1(.din(w_dff_B_KSKsdCZ91_1),.dout(w_dff_B_ugv3GUcQ4_1),.clk(gclk));
	jdff dff_B_F34WJs6U2_1(.din(w_dff_B_ugv3GUcQ4_1),.dout(w_dff_B_F34WJs6U2_1),.clk(gclk));
	jdff dff_B_qYY2eNcY6_1(.din(w_dff_B_F34WJs6U2_1),.dout(w_dff_B_qYY2eNcY6_1),.clk(gclk));
	jdff dff_B_WhrdeZgS6_1(.din(w_dff_B_qYY2eNcY6_1),.dout(w_dff_B_WhrdeZgS6_1),.clk(gclk));
	jdff dff_B_dqS2YwLH8_1(.din(w_dff_B_WhrdeZgS6_1),.dout(w_dff_B_dqS2YwLH8_1),.clk(gclk));
	jdff dff_B_DwhQ158Q2_1(.din(w_dff_B_dqS2YwLH8_1),.dout(w_dff_B_DwhQ158Q2_1),.clk(gclk));
	jdff dff_B_28FqjB0d4_1(.din(w_dff_B_DwhQ158Q2_1),.dout(w_dff_B_28FqjB0d4_1),.clk(gclk));
	jdff dff_B_LP409KKA4_1(.din(w_dff_B_28FqjB0d4_1),.dout(w_dff_B_LP409KKA4_1),.clk(gclk));
	jdff dff_B_XL4HHL9f7_1(.din(w_dff_B_LP409KKA4_1),.dout(w_dff_B_XL4HHL9f7_1),.clk(gclk));
	jdff dff_B_uSrom04Y5_1(.din(w_dff_B_XL4HHL9f7_1),.dout(w_dff_B_uSrom04Y5_1),.clk(gclk));
	jdff dff_A_OHWGpSNV7_0(.dout(w_n985_1[0]),.din(w_dff_A_OHWGpSNV7_0),.clk(gclk));
	jdff dff_A_h2N8nIye8_0(.dout(w_dff_A_OHWGpSNV7_0),.din(w_dff_A_h2N8nIye8_0),.clk(gclk));
	jdff dff_A_8eXgH3K64_0(.dout(w_dff_A_h2N8nIye8_0),.din(w_dff_A_8eXgH3K64_0),.clk(gclk));
	jdff dff_A_xP8nRnYM1_0(.dout(w_dff_A_8eXgH3K64_0),.din(w_dff_A_xP8nRnYM1_0),.clk(gclk));
	jdff dff_A_WhF8GNAk2_0(.dout(w_dff_A_xP8nRnYM1_0),.din(w_dff_A_WhF8GNAk2_0),.clk(gclk));
	jdff dff_A_EtEfJ8W07_0(.dout(w_dff_A_WhF8GNAk2_0),.din(w_dff_A_EtEfJ8W07_0),.clk(gclk));
	jdff dff_A_T9vIVRvM5_0(.dout(w_dff_A_EtEfJ8W07_0),.din(w_dff_A_T9vIVRvM5_0),.clk(gclk));
	jdff dff_A_YO0mP3XC1_2(.dout(w_n985_1[2]),.din(w_dff_A_YO0mP3XC1_2),.clk(gclk));
	jdff dff_A_YoNUvkDx4_2(.dout(w_dff_A_YO0mP3XC1_2),.din(w_dff_A_YoNUvkDx4_2),.clk(gclk));
	jdff dff_A_iBAILy4o7_2(.dout(w_dff_A_YoNUvkDx4_2),.din(w_dff_A_iBAILy4o7_2),.clk(gclk));
	jdff dff_A_feSVqn7k0_2(.dout(w_dff_A_iBAILy4o7_2),.din(w_dff_A_feSVqn7k0_2),.clk(gclk));
	jdff dff_A_ChpdGrbB6_2(.dout(w_dff_A_feSVqn7k0_2),.din(w_dff_A_ChpdGrbB6_2),.clk(gclk));
	jdff dff_A_dABCwaV04_2(.dout(w_dff_A_ChpdGrbB6_2),.din(w_dff_A_dABCwaV04_2),.clk(gclk));
	jdff dff_A_InRfc20D5_2(.dout(w_dff_A_dABCwaV04_2),.din(w_dff_A_InRfc20D5_2),.clk(gclk));
	jdff dff_A_0luYfXCa4_2(.dout(w_dff_A_InRfc20D5_2),.din(w_dff_A_0luYfXCa4_2),.clk(gclk));
	jdff dff_A_i3zcEiMj3_2(.dout(w_dff_A_0luYfXCa4_2),.din(w_dff_A_i3zcEiMj3_2),.clk(gclk));
	jdff dff_A_4QLG6wQk6_2(.dout(w_dff_A_i3zcEiMj3_2),.din(w_dff_A_4QLG6wQk6_2),.clk(gclk));
	jdff dff_A_gtJvAjE86_2(.dout(w_dff_A_4QLG6wQk6_2),.din(w_dff_A_gtJvAjE86_2),.clk(gclk));
	jdff dff_A_amNgEKYR2_2(.dout(w_dff_A_gtJvAjE86_2),.din(w_dff_A_amNgEKYR2_2),.clk(gclk));
	jdff dff_A_WXrBAOZO8_2(.dout(w_dff_A_amNgEKYR2_2),.din(w_dff_A_WXrBAOZO8_2),.clk(gclk));
	jdff dff_A_FhYieZXV1_2(.dout(w_dff_A_WXrBAOZO8_2),.din(w_dff_A_FhYieZXV1_2),.clk(gclk));
	jdff dff_A_6eZMbTnv8_2(.dout(w_dff_A_FhYieZXV1_2),.din(w_dff_A_6eZMbTnv8_2),.clk(gclk));
	jdff dff_A_VDJHXKIq1_2(.dout(w_dff_A_6eZMbTnv8_2),.din(w_dff_A_VDJHXKIq1_2),.clk(gclk));
	jdff dff_A_zRfb5UVR3_2(.dout(w_dff_A_VDJHXKIq1_2),.din(w_dff_A_zRfb5UVR3_2),.clk(gclk));
	jdff dff_A_dyh85Ttw8_2(.dout(w_dff_A_zRfb5UVR3_2),.din(w_dff_A_dyh85Ttw8_2),.clk(gclk));
	jdff dff_A_MLToMRuZ9_2(.dout(w_dff_A_dyh85Ttw8_2),.din(w_dff_A_MLToMRuZ9_2),.clk(gclk));
	jdff dff_A_aeKAGSCg7_1(.dout(w_n985_0[1]),.din(w_dff_A_aeKAGSCg7_1),.clk(gclk));
	jdff dff_A_pfKC3rsj5_1(.dout(w_dff_A_aeKAGSCg7_1),.din(w_dff_A_pfKC3rsj5_1),.clk(gclk));
	jdff dff_A_Jnk0oSli6_1(.dout(w_dff_A_pfKC3rsj5_1),.din(w_dff_A_Jnk0oSli6_1),.clk(gclk));
	jdff dff_A_9CdXQzzd2_1(.dout(w_dff_A_Jnk0oSli6_1),.din(w_dff_A_9CdXQzzd2_1),.clk(gclk));
	jdff dff_A_B34x5AsY1_1(.dout(w_dff_A_9CdXQzzd2_1),.din(w_dff_A_B34x5AsY1_1),.clk(gclk));
	jdff dff_A_OswyhW3j2_1(.dout(w_dff_A_B34x5AsY1_1),.din(w_dff_A_OswyhW3j2_1),.clk(gclk));
	jdff dff_A_rAQPOaZk1_1(.dout(w_dff_A_OswyhW3j2_1),.din(w_dff_A_rAQPOaZk1_1),.clk(gclk));
	jdff dff_A_snh6lWUk2_1(.dout(w_dff_A_rAQPOaZk1_1),.din(w_dff_A_snh6lWUk2_1),.clk(gclk));
	jdff dff_A_odiIjmux2_1(.dout(w_dff_A_snh6lWUk2_1),.din(w_dff_A_odiIjmux2_1),.clk(gclk));
	jdff dff_A_nvgoEXNm3_1(.dout(w_dff_A_odiIjmux2_1),.din(w_dff_A_nvgoEXNm3_1),.clk(gclk));
	jdff dff_A_aT01ZwOF8_1(.dout(w_dff_A_nvgoEXNm3_1),.din(w_dff_A_aT01ZwOF8_1),.clk(gclk));
	jdff dff_A_R2L2rZlr7_1(.dout(w_dff_A_aT01ZwOF8_1),.din(w_dff_A_R2L2rZlr7_1),.clk(gclk));
	jdff dff_A_4iqUQ62V3_1(.dout(w_dff_A_R2L2rZlr7_1),.din(w_dff_A_4iqUQ62V3_1),.clk(gclk));
	jdff dff_A_rKHVtsEn3_1(.dout(w_dff_A_4iqUQ62V3_1),.din(w_dff_A_rKHVtsEn3_1),.clk(gclk));
	jdff dff_A_Y0q6fX3z8_1(.dout(w_dff_A_rKHVtsEn3_1),.din(w_dff_A_Y0q6fX3z8_1),.clk(gclk));
	jdff dff_A_kNhOidYe1_1(.dout(w_dff_A_Y0q6fX3z8_1),.din(w_dff_A_kNhOidYe1_1),.clk(gclk));
	jdff dff_A_iYxEkZyg0_1(.dout(w_dff_A_kNhOidYe1_1),.din(w_dff_A_iYxEkZyg0_1),.clk(gclk));
	jdff dff_A_PqB0lklw9_2(.dout(w_n985_0[2]),.din(w_dff_A_PqB0lklw9_2),.clk(gclk));
	jdff dff_A_vWwPitHK1_2(.dout(w_dff_A_PqB0lklw9_2),.din(w_dff_A_vWwPitHK1_2),.clk(gclk));
	jdff dff_A_hpj13S168_2(.dout(w_dff_A_vWwPitHK1_2),.din(w_dff_A_hpj13S168_2),.clk(gclk));
	jdff dff_A_vqPZKqIW7_2(.dout(w_dff_A_hpj13S168_2),.din(w_dff_A_vqPZKqIW7_2),.clk(gclk));
	jdff dff_A_HMpgyEEf3_2(.dout(w_dff_A_vqPZKqIW7_2),.din(w_dff_A_HMpgyEEf3_2),.clk(gclk));
	jdff dff_A_w8nAFFtp9_2(.dout(w_dff_A_HMpgyEEf3_2),.din(w_dff_A_w8nAFFtp9_2),.clk(gclk));
	jdff dff_A_XPh3pkSs5_2(.dout(w_dff_A_w8nAFFtp9_2),.din(w_dff_A_XPh3pkSs5_2),.clk(gclk));
	jdff dff_A_YVBetRxS7_2(.dout(w_dff_A_XPh3pkSs5_2),.din(w_dff_A_YVBetRxS7_2),.clk(gclk));
	jdff dff_A_uSe7Axul1_2(.dout(w_dff_A_YVBetRxS7_2),.din(w_dff_A_uSe7Axul1_2),.clk(gclk));
	jdff dff_A_p0emwRUY2_2(.dout(w_dff_A_uSe7Axul1_2),.din(w_dff_A_p0emwRUY2_2),.clk(gclk));
	jdff dff_A_ICJEW9YY6_2(.dout(w_dff_A_p0emwRUY2_2),.din(w_dff_A_ICJEW9YY6_2),.clk(gclk));
	jdff dff_A_TzPdTV922_1(.dout(w_G1690_0[1]),.din(w_dff_A_TzPdTV922_1),.clk(gclk));
	jdff dff_A_jZQpmhwB0_2(.dout(w_G1689_0[2]),.din(w_dff_A_jZQpmhwB0_2),.clk(gclk));
	jdff dff_B_BsnuMHo72_1(.din(n1642),.dout(w_dff_B_BsnuMHo72_1),.clk(gclk));
	jdff dff_B_0OQA9ptp4_0(.din(n1649),.dout(w_dff_B_0OQA9ptp4_0),.clk(gclk));
	jdff dff_B_ZyxEP5N92_0(.din(w_dff_B_0OQA9ptp4_0),.dout(w_dff_B_ZyxEP5N92_0),.clk(gclk));
	jdff dff_B_OyDk8pw65_0(.din(w_dff_B_ZyxEP5N92_0),.dout(w_dff_B_OyDk8pw65_0),.clk(gclk));
	jdff dff_B_hQKoiH9Y0_0(.din(w_dff_B_OyDk8pw65_0),.dout(w_dff_B_hQKoiH9Y0_0),.clk(gclk));
	jdff dff_B_r7cCnYQ74_0(.din(w_dff_B_hQKoiH9Y0_0),.dout(w_dff_B_r7cCnYQ74_0),.clk(gclk));
	jdff dff_B_wS7Pabpk7_0(.din(w_dff_B_r7cCnYQ74_0),.dout(w_dff_B_wS7Pabpk7_0),.clk(gclk));
	jdff dff_B_eRCu8QB44_0(.din(w_dff_B_wS7Pabpk7_0),.dout(w_dff_B_eRCu8QB44_0),.clk(gclk));
	jdff dff_B_NCtyN3dR2_0(.din(w_dff_B_eRCu8QB44_0),.dout(w_dff_B_NCtyN3dR2_0),.clk(gclk));
	jdff dff_B_PpsFzXUk3_0(.din(w_dff_B_NCtyN3dR2_0),.dout(w_dff_B_PpsFzXUk3_0),.clk(gclk));
	jdff dff_B_v9lsnwlz1_0(.din(w_dff_B_PpsFzXUk3_0),.dout(w_dff_B_v9lsnwlz1_0),.clk(gclk));
	jdff dff_B_S72YKBWS7_0(.din(w_dff_B_v9lsnwlz1_0),.dout(w_dff_B_S72YKBWS7_0),.clk(gclk));
	jdff dff_B_twFnlQqg3_0(.din(w_dff_B_S72YKBWS7_0),.dout(w_dff_B_twFnlQqg3_0),.clk(gclk));
	jdff dff_B_JtyBBIX31_0(.din(w_dff_B_twFnlQqg3_0),.dout(w_dff_B_JtyBBIX31_0),.clk(gclk));
	jdff dff_B_moRuQVvE6_0(.din(w_dff_B_JtyBBIX31_0),.dout(w_dff_B_moRuQVvE6_0),.clk(gclk));
	jdff dff_B_Ohgyme1S1_0(.din(w_dff_B_moRuQVvE6_0),.dout(w_dff_B_Ohgyme1S1_0),.clk(gclk));
	jdff dff_B_6RFN7g056_0(.din(w_dff_B_Ohgyme1S1_0),.dout(w_dff_B_6RFN7g056_0),.clk(gclk));
	jdff dff_B_H6W0Emv19_0(.din(w_dff_B_6RFN7g056_0),.dout(w_dff_B_H6W0Emv19_0),.clk(gclk));
	jdff dff_B_CGcUBzOR8_0(.din(w_dff_B_H6W0Emv19_0),.dout(w_dff_B_CGcUBzOR8_0),.clk(gclk));
	jdff dff_B_bVOuko2y1_1(.din(n1646),.dout(w_dff_B_bVOuko2y1_1),.clk(gclk));
	jdff dff_B_U24SoQQf7_2(.din(n1634),.dout(w_dff_B_U24SoQQf7_2),.clk(gclk));
	jdff dff_B_oUZfakXc6_2(.din(w_dff_B_U24SoQQf7_2),.dout(w_dff_B_oUZfakXc6_2),.clk(gclk));
	jdff dff_B_JuqoCnrz3_2(.din(n1631),.dout(w_dff_B_JuqoCnrz3_2),.clk(gclk));
	jdff dff_B_OKfdq3cA1_1(.din(n1643),.dout(w_dff_B_OKfdq3cA1_1),.clk(gclk));
	jdff dff_B_8PX1GDoU5_1(.din(w_dff_B_OKfdq3cA1_1),.dout(w_dff_B_8PX1GDoU5_1),.clk(gclk));
	jdff dff_B_2r2ydSlc4_1(.din(w_dff_B_8PX1GDoU5_1),.dout(w_dff_B_2r2ydSlc4_1),.clk(gclk));
	jdff dff_B_hJTvTNBh9_1(.din(w_dff_B_2r2ydSlc4_1),.dout(w_dff_B_hJTvTNBh9_1),.clk(gclk));
	jdff dff_B_gdyVWrjk2_1(.din(w_dff_B_hJTvTNBh9_1),.dout(w_dff_B_gdyVWrjk2_1),.clk(gclk));
	jdff dff_B_TaKh9HbN9_1(.din(w_dff_B_gdyVWrjk2_1),.dout(w_dff_B_TaKh9HbN9_1),.clk(gclk));
	jdff dff_B_AZcMHsa48_1(.din(w_dff_B_TaKh9HbN9_1),.dout(w_dff_B_AZcMHsa48_1),.clk(gclk));
	jdff dff_B_6lxmEqr84_1(.din(w_dff_B_AZcMHsa48_1),.dout(w_dff_B_6lxmEqr84_1),.clk(gclk));
	jdff dff_B_NtIZYNf47_1(.din(w_dff_B_6lxmEqr84_1),.dout(w_dff_B_NtIZYNf47_1),.clk(gclk));
	jdff dff_B_B0icVx8h9_1(.din(w_dff_B_NtIZYNf47_1),.dout(w_dff_B_B0icVx8h9_1),.clk(gclk));
	jdff dff_B_kIFZwWzd7_1(.din(w_dff_B_B0icVx8h9_1),.dout(w_dff_B_kIFZwWzd7_1),.clk(gclk));
	jdff dff_B_2KSacEBF3_1(.din(w_dff_B_kIFZwWzd7_1),.dout(w_dff_B_2KSacEBF3_1),.clk(gclk));
	jdff dff_B_sLSg93yN4_1(.din(w_dff_B_2KSacEBF3_1),.dout(w_dff_B_sLSg93yN4_1),.clk(gclk));
	jdff dff_B_ZANhEngS8_1(.din(w_dff_B_sLSg93yN4_1),.dout(w_dff_B_ZANhEngS8_1),.clk(gclk));
	jdff dff_B_uYxTnCUy7_1(.din(w_dff_B_ZANhEngS8_1),.dout(w_dff_B_uYxTnCUy7_1),.clk(gclk));
	jdff dff_B_8uTCp8Hn8_1(.din(w_dff_B_uYxTnCUy7_1),.dout(w_dff_B_8uTCp8Hn8_1),.clk(gclk));
	jdff dff_B_NRIVh24E0_1(.din(w_dff_B_8uTCp8Hn8_1),.dout(w_dff_B_NRIVh24E0_1),.clk(gclk));
	jdff dff_B_1I29x71r3_1(.din(w_dff_B_NRIVh24E0_1),.dout(w_dff_B_1I29x71r3_1),.clk(gclk));
	jdff dff_B_dX64z8cV0_1(.din(w_dff_B_1I29x71r3_1),.dout(w_dff_B_dX64z8cV0_1),.clk(gclk));
	jdff dff_B_iNw3Vakc1_0(.din(n1628),.dout(w_dff_B_iNw3Vakc1_0),.clk(gclk));
	jdff dff_B_F6YrgLL71_0(.din(w_dff_B_iNw3Vakc1_0),.dout(w_dff_B_F6YrgLL71_0),.clk(gclk));
	jdff dff_B_Rc4dgdeP1_0(.din(w_dff_B_F6YrgLL71_0),.dout(w_dff_B_Rc4dgdeP1_0),.clk(gclk));
	jdff dff_B_DlpLbvfb8_0(.din(w_dff_B_Rc4dgdeP1_0),.dout(w_dff_B_DlpLbvfb8_0),.clk(gclk));
	jdff dff_B_rGm3yYio7_0(.din(w_dff_B_DlpLbvfb8_0),.dout(w_dff_B_rGm3yYio7_0),.clk(gclk));
	jdff dff_B_93RtKOiA9_0(.din(w_dff_B_rGm3yYio7_0),.dout(w_dff_B_93RtKOiA9_0),.clk(gclk));
	jdff dff_B_cSGC9RYB8_0(.din(w_dff_B_93RtKOiA9_0),.dout(w_dff_B_cSGC9RYB8_0),.clk(gclk));
	jdff dff_B_OMrgHnLd1_0(.din(w_dff_B_cSGC9RYB8_0),.dout(w_dff_B_OMrgHnLd1_0),.clk(gclk));
	jdff dff_B_qJzYmhjs5_0(.din(w_dff_B_OMrgHnLd1_0),.dout(w_dff_B_qJzYmhjs5_0),.clk(gclk));
	jdff dff_B_Stv8tSr94_0(.din(w_dff_B_qJzYmhjs5_0),.dout(w_dff_B_Stv8tSr94_0),.clk(gclk));
	jdff dff_B_rP4eNdoI2_0(.din(w_dff_B_Stv8tSr94_0),.dout(w_dff_B_rP4eNdoI2_0),.clk(gclk));
	jdff dff_B_1QiusGXx5_0(.din(w_dff_B_rP4eNdoI2_0),.dout(w_dff_B_1QiusGXx5_0),.clk(gclk));
	jdff dff_B_mUy9AMw66_0(.din(w_dff_B_1QiusGXx5_0),.dout(w_dff_B_mUy9AMw66_0),.clk(gclk));
	jdff dff_B_ZFPbteDe2_0(.din(w_dff_B_mUy9AMw66_0),.dout(w_dff_B_ZFPbteDe2_0),.clk(gclk));
	jdff dff_B_cvJSCxbs5_0(.din(w_dff_B_ZFPbteDe2_0),.dout(w_dff_B_cvJSCxbs5_0),.clk(gclk));
	jdff dff_B_Tya8Tj9E5_0(.din(w_dff_B_cvJSCxbs5_0),.dout(w_dff_B_Tya8Tj9E5_0),.clk(gclk));
	jdff dff_B_2tVAfDUS6_0(.din(w_dff_B_Tya8Tj9E5_0),.dout(w_dff_B_2tVAfDUS6_0),.clk(gclk));
	jdff dff_B_Shy0yNC95_0(.din(w_dff_B_2tVAfDUS6_0),.dout(w_dff_B_Shy0yNC95_0),.clk(gclk));
	jdff dff_B_MRWuuE6D0_0(.din(w_dff_B_Shy0yNC95_0),.dout(w_dff_B_MRWuuE6D0_0),.clk(gclk));
	jdff dff_A_FHG5wHSW6_1(.dout(w_n1609_0[1]),.din(w_dff_A_FHG5wHSW6_1),.clk(gclk));
	jdff dff_A_LU26bgDI7_1(.dout(w_dff_A_FHG5wHSW6_1),.din(w_dff_A_LU26bgDI7_1),.clk(gclk));
	jdff dff_A_sYZxVC6p4_1(.dout(w_dff_A_LU26bgDI7_1),.din(w_dff_A_sYZxVC6p4_1),.clk(gclk));
	jdff dff_A_26HXs43r8_1(.dout(w_dff_A_sYZxVC6p4_1),.din(w_dff_A_26HXs43r8_1),.clk(gclk));
	jdff dff_A_lZ7eUrRG4_1(.dout(w_dff_A_26HXs43r8_1),.din(w_dff_A_lZ7eUrRG4_1),.clk(gclk));
	jdff dff_A_FUVFASAc3_1(.dout(w_dff_A_lZ7eUrRG4_1),.din(w_dff_A_FUVFASAc3_1),.clk(gclk));
	jdff dff_A_m2doOAnp6_1(.dout(w_dff_A_FUVFASAc3_1),.din(w_dff_A_m2doOAnp6_1),.clk(gclk));
	jdff dff_A_SL8JSuej4_1(.dout(w_dff_A_m2doOAnp6_1),.din(w_dff_A_SL8JSuej4_1),.clk(gclk));
	jdff dff_A_OPVl9SYl6_1(.dout(w_dff_A_SL8JSuej4_1),.din(w_dff_A_OPVl9SYl6_1),.clk(gclk));
	jdff dff_A_9pWn6sQk9_1(.dout(w_dff_A_OPVl9SYl6_1),.din(w_dff_A_9pWn6sQk9_1),.clk(gclk));
	jdff dff_A_kAkLYPmA7_1(.dout(w_dff_A_9pWn6sQk9_1),.din(w_dff_A_kAkLYPmA7_1),.clk(gclk));
	jdff dff_A_bzrmhNfn7_1(.dout(w_dff_A_kAkLYPmA7_1),.din(w_dff_A_bzrmhNfn7_1),.clk(gclk));
	jdff dff_A_xoxhGbk60_1(.dout(w_dff_A_bzrmhNfn7_1),.din(w_dff_A_xoxhGbk60_1),.clk(gclk));
	jdff dff_A_UTf2MXfn7_1(.dout(w_dff_A_xoxhGbk60_1),.din(w_dff_A_UTf2MXfn7_1),.clk(gclk));
	jdff dff_A_ecD7gx984_1(.dout(w_dff_A_UTf2MXfn7_1),.din(w_dff_A_ecD7gx984_1),.clk(gclk));
	jdff dff_A_22JSAGlj9_1(.dout(w_dff_A_ecD7gx984_1),.din(w_dff_A_22JSAGlj9_1),.clk(gclk));
	jdff dff_A_6MWHxteX0_1(.dout(w_dff_A_22JSAGlj9_1),.din(w_dff_A_6MWHxteX0_1),.clk(gclk));
	jdff dff_A_CCd8nReW7_1(.dout(w_dff_A_6MWHxteX0_1),.din(w_dff_A_CCd8nReW7_1),.clk(gclk));
	jdff dff_A_bzIOoVfs3_1(.dout(w_dff_A_CCd8nReW7_1),.din(w_dff_A_bzIOoVfs3_1),.clk(gclk));
	jdff dff_A_8ibn2ThK1_1(.dout(w_dff_A_bzIOoVfs3_1),.din(w_dff_A_8ibn2ThK1_1),.clk(gclk));
	jdff dff_B_lUZDsqeU1_1(.din(n1392),.dout(w_dff_B_lUZDsqeU1_1),.clk(gclk));
	jdff dff_B_z42zrVKM5_1(.din(w_dff_B_lUZDsqeU1_1),.dout(w_dff_B_z42zrVKM5_1),.clk(gclk));
	jdff dff_B_QSnSHTIl6_1(.din(w_dff_B_z42zrVKM5_1),.dout(w_dff_B_QSnSHTIl6_1),.clk(gclk));
	jdff dff_B_EFsU1XA45_1(.din(w_dff_B_QSnSHTIl6_1),.dout(w_dff_B_EFsU1XA45_1),.clk(gclk));
	jdff dff_B_cKc2TOh76_1(.din(w_dff_B_EFsU1XA45_1),.dout(w_dff_B_cKc2TOh76_1),.clk(gclk));
	jdff dff_B_CQpW27lF9_1(.din(w_dff_B_cKc2TOh76_1),.dout(w_dff_B_CQpW27lF9_1),.clk(gclk));
	jdff dff_A_fgrJABZv7_1(.dout(w_n1447_0[1]),.din(w_dff_A_fgrJABZv7_1),.clk(gclk));
	jdff dff_B_YlSAaHFt4_1(.din(n1412),.dout(w_dff_B_YlSAaHFt4_1),.clk(gclk));
	jdff dff_B_F4g3du833_1(.din(w_dff_B_YlSAaHFt4_1),.dout(w_dff_B_F4g3du833_1),.clk(gclk));
	jdff dff_B_LBs5Rtdw0_1(.din(w_dff_B_F4g3du833_1),.dout(w_dff_B_LBs5Rtdw0_1),.clk(gclk));
	jdff dff_B_REGeQgUa0_1(.din(w_dff_B_LBs5Rtdw0_1),.dout(w_dff_B_REGeQgUa0_1),.clk(gclk));
	jdff dff_B_ZPyW40H24_1(.din(w_dff_B_REGeQgUa0_1),.dout(w_dff_B_ZPyW40H24_1),.clk(gclk));
	jdff dff_B_rfRIYaNb9_1(.din(w_dff_B_ZPyW40H24_1),.dout(w_dff_B_rfRIYaNb9_1),.clk(gclk));
	jdff dff_B_2aMxh9bk1_1(.din(w_dff_B_rfRIYaNb9_1),.dout(w_dff_B_2aMxh9bk1_1),.clk(gclk));
	jdff dff_B_0B84Cl4m5_1(.din(w_dff_B_2aMxh9bk1_1),.dout(w_dff_B_0B84Cl4m5_1),.clk(gclk));
	jdff dff_B_wBbD3bNt9_1(.din(w_dff_B_0B84Cl4m5_1),.dout(w_dff_B_wBbD3bNt9_1),.clk(gclk));
	jdff dff_B_d8pD8Ezv4_1(.din(w_dff_B_wBbD3bNt9_1),.dout(w_dff_B_d8pD8Ezv4_1),.clk(gclk));
	jdff dff_B_ANg88wro8_0(.din(n1443),.dout(w_dff_B_ANg88wro8_0),.clk(gclk));
	jdff dff_B_9GLwzPEr8_0(.din(n1440),.dout(w_dff_B_9GLwzPEr8_0),.clk(gclk));
	jdff dff_A_QtvilpXc4_1(.dout(w_n1438_0[1]),.din(w_dff_A_QtvilpXc4_1),.clk(gclk));
	jdff dff_A_uPM6mDAw0_1(.dout(w_dff_A_QtvilpXc4_1),.din(w_dff_A_uPM6mDAw0_1),.clk(gclk));
	jdff dff_A_KzB0g1Nb1_1(.dout(w_dff_A_uPM6mDAw0_1),.din(w_dff_A_KzB0g1Nb1_1),.clk(gclk));
	jdff dff_B_y9QNuL3z4_0(.din(n1437),.dout(w_dff_B_y9QNuL3z4_0),.clk(gclk));
	jdff dff_B_dFCMmpUR1_1(.din(n1427),.dout(w_dff_B_dFCMmpUR1_1),.clk(gclk));
	jdff dff_B_uHKiqOJY7_1(.din(n1428),.dout(w_dff_B_uHKiqOJY7_1),.clk(gclk));
	jdff dff_B_cUJPDF5T8_1(.din(w_dff_B_uHKiqOJY7_1),.dout(w_dff_B_cUJPDF5T8_1),.clk(gclk));
	jdff dff_B_76hbirnt5_1(.din(w_dff_B_cUJPDF5T8_1),.dout(w_dff_B_76hbirnt5_1),.clk(gclk));
	jdff dff_B_R5ODUbWW7_1(.din(w_dff_B_76hbirnt5_1),.dout(w_dff_B_R5ODUbWW7_1),.clk(gclk));
	jdff dff_B_JVbrCqGZ3_1(.din(w_dff_B_R5ODUbWW7_1),.dout(w_dff_B_JVbrCqGZ3_1),.clk(gclk));
	jdff dff_B_URvx2Jvn2_1(.din(w_dff_B_JVbrCqGZ3_1),.dout(w_dff_B_URvx2Jvn2_1),.clk(gclk));
	jdff dff_B_SIU56iQI0_1(.din(w_dff_B_URvx2Jvn2_1),.dout(w_dff_B_SIU56iQI0_1),.clk(gclk));
	jdff dff_B_BbDFpwmB6_1(.din(w_dff_B_SIU56iQI0_1),.dout(w_dff_B_BbDFpwmB6_1),.clk(gclk));
	jdff dff_B_7U2Armpn8_1(.din(w_dff_B_BbDFpwmB6_1),.dout(w_dff_B_7U2Armpn8_1),.clk(gclk));
	jdff dff_B_SQFxn9UY4_1(.din(w_dff_B_7U2Armpn8_1),.dout(w_dff_B_SQFxn9UY4_1),.clk(gclk));
	jdff dff_B_7J4yUeo43_1(.din(w_dff_B_SQFxn9UY4_1),.dout(w_dff_B_7J4yUeo43_1),.clk(gclk));
	jdff dff_B_CNapvRPK9_1(.din(n1414),.dout(w_dff_B_CNapvRPK9_1),.clk(gclk));
	jdff dff_B_9NzEBlA36_1(.din(w_dff_B_CNapvRPK9_1),.dout(w_dff_B_9NzEBlA36_1),.clk(gclk));
	jdff dff_B_ZqSJntMl5_1(.din(w_dff_B_9NzEBlA36_1),.dout(w_dff_B_ZqSJntMl5_1),.clk(gclk));
	jdff dff_B_vj4uRcAr3_1(.din(w_dff_B_ZqSJntMl5_1),.dout(w_dff_B_vj4uRcAr3_1),.clk(gclk));
	jdff dff_B_jPIh30mM3_1(.din(n1423),.dout(w_dff_B_jPIh30mM3_1),.clk(gclk));
	jdff dff_B_fXge62pK6_0(.din(n1422),.dout(w_dff_B_fXge62pK6_0),.clk(gclk));
	jdff dff_A_ChlsoDwO8_0(.dout(w_n1421_0[0]),.din(w_dff_A_ChlsoDwO8_0),.clk(gclk));
	jdff dff_A_0ay4vSmU3_0(.dout(w_dff_A_ChlsoDwO8_0),.din(w_dff_A_0ay4vSmU3_0),.clk(gclk));
	jdff dff_A_JXVu36Ka7_0(.dout(w_dff_A_0ay4vSmU3_0),.din(w_dff_A_JXVu36Ka7_0),.clk(gclk));
	jdff dff_B_AHQpbTXO6_1(.din(n1415),.dout(w_dff_B_AHQpbTXO6_1),.clk(gclk));
	jdff dff_A_C6FdzPPt8_1(.dout(w_n829_0[1]),.din(w_dff_A_C6FdzPPt8_1),.clk(gclk));
	jdff dff_A_w48cUdHX2_0(.dout(w_n614_1[0]),.din(w_dff_A_w48cUdHX2_0),.clk(gclk));
	jdff dff_A_EaANQjNV7_0(.dout(w_dff_A_w48cUdHX2_0),.din(w_dff_A_EaANQjNV7_0),.clk(gclk));
	jdff dff_A_aRyKXAax3_0(.dout(w_dff_A_EaANQjNV7_0),.din(w_dff_A_aRyKXAax3_0),.clk(gclk));
	jdff dff_A_TfB8AK0q8_0(.dout(w_dff_A_aRyKXAax3_0),.din(w_dff_A_TfB8AK0q8_0),.clk(gclk));
	jdff dff_A_pBW3DPRX8_0(.dout(w_dff_A_TfB8AK0q8_0),.din(w_dff_A_pBW3DPRX8_0),.clk(gclk));
	jdff dff_A_rxs2INgK8_2(.dout(w_n614_1[2]),.din(w_dff_A_rxs2INgK8_2),.clk(gclk));
	jdff dff_A_UQB2RqFo7_2(.dout(w_dff_A_rxs2INgK8_2),.din(w_dff_A_UQB2RqFo7_2),.clk(gclk));
	jdff dff_A_Tx2A3lWa6_2(.dout(w_dff_A_UQB2RqFo7_2),.din(w_dff_A_Tx2A3lWa6_2),.clk(gclk));
	jdff dff_A_J04wO39a1_2(.dout(w_dff_A_Tx2A3lWa6_2),.din(w_dff_A_J04wO39a1_2),.clk(gclk));
	jdff dff_A_H3wNa1iM6_2(.dout(w_dff_A_J04wO39a1_2),.din(w_dff_A_H3wNa1iM6_2),.clk(gclk));
	jdff dff_A_LOEMaROP6_2(.dout(w_dff_A_H3wNa1iM6_2),.din(w_dff_A_LOEMaROP6_2),.clk(gclk));
	jdff dff_A_QOi2xMeJ2_1(.dout(w_n828_0[1]),.din(w_dff_A_QOi2xMeJ2_1),.clk(gclk));
	jdff dff_A_cwgcIkMW2_1(.dout(w_dff_A_QOi2xMeJ2_1),.din(w_dff_A_cwgcIkMW2_1),.clk(gclk));
	jdff dff_A_EpDPndjc0_1(.dout(w_dff_A_cwgcIkMW2_1),.din(w_dff_A_EpDPndjc0_1),.clk(gclk));
	jdff dff_A_gO8VDvG40_1(.dout(w_dff_A_EpDPndjc0_1),.din(w_dff_A_gO8VDvG40_1),.clk(gclk));
	jdff dff_A_JP3Ip3nE2_1(.dout(w_dff_A_gO8VDvG40_1),.din(w_dff_A_JP3Ip3nE2_1),.clk(gclk));
	jdff dff_A_VnwMUdos2_1(.dout(w_dff_A_JP3Ip3nE2_1),.din(w_dff_A_VnwMUdos2_1),.clk(gclk));
	jdff dff_A_rwbuN3lF2_2(.dout(w_n828_0[2]),.din(w_dff_A_rwbuN3lF2_2),.clk(gclk));
	jdff dff_A_WutHriiW2_2(.dout(w_dff_A_rwbuN3lF2_2),.din(w_dff_A_WutHriiW2_2),.clk(gclk));
	jdff dff_B_xQFBRjFr0_2(.din(n787),.dout(w_dff_B_xQFBRjFr0_2),.clk(gclk));
	jdff dff_B_K3fr7C5p8_2(.din(w_dff_B_xQFBRjFr0_2),.dout(w_dff_B_K3fr7C5p8_2),.clk(gclk));
	jdff dff_B_NttktZYI2_2(.din(w_dff_B_K3fr7C5p8_2),.dout(w_dff_B_NttktZYI2_2),.clk(gclk));
	jdff dff_B_P4fo1Pmd8_2(.din(w_dff_B_NttktZYI2_2),.dout(w_dff_B_P4fo1Pmd8_2),.clk(gclk));
	jdff dff_B_BaqOPZ646_2(.din(w_dff_B_P4fo1Pmd8_2),.dout(w_dff_B_BaqOPZ646_2),.clk(gclk));
	jdff dff_B_S7yHHKqo3_2(.din(w_dff_B_BaqOPZ646_2),.dout(w_dff_B_S7yHHKqo3_2),.clk(gclk));
	jdff dff_B_HfrBjEFp6_2(.din(w_dff_B_S7yHHKqo3_2),.dout(w_dff_B_HfrBjEFp6_2),.clk(gclk));
	jdff dff_B_PJsAM0Am4_2(.din(w_dff_B_HfrBjEFp6_2),.dout(w_dff_B_PJsAM0Am4_2),.clk(gclk));
	jdff dff_B_tswFWHNN0_2(.din(w_dff_B_PJsAM0Am4_2),.dout(w_dff_B_tswFWHNN0_2),.clk(gclk));
	jdff dff_A_pdGcakNm7_1(.dout(w_n779_0[1]),.din(w_dff_A_pdGcakNm7_1),.clk(gclk));
	jdff dff_A_ffwLEjuB8_1(.dout(w_dff_A_pdGcakNm7_1),.din(w_dff_A_ffwLEjuB8_1),.clk(gclk));
	jdff dff_A_d3odaars2_1(.dout(w_dff_A_ffwLEjuB8_1),.din(w_dff_A_d3odaars2_1),.clk(gclk));
	jdff dff_A_esJnoely4_1(.dout(w_dff_A_d3odaars2_1),.din(w_dff_A_esJnoely4_1),.clk(gclk));
	jdff dff_A_HlIqDWum0_1(.dout(w_dff_A_esJnoely4_1),.din(w_dff_A_HlIqDWum0_1),.clk(gclk));
	jdff dff_A_hho9pabx0_1(.dout(w_dff_A_HlIqDWum0_1),.din(w_dff_A_hho9pabx0_1),.clk(gclk));
	jdff dff_A_wjyPR4Q55_1(.dout(w_dff_A_hho9pabx0_1),.din(w_dff_A_wjyPR4Q55_1),.clk(gclk));
	jdff dff_A_F0SmUnOV6_1(.dout(w_dff_A_wjyPR4Q55_1),.din(w_dff_A_F0SmUnOV6_1),.clk(gclk));
	jdff dff_A_Gghfwt0C2_1(.dout(w_dff_A_F0SmUnOV6_1),.din(w_dff_A_Gghfwt0C2_1),.clk(gclk));
	jdff dff_A_GfciHy3B3_1(.dout(w_dff_A_Gghfwt0C2_1),.din(w_dff_A_GfciHy3B3_1),.clk(gclk));
	jdff dff_A_LefhVn3Z6_1(.dout(w_dff_A_GfciHy3B3_1),.din(w_dff_A_LefhVn3Z6_1),.clk(gclk));
	jdff dff_A_WZyU70B86_1(.dout(w_dff_A_LefhVn3Z6_1),.din(w_dff_A_WZyU70B86_1),.clk(gclk));
	jdff dff_A_ySfB1G0n0_1(.dout(w_n636_1[1]),.din(w_dff_A_ySfB1G0n0_1),.clk(gclk));
	jdff dff_A_ADSSagpo0_1(.dout(w_dff_A_ySfB1G0n0_1),.din(w_dff_A_ADSSagpo0_1),.clk(gclk));
	jdff dff_A_K6f1eYEf2_2(.dout(w_n636_0[2]),.din(w_dff_A_K6f1eYEf2_2),.clk(gclk));
	jdff dff_A_BRclw7Kc3_0(.dout(w_n1411_0[0]),.din(w_dff_A_BRclw7Kc3_0),.clk(gclk));
	jdff dff_A_kiNFkwt71_0(.dout(w_dff_A_BRclw7Kc3_0),.din(w_dff_A_kiNFkwt71_0),.clk(gclk));
	jdff dff_A_jnlbi7kZ4_0(.dout(w_dff_A_kiNFkwt71_0),.din(w_dff_A_jnlbi7kZ4_0),.clk(gclk));
	jdff dff_A_Ru1gRn2Z3_0(.dout(w_dff_A_jnlbi7kZ4_0),.din(w_dff_A_Ru1gRn2Z3_0),.clk(gclk));
	jdff dff_A_jSszOj0K5_0(.dout(w_dff_A_Ru1gRn2Z3_0),.din(w_dff_A_jSszOj0K5_0),.clk(gclk));
	jdff dff_A_1HrCzaq51_0(.dout(w_dff_A_jSszOj0K5_0),.din(w_dff_A_1HrCzaq51_0),.clk(gclk));
	jdff dff_A_Kbxrl8Z16_0(.dout(w_dff_A_1HrCzaq51_0),.din(w_dff_A_Kbxrl8Z16_0),.clk(gclk));
	jdff dff_A_urhDNzTr3_0(.dout(w_dff_A_Kbxrl8Z16_0),.din(w_dff_A_urhDNzTr3_0),.clk(gclk));
	jdff dff_A_MMdQ1c6m6_0(.dout(w_dff_A_urhDNzTr3_0),.din(w_dff_A_MMdQ1c6m6_0),.clk(gclk));
	jdff dff_A_hIqyZcc48_0(.dout(w_dff_A_MMdQ1c6m6_0),.din(w_dff_A_hIqyZcc48_0),.clk(gclk));
	jdff dff_A_jIOBzIQ13_0(.dout(w_dff_A_hIqyZcc48_0),.din(w_dff_A_jIOBzIQ13_0),.clk(gclk));
	jdff dff_A_xyxMXKFh7_0(.dout(w_n1409_0[0]),.din(w_dff_A_xyxMXKFh7_0),.clk(gclk));
	jdff dff_B_AOf3PMd74_1(.din(n1405),.dout(w_dff_B_AOf3PMd74_1),.clk(gclk));
	jdff dff_B_RSBxnL4w9_0(.din(n1407),.dout(w_dff_B_RSBxnL4w9_0),.clk(gclk));
	jdff dff_B_fvTJbHeF9_0(.din(w_dff_B_RSBxnL4w9_0),.dout(w_dff_B_fvTJbHeF9_0),.clk(gclk));
	jdff dff_B_FcFEgFew3_0(.din(w_dff_B_fvTJbHeF9_0),.dout(w_dff_B_FcFEgFew3_0),.clk(gclk));
	jdff dff_B_9ODYf6pV6_0(.din(w_dff_B_FcFEgFew3_0),.dout(w_dff_B_9ODYf6pV6_0),.clk(gclk));
	jdff dff_A_aQ7HXJvB2_1(.dout(w_n968_0[1]),.din(w_dff_A_aQ7HXJvB2_1),.clk(gclk));
	jdff dff_A_MRlr7ald7_1(.dout(w_dff_A_aQ7HXJvB2_1),.din(w_dff_A_MRlr7ald7_1),.clk(gclk));
	jdff dff_A_J0qI5n7m6_1(.dout(w_dff_A_MRlr7ald7_1),.din(w_dff_A_J0qI5n7m6_1),.clk(gclk));
	jdff dff_A_ALpZQIjD5_1(.dout(w_dff_A_J0qI5n7m6_1),.din(w_dff_A_ALpZQIjD5_1),.clk(gclk));
	jdff dff_A_JjHPO06u2_1(.dout(w_dff_A_ALpZQIjD5_1),.din(w_dff_A_JjHPO06u2_1),.clk(gclk));
	jdff dff_B_6rqXqpJ01_2(.din(n968),.dout(w_dff_B_6rqXqpJ01_2),.clk(gclk));
	jdff dff_B_mwnP0hxW8_2(.din(w_dff_B_6rqXqpJ01_2),.dout(w_dff_B_mwnP0hxW8_2),.clk(gclk));
	jdff dff_B_KRKihJsA9_2(.din(w_dff_B_mwnP0hxW8_2),.dout(w_dff_B_KRKihJsA9_2),.clk(gclk));
	jdff dff_B_fGNxAou53_2(.din(w_dff_B_KRKihJsA9_2),.dout(w_dff_B_fGNxAou53_2),.clk(gclk));
	jdff dff_B_r2WXSA2G3_2(.din(w_dff_B_fGNxAou53_2),.dout(w_dff_B_r2WXSA2G3_2),.clk(gclk));
	jdff dff_B_x8jcFjAS6_0(.din(n1404),.dout(w_dff_B_x8jcFjAS6_0),.clk(gclk));
	jdff dff_B_fdXgcZAc6_0(.din(w_dff_B_x8jcFjAS6_0),.dout(w_dff_B_fdXgcZAc6_0),.clk(gclk));
	jdff dff_B_63HPZrNT6_1(.din(n1401),.dout(w_dff_B_63HPZrNT6_1),.clk(gclk));
	jdff dff_B_Qwk5WDrA8_1(.din(w_dff_B_63HPZrNT6_1),.dout(w_dff_B_Qwk5WDrA8_1),.clk(gclk));
	jdff dff_B_eM51dZqn7_1(.din(w_dff_B_Qwk5WDrA8_1),.dout(w_dff_B_eM51dZqn7_1),.clk(gclk));
	jdff dff_A_CmsnOfjB2_1(.dout(w_n651_0[1]),.din(w_dff_A_CmsnOfjB2_1),.clk(gclk));
	jdff dff_A_GOHXnMpZ8_1(.dout(w_dff_A_CmsnOfjB2_1),.din(w_dff_A_GOHXnMpZ8_1),.clk(gclk));
	jdff dff_A_QrUn5Y1q2_1(.dout(w_dff_A_GOHXnMpZ8_1),.din(w_dff_A_QrUn5Y1q2_1),.clk(gclk));
	jdff dff_A_CoR02alG1_2(.dout(w_n651_0[2]),.din(w_dff_A_CoR02alG1_2),.clk(gclk));
	jdff dff_A_oG4v0NJT1_2(.dout(w_dff_A_CoR02alG1_2),.din(w_dff_A_oG4v0NJT1_2),.clk(gclk));
	jdff dff_A_DF5FSiJD0_2(.dout(w_dff_A_oG4v0NJT1_2),.din(w_dff_A_DF5FSiJD0_2),.clk(gclk));
	jdff dff_A_rJR5CfaT1_2(.dout(w_dff_A_DF5FSiJD0_2),.din(w_dff_A_rJR5CfaT1_2),.clk(gclk));
	jdff dff_A_yikJDtD03_2(.dout(w_dff_A_rJR5CfaT1_2),.din(w_dff_A_yikJDtD03_2),.clk(gclk));
	jdff dff_A_Xkr6dqbD7_2(.dout(w_dff_A_yikJDtD03_2),.din(w_dff_A_Xkr6dqbD7_2),.clk(gclk));
	jdff dff_A_SSqurgJA3_2(.dout(w_dff_A_Xkr6dqbD7_2),.din(w_dff_A_SSqurgJA3_2),.clk(gclk));
	jdff dff_B_5tBr8GmK5_3(.din(n651),.dout(w_dff_B_5tBr8GmK5_3),.clk(gclk));
	jdff dff_A_466xwsJd9_0(.dout(w_n650_0[0]),.din(w_dff_A_466xwsJd9_0),.clk(gclk));
	jdff dff_A_3SyX6WOy6_0(.dout(w_dff_A_466xwsJd9_0),.din(w_dff_A_3SyX6WOy6_0),.clk(gclk));
	jdff dff_A_9ecManOQ7_0(.dout(w_dff_A_3SyX6WOy6_0),.din(w_dff_A_9ecManOQ7_0),.clk(gclk));
	jdff dff_A_L64PkMmi3_0(.dout(w_dff_A_9ecManOQ7_0),.din(w_dff_A_L64PkMmi3_0),.clk(gclk));
	jdff dff_A_9VMwjoTv1_0(.dout(w_dff_A_L64PkMmi3_0),.din(w_dff_A_9VMwjoTv1_0),.clk(gclk));
	jdff dff_A_eKYXsKcW3_0(.dout(w_dff_A_9VMwjoTv1_0),.din(w_dff_A_eKYXsKcW3_0),.clk(gclk));
	jdff dff_A_pDDuEHYq6_0(.dout(w_dff_A_eKYXsKcW3_0),.din(w_dff_A_pDDuEHYq6_0),.clk(gclk));
	jdff dff_A_38imH19D1_0(.dout(w_dff_A_pDDuEHYq6_0),.din(w_dff_A_38imH19D1_0),.clk(gclk));
	jdff dff_A_g83TBW6C0_0(.dout(w_dff_A_38imH19D1_0),.din(w_dff_A_g83TBW6C0_0),.clk(gclk));
	jdff dff_B_GtX4MKB26_1(.din(n1395),.dout(w_dff_B_GtX4MKB26_1),.clk(gclk));
	jdff dff_A_IA24yFJu7_1(.dout(w_n740_0[1]),.din(w_dff_A_IA24yFJu7_1),.clk(gclk));
	jdff dff_A_BkPpqbEr6_0(.dout(w_n739_1[0]),.din(w_dff_A_BkPpqbEr6_0),.clk(gclk));
	jdff dff_A_MQUS6LhM8_0(.dout(w_dff_A_BkPpqbEr6_0),.din(w_dff_A_MQUS6LhM8_0),.clk(gclk));
	jdff dff_A_OsDmPOrR7_0(.dout(w_dff_A_MQUS6LhM8_0),.din(w_dff_A_OsDmPOrR7_0),.clk(gclk));
	jdff dff_A_bqXPRDbF7_0(.dout(w_dff_A_OsDmPOrR7_0),.din(w_dff_A_bqXPRDbF7_0),.clk(gclk));
	jdff dff_A_AhheJNR09_0(.dout(w_dff_A_bqXPRDbF7_0),.din(w_dff_A_AhheJNR09_0),.clk(gclk));
	jdff dff_A_O7xdiAw80_0(.dout(w_dff_A_AhheJNR09_0),.din(w_dff_A_O7xdiAw80_0),.clk(gclk));
	jdff dff_A_ROPVd4b70_0(.dout(w_dff_A_O7xdiAw80_0),.din(w_dff_A_ROPVd4b70_0),.clk(gclk));
	jdff dff_A_NABcI0GJ6_0(.dout(w_dff_A_ROPVd4b70_0),.din(w_dff_A_NABcI0GJ6_0),.clk(gclk));
	jdff dff_A_mpgmD9Kb4_0(.dout(w_dff_A_NABcI0GJ6_0),.din(w_dff_A_mpgmD9Kb4_0),.clk(gclk));
	jdff dff_A_dkW0DJwa4_2(.dout(w_n739_0[2]),.din(w_dff_A_dkW0DJwa4_2),.clk(gclk));
	jdff dff_A_mkBWdZtU7_2(.dout(w_dff_A_dkW0DJwa4_2),.din(w_dff_A_mkBWdZtU7_2),.clk(gclk));
	jdff dff_A_zLgKIio29_2(.dout(w_dff_A_mkBWdZtU7_2),.din(w_dff_A_zLgKIio29_2),.clk(gclk));
	jdff dff_A_rIWb77up4_2(.dout(w_dff_A_zLgKIio29_2),.din(w_dff_A_rIWb77up4_2),.clk(gclk));
	jdff dff_A_edJapZXS5_2(.dout(w_dff_A_rIWb77up4_2),.din(w_dff_A_edJapZXS5_2),.clk(gclk));
	jdff dff_A_4o8dWzod0_2(.dout(w_n649_0[2]),.din(w_dff_A_4o8dWzod0_2),.clk(gclk));
	jdff dff_B_HkACRLua4_0(.din(n648),.dout(w_dff_B_HkACRLua4_0),.clk(gclk));
	jdff dff_B_EbanuIL94_1(.din(G323),.dout(w_dff_B_EbanuIL94_1),.clk(gclk));
	jdff dff_A_gIfxbOeB2_0(.dout(w_n640_1[0]),.din(w_dff_A_gIfxbOeB2_0),.clk(gclk));
	jdff dff_A_W8bNgbnM3_0(.dout(w_dff_A_gIfxbOeB2_0),.din(w_dff_A_W8bNgbnM3_0),.clk(gclk));
	jdff dff_A_KMn58kOm9_0(.dout(w_dff_A_W8bNgbnM3_0),.din(w_dff_A_KMn58kOm9_0),.clk(gclk));
	jdff dff_A_j9Cq96bD8_0(.dout(w_dff_A_KMn58kOm9_0),.din(w_dff_A_j9Cq96bD8_0),.clk(gclk));
	jdff dff_A_lXQfBWHf5_0(.dout(w_dff_A_j9Cq96bD8_0),.din(w_dff_A_lXQfBWHf5_0),.clk(gclk));
	jdff dff_A_Mrsvtuqe3_0(.dout(w_dff_A_lXQfBWHf5_0),.din(w_dff_A_Mrsvtuqe3_0),.clk(gclk));
	jdff dff_A_adanFM526_0(.dout(w_dff_A_Mrsvtuqe3_0),.din(w_dff_A_adanFM526_0),.clk(gclk));
	jdff dff_A_o3SGJcYE7_0(.dout(w_dff_A_adanFM526_0),.din(w_dff_A_o3SGJcYE7_0),.clk(gclk));
	jdff dff_A_3gixdF4m1_0(.dout(w_dff_A_o3SGJcYE7_0),.din(w_dff_A_3gixdF4m1_0),.clk(gclk));
	jdff dff_A_2UKq2RSX8_0(.dout(w_dff_A_3gixdF4m1_0),.din(w_dff_A_2UKq2RSX8_0),.clk(gclk));
	jdff dff_A_4qExMfTp2_0(.dout(w_dff_A_2UKq2RSX8_0),.din(w_dff_A_4qExMfTp2_0),.clk(gclk));
	jdff dff_A_5SPZsnnS9_0(.dout(w_n646_0[0]),.din(w_dff_A_5SPZsnnS9_0),.clk(gclk));
	jdff dff_A_XMc8XPuB1_0(.dout(w_dff_A_5SPZsnnS9_0),.din(w_dff_A_XMc8XPuB1_0),.clk(gclk));
	jdff dff_B_aa12GdHb2_0(.din(n644),.dout(w_dff_B_aa12GdHb2_0),.clk(gclk));
	jdff dff_B_lFMH0nP49_1(.din(G315),.dout(w_dff_B_lFMH0nP49_1),.clk(gclk));
	jdff dff_A_wCzkzTI42_1(.dout(w_n640_0[1]),.din(w_dff_A_wCzkzTI42_1),.clk(gclk));
	jdff dff_A_kMCd1Vpa5_2(.dout(w_n640_0[2]),.din(w_dff_A_kMCd1Vpa5_2),.clk(gclk));
	jdff dff_A_sXGtEOkU8_2(.dout(w_dff_A_kMCd1Vpa5_2),.din(w_dff_A_sXGtEOkU8_2),.clk(gclk));
	jdff dff_A_K8bEREo46_2(.dout(w_dff_A_sXGtEOkU8_2),.din(w_dff_A_K8bEREo46_2),.clk(gclk));
	jdff dff_A_OjVjRNuA3_2(.dout(w_dff_A_K8bEREo46_2),.din(w_dff_A_OjVjRNuA3_2),.clk(gclk));
	jdff dff_A_zlIap0zn3_2(.dout(w_dff_A_OjVjRNuA3_2),.din(w_dff_A_zlIap0zn3_2),.clk(gclk));
	jdff dff_A_FEP2jJOW5_2(.dout(w_dff_A_zlIap0zn3_2),.din(w_dff_A_FEP2jJOW5_2),.clk(gclk));
	jdff dff_A_3BiEFrMv1_2(.dout(w_dff_A_FEP2jJOW5_2),.din(w_dff_A_3BiEFrMv1_2),.clk(gclk));
	jdff dff_A_Uet3vZWn5_2(.dout(w_dff_A_3BiEFrMv1_2),.din(w_dff_A_Uet3vZWn5_2),.clk(gclk));
	jdff dff_A_8dmrSXMb2_2(.dout(w_dff_A_Uet3vZWn5_2),.din(w_dff_A_8dmrSXMb2_2),.clk(gclk));
	jdff dff_A_j7FfwYML2_2(.dout(w_dff_A_8dmrSXMb2_2),.din(w_dff_A_j7FfwYML2_2),.clk(gclk));
	jdff dff_A_SZza9EIx1_2(.dout(w_dff_A_j7FfwYML2_2),.din(w_dff_A_SZza9EIx1_2),.clk(gclk));
	jdff dff_B_8Vk4FzSE9_1(.din(n637),.dout(w_dff_B_8Vk4FzSE9_1),.clk(gclk));
	jdff dff_B_BVkNQ79x1_1(.din(G307),.dout(w_dff_B_BVkNQ79x1_1),.clk(gclk));
	jdff dff_B_1uHcbsMd7_0(.din(n1393),.dout(w_dff_B_1uHcbsMd7_0),.clk(gclk));
	jdff dff_B_TNEGyBiS4_0(.din(w_dff_B_1uHcbsMd7_0),.dout(w_dff_B_TNEGyBiS4_0),.clk(gclk));
	jdff dff_B_l1uAx0AP2_0(.din(w_dff_B_TNEGyBiS4_0),.dout(w_dff_B_l1uAx0AP2_0),.clk(gclk));
	jdff dff_A_TVYzYBxD9_0(.dout(w_n631_0[0]),.din(w_dff_A_TVYzYBxD9_0),.clk(gclk));
	jdff dff_A_MRAMZT0G8_0(.dout(w_dff_A_TVYzYBxD9_0),.din(w_dff_A_MRAMZT0G8_0),.clk(gclk));
	jdff dff_A_SNSIvQLJ8_0(.dout(w_dff_A_MRAMZT0G8_0),.din(w_dff_A_SNSIvQLJ8_0),.clk(gclk));
	jdff dff_A_71H4QDix5_1(.dout(w_n629_0[1]),.din(w_dff_A_71H4QDix5_1),.clk(gclk));
	jdff dff_A_A1l2JSGf8_1(.dout(w_dff_A_71H4QDix5_1),.din(w_dff_A_A1l2JSGf8_1),.clk(gclk));
	jdff dff_A_bAIxOVC57_1(.dout(w_dff_A_A1l2JSGf8_1),.din(w_dff_A_bAIxOVC57_1),.clk(gclk));
	jdff dff_A_ieu9LqiI2_1(.dout(w_n628_0[1]),.din(w_dff_A_ieu9LqiI2_1),.clk(gclk));
	jdff dff_B_sRRrq9fT4_0(.din(n627),.dout(w_dff_B_sRRrq9fT4_0),.clk(gclk));
	jdff dff_A_h4DbwCpQ5_0(.dout(w_n625_0[0]),.din(w_dff_A_h4DbwCpQ5_0),.clk(gclk));
	jdff dff_A_TV5Z6BNA5_2(.dout(w_n625_0[2]),.din(w_dff_A_TV5Z6BNA5_2),.clk(gclk));
	jdff dff_A_P6llDIia8_0(.dout(w_n623_0[0]),.din(w_dff_A_P6llDIia8_0),.clk(gclk));
	jdff dff_B_ow5BU3l15_0(.din(n616),.dout(w_dff_B_ow5BU3l15_0),.clk(gclk));
	jdff dff_A_rN5QuUBu0_0(.dout(w_G2174_0[0]),.din(w_dff_A_rN5QuUBu0_0),.clk(gclk));
	jdff dff_A_xnDHd5k14_0(.dout(w_dff_A_rN5QuUBu0_0),.din(w_dff_A_xnDHd5k14_0),.clk(gclk));
	jdff dff_A_U47ZbNnc1_0(.dout(w_dff_A_xnDHd5k14_0),.din(w_dff_A_U47ZbNnc1_0),.clk(gclk));
	jdff dff_A_VY8skPAt1_0(.dout(w_dff_A_U47ZbNnc1_0),.din(w_dff_A_VY8skPAt1_0),.clk(gclk));
	jdff dff_A_0yb5aQ5q4_0(.dout(w_dff_A_VY8skPAt1_0),.din(w_dff_A_0yb5aQ5q4_0),.clk(gclk));
	jdff dff_A_B9B5aRkE4_0(.dout(w_dff_A_0yb5aQ5q4_0),.din(w_dff_A_B9B5aRkE4_0),.clk(gclk));
	jdff dff_A_5wChciOM6_0(.dout(w_dff_A_B9B5aRkE4_0),.din(w_dff_A_5wChciOM6_0),.clk(gclk));
	jdff dff_A_ej0PMbLP8_0(.dout(w_dff_A_5wChciOM6_0),.din(w_dff_A_ej0PMbLP8_0),.clk(gclk));
	jdff dff_A_AYdZ9OPD3_0(.dout(w_dff_A_ej0PMbLP8_0),.din(w_dff_A_AYdZ9OPD3_0),.clk(gclk));
	jdff dff_A_DoYuYt3o0_0(.dout(w_dff_A_AYdZ9OPD3_0),.din(w_dff_A_DoYuYt3o0_0),.clk(gclk));
	jdff dff_A_FzmSQcjZ8_0(.dout(w_dff_A_DoYuYt3o0_0),.din(w_dff_A_FzmSQcjZ8_0),.clk(gclk));
	jdff dff_A_YFG3IsSo3_2(.dout(w_G2174_0[2]),.din(w_dff_A_YFG3IsSo3_2),.clk(gclk));
	jdff dff_A_eUw2U2AD1_2(.dout(w_dff_A_YFG3IsSo3_2),.din(w_dff_A_eUw2U2AD1_2),.clk(gclk));
	jdff dff_A_DNcLtVZT6_2(.dout(w_dff_A_eUw2U2AD1_2),.din(w_dff_A_DNcLtVZT6_2),.clk(gclk));
	jdff dff_A_DrSCtFhK1_2(.dout(w_dff_A_DNcLtVZT6_2),.din(w_dff_A_DrSCtFhK1_2),.clk(gclk));
	jdff dff_A_A3LqPYKu4_2(.dout(w_dff_A_DrSCtFhK1_2),.din(w_dff_A_A3LqPYKu4_2),.clk(gclk));
	jdff dff_A_3DUO5WVG8_2(.dout(w_dff_A_A3LqPYKu4_2),.din(w_dff_A_3DUO5WVG8_2),.clk(gclk));
	jdff dff_A_cChJUGIa0_2(.dout(w_dff_A_3DUO5WVG8_2),.din(w_dff_A_cChJUGIa0_2),.clk(gclk));
	jdff dff_A_TBhpKZhG1_2(.dout(w_dff_A_cChJUGIa0_2),.din(w_dff_A_TBhpKZhG1_2),.clk(gclk));
	jdff dff_B_Utw847178_1(.din(n711),.dout(w_dff_B_Utw847178_1),.clk(gclk));
	jdff dff_B_fIkYYlr24_1(.din(w_dff_B_Utw847178_1),.dout(w_dff_B_fIkYYlr24_1),.clk(gclk));
	jdff dff_B_q9lg12EA5_1(.din(w_dff_B_fIkYYlr24_1),.dout(w_dff_B_q9lg12EA5_1),.clk(gclk));
	jdff dff_B_gV0ujE1p6_1(.din(w_dff_B_q9lg12EA5_1),.dout(w_dff_B_gV0ujE1p6_1),.clk(gclk));
	jdff dff_B_3ZUXkE3q4_1(.din(w_dff_B_gV0ujE1p6_1),.dout(w_dff_B_3ZUXkE3q4_1),.clk(gclk));
	jdff dff_B_qOGmSgWp9_1(.din(w_dff_B_3ZUXkE3q4_1),.dout(w_dff_B_qOGmSgWp9_1),.clk(gclk));
	jdff dff_B_cNPK8Tiq9_1(.din(n712),.dout(w_dff_B_cNPK8Tiq9_1),.clk(gclk));
	jdff dff_B_0R7JY9iW9_1(.din(w_dff_B_cNPK8Tiq9_1),.dout(w_dff_B_0R7JY9iW9_1),.clk(gclk));
	jdff dff_B_efuL0FT03_1(.din(w_dff_B_0R7JY9iW9_1),.dout(w_dff_B_efuL0FT03_1),.clk(gclk));
	jdff dff_B_dt5rETtL5_1(.din(w_dff_B_efuL0FT03_1),.dout(w_dff_B_dt5rETtL5_1),.clk(gclk));
	jdff dff_B_B3RK3ujN2_1(.din(w_dff_B_dt5rETtL5_1),.dout(w_dff_B_B3RK3ujN2_1),.clk(gclk));
	jdff dff_B_mNPRY81a1_1(.din(n713),.dout(w_dff_B_mNPRY81a1_1),.clk(gclk));
	jdff dff_B_xkh3ej2l3_1(.din(w_dff_B_mNPRY81a1_1),.dout(w_dff_B_xkh3ej2l3_1),.clk(gclk));
	jdff dff_B_354K2EW42_1(.din(w_dff_B_xkh3ej2l3_1),.dout(w_dff_B_354K2EW42_1),.clk(gclk));
	jdff dff_B_xTDbuQrc6_1(.din(w_dff_B_354K2EW42_1),.dout(w_dff_B_xTDbuQrc6_1),.clk(gclk));
	jdff dff_A_fMv0x7dt0_0(.dout(w_n723_0[0]),.din(w_dff_A_fMv0x7dt0_0),.clk(gclk));
	jdff dff_A_KGO1f1I56_0(.dout(w_n621_2[0]),.din(w_dff_A_KGO1f1I56_0),.clk(gclk));
	jdff dff_A_s9lrbxa57_1(.dout(w_n721_0[1]),.din(w_dff_A_s9lrbxa57_1),.clk(gclk));
	jdff dff_A_rNSxHSxU8_1(.dout(w_dff_A_s9lrbxa57_1),.din(w_dff_A_rNSxHSxU8_1),.clk(gclk));
	jdff dff_A_p56n7AdR3_1(.dout(w_dff_A_rNSxHSxU8_1),.din(w_dff_A_p56n7AdR3_1),.clk(gclk));
	jdff dff_A_bbNVnxrp4_1(.dout(w_dff_A_p56n7AdR3_1),.din(w_dff_A_bbNVnxrp4_1),.clk(gclk));
	jdff dff_A_enNF7sed7_1(.dout(w_dff_A_bbNVnxrp4_1),.din(w_dff_A_enNF7sed7_1),.clk(gclk));
	jdff dff_A_IYre53nc7_1(.dout(w_dff_A_enNF7sed7_1),.din(w_dff_A_IYre53nc7_1),.clk(gclk));
	jdff dff_A_FYFbEOeg7_0(.dout(w_G358_0[0]),.din(w_dff_A_FYFbEOeg7_0),.clk(gclk));
	jdff dff_A_AT1Avun83_0(.dout(w_n388_1[0]),.din(w_dff_A_AT1Avun83_0),.clk(gclk));
	jdff dff_A_umPSBfAm7_1(.dout(w_n388_1[1]),.din(w_dff_A_umPSBfAm7_1),.clk(gclk));
	jdff dff_A_eUL5RS502_1(.dout(w_n717_0[1]),.din(w_dff_A_eUL5RS502_1),.clk(gclk));
	jdff dff_A_S2LToxqY5_1(.dout(w_dff_A_eUL5RS502_1),.din(w_dff_A_S2LToxqY5_1),.clk(gclk));
	jdff dff_A_d3P4bKgJ3_1(.dout(w_dff_A_S2LToxqY5_1),.din(w_dff_A_d3P4bKgJ3_1),.clk(gclk));
	jdff dff_A_VbcRc7wU1_2(.dout(w_n717_0[2]),.din(w_dff_A_VbcRc7wU1_2),.clk(gclk));
	jdff dff_A_YVKjARmo8_2(.dout(w_dff_A_VbcRc7wU1_2),.din(w_dff_A_YVKjARmo8_2),.clk(gclk));
	jdff dff_A_5N4U0R7P9_0(.dout(w_G348_0[0]),.din(w_dff_A_5N4U0R7P9_0),.clk(gclk));
	jdff dff_A_22LW2eOR1_0(.dout(w_G332_2[0]),.din(w_dff_A_22LW2eOR1_0),.clk(gclk));
	jdff dff_A_YUvWpXW59_0(.dout(w_n437_1[0]),.din(w_dff_A_YUvWpXW59_0),.clk(gclk));
	jdff dff_A_zQPB9WuL5_1(.dout(w_n437_1[1]),.din(w_dff_A_zQPB9WuL5_1),.clk(gclk));
	jdff dff_A_jbpgR47I0_0(.dout(w_G332_3[0]),.din(w_dff_A_jbpgR47I0_0),.clk(gclk));
	jdff dff_A_6hgNxPZ11_2(.dout(w_G332_3[2]),.din(w_dff_A_6hgNxPZ11_2),.clk(gclk));
	jdff dff_A_15kIWfyz3_0(.dout(w_n410_1[0]),.din(w_dff_A_15kIWfyz3_0),.clk(gclk));
	jdff dff_A_CyVrelK90_0(.dout(w_n614_2[0]),.din(w_dff_A_CyVrelK90_0),.clk(gclk));
	jdff dff_A_PexqyRIy5_0(.dout(w_dff_A_CyVrelK90_0),.din(w_dff_A_PexqyRIy5_0),.clk(gclk));
	jdff dff_A_pyxSFSNG2_0(.dout(w_dff_A_PexqyRIy5_0),.din(w_dff_A_pyxSFSNG2_0),.clk(gclk));
	jdff dff_A_HwhzBRUb9_1(.dout(w_n614_0[1]),.din(w_dff_A_HwhzBRUb9_1),.clk(gclk));
	jdff dff_A_uWtMHdEi7_1(.dout(w_dff_A_HwhzBRUb9_1),.din(w_dff_A_uWtMHdEi7_1),.clk(gclk));
	jdff dff_A_dFHUU87T3_2(.dout(w_n614_0[2]),.din(w_dff_A_dFHUU87T3_2),.clk(gclk));
	jdff dff_A_oIBi9uCt9_2(.dout(w_dff_A_dFHUU87T3_2),.din(w_dff_A_oIBi9uCt9_2),.clk(gclk));
	jdff dff_A_OpERxBMY3_2(.dout(w_dff_A_oIBi9uCt9_2),.din(w_dff_A_OpERxBMY3_2),.clk(gclk));
	jdff dff_A_dv9qDyKm0_2(.dout(w_dff_A_OpERxBMY3_2),.din(w_dff_A_dv9qDyKm0_2),.clk(gclk));
	jdff dff_B_2GSH3u6a3_1(.din(n610),.dout(w_dff_B_2GSH3u6a3_1),.clk(gclk));
	jdff dff_A_wdTD53Z07_0(.dout(w_G332_4[0]),.din(w_dff_A_wdTD53Z07_0),.clk(gclk));
	jdff dff_A_iJNkOBcs6_2(.dout(w_G332_1[2]),.din(w_dff_A_iJNkOBcs6_2),.clk(gclk));
	jdff dff_A_Q2Ystg7B1_1(.dout(w_G331_0[1]),.din(w_dff_A_Q2Ystg7B1_1),.clk(gclk));
	jdff dff_A_9zo8w2nC0_0(.dout(w_n1391_0[0]),.din(w_dff_A_9zo8w2nC0_0),.clk(gclk));
	jdff dff_A_2OpYfxyO8_0(.dout(w_dff_A_9zo8w2nC0_0),.din(w_dff_A_2OpYfxyO8_0),.clk(gclk));
	jdff dff_A_grOdrvAe0_0(.dout(w_dff_A_2OpYfxyO8_0),.din(w_dff_A_grOdrvAe0_0),.clk(gclk));
	jdff dff_A_gseW7AfT9_0(.dout(w_dff_A_grOdrvAe0_0),.din(w_dff_A_gseW7AfT9_0),.clk(gclk));
	jdff dff_A_PsI6B1CX7_0(.dout(w_dff_A_gseW7AfT9_0),.din(w_dff_A_PsI6B1CX7_0),.clk(gclk));
	jdff dff_A_gJrDnbTx0_0(.dout(w_dff_A_PsI6B1CX7_0),.din(w_dff_A_gJrDnbTx0_0),.clk(gclk));
	jdff dff_A_HBen2u2L4_0(.dout(w_dff_A_gJrDnbTx0_0),.din(w_dff_A_HBen2u2L4_0),.clk(gclk));
	jdff dff_B_JemMZoOb4_1(.din(n1389),.dout(w_dff_B_JemMZoOb4_1),.clk(gclk));
	jdff dff_B_l1aSVjxa3_1(.din(w_dff_B_JemMZoOb4_1),.dout(w_dff_B_l1aSVjxa3_1),.clk(gclk));
	jdff dff_A_229310Pj4_1(.dout(w_G4091_1[1]),.din(w_dff_A_229310Pj4_1),.clk(gclk));
	jdff dff_A_nEKMBtUX7_1(.dout(w_dff_A_229310Pj4_1),.din(w_dff_A_nEKMBtUX7_1),.clk(gclk));
	jdff dff_A_7pO45wdU2_1(.dout(w_dff_A_nEKMBtUX7_1),.din(w_dff_A_7pO45wdU2_1),.clk(gclk));
	jdff dff_A_fEPYXVYS3_1(.dout(w_dff_A_7pO45wdU2_1),.din(w_dff_A_fEPYXVYS3_1),.clk(gclk));
	jdff dff_A_XeoILYub2_1(.dout(w_dff_A_fEPYXVYS3_1),.din(w_dff_A_XeoILYub2_1),.clk(gclk));
	jdff dff_A_wDvfa1v54_1(.dout(w_dff_A_XeoILYub2_1),.din(w_dff_A_wDvfa1v54_1),.clk(gclk));
	jdff dff_A_Ps483HaZ6_1(.dout(w_dff_A_wDvfa1v54_1),.din(w_dff_A_Ps483HaZ6_1),.clk(gclk));
	jdff dff_A_viYBww8f6_1(.dout(w_dff_A_Ps483HaZ6_1),.din(w_dff_A_viYBww8f6_1),.clk(gclk));
	jdff dff_A_LuXkb1gQ3_1(.dout(w_dff_A_viYBww8f6_1),.din(w_dff_A_LuXkb1gQ3_1),.clk(gclk));
	jdff dff_A_c55wTJCO0_1(.dout(w_dff_A_LuXkb1gQ3_1),.din(w_dff_A_c55wTJCO0_1),.clk(gclk));
	jdff dff_A_lxZmYScW6_1(.dout(w_dff_A_c55wTJCO0_1),.din(w_dff_A_lxZmYScW6_1),.clk(gclk));
	jdff dff_A_H20UwY2C7_1(.dout(w_dff_A_lxZmYScW6_1),.din(w_dff_A_H20UwY2C7_1),.clk(gclk));
	jdff dff_A_v533jOmM9_1(.dout(w_dff_A_H20UwY2C7_1),.din(w_dff_A_v533jOmM9_1),.clk(gclk));
	jdff dff_A_W9shQgB82_1(.dout(w_dff_A_v533jOmM9_1),.din(w_dff_A_W9shQgB82_1),.clk(gclk));
	jdff dff_A_j6tD9JNz9_1(.dout(w_dff_A_W9shQgB82_1),.din(w_dff_A_j6tD9JNz9_1),.clk(gclk));
	jdff dff_A_YoCgkczG0_1(.dout(w_dff_A_j6tD9JNz9_1),.din(w_dff_A_YoCgkczG0_1),.clk(gclk));
	jdff dff_A_p4dN46MK3_1(.dout(w_dff_A_YoCgkczG0_1),.din(w_dff_A_p4dN46MK3_1),.clk(gclk));
	jdff dff_A_GBdJ8qxM0_1(.dout(w_dff_A_p4dN46MK3_1),.din(w_dff_A_GBdJ8qxM0_1),.clk(gclk));
	jdff dff_A_eI23THGf9_2(.dout(w_G4091_1[2]),.din(w_dff_A_eI23THGf9_2),.clk(gclk));
	jdff dff_A_gVNAxhYM2_2(.dout(w_dff_A_eI23THGf9_2),.din(w_dff_A_gVNAxhYM2_2),.clk(gclk));
	jdff dff_A_XYLxVUDh7_2(.dout(w_dff_A_gVNAxhYM2_2),.din(w_dff_A_XYLxVUDh7_2),.clk(gclk));
	jdff dff_A_drA0dc717_2(.dout(w_dff_A_XYLxVUDh7_2),.din(w_dff_A_drA0dc717_2),.clk(gclk));
	jdff dff_A_2GxEKn7v5_2(.dout(w_dff_A_drA0dc717_2),.din(w_dff_A_2GxEKn7v5_2),.clk(gclk));
	jdff dff_A_tlY3woxf6_2(.dout(w_dff_A_2GxEKn7v5_2),.din(w_dff_A_tlY3woxf6_2),.clk(gclk));
	jdff dff_A_zOM3h7rE3_2(.dout(w_dff_A_tlY3woxf6_2),.din(w_dff_A_zOM3h7rE3_2),.clk(gclk));
	jdff dff_A_KMxa9F4G3_2(.dout(w_dff_A_zOM3h7rE3_2),.din(w_dff_A_KMxa9F4G3_2),.clk(gclk));
	jdff dff_A_8ld0AhPF6_2(.dout(w_dff_A_KMxa9F4G3_2),.din(w_dff_A_8ld0AhPF6_2),.clk(gclk));
	jdff dff_A_U2nEUDmM9_2(.dout(w_dff_A_8ld0AhPF6_2),.din(w_dff_A_U2nEUDmM9_2),.clk(gclk));
	jdff dff_A_hcffjs9U1_0(.dout(w_n1383_0[0]),.din(w_dff_A_hcffjs9U1_0),.clk(gclk));
	jdff dff_A_ZDq3w5ma4_0(.dout(w_dff_A_hcffjs9U1_0),.din(w_dff_A_ZDq3w5ma4_0),.clk(gclk));
	jdff dff_B_7Zrzttfu0_1(.din(n1363),.dout(w_dff_B_7Zrzttfu0_1),.clk(gclk));
	jdff dff_B_hfwAfqic5_1(.din(w_dff_B_7Zrzttfu0_1),.dout(w_dff_B_hfwAfqic5_1),.clk(gclk));
	jdff dff_B_aN7DnGVD7_1(.din(n1376),.dout(w_dff_B_aN7DnGVD7_1),.clk(gclk));
	jdff dff_B_MNXlIaF17_1(.din(n1377),.dout(w_dff_B_MNXlIaF17_1),.clk(gclk));
	jdff dff_A_Fn8Bdpbb4_1(.dout(w_n426_0[1]),.din(w_dff_A_Fn8Bdpbb4_1),.clk(gclk));
	jdff dff_A_k31sob227_0(.dout(w_G503_1[0]),.din(w_dff_A_k31sob227_0),.clk(gclk));
	jdff dff_A_JKwks8bX3_0(.dout(w_dff_A_k31sob227_0),.din(w_dff_A_JKwks8bX3_0),.clk(gclk));
	jdff dff_A_86MfvnTh9_0(.dout(w_dff_A_JKwks8bX3_0),.din(w_dff_A_86MfvnTh9_0),.clk(gclk));
	jdff dff_A_Zlou7Hha4_0(.dout(w_dff_A_86MfvnTh9_0),.din(w_dff_A_Zlou7Hha4_0),.clk(gclk));
	jdff dff_A_0SmFqPbu6_1(.dout(w_G503_1[1]),.din(w_dff_A_0SmFqPbu6_1),.clk(gclk));
	jdff dff_A_wBrNA6kY6_1(.dout(w_G503_0[1]),.din(w_dff_A_wBrNA6kY6_1),.clk(gclk));
	jdff dff_A_vgOyOihe1_1(.dout(w_dff_A_wBrNA6kY6_1),.din(w_dff_A_vgOyOihe1_1),.clk(gclk));
	jdff dff_A_lS6kLNkC3_2(.dout(w_G503_0[2]),.din(w_dff_A_lS6kLNkC3_2),.clk(gclk));
	jdff dff_A_ABaQaqS04_2(.dout(w_dff_A_lS6kLNkC3_2),.din(w_dff_A_ABaQaqS04_2),.clk(gclk));
	jdff dff_A_F5NgWOo37_2(.dout(w_dff_A_ABaQaqS04_2),.din(w_dff_A_F5NgWOo37_2),.clk(gclk));
	jdff dff_A_pwLbgITt6_2(.dout(w_dff_A_F5NgWOo37_2),.din(w_dff_A_pwLbgITt6_2),.clk(gclk));
	jdff dff_A_Pix1T5Ii7_1(.dout(w_G324_1[1]),.din(w_dff_A_Pix1T5Ii7_1),.clk(gclk));
	jdff dff_A_2Z0K9zBT8_1(.dout(w_G324_0[1]),.din(w_dff_A_2Z0K9zBT8_1),.clk(gclk));
	jdff dff_B_5ZvWoKPI1_1(.din(n1368),.dout(w_dff_B_5ZvWoKPI1_1),.clk(gclk));
	jdff dff_B_a6IBdNjb5_1(.din(w_dff_B_5ZvWoKPI1_1),.dout(w_dff_B_a6IBdNjb5_1),.clk(gclk));
	jdff dff_A_oRe2HLmT5_2(.dout(w_n388_0[2]),.din(w_dff_A_oRe2HLmT5_2),.clk(gclk));
	jdff dff_B_l9V0R11f7_3(.din(n388),.dout(w_dff_B_l9V0R11f7_3),.clk(gclk));
	jdff dff_A_tiWIMtFl5_0(.dout(w_G534_1[0]),.din(w_dff_A_tiWIMtFl5_0),.clk(gclk));
	jdff dff_A_SyTGvP4b2_0(.dout(w_dff_A_tiWIMtFl5_0),.din(w_dff_A_SyTGvP4b2_0),.clk(gclk));
	jdff dff_A_YqbMMSiH2_0(.dout(w_dff_A_SyTGvP4b2_0),.din(w_dff_A_YqbMMSiH2_0),.clk(gclk));
	jdff dff_A_JNMCiPQM9_1(.dout(w_G534_1[1]),.din(w_dff_A_JNMCiPQM9_1),.clk(gclk));
	jdff dff_B_5j4gjsAx5_1(.din(n1364),.dout(w_dff_B_5j4gjsAx5_1),.clk(gclk));
	jdff dff_A_UjBQH0Zl5_1(.dout(w_G351_2[1]),.din(w_dff_A_UjBQH0Zl5_1),.clk(gclk));
	jdff dff_A_B8ChI9y29_1(.dout(w_G534_0[1]),.din(w_dff_A_B8ChI9y29_1),.clk(gclk));
	jdff dff_A_mVrS8o4v7_1(.dout(w_dff_A_B8ChI9y29_1),.din(w_dff_A_mVrS8o4v7_1),.clk(gclk));
	jdff dff_A_VeZtSxbX9_2(.dout(w_G534_0[2]),.din(w_dff_A_VeZtSxbX9_2),.clk(gclk));
	jdff dff_A_D7QHmD778_2(.dout(w_dff_A_VeZtSxbX9_2),.din(w_dff_A_D7QHmD778_2),.clk(gclk));
	jdff dff_A_Lm3Wb03d5_2(.dout(w_dff_A_D7QHmD778_2),.din(w_dff_A_Lm3Wb03d5_2),.clk(gclk));
	jdff dff_A_fMakeybT3_0(.dout(w_G351_1[0]),.din(w_dff_A_fMakeybT3_0),.clk(gclk));
	jdff dff_A_PQWTlDM18_2(.dout(w_n410_0[2]),.din(w_dff_A_PQWTlDM18_2),.clk(gclk));
	jdff dff_A_qVwVWVcQ5_1(.dout(w_G514_0[1]),.din(w_dff_A_qVwVWVcQ5_1),.clk(gclk));
	jdff dff_A_co0w1ynH1_2(.dout(w_G514_0[2]),.din(w_dff_A_co0w1ynH1_2),.clk(gclk));
	jdff dff_A_XxixcFjb6_2(.dout(w_dff_A_co0w1ynH1_2),.din(w_dff_A_XxixcFjb6_2),.clk(gclk));
	jdff dff_A_RkoxuewP3_1(.dout(w_G361_0[1]),.din(w_dff_A_RkoxuewP3_1),.clk(gclk));
	jdff dff_B_CKFMWMZG7_1(.din(n1354),.dout(w_dff_B_CKFMWMZG7_1),.clk(gclk));
	jdff dff_B_vc2CbMzP1_1(.din(w_dff_B_CKFMWMZG7_1),.dout(w_dff_B_vc2CbMzP1_1),.clk(gclk));
	jdff dff_B_B0WxHOIX3_1(.din(n1355),.dout(w_dff_B_B0WxHOIX3_1),.clk(gclk));
	jdff dff_B_nUiidziz7_1(.din(n378),.dout(w_dff_B_nUiidziz7_1),.clk(gclk));
	jdff dff_B_kgP3d0345_1(.din(n379),.dout(w_dff_B_kgP3d0345_1),.clk(gclk));
	jdff dff_A_ttX26wiQ4_0(.dout(w_G490_1[0]),.din(w_dff_A_ttX26wiQ4_0),.clk(gclk));
	jdff dff_A_4sasHgEi3_0(.dout(w_dff_A_ttX26wiQ4_0),.din(w_dff_A_4sasHgEi3_0),.clk(gclk));
	jdff dff_A_IGH3UTH66_0(.dout(w_dff_A_4sasHgEi3_0),.din(w_dff_A_IGH3UTH66_0),.clk(gclk));
	jdff dff_A_t3kZlWYQ2_1(.dout(w_G490_1[1]),.din(w_dff_A_t3kZlWYQ2_1),.clk(gclk));
	jdff dff_A_B9NRc5n21_1(.dout(w_dff_A_t3kZlWYQ2_1),.din(w_dff_A_B9NRc5n21_1),.clk(gclk));
	jdff dff_A_aEpA6uPn7_1(.dout(w_G490_0[1]),.din(w_dff_A_aEpA6uPn7_1),.clk(gclk));
	jdff dff_A_scUGrfox5_1(.dout(w_dff_A_aEpA6uPn7_1),.din(w_dff_A_scUGrfox5_1),.clk(gclk));
	jdff dff_A_fwBz1ci64_1(.dout(w_dff_A_scUGrfox5_1),.din(w_dff_A_fwBz1ci64_1),.clk(gclk));
	jdff dff_A_PYBRhA2j5_2(.dout(w_G490_0[2]),.din(w_dff_A_PYBRhA2j5_2),.clk(gclk));
	jdff dff_A_LvCUOXXt4_2(.dout(w_dff_A_PYBRhA2j5_2),.din(w_dff_A_LvCUOXXt4_2),.clk(gclk));
	jdff dff_A_SDo89qRs2_2(.dout(w_dff_A_LvCUOXXt4_2),.din(w_dff_A_SDo89qRs2_2),.clk(gclk));
	jdff dff_A_uICwoGZT6_0(.dout(w_G316_1[0]),.din(w_dff_A_uICwoGZT6_0),.clk(gclk));
	jdff dff_B_zavP2zuO7_1(.din(n365),.dout(w_dff_B_zavP2zuO7_1),.clk(gclk));
	jdff dff_B_niiqv8J41_1(.din(n367),.dout(w_dff_B_niiqv8J41_1),.clk(gclk));
	jdff dff_A_ISTEQ5Zl6_0(.dout(w_n362_0[0]),.din(w_dff_A_ISTEQ5Zl6_0),.clk(gclk));
	jdff dff_A_08cq8yE56_0(.dout(w_dff_A_ISTEQ5Zl6_0),.din(w_dff_A_08cq8yE56_0),.clk(gclk));
	jdff dff_A_xQReP0PA4_0(.dout(w_dff_A_08cq8yE56_0),.din(w_dff_A_xQReP0PA4_0),.clk(gclk));
	jdff dff_A_lOm9er0S6_0(.dout(w_G479_1[0]),.din(w_dff_A_lOm9er0S6_0),.clk(gclk));
	jdff dff_A_vcbZ96Yk7_0(.dout(w_dff_A_lOm9er0S6_0),.din(w_dff_A_vcbZ96Yk7_0),.clk(gclk));
	jdff dff_A_KXyZwOVb4_1(.dout(w_G479_0[1]),.din(w_dff_A_KXyZwOVb4_1),.clk(gclk));
	jdff dff_A_nQy1rt4A1_1(.dout(w_dff_A_KXyZwOVb4_1),.din(w_dff_A_nQy1rt4A1_1),.clk(gclk));
	jdff dff_A_Pxom4RSw4_1(.dout(w_dff_A_nQy1rt4A1_1),.din(w_dff_A_Pxom4RSw4_1),.clk(gclk));
	jdff dff_A_oa0EixC20_2(.dout(w_G479_0[2]),.din(w_dff_A_oa0EixC20_2),.clk(gclk));
	jdff dff_A_9PnPWOgg8_2(.dout(w_dff_A_oa0EixC20_2),.din(w_dff_A_9PnPWOgg8_2),.clk(gclk));
	jdff dff_A_DFmdfCgD2_2(.dout(w_dff_A_9PnPWOgg8_2),.din(w_dff_A_DFmdfCgD2_2),.clk(gclk));
	jdff dff_A_dltZK1Z17_0(.dout(w_G308_1[0]),.din(w_dff_A_dltZK1Z17_0),.clk(gclk));
	jdff dff_A_W0RigKhz8_0(.dout(w_G302_0[0]),.din(w_dff_A_W0RigKhz8_0),.clk(gclk));
	jdff dff_A_CapWvRY64_1(.dout(w_G302_0[1]),.din(w_dff_A_CapWvRY64_1),.clk(gclk));
	jdff dff_A_r1l9bUN20_0(.dout(w_n401_0[0]),.din(w_dff_A_r1l9bUN20_0),.clk(gclk));
	jdff dff_A_fPmmE3xD9_2(.dout(w_n401_0[2]),.din(w_dff_A_fPmmE3xD9_2),.clk(gclk));
	jdff dff_A_e4wCn9PN4_1(.dout(w_G293_0[1]),.din(w_dff_A_e4wCn9PN4_1),.clk(gclk));
	jdff dff_B_PWP6gSHG7_1(.din(n1349),.dout(w_dff_B_PWP6gSHG7_1),.clk(gclk));
	jdff dff_B_Ycv7c5LF4_1(.din(n1350),.dout(w_dff_B_Ycv7c5LF4_1),.clk(gclk));
	jdff dff_A_yvXDm0ym2_0(.dout(w_n437_0[0]),.din(w_dff_A_yvXDm0ym2_0),.clk(gclk));
	jdff dff_A_swV2kJDX7_2(.dout(w_n437_0[2]),.din(w_dff_A_swV2kJDX7_2),.clk(gclk));
	jdff dff_A_mrHgL0da5_2(.dout(w_dff_A_swV2kJDX7_2),.din(w_dff_A_mrHgL0da5_2),.clk(gclk));
	jdff dff_A_w0Ny0zwc1_0(.dout(w_G523_1[0]),.din(w_dff_A_w0Ny0zwc1_0),.clk(gclk));
	jdff dff_A_wIkX4I6r0_1(.dout(w_G523_0[1]),.din(w_dff_A_wIkX4I6r0_1),.clk(gclk));
	jdff dff_A_37sMpk473_1(.dout(w_dff_A_wIkX4I6r0_1),.din(w_dff_A_37sMpk473_1),.clk(gclk));
	jdff dff_A_rfAUD5jN9_1(.dout(w_dff_A_37sMpk473_1),.din(w_dff_A_rfAUD5jN9_1),.clk(gclk));
	jdff dff_A_pg6AqhMU6_2(.dout(w_G523_0[2]),.din(w_dff_A_pg6AqhMU6_2),.clk(gclk));
	jdff dff_A_8rATMYQt0_2(.dout(w_dff_A_pg6AqhMU6_2),.din(w_dff_A_8rATMYQt0_2),.clk(gclk));
	jdff dff_A_kjapD70J7_1(.dout(w_G341_2[1]),.din(w_dff_A_kjapD70J7_1),.clk(gclk));
	jdff dff_A_LHr0g24r7_2(.dout(w_G341_0[2]),.din(w_dff_A_LHr0g24r7_2),.clk(gclk));
	jdff dff_A_eIiTMP0c2_2(.dout(w_n746_0[2]),.din(w_dff_A_eIiTMP0c2_2),.clk(gclk));
	jdff dff_A_QYCTBoZC8_2(.dout(w_dff_A_eIiTMP0c2_2),.din(w_dff_A_QYCTBoZC8_2),.clk(gclk));
	jdff dff_A_af19hOMD6_2(.dout(w_dff_A_QYCTBoZC8_2),.din(w_dff_A_af19hOMD6_2),.clk(gclk));
	jdff dff_A_BZOLwxXs5_2(.dout(w_dff_A_af19hOMD6_2),.din(w_dff_A_BZOLwxXs5_2),.clk(gclk));
	jdff dff_A_3cWjdMqw2_2(.dout(w_dff_A_BZOLwxXs5_2),.din(w_dff_A_3cWjdMqw2_2),.clk(gclk));
	jdff dff_A_wfSd7gzC5_2(.dout(w_dff_A_3cWjdMqw2_2),.din(w_dff_A_wfSd7gzC5_2),.clk(gclk));
	jdff dff_A_OuQiUOlc6_2(.dout(w_dff_A_wfSd7gzC5_2),.din(w_dff_A_OuQiUOlc6_2),.clk(gclk));
	jdff dff_A_xkSxuZlZ0_2(.dout(w_dff_A_OuQiUOlc6_2),.din(w_dff_A_xkSxuZlZ0_2),.clk(gclk));
	jdff dff_A_7I1tCCSc0_2(.dout(w_dff_A_xkSxuZlZ0_2),.din(w_dff_A_7I1tCCSc0_2),.clk(gclk));
	jdff dff_A_ZBsC8Br30_2(.dout(w_dff_A_7I1tCCSc0_2),.din(w_dff_A_ZBsC8Br30_2),.clk(gclk));
	jdff dff_A_Hlfz5tLw4_2(.dout(w_dff_A_ZBsC8Br30_2),.din(w_dff_A_Hlfz5tLw4_2),.clk(gclk));
	jdff dff_A_64vyYzxK4_0(.dout(w_n1002_1[0]),.din(w_dff_A_64vyYzxK4_0),.clk(gclk));
	jdff dff_A_sEBCiPbv9_0(.dout(w_dff_A_64vyYzxK4_0),.din(w_dff_A_sEBCiPbv9_0),.clk(gclk));
	jdff dff_A_vVt0nama4_0(.dout(w_dff_A_sEBCiPbv9_0),.din(w_dff_A_vVt0nama4_0),.clk(gclk));
	jdff dff_A_nITTOkrd7_0(.dout(w_dff_A_vVt0nama4_0),.din(w_dff_A_nITTOkrd7_0),.clk(gclk));
	jdff dff_A_OPJm0w7Y9_0(.dout(w_dff_A_nITTOkrd7_0),.din(w_dff_A_OPJm0w7Y9_0),.clk(gclk));
	jdff dff_A_ayovNCNM2_0(.dout(w_dff_A_OPJm0w7Y9_0),.din(w_dff_A_ayovNCNM2_0),.clk(gclk));
	jdff dff_A_PTUN5wli3_2(.dout(w_n1002_1[2]),.din(w_dff_A_PTUN5wli3_2),.clk(gclk));
	jdff dff_A_r2h4RkPj9_2(.dout(w_dff_A_PTUN5wli3_2),.din(w_dff_A_r2h4RkPj9_2),.clk(gclk));
	jdff dff_A_RFaQ96J16_2(.dout(w_dff_A_r2h4RkPj9_2),.din(w_dff_A_RFaQ96J16_2),.clk(gclk));
	jdff dff_A_YOzNbAII1_2(.dout(w_dff_A_RFaQ96J16_2),.din(w_dff_A_YOzNbAII1_2),.clk(gclk));
	jdff dff_A_AY38Xu2F2_2(.dout(w_dff_A_YOzNbAII1_2),.din(w_dff_A_AY38Xu2F2_2),.clk(gclk));
	jdff dff_A_U7VDY1450_2(.dout(w_dff_A_AY38Xu2F2_2),.din(w_dff_A_U7VDY1450_2),.clk(gclk));
	jdff dff_A_pGhWEDCn9_2(.dout(w_dff_A_U7VDY1450_2),.din(w_dff_A_pGhWEDCn9_2),.clk(gclk));
	jdff dff_A_uB5ORrbZ4_2(.dout(w_dff_A_pGhWEDCn9_2),.din(w_dff_A_uB5ORrbZ4_2),.clk(gclk));
	jdff dff_A_CZaORwpN2_2(.dout(w_dff_A_uB5ORrbZ4_2),.din(w_dff_A_CZaORwpN2_2),.clk(gclk));
	jdff dff_A_pC2Mo1fT7_2(.dout(w_dff_A_CZaORwpN2_2),.din(w_dff_A_pC2Mo1fT7_2),.clk(gclk));
	jdff dff_A_khWV93EV6_2(.dout(w_dff_A_pC2Mo1fT7_2),.din(w_dff_A_khWV93EV6_2),.clk(gclk));
	jdff dff_A_b2z9rtlA0_2(.dout(w_dff_A_khWV93EV6_2),.din(w_dff_A_b2z9rtlA0_2),.clk(gclk));
	jdff dff_A_W6o0McAd1_2(.dout(w_dff_A_b2z9rtlA0_2),.din(w_dff_A_W6o0McAd1_2),.clk(gclk));
	jdff dff_A_8JDSD9gO1_2(.dout(w_dff_A_W6o0McAd1_2),.din(w_dff_A_8JDSD9gO1_2),.clk(gclk));
	jdff dff_A_TUGSEb6r3_2(.dout(w_dff_A_8JDSD9gO1_2),.din(w_dff_A_TUGSEb6r3_2),.clk(gclk));
	jdff dff_A_CdOctyaS7_2(.dout(w_dff_A_TUGSEb6r3_2),.din(w_dff_A_CdOctyaS7_2),.clk(gclk));
	jdff dff_A_KEAJMF1s8_2(.dout(w_dff_A_CdOctyaS7_2),.din(w_dff_A_KEAJMF1s8_2),.clk(gclk));
	jdff dff_A_IMnGiKEn7_2(.dout(w_dff_A_KEAJMF1s8_2),.din(w_dff_A_IMnGiKEn7_2),.clk(gclk));
	jdff dff_A_dk9yo68N9_1(.dout(w_n1002_0[1]),.din(w_dff_A_dk9yo68N9_1),.clk(gclk));
	jdff dff_A_04zl8Bxc6_1(.dout(w_dff_A_dk9yo68N9_1),.din(w_dff_A_04zl8Bxc6_1),.clk(gclk));
	jdff dff_A_gbA2SURq8_1(.dout(w_dff_A_04zl8Bxc6_1),.din(w_dff_A_gbA2SURq8_1),.clk(gclk));
	jdff dff_A_TVlTtE6r7_1(.dout(w_dff_A_gbA2SURq8_1),.din(w_dff_A_TVlTtE6r7_1),.clk(gclk));
	jdff dff_A_4ym3sVNQ8_1(.dout(w_dff_A_TVlTtE6r7_1),.din(w_dff_A_4ym3sVNQ8_1),.clk(gclk));
	jdff dff_A_Ag4lhDMZ7_1(.dout(w_dff_A_4ym3sVNQ8_1),.din(w_dff_A_Ag4lhDMZ7_1),.clk(gclk));
	jdff dff_A_kIlvUKcO3_1(.dout(w_dff_A_Ag4lhDMZ7_1),.din(w_dff_A_kIlvUKcO3_1),.clk(gclk));
	jdff dff_A_mtxJGkWf4_1(.dout(w_dff_A_kIlvUKcO3_1),.din(w_dff_A_mtxJGkWf4_1),.clk(gclk));
	jdff dff_A_3F0yJgCq5_1(.dout(w_dff_A_mtxJGkWf4_1),.din(w_dff_A_3F0yJgCq5_1),.clk(gclk));
	jdff dff_A_1yFmmmqE0_1(.dout(w_dff_A_3F0yJgCq5_1),.din(w_dff_A_1yFmmmqE0_1),.clk(gclk));
	jdff dff_A_51HlVrDt5_1(.dout(w_dff_A_1yFmmmqE0_1),.din(w_dff_A_51HlVrDt5_1),.clk(gclk));
	jdff dff_A_kNEKMNe02_1(.dout(w_dff_A_51HlVrDt5_1),.din(w_dff_A_kNEKMNe02_1),.clk(gclk));
	jdff dff_A_zI6r6zWP1_1(.dout(w_dff_A_kNEKMNe02_1),.din(w_dff_A_zI6r6zWP1_1),.clk(gclk));
	jdff dff_A_bIKN2Bid9_1(.dout(w_dff_A_zI6r6zWP1_1),.din(w_dff_A_bIKN2Bid9_1),.clk(gclk));
	jdff dff_A_f2ED1Poh3_1(.dout(w_dff_A_bIKN2Bid9_1),.din(w_dff_A_f2ED1Poh3_1),.clk(gclk));
	jdff dff_A_q4v7VrV62_1(.dout(w_dff_A_f2ED1Poh3_1),.din(w_dff_A_q4v7VrV62_1),.clk(gclk));
	jdff dff_A_HZx7zHi24_2(.dout(w_n1002_0[2]),.din(w_dff_A_HZx7zHi24_2),.clk(gclk));
	jdff dff_A_QtZZ1elG6_2(.dout(w_dff_A_HZx7zHi24_2),.din(w_dff_A_QtZZ1elG6_2),.clk(gclk));
	jdff dff_A_2P6TUELz8_2(.dout(w_dff_A_QtZZ1elG6_2),.din(w_dff_A_2P6TUELz8_2),.clk(gclk));
	jdff dff_A_vLjItTvK2_2(.dout(w_dff_A_2P6TUELz8_2),.din(w_dff_A_vLjItTvK2_2),.clk(gclk));
	jdff dff_A_ROOgjzFz8_2(.dout(w_dff_A_vLjItTvK2_2),.din(w_dff_A_ROOgjzFz8_2),.clk(gclk));
	jdff dff_A_5YMBjLyY9_2(.dout(w_dff_A_ROOgjzFz8_2),.din(w_dff_A_5YMBjLyY9_2),.clk(gclk));
	jdff dff_A_Amqs3Bit9_2(.dout(w_dff_A_5YMBjLyY9_2),.din(w_dff_A_Amqs3Bit9_2),.clk(gclk));
	jdff dff_B_6OeN7K636_1(.din(n1641),.dout(w_dff_B_6OeN7K636_1),.clk(gclk));
	jdff dff_B_1L6o6Cko8_1(.din(w_dff_B_6OeN7K636_1),.dout(w_dff_B_1L6o6Cko8_1),.clk(gclk));
	jdff dff_B_ImqgfV7J8_1(.din(w_dff_B_1L6o6Cko8_1),.dout(w_dff_B_ImqgfV7J8_1),.clk(gclk));
	jdff dff_B_EtkgiWtu9_1(.din(w_dff_B_ImqgfV7J8_1),.dout(w_dff_B_EtkgiWtu9_1),.clk(gclk));
	jdff dff_B_cGk6N2sD5_1(.din(w_dff_B_EtkgiWtu9_1),.dout(w_dff_B_cGk6N2sD5_1),.clk(gclk));
	jdff dff_B_S3mB3zSa6_1(.din(w_dff_B_cGk6N2sD5_1),.dout(w_dff_B_S3mB3zSa6_1),.clk(gclk));
	jdff dff_B_CJd9RD5S0_1(.din(w_dff_B_S3mB3zSa6_1),.dout(w_dff_B_CJd9RD5S0_1),.clk(gclk));
	jdff dff_B_uVr5f8oh2_1(.din(w_dff_B_CJd9RD5S0_1),.dout(w_dff_B_uVr5f8oh2_1),.clk(gclk));
	jdff dff_B_2wz2D0Pr1_1(.din(w_dff_B_uVr5f8oh2_1),.dout(w_dff_B_2wz2D0Pr1_1),.clk(gclk));
	jdff dff_B_8hrJ0wYW1_1(.din(w_dff_B_2wz2D0Pr1_1),.dout(w_dff_B_8hrJ0wYW1_1),.clk(gclk));
	jdff dff_B_R5F530526_1(.din(w_dff_B_8hrJ0wYW1_1),.dout(w_dff_B_R5F530526_1),.clk(gclk));
	jdff dff_B_souuacIB0_1(.din(w_dff_B_R5F530526_1),.dout(w_dff_B_souuacIB0_1),.clk(gclk));
	jdff dff_B_JRWM6lha9_1(.din(w_dff_B_souuacIB0_1),.dout(w_dff_B_JRWM6lha9_1),.clk(gclk));
	jdff dff_B_lyvI4CwF3_1(.din(w_dff_B_JRWM6lha9_1),.dout(w_dff_B_lyvI4CwF3_1),.clk(gclk));
	jdff dff_B_4GmtljTw5_1(.din(w_dff_B_lyvI4CwF3_1),.dout(w_dff_B_4GmtljTw5_1),.clk(gclk));
	jdff dff_B_76yLKDrR8_1(.din(w_dff_B_4GmtljTw5_1),.dout(w_dff_B_76yLKDrR8_1),.clk(gclk));
	jdff dff_B_Yx8Y5mBm5_1(.din(w_dff_B_76yLKDrR8_1),.dout(w_dff_B_Yx8Y5mBm5_1),.clk(gclk));
	jdff dff_B_jNzKA38i4_1(.din(w_dff_B_Yx8Y5mBm5_1),.dout(w_dff_B_jNzKA38i4_1),.clk(gclk));
	jdff dff_B_n3cs1FfX4_1(.din(w_dff_B_jNzKA38i4_1),.dout(w_dff_B_n3cs1FfX4_1),.clk(gclk));
	jdff dff_B_EhJkZzbA4_0(.din(n1600),.dout(w_dff_B_EhJkZzbA4_0),.clk(gclk));
	jdff dff_B_HS69KahT6_0(.din(w_dff_B_EhJkZzbA4_0),.dout(w_dff_B_HS69KahT6_0),.clk(gclk));
	jdff dff_B_ThUFz0mE9_0(.din(w_dff_B_HS69KahT6_0),.dout(w_dff_B_ThUFz0mE9_0),.clk(gclk));
	jdff dff_B_HnE2ciiS9_0(.din(w_dff_B_ThUFz0mE9_0),.dout(w_dff_B_HnE2ciiS9_0),.clk(gclk));
	jdff dff_B_93OsQDIC7_0(.din(w_dff_B_HnE2ciiS9_0),.dout(w_dff_B_93OsQDIC7_0),.clk(gclk));
	jdff dff_B_H20Gu3l83_0(.din(w_dff_B_93OsQDIC7_0),.dout(w_dff_B_H20Gu3l83_0),.clk(gclk));
	jdff dff_B_A7CSZ7zs0_0(.din(w_dff_B_H20Gu3l83_0),.dout(w_dff_B_A7CSZ7zs0_0),.clk(gclk));
	jdff dff_B_hj6k4AW68_0(.din(w_dff_B_A7CSZ7zs0_0),.dout(w_dff_B_hj6k4AW68_0),.clk(gclk));
	jdff dff_B_LtaItCx80_0(.din(w_dff_B_hj6k4AW68_0),.dout(w_dff_B_LtaItCx80_0),.clk(gclk));
	jdff dff_B_mBGTLlPb7_0(.din(w_dff_B_LtaItCx80_0),.dout(w_dff_B_mBGTLlPb7_0),.clk(gclk));
	jdff dff_B_hjTfYdzz3_0(.din(w_dff_B_mBGTLlPb7_0),.dout(w_dff_B_hjTfYdzz3_0),.clk(gclk));
	jdff dff_B_hmLUvkg22_0(.din(w_dff_B_hjTfYdzz3_0),.dout(w_dff_B_hmLUvkg22_0),.clk(gclk));
	jdff dff_B_CIp1uF8m0_0(.din(w_dff_B_hmLUvkg22_0),.dout(w_dff_B_CIp1uF8m0_0),.clk(gclk));
	jdff dff_B_tGGze2J71_0(.din(w_dff_B_CIp1uF8m0_0),.dout(w_dff_B_tGGze2J71_0),.clk(gclk));
	jdff dff_B_yCJCVwuc5_0(.din(w_dff_B_tGGze2J71_0),.dout(w_dff_B_yCJCVwuc5_0),.clk(gclk));
	jdff dff_B_2khqw2AR0_0(.din(w_dff_B_yCJCVwuc5_0),.dout(w_dff_B_2khqw2AR0_0),.clk(gclk));
	jdff dff_B_gQ3HQZ7w5_0(.din(w_dff_B_2khqw2AR0_0),.dout(w_dff_B_gQ3HQZ7w5_0),.clk(gclk));
	jdff dff_B_AsoKSNIU2_0(.din(w_dff_B_gQ3HQZ7w5_0),.dout(w_dff_B_AsoKSNIU2_0),.clk(gclk));
	jdff dff_B_88vVCwdc4_0(.din(w_dff_B_AsoKSNIU2_0),.dout(w_dff_B_88vVCwdc4_0),.clk(gclk));
	jdff dff_B_Qf1PQoZZ5_1(.din(n1540),.dout(w_dff_B_Qf1PQoZZ5_1),.clk(gclk));
	jdff dff_B_GncxnPhC1_1(.din(w_dff_B_Qf1PQoZZ5_1),.dout(w_dff_B_GncxnPhC1_1),.clk(gclk));
	jdff dff_B_c4GH5yc22_1(.din(w_dff_B_GncxnPhC1_1),.dout(w_dff_B_c4GH5yc22_1),.clk(gclk));
	jdff dff_B_6zxqdXAJ4_1(.din(w_dff_B_c4GH5yc22_1),.dout(w_dff_B_6zxqdXAJ4_1),.clk(gclk));
	jdff dff_B_mcGzYXIk5_1(.din(w_dff_B_6zxqdXAJ4_1),.dout(w_dff_B_mcGzYXIk5_1),.clk(gclk));
	jdff dff_B_L99eLpKe4_1(.din(w_dff_B_mcGzYXIk5_1),.dout(w_dff_B_L99eLpKe4_1),.clk(gclk));
	jdff dff_B_Jrysdmbr7_1(.din(w_dff_B_L99eLpKe4_1),.dout(w_dff_B_Jrysdmbr7_1),.clk(gclk));
	jdff dff_B_KSw97FQY9_1(.din(w_dff_B_Jrysdmbr7_1),.dout(w_dff_B_KSw97FQY9_1),.clk(gclk));
	jdff dff_B_pKrQqRjP2_0(.din(n1589),.dout(w_dff_B_pKrQqRjP2_0),.clk(gclk));
	jdff dff_B_5sQTU8zG9_0(.din(w_dff_B_pKrQqRjP2_0),.dout(w_dff_B_5sQTU8zG9_0),.clk(gclk));
	jdff dff_B_nhICFsvk8_1(.din(n1579),.dout(w_dff_B_nhICFsvk8_1),.clk(gclk));
	jdff dff_B_EtgMCAiT2_0(.din(n1586),.dout(w_dff_B_EtgMCAiT2_0),.clk(gclk));
	jdff dff_B_WVLqhli38_0(.din(w_dff_B_EtgMCAiT2_0),.dout(w_dff_B_WVLqhli38_0),.clk(gclk));
	jdff dff_B_0qPXDqtW9_0(.din(w_dff_B_WVLqhli38_0),.dout(w_dff_B_0qPXDqtW9_0),.clk(gclk));
	jdff dff_B_I3DZOT0N9_0(.din(n1584),.dout(w_dff_B_I3DZOT0N9_0),.clk(gclk));
	jdff dff_B_EVlwy7Ax0_1(.din(n1567),.dout(w_dff_B_EVlwy7Ax0_1),.clk(gclk));
	jdff dff_B_2MbpbnbB1_1(.din(w_dff_B_EVlwy7Ax0_1),.dout(w_dff_B_2MbpbnbB1_1),.clk(gclk));
	jdff dff_B_J2KV0Fnw6_1(.din(w_dff_B_2MbpbnbB1_1),.dout(w_dff_B_J2KV0Fnw6_1),.clk(gclk));
	jdff dff_B_0aGJ5bAa9_1(.din(w_dff_B_J2KV0Fnw6_1),.dout(w_dff_B_0aGJ5bAa9_1),.clk(gclk));
	jdff dff_B_1qJTC31r1_1(.din(w_dff_B_0aGJ5bAa9_1),.dout(w_dff_B_1qJTC31r1_1),.clk(gclk));
	jdff dff_B_2yjrLfHS5_1(.din(w_dff_B_1qJTC31r1_1),.dout(w_dff_B_2yjrLfHS5_1),.clk(gclk));
	jdff dff_B_YeW9ImRd9_1(.din(w_dff_B_2yjrLfHS5_1),.dout(w_dff_B_YeW9ImRd9_1),.clk(gclk));
	jdff dff_B_3KhERs6R8_1(.din(w_dff_B_YeW9ImRd9_1),.dout(w_dff_B_3KhERs6R8_1),.clk(gclk));
	jdff dff_B_1CoSnAiy8_1(.din(w_dff_B_3KhERs6R8_1),.dout(w_dff_B_1CoSnAiy8_1),.clk(gclk));
	jdff dff_B_XdrxUKX55_1(.din(w_dff_B_1CoSnAiy8_1),.dout(w_dff_B_XdrxUKX55_1),.clk(gclk));
	jdff dff_B_O9rHUWWP6_1(.din(w_dff_B_XdrxUKX55_1),.dout(w_dff_B_O9rHUWWP6_1),.clk(gclk));
	jdff dff_B_ybm314OY6_1(.din(w_dff_B_O9rHUWWP6_1),.dout(w_dff_B_ybm314OY6_1),.clk(gclk));
	jdff dff_B_wBB2siGO4_1(.din(w_dff_B_ybm314OY6_1),.dout(w_dff_B_wBB2siGO4_1),.clk(gclk));
	jdff dff_B_Pwv1sH3P1_1(.din(n1570),.dout(w_dff_B_Pwv1sH3P1_1),.clk(gclk));
	jdff dff_B_Y8zfDsM18_1(.din(w_dff_B_Pwv1sH3P1_1),.dout(w_dff_B_Y8zfDsM18_1),.clk(gclk));
	jdff dff_B_sMf275Oj5_1(.din(w_dff_B_Y8zfDsM18_1),.dout(w_dff_B_sMf275Oj5_1),.clk(gclk));
	jdff dff_B_CdlBZLKv8_1(.din(w_dff_B_sMf275Oj5_1),.dout(w_dff_B_CdlBZLKv8_1),.clk(gclk));
	jdff dff_B_TB6HaPrd4_1(.din(n1571),.dout(w_dff_B_TB6HaPrd4_1),.clk(gclk));
	jdff dff_B_6Th0vuFA4_1(.din(w_dff_B_TB6HaPrd4_1),.dout(w_dff_B_6Th0vuFA4_1),.clk(gclk));
	jdff dff_B_U2djDFY16_1(.din(w_dff_B_6Th0vuFA4_1),.dout(w_dff_B_U2djDFY16_1),.clk(gclk));
	jdff dff_B_2XTWqIPU0_1(.din(w_dff_B_U2djDFY16_1),.dout(w_dff_B_2XTWqIPU0_1),.clk(gclk));
	jdff dff_B_K30Kxw1G5_1(.din(w_dff_B_2XTWqIPU0_1),.dout(w_dff_B_K30Kxw1G5_1),.clk(gclk));
	jdff dff_B_To8vsBxy8_1(.din(w_dff_B_K30Kxw1G5_1),.dout(w_dff_B_To8vsBxy8_1),.clk(gclk));
	jdff dff_A_VeQVEag42_0(.dout(w_n855_0[0]),.din(w_dff_A_VeQVEag42_0),.clk(gclk));
	jdff dff_A_zx1Zjokm5_1(.dout(w_n853_0[1]),.din(w_dff_A_zx1Zjokm5_1),.clk(gclk));
	jdff dff_B_5bPD11Zu0_2(.din(n853),.dout(w_dff_B_5bPD11Zu0_2),.clk(gclk));
	jdff dff_B_8f7Rwor92_2(.din(w_dff_B_5bPD11Zu0_2),.dout(w_dff_B_8f7Rwor92_2),.clk(gclk));
	jdff dff_B_b8zsgBWp5_2(.din(w_dff_B_8f7Rwor92_2),.dout(w_dff_B_b8zsgBWp5_2),.clk(gclk));
	jdff dff_B_Ro7kTiWC3_2(.din(w_dff_B_b8zsgBWp5_2),.dout(w_dff_B_Ro7kTiWC3_2),.clk(gclk));
	jdff dff_A_xCxv6HKT2_0(.dout(w_n681_1[0]),.din(w_dff_A_xCxv6HKT2_0),.clk(gclk));
	jdff dff_A_HUQ0FT1o3_0(.dout(w_dff_A_xCxv6HKT2_0),.din(w_dff_A_HUQ0FT1o3_0),.clk(gclk));
	jdff dff_A_2Z8mXk8k5_0(.dout(w_dff_A_HUQ0FT1o3_0),.din(w_dff_A_2Z8mXk8k5_0),.clk(gclk));
	jdff dff_A_Z01nOi0E2_0(.dout(w_dff_A_2Z8mXk8k5_0),.din(w_dff_A_Z01nOi0E2_0),.clk(gclk));
	jdff dff_A_xySRvejU7_1(.dout(w_n681_1[1]),.din(w_dff_A_xySRvejU7_1),.clk(gclk));
	jdff dff_A_cq8EeuVL6_1(.dout(w_n1568_0[1]),.din(w_dff_A_cq8EeuVL6_1),.clk(gclk));
	jdff dff_B_Aqgco1yP8_1(.din(n1562),.dout(w_dff_B_Aqgco1yP8_1),.clk(gclk));
	jdff dff_B_R3AsyGgd0_0(.din(n1563),.dout(w_dff_B_R3AsyGgd0_0),.clk(gclk));
	jdff dff_B_2c3jPkB65_1(.din(n1557),.dout(w_dff_B_2c3jPkB65_1),.clk(gclk));
	jdff dff_A_kbnB72tY6_0(.dout(w_n1555_0[0]),.din(w_dff_A_kbnB72tY6_0),.clk(gclk));
	jdff dff_A_jvBsZeVC2_0(.dout(w_dff_A_kbnB72tY6_0),.din(w_dff_A_jvBsZeVC2_0),.clk(gclk));
	jdff dff_B_JwbTmWEP5_2(.din(n1553),.dout(w_dff_B_JwbTmWEP5_2),.clk(gclk));
	jdff dff_B_bV4ITsi30_2(.din(w_dff_B_JwbTmWEP5_2),.dout(w_dff_B_bV4ITsi30_2),.clk(gclk));
	jdff dff_B_PMsOGxPU2_2(.din(w_dff_B_bV4ITsi30_2),.dout(w_dff_B_PMsOGxPU2_2),.clk(gclk));
	jdff dff_B_o6QtMK7q2_2(.din(w_dff_B_PMsOGxPU2_2),.dout(w_dff_B_o6QtMK7q2_2),.clk(gclk));
	jdff dff_B_XU6W4ozn0_2(.din(w_dff_B_o6QtMK7q2_2),.dout(w_dff_B_XU6W4ozn0_2),.clk(gclk));
	jdff dff_B_Dy6tX2Yq7_2(.din(w_dff_B_XU6W4ozn0_2),.dout(w_dff_B_Dy6tX2Yq7_2),.clk(gclk));
	jdff dff_B_zwWypTr77_0(.din(n1551),.dout(w_dff_B_zwWypTr77_0),.clk(gclk));
	jdff dff_B_Owq66JFL6_0(.din(w_dff_B_zwWypTr77_0),.dout(w_dff_B_Owq66JFL6_0),.clk(gclk));
	jdff dff_B_ulmeB7oI0_0(.din(w_dff_B_Owq66JFL6_0),.dout(w_dff_B_ulmeB7oI0_0),.clk(gclk));
	jdff dff_B_yWXPpkU14_0(.din(n1550),.dout(w_dff_B_yWXPpkU14_0),.clk(gclk));
	jdff dff_B_Cxu0AvQP9_0(.din(w_dff_B_yWXPpkU14_0),.dout(w_dff_B_Cxu0AvQP9_0),.clk(gclk));
	jdff dff_B_SqxMVJQv9_0(.din(w_dff_B_Cxu0AvQP9_0),.dout(w_dff_B_SqxMVJQv9_0),.clk(gclk));
	jdff dff_B_SWU0Og0K2_0(.din(w_dff_B_SqxMVJQv9_0),.dout(w_dff_B_SWU0Og0K2_0),.clk(gclk));
	jdff dff_B_F6fTFBFL8_0(.din(w_dff_B_SWU0Og0K2_0),.dout(w_dff_B_F6fTFBFL8_0),.clk(gclk));
	jdff dff_A_3ja49RM29_2(.dout(w_n605_1[2]),.din(w_dff_A_3ja49RM29_2),.clk(gclk));
	jdff dff_A_wWqxvnFh5_2(.dout(w_dff_A_3ja49RM29_2),.din(w_dff_A_wWqxvnFh5_2),.clk(gclk));
	jdff dff_A_Gtb5rL9D6_2(.dout(w_dff_A_wWqxvnFh5_2),.din(w_dff_A_Gtb5rL9D6_2),.clk(gclk));
	jdff dff_A_RHBgMXWQ6_2(.dout(w_dff_A_Gtb5rL9D6_2),.din(w_dff_A_RHBgMXWQ6_2),.clk(gclk));
	jdff dff_A_aj8ithYg8_2(.dout(w_dff_A_RHBgMXWQ6_2),.din(w_dff_A_aj8ithYg8_2),.clk(gclk));
	jdff dff_A_S6JWOdGf1_2(.dout(w_dff_A_aj8ithYg8_2),.din(w_dff_A_S6JWOdGf1_2),.clk(gclk));
	jdff dff_A_WrZMAIQo0_2(.dout(w_dff_A_S6JWOdGf1_2),.din(w_dff_A_WrZMAIQo0_2),.clk(gclk));
	jdff dff_A_tc2FYKIM4_2(.dout(w_dff_A_WrZMAIQo0_2),.din(w_dff_A_tc2FYKIM4_2),.clk(gclk));
	jdff dff_A_OciTwPi61_2(.dout(w_dff_A_tc2FYKIM4_2),.din(w_dff_A_OciTwPi61_2),.clk(gclk));
	jdff dff_A_fHwo9xj71_2(.dout(w_dff_A_OciTwPi61_2),.din(w_dff_A_fHwo9xj71_2),.clk(gclk));
	jdff dff_A_jmPxkNvb8_2(.dout(w_dff_A_fHwo9xj71_2),.din(w_dff_A_jmPxkNvb8_2),.clk(gclk));
	jdff dff_A_YNBRqcRa7_2(.dout(w_dff_A_jmPxkNvb8_2),.din(w_dff_A_YNBRqcRa7_2),.clk(gclk));
	jdff dff_A_nHigQEHp3_1(.dout(w_n944_0[1]),.din(w_dff_A_nHigQEHp3_1),.clk(gclk));
	jdff dff_A_VEZ2Lyt87_1(.dout(w_dff_A_nHigQEHp3_1),.din(w_dff_A_VEZ2Lyt87_1),.clk(gclk));
	jdff dff_A_WC2N9Msk0_1(.dout(w_dff_A_VEZ2Lyt87_1),.din(w_dff_A_WC2N9Msk0_1),.clk(gclk));
	jdff dff_A_YAC9j1oB7_1(.dout(w_dff_A_WC2N9Msk0_1),.din(w_dff_A_YAC9j1oB7_1),.clk(gclk));
	jdff dff_A_Dl0Ry4UP1_1(.dout(w_dff_A_YAC9j1oB7_1),.din(w_dff_A_Dl0Ry4UP1_1),.clk(gclk));
	jdff dff_A_0MglTAon8_1(.dout(w_dff_A_Dl0Ry4UP1_1),.din(w_dff_A_0MglTAon8_1),.clk(gclk));
	jdff dff_A_y2HKCHyV4_1(.dout(w_dff_A_0MglTAon8_1),.din(w_dff_A_y2HKCHyV4_1),.clk(gclk));
	jdff dff_A_0EKC9WTT4_1(.dout(w_dff_A_y2HKCHyV4_1),.din(w_dff_A_0EKC9WTT4_1),.clk(gclk));
	jdff dff_A_IhjvjxkU8_1(.dout(w_dff_A_0EKC9WTT4_1),.din(w_dff_A_IhjvjxkU8_1),.clk(gclk));
	jdff dff_A_tpeqpbPU1_2(.dout(w_n930_0[2]),.din(w_dff_A_tpeqpbPU1_2),.clk(gclk));
	jdff dff_A_VbBdf96I2_2(.dout(w_dff_A_tpeqpbPU1_2),.din(w_dff_A_VbBdf96I2_2),.clk(gclk));
	jdff dff_A_swWSomix1_2(.dout(w_dff_A_VbBdf96I2_2),.din(w_dff_A_swWSomix1_2),.clk(gclk));
	jdff dff_A_4WZEEWt28_2(.dout(w_dff_A_swWSomix1_2),.din(w_dff_A_4WZEEWt28_2),.clk(gclk));
	jdff dff_A_ic1Sd5dt8_2(.dout(w_dff_A_4WZEEWt28_2),.din(w_dff_A_ic1Sd5dt8_2),.clk(gclk));
	jdff dff_A_cisqXhkJ5_2(.dout(w_dff_A_ic1Sd5dt8_2),.din(w_dff_A_cisqXhkJ5_2),.clk(gclk));
	jdff dff_A_Ad3UL6lH1_2(.dout(w_dff_A_cisqXhkJ5_2),.din(w_dff_A_Ad3UL6lH1_2),.clk(gclk));
	jdff dff_A_QjPZEWqj8_2(.dout(w_dff_A_Ad3UL6lH1_2),.din(w_dff_A_QjPZEWqj8_2),.clk(gclk));
	jdff dff_A_PFBHx6OY6_2(.dout(w_dff_A_QjPZEWqj8_2),.din(w_dff_A_PFBHx6OY6_2),.clk(gclk));
	jdff dff_B_blt8YHHv2_3(.din(n930),.dout(w_dff_B_blt8YHHv2_3),.clk(gclk));
	jdff dff_B_ue2FJvjL9_3(.din(w_dff_B_blt8YHHv2_3),.dout(w_dff_B_ue2FJvjL9_3),.clk(gclk));
	jdff dff_A_mWZi5Wvh4_1(.dout(w_n700_0[1]),.din(w_dff_A_mWZi5Wvh4_1),.clk(gclk));
	jdff dff_A_rt1CipLT7_1(.dout(w_dff_A_mWZi5Wvh4_1),.din(w_dff_A_rt1CipLT7_1),.clk(gclk));
	jdff dff_A_IMU7GyEl9_1(.dout(w_dff_A_rt1CipLT7_1),.din(w_dff_A_IMU7GyEl9_1),.clk(gclk));
	jdff dff_A_Bi2zBv3k9_0(.dout(w_n706_0[0]),.din(w_dff_A_Bi2zBv3k9_0),.clk(gclk));
	jdff dff_B_xyvvpyID3_1(.din(n701),.dout(w_dff_B_xyvvpyID3_1),.clk(gclk));
	jdff dff_B_QoISKYFR2_1(.din(w_dff_B_xyvvpyID3_1),.dout(w_dff_B_QoISKYFR2_1),.clk(gclk));
	jdff dff_B_Gw3mBlYD2_0(.din(n599),.dout(w_dff_B_Gw3mBlYD2_0),.clk(gclk));
	jdff dff_B_RdkYRMhY3_1(.din(G233),.dout(w_dff_B_RdkYRMhY3_1),.clk(gclk));
	jdff dff_B_8MNPYt2H8_2(.din(n702),.dout(w_dff_B_8MNPYt2H8_2),.clk(gclk));
	jdff dff_A_MVAVHnvF7_0(.dout(w_n604_0[0]),.din(w_dff_A_MVAVHnvF7_0),.clk(gclk));
	jdff dff_B_lJJhKMIC2_0(.din(n603),.dout(w_dff_B_lJJhKMIC2_0),.clk(gclk));
	jdff dff_B_OGZ3SmVF3_1(.din(G225),.dout(w_dff_B_OGZ3SmVF3_1),.clk(gclk));
	jdff dff_A_4PZcCC7F9_1(.dout(w_n928_0[1]),.din(w_dff_A_4PZcCC7F9_1),.clk(gclk));
	jdff dff_A_rU9nK9bv2_1(.dout(w_dff_A_4PZcCC7F9_1),.din(w_dff_A_rU9nK9bv2_1),.clk(gclk));
	jdff dff_A_N3VTAcw44_1(.dout(w_dff_A_rU9nK9bv2_1),.din(w_dff_A_N3VTAcw44_1),.clk(gclk));
	jdff dff_A_PcBj3BQH4_1(.dout(w_dff_A_N3VTAcw44_1),.din(w_dff_A_PcBj3BQH4_1),.clk(gclk));
	jdff dff_A_XcUoOKCH7_1(.dout(w_dff_A_PcBj3BQH4_1),.din(w_dff_A_XcUoOKCH7_1),.clk(gclk));
	jdff dff_A_X4NFrEQU5_1(.dout(w_dff_A_XcUoOKCH7_1),.din(w_dff_A_X4NFrEQU5_1),.clk(gclk));
	jdff dff_A_9kFtfxdw7_1(.dout(w_dff_A_X4NFrEQU5_1),.din(w_dff_A_9kFtfxdw7_1),.clk(gclk));
	jdff dff_A_Dt7atwku0_1(.dout(w_dff_A_9kFtfxdw7_1),.din(w_dff_A_Dt7atwku0_1),.clk(gclk));
	jdff dff_A_vb0eqkuN8_1(.dout(w_dff_A_Dt7atwku0_1),.din(w_dff_A_vb0eqkuN8_1),.clk(gclk));
	jdff dff_B_QCKE4Vj84_2(.din(n928),.dout(w_dff_B_QCKE4Vj84_2),.clk(gclk));
	jdff dff_B_njDmDYvj6_2(.din(w_dff_B_QCKE4Vj84_2),.dout(w_dff_B_njDmDYvj6_2),.clk(gclk));
	jdff dff_B_rI3rDfQO6_2(.din(w_dff_B_njDmDYvj6_2),.dout(w_dff_B_rI3rDfQO6_2),.clk(gclk));
	jdff dff_A_RcQxCNTJ4_0(.dout(w_n596_0[0]),.din(w_dff_A_RcQxCNTJ4_0),.clk(gclk));
	jdff dff_A_lJFZsVQE5_0(.dout(w_dff_A_RcQxCNTJ4_0),.din(w_dff_A_lJFZsVQE5_0),.clk(gclk));
	jdff dff_A_PEsInGMZ2_0(.dout(w_dff_A_lJFZsVQE5_0),.din(w_dff_A_PEsInGMZ2_0),.clk(gclk));
	jdff dff_A_qojEt2kH7_0(.dout(w_dff_A_PEsInGMZ2_0),.din(w_dff_A_qojEt2kH7_0),.clk(gclk));
	jdff dff_A_F0ZZ8ljA9_0(.dout(w_dff_A_qojEt2kH7_0),.din(w_dff_A_F0ZZ8ljA9_0),.clk(gclk));
	jdff dff_B_EBnxoP7t6_1(.din(n592),.dout(w_dff_B_EBnxoP7t6_1),.clk(gclk));
	jdff dff_B_eO5eMZRj6_1(.din(G209),.dout(w_dff_B_eO5eMZRj6_1),.clk(gclk));
	jdff dff_B_LWCDxLKe9_0(.din(n1544),.dout(w_dff_B_LWCDxLKe9_0),.clk(gclk));
	jdff dff_A_pEJMJpr07_0(.dout(w_n585_0[0]),.din(w_dff_A_pEJMJpr07_0),.clk(gclk));
	jdff dff_B_MniNMeSj0_0(.din(n584),.dout(w_dff_B_MniNMeSj0_0),.clk(gclk));
	jdff dff_B_zyEKpJaB5_0(.din(w_dff_B_MniNMeSj0_0),.dout(w_dff_B_zyEKpJaB5_0),.clk(gclk));
	jdff dff_A_1F8jFF1c1_0(.dout(w_n583_1[0]),.din(w_dff_A_1F8jFF1c1_0),.clk(gclk));
	jdff dff_A_qfSiuZc81_0(.dout(w_dff_A_1F8jFF1c1_0),.din(w_dff_A_qfSiuZc81_0),.clk(gclk));
	jdff dff_A_rBYzm1ut3_0(.dout(w_dff_A_qfSiuZc81_0),.din(w_dff_A_rBYzm1ut3_0),.clk(gclk));
	jdff dff_A_PDsN4Y8C0_0(.dout(w_n572_0[0]),.din(w_dff_A_PDsN4Y8C0_0),.clk(gclk));
	jdff dff_A_HNJiObHX0_0(.dout(w_dff_A_PDsN4Y8C0_0),.din(w_dff_A_HNJiObHX0_0),.clk(gclk));
	jdff dff_A_RbbxnHEB6_0(.dout(w_dff_A_HNJiObHX0_0),.din(w_dff_A_RbbxnHEB6_0),.clk(gclk));
	jdff dff_A_s3a2UhOY3_0(.dout(w_dff_A_RbbxnHEB6_0),.din(w_dff_A_s3a2UhOY3_0),.clk(gclk));
	jdff dff_A_rNtdnGCB4_1(.dout(w_n567_1[1]),.din(w_dff_A_rNtdnGCB4_1),.clk(gclk));
	jdff dff_A_Pi97kgwG7_1(.dout(w_n567_0[1]),.din(w_dff_A_Pi97kgwG7_1),.clk(gclk));
	jdff dff_A_bZmkYIdN2_1(.dout(w_dff_A_Pi97kgwG7_1),.din(w_dff_A_bZmkYIdN2_1),.clk(gclk));
	jdff dff_A_F5A5MZ505_1(.dout(w_dff_A_bZmkYIdN2_1),.din(w_dff_A_F5A5MZ505_1),.clk(gclk));
	jdff dff_A_ixbpSxxm4_0(.dout(w_n497_1[0]),.din(w_dff_A_ixbpSxxm4_0),.clk(gclk));
	jdff dff_A_Zn2BH9Cy0_0(.dout(w_n562_0[0]),.din(w_dff_A_Zn2BH9Cy0_0),.clk(gclk));
	jdff dff_A_M3mLHJYX1_0(.dout(w_dff_A_Zn2BH9Cy0_0),.din(w_dff_A_M3mLHJYX1_0),.clk(gclk));
	jdff dff_A_CtxohyMF6_0(.dout(w_dff_A_M3mLHJYX1_0),.din(w_dff_A_CtxohyMF6_0),.clk(gclk));
	jdff dff_A_PA9ynngi7_0(.dout(w_dff_A_CtxohyMF6_0),.din(w_dff_A_PA9ynngi7_0),.clk(gclk));
	jdff dff_A_0pE0wOE56_0(.dout(w_dff_A_PA9ynngi7_0),.din(w_dff_A_0pE0wOE56_0),.clk(gclk));
	jdff dff_B_TQvuXTWR4_2(.din(n562),.dout(w_dff_B_TQvuXTWR4_2),.clk(gclk));
	jdff dff_B_Vhp7DYjM5_2(.din(w_dff_B_TQvuXTWR4_2),.dout(w_dff_B_Vhp7DYjM5_2),.clk(gclk));
	jdff dff_A_Rzp9MT8F9_0(.dout(w_n561_0[0]),.din(w_dff_A_Rzp9MT8F9_0),.clk(gclk));
	jdff dff_A_VyHLCHxB8_1(.dout(w_n561_0[1]),.din(w_dff_A_VyHLCHxB8_1),.clk(gclk));
	jdff dff_A_giEofqP28_1(.dout(w_dff_A_VyHLCHxB8_1),.din(w_dff_A_giEofqP28_1),.clk(gclk));
	jdff dff_A_9OAdvTyj2_1(.dout(w_dff_A_giEofqP28_1),.din(w_dff_A_9OAdvTyj2_1),.clk(gclk));
	jdff dff_A_yfszB5K62_0(.dout(w_G1497_0[0]),.din(w_dff_A_yfszB5K62_0),.clk(gclk));
	jdff dff_A_a9ABx1MJ6_0(.dout(w_dff_A_yfszB5K62_0),.din(w_dff_A_a9ABx1MJ6_0),.clk(gclk));
	jdff dff_A_nXjwNtcd7_0(.dout(w_dff_A_a9ABx1MJ6_0),.din(w_dff_A_nXjwNtcd7_0),.clk(gclk));
	jdff dff_A_vaZlhGfN7_0(.dout(w_dff_A_nXjwNtcd7_0),.din(w_dff_A_vaZlhGfN7_0),.clk(gclk));
	jdff dff_A_G8o9lxgE4_0(.dout(w_dff_A_vaZlhGfN7_0),.din(w_dff_A_G8o9lxgE4_0),.clk(gclk));
	jdff dff_A_g5x9RPCW1_0(.dout(w_dff_A_G8o9lxgE4_0),.din(w_dff_A_g5x9RPCW1_0),.clk(gclk));
	jdff dff_A_cBTUSIlK9_0(.dout(w_dff_A_g5x9RPCW1_0),.din(w_dff_A_cBTUSIlK9_0),.clk(gclk));
	jdff dff_A_Kq47wWt17_0(.dout(w_dff_A_cBTUSIlK9_0),.din(w_dff_A_Kq47wWt17_0),.clk(gclk));
	jdff dff_A_cgE24JCS8_0(.dout(w_dff_A_Kq47wWt17_0),.din(w_dff_A_cgE24JCS8_0),.clk(gclk));
	jdff dff_A_IJB7r4Tb8_0(.dout(w_dff_A_cgE24JCS8_0),.din(w_dff_A_IJB7r4Tb8_0),.clk(gclk));
	jdff dff_A_3LWJ42QH3_0(.dout(w_dff_A_IJB7r4Tb8_0),.din(w_dff_A_3LWJ42QH3_0),.clk(gclk));
	jdff dff_A_QIPZdZ9U2_0(.dout(w_dff_A_3LWJ42QH3_0),.din(w_dff_A_QIPZdZ9U2_0),.clk(gclk));
	jdff dff_A_0YIluyBg5_2(.dout(w_G1497_0[2]),.din(w_dff_A_0YIluyBg5_2),.clk(gclk));
	jdff dff_A_x5RSzLg95_2(.dout(w_dff_A_0YIluyBg5_2),.din(w_dff_A_x5RSzLg95_2),.clk(gclk));
	jdff dff_A_KlZqlUxc6_2(.dout(w_dff_A_x5RSzLg95_2),.din(w_dff_A_KlZqlUxc6_2),.clk(gclk));
	jdff dff_A_tjtZVJ2u2_2(.dout(w_dff_A_KlZqlUxc6_2),.din(w_dff_A_tjtZVJ2u2_2),.clk(gclk));
	jdff dff_A_1N9g9ILt1_2(.dout(w_dff_A_tjtZVJ2u2_2),.din(w_dff_A_1N9g9ILt1_2),.clk(gclk));
	jdff dff_A_UwO2FDe47_2(.dout(w_dff_A_1N9g9ILt1_2),.din(w_dff_A_UwO2FDe47_2),.clk(gclk));
	jdff dff_A_0kENtmZp5_2(.dout(w_dff_A_UwO2FDe47_2),.din(w_dff_A_0kENtmZp5_2),.clk(gclk));
	jdff dff_A_017YlmjG8_2(.dout(w_dff_A_0kENtmZp5_2),.din(w_dff_A_017YlmjG8_2),.clk(gclk));
	jdff dff_A_GzSCvmyJ9_2(.dout(w_dff_A_017YlmjG8_2),.din(w_dff_A_GzSCvmyJ9_2),.clk(gclk));
	jdff dff_A_gmdSfpsv8_2(.dout(w_dff_A_GzSCvmyJ9_2),.din(w_dff_A_gmdSfpsv8_2),.clk(gclk));
	jdff dff_B_FboPHIRO5_1(.din(n675),.dout(w_dff_B_FboPHIRO5_1),.clk(gclk));
	jdff dff_B_RUghDjnJ6_1(.din(w_dff_B_FboPHIRO5_1),.dout(w_dff_B_RUghDjnJ6_1),.clk(gclk));
	jdff dff_B_hrQg93Qp0_1(.din(w_dff_B_RUghDjnJ6_1),.dout(w_dff_B_hrQg93Qp0_1),.clk(gclk));
	jdff dff_B_15CS6bYn4_1(.din(w_dff_B_hrQg93Qp0_1),.dout(w_dff_B_15CS6bYn4_1),.clk(gclk));
	jdff dff_B_T1NSR8jE9_1(.din(n676),.dout(w_dff_B_T1NSR8jE9_1),.clk(gclk));
	jdff dff_B_iF0KyPtM9_1(.din(w_dff_B_T1NSR8jE9_1),.dout(w_dff_B_iF0KyPtM9_1),.clk(gclk));
	jdff dff_B_tgCupd6O2_1(.din(w_dff_B_iF0KyPtM9_1),.dout(w_dff_B_tgCupd6O2_1),.clk(gclk));
	jdff dff_B_2VIl7vl08_1(.din(w_dff_B_tgCupd6O2_1),.dout(w_dff_B_2VIl7vl08_1),.clk(gclk));
	jdff dff_B_Uc3tdeoM0_1(.din(w_dff_B_2VIl7vl08_1),.dout(w_dff_B_Uc3tdeoM0_1),.clk(gclk));
	jdff dff_A_YAqQIAnL3_1(.dout(w_n691_0[1]),.din(w_dff_A_YAqQIAnL3_1),.clk(gclk));
	jdff dff_A_evSASmTu6_0(.dout(w_n689_0[0]),.din(w_dff_A_evSASmTu6_0),.clk(gclk));
	jdff dff_A_kGXM6RqT9_0(.dout(w_n687_0[0]),.din(w_dff_A_kGXM6RqT9_0),.clk(gclk));
	jdff dff_A_yuFEVChI9_1(.dout(w_n687_0[1]),.din(w_dff_A_yuFEVChI9_1),.clk(gclk));
	jdff dff_A_7pXUF9fR4_1(.dout(w_dff_A_yuFEVChI9_1),.din(w_dff_A_7pXUF9fR4_1),.clk(gclk));
	jdff dff_A_Plj7rlTI0_1(.dout(w_dff_A_7pXUF9fR4_1),.din(w_dff_A_Plj7rlTI0_1),.clk(gclk));
	jdff dff_A_qDDp2ip11_1(.dout(w_dff_A_Plj7rlTI0_1),.din(w_dff_A_qDDp2ip11_1),.clk(gclk));
	jdff dff_A_5IIaAJoR1_2(.dout(w_n571_0[2]),.din(w_dff_A_5IIaAJoR1_2),.clk(gclk));
	jdff dff_A_SRrG980J0_2(.dout(w_dff_A_5IIaAJoR1_2),.din(w_dff_A_SRrG980J0_2),.clk(gclk));
	jdff dff_A_gTlyjfpT1_2(.dout(w_dff_A_SRrG980J0_2),.din(w_dff_A_gTlyjfpT1_2),.clk(gclk));
	jdff dff_A_z8mKH3gn7_1(.dout(w_n569_0[1]),.din(w_dff_A_z8mKH3gn7_1),.clk(gclk));
	jdff dff_A_m1AaSk9P7_1(.dout(w_G280_0[1]),.din(w_dff_A_m1AaSk9P7_1),.clk(gclk));
	jdff dff_A_OkQ4V4ul0_0(.dout(w_n486_1[0]),.din(w_dff_A_OkQ4V4ul0_0),.clk(gclk));
	jdff dff_A_nMug4MFz8_0(.dout(w_n681_2[0]),.din(w_dff_A_nMug4MFz8_0),.clk(gclk));
	jdff dff_A_aNeRiGDk3_0(.dout(w_dff_A_nMug4MFz8_0),.din(w_dff_A_aNeRiGDk3_0),.clk(gclk));
	jdff dff_A_Q8688C4e3_1(.dout(w_n680_0[1]),.din(w_dff_A_Q8688C4e3_1),.clk(gclk));
	jdff dff_B_n06xFyHa9_2(.din(n680),.dout(w_dff_B_n06xFyHa9_2),.clk(gclk));
	jdff dff_A_quGm9qOq7_0(.dout(w_n451_1[0]),.din(w_dff_A_quGm9qOq7_0),.clk(gclk));
	jdff dff_A_R7x0xSWu1_1(.dout(w_n679_0[1]),.din(w_dff_A_R7x0xSWu1_1),.clk(gclk));
	jdff dff_A_y24sHRf73_1(.dout(w_dff_A_R7x0xSWu1_1),.din(w_dff_A_y24sHRf73_1),.clk(gclk));
	jdff dff_A_vDwub33C8_1(.dout(w_n678_0[1]),.din(w_dff_A_vDwub33C8_1),.clk(gclk));
	jdff dff_A_mMhdil6U0_1(.dout(w_dff_A_vDwub33C8_1),.din(w_dff_A_mMhdil6U0_1),.clk(gclk));
	jdff dff_A_AHYVuzOx6_1(.dout(w_dff_A_mMhdil6U0_1),.din(w_dff_A_AHYVuzOx6_1),.clk(gclk));
	jdff dff_B_sgRjECoX8_1(.din(n557),.dout(w_dff_B_sgRjECoX8_1),.clk(gclk));
	jdff dff_B_XMxOAZNd4_1(.din(G241),.dout(w_dff_B_XMxOAZNd4_1),.clk(gclk));
	jdff dff_B_udTWXWny9_2(.din(n1543),.dout(w_dff_B_udTWXWny9_2),.clk(gclk));
	jdff dff_B_UtgxsUNu9_2(.din(w_dff_B_udTWXWny9_2),.dout(w_dff_B_UtgxsUNu9_2),.clk(gclk));
	jdff dff_B_JPFUb9cB6_2(.din(w_dff_B_UtgxsUNu9_2),.dout(w_dff_B_JPFUb9cB6_2),.clk(gclk));
	jdff dff_B_tFhesDRj6_2(.din(w_dff_B_JPFUb9cB6_2),.dout(w_dff_B_tFhesDRj6_2),.clk(gclk));
	jdff dff_B_L9ZMFgnB6_2(.din(w_dff_B_tFhesDRj6_2),.dout(w_dff_B_L9ZMFgnB6_2),.clk(gclk));
	jdff dff_B_1pShMc1D2_2(.din(w_dff_B_L9ZMFgnB6_2),.dout(w_dff_B_1pShMc1D2_2),.clk(gclk));
	jdff dff_B_Dkqd5guL7_2(.din(w_dff_B_1pShMc1D2_2),.dout(w_dff_B_Dkqd5guL7_2),.clk(gclk));
	jdff dff_B_WknH7xHK3_2(.din(w_dff_B_Dkqd5guL7_2),.dout(w_dff_B_WknH7xHK3_2),.clk(gclk));
	jdff dff_B_Fg5lBWpv4_2(.din(w_dff_B_WknH7xHK3_2),.dout(w_dff_B_Fg5lBWpv4_2),.clk(gclk));
	jdff dff_B_kuwmshAL9_2(.din(w_dff_B_Fg5lBWpv4_2),.dout(w_dff_B_kuwmshAL9_2),.clk(gclk));
	jdff dff_A_Ysk3cZVl4_2(.dout(w_n583_0[2]),.din(w_dff_A_Ysk3cZVl4_2),.clk(gclk));
	jdff dff_A_dm6gyHFT9_2(.dout(w_dff_A_Ysk3cZVl4_2),.din(w_dff_A_dm6gyHFT9_2),.clk(gclk));
	jdff dff_A_TDrrSPXo7_2(.dout(w_dff_A_dm6gyHFT9_2),.din(w_dff_A_TDrrSPXo7_2),.clk(gclk));
	jdff dff_A_FskTuqoE1_2(.dout(w_dff_A_TDrrSPXo7_2),.din(w_dff_A_FskTuqoE1_2),.clk(gclk));
	jdff dff_A_legCigtL3_2(.dout(w_dff_A_FskTuqoE1_2),.din(w_dff_A_legCigtL3_2),.clk(gclk));
	jdff dff_A_gyPtAf1f2_1(.dout(w_n578_0[1]),.din(w_dff_A_gyPtAf1f2_1),.clk(gclk));
	jdff dff_A_Ssov5t7J6_1(.dout(w_dff_A_gyPtAf1f2_1),.din(w_dff_A_Ssov5t7J6_1),.clk(gclk));
	jdff dff_A_JScAPa3A8_1(.dout(w_dff_A_Ssov5t7J6_1),.din(w_dff_A_JScAPa3A8_1),.clk(gclk));
	jdff dff_A_HJZTXVlc5_1(.dout(w_dff_A_JScAPa3A8_1),.din(w_dff_A_HJZTXVlc5_1),.clk(gclk));
	jdff dff_A_5fld2Bhh1_1(.dout(w_dff_A_HJZTXVlc5_1),.din(w_dff_A_5fld2Bhh1_1),.clk(gclk));
	jdff dff_A_dkZK43yW7_1(.dout(w_dff_A_5fld2Bhh1_1),.din(w_dff_A_dkZK43yW7_1),.clk(gclk));
	jdff dff_A_H8aPmCPQ7_1(.dout(w_dff_A_dkZK43yW7_1),.din(w_dff_A_H8aPmCPQ7_1),.clk(gclk));
	jdff dff_B_SyGdP9t01_0(.din(n576),.dout(w_dff_B_SyGdP9t01_0),.clk(gclk));
	jdff dff_A_MVqbkzH00_0(.dout(w_G335_3[0]),.din(w_dff_A_MVqbkzH00_0),.clk(gclk));
	jdff dff_B_zXsy4sDE9_1(.din(G264),.dout(w_dff_B_zXsy4sDE9_1),.clk(gclk));
	jdff dff_A_E2vqs1Gz9_0(.dout(w_n473_1[0]),.din(w_dff_A_E2vqs1Gz9_0),.clk(gclk));
	jdff dff_A_Rx7my7XR1_0(.dout(w_dff_A_E2vqs1Gz9_0),.din(w_dff_A_Rx7my7XR1_0),.clk(gclk));
	jdff dff_A_F72lr6t99_1(.dout(w_n473_1[1]),.din(w_dff_A_F72lr6t99_1),.clk(gclk));
	jdff dff_A_OYI0EwiM0_1(.dout(w_n943_0[1]),.din(w_dff_A_OYI0EwiM0_1),.clk(gclk));
	jdff dff_A_SVbnN9s24_1(.dout(w_dff_A_OYI0EwiM0_1),.din(w_dff_A_SVbnN9s24_1),.clk(gclk));
	jdff dff_A_TlknoW6D7_1(.dout(w_dff_A_SVbnN9s24_1),.din(w_dff_A_TlknoW6D7_1),.clk(gclk));
	jdff dff_A_EmzmYA7F1_1(.dout(w_dff_A_TlknoW6D7_1),.din(w_dff_A_EmzmYA7F1_1),.clk(gclk));
	jdff dff_A_IsFo5hR41_1(.dout(w_dff_A_EmzmYA7F1_1),.din(w_dff_A_IsFo5hR41_1),.clk(gclk));
	jdff dff_A_FS1dtY4e7_1(.dout(w_dff_A_IsFo5hR41_1),.din(w_dff_A_FS1dtY4e7_1),.clk(gclk));
	jdff dff_A_bKObz1oh2_1(.dout(w_dff_A_FS1dtY4e7_1),.din(w_dff_A_bKObz1oh2_1),.clk(gclk));
	jdff dff_A_qdG8UMs30_1(.dout(w_dff_A_bKObz1oh2_1),.din(w_dff_A_qdG8UMs30_1),.clk(gclk));
	jdff dff_A_tTROXtQE4_1(.dout(w_dff_A_qdG8UMs30_1),.din(w_dff_A_tTROXtQE4_1),.clk(gclk));
	jdff dff_A_VaI15jXt6_1(.dout(w_dff_A_tTROXtQE4_1),.din(w_dff_A_VaI15jXt6_1),.clk(gclk));
	jdff dff_A_irDksPBB8_1(.dout(w_dff_A_VaI15jXt6_1),.din(w_dff_A_irDksPBB8_1),.clk(gclk));
	jdff dff_A_QjppZzxw4_1(.dout(w_dff_A_irDksPBB8_1),.din(w_dff_A_QjppZzxw4_1),.clk(gclk));
	jdff dff_A_2NXqZb9L5_1(.dout(w_n591_0[1]),.din(w_dff_A_2NXqZb9L5_1),.clk(gclk));
	jdff dff_A_0Rqlm6JO6_1(.dout(w_n590_0[1]),.din(w_dff_A_0Rqlm6JO6_1),.clk(gclk));
	jdff dff_A_BIFyI2Ba4_1(.dout(w_dff_A_0Rqlm6JO6_1),.din(w_dff_A_BIFyI2Ba4_1),.clk(gclk));
	jdff dff_B_jK6rhq0e3_0(.din(n589),.dout(w_dff_B_jK6rhq0e3_0),.clk(gclk));
	jdff dff_B_gwnaqesO9_1(.din(G217),.dout(w_dff_B_gwnaqesO9_1),.clk(gclk));
	jdff dff_A_f7lUCiew2_0(.dout(w_G335_4[0]),.din(w_dff_A_f7lUCiew2_0),.clk(gclk));
	jdff dff_A_giWd21D36_2(.dout(w_G335_1[2]),.din(w_dff_A_giWd21D36_2),.clk(gclk));
	jdff dff_A_8oKXciT03_1(.dout(w_n750_0[1]),.din(w_dff_A_8oKXciT03_1),.clk(gclk));
	jdff dff_A_T5WUaTeX7_1(.dout(w_dff_A_8oKXciT03_1),.din(w_dff_A_T5WUaTeX7_1),.clk(gclk));
	jdff dff_A_rqE1AeFv5_1(.dout(w_dff_A_T5WUaTeX7_1),.din(w_dff_A_rqE1AeFv5_1),.clk(gclk));
	jdff dff_A_J7TlupEE3_1(.dout(w_dff_A_rqE1AeFv5_1),.din(w_dff_A_J7TlupEE3_1),.clk(gclk));
	jdff dff_A_vyzf7wGv7_1(.dout(w_dff_A_J7TlupEE3_1),.din(w_dff_A_vyzf7wGv7_1),.clk(gclk));
	jdff dff_A_aW4fAWQe5_1(.dout(w_dff_A_vyzf7wGv7_1),.din(w_dff_A_aW4fAWQe5_1),.clk(gclk));
	jdff dff_A_8AIJ25oZ5_1(.dout(w_dff_A_aW4fAWQe5_1),.din(w_dff_A_8AIJ25oZ5_1),.clk(gclk));
	jdff dff_A_5Q8c7W6x3_1(.dout(w_dff_A_8AIJ25oZ5_1),.din(w_dff_A_5Q8c7W6x3_1),.clk(gclk));
	jdff dff_A_PWdd2DEy6_1(.dout(w_dff_A_5Q8c7W6x3_1),.din(w_dff_A_PWdd2DEy6_1),.clk(gclk));
	jdff dff_A_8PrYpk353_1(.dout(w_dff_A_PWdd2DEy6_1),.din(w_dff_A_8PrYpk353_1),.clk(gclk));
	jdff dff_A_S5lETVX55_1(.dout(w_dff_A_8PrYpk353_1),.din(w_dff_A_S5lETVX55_1),.clk(gclk));
	jdff dff_A_fiYCsWVX3_1(.dout(w_dff_A_S5lETVX55_1),.din(w_dff_A_fiYCsWVX3_1),.clk(gclk));
	jdff dff_A_s7dU7DEJ4_1(.dout(w_dff_A_fiYCsWVX3_1),.din(w_dff_A_s7dU7DEJ4_1),.clk(gclk));
	jdff dff_A_hQMLIAPg0_1(.dout(w_dff_A_s7dU7DEJ4_1),.din(w_dff_A_hQMLIAPg0_1),.clk(gclk));
	jdff dff_A_Xrkgt8Uq2_1(.dout(w_dff_A_hQMLIAPg0_1),.din(w_dff_A_Xrkgt8Uq2_1),.clk(gclk));
	jdff dff_A_QzXpiAQL1_1(.dout(w_dff_A_Xrkgt8Uq2_1),.din(w_dff_A_QzXpiAQL1_1),.clk(gclk));
	jdff dff_A_UfmvrRkC4_1(.dout(w_dff_A_QzXpiAQL1_1),.din(w_dff_A_UfmvrRkC4_1),.clk(gclk));
	jdff dff_A_hzxSu0t47_2(.dout(w_n750_0[2]),.din(w_dff_A_hzxSu0t47_2),.clk(gclk));
	jdff dff_A_PlNFSRZF0_2(.dout(w_dff_A_hzxSu0t47_2),.din(w_dff_A_PlNFSRZF0_2),.clk(gclk));
	jdff dff_A_WB2Uv4N09_2(.dout(w_dff_A_PlNFSRZF0_2),.din(w_dff_A_WB2Uv4N09_2),.clk(gclk));
	jdff dff_A_QuvMuqkL5_2(.dout(w_dff_A_WB2Uv4N09_2),.din(w_dff_A_QuvMuqkL5_2),.clk(gclk));
	jdff dff_A_pEF531yR7_2(.dout(w_dff_A_QuvMuqkL5_2),.din(w_dff_A_pEF531yR7_2),.clk(gclk));
	jdff dff_A_2Iy5PONt3_2(.dout(w_dff_A_pEF531yR7_2),.din(w_dff_A_2Iy5PONt3_2),.clk(gclk));
	jdff dff_A_v0uVrX126_2(.dout(w_dff_A_2Iy5PONt3_2),.din(w_dff_A_v0uVrX126_2),.clk(gclk));
	jdff dff_A_JuSmpmgD2_2(.dout(w_dff_A_v0uVrX126_2),.din(w_dff_A_JuSmpmgD2_2),.clk(gclk));
	jdff dff_A_HsNOgYfh5_2(.dout(w_G4091_2[2]),.din(w_dff_A_HsNOgYfh5_2),.clk(gclk));
	jdff dff_A_xthy18NE9_2(.dout(w_G4091_0[2]),.din(w_dff_A_xthy18NE9_2),.clk(gclk));
	jdff dff_A_t40zNYXZ9_2(.dout(w_dff_A_xthy18NE9_2),.din(w_dff_A_t40zNYXZ9_2),.clk(gclk));
	jdff dff_A_nQRxAP3K2_2(.dout(w_dff_A_t40zNYXZ9_2),.din(w_dff_A_nQRxAP3K2_2),.clk(gclk));
	jdff dff_A_K5oSnFpI3_2(.dout(w_dff_A_nQRxAP3K2_2),.din(w_dff_A_K5oSnFpI3_2),.clk(gclk));
	jdff dff_A_zpJyU6uJ7_2(.dout(w_dff_A_K5oSnFpI3_2),.din(w_dff_A_zpJyU6uJ7_2),.clk(gclk));
	jdff dff_A_GZprBdzv7_2(.dout(w_dff_A_zpJyU6uJ7_2),.din(w_dff_A_GZprBdzv7_2),.clk(gclk));
	jdff dff_A_EfOBnjDB0_2(.dout(w_dff_A_GZprBdzv7_2),.din(w_dff_A_EfOBnjDB0_2),.clk(gclk));
	jdff dff_A_Zs4y31Dq2_2(.dout(w_dff_A_EfOBnjDB0_2),.din(w_dff_A_Zs4y31Dq2_2),.clk(gclk));
	jdff dff_A_zg1pibig3_2(.dout(w_dff_A_Zs4y31Dq2_2),.din(w_dff_A_zg1pibig3_2),.clk(gclk));
	jdff dff_A_3geM0Cms6_2(.dout(w_dff_A_zg1pibig3_2),.din(w_dff_A_3geM0Cms6_2),.clk(gclk));
	jdff dff_A_txTqEs2L8_2(.dout(w_dff_A_3geM0Cms6_2),.din(w_dff_A_txTqEs2L8_2),.clk(gclk));
	jdff dff_A_HGT1TjPl5_2(.dout(w_dff_A_txTqEs2L8_2),.din(w_dff_A_HGT1TjPl5_2),.clk(gclk));
	jdff dff_A_1RahILR75_2(.dout(w_dff_A_HGT1TjPl5_2),.din(w_dff_A_1RahILR75_2),.clk(gclk));
	jdff dff_A_yg7oj4gc8_2(.dout(w_dff_A_1RahILR75_2),.din(w_dff_A_yg7oj4gc8_2),.clk(gclk));
	jdff dff_A_7NfPz0Xh7_2(.dout(w_dff_A_yg7oj4gc8_2),.din(w_dff_A_7NfPz0Xh7_2),.clk(gclk));
	jdff dff_A_DaipWDjI3_2(.dout(w_dff_A_7NfPz0Xh7_2),.din(w_dff_A_DaipWDjI3_2),.clk(gclk));
	jdff dff_A_2isySGdC3_2(.dout(w_dff_A_DaipWDjI3_2),.din(w_dff_A_2isySGdC3_2),.clk(gclk));
	jdff dff_A_4XKB28U33_2(.dout(w_dff_A_2isySGdC3_2),.din(w_dff_A_4XKB28U33_2),.clk(gclk));
	jdff dff_B_tFWjCfY76_2(.din(n1533),.dout(w_dff_B_tFWjCfY76_2),.clk(gclk));
	jdff dff_B_ypoCYK9M4_1(.din(n1526),.dout(w_dff_B_ypoCYK9M4_1),.clk(gclk));
	jdff dff_B_9VCie3KC0_1(.din(n1527),.dout(w_dff_B_9VCie3KC0_1),.clk(gclk));
	jdff dff_A_W71XNuJJ0_0(.dout(w_n486_0[0]),.din(w_dff_A_W71XNuJJ0_0),.clk(gclk));
	jdff dff_A_RIOyuKSd2_2(.dout(w_n486_0[2]),.din(w_dff_A_RIOyuKSd2_2),.clk(gclk));
	jdff dff_A_AYrARYnc4_2(.dout(w_dff_A_RIOyuKSd2_2),.din(w_dff_A_AYrARYnc4_2),.clk(gclk));
	jdff dff_A_tpZMpNCi1_0(.dout(w_G411_0[0]),.din(w_dff_A_tpZMpNCi1_0),.clk(gclk));
	jdff dff_A_IBV2KcPm6_0(.dout(w_dff_A_tpZMpNCi1_0),.din(w_dff_A_IBV2KcPm6_0),.clk(gclk));
	jdff dff_A_KdrmsbCd1_1(.dout(w_G411_0[1]),.din(w_dff_A_KdrmsbCd1_1),.clk(gclk));
	jdff dff_A_k47UJfMu3_1(.dout(w_G273_2[1]),.din(w_dff_A_k47UJfMu3_1),.clk(gclk));
	jdff dff_A_LzTv22fS0_2(.dout(w_G273_0[2]),.din(w_dff_A_LzTv22fS0_2),.clk(gclk));
	jdff dff_B_3IdeH9Np3_1(.din(n1518),.dout(w_dff_B_3IdeH9Np3_1),.clk(gclk));
	jdff dff_B_acLe9BB14_1(.din(w_dff_B_3IdeH9Np3_1),.dout(w_dff_B_acLe9BB14_1),.clk(gclk));
	jdff dff_A_BuHAXN7I3_2(.dout(w_n473_0[2]),.din(w_dff_A_BuHAXN7I3_2),.clk(gclk));
	jdff dff_A_cR87xW9l6_2(.dout(w_dff_A_BuHAXN7I3_2),.din(w_dff_A_cR87xW9l6_2),.clk(gclk));
	jdff dff_B_9tSn0Y3k1_3(.din(n473),.dout(w_dff_B_9tSn0Y3k1_3),.clk(gclk));
	jdff dff_B_hmWGLqJC7_1(.din(n1514),.dout(w_dff_B_hmWGLqJC7_1),.clk(gclk));
	jdff dff_A_AHWfAdJj2_1(.dout(w_G257_2[1]),.din(w_dff_A_AHWfAdJj2_1),.clk(gclk));
	jdff dff_A_EXVkxyFG1_0(.dout(w_G389_0[0]),.din(w_dff_A_EXVkxyFG1_0),.clk(gclk));
	jdff dff_A_8QLBYNJY8_0(.dout(w_dff_A_EXVkxyFG1_0),.din(w_dff_A_8QLBYNJY8_0),.clk(gclk));
	jdff dff_A_emFgZITx2_1(.dout(w_G389_0[1]),.din(w_dff_A_emFgZITx2_1),.clk(gclk));
	jdff dff_A_WQTppcFP4_0(.dout(w_G257_1[0]),.din(w_dff_A_WQTppcFP4_0),.clk(gclk));
	jdff dff_B_FBmqfDmr8_1(.din(n1507),.dout(w_dff_B_FBmqfDmr8_1),.clk(gclk));
	jdff dff_B_MuDZpq9d7_1(.din(n1508),.dout(w_dff_B_MuDZpq9d7_1),.clk(gclk));
	jdff dff_A_XBsqqt4V8_0(.dout(w_n451_0[0]),.din(w_dff_A_XBsqqt4V8_0),.clk(gclk));
	jdff dff_A_g7GwuWCI6_2(.dout(w_n451_0[2]),.din(w_dff_A_g7GwuWCI6_2),.clk(gclk));
	jdff dff_A_KKnWbrl30_2(.dout(w_dff_A_g7GwuWCI6_2),.din(w_dff_A_KKnWbrl30_2),.clk(gclk));
	jdff dff_A_epP7q5ez9_0(.dout(w_G400_1[0]),.din(w_dff_A_epP7q5ez9_0),.clk(gclk));
	jdff dff_A_GiVZV48h2_1(.dout(w_G400_0[1]),.din(w_dff_A_GiVZV48h2_1),.clk(gclk));
	jdff dff_A_3gDDM7YM7_1(.dout(w_dff_A_GiVZV48h2_1),.din(w_dff_A_3gDDM7YM7_1),.clk(gclk));
	jdff dff_A_2BKmGxKs5_2(.dout(w_G400_0[2]),.din(w_dff_A_2BKmGxKs5_2),.clk(gclk));
	jdff dff_A_tgC1v8gX3_2(.dout(w_dff_A_2BKmGxKs5_2),.din(w_dff_A_tgC1v8gX3_2),.clk(gclk));
	jdff dff_A_6TXoc7rK1_2(.dout(w_dff_A_tgC1v8gX3_2),.din(w_dff_A_6TXoc7rK1_2),.clk(gclk));
	jdff dff_A_Nvzu5XCg3_0(.dout(w_G265_2[0]),.din(w_dff_A_Nvzu5XCg3_0),.clk(gclk));
	jdff dff_A_VmEvoykn8_2(.dout(w_G265_0[2]),.din(w_dff_A_VmEvoykn8_2),.clk(gclk));
	jdff dff_B_TnDCwe8l9_1(.din(n1498),.dout(w_dff_B_TnDCwe8l9_1),.clk(gclk));
	jdff dff_B_0XVfhXz86_1(.din(n1499),.dout(w_dff_B_0XVfhXz86_1),.clk(gclk));
	jdff dff_A_hcaBnGNJ4_0(.dout(w_n497_0[0]),.din(w_dff_A_hcaBnGNJ4_0),.clk(gclk));
	jdff dff_A_dkRzf9Fo3_2(.dout(w_n497_0[2]),.din(w_dff_A_dkRzf9Fo3_2),.clk(gclk));
	jdff dff_A_aL3GOddb6_2(.dout(w_dff_A_dkRzf9Fo3_2),.din(w_dff_A_aL3GOddb6_2),.clk(gclk));
	jdff dff_A_6NnZ85746_0(.dout(w_G374_0[0]),.din(w_dff_A_6NnZ85746_0),.clk(gclk));
	jdff dff_A_uzHU8Ycj9_0(.dout(w_dff_A_6NnZ85746_0),.din(w_dff_A_uzHU8Ycj9_0),.clk(gclk));
	jdff dff_A_zxoV718G2_1(.dout(w_G374_0[1]),.din(w_dff_A_zxoV718G2_1),.clk(gclk));
	jdff dff_A_5f3YffZc9_0(.dout(w_G281_2[0]),.din(w_dff_A_5f3YffZc9_0),.clk(gclk));
	jdff dff_A_i4yijk0O8_2(.dout(w_G281_0[2]),.din(w_dff_A_i4yijk0O8_2),.clk(gclk));
	jdff dff_B_1P3BHLgR7_1(.din(n1463),.dout(w_dff_B_1P3BHLgR7_1),.clk(gclk));
	jdff dff_B_RzIglBOu5_1(.din(w_dff_B_1P3BHLgR7_1),.dout(w_dff_B_RzIglBOu5_1),.clk(gclk));
	jdff dff_B_9WJTBuJM3_1(.din(n1486),.dout(w_dff_B_9WJTBuJM3_1),.clk(gclk));
	jdff dff_B_Dbht9dBE8_1(.din(n1487),.dout(w_dff_B_Dbht9dBE8_1),.clk(gclk));
	jdff dff_A_EizV1JxL4_1(.dout(w_G210_1[1]),.din(w_dff_A_EizV1JxL4_1),.clk(gclk));
	jdff dff_A_cjga727m6_1(.dout(w_n543_0[1]),.din(w_dff_A_cjga727m6_1),.clk(gclk));
	jdff dff_A_DSYuGwNq6_0(.dout(w_G457_2[0]),.din(w_dff_A_DSYuGwNq6_0),.clk(gclk));
	jdff dff_A_utIED0WE2_0(.dout(w_G457_0[0]),.din(w_dff_A_utIED0WE2_0),.clk(gclk));
	jdff dff_A_yQ2rIpMw1_0(.dout(w_dff_A_utIED0WE2_0),.din(w_dff_A_yQ2rIpMw1_0),.clk(gclk));
	jdff dff_A_sWDiBuh02_0(.dout(w_dff_A_yQ2rIpMw1_0),.din(w_dff_A_sWDiBuh02_0),.clk(gclk));
	jdff dff_A_JUV4H6lN0_2(.dout(w_G457_0[2]),.din(w_dff_A_JUV4H6lN0_2),.clk(gclk));
	jdff dff_A_siA6kNFd3_2(.dout(w_dff_A_JUV4H6lN0_2),.din(w_dff_A_siA6kNFd3_2),.clk(gclk));
	jdff dff_A_TRyHePPu3_1(.dout(w_G210_2[1]),.din(w_dff_A_TRyHePPu3_1),.clk(gclk));
	jdff dff_A_UBKQ6Prb5_2(.dout(w_G210_0[2]),.din(w_dff_A_UBKQ6Prb5_2),.clk(gclk));
	jdff dff_B_VwSpmpmP0_1(.din(n1478),.dout(w_dff_B_VwSpmpmP0_1),.clk(gclk));
	jdff dff_B_ft2Gh3C70_1(.din(w_dff_B_VwSpmpmP0_1),.dout(w_dff_B_ft2Gh3C70_1),.clk(gclk));
	jdff dff_B_nQshTVjR8_2(.din(n509),.dout(w_dff_B_nQshTVjR8_2),.clk(gclk));
	jdff dff_A_Rg98vPlY4_0(.dout(w_G468_1[0]),.din(w_dff_A_Rg98vPlY4_0),.clk(gclk));
	jdff dff_A_vZnYrOku2_0(.dout(w_dff_A_Rg98vPlY4_0),.din(w_dff_A_vZnYrOku2_0),.clk(gclk));
	jdff dff_A_zPwGSvjv5_0(.dout(w_dff_A_vZnYrOku2_0),.din(w_dff_A_zPwGSvjv5_0),.clk(gclk));
	jdff dff_A_ePZeCHJY0_1(.dout(w_G468_1[1]),.din(w_dff_A_ePZeCHJY0_1),.clk(gclk));
	jdff dff_B_nEin9Box4_1(.din(n1474),.dout(w_dff_B_nEin9Box4_1),.clk(gclk));
	jdff dff_A_5rnoyF4a9_1(.dout(w_G218_2[1]),.din(w_dff_A_5rnoyF4a9_1),.clk(gclk));
	jdff dff_A_BKcFDSnW7_1(.dout(w_G468_0[1]),.din(w_dff_A_BKcFDSnW7_1),.clk(gclk));
	jdff dff_A_gU7880GW8_1(.dout(w_dff_A_BKcFDSnW7_1),.din(w_dff_A_gU7880GW8_1),.clk(gclk));
	jdff dff_A_3ddKH4RU8_2(.dout(w_G468_0[2]),.din(w_dff_A_3ddKH4RU8_2),.clk(gclk));
	jdff dff_A_EqCpre9Y7_2(.dout(w_dff_A_3ddKH4RU8_2),.din(w_dff_A_EqCpre9Y7_2),.clk(gclk));
	jdff dff_A_F12oIkZY4_2(.dout(w_dff_A_EqCpre9Y7_2),.din(w_dff_A_F12oIkZY4_2),.clk(gclk));
	jdff dff_A_7sPGyeUk4_0(.dout(w_G218_1[0]),.din(w_dff_A_7sPGyeUk4_0),.clk(gclk));
	jdff dff_B_XAClLi7a5_1(.din(n1468),.dout(w_dff_B_XAClLi7a5_1),.clk(gclk));
	jdff dff_B_ObJKJAL65_1(.din(w_dff_B_XAClLi7a5_1),.dout(w_dff_B_ObJKJAL65_1),.clk(gclk));
	jdff dff_B_VElSIzjE4_2(.din(n532),.dout(w_dff_B_VElSIzjE4_2),.clk(gclk));
	jdff dff_A_3BiR3btB8_0(.dout(w_G422_2[0]),.din(w_dff_A_3BiR3btB8_0),.clk(gclk));
	jdff dff_B_bhkwObJ23_1(.din(n1464),.dout(w_dff_B_bhkwObJ23_1),.clk(gclk));
	jdff dff_A_uazgisl77_1(.dout(w_G226_2[1]),.din(w_dff_A_uazgisl77_1),.clk(gclk));
	jdff dff_A_hmoDB3ZB7_0(.dout(w_G422_0[0]),.din(w_dff_A_hmoDB3ZB7_0),.clk(gclk));
	jdff dff_A_XJZbC1zp8_0(.dout(w_dff_A_hmoDB3ZB7_0),.din(w_dff_A_XJZbC1zp8_0),.clk(gclk));
	jdff dff_A_u7SX3Bg06_0(.dout(w_dff_A_XJZbC1zp8_0),.din(w_dff_A_u7SX3Bg06_0),.clk(gclk));
	jdff dff_A_VwRRsoqh0_2(.dout(w_G422_0[2]),.din(w_dff_A_VwRRsoqh0_2),.clk(gclk));
	jdff dff_A_3mpWkusM1_2(.dout(w_dff_A_VwRRsoqh0_2),.din(w_dff_A_3mpWkusM1_2),.clk(gclk));
	jdff dff_A_FkEO5EKi9_1(.dout(w_G251_4[1]),.din(w_dff_A_FkEO5EKi9_1),.clk(gclk));
	jdff dff_A_8ErAXYhy7_2(.dout(w_G251_4[2]),.din(w_dff_A_8ErAXYhy7_2),.clk(gclk));
	jdff dff_A_oh0mZN6n0_1(.dout(w_G251_1[1]),.din(w_dff_A_oh0mZN6n0_1),.clk(gclk));
	jdff dff_A_UvE4980e5_2(.dout(w_G251_1[2]),.din(w_dff_A_UvE4980e5_2),.clk(gclk));
	jdff dff_A_UIM1XxVP6_0(.dout(w_G226_1[0]),.din(w_dff_A_UIM1XxVP6_0),.clk(gclk));
	jdff dff_B_mmaQjxYO6_1(.din(n523),.dout(w_dff_B_mmaQjxYO6_1),.clk(gclk));
	jdff dff_B_Vte1rW7f8_1(.din(n524),.dout(w_dff_B_Vte1rW7f8_1),.clk(gclk));
	jdff dff_A_vBnwzuFg4_0(.dout(w_G446_1[0]),.din(w_dff_A_vBnwzuFg4_0),.clk(gclk));
	jdff dff_A_gbBNtmKH0_0(.dout(w_dff_A_vBnwzuFg4_0),.din(w_dff_A_gbBNtmKH0_0),.clk(gclk));
	jdff dff_A_etOclqIw0_0(.dout(w_dff_A_gbBNtmKH0_0),.din(w_dff_A_etOclqIw0_0),.clk(gclk));
	jdff dff_A_YeycLRNs9_0(.dout(w_dff_A_etOclqIw0_0),.din(w_dff_A_YeycLRNs9_0),.clk(gclk));
	jdff dff_A_sl8a1jJF6_1(.dout(w_G446_1[1]),.din(w_dff_A_sl8a1jJF6_1),.clk(gclk));
	jdff dff_A_5acy51VL2_1(.dout(w_dff_A_sl8a1jJF6_1),.din(w_dff_A_5acy51VL2_1),.clk(gclk));
	jdff dff_A_SLdMtM8b8_1(.dout(w_G446_0[1]),.din(w_dff_A_SLdMtM8b8_1),.clk(gclk));
	jdff dff_A_d3aCecw68_1(.dout(w_dff_A_SLdMtM8b8_1),.din(w_dff_A_d3aCecw68_1),.clk(gclk));
	jdff dff_A_YcZ4Jqcu3_1(.dout(w_dff_A_d3aCecw68_1),.din(w_dff_A_YcZ4Jqcu3_1),.clk(gclk));
	jdff dff_A_mw3Zve2w6_1(.dout(w_dff_A_YcZ4Jqcu3_1),.din(w_dff_A_mw3Zve2w6_1),.clk(gclk));
	jdff dff_A_Yi7meXIa0_2(.dout(w_G446_0[2]),.din(w_dff_A_Yi7meXIa0_2),.clk(gclk));
	jdff dff_A_tol8jPOT1_2(.dout(w_dff_A_Yi7meXIa0_2),.din(w_dff_A_tol8jPOT1_2),.clk(gclk));
	jdff dff_A_8xvh3C4x5_2(.dout(w_dff_A_tol8jPOT1_2),.din(w_dff_A_8xvh3C4x5_2),.clk(gclk));
	jdff dff_A_fLq7odAN5_2(.dout(w_dff_A_8xvh3C4x5_2),.din(w_dff_A_fLq7odAN5_2),.clk(gclk));
	jdff dff_A_Iri93B0L9_0(.dout(w_G206_0[0]),.din(w_dff_A_Iri93B0L9_0),.clk(gclk));
	jdff dff_B_cQGu051n7_1(.din(n1458),.dout(w_dff_B_cQGu051n7_1),.clk(gclk));
	jdff dff_B_gleghccY1_1(.din(n1459),.dout(w_dff_B_gleghccY1_1),.clk(gclk));
	jdff dff_A_WP939Db63_0(.dout(w_G242_1[0]),.din(w_dff_A_WP939Db63_0),.clk(gclk));
	jdff dff_A_m8xX8rCk2_1(.dout(w_G242_1[1]),.din(w_dff_A_m8xX8rCk2_1),.clk(gclk));
	jdff dff_A_cJfO8GK75_1(.dout(w_G242_0[1]),.din(w_dff_A_cJfO8GK75_1),.clk(gclk));
	jdff dff_A_hCUj84rT2_2(.dout(w_G242_0[2]),.din(w_dff_A_hCUj84rT2_2),.clk(gclk));
	jdff dff_A_DcYzTp8C6_2(.dout(w_G248_3[2]),.din(w_dff_A_DcYzTp8C6_2),.clk(gclk));
	jdff dff_A_eoHESROo4_1(.dout(w_n462_0[1]),.din(w_dff_A_eoHESROo4_1),.clk(gclk));
	jdff dff_A_yes0HgDd1_1(.dout(w_dff_A_eoHESROo4_1),.din(w_dff_A_yes0HgDd1_1),.clk(gclk));
	jdff dff_A_kgki6oiX8_1(.dout(w_dff_A_yes0HgDd1_1),.din(w_dff_A_kgki6oiX8_1),.clk(gclk));
	jdff dff_A_3aaz8XkD0_1(.dout(w_dff_A_kgki6oiX8_1),.din(w_dff_A_3aaz8XkD0_1),.clk(gclk));
	jdff dff_A_4vYs8wAb7_2(.dout(w_n462_0[2]),.din(w_dff_A_4vYs8wAb7_2),.clk(gclk));
	jdff dff_A_1TuDV9NO0_0(.dout(w_G435_1[0]),.din(w_dff_A_1TuDV9NO0_0),.clk(gclk));
	jdff dff_A_EgU4L2EN6_0(.dout(w_dff_A_1TuDV9NO0_0),.din(w_dff_A_EgU4L2EN6_0),.clk(gclk));
	jdff dff_A_ffFxNKV48_0(.dout(w_dff_A_EgU4L2EN6_0),.din(w_dff_A_ffFxNKV48_0),.clk(gclk));
	jdff dff_A_Jgsa7gf44_0(.dout(w_dff_A_ffFxNKV48_0),.din(w_dff_A_Jgsa7gf44_0),.clk(gclk));
	jdff dff_A_8PTPxEZU2_1(.dout(w_G435_1[1]),.din(w_dff_A_8PTPxEZU2_1),.clk(gclk));
	jdff dff_A_eMy77nlV4_1(.dout(w_G435_0[1]),.din(w_dff_A_eMy77nlV4_1),.clk(gclk));
	jdff dff_A_KBCP7C4J6_1(.dout(w_dff_A_eMy77nlV4_1),.din(w_dff_A_KBCP7C4J6_1),.clk(gclk));
	jdff dff_A_1UlOwWN55_2(.dout(w_G435_0[2]),.din(w_dff_A_1UlOwWN55_2),.clk(gclk));
	jdff dff_A_SAia8h8T3_2(.dout(w_dff_A_1UlOwWN55_2),.din(w_dff_A_SAia8h8T3_2),.clk(gclk));
	jdff dff_A_aieTzyUI2_2(.dout(w_dff_A_SAia8h8T3_2),.din(w_dff_A_aieTzyUI2_2),.clk(gclk));
	jdff dff_A_5srVuwcl4_2(.dout(w_dff_A_aieTzyUI2_2),.din(w_dff_A_5srVuwcl4_2),.clk(gclk));
	jdff dff_A_KEFDYI724_1(.dout(w_G251_0[1]),.din(w_dff_A_KEFDYI724_1),.clk(gclk));
	jdff dff_A_UWfb0VmV7_2(.dout(w_G251_0[2]),.din(w_dff_A_UWfb0VmV7_2),.clk(gclk));
	jdff dff_A_kc6Gp8Ba3_0(.dout(w_G234_2[0]),.din(w_dff_A_kc6Gp8Ba3_0),.clk(gclk));
	jdff dff_A_xxiY3hzF4_2(.dout(w_G234_0[2]),.din(w_dff_A_xxiY3hzF4_2),.clk(gclk));
	jdff dff_A_viGpsNUS2_0(.dout(w_G4092_1[0]),.din(w_dff_A_viGpsNUS2_0),.clk(gclk));
	jdff dff_A_73wzFBMd0_0(.dout(w_dff_A_viGpsNUS2_0),.din(w_dff_A_73wzFBMd0_0),.clk(gclk));
	jdff dff_A_eusntHHy5_0(.dout(w_dff_A_73wzFBMd0_0),.din(w_dff_A_eusntHHy5_0),.clk(gclk));
	jdff dff_A_ef7UMty77_0(.dout(w_dff_A_eusntHHy5_0),.din(w_dff_A_ef7UMty77_0),.clk(gclk));
	jdff dff_A_YSEkqc135_0(.dout(w_dff_A_ef7UMty77_0),.din(w_dff_A_YSEkqc135_0),.clk(gclk));
	jdff dff_A_BBXnGp3V1_0(.dout(w_dff_A_YSEkqc135_0),.din(w_dff_A_BBXnGp3V1_0),.clk(gclk));
	jdff dff_A_F0NkKZMh2_0(.dout(w_dff_A_BBXnGp3V1_0),.din(w_dff_A_F0NkKZMh2_0),.clk(gclk));
	jdff dff_A_xZchiVRd2_0(.dout(w_dff_A_F0NkKZMh2_0),.din(w_dff_A_xZchiVRd2_0),.clk(gclk));
	jdff dff_A_f6xoYpup5_0(.dout(w_dff_A_xZchiVRd2_0),.din(w_dff_A_f6xoYpup5_0),.clk(gclk));
	jdff dff_A_MpgP6oaC4_0(.dout(w_dff_A_f6xoYpup5_0),.din(w_dff_A_MpgP6oaC4_0),.clk(gclk));
	jdff dff_A_I4mWuMdI9_0(.dout(w_dff_A_MpgP6oaC4_0),.din(w_dff_A_I4mWuMdI9_0),.clk(gclk));
	jdff dff_A_X5iFbqWZ6_1(.dout(w_G4092_1[1]),.din(w_dff_A_X5iFbqWZ6_1),.clk(gclk));
	jdff dff_A_paExvVgh1_0(.dout(w_n999_1[0]),.din(w_dff_A_paExvVgh1_0),.clk(gclk));
	jdff dff_A_z9T9hpxY0_0(.dout(w_dff_A_paExvVgh1_0),.din(w_dff_A_z9T9hpxY0_0),.clk(gclk));
	jdff dff_A_UKZDXthg8_0(.dout(w_dff_A_z9T9hpxY0_0),.din(w_dff_A_UKZDXthg8_0),.clk(gclk));
	jdff dff_A_xmJ00wV22_0(.dout(w_dff_A_UKZDXthg8_0),.din(w_dff_A_xmJ00wV22_0),.clk(gclk));
	jdff dff_A_yV3IXiGf0_0(.dout(w_dff_A_xmJ00wV22_0),.din(w_dff_A_yV3IXiGf0_0),.clk(gclk));
	jdff dff_A_m54Pr7NK1_0(.dout(w_dff_A_yV3IXiGf0_0),.din(w_dff_A_m54Pr7NK1_0),.clk(gclk));
	jdff dff_A_WnuzEvYQ9_0(.dout(w_dff_A_m54Pr7NK1_0),.din(w_dff_A_WnuzEvYQ9_0),.clk(gclk));
	jdff dff_A_uA2oguuJ4_2(.dout(w_n999_1[2]),.din(w_dff_A_uA2oguuJ4_2),.clk(gclk));
	jdff dff_A_Z8XlFiam4_2(.dout(w_dff_A_uA2oguuJ4_2),.din(w_dff_A_Z8XlFiam4_2),.clk(gclk));
	jdff dff_A_V2vDih6Z4_2(.dout(w_dff_A_Z8XlFiam4_2),.din(w_dff_A_V2vDih6Z4_2),.clk(gclk));
	jdff dff_A_B3VACOQO5_2(.dout(w_dff_A_V2vDih6Z4_2),.din(w_dff_A_B3VACOQO5_2),.clk(gclk));
	jdff dff_A_YdI9tNGe6_2(.dout(w_dff_A_B3VACOQO5_2),.din(w_dff_A_YdI9tNGe6_2),.clk(gclk));
	jdff dff_A_25CNjiae8_2(.dout(w_dff_A_YdI9tNGe6_2),.din(w_dff_A_25CNjiae8_2),.clk(gclk));
	jdff dff_A_GA86mqIH2_2(.dout(w_dff_A_25CNjiae8_2),.din(w_dff_A_GA86mqIH2_2),.clk(gclk));
	jdff dff_A_OXYgzVS37_2(.dout(w_dff_A_GA86mqIH2_2),.din(w_dff_A_OXYgzVS37_2),.clk(gclk));
	jdff dff_A_rSPrbVlt1_2(.dout(w_dff_A_OXYgzVS37_2),.din(w_dff_A_rSPrbVlt1_2),.clk(gclk));
	jdff dff_A_P7dYRDUJ9_2(.dout(w_dff_A_rSPrbVlt1_2),.din(w_dff_A_P7dYRDUJ9_2),.clk(gclk));
	jdff dff_A_yj4tkaQ32_2(.dout(w_dff_A_P7dYRDUJ9_2),.din(w_dff_A_yj4tkaQ32_2),.clk(gclk));
	jdff dff_A_eqbKIpKc0_2(.dout(w_dff_A_yj4tkaQ32_2),.din(w_dff_A_eqbKIpKc0_2),.clk(gclk));
	jdff dff_A_NxKFlP6E5_2(.dout(w_dff_A_eqbKIpKc0_2),.din(w_dff_A_NxKFlP6E5_2),.clk(gclk));
	jdff dff_A_KpIEWaYu1_2(.dout(w_dff_A_NxKFlP6E5_2),.din(w_dff_A_KpIEWaYu1_2),.clk(gclk));
	jdff dff_A_cA8amEaP6_2(.dout(w_dff_A_KpIEWaYu1_2),.din(w_dff_A_cA8amEaP6_2),.clk(gclk));
	jdff dff_A_0IEw0WLI3_2(.dout(w_dff_A_cA8amEaP6_2),.din(w_dff_A_0IEw0WLI3_2),.clk(gclk));
	jdff dff_A_a9MBk0zK8_2(.dout(w_dff_A_0IEw0WLI3_2),.din(w_dff_A_a9MBk0zK8_2),.clk(gclk));
	jdff dff_A_jMDahzlB6_2(.dout(w_dff_A_a9MBk0zK8_2),.din(w_dff_A_jMDahzlB6_2),.clk(gclk));
	jdff dff_A_EYUNAq5J7_2(.dout(w_dff_A_jMDahzlB6_2),.din(w_dff_A_EYUNAq5J7_2),.clk(gclk));
	jdff dff_A_U9LGVDfH9_1(.dout(w_n999_0[1]),.din(w_dff_A_U9LGVDfH9_1),.clk(gclk));
	jdff dff_A_pqBhYW279_1(.dout(w_dff_A_U9LGVDfH9_1),.din(w_dff_A_pqBhYW279_1),.clk(gclk));
	jdff dff_A_1tJYaH7l4_1(.dout(w_dff_A_pqBhYW279_1),.din(w_dff_A_1tJYaH7l4_1),.clk(gclk));
	jdff dff_A_0x5ZJo1h4_1(.dout(w_dff_A_1tJYaH7l4_1),.din(w_dff_A_0x5ZJo1h4_1),.clk(gclk));
	jdff dff_A_8lB0GH520_1(.dout(w_dff_A_0x5ZJo1h4_1),.din(w_dff_A_8lB0GH520_1),.clk(gclk));
	jdff dff_A_CFa9rKFI5_1(.dout(w_dff_A_8lB0GH520_1),.din(w_dff_A_CFa9rKFI5_1),.clk(gclk));
	jdff dff_A_bmZURhFr1_1(.dout(w_dff_A_CFa9rKFI5_1),.din(w_dff_A_bmZURhFr1_1),.clk(gclk));
	jdff dff_A_Eri2EBMQ1_1(.dout(w_dff_A_bmZURhFr1_1),.din(w_dff_A_Eri2EBMQ1_1),.clk(gclk));
	jdff dff_A_ZCRpgCFQ0_1(.dout(w_dff_A_Eri2EBMQ1_1),.din(w_dff_A_ZCRpgCFQ0_1),.clk(gclk));
	jdff dff_A_IljkbICw2_1(.dout(w_dff_A_ZCRpgCFQ0_1),.din(w_dff_A_IljkbICw2_1),.clk(gclk));
	jdff dff_A_eK0j9ZaM5_1(.dout(w_dff_A_IljkbICw2_1),.din(w_dff_A_eK0j9ZaM5_1),.clk(gclk));
	jdff dff_A_UyraIZti2_1(.dout(w_dff_A_eK0j9ZaM5_1),.din(w_dff_A_UyraIZti2_1),.clk(gclk));
	jdff dff_A_KcEHa6Yr4_1(.dout(w_dff_A_UyraIZti2_1),.din(w_dff_A_KcEHa6Yr4_1),.clk(gclk));
	jdff dff_A_bH6cEhzw1_1(.dout(w_dff_A_KcEHa6Yr4_1),.din(w_dff_A_bH6cEhzw1_1),.clk(gclk));
	jdff dff_A_mOFV86Bz2_1(.dout(w_dff_A_bH6cEhzw1_1),.din(w_dff_A_mOFV86Bz2_1),.clk(gclk));
	jdff dff_A_1Ox31FK61_1(.dout(w_dff_A_mOFV86Bz2_1),.din(w_dff_A_1Ox31FK61_1),.clk(gclk));
	jdff dff_A_XUckKp2H8_1(.dout(w_dff_A_1Ox31FK61_1),.din(w_dff_A_XUckKp2H8_1),.clk(gclk));
	jdff dff_A_8Ep4cE458_2(.dout(w_n999_0[2]),.din(w_dff_A_8Ep4cE458_2),.clk(gclk));
	jdff dff_A_NBBAmwgZ2_2(.dout(w_dff_A_8Ep4cE458_2),.din(w_dff_A_NBBAmwgZ2_2),.clk(gclk));
	jdff dff_A_buy3CmPo8_2(.dout(w_dff_A_NBBAmwgZ2_2),.din(w_dff_A_buy3CmPo8_2),.clk(gclk));
	jdff dff_A_BFHhjxBJ5_2(.dout(w_dff_A_buy3CmPo8_2),.din(w_dff_A_BFHhjxBJ5_2),.clk(gclk));
	jdff dff_A_Dyiuatp05_2(.dout(w_dff_A_BFHhjxBJ5_2),.din(w_dff_A_Dyiuatp05_2),.clk(gclk));
	jdff dff_A_WAXdgUYi1_2(.dout(w_dff_A_Dyiuatp05_2),.din(w_dff_A_WAXdgUYi1_2),.clk(gclk));
	jdff dff_A_LCgryU6H4_2(.dout(w_dff_A_WAXdgUYi1_2),.din(w_dff_A_LCgryU6H4_2),.clk(gclk));
	jdff dff_A_mBeDuA271_2(.dout(w_dff_A_LCgryU6H4_2),.din(w_dff_A_mBeDuA271_2),.clk(gclk));
	jdff dff_A_XWAPLWbL5_2(.dout(w_dff_A_mBeDuA271_2),.din(w_dff_A_XWAPLWbL5_2),.clk(gclk));
	jdff dff_A_ui7oAtrb7_2(.dout(w_dff_A_XWAPLWbL5_2),.din(w_dff_A_ui7oAtrb7_2),.clk(gclk));
	jdff dff_A_9XPHNBBU0_2(.dout(w_dff_A_ui7oAtrb7_2),.din(w_dff_A_9XPHNBBU0_2),.clk(gclk));
	jdff dff_A_sIWnwDEh7_1(.dout(w_G1694_0[1]),.din(w_dff_A_sIWnwDEh7_1),.clk(gclk));
	jdff dff_A_FgyHJt2a3_2(.dout(w_G1691_0[2]),.din(w_dff_A_FgyHJt2a3_2),.clk(gclk));
	jdff dff_B_I4fAPK9e7_2(.din(n1624),.dout(w_dff_B_I4fAPK9e7_2),.clk(gclk));
	jdff dff_B_4H455TCA6_2(.din(w_dff_B_I4fAPK9e7_2),.dout(w_dff_B_4H455TCA6_2),.clk(gclk));
	jdff dff_B_ZZ47TlVM0_2(.din(w_dff_B_4H455TCA6_2),.dout(w_dff_B_ZZ47TlVM0_2),.clk(gclk));
	jdff dff_B_dRf9BErv4_2(.din(w_dff_B_ZZ47TlVM0_2),.dout(w_dff_B_dRf9BErv4_2),.clk(gclk));
	jdff dff_B_STXNS9JG9_2(.din(w_dff_B_dRf9BErv4_2),.dout(w_dff_B_STXNS9JG9_2),.clk(gclk));
	jdff dff_B_XASqlK6q9_2(.din(w_dff_B_STXNS9JG9_2),.dout(w_dff_B_XASqlK6q9_2),.clk(gclk));
	jdff dff_B_BlCSfxRv7_2(.din(w_dff_B_XASqlK6q9_2),.dout(w_dff_B_BlCSfxRv7_2),.clk(gclk));
	jdff dff_B_JUaKTUWs0_2(.din(w_dff_B_BlCSfxRv7_2),.dout(w_dff_B_JUaKTUWs0_2),.clk(gclk));
	jdff dff_B_82I58rjp0_2(.din(w_dff_B_JUaKTUWs0_2),.dout(w_dff_B_82I58rjp0_2),.clk(gclk));
	jdff dff_B_Mvh5p9V32_2(.din(w_dff_B_82I58rjp0_2),.dout(w_dff_B_Mvh5p9V32_2),.clk(gclk));
	jdff dff_B_D3YV7bYd5_2(.din(w_dff_B_Mvh5p9V32_2),.dout(w_dff_B_D3YV7bYd5_2),.clk(gclk));
	jdff dff_B_6zTa0c6n0_2(.din(w_dff_B_D3YV7bYd5_2),.dout(w_dff_B_6zTa0c6n0_2),.clk(gclk));
	jdff dff_B_F2GTTvIS0_2(.din(w_dff_B_6zTa0c6n0_2),.dout(w_dff_B_F2GTTvIS0_2),.clk(gclk));
	jdff dff_B_yjTMlEDO2_2(.din(w_dff_B_F2GTTvIS0_2),.dout(w_dff_B_yjTMlEDO2_2),.clk(gclk));
	jdff dff_B_xN6DHAUf0_2(.din(w_dff_B_yjTMlEDO2_2),.dout(w_dff_B_xN6DHAUf0_2),.clk(gclk));
	jdff dff_B_lzCdJ9k40_2(.din(w_dff_B_xN6DHAUf0_2),.dout(w_dff_B_lzCdJ9k40_2),.clk(gclk));
	jdff dff_B_nHxI0s1Y8_2(.din(w_dff_B_lzCdJ9k40_2),.dout(w_dff_B_nHxI0s1Y8_2),.clk(gclk));
	jdff dff_B_E3zpKwOW7_2(.din(w_dff_B_nHxI0s1Y8_2),.dout(w_dff_B_E3zpKwOW7_2),.clk(gclk));
	jdff dff_B_uOSiCRB66_2(.din(w_dff_B_E3zpKwOW7_2),.dout(w_dff_B_uOSiCRB66_2),.clk(gclk));
	jdff dff_B_yrnmnuY47_2(.din(w_dff_B_uOSiCRB66_2),.dout(w_dff_B_yrnmnuY47_2),.clk(gclk));
	jdff dff_B_YYSXf3Cw1_2(.din(w_dff_B_yrnmnuY47_2),.dout(w_dff_B_YYSXf3Cw1_2),.clk(gclk));
	jdff dff_B_Y8KiCjfk3_2(.din(w_dff_B_YYSXf3Cw1_2),.dout(w_dff_B_Y8KiCjfk3_2),.clk(gclk));
	jdff dff_B_qJRpuyjt6_2(.din(w_dff_B_Y8KiCjfk3_2),.dout(w_dff_B_qJRpuyjt6_2),.clk(gclk));
	jdff dff_B_SUr3R1MO3_2(.din(w_dff_B_qJRpuyjt6_2),.dout(w_dff_B_SUr3R1MO3_2),.clk(gclk));
	jdff dff_A_Er0lPOGE3_2(.dout(w_G137_3[2]),.din(w_dff_A_Er0lPOGE3_2),.clk(gclk));
	jdff dff_A_JSk4D0w16_2(.dout(w_dff_A_Er0lPOGE3_2),.din(w_dff_A_JSk4D0w16_2),.clk(gclk));
	jdff dff_A_0o1yUlot0_2(.dout(w_dff_A_JSk4D0w16_2),.din(w_dff_A_0o1yUlot0_2),.clk(gclk));
	jdff dff_A_eyin0HN03_2(.dout(w_dff_A_0o1yUlot0_2),.din(w_dff_A_eyin0HN03_2),.clk(gclk));
	jdff dff_A_gZs5dwrj8_2(.dout(w_dff_A_eyin0HN03_2),.din(w_dff_A_gZs5dwrj8_2),.clk(gclk));
	jdff dff_A_9UTA3UMW8_2(.dout(w_dff_A_gZs5dwrj8_2),.din(w_dff_A_9UTA3UMW8_2),.clk(gclk));
	jdff dff_A_ixkDvfLk6_2(.dout(w_dff_A_9UTA3UMW8_2),.din(w_dff_A_ixkDvfLk6_2),.clk(gclk));
	jdff dff_A_X7PDkg0r9_2(.dout(w_dff_A_ixkDvfLk6_2),.din(w_dff_A_X7PDkg0r9_2),.clk(gclk));
	jdff dff_A_aYbBW02x0_2(.dout(w_dff_A_X7PDkg0r9_2),.din(w_dff_A_aYbBW02x0_2),.clk(gclk));
	jdff dff_A_tTdMNgQg1_2(.dout(w_dff_A_aYbBW02x0_2),.din(w_dff_A_tTdMNgQg1_2),.clk(gclk));
	jdff dff_A_HiGLvP440_2(.dout(w_dff_A_tTdMNgQg1_2),.din(w_dff_A_HiGLvP440_2),.clk(gclk));
	jdff dff_A_8v3DeU6y5_2(.dout(w_dff_A_HiGLvP440_2),.din(w_dff_A_8v3DeU6y5_2),.clk(gclk));
	jdff dff_A_Ohp9CgnO1_2(.dout(w_dff_A_8v3DeU6y5_2),.din(w_dff_A_Ohp9CgnO1_2),.clk(gclk));
	jdff dff_A_eSsG7fWD5_2(.dout(w_dff_A_Ohp9CgnO1_2),.din(w_dff_A_eSsG7fWD5_2),.clk(gclk));
	jdff dff_A_ZGCSzzn94_2(.dout(w_dff_A_eSsG7fWD5_2),.din(w_dff_A_ZGCSzzn94_2),.clk(gclk));
	jdff dff_A_KZHb8zjT1_2(.dout(w_dff_A_ZGCSzzn94_2),.din(w_dff_A_KZHb8zjT1_2),.clk(gclk));
	jdff dff_A_KTxw2vow3_2(.dout(w_dff_A_KZHb8zjT1_2),.din(w_dff_A_KTxw2vow3_2),.clk(gclk));
	jdff dff_A_SRCD7BNj2_2(.dout(w_dff_A_KTxw2vow3_2),.din(w_dff_A_SRCD7BNj2_2),.clk(gclk));
	jdff dff_A_pKCtvoOt9_2(.dout(w_dff_A_SRCD7BNj2_2),.din(w_dff_A_pKCtvoOt9_2),.clk(gclk));
	jdff dff_A_o9V2RABJ1_2(.dout(w_dff_A_pKCtvoOt9_2),.din(w_dff_A_o9V2RABJ1_2),.clk(gclk));
	jdff dff_A_KOoTQLek9_2(.dout(w_dff_A_o9V2RABJ1_2),.din(w_dff_A_KOoTQLek9_2),.clk(gclk));
	jdff dff_A_IntbbyyG8_2(.dout(w_dff_A_KOoTQLek9_2),.din(w_dff_A_IntbbyyG8_2),.clk(gclk));
	jdff dff_A_vbqnXyDv5_2(.dout(w_dff_A_IntbbyyG8_2),.din(w_dff_A_vbqnXyDv5_2),.clk(gclk));
	jdff dff_A_URHU4IuH9_0(.dout(w_G137_0[0]),.din(w_dff_A_URHU4IuH9_0),.clk(gclk));
	jdff dff_A_uu1NyUgA1_0(.dout(w_dff_A_URHU4IuH9_0),.din(w_dff_A_uu1NyUgA1_0),.clk(gclk));
	jdff dff_A_aIBjR3T21_0(.dout(w_dff_A_uu1NyUgA1_0),.din(w_dff_A_aIBjR3T21_0),.clk(gclk));
	jdff dff_A_H8jccFVF9_0(.dout(w_dff_A_aIBjR3T21_0),.din(w_dff_A_H8jccFVF9_0),.clk(gclk));
	jdff dff_A_fFriHcp03_0(.dout(w_dff_A_H8jccFVF9_0),.din(w_dff_A_fFriHcp03_0),.clk(gclk));
	jdff dff_A_qiJpGME05_0(.dout(w_dff_A_fFriHcp03_0),.din(w_dff_A_qiJpGME05_0),.clk(gclk));
	jdff dff_A_tpzyB56f6_0(.dout(w_dff_A_qiJpGME05_0),.din(w_dff_A_tpzyB56f6_0),.clk(gclk));
	jdff dff_A_Tj6fM6md4_0(.dout(w_dff_A_tpzyB56f6_0),.din(w_dff_A_Tj6fM6md4_0),.clk(gclk));
	jdff dff_A_klsyIl0w4_0(.dout(w_dff_A_Tj6fM6md4_0),.din(w_dff_A_klsyIl0w4_0),.clk(gclk));
	jdff dff_A_XpyP0Agr4_0(.dout(w_dff_A_klsyIl0w4_0),.din(w_dff_A_XpyP0Agr4_0),.clk(gclk));
	jdff dff_A_EUchdzbn9_0(.dout(w_dff_A_XpyP0Agr4_0),.din(w_dff_A_EUchdzbn9_0),.clk(gclk));
	jdff dff_A_Z0RAvOnB2_0(.dout(w_dff_A_EUchdzbn9_0),.din(w_dff_A_Z0RAvOnB2_0),.clk(gclk));
	jdff dff_A_A9U70sOV4_0(.dout(w_dff_A_Z0RAvOnB2_0),.din(w_dff_A_A9U70sOV4_0),.clk(gclk));
	jdff dff_A_tbZV8FCz1_0(.dout(w_dff_A_A9U70sOV4_0),.din(w_dff_A_tbZV8FCz1_0),.clk(gclk));
	jdff dff_A_TqW5byGS9_0(.dout(w_dff_A_tbZV8FCz1_0),.din(w_dff_A_TqW5byGS9_0),.clk(gclk));
	jdff dff_A_w46tlnWm0_0(.dout(w_dff_A_TqW5byGS9_0),.din(w_dff_A_w46tlnWm0_0),.clk(gclk));
	jdff dff_A_EZFj4lep1_1(.dout(w_G137_0[1]),.din(w_dff_A_EZFj4lep1_1),.clk(gclk));
	jdff dff_A_DzxPqTsI9_1(.dout(w_dff_A_EZFj4lep1_1),.din(w_dff_A_DzxPqTsI9_1),.clk(gclk));
	jdff dff_A_EcQsoT9g3_1(.dout(w_dff_A_DzxPqTsI9_1),.din(w_dff_A_EcQsoT9g3_1),.clk(gclk));
	jdff dff_A_Nyiiwyuu1_1(.dout(w_dff_A_EcQsoT9g3_1),.din(w_dff_A_Nyiiwyuu1_1),.clk(gclk));
	jdff dff_A_R2AOgfTK1_1(.dout(w_dff_A_Nyiiwyuu1_1),.din(w_dff_A_R2AOgfTK1_1),.clk(gclk));
	jdff dff_A_CKvgTkiE3_1(.dout(w_dff_A_R2AOgfTK1_1),.din(w_dff_A_CKvgTkiE3_1),.clk(gclk));
	jdff dff_A_jvrLVt7O3_1(.dout(w_dff_A_CKvgTkiE3_1),.din(w_dff_A_jvrLVt7O3_1),.clk(gclk));
	jdff dff_A_gcqKeMoa8_1(.dout(w_dff_A_jvrLVt7O3_1),.din(w_dff_A_gcqKeMoa8_1),.clk(gclk));
	jdff dff_A_ggVqkWvU9_1(.dout(w_dff_A_gcqKeMoa8_1),.din(w_dff_A_ggVqkWvU9_1),.clk(gclk));
	jdff dff_A_i1Rasi4v5_1(.dout(w_dff_A_ggVqkWvU9_1),.din(w_dff_A_i1Rasi4v5_1),.clk(gclk));
	jdff dff_A_ZmlcfrZO8_1(.dout(w_dff_A_i1Rasi4v5_1),.din(w_dff_A_ZmlcfrZO8_1),.clk(gclk));
	jdff dff_A_EBC8N9T79_1(.dout(w_dff_A_js2yMspE4_0),.din(w_dff_A_EBC8N9T79_1),.clk(gclk));
	jdff dff_A_js2yMspE4_0(.dout(w_dff_A_ETMMXGaF0_0),.din(w_dff_A_js2yMspE4_0),.clk(gclk));
	jdff dff_A_ETMMXGaF0_0(.dout(w_dff_A_J4U27oSg2_0),.din(w_dff_A_ETMMXGaF0_0),.clk(gclk));
	jdff dff_A_J4U27oSg2_0(.dout(w_dff_A_yw8o5U4R2_0),.din(w_dff_A_J4U27oSg2_0),.clk(gclk));
	jdff dff_A_yw8o5U4R2_0(.dout(w_dff_A_tJc0cKRv9_0),.din(w_dff_A_yw8o5U4R2_0),.clk(gclk));
	jdff dff_A_tJc0cKRv9_0(.dout(w_dff_A_rZAseHNZ2_0),.din(w_dff_A_tJc0cKRv9_0),.clk(gclk));
	jdff dff_A_rZAseHNZ2_0(.dout(w_dff_A_VBTPSrG00_0),.din(w_dff_A_rZAseHNZ2_0),.clk(gclk));
	jdff dff_A_VBTPSrG00_0(.dout(w_dff_A_9fyArUqG1_0),.din(w_dff_A_VBTPSrG00_0),.clk(gclk));
	jdff dff_A_9fyArUqG1_0(.dout(w_dff_A_uvRscf898_0),.din(w_dff_A_9fyArUqG1_0),.clk(gclk));
	jdff dff_A_uvRscf898_0(.dout(w_dff_A_przgP03g2_0),.din(w_dff_A_uvRscf898_0),.clk(gclk));
	jdff dff_A_przgP03g2_0(.dout(w_dff_A_swLddxws3_0),.din(w_dff_A_przgP03g2_0),.clk(gclk));
	jdff dff_A_swLddxws3_0(.dout(w_dff_A_nam4BOlK4_0),.din(w_dff_A_swLddxws3_0),.clk(gclk));
	jdff dff_A_nam4BOlK4_0(.dout(w_dff_A_ohgHWyp62_0),.din(w_dff_A_nam4BOlK4_0),.clk(gclk));
	jdff dff_A_ohgHWyp62_0(.dout(w_dff_A_Nx0DBZ8l6_0),.din(w_dff_A_ohgHWyp62_0),.clk(gclk));
	jdff dff_A_Nx0DBZ8l6_0(.dout(w_dff_A_ovoHPIdI6_0),.din(w_dff_A_Nx0DBZ8l6_0),.clk(gclk));
	jdff dff_A_ovoHPIdI6_0(.dout(w_dff_A_vm0Sb9pr3_0),.din(w_dff_A_ovoHPIdI6_0),.clk(gclk));
	jdff dff_A_vm0Sb9pr3_0(.dout(w_dff_A_wb4zkTA16_0),.din(w_dff_A_vm0Sb9pr3_0),.clk(gclk));
	jdff dff_A_wb4zkTA16_0(.dout(w_dff_A_GPiQ5TuP8_0),.din(w_dff_A_wb4zkTA16_0),.clk(gclk));
	jdff dff_A_GPiQ5TuP8_0(.dout(w_dff_A_3Jvt1A2P3_0),.din(w_dff_A_GPiQ5TuP8_0),.clk(gclk));
	jdff dff_A_3Jvt1A2P3_0(.dout(w_dff_A_a8ceP99Q8_0),.din(w_dff_A_3Jvt1A2P3_0),.clk(gclk));
	jdff dff_A_a8ceP99Q8_0(.dout(w_dff_A_UIbrAWwd8_0),.din(w_dff_A_a8ceP99Q8_0),.clk(gclk));
	jdff dff_A_UIbrAWwd8_0(.dout(w_dff_A_fnZgtWOm9_0),.din(w_dff_A_UIbrAWwd8_0),.clk(gclk));
	jdff dff_A_fnZgtWOm9_0(.dout(w_dff_A_8VO7QJRY0_0),.din(w_dff_A_fnZgtWOm9_0),.clk(gclk));
	jdff dff_A_8VO7QJRY0_0(.dout(w_dff_A_8iXvTUpm7_0),.din(w_dff_A_8VO7QJRY0_0),.clk(gclk));
	jdff dff_A_8iXvTUpm7_0(.dout(w_dff_A_4dUJQMso6_0),.din(w_dff_A_8iXvTUpm7_0),.clk(gclk));
	jdff dff_A_4dUJQMso6_0(.dout(G144),.din(w_dff_A_4dUJQMso6_0),.clk(gclk));
	jdff dff_A_kk7cd6j65_1(.dout(w_dff_A_Afz9WXRJ5_0),.din(w_dff_A_kk7cd6j65_1),.clk(gclk));
	jdff dff_A_Afz9WXRJ5_0(.dout(w_dff_A_QTfMMhmG7_0),.din(w_dff_A_Afz9WXRJ5_0),.clk(gclk));
	jdff dff_A_QTfMMhmG7_0(.dout(w_dff_A_UwQjHgiN5_0),.din(w_dff_A_QTfMMhmG7_0),.clk(gclk));
	jdff dff_A_UwQjHgiN5_0(.dout(w_dff_A_6fDo3UPn2_0),.din(w_dff_A_UwQjHgiN5_0),.clk(gclk));
	jdff dff_A_6fDo3UPn2_0(.dout(w_dff_A_2ci3SdFX7_0),.din(w_dff_A_6fDo3UPn2_0),.clk(gclk));
	jdff dff_A_2ci3SdFX7_0(.dout(w_dff_A_cll7EyyK5_0),.din(w_dff_A_2ci3SdFX7_0),.clk(gclk));
	jdff dff_A_cll7EyyK5_0(.dout(w_dff_A_z3lprCox2_0),.din(w_dff_A_cll7EyyK5_0),.clk(gclk));
	jdff dff_A_z3lprCox2_0(.dout(w_dff_A_IjdktLEQ4_0),.din(w_dff_A_z3lprCox2_0),.clk(gclk));
	jdff dff_A_IjdktLEQ4_0(.dout(w_dff_A_QkR49ma34_0),.din(w_dff_A_IjdktLEQ4_0),.clk(gclk));
	jdff dff_A_QkR49ma34_0(.dout(w_dff_A_6KvwVae57_0),.din(w_dff_A_QkR49ma34_0),.clk(gclk));
	jdff dff_A_6KvwVae57_0(.dout(w_dff_A_ZDRkilbs7_0),.din(w_dff_A_6KvwVae57_0),.clk(gclk));
	jdff dff_A_ZDRkilbs7_0(.dout(w_dff_A_9J2KbRkJ1_0),.din(w_dff_A_ZDRkilbs7_0),.clk(gclk));
	jdff dff_A_9J2KbRkJ1_0(.dout(w_dff_A_erEWjDxi5_0),.din(w_dff_A_9J2KbRkJ1_0),.clk(gclk));
	jdff dff_A_erEWjDxi5_0(.dout(w_dff_A_WYboSFBI7_0),.din(w_dff_A_erEWjDxi5_0),.clk(gclk));
	jdff dff_A_WYboSFBI7_0(.dout(w_dff_A_51ysUhir2_0),.din(w_dff_A_WYboSFBI7_0),.clk(gclk));
	jdff dff_A_51ysUhir2_0(.dout(w_dff_A_OwtHNWEa3_0),.din(w_dff_A_51ysUhir2_0),.clk(gclk));
	jdff dff_A_OwtHNWEa3_0(.dout(w_dff_A_potMbMC38_0),.din(w_dff_A_OwtHNWEa3_0),.clk(gclk));
	jdff dff_A_potMbMC38_0(.dout(w_dff_A_gZb5bDv29_0),.din(w_dff_A_potMbMC38_0),.clk(gclk));
	jdff dff_A_gZb5bDv29_0(.dout(w_dff_A_8iW0Sl4i6_0),.din(w_dff_A_gZb5bDv29_0),.clk(gclk));
	jdff dff_A_8iW0Sl4i6_0(.dout(w_dff_A_dapypv925_0),.din(w_dff_A_8iW0Sl4i6_0),.clk(gclk));
	jdff dff_A_dapypv925_0(.dout(w_dff_A_oRvrw7KV7_0),.din(w_dff_A_dapypv925_0),.clk(gclk));
	jdff dff_A_oRvrw7KV7_0(.dout(w_dff_A_kKNB3afA4_0),.din(w_dff_A_oRvrw7KV7_0),.clk(gclk));
	jdff dff_A_kKNB3afA4_0(.dout(w_dff_A_A0f1L1Lt5_0),.din(w_dff_A_kKNB3afA4_0),.clk(gclk));
	jdff dff_A_A0f1L1Lt5_0(.dout(w_dff_A_afSXXLl07_0),.din(w_dff_A_A0f1L1Lt5_0),.clk(gclk));
	jdff dff_A_afSXXLl07_0(.dout(w_dff_A_TK4XX8yx8_0),.din(w_dff_A_afSXXLl07_0),.clk(gclk));
	jdff dff_A_TK4XX8yx8_0(.dout(G298),.din(w_dff_A_TK4XX8yx8_0),.clk(gclk));
	jdff dff_A_a27FDOlD2_1(.dout(w_dff_A_7kA1e56U5_0),.din(w_dff_A_a27FDOlD2_1),.clk(gclk));
	jdff dff_A_7kA1e56U5_0(.dout(w_dff_A_dpgSKpl85_0),.din(w_dff_A_7kA1e56U5_0),.clk(gclk));
	jdff dff_A_dpgSKpl85_0(.dout(w_dff_A_DMyUoc0k3_0),.din(w_dff_A_dpgSKpl85_0),.clk(gclk));
	jdff dff_A_DMyUoc0k3_0(.dout(w_dff_A_vXrsnBNS9_0),.din(w_dff_A_DMyUoc0k3_0),.clk(gclk));
	jdff dff_A_vXrsnBNS9_0(.dout(w_dff_A_FjUPWESn4_0),.din(w_dff_A_vXrsnBNS9_0),.clk(gclk));
	jdff dff_A_FjUPWESn4_0(.dout(w_dff_A_JlvJ4awX3_0),.din(w_dff_A_FjUPWESn4_0),.clk(gclk));
	jdff dff_A_JlvJ4awX3_0(.dout(w_dff_A_RfMBeTad3_0),.din(w_dff_A_JlvJ4awX3_0),.clk(gclk));
	jdff dff_A_RfMBeTad3_0(.dout(w_dff_A_lyYrReaj8_0),.din(w_dff_A_RfMBeTad3_0),.clk(gclk));
	jdff dff_A_lyYrReaj8_0(.dout(w_dff_A_p6NWMAvP8_0),.din(w_dff_A_lyYrReaj8_0),.clk(gclk));
	jdff dff_A_p6NWMAvP8_0(.dout(w_dff_A_ktLqLAGX5_0),.din(w_dff_A_p6NWMAvP8_0),.clk(gclk));
	jdff dff_A_ktLqLAGX5_0(.dout(w_dff_A_nsKCijmv8_0),.din(w_dff_A_ktLqLAGX5_0),.clk(gclk));
	jdff dff_A_nsKCijmv8_0(.dout(w_dff_A_LHIomuu80_0),.din(w_dff_A_nsKCijmv8_0),.clk(gclk));
	jdff dff_A_LHIomuu80_0(.dout(w_dff_A_6wFpFbRk4_0),.din(w_dff_A_LHIomuu80_0),.clk(gclk));
	jdff dff_A_6wFpFbRk4_0(.dout(w_dff_A_rcvUU5IZ6_0),.din(w_dff_A_6wFpFbRk4_0),.clk(gclk));
	jdff dff_A_rcvUU5IZ6_0(.dout(w_dff_A_8qSdgszb4_0),.din(w_dff_A_rcvUU5IZ6_0),.clk(gclk));
	jdff dff_A_8qSdgszb4_0(.dout(w_dff_A_yFexwtY77_0),.din(w_dff_A_8qSdgszb4_0),.clk(gclk));
	jdff dff_A_yFexwtY77_0(.dout(w_dff_A_xda3Vy0d6_0),.din(w_dff_A_yFexwtY77_0),.clk(gclk));
	jdff dff_A_xda3Vy0d6_0(.dout(w_dff_A_qzY6k9bV1_0),.din(w_dff_A_xda3Vy0d6_0),.clk(gclk));
	jdff dff_A_qzY6k9bV1_0(.dout(w_dff_A_LmZ0mUY13_0),.din(w_dff_A_qzY6k9bV1_0),.clk(gclk));
	jdff dff_A_LmZ0mUY13_0(.dout(w_dff_A_itLtmvNN7_0),.din(w_dff_A_LmZ0mUY13_0),.clk(gclk));
	jdff dff_A_itLtmvNN7_0(.dout(w_dff_A_ljAecS813_0),.din(w_dff_A_itLtmvNN7_0),.clk(gclk));
	jdff dff_A_ljAecS813_0(.dout(w_dff_A_xXPOArSh9_0),.din(w_dff_A_ljAecS813_0),.clk(gclk));
	jdff dff_A_xXPOArSh9_0(.dout(w_dff_A_jendyGrO6_0),.din(w_dff_A_xXPOArSh9_0),.clk(gclk));
	jdff dff_A_jendyGrO6_0(.dout(w_dff_A_f7A6Kc5N3_0),.din(w_dff_A_jendyGrO6_0),.clk(gclk));
	jdff dff_A_f7A6Kc5N3_0(.dout(w_dff_A_ZmdUGqAM2_0),.din(w_dff_A_f7A6Kc5N3_0),.clk(gclk));
	jdff dff_A_ZmdUGqAM2_0(.dout(G973),.din(w_dff_A_ZmdUGqAM2_0),.clk(gclk));
	jdff dff_A_x1fDTMpv4_1(.dout(w_dff_A_3eJkcZNv9_0),.din(w_dff_A_x1fDTMpv4_1),.clk(gclk));
	jdff dff_A_3eJkcZNv9_0(.dout(w_dff_A_X9tajY7k8_0),.din(w_dff_A_3eJkcZNv9_0),.clk(gclk));
	jdff dff_A_X9tajY7k8_0(.dout(w_dff_A_xA0mRPKS0_0),.din(w_dff_A_X9tajY7k8_0),.clk(gclk));
	jdff dff_A_xA0mRPKS0_0(.dout(w_dff_A_rLehVRFX3_0),.din(w_dff_A_xA0mRPKS0_0),.clk(gclk));
	jdff dff_A_rLehVRFX3_0(.dout(w_dff_A_etlAf4X79_0),.din(w_dff_A_rLehVRFX3_0),.clk(gclk));
	jdff dff_A_etlAf4X79_0(.dout(w_dff_A_64z72IBX9_0),.din(w_dff_A_etlAf4X79_0),.clk(gclk));
	jdff dff_A_64z72IBX9_0(.dout(w_dff_A_mh6W16JF8_0),.din(w_dff_A_64z72IBX9_0),.clk(gclk));
	jdff dff_A_mh6W16JF8_0(.dout(w_dff_A_Fm2SPi825_0),.din(w_dff_A_mh6W16JF8_0),.clk(gclk));
	jdff dff_A_Fm2SPi825_0(.dout(w_dff_A_Qp7NrPNx3_0),.din(w_dff_A_Fm2SPi825_0),.clk(gclk));
	jdff dff_A_Qp7NrPNx3_0(.dout(w_dff_A_ZJ9sOzGb5_0),.din(w_dff_A_Qp7NrPNx3_0),.clk(gclk));
	jdff dff_A_ZJ9sOzGb5_0(.dout(w_dff_A_oG8MZvNo1_0),.din(w_dff_A_ZJ9sOzGb5_0),.clk(gclk));
	jdff dff_A_oG8MZvNo1_0(.dout(w_dff_A_yguufseH2_0),.din(w_dff_A_oG8MZvNo1_0),.clk(gclk));
	jdff dff_A_yguufseH2_0(.dout(w_dff_A_9yPlCXyn4_0),.din(w_dff_A_yguufseH2_0),.clk(gclk));
	jdff dff_A_9yPlCXyn4_0(.dout(w_dff_A_Yo1dwklH7_0),.din(w_dff_A_9yPlCXyn4_0),.clk(gclk));
	jdff dff_A_Yo1dwklH7_0(.dout(w_dff_A_7BLirZBO5_0),.din(w_dff_A_Yo1dwklH7_0),.clk(gclk));
	jdff dff_A_7BLirZBO5_0(.dout(w_dff_A_oqmu97qb3_0),.din(w_dff_A_7BLirZBO5_0),.clk(gclk));
	jdff dff_A_oqmu97qb3_0(.dout(w_dff_A_MDSAPr0g9_0),.din(w_dff_A_oqmu97qb3_0),.clk(gclk));
	jdff dff_A_MDSAPr0g9_0(.dout(w_dff_A_e3wYAzRF4_0),.din(w_dff_A_MDSAPr0g9_0),.clk(gclk));
	jdff dff_A_e3wYAzRF4_0(.dout(w_dff_A_QoQM8ycS2_0),.din(w_dff_A_e3wYAzRF4_0),.clk(gclk));
	jdff dff_A_QoQM8ycS2_0(.dout(w_dff_A_FMf0Y2x02_0),.din(w_dff_A_QoQM8ycS2_0),.clk(gclk));
	jdff dff_A_FMf0Y2x02_0(.dout(w_dff_A_O69NHFZw0_0),.din(w_dff_A_FMf0Y2x02_0),.clk(gclk));
	jdff dff_A_O69NHFZw0_0(.dout(w_dff_A_EfjyputL3_0),.din(w_dff_A_O69NHFZw0_0),.clk(gclk));
	jdff dff_A_EfjyputL3_0(.dout(w_dff_A_RAJk3tgW3_0),.din(w_dff_A_EfjyputL3_0),.clk(gclk));
	jdff dff_A_RAJk3tgW3_0(.dout(w_dff_A_17NypG9V3_0),.din(w_dff_A_RAJk3tgW3_0),.clk(gclk));
	jdff dff_A_17NypG9V3_0(.dout(G594),.din(w_dff_A_17NypG9V3_0),.clk(gclk));
	jdff dff_A_Md6sOKZ80_1(.dout(w_dff_A_XvKxEYeb3_0),.din(w_dff_A_Md6sOKZ80_1),.clk(gclk));
	jdff dff_A_XvKxEYeb3_0(.dout(w_dff_A_i3XhF68D7_0),.din(w_dff_A_XvKxEYeb3_0),.clk(gclk));
	jdff dff_A_i3XhF68D7_0(.dout(w_dff_A_8xqEaYYx2_0),.din(w_dff_A_i3XhF68D7_0),.clk(gclk));
	jdff dff_A_8xqEaYYx2_0(.dout(w_dff_A_jtvLgiD99_0),.din(w_dff_A_8xqEaYYx2_0),.clk(gclk));
	jdff dff_A_jtvLgiD99_0(.dout(w_dff_A_iXZdZlzp7_0),.din(w_dff_A_jtvLgiD99_0),.clk(gclk));
	jdff dff_A_iXZdZlzp7_0(.dout(w_dff_A_XlzTt09d7_0),.din(w_dff_A_iXZdZlzp7_0),.clk(gclk));
	jdff dff_A_XlzTt09d7_0(.dout(w_dff_A_HktJ1QZd2_0),.din(w_dff_A_XlzTt09d7_0),.clk(gclk));
	jdff dff_A_HktJ1QZd2_0(.dout(w_dff_A_47HNa0811_0),.din(w_dff_A_HktJ1QZd2_0),.clk(gclk));
	jdff dff_A_47HNa0811_0(.dout(w_dff_A_syDUelsQ0_0),.din(w_dff_A_47HNa0811_0),.clk(gclk));
	jdff dff_A_syDUelsQ0_0(.dout(w_dff_A_152ntPtq1_0),.din(w_dff_A_syDUelsQ0_0),.clk(gclk));
	jdff dff_A_152ntPtq1_0(.dout(w_dff_A_IdCc1g4u1_0),.din(w_dff_A_152ntPtq1_0),.clk(gclk));
	jdff dff_A_IdCc1g4u1_0(.dout(w_dff_A_nMrDRXjR8_0),.din(w_dff_A_IdCc1g4u1_0),.clk(gclk));
	jdff dff_A_nMrDRXjR8_0(.dout(w_dff_A_1CQ8pp6U0_0),.din(w_dff_A_nMrDRXjR8_0),.clk(gclk));
	jdff dff_A_1CQ8pp6U0_0(.dout(w_dff_A_b7PLKkUf2_0),.din(w_dff_A_1CQ8pp6U0_0),.clk(gclk));
	jdff dff_A_b7PLKkUf2_0(.dout(w_dff_A_OPoYeikb9_0),.din(w_dff_A_b7PLKkUf2_0),.clk(gclk));
	jdff dff_A_OPoYeikb9_0(.dout(w_dff_A_0lGNWpoZ8_0),.din(w_dff_A_OPoYeikb9_0),.clk(gclk));
	jdff dff_A_0lGNWpoZ8_0(.dout(w_dff_A_orosTVSG8_0),.din(w_dff_A_0lGNWpoZ8_0),.clk(gclk));
	jdff dff_A_orosTVSG8_0(.dout(w_dff_A_Mb4puldy6_0),.din(w_dff_A_orosTVSG8_0),.clk(gclk));
	jdff dff_A_Mb4puldy6_0(.dout(w_dff_A_LRDgmMRD0_0),.din(w_dff_A_Mb4puldy6_0),.clk(gclk));
	jdff dff_A_LRDgmMRD0_0(.dout(w_dff_A_FJsbvNw90_0),.din(w_dff_A_LRDgmMRD0_0),.clk(gclk));
	jdff dff_A_FJsbvNw90_0(.dout(w_dff_A_DQmwjfCt4_0),.din(w_dff_A_FJsbvNw90_0),.clk(gclk));
	jdff dff_A_DQmwjfCt4_0(.dout(w_dff_A_HRGuZvis1_0),.din(w_dff_A_DQmwjfCt4_0),.clk(gclk));
	jdff dff_A_HRGuZvis1_0(.dout(w_dff_A_DCOAnzVo8_0),.din(w_dff_A_HRGuZvis1_0),.clk(gclk));
	jdff dff_A_DCOAnzVo8_0(.dout(w_dff_A_mybCOiNB9_0),.din(w_dff_A_DCOAnzVo8_0),.clk(gclk));
	jdff dff_A_mybCOiNB9_0(.dout(G599),.din(w_dff_A_mybCOiNB9_0),.clk(gclk));
	jdff dff_A_95yRjwe90_1(.dout(w_dff_A_NGnFQ2mj3_0),.din(w_dff_A_95yRjwe90_1),.clk(gclk));
	jdff dff_A_NGnFQ2mj3_0(.dout(w_dff_A_Df8ddHxv7_0),.din(w_dff_A_NGnFQ2mj3_0),.clk(gclk));
	jdff dff_A_Df8ddHxv7_0(.dout(w_dff_A_Q92jIBqk5_0),.din(w_dff_A_Df8ddHxv7_0),.clk(gclk));
	jdff dff_A_Q92jIBqk5_0(.dout(w_dff_A_NKYpk9oX1_0),.din(w_dff_A_Q92jIBqk5_0),.clk(gclk));
	jdff dff_A_NKYpk9oX1_0(.dout(w_dff_A_T0RH3nWO7_0),.din(w_dff_A_NKYpk9oX1_0),.clk(gclk));
	jdff dff_A_T0RH3nWO7_0(.dout(w_dff_A_zalk2Z9V1_0),.din(w_dff_A_T0RH3nWO7_0),.clk(gclk));
	jdff dff_A_zalk2Z9V1_0(.dout(w_dff_A_lpdgsik56_0),.din(w_dff_A_zalk2Z9V1_0),.clk(gclk));
	jdff dff_A_lpdgsik56_0(.dout(w_dff_A_YZTgR7Uj7_0),.din(w_dff_A_lpdgsik56_0),.clk(gclk));
	jdff dff_A_YZTgR7Uj7_0(.dout(w_dff_A_ZDRfD1Ay2_0),.din(w_dff_A_YZTgR7Uj7_0),.clk(gclk));
	jdff dff_A_ZDRfD1Ay2_0(.dout(w_dff_A_PNqNJOAs8_0),.din(w_dff_A_ZDRfD1Ay2_0),.clk(gclk));
	jdff dff_A_PNqNJOAs8_0(.dout(w_dff_A_kkFJ5V7M9_0),.din(w_dff_A_PNqNJOAs8_0),.clk(gclk));
	jdff dff_A_kkFJ5V7M9_0(.dout(w_dff_A_rEzTzose3_0),.din(w_dff_A_kkFJ5V7M9_0),.clk(gclk));
	jdff dff_A_rEzTzose3_0(.dout(w_dff_A_ONqr2cy19_0),.din(w_dff_A_rEzTzose3_0),.clk(gclk));
	jdff dff_A_ONqr2cy19_0(.dout(w_dff_A_K1mUvgZK7_0),.din(w_dff_A_ONqr2cy19_0),.clk(gclk));
	jdff dff_A_K1mUvgZK7_0(.dout(w_dff_A_hHnvlRYC9_0),.din(w_dff_A_K1mUvgZK7_0),.clk(gclk));
	jdff dff_A_hHnvlRYC9_0(.dout(w_dff_A_fKJnZX4L7_0),.din(w_dff_A_hHnvlRYC9_0),.clk(gclk));
	jdff dff_A_fKJnZX4L7_0(.dout(w_dff_A_DpPOdRXR4_0),.din(w_dff_A_fKJnZX4L7_0),.clk(gclk));
	jdff dff_A_DpPOdRXR4_0(.dout(w_dff_A_QpbcdHhU9_0),.din(w_dff_A_DpPOdRXR4_0),.clk(gclk));
	jdff dff_A_QpbcdHhU9_0(.dout(w_dff_A_0Jh4CTBc1_0),.din(w_dff_A_QpbcdHhU9_0),.clk(gclk));
	jdff dff_A_0Jh4CTBc1_0(.dout(w_dff_A_stYB7YaL3_0),.din(w_dff_A_0Jh4CTBc1_0),.clk(gclk));
	jdff dff_A_stYB7YaL3_0(.dout(w_dff_A_AGBLizWo8_0),.din(w_dff_A_stYB7YaL3_0),.clk(gclk));
	jdff dff_A_AGBLizWo8_0(.dout(w_dff_A_pK6j8JNo6_0),.din(w_dff_A_AGBLizWo8_0),.clk(gclk));
	jdff dff_A_pK6j8JNo6_0(.dout(w_dff_A_L1JQmsCW1_0),.din(w_dff_A_pK6j8JNo6_0),.clk(gclk));
	jdff dff_A_L1JQmsCW1_0(.dout(w_dff_A_xTZ1dCBt8_0),.din(w_dff_A_L1JQmsCW1_0),.clk(gclk));
	jdff dff_A_xTZ1dCBt8_0(.dout(G600),.din(w_dff_A_xTZ1dCBt8_0),.clk(gclk));
	jdff dff_A_AtXnEyBC7_1(.dout(w_dff_A_FouQWFaB4_0),.din(w_dff_A_AtXnEyBC7_1),.clk(gclk));
	jdff dff_A_FouQWFaB4_0(.dout(w_dff_A_5ZHZUS7M6_0),.din(w_dff_A_FouQWFaB4_0),.clk(gclk));
	jdff dff_A_5ZHZUS7M6_0(.dout(w_dff_A_GmgpDGDR2_0),.din(w_dff_A_5ZHZUS7M6_0),.clk(gclk));
	jdff dff_A_GmgpDGDR2_0(.dout(w_dff_A_PriqH0wm6_0),.din(w_dff_A_GmgpDGDR2_0),.clk(gclk));
	jdff dff_A_PriqH0wm6_0(.dout(w_dff_A_sMmzXXj41_0),.din(w_dff_A_PriqH0wm6_0),.clk(gclk));
	jdff dff_A_sMmzXXj41_0(.dout(w_dff_A_Wl47g9D92_0),.din(w_dff_A_sMmzXXj41_0),.clk(gclk));
	jdff dff_A_Wl47g9D92_0(.dout(w_dff_A_pu988qNr8_0),.din(w_dff_A_Wl47g9D92_0),.clk(gclk));
	jdff dff_A_pu988qNr8_0(.dout(w_dff_A_TiDgNwFx9_0),.din(w_dff_A_pu988qNr8_0),.clk(gclk));
	jdff dff_A_TiDgNwFx9_0(.dout(w_dff_A_qfXhWJqT3_0),.din(w_dff_A_TiDgNwFx9_0),.clk(gclk));
	jdff dff_A_qfXhWJqT3_0(.dout(w_dff_A_ucyWdUIR6_0),.din(w_dff_A_qfXhWJqT3_0),.clk(gclk));
	jdff dff_A_ucyWdUIR6_0(.dout(w_dff_A_e59Izlyj0_0),.din(w_dff_A_ucyWdUIR6_0),.clk(gclk));
	jdff dff_A_e59Izlyj0_0(.dout(w_dff_A_NCxwK95s0_0),.din(w_dff_A_e59Izlyj0_0),.clk(gclk));
	jdff dff_A_NCxwK95s0_0(.dout(w_dff_A_EHU2iTZ85_0),.din(w_dff_A_NCxwK95s0_0),.clk(gclk));
	jdff dff_A_EHU2iTZ85_0(.dout(w_dff_A_I3LmKJ0a0_0),.din(w_dff_A_EHU2iTZ85_0),.clk(gclk));
	jdff dff_A_I3LmKJ0a0_0(.dout(w_dff_A_RGgYilYt3_0),.din(w_dff_A_I3LmKJ0a0_0),.clk(gclk));
	jdff dff_A_RGgYilYt3_0(.dout(w_dff_A_jYc7f8nn5_0),.din(w_dff_A_RGgYilYt3_0),.clk(gclk));
	jdff dff_A_jYc7f8nn5_0(.dout(w_dff_A_Jo20Jtiw2_0),.din(w_dff_A_jYc7f8nn5_0),.clk(gclk));
	jdff dff_A_Jo20Jtiw2_0(.dout(w_dff_A_uoq4Zv620_0),.din(w_dff_A_Jo20Jtiw2_0),.clk(gclk));
	jdff dff_A_uoq4Zv620_0(.dout(w_dff_A_dhqS9DYw0_0),.din(w_dff_A_uoq4Zv620_0),.clk(gclk));
	jdff dff_A_dhqS9DYw0_0(.dout(w_dff_A_1EcuuRWd2_0),.din(w_dff_A_dhqS9DYw0_0),.clk(gclk));
	jdff dff_A_1EcuuRWd2_0(.dout(w_dff_A_tqaP1fcJ2_0),.din(w_dff_A_1EcuuRWd2_0),.clk(gclk));
	jdff dff_A_tqaP1fcJ2_0(.dout(w_dff_A_T6cWsFWg9_0),.din(w_dff_A_tqaP1fcJ2_0),.clk(gclk));
	jdff dff_A_T6cWsFWg9_0(.dout(w_dff_A_PFp8LOMS9_0),.din(w_dff_A_T6cWsFWg9_0),.clk(gclk));
	jdff dff_A_PFp8LOMS9_0(.dout(w_dff_A_eIIO9z1t3_0),.din(w_dff_A_PFp8LOMS9_0),.clk(gclk));
	jdff dff_A_eIIO9z1t3_0(.dout(G601),.din(w_dff_A_eIIO9z1t3_0),.clk(gclk));
	jdff dff_A_d5oFxJLf5_1(.dout(w_dff_A_quqgr5Ep4_0),.din(w_dff_A_d5oFxJLf5_1),.clk(gclk));
	jdff dff_A_quqgr5Ep4_0(.dout(w_dff_A_nDQWTRPm9_0),.din(w_dff_A_quqgr5Ep4_0),.clk(gclk));
	jdff dff_A_nDQWTRPm9_0(.dout(w_dff_A_IXPg4fPj5_0),.din(w_dff_A_nDQWTRPm9_0),.clk(gclk));
	jdff dff_A_IXPg4fPj5_0(.dout(w_dff_A_OT9aXnPz7_0),.din(w_dff_A_IXPg4fPj5_0),.clk(gclk));
	jdff dff_A_OT9aXnPz7_0(.dout(w_dff_A_bgBFMxfz9_0),.din(w_dff_A_OT9aXnPz7_0),.clk(gclk));
	jdff dff_A_bgBFMxfz9_0(.dout(w_dff_A_1CRCRvHU6_0),.din(w_dff_A_bgBFMxfz9_0),.clk(gclk));
	jdff dff_A_1CRCRvHU6_0(.dout(w_dff_A_4dYcBy0D5_0),.din(w_dff_A_1CRCRvHU6_0),.clk(gclk));
	jdff dff_A_4dYcBy0D5_0(.dout(w_dff_A_YZE2bGGd5_0),.din(w_dff_A_4dYcBy0D5_0),.clk(gclk));
	jdff dff_A_YZE2bGGd5_0(.dout(w_dff_A_Gf0si6rP2_0),.din(w_dff_A_YZE2bGGd5_0),.clk(gclk));
	jdff dff_A_Gf0si6rP2_0(.dout(w_dff_A_pu2G6fmg5_0),.din(w_dff_A_Gf0si6rP2_0),.clk(gclk));
	jdff dff_A_pu2G6fmg5_0(.dout(w_dff_A_y2EVG8CJ1_0),.din(w_dff_A_pu2G6fmg5_0),.clk(gclk));
	jdff dff_A_y2EVG8CJ1_0(.dout(w_dff_A_1H3gRmuE6_0),.din(w_dff_A_y2EVG8CJ1_0),.clk(gclk));
	jdff dff_A_1H3gRmuE6_0(.dout(w_dff_A_uLkpO3pV7_0),.din(w_dff_A_1H3gRmuE6_0),.clk(gclk));
	jdff dff_A_uLkpO3pV7_0(.dout(w_dff_A_rAJ53Wdx1_0),.din(w_dff_A_uLkpO3pV7_0),.clk(gclk));
	jdff dff_A_rAJ53Wdx1_0(.dout(w_dff_A_0HpOOd7h2_0),.din(w_dff_A_rAJ53Wdx1_0),.clk(gclk));
	jdff dff_A_0HpOOd7h2_0(.dout(w_dff_A_T8Kb0OIX8_0),.din(w_dff_A_0HpOOd7h2_0),.clk(gclk));
	jdff dff_A_T8Kb0OIX8_0(.dout(w_dff_A_scDPLGRk8_0),.din(w_dff_A_T8Kb0OIX8_0),.clk(gclk));
	jdff dff_A_scDPLGRk8_0(.dout(w_dff_A_7RWBD3Em3_0),.din(w_dff_A_scDPLGRk8_0),.clk(gclk));
	jdff dff_A_7RWBD3Em3_0(.dout(w_dff_A_AsPJgWuK7_0),.din(w_dff_A_7RWBD3Em3_0),.clk(gclk));
	jdff dff_A_AsPJgWuK7_0(.dout(w_dff_A_quc44TPB0_0),.din(w_dff_A_AsPJgWuK7_0),.clk(gclk));
	jdff dff_A_quc44TPB0_0(.dout(w_dff_A_YG3pGkx39_0),.din(w_dff_A_quc44TPB0_0),.clk(gclk));
	jdff dff_A_YG3pGkx39_0(.dout(w_dff_A_Q0csuqQ08_0),.din(w_dff_A_YG3pGkx39_0),.clk(gclk));
	jdff dff_A_Q0csuqQ08_0(.dout(w_dff_A_MEDAvAne0_0),.din(w_dff_A_Q0csuqQ08_0),.clk(gclk));
	jdff dff_A_MEDAvAne0_0(.dout(w_dff_A_YbC1Kx7X5_0),.din(w_dff_A_MEDAvAne0_0),.clk(gclk));
	jdff dff_A_YbC1Kx7X5_0(.dout(G602),.din(w_dff_A_YbC1Kx7X5_0),.clk(gclk));
	jdff dff_A_psklSFAO5_1(.dout(w_dff_A_syrspiJb8_0),.din(w_dff_A_psklSFAO5_1),.clk(gclk));
	jdff dff_A_syrspiJb8_0(.dout(w_dff_A_XSH3hame1_0),.din(w_dff_A_syrspiJb8_0),.clk(gclk));
	jdff dff_A_XSH3hame1_0(.dout(w_dff_A_K8z4jh8m4_0),.din(w_dff_A_XSH3hame1_0),.clk(gclk));
	jdff dff_A_K8z4jh8m4_0(.dout(w_dff_A_LLaQKBrF0_0),.din(w_dff_A_K8z4jh8m4_0),.clk(gclk));
	jdff dff_A_LLaQKBrF0_0(.dout(w_dff_A_eu9UKrS33_0),.din(w_dff_A_LLaQKBrF0_0),.clk(gclk));
	jdff dff_A_eu9UKrS33_0(.dout(w_dff_A_N57dancA2_0),.din(w_dff_A_eu9UKrS33_0),.clk(gclk));
	jdff dff_A_N57dancA2_0(.dout(w_dff_A_Xb1Xrrqc1_0),.din(w_dff_A_N57dancA2_0),.clk(gclk));
	jdff dff_A_Xb1Xrrqc1_0(.dout(w_dff_A_8byz53nP5_0),.din(w_dff_A_Xb1Xrrqc1_0),.clk(gclk));
	jdff dff_A_8byz53nP5_0(.dout(w_dff_A_ylQtX0ZS3_0),.din(w_dff_A_8byz53nP5_0),.clk(gclk));
	jdff dff_A_ylQtX0ZS3_0(.dout(w_dff_A_YZHKLBLI0_0),.din(w_dff_A_ylQtX0ZS3_0),.clk(gclk));
	jdff dff_A_YZHKLBLI0_0(.dout(w_dff_A_A0PZnddb2_0),.din(w_dff_A_YZHKLBLI0_0),.clk(gclk));
	jdff dff_A_A0PZnddb2_0(.dout(w_dff_A_3MCGZOZF1_0),.din(w_dff_A_A0PZnddb2_0),.clk(gclk));
	jdff dff_A_3MCGZOZF1_0(.dout(w_dff_A_9UjTvXEI2_0),.din(w_dff_A_3MCGZOZF1_0),.clk(gclk));
	jdff dff_A_9UjTvXEI2_0(.dout(w_dff_A_yx2royOW5_0),.din(w_dff_A_9UjTvXEI2_0),.clk(gclk));
	jdff dff_A_yx2royOW5_0(.dout(w_dff_A_5ommu2eA0_0),.din(w_dff_A_yx2royOW5_0),.clk(gclk));
	jdff dff_A_5ommu2eA0_0(.dout(w_dff_A_IdFX6uti6_0),.din(w_dff_A_5ommu2eA0_0),.clk(gclk));
	jdff dff_A_IdFX6uti6_0(.dout(w_dff_A_KoxbzP5h4_0),.din(w_dff_A_IdFX6uti6_0),.clk(gclk));
	jdff dff_A_KoxbzP5h4_0(.dout(w_dff_A_eOMRKb965_0),.din(w_dff_A_KoxbzP5h4_0),.clk(gclk));
	jdff dff_A_eOMRKb965_0(.dout(w_dff_A_UcSv1Yyw5_0),.din(w_dff_A_eOMRKb965_0),.clk(gclk));
	jdff dff_A_UcSv1Yyw5_0(.dout(w_dff_A_HMmeEGFG3_0),.din(w_dff_A_UcSv1Yyw5_0),.clk(gclk));
	jdff dff_A_HMmeEGFG3_0(.dout(w_dff_A_MX8T0eGB3_0),.din(w_dff_A_HMmeEGFG3_0),.clk(gclk));
	jdff dff_A_MX8T0eGB3_0(.dout(w_dff_A_cq4jRdSq2_0),.din(w_dff_A_MX8T0eGB3_0),.clk(gclk));
	jdff dff_A_cq4jRdSq2_0(.dout(w_dff_A_pvGf9Poj9_0),.din(w_dff_A_cq4jRdSq2_0),.clk(gclk));
	jdff dff_A_pvGf9Poj9_0(.dout(w_dff_A_1L88bpv31_0),.din(w_dff_A_pvGf9Poj9_0),.clk(gclk));
	jdff dff_A_1L88bpv31_0(.dout(G603),.din(w_dff_A_1L88bpv31_0),.clk(gclk));
	jdff dff_A_TwNsD2rL2_1(.dout(w_dff_A_zLtiV7Hl9_0),.din(w_dff_A_TwNsD2rL2_1),.clk(gclk));
	jdff dff_A_zLtiV7Hl9_0(.dout(w_dff_A_duLohmMZ1_0),.din(w_dff_A_zLtiV7Hl9_0),.clk(gclk));
	jdff dff_A_duLohmMZ1_0(.dout(w_dff_A_hjWfbfeb6_0),.din(w_dff_A_duLohmMZ1_0),.clk(gclk));
	jdff dff_A_hjWfbfeb6_0(.dout(w_dff_A_OSSPYYo76_0),.din(w_dff_A_hjWfbfeb6_0),.clk(gclk));
	jdff dff_A_OSSPYYo76_0(.dout(w_dff_A_E6ZTtMGZ3_0),.din(w_dff_A_OSSPYYo76_0),.clk(gclk));
	jdff dff_A_E6ZTtMGZ3_0(.dout(w_dff_A_0IPypipt7_0),.din(w_dff_A_E6ZTtMGZ3_0),.clk(gclk));
	jdff dff_A_0IPypipt7_0(.dout(w_dff_A_Z2xrnaVM5_0),.din(w_dff_A_0IPypipt7_0),.clk(gclk));
	jdff dff_A_Z2xrnaVM5_0(.dout(w_dff_A_Hg0nen860_0),.din(w_dff_A_Z2xrnaVM5_0),.clk(gclk));
	jdff dff_A_Hg0nen860_0(.dout(w_dff_A_XDf9c3wR6_0),.din(w_dff_A_Hg0nen860_0),.clk(gclk));
	jdff dff_A_XDf9c3wR6_0(.dout(w_dff_A_buoU9x751_0),.din(w_dff_A_XDf9c3wR6_0),.clk(gclk));
	jdff dff_A_buoU9x751_0(.dout(w_dff_A_h7ZSJErN6_0),.din(w_dff_A_buoU9x751_0),.clk(gclk));
	jdff dff_A_h7ZSJErN6_0(.dout(w_dff_A_g9BseHpq7_0),.din(w_dff_A_h7ZSJErN6_0),.clk(gclk));
	jdff dff_A_g9BseHpq7_0(.dout(w_dff_A_7xrpUrne1_0),.din(w_dff_A_g9BseHpq7_0),.clk(gclk));
	jdff dff_A_7xrpUrne1_0(.dout(w_dff_A_DZ7eClga0_0),.din(w_dff_A_7xrpUrne1_0),.clk(gclk));
	jdff dff_A_DZ7eClga0_0(.dout(w_dff_A_gWzVaXk65_0),.din(w_dff_A_DZ7eClga0_0),.clk(gclk));
	jdff dff_A_gWzVaXk65_0(.dout(w_dff_A_KZcGxfVS7_0),.din(w_dff_A_gWzVaXk65_0),.clk(gclk));
	jdff dff_A_KZcGxfVS7_0(.dout(w_dff_A_dv9B6CSK3_0),.din(w_dff_A_KZcGxfVS7_0),.clk(gclk));
	jdff dff_A_dv9B6CSK3_0(.dout(w_dff_A_LajfI1038_0),.din(w_dff_A_dv9B6CSK3_0),.clk(gclk));
	jdff dff_A_LajfI1038_0(.dout(w_dff_A_QeLeoSHx3_0),.din(w_dff_A_LajfI1038_0),.clk(gclk));
	jdff dff_A_QeLeoSHx3_0(.dout(w_dff_A_bPIA2cJk9_0),.din(w_dff_A_QeLeoSHx3_0),.clk(gclk));
	jdff dff_A_bPIA2cJk9_0(.dout(w_dff_A_CgEWVihV8_0),.din(w_dff_A_bPIA2cJk9_0),.clk(gclk));
	jdff dff_A_CgEWVihV8_0(.dout(w_dff_A_KflzC4fR3_0),.din(w_dff_A_CgEWVihV8_0),.clk(gclk));
	jdff dff_A_KflzC4fR3_0(.dout(w_dff_A_n19JPVCU6_0),.din(w_dff_A_KflzC4fR3_0),.clk(gclk));
	jdff dff_A_n19JPVCU6_0(.dout(w_dff_A_Egpwz42Y4_0),.din(w_dff_A_n19JPVCU6_0),.clk(gclk));
	jdff dff_A_Egpwz42Y4_0(.dout(G604),.din(w_dff_A_Egpwz42Y4_0),.clk(gclk));
	jdff dff_A_g9Y6z9mT9_1(.dout(w_dff_A_xoVR1WGa0_0),.din(w_dff_A_g9Y6z9mT9_1),.clk(gclk));
	jdff dff_A_xoVR1WGa0_0(.dout(w_dff_A_GbRR1pC52_0),.din(w_dff_A_xoVR1WGa0_0),.clk(gclk));
	jdff dff_A_GbRR1pC52_0(.dout(w_dff_A_SRYHYUhx9_0),.din(w_dff_A_GbRR1pC52_0),.clk(gclk));
	jdff dff_A_SRYHYUhx9_0(.dout(w_dff_A_2Bze2Tpt1_0),.din(w_dff_A_SRYHYUhx9_0),.clk(gclk));
	jdff dff_A_2Bze2Tpt1_0(.dout(w_dff_A_8qPQBUGx5_0),.din(w_dff_A_2Bze2Tpt1_0),.clk(gclk));
	jdff dff_A_8qPQBUGx5_0(.dout(w_dff_A_Anzu2NlP5_0),.din(w_dff_A_8qPQBUGx5_0),.clk(gclk));
	jdff dff_A_Anzu2NlP5_0(.dout(w_dff_A_Og5HVl4t3_0),.din(w_dff_A_Anzu2NlP5_0),.clk(gclk));
	jdff dff_A_Og5HVl4t3_0(.dout(w_dff_A_RKVFx3rx9_0),.din(w_dff_A_Og5HVl4t3_0),.clk(gclk));
	jdff dff_A_RKVFx3rx9_0(.dout(w_dff_A_oKhytRBm2_0),.din(w_dff_A_RKVFx3rx9_0),.clk(gclk));
	jdff dff_A_oKhytRBm2_0(.dout(w_dff_A_cj2SuduW6_0),.din(w_dff_A_oKhytRBm2_0),.clk(gclk));
	jdff dff_A_cj2SuduW6_0(.dout(w_dff_A_VAivyzf87_0),.din(w_dff_A_cj2SuduW6_0),.clk(gclk));
	jdff dff_A_VAivyzf87_0(.dout(w_dff_A_uP6xiXyD9_0),.din(w_dff_A_VAivyzf87_0),.clk(gclk));
	jdff dff_A_uP6xiXyD9_0(.dout(w_dff_A_nEF9ZX820_0),.din(w_dff_A_uP6xiXyD9_0),.clk(gclk));
	jdff dff_A_nEF9ZX820_0(.dout(w_dff_A_Y9Y79gPP0_0),.din(w_dff_A_nEF9ZX820_0),.clk(gclk));
	jdff dff_A_Y9Y79gPP0_0(.dout(w_dff_A_bA9IK4OQ6_0),.din(w_dff_A_Y9Y79gPP0_0),.clk(gclk));
	jdff dff_A_bA9IK4OQ6_0(.dout(w_dff_A_qR2bPC1j4_0),.din(w_dff_A_bA9IK4OQ6_0),.clk(gclk));
	jdff dff_A_qR2bPC1j4_0(.dout(w_dff_A_j646Whri1_0),.din(w_dff_A_qR2bPC1j4_0),.clk(gclk));
	jdff dff_A_j646Whri1_0(.dout(w_dff_A_9ekTT3Ee1_0),.din(w_dff_A_j646Whri1_0),.clk(gclk));
	jdff dff_A_9ekTT3Ee1_0(.dout(w_dff_A_CTxqaQiW0_0),.din(w_dff_A_9ekTT3Ee1_0),.clk(gclk));
	jdff dff_A_CTxqaQiW0_0(.dout(w_dff_A_9eDpmNFz8_0),.din(w_dff_A_CTxqaQiW0_0),.clk(gclk));
	jdff dff_A_9eDpmNFz8_0(.dout(w_dff_A_ArXhC84a1_0),.din(w_dff_A_9eDpmNFz8_0),.clk(gclk));
	jdff dff_A_ArXhC84a1_0(.dout(w_dff_A_FUPUOTjR9_0),.din(w_dff_A_ArXhC84a1_0),.clk(gclk));
	jdff dff_A_FUPUOTjR9_0(.dout(w_dff_A_K8MWOyGH7_0),.din(w_dff_A_FUPUOTjR9_0),.clk(gclk));
	jdff dff_A_K8MWOyGH7_0(.dout(w_dff_A_zQTFQxmk5_0),.din(w_dff_A_K8MWOyGH7_0),.clk(gclk));
	jdff dff_A_zQTFQxmk5_0(.dout(G611),.din(w_dff_A_zQTFQxmk5_0),.clk(gclk));
	jdff dff_A_wMjzKV3T2_1(.dout(w_dff_A_gmVc3HeH7_0),.din(w_dff_A_wMjzKV3T2_1),.clk(gclk));
	jdff dff_A_gmVc3HeH7_0(.dout(w_dff_A_YPmVzXo50_0),.din(w_dff_A_gmVc3HeH7_0),.clk(gclk));
	jdff dff_A_YPmVzXo50_0(.dout(w_dff_A_xqcHp5R21_0),.din(w_dff_A_YPmVzXo50_0),.clk(gclk));
	jdff dff_A_xqcHp5R21_0(.dout(w_dff_A_rVueodNB8_0),.din(w_dff_A_xqcHp5R21_0),.clk(gclk));
	jdff dff_A_rVueodNB8_0(.dout(w_dff_A_eHzjibSc4_0),.din(w_dff_A_rVueodNB8_0),.clk(gclk));
	jdff dff_A_eHzjibSc4_0(.dout(w_dff_A_5uZGPdgs1_0),.din(w_dff_A_eHzjibSc4_0),.clk(gclk));
	jdff dff_A_5uZGPdgs1_0(.dout(w_dff_A_HRzcRnuI6_0),.din(w_dff_A_5uZGPdgs1_0),.clk(gclk));
	jdff dff_A_HRzcRnuI6_0(.dout(w_dff_A_rLCtRtjC3_0),.din(w_dff_A_HRzcRnuI6_0),.clk(gclk));
	jdff dff_A_rLCtRtjC3_0(.dout(w_dff_A_XwsGc7vW0_0),.din(w_dff_A_rLCtRtjC3_0),.clk(gclk));
	jdff dff_A_XwsGc7vW0_0(.dout(w_dff_A_K6oDWatf0_0),.din(w_dff_A_XwsGc7vW0_0),.clk(gclk));
	jdff dff_A_K6oDWatf0_0(.dout(w_dff_A_Rshwbgwf2_0),.din(w_dff_A_K6oDWatf0_0),.clk(gclk));
	jdff dff_A_Rshwbgwf2_0(.dout(w_dff_A_QR3LTFu02_0),.din(w_dff_A_Rshwbgwf2_0),.clk(gclk));
	jdff dff_A_QR3LTFu02_0(.dout(w_dff_A_WBggRGbi8_0),.din(w_dff_A_QR3LTFu02_0),.clk(gclk));
	jdff dff_A_WBggRGbi8_0(.dout(w_dff_A_OeeRPS5c6_0),.din(w_dff_A_WBggRGbi8_0),.clk(gclk));
	jdff dff_A_OeeRPS5c6_0(.dout(w_dff_A_ZONYte9y6_0),.din(w_dff_A_OeeRPS5c6_0),.clk(gclk));
	jdff dff_A_ZONYte9y6_0(.dout(w_dff_A_V31Tc6V30_0),.din(w_dff_A_ZONYte9y6_0),.clk(gclk));
	jdff dff_A_V31Tc6V30_0(.dout(w_dff_A_H93WLYsM3_0),.din(w_dff_A_V31Tc6V30_0),.clk(gclk));
	jdff dff_A_H93WLYsM3_0(.dout(w_dff_A_xwm1JBI16_0),.din(w_dff_A_H93WLYsM3_0),.clk(gclk));
	jdff dff_A_xwm1JBI16_0(.dout(w_dff_A_Zx9bzyRT9_0),.din(w_dff_A_xwm1JBI16_0),.clk(gclk));
	jdff dff_A_Zx9bzyRT9_0(.dout(w_dff_A_zo4VTCwN4_0),.din(w_dff_A_Zx9bzyRT9_0),.clk(gclk));
	jdff dff_A_zo4VTCwN4_0(.dout(w_dff_A_TwlQBUXs8_0),.din(w_dff_A_zo4VTCwN4_0),.clk(gclk));
	jdff dff_A_TwlQBUXs8_0(.dout(w_dff_A_5ZZaC6uo4_0),.din(w_dff_A_TwlQBUXs8_0),.clk(gclk));
	jdff dff_A_5ZZaC6uo4_0(.dout(w_dff_A_ZcXqDxnv5_0),.din(w_dff_A_5ZZaC6uo4_0),.clk(gclk));
	jdff dff_A_ZcXqDxnv5_0(.dout(w_dff_A_uxhrSHau9_0),.din(w_dff_A_ZcXqDxnv5_0),.clk(gclk));
	jdff dff_A_uxhrSHau9_0(.dout(G612),.din(w_dff_A_uxhrSHau9_0),.clk(gclk));
	jdff dff_A_ngmk1eik7_2(.dout(w_dff_A_rCDjaHpI3_0),.din(w_dff_A_ngmk1eik7_2),.clk(gclk));
	jdff dff_A_rCDjaHpI3_0(.dout(w_dff_A_8Fp46olI2_0),.din(w_dff_A_rCDjaHpI3_0),.clk(gclk));
	jdff dff_A_8Fp46olI2_0(.dout(w_dff_A_D00HEcCH4_0),.din(w_dff_A_8Fp46olI2_0),.clk(gclk));
	jdff dff_A_D00HEcCH4_0(.dout(w_dff_A_gH1Kf8c15_0),.din(w_dff_A_D00HEcCH4_0),.clk(gclk));
	jdff dff_A_gH1Kf8c15_0(.dout(w_dff_A_8KpQHMKD2_0),.din(w_dff_A_gH1Kf8c15_0),.clk(gclk));
	jdff dff_A_8KpQHMKD2_0(.dout(w_dff_A_VLlphInN5_0),.din(w_dff_A_8KpQHMKD2_0),.clk(gclk));
	jdff dff_A_VLlphInN5_0(.dout(w_dff_A_sEYst0N12_0),.din(w_dff_A_VLlphInN5_0),.clk(gclk));
	jdff dff_A_sEYst0N12_0(.dout(w_dff_A_oDNmbRjH9_0),.din(w_dff_A_sEYst0N12_0),.clk(gclk));
	jdff dff_A_oDNmbRjH9_0(.dout(w_dff_A_ZnmBmKwa8_0),.din(w_dff_A_oDNmbRjH9_0),.clk(gclk));
	jdff dff_A_ZnmBmKwa8_0(.dout(w_dff_A_dpsqOQpb0_0),.din(w_dff_A_ZnmBmKwa8_0),.clk(gclk));
	jdff dff_A_dpsqOQpb0_0(.dout(w_dff_A_OjUtfoEE1_0),.din(w_dff_A_dpsqOQpb0_0),.clk(gclk));
	jdff dff_A_OjUtfoEE1_0(.dout(w_dff_A_9BfVnHtw1_0),.din(w_dff_A_OjUtfoEE1_0),.clk(gclk));
	jdff dff_A_9BfVnHtw1_0(.dout(w_dff_A_QQFFRuzS3_0),.din(w_dff_A_9BfVnHtw1_0),.clk(gclk));
	jdff dff_A_QQFFRuzS3_0(.dout(w_dff_A_px73EUeB5_0),.din(w_dff_A_QQFFRuzS3_0),.clk(gclk));
	jdff dff_A_px73EUeB5_0(.dout(w_dff_A_M5txvtd66_0),.din(w_dff_A_px73EUeB5_0),.clk(gclk));
	jdff dff_A_M5txvtd66_0(.dout(w_dff_A_haqALR7a5_0),.din(w_dff_A_M5txvtd66_0),.clk(gclk));
	jdff dff_A_haqALR7a5_0(.dout(w_dff_A_GMIVcFp51_0),.din(w_dff_A_haqALR7a5_0),.clk(gclk));
	jdff dff_A_GMIVcFp51_0(.dout(w_dff_A_VthD3EiR5_0),.din(w_dff_A_GMIVcFp51_0),.clk(gclk));
	jdff dff_A_VthD3EiR5_0(.dout(w_dff_A_Qo5xvpQj6_0),.din(w_dff_A_VthD3EiR5_0),.clk(gclk));
	jdff dff_A_Qo5xvpQj6_0(.dout(w_dff_A_b2JQRBmH9_0),.din(w_dff_A_Qo5xvpQj6_0),.clk(gclk));
	jdff dff_A_b2JQRBmH9_0(.dout(w_dff_A_ifWuJqJ83_0),.din(w_dff_A_b2JQRBmH9_0),.clk(gclk));
	jdff dff_A_ifWuJqJ83_0(.dout(w_dff_A_Zz5O4hms8_0),.din(w_dff_A_ifWuJqJ83_0),.clk(gclk));
	jdff dff_A_Zz5O4hms8_0(.dout(w_dff_A_3QCPLwDI3_0),.din(w_dff_A_Zz5O4hms8_0),.clk(gclk));
	jdff dff_A_3QCPLwDI3_0(.dout(w_dff_A_nNDblEMt0_0),.din(w_dff_A_3QCPLwDI3_0),.clk(gclk));
	jdff dff_A_nNDblEMt0_0(.dout(G810),.din(w_dff_A_nNDblEMt0_0),.clk(gclk));
	jdff dff_A_WaFIGnAa9_1(.dout(w_dff_A_93k3q9BE5_0),.din(w_dff_A_WaFIGnAa9_1),.clk(gclk));
	jdff dff_A_93k3q9BE5_0(.dout(w_dff_A_9hnNWfb10_0),.din(w_dff_A_93k3q9BE5_0),.clk(gclk));
	jdff dff_A_9hnNWfb10_0(.dout(w_dff_A_2sykZE7m1_0),.din(w_dff_A_9hnNWfb10_0),.clk(gclk));
	jdff dff_A_2sykZE7m1_0(.dout(w_dff_A_rNgubPbI6_0),.din(w_dff_A_2sykZE7m1_0),.clk(gclk));
	jdff dff_A_rNgubPbI6_0(.dout(w_dff_A_iVnlT7Q32_0),.din(w_dff_A_rNgubPbI6_0),.clk(gclk));
	jdff dff_A_iVnlT7Q32_0(.dout(w_dff_A_c9kx7tNO6_0),.din(w_dff_A_iVnlT7Q32_0),.clk(gclk));
	jdff dff_A_c9kx7tNO6_0(.dout(w_dff_A_SOLqzsQl7_0),.din(w_dff_A_c9kx7tNO6_0),.clk(gclk));
	jdff dff_A_SOLqzsQl7_0(.dout(w_dff_A_d7pt807o9_0),.din(w_dff_A_SOLqzsQl7_0),.clk(gclk));
	jdff dff_A_d7pt807o9_0(.dout(w_dff_A_ooIhtFkB7_0),.din(w_dff_A_d7pt807o9_0),.clk(gclk));
	jdff dff_A_ooIhtFkB7_0(.dout(w_dff_A_nZQSRnHI9_0),.din(w_dff_A_ooIhtFkB7_0),.clk(gclk));
	jdff dff_A_nZQSRnHI9_0(.dout(w_dff_A_QxlC37c31_0),.din(w_dff_A_nZQSRnHI9_0),.clk(gclk));
	jdff dff_A_QxlC37c31_0(.dout(w_dff_A_nJjLr0CU5_0),.din(w_dff_A_QxlC37c31_0),.clk(gclk));
	jdff dff_A_nJjLr0CU5_0(.dout(w_dff_A_tjkX94Uo2_0),.din(w_dff_A_nJjLr0CU5_0),.clk(gclk));
	jdff dff_A_tjkX94Uo2_0(.dout(w_dff_A_4ncXZcSP6_0),.din(w_dff_A_tjkX94Uo2_0),.clk(gclk));
	jdff dff_A_4ncXZcSP6_0(.dout(w_dff_A_ul7MAnSa8_0),.din(w_dff_A_4ncXZcSP6_0),.clk(gclk));
	jdff dff_A_ul7MAnSa8_0(.dout(w_dff_A_A9lO3CyH0_0),.din(w_dff_A_ul7MAnSa8_0),.clk(gclk));
	jdff dff_A_A9lO3CyH0_0(.dout(w_dff_A_tei56dez2_0),.din(w_dff_A_A9lO3CyH0_0),.clk(gclk));
	jdff dff_A_tei56dez2_0(.dout(w_dff_A_dbgaP0Rd6_0),.din(w_dff_A_tei56dez2_0),.clk(gclk));
	jdff dff_A_dbgaP0Rd6_0(.dout(w_dff_A_zIE918rM8_0),.din(w_dff_A_dbgaP0Rd6_0),.clk(gclk));
	jdff dff_A_zIE918rM8_0(.dout(w_dff_A_jHC6zbkX0_0),.din(w_dff_A_zIE918rM8_0),.clk(gclk));
	jdff dff_A_jHC6zbkX0_0(.dout(w_dff_A_yXCkIIaN8_0),.din(w_dff_A_jHC6zbkX0_0),.clk(gclk));
	jdff dff_A_yXCkIIaN8_0(.dout(w_dff_A_Kd84SJZL2_0),.din(w_dff_A_yXCkIIaN8_0),.clk(gclk));
	jdff dff_A_Kd84SJZL2_0(.dout(w_dff_A_XpduZ7gz3_0),.din(w_dff_A_Kd84SJZL2_0),.clk(gclk));
	jdff dff_A_XpduZ7gz3_0(.dout(w_dff_A_ZcQWVm3f9_0),.din(w_dff_A_XpduZ7gz3_0),.clk(gclk));
	jdff dff_A_ZcQWVm3f9_0(.dout(G848),.din(w_dff_A_ZcQWVm3f9_0),.clk(gclk));
	jdff dff_A_A8hVAlbl2_1(.dout(w_dff_A_KH2E4U4e4_0),.din(w_dff_A_A8hVAlbl2_1),.clk(gclk));
	jdff dff_A_KH2E4U4e4_0(.dout(w_dff_A_tkfU81ia3_0),.din(w_dff_A_KH2E4U4e4_0),.clk(gclk));
	jdff dff_A_tkfU81ia3_0(.dout(w_dff_A_nCnTvZXH7_0),.din(w_dff_A_tkfU81ia3_0),.clk(gclk));
	jdff dff_A_nCnTvZXH7_0(.dout(w_dff_A_92PqVcHB6_0),.din(w_dff_A_nCnTvZXH7_0),.clk(gclk));
	jdff dff_A_92PqVcHB6_0(.dout(w_dff_A_tNAYM1pR1_0),.din(w_dff_A_92PqVcHB6_0),.clk(gclk));
	jdff dff_A_tNAYM1pR1_0(.dout(w_dff_A_wVXn3hKW8_0),.din(w_dff_A_tNAYM1pR1_0),.clk(gclk));
	jdff dff_A_wVXn3hKW8_0(.dout(w_dff_A_rIPsPQuG7_0),.din(w_dff_A_wVXn3hKW8_0),.clk(gclk));
	jdff dff_A_rIPsPQuG7_0(.dout(w_dff_A_zgWqaAK52_0),.din(w_dff_A_rIPsPQuG7_0),.clk(gclk));
	jdff dff_A_zgWqaAK52_0(.dout(w_dff_A_dtvCJSli3_0),.din(w_dff_A_zgWqaAK52_0),.clk(gclk));
	jdff dff_A_dtvCJSli3_0(.dout(w_dff_A_yJayNhdq3_0),.din(w_dff_A_dtvCJSli3_0),.clk(gclk));
	jdff dff_A_yJayNhdq3_0(.dout(w_dff_A_2GEzOe1q2_0),.din(w_dff_A_yJayNhdq3_0),.clk(gclk));
	jdff dff_A_2GEzOe1q2_0(.dout(w_dff_A_L5oDVMKh8_0),.din(w_dff_A_2GEzOe1q2_0),.clk(gclk));
	jdff dff_A_L5oDVMKh8_0(.dout(w_dff_A_BowNEFNZ4_0),.din(w_dff_A_L5oDVMKh8_0),.clk(gclk));
	jdff dff_A_BowNEFNZ4_0(.dout(w_dff_A_VKRxySFe8_0),.din(w_dff_A_BowNEFNZ4_0),.clk(gclk));
	jdff dff_A_VKRxySFe8_0(.dout(w_dff_A_WLAFVOWO8_0),.din(w_dff_A_VKRxySFe8_0),.clk(gclk));
	jdff dff_A_WLAFVOWO8_0(.dout(w_dff_A_Bgsxl5rv3_0),.din(w_dff_A_WLAFVOWO8_0),.clk(gclk));
	jdff dff_A_Bgsxl5rv3_0(.dout(w_dff_A_QgrlKjMZ9_0),.din(w_dff_A_Bgsxl5rv3_0),.clk(gclk));
	jdff dff_A_QgrlKjMZ9_0(.dout(w_dff_A_9CvrZqXc7_0),.din(w_dff_A_QgrlKjMZ9_0),.clk(gclk));
	jdff dff_A_9CvrZqXc7_0(.dout(w_dff_A_cNkqUffv4_0),.din(w_dff_A_9CvrZqXc7_0),.clk(gclk));
	jdff dff_A_cNkqUffv4_0(.dout(w_dff_A_ajt3F2WD9_0),.din(w_dff_A_cNkqUffv4_0),.clk(gclk));
	jdff dff_A_ajt3F2WD9_0(.dout(w_dff_A_dqDyWFJM1_0),.din(w_dff_A_ajt3F2WD9_0),.clk(gclk));
	jdff dff_A_dqDyWFJM1_0(.dout(w_dff_A_UXRWSh954_0),.din(w_dff_A_dqDyWFJM1_0),.clk(gclk));
	jdff dff_A_UXRWSh954_0(.dout(w_dff_A_5VHLvVjS9_0),.din(w_dff_A_UXRWSh954_0),.clk(gclk));
	jdff dff_A_5VHLvVjS9_0(.dout(w_dff_A_yt3bbOY15_0),.din(w_dff_A_5VHLvVjS9_0),.clk(gclk));
	jdff dff_A_yt3bbOY15_0(.dout(G849),.din(w_dff_A_yt3bbOY15_0),.clk(gclk));
	jdff dff_A_6894XwHg4_1(.dout(w_dff_A_VUbwMfnm3_0),.din(w_dff_A_6894XwHg4_1),.clk(gclk));
	jdff dff_A_VUbwMfnm3_0(.dout(w_dff_A_zr9POrwW8_0),.din(w_dff_A_VUbwMfnm3_0),.clk(gclk));
	jdff dff_A_zr9POrwW8_0(.dout(w_dff_A_sMbWaRLX6_0),.din(w_dff_A_zr9POrwW8_0),.clk(gclk));
	jdff dff_A_sMbWaRLX6_0(.dout(w_dff_A_1XPA7sXR5_0),.din(w_dff_A_sMbWaRLX6_0),.clk(gclk));
	jdff dff_A_1XPA7sXR5_0(.dout(w_dff_A_kFXeJVb30_0),.din(w_dff_A_1XPA7sXR5_0),.clk(gclk));
	jdff dff_A_kFXeJVb30_0(.dout(w_dff_A_y2PETxVf7_0),.din(w_dff_A_kFXeJVb30_0),.clk(gclk));
	jdff dff_A_y2PETxVf7_0(.dout(w_dff_A_x4CznEat7_0),.din(w_dff_A_y2PETxVf7_0),.clk(gclk));
	jdff dff_A_x4CznEat7_0(.dout(w_dff_A_PRj8j7ey4_0),.din(w_dff_A_x4CznEat7_0),.clk(gclk));
	jdff dff_A_PRj8j7ey4_0(.dout(w_dff_A_FrficphV1_0),.din(w_dff_A_PRj8j7ey4_0),.clk(gclk));
	jdff dff_A_FrficphV1_0(.dout(w_dff_A_s5TIPeLb3_0),.din(w_dff_A_FrficphV1_0),.clk(gclk));
	jdff dff_A_s5TIPeLb3_0(.dout(w_dff_A_2kcw91Yq1_0),.din(w_dff_A_s5TIPeLb3_0),.clk(gclk));
	jdff dff_A_2kcw91Yq1_0(.dout(w_dff_A_8sfHadIK8_0),.din(w_dff_A_2kcw91Yq1_0),.clk(gclk));
	jdff dff_A_8sfHadIK8_0(.dout(w_dff_A_OSf0b74V5_0),.din(w_dff_A_8sfHadIK8_0),.clk(gclk));
	jdff dff_A_OSf0b74V5_0(.dout(w_dff_A_dRVYuHOA4_0),.din(w_dff_A_OSf0b74V5_0),.clk(gclk));
	jdff dff_A_dRVYuHOA4_0(.dout(w_dff_A_2M1msprE8_0),.din(w_dff_A_dRVYuHOA4_0),.clk(gclk));
	jdff dff_A_2M1msprE8_0(.dout(w_dff_A_gOzqewLt1_0),.din(w_dff_A_2M1msprE8_0),.clk(gclk));
	jdff dff_A_gOzqewLt1_0(.dout(w_dff_A_a5EILIGX6_0),.din(w_dff_A_gOzqewLt1_0),.clk(gclk));
	jdff dff_A_a5EILIGX6_0(.dout(w_dff_A_582nY0w96_0),.din(w_dff_A_a5EILIGX6_0),.clk(gclk));
	jdff dff_A_582nY0w96_0(.dout(w_dff_A_QMTVzXzd3_0),.din(w_dff_A_582nY0w96_0),.clk(gclk));
	jdff dff_A_QMTVzXzd3_0(.dout(w_dff_A_cIUchttw2_0),.din(w_dff_A_QMTVzXzd3_0),.clk(gclk));
	jdff dff_A_cIUchttw2_0(.dout(w_dff_A_C5aoSTNr3_0),.din(w_dff_A_cIUchttw2_0),.clk(gclk));
	jdff dff_A_C5aoSTNr3_0(.dout(w_dff_A_kIt2ysnS1_0),.din(w_dff_A_C5aoSTNr3_0),.clk(gclk));
	jdff dff_A_kIt2ysnS1_0(.dout(w_dff_A_5JgXSuOx1_0),.din(w_dff_A_kIt2ysnS1_0),.clk(gclk));
	jdff dff_A_5JgXSuOx1_0(.dout(w_dff_A_nKfqeR3a3_0),.din(w_dff_A_5JgXSuOx1_0),.clk(gclk));
	jdff dff_A_nKfqeR3a3_0(.dout(G850),.din(w_dff_A_nKfqeR3a3_0),.clk(gclk));
	jdff dff_A_HHWOph5b7_1(.dout(w_dff_A_ZAzv3gLz8_0),.din(w_dff_A_HHWOph5b7_1),.clk(gclk));
	jdff dff_A_ZAzv3gLz8_0(.dout(w_dff_A_Kels9HHA8_0),.din(w_dff_A_ZAzv3gLz8_0),.clk(gclk));
	jdff dff_A_Kels9HHA8_0(.dout(w_dff_A_LkcUbwPK6_0),.din(w_dff_A_Kels9HHA8_0),.clk(gclk));
	jdff dff_A_LkcUbwPK6_0(.dout(w_dff_A_B9sJDTNd5_0),.din(w_dff_A_LkcUbwPK6_0),.clk(gclk));
	jdff dff_A_B9sJDTNd5_0(.dout(w_dff_A_1DfwWTjw2_0),.din(w_dff_A_B9sJDTNd5_0),.clk(gclk));
	jdff dff_A_1DfwWTjw2_0(.dout(w_dff_A_C13xRN3G3_0),.din(w_dff_A_1DfwWTjw2_0),.clk(gclk));
	jdff dff_A_C13xRN3G3_0(.dout(w_dff_A_9h366wQY5_0),.din(w_dff_A_C13xRN3G3_0),.clk(gclk));
	jdff dff_A_9h366wQY5_0(.dout(w_dff_A_aHEwNMML6_0),.din(w_dff_A_9h366wQY5_0),.clk(gclk));
	jdff dff_A_aHEwNMML6_0(.dout(w_dff_A_rtXwMPxD3_0),.din(w_dff_A_aHEwNMML6_0),.clk(gclk));
	jdff dff_A_rtXwMPxD3_0(.dout(w_dff_A_0qSHGKcc8_0),.din(w_dff_A_rtXwMPxD3_0),.clk(gclk));
	jdff dff_A_0qSHGKcc8_0(.dout(w_dff_A_eDZD0ueg6_0),.din(w_dff_A_0qSHGKcc8_0),.clk(gclk));
	jdff dff_A_eDZD0ueg6_0(.dout(w_dff_A_48n1I4sP6_0),.din(w_dff_A_eDZD0ueg6_0),.clk(gclk));
	jdff dff_A_48n1I4sP6_0(.dout(w_dff_A_5VSxk5bT8_0),.din(w_dff_A_48n1I4sP6_0),.clk(gclk));
	jdff dff_A_5VSxk5bT8_0(.dout(w_dff_A_tlqG2zrB3_0),.din(w_dff_A_5VSxk5bT8_0),.clk(gclk));
	jdff dff_A_tlqG2zrB3_0(.dout(w_dff_A_hntE2EzT4_0),.din(w_dff_A_tlqG2zrB3_0),.clk(gclk));
	jdff dff_A_hntE2EzT4_0(.dout(w_dff_A_frLa6Gon1_0),.din(w_dff_A_hntE2EzT4_0),.clk(gclk));
	jdff dff_A_frLa6Gon1_0(.dout(w_dff_A_teqW8fCd1_0),.din(w_dff_A_frLa6Gon1_0),.clk(gclk));
	jdff dff_A_teqW8fCd1_0(.dout(w_dff_A_DrdRFazP4_0),.din(w_dff_A_teqW8fCd1_0),.clk(gclk));
	jdff dff_A_DrdRFazP4_0(.dout(w_dff_A_Wn06qBZI2_0),.din(w_dff_A_DrdRFazP4_0),.clk(gclk));
	jdff dff_A_Wn06qBZI2_0(.dout(w_dff_A_QnuJmDG62_0),.din(w_dff_A_Wn06qBZI2_0),.clk(gclk));
	jdff dff_A_QnuJmDG62_0(.dout(w_dff_A_6aFDZH2V1_0),.din(w_dff_A_QnuJmDG62_0),.clk(gclk));
	jdff dff_A_6aFDZH2V1_0(.dout(w_dff_A_MivsMC8G0_0),.din(w_dff_A_6aFDZH2V1_0),.clk(gclk));
	jdff dff_A_MivsMC8G0_0(.dout(w_dff_A_G6V5Phx14_0),.din(w_dff_A_MivsMC8G0_0),.clk(gclk));
	jdff dff_A_G6V5Phx14_0(.dout(w_dff_A_BBo1gajo5_0),.din(w_dff_A_G6V5Phx14_0),.clk(gclk));
	jdff dff_A_BBo1gajo5_0(.dout(G851),.din(w_dff_A_BBo1gajo5_0),.clk(gclk));
	jdff dff_A_YkzxoQtB2_2(.dout(w_dff_A_mmoyTtaK6_0),.din(w_dff_A_YkzxoQtB2_2),.clk(gclk));
	jdff dff_A_mmoyTtaK6_0(.dout(w_dff_A_UYGS9ZSh3_0),.din(w_dff_A_mmoyTtaK6_0),.clk(gclk));
	jdff dff_A_UYGS9ZSh3_0(.dout(w_dff_A_QmOblBJQ6_0),.din(w_dff_A_UYGS9ZSh3_0),.clk(gclk));
	jdff dff_A_QmOblBJQ6_0(.dout(w_dff_A_eP4zlPHi9_0),.din(w_dff_A_QmOblBJQ6_0),.clk(gclk));
	jdff dff_A_eP4zlPHi9_0(.dout(w_dff_A_odDFbvq47_0),.din(w_dff_A_eP4zlPHi9_0),.clk(gclk));
	jdff dff_A_odDFbvq47_0(.dout(w_dff_A_GykK2TQp8_0),.din(w_dff_A_odDFbvq47_0),.clk(gclk));
	jdff dff_A_GykK2TQp8_0(.dout(w_dff_A_kegSiuQZ0_0),.din(w_dff_A_GykK2TQp8_0),.clk(gclk));
	jdff dff_A_kegSiuQZ0_0(.dout(w_dff_A_LsPpmI8K4_0),.din(w_dff_A_kegSiuQZ0_0),.clk(gclk));
	jdff dff_A_LsPpmI8K4_0(.dout(w_dff_A_P7vfS4vW8_0),.din(w_dff_A_LsPpmI8K4_0),.clk(gclk));
	jdff dff_A_P7vfS4vW8_0(.dout(w_dff_A_wYl99yhY5_0),.din(w_dff_A_P7vfS4vW8_0),.clk(gclk));
	jdff dff_A_wYl99yhY5_0(.dout(w_dff_A_mdSwKMO74_0),.din(w_dff_A_wYl99yhY5_0),.clk(gclk));
	jdff dff_A_mdSwKMO74_0(.dout(w_dff_A_uZ27h9L10_0),.din(w_dff_A_mdSwKMO74_0),.clk(gclk));
	jdff dff_A_uZ27h9L10_0(.dout(w_dff_A_7dZeTwjs7_0),.din(w_dff_A_uZ27h9L10_0),.clk(gclk));
	jdff dff_A_7dZeTwjs7_0(.dout(w_dff_A_xdFoL6JW4_0),.din(w_dff_A_7dZeTwjs7_0),.clk(gclk));
	jdff dff_A_xdFoL6JW4_0(.dout(w_dff_A_J9zpjoO99_0),.din(w_dff_A_xdFoL6JW4_0),.clk(gclk));
	jdff dff_A_J9zpjoO99_0(.dout(w_dff_A_SpWTup9B5_0),.din(w_dff_A_J9zpjoO99_0),.clk(gclk));
	jdff dff_A_SpWTup9B5_0(.dout(w_dff_A_Iizw5isy6_0),.din(w_dff_A_SpWTup9B5_0),.clk(gclk));
	jdff dff_A_Iizw5isy6_0(.dout(w_dff_A_WW3mjIsK2_0),.din(w_dff_A_Iizw5isy6_0),.clk(gclk));
	jdff dff_A_WW3mjIsK2_0(.dout(w_dff_A_Qax9Srjc9_0),.din(w_dff_A_WW3mjIsK2_0),.clk(gclk));
	jdff dff_A_Qax9Srjc9_0(.dout(w_dff_A_bVqY3Jc39_0),.din(w_dff_A_Qax9Srjc9_0),.clk(gclk));
	jdff dff_A_bVqY3Jc39_0(.dout(w_dff_A_hdUwCm208_0),.din(w_dff_A_bVqY3Jc39_0),.clk(gclk));
	jdff dff_A_hdUwCm208_0(.dout(w_dff_A_Uo588KnT3_0),.din(w_dff_A_hdUwCm208_0),.clk(gclk));
	jdff dff_A_Uo588KnT3_0(.dout(w_dff_A_sMAmJ0391_0),.din(w_dff_A_Uo588KnT3_0),.clk(gclk));
	jdff dff_A_sMAmJ0391_0(.dout(w_dff_A_SYGTJskO0_0),.din(w_dff_A_sMAmJ0391_0),.clk(gclk));
	jdff dff_A_SYGTJskO0_0(.dout(G634),.din(w_dff_A_SYGTJskO0_0),.clk(gclk));
	jdff dff_A_gMoTHiyF2_2(.dout(w_dff_A_VTjsgKuU1_0),.din(w_dff_A_gMoTHiyF2_2),.clk(gclk));
	jdff dff_A_VTjsgKuU1_0(.dout(w_dff_A_b2ZEFNbE4_0),.din(w_dff_A_VTjsgKuU1_0),.clk(gclk));
	jdff dff_A_b2ZEFNbE4_0(.dout(w_dff_A_apAu1UK38_0),.din(w_dff_A_b2ZEFNbE4_0),.clk(gclk));
	jdff dff_A_apAu1UK38_0(.dout(w_dff_A_1xrwjf0X2_0),.din(w_dff_A_apAu1UK38_0),.clk(gclk));
	jdff dff_A_1xrwjf0X2_0(.dout(w_dff_A_D61E1PyV9_0),.din(w_dff_A_1xrwjf0X2_0),.clk(gclk));
	jdff dff_A_D61E1PyV9_0(.dout(w_dff_A_7QbUsl7H7_0),.din(w_dff_A_D61E1PyV9_0),.clk(gclk));
	jdff dff_A_7QbUsl7H7_0(.dout(w_dff_A_mdLjyh2k4_0),.din(w_dff_A_7QbUsl7H7_0),.clk(gclk));
	jdff dff_A_mdLjyh2k4_0(.dout(w_dff_A_VROJQ4Gx0_0),.din(w_dff_A_mdLjyh2k4_0),.clk(gclk));
	jdff dff_A_VROJQ4Gx0_0(.dout(w_dff_A_1sAMcDo47_0),.din(w_dff_A_VROJQ4Gx0_0),.clk(gclk));
	jdff dff_A_1sAMcDo47_0(.dout(w_dff_A_CijIXDxo4_0),.din(w_dff_A_1sAMcDo47_0),.clk(gclk));
	jdff dff_A_CijIXDxo4_0(.dout(w_dff_A_St6DHmPu7_0),.din(w_dff_A_CijIXDxo4_0),.clk(gclk));
	jdff dff_A_St6DHmPu7_0(.dout(w_dff_A_snPcbtFQ5_0),.din(w_dff_A_St6DHmPu7_0),.clk(gclk));
	jdff dff_A_snPcbtFQ5_0(.dout(w_dff_A_qyj4bKDl1_0),.din(w_dff_A_snPcbtFQ5_0),.clk(gclk));
	jdff dff_A_qyj4bKDl1_0(.dout(w_dff_A_FZlwYflm1_0),.din(w_dff_A_qyj4bKDl1_0),.clk(gclk));
	jdff dff_A_FZlwYflm1_0(.dout(w_dff_A_IcH8j55H2_0),.din(w_dff_A_FZlwYflm1_0),.clk(gclk));
	jdff dff_A_IcH8j55H2_0(.dout(w_dff_A_dGM0tJA56_0),.din(w_dff_A_IcH8j55H2_0),.clk(gclk));
	jdff dff_A_dGM0tJA56_0(.dout(w_dff_A_6CXnUImU7_0),.din(w_dff_A_dGM0tJA56_0),.clk(gclk));
	jdff dff_A_6CXnUImU7_0(.dout(w_dff_A_SHy3muHk4_0),.din(w_dff_A_6CXnUImU7_0),.clk(gclk));
	jdff dff_A_SHy3muHk4_0(.dout(w_dff_A_hwHC8ITx6_0),.din(w_dff_A_SHy3muHk4_0),.clk(gclk));
	jdff dff_A_hwHC8ITx6_0(.dout(w_dff_A_zmw4w8hz5_0),.din(w_dff_A_hwHC8ITx6_0),.clk(gclk));
	jdff dff_A_zmw4w8hz5_0(.dout(w_dff_A_sYxNjcml1_0),.din(w_dff_A_zmw4w8hz5_0),.clk(gclk));
	jdff dff_A_sYxNjcml1_0(.dout(w_dff_A_l5LsU9RF8_0),.din(w_dff_A_sYxNjcml1_0),.clk(gclk));
	jdff dff_A_l5LsU9RF8_0(.dout(w_dff_A_t8HbDwEf1_0),.din(w_dff_A_l5LsU9RF8_0),.clk(gclk));
	jdff dff_A_t8HbDwEf1_0(.dout(G815),.din(w_dff_A_t8HbDwEf1_0),.clk(gclk));
	jdff dff_A_YXrgNVZe8_2(.dout(w_dff_A_XBiahQiV1_0),.din(w_dff_A_YXrgNVZe8_2),.clk(gclk));
	jdff dff_A_XBiahQiV1_0(.dout(w_dff_A_VHUl1q965_0),.din(w_dff_A_XBiahQiV1_0),.clk(gclk));
	jdff dff_A_VHUl1q965_0(.dout(w_dff_A_5kJR66x03_0),.din(w_dff_A_VHUl1q965_0),.clk(gclk));
	jdff dff_A_5kJR66x03_0(.dout(w_dff_A_k8G3Iiji4_0),.din(w_dff_A_5kJR66x03_0),.clk(gclk));
	jdff dff_A_k8G3Iiji4_0(.dout(w_dff_A_SBLV8qSQ0_0),.din(w_dff_A_k8G3Iiji4_0),.clk(gclk));
	jdff dff_A_SBLV8qSQ0_0(.dout(w_dff_A_eu8hscUt3_0),.din(w_dff_A_SBLV8qSQ0_0),.clk(gclk));
	jdff dff_A_eu8hscUt3_0(.dout(w_dff_A_pD89C3Zv5_0),.din(w_dff_A_eu8hscUt3_0),.clk(gclk));
	jdff dff_A_pD89C3Zv5_0(.dout(w_dff_A_VlRmVwy42_0),.din(w_dff_A_pD89C3Zv5_0),.clk(gclk));
	jdff dff_A_VlRmVwy42_0(.dout(w_dff_A_YONZH3dx4_0),.din(w_dff_A_VlRmVwy42_0),.clk(gclk));
	jdff dff_A_YONZH3dx4_0(.dout(w_dff_A_DPkgoYry5_0),.din(w_dff_A_YONZH3dx4_0),.clk(gclk));
	jdff dff_A_DPkgoYry5_0(.dout(w_dff_A_dzQlXcd66_0),.din(w_dff_A_DPkgoYry5_0),.clk(gclk));
	jdff dff_A_dzQlXcd66_0(.dout(w_dff_A_Y0zh1ZFY3_0),.din(w_dff_A_dzQlXcd66_0),.clk(gclk));
	jdff dff_A_Y0zh1ZFY3_0(.dout(w_dff_A_MqYoul0z3_0),.din(w_dff_A_Y0zh1ZFY3_0),.clk(gclk));
	jdff dff_A_MqYoul0z3_0(.dout(w_dff_A_ClAPdzkd6_0),.din(w_dff_A_MqYoul0z3_0),.clk(gclk));
	jdff dff_A_ClAPdzkd6_0(.dout(w_dff_A_dtA90Sy32_0),.din(w_dff_A_ClAPdzkd6_0),.clk(gclk));
	jdff dff_A_dtA90Sy32_0(.dout(w_dff_A_VjPpPFTp6_0),.din(w_dff_A_dtA90Sy32_0),.clk(gclk));
	jdff dff_A_VjPpPFTp6_0(.dout(w_dff_A_ApezIZL96_0),.din(w_dff_A_VjPpPFTp6_0),.clk(gclk));
	jdff dff_A_ApezIZL96_0(.dout(w_dff_A_QSzkMrGA6_0),.din(w_dff_A_ApezIZL96_0),.clk(gclk));
	jdff dff_A_QSzkMrGA6_0(.dout(w_dff_A_tx9EFmX79_0),.din(w_dff_A_QSzkMrGA6_0),.clk(gclk));
	jdff dff_A_tx9EFmX79_0(.dout(w_dff_A_4onzlFIs1_0),.din(w_dff_A_tx9EFmX79_0),.clk(gclk));
	jdff dff_A_4onzlFIs1_0(.dout(w_dff_A_A8BHtBpx3_0),.din(w_dff_A_4onzlFIs1_0),.clk(gclk));
	jdff dff_A_A8BHtBpx3_0(.dout(w_dff_A_pSIcjSir7_0),.din(w_dff_A_A8BHtBpx3_0),.clk(gclk));
	jdff dff_A_pSIcjSir7_0(.dout(w_dff_A_ufMWgX2S9_0),.din(w_dff_A_pSIcjSir7_0),.clk(gclk));
	jdff dff_A_ufMWgX2S9_0(.dout(G845),.din(w_dff_A_ufMWgX2S9_0),.clk(gclk));
	jdff dff_A_1vhZ3Duu7_1(.dout(w_dff_A_xaBEhCvg3_0),.din(w_dff_A_1vhZ3Duu7_1),.clk(gclk));
	jdff dff_A_xaBEhCvg3_0(.dout(w_dff_A_pMzJ0rrY7_0),.din(w_dff_A_xaBEhCvg3_0),.clk(gclk));
	jdff dff_A_pMzJ0rrY7_0(.dout(w_dff_A_fO54PrRc4_0),.din(w_dff_A_pMzJ0rrY7_0),.clk(gclk));
	jdff dff_A_fO54PrRc4_0(.dout(w_dff_A_eWGuX4Hb2_0),.din(w_dff_A_fO54PrRc4_0),.clk(gclk));
	jdff dff_A_eWGuX4Hb2_0(.dout(w_dff_A_NR5x9ZaJ0_0),.din(w_dff_A_eWGuX4Hb2_0),.clk(gclk));
	jdff dff_A_NR5x9ZaJ0_0(.dout(w_dff_A_MWxkboMK8_0),.din(w_dff_A_NR5x9ZaJ0_0),.clk(gclk));
	jdff dff_A_MWxkboMK8_0(.dout(w_dff_A_UKXlgs5R2_0),.din(w_dff_A_MWxkboMK8_0),.clk(gclk));
	jdff dff_A_UKXlgs5R2_0(.dout(w_dff_A_uK8usMXv9_0),.din(w_dff_A_UKXlgs5R2_0),.clk(gclk));
	jdff dff_A_uK8usMXv9_0(.dout(w_dff_A_7dLbHxSa0_0),.din(w_dff_A_uK8usMXv9_0),.clk(gclk));
	jdff dff_A_7dLbHxSa0_0(.dout(w_dff_A_4aFYLfiw4_0),.din(w_dff_A_7dLbHxSa0_0),.clk(gclk));
	jdff dff_A_4aFYLfiw4_0(.dout(w_dff_A_OKojFEkQ4_0),.din(w_dff_A_4aFYLfiw4_0),.clk(gclk));
	jdff dff_A_OKojFEkQ4_0(.dout(w_dff_A_fbpJGHyl3_0),.din(w_dff_A_OKojFEkQ4_0),.clk(gclk));
	jdff dff_A_fbpJGHyl3_0(.dout(w_dff_A_FhDDhKGI1_0),.din(w_dff_A_fbpJGHyl3_0),.clk(gclk));
	jdff dff_A_FhDDhKGI1_0(.dout(w_dff_A_LHAumLIi6_0),.din(w_dff_A_FhDDhKGI1_0),.clk(gclk));
	jdff dff_A_LHAumLIi6_0(.dout(w_dff_A_HsLX4xME8_0),.din(w_dff_A_LHAumLIi6_0),.clk(gclk));
	jdff dff_A_HsLX4xME8_0(.dout(w_dff_A_CfemMX3W6_0),.din(w_dff_A_HsLX4xME8_0),.clk(gclk));
	jdff dff_A_CfemMX3W6_0(.dout(w_dff_A_i1NQu6Jo8_0),.din(w_dff_A_CfemMX3W6_0),.clk(gclk));
	jdff dff_A_i1NQu6Jo8_0(.dout(w_dff_A_x9aHuxnc3_0),.din(w_dff_A_i1NQu6Jo8_0),.clk(gclk));
	jdff dff_A_x9aHuxnc3_0(.dout(w_dff_A_RZLM3YlS2_0),.din(w_dff_A_x9aHuxnc3_0),.clk(gclk));
	jdff dff_A_RZLM3YlS2_0(.dout(w_dff_A_rRg7ndCF2_0),.din(w_dff_A_RZLM3YlS2_0),.clk(gclk));
	jdff dff_A_rRg7ndCF2_0(.dout(w_dff_A_2h9pkyBl4_0),.din(w_dff_A_rRg7ndCF2_0),.clk(gclk));
	jdff dff_A_2h9pkyBl4_0(.dout(w_dff_A_HCWGWcV32_0),.din(w_dff_A_2h9pkyBl4_0),.clk(gclk));
	jdff dff_A_HCWGWcV32_0(.dout(w_dff_A_blhjv9jP2_0),.din(w_dff_A_HCWGWcV32_0),.clk(gclk));
	jdff dff_A_blhjv9jP2_0(.dout(G847),.din(w_dff_A_blhjv9jP2_0),.clk(gclk));
	jdff dff_A_2BQXXCY79_1(.dout(w_dff_A_xRGig8377_0),.din(w_dff_A_2BQXXCY79_1),.clk(gclk));
	jdff dff_A_xRGig8377_0(.dout(w_dff_A_RIhUx2nw8_0),.din(w_dff_A_xRGig8377_0),.clk(gclk));
	jdff dff_A_RIhUx2nw8_0(.dout(w_dff_A_aJAoDH2g5_0),.din(w_dff_A_RIhUx2nw8_0),.clk(gclk));
	jdff dff_A_aJAoDH2g5_0(.dout(w_dff_A_xyljvqlp7_0),.din(w_dff_A_aJAoDH2g5_0),.clk(gclk));
	jdff dff_A_xyljvqlp7_0(.dout(w_dff_A_kYNBknzr6_0),.din(w_dff_A_xyljvqlp7_0),.clk(gclk));
	jdff dff_A_kYNBknzr6_0(.dout(w_dff_A_e4dVA2Wt2_0),.din(w_dff_A_kYNBknzr6_0),.clk(gclk));
	jdff dff_A_e4dVA2Wt2_0(.dout(w_dff_A_LAGxNsX03_0),.din(w_dff_A_e4dVA2Wt2_0),.clk(gclk));
	jdff dff_A_LAGxNsX03_0(.dout(w_dff_A_kgcAoagA8_0),.din(w_dff_A_LAGxNsX03_0),.clk(gclk));
	jdff dff_A_kgcAoagA8_0(.dout(w_dff_A_PBlo9OsH1_0),.din(w_dff_A_kgcAoagA8_0),.clk(gclk));
	jdff dff_A_PBlo9OsH1_0(.dout(w_dff_A_JM4zImIa8_0),.din(w_dff_A_PBlo9OsH1_0),.clk(gclk));
	jdff dff_A_JM4zImIa8_0(.dout(w_dff_A_iP1J6CzE5_0),.din(w_dff_A_JM4zImIa8_0),.clk(gclk));
	jdff dff_A_iP1J6CzE5_0(.dout(w_dff_A_MhWhCN8g5_0),.din(w_dff_A_iP1J6CzE5_0),.clk(gclk));
	jdff dff_A_MhWhCN8g5_0(.dout(w_dff_A_TEZCAOzt6_0),.din(w_dff_A_MhWhCN8g5_0),.clk(gclk));
	jdff dff_A_TEZCAOzt6_0(.dout(w_dff_A_ujoQjHiV7_0),.din(w_dff_A_TEZCAOzt6_0),.clk(gclk));
	jdff dff_A_ujoQjHiV7_0(.dout(w_dff_A_rN5FmHAw0_0),.din(w_dff_A_ujoQjHiV7_0),.clk(gclk));
	jdff dff_A_rN5FmHAw0_0(.dout(w_dff_A_aF6gTfrh1_0),.din(w_dff_A_rN5FmHAw0_0),.clk(gclk));
	jdff dff_A_aF6gTfrh1_0(.dout(w_dff_A_7gd1M7G10_0),.din(w_dff_A_aF6gTfrh1_0),.clk(gclk));
	jdff dff_A_7gd1M7G10_0(.dout(w_dff_A_jWpSByPW4_0),.din(w_dff_A_7gd1M7G10_0),.clk(gclk));
	jdff dff_A_jWpSByPW4_0(.dout(w_dff_A_0Xqw2c5Z1_0),.din(w_dff_A_jWpSByPW4_0),.clk(gclk));
	jdff dff_A_0Xqw2c5Z1_0(.dout(w_dff_A_zoN5m0oc5_0),.din(w_dff_A_0Xqw2c5Z1_0),.clk(gclk));
	jdff dff_A_zoN5m0oc5_0(.dout(w_dff_A_2Gpg6zHf6_0),.din(w_dff_A_zoN5m0oc5_0),.clk(gclk));
	jdff dff_A_2Gpg6zHf6_0(.dout(w_dff_A_xEoyoL3u4_0),.din(w_dff_A_2Gpg6zHf6_0),.clk(gclk));
	jdff dff_A_xEoyoL3u4_0(.dout(w_dff_A_4EYDmp5c0_0),.din(w_dff_A_xEoyoL3u4_0),.clk(gclk));
	jdff dff_A_4EYDmp5c0_0(.dout(w_dff_A_6BNVEGbH7_0),.din(w_dff_A_4EYDmp5c0_0),.clk(gclk));
	jdff dff_A_6BNVEGbH7_0(.dout(w_dff_A_XHnryFNT6_0),.din(w_dff_A_6BNVEGbH7_0),.clk(gclk));
	jdff dff_A_XHnryFNT6_0(.dout(G926),.din(w_dff_A_XHnryFNT6_0),.clk(gclk));
	jdff dff_A_RJ7IrVGd3_1(.dout(w_dff_A_EQ37yykE3_0),.din(w_dff_A_RJ7IrVGd3_1),.clk(gclk));
	jdff dff_A_EQ37yykE3_0(.dout(w_dff_A_VLt9xiM65_0),.din(w_dff_A_EQ37yykE3_0),.clk(gclk));
	jdff dff_A_VLt9xiM65_0(.dout(w_dff_A_DSCdIuQx6_0),.din(w_dff_A_VLt9xiM65_0),.clk(gclk));
	jdff dff_A_DSCdIuQx6_0(.dout(w_dff_A_iApKW7MT5_0),.din(w_dff_A_DSCdIuQx6_0),.clk(gclk));
	jdff dff_A_iApKW7MT5_0(.dout(w_dff_A_CUKLLEQw9_0),.din(w_dff_A_iApKW7MT5_0),.clk(gclk));
	jdff dff_A_CUKLLEQw9_0(.dout(w_dff_A_o0AZu8551_0),.din(w_dff_A_CUKLLEQw9_0),.clk(gclk));
	jdff dff_A_o0AZu8551_0(.dout(w_dff_A_qR4tpdR63_0),.din(w_dff_A_o0AZu8551_0),.clk(gclk));
	jdff dff_A_qR4tpdR63_0(.dout(w_dff_A_Y78l4tbm7_0),.din(w_dff_A_qR4tpdR63_0),.clk(gclk));
	jdff dff_A_Y78l4tbm7_0(.dout(w_dff_A_t0iMmbE84_0),.din(w_dff_A_Y78l4tbm7_0),.clk(gclk));
	jdff dff_A_t0iMmbE84_0(.dout(w_dff_A_aprY7Hxz7_0),.din(w_dff_A_t0iMmbE84_0),.clk(gclk));
	jdff dff_A_aprY7Hxz7_0(.dout(w_dff_A_T6rcURAQ7_0),.din(w_dff_A_aprY7Hxz7_0),.clk(gclk));
	jdff dff_A_T6rcURAQ7_0(.dout(w_dff_A_cSNB2yKf2_0),.din(w_dff_A_T6rcURAQ7_0),.clk(gclk));
	jdff dff_A_cSNB2yKf2_0(.dout(w_dff_A_IgglOpA07_0),.din(w_dff_A_cSNB2yKf2_0),.clk(gclk));
	jdff dff_A_IgglOpA07_0(.dout(w_dff_A_9kxFLE7j3_0),.din(w_dff_A_IgglOpA07_0),.clk(gclk));
	jdff dff_A_9kxFLE7j3_0(.dout(w_dff_A_l8NvcR8K1_0),.din(w_dff_A_9kxFLE7j3_0),.clk(gclk));
	jdff dff_A_l8NvcR8K1_0(.dout(w_dff_A_CSYG8x4H4_0),.din(w_dff_A_l8NvcR8K1_0),.clk(gclk));
	jdff dff_A_CSYG8x4H4_0(.dout(w_dff_A_pHJ7DrXq5_0),.din(w_dff_A_CSYG8x4H4_0),.clk(gclk));
	jdff dff_A_pHJ7DrXq5_0(.dout(w_dff_A_rpGTnU5z4_0),.din(w_dff_A_pHJ7DrXq5_0),.clk(gclk));
	jdff dff_A_rpGTnU5z4_0(.dout(w_dff_A_2Hrmf9zX9_0),.din(w_dff_A_rpGTnU5z4_0),.clk(gclk));
	jdff dff_A_2Hrmf9zX9_0(.dout(w_dff_A_0yDnFnFU8_0),.din(w_dff_A_2Hrmf9zX9_0),.clk(gclk));
	jdff dff_A_0yDnFnFU8_0(.dout(w_dff_A_ORSg5U0o0_0),.din(w_dff_A_0yDnFnFU8_0),.clk(gclk));
	jdff dff_A_ORSg5U0o0_0(.dout(w_dff_A_hxUxrhRC9_0),.din(w_dff_A_ORSg5U0o0_0),.clk(gclk));
	jdff dff_A_hxUxrhRC9_0(.dout(w_dff_A_Fl09Z4x47_0),.din(w_dff_A_hxUxrhRC9_0),.clk(gclk));
	jdff dff_A_Fl09Z4x47_0(.dout(w_dff_A_ReZpeQio9_0),.din(w_dff_A_Fl09Z4x47_0),.clk(gclk));
	jdff dff_A_ReZpeQio9_0(.dout(w_dff_A_hwsWkcta6_0),.din(w_dff_A_ReZpeQio9_0),.clk(gclk));
	jdff dff_A_hwsWkcta6_0(.dout(G923),.din(w_dff_A_hwsWkcta6_0),.clk(gclk));
	jdff dff_A_88VaWVqO6_1(.dout(w_dff_A_KafEuoPR1_0),.din(w_dff_A_88VaWVqO6_1),.clk(gclk));
	jdff dff_A_KafEuoPR1_0(.dout(w_dff_A_y8BZduW51_0),.din(w_dff_A_KafEuoPR1_0),.clk(gclk));
	jdff dff_A_y8BZduW51_0(.dout(w_dff_A_0otdT7wu5_0),.din(w_dff_A_y8BZduW51_0),.clk(gclk));
	jdff dff_A_0otdT7wu5_0(.dout(w_dff_A_wi4BtpDo2_0),.din(w_dff_A_0otdT7wu5_0),.clk(gclk));
	jdff dff_A_wi4BtpDo2_0(.dout(w_dff_A_EOmIOPxI8_0),.din(w_dff_A_wi4BtpDo2_0),.clk(gclk));
	jdff dff_A_EOmIOPxI8_0(.dout(w_dff_A_rJwRTXNY3_0),.din(w_dff_A_EOmIOPxI8_0),.clk(gclk));
	jdff dff_A_rJwRTXNY3_0(.dout(w_dff_A_2pBZzS9a0_0),.din(w_dff_A_rJwRTXNY3_0),.clk(gclk));
	jdff dff_A_2pBZzS9a0_0(.dout(w_dff_A_OZjfciZ72_0),.din(w_dff_A_2pBZzS9a0_0),.clk(gclk));
	jdff dff_A_OZjfciZ72_0(.dout(w_dff_A_SlnPlGr07_0),.din(w_dff_A_OZjfciZ72_0),.clk(gclk));
	jdff dff_A_SlnPlGr07_0(.dout(w_dff_A_k3fXH3ul1_0),.din(w_dff_A_SlnPlGr07_0),.clk(gclk));
	jdff dff_A_k3fXH3ul1_0(.dout(w_dff_A_RiZrk0bw3_0),.din(w_dff_A_k3fXH3ul1_0),.clk(gclk));
	jdff dff_A_RiZrk0bw3_0(.dout(w_dff_A_DNyaSlRn9_0),.din(w_dff_A_RiZrk0bw3_0),.clk(gclk));
	jdff dff_A_DNyaSlRn9_0(.dout(w_dff_A_4Gw6z5kt8_0),.din(w_dff_A_DNyaSlRn9_0),.clk(gclk));
	jdff dff_A_4Gw6z5kt8_0(.dout(w_dff_A_X9B1OuZc4_0),.din(w_dff_A_4Gw6z5kt8_0),.clk(gclk));
	jdff dff_A_X9B1OuZc4_0(.dout(w_dff_A_2VIMb5Cm1_0),.din(w_dff_A_X9B1OuZc4_0),.clk(gclk));
	jdff dff_A_2VIMb5Cm1_0(.dout(w_dff_A_cYzohbvw3_0),.din(w_dff_A_2VIMb5Cm1_0),.clk(gclk));
	jdff dff_A_cYzohbvw3_0(.dout(w_dff_A_FsVl5IM42_0),.din(w_dff_A_cYzohbvw3_0),.clk(gclk));
	jdff dff_A_FsVl5IM42_0(.dout(w_dff_A_INu8qnWm9_0),.din(w_dff_A_FsVl5IM42_0),.clk(gclk));
	jdff dff_A_INu8qnWm9_0(.dout(w_dff_A_8mtilUTZ5_0),.din(w_dff_A_INu8qnWm9_0),.clk(gclk));
	jdff dff_A_8mtilUTZ5_0(.dout(w_dff_A_PqAGtkmO5_0),.din(w_dff_A_8mtilUTZ5_0),.clk(gclk));
	jdff dff_A_PqAGtkmO5_0(.dout(w_dff_A_anoYIH2a4_0),.din(w_dff_A_PqAGtkmO5_0),.clk(gclk));
	jdff dff_A_anoYIH2a4_0(.dout(w_dff_A_mrfNQf350_0),.din(w_dff_A_anoYIH2a4_0),.clk(gclk));
	jdff dff_A_mrfNQf350_0(.dout(w_dff_A_JQf7NqGh5_0),.din(w_dff_A_mrfNQf350_0),.clk(gclk));
	jdff dff_A_JQf7NqGh5_0(.dout(w_dff_A_FjF4b82V7_0),.din(w_dff_A_JQf7NqGh5_0),.clk(gclk));
	jdff dff_A_FjF4b82V7_0(.dout(w_dff_A_jwap2BjM8_0),.din(w_dff_A_FjF4b82V7_0),.clk(gclk));
	jdff dff_A_jwap2BjM8_0(.dout(G921),.din(w_dff_A_jwap2BjM8_0),.clk(gclk));
	jdff dff_A_QSbbVJ567_1(.dout(w_dff_A_QaZHnHBu1_0),.din(w_dff_A_QSbbVJ567_1),.clk(gclk));
	jdff dff_A_QaZHnHBu1_0(.dout(w_dff_A_b0Q9CeWZ6_0),.din(w_dff_A_QaZHnHBu1_0),.clk(gclk));
	jdff dff_A_b0Q9CeWZ6_0(.dout(w_dff_A_q8qnf7pK3_0),.din(w_dff_A_b0Q9CeWZ6_0),.clk(gclk));
	jdff dff_A_q8qnf7pK3_0(.dout(w_dff_A_JlJcvdNA9_0),.din(w_dff_A_q8qnf7pK3_0),.clk(gclk));
	jdff dff_A_JlJcvdNA9_0(.dout(w_dff_A_TWurAjsC4_0),.din(w_dff_A_JlJcvdNA9_0),.clk(gclk));
	jdff dff_A_TWurAjsC4_0(.dout(w_dff_A_Cc5q8fmD4_0),.din(w_dff_A_TWurAjsC4_0),.clk(gclk));
	jdff dff_A_Cc5q8fmD4_0(.dout(w_dff_A_a3SwUa8v9_0),.din(w_dff_A_Cc5q8fmD4_0),.clk(gclk));
	jdff dff_A_a3SwUa8v9_0(.dout(w_dff_A_T8pQasFM0_0),.din(w_dff_A_a3SwUa8v9_0),.clk(gclk));
	jdff dff_A_T8pQasFM0_0(.dout(w_dff_A_cenyqIl21_0),.din(w_dff_A_T8pQasFM0_0),.clk(gclk));
	jdff dff_A_cenyqIl21_0(.dout(w_dff_A_MmF2BjKi5_0),.din(w_dff_A_cenyqIl21_0),.clk(gclk));
	jdff dff_A_MmF2BjKi5_0(.dout(w_dff_A_aCTppGsN4_0),.din(w_dff_A_MmF2BjKi5_0),.clk(gclk));
	jdff dff_A_aCTppGsN4_0(.dout(w_dff_A_fEsJgHJk9_0),.din(w_dff_A_aCTppGsN4_0),.clk(gclk));
	jdff dff_A_fEsJgHJk9_0(.dout(w_dff_A_TW6FMMtF0_0),.din(w_dff_A_fEsJgHJk9_0),.clk(gclk));
	jdff dff_A_TW6FMMtF0_0(.dout(w_dff_A_L5WsDwWb4_0),.din(w_dff_A_TW6FMMtF0_0),.clk(gclk));
	jdff dff_A_L5WsDwWb4_0(.dout(w_dff_A_kIj1TW136_0),.din(w_dff_A_L5WsDwWb4_0),.clk(gclk));
	jdff dff_A_kIj1TW136_0(.dout(w_dff_A_Es77KwOD5_0),.din(w_dff_A_kIj1TW136_0),.clk(gclk));
	jdff dff_A_Es77KwOD5_0(.dout(w_dff_A_ZvSmXE3U3_0),.din(w_dff_A_Es77KwOD5_0),.clk(gclk));
	jdff dff_A_ZvSmXE3U3_0(.dout(w_dff_A_YhyW6Jog0_0),.din(w_dff_A_ZvSmXE3U3_0),.clk(gclk));
	jdff dff_A_YhyW6Jog0_0(.dout(w_dff_A_j5E0o9H89_0),.din(w_dff_A_YhyW6Jog0_0),.clk(gclk));
	jdff dff_A_j5E0o9H89_0(.dout(w_dff_A_cXT5Wqs20_0),.din(w_dff_A_j5E0o9H89_0),.clk(gclk));
	jdff dff_A_cXT5Wqs20_0(.dout(w_dff_A_0VjhFhUN5_0),.din(w_dff_A_cXT5Wqs20_0),.clk(gclk));
	jdff dff_A_0VjhFhUN5_0(.dout(w_dff_A_qjYREwnY3_0),.din(w_dff_A_0VjhFhUN5_0),.clk(gclk));
	jdff dff_A_qjYREwnY3_0(.dout(w_dff_A_DesNHXqO3_0),.din(w_dff_A_qjYREwnY3_0),.clk(gclk));
	jdff dff_A_DesNHXqO3_0(.dout(w_dff_A_oROOZXXm2_0),.din(w_dff_A_DesNHXqO3_0),.clk(gclk));
	jdff dff_A_oROOZXXm2_0(.dout(w_dff_A_vqllTW0F0_0),.din(w_dff_A_oROOZXXm2_0),.clk(gclk));
	jdff dff_A_vqllTW0F0_0(.dout(G892),.din(w_dff_A_vqllTW0F0_0),.clk(gclk));
	jdff dff_A_QFHYc7Fj1_1(.dout(w_dff_A_PMZF4mUi7_0),.din(w_dff_A_QFHYc7Fj1_1),.clk(gclk));
	jdff dff_A_PMZF4mUi7_0(.dout(w_dff_A_uMG66Qip9_0),.din(w_dff_A_PMZF4mUi7_0),.clk(gclk));
	jdff dff_A_uMG66Qip9_0(.dout(w_dff_A_tBtDY7Dj9_0),.din(w_dff_A_uMG66Qip9_0),.clk(gclk));
	jdff dff_A_tBtDY7Dj9_0(.dout(w_dff_A_8tU4DtWU5_0),.din(w_dff_A_tBtDY7Dj9_0),.clk(gclk));
	jdff dff_A_8tU4DtWU5_0(.dout(w_dff_A_czryexAs0_0),.din(w_dff_A_8tU4DtWU5_0),.clk(gclk));
	jdff dff_A_czryexAs0_0(.dout(w_dff_A_NU64LTm80_0),.din(w_dff_A_czryexAs0_0),.clk(gclk));
	jdff dff_A_NU64LTm80_0(.dout(w_dff_A_OZfb0iRl5_0),.din(w_dff_A_NU64LTm80_0),.clk(gclk));
	jdff dff_A_OZfb0iRl5_0(.dout(w_dff_A_jquXzVdc4_0),.din(w_dff_A_OZfb0iRl5_0),.clk(gclk));
	jdff dff_A_jquXzVdc4_0(.dout(w_dff_A_IT3xMGJ89_0),.din(w_dff_A_jquXzVdc4_0),.clk(gclk));
	jdff dff_A_IT3xMGJ89_0(.dout(w_dff_A_FyGmX1Lx0_0),.din(w_dff_A_IT3xMGJ89_0),.clk(gclk));
	jdff dff_A_FyGmX1Lx0_0(.dout(w_dff_A_t4BVRV3q9_0),.din(w_dff_A_FyGmX1Lx0_0),.clk(gclk));
	jdff dff_A_t4BVRV3q9_0(.dout(w_dff_A_KEWsQdWT0_0),.din(w_dff_A_t4BVRV3q9_0),.clk(gclk));
	jdff dff_A_KEWsQdWT0_0(.dout(w_dff_A_fBF1V4431_0),.din(w_dff_A_KEWsQdWT0_0),.clk(gclk));
	jdff dff_A_fBF1V4431_0(.dout(w_dff_A_02EqBpfb9_0),.din(w_dff_A_fBF1V4431_0),.clk(gclk));
	jdff dff_A_02EqBpfb9_0(.dout(w_dff_A_yovzNn3U8_0),.din(w_dff_A_02EqBpfb9_0),.clk(gclk));
	jdff dff_A_yovzNn3U8_0(.dout(w_dff_A_9u5Ufmuo3_0),.din(w_dff_A_yovzNn3U8_0),.clk(gclk));
	jdff dff_A_9u5Ufmuo3_0(.dout(w_dff_A_pYnQYhqq5_0),.din(w_dff_A_9u5Ufmuo3_0),.clk(gclk));
	jdff dff_A_pYnQYhqq5_0(.dout(w_dff_A_4fMweFG82_0),.din(w_dff_A_pYnQYhqq5_0),.clk(gclk));
	jdff dff_A_4fMweFG82_0(.dout(w_dff_A_ndtvTD3M6_0),.din(w_dff_A_4fMweFG82_0),.clk(gclk));
	jdff dff_A_ndtvTD3M6_0(.dout(w_dff_A_XH45lJcj2_0),.din(w_dff_A_ndtvTD3M6_0),.clk(gclk));
	jdff dff_A_XH45lJcj2_0(.dout(w_dff_A_Rrs8FY0R6_0),.din(w_dff_A_XH45lJcj2_0),.clk(gclk));
	jdff dff_A_Rrs8FY0R6_0(.dout(w_dff_A_ShDWRVng2_0),.din(w_dff_A_Rrs8FY0R6_0),.clk(gclk));
	jdff dff_A_ShDWRVng2_0(.dout(w_dff_A_9UtbIp9q9_0),.din(w_dff_A_ShDWRVng2_0),.clk(gclk));
	jdff dff_A_9UtbIp9q9_0(.dout(w_dff_A_MikKOYaC1_0),.din(w_dff_A_9UtbIp9q9_0),.clk(gclk));
	jdff dff_A_MikKOYaC1_0(.dout(w_dff_A_aTsBRGqL6_0),.din(w_dff_A_MikKOYaC1_0),.clk(gclk));
	jdff dff_A_aTsBRGqL6_0(.dout(G887),.din(w_dff_A_aTsBRGqL6_0),.clk(gclk));
	jdff dff_A_0OPq6GU27_1(.dout(w_dff_A_ISi2XYXx9_0),.din(w_dff_A_0OPq6GU27_1),.clk(gclk));
	jdff dff_A_ISi2XYXx9_0(.dout(w_dff_A_XuQgYQ138_0),.din(w_dff_A_ISi2XYXx9_0),.clk(gclk));
	jdff dff_A_XuQgYQ138_0(.dout(w_dff_A_UBTHxJvq6_0),.din(w_dff_A_XuQgYQ138_0),.clk(gclk));
	jdff dff_A_UBTHxJvq6_0(.dout(w_dff_A_bhTwe7ii2_0),.din(w_dff_A_UBTHxJvq6_0),.clk(gclk));
	jdff dff_A_bhTwe7ii2_0(.dout(w_dff_A_0Drf1Qww0_0),.din(w_dff_A_bhTwe7ii2_0),.clk(gclk));
	jdff dff_A_0Drf1Qww0_0(.dout(w_dff_A_EbAhbqOP8_0),.din(w_dff_A_0Drf1Qww0_0),.clk(gclk));
	jdff dff_A_EbAhbqOP8_0(.dout(w_dff_A_sGW2EcJY2_0),.din(w_dff_A_EbAhbqOP8_0),.clk(gclk));
	jdff dff_A_sGW2EcJY2_0(.dout(w_dff_A_nH53o9AR5_0),.din(w_dff_A_sGW2EcJY2_0),.clk(gclk));
	jdff dff_A_nH53o9AR5_0(.dout(w_dff_A_uOnF7NKK8_0),.din(w_dff_A_nH53o9AR5_0),.clk(gclk));
	jdff dff_A_uOnF7NKK8_0(.dout(w_dff_A_PiVhECcY8_0),.din(w_dff_A_uOnF7NKK8_0),.clk(gclk));
	jdff dff_A_PiVhECcY8_0(.dout(w_dff_A_fV546wwq1_0),.din(w_dff_A_PiVhECcY8_0),.clk(gclk));
	jdff dff_A_fV546wwq1_0(.dout(w_dff_A_zUyqGHW02_0),.din(w_dff_A_fV546wwq1_0),.clk(gclk));
	jdff dff_A_zUyqGHW02_0(.dout(w_dff_A_v0fWeeZW3_0),.din(w_dff_A_zUyqGHW02_0),.clk(gclk));
	jdff dff_A_v0fWeeZW3_0(.dout(w_dff_A_7ujRWc1N2_0),.din(w_dff_A_v0fWeeZW3_0),.clk(gclk));
	jdff dff_A_7ujRWc1N2_0(.dout(w_dff_A_3GxMm94q8_0),.din(w_dff_A_7ujRWc1N2_0),.clk(gclk));
	jdff dff_A_3GxMm94q8_0(.dout(w_dff_A_EDVHbBsq2_0),.din(w_dff_A_3GxMm94q8_0),.clk(gclk));
	jdff dff_A_EDVHbBsq2_0(.dout(w_dff_A_BVvSRfeC8_0),.din(w_dff_A_EDVHbBsq2_0),.clk(gclk));
	jdff dff_A_BVvSRfeC8_0(.dout(w_dff_A_abvTzoZR6_0),.din(w_dff_A_BVvSRfeC8_0),.clk(gclk));
	jdff dff_A_abvTzoZR6_0(.dout(w_dff_A_zymTnHTE3_0),.din(w_dff_A_abvTzoZR6_0),.clk(gclk));
	jdff dff_A_zymTnHTE3_0(.dout(w_dff_A_7p8fuMN78_0),.din(w_dff_A_zymTnHTE3_0),.clk(gclk));
	jdff dff_A_7p8fuMN78_0(.dout(w_dff_A_VDEYP1cj6_0),.din(w_dff_A_7p8fuMN78_0),.clk(gclk));
	jdff dff_A_VDEYP1cj6_0(.dout(w_dff_A_gs9mOI0f8_0),.din(w_dff_A_VDEYP1cj6_0),.clk(gclk));
	jdff dff_A_gs9mOI0f8_0(.dout(w_dff_A_WmsrZvsf4_0),.din(w_dff_A_gs9mOI0f8_0),.clk(gclk));
	jdff dff_A_WmsrZvsf4_0(.dout(w_dff_A_QpbmHz4K1_0),.din(w_dff_A_WmsrZvsf4_0),.clk(gclk));
	jdff dff_A_QpbmHz4K1_0(.dout(G606),.din(w_dff_A_QpbmHz4K1_0),.clk(gclk));
	jdff dff_A_9LMyKtbq7_2(.dout(w_dff_A_LeX4LYJX0_0),.din(w_dff_A_9LMyKtbq7_2),.clk(gclk));
	jdff dff_A_LeX4LYJX0_0(.dout(w_dff_A_31sOqvSO5_0),.din(w_dff_A_LeX4LYJX0_0),.clk(gclk));
	jdff dff_A_31sOqvSO5_0(.dout(w_dff_A_feVftU9h6_0),.din(w_dff_A_31sOqvSO5_0),.clk(gclk));
	jdff dff_A_feVftU9h6_0(.dout(w_dff_A_xUGPZ3vK8_0),.din(w_dff_A_feVftU9h6_0),.clk(gclk));
	jdff dff_A_xUGPZ3vK8_0(.dout(w_dff_A_Mu1m9N2G5_0),.din(w_dff_A_xUGPZ3vK8_0),.clk(gclk));
	jdff dff_A_Mu1m9N2G5_0(.dout(w_dff_A_QvVAdbMb9_0),.din(w_dff_A_Mu1m9N2G5_0),.clk(gclk));
	jdff dff_A_QvVAdbMb9_0(.dout(w_dff_A_mz4tHFXy9_0),.din(w_dff_A_QvVAdbMb9_0),.clk(gclk));
	jdff dff_A_mz4tHFXy9_0(.dout(w_dff_A_ankZ8yng9_0),.din(w_dff_A_mz4tHFXy9_0),.clk(gclk));
	jdff dff_A_ankZ8yng9_0(.dout(w_dff_A_tQw9pSRx5_0),.din(w_dff_A_ankZ8yng9_0),.clk(gclk));
	jdff dff_A_tQw9pSRx5_0(.dout(w_dff_A_5D6J6niT6_0),.din(w_dff_A_tQw9pSRx5_0),.clk(gclk));
	jdff dff_A_5D6J6niT6_0(.dout(w_dff_A_4hyGW6N78_0),.din(w_dff_A_5D6J6niT6_0),.clk(gclk));
	jdff dff_A_4hyGW6N78_0(.dout(w_dff_A_HSU2GkO85_0),.din(w_dff_A_4hyGW6N78_0),.clk(gclk));
	jdff dff_A_HSU2GkO85_0(.dout(w_dff_A_rmPzrKzX1_0),.din(w_dff_A_HSU2GkO85_0),.clk(gclk));
	jdff dff_A_rmPzrKzX1_0(.dout(w_dff_A_8LjF2bIZ4_0),.din(w_dff_A_rmPzrKzX1_0),.clk(gclk));
	jdff dff_A_8LjF2bIZ4_0(.dout(w_dff_A_Qq1VabVP3_0),.din(w_dff_A_8LjF2bIZ4_0),.clk(gclk));
	jdff dff_A_Qq1VabVP3_0(.dout(w_dff_A_J8ETL6sl0_0),.din(w_dff_A_Qq1VabVP3_0),.clk(gclk));
	jdff dff_A_J8ETL6sl0_0(.dout(w_dff_A_pKy6pIv48_0),.din(w_dff_A_J8ETL6sl0_0),.clk(gclk));
	jdff dff_A_pKy6pIv48_0(.dout(w_dff_A_gYQTGHsH9_0),.din(w_dff_A_pKy6pIv48_0),.clk(gclk));
	jdff dff_A_gYQTGHsH9_0(.dout(w_dff_A_omIm2yxE2_0),.din(w_dff_A_gYQTGHsH9_0),.clk(gclk));
	jdff dff_A_omIm2yxE2_0(.dout(w_dff_A_IAowf1US3_0),.din(w_dff_A_omIm2yxE2_0),.clk(gclk));
	jdff dff_A_IAowf1US3_0(.dout(w_dff_A_JmMCQgqB9_0),.din(w_dff_A_IAowf1US3_0),.clk(gclk));
	jdff dff_A_JmMCQgqB9_0(.dout(w_dff_A_OotEsjpD2_0),.din(w_dff_A_JmMCQgqB9_0),.clk(gclk));
	jdff dff_A_OotEsjpD2_0(.dout(G656),.din(w_dff_A_OotEsjpD2_0),.clk(gclk));
	jdff dff_A_4FDeHSQK4_2(.dout(w_dff_A_53F08RXh9_0),.din(w_dff_A_4FDeHSQK4_2),.clk(gclk));
	jdff dff_A_53F08RXh9_0(.dout(w_dff_A_bwvFUUO72_0),.din(w_dff_A_53F08RXh9_0),.clk(gclk));
	jdff dff_A_bwvFUUO72_0(.dout(w_dff_A_A5EdTfQo3_0),.din(w_dff_A_bwvFUUO72_0),.clk(gclk));
	jdff dff_A_A5EdTfQo3_0(.dout(w_dff_A_ZFRSGBK33_0),.din(w_dff_A_A5EdTfQo3_0),.clk(gclk));
	jdff dff_A_ZFRSGBK33_0(.dout(w_dff_A_zWCgwJ4T9_0),.din(w_dff_A_ZFRSGBK33_0),.clk(gclk));
	jdff dff_A_zWCgwJ4T9_0(.dout(w_dff_A_YfNqVm6O9_0),.din(w_dff_A_zWCgwJ4T9_0),.clk(gclk));
	jdff dff_A_YfNqVm6O9_0(.dout(w_dff_A_5gVsKW0k9_0),.din(w_dff_A_YfNqVm6O9_0),.clk(gclk));
	jdff dff_A_5gVsKW0k9_0(.dout(w_dff_A_QrXXHDQH4_0),.din(w_dff_A_5gVsKW0k9_0),.clk(gclk));
	jdff dff_A_QrXXHDQH4_0(.dout(w_dff_A_xl3S76Rj6_0),.din(w_dff_A_QrXXHDQH4_0),.clk(gclk));
	jdff dff_A_xl3S76Rj6_0(.dout(w_dff_A_2RrXjq8U9_0),.din(w_dff_A_xl3S76Rj6_0),.clk(gclk));
	jdff dff_A_2RrXjq8U9_0(.dout(w_dff_A_gvcGSg713_0),.din(w_dff_A_2RrXjq8U9_0),.clk(gclk));
	jdff dff_A_gvcGSg713_0(.dout(w_dff_A_dOowzlRw3_0),.din(w_dff_A_gvcGSg713_0),.clk(gclk));
	jdff dff_A_dOowzlRw3_0(.dout(w_dff_A_aWPlizYh8_0),.din(w_dff_A_dOowzlRw3_0),.clk(gclk));
	jdff dff_A_aWPlizYh8_0(.dout(w_dff_A_s0gU8yuk9_0),.din(w_dff_A_aWPlizYh8_0),.clk(gclk));
	jdff dff_A_s0gU8yuk9_0(.dout(w_dff_A_aAet1x6W0_0),.din(w_dff_A_s0gU8yuk9_0),.clk(gclk));
	jdff dff_A_aAet1x6W0_0(.dout(w_dff_A_YnBY93x42_0),.din(w_dff_A_aAet1x6W0_0),.clk(gclk));
	jdff dff_A_YnBY93x42_0(.dout(w_dff_A_WmY2AXVv1_0),.din(w_dff_A_YnBY93x42_0),.clk(gclk));
	jdff dff_A_WmY2AXVv1_0(.dout(w_dff_A_4e7QblSY1_0),.din(w_dff_A_WmY2AXVv1_0),.clk(gclk));
	jdff dff_A_4e7QblSY1_0(.dout(w_dff_A_GgJPlDrh0_0),.din(w_dff_A_4e7QblSY1_0),.clk(gclk));
	jdff dff_A_GgJPlDrh0_0(.dout(w_dff_A_Q7wGKW2c0_0),.din(w_dff_A_GgJPlDrh0_0),.clk(gclk));
	jdff dff_A_Q7wGKW2c0_0(.dout(w_dff_A_aXxieiC35_0),.din(w_dff_A_Q7wGKW2c0_0),.clk(gclk));
	jdff dff_A_aXxieiC35_0(.dout(w_dff_A_4tE1sT3T7_0),.din(w_dff_A_aXxieiC35_0),.clk(gclk));
	jdff dff_A_4tE1sT3T7_0(.dout(w_dff_A_v0aZb5kz5_0),.din(w_dff_A_4tE1sT3T7_0),.clk(gclk));
	jdff dff_A_v0aZb5kz5_0(.dout(G809),.din(w_dff_A_v0aZb5kz5_0),.clk(gclk));
	jdff dff_A_uN1e9ym35_1(.dout(w_dff_A_DDE8BJzV5_0),.din(w_dff_A_uN1e9ym35_1),.clk(gclk));
	jdff dff_A_DDE8BJzV5_0(.dout(w_dff_A_TSonxKRY3_0),.din(w_dff_A_DDE8BJzV5_0),.clk(gclk));
	jdff dff_A_TSonxKRY3_0(.dout(w_dff_A_rCza6zCY6_0),.din(w_dff_A_TSonxKRY3_0),.clk(gclk));
	jdff dff_A_rCza6zCY6_0(.dout(w_dff_A_khmZ2pxx1_0),.din(w_dff_A_rCza6zCY6_0),.clk(gclk));
	jdff dff_A_khmZ2pxx1_0(.dout(w_dff_A_XngQgKQy3_0),.din(w_dff_A_khmZ2pxx1_0),.clk(gclk));
	jdff dff_A_XngQgKQy3_0(.dout(w_dff_A_7fnFMIBm4_0),.din(w_dff_A_XngQgKQy3_0),.clk(gclk));
	jdff dff_A_7fnFMIBm4_0(.dout(w_dff_A_AIDI0fd23_0),.din(w_dff_A_7fnFMIBm4_0),.clk(gclk));
	jdff dff_A_AIDI0fd23_0(.dout(w_dff_A_KgGs29KD8_0),.din(w_dff_A_AIDI0fd23_0),.clk(gclk));
	jdff dff_A_KgGs29KD8_0(.dout(w_dff_A_wEa3E1EL0_0),.din(w_dff_A_KgGs29KD8_0),.clk(gclk));
	jdff dff_A_wEa3E1EL0_0(.dout(w_dff_A_LKZzLQPY9_0),.din(w_dff_A_wEa3E1EL0_0),.clk(gclk));
	jdff dff_A_LKZzLQPY9_0(.dout(w_dff_A_e0xTxuDQ8_0),.din(w_dff_A_LKZzLQPY9_0),.clk(gclk));
	jdff dff_A_e0xTxuDQ8_0(.dout(w_dff_A_DqdAE0c33_0),.din(w_dff_A_e0xTxuDQ8_0),.clk(gclk));
	jdff dff_A_DqdAE0c33_0(.dout(w_dff_A_gbRStlEe3_0),.din(w_dff_A_DqdAE0c33_0),.clk(gclk));
	jdff dff_A_gbRStlEe3_0(.dout(w_dff_A_Zpg4qWUR8_0),.din(w_dff_A_gbRStlEe3_0),.clk(gclk));
	jdff dff_A_Zpg4qWUR8_0(.dout(w_dff_A_PDyuMfC12_0),.din(w_dff_A_Zpg4qWUR8_0),.clk(gclk));
	jdff dff_A_PDyuMfC12_0(.dout(w_dff_A_Zqu5CR5b2_0),.din(w_dff_A_PDyuMfC12_0),.clk(gclk));
	jdff dff_A_Zqu5CR5b2_0(.dout(w_dff_A_drXXU6Wl0_0),.din(w_dff_A_Zqu5CR5b2_0),.clk(gclk));
	jdff dff_A_drXXU6Wl0_0(.dout(w_dff_A_r8wfL2rL3_0),.din(w_dff_A_drXXU6Wl0_0),.clk(gclk));
	jdff dff_A_r8wfL2rL3_0(.dout(w_dff_A_x6ak8e884_0),.din(w_dff_A_r8wfL2rL3_0),.clk(gclk));
	jdff dff_A_x6ak8e884_0(.dout(w_dff_A_Gp1Zj1qL1_0),.din(w_dff_A_x6ak8e884_0),.clk(gclk));
	jdff dff_A_Gp1Zj1qL1_0(.dout(w_dff_A_dBzxZnWH7_0),.din(w_dff_A_Gp1Zj1qL1_0),.clk(gclk));
	jdff dff_A_dBzxZnWH7_0(.dout(w_dff_A_OES7JWNi8_0),.din(w_dff_A_dBzxZnWH7_0),.clk(gclk));
	jdff dff_A_OES7JWNi8_0(.dout(w_dff_A_6Vlmlz5H5_0),.din(w_dff_A_OES7JWNi8_0),.clk(gclk));
	jdff dff_A_6Vlmlz5H5_0(.dout(w_dff_A_9RerqaJa3_0),.din(w_dff_A_6Vlmlz5H5_0),.clk(gclk));
	jdff dff_A_9RerqaJa3_0(.dout(w_dff_A_EikSB4526_0),.din(w_dff_A_9RerqaJa3_0),.clk(gclk));
	jdff dff_A_EikSB4526_0(.dout(G993),.din(w_dff_A_EikSB4526_0),.clk(gclk));
	jdff dff_A_NnNpN7LE0_1(.dout(w_dff_A_98i8w2QX4_0),.din(w_dff_A_NnNpN7LE0_1),.clk(gclk));
	jdff dff_A_98i8w2QX4_0(.dout(w_dff_A_9dYQ0MBV4_0),.din(w_dff_A_98i8w2QX4_0),.clk(gclk));
	jdff dff_A_9dYQ0MBV4_0(.dout(w_dff_A_DhBOJ4mI0_0),.din(w_dff_A_9dYQ0MBV4_0),.clk(gclk));
	jdff dff_A_DhBOJ4mI0_0(.dout(w_dff_A_NOiHHKfc2_0),.din(w_dff_A_DhBOJ4mI0_0),.clk(gclk));
	jdff dff_A_NOiHHKfc2_0(.dout(w_dff_A_VTOlczNQ1_0),.din(w_dff_A_NOiHHKfc2_0),.clk(gclk));
	jdff dff_A_VTOlczNQ1_0(.dout(w_dff_A_KhdQQ4Ov4_0),.din(w_dff_A_VTOlczNQ1_0),.clk(gclk));
	jdff dff_A_KhdQQ4Ov4_0(.dout(w_dff_A_ZiODlsO86_0),.din(w_dff_A_KhdQQ4Ov4_0),.clk(gclk));
	jdff dff_A_ZiODlsO86_0(.dout(w_dff_A_jDwPP2oX9_0),.din(w_dff_A_ZiODlsO86_0),.clk(gclk));
	jdff dff_A_jDwPP2oX9_0(.dout(w_dff_A_wGH08fmO7_0),.din(w_dff_A_jDwPP2oX9_0),.clk(gclk));
	jdff dff_A_wGH08fmO7_0(.dout(w_dff_A_Ym82e2Zy0_0),.din(w_dff_A_wGH08fmO7_0),.clk(gclk));
	jdff dff_A_Ym82e2Zy0_0(.dout(w_dff_A_yseIjvsq8_0),.din(w_dff_A_Ym82e2Zy0_0),.clk(gclk));
	jdff dff_A_yseIjvsq8_0(.dout(w_dff_A_IlsbZwWv8_0),.din(w_dff_A_yseIjvsq8_0),.clk(gclk));
	jdff dff_A_IlsbZwWv8_0(.dout(w_dff_A_BoRetuJU2_0),.din(w_dff_A_IlsbZwWv8_0),.clk(gclk));
	jdff dff_A_BoRetuJU2_0(.dout(w_dff_A_DaNirjya4_0),.din(w_dff_A_BoRetuJU2_0),.clk(gclk));
	jdff dff_A_DaNirjya4_0(.dout(w_dff_A_NxuwoN3R6_0),.din(w_dff_A_DaNirjya4_0),.clk(gclk));
	jdff dff_A_NxuwoN3R6_0(.dout(w_dff_A_Cm3wGoB99_0),.din(w_dff_A_NxuwoN3R6_0),.clk(gclk));
	jdff dff_A_Cm3wGoB99_0(.dout(w_dff_A_Qc4MAacK3_0),.din(w_dff_A_Cm3wGoB99_0),.clk(gclk));
	jdff dff_A_Qc4MAacK3_0(.dout(w_dff_A_sJAmPAgd3_0),.din(w_dff_A_Qc4MAacK3_0),.clk(gclk));
	jdff dff_A_sJAmPAgd3_0(.dout(w_dff_A_RXmgIt4l6_0),.din(w_dff_A_sJAmPAgd3_0),.clk(gclk));
	jdff dff_A_RXmgIt4l6_0(.dout(w_dff_A_T7iJOIGc1_0),.din(w_dff_A_RXmgIt4l6_0),.clk(gclk));
	jdff dff_A_T7iJOIGc1_0(.dout(w_dff_A_VHaoAV704_0),.din(w_dff_A_T7iJOIGc1_0),.clk(gclk));
	jdff dff_A_VHaoAV704_0(.dout(w_dff_A_SEL3KXPi7_0),.din(w_dff_A_VHaoAV704_0),.clk(gclk));
	jdff dff_A_SEL3KXPi7_0(.dout(w_dff_A_rMQA6tWD0_0),.din(w_dff_A_SEL3KXPi7_0),.clk(gclk));
	jdff dff_A_rMQA6tWD0_0(.dout(w_dff_A_75qgGpF97_0),.din(w_dff_A_rMQA6tWD0_0),.clk(gclk));
	jdff dff_A_75qgGpF97_0(.dout(w_dff_A_6pcevl1s5_0),.din(w_dff_A_75qgGpF97_0),.clk(gclk));
	jdff dff_A_6pcevl1s5_0(.dout(G978),.din(w_dff_A_6pcevl1s5_0),.clk(gclk));
	jdff dff_A_2LtSmUnw2_1(.dout(w_dff_A_DCEKpMZe3_0),.din(w_dff_A_2LtSmUnw2_1),.clk(gclk));
	jdff dff_A_DCEKpMZe3_0(.dout(w_dff_A_0RrCnvrw0_0),.din(w_dff_A_DCEKpMZe3_0),.clk(gclk));
	jdff dff_A_0RrCnvrw0_0(.dout(w_dff_A_ucFluxaL0_0),.din(w_dff_A_0RrCnvrw0_0),.clk(gclk));
	jdff dff_A_ucFluxaL0_0(.dout(w_dff_A_JFZVaWzo0_0),.din(w_dff_A_ucFluxaL0_0),.clk(gclk));
	jdff dff_A_JFZVaWzo0_0(.dout(w_dff_A_xGJ73V7C3_0),.din(w_dff_A_JFZVaWzo0_0),.clk(gclk));
	jdff dff_A_xGJ73V7C3_0(.dout(w_dff_A_hXk3t87U7_0),.din(w_dff_A_xGJ73V7C3_0),.clk(gclk));
	jdff dff_A_hXk3t87U7_0(.dout(w_dff_A_lvOqVOJH5_0),.din(w_dff_A_hXk3t87U7_0),.clk(gclk));
	jdff dff_A_lvOqVOJH5_0(.dout(w_dff_A_Dj34yWJ18_0),.din(w_dff_A_lvOqVOJH5_0),.clk(gclk));
	jdff dff_A_Dj34yWJ18_0(.dout(w_dff_A_KRYBHC5Y6_0),.din(w_dff_A_Dj34yWJ18_0),.clk(gclk));
	jdff dff_A_KRYBHC5Y6_0(.dout(w_dff_A_4u9beA0C5_0),.din(w_dff_A_KRYBHC5Y6_0),.clk(gclk));
	jdff dff_A_4u9beA0C5_0(.dout(w_dff_A_w4d3SPld0_0),.din(w_dff_A_4u9beA0C5_0),.clk(gclk));
	jdff dff_A_w4d3SPld0_0(.dout(w_dff_A_ARXar45I3_0),.din(w_dff_A_w4d3SPld0_0),.clk(gclk));
	jdff dff_A_ARXar45I3_0(.dout(w_dff_A_SkSXS6uy7_0),.din(w_dff_A_ARXar45I3_0),.clk(gclk));
	jdff dff_A_SkSXS6uy7_0(.dout(w_dff_A_jiEc8ZSq2_0),.din(w_dff_A_SkSXS6uy7_0),.clk(gclk));
	jdff dff_A_jiEc8ZSq2_0(.dout(w_dff_A_XQ7Z9yFc3_0),.din(w_dff_A_jiEc8ZSq2_0),.clk(gclk));
	jdff dff_A_XQ7Z9yFc3_0(.dout(w_dff_A_9dvFI3ha0_0),.din(w_dff_A_XQ7Z9yFc3_0),.clk(gclk));
	jdff dff_A_9dvFI3ha0_0(.dout(w_dff_A_4Wv4Koqv0_0),.din(w_dff_A_9dvFI3ha0_0),.clk(gclk));
	jdff dff_A_4Wv4Koqv0_0(.dout(w_dff_A_XGyd3ihA6_0),.din(w_dff_A_4Wv4Koqv0_0),.clk(gclk));
	jdff dff_A_XGyd3ihA6_0(.dout(w_dff_A_UhiWgx794_0),.din(w_dff_A_XGyd3ihA6_0),.clk(gclk));
	jdff dff_A_UhiWgx794_0(.dout(w_dff_A_94BZuozg1_0),.din(w_dff_A_UhiWgx794_0),.clk(gclk));
	jdff dff_A_94BZuozg1_0(.dout(w_dff_A_prXiWfPG5_0),.din(w_dff_A_94BZuozg1_0),.clk(gclk));
	jdff dff_A_prXiWfPG5_0(.dout(w_dff_A_oW37fLM99_0),.din(w_dff_A_prXiWfPG5_0),.clk(gclk));
	jdff dff_A_oW37fLM99_0(.dout(w_dff_A_PRPlMr0e0_0),.din(w_dff_A_oW37fLM99_0),.clk(gclk));
	jdff dff_A_PRPlMr0e0_0(.dout(w_dff_A_7XjXvFRw8_0),.din(w_dff_A_PRPlMr0e0_0),.clk(gclk));
	jdff dff_A_7XjXvFRw8_0(.dout(w_dff_A_0kCIwMLz2_0),.din(w_dff_A_7XjXvFRw8_0),.clk(gclk));
	jdff dff_A_0kCIwMLz2_0(.dout(G949),.din(w_dff_A_0kCIwMLz2_0),.clk(gclk));
	jdff dff_A_bhCkHx8o1_1(.dout(w_dff_A_zLAD9MAs6_0),.din(w_dff_A_bhCkHx8o1_1),.clk(gclk));
	jdff dff_A_zLAD9MAs6_0(.dout(w_dff_A_b6PyrG9D0_0),.din(w_dff_A_zLAD9MAs6_0),.clk(gclk));
	jdff dff_A_b6PyrG9D0_0(.dout(w_dff_A_lvAjtu2Q0_0),.din(w_dff_A_b6PyrG9D0_0),.clk(gclk));
	jdff dff_A_lvAjtu2Q0_0(.dout(w_dff_A_T2xVdAGo9_0),.din(w_dff_A_lvAjtu2Q0_0),.clk(gclk));
	jdff dff_A_T2xVdAGo9_0(.dout(w_dff_A_jixHMTo23_0),.din(w_dff_A_T2xVdAGo9_0),.clk(gclk));
	jdff dff_A_jixHMTo23_0(.dout(w_dff_A_mECcdmDu5_0),.din(w_dff_A_jixHMTo23_0),.clk(gclk));
	jdff dff_A_mECcdmDu5_0(.dout(w_dff_A_FNhYLUNV5_0),.din(w_dff_A_mECcdmDu5_0),.clk(gclk));
	jdff dff_A_FNhYLUNV5_0(.dout(w_dff_A_8OQW41Jt0_0),.din(w_dff_A_FNhYLUNV5_0),.clk(gclk));
	jdff dff_A_8OQW41Jt0_0(.dout(w_dff_A_7yVhsTkT7_0),.din(w_dff_A_8OQW41Jt0_0),.clk(gclk));
	jdff dff_A_7yVhsTkT7_0(.dout(w_dff_A_AY4Qnx3m1_0),.din(w_dff_A_7yVhsTkT7_0),.clk(gclk));
	jdff dff_A_AY4Qnx3m1_0(.dout(w_dff_A_2KyOlAVx1_0),.din(w_dff_A_AY4Qnx3m1_0),.clk(gclk));
	jdff dff_A_2KyOlAVx1_0(.dout(w_dff_A_cGMDKwWw0_0),.din(w_dff_A_2KyOlAVx1_0),.clk(gclk));
	jdff dff_A_cGMDKwWw0_0(.dout(w_dff_A_b697pHxQ3_0),.din(w_dff_A_cGMDKwWw0_0),.clk(gclk));
	jdff dff_A_b697pHxQ3_0(.dout(w_dff_A_XwvzxxTH2_0),.din(w_dff_A_b697pHxQ3_0),.clk(gclk));
	jdff dff_A_XwvzxxTH2_0(.dout(w_dff_A_QEI5p7Ym3_0),.din(w_dff_A_XwvzxxTH2_0),.clk(gclk));
	jdff dff_A_QEI5p7Ym3_0(.dout(w_dff_A_i89gtJ4S1_0),.din(w_dff_A_QEI5p7Ym3_0),.clk(gclk));
	jdff dff_A_i89gtJ4S1_0(.dout(w_dff_A_hkTJ0VYW7_0),.din(w_dff_A_i89gtJ4S1_0),.clk(gclk));
	jdff dff_A_hkTJ0VYW7_0(.dout(w_dff_A_frv7p8y58_0),.din(w_dff_A_hkTJ0VYW7_0),.clk(gclk));
	jdff dff_A_frv7p8y58_0(.dout(w_dff_A_pX3Q8Uax0_0),.din(w_dff_A_frv7p8y58_0),.clk(gclk));
	jdff dff_A_pX3Q8Uax0_0(.dout(w_dff_A_X8Oysb7a4_0),.din(w_dff_A_pX3Q8Uax0_0),.clk(gclk));
	jdff dff_A_X8Oysb7a4_0(.dout(w_dff_A_SJshBxdt8_0),.din(w_dff_A_X8Oysb7a4_0),.clk(gclk));
	jdff dff_A_SJshBxdt8_0(.dout(w_dff_A_wgAF5rYA2_0),.din(w_dff_A_SJshBxdt8_0),.clk(gclk));
	jdff dff_A_wgAF5rYA2_0(.dout(w_dff_A_nCKnPfb64_0),.din(w_dff_A_wgAF5rYA2_0),.clk(gclk));
	jdff dff_A_nCKnPfb64_0(.dout(w_dff_A_CGUXvuJH3_0),.din(w_dff_A_nCKnPfb64_0),.clk(gclk));
	jdff dff_A_CGUXvuJH3_0(.dout(w_dff_A_SZHdqKEr8_0),.din(w_dff_A_CGUXvuJH3_0),.clk(gclk));
	jdff dff_A_SZHdqKEr8_0(.dout(G939),.din(w_dff_A_SZHdqKEr8_0),.clk(gclk));
	jdff dff_A_RvDEgF9N8_1(.dout(w_dff_A_IznpfcOq9_0),.din(w_dff_A_RvDEgF9N8_1),.clk(gclk));
	jdff dff_A_IznpfcOq9_0(.dout(w_dff_A_uC2juEjC4_0),.din(w_dff_A_IznpfcOq9_0),.clk(gclk));
	jdff dff_A_uC2juEjC4_0(.dout(w_dff_A_BEDOENFC3_0),.din(w_dff_A_uC2juEjC4_0),.clk(gclk));
	jdff dff_A_BEDOENFC3_0(.dout(w_dff_A_QjCXCqBQ4_0),.din(w_dff_A_BEDOENFC3_0),.clk(gclk));
	jdff dff_A_QjCXCqBQ4_0(.dout(w_dff_A_o8QopJDN1_0),.din(w_dff_A_QjCXCqBQ4_0),.clk(gclk));
	jdff dff_A_o8QopJDN1_0(.dout(w_dff_A_vKCqEmq32_0),.din(w_dff_A_o8QopJDN1_0),.clk(gclk));
	jdff dff_A_vKCqEmq32_0(.dout(w_dff_A_zqgyP5oj2_0),.din(w_dff_A_vKCqEmq32_0),.clk(gclk));
	jdff dff_A_zqgyP5oj2_0(.dout(w_dff_A_Mm1v7Vpq4_0),.din(w_dff_A_zqgyP5oj2_0),.clk(gclk));
	jdff dff_A_Mm1v7Vpq4_0(.dout(w_dff_A_SEvXjhlY9_0),.din(w_dff_A_Mm1v7Vpq4_0),.clk(gclk));
	jdff dff_A_SEvXjhlY9_0(.dout(w_dff_A_aV8lqEBR2_0),.din(w_dff_A_SEvXjhlY9_0),.clk(gclk));
	jdff dff_A_aV8lqEBR2_0(.dout(w_dff_A_gtfNUY6z8_0),.din(w_dff_A_aV8lqEBR2_0),.clk(gclk));
	jdff dff_A_gtfNUY6z8_0(.dout(w_dff_A_WgVb8MiY2_0),.din(w_dff_A_gtfNUY6z8_0),.clk(gclk));
	jdff dff_A_WgVb8MiY2_0(.dout(w_dff_A_utU4WP8j4_0),.din(w_dff_A_WgVb8MiY2_0),.clk(gclk));
	jdff dff_A_utU4WP8j4_0(.dout(w_dff_A_wYt4UxtS9_0),.din(w_dff_A_utU4WP8j4_0),.clk(gclk));
	jdff dff_A_wYt4UxtS9_0(.dout(w_dff_A_LChqDAVs6_0),.din(w_dff_A_wYt4UxtS9_0),.clk(gclk));
	jdff dff_A_LChqDAVs6_0(.dout(w_dff_A_WFQUi4jm7_0),.din(w_dff_A_LChqDAVs6_0),.clk(gclk));
	jdff dff_A_WFQUi4jm7_0(.dout(w_dff_A_fh5MCp210_0),.din(w_dff_A_WFQUi4jm7_0),.clk(gclk));
	jdff dff_A_fh5MCp210_0(.dout(w_dff_A_3BRew9G51_0),.din(w_dff_A_fh5MCp210_0),.clk(gclk));
	jdff dff_A_3BRew9G51_0(.dout(w_dff_A_7voMf0we2_0),.din(w_dff_A_3BRew9G51_0),.clk(gclk));
	jdff dff_A_7voMf0we2_0(.dout(w_dff_A_aMG0QwnA1_0),.din(w_dff_A_7voMf0we2_0),.clk(gclk));
	jdff dff_A_aMG0QwnA1_0(.dout(w_dff_A_rhrrGLpy9_0),.din(w_dff_A_aMG0QwnA1_0),.clk(gclk));
	jdff dff_A_rhrrGLpy9_0(.dout(w_dff_A_6ajUOm4r9_0),.din(w_dff_A_rhrrGLpy9_0),.clk(gclk));
	jdff dff_A_6ajUOm4r9_0(.dout(w_dff_A_OCYlJY7m3_0),.din(w_dff_A_6ajUOm4r9_0),.clk(gclk));
	jdff dff_A_OCYlJY7m3_0(.dout(w_dff_A_uHcHn3hs4_0),.din(w_dff_A_OCYlJY7m3_0),.clk(gclk));
	jdff dff_A_uHcHn3hs4_0(.dout(w_dff_A_qZ1mA9zs2_0),.din(w_dff_A_uHcHn3hs4_0),.clk(gclk));
	jdff dff_A_qZ1mA9zs2_0(.dout(G889),.din(w_dff_A_qZ1mA9zs2_0),.clk(gclk));
	jdff dff_A_T8dVu50g8_1(.dout(w_dff_A_zCnTskqc8_0),.din(w_dff_A_T8dVu50g8_1),.clk(gclk));
	jdff dff_A_zCnTskqc8_0(.dout(w_dff_A_gHTbkyaV1_0),.din(w_dff_A_zCnTskqc8_0),.clk(gclk));
	jdff dff_A_gHTbkyaV1_0(.dout(w_dff_A_olhd6I4n0_0),.din(w_dff_A_gHTbkyaV1_0),.clk(gclk));
	jdff dff_A_olhd6I4n0_0(.dout(w_dff_A_wPRKyTpU9_0),.din(w_dff_A_olhd6I4n0_0),.clk(gclk));
	jdff dff_A_wPRKyTpU9_0(.dout(w_dff_A_Hx7mchhX6_0),.din(w_dff_A_wPRKyTpU9_0),.clk(gclk));
	jdff dff_A_Hx7mchhX6_0(.dout(w_dff_A_FNdUpmAq0_0),.din(w_dff_A_Hx7mchhX6_0),.clk(gclk));
	jdff dff_A_FNdUpmAq0_0(.dout(w_dff_A_JpvWkjLX2_0),.din(w_dff_A_FNdUpmAq0_0),.clk(gclk));
	jdff dff_A_JpvWkjLX2_0(.dout(w_dff_A_6kbN3b4b6_0),.din(w_dff_A_JpvWkjLX2_0),.clk(gclk));
	jdff dff_A_6kbN3b4b6_0(.dout(w_dff_A_9TxPnvMs2_0),.din(w_dff_A_6kbN3b4b6_0),.clk(gclk));
	jdff dff_A_9TxPnvMs2_0(.dout(w_dff_A_jyClKqdg3_0),.din(w_dff_A_9TxPnvMs2_0),.clk(gclk));
	jdff dff_A_jyClKqdg3_0(.dout(w_dff_A_C72m2Eqj5_0),.din(w_dff_A_jyClKqdg3_0),.clk(gclk));
	jdff dff_A_C72m2Eqj5_0(.dout(w_dff_A_GUGD6aYS7_0),.din(w_dff_A_C72m2Eqj5_0),.clk(gclk));
	jdff dff_A_GUGD6aYS7_0(.dout(w_dff_A_tqigecYc7_0),.din(w_dff_A_GUGD6aYS7_0),.clk(gclk));
	jdff dff_A_tqigecYc7_0(.dout(w_dff_A_ECmDm9Ct1_0),.din(w_dff_A_tqigecYc7_0),.clk(gclk));
	jdff dff_A_ECmDm9Ct1_0(.dout(w_dff_A_iCCmfY0J1_0),.din(w_dff_A_ECmDm9Ct1_0),.clk(gclk));
	jdff dff_A_iCCmfY0J1_0(.dout(w_dff_A_eM0jEiUq3_0),.din(w_dff_A_iCCmfY0J1_0),.clk(gclk));
	jdff dff_A_eM0jEiUq3_0(.dout(w_dff_A_4wD3UChI2_0),.din(w_dff_A_eM0jEiUq3_0),.clk(gclk));
	jdff dff_A_4wD3UChI2_0(.dout(w_dff_A_6cuahdtq3_0),.din(w_dff_A_4wD3UChI2_0),.clk(gclk));
	jdff dff_A_6cuahdtq3_0(.dout(w_dff_A_bARsrghJ2_0),.din(w_dff_A_6cuahdtq3_0),.clk(gclk));
	jdff dff_A_bARsrghJ2_0(.dout(w_dff_A_bYhM0UFD5_0),.din(w_dff_A_bARsrghJ2_0),.clk(gclk));
	jdff dff_A_bYhM0UFD5_0(.dout(w_dff_A_2ntibkXR3_0),.din(w_dff_A_bYhM0UFD5_0),.clk(gclk));
	jdff dff_A_2ntibkXR3_0(.dout(w_dff_A_cgYWLNPD1_0),.din(w_dff_A_2ntibkXR3_0),.clk(gclk));
	jdff dff_A_cgYWLNPD1_0(.dout(w_dff_A_HVpuMc0R9_0),.din(w_dff_A_cgYWLNPD1_0),.clk(gclk));
	jdff dff_A_HVpuMc0R9_0(.dout(w_dff_A_ThLUgkNN4_0),.din(w_dff_A_HVpuMc0R9_0),.clk(gclk));
	jdff dff_A_ThLUgkNN4_0(.dout(G593),.din(w_dff_A_ThLUgkNN4_0),.clk(gclk));
	jdff dff_A_tjW8NLMX1_2(.dout(w_dff_A_H9TNAipS8_0),.din(w_dff_A_tjW8NLMX1_2),.clk(gclk));
	jdff dff_A_H9TNAipS8_0(.dout(w_dff_A_sil2BaHk4_0),.din(w_dff_A_H9TNAipS8_0),.clk(gclk));
	jdff dff_A_sil2BaHk4_0(.dout(w_dff_A_VLwvdYqM6_0),.din(w_dff_A_sil2BaHk4_0),.clk(gclk));
	jdff dff_A_VLwvdYqM6_0(.dout(w_dff_A_rX4nh5r81_0),.din(w_dff_A_VLwvdYqM6_0),.clk(gclk));
	jdff dff_A_rX4nh5r81_0(.dout(w_dff_A_vch1eA7O4_0),.din(w_dff_A_rX4nh5r81_0),.clk(gclk));
	jdff dff_A_vch1eA7O4_0(.dout(w_dff_A_7Uklk3uY4_0),.din(w_dff_A_vch1eA7O4_0),.clk(gclk));
	jdff dff_A_7Uklk3uY4_0(.dout(w_dff_A_hl8XfH9q8_0),.din(w_dff_A_7Uklk3uY4_0),.clk(gclk));
	jdff dff_A_hl8XfH9q8_0(.dout(w_dff_A_dY4JM8Ma9_0),.din(w_dff_A_hl8XfH9q8_0),.clk(gclk));
	jdff dff_A_dY4JM8Ma9_0(.dout(w_dff_A_GZ03g1l60_0),.din(w_dff_A_dY4JM8Ma9_0),.clk(gclk));
	jdff dff_A_GZ03g1l60_0(.dout(w_dff_A_gWiapdnz4_0),.din(w_dff_A_GZ03g1l60_0),.clk(gclk));
	jdff dff_A_gWiapdnz4_0(.dout(w_dff_A_jDBS4Kto3_0),.din(w_dff_A_gWiapdnz4_0),.clk(gclk));
	jdff dff_A_jDBS4Kto3_0(.dout(w_dff_A_P93ZEZVW4_0),.din(w_dff_A_jDBS4Kto3_0),.clk(gclk));
	jdff dff_A_P93ZEZVW4_0(.dout(w_dff_A_lg3M9YNX1_0),.din(w_dff_A_P93ZEZVW4_0),.clk(gclk));
	jdff dff_A_lg3M9YNX1_0(.dout(w_dff_A_qXoz65Xu8_0),.din(w_dff_A_lg3M9YNX1_0),.clk(gclk));
	jdff dff_A_qXoz65Xu8_0(.dout(w_dff_A_XUmZkIFP7_0),.din(w_dff_A_qXoz65Xu8_0),.clk(gclk));
	jdff dff_A_XUmZkIFP7_0(.dout(w_dff_A_AQvfuaaX8_0),.din(w_dff_A_XUmZkIFP7_0),.clk(gclk));
	jdff dff_A_AQvfuaaX8_0(.dout(w_dff_A_kg737fNl7_0),.din(w_dff_A_AQvfuaaX8_0),.clk(gclk));
	jdff dff_A_kg737fNl7_0(.dout(w_dff_A_SNaRIK6p4_0),.din(w_dff_A_kg737fNl7_0),.clk(gclk));
	jdff dff_A_SNaRIK6p4_0(.dout(w_dff_A_Wkobyo4c0_0),.din(w_dff_A_SNaRIK6p4_0),.clk(gclk));
	jdff dff_A_Wkobyo4c0_0(.dout(w_dff_A_6aUo4ehg0_0),.din(w_dff_A_Wkobyo4c0_0),.clk(gclk));
	jdff dff_A_6aUo4ehg0_0(.dout(w_dff_A_kxfuJvZt2_0),.din(w_dff_A_6aUo4ehg0_0),.clk(gclk));
	jdff dff_A_kxfuJvZt2_0(.dout(G636),.din(w_dff_A_kxfuJvZt2_0),.clk(gclk));
	jdff dff_A_uZFyizaT3_2(.dout(w_dff_A_Iup5Etr22_0),.din(w_dff_A_uZFyizaT3_2),.clk(gclk));
	jdff dff_A_Iup5Etr22_0(.dout(w_dff_A_zEyb8kbB2_0),.din(w_dff_A_Iup5Etr22_0),.clk(gclk));
	jdff dff_A_zEyb8kbB2_0(.dout(w_dff_A_KMKmbzve9_0),.din(w_dff_A_zEyb8kbB2_0),.clk(gclk));
	jdff dff_A_KMKmbzve9_0(.dout(w_dff_A_tCRS59BQ5_0),.din(w_dff_A_KMKmbzve9_0),.clk(gclk));
	jdff dff_A_tCRS59BQ5_0(.dout(w_dff_A_3A0r1Zwr9_0),.din(w_dff_A_tCRS59BQ5_0),.clk(gclk));
	jdff dff_A_3A0r1Zwr9_0(.dout(w_dff_A_ynd2r14n7_0),.din(w_dff_A_3A0r1Zwr9_0),.clk(gclk));
	jdff dff_A_ynd2r14n7_0(.dout(w_dff_A_9QrrjaJT4_0),.din(w_dff_A_ynd2r14n7_0),.clk(gclk));
	jdff dff_A_9QrrjaJT4_0(.dout(w_dff_A_ozVDdAKz4_0),.din(w_dff_A_9QrrjaJT4_0),.clk(gclk));
	jdff dff_A_ozVDdAKz4_0(.dout(w_dff_A_3oAHYtvh7_0),.din(w_dff_A_ozVDdAKz4_0),.clk(gclk));
	jdff dff_A_3oAHYtvh7_0(.dout(w_dff_A_O0EBbhyD2_0),.din(w_dff_A_3oAHYtvh7_0),.clk(gclk));
	jdff dff_A_O0EBbhyD2_0(.dout(w_dff_A_SgG66Y1N3_0),.din(w_dff_A_O0EBbhyD2_0),.clk(gclk));
	jdff dff_A_SgG66Y1N3_0(.dout(w_dff_A_FR8mPSDU0_0),.din(w_dff_A_SgG66Y1N3_0),.clk(gclk));
	jdff dff_A_FR8mPSDU0_0(.dout(w_dff_A_EZgT09lv2_0),.din(w_dff_A_FR8mPSDU0_0),.clk(gclk));
	jdff dff_A_EZgT09lv2_0(.dout(w_dff_A_mdVCiKD18_0),.din(w_dff_A_EZgT09lv2_0),.clk(gclk));
	jdff dff_A_mdVCiKD18_0(.dout(w_dff_A_pLRXoKy13_0),.din(w_dff_A_mdVCiKD18_0),.clk(gclk));
	jdff dff_A_pLRXoKy13_0(.dout(w_dff_A_ilRRf97M4_0),.din(w_dff_A_pLRXoKy13_0),.clk(gclk));
	jdff dff_A_ilRRf97M4_0(.dout(w_dff_A_A3p5oRWj4_0),.din(w_dff_A_ilRRf97M4_0),.clk(gclk));
	jdff dff_A_A3p5oRWj4_0(.dout(w_dff_A_oHAqSUbo6_0),.din(w_dff_A_A3p5oRWj4_0),.clk(gclk));
	jdff dff_A_oHAqSUbo6_0(.dout(w_dff_A_xrM4FbYP1_0),.din(w_dff_A_oHAqSUbo6_0),.clk(gclk));
	jdff dff_A_xrM4FbYP1_0(.dout(w_dff_A_10oEFGMw0_0),.din(w_dff_A_xrM4FbYP1_0),.clk(gclk));
	jdff dff_A_10oEFGMw0_0(.dout(w_dff_A_IDmsZhwS0_0),.din(w_dff_A_10oEFGMw0_0),.clk(gclk));
	jdff dff_A_IDmsZhwS0_0(.dout(G704),.din(w_dff_A_IDmsZhwS0_0),.clk(gclk));
	jdff dff_A_aInYLOFA7_2(.dout(w_dff_A_ZzjTEjGE7_0),.din(w_dff_A_aInYLOFA7_2),.clk(gclk));
	jdff dff_A_ZzjTEjGE7_0(.dout(w_dff_A_hvGCZTZv2_0),.din(w_dff_A_ZzjTEjGE7_0),.clk(gclk));
	jdff dff_A_hvGCZTZv2_0(.dout(w_dff_A_dk8TRHFN4_0),.din(w_dff_A_hvGCZTZv2_0),.clk(gclk));
	jdff dff_A_dk8TRHFN4_0(.dout(w_dff_A_3Ga9Nzbe8_0),.din(w_dff_A_dk8TRHFN4_0),.clk(gclk));
	jdff dff_A_3Ga9Nzbe8_0(.dout(w_dff_A_DBBTDaqh3_0),.din(w_dff_A_3Ga9Nzbe8_0),.clk(gclk));
	jdff dff_A_DBBTDaqh3_0(.dout(w_dff_A_ACcmO2X72_0),.din(w_dff_A_DBBTDaqh3_0),.clk(gclk));
	jdff dff_A_ACcmO2X72_0(.dout(w_dff_A_ORXd5Uni3_0),.din(w_dff_A_ACcmO2X72_0),.clk(gclk));
	jdff dff_A_ORXd5Uni3_0(.dout(w_dff_A_qkeM14Wh7_0),.din(w_dff_A_ORXd5Uni3_0),.clk(gclk));
	jdff dff_A_qkeM14Wh7_0(.dout(w_dff_A_HeTKmtDF6_0),.din(w_dff_A_qkeM14Wh7_0),.clk(gclk));
	jdff dff_A_HeTKmtDF6_0(.dout(w_dff_A_aWji6Cq39_0),.din(w_dff_A_HeTKmtDF6_0),.clk(gclk));
	jdff dff_A_aWji6Cq39_0(.dout(w_dff_A_uuD7Po8Z1_0),.din(w_dff_A_aWji6Cq39_0),.clk(gclk));
	jdff dff_A_uuD7Po8Z1_0(.dout(w_dff_A_5GOF8sjO1_0),.din(w_dff_A_uuD7Po8Z1_0),.clk(gclk));
	jdff dff_A_5GOF8sjO1_0(.dout(w_dff_A_4GQM5DdY2_0),.din(w_dff_A_5GOF8sjO1_0),.clk(gclk));
	jdff dff_A_4GQM5DdY2_0(.dout(w_dff_A_ry4Va7jZ7_0),.din(w_dff_A_4GQM5DdY2_0),.clk(gclk));
	jdff dff_A_ry4Va7jZ7_0(.dout(w_dff_A_DIqvilCI7_0),.din(w_dff_A_ry4Va7jZ7_0),.clk(gclk));
	jdff dff_A_DIqvilCI7_0(.dout(w_dff_A_a4WbtcNh0_0),.din(w_dff_A_DIqvilCI7_0),.clk(gclk));
	jdff dff_A_a4WbtcNh0_0(.dout(w_dff_A_TvK4fqcj2_0),.din(w_dff_A_a4WbtcNh0_0),.clk(gclk));
	jdff dff_A_TvK4fqcj2_0(.dout(w_dff_A_w9GpjKFG1_0),.din(w_dff_A_TvK4fqcj2_0),.clk(gclk));
	jdff dff_A_w9GpjKFG1_0(.dout(w_dff_A_g32NSzLX6_0),.din(w_dff_A_w9GpjKFG1_0),.clk(gclk));
	jdff dff_A_g32NSzLX6_0(.dout(w_dff_A_IFl1JOmu2_0),.din(w_dff_A_g32NSzLX6_0),.clk(gclk));
	jdff dff_A_IFl1JOmu2_0(.dout(w_dff_A_Hq8CUuOH4_0),.din(w_dff_A_IFl1JOmu2_0),.clk(gclk));
	jdff dff_A_Hq8CUuOH4_0(.dout(G717),.din(w_dff_A_Hq8CUuOH4_0),.clk(gclk));
	jdff dff_A_1RnTGjF92_2(.dout(w_dff_A_XpeFdbpX0_0),.din(w_dff_A_1RnTGjF92_2),.clk(gclk));
	jdff dff_A_XpeFdbpX0_0(.dout(w_dff_A_qXnvJGO68_0),.din(w_dff_A_XpeFdbpX0_0),.clk(gclk));
	jdff dff_A_qXnvJGO68_0(.dout(w_dff_A_hPdSzwCK3_0),.din(w_dff_A_qXnvJGO68_0),.clk(gclk));
	jdff dff_A_hPdSzwCK3_0(.dout(w_dff_A_Aw2K0WOu6_0),.din(w_dff_A_hPdSzwCK3_0),.clk(gclk));
	jdff dff_A_Aw2K0WOu6_0(.dout(w_dff_A_Lim1RbxU1_0),.din(w_dff_A_Aw2K0WOu6_0),.clk(gclk));
	jdff dff_A_Lim1RbxU1_0(.dout(w_dff_A_gVqOoBCH6_0),.din(w_dff_A_Lim1RbxU1_0),.clk(gclk));
	jdff dff_A_gVqOoBCH6_0(.dout(w_dff_A_clBYr3K46_0),.din(w_dff_A_gVqOoBCH6_0),.clk(gclk));
	jdff dff_A_clBYr3K46_0(.dout(w_dff_A_k5oBvWcm8_0),.din(w_dff_A_clBYr3K46_0),.clk(gclk));
	jdff dff_A_k5oBvWcm8_0(.dout(w_dff_A_nV9mWPoL6_0),.din(w_dff_A_k5oBvWcm8_0),.clk(gclk));
	jdff dff_A_nV9mWPoL6_0(.dout(w_dff_A_vgpmPwJH4_0),.din(w_dff_A_nV9mWPoL6_0),.clk(gclk));
	jdff dff_A_vgpmPwJH4_0(.dout(w_dff_A_tagrcOs30_0),.din(w_dff_A_vgpmPwJH4_0),.clk(gclk));
	jdff dff_A_tagrcOs30_0(.dout(w_dff_A_IQ12Qa1e2_0),.din(w_dff_A_tagrcOs30_0),.clk(gclk));
	jdff dff_A_IQ12Qa1e2_0(.dout(w_dff_A_UWdADaUp5_0),.din(w_dff_A_IQ12Qa1e2_0),.clk(gclk));
	jdff dff_A_UWdADaUp5_0(.dout(w_dff_A_Hk7d1xco6_0),.din(w_dff_A_UWdADaUp5_0),.clk(gclk));
	jdff dff_A_Hk7d1xco6_0(.dout(w_dff_A_G54k42aC6_0),.din(w_dff_A_Hk7d1xco6_0),.clk(gclk));
	jdff dff_A_G54k42aC6_0(.dout(w_dff_A_heO1fFTY3_0),.din(w_dff_A_G54k42aC6_0),.clk(gclk));
	jdff dff_A_heO1fFTY3_0(.dout(w_dff_A_zDmiktN89_0),.din(w_dff_A_heO1fFTY3_0),.clk(gclk));
	jdff dff_A_zDmiktN89_0(.dout(w_dff_A_4u5QF0U34_0),.din(w_dff_A_zDmiktN89_0),.clk(gclk));
	jdff dff_A_4u5QF0U34_0(.dout(w_dff_A_HVzwcJTv6_0),.din(w_dff_A_4u5QF0U34_0),.clk(gclk));
	jdff dff_A_HVzwcJTv6_0(.dout(w_dff_A_WK95aYuy6_0),.din(w_dff_A_HVzwcJTv6_0),.clk(gclk));
	jdff dff_A_WK95aYuy6_0(.dout(w_dff_A_dU76sXvb9_0),.din(w_dff_A_WK95aYuy6_0),.clk(gclk));
	jdff dff_A_dU76sXvb9_0(.dout(w_dff_A_jHzqXZsV3_0),.din(w_dff_A_dU76sXvb9_0),.clk(gclk));
	jdff dff_A_jHzqXZsV3_0(.dout(G820),.din(w_dff_A_jHzqXZsV3_0),.clk(gclk));
	jdff dff_A_MTvHxVse2_2(.dout(w_dff_A_hBJW0UE92_0),.din(w_dff_A_MTvHxVse2_2),.clk(gclk));
	jdff dff_A_hBJW0UE92_0(.dout(w_dff_A_dy8GyFLw3_0),.din(w_dff_A_hBJW0UE92_0),.clk(gclk));
	jdff dff_A_dy8GyFLw3_0(.dout(w_dff_A_iPZrgL0e7_0),.din(w_dff_A_dy8GyFLw3_0),.clk(gclk));
	jdff dff_A_iPZrgL0e7_0(.dout(w_dff_A_vYlvHLsT8_0),.din(w_dff_A_iPZrgL0e7_0),.clk(gclk));
	jdff dff_A_vYlvHLsT8_0(.dout(w_dff_A_GaaDZ0Cp9_0),.din(w_dff_A_vYlvHLsT8_0),.clk(gclk));
	jdff dff_A_GaaDZ0Cp9_0(.dout(w_dff_A_T47ab6ca4_0),.din(w_dff_A_GaaDZ0Cp9_0),.clk(gclk));
	jdff dff_A_T47ab6ca4_0(.dout(w_dff_A_jYjs7tBs0_0),.din(w_dff_A_T47ab6ca4_0),.clk(gclk));
	jdff dff_A_jYjs7tBs0_0(.dout(w_dff_A_8hUwGXOE5_0),.din(w_dff_A_jYjs7tBs0_0),.clk(gclk));
	jdff dff_A_8hUwGXOE5_0(.dout(w_dff_A_v7nK7nE98_0),.din(w_dff_A_8hUwGXOE5_0),.clk(gclk));
	jdff dff_A_v7nK7nE98_0(.dout(w_dff_A_wrw7TbOF9_0),.din(w_dff_A_v7nK7nE98_0),.clk(gclk));
	jdff dff_A_wrw7TbOF9_0(.dout(w_dff_A_wztYHFfo8_0),.din(w_dff_A_wrw7TbOF9_0),.clk(gclk));
	jdff dff_A_wztYHFfo8_0(.dout(w_dff_A_UAx68KMz9_0),.din(w_dff_A_wztYHFfo8_0),.clk(gclk));
	jdff dff_A_UAx68KMz9_0(.dout(w_dff_A_Vl0CtV079_0),.din(w_dff_A_UAx68KMz9_0),.clk(gclk));
	jdff dff_A_Vl0CtV079_0(.dout(w_dff_A_2cPrXCWR7_0),.din(w_dff_A_Vl0CtV079_0),.clk(gclk));
	jdff dff_A_2cPrXCWR7_0(.dout(w_dff_A_F84Qf7T07_0),.din(w_dff_A_2cPrXCWR7_0),.clk(gclk));
	jdff dff_A_F84Qf7T07_0(.dout(w_dff_A_CyKOGwFh5_0),.din(w_dff_A_F84Qf7T07_0),.clk(gclk));
	jdff dff_A_CyKOGwFh5_0(.dout(w_dff_A_IdE90A2W3_0),.din(w_dff_A_CyKOGwFh5_0),.clk(gclk));
	jdff dff_A_IdE90A2W3_0(.dout(w_dff_A_AbukKjR94_0),.din(w_dff_A_IdE90A2W3_0),.clk(gclk));
	jdff dff_A_AbukKjR94_0(.dout(w_dff_A_nRVSS5K52_0),.din(w_dff_A_AbukKjR94_0),.clk(gclk));
	jdff dff_A_nRVSS5K52_0(.dout(w_dff_A_uxirQxCC7_0),.din(w_dff_A_nRVSS5K52_0),.clk(gclk));
	jdff dff_A_uxirQxCC7_0(.dout(G639),.din(w_dff_A_uxirQxCC7_0),.clk(gclk));
	jdff dff_A_QgILRn1A0_2(.dout(w_dff_A_rJEdO5Bd8_0),.din(w_dff_A_QgILRn1A0_2),.clk(gclk));
	jdff dff_A_rJEdO5Bd8_0(.dout(w_dff_A_ONVyIf2B8_0),.din(w_dff_A_rJEdO5Bd8_0),.clk(gclk));
	jdff dff_A_ONVyIf2B8_0(.dout(w_dff_A_Diyd9NdS1_0),.din(w_dff_A_ONVyIf2B8_0),.clk(gclk));
	jdff dff_A_Diyd9NdS1_0(.dout(w_dff_A_YFEfdFOq8_0),.din(w_dff_A_Diyd9NdS1_0),.clk(gclk));
	jdff dff_A_YFEfdFOq8_0(.dout(w_dff_A_nsDddu9i0_0),.din(w_dff_A_YFEfdFOq8_0),.clk(gclk));
	jdff dff_A_nsDddu9i0_0(.dout(w_dff_A_WwWJaJPh2_0),.din(w_dff_A_nsDddu9i0_0),.clk(gclk));
	jdff dff_A_WwWJaJPh2_0(.dout(w_dff_A_H7AXLq781_0),.din(w_dff_A_WwWJaJPh2_0),.clk(gclk));
	jdff dff_A_H7AXLq781_0(.dout(w_dff_A_GGInvWlw1_0),.din(w_dff_A_H7AXLq781_0),.clk(gclk));
	jdff dff_A_GGInvWlw1_0(.dout(w_dff_A_mPbDdSW04_0),.din(w_dff_A_GGInvWlw1_0),.clk(gclk));
	jdff dff_A_mPbDdSW04_0(.dout(w_dff_A_mAjVKfb88_0),.din(w_dff_A_mPbDdSW04_0),.clk(gclk));
	jdff dff_A_mAjVKfb88_0(.dout(w_dff_A_JxsdCr5v8_0),.din(w_dff_A_mAjVKfb88_0),.clk(gclk));
	jdff dff_A_JxsdCr5v8_0(.dout(w_dff_A_mG9LsSU07_0),.din(w_dff_A_JxsdCr5v8_0),.clk(gclk));
	jdff dff_A_mG9LsSU07_0(.dout(w_dff_A_ceylxuyL0_0),.din(w_dff_A_mG9LsSU07_0),.clk(gclk));
	jdff dff_A_ceylxuyL0_0(.dout(w_dff_A_Qw3y8sc13_0),.din(w_dff_A_ceylxuyL0_0),.clk(gclk));
	jdff dff_A_Qw3y8sc13_0(.dout(w_dff_A_H7WRDg3Q7_0),.din(w_dff_A_Qw3y8sc13_0),.clk(gclk));
	jdff dff_A_H7WRDg3Q7_0(.dout(w_dff_A_Rfx2JrZF2_0),.din(w_dff_A_H7WRDg3Q7_0),.clk(gclk));
	jdff dff_A_Rfx2JrZF2_0(.dout(w_dff_A_0CYqhtmb9_0),.din(w_dff_A_Rfx2JrZF2_0),.clk(gclk));
	jdff dff_A_0CYqhtmb9_0(.dout(w_dff_A_FsE5HE270_0),.din(w_dff_A_0CYqhtmb9_0),.clk(gclk));
	jdff dff_A_FsE5HE270_0(.dout(w_dff_A_M1KVHirV2_0),.din(w_dff_A_FsE5HE270_0),.clk(gclk));
	jdff dff_A_M1KVHirV2_0(.dout(w_dff_A_aZo1DHpL7_0),.din(w_dff_A_M1KVHirV2_0),.clk(gclk));
	jdff dff_A_aZo1DHpL7_0(.dout(G673),.din(w_dff_A_aZo1DHpL7_0),.clk(gclk));
	jdff dff_A_0GmzN7ei2_2(.dout(w_dff_A_duon9KZm0_0),.din(w_dff_A_0GmzN7ei2_2),.clk(gclk));
	jdff dff_A_duon9KZm0_0(.dout(w_dff_A_zAKwyIc84_0),.din(w_dff_A_duon9KZm0_0),.clk(gclk));
	jdff dff_A_zAKwyIc84_0(.dout(w_dff_A_mBPgKd0S5_0),.din(w_dff_A_zAKwyIc84_0),.clk(gclk));
	jdff dff_A_mBPgKd0S5_0(.dout(w_dff_A_SLtzBcl09_0),.din(w_dff_A_mBPgKd0S5_0),.clk(gclk));
	jdff dff_A_SLtzBcl09_0(.dout(w_dff_A_ekZ0o5Kc1_0),.din(w_dff_A_SLtzBcl09_0),.clk(gclk));
	jdff dff_A_ekZ0o5Kc1_0(.dout(w_dff_A_tjAcEdqW8_0),.din(w_dff_A_ekZ0o5Kc1_0),.clk(gclk));
	jdff dff_A_tjAcEdqW8_0(.dout(w_dff_A_R6i15A043_0),.din(w_dff_A_tjAcEdqW8_0),.clk(gclk));
	jdff dff_A_R6i15A043_0(.dout(w_dff_A_UUGW9Jqa0_0),.din(w_dff_A_R6i15A043_0),.clk(gclk));
	jdff dff_A_UUGW9Jqa0_0(.dout(w_dff_A_VNKoP4VG1_0),.din(w_dff_A_UUGW9Jqa0_0),.clk(gclk));
	jdff dff_A_VNKoP4VG1_0(.dout(w_dff_A_6kqBOXer0_0),.din(w_dff_A_VNKoP4VG1_0),.clk(gclk));
	jdff dff_A_6kqBOXer0_0(.dout(w_dff_A_kH2wlUKi1_0),.din(w_dff_A_6kqBOXer0_0),.clk(gclk));
	jdff dff_A_kH2wlUKi1_0(.dout(w_dff_A_LbLNEQLS3_0),.din(w_dff_A_kH2wlUKi1_0),.clk(gclk));
	jdff dff_A_LbLNEQLS3_0(.dout(w_dff_A_10js08Js5_0),.din(w_dff_A_LbLNEQLS3_0),.clk(gclk));
	jdff dff_A_10js08Js5_0(.dout(w_dff_A_eeOB5FER8_0),.din(w_dff_A_10js08Js5_0),.clk(gclk));
	jdff dff_A_eeOB5FER8_0(.dout(w_dff_A_NyySJDko3_0),.din(w_dff_A_eeOB5FER8_0),.clk(gclk));
	jdff dff_A_NyySJDko3_0(.dout(w_dff_A_6JavPM1P1_0),.din(w_dff_A_NyySJDko3_0),.clk(gclk));
	jdff dff_A_6JavPM1P1_0(.dout(w_dff_A_A89uGD5j2_0),.din(w_dff_A_6JavPM1P1_0),.clk(gclk));
	jdff dff_A_A89uGD5j2_0(.dout(w_dff_A_TU3vFcyh3_0),.din(w_dff_A_A89uGD5j2_0),.clk(gclk));
	jdff dff_A_TU3vFcyh3_0(.dout(w_dff_A_ck8ovaT59_0),.din(w_dff_A_TU3vFcyh3_0),.clk(gclk));
	jdff dff_A_ck8ovaT59_0(.dout(w_dff_A_VTUk3OHL6_0),.din(w_dff_A_ck8ovaT59_0),.clk(gclk));
	jdff dff_A_VTUk3OHL6_0(.dout(G707),.din(w_dff_A_VTUk3OHL6_0),.clk(gclk));
	jdff dff_A_0tDgTm6S3_2(.dout(w_dff_A_jzhstoLj0_0),.din(w_dff_A_0tDgTm6S3_2),.clk(gclk));
	jdff dff_A_jzhstoLj0_0(.dout(w_dff_A_nUx6zhfL5_0),.din(w_dff_A_jzhstoLj0_0),.clk(gclk));
	jdff dff_A_nUx6zhfL5_0(.dout(w_dff_A_XjufneCv9_0),.din(w_dff_A_nUx6zhfL5_0),.clk(gclk));
	jdff dff_A_XjufneCv9_0(.dout(w_dff_A_UvBoPF852_0),.din(w_dff_A_XjufneCv9_0),.clk(gclk));
	jdff dff_A_UvBoPF852_0(.dout(w_dff_A_hjuMrogZ7_0),.din(w_dff_A_UvBoPF852_0),.clk(gclk));
	jdff dff_A_hjuMrogZ7_0(.dout(w_dff_A_R8kemgtX8_0),.din(w_dff_A_hjuMrogZ7_0),.clk(gclk));
	jdff dff_A_R8kemgtX8_0(.dout(w_dff_A_r3H9kFdA5_0),.din(w_dff_A_R8kemgtX8_0),.clk(gclk));
	jdff dff_A_r3H9kFdA5_0(.dout(w_dff_A_6DdDNP5z0_0),.din(w_dff_A_r3H9kFdA5_0),.clk(gclk));
	jdff dff_A_6DdDNP5z0_0(.dout(w_dff_A_8vrG5R2g8_0),.din(w_dff_A_6DdDNP5z0_0),.clk(gclk));
	jdff dff_A_8vrG5R2g8_0(.dout(w_dff_A_gs3auYyT9_0),.din(w_dff_A_8vrG5R2g8_0),.clk(gclk));
	jdff dff_A_gs3auYyT9_0(.dout(w_dff_A_GakBwCVH6_0),.din(w_dff_A_gs3auYyT9_0),.clk(gclk));
	jdff dff_A_GakBwCVH6_0(.dout(w_dff_A_qo3XzztQ9_0),.din(w_dff_A_GakBwCVH6_0),.clk(gclk));
	jdff dff_A_qo3XzztQ9_0(.dout(w_dff_A_YLapVxBp0_0),.din(w_dff_A_qo3XzztQ9_0),.clk(gclk));
	jdff dff_A_YLapVxBp0_0(.dout(w_dff_A_lSmte0YH2_0),.din(w_dff_A_YLapVxBp0_0),.clk(gclk));
	jdff dff_A_lSmte0YH2_0(.dout(w_dff_A_tQ2AxIQU9_0),.din(w_dff_A_lSmte0YH2_0),.clk(gclk));
	jdff dff_A_tQ2AxIQU9_0(.dout(w_dff_A_OP2lL9df7_0),.din(w_dff_A_tQ2AxIQU9_0),.clk(gclk));
	jdff dff_A_OP2lL9df7_0(.dout(w_dff_A_ZwzSGMdN1_0),.din(w_dff_A_OP2lL9df7_0),.clk(gclk));
	jdff dff_A_ZwzSGMdN1_0(.dout(w_dff_A_YZcJYF1H1_0),.din(w_dff_A_ZwzSGMdN1_0),.clk(gclk));
	jdff dff_A_YZcJYF1H1_0(.dout(w_dff_A_q4ijwy397_0),.din(w_dff_A_YZcJYF1H1_0),.clk(gclk));
	jdff dff_A_q4ijwy397_0(.dout(w_dff_A_WmIreB3a9_0),.din(w_dff_A_q4ijwy397_0),.clk(gclk));
	jdff dff_A_WmIreB3a9_0(.dout(G715),.din(w_dff_A_WmIreB3a9_0),.clk(gclk));
	jdff dff_A_MDA1CyFJ0_2(.dout(w_dff_A_lOytSnZh2_0),.din(w_dff_A_MDA1CyFJ0_2),.clk(gclk));
	jdff dff_A_lOytSnZh2_0(.dout(w_dff_A_Vwr0DdND6_0),.din(w_dff_A_lOytSnZh2_0),.clk(gclk));
	jdff dff_A_Vwr0DdND6_0(.dout(w_dff_A_EcwGGLiT4_0),.din(w_dff_A_Vwr0DdND6_0),.clk(gclk));
	jdff dff_A_EcwGGLiT4_0(.dout(w_dff_A_kEeA7pO89_0),.din(w_dff_A_EcwGGLiT4_0),.clk(gclk));
	jdff dff_A_kEeA7pO89_0(.dout(w_dff_A_EjAI1DBK7_0),.din(w_dff_A_kEeA7pO89_0),.clk(gclk));
	jdff dff_A_EjAI1DBK7_0(.dout(w_dff_A_080ubyZE2_0),.din(w_dff_A_EjAI1DBK7_0),.clk(gclk));
	jdff dff_A_080ubyZE2_0(.dout(w_dff_A_ZJmhIdV58_0),.din(w_dff_A_080ubyZE2_0),.clk(gclk));
	jdff dff_A_ZJmhIdV58_0(.dout(w_dff_A_rKaC1NUK0_0),.din(w_dff_A_ZJmhIdV58_0),.clk(gclk));
	jdff dff_A_rKaC1NUK0_0(.dout(w_dff_A_l4kRRui19_0),.din(w_dff_A_rKaC1NUK0_0),.clk(gclk));
	jdff dff_A_l4kRRui19_0(.dout(w_dff_A_KrnvwBLl7_0),.din(w_dff_A_l4kRRui19_0),.clk(gclk));
	jdff dff_A_KrnvwBLl7_0(.dout(w_dff_A_ag3fLpp56_0),.din(w_dff_A_KrnvwBLl7_0),.clk(gclk));
	jdff dff_A_ag3fLpp56_0(.dout(w_dff_A_Ax5Uy56q6_0),.din(w_dff_A_ag3fLpp56_0),.clk(gclk));
	jdff dff_A_Ax5Uy56q6_0(.dout(w_dff_A_Hv0zqIUP4_0),.din(w_dff_A_Ax5Uy56q6_0),.clk(gclk));
	jdff dff_A_Hv0zqIUP4_0(.dout(w_dff_A_YOg9rkaN6_0),.din(w_dff_A_Hv0zqIUP4_0),.clk(gclk));
	jdff dff_A_YOg9rkaN6_0(.dout(w_dff_A_nPJjfh300_0),.din(w_dff_A_YOg9rkaN6_0),.clk(gclk));
	jdff dff_A_nPJjfh300_0(.dout(w_dff_A_1XsTjUlC5_0),.din(w_dff_A_nPJjfh300_0),.clk(gclk));
	jdff dff_A_1XsTjUlC5_0(.dout(G598),.din(w_dff_A_1XsTjUlC5_0),.clk(gclk));
	jdff dff_A_JI54GYgt8_2(.dout(w_dff_A_w0BV9Hwn9_0),.din(w_dff_A_JI54GYgt8_2),.clk(gclk));
	jdff dff_A_w0BV9Hwn9_0(.dout(w_dff_A_JRxSQKDk0_0),.din(w_dff_A_w0BV9Hwn9_0),.clk(gclk));
	jdff dff_A_JRxSQKDk0_0(.dout(w_dff_A_eh6D1e7U1_0),.din(w_dff_A_JRxSQKDk0_0),.clk(gclk));
	jdff dff_A_eh6D1e7U1_0(.dout(w_dff_A_BTHJQcXM5_0),.din(w_dff_A_eh6D1e7U1_0),.clk(gclk));
	jdff dff_A_BTHJQcXM5_0(.dout(w_dff_A_cDVLQgpE8_0),.din(w_dff_A_BTHJQcXM5_0),.clk(gclk));
	jdff dff_A_cDVLQgpE8_0(.dout(w_dff_A_sbTycoJG4_0),.din(w_dff_A_cDVLQgpE8_0),.clk(gclk));
	jdff dff_A_sbTycoJG4_0(.dout(w_dff_A_jQYkZMLj8_0),.din(w_dff_A_sbTycoJG4_0),.clk(gclk));
	jdff dff_A_jQYkZMLj8_0(.dout(w_dff_A_6FLfHyDC3_0),.din(w_dff_A_jQYkZMLj8_0),.clk(gclk));
	jdff dff_A_6FLfHyDC3_0(.dout(w_dff_A_1M0IZtja1_0),.din(w_dff_A_6FLfHyDC3_0),.clk(gclk));
	jdff dff_A_1M0IZtja1_0(.dout(w_dff_A_XiVTC9CX2_0),.din(w_dff_A_1M0IZtja1_0),.clk(gclk));
	jdff dff_A_XiVTC9CX2_0(.dout(w_dff_A_khFTa7cK8_0),.din(w_dff_A_XiVTC9CX2_0),.clk(gclk));
	jdff dff_A_khFTa7cK8_0(.dout(w_dff_A_gfIZ3ys35_0),.din(w_dff_A_khFTa7cK8_0),.clk(gclk));
	jdff dff_A_gfIZ3ys35_0(.dout(w_dff_A_5o39kAha7_0),.din(w_dff_A_gfIZ3ys35_0),.clk(gclk));
	jdff dff_A_5o39kAha7_0(.dout(w_dff_A_SM6zpNTd5_0),.din(w_dff_A_5o39kAha7_0),.clk(gclk));
	jdff dff_A_SM6zpNTd5_0(.dout(w_dff_A_8Uh82O9k9_0),.din(w_dff_A_SM6zpNTd5_0),.clk(gclk));
	jdff dff_A_8Uh82O9k9_0(.dout(w_dff_A_vhiEA8VD0_0),.din(w_dff_A_8Uh82O9k9_0),.clk(gclk));
	jdff dff_A_vhiEA8VD0_0(.dout(G610),.din(w_dff_A_vhiEA8VD0_0),.clk(gclk));
	jdff dff_A_QgbmpZht9_2(.dout(w_dff_A_GMILkGLM9_0),.din(w_dff_A_QgbmpZht9_2),.clk(gclk));
	jdff dff_A_GMILkGLM9_0(.dout(w_dff_A_VlpjscMX6_0),.din(w_dff_A_GMILkGLM9_0),.clk(gclk));
	jdff dff_A_VlpjscMX6_0(.dout(w_dff_A_yKboFWFA5_0),.din(w_dff_A_VlpjscMX6_0),.clk(gclk));
	jdff dff_A_yKboFWFA5_0(.dout(w_dff_A_KX9Tqpgr0_0),.din(w_dff_A_yKboFWFA5_0),.clk(gclk));
	jdff dff_A_KX9Tqpgr0_0(.dout(w_dff_A_NsyMePNK7_0),.din(w_dff_A_KX9Tqpgr0_0),.clk(gclk));
	jdff dff_A_NsyMePNK7_0(.dout(w_dff_A_VjAGNj3F7_0),.din(w_dff_A_NsyMePNK7_0),.clk(gclk));
	jdff dff_A_VjAGNj3F7_0(.dout(w_dff_A_moX6JpjN0_0),.din(w_dff_A_VjAGNj3F7_0),.clk(gclk));
	jdff dff_A_moX6JpjN0_0(.dout(w_dff_A_Lr7p19I87_0),.din(w_dff_A_moX6JpjN0_0),.clk(gclk));
	jdff dff_A_Lr7p19I87_0(.dout(w_dff_A_mL4SnxAD9_0),.din(w_dff_A_Lr7p19I87_0),.clk(gclk));
	jdff dff_A_mL4SnxAD9_0(.dout(w_dff_A_wDWFw27g5_0),.din(w_dff_A_mL4SnxAD9_0),.clk(gclk));
	jdff dff_A_wDWFw27g5_0(.dout(w_dff_A_HmxKfANZ3_0),.din(w_dff_A_wDWFw27g5_0),.clk(gclk));
	jdff dff_A_HmxKfANZ3_0(.dout(w_dff_A_mz0dJCbt9_0),.din(w_dff_A_HmxKfANZ3_0),.clk(gclk));
	jdff dff_A_mz0dJCbt9_0(.dout(w_dff_A_GULorWJ72_0),.din(w_dff_A_mz0dJCbt9_0),.clk(gclk));
	jdff dff_A_GULorWJ72_0(.dout(w_dff_A_iQdzLS0R2_0),.din(w_dff_A_GULorWJ72_0),.clk(gclk));
	jdff dff_A_iQdzLS0R2_0(.dout(G588),.din(w_dff_A_iQdzLS0R2_0),.clk(gclk));
	jdff dff_A_0OgvtRqK7_2(.dout(w_dff_A_cSb0UA0b2_0),.din(w_dff_A_0OgvtRqK7_2),.clk(gclk));
	jdff dff_A_cSb0UA0b2_0(.dout(w_dff_A_XcHrV9VL9_0),.din(w_dff_A_cSb0UA0b2_0),.clk(gclk));
	jdff dff_A_XcHrV9VL9_0(.dout(w_dff_A_4jSMUs2g9_0),.din(w_dff_A_XcHrV9VL9_0),.clk(gclk));
	jdff dff_A_4jSMUs2g9_0(.dout(w_dff_A_oUSY9uU15_0),.din(w_dff_A_4jSMUs2g9_0),.clk(gclk));
	jdff dff_A_oUSY9uU15_0(.dout(w_dff_A_Vaw4VKmV6_0),.din(w_dff_A_oUSY9uU15_0),.clk(gclk));
	jdff dff_A_Vaw4VKmV6_0(.dout(w_dff_A_juh1xyHG3_0),.din(w_dff_A_Vaw4VKmV6_0),.clk(gclk));
	jdff dff_A_juh1xyHG3_0(.dout(w_dff_A_Q0wTUQkw1_0),.din(w_dff_A_juh1xyHG3_0),.clk(gclk));
	jdff dff_A_Q0wTUQkw1_0(.dout(w_dff_A_kbJX1bYZ4_0),.din(w_dff_A_Q0wTUQkw1_0),.clk(gclk));
	jdff dff_A_kbJX1bYZ4_0(.dout(w_dff_A_H7nS2ORk9_0),.din(w_dff_A_kbJX1bYZ4_0),.clk(gclk));
	jdff dff_A_H7nS2ORk9_0(.dout(w_dff_A_1zcunMHv4_0),.din(w_dff_A_H7nS2ORk9_0),.clk(gclk));
	jdff dff_A_1zcunMHv4_0(.dout(w_dff_A_6EvOP3fu0_0),.din(w_dff_A_1zcunMHv4_0),.clk(gclk));
	jdff dff_A_6EvOP3fu0_0(.dout(w_dff_A_wqiLaPqg7_0),.din(w_dff_A_6EvOP3fu0_0),.clk(gclk));
	jdff dff_A_wqiLaPqg7_0(.dout(w_dff_A_yzKXFTsU4_0),.din(w_dff_A_wqiLaPqg7_0),.clk(gclk));
	jdff dff_A_yzKXFTsU4_0(.dout(w_dff_A_OpiAFAgk7_0),.din(w_dff_A_yzKXFTsU4_0),.clk(gclk));
	jdff dff_A_OpiAFAgk7_0(.dout(w_dff_A_8yGStRn20_0),.din(w_dff_A_OpiAFAgk7_0),.clk(gclk));
	jdff dff_A_8yGStRn20_0(.dout(w_dff_A_RaNgJZ0x9_0),.din(w_dff_A_8yGStRn20_0),.clk(gclk));
	jdff dff_A_RaNgJZ0x9_0(.dout(G615),.din(w_dff_A_RaNgJZ0x9_0),.clk(gclk));
	jdff dff_A_WZtzsak76_2(.dout(w_dff_A_cT7U8lKk6_0),.din(w_dff_A_WZtzsak76_2),.clk(gclk));
	jdff dff_A_cT7U8lKk6_0(.dout(w_dff_A_suS6PqyK1_0),.din(w_dff_A_cT7U8lKk6_0),.clk(gclk));
	jdff dff_A_suS6PqyK1_0(.dout(w_dff_A_PInrur1m3_0),.din(w_dff_A_suS6PqyK1_0),.clk(gclk));
	jdff dff_A_PInrur1m3_0(.dout(w_dff_A_neArHU5K6_0),.din(w_dff_A_PInrur1m3_0),.clk(gclk));
	jdff dff_A_neArHU5K6_0(.dout(w_dff_A_50ZKOalW7_0),.din(w_dff_A_neArHU5K6_0),.clk(gclk));
	jdff dff_A_50ZKOalW7_0(.dout(w_dff_A_27h0MhW31_0),.din(w_dff_A_50ZKOalW7_0),.clk(gclk));
	jdff dff_A_27h0MhW31_0(.dout(w_dff_A_kMTM2Ou99_0),.din(w_dff_A_27h0MhW31_0),.clk(gclk));
	jdff dff_A_kMTM2Ou99_0(.dout(w_dff_A_bJc3GcsB8_0),.din(w_dff_A_kMTM2Ou99_0),.clk(gclk));
	jdff dff_A_bJc3GcsB8_0(.dout(w_dff_A_jm0biYLj5_0),.din(w_dff_A_bJc3GcsB8_0),.clk(gclk));
	jdff dff_A_jm0biYLj5_0(.dout(w_dff_A_JytWYUNK9_0),.din(w_dff_A_jm0biYLj5_0),.clk(gclk));
	jdff dff_A_JytWYUNK9_0(.dout(w_dff_A_Z2F8HuOt0_0),.din(w_dff_A_JytWYUNK9_0),.clk(gclk));
	jdff dff_A_Z2F8HuOt0_0(.dout(w_dff_A_WNgr8LQn6_0),.din(w_dff_A_Z2F8HuOt0_0),.clk(gclk));
	jdff dff_A_WNgr8LQn6_0(.dout(w_dff_A_os8tY1mZ1_0),.din(w_dff_A_WNgr8LQn6_0),.clk(gclk));
	jdff dff_A_os8tY1mZ1_0(.dout(w_dff_A_jZmj1A6T9_0),.din(w_dff_A_os8tY1mZ1_0),.clk(gclk));
	jdff dff_A_jZmj1A6T9_0(.dout(w_dff_A_x1YibhHq6_0),.din(w_dff_A_jZmj1A6T9_0),.clk(gclk));
	jdff dff_A_x1YibhHq6_0(.dout(w_dff_A_eLgRMScw4_0),.din(w_dff_A_x1YibhHq6_0),.clk(gclk));
	jdff dff_A_eLgRMScw4_0(.dout(G626),.din(w_dff_A_eLgRMScw4_0),.clk(gclk));
	jdff dff_A_aqgWgVCw7_2(.dout(w_dff_A_O1rFA57x9_0),.din(w_dff_A_aqgWgVCw7_2),.clk(gclk));
	jdff dff_A_O1rFA57x9_0(.dout(w_dff_A_7PQ4g2Kp1_0),.din(w_dff_A_O1rFA57x9_0),.clk(gclk));
	jdff dff_A_7PQ4g2Kp1_0(.dout(w_dff_A_9Qe5Fee53_0),.din(w_dff_A_7PQ4g2Kp1_0),.clk(gclk));
	jdff dff_A_9Qe5Fee53_0(.dout(w_dff_A_4ToV2gLw2_0),.din(w_dff_A_9Qe5Fee53_0),.clk(gclk));
	jdff dff_A_4ToV2gLw2_0(.dout(w_dff_A_VfvOAFy55_0),.din(w_dff_A_4ToV2gLw2_0),.clk(gclk));
	jdff dff_A_VfvOAFy55_0(.dout(w_dff_A_XbPDiyvr6_0),.din(w_dff_A_VfvOAFy55_0),.clk(gclk));
	jdff dff_A_XbPDiyvr6_0(.dout(w_dff_A_MC29mWjU4_0),.din(w_dff_A_XbPDiyvr6_0),.clk(gclk));
	jdff dff_A_MC29mWjU4_0(.dout(w_dff_A_h5ic0Zw61_0),.din(w_dff_A_MC29mWjU4_0),.clk(gclk));
	jdff dff_A_h5ic0Zw61_0(.dout(w_dff_A_Lav6XARH1_0),.din(w_dff_A_h5ic0Zw61_0),.clk(gclk));
	jdff dff_A_Lav6XARH1_0(.dout(w_dff_A_YHyRqu6v2_0),.din(w_dff_A_Lav6XARH1_0),.clk(gclk));
	jdff dff_A_YHyRqu6v2_0(.dout(w_dff_A_E98IyfpV3_0),.din(w_dff_A_YHyRqu6v2_0),.clk(gclk));
	jdff dff_A_E98IyfpV3_0(.dout(w_dff_A_HzqF36XT4_0),.din(w_dff_A_E98IyfpV3_0),.clk(gclk));
	jdff dff_A_HzqF36XT4_0(.dout(w_dff_A_XZoiT8XU2_0),.din(w_dff_A_HzqF36XT4_0),.clk(gclk));
	jdff dff_A_XZoiT8XU2_0(.dout(w_dff_A_Z16LTNoq6_0),.din(w_dff_A_XZoiT8XU2_0),.clk(gclk));
	jdff dff_A_Z16LTNoq6_0(.dout(G632),.din(w_dff_A_Z16LTNoq6_0),.clk(gclk));
	jdff dff_A_ExzIBIS38_1(.dout(w_dff_A_dtNI1rGH3_0),.din(w_dff_A_ExzIBIS38_1),.clk(gclk));
	jdff dff_A_dtNI1rGH3_0(.dout(w_dff_A_FNDp067N1_0),.din(w_dff_A_dtNI1rGH3_0),.clk(gclk));
	jdff dff_A_FNDp067N1_0(.dout(w_dff_A_xV7j1vtZ2_0),.din(w_dff_A_FNDp067N1_0),.clk(gclk));
	jdff dff_A_xV7j1vtZ2_0(.dout(w_dff_A_Mbdo1fJG4_0),.din(w_dff_A_xV7j1vtZ2_0),.clk(gclk));
	jdff dff_A_Mbdo1fJG4_0(.dout(w_dff_A_FwPVKu9g9_0),.din(w_dff_A_Mbdo1fJG4_0),.clk(gclk));
	jdff dff_A_FwPVKu9g9_0(.dout(w_dff_A_vV9WBLU51_0),.din(w_dff_A_FwPVKu9g9_0),.clk(gclk));
	jdff dff_A_vV9WBLU51_0(.dout(w_dff_A_7IbmsY3R9_0),.din(w_dff_A_vV9WBLU51_0),.clk(gclk));
	jdff dff_A_7IbmsY3R9_0(.dout(w_dff_A_3TYXNsXY0_0),.din(w_dff_A_7IbmsY3R9_0),.clk(gclk));
	jdff dff_A_3TYXNsXY0_0(.dout(w_dff_A_1wyZqhUV3_0),.din(w_dff_A_3TYXNsXY0_0),.clk(gclk));
	jdff dff_A_1wyZqhUV3_0(.dout(w_dff_A_4w8sKzXo0_0),.din(w_dff_A_1wyZqhUV3_0),.clk(gclk));
	jdff dff_A_4w8sKzXo0_0(.dout(w_dff_A_NJ3Sotag4_0),.din(w_dff_A_4w8sKzXo0_0),.clk(gclk));
	jdff dff_A_NJ3Sotag4_0(.dout(w_dff_A_DbYTJV8b8_0),.din(w_dff_A_NJ3Sotag4_0),.clk(gclk));
	jdff dff_A_DbYTJV8b8_0(.dout(w_dff_A_hQ1JA2t21_0),.din(w_dff_A_DbYTJV8b8_0),.clk(gclk));
	jdff dff_A_hQ1JA2t21_0(.dout(w_dff_A_1ur4pzOk2_0),.din(w_dff_A_hQ1JA2t21_0),.clk(gclk));
	jdff dff_A_1ur4pzOk2_0(.dout(w_dff_A_R0NBYpVr0_0),.din(w_dff_A_1ur4pzOk2_0),.clk(gclk));
	jdff dff_A_R0NBYpVr0_0(.dout(w_dff_A_hmiUOb7Z4_0),.din(w_dff_A_R0NBYpVr0_0),.clk(gclk));
	jdff dff_A_hmiUOb7Z4_0(.dout(w_dff_A_ow0Cb9UT8_0),.din(w_dff_A_hmiUOb7Z4_0),.clk(gclk));
	jdff dff_A_ow0Cb9UT8_0(.dout(w_dff_A_cvczcfHv9_0),.din(w_dff_A_ow0Cb9UT8_0),.clk(gclk));
	jdff dff_A_cvczcfHv9_0(.dout(w_dff_A_m0IDceCV9_0),.din(w_dff_A_cvczcfHv9_0),.clk(gclk));
	jdff dff_A_m0IDceCV9_0(.dout(w_dff_A_sinQH8b84_0),.din(w_dff_A_m0IDceCV9_0),.clk(gclk));
	jdff dff_A_sinQH8b84_0(.dout(G1002),.din(w_dff_A_sinQH8b84_0),.clk(gclk));
	jdff dff_A_eF25cZUD2_1(.dout(w_dff_A_NT17urFK9_0),.din(w_dff_A_eF25cZUD2_1),.clk(gclk));
	jdff dff_A_NT17urFK9_0(.dout(w_dff_A_IxLx04z91_0),.din(w_dff_A_NT17urFK9_0),.clk(gclk));
	jdff dff_A_IxLx04z91_0(.dout(w_dff_A_5wUPmnbG6_0),.din(w_dff_A_IxLx04z91_0),.clk(gclk));
	jdff dff_A_5wUPmnbG6_0(.dout(w_dff_A_icRxBarg5_0),.din(w_dff_A_5wUPmnbG6_0),.clk(gclk));
	jdff dff_A_icRxBarg5_0(.dout(w_dff_A_Mam7M0j77_0),.din(w_dff_A_icRxBarg5_0),.clk(gclk));
	jdff dff_A_Mam7M0j77_0(.dout(w_dff_A_qRNFJs2l4_0),.din(w_dff_A_Mam7M0j77_0),.clk(gclk));
	jdff dff_A_qRNFJs2l4_0(.dout(w_dff_A_2UFy3Wgo0_0),.din(w_dff_A_qRNFJs2l4_0),.clk(gclk));
	jdff dff_A_2UFy3Wgo0_0(.dout(w_dff_A_KpDxxA5a9_0),.din(w_dff_A_2UFy3Wgo0_0),.clk(gclk));
	jdff dff_A_KpDxxA5a9_0(.dout(w_dff_A_RmcJZGW83_0),.din(w_dff_A_KpDxxA5a9_0),.clk(gclk));
	jdff dff_A_RmcJZGW83_0(.dout(w_dff_A_l1OlhjxF7_0),.din(w_dff_A_RmcJZGW83_0),.clk(gclk));
	jdff dff_A_l1OlhjxF7_0(.dout(w_dff_A_2zAfa6a85_0),.din(w_dff_A_l1OlhjxF7_0),.clk(gclk));
	jdff dff_A_2zAfa6a85_0(.dout(w_dff_A_B4Pxk3qv3_0),.din(w_dff_A_2zAfa6a85_0),.clk(gclk));
	jdff dff_A_B4Pxk3qv3_0(.dout(w_dff_A_j1qw7Aax9_0),.din(w_dff_A_B4Pxk3qv3_0),.clk(gclk));
	jdff dff_A_j1qw7Aax9_0(.dout(w_dff_A_ZL6gaiFr9_0),.din(w_dff_A_j1qw7Aax9_0),.clk(gclk));
	jdff dff_A_ZL6gaiFr9_0(.dout(w_dff_A_zAWVk2s33_0),.din(w_dff_A_ZL6gaiFr9_0),.clk(gclk));
	jdff dff_A_zAWVk2s33_0(.dout(w_dff_A_Yw9bDhUO8_0),.din(w_dff_A_zAWVk2s33_0),.clk(gclk));
	jdff dff_A_Yw9bDhUO8_0(.dout(w_dff_A_Zi4ClYjW8_0),.din(w_dff_A_Yw9bDhUO8_0),.clk(gclk));
	jdff dff_A_Zi4ClYjW8_0(.dout(w_dff_A_aIZ3bLTn5_0),.din(w_dff_A_Zi4ClYjW8_0),.clk(gclk));
	jdff dff_A_aIZ3bLTn5_0(.dout(w_dff_A_tv8cw3Th2_0),.din(w_dff_A_aIZ3bLTn5_0),.clk(gclk));
	jdff dff_A_tv8cw3Th2_0(.dout(w_dff_A_Tz0ymolQ7_0),.din(w_dff_A_tv8cw3Th2_0),.clk(gclk));
	jdff dff_A_Tz0ymolQ7_0(.dout(G1004),.din(w_dff_A_Tz0ymolQ7_0),.clk(gclk));
	jdff dff_A_mfoVLXEC9_2(.dout(w_dff_A_agD0E8LR5_0),.din(w_dff_A_mfoVLXEC9_2),.clk(gclk));
	jdff dff_A_agD0E8LR5_0(.dout(w_dff_A_eEYs9Fey2_0),.din(w_dff_A_agD0E8LR5_0),.clk(gclk));
	jdff dff_A_eEYs9Fey2_0(.dout(w_dff_A_4gBT5zXA3_0),.din(w_dff_A_eEYs9Fey2_0),.clk(gclk));
	jdff dff_A_4gBT5zXA3_0(.dout(w_dff_A_EP4GlbTC9_0),.din(w_dff_A_4gBT5zXA3_0),.clk(gclk));
	jdff dff_A_EP4GlbTC9_0(.dout(w_dff_A_eBdOUDx58_0),.din(w_dff_A_EP4GlbTC9_0),.clk(gclk));
	jdff dff_A_eBdOUDx58_0(.dout(w_dff_A_bgH74ekf0_0),.din(w_dff_A_eBdOUDx58_0),.clk(gclk));
	jdff dff_A_bgH74ekf0_0(.dout(w_dff_A_T5NmPRPy0_0),.din(w_dff_A_bgH74ekf0_0),.clk(gclk));
	jdff dff_A_T5NmPRPy0_0(.dout(w_dff_A_oMBoHOQK8_0),.din(w_dff_A_T5NmPRPy0_0),.clk(gclk));
	jdff dff_A_oMBoHOQK8_0(.dout(w_dff_A_BzwpgGgq8_0),.din(w_dff_A_oMBoHOQK8_0),.clk(gclk));
	jdff dff_A_BzwpgGgq8_0(.dout(w_dff_A_PjLHKwBi4_0),.din(w_dff_A_BzwpgGgq8_0),.clk(gclk));
	jdff dff_A_PjLHKwBi4_0(.dout(w_dff_A_PXBX8FA26_0),.din(w_dff_A_PjLHKwBi4_0),.clk(gclk));
	jdff dff_A_PXBX8FA26_0(.dout(G591),.din(w_dff_A_PXBX8FA26_0),.clk(gclk));
	jdff dff_A_qJmjJP2c4_2(.dout(w_dff_A_qXRAtiND2_0),.din(w_dff_A_qJmjJP2c4_2),.clk(gclk));
	jdff dff_A_qXRAtiND2_0(.dout(w_dff_A_Jbk10W3U2_0),.din(w_dff_A_qXRAtiND2_0),.clk(gclk));
	jdff dff_A_Jbk10W3U2_0(.dout(w_dff_A_RHWDoGBm5_0),.din(w_dff_A_Jbk10W3U2_0),.clk(gclk));
	jdff dff_A_RHWDoGBm5_0(.dout(w_dff_A_2mJQbMZB9_0),.din(w_dff_A_RHWDoGBm5_0),.clk(gclk));
	jdff dff_A_2mJQbMZB9_0(.dout(w_dff_A_fyVjTgFU0_0),.din(w_dff_A_2mJQbMZB9_0),.clk(gclk));
	jdff dff_A_fyVjTgFU0_0(.dout(w_dff_A_kIpIJOjR6_0),.din(w_dff_A_fyVjTgFU0_0),.clk(gclk));
	jdff dff_A_kIpIJOjR6_0(.dout(w_dff_A_jyJCDh204_0),.din(w_dff_A_kIpIJOjR6_0),.clk(gclk));
	jdff dff_A_jyJCDh204_0(.dout(w_dff_A_aM6fNRj28_0),.din(w_dff_A_jyJCDh204_0),.clk(gclk));
	jdff dff_A_aM6fNRj28_0(.dout(w_dff_A_v4gygKSV0_0),.din(w_dff_A_aM6fNRj28_0),.clk(gclk));
	jdff dff_A_v4gygKSV0_0(.dout(w_dff_A_KTkZyOXT9_0),.din(w_dff_A_v4gygKSV0_0),.clk(gclk));
	jdff dff_A_KTkZyOXT9_0(.dout(w_dff_A_k4ucQ4pX3_0),.din(w_dff_A_KTkZyOXT9_0),.clk(gclk));
	jdff dff_A_k4ucQ4pX3_0(.dout(G618),.din(w_dff_A_k4ucQ4pX3_0),.clk(gclk));
	jdff dff_A_yfLRIfqS6_2(.dout(w_dff_A_1xgzYpP76_0),.din(w_dff_A_yfLRIfqS6_2),.clk(gclk));
	jdff dff_A_1xgzYpP76_0(.dout(w_dff_A_zPAqavb28_0),.din(w_dff_A_1xgzYpP76_0),.clk(gclk));
	jdff dff_A_zPAqavb28_0(.dout(w_dff_A_FNI2N5oB0_0),.din(w_dff_A_zPAqavb28_0),.clk(gclk));
	jdff dff_A_FNI2N5oB0_0(.dout(w_dff_A_qxSqAmE30_0),.din(w_dff_A_FNI2N5oB0_0),.clk(gclk));
	jdff dff_A_qxSqAmE30_0(.dout(w_dff_A_5kmgiiRM4_0),.din(w_dff_A_qxSqAmE30_0),.clk(gclk));
	jdff dff_A_5kmgiiRM4_0(.dout(w_dff_A_fZpHNZqr8_0),.din(w_dff_A_5kmgiiRM4_0),.clk(gclk));
	jdff dff_A_fZpHNZqr8_0(.dout(w_dff_A_1O928NQu3_0),.din(w_dff_A_fZpHNZqr8_0),.clk(gclk));
	jdff dff_A_1O928NQu3_0(.dout(w_dff_A_C6KvVvRw4_0),.din(w_dff_A_1O928NQu3_0),.clk(gclk));
	jdff dff_A_C6KvVvRw4_0(.dout(w_dff_A_NzqAHX8J0_0),.din(w_dff_A_C6KvVvRw4_0),.clk(gclk));
	jdff dff_A_NzqAHX8J0_0(.dout(w_dff_A_xhWMExsS6_0),.din(w_dff_A_NzqAHX8J0_0),.clk(gclk));
	jdff dff_A_xhWMExsS6_0(.dout(w_dff_A_D0YIkcmq8_0),.din(w_dff_A_xhWMExsS6_0),.clk(gclk));
	jdff dff_A_D0YIkcmq8_0(.dout(G621),.din(w_dff_A_D0YIkcmq8_0),.clk(gclk));
	jdff dff_A_pW3zWuB61_2(.dout(w_dff_A_iuhgNjMk9_0),.din(w_dff_A_pW3zWuB61_2),.clk(gclk));
	jdff dff_A_iuhgNjMk9_0(.dout(w_dff_A_0btv8qbN4_0),.din(w_dff_A_iuhgNjMk9_0),.clk(gclk));
	jdff dff_A_0btv8qbN4_0(.dout(w_dff_A_Fvk6Rn4J5_0),.din(w_dff_A_0btv8qbN4_0),.clk(gclk));
	jdff dff_A_Fvk6Rn4J5_0(.dout(w_dff_A_ucJdm4dT2_0),.din(w_dff_A_Fvk6Rn4J5_0),.clk(gclk));
	jdff dff_A_ucJdm4dT2_0(.dout(w_dff_A_qkcwqVzg9_0),.din(w_dff_A_ucJdm4dT2_0),.clk(gclk));
	jdff dff_A_qkcwqVzg9_0(.dout(w_dff_A_dFplCsJf4_0),.din(w_dff_A_qkcwqVzg9_0),.clk(gclk));
	jdff dff_A_dFplCsJf4_0(.dout(w_dff_A_8JPelck91_0),.din(w_dff_A_dFplCsJf4_0),.clk(gclk));
	jdff dff_A_8JPelck91_0(.dout(w_dff_A_PRTB8Ws46_0),.din(w_dff_A_8JPelck91_0),.clk(gclk));
	jdff dff_A_PRTB8Ws46_0(.dout(w_dff_A_U2gk24EX5_0),.din(w_dff_A_PRTB8Ws46_0),.clk(gclk));
	jdff dff_A_U2gk24EX5_0(.dout(w_dff_A_TDcCbFpz4_0),.din(w_dff_A_U2gk24EX5_0),.clk(gclk));
	jdff dff_A_TDcCbFpz4_0(.dout(w_dff_A_jytQ3geU6_0),.din(w_dff_A_TDcCbFpz4_0),.clk(gclk));
	jdff dff_A_jytQ3geU6_0(.dout(G629),.din(w_dff_A_jytQ3geU6_0),.clk(gclk));
	jdff dff_A_St9eEOx71_1(.dout(w_dff_A_28mVbJ1Z5_0),.din(w_dff_A_St9eEOx71_1),.clk(gclk));
	jdff dff_A_28mVbJ1Z5_0(.dout(w_dff_A_goPkPOBL5_0),.din(w_dff_A_28mVbJ1Z5_0),.clk(gclk));
	jdff dff_A_goPkPOBL5_0(.dout(w_dff_A_b7hYGBal6_0),.din(w_dff_A_goPkPOBL5_0),.clk(gclk));
	jdff dff_A_b7hYGBal6_0(.dout(w_dff_A_YlYZW9CP0_0),.din(w_dff_A_b7hYGBal6_0),.clk(gclk));
	jdff dff_A_YlYZW9CP0_0(.dout(w_dff_A_54xN6qlU2_0),.din(w_dff_A_YlYZW9CP0_0),.clk(gclk));
	jdff dff_A_54xN6qlU2_0(.dout(w_dff_A_1EkmCJbj1_0),.din(w_dff_A_54xN6qlU2_0),.clk(gclk));
	jdff dff_A_1EkmCJbj1_0(.dout(w_dff_A_dhvbG9Hp7_0),.din(w_dff_A_1EkmCJbj1_0),.clk(gclk));
	jdff dff_A_dhvbG9Hp7_0(.dout(w_dff_A_Toz8Cyf38_0),.din(w_dff_A_dhvbG9Hp7_0),.clk(gclk));
	jdff dff_A_Toz8Cyf38_0(.dout(w_dff_A_9z8b24NF3_0),.din(w_dff_A_Toz8Cyf38_0),.clk(gclk));
	jdff dff_A_9z8b24NF3_0(.dout(w_dff_A_Oi2rYkvS8_0),.din(w_dff_A_9z8b24NF3_0),.clk(gclk));
	jdff dff_A_Oi2rYkvS8_0(.dout(w_dff_A_TZIFYD3p2_0),.din(w_dff_A_Oi2rYkvS8_0),.clk(gclk));
	jdff dff_A_TZIFYD3p2_0(.dout(w_dff_A_3B1wfRkm1_0),.din(w_dff_A_TZIFYD3p2_0),.clk(gclk));
	jdff dff_A_3B1wfRkm1_0(.dout(w_dff_A_zkPkpbQs3_0),.din(w_dff_A_3B1wfRkm1_0),.clk(gclk));
	jdff dff_A_zkPkpbQs3_0(.dout(w_dff_A_kQaVA9b58_0),.din(w_dff_A_zkPkpbQs3_0),.clk(gclk));
	jdff dff_A_kQaVA9b58_0(.dout(w_dff_A_080eNj162_0),.din(w_dff_A_kQaVA9b58_0),.clk(gclk));
	jdff dff_A_080eNj162_0(.dout(w_dff_A_gbqxKkWf3_0),.din(w_dff_A_080eNj162_0),.clk(gclk));
	jdff dff_A_gbqxKkWf3_0(.dout(w_dff_A_mWCct4wI7_0),.din(w_dff_A_gbqxKkWf3_0),.clk(gclk));
	jdff dff_A_mWCct4wI7_0(.dout(w_dff_A_7peJnpA54_0),.din(w_dff_A_mWCct4wI7_0),.clk(gclk));
	jdff dff_A_7peJnpA54_0(.dout(G822),.din(w_dff_A_7peJnpA54_0),.clk(gclk));
	jdff dff_A_YdqD4BPM6_1(.dout(w_dff_A_HTJ3dgCR4_0),.din(w_dff_A_YdqD4BPM6_1),.clk(gclk));
	jdff dff_A_HTJ3dgCR4_0(.dout(w_dff_A_uZRmZeWc7_0),.din(w_dff_A_HTJ3dgCR4_0),.clk(gclk));
	jdff dff_A_uZRmZeWc7_0(.dout(w_dff_A_5NiqtKD21_0),.din(w_dff_A_uZRmZeWc7_0),.clk(gclk));
	jdff dff_A_5NiqtKD21_0(.dout(w_dff_A_ZbxeuFVB9_0),.din(w_dff_A_5NiqtKD21_0),.clk(gclk));
	jdff dff_A_ZbxeuFVB9_0(.dout(w_dff_A_v6c3OxBq7_0),.din(w_dff_A_ZbxeuFVB9_0),.clk(gclk));
	jdff dff_A_v6c3OxBq7_0(.dout(w_dff_A_IaM5GIxE4_0),.din(w_dff_A_v6c3OxBq7_0),.clk(gclk));
	jdff dff_A_IaM5GIxE4_0(.dout(w_dff_A_mX0o1eqC2_0),.din(w_dff_A_IaM5GIxE4_0),.clk(gclk));
	jdff dff_A_mX0o1eqC2_0(.dout(w_dff_A_zqHrxjU17_0),.din(w_dff_A_mX0o1eqC2_0),.clk(gclk));
	jdff dff_A_zqHrxjU17_0(.dout(w_dff_A_kq9v8JyC2_0),.din(w_dff_A_zqHrxjU17_0),.clk(gclk));
	jdff dff_A_kq9v8JyC2_0(.dout(w_dff_A_JwpVFd7m3_0),.din(w_dff_A_kq9v8JyC2_0),.clk(gclk));
	jdff dff_A_JwpVFd7m3_0(.dout(w_dff_A_wEb8cgZo2_0),.din(w_dff_A_JwpVFd7m3_0),.clk(gclk));
	jdff dff_A_wEb8cgZo2_0(.dout(w_dff_A_mmNzRu3N0_0),.din(w_dff_A_wEb8cgZo2_0),.clk(gclk));
	jdff dff_A_mmNzRu3N0_0(.dout(w_dff_A_wwsAQM7y3_0),.din(w_dff_A_mmNzRu3N0_0),.clk(gclk));
	jdff dff_A_wwsAQM7y3_0(.dout(w_dff_A_WRqjnmJp9_0),.din(w_dff_A_wwsAQM7y3_0),.clk(gclk));
	jdff dff_A_WRqjnmJp9_0(.dout(w_dff_A_Y9r4UMe27_0),.din(w_dff_A_WRqjnmJp9_0),.clk(gclk));
	jdff dff_A_Y9r4UMe27_0(.dout(w_dff_A_RD1lG3ow5_0),.din(w_dff_A_Y9r4UMe27_0),.clk(gclk));
	jdff dff_A_RD1lG3ow5_0(.dout(w_dff_A_ltiR10Xa4_0),.din(w_dff_A_RD1lG3ow5_0),.clk(gclk));
	jdff dff_A_ltiR10Xa4_0(.dout(G838),.din(w_dff_A_ltiR10Xa4_0),.clk(gclk));
	jdff dff_A_CnsGiYrK3_1(.dout(w_dff_A_83EKGves6_0),.din(w_dff_A_CnsGiYrK3_1),.clk(gclk));
	jdff dff_A_83EKGves6_0(.dout(w_dff_A_vJPsZl701_0),.din(w_dff_A_83EKGves6_0),.clk(gclk));
	jdff dff_A_vJPsZl701_0(.dout(w_dff_A_y2Xoglld7_0),.din(w_dff_A_vJPsZl701_0),.clk(gclk));
	jdff dff_A_y2Xoglld7_0(.dout(w_dff_A_8SvZ74Qm2_0),.din(w_dff_A_y2Xoglld7_0),.clk(gclk));
	jdff dff_A_8SvZ74Qm2_0(.dout(w_dff_A_pOp9XGEc4_0),.din(w_dff_A_8SvZ74Qm2_0),.clk(gclk));
	jdff dff_A_pOp9XGEc4_0(.dout(w_dff_A_C6CLZAK44_0),.din(w_dff_A_pOp9XGEc4_0),.clk(gclk));
	jdff dff_A_C6CLZAK44_0(.dout(w_dff_A_fq9BW8Aj6_0),.din(w_dff_A_C6CLZAK44_0),.clk(gclk));
	jdff dff_A_fq9BW8Aj6_0(.dout(w_dff_A_UlaYkN8l8_0),.din(w_dff_A_fq9BW8Aj6_0),.clk(gclk));
	jdff dff_A_UlaYkN8l8_0(.dout(w_dff_A_DhcYCfRX8_0),.din(w_dff_A_UlaYkN8l8_0),.clk(gclk));
	jdff dff_A_DhcYCfRX8_0(.dout(w_dff_A_4llKW2k82_0),.din(w_dff_A_DhcYCfRX8_0),.clk(gclk));
	jdff dff_A_4llKW2k82_0(.dout(w_dff_A_Z9I3IhsS7_0),.din(w_dff_A_4llKW2k82_0),.clk(gclk));
	jdff dff_A_Z9I3IhsS7_0(.dout(w_dff_A_uy0SWKff0_0),.din(w_dff_A_Z9I3IhsS7_0),.clk(gclk));
	jdff dff_A_uy0SWKff0_0(.dout(w_dff_A_eaUrWHnD8_0),.din(w_dff_A_uy0SWKff0_0),.clk(gclk));
	jdff dff_A_eaUrWHnD8_0(.dout(w_dff_A_LbwBuooE3_0),.din(w_dff_A_eaUrWHnD8_0),.clk(gclk));
	jdff dff_A_LbwBuooE3_0(.dout(w_dff_A_SwDsi6jB6_0),.din(w_dff_A_LbwBuooE3_0),.clk(gclk));
	jdff dff_A_SwDsi6jB6_0(.dout(w_dff_A_NXQF4HCr1_0),.din(w_dff_A_SwDsi6jB6_0),.clk(gclk));
	jdff dff_A_NXQF4HCr1_0(.dout(w_dff_A_yjsLMZjX3_0),.din(w_dff_A_NXQF4HCr1_0),.clk(gclk));
	jdff dff_A_yjsLMZjX3_0(.dout(G861),.din(w_dff_A_yjsLMZjX3_0),.clk(gclk));
	jdff dff_A_k5yPLMrJ3_1(.dout(w_dff_A_fvq3IfaD1_0),.din(w_dff_A_k5yPLMrJ3_1),.clk(gclk));
	jdff dff_A_fvq3IfaD1_0(.dout(w_dff_A_k6II2E9H3_0),.din(w_dff_A_fvq3IfaD1_0),.clk(gclk));
	jdff dff_A_k6II2E9H3_0(.dout(w_dff_A_sa7mXR8O1_0),.din(w_dff_A_k6II2E9H3_0),.clk(gclk));
	jdff dff_A_sa7mXR8O1_0(.dout(w_dff_A_aINk9Eez8_0),.din(w_dff_A_sa7mXR8O1_0),.clk(gclk));
	jdff dff_A_aINk9Eez8_0(.dout(w_dff_A_JFc5wbhj1_0),.din(w_dff_A_aINk9Eez8_0),.clk(gclk));
	jdff dff_A_JFc5wbhj1_0(.dout(w_dff_A_kwa8IYkA3_0),.din(w_dff_A_JFc5wbhj1_0),.clk(gclk));
	jdff dff_A_kwa8IYkA3_0(.dout(G623),.din(w_dff_A_kwa8IYkA3_0),.clk(gclk));
	jdff dff_A_GvPDbonV7_2(.dout(w_dff_A_nOSyCAkd3_0),.din(w_dff_A_GvPDbonV7_2),.clk(gclk));
	jdff dff_A_nOSyCAkd3_0(.dout(w_dff_A_jU9lzuWV8_0),.din(w_dff_A_nOSyCAkd3_0),.clk(gclk));
	jdff dff_A_jU9lzuWV8_0(.dout(w_dff_A_PKIvM7vx3_0),.din(w_dff_A_jU9lzuWV8_0),.clk(gclk));
	jdff dff_A_PKIvM7vx3_0(.dout(w_dff_A_ZQ72ZoxQ3_0),.din(w_dff_A_PKIvM7vx3_0),.clk(gclk));
	jdff dff_A_ZQ72ZoxQ3_0(.dout(w_dff_A_cviQh5KU4_0),.din(w_dff_A_ZQ72ZoxQ3_0),.clk(gclk));
	jdff dff_A_cviQh5KU4_0(.dout(w_dff_A_Ynk9Rojw0_0),.din(w_dff_A_cviQh5KU4_0),.clk(gclk));
	jdff dff_A_Ynk9Rojw0_0(.dout(w_dff_A_8BGQ4quh3_0),.din(w_dff_A_Ynk9Rojw0_0),.clk(gclk));
	jdff dff_A_8BGQ4quh3_0(.dout(w_dff_A_WXGd0sNX2_0),.din(w_dff_A_8BGQ4quh3_0),.clk(gclk));
	jdff dff_A_WXGd0sNX2_0(.dout(w_dff_A_3Wg9Z3FU3_0),.din(w_dff_A_WXGd0sNX2_0),.clk(gclk));
	jdff dff_A_3Wg9Z3FU3_0(.dout(w_dff_A_Ic59kQtS7_0),.din(w_dff_A_3Wg9Z3FU3_0),.clk(gclk));
	jdff dff_A_Ic59kQtS7_0(.dout(w_dff_A_BWxXN7Q49_0),.din(w_dff_A_Ic59kQtS7_0),.clk(gclk));
	jdff dff_A_BWxXN7Q49_0(.dout(w_dff_A_599oNvDw3_0),.din(w_dff_A_BWxXN7Q49_0),.clk(gclk));
	jdff dff_A_599oNvDw3_0(.dout(w_dff_A_wDus7Xlx0_0),.din(w_dff_A_599oNvDw3_0),.clk(gclk));
	jdff dff_A_wDus7Xlx0_0(.dout(w_dff_A_zizyxwgW1_0),.din(w_dff_A_wDus7Xlx0_0),.clk(gclk));
	jdff dff_A_zizyxwgW1_0(.dout(G722),.din(w_dff_A_zizyxwgW1_0),.clk(gclk));
	jdff dff_A_ZffOHOwP8_1(.dout(w_dff_A_oW5c9Yys4_0),.din(w_dff_A_ZffOHOwP8_1),.clk(gclk));
	jdff dff_A_oW5c9Yys4_0(.dout(w_dff_A_aoX9PM4h8_0),.din(w_dff_A_oW5c9Yys4_0),.clk(gclk));
	jdff dff_A_aoX9PM4h8_0(.dout(w_dff_A_l1oc758E6_0),.din(w_dff_A_aoX9PM4h8_0),.clk(gclk));
	jdff dff_A_l1oc758E6_0(.dout(w_dff_A_5fYMrykJ1_0),.din(w_dff_A_l1oc758E6_0),.clk(gclk));
	jdff dff_A_5fYMrykJ1_0(.dout(w_dff_A_GINYGC9z5_0),.din(w_dff_A_5fYMrykJ1_0),.clk(gclk));
	jdff dff_A_GINYGC9z5_0(.dout(w_dff_A_A6p88IdL0_0),.din(w_dff_A_GINYGC9z5_0),.clk(gclk));
	jdff dff_A_A6p88IdL0_0(.dout(w_dff_A_0QIqRIev7_0),.din(w_dff_A_A6p88IdL0_0),.clk(gclk));
	jdff dff_A_0QIqRIev7_0(.dout(w_dff_A_p4Ml6w9n1_0),.din(w_dff_A_0QIqRIev7_0),.clk(gclk));
	jdff dff_A_p4Ml6w9n1_0(.dout(w_dff_A_p2ELthUi3_0),.din(w_dff_A_p4Ml6w9n1_0),.clk(gclk));
	jdff dff_A_p2ELthUi3_0(.dout(w_dff_A_U0md0XSE7_0),.din(w_dff_A_p2ELthUi3_0),.clk(gclk));
	jdff dff_A_U0md0XSE7_0(.dout(w_dff_A_8CNkI0eU4_0),.din(w_dff_A_U0md0XSE7_0),.clk(gclk));
	jdff dff_A_8CNkI0eU4_0(.dout(G832),.din(w_dff_A_8CNkI0eU4_0),.clk(gclk));
	jdff dff_A_msTcj59W3_1(.dout(w_dff_A_G5MbsiEP4_0),.din(w_dff_A_msTcj59W3_1),.clk(gclk));
	jdff dff_A_G5MbsiEP4_0(.dout(w_dff_A_bOsgKylV9_0),.din(w_dff_A_G5MbsiEP4_0),.clk(gclk));
	jdff dff_A_bOsgKylV9_0(.dout(w_dff_A_30rWTXLk2_0),.din(w_dff_A_bOsgKylV9_0),.clk(gclk));
	jdff dff_A_30rWTXLk2_0(.dout(w_dff_A_6X6SDLcT4_0),.din(w_dff_A_30rWTXLk2_0),.clk(gclk));
	jdff dff_A_6X6SDLcT4_0(.dout(w_dff_A_jUpFiyuG7_0),.din(w_dff_A_6X6SDLcT4_0),.clk(gclk));
	jdff dff_A_jUpFiyuG7_0(.dout(w_dff_A_ZTjhmtnF4_0),.din(w_dff_A_jUpFiyuG7_0),.clk(gclk));
	jdff dff_A_ZTjhmtnF4_0(.dout(w_dff_A_kFPYv3nn6_0),.din(w_dff_A_ZTjhmtnF4_0),.clk(gclk));
	jdff dff_A_kFPYv3nn6_0(.dout(w_dff_A_sNo9Dghe2_0),.din(w_dff_A_kFPYv3nn6_0),.clk(gclk));
	jdff dff_A_sNo9Dghe2_0(.dout(w_dff_A_HiM0Gdkd7_0),.din(w_dff_A_sNo9Dghe2_0),.clk(gclk));
	jdff dff_A_HiM0Gdkd7_0(.dout(w_dff_A_oTtU9Rbv7_0),.din(w_dff_A_HiM0Gdkd7_0),.clk(gclk));
	jdff dff_A_oTtU9Rbv7_0(.dout(w_dff_A_SWTTSma93_0),.din(w_dff_A_oTtU9Rbv7_0),.clk(gclk));
	jdff dff_A_SWTTSma93_0(.dout(w_dff_A_0XJcPhsN7_0),.din(w_dff_A_SWTTSma93_0),.clk(gclk));
	jdff dff_A_0XJcPhsN7_0(.dout(w_dff_A_tkE1fDqo8_0),.din(w_dff_A_0XJcPhsN7_0),.clk(gclk));
	jdff dff_A_tkE1fDqo8_0(.dout(G834),.din(w_dff_A_tkE1fDqo8_0),.clk(gclk));
	jdff dff_A_DncwKVdg0_1(.dout(w_dff_A_tnnEG8Ec3_0),.din(w_dff_A_DncwKVdg0_1),.clk(gclk));
	jdff dff_A_tnnEG8Ec3_0(.dout(w_dff_A_9RApjLTs8_0),.din(w_dff_A_tnnEG8Ec3_0),.clk(gclk));
	jdff dff_A_9RApjLTs8_0(.dout(w_dff_A_vGznwiUd3_0),.din(w_dff_A_9RApjLTs8_0),.clk(gclk));
	jdff dff_A_vGznwiUd3_0(.dout(w_dff_A_2ITdwgpn3_0),.din(w_dff_A_vGznwiUd3_0),.clk(gclk));
	jdff dff_A_2ITdwgpn3_0(.dout(w_dff_A_NLL83CuD4_0),.din(w_dff_A_2ITdwgpn3_0),.clk(gclk));
	jdff dff_A_NLL83CuD4_0(.dout(w_dff_A_ncehto3S7_0),.din(w_dff_A_NLL83CuD4_0),.clk(gclk));
	jdff dff_A_ncehto3S7_0(.dout(w_dff_A_kas13WDr1_0),.din(w_dff_A_ncehto3S7_0),.clk(gclk));
	jdff dff_A_kas13WDr1_0(.dout(w_dff_A_XHruMOpB4_0),.din(w_dff_A_kas13WDr1_0),.clk(gclk));
	jdff dff_A_XHruMOpB4_0(.dout(w_dff_A_r1SwHZWk8_0),.din(w_dff_A_XHruMOpB4_0),.clk(gclk));
	jdff dff_A_r1SwHZWk8_0(.dout(w_dff_A_Sq7VWW7F2_0),.din(w_dff_A_r1SwHZWk8_0),.clk(gclk));
	jdff dff_A_Sq7VWW7F2_0(.dout(w_dff_A_duDx3le64_0),.din(w_dff_A_Sq7VWW7F2_0),.clk(gclk));
	jdff dff_A_duDx3le64_0(.dout(w_dff_A_DL6aqxX38_0),.din(w_dff_A_duDx3le64_0),.clk(gclk));
	jdff dff_A_DL6aqxX38_0(.dout(w_dff_A_eFrnj7hA1_0),.din(w_dff_A_DL6aqxX38_0),.clk(gclk));
	jdff dff_A_eFrnj7hA1_0(.dout(w_dff_A_NVcIuwAK2_0),.din(w_dff_A_eFrnj7hA1_0),.clk(gclk));
	jdff dff_A_NVcIuwAK2_0(.dout(w_dff_A_8Sppg9R88_0),.din(w_dff_A_NVcIuwAK2_0),.clk(gclk));
	jdff dff_A_8Sppg9R88_0(.dout(G836),.din(w_dff_A_8Sppg9R88_0),.clk(gclk));
	jdff dff_A_8TrmV4bo1_2(.dout(w_dff_A_fzwUM4R65_0),.din(w_dff_A_8TrmV4bo1_2),.clk(gclk));
	jdff dff_A_fzwUM4R65_0(.dout(w_dff_A_0TgI2VJp1_0),.din(w_dff_A_fzwUM4R65_0),.clk(gclk));
	jdff dff_A_0TgI2VJp1_0(.dout(w_dff_A_exINZv4C0_0),.din(w_dff_A_0TgI2VJp1_0),.clk(gclk));
	jdff dff_A_exINZv4C0_0(.dout(w_dff_A_FUM9BEya1_0),.din(w_dff_A_exINZv4C0_0),.clk(gclk));
	jdff dff_A_FUM9BEya1_0(.dout(w_dff_A_TRWfubfV1_0),.din(w_dff_A_FUM9BEya1_0),.clk(gclk));
	jdff dff_A_TRWfubfV1_0(.dout(w_dff_A_XH9IXdoh1_0),.din(w_dff_A_TRWfubfV1_0),.clk(gclk));
	jdff dff_A_XH9IXdoh1_0(.dout(w_dff_A_C4theoMg4_0),.din(w_dff_A_XH9IXdoh1_0),.clk(gclk));
	jdff dff_A_C4theoMg4_0(.dout(w_dff_A_lfP9KjOp0_0),.din(w_dff_A_C4theoMg4_0),.clk(gclk));
	jdff dff_A_lfP9KjOp0_0(.dout(w_dff_A_IGWmh2l21_0),.din(w_dff_A_lfP9KjOp0_0),.clk(gclk));
	jdff dff_A_IGWmh2l21_0(.dout(w_dff_A_yOj7mIoi4_0),.din(w_dff_A_IGWmh2l21_0),.clk(gclk));
	jdff dff_A_yOj7mIoi4_0(.dout(w_dff_A_oqpB9X5S2_0),.din(w_dff_A_yOj7mIoi4_0),.clk(gclk));
	jdff dff_A_oqpB9X5S2_0(.dout(w_dff_A_gdq1cazK1_0),.din(w_dff_A_oqpB9X5S2_0),.clk(gclk));
	jdff dff_A_gdq1cazK1_0(.dout(w_dff_A_6MRdUHit8_0),.din(w_dff_A_gdq1cazK1_0),.clk(gclk));
	jdff dff_A_6MRdUHit8_0(.dout(w_dff_A_NrW5qRyb0_0),.din(w_dff_A_6MRdUHit8_0),.clk(gclk));
	jdff dff_A_NrW5qRyb0_0(.dout(G859),.din(w_dff_A_NrW5qRyb0_0),.clk(gclk));
	jdff dff_A_IXVtm8zU8_1(.dout(w_dff_A_mB5v21pN5_0),.din(w_dff_A_IXVtm8zU8_1),.clk(gclk));
	jdff dff_A_mB5v21pN5_0(.dout(w_dff_A_sTsNouiN8_0),.din(w_dff_A_mB5v21pN5_0),.clk(gclk));
	jdff dff_A_sTsNouiN8_0(.dout(w_dff_A_S4my90vB1_0),.din(w_dff_A_sTsNouiN8_0),.clk(gclk));
	jdff dff_A_S4my90vB1_0(.dout(w_dff_A_cwFEfvcJ1_0),.din(w_dff_A_S4my90vB1_0),.clk(gclk));
	jdff dff_A_cwFEfvcJ1_0(.dout(w_dff_A_EoNNZtM72_0),.din(w_dff_A_cwFEfvcJ1_0),.clk(gclk));
	jdff dff_A_EoNNZtM72_0(.dout(w_dff_A_rlLH4CzB7_0),.din(w_dff_A_EoNNZtM72_0),.clk(gclk));
	jdff dff_A_rlLH4CzB7_0(.dout(w_dff_A_DXI2DKSU4_0),.din(w_dff_A_rlLH4CzB7_0),.clk(gclk));
	jdff dff_A_DXI2DKSU4_0(.dout(w_dff_A_8aLZA2Wn5_0),.din(w_dff_A_DXI2DKSU4_0),.clk(gclk));
	jdff dff_A_8aLZA2Wn5_0(.dout(w_dff_A_hEMT2bfT0_0),.din(w_dff_A_8aLZA2Wn5_0),.clk(gclk));
	jdff dff_A_hEMT2bfT0_0(.dout(G871),.din(w_dff_A_hEMT2bfT0_0),.clk(gclk));
	jdff dff_A_NIZhYMSx1_1(.dout(w_dff_A_jFbfgyKv5_0),.din(w_dff_A_NIZhYMSx1_1),.clk(gclk));
	jdff dff_A_jFbfgyKv5_0(.dout(w_dff_A_eh8TOSl19_0),.din(w_dff_A_jFbfgyKv5_0),.clk(gclk));
	jdff dff_A_eh8TOSl19_0(.dout(w_dff_A_1bpmZKHO7_0),.din(w_dff_A_eh8TOSl19_0),.clk(gclk));
	jdff dff_A_1bpmZKHO7_0(.dout(w_dff_A_8NmM8OaC8_0),.din(w_dff_A_1bpmZKHO7_0),.clk(gclk));
	jdff dff_A_8NmM8OaC8_0(.dout(w_dff_A_GfU1i5mF8_0),.din(w_dff_A_8NmM8OaC8_0),.clk(gclk));
	jdff dff_A_GfU1i5mF8_0(.dout(w_dff_A_vnlUsT7q5_0),.din(w_dff_A_GfU1i5mF8_0),.clk(gclk));
	jdff dff_A_vnlUsT7q5_0(.dout(w_dff_A_eqLJrOBc0_0),.din(w_dff_A_vnlUsT7q5_0),.clk(gclk));
	jdff dff_A_eqLJrOBc0_0(.dout(w_dff_A_gd9cEWXz6_0),.din(w_dff_A_eqLJrOBc0_0),.clk(gclk));
	jdff dff_A_gd9cEWXz6_0(.dout(w_dff_A_MXURVI2L3_0),.din(w_dff_A_gd9cEWXz6_0),.clk(gclk));
	jdff dff_A_MXURVI2L3_0(.dout(w_dff_A_TSBzS8134_0),.din(w_dff_A_MXURVI2L3_0),.clk(gclk));
	jdff dff_A_TSBzS8134_0(.dout(w_dff_A_o2n5yBar4_0),.din(w_dff_A_TSBzS8134_0),.clk(gclk));
	jdff dff_A_o2n5yBar4_0(.dout(G873),.din(w_dff_A_o2n5yBar4_0),.clk(gclk));
	jdff dff_A_wxyThvto1_1(.dout(w_dff_A_Oq0L4EC19_0),.din(w_dff_A_wxyThvto1_1),.clk(gclk));
	jdff dff_A_Oq0L4EC19_0(.dout(w_dff_A_fXrKLlaH6_0),.din(w_dff_A_Oq0L4EC19_0),.clk(gclk));
	jdff dff_A_fXrKLlaH6_0(.dout(w_dff_A_T4RqAqNP5_0),.din(w_dff_A_fXrKLlaH6_0),.clk(gclk));
	jdff dff_A_T4RqAqNP5_0(.dout(w_dff_A_DJcXeLtS2_0),.din(w_dff_A_T4RqAqNP5_0),.clk(gclk));
	jdff dff_A_DJcXeLtS2_0(.dout(w_dff_A_VNLv3DNN9_0),.din(w_dff_A_DJcXeLtS2_0),.clk(gclk));
	jdff dff_A_VNLv3DNN9_0(.dout(w_dff_A_4PTJZ3kK0_0),.din(w_dff_A_VNLv3DNN9_0),.clk(gclk));
	jdff dff_A_4PTJZ3kK0_0(.dout(w_dff_A_TP6gSsnx5_0),.din(w_dff_A_4PTJZ3kK0_0),.clk(gclk));
	jdff dff_A_TP6gSsnx5_0(.dout(w_dff_A_gbDFa50o7_0),.din(w_dff_A_TP6gSsnx5_0),.clk(gclk));
	jdff dff_A_gbDFa50o7_0(.dout(w_dff_A_KRg67GBY7_0),.din(w_dff_A_gbDFa50o7_0),.clk(gclk));
	jdff dff_A_KRg67GBY7_0(.dout(w_dff_A_7ghoOdvN1_0),.din(w_dff_A_KRg67GBY7_0),.clk(gclk));
	jdff dff_A_7ghoOdvN1_0(.dout(w_dff_A_ZL9nOHXE2_0),.din(w_dff_A_7ghoOdvN1_0),.clk(gclk));
	jdff dff_A_ZL9nOHXE2_0(.dout(w_dff_A_ohaO0QbP3_0),.din(w_dff_A_ZL9nOHXE2_0),.clk(gclk));
	jdff dff_A_ohaO0QbP3_0(.dout(G875),.din(w_dff_A_ohaO0QbP3_0),.clk(gclk));
	jdff dff_A_y2fvlRfV5_1(.dout(w_dff_A_LnYSCbXn9_0),.din(w_dff_A_y2fvlRfV5_1),.clk(gclk));
	jdff dff_A_LnYSCbXn9_0(.dout(w_dff_A_f6lpTfON3_0),.din(w_dff_A_LnYSCbXn9_0),.clk(gclk));
	jdff dff_A_f6lpTfON3_0(.dout(w_dff_A_CciD38DR3_0),.din(w_dff_A_f6lpTfON3_0),.clk(gclk));
	jdff dff_A_CciD38DR3_0(.dout(w_dff_A_LrwxJvo53_0),.din(w_dff_A_CciD38DR3_0),.clk(gclk));
	jdff dff_A_LrwxJvo53_0(.dout(w_dff_A_eNXeGQas8_0),.din(w_dff_A_LrwxJvo53_0),.clk(gclk));
	jdff dff_A_eNXeGQas8_0(.dout(w_dff_A_o6GTmLG27_0),.din(w_dff_A_eNXeGQas8_0),.clk(gclk));
	jdff dff_A_o6GTmLG27_0(.dout(w_dff_A_PFpfjHWI0_0),.din(w_dff_A_o6GTmLG27_0),.clk(gclk));
	jdff dff_A_PFpfjHWI0_0(.dout(w_dff_A_kuafdsuF8_0),.din(w_dff_A_PFpfjHWI0_0),.clk(gclk));
	jdff dff_A_kuafdsuF8_0(.dout(w_dff_A_SHCZbjsl4_0),.din(w_dff_A_kuafdsuF8_0),.clk(gclk));
	jdff dff_A_SHCZbjsl4_0(.dout(w_dff_A_miEUHJyN4_0),.din(w_dff_A_SHCZbjsl4_0),.clk(gclk));
	jdff dff_A_miEUHJyN4_0(.dout(w_dff_A_I8dm8M1B8_0),.din(w_dff_A_miEUHJyN4_0),.clk(gclk));
	jdff dff_A_I8dm8M1B8_0(.dout(w_dff_A_vvM4LYCS8_0),.din(w_dff_A_I8dm8M1B8_0),.clk(gclk));
	jdff dff_A_vvM4LYCS8_0(.dout(w_dff_A_N3gyNNC57_0),.din(w_dff_A_vvM4LYCS8_0),.clk(gclk));
	jdff dff_A_N3gyNNC57_0(.dout(G877),.din(w_dff_A_N3gyNNC57_0),.clk(gclk));
	jdff dff_A_hy3XRMt16_1(.dout(w_dff_A_nlJ6vhn78_0),.din(w_dff_A_hy3XRMt16_1),.clk(gclk));
	jdff dff_A_nlJ6vhn78_0(.dout(w_dff_A_YgsIYrS27_0),.din(w_dff_A_nlJ6vhn78_0),.clk(gclk));
	jdff dff_A_YgsIYrS27_0(.dout(w_dff_A_sVtdwruG0_0),.din(w_dff_A_YgsIYrS27_0),.clk(gclk));
	jdff dff_A_sVtdwruG0_0(.dout(w_dff_A_TvKM6GDk6_0),.din(w_dff_A_sVtdwruG0_0),.clk(gclk));
	jdff dff_A_TvKM6GDk6_0(.dout(w_dff_A_By65h7ve9_0),.din(w_dff_A_TvKM6GDk6_0),.clk(gclk));
	jdff dff_A_By65h7ve9_0(.dout(w_dff_A_q2ep5t2e9_0),.din(w_dff_A_By65h7ve9_0),.clk(gclk));
	jdff dff_A_q2ep5t2e9_0(.dout(w_dff_A_6pvA1WnF9_0),.din(w_dff_A_q2ep5t2e9_0),.clk(gclk));
	jdff dff_A_6pvA1WnF9_0(.dout(w_dff_A_ZG5ktrdT5_0),.din(w_dff_A_6pvA1WnF9_0),.clk(gclk));
	jdff dff_A_ZG5ktrdT5_0(.dout(w_dff_A_EKkAAozQ3_0),.din(w_dff_A_ZG5ktrdT5_0),.clk(gclk));
	jdff dff_A_EKkAAozQ3_0(.dout(w_dff_A_LqGWjEKb4_0),.din(w_dff_A_EKkAAozQ3_0),.clk(gclk));
	jdff dff_A_LqGWjEKb4_0(.dout(w_dff_A_yyBRG0eW2_0),.din(w_dff_A_LqGWjEKb4_0),.clk(gclk));
	jdff dff_A_yyBRG0eW2_0(.dout(w_dff_A_3cu7Ywe51_0),.din(w_dff_A_yyBRG0eW2_0),.clk(gclk));
	jdff dff_A_3cu7Ywe51_0(.dout(w_dff_A_wBIAyGJL9_0),.din(w_dff_A_3cu7Ywe51_0),.clk(gclk));
	jdff dff_A_wBIAyGJL9_0(.dout(w_dff_A_ocAGjrj65_0),.din(w_dff_A_wBIAyGJL9_0),.clk(gclk));
	jdff dff_A_ocAGjrj65_0(.dout(w_dff_A_lavgTu5v9_0),.din(w_dff_A_ocAGjrj65_0),.clk(gclk));
	jdff dff_A_lavgTu5v9_0(.dout(w_dff_A_z2no7W9H4_0),.din(w_dff_A_lavgTu5v9_0),.clk(gclk));
	jdff dff_A_z2no7W9H4_0(.dout(G998),.din(w_dff_A_z2no7W9H4_0),.clk(gclk));
	jdff dff_A_yV3M3vWw4_1(.dout(w_dff_A_nxPx0cIa5_0),.din(w_dff_A_yV3M3vWw4_1),.clk(gclk));
	jdff dff_A_nxPx0cIa5_0(.dout(w_dff_A_5kYh2G7x1_0),.din(w_dff_A_nxPx0cIa5_0),.clk(gclk));
	jdff dff_A_5kYh2G7x1_0(.dout(w_dff_A_T8lqoWCL7_0),.din(w_dff_A_5kYh2G7x1_0),.clk(gclk));
	jdff dff_A_T8lqoWCL7_0(.dout(w_dff_A_Ypktngn25_0),.din(w_dff_A_T8lqoWCL7_0),.clk(gclk));
	jdff dff_A_Ypktngn25_0(.dout(w_dff_A_slSZQgGt1_0),.din(w_dff_A_Ypktngn25_0),.clk(gclk));
	jdff dff_A_slSZQgGt1_0(.dout(w_dff_A_l5VXW8zM2_0),.din(w_dff_A_slSZQgGt1_0),.clk(gclk));
	jdff dff_A_l5VXW8zM2_0(.dout(w_dff_A_4hkbVbUF9_0),.din(w_dff_A_l5VXW8zM2_0),.clk(gclk));
	jdff dff_A_4hkbVbUF9_0(.dout(w_dff_A_4Hk71Rpv7_0),.din(w_dff_A_4hkbVbUF9_0),.clk(gclk));
	jdff dff_A_4Hk71Rpv7_0(.dout(w_dff_A_wcunGtT17_0),.din(w_dff_A_4Hk71Rpv7_0),.clk(gclk));
	jdff dff_A_wcunGtT17_0(.dout(w_dff_A_njRTuOBR8_0),.din(w_dff_A_wcunGtT17_0),.clk(gclk));
	jdff dff_A_njRTuOBR8_0(.dout(w_dff_A_slk0RpSk6_0),.din(w_dff_A_njRTuOBR8_0),.clk(gclk));
	jdff dff_A_slk0RpSk6_0(.dout(w_dff_A_pfBskIu99_0),.din(w_dff_A_slk0RpSk6_0),.clk(gclk));
	jdff dff_A_pfBskIu99_0(.dout(w_dff_A_OhDAgSNI0_0),.din(w_dff_A_pfBskIu99_0),.clk(gclk));
	jdff dff_A_OhDAgSNI0_0(.dout(w_dff_A_PIs04hum8_0),.din(w_dff_A_OhDAgSNI0_0),.clk(gclk));
	jdff dff_A_PIs04hum8_0(.dout(w_dff_A_8LmpDHTm3_0),.din(w_dff_A_PIs04hum8_0),.clk(gclk));
	jdff dff_A_8LmpDHTm3_0(.dout(w_dff_A_A6MBRDD45_0),.din(w_dff_A_8LmpDHTm3_0),.clk(gclk));
	jdff dff_A_A6MBRDD45_0(.dout(w_dff_A_DHHKKRtK9_0),.din(w_dff_A_A6MBRDD45_0),.clk(gclk));
	jdff dff_A_DHHKKRtK9_0(.dout(w_dff_A_wcbljaey5_0),.din(w_dff_A_DHHKKRtK9_0),.clk(gclk));
	jdff dff_A_wcbljaey5_0(.dout(G1000),.din(w_dff_A_wcbljaey5_0),.clk(gclk));
	jdff dff_A_rzj3Gxf21_2(.dout(w_dff_A_S48jCoEZ7_0),.din(w_dff_A_rzj3Gxf21_2),.clk(gclk));
	jdff dff_A_S48jCoEZ7_0(.dout(w_dff_A_436cEISi1_0),.din(w_dff_A_S48jCoEZ7_0),.clk(gclk));
	jdff dff_A_436cEISi1_0(.dout(w_dff_A_MX9ZfvsT3_0),.din(w_dff_A_436cEISi1_0),.clk(gclk));
	jdff dff_A_MX9ZfvsT3_0(.dout(w_dff_A_KSpr5fVE0_0),.din(w_dff_A_MX9ZfvsT3_0),.clk(gclk));
	jdff dff_A_KSpr5fVE0_0(.dout(G575),.din(w_dff_A_KSpr5fVE0_0),.clk(gclk));
	jdff dff_A_OurWUoh22_2(.dout(w_dff_A_a4YtDaw40_0),.din(w_dff_A_OurWUoh22_2),.clk(gclk));
	jdff dff_A_a4YtDaw40_0(.dout(w_dff_A_6pYyqoxk1_0),.din(w_dff_A_a4YtDaw40_0),.clk(gclk));
	jdff dff_A_6pYyqoxk1_0(.dout(w_dff_A_ThUQVMEj6_0),.din(w_dff_A_6pYyqoxk1_0),.clk(gclk));
	jdff dff_A_ThUQVMEj6_0(.dout(w_dff_A_SHcAE3dZ9_0),.din(w_dff_A_ThUQVMEj6_0),.clk(gclk));
	jdff dff_A_SHcAE3dZ9_0(.dout(w_dff_A_GT0N0tKO8_0),.din(w_dff_A_SHcAE3dZ9_0),.clk(gclk));
	jdff dff_A_GT0N0tKO8_0(.dout(w_dff_A_P9zOJhhd5_0),.din(w_dff_A_GT0N0tKO8_0),.clk(gclk));
	jdff dff_A_P9zOJhhd5_0(.dout(w_dff_A_M4wuqmaJ9_0),.din(w_dff_A_P9zOJhhd5_0),.clk(gclk));
	jdff dff_A_M4wuqmaJ9_0(.dout(G585),.din(w_dff_A_M4wuqmaJ9_0),.clk(gclk));
	jdff dff_A_CdLv686k3_2(.dout(w_dff_A_wVnRgiAg5_0),.din(w_dff_A_CdLv686k3_2),.clk(gclk));
	jdff dff_A_wVnRgiAg5_0(.dout(w_dff_A_Rv1xzE9Q1_0),.din(w_dff_A_wVnRgiAg5_0),.clk(gclk));
	jdff dff_A_Rv1xzE9Q1_0(.dout(w_dff_A_t8FSO4NZ3_0),.din(w_dff_A_Rv1xzE9Q1_0),.clk(gclk));
	jdff dff_A_t8FSO4NZ3_0(.dout(w_dff_A_qvkchFAl0_0),.din(w_dff_A_t8FSO4NZ3_0),.clk(gclk));
	jdff dff_A_qvkchFAl0_0(.dout(w_dff_A_IBXzG8LL3_0),.din(w_dff_A_qvkchFAl0_0),.clk(gclk));
	jdff dff_A_IBXzG8LL3_0(.dout(w_dff_A_Am64hqcN0_0),.din(w_dff_A_IBXzG8LL3_0),.clk(gclk));
	jdff dff_A_Am64hqcN0_0(.dout(w_dff_A_XBItEODN1_0),.din(w_dff_A_Am64hqcN0_0),.clk(gclk));
	jdff dff_A_XBItEODN1_0(.dout(w_dff_A_YY3Ejfev2_0),.din(w_dff_A_XBItEODN1_0),.clk(gclk));
	jdff dff_A_YY3Ejfev2_0(.dout(w_dff_A_xvs258ej6_0),.din(w_dff_A_YY3Ejfev2_0),.clk(gclk));
	jdff dff_A_xvs258ej6_0(.dout(w_dff_A_pAvuaBLZ7_0),.din(w_dff_A_xvs258ej6_0),.clk(gclk));
	jdff dff_A_pAvuaBLZ7_0(.dout(w_dff_A_yYjyoZsI5_0),.din(w_dff_A_pAvuaBLZ7_0),.clk(gclk));
	jdff dff_A_yYjyoZsI5_0(.dout(w_dff_A_W6VhlTt27_0),.din(w_dff_A_yYjyoZsI5_0),.clk(gclk));
	jdff dff_A_W6VhlTt27_0(.dout(w_dff_A_wuqM8eDK6_0),.din(w_dff_A_W6VhlTt27_0),.clk(gclk));
	jdff dff_A_wuqM8eDK6_0(.dout(G661),.din(w_dff_A_wuqM8eDK6_0),.clk(gclk));
	jdff dff_A_eISRmwvG1_2(.dout(w_dff_A_DuJnvwwJ7_0),.din(w_dff_A_eISRmwvG1_2),.clk(gclk));
	jdff dff_A_DuJnvwwJ7_0(.dout(w_dff_A_IhZ6kUNN7_0),.din(w_dff_A_DuJnvwwJ7_0),.clk(gclk));
	jdff dff_A_IhZ6kUNN7_0(.dout(w_dff_A_79epYESg6_0),.din(w_dff_A_IhZ6kUNN7_0),.clk(gclk));
	jdff dff_A_79epYESg6_0(.dout(w_dff_A_xNo22IQ48_0),.din(w_dff_A_79epYESg6_0),.clk(gclk));
	jdff dff_A_xNo22IQ48_0(.dout(w_dff_A_mbfguTpo1_0),.din(w_dff_A_xNo22IQ48_0),.clk(gclk));
	jdff dff_A_mbfguTpo1_0(.dout(w_dff_A_TyWnQ3Gf6_0),.din(w_dff_A_mbfguTpo1_0),.clk(gclk));
	jdff dff_A_TyWnQ3Gf6_0(.dout(w_dff_A_qtOORKx37_0),.din(w_dff_A_TyWnQ3Gf6_0),.clk(gclk));
	jdff dff_A_qtOORKx37_0(.dout(w_dff_A_iIR2E4HM4_0),.din(w_dff_A_qtOORKx37_0),.clk(gclk));
	jdff dff_A_iIR2E4HM4_0(.dout(w_dff_A_vo6ZiUby3_0),.din(w_dff_A_iIR2E4HM4_0),.clk(gclk));
	jdff dff_A_vo6ZiUby3_0(.dout(w_dff_A_55iAiWu90_0),.din(w_dff_A_vo6ZiUby3_0),.clk(gclk));
	jdff dff_A_55iAiWu90_0(.dout(w_dff_A_3oMyx8CQ1_0),.din(w_dff_A_55iAiWu90_0),.clk(gclk));
	jdff dff_A_3oMyx8CQ1_0(.dout(w_dff_A_z9amqPRY5_0),.din(w_dff_A_3oMyx8CQ1_0),.clk(gclk));
	jdff dff_A_z9amqPRY5_0(.dout(w_dff_A_GzH6xKpN8_0),.din(w_dff_A_z9amqPRY5_0),.clk(gclk));
	jdff dff_A_GzH6xKpN8_0(.dout(G693),.din(w_dff_A_GzH6xKpN8_0),.clk(gclk));
	jdff dff_A_pbgvSBrL9_2(.dout(w_dff_A_yXroYVSS5_0),.din(w_dff_A_pbgvSBrL9_2),.clk(gclk));
	jdff dff_A_yXroYVSS5_0(.dout(w_dff_A_GCfkkTRs0_0),.din(w_dff_A_yXroYVSS5_0),.clk(gclk));
	jdff dff_A_GCfkkTRs0_0(.dout(w_dff_A_v7RLv10f3_0),.din(w_dff_A_GCfkkTRs0_0),.clk(gclk));
	jdff dff_A_v7RLv10f3_0(.dout(w_dff_A_vMTtlUYk2_0),.din(w_dff_A_v7RLv10f3_0),.clk(gclk));
	jdff dff_A_vMTtlUYk2_0(.dout(w_dff_A_wFZsi1fI6_0),.din(w_dff_A_vMTtlUYk2_0),.clk(gclk));
	jdff dff_A_wFZsi1fI6_0(.dout(w_dff_A_BhPHxHby8_0),.din(w_dff_A_wFZsi1fI6_0),.clk(gclk));
	jdff dff_A_BhPHxHby8_0(.dout(G747),.din(w_dff_A_BhPHxHby8_0),.clk(gclk));
	jdff dff_A_eFLyZN3r9_2(.dout(w_dff_A_qO2PfSKg0_0),.din(w_dff_A_eFLyZN3r9_2),.clk(gclk));
	jdff dff_A_qO2PfSKg0_0(.dout(w_dff_A_YYQfVngw2_0),.din(w_dff_A_qO2PfSKg0_0),.clk(gclk));
	jdff dff_A_YYQfVngw2_0(.dout(w_dff_A_tFBjUQuU0_0),.din(w_dff_A_YYQfVngw2_0),.clk(gclk));
	jdff dff_A_tFBjUQuU0_0(.dout(w_dff_A_iB1mXwn10_0),.din(w_dff_A_tFBjUQuU0_0),.clk(gclk));
	jdff dff_A_iB1mXwn10_0(.dout(w_dff_A_Sxr1TNJc6_0),.din(w_dff_A_iB1mXwn10_0),.clk(gclk));
	jdff dff_A_Sxr1TNJc6_0(.dout(w_dff_A_aU2zvkL33_0),.din(w_dff_A_Sxr1TNJc6_0),.clk(gclk));
	jdff dff_A_aU2zvkL33_0(.dout(w_dff_A_MrPJLRpt8_0),.din(w_dff_A_aU2zvkL33_0),.clk(gclk));
	jdff dff_A_MrPJLRpt8_0(.dout(w_dff_A_QTOLHuFS9_0),.din(w_dff_A_MrPJLRpt8_0),.clk(gclk));
	jdff dff_A_QTOLHuFS9_0(.dout(G752),.din(w_dff_A_QTOLHuFS9_0),.clk(gclk));
	jdff dff_A_SmweK2rc4_2(.dout(w_dff_A_kCf0gnem7_0),.din(w_dff_A_SmweK2rc4_2),.clk(gclk));
	jdff dff_A_kCf0gnem7_0(.dout(w_dff_A_mncjqRI36_0),.din(w_dff_A_kCf0gnem7_0),.clk(gclk));
	jdff dff_A_mncjqRI36_0(.dout(w_dff_A_J6oIVXMM4_0),.din(w_dff_A_mncjqRI36_0),.clk(gclk));
	jdff dff_A_J6oIVXMM4_0(.dout(w_dff_A_wv7nFki81_0),.din(w_dff_A_J6oIVXMM4_0),.clk(gclk));
	jdff dff_A_wv7nFki81_0(.dout(w_dff_A_D4g7LYgi0_0),.din(w_dff_A_wv7nFki81_0),.clk(gclk));
	jdff dff_A_D4g7LYgi0_0(.dout(w_dff_A_XyJRopmA2_0),.din(w_dff_A_D4g7LYgi0_0),.clk(gclk));
	jdff dff_A_XyJRopmA2_0(.dout(w_dff_A_7oUpz2pl4_0),.din(w_dff_A_XyJRopmA2_0),.clk(gclk));
	jdff dff_A_7oUpz2pl4_0(.dout(w_dff_A_11VyRUfz4_0),.din(w_dff_A_7oUpz2pl4_0),.clk(gclk));
	jdff dff_A_11VyRUfz4_0(.dout(w_dff_A_vNTKL5wL6_0),.din(w_dff_A_11VyRUfz4_0),.clk(gclk));
	jdff dff_A_vNTKL5wL6_0(.dout(G757),.din(w_dff_A_vNTKL5wL6_0),.clk(gclk));
	jdff dff_A_19H5GxO39_2(.dout(w_dff_A_CkplTEF39_0),.din(w_dff_A_19H5GxO39_2),.clk(gclk));
	jdff dff_A_CkplTEF39_0(.dout(w_dff_A_VpQ895LF5_0),.din(w_dff_A_CkplTEF39_0),.clk(gclk));
	jdff dff_A_VpQ895LF5_0(.dout(w_dff_A_LPzmIaxm7_0),.din(w_dff_A_VpQ895LF5_0),.clk(gclk));
	jdff dff_A_LPzmIaxm7_0(.dout(w_dff_A_T98IUh9p5_0),.din(w_dff_A_LPzmIaxm7_0),.clk(gclk));
	jdff dff_A_T98IUh9p5_0(.dout(w_dff_A_kEinjJWw5_0),.din(w_dff_A_T98IUh9p5_0),.clk(gclk));
	jdff dff_A_kEinjJWw5_0(.dout(w_dff_A_p35Tfkqo2_0),.din(w_dff_A_kEinjJWw5_0),.clk(gclk));
	jdff dff_A_p35Tfkqo2_0(.dout(w_dff_A_CF4nTgrd4_0),.din(w_dff_A_p35Tfkqo2_0),.clk(gclk));
	jdff dff_A_CF4nTgrd4_0(.dout(w_dff_A_333Bxx204_0),.din(w_dff_A_CF4nTgrd4_0),.clk(gclk));
	jdff dff_A_333Bxx204_0(.dout(w_dff_A_vIISzsln7_0),.din(w_dff_A_333Bxx204_0),.clk(gclk));
	jdff dff_A_vIISzsln7_0(.dout(w_dff_A_vXSVgGy34_0),.din(w_dff_A_vIISzsln7_0),.clk(gclk));
	jdff dff_A_vXSVgGy34_0(.dout(G762),.din(w_dff_A_vXSVgGy34_0),.clk(gclk));
	jdff dff_A_pYaVT0Rd8_2(.dout(w_dff_A_Pf47elGq7_0),.din(w_dff_A_pYaVT0Rd8_2),.clk(gclk));
	jdff dff_A_Pf47elGq7_0(.dout(w_dff_A_Cq73wuwD4_0),.din(w_dff_A_Pf47elGq7_0),.clk(gclk));
	jdff dff_A_Cq73wuwD4_0(.dout(w_dff_A_gJojppiQ8_0),.din(w_dff_A_Cq73wuwD4_0),.clk(gclk));
	jdff dff_A_gJojppiQ8_0(.dout(w_dff_A_RbW9zctz4_0),.din(w_dff_A_gJojppiQ8_0),.clk(gclk));
	jdff dff_A_RbW9zctz4_0(.dout(w_dff_A_6l2Ydi907_0),.din(w_dff_A_RbW9zctz4_0),.clk(gclk));
	jdff dff_A_6l2Ydi907_0(.dout(w_dff_A_05xG1v6s4_0),.din(w_dff_A_6l2Ydi907_0),.clk(gclk));
	jdff dff_A_05xG1v6s4_0(.dout(G787),.din(w_dff_A_05xG1v6s4_0),.clk(gclk));
	jdff dff_A_zWQ5oN7u7_2(.dout(w_dff_A_kZqLK9Oe2_0),.din(w_dff_A_zWQ5oN7u7_2),.clk(gclk));
	jdff dff_A_kZqLK9Oe2_0(.dout(w_dff_A_RrjdQ1Ie4_0),.din(w_dff_A_kZqLK9Oe2_0),.clk(gclk));
	jdff dff_A_RrjdQ1Ie4_0(.dout(w_dff_A_f81B8eNJ3_0),.din(w_dff_A_RrjdQ1Ie4_0),.clk(gclk));
	jdff dff_A_f81B8eNJ3_0(.dout(w_dff_A_Xjvw3LUK6_0),.din(w_dff_A_f81B8eNJ3_0),.clk(gclk));
	jdff dff_A_Xjvw3LUK6_0(.dout(w_dff_A_0DkL6X2v5_0),.din(w_dff_A_Xjvw3LUK6_0),.clk(gclk));
	jdff dff_A_0DkL6X2v5_0(.dout(w_dff_A_UHprJJi11_0),.din(w_dff_A_0DkL6X2v5_0),.clk(gclk));
	jdff dff_A_UHprJJi11_0(.dout(w_dff_A_bZ7fGTv52_0),.din(w_dff_A_UHprJJi11_0),.clk(gclk));
	jdff dff_A_bZ7fGTv52_0(.dout(w_dff_A_cxwBHQIU5_0),.din(w_dff_A_bZ7fGTv52_0),.clk(gclk));
	jdff dff_A_cxwBHQIU5_0(.dout(G792),.din(w_dff_A_cxwBHQIU5_0),.clk(gclk));
	jdff dff_A_3Phyc5ei6_2(.dout(w_dff_A_fbbGPwTf2_0),.din(w_dff_A_3Phyc5ei6_2),.clk(gclk));
	jdff dff_A_fbbGPwTf2_0(.dout(w_dff_A_OSuH9g8x7_0),.din(w_dff_A_fbbGPwTf2_0),.clk(gclk));
	jdff dff_A_OSuH9g8x7_0(.dout(w_dff_A_Gv1QOu920_0),.din(w_dff_A_OSuH9g8x7_0),.clk(gclk));
	jdff dff_A_Gv1QOu920_0(.dout(w_dff_A_ZTMCKfLC4_0),.din(w_dff_A_Gv1QOu920_0),.clk(gclk));
	jdff dff_A_ZTMCKfLC4_0(.dout(w_dff_A_N6lVp1zz8_0),.din(w_dff_A_ZTMCKfLC4_0),.clk(gclk));
	jdff dff_A_N6lVp1zz8_0(.dout(w_dff_A_ezaOVLRV0_0),.din(w_dff_A_N6lVp1zz8_0),.clk(gclk));
	jdff dff_A_ezaOVLRV0_0(.dout(w_dff_A_bmrWEQNl7_0),.din(w_dff_A_ezaOVLRV0_0),.clk(gclk));
	jdff dff_A_bmrWEQNl7_0(.dout(w_dff_A_xHk89ZmV2_0),.din(w_dff_A_bmrWEQNl7_0),.clk(gclk));
	jdff dff_A_xHk89ZmV2_0(.dout(w_dff_A_i4XbFAfI4_0),.din(w_dff_A_xHk89ZmV2_0),.clk(gclk));
	jdff dff_A_i4XbFAfI4_0(.dout(G797),.din(w_dff_A_i4XbFAfI4_0),.clk(gclk));
	jdff dff_A_kR71S9B18_2(.dout(w_dff_A_aCA6XL235_0),.din(w_dff_A_kR71S9B18_2),.clk(gclk));
	jdff dff_A_aCA6XL235_0(.dout(w_dff_A_TakHbnji0_0),.din(w_dff_A_aCA6XL235_0),.clk(gclk));
	jdff dff_A_TakHbnji0_0(.dout(w_dff_A_QJtBWF2X1_0),.din(w_dff_A_TakHbnji0_0),.clk(gclk));
	jdff dff_A_QJtBWF2X1_0(.dout(w_dff_A_KW4ljHCu3_0),.din(w_dff_A_QJtBWF2X1_0),.clk(gclk));
	jdff dff_A_KW4ljHCu3_0(.dout(w_dff_A_Ru72osg75_0),.din(w_dff_A_KW4ljHCu3_0),.clk(gclk));
	jdff dff_A_Ru72osg75_0(.dout(w_dff_A_IenheodB6_0),.din(w_dff_A_Ru72osg75_0),.clk(gclk));
	jdff dff_A_IenheodB6_0(.dout(w_dff_A_MCNNZQST9_0),.din(w_dff_A_IenheodB6_0),.clk(gclk));
	jdff dff_A_MCNNZQST9_0(.dout(w_dff_A_Lwtw3oUA6_0),.din(w_dff_A_MCNNZQST9_0),.clk(gclk));
	jdff dff_A_Lwtw3oUA6_0(.dout(w_dff_A_vBUBildu3_0),.din(w_dff_A_Lwtw3oUA6_0),.clk(gclk));
	jdff dff_A_vBUBildu3_0(.dout(w_dff_A_T5KTvmcx1_0),.din(w_dff_A_vBUBildu3_0),.clk(gclk));
	jdff dff_A_T5KTvmcx1_0(.dout(G802),.din(w_dff_A_T5KTvmcx1_0),.clk(gclk));
	jdff dff_A_K4P7N6hP0_2(.dout(w_dff_A_EMuOqUc83_0),.din(w_dff_A_K4P7N6hP0_2),.clk(gclk));
	jdff dff_A_EMuOqUc83_0(.dout(w_dff_A_I0icv16C9_0),.din(w_dff_A_EMuOqUc83_0),.clk(gclk));
	jdff dff_A_I0icv16C9_0(.dout(w_dff_A_AqOhtOe31_0),.din(w_dff_A_I0icv16C9_0),.clk(gclk));
	jdff dff_A_AqOhtOe31_0(.dout(w_dff_A_rRZTnKA65_0),.din(w_dff_A_AqOhtOe31_0),.clk(gclk));
	jdff dff_A_rRZTnKA65_0(.dout(w_dff_A_AkyEd3kP8_0),.din(w_dff_A_rRZTnKA65_0),.clk(gclk));
	jdff dff_A_AkyEd3kP8_0(.dout(G642),.din(w_dff_A_AkyEd3kP8_0),.clk(gclk));
	jdff dff_A_ezoq8C9i9_2(.dout(w_dff_A_r7ofSOrF0_0),.din(w_dff_A_ezoq8C9i9_2),.clk(gclk));
	jdff dff_A_r7ofSOrF0_0(.dout(w_dff_A_JfKnqpVd0_0),.din(w_dff_A_r7ofSOrF0_0),.clk(gclk));
	jdff dff_A_JfKnqpVd0_0(.dout(w_dff_A_gkw2YFHw9_0),.din(w_dff_A_JfKnqpVd0_0),.clk(gclk));
	jdff dff_A_gkw2YFHw9_0(.dout(w_dff_A_HwHOl2M93_0),.din(w_dff_A_gkw2YFHw9_0),.clk(gclk));
	jdff dff_A_HwHOl2M93_0(.dout(w_dff_A_8bQOTEfo0_0),.din(w_dff_A_HwHOl2M93_0),.clk(gclk));
	jdff dff_A_8bQOTEfo0_0(.dout(w_dff_A_taEuKB0R6_0),.din(w_dff_A_8bQOTEfo0_0),.clk(gclk));
	jdff dff_A_taEuKB0R6_0(.dout(w_dff_A_w2qqhGHj4_0),.din(w_dff_A_taEuKB0R6_0),.clk(gclk));
	jdff dff_A_w2qqhGHj4_0(.dout(w_dff_A_8Xgfz7I19_0),.din(w_dff_A_w2qqhGHj4_0),.clk(gclk));
	jdff dff_A_8Xgfz7I19_0(.dout(w_dff_A_3St8Wg039_0),.din(w_dff_A_8Xgfz7I19_0),.clk(gclk));
	jdff dff_A_3St8Wg039_0(.dout(G664),.din(w_dff_A_3St8Wg039_0),.clk(gclk));
	jdff dff_A_gnv61TFV1_2(.dout(w_dff_A_mMfZiepW4_0),.din(w_dff_A_gnv61TFV1_2),.clk(gclk));
	jdff dff_A_mMfZiepW4_0(.dout(w_dff_A_CkU8mcFC0_0),.din(w_dff_A_mMfZiepW4_0),.clk(gclk));
	jdff dff_A_CkU8mcFC0_0(.dout(w_dff_A_9SL0YjeN3_0),.din(w_dff_A_CkU8mcFC0_0),.clk(gclk));
	jdff dff_A_9SL0YjeN3_0(.dout(w_dff_A_lH1SOfWF7_0),.din(w_dff_A_9SL0YjeN3_0),.clk(gclk));
	jdff dff_A_lH1SOfWF7_0(.dout(w_dff_A_GkkDKFhC6_0),.din(w_dff_A_lH1SOfWF7_0),.clk(gclk));
	jdff dff_A_GkkDKFhC6_0(.dout(w_dff_A_ezHOAA2O4_0),.din(w_dff_A_GkkDKFhC6_0),.clk(gclk));
	jdff dff_A_ezHOAA2O4_0(.dout(w_dff_A_gC63kOGS8_0),.din(w_dff_A_ezHOAA2O4_0),.clk(gclk));
	jdff dff_A_gC63kOGS8_0(.dout(w_dff_A_QTUfGkKg6_0),.din(w_dff_A_gC63kOGS8_0),.clk(gclk));
	jdff dff_A_QTUfGkKg6_0(.dout(G667),.din(w_dff_A_QTUfGkKg6_0),.clk(gclk));
	jdff dff_A_rJmF9iXA4_2(.dout(w_dff_A_wuCNB4UR3_0),.din(w_dff_A_rJmF9iXA4_2),.clk(gclk));
	jdff dff_A_wuCNB4UR3_0(.dout(w_dff_A_CUGWhDlB8_0),.din(w_dff_A_wuCNB4UR3_0),.clk(gclk));
	jdff dff_A_CUGWhDlB8_0(.dout(w_dff_A_j4GLjSqq9_0),.din(w_dff_A_CUGWhDlB8_0),.clk(gclk));
	jdff dff_A_j4GLjSqq9_0(.dout(w_dff_A_eva3bVmB9_0),.din(w_dff_A_j4GLjSqq9_0),.clk(gclk));
	jdff dff_A_eva3bVmB9_0(.dout(w_dff_A_jRtr63dN5_0),.din(w_dff_A_eva3bVmB9_0),.clk(gclk));
	jdff dff_A_jRtr63dN5_0(.dout(w_dff_A_IpUQfIyO6_0),.din(w_dff_A_jRtr63dN5_0),.clk(gclk));
	jdff dff_A_IpUQfIyO6_0(.dout(w_dff_A_roGkLfMO2_0),.din(w_dff_A_IpUQfIyO6_0),.clk(gclk));
	jdff dff_A_roGkLfMO2_0(.dout(G670),.din(w_dff_A_roGkLfMO2_0),.clk(gclk));
	jdff dff_A_Ox1Xngjw7_2(.dout(w_dff_A_CI8vtukZ7_0),.din(w_dff_A_Ox1Xngjw7_2),.clk(gclk));
	jdff dff_A_CI8vtukZ7_0(.dout(w_dff_A_fSKr5kwp3_0),.din(w_dff_A_CI8vtukZ7_0),.clk(gclk));
	jdff dff_A_fSKr5kwp3_0(.dout(w_dff_A_LVci0KQs4_0),.din(w_dff_A_fSKr5kwp3_0),.clk(gclk));
	jdff dff_A_LVci0KQs4_0(.dout(w_dff_A_EFKPCJSO0_0),.din(w_dff_A_LVci0KQs4_0),.clk(gclk));
	jdff dff_A_EFKPCJSO0_0(.dout(w_dff_A_8A0phuLi9_0),.din(w_dff_A_EFKPCJSO0_0),.clk(gclk));
	jdff dff_A_8A0phuLi9_0(.dout(G676),.din(w_dff_A_8A0phuLi9_0),.clk(gclk));
	jdff dff_A_McN35ANS3_2(.dout(w_dff_A_BosRwV852_0),.din(w_dff_A_McN35ANS3_2),.clk(gclk));
	jdff dff_A_BosRwV852_0(.dout(w_dff_A_qlzsTmU16_0),.din(w_dff_A_BosRwV852_0),.clk(gclk));
	jdff dff_A_qlzsTmU16_0(.dout(w_dff_A_W79NsMZG5_0),.din(w_dff_A_qlzsTmU16_0),.clk(gclk));
	jdff dff_A_W79NsMZG5_0(.dout(w_dff_A_6txG9rdT9_0),.din(w_dff_A_W79NsMZG5_0),.clk(gclk));
	jdff dff_A_6txG9rdT9_0(.dout(w_dff_A_kzKdnUt37_0),.din(w_dff_A_6txG9rdT9_0),.clk(gclk));
	jdff dff_A_kzKdnUt37_0(.dout(w_dff_A_2NJkJHVQ0_0),.din(w_dff_A_kzKdnUt37_0),.clk(gclk));
	jdff dff_A_2NJkJHVQ0_0(.dout(w_dff_A_qWXZYGSi6_0),.din(w_dff_A_2NJkJHVQ0_0),.clk(gclk));
	jdff dff_A_qWXZYGSi6_0(.dout(w_dff_A_o0iUeAoK2_0),.din(w_dff_A_qWXZYGSi6_0),.clk(gclk));
	jdff dff_A_o0iUeAoK2_0(.dout(w_dff_A_5qvAay5z2_0),.din(w_dff_A_o0iUeAoK2_0),.clk(gclk));
	jdff dff_A_5qvAay5z2_0(.dout(G696),.din(w_dff_A_5qvAay5z2_0),.clk(gclk));
	jdff dff_A_EEV2iFkR2_2(.dout(w_dff_A_t7TnUSKN7_0),.din(w_dff_A_EEV2iFkR2_2),.clk(gclk));
	jdff dff_A_t7TnUSKN7_0(.dout(w_dff_A_1fQoPR9M5_0),.din(w_dff_A_t7TnUSKN7_0),.clk(gclk));
	jdff dff_A_1fQoPR9M5_0(.dout(w_dff_A_fiJjTg9N5_0),.din(w_dff_A_1fQoPR9M5_0),.clk(gclk));
	jdff dff_A_fiJjTg9N5_0(.dout(w_dff_A_zW4POg2M2_0),.din(w_dff_A_fiJjTg9N5_0),.clk(gclk));
	jdff dff_A_zW4POg2M2_0(.dout(w_dff_A_U8jJeBae8_0),.din(w_dff_A_zW4POg2M2_0),.clk(gclk));
	jdff dff_A_U8jJeBae8_0(.dout(w_dff_A_mC2kIqIz9_0),.din(w_dff_A_U8jJeBae8_0),.clk(gclk));
	jdff dff_A_mC2kIqIz9_0(.dout(w_dff_A_k1mwG7fn4_0),.din(w_dff_A_mC2kIqIz9_0),.clk(gclk));
	jdff dff_A_k1mwG7fn4_0(.dout(w_dff_A_hP4eKqU42_0),.din(w_dff_A_k1mwG7fn4_0),.clk(gclk));
	jdff dff_A_hP4eKqU42_0(.dout(G699),.din(w_dff_A_hP4eKqU42_0),.clk(gclk));
	jdff dff_A_x965G86B7_2(.dout(w_dff_A_zXf9E0Og1_0),.din(w_dff_A_x965G86B7_2),.clk(gclk));
	jdff dff_A_zXf9E0Og1_0(.dout(w_dff_A_70xlT3x62_0),.din(w_dff_A_zXf9E0Og1_0),.clk(gclk));
	jdff dff_A_70xlT3x62_0(.dout(w_dff_A_Lm8y4DcO9_0),.din(w_dff_A_70xlT3x62_0),.clk(gclk));
	jdff dff_A_Lm8y4DcO9_0(.dout(w_dff_A_a06eyMM67_0),.din(w_dff_A_Lm8y4DcO9_0),.clk(gclk));
	jdff dff_A_a06eyMM67_0(.dout(w_dff_A_eeeVtZlV6_0),.din(w_dff_A_a06eyMM67_0),.clk(gclk));
	jdff dff_A_eeeVtZlV6_0(.dout(w_dff_A_3r2jDFcY2_0),.din(w_dff_A_eeeVtZlV6_0),.clk(gclk));
	jdff dff_A_3r2jDFcY2_0(.dout(w_dff_A_w55egnzk1_0),.din(w_dff_A_3r2jDFcY2_0),.clk(gclk));
	jdff dff_A_w55egnzk1_0(.dout(G702),.din(w_dff_A_w55egnzk1_0),.clk(gclk));
	jdff dff_A_YIjMVBcl3_2(.dout(w_dff_A_YDP4YiCG6_0),.din(w_dff_A_YIjMVBcl3_2),.clk(gclk));
	jdff dff_A_YDP4YiCG6_0(.dout(w_dff_A_BX6lASSb2_0),.din(w_dff_A_YDP4YiCG6_0),.clk(gclk));
	jdff dff_A_BX6lASSb2_0(.dout(w_dff_A_K6m8maJW8_0),.din(w_dff_A_BX6lASSb2_0),.clk(gclk));
	jdff dff_A_K6m8maJW8_0(.dout(w_dff_A_KrXez6WB0_0),.din(w_dff_A_K6m8maJW8_0),.clk(gclk));
	jdff dff_A_KrXez6WB0_0(.dout(G818),.din(w_dff_A_KrXez6WB0_0),.clk(gclk));
	jdff dff_A_VUuDR6GP3_2(.dout(w_dff_A_2UUTflwp7_0),.din(w_dff_A_VUuDR6GP3_2),.clk(gclk));
	jdff dff_A_2UUTflwp7_0(.dout(w_dff_A_AqNe3o8C0_0),.din(w_dff_A_2UUTflwp7_0),.clk(gclk));
	jdff dff_A_AqNe3o8C0_0(.dout(w_dff_A_cJHUWzDP6_0),.din(w_dff_A_AqNe3o8C0_0),.clk(gclk));
	jdff dff_A_cJHUWzDP6_0(.dout(w_dff_A_ZQGg0kSb7_0),.din(w_dff_A_cJHUWzDP6_0),.clk(gclk));
	jdff dff_A_ZQGg0kSb7_0(.dout(w_dff_A_UJdi8eDm4_0),.din(w_dff_A_ZQGg0kSb7_0),.clk(gclk));
	jdff dff_A_UJdi8eDm4_0(.dout(w_dff_A_cRGRjQb90_0),.din(w_dff_A_UJdi8eDm4_0),.clk(gclk));
	jdff dff_A_cRGRjQb90_0(.dout(w_dff_A_jx2THHHv0_0),.din(w_dff_A_cRGRjQb90_0),.clk(gclk));
	jdff dff_A_jx2THHHv0_0(.dout(w_dff_A_55bRIRtq1_0),.din(w_dff_A_jx2THHHv0_0),.clk(gclk));
	jdff dff_A_55bRIRtq1_0(.dout(G813),.din(w_dff_A_55bRIRtq1_0),.clk(gclk));
	jdff dff_A_dRifuz8t7_1(.dout(w_dff_A_Lj2wljKi8_0),.din(w_dff_A_dRifuz8t7_1),.clk(gclk));
	jdff dff_A_Lj2wljKi8_0(.dout(w_dff_A_n9v9kLba2_0),.din(w_dff_A_Lj2wljKi8_0),.clk(gclk));
	jdff dff_A_n9v9kLba2_0(.dout(w_dff_A_L1aXTwpM2_0),.din(w_dff_A_n9v9kLba2_0),.clk(gclk));
	jdff dff_A_L1aXTwpM2_0(.dout(w_dff_A_5hZJmb488_0),.din(w_dff_A_L1aXTwpM2_0),.clk(gclk));
	jdff dff_A_5hZJmb488_0(.dout(G824),.din(w_dff_A_5hZJmb488_0),.clk(gclk));
	jdff dff_A_8Pa9YStv0_1(.dout(w_dff_A_8FDlU7Z94_0),.din(w_dff_A_8Pa9YStv0_1),.clk(gclk));
	jdff dff_A_8FDlU7Z94_0(.dout(w_dff_A_YA723v3U1_0),.din(w_dff_A_8FDlU7Z94_0),.clk(gclk));
	jdff dff_A_YA723v3U1_0(.dout(w_dff_A_dKnmV6xp3_0),.din(w_dff_A_YA723v3U1_0),.clk(gclk));
	jdff dff_A_dKnmV6xp3_0(.dout(w_dff_A_4f4smzWv7_0),.din(w_dff_A_dKnmV6xp3_0),.clk(gclk));
	jdff dff_A_4f4smzWv7_0(.dout(w_dff_A_r2WU4mxa7_0),.din(w_dff_A_4f4smzWv7_0),.clk(gclk));
	jdff dff_A_r2WU4mxa7_0(.dout(w_dff_A_0eCZVfks5_0),.din(w_dff_A_r2WU4mxa7_0),.clk(gclk));
	jdff dff_A_0eCZVfks5_0(.dout(w_dff_A_unZc6zDF5_0),.din(w_dff_A_0eCZVfks5_0),.clk(gclk));
	jdff dff_A_unZc6zDF5_0(.dout(G826),.din(w_dff_A_unZc6zDF5_0),.clk(gclk));
	jdff dff_A_WWL5M9oO4_1(.dout(w_dff_A_MwQ62wHi0_0),.din(w_dff_A_WWL5M9oO4_1),.clk(gclk));
	jdff dff_A_MwQ62wHi0_0(.dout(w_dff_A_bXXqA2gj0_0),.din(w_dff_A_MwQ62wHi0_0),.clk(gclk));
	jdff dff_A_bXXqA2gj0_0(.dout(w_dff_A_vQzWbjcD8_0),.din(w_dff_A_bXXqA2gj0_0),.clk(gclk));
	jdff dff_A_vQzWbjcD8_0(.dout(w_dff_A_89pAjEOo2_0),.din(w_dff_A_vQzWbjcD8_0),.clk(gclk));
	jdff dff_A_89pAjEOo2_0(.dout(w_dff_A_Z6Md5XyQ1_0),.din(w_dff_A_89pAjEOo2_0),.clk(gclk));
	jdff dff_A_Z6Md5XyQ1_0(.dout(w_dff_A_V6uqVzyG3_0),.din(w_dff_A_Z6Md5XyQ1_0),.clk(gclk));
	jdff dff_A_V6uqVzyG3_0(.dout(w_dff_A_L7SR8ykS2_0),.din(w_dff_A_V6uqVzyG3_0),.clk(gclk));
	jdff dff_A_L7SR8ykS2_0(.dout(G828),.din(w_dff_A_L7SR8ykS2_0),.clk(gclk));
	jdff dff_A_mLyNlAgr2_1(.dout(w_dff_A_mraoG5du0_0),.din(w_dff_A_mLyNlAgr2_1),.clk(gclk));
	jdff dff_A_mraoG5du0_0(.dout(w_dff_A_YEawgPrx4_0),.din(w_dff_A_mraoG5du0_0),.clk(gclk));
	jdff dff_A_YEawgPrx4_0(.dout(w_dff_A_B7gsoJio3_0),.din(w_dff_A_YEawgPrx4_0),.clk(gclk));
	jdff dff_A_B7gsoJio3_0(.dout(w_dff_A_uV8eFwMf2_0),.din(w_dff_A_B7gsoJio3_0),.clk(gclk));
	jdff dff_A_uV8eFwMf2_0(.dout(w_dff_A_nGiSCrPh2_0),.din(w_dff_A_uV8eFwMf2_0),.clk(gclk));
	jdff dff_A_nGiSCrPh2_0(.dout(w_dff_A_8Ynurn2G0_0),.din(w_dff_A_nGiSCrPh2_0),.clk(gclk));
	jdff dff_A_8Ynurn2G0_0(.dout(w_dff_A_gxQ3cpsS0_0),.din(w_dff_A_8Ynurn2G0_0),.clk(gclk));
	jdff dff_A_gxQ3cpsS0_0(.dout(w_dff_A_aljJRhok0_0),.din(w_dff_A_gxQ3cpsS0_0),.clk(gclk));
	jdff dff_A_aljJRhok0_0(.dout(G830),.din(w_dff_A_aljJRhok0_0),.clk(gclk));
	jdff dff_A_dWiR3lKc9_2(.dout(w_dff_A_REBnqDrA5_0),.din(w_dff_A_dWiR3lKc9_2),.clk(gclk));
	jdff dff_A_REBnqDrA5_0(.dout(w_dff_A_sKBWvyPh9_0),.din(w_dff_A_REBnqDrA5_0),.clk(gclk));
	jdff dff_A_sKBWvyPh9_0(.dout(w_dff_A_5ToOHbWm8_0),.din(w_dff_A_sKBWvyPh9_0),.clk(gclk));
	jdff dff_A_5ToOHbWm8_0(.dout(w_dff_A_LoIhxFRI9_0),.din(w_dff_A_5ToOHbWm8_0),.clk(gclk));
	jdff dff_A_LoIhxFRI9_0(.dout(w_dff_A_2HMndqNF9_0),.din(w_dff_A_LoIhxFRI9_0),.clk(gclk));
	jdff dff_A_2HMndqNF9_0(.dout(w_dff_A_WS56Qo9Z5_0),.din(w_dff_A_2HMndqNF9_0),.clk(gclk));
	jdff dff_A_WS56Qo9Z5_0(.dout(w_dff_A_6UAEFGew6_0),.din(w_dff_A_WS56Qo9Z5_0),.clk(gclk));
	jdff dff_A_6UAEFGew6_0(.dout(w_dff_A_SYj6CJqL4_0),.din(w_dff_A_6UAEFGew6_0),.clk(gclk));
	jdff dff_A_SYj6CJqL4_0(.dout(w_dff_A_hV5cQzcV5_0),.din(w_dff_A_SYj6CJqL4_0),.clk(gclk));
	jdff dff_A_hV5cQzcV5_0(.dout(w_dff_A_eyz1tPcM8_0),.din(w_dff_A_hV5cQzcV5_0),.clk(gclk));
	jdff dff_A_eyz1tPcM8_0(.dout(w_dff_A_oe773Z964_0),.din(w_dff_A_eyz1tPcM8_0),.clk(gclk));
	jdff dff_A_oe773Z964_0(.dout(w_dff_A_HBm8Pqso5_0),.din(w_dff_A_oe773Z964_0),.clk(gclk));
	jdff dff_A_HBm8Pqso5_0(.dout(w_dff_A_WPtnuktD0_0),.din(w_dff_A_HBm8Pqso5_0),.clk(gclk));
	jdff dff_A_WPtnuktD0_0(.dout(w_dff_A_3ikstzRv4_0),.din(w_dff_A_WPtnuktD0_0),.clk(gclk));
	jdff dff_A_3ikstzRv4_0(.dout(w_dff_A_5gC9Os1p4_0),.din(w_dff_A_3ikstzRv4_0),.clk(gclk));
	jdff dff_A_5gC9Os1p4_0(.dout(G854),.din(w_dff_A_5gC9Os1p4_0),.clk(gclk));
	jdff dff_A_YbUu0rt76_1(.dout(w_dff_A_uMJxHwHR9_0),.din(w_dff_A_YbUu0rt76_1),.clk(gclk));
	jdff dff_A_uMJxHwHR9_0(.dout(w_dff_A_ELEPugdY3_0),.din(w_dff_A_uMJxHwHR9_0),.clk(gclk));
	jdff dff_A_ELEPugdY3_0(.dout(w_dff_A_Cn3iv0w64_0),.din(w_dff_A_ELEPugdY3_0),.clk(gclk));
	jdff dff_A_Cn3iv0w64_0(.dout(G863),.din(w_dff_A_Cn3iv0w64_0),.clk(gclk));
	jdff dff_A_jFPW27Js2_1(.dout(w_dff_A_XD6j3chI0_0),.din(w_dff_A_jFPW27Js2_1),.clk(gclk));
	jdff dff_A_XD6j3chI0_0(.dout(w_dff_A_z6FqgfEj7_0),.din(w_dff_A_XD6j3chI0_0),.clk(gclk));
	jdff dff_A_z6FqgfEj7_0(.dout(w_dff_A_LFRXAEMs0_0),.din(w_dff_A_z6FqgfEj7_0),.clk(gclk));
	jdff dff_A_LFRXAEMs0_0(.dout(w_dff_A_EMv9EHTg6_0),.din(w_dff_A_LFRXAEMs0_0),.clk(gclk));
	jdff dff_A_EMv9EHTg6_0(.dout(G865),.din(w_dff_A_EMv9EHTg6_0),.clk(gclk));
	jdff dff_A_yZxRu1CP2_1(.dout(w_dff_A_t0UT0z536_0),.din(w_dff_A_yZxRu1CP2_1),.clk(gclk));
	jdff dff_A_t0UT0z536_0(.dout(w_dff_A_wyGvadyG9_0),.din(w_dff_A_t0UT0z536_0),.clk(gclk));
	jdff dff_A_wyGvadyG9_0(.dout(w_dff_A_8R4oR8H47_0),.din(w_dff_A_wyGvadyG9_0),.clk(gclk));
	jdff dff_A_8R4oR8H47_0(.dout(w_dff_A_JPMgzgEx2_0),.din(w_dff_A_8R4oR8H47_0),.clk(gclk));
	jdff dff_A_JPMgzgEx2_0(.dout(w_dff_A_Q7zqQz1Q8_0),.din(w_dff_A_JPMgzgEx2_0),.clk(gclk));
	jdff dff_A_Q7zqQz1Q8_0(.dout(w_dff_A_CR2Xnq2k7_0),.din(w_dff_A_Q7zqQz1Q8_0),.clk(gclk));
	jdff dff_A_CR2Xnq2k7_0(.dout(G867),.din(w_dff_A_CR2Xnq2k7_0),.clk(gclk));
	jdff dff_A_3kPjIFex3_1(.dout(w_dff_A_asAFbCei9_0),.din(w_dff_A_3kPjIFex3_1),.clk(gclk));
	jdff dff_A_asAFbCei9_0(.dout(w_dff_A_cCdNDXPH6_0),.din(w_dff_A_asAFbCei9_0),.clk(gclk));
	jdff dff_A_cCdNDXPH6_0(.dout(w_dff_A_XvoRUMQB7_0),.din(w_dff_A_cCdNDXPH6_0),.clk(gclk));
	jdff dff_A_XvoRUMQB7_0(.dout(w_dff_A_XErBjIMI5_0),.din(w_dff_A_XvoRUMQB7_0),.clk(gclk));
	jdff dff_A_XErBjIMI5_0(.dout(w_dff_A_LUW5uCGe2_0),.din(w_dff_A_XErBjIMI5_0),.clk(gclk));
	jdff dff_A_LUW5uCGe2_0(.dout(w_dff_A_c6BudVkf4_0),.din(w_dff_A_LUW5uCGe2_0),.clk(gclk));
	jdff dff_A_c6BudVkf4_0(.dout(w_dff_A_c349SEMu3_0),.din(w_dff_A_c6BudVkf4_0),.clk(gclk));
	jdff dff_A_c349SEMu3_0(.dout(G869),.din(w_dff_A_c349SEMu3_0),.clk(gclk));
	jdff dff_A_nWpQUXif7_2(.dout(w_dff_A_qnQCP2FW6_0),.din(w_dff_A_nWpQUXif7_2),.clk(gclk));
	jdff dff_A_qnQCP2FW6_0(.dout(w_dff_A_w46jqcqI5_0),.din(w_dff_A_qnQCP2FW6_0),.clk(gclk));
	jdff dff_A_w46jqcqI5_0(.dout(G712),.din(w_dff_A_w46jqcqI5_0),.clk(gclk));
	jdff dff_A_wC6dLpOY8_2(.dout(w_dff_A_DJoEsS8a5_0),.din(w_dff_A_wC6dLpOY8_2),.clk(gclk));
	jdff dff_A_DJoEsS8a5_0(.dout(w_dff_A_ZDnS8Dex4_0),.din(w_dff_A_DJoEsS8a5_0),.clk(gclk));
	jdff dff_A_ZDnS8Dex4_0(.dout(G727),.din(w_dff_A_ZDnS8Dex4_0),.clk(gclk));
	jdff dff_A_aOg13yvN6_2(.dout(w_dff_A_BoKCrHaW0_0),.din(w_dff_A_aOg13yvN6_2),.clk(gclk));
	jdff dff_A_BoKCrHaW0_0(.dout(w_dff_A_iJi8hbqm4_0),.din(w_dff_A_BoKCrHaW0_0),.clk(gclk));
	jdff dff_A_iJi8hbqm4_0(.dout(w_dff_A_jjn7m34c5_0),.din(w_dff_A_iJi8hbqm4_0),.clk(gclk));
	jdff dff_A_jjn7m34c5_0(.dout(G732),.din(w_dff_A_jjn7m34c5_0),.clk(gclk));
	jdff dff_A_Gz7SUmwg3_2(.dout(w_dff_A_vR67JDpJ5_0),.din(w_dff_A_Gz7SUmwg3_2),.clk(gclk));
	jdff dff_A_vR67JDpJ5_0(.dout(w_dff_A_gKNKnbk48_0),.din(w_dff_A_vR67JDpJ5_0),.clk(gclk));
	jdff dff_A_gKNKnbk48_0(.dout(w_dff_A_WOszV7J96_0),.din(w_dff_A_gKNKnbk48_0),.clk(gclk));
	jdff dff_A_WOszV7J96_0(.dout(G737),.din(w_dff_A_WOszV7J96_0),.clk(gclk));
	jdff dff_A_Kj9RkwBZ2_2(.dout(w_dff_A_YAt4ZZqV2_0),.din(w_dff_A_Kj9RkwBZ2_2),.clk(gclk));
	jdff dff_A_YAt4ZZqV2_0(.dout(w_dff_A_en51KzfX7_0),.din(w_dff_A_YAt4ZZqV2_0),.clk(gclk));
	jdff dff_A_en51KzfX7_0(.dout(w_dff_A_5aBGWT594_0),.din(w_dff_A_en51KzfX7_0),.clk(gclk));
	jdff dff_A_5aBGWT594_0(.dout(w_dff_A_SC7UKnfq8_0),.din(w_dff_A_5aBGWT594_0),.clk(gclk));
	jdff dff_A_SC7UKnfq8_0(.dout(G742),.din(w_dff_A_SC7UKnfq8_0),.clk(gclk));
	jdff dff_A_r913b9Tx0_2(.dout(w_dff_A_MyLslFcV2_0),.din(w_dff_A_r913b9Tx0_2),.clk(gclk));
	jdff dff_A_MyLslFcV2_0(.dout(w_dff_A_KyIDrp7O3_0),.din(w_dff_A_MyLslFcV2_0),.clk(gclk));
	jdff dff_A_KyIDrp7O3_0(.dout(w_dff_A_MUyDFMxZ5_0),.din(w_dff_A_KyIDrp7O3_0),.clk(gclk));
	jdff dff_A_MUyDFMxZ5_0(.dout(G772),.din(w_dff_A_MUyDFMxZ5_0),.clk(gclk));
	jdff dff_A_B7zzNCht4_2(.dout(w_dff_A_gzPPoZzQ1_0),.din(w_dff_A_B7zzNCht4_2),.clk(gclk));
	jdff dff_A_gzPPoZzQ1_0(.dout(w_dff_A_Pb2PdW7y6_0),.din(w_dff_A_gzPPoZzQ1_0),.clk(gclk));
	jdff dff_A_Pb2PdW7y6_0(.dout(w_dff_A_3L2PEZOQ6_0),.din(w_dff_A_Pb2PdW7y6_0),.clk(gclk));
	jdff dff_A_3L2PEZOQ6_0(.dout(G777),.din(w_dff_A_3L2PEZOQ6_0),.clk(gclk));
	jdff dff_A_zAFhLVgo8_2(.dout(w_dff_A_PHqc0E8t0_0),.din(w_dff_A_zAFhLVgo8_2),.clk(gclk));
	jdff dff_A_PHqc0E8t0_0(.dout(w_dff_A_qPJeZuC07_0),.din(w_dff_A_PHqc0E8t0_0),.clk(gclk));
	jdff dff_A_qPJeZuC07_0(.dout(w_dff_A_qmraD4Nd5_0),.din(w_dff_A_qPJeZuC07_0),.clk(gclk));
	jdff dff_A_qmraD4Nd5_0(.dout(w_dff_A_btpGjl9F0_0),.din(w_dff_A_qmraD4Nd5_0),.clk(gclk));
	jdff dff_A_btpGjl9F0_0(.dout(G782),.din(w_dff_A_btpGjl9F0_0),.clk(gclk));
	jdff dff_A_IHkscreG0_2(.dout(w_dff_A_vvc2VZZb5_0),.din(w_dff_A_IHkscreG0_2),.clk(gclk));
	jdff dff_A_vvc2VZZb5_0(.dout(w_dff_A_AcozqTrH7_0),.din(w_dff_A_vvc2VZZb5_0),.clk(gclk));
	jdff dff_A_AcozqTrH7_0(.dout(w_dff_A_Po0WJqnD9_0),.din(w_dff_A_AcozqTrH7_0),.clk(gclk));
	jdff dff_A_Po0WJqnD9_0(.dout(G645),.din(w_dff_A_Po0WJqnD9_0),.clk(gclk));
	jdff dff_A_waPH8W0z0_2(.dout(w_dff_A_W3CeAKtQ5_0),.din(w_dff_A_waPH8W0z0_2),.clk(gclk));
	jdff dff_A_W3CeAKtQ5_0(.dout(w_dff_A_8F4EYnfM6_0),.din(w_dff_A_W3CeAKtQ5_0),.clk(gclk));
	jdff dff_A_8F4EYnfM6_0(.dout(G648),.din(w_dff_A_8F4EYnfM6_0),.clk(gclk));
	jdff dff_A_Ma7drrNq3_2(.dout(w_dff_A_To0ayZgd9_0),.din(w_dff_A_Ma7drrNq3_2),.clk(gclk));
	jdff dff_A_To0ayZgd9_0(.dout(w_dff_A_4p4Wrc8s2_0),.din(w_dff_A_To0ayZgd9_0),.clk(gclk));
	jdff dff_A_4p4Wrc8s2_0(.dout(G651),.din(w_dff_A_4p4Wrc8s2_0),.clk(gclk));
	jdff dff_A_CSW3oR7E2_2(.dout(w_dff_A_ZApLNaRm5_0),.din(w_dff_A_CSW3oR7E2_2),.clk(gclk));
	jdff dff_A_ZApLNaRm5_0(.dout(G654),.din(w_dff_A_ZApLNaRm5_0),.clk(gclk));
	jdff dff_A_jCh5PqgI7_2(.dout(w_dff_A_LQ1RT4Xg3_0),.din(w_dff_A_jCh5PqgI7_2),.clk(gclk));
	jdff dff_A_LQ1RT4Xg3_0(.dout(w_dff_A_1TfznRbi4_0),.din(w_dff_A_LQ1RT4Xg3_0),.clk(gclk));
	jdff dff_A_1TfznRbi4_0(.dout(w_dff_A_yIsjDxSq4_0),.din(w_dff_A_1TfznRbi4_0),.clk(gclk));
	jdff dff_A_yIsjDxSq4_0(.dout(G679),.din(w_dff_A_yIsjDxSq4_0),.clk(gclk));
	jdff dff_A_QI9HYEpX5_2(.dout(w_dff_A_TD904Lgl4_0),.din(w_dff_A_QI9HYEpX5_2),.clk(gclk));
	jdff dff_A_TD904Lgl4_0(.dout(w_dff_A_6eNES9vT4_0),.din(w_dff_A_TD904Lgl4_0),.clk(gclk));
	jdff dff_A_6eNES9vT4_0(.dout(G682),.din(w_dff_A_6eNES9vT4_0),.clk(gclk));
	jdff dff_A_MbjnhRRh3_2(.dout(w_dff_A_qARrPKVs1_0),.din(w_dff_A_MbjnhRRh3_2),.clk(gclk));
	jdff dff_A_qARrPKVs1_0(.dout(w_dff_A_seMwHF2r9_0),.din(w_dff_A_qARrPKVs1_0),.clk(gclk));
	jdff dff_A_seMwHF2r9_0(.dout(G685),.din(w_dff_A_seMwHF2r9_0),.clk(gclk));
	jdff dff_A_j5GasjKW1_2(.dout(w_dff_A_rwYucOoo7_0),.din(w_dff_A_j5GasjKW1_2),.clk(gclk));
	jdff dff_A_rwYucOoo7_0(.dout(G688),.din(w_dff_A_rwYucOoo7_0),.clk(gclk));
	jdff dff_A_JuKIKgog1_2(.dout(w_dff_A_xoyA0ozh6_0),.din(w_dff_A_JuKIKgog1_2),.clk(gclk));
	jdff dff_A_xoyA0ozh6_0(.dout(w_dff_A_YZNLLjuP3_0),.din(w_dff_A_xoyA0ozh6_0),.clk(gclk));
	jdff dff_A_YZNLLjuP3_0(.dout(w_dff_A_novSlxr97_0),.din(w_dff_A_YZNLLjuP3_0),.clk(gclk));
	jdff dff_A_novSlxr97_0(.dout(G843),.din(w_dff_A_novSlxr97_0),.clk(gclk));
	jdff dff_A_fExTKHZC7_2(.dout(w_dff_A_udOtkEGA8_0),.din(w_dff_A_fExTKHZC7_2),.clk(gclk));
	jdff dff_A_udOtkEGA8_0(.dout(w_dff_A_lIrjR9Jj0_0),.din(w_dff_A_udOtkEGA8_0),.clk(gclk));
	jdff dff_A_lIrjR9Jj0_0(.dout(w_dff_A_0Qtxkv1O2_0),.din(w_dff_A_lIrjR9Jj0_0),.clk(gclk));
	jdff dff_A_0Qtxkv1O2_0(.dout(G882),.din(w_dff_A_0Qtxkv1O2_0),.clk(gclk));
	jdff dff_A_1182Ow2c0_2(.dout(G767),.din(w_dff_A_1182Ow2c0_2),.clk(gclk));
	jdff dff_A_GtGQe1WM9_2(.dout(G807),.din(w_dff_A_GtGQe1WM9_2),.clk(gclk));
endmodule

