// Benchmark "c1908" written by ABC on Wed May 27 22:07:08 2020

module rf_c1908 ( 
    G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
    G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234, G237,
    G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n158, n159, n160,
    n161, n162, n163, n164, n166, n167, n168, n169, n171, n172, n173, n174,
    n175, n176, n177, n179, n180, n181, n182, n183, n184, n185, n186, n188,
    n189, n190, n192, n193, n195, n196, n197, n198, n199, n200, n202, n204,
    n205, n207, n208, n209, n210, n212, n213, n215, n216, n217, n218, n219,
    n220, n222, n224, n225, n226, n228, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n345,
    n346, n347, n348, n349, n350, n351, n352, n354, n355, n356, n357, n358,
    n359, n360, n361, n363, n364, n365, n366, n367, n368, n369, n370, n372,
    n373, n374, n375, n376, n377, n378, n380, n381, n382, n383, n384, n386,
    n387, n388, n389, n390, n391, n392, n394, n395, n396, n397, n398, n399,
    n400, n401;
  jnot g000(.din(G146), .dout(n58));
  jxor g001(.dina(G140), .dinb(G125), .dout(n59));
  jxor g002(.dina(n59), .dinb(n58), .dout(n60));
  jnot g003(.din(G953), .dout(n61));
  jand g004(.dina(n61), .dinb(G234), .dout(n62));
  jand g005(.dina(n62), .dinb(G221), .dout(n63));
  jxor g006(.dina(n63), .dinb(G137), .dout(n64));
  jxor g007(.dina(G128), .dinb(G119), .dout(n65));
  jxor g008(.dina(n65), .dinb(n64), .dout(n66));
  jxor g009(.dina(n66), .dinb(G110), .dout(n67));
  jxor g010(.dina(n67), .dinb(n60), .dout(n68));
  jor  g011(.dina(n68), .dinb(G902), .dout(n69));
  jnot g012(.din(G902), .dout(n70));
  jand g013(.dina(n70), .dinb(G234), .dout(n71));
  jnot g014(.din(n71), .dout(n72));
  jand g015(.dina(n72), .dinb(G217), .dout(n73));
  jxor g016(.dina(n73), .dinb(n69), .dout(n74));
  jnot g017(.din(G134), .dout(n75));
  jxor g018(.dina(G137), .dinb(n75), .dout(n76));
  jnot g019(.din(G131), .dout(n77));
  jxor g020(.dina(G146), .dinb(G143), .dout(n78));
  jxor g021(.dina(n78), .dinb(G128), .dout(n79));
  jxor g022(.dina(n79), .dinb(n77), .dout(n80));
  jxor g023(.dina(n80), .dinb(n76), .dout(n81));
  jnot g024(.din(G113), .dout(n82));
  jxor g025(.dina(G119), .dinb(G116), .dout(n83));
  jxor g026(.dina(n83), .dinb(n82), .dout(n84));
  jnot g027(.din(G210), .dout(n85));
  jor  g028(.dina(G953), .dinb(G237), .dout(n86));
  jor  g029(.dina(n86), .dinb(n85), .dout(n87));
  jxor g030(.dina(n87), .dinb(G101), .dout(n88));
  jxor g031(.dina(n88), .dinb(n84), .dout(n89));
  jxor g032(.dina(n89), .dinb(n81), .dout(n90));
  jand g033(.dina(n90), .dinb(n70), .dout(n91));
  jxor g034(.dina(n91), .dinb(G472), .dout(n92));
  jand g035(.dina(n92), .dinb(n74), .dout(n93));
  jor  g036(.dina(G902), .dinb(G237), .dout(n94));
  jand g037(.dina(n94), .dinb(G214), .dout(n95));
  jnot g038(.din(n95), .dout(n96));
  jand g039(.dina(n94), .dinb(G210), .dout(n97));
  jnot g040(.din(G110), .dout(n98));
  jxor g041(.dina(G122), .dinb(n98), .dout(n99));
  jxor g042(.dina(G107), .dinb(G104), .dout(n100));
  jxor g043(.dina(n100), .dinb(G101), .dout(n101));
  jxor g044(.dina(n101), .dinb(n84), .dout(n102));
  jxor g045(.dina(n102), .dinb(n99), .dout(n103));
  jand g046(.dina(n61), .dinb(G224), .dout(n104));
  jxor g047(.dina(n79), .dinb(G125), .dout(n105));
  jxor g048(.dina(n105), .dinb(n104), .dout(n106));
  jxor g049(.dina(n106), .dinb(n103), .dout(n107));
  jand g050(.dina(n107), .dinb(n70), .dout(n108));
  jxor g051(.dina(n108), .dinb(n97), .dout(n109));
  jand g052(.dina(n109), .dinb(n96), .dout(n110));
  jnot g053(.din(G221), .dout(n111));
  jor  g054(.dina(n71), .dinb(n111), .dout(n112));
  jxor g055(.dina(G140), .dinb(G110), .dout(n113));
  jand g056(.dina(n61), .dinb(G227), .dout(n114));
  jxor g057(.dina(n114), .dinb(n101), .dout(n115));
  jxor g058(.dina(n115), .dinb(n113), .dout(n116));
  jxor g059(.dina(n116), .dinb(n81), .dout(n117));
  jand g060(.dina(n117), .dinb(n70), .dout(n118));
  jxor g061(.dina(n118), .dinb(G469), .dout(n119));
  jand g062(.dina(n119), .dinb(n112), .dout(n120));
  jand g063(.dina(n120), .dinb(n110), .dout(n121));
  jand g064(.dina(n121), .dinb(n93), .dout(n122));
  jnot g065(.din(G478), .dout(n123));
  jxor g066(.dina(G143), .dinb(G128), .dout(n124));
  jand g067(.dina(n62), .dinb(G217), .dout(n125));
  jxor g068(.dina(G122), .dinb(G116), .dout(n126));
  jxor g069(.dina(G134), .dinb(G107), .dout(n127));
  jxor g070(.dina(n127), .dinb(n126), .dout(n128));
  jxor g071(.dina(n128), .dinb(n125), .dout(n129));
  jxor g072(.dina(n129), .dinb(n124), .dout(n130));
  jand g073(.dina(n130), .dinb(n70), .dout(n131));
  jxor g074(.dina(n131), .dinb(n123), .dout(n132));
  jnot g075(.din(G475), .dout(n133));
  jxor g076(.dina(G143), .dinb(n77), .dout(n134));
  jxor g077(.dina(G122), .dinb(n82), .dout(n135));
  jxor g078(.dina(n135), .dinb(G104), .dout(n136));
  jnot g079(.din(G214), .dout(n137));
  jor  g080(.dina(n86), .dinb(n137), .dout(n138));
  jxor g081(.dina(n138), .dinb(n60), .dout(n139));
  jxor g082(.dina(n139), .dinb(n136), .dout(n140));
  jxor g083(.dina(n140), .dinb(n134), .dout(n141));
  jand g084(.dina(n141), .dinb(n70), .dout(n142));
  jxor g085(.dina(n142), .dinb(n133), .dout(n143));
  jand g086(.dina(n143), .dinb(n132), .dout(n144));
  jor  g087(.dina(n61), .dinb(G898), .dout(n145));
  jand g088(.dina(G237), .dinb(G234), .dout(n146));
  jor  g089(.dina(n146), .dinb(n70), .dout(n147));
  jor  g090(.dina(n147), .dinb(n145), .dout(n148));
  jnot g091(.din(n146), .dout(n149));
  jand g092(.dina(n61), .dinb(G952), .dout(n150));
  jand g093(.dina(n150), .dinb(n149), .dout(n151));
  jnot g094(.din(n151), .dout(n152));
  jand g095(.dina(n152), .dinb(n148), .dout(n153));
  jnot g096(.din(n153), .dout(n154));
  jand g097(.dina(n154), .dinb(n144), .dout(n155));
  jand g098(.dina(n155), .dinb(n122), .dout(n156));
  jxor g099(.dina(n156), .dinb(G101), .dout(G3));
  jnot g100(.din(n92), .dout(n158));
  jand g101(.dina(n158), .dinb(n74), .dout(n159));
  jand g102(.dina(n159), .dinb(n121), .dout(n160));
  jxor g103(.dina(n142), .dinb(G475), .dout(n161));
  jand g104(.dina(n161), .dinb(n132), .dout(n162));
  jand g105(.dina(n162), .dinb(n154), .dout(n163));
  jand g106(.dina(n163), .dinb(n160), .dout(n164));
  jxor g107(.dina(n164), .dinb(G104), .dout(G6));
  jxor g108(.dina(n131), .dinb(G478), .dout(n166));
  jand g109(.dina(n143), .dinb(n166), .dout(n167));
  jand g110(.dina(n167), .dinb(n154), .dout(n168));
  jand g111(.dina(n168), .dinb(n160), .dout(n169));
  jxor g112(.dina(n169), .dinb(G107), .dout(G9));
  jnot g113(.din(n60), .dout(n171));
  jxor g114(.dina(n67), .dinb(n171), .dout(n172));
  jand g115(.dina(n172), .dinb(n70), .dout(n173));
  jxor g116(.dina(n73), .dinb(n173), .dout(n174));
  jand g117(.dina(n158), .dinb(n174), .dout(n175));
  jand g118(.dina(n175), .dinb(n155), .dout(n176));
  jand g119(.dina(n176), .dinb(n121), .dout(n177));
  jxor g120(.dina(n177), .dinb(G110), .dout(G12));
  jand g121(.dina(n92), .dinb(n174), .dout(n179));
  jand g122(.dina(n179), .dinb(n121), .dout(n180));
  jor  g123(.dina(n61), .dinb(G900), .dout(n181));
  jor  g124(.dina(n181), .dinb(n147), .dout(n182));
  jand g125(.dina(n182), .dinb(n152), .dout(n183));
  jnot g126(.din(n183), .dout(n184));
  jand g127(.dina(n184), .dinb(n167), .dout(n185));
  jand g128(.dina(n185), .dinb(n180), .dout(n186));
  jxor g129(.dina(n186), .dinb(G128), .dout(G30));
  jand g130(.dina(n161), .dinb(n166), .dout(n188));
  jand g131(.dina(n188), .dinb(n184), .dout(n189));
  jand g132(.dina(n189), .dinb(n122), .dout(n190));
  jxor g133(.dina(n190), .dinb(G143), .dout(G45));
  jand g134(.dina(n184), .dinb(n162), .dout(n192));
  jand g135(.dina(n192), .dinb(n180), .dout(n193));
  jxor g136(.dina(n193), .dinb(G146), .dout(G48));
  jnot g137(.din(G469), .dout(n195));
  jxor g138(.dina(n118), .dinb(n195), .dout(n196));
  jand g139(.dina(n196), .dinb(n112), .dout(n197));
  jand g140(.dina(n197), .dinb(n110), .dout(n198));
  jand g141(.dina(n198), .dinb(n93), .dout(n199));
  jand g142(.dina(n199), .dinb(n163), .dout(n200));
  jxor g143(.dina(n200), .dinb(G113), .dout(G15));
  jand g144(.dina(n199), .dinb(n168), .dout(n202));
  jxor g145(.dina(n202), .dinb(G116), .dout(G18));
  jand g146(.dina(n198), .dinb(n179), .dout(n204));
  jand g147(.dina(n204), .dinb(n155), .dout(n205));
  jxor g148(.dina(n205), .dinb(G119), .dout(G21));
  jand g149(.dina(n197), .dinb(n159), .dout(n207));
  jand g150(.dina(n154), .dinb(n110), .dout(n208));
  jand g151(.dina(n208), .dinb(n188), .dout(n209));
  jand g152(.dina(n209), .dinb(n207), .dout(n210));
  jxor g153(.dina(n210), .dinb(G122), .dout(G24));
  jand g154(.dina(n192), .dinb(n175), .dout(n212));
  jand g155(.dina(n212), .dinb(n198), .dout(n213));
  jxor g156(.dina(n213), .dinb(G125), .dout(G27));
  jnot g157(.din(n97), .dout(n215));
  jxor g158(.dina(n108), .dinb(n215), .dout(n216));
  jand g159(.dina(n216), .dinb(n96), .dout(n217));
  jand g160(.dina(n217), .dinb(n120), .dout(n218));
  jand g161(.dina(n218), .dinb(n93), .dout(n219));
  jand g162(.dina(n219), .dinb(n192), .dout(n220));
  jxor g163(.dina(n220), .dinb(G131), .dout(G33));
  jand g164(.dina(n219), .dinb(n185), .dout(n222));
  jxor g165(.dina(n222), .dinb(G134), .dout(G36));
  jand g166(.dina(n184), .dinb(n144), .dout(n224));
  jand g167(.dina(n224), .dinb(n179), .dout(n225));
  jand g168(.dina(n225), .dinb(n218), .dout(n226));
  jxor g169(.dina(n226), .dinb(G137), .dout(G39));
  jand g170(.dina(n218), .dinb(n212), .dout(n228));
  jxor g171(.dina(n228), .dinb(G140), .dout(G42));
  jor  g172(.dina(n177), .dinb(n169), .dout(n230));
  jor  g173(.dina(n202), .dinb(n164), .dout(n231));
  jor  g174(.dina(n231), .dinb(n230), .dout(n232));
  jor  g175(.dina(n205), .dinb(n156), .dout(n233));
  jor  g176(.dina(n210), .dinb(n200), .dout(n234));
  jor  g177(.dina(n234), .dinb(n233), .dout(n235));
  jor  g178(.dina(n235), .dinb(n232), .dout(n236));
  jor  g179(.dina(n220), .dinb(n193), .dout(n237));
  jor  g180(.dina(n222), .dinb(n186), .dout(n238));
  jor  g181(.dina(n238), .dinb(n237), .dout(n239));
  jor  g182(.dina(n228), .dinb(n190), .dout(n240));
  jor  g183(.dina(n226), .dinb(n213), .dout(n241));
  jor  g184(.dina(n241), .dinb(n240), .dout(n242));
  jor  g185(.dina(n242), .dinb(n239), .dout(n243));
  jor  g186(.dina(n243), .dinb(n236), .dout(n244));
  jor  g187(.dina(n218), .dinb(n198), .dout(n245));
  jand g188(.dina(n245), .dinb(n144), .dout(n246));
  jand g189(.dina(n217), .dinb(n197), .dout(n247));
  jxor g190(.dina(n143), .dinb(n132), .dout(n248));
  jand g191(.dina(n248), .dinb(n247), .dout(n249));
  jor  g192(.dina(n249), .dinb(n246), .dout(n250));
  jand g193(.dina(n250), .dinb(n159), .dout(n251));
  jand g194(.dina(n217), .dinb(n144), .dout(n252));
  jor  g195(.dina(n92), .dinb(n174), .dout(n253));
  jor  g196(.dina(n158), .dinb(n74), .dout(n254));
  jand g197(.dina(n197), .dinb(n254), .dout(n255));
  jand g198(.dina(n255), .dinb(n253), .dout(n256));
  jand g199(.dina(n256), .dinb(n252), .dout(n257));
  jor  g200(.dina(n257), .dinb(n251), .dout(n258));
  jand g201(.dina(n258), .dinb(n151), .dout(n259));
  jxor g202(.dina(n112), .dinb(n96), .dout(n260));
  jand g203(.dina(n260), .dinb(n151), .dout(n261));
  jand g204(.dina(n261), .dinb(n196), .dout(n262));
  jand g205(.dina(n262), .dinb(n216), .dout(n263));
  jand g206(.dina(n159), .dinb(n144), .dout(n264));
  jand g207(.dina(n264), .dinb(n263), .dout(n265));
  jor  g208(.dina(n265), .dinb(n259), .dout(n266));
  jor  g209(.dina(n266), .dinb(n244), .dout(n267));
  jand g210(.dina(n267), .dinb(G952), .dout(n268));
  jand g211(.dina(n252), .dinb(n207), .dout(n269));
  jor  g212(.dina(n269), .dinb(G953), .dout(n270));
  jor  g213(.dina(n270), .dinb(n268), .dout(G75));
  jnot g214(.din(n107), .dout(n272));
  jor  g215(.dina(n216), .dinb(n95), .dout(n273));
  jnot g216(.din(n112), .dout(n274));
  jor  g217(.dina(n196), .dinb(n274), .dout(n275));
  jor  g218(.dina(n275), .dinb(n273), .dout(n276));
  jor  g219(.dina(n253), .dinb(n276), .dout(n277));
  jnot g220(.din(n168), .dout(n278));
  jor  g221(.dina(n278), .dinb(n277), .dout(n279));
  jor  g222(.dina(n161), .dinb(n166), .dout(n280));
  jor  g223(.dina(n153), .dinb(n280), .dout(n281));
  jor  g224(.dina(n92), .dinb(n74), .dout(n282));
  jor  g225(.dina(n282), .dinb(n281), .dout(n283));
  jor  g226(.dina(n283), .dinb(n276), .dout(n284));
  jand g227(.dina(n284), .dinb(n279), .dout(n285));
  jnot g228(.din(n163), .dout(n286));
  jor  g229(.dina(n286), .dinb(n277), .dout(n287));
  jor  g230(.dina(n158), .dinb(n174), .dout(n288));
  jor  g231(.dina(n119), .dinb(n274), .dout(n289));
  jor  g232(.dina(n289), .dinb(n273), .dout(n290));
  jor  g233(.dina(n290), .dinb(n288), .dout(n291));
  jor  g234(.dina(n291), .dinb(n278), .dout(n292));
  jand g235(.dina(n292), .dinb(n287), .dout(n293));
  jand g236(.dina(n293), .dinb(n285), .dout(n294));
  jor  g237(.dina(n276), .dinb(n288), .dout(n295));
  jor  g238(.dina(n281), .dinb(n295), .dout(n296));
  jor  g239(.dina(n290), .dinb(n254), .dout(n297));
  jor  g240(.dina(n297), .dinb(n281), .dout(n298));
  jand g241(.dina(n298), .dinb(n296), .dout(n299));
  jor  g242(.dina(n291), .dinb(n286), .dout(n300));
  jor  g243(.dina(n289), .dinb(n253), .dout(n301));
  jnot g244(.din(n188), .dout(n302));
  jor  g245(.dina(n153), .dinb(n273), .dout(n303));
  jor  g246(.dina(n303), .dinb(n302), .dout(n304));
  jor  g247(.dina(n304), .dinb(n301), .dout(n305));
  jand g248(.dina(n305), .dinb(n300), .dout(n306));
  jand g249(.dina(n306), .dinb(n299), .dout(n307));
  jand g250(.dina(n307), .dinb(n294), .dout(n308));
  jor  g251(.dina(n254), .dinb(n276), .dout(n309));
  jor  g252(.dina(n143), .dinb(n166), .dout(n310));
  jor  g253(.dina(n183), .dinb(n310), .dout(n311));
  jor  g254(.dina(n311), .dinb(n309), .dout(n312));
  jor  g255(.dina(n109), .dinb(n95), .dout(n313));
  jor  g256(.dina(n313), .dinb(n275), .dout(n314));
  jor  g257(.dina(n314), .dinb(n288), .dout(n315));
  jor  g258(.dina(n315), .dinb(n311), .dout(n316));
  jand g259(.dina(n316), .dinb(n312), .dout(n317));
  jnot g260(.din(n185), .dout(n318));
  jor  g261(.dina(n318), .dinb(n309), .dout(n319));
  jor  g262(.dina(n315), .dinb(n318), .dout(n320));
  jand g263(.dina(n320), .dinb(n319), .dout(n321));
  jand g264(.dina(n321), .dinb(n317), .dout(n322));
  jnot g265(.din(n189), .dout(n323));
  jor  g266(.dina(n323), .dinb(n295), .dout(n324));
  jor  g267(.dina(n311), .dinb(n282), .dout(n325));
  jor  g268(.dina(n314), .dinb(n325), .dout(n326));
  jand g269(.dina(n326), .dinb(n324), .dout(n327));
  jor  g270(.dina(n325), .dinb(n290), .dout(n328));
  jor  g271(.dina(n183), .dinb(n280), .dout(n329));
  jor  g272(.dina(n329), .dinb(n254), .dout(n330));
  jor  g273(.dina(n330), .dinb(n314), .dout(n331));
  jand g274(.dina(n331), .dinb(n328), .dout(n332));
  jand g275(.dina(n332), .dinb(n327), .dout(n333));
  jand g276(.dina(n333), .dinb(n322), .dout(n334));
  jand g277(.dina(n334), .dinb(n308), .dout(n335));
  jand g278(.dina(G902), .dinb(G210), .dout(n336));
  jnot g279(.din(n336), .dout(n337));
  jor  g280(.dina(n337), .dinb(n335), .dout(n338));
  jor  g281(.dina(n338), .dinb(n272), .dout(n339));
  jor  g282(.dina(n61), .dinb(G952), .dout(n340));
  jand g283(.dina(n336), .dinb(n244), .dout(n341));
  jor  g284(.dina(n341), .dinb(n107), .dout(n342));
  jand g285(.dina(n342), .dinb(n340), .dout(n343));
  jand g286(.dina(n343), .dinb(n339), .dout(G51));
  jnot g287(.din(n117), .dout(n345));
  jand g288(.dina(G902), .dinb(G469), .dout(n346));
  jnot g289(.din(n346), .dout(n347));
  jor  g290(.dina(n347), .dinb(n335), .dout(n348));
  jor  g291(.dina(n348), .dinb(n345), .dout(n349));
  jand g292(.dina(n346), .dinb(n244), .dout(n350));
  jor  g293(.dina(n350), .dinb(n117), .dout(n351));
  jand g294(.dina(n351), .dinb(n340), .dout(n352));
  jand g295(.dina(n352), .dinb(n349), .dout(G54));
  jnot g296(.din(n141), .dout(n354));
  jand g297(.dina(G902), .dinb(G475), .dout(n355));
  jnot g298(.din(n355), .dout(n356));
  jor  g299(.dina(n356), .dinb(n335), .dout(n357));
  jor  g300(.dina(n357), .dinb(n354), .dout(n358));
  jand g301(.dina(n355), .dinb(n244), .dout(n359));
  jor  g302(.dina(n359), .dinb(n141), .dout(n360));
  jand g303(.dina(n360), .dinb(n340), .dout(n361));
  jand g304(.dina(n361), .dinb(n358), .dout(G60));
  jnot g305(.din(n130), .dout(n363));
  jand g306(.dina(G902), .dinb(G478), .dout(n364));
  jnot g307(.din(n364), .dout(n365));
  jor  g308(.dina(n365), .dinb(n335), .dout(n366));
  jor  g309(.dina(n366), .dinb(n363), .dout(n367));
  jand g310(.dina(n364), .dinb(n244), .dout(n368));
  jor  g311(.dina(n368), .dinb(n130), .dout(n369));
  jand g312(.dina(n369), .dinb(n340), .dout(n370));
  jand g313(.dina(n370), .dinb(n367), .dout(G63));
  jand g314(.dina(G902), .dinb(G217), .dout(n372));
  jand g315(.dina(n372), .dinb(n244), .dout(n373));
  jor  g316(.dina(n373), .dinb(n172), .dout(n374));
  jnot g317(.din(n372), .dout(n375));
  jor  g318(.dina(n375), .dinb(n335), .dout(n376));
  jor  g319(.dina(n376), .dinb(n68), .dout(n377));
  jand g320(.dina(n377), .dinb(n340), .dout(n378));
  jand g321(.dina(n378), .dinb(n374), .dout(G66));
  jnot g322(.din(n145), .dout(n380));
  jor  g323(.dina(n308), .dinb(G953), .dout(n381));
  jor  g324(.dina(n61), .dinb(G224), .dout(n382));
  jand g325(.dina(n382), .dinb(n381), .dout(n383));
  jxor g326(.dina(n383), .dinb(n103), .dout(n384));
  jor  g327(.dina(n384), .dinb(n380), .dout(G69));
  jor  g328(.dina(n334), .dinb(G953), .dout(n386));
  jor  g329(.dina(n61), .dinb(G227), .dout(n387));
  jand g330(.dina(n387), .dinb(n181), .dout(n388));
  jand g331(.dina(n388), .dinb(n386), .dout(n389));
  jnot g332(.din(n181), .dout(n390));
  jxor g333(.dina(n81), .dinb(n59), .dout(n391));
  jor  g334(.dina(n391), .dinb(n390), .dout(n392));
  jxor g335(.dina(n392), .dinb(n389), .dout(G72));
  jnot g336(.din(n90), .dout(n394));
  jand g337(.dina(G902), .dinb(G472), .dout(n395));
  jnot g338(.din(n395), .dout(n396));
  jor  g339(.dina(n396), .dinb(n335), .dout(n397));
  jor  g340(.dina(n397), .dinb(n394), .dout(n398));
  jand g341(.dina(n395), .dinb(n244), .dout(n399));
  jor  g342(.dina(n399), .dinb(n90), .dout(n400));
  jand g343(.dina(n400), .dinb(n340), .dout(n401));
  jand g344(.dina(n401), .dinb(n398), .dout(G57));
endmodule


