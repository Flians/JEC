/*

c499:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jdff: 435
	jor: 10
	jand: 61

Summary:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jdff: 435
	jor: 10
	jand: 61
*/

module c499(gclk, Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9, Gid10, Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19, Gid20, Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29, Gid30, Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr, God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10, God11, God12, God13, God14, God15, God16, God17, God18, God19, God20, God21, God22, God23, God24, God25, God26, God27, God28, God29, God30, God31);
	input gclk;
	input Gid0;
	input Gid1;
	input Gid2;
	input Gid3;
	input Gid4;
	input Gid5;
	input Gid6;
	input Gid7;
	input Gid8;
	input Gid9;
	input Gid10;
	input Gid11;
	input Gid12;
	input Gid13;
	input Gid14;
	input Gid15;
	input Gid16;
	input Gid17;
	input Gid18;
	input Gid19;
	input Gid20;
	input Gid21;
	input Gid22;
	input Gid23;
	input Gid24;
	input Gid25;
	input Gid26;
	input Gid27;
	input Gid28;
	input Gid29;
	input Gid30;
	input Gid31;
	input Gic0;
	input Gic1;
	input Gic2;
	input Gic3;
	input Gic4;
	input Gic5;
	input Gic6;
	input Gic7;
	input Gr;
	output God0;
	output God1;
	output God2;
	output God3;
	output God4;
	output God5;
	output God6;
	output God7;
	output God8;
	output God9;
	output God10;
	output God11;
	output God12;
	output God13;
	output God14;
	output God15;
	output God16;
	output God17;
	output God18;
	output God19;
	output God20;
	output God21;
	output God22;
	output God23;
	output God24;
	output God25;
	output God26;
	output God27;
	output God28;
	output God29;
	output God30;
	output God31;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n178;
	wire n179;
	wire n181;
	wire n182;
	wire n184;
	wire n185;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n192;
	wire n194;
	wire n196;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n204;
	wire n206;
	wire n208;
	wire n210;
	wire n211;
	wire n212;
	wire n214;
	wire n216;
	wire n218;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n233;
	wire n235;
	wire n237;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n244;
	wire n246;
	wire n248;
	wire n250;
	wire n251;
	wire n252;
	wire n254;
	wire n256;
	wire n258;
	wire n260;
	wire n261;
	wire n263;
	wire n265;
	wire n267;
	wire[2:0] w_Gid0_0;
	wire[2:0] w_Gid1_0;
	wire[2:0] w_Gid2_0;
	wire[2:0] w_Gid3_0;
	wire[2:0] w_Gid4_0;
	wire[2:0] w_Gid5_0;
	wire[2:0] w_Gid6_0;
	wire[2:0] w_Gid7_0;
	wire[2:0] w_Gid8_0;
	wire[2:0] w_Gid9_0;
	wire[2:0] w_Gid10_0;
	wire[2:0] w_Gid11_0;
	wire[2:0] w_Gid12_0;
	wire[2:0] w_Gid13_0;
	wire[2:0] w_Gid14_0;
	wire[2:0] w_Gid15_0;
	wire[2:0] w_Gid16_0;
	wire[2:0] w_Gid17_0;
	wire[2:0] w_Gid18_0;
	wire[2:0] w_Gid19_0;
	wire[2:0] w_Gid20_0;
	wire[2:0] w_Gid21_0;
	wire[2:0] w_Gid22_0;
	wire[2:0] w_Gid23_0;
	wire[2:0] w_Gid24_0;
	wire[2:0] w_Gid25_0;
	wire[2:0] w_Gid26_0;
	wire[2:0] w_Gid27_0;
	wire[2:0] w_Gid28_0;
	wire[2:0] w_Gid29_0;
	wire[2:0] w_Gid30_0;
	wire[2:0] w_Gid31_0;
	wire[2:0] w_n74_0;
	wire[2:0] w_n74_1;
	wire[2:0] w_n74_2;
	wire[1:0] w_n74_3;
	wire[1:0] w_n78_0;
	wire[1:0] w_n85_0;
	wire[2:0] w_n87_0;
	wire[1:0] w_n87_1;
	wire[2:0] w_n88_0;
	wire[2:0] w_n88_1;
	wire[1:0] w_n93_0;
	wire[1:0] w_n97_0;
	wire[2:0] w_n102_0;
	wire[1:0] w_n102_1;
	wire[1:0] w_n107_0;
	wire[1:0] w_n111_0;
	wire[2:0] w_n116_0;
	wire[1:0] w_n116_1;
	wire[2:0] w_n117_0;
	wire[2:0] w_n117_1;
	wire[1:0] w_n118_0;
	wire[2:0] w_n126_0;
	wire[1:0] w_n126_1;
	wire[2:0] w_n127_0;
	wire[2:0] w_n127_1;
	wire[2:0] w_n135_0;
	wire[1:0] w_n135_1;
	wire[1:0] w_n141_0;
	wire[1:0] w_n145_0;
	wire[2:0] w_n150_0;
	wire[1:0] w_n150_1;
	wire[2:0] w_n159_0;
	wire[1:0] w_n159_1;
	wire[2:0] w_n167_0;
	wire[1:0] w_n167_1;
	wire[2:0] w_n173_0;
	wire[1:0] w_n174_0;
	wire[2:0] w_n175_0;
	wire[1:0] w_n175_1;
	wire[2:0] w_n178_0;
	wire[2:0] w_n178_1;
	wire[2:0] w_n181_0;
	wire[2:0] w_n181_1;
	wire[2:0] w_n184_0;
	wire[2:0] w_n184_1;
	wire[2:0] w_n187_0;
	wire[2:0] w_n187_1;
	wire[1:0] w_n188_0;
	wire[2:0] w_n189_0;
	wire[1:0] w_n189_1;
	wire[2:0] w_n198_0;
	wire[2:0] w_n198_1;
	wire[1:0] w_n199_0;
	wire[2:0] w_n201_0;
	wire[1:0] w_n201_1;
	wire[2:0] w_n211_0;
	wire[1:0] w_n211_1;
	wire[1:0] w_n220_0;
	wire[1:0] w_n228_0;
	wire[1:0] w_n229_0;
	wire[2:0] w_n230_0;
	wire[1:0] w_n230_1;
	wire[1:0] w_n240_0;
	wire[2:0] w_n241_0;
	wire[1:0] w_n241_1;
	wire[1:0] w_n250_0;
	wire[2:0] w_n251_0;
	wire[1:0] w_n251_1;
	wire[2:0] w_n260_0;
	wire[1:0] w_n260_1;
	wire w_dff_B_zLnaYhAk3_1;
	wire w_dff_A_ncZ1c8Jf5_1;
	wire w_dff_A_2EossxO28_2;
	wire w_dff_A_CPfiQIe21_1;
	wire w_dff_A_VQyutGvp7_2;
	wire w_dff_A_KPVIS0wL0_1;
	wire w_dff_A_ziY5YhhM6_2;
	wire w_dff_A_vaNRwcjV5_1;
	wire w_dff_A_aj31bKFg6_1;
	wire w_dff_A_168aCpzU1_1;
	wire w_dff_A_ihKwuW0B4_2;
	wire w_dff_A_waxZHvun6_1;
	wire w_dff_A_HzqdGCER1_1;
	wire w_dff_A_p63vZo0A3_0;
	wire w_dff_A_vfU1zxwq9_0;
	wire w_dff_A_ZytrEjEw0_0;
	wire w_dff_A_yGPBCphy2_0;
	wire w_dff_A_DZ809y9N7_1;
	wire w_dff_A_mwPam5KB4_1;
	wire w_dff_A_VAVyDwbQ9_1;
	wire w_dff_A_qcxs7akv1_1;
	wire w_dff_A_hCqw5WZ39_0;
	wire w_dff_A_WoHjTkUS1_0;
	wire w_dff_A_iOAy8MW69_0;
	wire w_dff_A_TSQ0bVc40_0;
	wire w_dff_A_hDtm3F0v9_1;
	wire w_dff_A_sptfIzyr5_1;
	wire w_dff_A_ueGalGHp5_1;
	wire w_dff_A_0jOseWON2_1;
	wire w_dff_A_04w2cuD38_0;
	wire w_dff_A_m0akYXC16_0;
	wire w_dff_A_3fiVKfNN5_0;
	wire w_dff_A_8NCA6Alt8_0;
	wire w_dff_A_RVMOrcW43_1;
	wire w_dff_A_OHfnjzZ42_1;
	wire w_dff_A_m1bX7gt12_1;
	wire w_dff_A_VhyRl4SB1_1;
	wire w_dff_B_1JtBnWzE5_2;
	wire w_dff_B_9Qw26Ghh9_2;
	wire w_dff_A_oCzz8iJF7_0;
	wire w_dff_A_q1wejxtZ8_0;
	wire w_dff_A_hL8dYl2p6_0;
	wire w_dff_A_kYT75gjZ8_2;
	wire w_dff_A_yzQk7i3X5_2;
	wire w_dff_A_xj9ez3eS0_2;
	wire w_dff_A_5y2hzcLU2_0;
	wire w_dff_A_qYZoe9lW8_0;
	wire w_dff_A_hUNFsei67_0;
	wire w_dff_A_dqc5tMAp0_0;
	wire w_dff_A_gWkHxOwb2_1;
	wire w_dff_A_RLoADiQL6_1;
	wire w_dff_A_NGNee5407_1;
	wire w_dff_A_z3kZ9A2m7_1;
	wire w_dff_B_LnPM9yPY5_1;
	wire w_dff_A_iovCjw1W2_0;
	wire w_dff_A_NiL0Jq5Y6_0;
	wire w_dff_A_tAhxaWUj3_0;
	wire w_dff_A_xvIr2wzL9_2;
	wire w_dff_A_xXqfDksf7_2;
	wire w_dff_A_WSh7d3nm1_2;
	wire w_dff_A_2ryBKwmj2_1;
	wire w_dff_A_qn4MyplS4_1;
	wire w_dff_A_liH1Uy9H7_1;
	wire w_dff_A_HVPAQLgR8_1;
	wire w_dff_A_sP1QHHi05_2;
	wire w_dff_A_dvobQml51_2;
	wire w_dff_A_NtPfuvxQ8_2;
	wire w_dff_A_AECdvskk8_2;
	wire w_dff_A_Ljjz6T0o5_0;
	wire w_dff_A_e9yoTzR81_1;
	wire w_dff_A_y9e5IHdq7_1;
	wire w_dff_A_jq3AilBr5_1;
	wire w_dff_A_GKF9Xxt81_1;
	wire w_dff_A_XoLKLvV84_2;
	wire w_dff_A_4B65W6kT7_2;
	wire w_dff_A_dz94ukJp1_2;
	wire w_dff_A_zfN8Qyt76_2;
	wire w_dff_A_YUTr4cZx2_1;
	wire w_dff_A_Ck6uPS2X6_1;
	wire w_dff_A_1iTlczd10_1;
	wire w_dff_A_mxBeo0iR1_1;
	wire w_dff_A_rijR7ckf2_1;
	wire w_dff_A_0t9hgo6Z4_2;
	wire w_dff_A_RvJvErBH1_2;
	wire w_dff_A_WMoCnv7L8_2;
	wire w_dff_A_BAk5pbYc4_2;
	wire w_dff_A_e0deb75v8_0;
	wire w_dff_B_e93qed7n2_1;
	wire w_dff_A_Zixou12u7_1;
	wire w_dff_A_FREWL7EQ4_0;
	wire w_dff_A_r5mUtZ1w0_0;
	wire w_dff_A_jXuuHFic2_0;
	wire w_dff_A_hqdBNAVq0_0;
	wire w_dff_A_LkmloUJ54_0;
	wire w_dff_A_KMUGUlvE4_0;
	wire w_dff_A_0XgOS5ZN1_0;
	wire w_dff_A_Qaj5Waxr0_0;
	wire w_dff_A_5ycgIj5v7_0;
	wire w_dff_A_T3t3nIWk8_0;
	wire w_dff_A_rvnDP1ph8_0;
	wire w_dff_A_Cc9KnMvu6_0;
	wire w_dff_A_BFT77zb42_0;
	wire w_dff_A_74wVKOLo1_0;
	wire w_dff_A_99MEHm830_0;
	wire w_dff_A_FCiKgdIT2_0;
	wire w_dff_A_vXuNS80w5_0;
	wire w_dff_A_yf9aZ6Bo5_0;
	wire w_dff_A_qJXJclC73_0;
	wire w_dff_A_66aYhiXR7_0;
	wire w_dff_A_CHas1LHi4_0;
	wire w_dff_A_fG3UcLW36_0;
	wire w_dff_A_mCVYHet33_2;
	wire w_dff_A_aE84ATNk0_2;
	wire w_dff_A_up7CYHIQ2_2;
	wire w_dff_A_s6EPuhFG3_1;
	wire w_dff_A_q1Tmkjhg8_0;
	wire w_dff_A_WoMNUxuA9_0;
	wire w_dff_A_jTuDcu4A1_0;
	wire w_dff_A_sJKUTsoZ6_0;
	wire w_dff_A_zTXQJi4O2_0;
	wire w_dff_A_MDHdZqXY2_0;
	wire w_dff_A_zGVrZsi95_0;
	wire w_dff_A_l6x9zAjl7_0;
	wire w_dff_A_7tleaXJX8_0;
	wire w_dff_A_ZLw59waI6_0;
	wire w_dff_A_pbkv4RCK0_0;
	wire w_dff_A_h6BO7UyX8_0;
	wire w_dff_A_os3UQUEN7_0;
	wire w_dff_A_BUgum97z5_0;
	wire w_dff_A_8iHpVQn43_0;
	wire w_dff_A_QVqaKatW4_0;
	wire w_dff_A_go8BBj3z6_0;
	wire w_dff_A_4I3nMOGK9_0;
	wire w_dff_A_F9swWSKi8_0;
	wire w_dff_B_aiquepbI0_2;
	wire w_dff_B_XdS5RqLz8_2;
	wire w_dff_A_duyvdjvf5_0;
	wire w_dff_A_VOoJv4I02_0;
	wire w_dff_A_JXsgy0qd6_0;
	wire w_dff_A_ataSTmQa3_2;
	wire w_dff_A_h8aYYNzM2_2;
	wire w_dff_A_m0QOCOpM9_2;
	wire w_dff_A_L009HIxL8_1;
	wire w_dff_A_obwLJFET9_0;
	wire w_dff_A_38vUVyGS0_0;
	wire w_dff_A_tyNC6W9l4_0;
	wire w_dff_A_pgv0ZQTQ7_0;
	wire w_dff_A_rZIop5ca6_0;
	wire w_dff_A_LBLWlta38_0;
	wire w_dff_A_hO6pMVH44_0;
	wire w_dff_A_XSgzrLmB4_0;
	wire w_dff_A_WcyjloGZ2_0;
	wire w_dff_A_cFjvw5JH8_0;
	wire w_dff_A_7H716H7I0_0;
	wire w_dff_A_l67q1CMO8_0;
	wire w_dff_A_E1bn7CGa6_0;
	wire w_dff_A_t825I58D2_0;
	wire w_dff_A_juBNwpGl8_0;
	wire w_dff_A_JIjB9Fy70_0;
	wire w_dff_A_UadGAP8n7_0;
	wire w_dff_A_CB67CI6b8_0;
	wire w_dff_A_zjbSdnLV9_0;
	wire w_dff_A_0Rjp8F4g1_0;
	wire w_dff_A_kh98CfO54_0;
	wire w_dff_A_GKKIGPxi3_0;
	wire w_dff_A_CTXqkuQH4_0;
	wire w_dff_A_ohLGYgoh5_0;
	wire w_dff_A_jV3smZcq9_0;
	wire w_dff_A_imCf9JM81_0;
	wire w_dff_A_vyKRC8Fd8_0;
	wire w_dff_A_NEp2ucVn4_0;
	wire w_dff_A_OvZnt1XA4_0;
	wire w_dff_A_i4agnnAC7_0;
	wire w_dff_A_TCzJcbbe7_0;
	wire w_dff_A_EKLPA0jg1_0;
	wire w_dff_A_CFZSfiML6_0;
	wire w_dff_A_GYa4Asfj9_0;
	wire w_dff_A_NDFosJTS4_0;
	wire w_dff_A_kFHIGF7R9_0;
	wire w_dff_A_kFK45YSH2_0;
	wire w_dff_A_icOdlJz91_0;
	wire w_dff_A_1A0bEObr3_0;
	wire w_dff_A_OZgTqKq69_0;
	wire w_dff_A_NwoNFBMR4_0;
	wire w_dff_A_LMa73EUp2_0;
	wire w_dff_A_gwDqsdTV1_0;
	wire w_dff_A_8X8tpmhG6_0;
	wire w_dff_A_uVzoXuKk8_0;
	wire w_dff_A_A8v23lbd1_0;
	wire w_dff_A_y2iRngSq2_0;
	wire w_dff_A_cU4WwANM7_0;
	wire w_dff_A_qlllOe9G5_0;
	wire w_dff_A_AaSaQZxW2_0;
	wire w_dff_A_uPXwmlmu1_0;
	wire w_dff_A_WSkG8AvX5_0;
	wire w_dff_A_tuZS5JXj2_0;
	wire w_dff_A_S9zK4OwL6_0;
	wire w_dff_A_nUxSZ8Jt8_0;
	wire w_dff_A_nzoEoApV7_0;
	wire w_dff_A_2HhnoT8C7_0;
	wire w_dff_A_VEDrPZW67_0;
	wire w_dff_A_ZCxqcaoc6_0;
	wire w_dff_A_LvZR9Phi7_0;
	wire w_dff_A_PsBjJkkA1_0;
	wire w_dff_A_1mS88ppG6_0;
	wire w_dff_A_aVmEZv8P6_0;
	wire w_dff_A_MyJEfLPR1_0;
	wire w_dff_A_WYgMBVAS8_0;
	wire w_dff_A_YH47ltTr5_0;
	wire w_dff_A_GD61wjyg1_0;
	wire w_dff_A_PZmG05BB1_0;
	wire w_dff_A_IIherzhR4_0;
	wire w_dff_A_fovtXY267_0;
	wire w_dff_A_kbJT9drN5_0;
	wire w_dff_A_x5dBkqh31_0;
	wire w_dff_A_utaxoCqY8_0;
	wire w_dff_A_NklgPUGx9_0;
	wire w_dff_A_xUdDCLmE0_0;
	wire w_dff_A_PXjVvBEB9_0;
	wire w_dff_A_DpSR2YLJ5_0;
	wire w_dff_A_X9qv8aYt1_0;
	wire w_dff_A_4mvnpGSs4_0;
	wire w_dff_A_M2PaOgjg4_1;
	wire w_dff_A_gTU0I0Kb0_0;
	wire w_dff_A_WIs0Z4UN8_0;
	wire w_dff_A_u4wlr4fZ6_0;
	wire w_dff_A_GXgv57cO7_0;
	wire w_dff_A_wYwrtSa60_0;
	wire w_dff_A_bz7dgpLW0_0;
	wire w_dff_A_Gimmhwj84_0;
	wire w_dff_A_jdzJNB5P9_0;
	wire w_dff_A_krzVkPLu8_0;
	wire w_dff_A_ZVPfoTQT1_0;
	wire w_dff_A_T3PkQYSn8_0;
	wire w_dff_A_18CUV6Ru3_0;
	wire w_dff_A_6pVS6k936_0;
	wire w_dff_A_lzsodhkK0_0;
	wire w_dff_A_Twi8rjzG3_0;
	wire w_dff_A_DXylPXA64_0;
	wire w_dff_A_mAXnUtDa9_0;
	wire w_dff_A_BdHwYyGn0_0;
	wire w_dff_A_punfCYko1_0;
	wire w_dff_A_p6PpfRME7_0;
	wire w_dff_A_hAeLU9z48_0;
	wire w_dff_A_etOMWfyO9_0;
	wire w_dff_A_0XO7gUnA1_0;
	wire w_dff_A_QZnDrBzG9_0;
	wire w_dff_A_7tTQfzcv2_0;
	wire w_dff_A_SFMbC9eO1_0;
	wire w_dff_A_vwehtSZr8_0;
	wire w_dff_A_oXRTpgMH9_0;
	wire w_dff_A_s8PsiCvj2_0;
	wire w_dff_A_dfvbAn5o2_0;
	wire w_dff_A_13ziitp32_0;
	wire w_dff_A_Os2y9z362_0;
	wire w_dff_A_CDr5DGOV4_0;
	wire w_dff_A_P2zTSOq49_0;
	wire w_dff_A_wOEwAWjA8_0;
	wire w_dff_A_3Cq1DJl64_0;
	wire w_dff_A_ZKCrxvLZ9_0;
	wire w_dff_A_gOsP3EXH8_0;
	wire w_dff_A_h0Czj1or7_0;
	wire w_dff_A_VTLfBYCw0_0;
	wire w_dff_A_zgVfTEFh7_0;
	wire w_dff_A_RBWBVSMS7_0;
	wire w_dff_A_S6plSNAH6_0;
	wire w_dff_A_xnV2Ju8e4_0;
	wire w_dff_A_xV84ZD570_0;
	wire w_dff_A_4M3YrL6v0_0;
	wire w_dff_A_OspzlrJ09_0;
	wire w_dff_A_TrPnLkSF3_0;
	wire w_dff_A_PTACoQEj3_0;
	wire w_dff_A_43cg13IY7_0;
	wire w_dff_A_mxq1je1t2_0;
	wire w_dff_A_mS1eXdau5_0;
	wire w_dff_A_nFVETzrZ4_0;
	wire w_dff_A_g4RbweXX6_0;
	wire w_dff_A_ig0ght1b3_0;
	wire w_dff_A_Ouy2aaX18_0;
	wire w_dff_A_Ad33Ftai6_0;
	wire w_dff_A_90WTBUTz0_0;
	wire w_dff_A_cp8oMZvJ2_0;
	wire w_dff_A_uELTC4HS0_0;
	wire w_dff_A_ZZzWmknK8_0;
	wire w_dff_A_5nAuIPLh2_0;
	wire w_dff_A_K3RS4MwB4_0;
	wire w_dff_A_OreutxFh6_0;
	wire w_dff_A_onmFFsOP8_0;
	wire w_dff_A_Qia66mh76_0;
	wire w_dff_A_l2Fdh7NJ8_0;
	wire w_dff_A_FrWsUU4w4_0;
	wire w_dff_A_vZQsEkA11_0;
	wire w_dff_A_5G4NSmpD5_0;
	wire w_dff_A_GCEXWUqS2_0;
	wire w_dff_A_9nHm4XVh8_0;
	wire w_dff_A_ISqqhTi83_0;
	wire w_dff_A_ncqyS2lK9_0;
	wire w_dff_A_zbYCkq4b8_0;
	wire w_dff_A_CpdxpCqa6_0;
	wire w_dff_A_2UAWJVpw0_0;
	wire w_dff_A_dMhJLwUS9_0;
	wire w_dff_A_F4KuuzIG1_0;
	wire w_dff_A_WS4T4fbu6_1;
	wire w_dff_A_SUWXhwpU6_1;
	wire w_dff_A_zFNKhXHj5_1;
	wire w_dff_A_Gp5oCYap9_1;
	wire w_dff_A_mezL70Ep5_2;
	wire w_dff_A_mvPXw4ex2_2;
	wire w_dff_A_kSrOh2pl4_2;
	wire w_dff_A_KfhzSFjL0_2;
	wire w_dff_A_SrQ33Zs43_1;
	wire w_dff_A_ayBzVqxe7_0;
	wire w_dff_A_OsCJGy7G5_0;
	wire w_dff_A_hDykUPTt6_0;
	wire w_dff_A_YOr88fZs6_0;
	wire w_dff_A_9Hicxlfj6_0;
	wire w_dff_A_S5kaVC0d6_0;
	wire w_dff_A_r5f02Pg75_0;
	wire w_dff_A_27OZu5vy8_0;
	wire w_dff_A_udL76qcW8_0;
	wire w_dff_A_XsVLztRM6_0;
	wire w_dff_A_pAWR0Zxn2_0;
	wire w_dff_A_G3o4Gvh99_0;
	wire w_dff_A_tB46nrLl9_0;
	wire w_dff_A_xsUikkql9_0;
	wire w_dff_A_MgOuSpVs7_0;
	wire w_dff_A_LG73gyN70_0;
	wire w_dff_A_beARBm5V2_0;
	wire w_dff_A_fqWoQ2uE2_0;
	wire w_dff_A_mHsqquK34_0;
	wire w_dff_A_6EJUutyz5_0;
	wire w_dff_A_dlCRRlbm7_0;
	wire w_dff_A_3MpTAxUU5_0;
	wire w_dff_A_MevaaZEz8_0;
	wire w_dff_A_Ae7ctVL45_0;
	wire w_dff_A_WBqiegTa1_0;
	wire w_dff_A_pqxqYhxx6_0;
	wire w_dff_A_1TtFD5TO2_0;
	wire w_dff_A_wBNhqVY15_0;
	wire w_dff_A_h3OHrec87_0;
	wire w_dff_A_XdLnXq9U9_0;
	wire w_dff_A_aPbx6nzc7_0;
	wire w_dff_A_RZklojRm9_0;
	wire w_dff_A_sFEORtIR9_0;
	wire w_dff_A_uRBDuVzz8_0;
	wire w_dff_A_fQ2piNSh3_0;
	wire w_dff_A_eC98ewXI3_0;
	wire w_dff_A_tJ5moZB72_0;
	wire w_dff_A_iY7kSZQQ6_0;
	wire w_dff_A_31zVupeu1_0;
	wire w_dff_A_njhaywae7_0;
	wire w_dff_A_3vEXTt2O5_0;
	wire w_dff_A_pvZffa4Y3_0;
	wire w_dff_A_wV9dlqrx8_0;
	wire w_dff_A_OsoCbngY1_0;
	wire w_dff_A_J9Y53Guw0_0;
	wire w_dff_A_qdaMsgC00_0;
	wire w_dff_A_qYOVCnRs3_0;
	wire w_dff_A_JDbXe0Kk6_0;
	wire w_dff_A_fp8Lhak87_0;
	wire w_dff_A_DqsI2tef5_0;
	wire w_dff_A_5Id62eyV1_0;
	wire w_dff_A_RPzDK8EP9_0;
	wire w_dff_A_DqR24QHW6_0;
	wire w_dff_A_eofqEATT6_0;
	wire w_dff_A_u9t5AbKR6_0;
	wire w_dff_A_VU4fVyCB1_0;
	wire w_dff_A_GhMeJAU66_0;
	wire w_dff_A_7sIksdo32_0;
	wire w_dff_A_A4MTaJyG7_0;
	wire w_dff_A_T6jDC0ny1_0;
	wire w_dff_A_Y6aytHgg7_0;
	wire w_dff_A_tgBk6IEc0_0;
	wire w_dff_A_lMuE5vKe9_0;
	wire w_dff_A_FRBlaDhn3_0;
	wire w_dff_A_ifgivyBk4_0;
	wire w_dff_A_uA7972LX0_0;
	wire w_dff_A_u7SSCR2M0_0;
	wire w_dff_A_qtAlqtt74_0;
	wire w_dff_A_LWqr1tJp3_0;
	wire w_dff_A_Ly6vFl2o1_0;
	wire w_dff_A_CEkfR8YQ4_0;
	wire w_dff_A_o9mQOxpV7_0;
	wire w_dff_A_Ny2axnXR6_0;
	wire w_dff_A_G30zSihx9_0;
	wire w_dff_A_4i5VYRsY1_0;
	wire w_dff_A_goQn8Qyb4_0;
	wire w_dff_A_iNp35z6R9_0;
	wire w_dff_A_maScKN3y1_0;
	wire w_dff_A_OAFdzDG37_0;
	wire w_dff_A_MjaR1rzo9_0;
	wire w_dff_A_ACiX3UiA0_0;
	wire w_dff_A_VYfUQqX12_0;
	wire w_dff_A_pUeDmXg80_0;
	wire w_dff_A_gKkyzRf58_0;
	wire w_dff_A_mlCME7o44_0;
	wire w_dff_A_RLZnhZwo1_0;
	wire w_dff_A_ZfYRbZaL8_0;
	wire w_dff_A_H7x4cxRG7_0;
	wire w_dff_A_iqB6IdW90_0;
	wire w_dff_A_FyydgOjX7_0;
	wire w_dff_A_k8h9TTbj5_0;
	wire w_dff_A_dVSuBviO3_0;
	wire w_dff_A_YH8VLY5L1_0;
	wire w_dff_A_fbqP6Ep64_0;
	wire w_dff_A_GaRLcLru9_0;
	wire w_dff_A_fEzr8Q1O8_0;
	wire w_dff_A_GOwmHF5K7_0;
	wire w_dff_A_oG4BV4si9_0;
	wire w_dff_A_Qonvgfhz0_0;
	wire w_dff_A_iNlfX4sN5_0;
	wire w_dff_A_19OnYZKV4_0;
	wire w_dff_A_N5d65ejs1_0;
	wire w_dff_A_vbE2pn4c1_0;
	wire w_dff_A_rjQt1ruS5_0;
	wire w_dff_A_FXMUWy943_0;
	wire w_dff_A_LhFtLdlN9_0;
	wire w_dff_A_YxFBohNB7_0;
	wire w_dff_A_J0Mz2ybJ0_0;
	wire w_dff_A_l7uWztIC1_0;
	wire w_dff_A_swupLrXb5_0;
	wire w_dff_A_SYOKoGYC8_0;
	wire w_dff_A_imZhQM7P7_0;
	wire w_dff_A_KzaP0acl2_0;
	wire w_dff_A_rlQwKjD73_0;
	wire w_dff_A_bSYgqp1s3_0;
	wire w_dff_A_eYIyeTjg8_0;
	wire w_dff_A_SymbD6mv0_2;
	wire w_dff_A_3D6ctpqb9_2;
	wire w_dff_A_GMwuJEWF7_2;
	wire w_dff_A_nxTxlJCZ9_2;
	wire w_dff_A_GU7KRKHU2_2;
	wire w_dff_A_GLtL4owQ8_2;
	wire w_dff_A_p1uJu0Ob8_2;
	wire w_dff_A_VEiGf8yR7_2;
	jnot g000(.din(Gic0),.dout(n73),.clk(gclk));
	jnot g001(.din(Gr),.dout(n74),.clk(gclk));
	jor g002(.dina(w_n74_3[1]),.dinb(n73),.dout(n75),.clk(gclk));
	jxor g003(.dina(w_Gid17_0[2]),.dinb(w_Gid16_0[2]),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_Gid19_0[2]),.dinb(w_Gid18_0[2]),.dout(n77),.clk(gclk));
	jxor g005(.dina(n77),.dinb(n76),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_n78_0[1]),.dinb(n75),.dout(n79),.clk(gclk));
	jxor g007(.dina(w_Gid4_0[2]),.dinb(w_Gid0_0[2]),.dout(n80),.clk(gclk));
	jxor g008(.dina(w_Gid12_0[2]),.dinb(w_Gid8_0[2]),.dout(n81),.clk(gclk));
	jxor g009(.dina(n81),.dinb(n80),.dout(n82),.clk(gclk));
	jxor g010(.dina(w_Gid21_0[2]),.dinb(w_Gid20_0[2]),.dout(n83),.clk(gclk));
	jxor g011(.dina(w_Gid23_0[2]),.dinb(w_Gid22_0[2]),.dout(n84),.clk(gclk));
	jxor g012(.dina(n84),.dinb(n83),.dout(n85),.clk(gclk));
	jxor g013(.dina(w_n85_0[1]),.dinb(n82),.dout(n86),.clk(gclk));
	jxor g014(.dina(n86),.dinb(n79),.dout(n87),.clk(gclk));
	jnot g015(.din(w_n87_1[1]),.dout(n88),.clk(gclk));
	jnot g016(.din(Gic7),.dout(n89),.clk(gclk));
	jor g017(.dina(w_n74_3[0]),.dinb(n89),.dout(n90),.clk(gclk));
	jxor g018(.dina(w_Gid5_0[2]),.dinb(w_Gid4_0[1]),.dout(n91),.clk(gclk));
	jxor g019(.dina(w_Gid7_0[2]),.dinb(w_Gid6_0[2]),.dout(n92),.clk(gclk));
	jxor g020(.dina(n92),.dinb(n91),.dout(n93),.clk(gclk));
	jxor g021(.dina(w_n93_0[1]),.dinb(n90),.dout(n94),.clk(gclk));
	jxor g022(.dina(w_Gid13_0[2]),.dinb(w_Gid12_0[1]),.dout(n95),.clk(gclk));
	jxor g023(.dina(w_Gid15_0[2]),.dinb(w_Gid14_0[2]),.dout(n96),.clk(gclk));
	jxor g024(.dina(n96),.dinb(n95),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_Gid23_0[1]),.dinb(w_Gid19_0[1]),.dout(n98),.clk(gclk));
	jxor g026(.dina(w_Gid31_0[2]),.dinb(w_Gid27_0[2]),.dout(n99),.clk(gclk));
	jxor g027(.dina(n99),.dinb(n98),.dout(n100),.clk(gclk));
	jxor g028(.dina(n100),.dinb(w_n97_0[1]),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n94),.dout(n102),.clk(gclk));
	jnot g030(.din(Gic6),.dout(n103),.clk(gclk));
	jor g031(.dina(w_n74_2[2]),.dinb(n103),.dout(n104),.clk(gclk));
	jxor g032(.dina(w_Gid1_0[2]),.dinb(w_Gid0_0[1]),.dout(n105),.clk(gclk));
	jxor g033(.dina(w_Gid3_0[2]),.dinb(w_Gid2_0[2]),.dout(n106),.clk(gclk));
	jxor g034(.dina(n106),.dinb(n105),.dout(n107),.clk(gclk));
	jxor g035(.dina(w_n107_0[1]),.dinb(n104),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_Gid9_0[2]),.dinb(w_Gid8_0[1]),.dout(n109),.clk(gclk));
	jxor g037(.dina(w_Gid11_0[2]),.dinb(w_Gid10_0[2]),.dout(n110),.clk(gclk));
	jxor g038(.dina(n110),.dinb(n109),.dout(n111),.clk(gclk));
	jxor g039(.dina(w_Gid22_0[1]),.dinb(w_Gid18_0[1]),.dout(n112),.clk(gclk));
	jxor g040(.dina(w_Gid30_0[2]),.dinb(w_Gid26_0[2]),.dout(n113),.clk(gclk));
	jxor g041(.dina(n113),.dinb(n112),.dout(n114),.clk(gclk));
	jxor g042(.dina(n114),.dinb(w_n111_0[1]),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(n108),.dout(n116),.clk(gclk));
	jnot g044(.din(w_n116_1[1]),.dout(n117),.clk(gclk));
	jand g045(.dina(w_n117_1[2]),.dinb(w_n102_1[1]),.dout(n118),.clk(gclk));
	jnot g046(.din(Gic4),.dout(n119),.clk(gclk));
	jor g047(.dina(w_n74_2[1]),.dinb(n119),.dout(n120),.clk(gclk));
	jxor g048(.dina(n120),.dinb(w_n93_0[0]),.dout(n121),.clk(gclk));
	jxor g049(.dina(w_Gid20_0[1]),.dinb(w_Gid16_0[1]),.dout(n122),.clk(gclk));
	jxor g050(.dina(w_Gid28_0[2]),.dinb(w_Gid24_0[2]),.dout(n123),.clk(gclk));
	jxor g051(.dina(n123),.dinb(n122),.dout(n124),.clk(gclk));
	jxor g052(.dina(n124),.dinb(w_n107_0[0]),.dout(n125),.clk(gclk));
	jxor g053(.dina(n125),.dinb(n121),.dout(n126),.clk(gclk));
	jnot g054(.din(w_n126_1[1]),.dout(n127),.clk(gclk));
	jnot g055(.din(Gic5),.dout(n128),.clk(gclk));
	jor g056(.dina(w_n74_2[0]),.dinb(n128),.dout(n129),.clk(gclk));
	jxor g057(.dina(n129),.dinb(w_n97_0[0]),.dout(n130),.clk(gclk));
	jxor g058(.dina(w_Gid21_0[1]),.dinb(w_Gid17_0[1]),.dout(n131),.clk(gclk));
	jxor g059(.dina(w_Gid29_0[2]),.dinb(w_Gid25_0[2]),.dout(n132),.clk(gclk));
	jxor g060(.dina(n132),.dinb(n131),.dout(n133),.clk(gclk));
	jxor g061(.dina(n133),.dinb(w_n111_0[0]),.dout(n134),.clk(gclk));
	jxor g062(.dina(n134),.dinb(n130),.dout(n135),.clk(gclk));
	jand g063(.dina(w_n135_1[1]),.dinb(w_n127_1[2]),.dout(n136),.clk(gclk));
	jnot g064(.din(Gic1),.dout(n137),.clk(gclk));
	jor g065(.dina(w_n74_1[2]),.dinb(n137),.dout(n138),.clk(gclk));
	jxor g066(.dina(w_Gid29_0[1]),.dinb(w_Gid28_0[1]),.dout(n139),.clk(gclk));
	jxor g067(.dina(w_Gid31_0[1]),.dinb(w_Gid30_0[1]),.dout(n140),.clk(gclk));
	jxor g068(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g069(.dina(w_n141_0[1]),.dinb(n138),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_Gid25_0[1]),.dinb(w_Gid24_0[1]),.dout(n143),.clk(gclk));
	jxor g071(.dina(w_Gid27_0[1]),.dinb(w_Gid26_0[1]),.dout(n144),.clk(gclk));
	jxor g072(.dina(n144),.dinb(n143),.dout(n145),.clk(gclk));
	jxor g073(.dina(w_Gid5_0[1]),.dinb(w_Gid1_0[1]),.dout(n146),.clk(gclk));
	jxor g074(.dina(w_Gid13_0[1]),.dinb(w_Gid9_0[1]),.dout(n147),.clk(gclk));
	jxor g075(.dina(n147),.dinb(n146),.dout(n148),.clk(gclk));
	jxor g076(.dina(n148),.dinb(w_n145_0[1]),.dout(n149),.clk(gclk));
	jxor g077(.dina(n149),.dinb(n142),.dout(n150),.clk(gclk));
	jxor g078(.dina(w_n150_1[1]),.dinb(w_n87_1[0]),.dout(n151),.clk(gclk));
	jnot g079(.din(Gic3),.dout(n152),.clk(gclk));
	jor g080(.dina(w_n74_1[1]),.dinb(n152),.dout(n153),.clk(gclk));
	jxor g081(.dina(n153),.dinb(w_n85_0[0]),.dout(n154),.clk(gclk));
	jxor g082(.dina(w_Gid7_0[1]),.dinb(w_Gid3_0[1]),.dout(n155),.clk(gclk));
	jxor g083(.dina(w_Gid15_0[1]),.dinb(w_Gid11_0[1]),.dout(n156),.clk(gclk));
	jxor g084(.dina(n156),.dinb(n155),.dout(n157),.clk(gclk));
	jxor g085(.dina(n157),.dinb(w_n141_0[0]),.dout(n158),.clk(gclk));
	jxor g086(.dina(n158),.dinb(n154),.dout(n159),.clk(gclk));
	jnot g087(.din(Gic2),.dout(n160),.clk(gclk));
	jor g088(.dina(w_n74_1[0]),.dinb(n160),.dout(n161),.clk(gclk));
	jxor g089(.dina(n161),.dinb(w_n78_0[0]),.dout(n162),.clk(gclk));
	jxor g090(.dina(w_Gid6_0[1]),.dinb(w_Gid2_0[1]),.dout(n163),.clk(gclk));
	jxor g091(.dina(w_Gid14_0[1]),.dinb(w_Gid10_0[1]),.dout(n164),.clk(gclk));
	jxor g092(.dina(n164),.dinb(n163),.dout(n165),.clk(gclk));
	jxor g093(.dina(n165),.dinb(w_n145_0[0]),.dout(n166),.clk(gclk));
	jxor g094(.dina(n166),.dinb(n162),.dout(n167),.clk(gclk));
	jand g095(.dina(w_n167_1[1]),.dinb(w_n159_1[1]),.dout(n168),.clk(gclk));
	jand g096(.dina(n168),.dinb(n151),.dout(n169),.clk(gclk));
	jxor g097(.dina(w_n167_1[0]),.dinb(w_n159_1[0]),.dout(n170),.clk(gclk));
	jand g098(.dina(w_n150_1[0]),.dinb(w_n87_0[2]),.dout(n171),.clk(gclk));
	jand g099(.dina(n171),.dinb(n170),.dout(n172),.clk(gclk));
	jor g100(.dina(n172),.dinb(n169),.dout(n173),.clk(gclk));
	jand g101(.dina(w_n173_0[2]),.dinb(w_dff_B_zLnaYhAk3_1),.dout(n174),.clk(gclk));
	jand g102(.dina(w_n174_0[1]),.dinb(w_n118_0[1]),.dout(n175),.clk(gclk));
	jand g103(.dina(w_n175_1[1]),.dinb(w_n88_1[2]),.dout(n176),.clk(gclk));
	jxor g104(.dina(n176),.dinb(w_Gid0_0[0]),.dout(God0),.clk(gclk));
	jnot g105(.din(w_n150_0[2]),.dout(n178),.clk(gclk));
	jand g106(.dina(w_n175_1[0]),.dinb(w_n178_1[2]),.dout(n179),.clk(gclk));
	jxor g107(.dina(n179),.dinb(w_Gid1_0[0]),.dout(God1),.clk(gclk));
	jnot g108(.din(w_n167_0[2]),.dout(n181),.clk(gclk));
	jand g109(.dina(w_n175_0[2]),.dinb(w_n181_1[2]),.dout(n182),.clk(gclk));
	jxor g110(.dina(n182),.dinb(w_Gid2_0[0]),.dout(God2),.clk(gclk));
	jnot g111(.din(w_n159_0[2]),.dout(n184),.clk(gclk));
	jand g112(.dina(w_n175_0[1]),.dinb(w_n184_1[2]),.dout(n185),.clk(gclk));
	jxor g113(.dina(n185),.dinb(w_Gid3_0[0]),.dout(God3),.clk(gclk));
	jnot g114(.din(w_n102_1[0]),.dout(n187),.clk(gclk));
	jand g115(.dina(w_n116_1[0]),.dinb(w_n187_1[2]),.dout(n188),.clk(gclk));
	jand g116(.dina(w_n188_0[1]),.dinb(w_n174_0[0]),.dout(n189),.clk(gclk));
	jand g117(.dina(w_n189_1[1]),.dinb(w_n88_1[1]),.dout(n190),.clk(gclk));
	jxor g118(.dina(n190),.dinb(w_Gid4_0[0]),.dout(God4),.clk(gclk));
	jand g119(.dina(w_n189_1[0]),.dinb(w_n178_1[1]),.dout(n192),.clk(gclk));
	jxor g120(.dina(n192),.dinb(w_Gid5_0[0]),.dout(God5),.clk(gclk));
	jand g121(.dina(w_n189_0[2]),.dinb(w_n181_1[1]),.dout(n194),.clk(gclk));
	jxor g122(.dina(n194),.dinb(w_Gid6_0[0]),.dout(God6),.clk(gclk));
	jand g123(.dina(w_n189_0[1]),.dinb(w_n184_1[1]),.dout(n196),.clk(gclk));
	jxor g124(.dina(n196),.dinb(w_Gid7_0[0]),.dout(God7),.clk(gclk));
	jnot g125(.din(w_n135_1[0]),.dout(n198),.clk(gclk));
	jand g126(.dina(w_n198_1[2]),.dinb(w_n126_1[0]),.dout(n199),.clk(gclk));
	jand g127(.dina(w_n199_0[1]),.dinb(w_n118_0[0]),.dout(n200),.clk(gclk));
	jand g128(.dina(n200),.dinb(w_n173_0[1]),.dout(n201),.clk(gclk));
	jand g129(.dina(w_n201_1[1]),.dinb(w_n88_1[0]),.dout(n202),.clk(gclk));
	jxor g130(.dina(n202),.dinb(w_Gid8_0[0]),.dout(w_dff_A_SymbD6mv0_2),.clk(gclk));
	jand g131(.dina(w_n201_1[0]),.dinb(w_n178_1[0]),.dout(n204),.clk(gclk));
	jxor g132(.dina(n204),.dinb(w_Gid9_0[0]),.dout(w_dff_A_3D6ctpqb9_2),.clk(gclk));
	jand g133(.dina(w_n201_0[2]),.dinb(w_n181_1[0]),.dout(n206),.clk(gclk));
	jxor g134(.dina(n206),.dinb(w_Gid10_0[0]),.dout(w_dff_A_GMwuJEWF7_2),.clk(gclk));
	jand g135(.dina(w_n201_0[1]),.dinb(w_n184_1[0]),.dout(n208),.clk(gclk));
	jxor g136(.dina(n208),.dinb(w_Gid11_0[0]),.dout(w_dff_A_nxTxlJCZ9_2),.clk(gclk));
	jand g137(.dina(w_n199_0[0]),.dinb(w_n188_0[0]),.dout(n210),.clk(gclk));
	jand g138(.dina(n210),.dinb(w_n173_0[0]),.dout(n211),.clk(gclk));
	jand g139(.dina(w_n211_1[1]),.dinb(w_n88_0[2]),.dout(n212),.clk(gclk));
	jxor g140(.dina(n212),.dinb(w_Gid12_0[0]),.dout(w_dff_A_GU7KRKHU2_2),.clk(gclk));
	jand g141(.dina(w_n211_1[0]),.dinb(w_n178_0[2]),.dout(n214),.clk(gclk));
	jxor g142(.dina(n214),.dinb(w_Gid13_0[0]),.dout(w_dff_A_GLtL4owQ8_2),.clk(gclk));
	jand g143(.dina(w_n211_0[2]),.dinb(w_n181_0[2]),.dout(n216),.clk(gclk));
	jxor g144(.dina(n216),.dinb(w_Gid14_0[0]),.dout(w_dff_A_p1uJu0Ob8_2),.clk(gclk));
	jand g145(.dina(w_n211_0[1]),.dinb(w_n184_0[2]),.dout(n218),.clk(gclk));
	jxor g146(.dina(n218),.dinb(w_Gid15_0[0]),.dout(w_dff_A_VEiGf8yR7_2),.clk(gclk));
	jand g147(.dina(w_n150_0[1]),.dinb(w_n88_0[1]),.dout(n220),.clk(gclk));
	jand g148(.dina(w_n181_0[1]),.dinb(w_n159_0[1]),.dout(n221),.clk(gclk));
	jxor g149(.dina(w_n116_0[2]),.dinb(w_n102_0[2]),.dout(n222),.clk(gclk));
	jand g150(.dina(w_n135_0[2]),.dinb(w_n126_0[2]),.dout(n223),.clk(gclk));
	jand g151(.dina(n223),.dinb(n222),.dout(n224),.clk(gclk));
	jxor g152(.dina(w_n135_0[1]),.dinb(w_n126_0[1]),.dout(n225),.clk(gclk));
	jand g153(.dina(w_n116_0[1]),.dinb(w_n102_0[1]),.dout(n226),.clk(gclk));
	jand g154(.dina(n226),.dinb(n225),.dout(n227),.clk(gclk));
	jor g155(.dina(n227),.dinb(n224),.dout(n228),.clk(gclk));
	jand g156(.dina(w_n228_0[1]),.dinb(w_dff_B_LnPM9yPY5_1),.dout(n229),.clk(gclk));
	jand g157(.dina(w_n229_0[1]),.dinb(w_n220_0[1]),.dout(n230),.clk(gclk));
	jand g158(.dina(w_n230_1[1]),.dinb(w_n127_1[1]),.dout(n231),.clk(gclk));
	jxor g159(.dina(n231),.dinb(w_Gid16_0[0]),.dout(God16),.clk(gclk));
	jand g160(.dina(w_n230_1[0]),.dinb(w_n198_1[1]),.dout(n233),.clk(gclk));
	jxor g161(.dina(n233),.dinb(w_Gid17_0[0]),.dout(God17),.clk(gclk));
	jand g162(.dina(w_n230_0[2]),.dinb(w_n117_1[1]),.dout(n235),.clk(gclk));
	jxor g163(.dina(n235),.dinb(w_Gid18_0[0]),.dout(God18),.clk(gclk));
	jand g164(.dina(w_n230_0[1]),.dinb(w_n187_1[1]),.dout(n237),.clk(gclk));
	jxor g165(.dina(n237),.dinb(w_Gid19_0[0]),.dout(God19),.clk(gclk));
	jand g166(.dina(w_n167_0[1]),.dinb(w_n184_0[1]),.dout(n239),.clk(gclk));
	jand g167(.dina(w_n228_0[0]),.dinb(w_dff_B_e93qed7n2_1),.dout(n240),.clk(gclk));
	jand g168(.dina(w_n240_0[1]),.dinb(w_n220_0[0]),.dout(n241),.clk(gclk));
	jand g169(.dina(w_n241_1[1]),.dinb(w_n127_1[0]),.dout(n242),.clk(gclk));
	jxor g170(.dina(n242),.dinb(w_Gid20_0[0]),.dout(God20),.clk(gclk));
	jand g171(.dina(w_n241_1[0]),.dinb(w_n198_1[0]),.dout(n244),.clk(gclk));
	jxor g172(.dina(n244),.dinb(w_Gid21_0[0]),.dout(God21),.clk(gclk));
	jand g173(.dina(w_n241_0[2]),.dinb(w_n117_1[0]),.dout(n246),.clk(gclk));
	jxor g174(.dina(n246),.dinb(w_Gid22_0[0]),.dout(God22),.clk(gclk));
	jand g175(.dina(w_n241_0[1]),.dinb(w_n187_1[0]),.dout(n248),.clk(gclk));
	jxor g176(.dina(n248),.dinb(w_Gid23_0[0]),.dout(God23),.clk(gclk));
	jand g177(.dina(w_n178_0[1]),.dinb(w_n87_0[1]),.dout(n250),.clk(gclk));
	jand g178(.dina(w_n229_0[0]),.dinb(w_n250_0[1]),.dout(n251),.clk(gclk));
	jand g179(.dina(w_n251_1[1]),.dinb(w_n127_0[2]),.dout(n252),.clk(gclk));
	jxor g180(.dina(n252),.dinb(w_Gid24_0[0]),.dout(God24),.clk(gclk));
	jand g181(.dina(w_n251_1[0]),.dinb(w_n198_0[2]),.dout(n254),.clk(gclk));
	jxor g182(.dina(n254),.dinb(w_Gid25_0[0]),.dout(God25),.clk(gclk));
	jand g183(.dina(w_n251_0[2]),.dinb(w_n117_0[2]),.dout(n256),.clk(gclk));
	jxor g184(.dina(n256),.dinb(w_Gid26_0[0]),.dout(God26),.clk(gclk));
	jand g185(.dina(w_n251_0[1]),.dinb(w_n187_0[2]),.dout(n258),.clk(gclk));
	jxor g186(.dina(n258),.dinb(w_Gid27_0[0]),.dout(God27),.clk(gclk));
	jand g187(.dina(w_n240_0[0]),.dinb(w_n250_0[0]),.dout(n260),.clk(gclk));
	jand g188(.dina(w_n260_1[1]),.dinb(w_n127_0[1]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_Gid28_0[0]),.dout(God28),.clk(gclk));
	jand g190(.dina(w_n260_1[0]),.dinb(w_n198_0[1]),.dout(n263),.clk(gclk));
	jxor g191(.dina(n263),.dinb(w_Gid29_0[0]),.dout(God29),.clk(gclk));
	jand g192(.dina(w_n260_0[2]),.dinb(w_n117_0[1]),.dout(n265),.clk(gclk));
	jxor g193(.dina(n265),.dinb(w_Gid30_0[0]),.dout(God30),.clk(gclk));
	jand g194(.dina(w_n260_0[1]),.dinb(w_n187_0[1]),.dout(n267),.clk(gclk));
	jxor g195(.dina(n267),.dinb(w_Gid31_0[0]),.dout(God31),.clk(gclk));
	jspl3 jspl3_w_Gid0_0(.douta(w_dff_A_PTACoQEj3_0),.doutb(w_Gid0_0[1]),.doutc(w_Gid0_0[2]),.din(Gid0));
	jspl3 jspl3_w_Gid1_0(.douta(w_dff_A_zjbSdnLV9_0),.doutb(w_Gid1_0[1]),.doutc(w_Gid1_0[2]),.din(Gid1));
	jspl3 jspl3_w_Gid2_0(.douta(w_dff_A_qJXJclC73_0),.doutb(w_Gid2_0[1]),.doutc(w_Gid2_0[2]),.din(Gid2));
	jspl3 jspl3_w_Gid3_0(.douta(w_dff_A_F9swWSKi8_0),.doutb(w_Gid3_0[1]),.doutc(w_Gid3_0[2]),.din(Gid3));
	jspl3 jspl3_w_Gid4_0(.douta(w_dff_A_eYIyeTjg8_0),.doutb(w_Gid4_0[1]),.doutc(w_Gid4_0[2]),.din(Gid4));
	jspl3 jspl3_w_Gid5_0(.douta(w_dff_A_LhFtLdlN9_0),.doutb(w_Gid5_0[1]),.doutc(w_Gid5_0[2]),.din(Gid5));
	jspl3 jspl3_w_Gid6_0(.douta(w_dff_A_fEzr8Q1O8_0),.doutb(w_Gid6_0[1]),.doutc(w_Gid6_0[2]),.din(Gid6));
	jspl3 jspl3_w_Gid7_0(.douta(w_dff_A_RLZnhZwo1_0),.doutb(w_Gid7_0[1]),.doutc(w_Gid7_0[2]),.din(Gid7));
	jspl3 jspl3_w_Gid8_0(.douta(w_dff_A_h0Czj1or7_0),.doutb(w_Gid8_0[1]),.doutc(w_Gid8_0[2]),.din(Gid8));
	jspl3 jspl3_w_Gid9_0(.douta(w_dff_A_WcyjloGZ2_0),.doutb(w_Gid9_0[1]),.doutc(w_Gid9_0[2]),.din(Gid9));
	jspl3 jspl3_w_Gid10_0(.douta(w_dff_A_5ycgIj5v7_0),.doutb(w_Gid10_0[1]),.doutc(w_Gid10_0[2]),.din(Gid10));
	jspl3 jspl3_w_Gid11_0(.douta(w_dff_A_7tleaXJX8_0),.doutb(w_Gid11_0[1]),.doutc(w_Gid11_0[2]),.din(Gid11));
	jspl3 jspl3_w_Gid12_0(.douta(w_dff_A_goQn8Qyb4_0),.doutb(w_Gid12_0[1]),.doutc(w_Gid12_0[2]),.din(Gid12));
	jspl3 jspl3_w_Gid13_0(.douta(w_dff_A_u7SSCR2M0_0),.doutb(w_Gid13_0[1]),.doutc(w_Gid13_0[2]),.din(Gid13));
	jspl3 jspl3_w_Gid14_0(.douta(w_dff_A_7sIksdo32_0),.doutb(w_Gid14_0[1]),.doutc(w_Gid14_0[2]),.din(Gid14));
	jspl3 jspl3_w_Gid15_0(.douta(w_dff_A_fp8Lhak87_0),.doutb(w_Gid15_0[1]),.doutc(w_Gid15_0[2]),.din(Gid15));
	jspl3 jspl3_w_Gid16_0(.douta(w_dff_A_F4KuuzIG1_0),.doutb(w_Gid16_0[1]),.doutc(w_Gid16_0[2]),.din(Gid16));
	jspl3 jspl3_w_Gid17_0(.douta(w_dff_A_vZQsEkA11_0),.doutb(w_Gid17_0[1]),.doutc(w_Gid17_0[2]),.din(Gid17));
	jspl3 jspl3_w_Gid18_0(.douta(w_dff_A_cp8oMZvJ2_0),.doutb(w_Gid18_0[1]),.doutc(w_Gid18_0[2]),.din(Gid18));
	jspl3 jspl3_w_Gid19_0(.douta(w_dff_A_njhaywae7_0),.doutb(w_Gid19_0[1]),.doutc(w_Gid19_0[2]),.din(Gid19));
	jspl3 jspl3_w_Gid20_0(.douta(w_dff_A_dfvbAn5o2_0),.doutb(w_Gid20_0[1]),.doutc(w_Gid20_0[2]),.din(Gid20));
	jspl3 jspl3_w_Gid21_0(.douta(w_dff_A_p6PpfRME7_0),.doutb(w_Gid21_0[1]),.doutc(w_Gid21_0[2]),.din(Gid21));
	jspl3 jspl3_w_Gid22_0(.douta(w_dff_A_ZVPfoTQT1_0),.doutb(w_Gid22_0[1]),.doutc(w_Gid22_0[2]),.din(Gid22));
	jspl3 jspl3_w_Gid23_0(.douta(w_dff_A_XdLnXq9U9_0),.doutb(w_Gid23_0[1]),.doutc(w_Gid23_0[2]),.din(Gid23));
	jspl3 jspl3_w_Gid24_0(.douta(w_dff_A_qlllOe9G5_0),.doutb(w_Gid24_0[1]),.doutc(w_Gid24_0[2]),.din(Gid24));
	jspl3 jspl3_w_Gid25_0(.douta(w_dff_A_1A0bEObr3_0),.doutb(w_Gid25_0[1]),.doutc(w_Gid25_0[2]),.din(Gid25));
	jspl3 jspl3_w_Gid26_0(.douta(w_dff_A_OvZnt1XA4_0),.doutb(w_Gid26_0[1]),.doutc(w_Gid26_0[2]),.din(Gid26));
	jspl3 jspl3_w_Gid27_0(.douta(w_dff_A_6EJUutyz5_0),.doutb(w_Gid27_0[1]),.doutc(w_Gid27_0[2]),.din(Gid27));
	jspl3 jspl3_w_Gid28_0(.douta(w_dff_A_4mvnpGSs4_0),.doutb(w_Gid28_0[1]),.doutc(w_Gid28_0[2]),.din(Gid28));
	jspl3 jspl3_w_Gid29_0(.douta(w_dff_A_IIherzhR4_0),.doutb(w_Gid29_0[1]),.doutc(w_Gid29_0[2]),.din(Gid29));
	jspl3 jspl3_w_Gid30_0(.douta(w_dff_A_ZCxqcaoc6_0),.doutb(w_Gid30_0[1]),.doutc(w_Gid30_0[2]),.din(Gid30));
	jspl3 jspl3_w_Gid31_0(.douta(w_dff_A_XsVLztRM6_0),.doutb(w_Gid31_0[1]),.doutc(w_Gid31_0[2]),.din(Gid31));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl3 jspl3_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.doutc(w_n74_1[2]),.din(w_n74_0[0]));
	jspl3 jspl3_w_n74_2(.douta(w_n74_2[0]),.doutb(w_n74_2[1]),.doutc(w_n74_2[2]),.din(w_n74_0[1]));
	jspl jspl_w_n74_3(.douta(w_n74_3[0]),.doutb(w_n74_3[1]),.din(w_n74_0[2]));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl3 jspl3_w_n87_0(.douta(w_n87_0[0]),.doutb(w_dff_A_M2PaOgjg4_1),.doutc(w_n87_0[2]),.din(n87));
	jspl jspl_w_n87_1(.douta(w_n87_1[0]),.doutb(w_n87_1[1]),.din(w_n87_0[0]));
	jspl3 jspl3_w_n88_0(.douta(w_dff_A_hL8dYl2p6_0),.doutb(w_n88_0[1]),.doutc(w_dff_A_xj9ez3eS0_2),.din(n88));
	jspl3 jspl3_w_n88_1(.douta(w_n88_1[0]),.doutb(w_dff_A_ncZ1c8Jf5_1),.doutc(w_dff_A_2EossxO28_2),.din(w_n88_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl3 jspl3_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.doutc(w_n102_0[2]),.din(n102));
	jspl jspl_w_n102_1(.douta(w_n102_1[0]),.doutb(w_dff_A_SrQ33Zs43_1),.din(w_n102_0[0]));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.doutc(w_n116_0[2]),.din(n116));
	jspl jspl_w_n116_1(.douta(w_dff_A_e0deb75v8_0),.doutb(w_n116_1[1]),.din(w_n116_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_rijR7ckf2_1),.doutc(w_dff_A_BAk5pbYc4_2),.din(n117));
	jspl3 jspl3_w_n117_1(.douta(w_dff_A_8NCA6Alt8_0),.doutb(w_dff_A_VhyRl4SB1_1),.doutc(w_n117_1[2]),.din(w_n117_0[0]));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_dff_A_aj31bKFg6_1),.din(n118));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl jspl_w_n126_1(.douta(w_dff_A_Ljjz6T0o5_0),.doutb(w_n126_1[1]),.din(w_n126_0[0]));
	jspl3 jspl3_w_n127_0(.douta(w_n127_0[0]),.doutb(w_dff_A_HVPAQLgR8_1),.doutc(w_dff_A_AECdvskk8_2),.din(n127));
	jspl3 jspl3_w_n127_1(.douta(w_dff_A_yGPBCphy2_0),.doutb(w_dff_A_qcxs7akv1_1),.doutc(w_n127_1[2]),.din(w_n127_0[0]));
	jspl3 jspl3_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.doutc(w_n135_0[2]),.din(n135));
	jspl jspl_w_n135_1(.douta(w_n135_1[0]),.doutb(w_dff_A_YUTr4cZx2_1),.din(w_n135_0[0]));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl3 jspl3_w_n150_0(.douta(w_n150_0[0]),.doutb(w_dff_A_L009HIxL8_1),.doutc(w_n150_0[2]),.din(n150));
	jspl jspl_w_n150_1(.douta(w_n150_1[0]),.doutb(w_n150_1[1]),.din(w_n150_0[0]));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_dff_A_s6EPuhFG3_1),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_dff_A_Zixou12u7_1),.doutc(w_n167_0[2]),.din(n167));
	jspl jspl_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.din(n174));
	jspl3 jspl3_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.doutc(w_n175_0[2]),.din(n175));
	jspl jspl_w_n175_1(.douta(w_n175_1[0]),.doutb(w_n175_1[1]),.din(w_n175_0[0]));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_JXsgy0qd6_0),.doutb(w_n178_0[1]),.doutc(w_dff_A_m0QOCOpM9_2),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_dff_A_CPfiQIe21_1),.doutc(w_dff_A_VQyutGvp7_2),.din(w_n178_0[0]));
	jspl3 jspl3_w_n181_0(.douta(w_dff_A_tAhxaWUj3_0),.doutb(w_n181_0[1]),.doutc(w_dff_A_WSh7d3nm1_2),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_dff_A_KPVIS0wL0_1),.doutc(w_dff_A_ziY5YhhM6_2),.din(w_n181_0[0]));
	jspl3 jspl3_w_n184_0(.douta(w_dff_A_fG3UcLW36_0),.doutb(w_n184_0[1]),.doutc(w_dff_A_up7CYHIQ2_2),.din(n184));
	jspl3 jspl3_w_n184_1(.douta(w_n184_1[0]),.doutb(w_dff_A_168aCpzU1_1),.doutc(w_dff_A_ihKwuW0B4_2),.din(w_n184_0[0]));
	jspl3 jspl3_w_n187_0(.douta(w_n187_0[0]),.doutb(w_dff_A_Gp5oCYap9_1),.doutc(w_dff_A_KfhzSFjL0_2),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_dff_A_dqc5tMAp0_0),.doutb(w_dff_A_z3kZ9A2m7_1),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_dff_A_HzqdGCER1_1),.din(n188));
	jspl3 jspl3_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.doutc(w_n189_0[2]),.din(n189));
	jspl jspl_w_n189_1(.douta(w_n189_1[0]),.doutb(w_n189_1[1]),.din(w_n189_0[0]));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_dff_A_GKF9Xxt81_1),.doutc(w_dff_A_zfN8Qyt76_2),.din(n198));
	jspl3 jspl3_w_n198_1(.douta(w_dff_A_TSQ0bVc40_0),.doutb(w_dff_A_0jOseWON2_1),.doutc(w_n198_1[2]),.din(w_n198_0[0]));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl3 jspl3_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.doutc(w_n201_0[2]),.din(n201));
	jspl jspl_w_n201_1(.douta(w_n201_1[0]),.doutb(w_n201_1[1]),.din(w_n201_0[0]));
	jspl3 jspl3_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.doutc(w_n211_0[2]),.din(n211));
	jspl jspl_w_n211_1(.douta(w_n211_1[0]),.doutb(w_n211_1[1]),.din(w_n211_0[0]));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(w_dff_B_9Qw26Ghh9_2));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.din(n229));
	jspl3 jspl3_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.doutc(w_n230_0[2]),.din(n230));
	jspl jspl_w_n230_1(.douta(w_n230_1[0]),.doutb(w_n230_1[1]),.din(w_n230_0[0]));
	jspl jspl_w_n240_0(.douta(w_n240_0[0]),.doutb(w_n240_0[1]),.din(n240));
	jspl3 jspl3_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.doutc(w_n241_0[2]),.din(n241));
	jspl jspl_w_n241_1(.douta(w_n241_1[0]),.doutb(w_n241_1[1]),.din(w_n241_0[0]));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(w_dff_B_XdS5RqLz8_2));
	jspl3 jspl3_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.doutc(w_n251_0[2]),.din(n251));
	jspl jspl_w_n251_1(.douta(w_n251_1[0]),.doutb(w_n251_1[1]),.din(w_n251_0[0]));
	jspl3 jspl3_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.doutc(w_n260_0[2]),.din(n260));
	jspl jspl_w_n260_1(.douta(w_n260_1[0]),.doutb(w_n260_1[1]),.din(w_n260_0[0]));
	jdff dff_B_zLnaYhAk3_1(.din(n136),.dout(w_dff_B_zLnaYhAk3_1),.clk(gclk));
	jdff dff_A_ncZ1c8Jf5_1(.dout(w_n88_1[1]),.din(w_dff_A_ncZ1c8Jf5_1),.clk(gclk));
	jdff dff_A_2EossxO28_2(.dout(w_n88_1[2]),.din(w_dff_A_2EossxO28_2),.clk(gclk));
	jdff dff_A_CPfiQIe21_1(.dout(w_n178_1[1]),.din(w_dff_A_CPfiQIe21_1),.clk(gclk));
	jdff dff_A_VQyutGvp7_2(.dout(w_n178_1[2]),.din(w_dff_A_VQyutGvp7_2),.clk(gclk));
	jdff dff_A_KPVIS0wL0_1(.dout(w_n181_1[1]),.din(w_dff_A_KPVIS0wL0_1),.clk(gclk));
	jdff dff_A_ziY5YhhM6_2(.dout(w_n181_1[2]),.din(w_dff_A_ziY5YhhM6_2),.clk(gclk));
	jdff dff_A_vaNRwcjV5_1(.dout(w_n118_0[1]),.din(w_dff_A_vaNRwcjV5_1),.clk(gclk));
	jdff dff_A_aj31bKFg6_1(.dout(w_dff_A_vaNRwcjV5_1),.din(w_dff_A_aj31bKFg6_1),.clk(gclk));
	jdff dff_A_168aCpzU1_1(.dout(w_n184_1[1]),.din(w_dff_A_168aCpzU1_1),.clk(gclk));
	jdff dff_A_ihKwuW0B4_2(.dout(w_n184_1[2]),.din(w_dff_A_ihKwuW0B4_2),.clk(gclk));
	jdff dff_A_waxZHvun6_1(.dout(w_n188_0[1]),.din(w_dff_A_waxZHvun6_1),.clk(gclk));
	jdff dff_A_HzqdGCER1_1(.dout(w_dff_A_waxZHvun6_1),.din(w_dff_A_HzqdGCER1_1),.clk(gclk));
	jdff dff_A_p63vZo0A3_0(.dout(w_n127_1[0]),.din(w_dff_A_p63vZo0A3_0),.clk(gclk));
	jdff dff_A_vfU1zxwq9_0(.dout(w_dff_A_p63vZo0A3_0),.din(w_dff_A_vfU1zxwq9_0),.clk(gclk));
	jdff dff_A_ZytrEjEw0_0(.dout(w_dff_A_vfU1zxwq9_0),.din(w_dff_A_ZytrEjEw0_0),.clk(gclk));
	jdff dff_A_yGPBCphy2_0(.dout(w_dff_A_ZytrEjEw0_0),.din(w_dff_A_yGPBCphy2_0),.clk(gclk));
	jdff dff_A_DZ809y9N7_1(.dout(w_n127_1[1]),.din(w_dff_A_DZ809y9N7_1),.clk(gclk));
	jdff dff_A_mwPam5KB4_1(.dout(w_dff_A_DZ809y9N7_1),.din(w_dff_A_mwPam5KB4_1),.clk(gclk));
	jdff dff_A_VAVyDwbQ9_1(.dout(w_dff_A_mwPam5KB4_1),.din(w_dff_A_VAVyDwbQ9_1),.clk(gclk));
	jdff dff_A_qcxs7akv1_1(.dout(w_dff_A_VAVyDwbQ9_1),.din(w_dff_A_qcxs7akv1_1),.clk(gclk));
	jdff dff_A_hCqw5WZ39_0(.dout(w_n198_1[0]),.din(w_dff_A_hCqw5WZ39_0),.clk(gclk));
	jdff dff_A_WoHjTkUS1_0(.dout(w_dff_A_hCqw5WZ39_0),.din(w_dff_A_WoHjTkUS1_0),.clk(gclk));
	jdff dff_A_iOAy8MW69_0(.dout(w_dff_A_WoHjTkUS1_0),.din(w_dff_A_iOAy8MW69_0),.clk(gclk));
	jdff dff_A_TSQ0bVc40_0(.dout(w_dff_A_iOAy8MW69_0),.din(w_dff_A_TSQ0bVc40_0),.clk(gclk));
	jdff dff_A_hDtm3F0v9_1(.dout(w_n198_1[1]),.din(w_dff_A_hDtm3F0v9_1),.clk(gclk));
	jdff dff_A_sptfIzyr5_1(.dout(w_dff_A_hDtm3F0v9_1),.din(w_dff_A_sptfIzyr5_1),.clk(gclk));
	jdff dff_A_ueGalGHp5_1(.dout(w_dff_A_sptfIzyr5_1),.din(w_dff_A_ueGalGHp5_1),.clk(gclk));
	jdff dff_A_0jOseWON2_1(.dout(w_dff_A_ueGalGHp5_1),.din(w_dff_A_0jOseWON2_1),.clk(gclk));
	jdff dff_A_04w2cuD38_0(.dout(w_n117_1[0]),.din(w_dff_A_04w2cuD38_0),.clk(gclk));
	jdff dff_A_m0akYXC16_0(.dout(w_dff_A_04w2cuD38_0),.din(w_dff_A_m0akYXC16_0),.clk(gclk));
	jdff dff_A_3fiVKfNN5_0(.dout(w_dff_A_m0akYXC16_0),.din(w_dff_A_3fiVKfNN5_0),.clk(gclk));
	jdff dff_A_8NCA6Alt8_0(.dout(w_dff_A_3fiVKfNN5_0),.din(w_dff_A_8NCA6Alt8_0),.clk(gclk));
	jdff dff_A_RVMOrcW43_1(.dout(w_n117_1[1]),.din(w_dff_A_RVMOrcW43_1),.clk(gclk));
	jdff dff_A_OHfnjzZ42_1(.dout(w_dff_A_RVMOrcW43_1),.din(w_dff_A_OHfnjzZ42_1),.clk(gclk));
	jdff dff_A_m1bX7gt12_1(.dout(w_dff_A_OHfnjzZ42_1),.din(w_dff_A_m1bX7gt12_1),.clk(gclk));
	jdff dff_A_VhyRl4SB1_1(.dout(w_dff_A_m1bX7gt12_1),.din(w_dff_A_VhyRl4SB1_1),.clk(gclk));
	jdff dff_B_1JtBnWzE5_2(.din(n220),.dout(w_dff_B_1JtBnWzE5_2),.clk(gclk));
	jdff dff_B_9Qw26Ghh9_2(.din(w_dff_B_1JtBnWzE5_2),.dout(w_dff_B_9Qw26Ghh9_2),.clk(gclk));
	jdff dff_A_oCzz8iJF7_0(.dout(w_n88_0[0]),.din(w_dff_A_oCzz8iJF7_0),.clk(gclk));
	jdff dff_A_q1wejxtZ8_0(.dout(w_dff_A_oCzz8iJF7_0),.din(w_dff_A_q1wejxtZ8_0),.clk(gclk));
	jdff dff_A_hL8dYl2p6_0(.dout(w_dff_A_q1wejxtZ8_0),.din(w_dff_A_hL8dYl2p6_0),.clk(gclk));
	jdff dff_A_kYT75gjZ8_2(.dout(w_n88_0[2]),.din(w_dff_A_kYT75gjZ8_2),.clk(gclk));
	jdff dff_A_yzQk7i3X5_2(.dout(w_dff_A_kYT75gjZ8_2),.din(w_dff_A_yzQk7i3X5_2),.clk(gclk));
	jdff dff_A_xj9ez3eS0_2(.dout(w_dff_A_yzQk7i3X5_2),.din(w_dff_A_xj9ez3eS0_2),.clk(gclk));
	jdff dff_A_5y2hzcLU2_0(.dout(w_n187_1[0]),.din(w_dff_A_5y2hzcLU2_0),.clk(gclk));
	jdff dff_A_qYZoe9lW8_0(.dout(w_dff_A_5y2hzcLU2_0),.din(w_dff_A_qYZoe9lW8_0),.clk(gclk));
	jdff dff_A_hUNFsei67_0(.dout(w_dff_A_qYZoe9lW8_0),.din(w_dff_A_hUNFsei67_0),.clk(gclk));
	jdff dff_A_dqc5tMAp0_0(.dout(w_dff_A_hUNFsei67_0),.din(w_dff_A_dqc5tMAp0_0),.clk(gclk));
	jdff dff_A_gWkHxOwb2_1(.dout(w_n187_1[1]),.din(w_dff_A_gWkHxOwb2_1),.clk(gclk));
	jdff dff_A_RLoADiQL6_1(.dout(w_dff_A_gWkHxOwb2_1),.din(w_dff_A_RLoADiQL6_1),.clk(gclk));
	jdff dff_A_NGNee5407_1(.dout(w_dff_A_RLoADiQL6_1),.din(w_dff_A_NGNee5407_1),.clk(gclk));
	jdff dff_A_z3kZ9A2m7_1(.dout(w_dff_A_NGNee5407_1),.din(w_dff_A_z3kZ9A2m7_1),.clk(gclk));
	jdff dff_B_LnPM9yPY5_1(.din(n221),.dout(w_dff_B_LnPM9yPY5_1),.clk(gclk));
	jdff dff_A_iovCjw1W2_0(.dout(w_n181_0[0]),.din(w_dff_A_iovCjw1W2_0),.clk(gclk));
	jdff dff_A_NiL0Jq5Y6_0(.dout(w_dff_A_iovCjw1W2_0),.din(w_dff_A_NiL0Jq5Y6_0),.clk(gclk));
	jdff dff_A_tAhxaWUj3_0(.dout(w_dff_A_NiL0Jq5Y6_0),.din(w_dff_A_tAhxaWUj3_0),.clk(gclk));
	jdff dff_A_xvIr2wzL9_2(.dout(w_n181_0[2]),.din(w_dff_A_xvIr2wzL9_2),.clk(gclk));
	jdff dff_A_xXqfDksf7_2(.dout(w_dff_A_xvIr2wzL9_2),.din(w_dff_A_xXqfDksf7_2),.clk(gclk));
	jdff dff_A_WSh7d3nm1_2(.dout(w_dff_A_xXqfDksf7_2),.din(w_dff_A_WSh7d3nm1_2),.clk(gclk));
	jdff dff_A_2ryBKwmj2_1(.dout(w_n127_0[1]),.din(w_dff_A_2ryBKwmj2_1),.clk(gclk));
	jdff dff_A_qn4MyplS4_1(.dout(w_dff_A_2ryBKwmj2_1),.din(w_dff_A_qn4MyplS4_1),.clk(gclk));
	jdff dff_A_liH1Uy9H7_1(.dout(w_dff_A_qn4MyplS4_1),.din(w_dff_A_liH1Uy9H7_1),.clk(gclk));
	jdff dff_A_HVPAQLgR8_1(.dout(w_dff_A_liH1Uy9H7_1),.din(w_dff_A_HVPAQLgR8_1),.clk(gclk));
	jdff dff_A_sP1QHHi05_2(.dout(w_n127_0[2]),.din(w_dff_A_sP1QHHi05_2),.clk(gclk));
	jdff dff_A_dvobQml51_2(.dout(w_dff_A_sP1QHHi05_2),.din(w_dff_A_dvobQml51_2),.clk(gclk));
	jdff dff_A_NtPfuvxQ8_2(.dout(w_dff_A_dvobQml51_2),.din(w_dff_A_NtPfuvxQ8_2),.clk(gclk));
	jdff dff_A_AECdvskk8_2(.dout(w_dff_A_NtPfuvxQ8_2),.din(w_dff_A_AECdvskk8_2),.clk(gclk));
	jdff dff_A_Ljjz6T0o5_0(.dout(w_n126_1[0]),.din(w_dff_A_Ljjz6T0o5_0),.clk(gclk));
	jdff dff_A_e9yoTzR81_1(.dout(w_n198_0[1]),.din(w_dff_A_e9yoTzR81_1),.clk(gclk));
	jdff dff_A_y9e5IHdq7_1(.dout(w_dff_A_e9yoTzR81_1),.din(w_dff_A_y9e5IHdq7_1),.clk(gclk));
	jdff dff_A_jq3AilBr5_1(.dout(w_dff_A_y9e5IHdq7_1),.din(w_dff_A_jq3AilBr5_1),.clk(gclk));
	jdff dff_A_GKF9Xxt81_1(.dout(w_dff_A_jq3AilBr5_1),.din(w_dff_A_GKF9Xxt81_1),.clk(gclk));
	jdff dff_A_XoLKLvV84_2(.dout(w_n198_0[2]),.din(w_dff_A_XoLKLvV84_2),.clk(gclk));
	jdff dff_A_4B65W6kT7_2(.dout(w_dff_A_XoLKLvV84_2),.din(w_dff_A_4B65W6kT7_2),.clk(gclk));
	jdff dff_A_dz94ukJp1_2(.dout(w_dff_A_4B65W6kT7_2),.din(w_dff_A_dz94ukJp1_2),.clk(gclk));
	jdff dff_A_zfN8Qyt76_2(.dout(w_dff_A_dz94ukJp1_2),.din(w_dff_A_zfN8Qyt76_2),.clk(gclk));
	jdff dff_A_YUTr4cZx2_1(.dout(w_n135_1[1]),.din(w_dff_A_YUTr4cZx2_1),.clk(gclk));
	jdff dff_A_Ck6uPS2X6_1(.dout(w_n117_0[1]),.din(w_dff_A_Ck6uPS2X6_1),.clk(gclk));
	jdff dff_A_1iTlczd10_1(.dout(w_dff_A_Ck6uPS2X6_1),.din(w_dff_A_1iTlczd10_1),.clk(gclk));
	jdff dff_A_mxBeo0iR1_1(.dout(w_dff_A_1iTlczd10_1),.din(w_dff_A_mxBeo0iR1_1),.clk(gclk));
	jdff dff_A_rijR7ckf2_1(.dout(w_dff_A_mxBeo0iR1_1),.din(w_dff_A_rijR7ckf2_1),.clk(gclk));
	jdff dff_A_0t9hgo6Z4_2(.dout(w_n117_0[2]),.din(w_dff_A_0t9hgo6Z4_2),.clk(gclk));
	jdff dff_A_RvJvErBH1_2(.dout(w_dff_A_0t9hgo6Z4_2),.din(w_dff_A_RvJvErBH1_2),.clk(gclk));
	jdff dff_A_WMoCnv7L8_2(.dout(w_dff_A_RvJvErBH1_2),.din(w_dff_A_WMoCnv7L8_2),.clk(gclk));
	jdff dff_A_BAk5pbYc4_2(.dout(w_dff_A_WMoCnv7L8_2),.din(w_dff_A_BAk5pbYc4_2),.clk(gclk));
	jdff dff_A_e0deb75v8_0(.dout(w_n116_1[0]),.din(w_dff_A_e0deb75v8_0),.clk(gclk));
	jdff dff_B_e93qed7n2_1(.din(n239),.dout(w_dff_B_e93qed7n2_1),.clk(gclk));
	jdff dff_A_Zixou12u7_1(.dout(w_n167_0[1]),.din(w_dff_A_Zixou12u7_1),.clk(gclk));
	jdff dff_A_FREWL7EQ4_0(.dout(w_Gid10_0[0]),.din(w_dff_A_FREWL7EQ4_0),.clk(gclk));
	jdff dff_A_r5mUtZ1w0_0(.dout(w_dff_A_FREWL7EQ4_0),.din(w_dff_A_r5mUtZ1w0_0),.clk(gclk));
	jdff dff_A_jXuuHFic2_0(.dout(w_dff_A_r5mUtZ1w0_0),.din(w_dff_A_jXuuHFic2_0),.clk(gclk));
	jdff dff_A_hqdBNAVq0_0(.dout(w_dff_A_jXuuHFic2_0),.din(w_dff_A_hqdBNAVq0_0),.clk(gclk));
	jdff dff_A_LkmloUJ54_0(.dout(w_dff_A_hqdBNAVq0_0),.din(w_dff_A_LkmloUJ54_0),.clk(gclk));
	jdff dff_A_KMUGUlvE4_0(.dout(w_dff_A_LkmloUJ54_0),.din(w_dff_A_KMUGUlvE4_0),.clk(gclk));
	jdff dff_A_0XgOS5ZN1_0(.dout(w_dff_A_KMUGUlvE4_0),.din(w_dff_A_0XgOS5ZN1_0),.clk(gclk));
	jdff dff_A_Qaj5Waxr0_0(.dout(w_dff_A_0XgOS5ZN1_0),.din(w_dff_A_Qaj5Waxr0_0),.clk(gclk));
	jdff dff_A_5ycgIj5v7_0(.dout(w_dff_A_Qaj5Waxr0_0),.din(w_dff_A_5ycgIj5v7_0),.clk(gclk));
	jdff dff_A_T3t3nIWk8_0(.dout(w_Gid2_0[0]),.din(w_dff_A_T3t3nIWk8_0),.clk(gclk));
	jdff dff_A_rvnDP1ph8_0(.dout(w_dff_A_T3t3nIWk8_0),.din(w_dff_A_rvnDP1ph8_0),.clk(gclk));
	jdff dff_A_Cc9KnMvu6_0(.dout(w_dff_A_rvnDP1ph8_0),.din(w_dff_A_Cc9KnMvu6_0),.clk(gclk));
	jdff dff_A_BFT77zb42_0(.dout(w_dff_A_Cc9KnMvu6_0),.din(w_dff_A_BFT77zb42_0),.clk(gclk));
	jdff dff_A_74wVKOLo1_0(.dout(w_dff_A_BFT77zb42_0),.din(w_dff_A_74wVKOLo1_0),.clk(gclk));
	jdff dff_A_99MEHm830_0(.dout(w_dff_A_74wVKOLo1_0),.din(w_dff_A_99MEHm830_0),.clk(gclk));
	jdff dff_A_FCiKgdIT2_0(.dout(w_dff_A_99MEHm830_0),.din(w_dff_A_FCiKgdIT2_0),.clk(gclk));
	jdff dff_A_vXuNS80w5_0(.dout(w_dff_A_FCiKgdIT2_0),.din(w_dff_A_vXuNS80w5_0),.clk(gclk));
	jdff dff_A_yf9aZ6Bo5_0(.dout(w_dff_A_vXuNS80w5_0),.din(w_dff_A_yf9aZ6Bo5_0),.clk(gclk));
	jdff dff_A_qJXJclC73_0(.dout(w_dff_A_yf9aZ6Bo5_0),.din(w_dff_A_qJXJclC73_0),.clk(gclk));
	jdff dff_A_66aYhiXR7_0(.dout(w_n184_0[0]),.din(w_dff_A_66aYhiXR7_0),.clk(gclk));
	jdff dff_A_CHas1LHi4_0(.dout(w_dff_A_66aYhiXR7_0),.din(w_dff_A_CHas1LHi4_0),.clk(gclk));
	jdff dff_A_fG3UcLW36_0(.dout(w_dff_A_CHas1LHi4_0),.din(w_dff_A_fG3UcLW36_0),.clk(gclk));
	jdff dff_A_mCVYHet33_2(.dout(w_n184_0[2]),.din(w_dff_A_mCVYHet33_2),.clk(gclk));
	jdff dff_A_aE84ATNk0_2(.dout(w_dff_A_mCVYHet33_2),.din(w_dff_A_aE84ATNk0_2),.clk(gclk));
	jdff dff_A_up7CYHIQ2_2(.dout(w_dff_A_aE84ATNk0_2),.din(w_dff_A_up7CYHIQ2_2),.clk(gclk));
	jdff dff_A_s6EPuhFG3_1(.dout(w_n159_0[1]),.din(w_dff_A_s6EPuhFG3_1),.clk(gclk));
	jdff dff_A_q1Tmkjhg8_0(.dout(w_Gid11_0[0]),.din(w_dff_A_q1Tmkjhg8_0),.clk(gclk));
	jdff dff_A_WoMNUxuA9_0(.dout(w_dff_A_q1Tmkjhg8_0),.din(w_dff_A_WoMNUxuA9_0),.clk(gclk));
	jdff dff_A_jTuDcu4A1_0(.dout(w_dff_A_WoMNUxuA9_0),.din(w_dff_A_jTuDcu4A1_0),.clk(gclk));
	jdff dff_A_sJKUTsoZ6_0(.dout(w_dff_A_jTuDcu4A1_0),.din(w_dff_A_sJKUTsoZ6_0),.clk(gclk));
	jdff dff_A_zTXQJi4O2_0(.dout(w_dff_A_sJKUTsoZ6_0),.din(w_dff_A_zTXQJi4O2_0),.clk(gclk));
	jdff dff_A_MDHdZqXY2_0(.dout(w_dff_A_zTXQJi4O2_0),.din(w_dff_A_MDHdZqXY2_0),.clk(gclk));
	jdff dff_A_zGVrZsi95_0(.dout(w_dff_A_MDHdZqXY2_0),.din(w_dff_A_zGVrZsi95_0),.clk(gclk));
	jdff dff_A_l6x9zAjl7_0(.dout(w_dff_A_zGVrZsi95_0),.din(w_dff_A_l6x9zAjl7_0),.clk(gclk));
	jdff dff_A_7tleaXJX8_0(.dout(w_dff_A_l6x9zAjl7_0),.din(w_dff_A_7tleaXJX8_0),.clk(gclk));
	jdff dff_A_ZLw59waI6_0(.dout(w_Gid3_0[0]),.din(w_dff_A_ZLw59waI6_0),.clk(gclk));
	jdff dff_A_pbkv4RCK0_0(.dout(w_dff_A_ZLw59waI6_0),.din(w_dff_A_pbkv4RCK0_0),.clk(gclk));
	jdff dff_A_h6BO7UyX8_0(.dout(w_dff_A_pbkv4RCK0_0),.din(w_dff_A_h6BO7UyX8_0),.clk(gclk));
	jdff dff_A_os3UQUEN7_0(.dout(w_dff_A_h6BO7UyX8_0),.din(w_dff_A_os3UQUEN7_0),.clk(gclk));
	jdff dff_A_BUgum97z5_0(.dout(w_dff_A_os3UQUEN7_0),.din(w_dff_A_BUgum97z5_0),.clk(gclk));
	jdff dff_A_8iHpVQn43_0(.dout(w_dff_A_BUgum97z5_0),.din(w_dff_A_8iHpVQn43_0),.clk(gclk));
	jdff dff_A_QVqaKatW4_0(.dout(w_dff_A_8iHpVQn43_0),.din(w_dff_A_QVqaKatW4_0),.clk(gclk));
	jdff dff_A_go8BBj3z6_0(.dout(w_dff_A_QVqaKatW4_0),.din(w_dff_A_go8BBj3z6_0),.clk(gclk));
	jdff dff_A_4I3nMOGK9_0(.dout(w_dff_A_go8BBj3z6_0),.din(w_dff_A_4I3nMOGK9_0),.clk(gclk));
	jdff dff_A_F9swWSKi8_0(.dout(w_dff_A_4I3nMOGK9_0),.din(w_dff_A_F9swWSKi8_0),.clk(gclk));
	jdff dff_B_aiquepbI0_2(.din(n250),.dout(w_dff_B_aiquepbI0_2),.clk(gclk));
	jdff dff_B_XdS5RqLz8_2(.din(w_dff_B_aiquepbI0_2),.dout(w_dff_B_XdS5RqLz8_2),.clk(gclk));
	jdff dff_A_duyvdjvf5_0(.dout(w_n178_0[0]),.din(w_dff_A_duyvdjvf5_0),.clk(gclk));
	jdff dff_A_VOoJv4I02_0(.dout(w_dff_A_duyvdjvf5_0),.din(w_dff_A_VOoJv4I02_0),.clk(gclk));
	jdff dff_A_JXsgy0qd6_0(.dout(w_dff_A_VOoJv4I02_0),.din(w_dff_A_JXsgy0qd6_0),.clk(gclk));
	jdff dff_A_ataSTmQa3_2(.dout(w_n178_0[2]),.din(w_dff_A_ataSTmQa3_2),.clk(gclk));
	jdff dff_A_h8aYYNzM2_2(.dout(w_dff_A_ataSTmQa3_2),.din(w_dff_A_h8aYYNzM2_2),.clk(gclk));
	jdff dff_A_m0QOCOpM9_2(.dout(w_dff_A_h8aYYNzM2_2),.din(w_dff_A_m0QOCOpM9_2),.clk(gclk));
	jdff dff_A_L009HIxL8_1(.dout(w_n150_0[1]),.din(w_dff_A_L009HIxL8_1),.clk(gclk));
	jdff dff_A_obwLJFET9_0(.dout(w_Gid9_0[0]),.din(w_dff_A_obwLJFET9_0),.clk(gclk));
	jdff dff_A_38vUVyGS0_0(.dout(w_dff_A_obwLJFET9_0),.din(w_dff_A_38vUVyGS0_0),.clk(gclk));
	jdff dff_A_tyNC6W9l4_0(.dout(w_dff_A_38vUVyGS0_0),.din(w_dff_A_tyNC6W9l4_0),.clk(gclk));
	jdff dff_A_pgv0ZQTQ7_0(.dout(w_dff_A_tyNC6W9l4_0),.din(w_dff_A_pgv0ZQTQ7_0),.clk(gclk));
	jdff dff_A_rZIop5ca6_0(.dout(w_dff_A_pgv0ZQTQ7_0),.din(w_dff_A_rZIop5ca6_0),.clk(gclk));
	jdff dff_A_LBLWlta38_0(.dout(w_dff_A_rZIop5ca6_0),.din(w_dff_A_LBLWlta38_0),.clk(gclk));
	jdff dff_A_hO6pMVH44_0(.dout(w_dff_A_LBLWlta38_0),.din(w_dff_A_hO6pMVH44_0),.clk(gclk));
	jdff dff_A_XSgzrLmB4_0(.dout(w_dff_A_hO6pMVH44_0),.din(w_dff_A_XSgzrLmB4_0),.clk(gclk));
	jdff dff_A_WcyjloGZ2_0(.dout(w_dff_A_XSgzrLmB4_0),.din(w_dff_A_WcyjloGZ2_0),.clk(gclk));
	jdff dff_A_cFjvw5JH8_0(.dout(w_Gid1_0[0]),.din(w_dff_A_cFjvw5JH8_0),.clk(gclk));
	jdff dff_A_7H716H7I0_0(.dout(w_dff_A_cFjvw5JH8_0),.din(w_dff_A_7H716H7I0_0),.clk(gclk));
	jdff dff_A_l67q1CMO8_0(.dout(w_dff_A_7H716H7I0_0),.din(w_dff_A_l67q1CMO8_0),.clk(gclk));
	jdff dff_A_E1bn7CGa6_0(.dout(w_dff_A_l67q1CMO8_0),.din(w_dff_A_E1bn7CGa6_0),.clk(gclk));
	jdff dff_A_t825I58D2_0(.dout(w_dff_A_E1bn7CGa6_0),.din(w_dff_A_t825I58D2_0),.clk(gclk));
	jdff dff_A_juBNwpGl8_0(.dout(w_dff_A_t825I58D2_0),.din(w_dff_A_juBNwpGl8_0),.clk(gclk));
	jdff dff_A_JIjB9Fy70_0(.dout(w_dff_A_juBNwpGl8_0),.din(w_dff_A_JIjB9Fy70_0),.clk(gclk));
	jdff dff_A_UadGAP8n7_0(.dout(w_dff_A_JIjB9Fy70_0),.din(w_dff_A_UadGAP8n7_0),.clk(gclk));
	jdff dff_A_CB67CI6b8_0(.dout(w_dff_A_UadGAP8n7_0),.din(w_dff_A_CB67CI6b8_0),.clk(gclk));
	jdff dff_A_zjbSdnLV9_0(.dout(w_dff_A_CB67CI6b8_0),.din(w_dff_A_zjbSdnLV9_0),.clk(gclk));
	jdff dff_A_0Rjp8F4g1_0(.dout(w_Gid26_0[0]),.din(w_dff_A_0Rjp8F4g1_0),.clk(gclk));
	jdff dff_A_kh98CfO54_0(.dout(w_dff_A_0Rjp8F4g1_0),.din(w_dff_A_kh98CfO54_0),.clk(gclk));
	jdff dff_A_GKKIGPxi3_0(.dout(w_dff_A_kh98CfO54_0),.din(w_dff_A_GKKIGPxi3_0),.clk(gclk));
	jdff dff_A_CTXqkuQH4_0(.dout(w_dff_A_GKKIGPxi3_0),.din(w_dff_A_CTXqkuQH4_0),.clk(gclk));
	jdff dff_A_ohLGYgoh5_0(.dout(w_dff_A_CTXqkuQH4_0),.din(w_dff_A_ohLGYgoh5_0),.clk(gclk));
	jdff dff_A_jV3smZcq9_0(.dout(w_dff_A_ohLGYgoh5_0),.din(w_dff_A_jV3smZcq9_0),.clk(gclk));
	jdff dff_A_imCf9JM81_0(.dout(w_dff_A_jV3smZcq9_0),.din(w_dff_A_imCf9JM81_0),.clk(gclk));
	jdff dff_A_vyKRC8Fd8_0(.dout(w_dff_A_imCf9JM81_0),.din(w_dff_A_vyKRC8Fd8_0),.clk(gclk));
	jdff dff_A_NEp2ucVn4_0(.dout(w_dff_A_vyKRC8Fd8_0),.din(w_dff_A_NEp2ucVn4_0),.clk(gclk));
	jdff dff_A_OvZnt1XA4_0(.dout(w_dff_A_NEp2ucVn4_0),.din(w_dff_A_OvZnt1XA4_0),.clk(gclk));
	jdff dff_A_i4agnnAC7_0(.dout(w_Gid25_0[0]),.din(w_dff_A_i4agnnAC7_0),.clk(gclk));
	jdff dff_A_TCzJcbbe7_0(.dout(w_dff_A_i4agnnAC7_0),.din(w_dff_A_TCzJcbbe7_0),.clk(gclk));
	jdff dff_A_EKLPA0jg1_0(.dout(w_dff_A_TCzJcbbe7_0),.din(w_dff_A_EKLPA0jg1_0),.clk(gclk));
	jdff dff_A_CFZSfiML6_0(.dout(w_dff_A_EKLPA0jg1_0),.din(w_dff_A_CFZSfiML6_0),.clk(gclk));
	jdff dff_A_GYa4Asfj9_0(.dout(w_dff_A_CFZSfiML6_0),.din(w_dff_A_GYa4Asfj9_0),.clk(gclk));
	jdff dff_A_NDFosJTS4_0(.dout(w_dff_A_GYa4Asfj9_0),.din(w_dff_A_NDFosJTS4_0),.clk(gclk));
	jdff dff_A_kFHIGF7R9_0(.dout(w_dff_A_NDFosJTS4_0),.din(w_dff_A_kFHIGF7R9_0),.clk(gclk));
	jdff dff_A_kFK45YSH2_0(.dout(w_dff_A_kFHIGF7R9_0),.din(w_dff_A_kFK45YSH2_0),.clk(gclk));
	jdff dff_A_icOdlJz91_0(.dout(w_dff_A_kFK45YSH2_0),.din(w_dff_A_icOdlJz91_0),.clk(gclk));
	jdff dff_A_1A0bEObr3_0(.dout(w_dff_A_icOdlJz91_0),.din(w_dff_A_1A0bEObr3_0),.clk(gclk));
	jdff dff_A_OZgTqKq69_0(.dout(w_Gid24_0[0]),.din(w_dff_A_OZgTqKq69_0),.clk(gclk));
	jdff dff_A_NwoNFBMR4_0(.dout(w_dff_A_OZgTqKq69_0),.din(w_dff_A_NwoNFBMR4_0),.clk(gclk));
	jdff dff_A_LMa73EUp2_0(.dout(w_dff_A_NwoNFBMR4_0),.din(w_dff_A_LMa73EUp2_0),.clk(gclk));
	jdff dff_A_gwDqsdTV1_0(.dout(w_dff_A_LMa73EUp2_0),.din(w_dff_A_gwDqsdTV1_0),.clk(gclk));
	jdff dff_A_8X8tpmhG6_0(.dout(w_dff_A_gwDqsdTV1_0),.din(w_dff_A_8X8tpmhG6_0),.clk(gclk));
	jdff dff_A_uVzoXuKk8_0(.dout(w_dff_A_8X8tpmhG6_0),.din(w_dff_A_uVzoXuKk8_0),.clk(gclk));
	jdff dff_A_A8v23lbd1_0(.dout(w_dff_A_uVzoXuKk8_0),.din(w_dff_A_A8v23lbd1_0),.clk(gclk));
	jdff dff_A_y2iRngSq2_0(.dout(w_dff_A_A8v23lbd1_0),.din(w_dff_A_y2iRngSq2_0),.clk(gclk));
	jdff dff_A_cU4WwANM7_0(.dout(w_dff_A_y2iRngSq2_0),.din(w_dff_A_cU4WwANM7_0),.clk(gclk));
	jdff dff_A_qlllOe9G5_0(.dout(w_dff_A_cU4WwANM7_0),.din(w_dff_A_qlllOe9G5_0),.clk(gclk));
	jdff dff_A_AaSaQZxW2_0(.dout(w_Gid30_0[0]),.din(w_dff_A_AaSaQZxW2_0),.clk(gclk));
	jdff dff_A_uPXwmlmu1_0(.dout(w_dff_A_AaSaQZxW2_0),.din(w_dff_A_uPXwmlmu1_0),.clk(gclk));
	jdff dff_A_WSkG8AvX5_0(.dout(w_dff_A_uPXwmlmu1_0),.din(w_dff_A_WSkG8AvX5_0),.clk(gclk));
	jdff dff_A_tuZS5JXj2_0(.dout(w_dff_A_WSkG8AvX5_0),.din(w_dff_A_tuZS5JXj2_0),.clk(gclk));
	jdff dff_A_S9zK4OwL6_0(.dout(w_dff_A_tuZS5JXj2_0),.din(w_dff_A_S9zK4OwL6_0),.clk(gclk));
	jdff dff_A_nUxSZ8Jt8_0(.dout(w_dff_A_S9zK4OwL6_0),.din(w_dff_A_nUxSZ8Jt8_0),.clk(gclk));
	jdff dff_A_nzoEoApV7_0(.dout(w_dff_A_nUxSZ8Jt8_0),.din(w_dff_A_nzoEoApV7_0),.clk(gclk));
	jdff dff_A_2HhnoT8C7_0(.dout(w_dff_A_nzoEoApV7_0),.din(w_dff_A_2HhnoT8C7_0),.clk(gclk));
	jdff dff_A_VEDrPZW67_0(.dout(w_dff_A_2HhnoT8C7_0),.din(w_dff_A_VEDrPZW67_0),.clk(gclk));
	jdff dff_A_ZCxqcaoc6_0(.dout(w_dff_A_VEDrPZW67_0),.din(w_dff_A_ZCxqcaoc6_0),.clk(gclk));
	jdff dff_A_LvZR9Phi7_0(.dout(w_Gid29_0[0]),.din(w_dff_A_LvZR9Phi7_0),.clk(gclk));
	jdff dff_A_PsBjJkkA1_0(.dout(w_dff_A_LvZR9Phi7_0),.din(w_dff_A_PsBjJkkA1_0),.clk(gclk));
	jdff dff_A_1mS88ppG6_0(.dout(w_dff_A_PsBjJkkA1_0),.din(w_dff_A_1mS88ppG6_0),.clk(gclk));
	jdff dff_A_aVmEZv8P6_0(.dout(w_dff_A_1mS88ppG6_0),.din(w_dff_A_aVmEZv8P6_0),.clk(gclk));
	jdff dff_A_MyJEfLPR1_0(.dout(w_dff_A_aVmEZv8P6_0),.din(w_dff_A_MyJEfLPR1_0),.clk(gclk));
	jdff dff_A_WYgMBVAS8_0(.dout(w_dff_A_MyJEfLPR1_0),.din(w_dff_A_WYgMBVAS8_0),.clk(gclk));
	jdff dff_A_YH47ltTr5_0(.dout(w_dff_A_WYgMBVAS8_0),.din(w_dff_A_YH47ltTr5_0),.clk(gclk));
	jdff dff_A_GD61wjyg1_0(.dout(w_dff_A_YH47ltTr5_0),.din(w_dff_A_GD61wjyg1_0),.clk(gclk));
	jdff dff_A_PZmG05BB1_0(.dout(w_dff_A_GD61wjyg1_0),.din(w_dff_A_PZmG05BB1_0),.clk(gclk));
	jdff dff_A_IIherzhR4_0(.dout(w_dff_A_PZmG05BB1_0),.din(w_dff_A_IIherzhR4_0),.clk(gclk));
	jdff dff_A_fovtXY267_0(.dout(w_Gid28_0[0]),.din(w_dff_A_fovtXY267_0),.clk(gclk));
	jdff dff_A_kbJT9drN5_0(.dout(w_dff_A_fovtXY267_0),.din(w_dff_A_kbJT9drN5_0),.clk(gclk));
	jdff dff_A_x5dBkqh31_0(.dout(w_dff_A_kbJT9drN5_0),.din(w_dff_A_x5dBkqh31_0),.clk(gclk));
	jdff dff_A_utaxoCqY8_0(.dout(w_dff_A_x5dBkqh31_0),.din(w_dff_A_utaxoCqY8_0),.clk(gclk));
	jdff dff_A_NklgPUGx9_0(.dout(w_dff_A_utaxoCqY8_0),.din(w_dff_A_NklgPUGx9_0),.clk(gclk));
	jdff dff_A_xUdDCLmE0_0(.dout(w_dff_A_NklgPUGx9_0),.din(w_dff_A_xUdDCLmE0_0),.clk(gclk));
	jdff dff_A_PXjVvBEB9_0(.dout(w_dff_A_xUdDCLmE0_0),.din(w_dff_A_PXjVvBEB9_0),.clk(gclk));
	jdff dff_A_DpSR2YLJ5_0(.dout(w_dff_A_PXjVvBEB9_0),.din(w_dff_A_DpSR2YLJ5_0),.clk(gclk));
	jdff dff_A_X9qv8aYt1_0(.dout(w_dff_A_DpSR2YLJ5_0),.din(w_dff_A_X9qv8aYt1_0),.clk(gclk));
	jdff dff_A_4mvnpGSs4_0(.dout(w_dff_A_X9qv8aYt1_0),.din(w_dff_A_4mvnpGSs4_0),.clk(gclk));
	jdff dff_A_M2PaOgjg4_1(.dout(w_n87_0[1]),.din(w_dff_A_M2PaOgjg4_1),.clk(gclk));
	jdff dff_A_gTU0I0Kb0_0(.dout(w_Gid22_0[0]),.din(w_dff_A_gTU0I0Kb0_0),.clk(gclk));
	jdff dff_A_WIs0Z4UN8_0(.dout(w_dff_A_gTU0I0Kb0_0),.din(w_dff_A_WIs0Z4UN8_0),.clk(gclk));
	jdff dff_A_u4wlr4fZ6_0(.dout(w_dff_A_WIs0Z4UN8_0),.din(w_dff_A_u4wlr4fZ6_0),.clk(gclk));
	jdff dff_A_GXgv57cO7_0(.dout(w_dff_A_u4wlr4fZ6_0),.din(w_dff_A_GXgv57cO7_0),.clk(gclk));
	jdff dff_A_wYwrtSa60_0(.dout(w_dff_A_GXgv57cO7_0),.din(w_dff_A_wYwrtSa60_0),.clk(gclk));
	jdff dff_A_bz7dgpLW0_0(.dout(w_dff_A_wYwrtSa60_0),.din(w_dff_A_bz7dgpLW0_0),.clk(gclk));
	jdff dff_A_Gimmhwj84_0(.dout(w_dff_A_bz7dgpLW0_0),.din(w_dff_A_Gimmhwj84_0),.clk(gclk));
	jdff dff_A_jdzJNB5P9_0(.dout(w_dff_A_Gimmhwj84_0),.din(w_dff_A_jdzJNB5P9_0),.clk(gclk));
	jdff dff_A_krzVkPLu8_0(.dout(w_dff_A_jdzJNB5P9_0),.din(w_dff_A_krzVkPLu8_0),.clk(gclk));
	jdff dff_A_ZVPfoTQT1_0(.dout(w_dff_A_krzVkPLu8_0),.din(w_dff_A_ZVPfoTQT1_0),.clk(gclk));
	jdff dff_A_T3PkQYSn8_0(.dout(w_Gid21_0[0]),.din(w_dff_A_T3PkQYSn8_0),.clk(gclk));
	jdff dff_A_18CUV6Ru3_0(.dout(w_dff_A_T3PkQYSn8_0),.din(w_dff_A_18CUV6Ru3_0),.clk(gclk));
	jdff dff_A_6pVS6k936_0(.dout(w_dff_A_18CUV6Ru3_0),.din(w_dff_A_6pVS6k936_0),.clk(gclk));
	jdff dff_A_lzsodhkK0_0(.dout(w_dff_A_6pVS6k936_0),.din(w_dff_A_lzsodhkK0_0),.clk(gclk));
	jdff dff_A_Twi8rjzG3_0(.dout(w_dff_A_lzsodhkK0_0),.din(w_dff_A_Twi8rjzG3_0),.clk(gclk));
	jdff dff_A_DXylPXA64_0(.dout(w_dff_A_Twi8rjzG3_0),.din(w_dff_A_DXylPXA64_0),.clk(gclk));
	jdff dff_A_mAXnUtDa9_0(.dout(w_dff_A_DXylPXA64_0),.din(w_dff_A_mAXnUtDa9_0),.clk(gclk));
	jdff dff_A_BdHwYyGn0_0(.dout(w_dff_A_mAXnUtDa9_0),.din(w_dff_A_BdHwYyGn0_0),.clk(gclk));
	jdff dff_A_punfCYko1_0(.dout(w_dff_A_BdHwYyGn0_0),.din(w_dff_A_punfCYko1_0),.clk(gclk));
	jdff dff_A_p6PpfRME7_0(.dout(w_dff_A_punfCYko1_0),.din(w_dff_A_p6PpfRME7_0),.clk(gclk));
	jdff dff_A_hAeLU9z48_0(.dout(w_Gid20_0[0]),.din(w_dff_A_hAeLU9z48_0),.clk(gclk));
	jdff dff_A_etOMWfyO9_0(.dout(w_dff_A_hAeLU9z48_0),.din(w_dff_A_etOMWfyO9_0),.clk(gclk));
	jdff dff_A_0XO7gUnA1_0(.dout(w_dff_A_etOMWfyO9_0),.din(w_dff_A_0XO7gUnA1_0),.clk(gclk));
	jdff dff_A_QZnDrBzG9_0(.dout(w_dff_A_0XO7gUnA1_0),.din(w_dff_A_QZnDrBzG9_0),.clk(gclk));
	jdff dff_A_7tTQfzcv2_0(.dout(w_dff_A_QZnDrBzG9_0),.din(w_dff_A_7tTQfzcv2_0),.clk(gclk));
	jdff dff_A_SFMbC9eO1_0(.dout(w_dff_A_7tTQfzcv2_0),.din(w_dff_A_SFMbC9eO1_0),.clk(gclk));
	jdff dff_A_vwehtSZr8_0(.dout(w_dff_A_SFMbC9eO1_0),.din(w_dff_A_vwehtSZr8_0),.clk(gclk));
	jdff dff_A_oXRTpgMH9_0(.dout(w_dff_A_vwehtSZr8_0),.din(w_dff_A_oXRTpgMH9_0),.clk(gclk));
	jdff dff_A_s8PsiCvj2_0(.dout(w_dff_A_oXRTpgMH9_0),.din(w_dff_A_s8PsiCvj2_0),.clk(gclk));
	jdff dff_A_dfvbAn5o2_0(.dout(w_dff_A_s8PsiCvj2_0),.din(w_dff_A_dfvbAn5o2_0),.clk(gclk));
	jdff dff_A_13ziitp32_0(.dout(w_Gid8_0[0]),.din(w_dff_A_13ziitp32_0),.clk(gclk));
	jdff dff_A_Os2y9z362_0(.dout(w_dff_A_13ziitp32_0),.din(w_dff_A_Os2y9z362_0),.clk(gclk));
	jdff dff_A_CDr5DGOV4_0(.dout(w_dff_A_Os2y9z362_0),.din(w_dff_A_CDr5DGOV4_0),.clk(gclk));
	jdff dff_A_P2zTSOq49_0(.dout(w_dff_A_CDr5DGOV4_0),.din(w_dff_A_P2zTSOq49_0),.clk(gclk));
	jdff dff_A_wOEwAWjA8_0(.dout(w_dff_A_P2zTSOq49_0),.din(w_dff_A_wOEwAWjA8_0),.clk(gclk));
	jdff dff_A_3Cq1DJl64_0(.dout(w_dff_A_wOEwAWjA8_0),.din(w_dff_A_3Cq1DJl64_0),.clk(gclk));
	jdff dff_A_ZKCrxvLZ9_0(.dout(w_dff_A_3Cq1DJl64_0),.din(w_dff_A_ZKCrxvLZ9_0),.clk(gclk));
	jdff dff_A_gOsP3EXH8_0(.dout(w_dff_A_ZKCrxvLZ9_0),.din(w_dff_A_gOsP3EXH8_0),.clk(gclk));
	jdff dff_A_h0Czj1or7_0(.dout(w_dff_A_gOsP3EXH8_0),.din(w_dff_A_h0Czj1or7_0),.clk(gclk));
	jdff dff_A_VTLfBYCw0_0(.dout(w_Gid0_0[0]),.din(w_dff_A_VTLfBYCw0_0),.clk(gclk));
	jdff dff_A_zgVfTEFh7_0(.dout(w_dff_A_VTLfBYCw0_0),.din(w_dff_A_zgVfTEFh7_0),.clk(gclk));
	jdff dff_A_RBWBVSMS7_0(.dout(w_dff_A_zgVfTEFh7_0),.din(w_dff_A_RBWBVSMS7_0),.clk(gclk));
	jdff dff_A_S6plSNAH6_0(.dout(w_dff_A_RBWBVSMS7_0),.din(w_dff_A_S6plSNAH6_0),.clk(gclk));
	jdff dff_A_xnV2Ju8e4_0(.dout(w_dff_A_S6plSNAH6_0),.din(w_dff_A_xnV2Ju8e4_0),.clk(gclk));
	jdff dff_A_xV84ZD570_0(.dout(w_dff_A_xnV2Ju8e4_0),.din(w_dff_A_xV84ZD570_0),.clk(gclk));
	jdff dff_A_4M3YrL6v0_0(.dout(w_dff_A_xV84ZD570_0),.din(w_dff_A_4M3YrL6v0_0),.clk(gclk));
	jdff dff_A_OspzlrJ09_0(.dout(w_dff_A_4M3YrL6v0_0),.din(w_dff_A_OspzlrJ09_0),.clk(gclk));
	jdff dff_A_TrPnLkSF3_0(.dout(w_dff_A_OspzlrJ09_0),.din(w_dff_A_TrPnLkSF3_0),.clk(gclk));
	jdff dff_A_PTACoQEj3_0(.dout(w_dff_A_TrPnLkSF3_0),.din(w_dff_A_PTACoQEj3_0),.clk(gclk));
	jdff dff_A_43cg13IY7_0(.dout(w_Gid18_0[0]),.din(w_dff_A_43cg13IY7_0),.clk(gclk));
	jdff dff_A_mxq1je1t2_0(.dout(w_dff_A_43cg13IY7_0),.din(w_dff_A_mxq1je1t2_0),.clk(gclk));
	jdff dff_A_mS1eXdau5_0(.dout(w_dff_A_mxq1je1t2_0),.din(w_dff_A_mS1eXdau5_0),.clk(gclk));
	jdff dff_A_nFVETzrZ4_0(.dout(w_dff_A_mS1eXdau5_0),.din(w_dff_A_nFVETzrZ4_0),.clk(gclk));
	jdff dff_A_g4RbweXX6_0(.dout(w_dff_A_nFVETzrZ4_0),.din(w_dff_A_g4RbweXX6_0),.clk(gclk));
	jdff dff_A_ig0ght1b3_0(.dout(w_dff_A_g4RbweXX6_0),.din(w_dff_A_ig0ght1b3_0),.clk(gclk));
	jdff dff_A_Ouy2aaX18_0(.dout(w_dff_A_ig0ght1b3_0),.din(w_dff_A_Ouy2aaX18_0),.clk(gclk));
	jdff dff_A_Ad33Ftai6_0(.dout(w_dff_A_Ouy2aaX18_0),.din(w_dff_A_Ad33Ftai6_0),.clk(gclk));
	jdff dff_A_90WTBUTz0_0(.dout(w_dff_A_Ad33Ftai6_0),.din(w_dff_A_90WTBUTz0_0),.clk(gclk));
	jdff dff_A_cp8oMZvJ2_0(.dout(w_dff_A_90WTBUTz0_0),.din(w_dff_A_cp8oMZvJ2_0),.clk(gclk));
	jdff dff_A_uELTC4HS0_0(.dout(w_Gid17_0[0]),.din(w_dff_A_uELTC4HS0_0),.clk(gclk));
	jdff dff_A_ZZzWmknK8_0(.dout(w_dff_A_uELTC4HS0_0),.din(w_dff_A_ZZzWmknK8_0),.clk(gclk));
	jdff dff_A_5nAuIPLh2_0(.dout(w_dff_A_ZZzWmknK8_0),.din(w_dff_A_5nAuIPLh2_0),.clk(gclk));
	jdff dff_A_K3RS4MwB4_0(.dout(w_dff_A_5nAuIPLh2_0),.din(w_dff_A_K3RS4MwB4_0),.clk(gclk));
	jdff dff_A_OreutxFh6_0(.dout(w_dff_A_K3RS4MwB4_0),.din(w_dff_A_OreutxFh6_0),.clk(gclk));
	jdff dff_A_onmFFsOP8_0(.dout(w_dff_A_OreutxFh6_0),.din(w_dff_A_onmFFsOP8_0),.clk(gclk));
	jdff dff_A_Qia66mh76_0(.dout(w_dff_A_onmFFsOP8_0),.din(w_dff_A_Qia66mh76_0),.clk(gclk));
	jdff dff_A_l2Fdh7NJ8_0(.dout(w_dff_A_Qia66mh76_0),.din(w_dff_A_l2Fdh7NJ8_0),.clk(gclk));
	jdff dff_A_FrWsUU4w4_0(.dout(w_dff_A_l2Fdh7NJ8_0),.din(w_dff_A_FrWsUU4w4_0),.clk(gclk));
	jdff dff_A_vZQsEkA11_0(.dout(w_dff_A_FrWsUU4w4_0),.din(w_dff_A_vZQsEkA11_0),.clk(gclk));
	jdff dff_A_5G4NSmpD5_0(.dout(w_Gid16_0[0]),.din(w_dff_A_5G4NSmpD5_0),.clk(gclk));
	jdff dff_A_GCEXWUqS2_0(.dout(w_dff_A_5G4NSmpD5_0),.din(w_dff_A_GCEXWUqS2_0),.clk(gclk));
	jdff dff_A_9nHm4XVh8_0(.dout(w_dff_A_GCEXWUqS2_0),.din(w_dff_A_9nHm4XVh8_0),.clk(gclk));
	jdff dff_A_ISqqhTi83_0(.dout(w_dff_A_9nHm4XVh8_0),.din(w_dff_A_ISqqhTi83_0),.clk(gclk));
	jdff dff_A_ncqyS2lK9_0(.dout(w_dff_A_ISqqhTi83_0),.din(w_dff_A_ncqyS2lK9_0),.clk(gclk));
	jdff dff_A_zbYCkq4b8_0(.dout(w_dff_A_ncqyS2lK9_0),.din(w_dff_A_zbYCkq4b8_0),.clk(gclk));
	jdff dff_A_CpdxpCqa6_0(.dout(w_dff_A_zbYCkq4b8_0),.din(w_dff_A_CpdxpCqa6_0),.clk(gclk));
	jdff dff_A_2UAWJVpw0_0(.dout(w_dff_A_CpdxpCqa6_0),.din(w_dff_A_2UAWJVpw0_0),.clk(gclk));
	jdff dff_A_dMhJLwUS9_0(.dout(w_dff_A_2UAWJVpw0_0),.din(w_dff_A_dMhJLwUS9_0),.clk(gclk));
	jdff dff_A_F4KuuzIG1_0(.dout(w_dff_A_dMhJLwUS9_0),.din(w_dff_A_F4KuuzIG1_0),.clk(gclk));
	jdff dff_A_WS4T4fbu6_1(.dout(w_n187_0[1]),.din(w_dff_A_WS4T4fbu6_1),.clk(gclk));
	jdff dff_A_SUWXhwpU6_1(.dout(w_dff_A_WS4T4fbu6_1),.din(w_dff_A_SUWXhwpU6_1),.clk(gclk));
	jdff dff_A_zFNKhXHj5_1(.dout(w_dff_A_SUWXhwpU6_1),.din(w_dff_A_zFNKhXHj5_1),.clk(gclk));
	jdff dff_A_Gp5oCYap9_1(.dout(w_dff_A_zFNKhXHj5_1),.din(w_dff_A_Gp5oCYap9_1),.clk(gclk));
	jdff dff_A_mezL70Ep5_2(.dout(w_n187_0[2]),.din(w_dff_A_mezL70Ep5_2),.clk(gclk));
	jdff dff_A_mvPXw4ex2_2(.dout(w_dff_A_mezL70Ep5_2),.din(w_dff_A_mvPXw4ex2_2),.clk(gclk));
	jdff dff_A_kSrOh2pl4_2(.dout(w_dff_A_mvPXw4ex2_2),.din(w_dff_A_kSrOh2pl4_2),.clk(gclk));
	jdff dff_A_KfhzSFjL0_2(.dout(w_dff_A_kSrOh2pl4_2),.din(w_dff_A_KfhzSFjL0_2),.clk(gclk));
	jdff dff_A_SrQ33Zs43_1(.dout(w_n102_1[1]),.din(w_dff_A_SrQ33Zs43_1),.clk(gclk));
	jdff dff_A_ayBzVqxe7_0(.dout(w_Gid31_0[0]),.din(w_dff_A_ayBzVqxe7_0),.clk(gclk));
	jdff dff_A_OsCJGy7G5_0(.dout(w_dff_A_ayBzVqxe7_0),.din(w_dff_A_OsCJGy7G5_0),.clk(gclk));
	jdff dff_A_hDykUPTt6_0(.dout(w_dff_A_OsCJGy7G5_0),.din(w_dff_A_hDykUPTt6_0),.clk(gclk));
	jdff dff_A_YOr88fZs6_0(.dout(w_dff_A_hDykUPTt6_0),.din(w_dff_A_YOr88fZs6_0),.clk(gclk));
	jdff dff_A_9Hicxlfj6_0(.dout(w_dff_A_YOr88fZs6_0),.din(w_dff_A_9Hicxlfj6_0),.clk(gclk));
	jdff dff_A_S5kaVC0d6_0(.dout(w_dff_A_9Hicxlfj6_0),.din(w_dff_A_S5kaVC0d6_0),.clk(gclk));
	jdff dff_A_r5f02Pg75_0(.dout(w_dff_A_S5kaVC0d6_0),.din(w_dff_A_r5f02Pg75_0),.clk(gclk));
	jdff dff_A_27OZu5vy8_0(.dout(w_dff_A_r5f02Pg75_0),.din(w_dff_A_27OZu5vy8_0),.clk(gclk));
	jdff dff_A_udL76qcW8_0(.dout(w_dff_A_27OZu5vy8_0),.din(w_dff_A_udL76qcW8_0),.clk(gclk));
	jdff dff_A_XsVLztRM6_0(.dout(w_dff_A_udL76qcW8_0),.din(w_dff_A_XsVLztRM6_0),.clk(gclk));
	jdff dff_A_pAWR0Zxn2_0(.dout(w_Gid27_0[0]),.din(w_dff_A_pAWR0Zxn2_0),.clk(gclk));
	jdff dff_A_G3o4Gvh99_0(.dout(w_dff_A_pAWR0Zxn2_0),.din(w_dff_A_G3o4Gvh99_0),.clk(gclk));
	jdff dff_A_tB46nrLl9_0(.dout(w_dff_A_G3o4Gvh99_0),.din(w_dff_A_tB46nrLl9_0),.clk(gclk));
	jdff dff_A_xsUikkql9_0(.dout(w_dff_A_tB46nrLl9_0),.din(w_dff_A_xsUikkql9_0),.clk(gclk));
	jdff dff_A_MgOuSpVs7_0(.dout(w_dff_A_xsUikkql9_0),.din(w_dff_A_MgOuSpVs7_0),.clk(gclk));
	jdff dff_A_LG73gyN70_0(.dout(w_dff_A_MgOuSpVs7_0),.din(w_dff_A_LG73gyN70_0),.clk(gclk));
	jdff dff_A_beARBm5V2_0(.dout(w_dff_A_LG73gyN70_0),.din(w_dff_A_beARBm5V2_0),.clk(gclk));
	jdff dff_A_fqWoQ2uE2_0(.dout(w_dff_A_beARBm5V2_0),.din(w_dff_A_fqWoQ2uE2_0),.clk(gclk));
	jdff dff_A_mHsqquK34_0(.dout(w_dff_A_fqWoQ2uE2_0),.din(w_dff_A_mHsqquK34_0),.clk(gclk));
	jdff dff_A_6EJUutyz5_0(.dout(w_dff_A_mHsqquK34_0),.din(w_dff_A_6EJUutyz5_0),.clk(gclk));
	jdff dff_A_dlCRRlbm7_0(.dout(w_Gid23_0[0]),.din(w_dff_A_dlCRRlbm7_0),.clk(gclk));
	jdff dff_A_3MpTAxUU5_0(.dout(w_dff_A_dlCRRlbm7_0),.din(w_dff_A_3MpTAxUU5_0),.clk(gclk));
	jdff dff_A_MevaaZEz8_0(.dout(w_dff_A_3MpTAxUU5_0),.din(w_dff_A_MevaaZEz8_0),.clk(gclk));
	jdff dff_A_Ae7ctVL45_0(.dout(w_dff_A_MevaaZEz8_0),.din(w_dff_A_Ae7ctVL45_0),.clk(gclk));
	jdff dff_A_WBqiegTa1_0(.dout(w_dff_A_Ae7ctVL45_0),.din(w_dff_A_WBqiegTa1_0),.clk(gclk));
	jdff dff_A_pqxqYhxx6_0(.dout(w_dff_A_WBqiegTa1_0),.din(w_dff_A_pqxqYhxx6_0),.clk(gclk));
	jdff dff_A_1TtFD5TO2_0(.dout(w_dff_A_pqxqYhxx6_0),.din(w_dff_A_1TtFD5TO2_0),.clk(gclk));
	jdff dff_A_wBNhqVY15_0(.dout(w_dff_A_1TtFD5TO2_0),.din(w_dff_A_wBNhqVY15_0),.clk(gclk));
	jdff dff_A_h3OHrec87_0(.dout(w_dff_A_wBNhqVY15_0),.din(w_dff_A_h3OHrec87_0),.clk(gclk));
	jdff dff_A_XdLnXq9U9_0(.dout(w_dff_A_h3OHrec87_0),.din(w_dff_A_XdLnXq9U9_0),.clk(gclk));
	jdff dff_A_aPbx6nzc7_0(.dout(w_Gid19_0[0]),.din(w_dff_A_aPbx6nzc7_0),.clk(gclk));
	jdff dff_A_RZklojRm9_0(.dout(w_dff_A_aPbx6nzc7_0),.din(w_dff_A_RZklojRm9_0),.clk(gclk));
	jdff dff_A_sFEORtIR9_0(.dout(w_dff_A_RZklojRm9_0),.din(w_dff_A_sFEORtIR9_0),.clk(gclk));
	jdff dff_A_uRBDuVzz8_0(.dout(w_dff_A_sFEORtIR9_0),.din(w_dff_A_uRBDuVzz8_0),.clk(gclk));
	jdff dff_A_fQ2piNSh3_0(.dout(w_dff_A_uRBDuVzz8_0),.din(w_dff_A_fQ2piNSh3_0),.clk(gclk));
	jdff dff_A_eC98ewXI3_0(.dout(w_dff_A_fQ2piNSh3_0),.din(w_dff_A_eC98ewXI3_0),.clk(gclk));
	jdff dff_A_tJ5moZB72_0(.dout(w_dff_A_eC98ewXI3_0),.din(w_dff_A_tJ5moZB72_0),.clk(gclk));
	jdff dff_A_iY7kSZQQ6_0(.dout(w_dff_A_tJ5moZB72_0),.din(w_dff_A_iY7kSZQQ6_0),.clk(gclk));
	jdff dff_A_31zVupeu1_0(.dout(w_dff_A_iY7kSZQQ6_0),.din(w_dff_A_31zVupeu1_0),.clk(gclk));
	jdff dff_A_njhaywae7_0(.dout(w_dff_A_31zVupeu1_0),.din(w_dff_A_njhaywae7_0),.clk(gclk));
	jdff dff_A_3vEXTt2O5_0(.dout(w_Gid15_0[0]),.din(w_dff_A_3vEXTt2O5_0),.clk(gclk));
	jdff dff_A_pvZffa4Y3_0(.dout(w_dff_A_3vEXTt2O5_0),.din(w_dff_A_pvZffa4Y3_0),.clk(gclk));
	jdff dff_A_wV9dlqrx8_0(.dout(w_dff_A_pvZffa4Y3_0),.din(w_dff_A_wV9dlqrx8_0),.clk(gclk));
	jdff dff_A_OsoCbngY1_0(.dout(w_dff_A_wV9dlqrx8_0),.din(w_dff_A_OsoCbngY1_0),.clk(gclk));
	jdff dff_A_J9Y53Guw0_0(.dout(w_dff_A_OsoCbngY1_0),.din(w_dff_A_J9Y53Guw0_0),.clk(gclk));
	jdff dff_A_qdaMsgC00_0(.dout(w_dff_A_J9Y53Guw0_0),.din(w_dff_A_qdaMsgC00_0),.clk(gclk));
	jdff dff_A_qYOVCnRs3_0(.dout(w_dff_A_qdaMsgC00_0),.din(w_dff_A_qYOVCnRs3_0),.clk(gclk));
	jdff dff_A_JDbXe0Kk6_0(.dout(w_dff_A_qYOVCnRs3_0),.din(w_dff_A_JDbXe0Kk6_0),.clk(gclk));
	jdff dff_A_fp8Lhak87_0(.dout(w_dff_A_JDbXe0Kk6_0),.din(w_dff_A_fp8Lhak87_0),.clk(gclk));
	jdff dff_A_DqsI2tef5_0(.dout(w_Gid14_0[0]),.din(w_dff_A_DqsI2tef5_0),.clk(gclk));
	jdff dff_A_5Id62eyV1_0(.dout(w_dff_A_DqsI2tef5_0),.din(w_dff_A_5Id62eyV1_0),.clk(gclk));
	jdff dff_A_RPzDK8EP9_0(.dout(w_dff_A_5Id62eyV1_0),.din(w_dff_A_RPzDK8EP9_0),.clk(gclk));
	jdff dff_A_DqR24QHW6_0(.dout(w_dff_A_RPzDK8EP9_0),.din(w_dff_A_DqR24QHW6_0),.clk(gclk));
	jdff dff_A_eofqEATT6_0(.dout(w_dff_A_DqR24QHW6_0),.din(w_dff_A_eofqEATT6_0),.clk(gclk));
	jdff dff_A_u9t5AbKR6_0(.dout(w_dff_A_eofqEATT6_0),.din(w_dff_A_u9t5AbKR6_0),.clk(gclk));
	jdff dff_A_VU4fVyCB1_0(.dout(w_dff_A_u9t5AbKR6_0),.din(w_dff_A_VU4fVyCB1_0),.clk(gclk));
	jdff dff_A_GhMeJAU66_0(.dout(w_dff_A_VU4fVyCB1_0),.din(w_dff_A_GhMeJAU66_0),.clk(gclk));
	jdff dff_A_7sIksdo32_0(.dout(w_dff_A_GhMeJAU66_0),.din(w_dff_A_7sIksdo32_0),.clk(gclk));
	jdff dff_A_A4MTaJyG7_0(.dout(w_Gid13_0[0]),.din(w_dff_A_A4MTaJyG7_0),.clk(gclk));
	jdff dff_A_T6jDC0ny1_0(.dout(w_dff_A_A4MTaJyG7_0),.din(w_dff_A_T6jDC0ny1_0),.clk(gclk));
	jdff dff_A_Y6aytHgg7_0(.dout(w_dff_A_T6jDC0ny1_0),.din(w_dff_A_Y6aytHgg7_0),.clk(gclk));
	jdff dff_A_tgBk6IEc0_0(.dout(w_dff_A_Y6aytHgg7_0),.din(w_dff_A_tgBk6IEc0_0),.clk(gclk));
	jdff dff_A_lMuE5vKe9_0(.dout(w_dff_A_tgBk6IEc0_0),.din(w_dff_A_lMuE5vKe9_0),.clk(gclk));
	jdff dff_A_FRBlaDhn3_0(.dout(w_dff_A_lMuE5vKe9_0),.din(w_dff_A_FRBlaDhn3_0),.clk(gclk));
	jdff dff_A_ifgivyBk4_0(.dout(w_dff_A_FRBlaDhn3_0),.din(w_dff_A_ifgivyBk4_0),.clk(gclk));
	jdff dff_A_uA7972LX0_0(.dout(w_dff_A_ifgivyBk4_0),.din(w_dff_A_uA7972LX0_0),.clk(gclk));
	jdff dff_A_u7SSCR2M0_0(.dout(w_dff_A_uA7972LX0_0),.din(w_dff_A_u7SSCR2M0_0),.clk(gclk));
	jdff dff_A_qtAlqtt74_0(.dout(w_Gid12_0[0]),.din(w_dff_A_qtAlqtt74_0),.clk(gclk));
	jdff dff_A_LWqr1tJp3_0(.dout(w_dff_A_qtAlqtt74_0),.din(w_dff_A_LWqr1tJp3_0),.clk(gclk));
	jdff dff_A_Ly6vFl2o1_0(.dout(w_dff_A_LWqr1tJp3_0),.din(w_dff_A_Ly6vFl2o1_0),.clk(gclk));
	jdff dff_A_CEkfR8YQ4_0(.dout(w_dff_A_Ly6vFl2o1_0),.din(w_dff_A_CEkfR8YQ4_0),.clk(gclk));
	jdff dff_A_o9mQOxpV7_0(.dout(w_dff_A_CEkfR8YQ4_0),.din(w_dff_A_o9mQOxpV7_0),.clk(gclk));
	jdff dff_A_Ny2axnXR6_0(.dout(w_dff_A_o9mQOxpV7_0),.din(w_dff_A_Ny2axnXR6_0),.clk(gclk));
	jdff dff_A_G30zSihx9_0(.dout(w_dff_A_Ny2axnXR6_0),.din(w_dff_A_G30zSihx9_0),.clk(gclk));
	jdff dff_A_4i5VYRsY1_0(.dout(w_dff_A_G30zSihx9_0),.din(w_dff_A_4i5VYRsY1_0),.clk(gclk));
	jdff dff_A_goQn8Qyb4_0(.dout(w_dff_A_4i5VYRsY1_0),.din(w_dff_A_goQn8Qyb4_0),.clk(gclk));
	jdff dff_A_iNp35z6R9_0(.dout(w_Gid7_0[0]),.din(w_dff_A_iNp35z6R9_0),.clk(gclk));
	jdff dff_A_maScKN3y1_0(.dout(w_dff_A_iNp35z6R9_0),.din(w_dff_A_maScKN3y1_0),.clk(gclk));
	jdff dff_A_OAFdzDG37_0(.dout(w_dff_A_maScKN3y1_0),.din(w_dff_A_OAFdzDG37_0),.clk(gclk));
	jdff dff_A_MjaR1rzo9_0(.dout(w_dff_A_OAFdzDG37_0),.din(w_dff_A_MjaR1rzo9_0),.clk(gclk));
	jdff dff_A_ACiX3UiA0_0(.dout(w_dff_A_MjaR1rzo9_0),.din(w_dff_A_ACiX3UiA0_0),.clk(gclk));
	jdff dff_A_VYfUQqX12_0(.dout(w_dff_A_ACiX3UiA0_0),.din(w_dff_A_VYfUQqX12_0),.clk(gclk));
	jdff dff_A_pUeDmXg80_0(.dout(w_dff_A_VYfUQqX12_0),.din(w_dff_A_pUeDmXg80_0),.clk(gclk));
	jdff dff_A_gKkyzRf58_0(.dout(w_dff_A_pUeDmXg80_0),.din(w_dff_A_gKkyzRf58_0),.clk(gclk));
	jdff dff_A_mlCME7o44_0(.dout(w_dff_A_gKkyzRf58_0),.din(w_dff_A_mlCME7o44_0),.clk(gclk));
	jdff dff_A_RLZnhZwo1_0(.dout(w_dff_A_mlCME7o44_0),.din(w_dff_A_RLZnhZwo1_0),.clk(gclk));
	jdff dff_A_ZfYRbZaL8_0(.dout(w_Gid6_0[0]),.din(w_dff_A_ZfYRbZaL8_0),.clk(gclk));
	jdff dff_A_H7x4cxRG7_0(.dout(w_dff_A_ZfYRbZaL8_0),.din(w_dff_A_H7x4cxRG7_0),.clk(gclk));
	jdff dff_A_iqB6IdW90_0(.dout(w_dff_A_H7x4cxRG7_0),.din(w_dff_A_iqB6IdW90_0),.clk(gclk));
	jdff dff_A_FyydgOjX7_0(.dout(w_dff_A_iqB6IdW90_0),.din(w_dff_A_FyydgOjX7_0),.clk(gclk));
	jdff dff_A_k8h9TTbj5_0(.dout(w_dff_A_FyydgOjX7_0),.din(w_dff_A_k8h9TTbj5_0),.clk(gclk));
	jdff dff_A_dVSuBviO3_0(.dout(w_dff_A_k8h9TTbj5_0),.din(w_dff_A_dVSuBviO3_0),.clk(gclk));
	jdff dff_A_YH8VLY5L1_0(.dout(w_dff_A_dVSuBviO3_0),.din(w_dff_A_YH8VLY5L1_0),.clk(gclk));
	jdff dff_A_fbqP6Ep64_0(.dout(w_dff_A_YH8VLY5L1_0),.din(w_dff_A_fbqP6Ep64_0),.clk(gclk));
	jdff dff_A_GaRLcLru9_0(.dout(w_dff_A_fbqP6Ep64_0),.din(w_dff_A_GaRLcLru9_0),.clk(gclk));
	jdff dff_A_fEzr8Q1O8_0(.dout(w_dff_A_GaRLcLru9_0),.din(w_dff_A_fEzr8Q1O8_0),.clk(gclk));
	jdff dff_A_GOwmHF5K7_0(.dout(w_Gid5_0[0]),.din(w_dff_A_GOwmHF5K7_0),.clk(gclk));
	jdff dff_A_oG4BV4si9_0(.dout(w_dff_A_GOwmHF5K7_0),.din(w_dff_A_oG4BV4si9_0),.clk(gclk));
	jdff dff_A_Qonvgfhz0_0(.dout(w_dff_A_oG4BV4si9_0),.din(w_dff_A_Qonvgfhz0_0),.clk(gclk));
	jdff dff_A_iNlfX4sN5_0(.dout(w_dff_A_Qonvgfhz0_0),.din(w_dff_A_iNlfX4sN5_0),.clk(gclk));
	jdff dff_A_19OnYZKV4_0(.dout(w_dff_A_iNlfX4sN5_0),.din(w_dff_A_19OnYZKV4_0),.clk(gclk));
	jdff dff_A_N5d65ejs1_0(.dout(w_dff_A_19OnYZKV4_0),.din(w_dff_A_N5d65ejs1_0),.clk(gclk));
	jdff dff_A_vbE2pn4c1_0(.dout(w_dff_A_N5d65ejs1_0),.din(w_dff_A_vbE2pn4c1_0),.clk(gclk));
	jdff dff_A_rjQt1ruS5_0(.dout(w_dff_A_vbE2pn4c1_0),.din(w_dff_A_rjQt1ruS5_0),.clk(gclk));
	jdff dff_A_FXMUWy943_0(.dout(w_dff_A_rjQt1ruS5_0),.din(w_dff_A_FXMUWy943_0),.clk(gclk));
	jdff dff_A_LhFtLdlN9_0(.dout(w_dff_A_FXMUWy943_0),.din(w_dff_A_LhFtLdlN9_0),.clk(gclk));
	jdff dff_A_YxFBohNB7_0(.dout(w_Gid4_0[0]),.din(w_dff_A_YxFBohNB7_0),.clk(gclk));
	jdff dff_A_J0Mz2ybJ0_0(.dout(w_dff_A_YxFBohNB7_0),.din(w_dff_A_J0Mz2ybJ0_0),.clk(gclk));
	jdff dff_A_l7uWztIC1_0(.dout(w_dff_A_J0Mz2ybJ0_0),.din(w_dff_A_l7uWztIC1_0),.clk(gclk));
	jdff dff_A_swupLrXb5_0(.dout(w_dff_A_l7uWztIC1_0),.din(w_dff_A_swupLrXb5_0),.clk(gclk));
	jdff dff_A_SYOKoGYC8_0(.dout(w_dff_A_swupLrXb5_0),.din(w_dff_A_SYOKoGYC8_0),.clk(gclk));
	jdff dff_A_imZhQM7P7_0(.dout(w_dff_A_SYOKoGYC8_0),.din(w_dff_A_imZhQM7P7_0),.clk(gclk));
	jdff dff_A_KzaP0acl2_0(.dout(w_dff_A_imZhQM7P7_0),.din(w_dff_A_KzaP0acl2_0),.clk(gclk));
	jdff dff_A_rlQwKjD73_0(.dout(w_dff_A_KzaP0acl2_0),.din(w_dff_A_rlQwKjD73_0),.clk(gclk));
	jdff dff_A_bSYgqp1s3_0(.dout(w_dff_A_rlQwKjD73_0),.din(w_dff_A_bSYgqp1s3_0),.clk(gclk));
	jdff dff_A_eYIyeTjg8_0(.dout(w_dff_A_bSYgqp1s3_0),.din(w_dff_A_eYIyeTjg8_0),.clk(gclk));
	jdff dff_A_SymbD6mv0_2(.dout(God8),.din(w_dff_A_SymbD6mv0_2),.clk(gclk));
	jdff dff_A_3D6ctpqb9_2(.dout(God9),.din(w_dff_A_3D6ctpqb9_2),.clk(gclk));
	jdff dff_A_GMwuJEWF7_2(.dout(God10),.din(w_dff_A_GMwuJEWF7_2),.clk(gclk));
	jdff dff_A_nxTxlJCZ9_2(.dout(God11),.din(w_dff_A_nxTxlJCZ9_2),.clk(gclk));
	jdff dff_A_GU7KRKHU2_2(.dout(God12),.din(w_dff_A_GU7KRKHU2_2),.clk(gclk));
	jdff dff_A_GLtL4owQ8_2(.dout(God13),.din(w_dff_A_GLtL4owQ8_2),.clk(gclk));
	jdff dff_A_p1uJu0Ob8_2(.dout(God14),.din(w_dff_A_p1uJu0Ob8_2),.clk(gclk));
	jdff dff_A_VEiGf8yR7_2(.dout(God15),.din(w_dff_A_VEiGf8yR7_2),.clk(gclk));
endmodule

