/*
rf_c432:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jdff: 1153
	jand: 111
	jor: 110

Summary:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jdff: 1153
	jand: 111
	jor: 110

The maximum logic level gap of any gate:
	rf_c432: 8
*/

module rf_c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n43;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n150;
	wire n151;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n217;
	wire n218;
	wire n219;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n235;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n244;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n262;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G4gat_0;
	wire [2:0] w_G8gat_0;
	wire [2:0] w_G11gat_0;
	wire [2:0] w_G14gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G21gat_0;
	wire [1:0] w_G21gat_1;
	wire [1:0] w_G24gat_0;
	wire [1:0] w_G27gat_0;
	wire [1:0] w_G30gat_0;
	wire [2:0] w_G34gat_0;
	wire [2:0] w_G37gat_0;
	wire [1:0] w_G40gat_0;
	wire [2:0] w_G43gat_0;
	wire [1:0] w_G43gat_1;
	wire [1:0] w_G47gat_0;
	wire [2:0] w_G50gat_0;
	wire [1:0] w_G53gat_0;
	wire [2:0] w_G56gat_0;
	wire [2:0] w_G60gat_0;
	wire [2:0] w_G63gat_0;
	wire [1:0] w_G66gat_0;
	wire [2:0] w_G69gat_0;
	wire [2:0] w_G73gat_0;
	wire [1:0] w_G76gat_0;
	wire [1:0] w_G79gat_0;
	wire [2:0] w_G82gat_0;
	wire [2:0] w_G86gat_0;
	wire [1:0] w_G86gat_1;
	wire [2:0] w_G89gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G95gat_0;
	wire [2:0] w_G99gat_0;
	wire [2:0] w_G102gat_0;
	wire [1:0] w_G105gat_0;
	wire [2:0] w_G108gat_0;
	wire [2:0] w_G112gat_0;
	wire [1:0] w_G115gat_0;
	wire [2:0] w_G223gat_0;
	wire [2:0] w_G223gat_1;
	wire [2:0] w_G223gat_2;
	wire [1:0] w_G223gat_3;
	wire G223gat_fa_;
	wire [2:0] w_G329gat_0;
	wire [2:0] w_G329gat_1;
	wire [2:0] w_G329gat_2;
	wire [2:0] w_G329gat_3;
	wire [2:0] w_G329gat_4;
	wire [2:0] w_G329gat_5;
	wire w_G329gat_6;
	wire G329gat_fa_;
	wire [2:0] w_G370gat_0;
	wire [2:0] w_G370gat_1;
	wire w_G370gat_2;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire [1:0] w_n43_0;
	wire [1:0] w_n44_0;
	wire [1:0] w_n47_0;
	wire [1:0] w_n52_0;
	wire [1:0] w_n53_0;
	wire [1:0] w_n56_0;
	wire [1:0] w_n58_0;
	wire [1:0] w_n61_0;
	wire [1:0] w_n63_0;
	wire [1:0] w_n69_0;
	wire [1:0] w_n71_0;
	wire [1:0] w_n72_0;
	wire [1:0] w_n73_0;
	wire [1:0] w_n77_0;
	wire [1:0] w_n78_0;
	wire [1:0] w_n79_0;
	wire [1:0] w_n82_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n87_0;
	wire [1:0] w_n89_0;
	wire [2:0] w_n94_0;
	wire [2:0] w_n94_1;
	wire [2:0] w_n94_2;
	wire [2:0] w_n94_3;
	wire [1:0] w_n94_4;
	wire [1:0] w_n96_0;
	wire [1:0] w_n98_0;
	wire [1:0] w_n100_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n109_0;
	wire [2:0] w_n114_0;
	wire [1:0] w_n115_0;
	wire [1:0] w_n119_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n123_0;
	wire [2:0] w_n126_0;
	wire [1:0] w_n128_0;
	wire [2:0] w_n130_0;
	wire [1:0] w_n132_0;
	wire [1:0] w_n139_0;
	wire [1:0] w_n141_0;
	wire [1:0] w_n142_0;
	wire [1:0] w_n145_0;
	wire [1:0] w_n146_0;
	wire [1:0] w_n147_0;
	wire [1:0] w_n150_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n154_0;
	wire [1:0] w_n156_0;
	wire [1:0] w_n159_0;
	wire [1:0] w_n164_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n174_0;
	wire [1:0] w_n177_0;
	wire [2:0] w_n182_0;
	wire [2:0] w_n182_1;
	wire [2:0] w_n182_2;
	wire [1:0] w_n182_3;
	wire [1:0] w_n184_0;
	wire [1:0] w_n188_0;
	wire [1:0] w_n191_0;
	wire [1:0] w_n193_0;
	wire [1:0] w_n197_0;
	wire [1:0] w_n198_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n217_0;
	wire [1:0] w_n219_0;
	wire [1:0] w_n222_0;
	wire [1:0] w_n224_0;
	wire [1:0] w_n231_0;
	wire [1:0] w_n254_0;
	wire [1:0] w_n260_0;
	wire [2:0] w_n271_0;
	wire [2:0] w_n271_1;
	wire [2:0] w_n271_2;
	wire [1:0] w_n271_3;
	wire [1:0] w_n274_0;
	wire [1:0] w_n281_0;
	wire [1:0] w_n283_0;
	wire [1:0] w_n286_0;
	wire [1:0] w_n290_0;
	wire [1:0] w_n293_0;
	wire [1:0] w_n296_0;
	wire [1:0] w_n303_0;
	wire [1:0] w_n305_0;
	wire [1:0] w_n313_0;
	wire [1:0] w_n314_0;
	wire [2:0] w_n317_0;
	wire [1:0] w_n319_0;
	wire w_dff_B_95uf8pzk0_1;
	wire w_dff_B_letGXm1p6_1;
	wire w_dff_B_TBCYFE2o0_1;
	wire w_dff_B_pTm7TwKv4_0;
	wire w_dff_B_ZFViDVo62_0;
	wire w_dff_B_M4uKZ33d6_0;
	wire w_dff_B_BzQbd4wn1_0;
	wire w_dff_B_2aQgTpKd8_0;
	wire w_dff_B_zqiK0Xpw6_1;
	wire w_dff_A_ap4p4pgH8_0;
	wire w_dff_B_Zb5l6RDP0_0;
	wire w_dff_B_XihP7rBk7_0;
	wire w_dff_B_tm2ksOGf1_0;
	wire w_dff_B_mKHebEnU9_0;
	wire w_dff_B_TNL17A3L5_0;
	wire w_dff_A_bhTq7Q2L7_0;
	wire w_dff_B_RIYvRidS5_1;
	wire w_dff_B_LSjvtylg8_0;
	wire w_dff_B_MqE7YZoz4_0;
	wire w_dff_B_ZTCuf4J51_0;
	wire w_dff_B_KlpllYaD6_0;
	wire w_dff_B_DkoggYqW3_0;
	wire w_dff_A_lUbJeBKw1_0;
	wire w_dff_A_Ht0QTSse1_0;
	wire w_dff_A_qS4YkDag0_0;
	wire w_dff_A_DxhtPWx42_0;
	wire w_dff_A_Y6V6tujw5_0;
	wire w_dff_A_YbFHvBUL5_0;
	wire w_dff_A_ww5EVM0P1_0;
	wire w_dff_B_61851nHU8_1;
	wire w_dff_B_Vy3M2GSb4_1;
	wire w_dff_B_lsmVxR8I6_1;
	wire w_dff_B_OGRnpnlf3_1;
	wire w_dff_B_IOwF4Glq7_1;
	wire w_dff_B_63lnhOn55_1;
	wire w_dff_B_sMrOjCU75_1;
	wire w_dff_B_sFDJB6s57_1;
	wire w_dff_B_ZAn4Sgqp9_1;
	wire w_dff_B_P06ILHvw6_1;
	wire w_dff_B_zZX3Faph4_1;
	wire w_dff_B_XaagROtF9_1;
	wire w_dff_B_QEnaAqci1_1;
	wire w_dff_B_EYcpcktT1_1;
	wire w_dff_B_s5oZxAZy6_1;
	wire w_dff_B_Y3tVv5mi2_1;
	wire w_dff_B_4EwAZuwG0_1;
	wire w_dff_B_bPVohXzw7_1;
	wire w_dff_B_XMUnQGRf5_1;
	wire w_dff_B_XvNhl9Hs3_1;
	wire w_dff_B_87glUefm9_1;
	wire w_dff_B_l5MATZEJ2_1;
	wire w_dff_B_vCzdesii0_1;
	wire w_dff_B_jfxZeJNT7_1;
	wire w_dff_B_erZJyVKo4_1;
	wire w_dff_B_RwErxWos9_1;
	wire w_dff_B_eADzKhT00_1;
	wire w_dff_B_zDm1Bszp8_0;
	wire w_dff_B_yx1vB4yl4_0;
	wire w_dff_B_Gh5mMvPZ6_0;
	wire w_dff_A_YvsfF6k72_1;
	wire w_dff_A_yqcP8mIO8_1;
	wire w_dff_A_p4YkqInR2_1;
	wire w_dff_A_wfABZNCu4_1;
	wire w_dff_A_nu4IWkEs7_1;
	wire w_dff_A_ZkBAqm027_1;
	wire w_dff_B_Vhe6vJ0b1_1;
	wire w_dff_B_tXGSSCjs9_0;
	wire w_dff_B_V4QtIwkQ2_0;
	wire w_dff_B_rnzU1YTc2_0;
	wire w_dff_B_wszG0AMj8_0;
	wire w_dff_B_sJNE8zIO8_0;
	wire w_dff_B_a1rqcxTg0_1;
	wire w_dff_B_qUUUr8lb5_0;
	wire w_dff_B_maInDkaC0_0;
	wire w_dff_B_39ayU2Sl8_0;
	wire w_dff_B_iR4wkDcl9_0;
	wire w_dff_A_3WSsRxUf9_0;
	wire w_dff_A_se6up4Ss9_0;
	wire w_dff_A_cHk6rDJq0_0;
	wire w_dff_A_jCNboXfa1_0;
	wire w_dff_A_IMLsThk60_0;
	wire w_dff_A_GzvYsrTd6_0;
	wire w_dff_A_SKKqbJ652_0;
	wire w_dff_A_8zBGWutK1_0;
	wire w_dff_A_jT2p71gI7_0;
	wire w_dff_A_SXoqwkCD7_0;
	wire w_dff_A_k33Srw5y6_0;
	wire w_dff_A_kM1VUIek2_0;
	wire w_dff_A_eb3iF4Np2_0;
	wire w_dff_A_nC1hyU7V1_0;
	wire w_dff_A_Ux3zMEJf2_0;
	wire w_dff_A_BJy6mq5s7_0;
	wire w_dff_A_q8Bkd44h3_0;
	wire w_dff_A_tVDtwLTa1_0;
	wire w_dff_B_akSLQiSm2_0;
	wire w_dff_B_LBaWGVAn0_0;
	wire w_dff_B_5AGmBoIP4_0;
	wire w_dff_B_kauUpNH26_0;
	wire w_dff_B_Cje7cwRF8_0;
	wire w_dff_B_uXF6yqlK1_0;
	wire w_dff_B_moVH5SBR5_1;
	wire w_dff_B_0pCmD9204_1;
	wire w_dff_B_WWvHWYd57_1;
	wire w_dff_A_ux7bgzkJ7_0;
	wire w_dff_A_IPNqJfBU6_0;
	wire w_dff_A_KxMR96IR3_0;
	wire w_dff_A_cNOtW5Mx9_0;
	wire w_dff_A_qOv4CHeU1_0;
	wire w_dff_A_6c6mhX8v0_0;
	wire w_dff_A_fDii76br6_0;
	wire w_dff_A_zpHB0f9z4_0;
	wire w_dff_A_llTFJ1Qm0_0;
	wire w_dff_A_ybiPwF451_0;
	wire w_dff_A_UrpyTP039_0;
	wire w_dff_B_T3Is5w2W2_2;
	wire w_dff_B_pKTwd5Z91_2;
	wire w_dff_B_CqtvmWDt2_2;
	wire w_dff_B_08764Txh0_2;
	wire w_dff_B_pXtP3Vtx6_2;
	wire w_dff_B_eKkeObvC3_2;
	wire w_dff_B_OJgdGmN87_2;
	wire w_dff_B_pSVPQ7HT1_2;
	wire w_dff_B_t92uup1W4_2;
	wire w_dff_B_vlqbdS308_2;
	wire w_dff_B_jnVQKEtB0_2;
	wire w_dff_B_6aDjtOHo2_2;
	wire w_dff_B_12btdkct8_2;
	wire w_dff_B_gbWZni8G5_2;
	wire w_dff_A_Grp4gKbN7_0;
	wire w_dff_A_ITG7dhPe3_0;
	wire w_dff_A_rOAgBkxG5_0;
	wire w_dff_A_e8bdT4yK3_0;
	wire w_dff_A_SDe99cyn0_0;
	wire w_dff_A_e8PApaLy4_0;
	wire w_dff_A_KHl453nB9_0;
	wire w_dff_A_Jz1BAu5o4_0;
	wire w_dff_A_W99BY7sm6_0;
	wire w_dff_A_8UNSU2Zm8_0;
	wire w_dff_A_vo7ecOzY8_0;
	wire w_dff_A_cNYE0Rxi5_0;
	wire w_dff_A_oM79tBM66_0;
	wire w_dff_A_JO4lQiNv4_0;
	wire w_dff_A_AvwkGZtH5_0;
	wire w_dff_A_9KkDxQ5a3_1;
	wire w_dff_A_d8smjoO24_1;
	wire w_dff_A_iYCqwx7Q1_1;
	wire w_dff_A_LmDCxI092_1;
	wire w_dff_A_RzoDSxuh6_0;
	wire w_dff_A_87mnJcZt7_0;
	wire w_dff_A_Cn4HUcMZ8_0;
	wire w_dff_A_4WHONs2a7_0;
	wire w_dff_A_tf2Eq1HF3_0;
	wire w_dff_A_5dQwUhWN5_0;
	wire w_dff_A_XVPZIjSM2_0;
	wire w_dff_A_bKBSNtxC2_0;
	wire w_dff_A_hQecb5Yc4_0;
	wire w_dff_A_GYxAzLjh8_0;
	wire w_dff_A_zSHVQ4E95_0;
	wire w_dff_B_nMRYpbD35_2;
	wire w_dff_B_vCdUxLIY4_2;
	wire w_dff_B_ZIWcIQdJ4_2;
	wire w_dff_B_JyJZ34XK2_2;
	wire w_dff_B_zRU6HOQA3_2;
	wire w_dff_B_qAJHj5iF4_2;
	wire w_dff_B_Z2zh11bp5_2;
	wire w_dff_B_fgU23e0C8_2;
	wire w_dff_A_8xMlCICc9_0;
	wire w_dff_A_n85eMn4U7_0;
	wire w_dff_A_hP8Jo5fs6_0;
	wire w_dff_A_3GJcADem5_0;
	wire w_dff_A_ayoFeQod0_0;
	wire w_dff_A_qpPAXIMO3_0;
	wire w_dff_A_wXmZkkXC5_0;
	wire w_dff_A_Ztxnv9k10_0;
	wire w_dff_A_hzillUTC0_0;
	wire w_dff_A_OybFytYO1_0;
	wire w_dff_A_kwAPfovI5_0;
	wire w_dff_A_T4MwwXy39_0;
	wire w_dff_A_0iTrAXob9_0;
	wire w_dff_A_piB35lYS0_0;
	wire w_dff_A_kYFkFj4w9_0;
	wire w_dff_A_pXpSgiNB9_0;
	wire w_dff_A_y6Ii1q5d4_0;
	wire w_dff_A_KA6riDI94_0;
	wire w_dff_A_flqTqVj67_0;
	wire w_dff_A_diYIX76x0_0;
	wire w_dff_B_lnn5Uzfq6_1;
	wire w_dff_B_U98fcXty5_1;
	wire w_dff_B_xlcXHhRu7_1;
	wire w_dff_B_efK2R0bh5_1;
	wire w_dff_B_X67VoH9R1_1;
	wire w_dff_B_TGwtTXDD7_1;
	wire w_dff_B_00zlxIno6_1;
	wire w_dff_B_6KJG3Flh1_1;
	wire w_dff_B_fALiyNYM4_1;
	wire w_dff_B_z1LzTmC00_1;
	wire w_dff_B_B01hDh9Y3_1;
	wire w_dff_B_o98iBe3S6_1;
	wire w_dff_B_xElPkw5s0_1;
	wire w_dff_B_W5Y98niU1_1;
	wire w_dff_B_1hD0ELZz5_1;
	wire w_dff_B_L28FJEj32_1;
	wire w_dff_B_bUzvdw0K2_1;
	wire w_dff_B_AXbgqMsT7_1;
	wire w_dff_B_EGEo9Tis2_1;
	wire w_dff_B_krtebK9K0_1;
	wire w_dff_B_qitdhjvU1_1;
	wire w_dff_B_YrtmM10h8_1;
	wire w_dff_B_HmraLxQV5_1;
	wire w_dff_B_A6mZnrIx9_1;
	wire w_dff_B_IRfLmUY64_1;
	wire w_dff_B_dpOwkNU81_1;
	wire w_dff_A_TpSj3xwa4_0;
	wire w_dff_A_cnwC30Rj0_0;
	wire w_dff_A_YUca2dnA6_0;
	wire w_dff_A_nyA0KeG70_0;
	wire w_dff_A_87Dcb33u9_0;
	wire w_dff_A_QRl0R2Rj7_0;
	wire w_dff_A_hNQMmCzg6_0;
	wire w_dff_A_LLwNLMZU3_0;
	wire w_dff_A_zSyOxV917_0;
	wire w_dff_A_I6lDnbCy9_0;
	wire w_dff_A_aSyy6zo64_0;
	wire w_dff_A_aNyeiOYG6_0;
	wire w_dff_A_Srj0DVv62_0;
	wire w_dff_A_7g9FVgZL0_0;
	wire w_dff_A_X0N0VDcb5_0;
	wire w_dff_A_ZqZMyaQl6_1;
	wire w_dff_A_aTIWMwVj2_1;
	wire w_dff_A_le4NPD2O9_1;
	wire w_dff_A_ybQYTo8r8_1;
	wire w_dff_A_pLdptZsi5_1;
	wire w_dff_A_QL7Q4aix8_1;
	wire w_dff_A_vkziZMf91_1;
	wire w_dff_A_8zERPKfg0_1;
	wire w_dff_A_WxUBDYyB5_1;
	wire w_dff_A_GCO729jO1_1;
	wire w_dff_A_Sg2vU5sp9_1;
	wire w_dff_A_n2X8c3xd3_1;
	wire w_dff_A_bQX8fFmd2_1;
	wire w_dff_A_FukfDVB72_1;
	wire w_dff_A_IVEt6Yi41_1;
	wire w_dff_A_rnL2bv6w1_1;
	wire w_dff_A_9zWOeDKj4_1;
	wire w_dff_A_PX4wzWm83_1;
	wire w_dff_A_F43mayrn8_1;
	wire w_dff_A_reYrKxhI4_1;
	wire w_dff_A_5O11Kk6m7_0;
	wire w_dff_A_jHfTwugk2_0;
	wire w_dff_A_Z39AWxCp2_0;
	wire w_dff_A_QncNGc8c7_0;
	wire w_dff_A_OnOWwz199_0;
	wire w_dff_A_mutchN9n9_0;
	wire w_dff_B_5na9E6hu8_2;
	wire w_dff_B_lldkz9KD6_2;
	wire w_dff_B_eXp3ymoj3_2;
	wire w_dff_B_w50sHWmX1_2;
	wire w_dff_B_momk3OCZ7_2;
	wire w_dff_B_VPnhVvQf6_2;
	wire w_dff_B_i7T2ylon8_2;
	wire w_dff_B_Hg1wGNpr9_2;
	wire w_dff_B_XQEDxvVJ3_2;
	wire w_dff_B_8WWWUYmp0_2;
	wire w_dff_B_pPgTgPVb9_2;
	wire w_dff_B_b3BVX2oY0_2;
	wire w_dff_B_uUvTNaPX9_2;
	wire w_dff_A_2VNDQKNF4_0;
	wire w_dff_A_VRPZQ8vi8_0;
	wire w_dff_A_K0v8OTU29_0;
	wire w_dff_A_6O5rJf7T4_0;
	wire w_dff_A_6cl3ISZv3_0;
	wire w_dff_A_dLTShI6e4_0;
	wire w_dff_A_lEY5TJhc5_0;
	wire w_dff_A_YSebzq7q0_0;
	wire w_dff_A_EPWGFcJD8_0;
	wire w_dff_A_IVYwyVLb4_0;
	wire w_dff_A_TNf5Xzci9_0;
	wire w_dff_A_SRzfEq2P7_0;
	wire w_dff_A_Sa2BPSPj2_0;
	wire w_dff_A_ZNR42zaU9_0;
	wire w_dff_A_RlohIgWY0_0;
	wire w_dff_A_8YKBPe6X5_0;
	wire w_dff_A_Xs0xBlaI4_0;
	wire w_dff_A_xMwM09Dw7_0;
	wire w_dff_A_ec6FnCUB3_0;
	wire w_dff_A_hTvL5vzG1_0;
	wire w_dff_A_83dePEjo1_1;
	wire w_dff_A_2kmHN2nr2_1;
	wire w_dff_A_bICRxTcp6_1;
	wire w_dff_A_A6pcBdQW9_1;
	wire w_dff_A_dqA1iTsp5_1;
	wire w_dff_A_2p6TzBdR0_1;
	wire w_dff_A_nOdvEM2O8_1;
	wire w_dff_A_lem8xaPx7_1;
	wire w_dff_A_w29xGCwv0_1;
	wire w_dff_A_EyvGYo8f4_1;
	wire w_dff_A_rNyqQz2R0_1;
	wire w_dff_A_ZkEt66zK0_1;
	wire w_dff_A_b8m4tGwy5_1;
	wire w_dff_A_Cja6zkSj7_1;
	wire w_dff_A_lzEL013z8_0;
	wire w_dff_A_HitMEIcW0_0;
	wire w_dff_A_Z1SZBG4I3_0;
	wire w_dff_A_vgxR4BZu9_0;
	wire w_dff_A_OcK3Z1p87_0;
	wire w_dff_A_kJY4IHWD0_0;
	wire w_dff_A_VlCqvEiy4_0;
	wire w_dff_A_3UtBEZuj6_0;
	wire w_dff_A_fHwwK6F40_0;
	wire w_dff_A_UKVnAVN40_0;
	wire w_dff_A_gGr99vMR6_0;
	wire w_dff_A_0CyklLM18_0;
	wire w_dff_B_qUqSm9GJ4_2;
	wire w_dff_B_7fuvmvCx4_2;
	wire w_dff_B_az7TCeYd7_2;
	wire w_dff_B_7RL1TIQc5_2;
	wire w_dff_B_SVdhd0Dc8_2;
	wire w_dff_B_0MyRwGPc8_2;
	wire w_dff_B_D9yHKpXV5_2;
	wire w_dff_B_np3gfNno3_2;
	wire w_dff_B_XoQwXwxj0_2;
	wire w_dff_B_BAQRRF1l2_2;
	wire w_dff_B_5VtNxWne5_2;
	wire w_dff_B_XBhqH1475_2;
	wire w_dff_B_fyrZXCvG0_2;
	wire w_dff_A_P4E9OfrU2_0;
	wire w_dff_A_NfnO9f7r4_0;
	wire w_dff_A_oF9666GH5_0;
	wire w_dff_A_TMJ6cU6F7_0;
	wire w_dff_A_q40O1sGG4_0;
	wire w_dff_A_KdSzsY7L4_0;
	wire w_dff_A_TDSvuKZa7_0;
	wire w_dff_A_Z0zALdGJ2_0;
	wire w_dff_A_14tCVaq02_0;
	wire w_dff_A_9ASsQCif4_0;
	wire w_dff_A_Yb4EtMYG4_0;
	wire w_dff_A_AOjEDhQx8_0;
	wire w_dff_A_NeiQxvBq5_0;
	wire w_dff_A_O0PhjXJJ1_0;
	wire w_dff_A_3DkbUKqV4_0;
	wire w_dff_A_q4PeoTyl5_0;
	wire w_dff_A_32hI6N2n9_0;
	wire w_dff_A_IYUO0ecr1_0;
	wire w_dff_A_11nRX98N3_0;
	wire w_dff_A_T30xqLpp4_0;
	wire w_dff_A_2gpDt1rw1_1;
	wire w_dff_A_z4WWpocZ0_1;
	wire w_dff_A_BiEMJDwr2_1;
	wire w_dff_A_x3s1wrdr0_1;
	wire w_dff_A_CUXDsklJ4_1;
	wire w_dff_A_9Jbz5w6N9_1;
	wire w_dff_A_s6t7iNYI6_1;
	wire w_dff_B_4QZ46xG08_0;
	wire w_dff_B_b6nSR68a2_0;
	wire w_dff_B_NJHj4LJQ3_0;
	wire w_dff_B_cylbLnVE1_0;
	wire w_dff_B_0xlbnkxf7_0;
	wire w_dff_A_kkuwY2iN0_0;
	wire w_dff_A_xEo5DSXc0_0;
	wire w_dff_A_JxBinVoZ4_0;
	wire w_dff_A_nUTgCvt80_0;
	wire w_dff_A_r7iu4eT31_0;
	wire w_dff_A_PZtx4D5a9_0;
	wire w_dff_A_D1zSyuGG8_0;
	wire w_dff_A_4WhcggbI7_0;
	wire w_dff_A_6VDJmKIe8_0;
	wire w_dff_A_AGZU92X91_0;
	wire w_dff_A_7EfEMMAw2_0;
	wire w_dff_A_gn9Dwxgk1_0;
	wire w_dff_A_nbLpy6kM5_0;
	wire w_dff_A_JYv7xi7H3_0;
	wire w_dff_A_Y4jSUqGe3_0;
	wire w_dff_A_1xfANVUj8_0;
	wire w_dff_A_wYFRCQu26_0;
	wire w_dff_A_CHVy6Qct6_0;
	wire w_dff_A_NztlICNx4_0;
	wire w_dff_A_K70pXfwm2_0;
	wire w_dff_A_rhgUzpww6_0;
	wire w_dff_A_lPudnZzQ4_0;
	wire w_dff_A_Tqzg5ZiU4_0;
	wire w_dff_A_is7xcMgr9_0;
	wire w_dff_A_ZSidA31H8_0;
	wire w_dff_A_AdleOg1T4_0;
	wire w_dff_A_2kr83mvm7_0;
	wire w_dff_A_7YB8gEZS0_0;
	wire w_dff_A_72YPSi479_0;
	wire w_dff_A_g7Y78fgg7_0;
	wire w_dff_A_ijzhXmIl2_0;
	wire w_dff_A_5mq645bi0_0;
	wire w_dff_A_vOdb2YxJ8_0;
	wire w_dff_A_Rp8YjN2A0_0;
	wire w_dff_A_wXz8MI1r6_0;
	wire w_dff_A_iPjsRmrz4_0;
	wire w_dff_A_Qiowc9UD7_0;
	wire w_dff_A_eS2VW7jv4_0;
	wire w_dff_A_OYC4wMHD3_0;
	wire w_dff_A_rvv8PztO5_0;
	wire w_dff_A_39boRS979_0;
	wire w_dff_A_NvpKZUwL4_0;
	wire w_dff_A_ySeg3elV5_0;
	wire w_dff_A_CfgtonVu2_0;
	wire w_dff_A_ajlO7iq04_0;
	wire w_dff_B_TULCKkIv7_1;
	wire w_dff_A_lOfZMnf54_0;
	wire w_dff_A_n6hXZ9SH3_0;
	wire w_dff_A_jUYZU3kF9_0;
	wire w_dff_A_gevSWNzF0_0;
	wire w_dff_A_6BGROkuE9_0;
	wire w_dff_A_eV97XeUj9_0;
	wire w_dff_A_Kf3ddpAR8_0;
	wire w_dff_A_AC3V1HOO4_0;
	wire w_dff_A_WE7qvhvl3_0;
	wire w_dff_A_VMbfIxYJ9_0;
	wire w_dff_A_Iyn24Ir93_0;
	wire w_dff_A_1NHobVf29_0;
	wire w_dff_B_OOZQruHx0_1;
	wire w_dff_B_c5c18Uis1_1;
	wire w_dff_B_PVqFOUhM9_1;
	wire w_dff_B_sgkt7iPm9_1;
	wire w_dff_B_5SkpzC2A4_1;
	wire w_dff_B_vuzsV2FC6_1;
	wire w_dff_A_nC9RLLDY4_0;
	wire w_dff_A_fSU0j8Yn2_0;
	wire w_dff_A_5UjwFNuN8_0;
	wire w_dff_A_I0B4DkU05_0;
	wire w_dff_B_DacFIcBk5_2;
	wire w_dff_B_i2Sflq2H1_0;
	wire w_dff_B_SlHUmUsE1_0;
	wire w_dff_B_nQ6YaW0S4_0;
	wire w_dff_B_i8ozyrsk5_0;
	wire w_dff_A_mIghtVWN7_0;
	wire w_dff_A_U6hHS9oy6_0;
	wire w_dff_A_3A1so0WA4_0;
	wire w_dff_A_M2mwOCZz0_0;
	wire w_dff_A_2TjCq7Hh6_0;
	wire w_dff_A_P8mWUwpS3_0;
	wire w_dff_A_X4qN0ZtE2_0;
	wire w_dff_A_ZnHftyNV4_0;
	wire w_dff_A_9cQavNd13_0;
	wire w_dff_A_pbaOLV8f9_0;
	wire w_dff_A_Ar5obENu8_0;
	wire w_dff_A_3fWF9Vay3_0;
	wire w_dff_A_X9fM55LS2_0;
	wire w_dff_A_5Q738wrw6_0;
	wire w_dff_A_DATfAEHS4_0;
	wire w_dff_A_gVjaJtsn2_0;
	wire w_dff_A_bRsrjABE0_0;
	wire w_dff_A_ZOGdPGs42_0;
	wire w_dff_A_upZOs5PZ5_0;
	wire w_dff_A_BdUgGSAh2_0;
	wire w_dff_A_Nc2x7Jwl2_0;
	wire w_dff_A_1mU1ZLEm8_0;
	wire w_dff_A_nl7IyFXG9_0;
	wire w_dff_B_ih3E6Wpi6_2;
	wire w_dff_B_D617FD3g6_2;
	wire w_dff_B_TAsBmQD71_2;
	wire w_dff_B_m9OscV3G6_2;
	wire w_dff_B_0C65iaNx5_2;
	wire w_dff_B_f4x8NmUE9_2;
	wire w_dff_B_6g7kN7jm8_2;
	wire w_dff_B_MybpwxhO4_2;
	wire w_dff_B_Rv3whGh50_2;
	wire w_dff_B_ujhZzmE93_2;
	wire w_dff_B_p9htagI23_2;
	wire w_dff_B_7tnf8wmb0_2;
	wire w_dff_B_IR8Bvya77_2;
	wire w_dff_B_ynVHqGdP0_2;
	wire w_dff_A_3OPq8lC90_0;
	wire w_dff_A_qLM8c9x33_0;
	wire w_dff_A_K8uVWCHg2_0;
	wire w_dff_A_wQUjB8Sy9_0;
	wire w_dff_A_dLf5Wvxq3_0;
	wire w_dff_A_3QiR7ewA2_0;
	wire w_dff_A_iWa6xviI8_0;
	wire w_dff_A_eklnG9MQ6_0;
	wire w_dff_A_GBFYKOkz5_0;
	wire w_dff_A_c63E0tea8_0;
	wire w_dff_A_qMmAYXyr9_0;
	wire w_dff_A_qahQb5Qc7_0;
	wire w_dff_A_FT22x3K41_0;
	wire w_dff_A_FjkyvDqN9_0;
	wire w_dff_A_IcPR62ao3_0;
	wire w_dff_A_dMFpHtVm4_1;
	wire w_dff_A_7bWL3VEH3_1;
	wire w_dff_A_3vDhBz6t5_1;
	wire w_dff_A_d05E4w361_1;
	wire w_dff_A_2wwBRVl54_1;
	wire w_dff_A_iswuUbvY4_1;
	wire w_dff_A_wSS7Uavd7_0;
	wire w_dff_A_ahDzLQV77_0;
	wire w_dff_A_tyBqzzah5_0;
	wire w_dff_A_lkFuCNfX4_0;
	wire w_dff_A_YbFSinoe7_0;
	wire w_dff_A_t3Hryi672_0;
	wire w_dff_A_yj0eJcbk9_0;
	wire w_dff_A_iS7P584Y7_0;
	wire w_dff_A_R5mgsJEh5_0;
	wire w_dff_A_KNtmxcGp2_0;
	wire w_dff_A_FP4D0iMU9_0;
	wire w_dff_A_b787DLJQ7_0;
	wire w_dff_B_3suSYngp4_2;
	wire w_dff_B_ryLnhs7O7_2;
	wire w_dff_B_nck2wWvV9_2;
	wire w_dff_B_SgbJxtLR8_2;
	wire w_dff_B_1bgoMqsc2_2;
	wire w_dff_B_4737DIKd2_2;
	wire w_dff_B_oJ0khUTh6_2;
	wire w_dff_A_CBhlU5Vi0_0;
	wire w_dff_A_Rhp8TIeZ8_0;
	wire w_dff_A_hqIttyzW7_0;
	wire w_dff_A_ggH5p7q20_0;
	wire w_dff_A_4LvNKKTI7_0;
	wire w_dff_A_2Aj9k8949_0;
	wire w_dff_A_WvQViioJ4_0;
	wire w_dff_A_36KIvm9k9_0;
	wire w_dff_A_rrQ8oGqq8_0;
	wire w_dff_A_grHjRU1c6_0;
	wire w_dff_A_38u79YLn2_0;
	wire w_dff_A_Ip7mFw6K8_0;
	wire w_dff_A_ylJ6p2Hj3_0;
	wire w_dff_A_lpLg8iFg3_0;
	wire w_dff_A_tbpptluP1_0;
	wire w_dff_A_MxJo78O71_0;
	wire w_dff_A_LPShTF3E9_0;
	wire w_dff_A_YLc1MDH15_0;
	wire w_dff_A_TfSFkQUk7_0;
	wire w_dff_A_4L7SPVuI9_0;
	wire w_dff_A_qKQ1EjVd3_1;
	wire w_dff_A_CWr6yg7X2_1;
	wire w_dff_A_OPhQx6q53_1;
	wire w_dff_A_YDMdgSf06_1;
	wire w_dff_A_NHH8y1P76_0;
	wire w_dff_A_dy9ywEpf3_0;
	wire w_dff_A_4Yn67P8E2_0;
	wire w_dff_A_36qhM1LE6_0;
	wire w_dff_A_rqGOiAIo8_0;
	wire w_dff_A_jggaCk2R5_0;
	wire w_dff_A_TH3VM6Wq8_0;
	wire w_dff_B_L8xAIm631_1;
	wire w_dff_B_5HVIxTto7_1;
	wire w_dff_A_KvN69eRv0_0;
	wire w_dff_A_8qC8Bxil9_0;
	wire w_dff_A_Ahft7AOV4_0;
	wire w_dff_A_EvMmlDyf5_0;
	wire w_dff_A_0KBaRO998_0;
	wire w_dff_A_HxjKhfpm3_0;
	wire w_dff_A_FYfj79HQ6_0;
	wire w_dff_A_nqUp2RTk9_0;
	wire w_dff_A_5TRk2knt2_0;
	wire w_dff_A_55IHtMGb3_0;
	wire w_dff_A_ikW0gD047_0;
	wire w_dff_A_rvw2qnGv6_1;
	wire w_dff_A_LzYGizPC2_1;
	wire w_dff_A_SrzJZZRR9_1;
	wire w_dff_A_8EMDDm7r3_1;
	wire w_dff_A_Ss3t7B913_1;
	wire w_dff_B_esKR7kkk1_3;
	wire w_dff_B_yQY2moTH4_3;
	wire w_dff_B_oeXp4PmU3_3;
	wire w_dff_B_ttlJSbP61_3;
	wire w_dff_B_Qfl55UKq8_3;
	wire w_dff_B_mKkf82ms6_3;
	wire w_dff_B_duBsfNaE5_3;
	wire w_dff_A_hnpq7YPZ0_0;
	wire w_dff_A_6ZzR6NVO8_0;
	wire w_dff_A_IhUCNGIH8_0;
	wire w_dff_A_yaCqGn8t2_0;
	wire w_dff_A_unDrCpin6_0;
	wire w_dff_A_alPvvsFh2_0;
	wire w_dff_A_Mr5eIYlc5_0;
	wire w_dff_A_6wYury1T2_0;
	wire w_dff_A_vz536jsF4_1;
	wire w_dff_A_zOFjjEo51_1;
	wire w_dff_A_OjvD6dLG8_1;
	wire w_dff_A_JjBEHFzh0_1;
	wire w_dff_A_GIjglU9u6_1;
	wire w_dff_A_elrsTPmC6_1;
	wire w_dff_A_gzX4iWzT6_1;
	wire w_dff_A_wf3DvDfL8_1;
	wire w_dff_A_WHh6n79A7_1;
	wire w_dff_A_LSGuI2nP5_1;
	wire w_dff_A_MIwgaU5U1_1;
	wire w_dff_A_BmWdvScP5_1;
	wire w_dff_A_ylkeI8A80_1;
	wire w_dff_A_P90YzDTl9_2;
	wire w_dff_A_kkPlUJ2S0_2;
	wire w_dff_A_boGCpCYk7_2;
	wire w_dff_A_r0km9SAv1_2;
	wire w_dff_A_cbe27X4j3_2;
	wire w_dff_A_FtHp9jB85_2;
	wire w_dff_A_1cc9wIDL4_2;
	wire w_dff_A_2S56qNHh7_2;
	wire w_dff_A_ngVAlWUj2_2;
	wire w_dff_A_1LyjpzAE0_2;
	wire w_dff_A_8bhxMlF20_2;
	wire w_dff_A_CgRXMc1o9_2;
	wire w_dff_A_8CzVoGhG7_2;
	wire w_dff_A_pCSGokb38_0;
	wire w_dff_A_IWZY9deA1_0;
	wire w_dff_A_Qx3ogJgN7_0;
	wire w_dff_A_xCyHPCLS3_0;
	wire w_dff_A_dRSkMPP55_0;
	wire w_dff_A_nFqf8QzF1_0;
	wire w_dff_A_2zuZ6jFB0_0;
	wire w_dff_A_D64y7Lok3_0;
	wire w_dff_A_nfY9ctfx9_0;
	wire w_dff_A_6DMYWMBQ7_0;
	wire w_dff_A_QLBicpOR7_0;
	wire w_dff_A_C7ESVwgH7_1;
	wire w_dff_A_SNot2wgA3_1;
	wire w_dff_A_p5ML6ha55_1;
	wire w_dff_A_sgt5feMI3_1;
	wire w_dff_A_u7RDWOiz3_1;
	wire w_dff_B_7iFtbWKM7_3;
	wire w_dff_B_uckc6IQQ9_3;
	wire w_dff_B_GtsIZzQw2_3;
	wire w_dff_B_QL9zLZh95_3;
	wire w_dff_B_C9hIiv3k6_3;
	wire w_dff_B_DnfFyvX56_3;
	wire w_dff_B_SWO0A4BS1_3;
	wire w_dff_A_kcobK8Is2_0;
	wire w_dff_A_CQM9eZFe7_0;
	wire w_dff_A_slPQWZ2C3_0;
	wire w_dff_A_TFALbzua9_0;
	wire w_dff_A_9EKSZZo06_0;
	wire w_dff_A_cjXAEE6s3_0;
	wire w_dff_A_BtYnkijl0_0;
	wire w_dff_A_zpvm1eo74_0;
	wire w_dff_A_yvnGjsRs8_1;
	wire w_dff_A_rw8qT8P43_1;
	wire w_dff_A_jlDVpJ7x8_1;
	wire w_dff_A_bOKXQDzp5_1;
	wire w_dff_A_ve1rEFdc6_1;
	wire w_dff_A_sVMokOZU3_1;
	wire w_dff_A_KFc4OUjj6_1;
	wire w_dff_A_GPzwGosk0_1;
	wire w_dff_A_lRCmjHhC6_1;
	wire w_dff_A_0xwpSxdc4_1;
	wire w_dff_A_4OjroygO6_1;
	wire w_dff_A_xsWauW9u4_1;
	wire w_dff_A_3RY14p7Q2_1;
	wire w_dff_A_ABVZFhL37_2;
	wire w_dff_A_zuVWxMWC9_2;
	wire w_dff_A_WNcFqDLe9_2;
	wire w_dff_A_fzOGFt1a7_2;
	wire w_dff_A_ubA3NRgw2_2;
	wire w_dff_A_OOhARacv6_2;
	wire w_dff_A_hE7n0a4I7_2;
	wire w_dff_A_UoDmrJph5_2;
	wire w_dff_A_zIohYmyg3_2;
	wire w_dff_A_Bq1laqnH5_2;
	wire w_dff_A_RsgW4ij96_2;
	wire w_dff_A_ktF3Za192_2;
	wire w_dff_A_kTePh0YY1_2;
	wire w_dff_B_rsRN4gi21_0;
	wire w_dff_A_DD2EwS6E1_1;
	wire w_dff_A_3mO9yJA19_1;
	wire w_dff_A_GqZtSLYu0_1;
	wire w_dff_A_LNLRBGh42_1;
	wire w_dff_A_0GVK19w73_1;
	wire w_dff_A_EUSJa4NQ3_0;
	wire w_dff_A_UzJrRbZe3_0;
	wire w_dff_A_vFgpuMpX8_0;
	wire w_dff_A_jJt15PHk3_0;
	wire w_dff_A_gObTqNUE4_0;
	wire w_dff_A_jE8scXq03_0;
	wire w_dff_A_qyEOFRol2_0;
	wire w_dff_A_RezMjxAs2_0;
	wire w_dff_A_s2sk7ri67_0;
	wire w_dff_A_0Hp699qs0_0;
	wire w_dff_A_4bkjgAZJ1_0;
	wire w_dff_A_cENlmcPz9_0;
	wire w_dff_A_7wffRQjy9_0;
	wire w_dff_B_Fv6m2CzD8_1;
	wire w_dff_B_TmclbHEC8_1;
	wire w_dff_B_KBCDqDzO1_1;
	wire w_dff_B_YhorwD8j4_1;
	wire w_dff_B_wKH6W4uK7_1;
	wire w_dff_B_aokus66T8_1;
	wire w_dff_B_u6r39nYs8_1;
	wire w_dff_A_it2qwHqH0_0;
	wire w_dff_A_qwn3zPLH3_0;
	wire w_dff_A_cyDwvHrD6_0;
	wire w_dff_A_wHUrBUHx2_0;
	wire w_dff_A_tm1iovNG2_0;
	wire w_dff_A_fOcwSh3o6_0;
	wire w_dff_A_ECDtJwif4_0;
	wire w_dff_A_2GhpTHQo1_0;
	wire w_dff_A_2S4R9faL7_0;
	wire w_dff_A_ODmWjlRV5_0;
	wire w_dff_A_rd3Fba8s6_0;
	wire w_dff_A_tko4XCxQ2_0;
	wire w_dff_A_tKksQxqR6_0;
	wire w_dff_A_KEyb8s4Y9_1;
	wire w_dff_A_U5B2XVT57_1;
	wire w_dff_A_tgiBVSHu4_1;
	wire w_dff_A_eucTybFG0_1;
	wire w_dff_A_dyrbwCaQ3_1;
	wire w_dff_A_zPHajorB1_1;
	wire w_dff_A_0r1rFZJN2_1;
	wire w_dff_A_gtyfAx5u2_1;
	wire w_dff_A_lyQsZuTS8_0;
	wire w_dff_A_8PsZVu7s4_0;
	wire w_dff_A_4x2ufxxD8_0;
	wire w_dff_A_5P6RYtYA6_0;
	wire w_dff_A_z7doHYr38_0;
	wire w_dff_A_bU20rqy65_0;
	wire w_dff_A_O709u4Bz7_0;
	wire w_dff_A_2iAQPlyp8_0;
	wire w_dff_A_hiYXJa653_0;
	wire w_dff_A_ZkJX8wsO7_0;
	wire w_dff_A_O1gGKJgq3_0;
	wire w_dff_A_w1nJKGU09_0;
	wire w_dff_A_GsPdezS24_0;
	wire w_dff_A_EZTCzFBR7_0;
	wire w_dff_A_hAAFYBmp5_0;
	wire w_dff_A_kAASZgl22_0;
	wire w_dff_A_XCqU0mN41_0;
	wire w_dff_A_ay6l1FQL0_0;
	wire w_dff_A_doOqM7bH5_0;
	wire w_dff_A_Ctzd03QN7_0;
	wire w_dff_A_kTjO4ryG8_0;
	wire w_dff_A_2Esfz2Cc2_2;
	wire w_dff_A_kA7UKfZ70_2;
	wire w_dff_A_FNMcSjCE6_2;
	wire w_dff_A_Sf7DTXvw4_2;
	wire w_dff_A_IodsmCM40_2;
	wire w_dff_A_OGXhtmPX5_2;
	wire w_dff_A_PJ5ac82i5_2;
	wire w_dff_A_HLRxu9hC8_2;
	wire w_dff_A_pdZLw88M9_0;
	wire w_dff_A_3T5QZSFe4_0;
	wire w_dff_A_Ix1wpVIR0_0;
	wire w_dff_A_QAVbQ8KG3_0;
	wire w_dff_A_ousPHLrB5_0;
	wire w_dff_A_riHUICMo6_0;
	wire w_dff_A_1BCrSjlV2_0;
	wire w_dff_A_ad8fcmtR1_0;
	wire w_dff_A_XH5Xx23o7_0;
	wire w_dff_A_MJcv7u0l3_0;
	wire w_dff_A_Klo8Z9nq0_0;
	wire w_dff_B_vbNPuuRj4_2;
	wire w_dff_B_wXu0phGn4_2;
	wire w_dff_B_TC71sZVX0_2;
	wire w_dff_B_riSjZN5b5_2;
	wire w_dff_B_yXinODag7_2;
	wire w_dff_B_Qo2yRTwU3_2;
	wire w_dff_B_Qpnbjv8i6_2;
	wire w_dff_A_1jLi4RYx1_0;
	wire w_dff_A_hdwRdQAI2_0;
	wire w_dff_A_I0FAqYFk4_0;
	wire w_dff_A_RPQm22uG9_0;
	wire w_dff_A_ToZX8LuQ5_0;
	wire w_dff_A_Eqvtuz0k7_0;
	wire w_dff_A_9Iq4itu71_0;
	wire w_dff_A_hgpJNaHG9_0;
	wire w_dff_A_GEyPZXY59_0;
	wire w_dff_A_85mXJdqJ6_0;
	wire w_dff_A_XiE6s5Pe4_0;
	wire w_dff_A_OxhLI8F16_0;
	wire w_dff_A_Uf4wyVZi1_0;
	wire w_dff_A_bmHSz2Tj0_1;
	wire w_dff_A_qlobzmpw6_1;
	wire w_dff_A_R441xY9b2_1;
	wire w_dff_A_V0yOCIhw4_1;
	wire w_dff_A_gGJtaM9k0_1;
	wire w_dff_A_bRpoo7C77_1;
	wire w_dff_A_0C47CxO73_1;
	wire w_dff_A_LFlt7WTf2_1;
	wire w_dff_B_FIU4XNhX5_1;
	wire w_dff_B_E79sbgNT4_1;
	wire w_dff_B_sox4Yx8h2_1;
	wire w_dff_B_BH8cCgRW1_1;
	wire w_dff_B_1PvCAizf9_1;
	wire w_dff_B_IY29OhhM2_1;
	wire w_dff_B_4aXRGgFB2_1;
	wire w_dff_A_Bl0vePuy3_0;
	wire w_dff_A_WPByknKX0_0;
	wire w_dff_A_psbqyxzE7_0;
	wire w_dff_A_vAiuKXTl7_0;
	wire w_dff_A_YDBVrOPt0_0;
	wire w_dff_A_KHOofYdl2_0;
	wire w_dff_A_BlT9XUv15_0;
	wire w_dff_A_4MmouBb57_0;
	wire w_dff_A_ryZQ9wY16_1;
	wire w_dff_A_NzIrbV8u5_1;
	wire w_dff_A_NumHLs2G7_1;
	wire w_dff_A_mZHBZK701_1;
	wire w_dff_A_70pygJTa6_1;
	wire w_dff_A_PNlwz2hy0_1;
	wire w_dff_A_5DxUnceN5_1;
	wire w_dff_A_u0Reuen91_1;
	wire w_dff_A_3S0Noii19_1;
	wire w_dff_A_HOdmcer34_1;
	wire w_dff_A_Js6aPtXj6_1;
	wire w_dff_A_ixIbOInX5_1;
	wire w_dff_A_3q3Udb6f2_1;
	wire w_dff_A_3WhSAtBC6_0;
	wire w_dff_A_C4yHK1bg7_0;
	wire w_dff_A_OHNi3BtC2_0;
	wire w_dff_A_tmvUf1fZ7_0;
	wire w_dff_A_vry5MGvC5_0;
	wire w_dff_A_FycskBfx6_0;
	wire w_dff_A_WYcYWevu1_0;
	wire w_dff_A_bNclPy5R3_0;
	wire w_dff_A_SBDThDsY3_0;
	wire w_dff_A_buxUTz049_0;
	wire w_dff_A_QQALszhd2_0;
	wire w_dff_B_3SWlJP7U6_2;
	wire w_dff_B_H7EoF3O72_2;
	wire w_dff_B_f6U0AA6u9_2;
	wire w_dff_B_jiu8K6Mv4_2;
	wire w_dff_B_h5wiugK65_2;
	wire w_dff_B_0L1AhYIW6_2;
	wire w_dff_B_zzOnSQo75_2;
	wire w_dff_A_pKoZdVtq3_0;
	wire w_dff_A_LBmYrF4v2_0;
	wire w_dff_A_vkLkEUDb0_0;
	wire w_dff_A_8nGOXfmL3_0;
	wire w_dff_A_tckeineN2_0;
	wire w_dff_A_V0OZ0ex87_0;
	wire w_dff_A_RAQ7soBi6_0;
	wire w_dff_A_3gY0AY0h1_0;
	wire w_dff_A_stDXda203_0;
	wire w_dff_A_4wrPObSd0_0;
	wire w_dff_A_inT0k7Z87_0;
	wire w_dff_A_5z3gmTeW9_0;
	wire w_dff_A_BF8gCdAp4_0;
	wire w_dff_A_MGDYFj995_1;
	wire w_dff_A_2T4XnEqm3_1;
	wire w_dff_A_Gm0vMFkY0_1;
	wire w_dff_A_n64ETrL61_1;
	wire w_dff_A_s1VW2A2j8_1;
	wire w_dff_A_mPsWAnai9_1;
	wire w_dff_A_iXdroaPO2_1;
	wire w_dff_A_6l4mxBtJ8_1;
	wire w_dff_A_ZAq4GogY7_0;
	wire w_dff_A_Zjd3FBVm9_0;
	wire w_dff_A_hP8e5VEY4_0;
	wire w_dff_A_E5jsua8o5_0;
	wire w_dff_A_x77Iu3pY1_0;
	wire w_dff_A_F1VAy6oj4_0;
	wire w_dff_B_1g27YgFr7_1;
	wire w_dff_B_7jHgBMXL3_1;
	wire w_dff_A_YS5WvG4O8_0;
	wire w_dff_A_RdscfmSd6_0;
	wire w_dff_A_vs4Yte5a6_0;
	wire w_dff_A_McmLrzke5_0;
	wire w_dff_A_TTdqR00b8_0;
	wire w_dff_A_vcoSxdJH7_0;
	wire w_dff_A_FNBBFI7k1_0;
	wire w_dff_A_egyvezmP1_0;
	wire w_dff_A_KAqRUqc41_0;
	wire w_dff_A_tNomMc159_0;
	wire w_dff_A_xxDRcru73_0;
	wire w_dff_A_t6pyZeN27_0;
	wire w_dff_A_0tDbL01y9_0;
	wire w_dff_A_QgsUMgbR2_0;
	wire w_dff_A_zSvERz9r7_0;
	wire w_dff_A_D8HQEZDm7_0;
	wire w_dff_A_VUMppq5o2_0;
	wire w_dff_A_PftCV0974_0;
	wire w_dff_A_H77QyUzX6_0;
	wire w_dff_A_ikqDVpKe9_0;
	wire w_dff_A_6IvXc7H93_0;
	wire w_dff_A_IEeZPfcm7_0;
	wire w_dff_A_E3m0gHHM1_0;
	wire w_dff_A_0iX5VOvF3_0;
	wire w_dff_A_0KSjwQtd3_0;
	wire w_dff_A_tJBtmbww6_0;
	wire w_dff_A_KIGRHkPL2_0;
	wire w_dff_A_3oa89vUu6_0;
	wire w_dff_A_CAjglNfV7_0;
	wire w_dff_A_OU2Z0wSZ9_0;
	wire w_dff_A_LbP9gmM75_0;
	wire w_dff_A_qKygx8oj3_0;
	wire w_dff_A_H49QXB351_0;
	wire w_dff_A_DQdR1sTx9_0;
	wire w_dff_A_0WKc5XU48_0;
	wire w_dff_A_1eDK6lYR9_0;
	wire w_dff_A_b8Ik8HGI4_0;
	wire w_dff_A_d4CkhFFo4_0;
	wire w_dff_A_Km5hpih89_0;
	wire w_dff_A_p5hPemGS8_0;
	wire w_dff_A_wgydJpYc2_0;
	wire w_dff_A_Fevppzgi7_0;
	wire w_dff_A_4rThsRKZ8_0;
	wire w_dff_A_mjNe2c9q6_0;
	wire w_dff_A_UN8sB5N10_0;
	wire w_dff_A_cQUYckR48_0;
	wire w_dff_A_vyhN0RL21_0;
	wire w_dff_A_XmSAc9Y30_0;
	wire w_dff_A_nPf3tF7K5_0;
	wire w_dff_A_im35mc7u0_0;
	wire w_dff_A_ibEiz88q1_0;
	wire w_dff_A_NQDn57kM7_0;
	wire w_dff_A_k8AqYqB49_0;
	wire w_dff_A_UEpzuz7S1_0;
	wire w_dff_A_9tiFhrMz9_0;
	wire w_dff_B_N7AGX4IP8_2;
	wire w_dff_B_6G06KosA9_2;
	wire w_dff_B_KOAIJrsW4_2;
	wire w_dff_B_B4a7me5l3_2;
	wire w_dff_B_fHVpo0DQ5_2;
	wire w_dff_B_YCdv7NHY3_2;
	wire w_dff_B_R69DaiPJ4_2;
	wire w_dff_A_68eKiuOq4_0;
	wire w_dff_A_7s7x76Wm0_0;
	wire w_dff_A_5VbRwkNE8_0;
	wire w_dff_A_DyW161X97_0;
	wire w_dff_A_W2PdFSHR5_0;
	wire w_dff_A_D6w4JkDp7_0;
	wire w_dff_A_8JH5ryuG1_0;
	wire w_dff_A_bNWg9gOY3_0;
	wire w_dff_A_5LwtncGv2_0;
	wire w_dff_A_SY7nT9p57_0;
	wire w_dff_A_qDDjToK53_0;
	wire w_dff_A_MEWjSqDL2_0;
	wire w_dff_A_y0ynk3B09_0;
	wire w_dff_A_aPcuxAQt9_1;
	wire w_dff_A_j4NiqdiA4_1;
	wire w_dff_A_ggz7T9v59_1;
	wire w_dff_A_QceUSftn8_1;
	wire w_dff_A_q5xRitIL5_1;
	wire w_dff_A_tXyKoq2u0_1;
	wire w_dff_A_PidPrwjK1_1;
	wire w_dff_A_nAPqZLqT6_1;
	wire w_dff_A_gJ6hF6OQ1_1;
	wire w_dff_A_SqMnunAP0_1;
	wire w_dff_A_x8GueNsS5_1;
	wire w_dff_A_69bqsicp0_1;
	wire w_dff_A_VEwuRhUd5_1;
	wire w_dff_A_8uzRIjdi1_1;
	wire w_dff_B_psk07u3V0_1;
	wire w_dff_B_oqycvCM21_1;
	wire w_dff_A_MMSOLrkf9_0;
	wire w_dff_A_EmbrQ3OK4_0;
	wire w_dff_A_5EwA2DpY9_0;
	wire w_dff_A_sSsn89L83_0;
	wire w_dff_A_5ABIk3ha6_0;
	wire w_dff_A_Rd3Iqsut7_0;
	wire w_dff_A_B0KcFS5N3_0;
	wire w_dff_A_OXR4KdRt3_2;
	wire w_dff_A_HGZVjoyq2_0;
	wire w_dff_A_y3JgxNnQ8_0;
	wire w_dff_A_xSbHDy8M1_0;
	wire w_dff_A_Zh6Zzmpx9_0;
	wire w_dff_A_GHmMaPQz1_0;
	wire w_dff_A_zxg6pJ4q5_0;
	wire w_dff_A_KlkLvP1s6_0;
	wire w_dff_A_l6Ex0cdx4_0;
	wire w_dff_A_wQCdnG0t0_0;
	wire w_dff_A_unlN3uPJ9_0;
	wire w_dff_A_qMJdKDQo4_0;
	wire w_dff_A_A24A1gXq5_1;
	wire w_dff_A_poMtGWKM2_0;
	wire w_dff_A_BGrAfOEQ2_0;
	wire w_dff_A_KOnpoR7X3_0;
	wire w_dff_A_xyIwAmPi0_0;
	wire w_dff_A_0ee1nJSj0_0;
	wire w_dff_A_mXeuhKAh9_0;
	wire w_dff_A_WiEggLot0_0;
	wire w_dff_A_k2SMsEB40_0;
	wire w_dff_A_Pdt8fVrR5_0;
	wire w_dff_A_Xslwsn9A7_0;
	wire w_dff_A_VTHH7CAn5_0;
	wire w_dff_A_wx4vqfXc1_1;
	wire w_dff_A_OtuWHIYh9_0;
	wire w_dff_A_CQZXVABP2_0;
	wire w_dff_A_t8svVLG17_0;
	wire w_dff_A_4DJWQcyM2_0;
	wire w_dff_A_Gj9lJwna2_0;
	wire w_dff_A_fsi7MOdP6_0;
	wire w_dff_A_MpS27uXT9_0;
	wire w_dff_A_LTw6E6Ql5_2;
	wire w_dff_A_b7HwALh75_0;
	wire w_dff_A_tUTfemSi8_0;
	wire w_dff_A_1qWtbnpy2_0;
	wire w_dff_A_ZnTlYI2p8_0;
	wire w_dff_A_bmwWrFaJ6_0;
	wire w_dff_A_SbywBC6r8_0;
	wire w_dff_A_2oG41Q1J2_0;
	wire w_dff_A_368eFpuS7_0;
	wire w_dff_A_EeKppYKU2_0;
	wire w_dff_A_e8Vraddr0_0;
	wire w_dff_A_XquBIlvv5_0;
	wire w_dff_A_o0bLKkPz9_1;
	wire w_dff_A_sxEaZZfL4_0;
	wire w_dff_A_3uv68hd12_0;
	wire w_dff_A_tMi8ojkN1_0;
	wire w_dff_A_gOAH3kGN4_0;
	wire w_dff_A_1NtzMFup5_0;
	wire w_dff_A_saW5UnnJ7_0;
	wire w_dff_A_Z5ttAmgn2_0;
	wire w_dff_A_WgCxUncS6_2;
	wire w_dff_A_zpHSg7Vy4_0;
	wire w_dff_A_LL1rQsT87_0;
	wire w_dff_A_KVTmalWt2_0;
	wire w_dff_A_5OMAOq8G4_0;
	wire w_dff_A_UoMNT9Qa5_0;
	wire w_dff_A_C4ohPfNl4_0;
	wire w_dff_A_iUHYDX1B0_0;
	wire w_dff_A_PWJzbRI75_0;
	wire w_dff_A_2ulqc1dc6_0;
	wire w_dff_A_KjHMfl831_0;
	wire w_dff_A_VjTQ0GMX3_0;
	wire w_dff_A_uTzSJXu04_1;
	wire w_dff_A_fBEA9jxP0_0;
	wire w_dff_A_OLfa3rfG0_0;
	wire w_dff_A_5EXQ7Kn36_0;
	wire w_dff_A_zK5BxrtN3_0;
	wire w_dff_A_isRDBUU88_0;
	wire w_dff_A_dvRx08Gc4_0;
	wire w_dff_A_Ge8B9hJt4_0;
	wire w_dff_A_4g578riZ3_2;
	wire w_dff_A_BWUVzlYy0_0;
	wire w_dff_A_iqYffsIx4_0;
	wire w_dff_A_7HGOLgLQ0_0;
	wire w_dff_A_8un81v9g3_0;
	wire w_dff_A_QQxypFdR7_0;
	wire w_dff_A_cOVi5QN32_0;
	wire w_dff_A_38LifaDN7_0;
	wire w_dff_A_zy3GkgzL0_0;
	wire w_dff_A_VMN1DwnB5_0;
	wire w_dff_A_IO7KywT24_0;
	wire w_dff_A_HZbKt9s03_0;
	wire w_dff_A_U0O983TN1_1;
	wire w_dff_A_9XmdiHfa7_0;
	wire w_dff_A_kxm4TQ1o1_0;
	wire w_dff_A_9EIHA2mN8_0;
	wire w_dff_A_3ykacEbC4_0;
	wire w_dff_A_wAnMmerE8_1;
	wire w_dff_A_xghP78uJ2_1;
	wire w_dff_A_Pjmk4a686_2;
	wire w_dff_A_rMRatPpU3_0;
	wire w_dff_A_vKMgwbGJ8_0;
	wire w_dff_A_msD5FqKo8_0;
	wire w_dff_A_9KzMed2U8_0;
	wire w_dff_A_baAoJW3O6_0;
	wire w_dff_A_N4JjRjiX8_0;
	wire w_dff_A_iK9sgUV75_1;
	wire w_dff_A_DbMQvbvi3_0;
	wire w_dff_A_KSeK94Xh3_0;
	wire w_dff_A_RUCOTxEn2_0;
	wire w_dff_A_yjFjDUBe5_0;
	wire w_dff_A_nAqjQpYU9_0;
	wire w_dff_A_IAVnKPJE6_0;
	wire w_dff_A_xXeOIwou4_0;
	wire w_dff_A_eny0RcZF5_2;
	wire w_dff_A_cjWThgh89_0;
	wire w_dff_A_KRiWLSeP7_0;
	wire w_dff_A_thtnU7wY1_0;
	wire w_dff_A_PSEeBRYd0_0;
	wire w_dff_A_jrm4zwtG2_0;
	wire w_dff_A_n9yPRBbA0_0;
	wire w_dff_A_YqfOQ8zT2_0;
	wire w_dff_A_s83XpgJt9_0;
	wire w_dff_A_ZFI4vkSL7_0;
	wire w_dff_A_mtSJ8G1E7_0;
	wire w_dff_A_MQd5T3JC6_0;
	wire w_dff_A_scHdCel47_1;
	wire w_dff_A_vq767C681_1;
	wire w_dff_A_8fNpvyNO4_0;
	wire w_dff_A_DMrYvpqC1_1;
	wire w_dff_A_G8whc0Pr5_1;
	wire w_dff_A_JHlZvLiu2_1;
	wire w_dff_A_y1wdbJ7V5_1;
	wire w_dff_A_RTUJgqj54_1;
	wire w_dff_A_rZNTymzR4_1;
	wire w_dff_A_YrRtR3Ve0_1;
	wire w_dff_A_7hgsGo9G1_1;
	wire w_dff_A_iYOw4pOk9_2;
	wire w_dff_A_a5LUy0Jh0_0;
	wire w_dff_A_lmUF8aNa7_0;
	wire w_dff_A_9aYZ00BV6_0;
	wire w_dff_A_58tyhiZ74_0;
	wire w_dff_A_1S6iYLtK3_0;
	wire w_dff_A_kmbyvGTf0_0;
	wire w_dff_A_WsAkDPUO5_0;
	wire w_dff_A_JODcJSlN7_0;
	wire w_dff_A_RgKDmBCP5_0;
	wire w_dff_A_3N6aZG4V1_0;
	wire w_dff_A_Z8LXqTPZ1_0;
	wire w_dff_A_PUZJsGRG5_0;
	wire w_dff_A_Vr9TnkqD2_0;
	wire w_dff_A_jdyjcmOa7_0;
	wire w_dff_A_E9ik2gEm3_0;
	wire w_dff_A_g0XFfzZl5_0;
	wire w_dff_A_st7JVpjz6_0;
	wire w_dff_A_gp6QfW5O2_0;
	wire w_dff_A_retoFnjf2_0;
	wire w_dff_A_pN3ggmc15_0;
	wire w_dff_A_I6MPMl0M1_0;
	wire w_dff_A_j00AEJWg8_0;
	wire w_dff_A_nGIOe9D07_0;
	wire w_dff_A_F2J5LdON6_0;
	wire w_dff_A_AcISA6RU7_2;
	wire w_dff_A_tkBIfQCV9_1;
	wire w_dff_A_YC0wFypt7_1;
	wire w_dff_A_HMT7AyUD1_1;
	wire w_dff_A_rIMszMo84_1;
	wire w_dff_A_B6clcUBo2_1;
	wire w_dff_A_5HP8BIJ01_1;
	wire w_dff_A_fDZDKLkV4_1;
	wire w_dff_A_y6qefsw96_1;
	wire w_dff_A_R2AnmVBV4_1;
	wire w_dff_A_lxZPLhBu6_1;
	wire w_dff_A_KdNP7kkJ2_1;
	wire w_dff_A_0Re8soi95_1;
	wire w_dff_A_2gHoIhD52_1;
	wire w_dff_A_wxwzoTvF1_1;
	wire w_dff_A_PYJI8UMC6_1;
	wire w_dff_A_MaxiYCp89_2;
	wire w_dff_A_4a1iUSTY4_0;
	wire w_dff_A_RxCxpIGD6_0;
	wire w_dff_A_QWADezyW3_0;
	wire w_dff_A_uL6REXsy7_0;
	wire w_dff_A_NAzGTNyg9_0;
	wire w_dff_A_G2P8yfdL6_0;
	wire w_dff_A_auaaU9JO5_0;
	wire w_dff_A_Z928laBU1_0;
	wire w_dff_A_iTGutd682_0;
	wire w_dff_A_h0b9DVmg1_0;
	wire w_dff_A_7RCADPY52_0;
	wire w_dff_A_VWaVx4QM1_0;
	wire w_dff_A_51UUfiLp3_0;
	wire w_dff_A_CKJaqjPo3_0;
	wire w_dff_A_sgcmtF7V4_0;
	wire w_dff_A_okGHrDh63_0;
	wire w_dff_A_B9DHgZ8K7_0;
	wire w_dff_A_cjO7Z7sD3_0;
	wire w_dff_A_GlggAXEA0_0;
	wire w_dff_A_R3l9X8Gn8_1;
	wire w_dff_A_Gw6NYGQ52_0;
	wire w_dff_A_4ifcTakD8_0;
	wire w_dff_A_qQXOIv9C2_0;
	wire w_dff_A_BWbWi0ka0_0;
	wire w_dff_A_w4Gaq2Dg0_0;
	wire w_dff_A_0k8GlC1P6_0;
	wire w_dff_A_QsnA1HsA9_0;
	wire w_dff_A_FJfEB19U4_0;
	wire w_dff_A_CfF1bmPV9_0;
	wire w_dff_A_4ZYY7OJs4_0;
	wire w_dff_A_ALrhgiIh9_0;
	wire w_dff_A_zl0zYyGv5_0;
	wire w_dff_A_cgYnHa567_1;
	wire w_dff_A_KJlCgD6r5_0;
	wire w_dff_A_FiOshWDZ9_0;
	wire w_dff_A_wAmORMbX5_0;
	wire w_dff_A_ZswGhIHK6_0;
	wire w_dff_A_vrpEtuVb5_0;
	wire w_dff_A_RCUy6P1j0_1;
	wire w_dff_A_9J82KA3Q7_0;
	jnot g000(.din(w_G76gat_0[1]),.dout(n43),.clk(gclk));
	jand g001(.dina(w_G82gat_0[2]),.dinb(w_n43_0[1]),.dout(n44),.clk(gclk));
	jnot g002(.din(w_G24gat_0[1]),.dout(n45),.clk(gclk));
	jand g003(.dina(w_G30gat_0[1]),.dinb(n45),.dout(n46),.clk(gclk));
	jnot g004(.din(w_G11gat_0[2]),.dout(n47),.clk(gclk));
	jand g005(.dina(w_G17gat_0[2]),.dinb(w_n47_0[1]),.dout(n48),.clk(gclk));
	jor g006(.dina(n48),.dinb(n46),.dout(n49),.clk(gclk));
	jor g007(.dina(n49),.dinb(w_n44_0[1]),.dout(n50),.clk(gclk));
	jnot g008(.din(w_G37gat_0[2]),.dout(n51),.clk(gclk));
	jand g009(.dina(w_G43gat_1[1]),.dinb(n51),.dout(n52),.clk(gclk));
	jnot g010(.din(w_G63gat_0[2]),.dout(n53),.clk(gclk));
	jand g011(.dina(w_G69gat_0[2]),.dinb(w_n53_0[1]),.dout(n54),.clk(gclk));
	jor g012(.dina(n54),.dinb(w_n52_0[1]),.dout(n55),.clk(gclk));
	jnot g013(.din(w_G102gat_0[2]),.dout(n56),.clk(gclk));
	jand g014(.dina(w_G108gat_0[2]),.dinb(w_n56_0[1]),.dout(n57),.clk(gclk));
	jnot g015(.din(w_G50gat_0[2]),.dout(n58),.clk(gclk));
	jand g016(.dina(w_G56gat_0[2]),.dinb(w_n58_0[1]),.dout(n59),.clk(gclk));
	jor g017(.dina(n59),.dinb(n57),.dout(n60),.clk(gclk));
	jnot g018(.din(w_G89gat_0[2]),.dout(n61),.clk(gclk));
	jand g019(.dina(w_G95gat_0[2]),.dinb(w_n61_0[1]),.dout(n62),.clk(gclk));
	jnot g020(.din(w_G1gat_0[2]),.dout(n63),.clk(gclk));
	jand g021(.dina(w_G4gat_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jor g022(.dina(n64),.dinb(n62),.dout(n65),.clk(gclk));
	jor g023(.dina(n65),.dinb(n60),.dout(n66),.clk(gclk));
	jor g024(.dina(n66),.dinb(w_dff_B_oqycvCM21_1),.dout(n67),.clk(gclk));
	jor g025(.dina(n67),.dinb(w_dff_B_psk07u3V0_1),.dout(G223gat_fa_),.clk(gclk));
	jnot g026(.din(w_G112gat_0[2]),.dout(n69),.clk(gclk));
	jnot g027(.din(w_n44_0[0]),.dout(n70),.clk(gclk));
	jnot g028(.din(w_G30gat_0[0]),.dout(n71),.clk(gclk));
	jor g029(.dina(w_n71_0[1]),.dinb(w_G24gat_0[0]),.dout(n72),.clk(gclk));
	jnot g030(.din(w_G17gat_0[1]),.dout(n73),.clk(gclk));
	jor g031(.dina(w_n73_0[1]),.dinb(w_G11gat_0[1]),.dout(n74),.clk(gclk));
	jand g032(.dina(n74),.dinb(w_n72_0[1]),.dout(n75),.clk(gclk));
	jand g033(.dina(n75),.dinb(n70),.dout(n76),.clk(gclk));
	jnot g034(.din(w_G43gat_1[0]),.dout(n77),.clk(gclk));
	jor g035(.dina(w_n77_0[1]),.dinb(w_G37gat_0[1]),.dout(n78),.clk(gclk));
	jnot g036(.din(w_G69gat_0[1]),.dout(n79),.clk(gclk));
	jor g037(.dina(w_n79_0[1]),.dinb(w_G63gat_0[1]),.dout(n80),.clk(gclk));
	jand g038(.dina(n80),.dinb(w_n78_0[1]),.dout(n81),.clk(gclk));
	jnot g039(.din(w_G108gat_0[1]),.dout(n82),.clk(gclk));
	jor g040(.dina(w_n82_0[1]),.dinb(w_G102gat_0[1]),.dout(n83),.clk(gclk));
	jnot g041(.din(w_G56gat_0[1]),.dout(n84),.clk(gclk));
	jor g042(.dina(w_n84_0[1]),.dinb(w_G50gat_0[1]),.dout(n85),.clk(gclk));
	jand g043(.dina(n85),.dinb(n83),.dout(n86),.clk(gclk));
	jnot g044(.din(w_G95gat_0[1]),.dout(n87),.clk(gclk));
	jor g045(.dina(w_n87_0[1]),.dinb(w_G89gat_0[1]),.dout(n88),.clk(gclk));
	jnot g046(.din(w_G4gat_0[1]),.dout(n89),.clk(gclk));
	jor g047(.dina(w_n89_0[1]),.dinb(w_G1gat_0[1]),.dout(n90),.clk(gclk));
	jand g048(.dina(n90),.dinb(n88),.dout(n91),.clk(gclk));
	jand g049(.dina(n91),.dinb(n86),.dout(n92),.clk(gclk));
	jand g050(.dina(n92),.dinb(w_dff_B_7jHgBMXL3_1),.dout(n93),.clk(gclk));
	jand g051(.dina(n93),.dinb(w_dff_B_1g27YgFr7_1),.dout(n94),.clk(gclk));
	jor g052(.dina(w_n94_4[1]),.dinb(w_n56_0[0]),.dout(n95),.clk(gclk));
	jand g053(.dina(n95),.dinb(w_G108gat_0[0]),.dout(n96),.clk(gclk));
	jand g054(.dina(w_n96_0[1]),.dinb(w_n69_0[1]),.dout(n97),.clk(gclk));
	jnot g055(.din(w_G8gat_0[2]),.dout(n98),.clk(gclk));
	jor g056(.dina(w_n94_4[0]),.dinb(w_n63_0[0]),.dout(n99),.clk(gclk));
	jand g057(.dina(n99),.dinb(w_G4gat_0[0]),.dout(n100),.clk(gclk));
	jand g058(.dina(w_n100_0[1]),.dinb(w_n98_0[1]),.dout(n101),.clk(gclk));
	jor g059(.dina(n101),.dinb(n97),.dout(n102),.clk(gclk));
	jnot g060(.din(w_G99gat_0[2]),.dout(n103),.clk(gclk));
	jor g061(.dina(w_n94_3[2]),.dinb(w_n61_0[0]),.dout(n104),.clk(gclk));
	jand g062(.dina(n104),.dinb(w_G95gat_0[0]),.dout(n105),.clk(gclk));
	jand g063(.dina(n105),.dinb(w_dff_B_4aXRGgFB2_1),.dout(n106),.clk(gclk));
	jnot g064(.din(w_G73gat_0[2]),.dout(n107),.clk(gclk));
	jor g065(.dina(w_n94_3[1]),.dinb(w_n53_0[0]),.dout(n108),.clk(gclk));
	jand g066(.dina(n108),.dinb(w_G69gat_0[0]),.dout(n109),.clk(gclk));
	jand g067(.dina(w_n109_0[1]),.dinb(w_n107_0[1]),.dout(n110),.clk(gclk));
	jor g068(.dina(n110),.dinb(n106),.dout(n111),.clk(gclk));
	jor g069(.dina(n111),.dinb(n102),.dout(n112),.clk(gclk));
	jxor g070(.dina(w_n94_3[0]),.dinb(w_n72_0[0]),.dout(n113),.clk(gclk));
	jor g071(.dina(n113),.dinb(w_n71_0[0]),.dout(n114),.clk(gclk));
	jor g072(.dina(w_n114_0[2]),.dinb(w_G34gat_0[2]),.dout(n115),.clk(gclk));
	jnot g073(.din(w_n115_0[1]),.dout(n116),.clk(gclk));
	jnot g074(.din(w_G60gat_0[2]),.dout(n117),.clk(gclk));
	jor g075(.dina(w_n94_2[2]),.dinb(w_n58_0[0]),.dout(n118),.clk(gclk));
	jand g076(.dina(n118),.dinb(w_G56gat_0[0]),.dout(n119),.clk(gclk));
	jand g077(.dina(w_n119_0[1]),.dinb(w_dff_B_u6r39nYs8_1),.dout(n120),.clk(gclk));
	jxor g078(.dina(w_n94_2[1]),.dinb(w_n52_0[0]),.dout(n121),.clk(gclk));
	jnot g079(.din(w_G47gat_0[1]),.dout(n122),.clk(gclk));
	jand g080(.dina(n122),.dinb(w_G43gat_0[2]),.dout(n123),.clk(gclk));
	jand g081(.dina(w_n123_0[1]),.dinb(w_n121_0[1]),.dout(n124),.clk(gclk));
	jor g082(.dina(w_dff_B_rsRN4gi21_0),.dinb(n120),.dout(n125),.clk(gclk));
	jnot g083(.din(w_G86gat_1[1]),.dout(n126),.clk(gclk));
	jor g084(.dina(w_n94_2[0]),.dinb(w_n43_0[0]),.dout(n127),.clk(gclk));
	jand g085(.dina(n127),.dinb(w_G82gat_0[1]),.dout(n128),.clk(gclk));
	jand g086(.dina(w_n128_0[1]),.dinb(w_n126_0[2]),.dout(n129),.clk(gclk));
	jnot g087(.din(w_G21gat_1[1]),.dout(n130),.clk(gclk));
	jor g088(.dina(w_n94_1[2]),.dinb(w_n47_0[0]),.dout(n131),.clk(gclk));
	jand g089(.dina(n131),.dinb(w_G17gat_0[0]),.dout(n132),.clk(gclk));
	jand g090(.dina(w_n132_0[1]),.dinb(w_n130_0[2]),.dout(n133),.clk(gclk));
	jor g091(.dina(n133),.dinb(n129),.dout(n134),.clk(gclk));
	jor g092(.dina(n134),.dinb(n125),.dout(n135),.clk(gclk));
	jor g093(.dina(n135),.dinb(w_dff_B_5HVIxTto7_1),.dout(n136),.clk(gclk));
	jor g094(.dina(n136),.dinb(w_dff_B_L8xAIm631_1),.dout(G329gat_fa_),.clk(gclk));
	jand g095(.dina(w_G223gat_3[1]),.dinb(w_G89gat_0[0]),.dout(n138),.clk(gclk));
	jor g096(.dina(n138),.dinb(w_n87_0[0]),.dout(n139),.clk(gclk));
	jand g097(.dina(w_G329gat_6),.dinb(w_G99gat_0[1]),.dout(n140),.clk(gclk));
	jor g098(.dina(n140),.dinb(w_n139_0[1]),.dout(n141),.clk(gclk));
	jor g099(.dina(w_n141_0[1]),.dinb(w_G105gat_0[1]),.dout(n142),.clk(gclk));
	jnot g100(.din(w_n142_0[1]),.dout(n143),.clk(gclk));
	jand g101(.dina(w_G223gat_3[0]),.dinb(w_G50gat_0[0]),.dout(n144),.clk(gclk));
	jor g102(.dina(n144),.dinb(w_n84_0[0]),.dout(n145),.clk(gclk));
	jor g103(.dina(w_n145_0[1]),.dinb(w_G60gat_0[1]),.dout(n146),.clk(gclk));
	jand g104(.dina(w_G329gat_5[2]),.dinb(w_n146_0[1]),.dout(n147),.clk(gclk));
	jnot g105(.din(w_n147_0[1]),.dout(n148),.clk(gclk));
	jnot g106(.din(w_G66gat_0[1]),.dout(n150),.clk(gclk));
	jand g107(.dina(w_n119_0[0]),.dinb(w_n150_0[1]),.dout(n151),.clk(gclk));
	jand g108(.dina(w_n151_0[1]),.dinb(n148),.dout(n153),.clk(gclk));
	jnot g109(.din(w_G79gat_0[1]),.dout(n154),.clk(gclk));
	jand g110(.dina(w_G223gat_2[2]),.dinb(w_G102gat_0[0]),.dout(n155),.clk(gclk));
	jor g111(.dina(n155),.dinb(w_n82_0[0]),.dout(n156),.clk(gclk));
	jor g112(.dina(w_n156_0[1]),.dinb(w_G112gat_0[1]),.dout(n157),.clk(gclk));
	jand g113(.dina(w_G223gat_2[1]),.dinb(w_G1gat_0[0]),.dout(n158),.clk(gclk));
	jor g114(.dina(n158),.dinb(w_n89_0[0]),.dout(n159),.clk(gclk));
	jor g115(.dina(w_n159_0[1]),.dinb(w_G8gat_0[1]),.dout(n160),.clk(gclk));
	jand g116(.dina(n160),.dinb(n157),.dout(n161),.clk(gclk));
	jor g117(.dina(w_n139_0[0]),.dinb(w_G99gat_0[0]),.dout(n162),.clk(gclk));
	jand g118(.dina(w_G223gat_2[0]),.dinb(w_G63gat_0[0]),.dout(n163),.clk(gclk));
	jor g119(.dina(n163),.dinb(w_n79_0[0]),.dout(n164),.clk(gclk));
	jor g120(.dina(w_n164_0[1]),.dinb(w_G73gat_0[1]),.dout(n165),.clk(gclk));
	jand g121(.dina(n165),.dinb(n162),.dout(n166),.clk(gclk));
	jand g122(.dina(n166),.dinb(n161),.dout(n167),.clk(gclk));
	jxor g123(.dina(w_n94_1[1]),.dinb(w_n78_0[0]),.dout(n168),.clk(gclk));
	jnot g124(.din(w_n123_0[0]),.dout(n169),.clk(gclk));
	jor g125(.dina(w_dff_B_i8ozyrsk5_0),.dinb(n168),.dout(n170),.clk(gclk));
	jand g126(.dina(w_n170_0[1]),.dinb(w_n146_0[0]),.dout(n171),.clk(gclk));
	jnot g127(.din(w_G82gat_0[0]),.dout(n172),.clk(gclk));
	jand g128(.dina(w_G223gat_1[2]),.dinb(w_G76gat_0[0]),.dout(n173),.clk(gclk));
	jor g129(.dina(n173),.dinb(w_dff_B_vuzsV2FC6_1),.dout(n174),.clk(gclk));
	jor g130(.dina(w_n174_0[1]),.dinb(w_G86gat_1[0]),.dout(n175),.clk(gclk));
	jand g131(.dina(w_G223gat_1[1]),.dinb(w_G11gat_0[0]),.dout(n176),.clk(gclk));
	jor g132(.dina(n176),.dinb(w_n73_0[0]),.dout(n177),.clk(gclk));
	jor g133(.dina(w_n177_0[1]),.dinb(w_G21gat_1[0]),.dout(n178),.clk(gclk));
	jand g134(.dina(n178),.dinb(n175),.dout(n179),.clk(gclk));
	jand g135(.dina(n179),.dinb(n171),.dout(n180),.clk(gclk));
	jand g136(.dina(n180),.dinb(w_n115_0[0]),.dout(n181),.clk(gclk));
	jand g137(.dina(n181),.dinb(w_dff_B_TULCKkIv7_1),.dout(n182),.clk(gclk));
	jor g138(.dina(w_n182_3[1]),.dinb(w_n107_0[0]),.dout(n183),.clk(gclk));
	jand g139(.dina(n183),.dinb(w_n109_0[0]),.dout(n184),.clk(gclk));
	jand g140(.dina(w_n184_0[1]),.dinb(w_n154_0[1]),.dout(n185),.clk(gclk));
	jor g141(.dina(n185),.dinb(n153),.dout(n186),.clk(gclk));
	jor g142(.dina(n186),.dinb(n143),.dout(n187),.clk(gclk));
	jand g143(.dina(w_G329gat_5[1]),.dinb(w_n170_0[0]),.dout(n188),.clk(gclk));
	jnot g144(.din(w_n188_0[1]),.dout(n189),.clk(gclk));
	jnot g145(.din(w_G53gat_0[1]),.dout(n191),.clk(gclk));
	jand g146(.dina(w_n191_0[1]),.dinb(w_G43gat_0[1]),.dout(n192),.clk(gclk));
	jand g147(.dina(w_dff_B_0xlbnkxf7_0),.dinb(w_n121_0[0]),.dout(n193),.clk(gclk));
	jand g148(.dina(w_n193_0[1]),.dinb(n189),.dout(n195),.clk(gclk));
	jor g149(.dina(w_n182_3[0]),.dinb(w_n130_0[1]),.dout(n196),.clk(gclk));
	jand g150(.dina(n196),.dinb(w_n132_0[0]),.dout(n197),.clk(gclk));
	jnot g151(.din(w_G27gat_0[1]),.dout(n198),.clk(gclk));
	jor g152(.dina(w_G329gat_5[0]),.dinb(w_G21gat_0[2]),.dout(n199),.clk(gclk));
	jand g153(.dina(n199),.dinb(w_n198_0[1]),.dout(n200),.clk(gclk));
	jand g154(.dina(n200),.dinb(w_n197_0[1]),.dout(n201),.clk(gclk));
	jor g155(.dina(n201),.dinb(n195),.dout(n202),.clk(gclk));
	jor g156(.dina(w_n182_2[2]),.dinb(w_n126_0[1]),.dout(n203),.clk(gclk));
	jand g157(.dina(n203),.dinb(w_n128_0[0]),.dout(n204),.clk(gclk));
	jnot g158(.din(w_G92gat_0[2]),.dout(n205),.clk(gclk));
	jor g159(.dina(w_G329gat_4[2]),.dinb(w_G86gat_0[2]),.dout(n206),.clk(gclk));
	jand g160(.dina(n206),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jand g161(.dina(n207),.dinb(w_n204_0[1]),.dout(n208),.clk(gclk));
	jnot g162(.din(w_G14gat_0[2]),.dout(n209),.clk(gclk));
	jor g163(.dina(w_n182_2[1]),.dinb(w_n98_0[0]),.dout(n210),.clk(gclk));
	jand g164(.dina(n210),.dinb(w_n100_0[0]),.dout(n211),.clk(gclk));
	jand g165(.dina(n211),.dinb(w_dff_B_dpOwkNU81_1),.dout(n212),.clk(gclk));
	jor g166(.dina(n212),.dinb(n208),.dout(n213),.clk(gclk));
	jnot g167(.din(w_G34gat_0[1]),.dout(n214),.clk(gclk));
	jor g168(.dina(w_n182_2[0]),.dinb(w_dff_B_o98iBe3S6_1),.dout(n215),.clk(gclk));
	jnot g169(.din(w_G40gat_0[1]),.dout(n217),.clk(gclk));
	jnot g170(.din(w_n114_0[1]),.dout(n218),.clk(gclk));
	jand g171(.dina(n218),.dinb(w_n217_0[1]),.dout(n219),.clk(gclk));
	jand g172(.dina(w_n219_0[1]),.dinb(n215),.dout(n221),.clk(gclk));
	jnot g173(.din(w_G115gat_0[1]),.dout(n222),.clk(gclk));
	jor g174(.dina(w_n182_1[2]),.dinb(w_n69_0[0]),.dout(n223),.clk(gclk));
	jand g175(.dina(n223),.dinb(w_n96_0[0]),.dout(n224),.clk(gclk));
	jand g176(.dina(w_n224_0[1]),.dinb(w_n222_0[1]),.dout(n225),.clk(gclk));
	jor g177(.dina(n225),.dinb(w_dff_B_WWvHWYd57_1),.dout(n226),.clk(gclk));
	jor g178(.dina(n226),.dinb(n213),.dout(n227),.clk(gclk));
	jor g179(.dina(n227),.dinb(w_dff_B_0pCmD9204_1),.dout(n228),.clk(gclk));
	jor g180(.dina(n228),.dinb(w_dff_B_moVH5SBR5_1),.dout(G370gat_fa_),.clk(gclk));
	jand g181(.dina(w_G329gat_4[1]),.dinb(w_G8gat_0[0]),.dout(n230),.clk(gclk));
	jor g182(.dina(n230),.dinb(w_n159_0[0]),.dout(n231),.clk(gclk));
	jand g183(.dina(w_G370gat_2),.dinb(w_G14gat_0[1]),.dout(n232),.clk(gclk));
	jor g184(.dina(n232),.dinb(w_n231_0[1]),.dout(n233),.clk(gclk));
	jnot g185(.din(w_n151_0[0]),.dout(n235),.clk(gclk));
	jor g186(.dina(w_dff_B_iR4wkDcl9_0),.dinb(w_n147_0[0]),.dout(n237),.clk(gclk));
	jand g187(.dina(w_G329gat_4[0]),.dinb(w_G73gat_0[0]),.dout(n238),.clk(gclk));
	jor g188(.dina(n238),.dinb(w_n164_0[0]),.dout(n239),.clk(gclk));
	jor g189(.dina(n239),.dinb(w_G79gat_0[0]),.dout(n240),.clk(gclk));
	jand g190(.dina(n240),.dinb(w_dff_B_a1rqcxTg0_1),.dout(n241),.clk(gclk));
	jand g191(.dina(n241),.dinb(w_n142_0[0]),.dout(n242),.clk(gclk));
	jnot g192(.din(w_n193_0[0]),.dout(n244),.clk(gclk));
	jor g193(.dina(w_dff_B_sJNE8zIO8_0),.dinb(w_n188_0[0]),.dout(n246),.clk(gclk));
	jand g194(.dina(w_G329gat_3[2]),.dinb(w_G21gat_0[1]),.dout(n247),.clk(gclk));
	jor g195(.dina(n247),.dinb(w_n177_0[0]),.dout(n248),.clk(gclk));
	jand g196(.dina(w_n182_1[1]),.dinb(w_n130_0[0]),.dout(n249),.clk(gclk));
	jor g197(.dina(n249),.dinb(w_G27gat_0[0]),.dout(n250),.clk(gclk));
	jor g198(.dina(n250),.dinb(n248),.dout(n251),.clk(gclk));
	jand g199(.dina(n251),.dinb(w_dff_B_Vhe6vJ0b1_1),.dout(n252),.clk(gclk));
	jand g200(.dina(w_G329gat_3[1]),.dinb(w_G86gat_0[1]),.dout(n253),.clk(gclk));
	jor g201(.dina(n253),.dinb(w_n174_0[0]),.dout(n254),.clk(gclk));
	jand g202(.dina(w_n182_1[0]),.dinb(w_n126_0[0]),.dout(n255),.clk(gclk));
	jor g203(.dina(n255),.dinb(w_G92gat_0[1]),.dout(n256),.clk(gclk));
	jor g204(.dina(n256),.dinb(w_n254_0[1]),.dout(n257),.clk(gclk));
	jor g205(.dina(w_n231_0[0]),.dinb(w_G14gat_0[0]),.dout(n258),.clk(gclk));
	jand g206(.dina(n258),.dinb(n257),.dout(n259),.clk(gclk));
	jand g207(.dina(w_G329gat_3[0]),.dinb(w_G34gat_0[0]),.dout(n260),.clk(gclk));
	jnot g208(.din(w_n219_0[0]),.dout(n262),.clk(gclk));
	jor g209(.dina(w_dff_B_Gh5mMvPZ6_0),.dinb(w_n260_0[1]),.dout(n264),.clk(gclk));
	jand g210(.dina(w_G329gat_2[2]),.dinb(w_G112gat_0[0]),.dout(n265),.clk(gclk));
	jor g211(.dina(n265),.dinb(w_n156_0[0]),.dout(n266),.clk(gclk));
	jor g212(.dina(n266),.dinb(w_G115gat_0[0]),.dout(n267),.clk(gclk));
	jand g213(.dina(n267),.dinb(w_dff_B_eADzKhT00_1),.dout(n268),.clk(gclk));
	jand g214(.dina(n268),.dinb(n259),.dout(n269),.clk(gclk));
	jand g215(.dina(n269),.dinb(w_dff_B_RwErxWos9_1),.dout(n270),.clk(gclk));
	jand g216(.dina(n270),.dinb(w_dff_B_erZJyVKo4_1),.dout(n271),.clk(gclk));
	jor g217(.dina(w_n271_3[1]),.dinb(w_n150_0[0]),.dout(n272),.clk(gclk));
	jand g218(.dina(w_G329gat_2[1]),.dinb(w_G60gat_0[0]),.dout(n273),.clk(gclk));
	jor g219(.dina(n273),.dinb(w_n145_0[0]),.dout(n274),.clk(gclk));
	jnot g220(.din(w_n274_0[1]),.dout(n275),.clk(gclk));
	jand g221(.dina(w_dff_B_2aQgTpKd8_0),.dinb(n272),.dout(n276),.clk(gclk));
	jor g222(.dina(w_n271_3[0]),.dinb(w_n191_0[0]),.dout(n277),.clk(gclk));
	jand g223(.dina(w_G329gat_2[0]),.dinb(w_G47gat_0[0]),.dout(n278),.clk(gclk));
	jand g224(.dina(w_G223gat_1[0]),.dinb(w_G37gat_0[0]),.dout(n279),.clk(gclk));
	jor g225(.dina(n279),.dinb(w_n77_0[0]),.dout(n280),.clk(gclk));
	jor g226(.dina(w_dff_B_uXF6yqlK1_0),.dinb(n278),.dout(n281),.clk(gclk));
	jnot g227(.din(w_n281_0[1]),.dout(n282),.clk(gclk));
	jand g228(.dina(w_dff_B_DkoggYqW3_0),.dinb(n277),.dout(n283),.clk(gclk));
	jor g229(.dina(w_n283_0[1]),.dinb(n276),.dout(n284),.clk(gclk));
	jor g230(.dina(w_n271_2[2]),.dinb(w_n198_0[0]),.dout(n285),.clk(gclk));
	jand g231(.dina(n285),.dinb(w_n197_0[0]),.dout(n286),.clk(gclk));
	jor g232(.dina(w_n271_2[1]),.dinb(w_n217_0[0]),.dout(n287),.clk(gclk));
	jor g233(.dina(w_n114_0[0]),.dinb(w_n260_0[0]),.dout(n290),.clk(gclk));
	jnot g234(.din(w_n290_0[1]),.dout(n291),.clk(gclk));
	jand g235(.dina(w_dff_B_TNL17A3L5_0),.dinb(n287),.dout(n292),.clk(gclk));
	jor g236(.dina(n292),.dinb(w_n286_0[1]),.dout(n293),.clk(gclk));
	jor g237(.dina(w_n293_0[1]),.dinb(n284),.dout(G430gat_fa_),.clk(gclk));
	jor g238(.dina(w_n271_2[0]),.dinb(w_n205_0[0]),.dout(n295),.clk(gclk));
	jand g239(.dina(n295),.dinb(w_n204_0[0]),.dout(n296),.clk(gclk));
	jor g240(.dina(w_n271_1[2]),.dinb(w_n222_0[0]),.dout(n297),.clk(gclk));
	jand g241(.dina(n297),.dinb(w_n224_0[0]),.dout(n298),.clk(gclk));
	jor g242(.dina(n298),.dinb(w_n296_0[1]),.dout(n299),.clk(gclk));
	jnot g243(.din(w_n141_0[0]),.dout(n300),.clk(gclk));
	jnot g244(.din(w_G105gat_0[0]),.dout(n301),.clk(gclk));
	jor g245(.dina(w_n271_1[1]),.dinb(w_dff_B_jfxZeJNT7_1),.dout(n302),.clk(gclk));
	jand g246(.dina(n302),.dinb(w_dff_B_IOwF4Glq7_1),.dout(n303),.clk(gclk));
	jor g247(.dina(w_n271_1[0]),.dinb(w_n154_0[0]),.dout(n304),.clk(gclk));
	jand g248(.dina(n304),.dinb(w_n184_0[0]),.dout(n305),.clk(gclk));
	jor g249(.dina(w_n305_0[1]),.dinb(w_n303_0[1]),.dout(n306),.clk(gclk));
	jor g250(.dina(n306),.dinb(n299),.dout(n307),.clk(gclk));
	jor g251(.dina(n307),.dinb(w_G430gat_0),.dout(n308),.clk(gclk));
	jand g252(.dina(n308),.dinb(w_dff_B_TBCYFE2o0_1),.dout(G421gat),.clk(gclk));
	jand g253(.dina(w_G370gat_1[2]),.dinb(w_G66gat_0[0]),.dout(n310),.clk(gclk));
	jor g254(.dina(w_n274_0[0]),.dinb(n310),.dout(n311),.clk(gclk));
	jand g255(.dina(w_G370gat_1[1]),.dinb(w_G53gat_0[0]),.dout(n312),.clk(gclk));
	jor g256(.dina(w_n281_0[0]),.dinb(n312),.dout(n313),.clk(gclk));
	jand g257(.dina(w_n313_0[1]),.dinb(n311),.dout(n314),.clk(gclk));
	jand g258(.dina(w_n296_0[0]),.dinb(w_n314_0[1]),.dout(n315),.clk(gclk));
	jand g259(.dina(w_G370gat_1[0]),.dinb(w_G40gat_0[0]),.dout(n316),.clk(gclk));
	jor g260(.dina(w_n290_0[0]),.dinb(n316),.dout(n317),.clk(gclk));
	jand g261(.dina(w_n305_0[0]),.dinb(w_n317_0[2]),.dout(n318),.clk(gclk));
	jand g262(.dina(n318),.dinb(w_n314_0[0]),.dout(n319),.clk(gclk));
	jor g263(.dina(w_n319_0[1]),.dinb(w_n293_0[0]),.dout(n320),.clk(gclk));
	jor g264(.dina(n320),.dinb(w_dff_B_zqiK0Xpw6_1),.dout(G431gat),.clk(gclk));
	jand g265(.dina(w_G370gat_0[2]),.dinb(w_G92gat_0[0]),.dout(n322),.clk(gclk));
	jor g266(.dina(n322),.dinb(w_n254_0[0]),.dout(n323),.clk(gclk));
	jand g267(.dina(n323),.dinb(w_n313_0[0]),.dout(n324),.clk(gclk));
	jand g268(.dina(w_n303_0[0]),.dinb(w_n317_0[1]),.dout(n325),.clk(gclk));
	jand g269(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jand g270(.dina(w_n317_0[0]),.dinb(w_n283_0[0]),.dout(n327),.clk(gclk));
	jor g271(.dina(n327),.dinb(w_n286_0[0]),.dout(n328),.clk(gclk));
	jor g272(.dina(n328),.dinb(w_n319_0[0]),.dout(n329),.clk(gclk));
	jor g273(.dina(n329),.dinb(w_dff_B_RIYvRidS5_1),.dout(G432gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_qMJdKDQo4_0),.doutb(w_dff_A_A24A1gXq5_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_dff_A_B0KcFS5N3_0),.doutb(w_G4gat_0[1]),.doutc(w_dff_A_OXR4KdRt3_2),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_BF8gCdAp4_0),.doutb(w_dff_A_6l4mxBtJ8_1),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G11gat_0(.douta(w_dff_A_MQd5T3JC6_0),.doutb(w_dff_A_scHdCel47_1),.doutc(w_G11gat_0[2]),.din(G11gat));
	jspl3 jspl3_w_G14gat_0(.douta(w_dff_A_X0N0VDcb5_0),.doutb(w_dff_A_reYrKxhI4_1),.doutc(w_G14gat_0[2]),.din(G14gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_dff_A_xXeOIwou4_0),.doutb(w_G17gat_0[1]),.doutc(w_dff_A_eny0RcZF5_2),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_G21gat_0[0]),.doutb(w_dff_A_ylkeI8A80_1),.doutc(w_dff_A_8CzVoGhG7_2),.din(G21gat));
	jspl jspl_w_G21gat_1(.douta(w_dff_A_6wYury1T2_0),.doutb(w_G21gat_1[1]),.din(w_G21gat_0[0]));
	jspl jspl_w_G24gat_0(.douta(w_dff_A_8fNpvyNO4_0),.doutb(w_G24gat_0[1]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_dff_A_O0PhjXJJ1_0),.doutb(w_G27gat_0[1]),.din(G27gat));
	jspl jspl_w_G30gat_0(.douta(w_G30gat_0[0]),.doutb(w_dff_A_vq767C681_1),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_dff_A_kTjO4ryG8_0),.doutb(w_G34gat_0[1]),.doutc(w_dff_A_HLRxu9hC8_2),.din(G34gat));
	jspl3 jspl3_w_G37gat_0(.douta(w_dff_A_N4JjRjiX8_0),.doutb(w_dff_A_iK9sgUV75_1),.doutc(w_G37gat_0[2]),.din(G37gat));
	jspl jspl_w_G40gat_0(.douta(w_dff_A_diYIX76x0_0),.doutb(w_G40gat_0[1]),.din(G40gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_G43gat_0[0]),.doutb(w_dff_A_xghP78uJ2_1),.doutc(w_dff_A_Pjmk4a686_2),.din(G43gat));
	jspl jspl_w_G43gat_1(.douta(w_G43gat_1[0]),.doutb(w_dff_A_wAnMmerE8_1),.din(w_G43gat_0[0]));
	jspl jspl_w_G47gat_0(.douta(w_dff_A_7wffRQjy9_0),.doutb(w_G47gat_0[1]),.din(G47gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_dff_A_XquBIlvv5_0),.doutb(w_dff_A_o0bLKkPz9_1),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_dff_A_OYC4wMHD3_0),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_dff_A_MpS27uXT9_0),.doutb(w_G56gat_0[1]),.doutc(w_dff_A_LTw6E6Ql5_2),.din(G56gat));
	jspl3 jspl3_w_G60gat_0(.douta(w_dff_A_tKksQxqR6_0),.doutb(w_dff_A_gtyfAx5u2_1),.doutc(w_G60gat_0[2]),.din(G60gat));
	jspl3 jspl3_w_G63gat_0(.douta(w_dff_A_HZbKt9s03_0),.doutb(w_dff_A_U0O983TN1_1),.doutc(w_G63gat_0[2]),.din(G63gat));
	jspl jspl_w_G66gat_0(.douta(w_dff_A_4L7SPVuI9_0),.doutb(w_G66gat_0[1]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_dff_A_Ge8B9hJt4_0),.doutb(w_G69gat_0[1]),.doutc(w_dff_A_4g578riZ3_2),.din(G69gat));
	jspl3 jspl3_w_G73gat_0(.douta(w_dff_A_Uf4wyVZi1_0),.doutb(w_dff_A_LFlt7WTf2_1),.doutc(w_G73gat_0[2]),.din(G73gat));
	jspl jspl_w_G76gat_0(.douta(w_dff_A_Z8LXqTPZ1_0),.doutb(w_G76gat_0[1]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_dff_A_IcPR62ao3_0),.doutb(w_G79gat_0[1]),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_G82gat_0[0]),.doutb(w_dff_A_7hgsGo9G1_1),.doutc(w_dff_A_iYOw4pOk9_2),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_dff_A_3RY14p7Q2_1),.doutc(w_dff_A_kTePh0YY1_2),.din(G86gat));
	jspl jspl_w_G86gat_1(.douta(w_dff_A_zpvm1eo74_0),.doutb(w_G86gat_1[1]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G89gat_0(.douta(w_dff_A_VTHH7CAn5_0),.doutb(w_dff_A_wx4vqfXc1_1),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_hTvL5vzG1_0),.doutb(w_dff_A_Cja6zkSj7_1),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_dff_A_F2J5LdON6_0),.doutb(w_G95gat_0[1]),.doutc(w_dff_A_AcISA6RU7_2),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_4MmouBb57_0),.doutb(w_dff_A_3q3Udb6f2_1),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl3 jspl3_w_G102gat_0(.douta(w_dff_A_VjTQ0GMX3_0),.doutb(w_dff_A_uTzSJXu04_1),.doutc(w_G102gat_0[2]),.din(G102gat));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_dff_A_PYJI8UMC6_1),.din(G105gat));
	jspl3 jspl3_w_G108gat_0(.douta(w_dff_A_Z5ttAmgn2_0),.doutb(w_G108gat_0[1]),.doutc(w_dff_A_WgCxUncS6_2),.din(G108gat));
	jspl3 jspl3_w_G112gat_0(.douta(w_dff_A_y0ynk3B09_0),.doutb(w_dff_A_nAPqZLqT6_1),.doutc(w_G112gat_0[2]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_dff_A_AvwkGZtH5_0),.doutb(w_G115gat_0[1]),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(w_dff_A_MaxiYCp89_2),.din(w_G223gat_0[2]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl3 jspl3_w_G329gat_4(.douta(w_G329gat_4[0]),.doutb(w_G329gat_4[1]),.doutc(w_G329gat_4[2]),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G329gat_5(.douta(w_G329gat_5[0]),.doutb(w_G329gat_5[1]),.doutc(w_G329gat_5[2]),.din(w_G329gat_1[1]));
	jspl jspl_w_G329gat_6(.douta(w_G329gat_6),.doutb(w_dff_A_R3l9X8Gn8_1),.din(w_G329gat_1[2]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_G370gat_1[2]),.din(w_G370gat_0[0]));
	jspl jspl_w_G370gat_2(.douta(w_G370gat_2),.doutb(w_dff_A_cgYnHa567_1),.din(w_G370gat_0[1]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(w_dff_A_RCUy6P1j0_1),.din(G430gat_fa_));
	jspl jspl_w_n43_0(.douta(w_dff_A_1S6iYLtK3_0),.doutb(w_n43_0[1]),.din(n43));
	jspl jspl_w_n44_0(.douta(w_n44_0[0]),.doutb(w_dff_A_DMrYvpqC1_1),.din(n44));
	jspl jspl_w_n47_0(.douta(w_dff_A_jrm4zwtG2_0),.doutb(w_n47_0[1]),.din(n47));
	jspl jspl_w_n52_0(.douta(w_dff_A_3ykacEbC4_0),.doutb(w_n52_0[1]),.din(n52));
	jspl jspl_w_n53_0(.douta(w_dff_A_QQxypFdR7_0),.doutb(w_n53_0[1]),.din(n53));
	jspl jspl_w_n56_0(.douta(w_dff_A_UoMNT9Qa5_0),.doutb(w_n56_0[1]),.din(n56));
	jspl jspl_w_n58_0(.douta(w_dff_A_bmwWrFaJ6_0),.doutb(w_n58_0[1]),.din(n58));
	jspl jspl_w_n61_0(.douta(w_dff_A_0ee1nJSj0_0),.doutb(w_n61_0[1]),.din(n61));
	jspl jspl_w_n63_0(.douta(w_dff_A_GHmMaPQz1_0),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n69_0(.douta(w_dff_A_9tiFhrMz9_0),.doutb(w_n69_0[1]),.din(w_dff_B_R69DaiPJ4_2));
	jspl jspl_w_n71_0(.douta(w_dff_A_im35mc7u0_0),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n72_0(.douta(w_dff_A_mjNe2c9q6_0),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n73_0(.douta(w_dff_A_p5hPemGS8_0),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n77_0(.douta(w_dff_A_DQdR1sTx9_0),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_dff_A_3oa89vUu6_0),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n79_0(.douta(w_dff_A_0iX5VOvF3_0),.doutb(w_n79_0[1]),.din(n79));
	jspl jspl_w_n82_0(.douta(w_dff_A_PftCV0974_0),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_dff_A_t6pyZeN27_0),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n87_0(.douta(w_dff_A_st7JVpjz6_0),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_dff_A_vcoSxdJH7_0),.doutb(w_n89_0[1]),.din(n89));
	jspl3 jspl3_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl3 jspl3_w_n94_1(.douta(w_n94_1[0]),.doutb(w_n94_1[1]),.doutc(w_n94_1[2]),.din(w_n94_0[0]));
	jspl3 jspl3_w_n94_2(.douta(w_n94_2[0]),.doutb(w_n94_2[1]),.doutc(w_n94_2[2]),.din(w_n94_0[1]));
	jspl3 jspl3_w_n94_3(.douta(w_n94_3[0]),.doutb(w_n94_3[1]),.doutc(w_n94_3[2]),.din(w_n94_0[2]));
	jspl jspl_w_n94_4(.douta(w_n94_4[0]),.doutb(w_n94_4[1]),.din(w_n94_1[0]));
	jspl jspl_w_n96_0(.douta(w_dff_A_F1VAy6oj4_0),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_dff_A_QQALszhd2_0),.doutb(w_n98_0[1]),.din(w_dff_B_zzOnSQo75_2));
	jspl jspl_w_n100_0(.douta(w_dff_A_FycskBfx6_0),.doutb(w_n100_0[1]),.din(n100));
	jspl jspl_w_n107_0(.douta(w_dff_A_Klo8Z9nq0_0),.doutb(w_n107_0[1]),.din(w_dff_B_Qpnbjv8i6_2));
	jspl jspl_w_n109_0(.douta(w_dff_A_riHUICMo6_0),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n114_0(.douta(w_dff_A_2iAQPlyp8_0),.doutb(w_n114_0[1]),.doutc(w_n114_0[2]),.din(n114));
	jspl jspl_w_n115_0(.douta(w_dff_A_8PsZVu7s4_0),.doutb(w_n115_0[1]),.din(n115));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n123_0(.douta(w_n123_0[0]),.doutb(w_dff_A_0GVK19w73_1),.din(n123));
	jspl3 jspl3_w_n126_0(.douta(w_dff_A_QLBicpOR7_0),.doutb(w_dff_A_u7RDWOiz3_1),.doutc(w_n126_0[2]),.din(w_dff_B_SWO0A4BS1_3));
	jspl jspl_w_n128_0(.douta(w_dff_A_nFqf8QzF1_0),.doutb(w_n128_0[1]),.din(n128));
	jspl3 jspl3_w_n130_0(.douta(w_dff_A_ikW0gD047_0),.doutb(w_dff_A_Ss3t7B913_1),.doutc(w_n130_0[2]),.din(w_dff_B_duBsfNaE5_3));
	jspl jspl_w_n132_0(.douta(w_dff_A_HxjKhfpm3_0),.doutb(w_n132_0[1]),.din(n132));
	jspl jspl_w_n139_0(.douta(w_n139_0[0]),.doutb(w_dff_A_8uzRIjdi1_1),.din(n139));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_dff_A_TH3VM6Wq8_0),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n145_0(.douta(w_dff_A_jggaCk2R5_0),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_YDMdgSf06_1),.din(n146));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl jspl_w_n150_0(.douta(w_dff_A_b787DLJQ7_0),.doutb(w_n150_0[1]),.din(w_dff_B_oJ0khUTh6_2));
	jspl jspl_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_iswuUbvY4_1),.din(n151));
	jspl jspl_w_n154_0(.douta(w_dff_A_nl7IyFXG9_0),.doutb(w_n154_0[1]),.din(w_dff_B_ynVHqGdP0_2));
	jspl jspl_w_n156_0(.douta(w_dff_A_ZOGdPGs42_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n159_0(.douta(w_dff_A_3fWF9Vay3_0),.doutb(w_n159_0[1]),.din(n159));
	jspl jspl_w_n164_0(.douta(w_dff_A_P8mWUwpS3_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n170_0(.douta(w_dff_A_I0B4DkU05_0),.doutb(w_n170_0[1]),.din(w_dff_B_DacFIcBk5_2));
	jspl jspl_w_n174_0(.douta(w_dff_A_1NHobVf29_0),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n177_0(.douta(w_dff_A_eV97XeUj9_0),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n182_2(.douta(w_n182_2[0]),.doutb(w_n182_2[1]),.doutc(w_n182_2[2]),.din(w_n182_0[1]));
	jspl jspl_w_n182_3(.douta(w_n182_3[0]),.doutb(w_n182_3[1]),.din(w_n182_0[2]));
	jspl jspl_w_n184_0(.douta(w_dff_A_ajlO7iq04_0),.doutb(w_n184_0[1]),.din(n184));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n191_0(.douta(w_dff_A_NztlICNx4_0),.doutb(w_n191_0[1]),.din(n191));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_dff_A_s6t7iNYI6_1),.din(n193));
	jspl jspl_w_n197_0(.douta(w_dff_A_T30xqLpp4_0),.doutb(w_n197_0[1]),.din(n197));
	jspl jspl_w_n198_0(.douta(w_dff_A_0CyklLM18_0),.doutb(w_n198_0[1]),.din(w_dff_B_fyrZXCvG0_2));
	jspl jspl_w_n204_0(.douta(w_dff_A_kJY4IHWD0_0),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n205_0(.douta(w_dff_A_mutchN9n9_0),.doutb(w_n205_0[1]),.din(w_dff_B_uUvTNaPX9_2));
	jspl jspl_w_n217_0(.douta(w_dff_A_zSHVQ4E95_0),.doutb(w_n217_0[1]),.din(w_dff_B_fgU23e0C8_2));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_dff_A_LmDCxI092_1),.din(n219));
	jspl jspl_w_n222_0(.douta(w_dff_A_UrpyTP039_0),.doutb(w_n222_0[1]),.din(w_dff_B_gbWZni8G5_2));
	jspl jspl_w_n224_0(.douta(w_dff_A_6c6mhX8v0_0),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_dff_A_ZkBAqm027_1),.din(n231));
	jspl jspl_w_n254_0(.douta(w_dff_A_kM1VUIek2_0),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_n271_1[0]),.doutb(w_n271_1[1]),.doutc(w_n271_1[2]),.din(w_n271_0[0]));
	jspl3 jspl3_w_n271_2(.douta(w_n271_2[0]),.doutb(w_n271_2[1]),.doutc(w_n271_2[2]),.din(w_n271_0[1]));
	jspl jspl_w_n271_3(.douta(w_n271_3[0]),.doutb(w_n271_3[1]),.din(w_n271_0[2]));
	jspl jspl_w_n274_0(.douta(w_dff_A_ww5EVM0P1_0),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n281_0(.douta(w_dff_A_tVDtwLTa1_0),.doutb(w_n281_0[1]),.din(n281));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.din(n283));
	jspl jspl_w_n286_0(.douta(w_dff_A_lUbJeBKw1_0),.doutb(w_n286_0[1]),.din(n286));
	jspl jspl_w_n290_0(.douta(w_dff_A_GzvYsrTd6_0),.doutb(w_n290_0[1]),.din(n290));
	jspl jspl_w_n293_0(.douta(w_dff_A_ap4p4pgH8_0),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n296_0(.douta(w_dff_A_bhTq7Q2L7_0),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(n305));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.din(n314));
	jspl3 jspl3_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.doutc(w_n317_0[2]),.din(n317));
	jspl jspl_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.din(n319));
	jdff dff_B_95uf8pzk0_1(.din(n233),.dout(w_dff_B_95uf8pzk0_1),.clk(gclk));
	jdff dff_B_letGXm1p6_1(.din(w_dff_B_95uf8pzk0_1),.dout(w_dff_B_letGXm1p6_1),.clk(gclk));
	jdff dff_B_TBCYFE2o0_1(.din(w_dff_B_letGXm1p6_1),.dout(w_dff_B_TBCYFE2o0_1),.clk(gclk));
	jdff dff_B_pTm7TwKv4_0(.din(n275),.dout(w_dff_B_pTm7TwKv4_0),.clk(gclk));
	jdff dff_B_ZFViDVo62_0(.din(w_dff_B_pTm7TwKv4_0),.dout(w_dff_B_ZFViDVo62_0),.clk(gclk));
	jdff dff_B_M4uKZ33d6_0(.din(w_dff_B_ZFViDVo62_0),.dout(w_dff_B_M4uKZ33d6_0),.clk(gclk));
	jdff dff_B_BzQbd4wn1_0(.din(w_dff_B_M4uKZ33d6_0),.dout(w_dff_B_BzQbd4wn1_0),.clk(gclk));
	jdff dff_B_2aQgTpKd8_0(.din(w_dff_B_BzQbd4wn1_0),.dout(w_dff_B_2aQgTpKd8_0),.clk(gclk));
	jdff dff_B_zqiK0Xpw6_1(.din(n315),.dout(w_dff_B_zqiK0Xpw6_1),.clk(gclk));
	jdff dff_A_ap4p4pgH8_0(.dout(w_n293_0[0]),.din(w_dff_A_ap4p4pgH8_0),.clk(gclk));
	jdff dff_B_Zb5l6RDP0_0(.din(n291),.dout(w_dff_B_Zb5l6RDP0_0),.clk(gclk));
	jdff dff_B_XihP7rBk7_0(.din(w_dff_B_Zb5l6RDP0_0),.dout(w_dff_B_XihP7rBk7_0),.clk(gclk));
	jdff dff_B_tm2ksOGf1_0(.din(w_dff_B_XihP7rBk7_0),.dout(w_dff_B_tm2ksOGf1_0),.clk(gclk));
	jdff dff_B_mKHebEnU9_0(.din(w_dff_B_tm2ksOGf1_0),.dout(w_dff_B_mKHebEnU9_0),.clk(gclk));
	jdff dff_B_TNL17A3L5_0(.din(w_dff_B_mKHebEnU9_0),.dout(w_dff_B_TNL17A3L5_0),.clk(gclk));
	jdff dff_A_bhTq7Q2L7_0(.dout(w_n296_0[0]),.din(w_dff_A_bhTq7Q2L7_0),.clk(gclk));
	jdff dff_B_RIYvRidS5_1(.din(n326),.dout(w_dff_B_RIYvRidS5_1),.clk(gclk));
	jdff dff_B_LSjvtylg8_0(.din(n282),.dout(w_dff_B_LSjvtylg8_0),.clk(gclk));
	jdff dff_B_MqE7YZoz4_0(.din(w_dff_B_LSjvtylg8_0),.dout(w_dff_B_MqE7YZoz4_0),.clk(gclk));
	jdff dff_B_ZTCuf4J51_0(.din(w_dff_B_MqE7YZoz4_0),.dout(w_dff_B_ZTCuf4J51_0),.clk(gclk));
	jdff dff_B_KlpllYaD6_0(.din(w_dff_B_ZTCuf4J51_0),.dout(w_dff_B_KlpllYaD6_0),.clk(gclk));
	jdff dff_B_DkoggYqW3_0(.din(w_dff_B_KlpllYaD6_0),.dout(w_dff_B_DkoggYqW3_0),.clk(gclk));
	jdff dff_A_lUbJeBKw1_0(.dout(w_n286_0[0]),.din(w_dff_A_lUbJeBKw1_0),.clk(gclk));
	jdff dff_A_Ht0QTSse1_0(.dout(w_n274_0[0]),.din(w_dff_A_Ht0QTSse1_0),.clk(gclk));
	jdff dff_A_qS4YkDag0_0(.dout(w_dff_A_Ht0QTSse1_0),.din(w_dff_A_qS4YkDag0_0),.clk(gclk));
	jdff dff_A_DxhtPWx42_0(.dout(w_dff_A_qS4YkDag0_0),.din(w_dff_A_DxhtPWx42_0),.clk(gclk));
	jdff dff_A_Y6V6tujw5_0(.dout(w_dff_A_DxhtPWx42_0),.din(w_dff_A_Y6V6tujw5_0),.clk(gclk));
	jdff dff_A_YbFHvBUL5_0(.dout(w_dff_A_Y6V6tujw5_0),.din(w_dff_A_YbFHvBUL5_0),.clk(gclk));
	jdff dff_A_ww5EVM0P1_0(.dout(w_dff_A_YbFHvBUL5_0),.din(w_dff_A_ww5EVM0P1_0),.clk(gclk));
	jdff dff_B_61851nHU8_1(.din(n300),.dout(w_dff_B_61851nHU8_1),.clk(gclk));
	jdff dff_B_Vy3M2GSb4_1(.din(w_dff_B_61851nHU8_1),.dout(w_dff_B_Vy3M2GSb4_1),.clk(gclk));
	jdff dff_B_lsmVxR8I6_1(.din(w_dff_B_Vy3M2GSb4_1),.dout(w_dff_B_lsmVxR8I6_1),.clk(gclk));
	jdff dff_B_OGRnpnlf3_1(.din(w_dff_B_lsmVxR8I6_1),.dout(w_dff_B_OGRnpnlf3_1),.clk(gclk));
	jdff dff_B_IOwF4Glq7_1(.din(w_dff_B_OGRnpnlf3_1),.dout(w_dff_B_IOwF4Glq7_1),.clk(gclk));
	jdff dff_B_63lnhOn55_1(.din(n301),.dout(w_dff_B_63lnhOn55_1),.clk(gclk));
	jdff dff_B_sMrOjCU75_1(.din(w_dff_B_63lnhOn55_1),.dout(w_dff_B_sMrOjCU75_1),.clk(gclk));
	jdff dff_B_sFDJB6s57_1(.din(w_dff_B_sMrOjCU75_1),.dout(w_dff_B_sFDJB6s57_1),.clk(gclk));
	jdff dff_B_ZAn4Sgqp9_1(.din(w_dff_B_sFDJB6s57_1),.dout(w_dff_B_ZAn4Sgqp9_1),.clk(gclk));
	jdff dff_B_P06ILHvw6_1(.din(w_dff_B_ZAn4Sgqp9_1),.dout(w_dff_B_P06ILHvw6_1),.clk(gclk));
	jdff dff_B_zZX3Faph4_1(.din(w_dff_B_P06ILHvw6_1),.dout(w_dff_B_zZX3Faph4_1),.clk(gclk));
	jdff dff_B_XaagROtF9_1(.din(w_dff_B_zZX3Faph4_1),.dout(w_dff_B_XaagROtF9_1),.clk(gclk));
	jdff dff_B_QEnaAqci1_1(.din(w_dff_B_XaagROtF9_1),.dout(w_dff_B_QEnaAqci1_1),.clk(gclk));
	jdff dff_B_EYcpcktT1_1(.din(w_dff_B_QEnaAqci1_1),.dout(w_dff_B_EYcpcktT1_1),.clk(gclk));
	jdff dff_B_s5oZxAZy6_1(.din(w_dff_B_EYcpcktT1_1),.dout(w_dff_B_s5oZxAZy6_1),.clk(gclk));
	jdff dff_B_Y3tVv5mi2_1(.din(w_dff_B_s5oZxAZy6_1),.dout(w_dff_B_Y3tVv5mi2_1),.clk(gclk));
	jdff dff_B_4EwAZuwG0_1(.din(w_dff_B_Y3tVv5mi2_1),.dout(w_dff_B_4EwAZuwG0_1),.clk(gclk));
	jdff dff_B_bPVohXzw7_1(.din(w_dff_B_4EwAZuwG0_1),.dout(w_dff_B_bPVohXzw7_1),.clk(gclk));
	jdff dff_B_XMUnQGRf5_1(.din(w_dff_B_bPVohXzw7_1),.dout(w_dff_B_XMUnQGRf5_1),.clk(gclk));
	jdff dff_B_XvNhl9Hs3_1(.din(w_dff_B_XMUnQGRf5_1),.dout(w_dff_B_XvNhl9Hs3_1),.clk(gclk));
	jdff dff_B_87glUefm9_1(.din(w_dff_B_XvNhl9Hs3_1),.dout(w_dff_B_87glUefm9_1),.clk(gclk));
	jdff dff_B_l5MATZEJ2_1(.din(w_dff_B_87glUefm9_1),.dout(w_dff_B_l5MATZEJ2_1),.clk(gclk));
	jdff dff_B_vCzdesii0_1(.din(w_dff_B_l5MATZEJ2_1),.dout(w_dff_B_vCzdesii0_1),.clk(gclk));
	jdff dff_B_jfxZeJNT7_1(.din(w_dff_B_vCzdesii0_1),.dout(w_dff_B_jfxZeJNT7_1),.clk(gclk));
	jdff dff_B_erZJyVKo4_1(.din(n242),.dout(w_dff_B_erZJyVKo4_1),.clk(gclk));
	jdff dff_B_RwErxWos9_1(.din(n252),.dout(w_dff_B_RwErxWos9_1),.clk(gclk));
	jdff dff_B_eADzKhT00_1(.din(n264),.dout(w_dff_B_eADzKhT00_1),.clk(gclk));
	jdff dff_B_zDm1Bszp8_0(.din(n262),.dout(w_dff_B_zDm1Bszp8_0),.clk(gclk));
	jdff dff_B_yx1vB4yl4_0(.din(w_dff_B_zDm1Bszp8_0),.dout(w_dff_B_yx1vB4yl4_0),.clk(gclk));
	jdff dff_B_Gh5mMvPZ6_0(.din(w_dff_B_yx1vB4yl4_0),.dout(w_dff_B_Gh5mMvPZ6_0),.clk(gclk));
	jdff dff_A_YvsfF6k72_1(.dout(w_n231_0[1]),.din(w_dff_A_YvsfF6k72_1),.clk(gclk));
	jdff dff_A_yqcP8mIO8_1(.dout(w_dff_A_YvsfF6k72_1),.din(w_dff_A_yqcP8mIO8_1),.clk(gclk));
	jdff dff_A_p4YkqInR2_1(.dout(w_dff_A_yqcP8mIO8_1),.din(w_dff_A_p4YkqInR2_1),.clk(gclk));
	jdff dff_A_wfABZNCu4_1(.dout(w_dff_A_p4YkqInR2_1),.din(w_dff_A_wfABZNCu4_1),.clk(gclk));
	jdff dff_A_nu4IWkEs7_1(.dout(w_dff_A_wfABZNCu4_1),.din(w_dff_A_nu4IWkEs7_1),.clk(gclk));
	jdff dff_A_ZkBAqm027_1(.dout(w_dff_A_nu4IWkEs7_1),.din(w_dff_A_ZkBAqm027_1),.clk(gclk));
	jdff dff_B_Vhe6vJ0b1_1(.din(n246),.dout(w_dff_B_Vhe6vJ0b1_1),.clk(gclk));
	jdff dff_B_tXGSSCjs9_0(.din(n244),.dout(w_dff_B_tXGSSCjs9_0),.clk(gclk));
	jdff dff_B_V4QtIwkQ2_0(.din(w_dff_B_tXGSSCjs9_0),.dout(w_dff_B_V4QtIwkQ2_0),.clk(gclk));
	jdff dff_B_rnzU1YTc2_0(.din(w_dff_B_V4QtIwkQ2_0),.dout(w_dff_B_rnzU1YTc2_0),.clk(gclk));
	jdff dff_B_wszG0AMj8_0(.din(w_dff_B_rnzU1YTc2_0),.dout(w_dff_B_wszG0AMj8_0),.clk(gclk));
	jdff dff_B_sJNE8zIO8_0(.din(w_dff_B_wszG0AMj8_0),.dout(w_dff_B_sJNE8zIO8_0),.clk(gclk));
	jdff dff_B_a1rqcxTg0_1(.din(n237),.dout(w_dff_B_a1rqcxTg0_1),.clk(gclk));
	jdff dff_B_qUUUr8lb5_0(.din(n235),.dout(w_dff_B_qUUUr8lb5_0),.clk(gclk));
	jdff dff_B_maInDkaC0_0(.din(w_dff_B_qUUUr8lb5_0),.dout(w_dff_B_maInDkaC0_0),.clk(gclk));
	jdff dff_B_39ayU2Sl8_0(.din(w_dff_B_maInDkaC0_0),.dout(w_dff_B_39ayU2Sl8_0),.clk(gclk));
	jdff dff_B_iR4wkDcl9_0(.din(w_dff_B_39ayU2Sl8_0),.dout(w_dff_B_iR4wkDcl9_0),.clk(gclk));
	jdff dff_A_3WSsRxUf9_0(.dout(w_n290_0[0]),.din(w_dff_A_3WSsRxUf9_0),.clk(gclk));
	jdff dff_A_se6up4Ss9_0(.dout(w_dff_A_3WSsRxUf9_0),.din(w_dff_A_se6up4Ss9_0),.clk(gclk));
	jdff dff_A_cHk6rDJq0_0(.dout(w_dff_A_se6up4Ss9_0),.din(w_dff_A_cHk6rDJq0_0),.clk(gclk));
	jdff dff_A_jCNboXfa1_0(.dout(w_dff_A_cHk6rDJq0_0),.din(w_dff_A_jCNboXfa1_0),.clk(gclk));
	jdff dff_A_IMLsThk60_0(.dout(w_dff_A_jCNboXfa1_0),.din(w_dff_A_IMLsThk60_0),.clk(gclk));
	jdff dff_A_GzvYsrTd6_0(.dout(w_dff_A_IMLsThk60_0),.din(w_dff_A_GzvYsrTd6_0),.clk(gclk));
	jdff dff_A_SKKqbJ652_0(.dout(w_n254_0[0]),.din(w_dff_A_SKKqbJ652_0),.clk(gclk));
	jdff dff_A_8zBGWutK1_0(.dout(w_dff_A_SKKqbJ652_0),.din(w_dff_A_8zBGWutK1_0),.clk(gclk));
	jdff dff_A_jT2p71gI7_0(.dout(w_dff_A_8zBGWutK1_0),.din(w_dff_A_jT2p71gI7_0),.clk(gclk));
	jdff dff_A_SXoqwkCD7_0(.dout(w_dff_A_jT2p71gI7_0),.din(w_dff_A_SXoqwkCD7_0),.clk(gclk));
	jdff dff_A_k33Srw5y6_0(.dout(w_dff_A_SXoqwkCD7_0),.din(w_dff_A_k33Srw5y6_0),.clk(gclk));
	jdff dff_A_kM1VUIek2_0(.dout(w_dff_A_k33Srw5y6_0),.din(w_dff_A_kM1VUIek2_0),.clk(gclk));
	jdff dff_A_eb3iF4Np2_0(.dout(w_n281_0[0]),.din(w_dff_A_eb3iF4Np2_0),.clk(gclk));
	jdff dff_A_nC1hyU7V1_0(.dout(w_dff_A_eb3iF4Np2_0),.din(w_dff_A_nC1hyU7V1_0),.clk(gclk));
	jdff dff_A_Ux3zMEJf2_0(.dout(w_dff_A_nC1hyU7V1_0),.din(w_dff_A_Ux3zMEJf2_0),.clk(gclk));
	jdff dff_A_BJy6mq5s7_0(.dout(w_dff_A_Ux3zMEJf2_0),.din(w_dff_A_BJy6mq5s7_0),.clk(gclk));
	jdff dff_A_q8Bkd44h3_0(.dout(w_dff_A_BJy6mq5s7_0),.din(w_dff_A_q8Bkd44h3_0),.clk(gclk));
	jdff dff_A_tVDtwLTa1_0(.dout(w_dff_A_q8Bkd44h3_0),.din(w_dff_A_tVDtwLTa1_0),.clk(gclk));
	jdff dff_B_akSLQiSm2_0(.din(n280),.dout(w_dff_B_akSLQiSm2_0),.clk(gclk));
	jdff dff_B_LBaWGVAn0_0(.din(w_dff_B_akSLQiSm2_0),.dout(w_dff_B_LBaWGVAn0_0),.clk(gclk));
	jdff dff_B_5AGmBoIP4_0(.din(w_dff_B_LBaWGVAn0_0),.dout(w_dff_B_5AGmBoIP4_0),.clk(gclk));
	jdff dff_B_kauUpNH26_0(.din(w_dff_B_5AGmBoIP4_0),.dout(w_dff_B_kauUpNH26_0),.clk(gclk));
	jdff dff_B_Cje7cwRF8_0(.din(w_dff_B_kauUpNH26_0),.dout(w_dff_B_Cje7cwRF8_0),.clk(gclk));
	jdff dff_B_uXF6yqlK1_0(.din(w_dff_B_Cje7cwRF8_0),.dout(w_dff_B_uXF6yqlK1_0),.clk(gclk));
	jdff dff_B_moVH5SBR5_1(.din(n187),.dout(w_dff_B_moVH5SBR5_1),.clk(gclk));
	jdff dff_B_0pCmD9204_1(.din(n202),.dout(w_dff_B_0pCmD9204_1),.clk(gclk));
	jdff dff_B_WWvHWYd57_1(.din(n221),.dout(w_dff_B_WWvHWYd57_1),.clk(gclk));
	jdff dff_A_ux7bgzkJ7_0(.dout(w_n224_0[0]),.din(w_dff_A_ux7bgzkJ7_0),.clk(gclk));
	jdff dff_A_IPNqJfBU6_0(.dout(w_dff_A_ux7bgzkJ7_0),.din(w_dff_A_IPNqJfBU6_0),.clk(gclk));
	jdff dff_A_KxMR96IR3_0(.dout(w_dff_A_IPNqJfBU6_0),.din(w_dff_A_KxMR96IR3_0),.clk(gclk));
	jdff dff_A_cNOtW5Mx9_0(.dout(w_dff_A_KxMR96IR3_0),.din(w_dff_A_cNOtW5Mx9_0),.clk(gclk));
	jdff dff_A_qOv4CHeU1_0(.dout(w_dff_A_cNOtW5Mx9_0),.din(w_dff_A_qOv4CHeU1_0),.clk(gclk));
	jdff dff_A_6c6mhX8v0_0(.dout(w_dff_A_qOv4CHeU1_0),.din(w_dff_A_6c6mhX8v0_0),.clk(gclk));
	jdff dff_A_fDii76br6_0(.dout(w_n222_0[0]),.din(w_dff_A_fDii76br6_0),.clk(gclk));
	jdff dff_A_zpHB0f9z4_0(.dout(w_dff_A_fDii76br6_0),.din(w_dff_A_zpHB0f9z4_0),.clk(gclk));
	jdff dff_A_llTFJ1Qm0_0(.dout(w_dff_A_zpHB0f9z4_0),.din(w_dff_A_llTFJ1Qm0_0),.clk(gclk));
	jdff dff_A_ybiPwF451_0(.dout(w_dff_A_llTFJ1Qm0_0),.din(w_dff_A_ybiPwF451_0),.clk(gclk));
	jdff dff_A_UrpyTP039_0(.dout(w_dff_A_ybiPwF451_0),.din(w_dff_A_UrpyTP039_0),.clk(gclk));
	jdff dff_B_T3Is5w2W2_2(.din(n222),.dout(w_dff_B_T3Is5w2W2_2),.clk(gclk));
	jdff dff_B_pKTwd5Z91_2(.din(w_dff_B_T3Is5w2W2_2),.dout(w_dff_B_pKTwd5Z91_2),.clk(gclk));
	jdff dff_B_CqtvmWDt2_2(.din(w_dff_B_pKTwd5Z91_2),.dout(w_dff_B_CqtvmWDt2_2),.clk(gclk));
	jdff dff_B_08764Txh0_2(.din(w_dff_B_CqtvmWDt2_2),.dout(w_dff_B_08764Txh0_2),.clk(gclk));
	jdff dff_B_pXtP3Vtx6_2(.din(w_dff_B_08764Txh0_2),.dout(w_dff_B_pXtP3Vtx6_2),.clk(gclk));
	jdff dff_B_eKkeObvC3_2(.din(w_dff_B_pXtP3Vtx6_2),.dout(w_dff_B_eKkeObvC3_2),.clk(gclk));
	jdff dff_B_OJgdGmN87_2(.din(w_dff_B_eKkeObvC3_2),.dout(w_dff_B_OJgdGmN87_2),.clk(gclk));
	jdff dff_B_pSVPQ7HT1_2(.din(w_dff_B_OJgdGmN87_2),.dout(w_dff_B_pSVPQ7HT1_2),.clk(gclk));
	jdff dff_B_t92uup1W4_2(.din(w_dff_B_pSVPQ7HT1_2),.dout(w_dff_B_t92uup1W4_2),.clk(gclk));
	jdff dff_B_vlqbdS308_2(.din(w_dff_B_t92uup1W4_2),.dout(w_dff_B_vlqbdS308_2),.clk(gclk));
	jdff dff_B_jnVQKEtB0_2(.din(w_dff_B_vlqbdS308_2),.dout(w_dff_B_jnVQKEtB0_2),.clk(gclk));
	jdff dff_B_6aDjtOHo2_2(.din(w_dff_B_jnVQKEtB0_2),.dout(w_dff_B_6aDjtOHo2_2),.clk(gclk));
	jdff dff_B_12btdkct8_2(.din(w_dff_B_6aDjtOHo2_2),.dout(w_dff_B_12btdkct8_2),.clk(gclk));
	jdff dff_B_gbWZni8G5_2(.din(w_dff_B_12btdkct8_2),.dout(w_dff_B_gbWZni8G5_2),.clk(gclk));
	jdff dff_A_Grp4gKbN7_0(.dout(w_G115gat_0[0]),.din(w_dff_A_Grp4gKbN7_0),.clk(gclk));
	jdff dff_A_ITG7dhPe3_0(.dout(w_dff_A_Grp4gKbN7_0),.din(w_dff_A_ITG7dhPe3_0),.clk(gclk));
	jdff dff_A_rOAgBkxG5_0(.dout(w_dff_A_ITG7dhPe3_0),.din(w_dff_A_rOAgBkxG5_0),.clk(gclk));
	jdff dff_A_e8bdT4yK3_0(.dout(w_dff_A_rOAgBkxG5_0),.din(w_dff_A_e8bdT4yK3_0),.clk(gclk));
	jdff dff_A_SDe99cyn0_0(.dout(w_dff_A_e8bdT4yK3_0),.din(w_dff_A_SDe99cyn0_0),.clk(gclk));
	jdff dff_A_e8PApaLy4_0(.dout(w_dff_A_SDe99cyn0_0),.din(w_dff_A_e8PApaLy4_0),.clk(gclk));
	jdff dff_A_KHl453nB9_0(.dout(w_dff_A_e8PApaLy4_0),.din(w_dff_A_KHl453nB9_0),.clk(gclk));
	jdff dff_A_Jz1BAu5o4_0(.dout(w_dff_A_KHl453nB9_0),.din(w_dff_A_Jz1BAu5o4_0),.clk(gclk));
	jdff dff_A_W99BY7sm6_0(.dout(w_dff_A_Jz1BAu5o4_0),.din(w_dff_A_W99BY7sm6_0),.clk(gclk));
	jdff dff_A_8UNSU2Zm8_0(.dout(w_dff_A_W99BY7sm6_0),.din(w_dff_A_8UNSU2Zm8_0),.clk(gclk));
	jdff dff_A_vo7ecOzY8_0(.dout(w_dff_A_8UNSU2Zm8_0),.din(w_dff_A_vo7ecOzY8_0),.clk(gclk));
	jdff dff_A_cNYE0Rxi5_0(.dout(w_dff_A_vo7ecOzY8_0),.din(w_dff_A_cNYE0Rxi5_0),.clk(gclk));
	jdff dff_A_oM79tBM66_0(.dout(w_dff_A_cNYE0Rxi5_0),.din(w_dff_A_oM79tBM66_0),.clk(gclk));
	jdff dff_A_JO4lQiNv4_0(.dout(w_dff_A_oM79tBM66_0),.din(w_dff_A_JO4lQiNv4_0),.clk(gclk));
	jdff dff_A_AvwkGZtH5_0(.dout(w_dff_A_JO4lQiNv4_0),.din(w_dff_A_AvwkGZtH5_0),.clk(gclk));
	jdff dff_A_9KkDxQ5a3_1(.dout(w_n219_0[1]),.din(w_dff_A_9KkDxQ5a3_1),.clk(gclk));
	jdff dff_A_d8smjoO24_1(.dout(w_dff_A_9KkDxQ5a3_1),.din(w_dff_A_d8smjoO24_1),.clk(gclk));
	jdff dff_A_iYCqwx7Q1_1(.dout(w_dff_A_d8smjoO24_1),.din(w_dff_A_iYCqwx7Q1_1),.clk(gclk));
	jdff dff_A_LmDCxI092_1(.dout(w_dff_A_iYCqwx7Q1_1),.din(w_dff_A_LmDCxI092_1),.clk(gclk));
	jdff dff_A_RzoDSxuh6_0(.dout(w_n217_0[0]),.din(w_dff_A_RzoDSxuh6_0),.clk(gclk));
	jdff dff_A_87mnJcZt7_0(.dout(w_dff_A_RzoDSxuh6_0),.din(w_dff_A_87mnJcZt7_0),.clk(gclk));
	jdff dff_A_Cn4HUcMZ8_0(.dout(w_dff_A_87mnJcZt7_0),.din(w_dff_A_Cn4HUcMZ8_0),.clk(gclk));
	jdff dff_A_4WHONs2a7_0(.dout(w_dff_A_Cn4HUcMZ8_0),.din(w_dff_A_4WHONs2a7_0),.clk(gclk));
	jdff dff_A_tf2Eq1HF3_0(.dout(w_dff_A_4WHONs2a7_0),.din(w_dff_A_tf2Eq1HF3_0),.clk(gclk));
	jdff dff_A_5dQwUhWN5_0(.dout(w_dff_A_tf2Eq1HF3_0),.din(w_dff_A_5dQwUhWN5_0),.clk(gclk));
	jdff dff_A_XVPZIjSM2_0(.dout(w_dff_A_5dQwUhWN5_0),.din(w_dff_A_XVPZIjSM2_0),.clk(gclk));
	jdff dff_A_bKBSNtxC2_0(.dout(w_dff_A_XVPZIjSM2_0),.din(w_dff_A_bKBSNtxC2_0),.clk(gclk));
	jdff dff_A_hQecb5Yc4_0(.dout(w_dff_A_bKBSNtxC2_0),.din(w_dff_A_hQecb5Yc4_0),.clk(gclk));
	jdff dff_A_GYxAzLjh8_0(.dout(w_dff_A_hQecb5Yc4_0),.din(w_dff_A_GYxAzLjh8_0),.clk(gclk));
	jdff dff_A_zSHVQ4E95_0(.dout(w_dff_A_GYxAzLjh8_0),.din(w_dff_A_zSHVQ4E95_0),.clk(gclk));
	jdff dff_B_nMRYpbD35_2(.din(n217),.dout(w_dff_B_nMRYpbD35_2),.clk(gclk));
	jdff dff_B_vCdUxLIY4_2(.din(w_dff_B_nMRYpbD35_2),.dout(w_dff_B_vCdUxLIY4_2),.clk(gclk));
	jdff dff_B_ZIWcIQdJ4_2(.din(w_dff_B_vCdUxLIY4_2),.dout(w_dff_B_ZIWcIQdJ4_2),.clk(gclk));
	jdff dff_B_JyJZ34XK2_2(.din(w_dff_B_ZIWcIQdJ4_2),.dout(w_dff_B_JyJZ34XK2_2),.clk(gclk));
	jdff dff_B_zRU6HOQA3_2(.din(w_dff_B_JyJZ34XK2_2),.dout(w_dff_B_zRU6HOQA3_2),.clk(gclk));
	jdff dff_B_qAJHj5iF4_2(.din(w_dff_B_zRU6HOQA3_2),.dout(w_dff_B_qAJHj5iF4_2),.clk(gclk));
	jdff dff_B_Z2zh11bp5_2(.din(w_dff_B_qAJHj5iF4_2),.dout(w_dff_B_Z2zh11bp5_2),.clk(gclk));
	jdff dff_B_fgU23e0C8_2(.din(w_dff_B_Z2zh11bp5_2),.dout(w_dff_B_fgU23e0C8_2),.clk(gclk));
	jdff dff_A_8xMlCICc9_0(.dout(w_G40gat_0[0]),.din(w_dff_A_8xMlCICc9_0),.clk(gclk));
	jdff dff_A_n85eMn4U7_0(.dout(w_dff_A_8xMlCICc9_0),.din(w_dff_A_n85eMn4U7_0),.clk(gclk));
	jdff dff_A_hP8Jo5fs6_0(.dout(w_dff_A_n85eMn4U7_0),.din(w_dff_A_hP8Jo5fs6_0),.clk(gclk));
	jdff dff_A_3GJcADem5_0(.dout(w_dff_A_hP8Jo5fs6_0),.din(w_dff_A_3GJcADem5_0),.clk(gclk));
	jdff dff_A_ayoFeQod0_0(.dout(w_dff_A_3GJcADem5_0),.din(w_dff_A_ayoFeQod0_0),.clk(gclk));
	jdff dff_A_qpPAXIMO3_0(.dout(w_dff_A_ayoFeQod0_0),.din(w_dff_A_qpPAXIMO3_0),.clk(gclk));
	jdff dff_A_wXmZkkXC5_0(.dout(w_dff_A_qpPAXIMO3_0),.din(w_dff_A_wXmZkkXC5_0),.clk(gclk));
	jdff dff_A_Ztxnv9k10_0(.dout(w_dff_A_wXmZkkXC5_0),.din(w_dff_A_Ztxnv9k10_0),.clk(gclk));
	jdff dff_A_hzillUTC0_0(.dout(w_dff_A_Ztxnv9k10_0),.din(w_dff_A_hzillUTC0_0),.clk(gclk));
	jdff dff_A_OybFytYO1_0(.dout(w_dff_A_hzillUTC0_0),.din(w_dff_A_OybFytYO1_0),.clk(gclk));
	jdff dff_A_kwAPfovI5_0(.dout(w_dff_A_OybFytYO1_0),.din(w_dff_A_kwAPfovI5_0),.clk(gclk));
	jdff dff_A_T4MwwXy39_0(.dout(w_dff_A_kwAPfovI5_0),.din(w_dff_A_T4MwwXy39_0),.clk(gclk));
	jdff dff_A_0iTrAXob9_0(.dout(w_dff_A_T4MwwXy39_0),.din(w_dff_A_0iTrAXob9_0),.clk(gclk));
	jdff dff_A_piB35lYS0_0(.dout(w_dff_A_0iTrAXob9_0),.din(w_dff_A_piB35lYS0_0),.clk(gclk));
	jdff dff_A_kYFkFj4w9_0(.dout(w_dff_A_piB35lYS0_0),.din(w_dff_A_kYFkFj4w9_0),.clk(gclk));
	jdff dff_A_pXpSgiNB9_0(.dout(w_dff_A_kYFkFj4w9_0),.din(w_dff_A_pXpSgiNB9_0),.clk(gclk));
	jdff dff_A_y6Ii1q5d4_0(.dout(w_dff_A_pXpSgiNB9_0),.din(w_dff_A_y6Ii1q5d4_0),.clk(gclk));
	jdff dff_A_KA6riDI94_0(.dout(w_dff_A_y6Ii1q5d4_0),.din(w_dff_A_KA6riDI94_0),.clk(gclk));
	jdff dff_A_flqTqVj67_0(.dout(w_dff_A_KA6riDI94_0),.din(w_dff_A_flqTqVj67_0),.clk(gclk));
	jdff dff_A_diYIX76x0_0(.dout(w_dff_A_flqTqVj67_0),.din(w_dff_A_diYIX76x0_0),.clk(gclk));
	jdff dff_B_lnn5Uzfq6_1(.din(n214),.dout(w_dff_B_lnn5Uzfq6_1),.clk(gclk));
	jdff dff_B_U98fcXty5_1(.din(w_dff_B_lnn5Uzfq6_1),.dout(w_dff_B_U98fcXty5_1),.clk(gclk));
	jdff dff_B_xlcXHhRu7_1(.din(w_dff_B_U98fcXty5_1),.dout(w_dff_B_xlcXHhRu7_1),.clk(gclk));
	jdff dff_B_efK2R0bh5_1(.din(w_dff_B_xlcXHhRu7_1),.dout(w_dff_B_efK2R0bh5_1),.clk(gclk));
	jdff dff_B_X67VoH9R1_1(.din(w_dff_B_efK2R0bh5_1),.dout(w_dff_B_X67VoH9R1_1),.clk(gclk));
	jdff dff_B_TGwtTXDD7_1(.din(w_dff_B_X67VoH9R1_1),.dout(w_dff_B_TGwtTXDD7_1),.clk(gclk));
	jdff dff_B_00zlxIno6_1(.din(w_dff_B_TGwtTXDD7_1),.dout(w_dff_B_00zlxIno6_1),.clk(gclk));
	jdff dff_B_6KJG3Flh1_1(.din(w_dff_B_00zlxIno6_1),.dout(w_dff_B_6KJG3Flh1_1),.clk(gclk));
	jdff dff_B_fALiyNYM4_1(.din(w_dff_B_6KJG3Flh1_1),.dout(w_dff_B_fALiyNYM4_1),.clk(gclk));
	jdff dff_B_z1LzTmC00_1(.din(w_dff_B_fALiyNYM4_1),.dout(w_dff_B_z1LzTmC00_1),.clk(gclk));
	jdff dff_B_B01hDh9Y3_1(.din(w_dff_B_z1LzTmC00_1),.dout(w_dff_B_B01hDh9Y3_1),.clk(gclk));
	jdff dff_B_o98iBe3S6_1(.din(w_dff_B_B01hDh9Y3_1),.dout(w_dff_B_o98iBe3S6_1),.clk(gclk));
	jdff dff_B_xElPkw5s0_1(.din(n209),.dout(w_dff_B_xElPkw5s0_1),.clk(gclk));
	jdff dff_B_W5Y98niU1_1(.din(w_dff_B_xElPkw5s0_1),.dout(w_dff_B_W5Y98niU1_1),.clk(gclk));
	jdff dff_B_1hD0ELZz5_1(.din(w_dff_B_W5Y98niU1_1),.dout(w_dff_B_1hD0ELZz5_1),.clk(gclk));
	jdff dff_B_L28FJEj32_1(.din(w_dff_B_1hD0ELZz5_1),.dout(w_dff_B_L28FJEj32_1),.clk(gclk));
	jdff dff_B_bUzvdw0K2_1(.din(w_dff_B_L28FJEj32_1),.dout(w_dff_B_bUzvdw0K2_1),.clk(gclk));
	jdff dff_B_AXbgqMsT7_1(.din(w_dff_B_bUzvdw0K2_1),.dout(w_dff_B_AXbgqMsT7_1),.clk(gclk));
	jdff dff_B_EGEo9Tis2_1(.din(w_dff_B_AXbgqMsT7_1),.dout(w_dff_B_EGEo9Tis2_1),.clk(gclk));
	jdff dff_B_krtebK9K0_1(.din(w_dff_B_EGEo9Tis2_1),.dout(w_dff_B_krtebK9K0_1),.clk(gclk));
	jdff dff_B_qitdhjvU1_1(.din(w_dff_B_krtebK9K0_1),.dout(w_dff_B_qitdhjvU1_1),.clk(gclk));
	jdff dff_B_YrtmM10h8_1(.din(w_dff_B_qitdhjvU1_1),.dout(w_dff_B_YrtmM10h8_1),.clk(gclk));
	jdff dff_B_HmraLxQV5_1(.din(w_dff_B_YrtmM10h8_1),.dout(w_dff_B_HmraLxQV5_1),.clk(gclk));
	jdff dff_B_A6mZnrIx9_1(.din(w_dff_B_HmraLxQV5_1),.dout(w_dff_B_A6mZnrIx9_1),.clk(gclk));
	jdff dff_B_IRfLmUY64_1(.din(w_dff_B_A6mZnrIx9_1),.dout(w_dff_B_IRfLmUY64_1),.clk(gclk));
	jdff dff_B_dpOwkNU81_1(.din(w_dff_B_IRfLmUY64_1),.dout(w_dff_B_dpOwkNU81_1),.clk(gclk));
	jdff dff_A_TpSj3xwa4_0(.dout(w_G14gat_0[0]),.din(w_dff_A_TpSj3xwa4_0),.clk(gclk));
	jdff dff_A_cnwC30Rj0_0(.dout(w_dff_A_TpSj3xwa4_0),.din(w_dff_A_cnwC30Rj0_0),.clk(gclk));
	jdff dff_A_YUca2dnA6_0(.dout(w_dff_A_cnwC30Rj0_0),.din(w_dff_A_YUca2dnA6_0),.clk(gclk));
	jdff dff_A_nyA0KeG70_0(.dout(w_dff_A_YUca2dnA6_0),.din(w_dff_A_nyA0KeG70_0),.clk(gclk));
	jdff dff_A_87Dcb33u9_0(.dout(w_dff_A_nyA0KeG70_0),.din(w_dff_A_87Dcb33u9_0),.clk(gclk));
	jdff dff_A_QRl0R2Rj7_0(.dout(w_dff_A_87Dcb33u9_0),.din(w_dff_A_QRl0R2Rj7_0),.clk(gclk));
	jdff dff_A_hNQMmCzg6_0(.dout(w_dff_A_QRl0R2Rj7_0),.din(w_dff_A_hNQMmCzg6_0),.clk(gclk));
	jdff dff_A_LLwNLMZU3_0(.dout(w_dff_A_hNQMmCzg6_0),.din(w_dff_A_LLwNLMZU3_0),.clk(gclk));
	jdff dff_A_zSyOxV917_0(.dout(w_dff_A_LLwNLMZU3_0),.din(w_dff_A_zSyOxV917_0),.clk(gclk));
	jdff dff_A_I6lDnbCy9_0(.dout(w_dff_A_zSyOxV917_0),.din(w_dff_A_I6lDnbCy9_0),.clk(gclk));
	jdff dff_A_aSyy6zo64_0(.dout(w_dff_A_I6lDnbCy9_0),.din(w_dff_A_aSyy6zo64_0),.clk(gclk));
	jdff dff_A_aNyeiOYG6_0(.dout(w_dff_A_aSyy6zo64_0),.din(w_dff_A_aNyeiOYG6_0),.clk(gclk));
	jdff dff_A_Srj0DVv62_0(.dout(w_dff_A_aNyeiOYG6_0),.din(w_dff_A_Srj0DVv62_0),.clk(gclk));
	jdff dff_A_7g9FVgZL0_0(.dout(w_dff_A_Srj0DVv62_0),.din(w_dff_A_7g9FVgZL0_0),.clk(gclk));
	jdff dff_A_X0N0VDcb5_0(.dout(w_dff_A_7g9FVgZL0_0),.din(w_dff_A_X0N0VDcb5_0),.clk(gclk));
	jdff dff_A_ZqZMyaQl6_1(.dout(w_G14gat_0[1]),.din(w_dff_A_ZqZMyaQl6_1),.clk(gclk));
	jdff dff_A_aTIWMwVj2_1(.dout(w_dff_A_ZqZMyaQl6_1),.din(w_dff_A_aTIWMwVj2_1),.clk(gclk));
	jdff dff_A_le4NPD2O9_1(.dout(w_dff_A_aTIWMwVj2_1),.din(w_dff_A_le4NPD2O9_1),.clk(gclk));
	jdff dff_A_ybQYTo8r8_1(.dout(w_dff_A_le4NPD2O9_1),.din(w_dff_A_ybQYTo8r8_1),.clk(gclk));
	jdff dff_A_pLdptZsi5_1(.dout(w_dff_A_ybQYTo8r8_1),.din(w_dff_A_pLdptZsi5_1),.clk(gclk));
	jdff dff_A_QL7Q4aix8_1(.dout(w_dff_A_pLdptZsi5_1),.din(w_dff_A_QL7Q4aix8_1),.clk(gclk));
	jdff dff_A_vkziZMf91_1(.dout(w_dff_A_QL7Q4aix8_1),.din(w_dff_A_vkziZMf91_1),.clk(gclk));
	jdff dff_A_8zERPKfg0_1(.dout(w_dff_A_vkziZMf91_1),.din(w_dff_A_8zERPKfg0_1),.clk(gclk));
	jdff dff_A_WxUBDYyB5_1(.dout(w_dff_A_8zERPKfg0_1),.din(w_dff_A_WxUBDYyB5_1),.clk(gclk));
	jdff dff_A_GCO729jO1_1(.dout(w_dff_A_WxUBDYyB5_1),.din(w_dff_A_GCO729jO1_1),.clk(gclk));
	jdff dff_A_Sg2vU5sp9_1(.dout(w_dff_A_GCO729jO1_1),.din(w_dff_A_Sg2vU5sp9_1),.clk(gclk));
	jdff dff_A_n2X8c3xd3_1(.dout(w_dff_A_Sg2vU5sp9_1),.din(w_dff_A_n2X8c3xd3_1),.clk(gclk));
	jdff dff_A_bQX8fFmd2_1(.dout(w_dff_A_n2X8c3xd3_1),.din(w_dff_A_bQX8fFmd2_1),.clk(gclk));
	jdff dff_A_FukfDVB72_1(.dout(w_dff_A_bQX8fFmd2_1),.din(w_dff_A_FukfDVB72_1),.clk(gclk));
	jdff dff_A_IVEt6Yi41_1(.dout(w_dff_A_FukfDVB72_1),.din(w_dff_A_IVEt6Yi41_1),.clk(gclk));
	jdff dff_A_rnL2bv6w1_1(.dout(w_dff_A_IVEt6Yi41_1),.din(w_dff_A_rnL2bv6w1_1),.clk(gclk));
	jdff dff_A_9zWOeDKj4_1(.dout(w_dff_A_rnL2bv6w1_1),.din(w_dff_A_9zWOeDKj4_1),.clk(gclk));
	jdff dff_A_PX4wzWm83_1(.dout(w_dff_A_9zWOeDKj4_1),.din(w_dff_A_PX4wzWm83_1),.clk(gclk));
	jdff dff_A_F43mayrn8_1(.dout(w_dff_A_PX4wzWm83_1),.din(w_dff_A_F43mayrn8_1),.clk(gclk));
	jdff dff_A_reYrKxhI4_1(.dout(w_dff_A_F43mayrn8_1),.din(w_dff_A_reYrKxhI4_1),.clk(gclk));
	jdff dff_A_5O11Kk6m7_0(.dout(w_n205_0[0]),.din(w_dff_A_5O11Kk6m7_0),.clk(gclk));
	jdff dff_A_jHfTwugk2_0(.dout(w_dff_A_5O11Kk6m7_0),.din(w_dff_A_jHfTwugk2_0),.clk(gclk));
	jdff dff_A_Z39AWxCp2_0(.dout(w_dff_A_jHfTwugk2_0),.din(w_dff_A_Z39AWxCp2_0),.clk(gclk));
	jdff dff_A_QncNGc8c7_0(.dout(w_dff_A_Z39AWxCp2_0),.din(w_dff_A_QncNGc8c7_0),.clk(gclk));
	jdff dff_A_OnOWwz199_0(.dout(w_dff_A_QncNGc8c7_0),.din(w_dff_A_OnOWwz199_0),.clk(gclk));
	jdff dff_A_mutchN9n9_0(.dout(w_dff_A_OnOWwz199_0),.din(w_dff_A_mutchN9n9_0),.clk(gclk));
	jdff dff_B_5na9E6hu8_2(.din(n205),.dout(w_dff_B_5na9E6hu8_2),.clk(gclk));
	jdff dff_B_lldkz9KD6_2(.din(w_dff_B_5na9E6hu8_2),.dout(w_dff_B_lldkz9KD6_2),.clk(gclk));
	jdff dff_B_eXp3ymoj3_2(.din(w_dff_B_lldkz9KD6_2),.dout(w_dff_B_eXp3ymoj3_2),.clk(gclk));
	jdff dff_B_w50sHWmX1_2(.din(w_dff_B_eXp3ymoj3_2),.dout(w_dff_B_w50sHWmX1_2),.clk(gclk));
	jdff dff_B_momk3OCZ7_2(.din(w_dff_B_w50sHWmX1_2),.dout(w_dff_B_momk3OCZ7_2),.clk(gclk));
	jdff dff_B_VPnhVvQf6_2(.din(w_dff_B_momk3OCZ7_2),.dout(w_dff_B_VPnhVvQf6_2),.clk(gclk));
	jdff dff_B_i7T2ylon8_2(.din(w_dff_B_VPnhVvQf6_2),.dout(w_dff_B_i7T2ylon8_2),.clk(gclk));
	jdff dff_B_Hg1wGNpr9_2(.din(w_dff_B_i7T2ylon8_2),.dout(w_dff_B_Hg1wGNpr9_2),.clk(gclk));
	jdff dff_B_XQEDxvVJ3_2(.din(w_dff_B_Hg1wGNpr9_2),.dout(w_dff_B_XQEDxvVJ3_2),.clk(gclk));
	jdff dff_B_8WWWUYmp0_2(.din(w_dff_B_XQEDxvVJ3_2),.dout(w_dff_B_8WWWUYmp0_2),.clk(gclk));
	jdff dff_B_pPgTgPVb9_2(.din(w_dff_B_8WWWUYmp0_2),.dout(w_dff_B_pPgTgPVb9_2),.clk(gclk));
	jdff dff_B_b3BVX2oY0_2(.din(w_dff_B_pPgTgPVb9_2),.dout(w_dff_B_b3BVX2oY0_2),.clk(gclk));
	jdff dff_B_uUvTNaPX9_2(.din(w_dff_B_b3BVX2oY0_2),.dout(w_dff_B_uUvTNaPX9_2),.clk(gclk));
	jdff dff_A_2VNDQKNF4_0(.dout(w_G92gat_0[0]),.din(w_dff_A_2VNDQKNF4_0),.clk(gclk));
	jdff dff_A_VRPZQ8vi8_0(.dout(w_dff_A_2VNDQKNF4_0),.din(w_dff_A_VRPZQ8vi8_0),.clk(gclk));
	jdff dff_A_K0v8OTU29_0(.dout(w_dff_A_VRPZQ8vi8_0),.din(w_dff_A_K0v8OTU29_0),.clk(gclk));
	jdff dff_A_6O5rJf7T4_0(.dout(w_dff_A_K0v8OTU29_0),.din(w_dff_A_6O5rJf7T4_0),.clk(gclk));
	jdff dff_A_6cl3ISZv3_0(.dout(w_dff_A_6O5rJf7T4_0),.din(w_dff_A_6cl3ISZv3_0),.clk(gclk));
	jdff dff_A_dLTShI6e4_0(.dout(w_dff_A_6cl3ISZv3_0),.din(w_dff_A_dLTShI6e4_0),.clk(gclk));
	jdff dff_A_lEY5TJhc5_0(.dout(w_dff_A_dLTShI6e4_0),.din(w_dff_A_lEY5TJhc5_0),.clk(gclk));
	jdff dff_A_YSebzq7q0_0(.dout(w_dff_A_lEY5TJhc5_0),.din(w_dff_A_YSebzq7q0_0),.clk(gclk));
	jdff dff_A_EPWGFcJD8_0(.dout(w_dff_A_YSebzq7q0_0),.din(w_dff_A_EPWGFcJD8_0),.clk(gclk));
	jdff dff_A_IVYwyVLb4_0(.dout(w_dff_A_EPWGFcJD8_0),.din(w_dff_A_IVYwyVLb4_0),.clk(gclk));
	jdff dff_A_TNf5Xzci9_0(.dout(w_dff_A_IVYwyVLb4_0),.din(w_dff_A_TNf5Xzci9_0),.clk(gclk));
	jdff dff_A_SRzfEq2P7_0(.dout(w_dff_A_TNf5Xzci9_0),.din(w_dff_A_SRzfEq2P7_0),.clk(gclk));
	jdff dff_A_Sa2BPSPj2_0(.dout(w_dff_A_SRzfEq2P7_0),.din(w_dff_A_Sa2BPSPj2_0),.clk(gclk));
	jdff dff_A_ZNR42zaU9_0(.dout(w_dff_A_Sa2BPSPj2_0),.din(w_dff_A_ZNR42zaU9_0),.clk(gclk));
	jdff dff_A_RlohIgWY0_0(.dout(w_dff_A_ZNR42zaU9_0),.din(w_dff_A_RlohIgWY0_0),.clk(gclk));
	jdff dff_A_8YKBPe6X5_0(.dout(w_dff_A_RlohIgWY0_0),.din(w_dff_A_8YKBPe6X5_0),.clk(gclk));
	jdff dff_A_Xs0xBlaI4_0(.dout(w_dff_A_8YKBPe6X5_0),.din(w_dff_A_Xs0xBlaI4_0),.clk(gclk));
	jdff dff_A_xMwM09Dw7_0(.dout(w_dff_A_Xs0xBlaI4_0),.din(w_dff_A_xMwM09Dw7_0),.clk(gclk));
	jdff dff_A_ec6FnCUB3_0(.dout(w_dff_A_xMwM09Dw7_0),.din(w_dff_A_ec6FnCUB3_0),.clk(gclk));
	jdff dff_A_hTvL5vzG1_0(.dout(w_dff_A_ec6FnCUB3_0),.din(w_dff_A_hTvL5vzG1_0),.clk(gclk));
	jdff dff_A_83dePEjo1_1(.dout(w_G92gat_0[1]),.din(w_dff_A_83dePEjo1_1),.clk(gclk));
	jdff dff_A_2kmHN2nr2_1(.dout(w_dff_A_83dePEjo1_1),.din(w_dff_A_2kmHN2nr2_1),.clk(gclk));
	jdff dff_A_bICRxTcp6_1(.dout(w_dff_A_2kmHN2nr2_1),.din(w_dff_A_bICRxTcp6_1),.clk(gclk));
	jdff dff_A_A6pcBdQW9_1(.dout(w_dff_A_bICRxTcp6_1),.din(w_dff_A_A6pcBdQW9_1),.clk(gclk));
	jdff dff_A_dqA1iTsp5_1(.dout(w_dff_A_A6pcBdQW9_1),.din(w_dff_A_dqA1iTsp5_1),.clk(gclk));
	jdff dff_A_2p6TzBdR0_1(.dout(w_dff_A_dqA1iTsp5_1),.din(w_dff_A_2p6TzBdR0_1),.clk(gclk));
	jdff dff_A_nOdvEM2O8_1(.dout(w_dff_A_2p6TzBdR0_1),.din(w_dff_A_nOdvEM2O8_1),.clk(gclk));
	jdff dff_A_lem8xaPx7_1(.dout(w_dff_A_nOdvEM2O8_1),.din(w_dff_A_lem8xaPx7_1),.clk(gclk));
	jdff dff_A_w29xGCwv0_1(.dout(w_dff_A_lem8xaPx7_1),.din(w_dff_A_w29xGCwv0_1),.clk(gclk));
	jdff dff_A_EyvGYo8f4_1(.dout(w_dff_A_w29xGCwv0_1),.din(w_dff_A_EyvGYo8f4_1),.clk(gclk));
	jdff dff_A_rNyqQz2R0_1(.dout(w_dff_A_EyvGYo8f4_1),.din(w_dff_A_rNyqQz2R0_1),.clk(gclk));
	jdff dff_A_ZkEt66zK0_1(.dout(w_dff_A_rNyqQz2R0_1),.din(w_dff_A_ZkEt66zK0_1),.clk(gclk));
	jdff dff_A_b8m4tGwy5_1(.dout(w_dff_A_ZkEt66zK0_1),.din(w_dff_A_b8m4tGwy5_1),.clk(gclk));
	jdff dff_A_Cja6zkSj7_1(.dout(w_dff_A_b8m4tGwy5_1),.din(w_dff_A_Cja6zkSj7_1),.clk(gclk));
	jdff dff_A_lzEL013z8_0(.dout(w_n204_0[0]),.din(w_dff_A_lzEL013z8_0),.clk(gclk));
	jdff dff_A_HitMEIcW0_0(.dout(w_dff_A_lzEL013z8_0),.din(w_dff_A_HitMEIcW0_0),.clk(gclk));
	jdff dff_A_Z1SZBG4I3_0(.dout(w_dff_A_HitMEIcW0_0),.din(w_dff_A_Z1SZBG4I3_0),.clk(gclk));
	jdff dff_A_vgxR4BZu9_0(.dout(w_dff_A_Z1SZBG4I3_0),.din(w_dff_A_vgxR4BZu9_0),.clk(gclk));
	jdff dff_A_OcK3Z1p87_0(.dout(w_dff_A_vgxR4BZu9_0),.din(w_dff_A_OcK3Z1p87_0),.clk(gclk));
	jdff dff_A_kJY4IHWD0_0(.dout(w_dff_A_OcK3Z1p87_0),.din(w_dff_A_kJY4IHWD0_0),.clk(gclk));
	jdff dff_A_VlCqvEiy4_0(.dout(w_n198_0[0]),.din(w_dff_A_VlCqvEiy4_0),.clk(gclk));
	jdff dff_A_3UtBEZuj6_0(.dout(w_dff_A_VlCqvEiy4_0),.din(w_dff_A_3UtBEZuj6_0),.clk(gclk));
	jdff dff_A_fHwwK6F40_0(.dout(w_dff_A_3UtBEZuj6_0),.din(w_dff_A_fHwwK6F40_0),.clk(gclk));
	jdff dff_A_UKVnAVN40_0(.dout(w_dff_A_fHwwK6F40_0),.din(w_dff_A_UKVnAVN40_0),.clk(gclk));
	jdff dff_A_gGr99vMR6_0(.dout(w_dff_A_UKVnAVN40_0),.din(w_dff_A_gGr99vMR6_0),.clk(gclk));
	jdff dff_A_0CyklLM18_0(.dout(w_dff_A_gGr99vMR6_0),.din(w_dff_A_0CyklLM18_0),.clk(gclk));
	jdff dff_B_qUqSm9GJ4_2(.din(n198),.dout(w_dff_B_qUqSm9GJ4_2),.clk(gclk));
	jdff dff_B_7fuvmvCx4_2(.din(w_dff_B_qUqSm9GJ4_2),.dout(w_dff_B_7fuvmvCx4_2),.clk(gclk));
	jdff dff_B_az7TCeYd7_2(.din(w_dff_B_7fuvmvCx4_2),.dout(w_dff_B_az7TCeYd7_2),.clk(gclk));
	jdff dff_B_7RL1TIQc5_2(.din(w_dff_B_az7TCeYd7_2),.dout(w_dff_B_7RL1TIQc5_2),.clk(gclk));
	jdff dff_B_SVdhd0Dc8_2(.din(w_dff_B_7RL1TIQc5_2),.dout(w_dff_B_SVdhd0Dc8_2),.clk(gclk));
	jdff dff_B_0MyRwGPc8_2(.din(w_dff_B_SVdhd0Dc8_2),.dout(w_dff_B_0MyRwGPc8_2),.clk(gclk));
	jdff dff_B_D9yHKpXV5_2(.din(w_dff_B_0MyRwGPc8_2),.dout(w_dff_B_D9yHKpXV5_2),.clk(gclk));
	jdff dff_B_np3gfNno3_2(.din(w_dff_B_D9yHKpXV5_2),.dout(w_dff_B_np3gfNno3_2),.clk(gclk));
	jdff dff_B_XoQwXwxj0_2(.din(w_dff_B_np3gfNno3_2),.dout(w_dff_B_XoQwXwxj0_2),.clk(gclk));
	jdff dff_B_BAQRRF1l2_2(.din(w_dff_B_XoQwXwxj0_2),.dout(w_dff_B_BAQRRF1l2_2),.clk(gclk));
	jdff dff_B_5VtNxWne5_2(.din(w_dff_B_BAQRRF1l2_2),.dout(w_dff_B_5VtNxWne5_2),.clk(gclk));
	jdff dff_B_XBhqH1475_2(.din(w_dff_B_5VtNxWne5_2),.dout(w_dff_B_XBhqH1475_2),.clk(gclk));
	jdff dff_B_fyrZXCvG0_2(.din(w_dff_B_XBhqH1475_2),.dout(w_dff_B_fyrZXCvG0_2),.clk(gclk));
	jdff dff_A_P4E9OfrU2_0(.dout(w_G27gat_0[0]),.din(w_dff_A_P4E9OfrU2_0),.clk(gclk));
	jdff dff_A_NfnO9f7r4_0(.dout(w_dff_A_P4E9OfrU2_0),.din(w_dff_A_NfnO9f7r4_0),.clk(gclk));
	jdff dff_A_oF9666GH5_0(.dout(w_dff_A_NfnO9f7r4_0),.din(w_dff_A_oF9666GH5_0),.clk(gclk));
	jdff dff_A_TMJ6cU6F7_0(.dout(w_dff_A_oF9666GH5_0),.din(w_dff_A_TMJ6cU6F7_0),.clk(gclk));
	jdff dff_A_q40O1sGG4_0(.dout(w_dff_A_TMJ6cU6F7_0),.din(w_dff_A_q40O1sGG4_0),.clk(gclk));
	jdff dff_A_KdSzsY7L4_0(.dout(w_dff_A_q40O1sGG4_0),.din(w_dff_A_KdSzsY7L4_0),.clk(gclk));
	jdff dff_A_TDSvuKZa7_0(.dout(w_dff_A_KdSzsY7L4_0),.din(w_dff_A_TDSvuKZa7_0),.clk(gclk));
	jdff dff_A_Z0zALdGJ2_0(.dout(w_dff_A_TDSvuKZa7_0),.din(w_dff_A_Z0zALdGJ2_0),.clk(gclk));
	jdff dff_A_14tCVaq02_0(.dout(w_dff_A_Z0zALdGJ2_0),.din(w_dff_A_14tCVaq02_0),.clk(gclk));
	jdff dff_A_9ASsQCif4_0(.dout(w_dff_A_14tCVaq02_0),.din(w_dff_A_9ASsQCif4_0),.clk(gclk));
	jdff dff_A_Yb4EtMYG4_0(.dout(w_dff_A_9ASsQCif4_0),.din(w_dff_A_Yb4EtMYG4_0),.clk(gclk));
	jdff dff_A_AOjEDhQx8_0(.dout(w_dff_A_Yb4EtMYG4_0),.din(w_dff_A_AOjEDhQx8_0),.clk(gclk));
	jdff dff_A_NeiQxvBq5_0(.dout(w_dff_A_AOjEDhQx8_0),.din(w_dff_A_NeiQxvBq5_0),.clk(gclk));
	jdff dff_A_O0PhjXJJ1_0(.dout(w_dff_A_NeiQxvBq5_0),.din(w_dff_A_O0PhjXJJ1_0),.clk(gclk));
	jdff dff_A_3DkbUKqV4_0(.dout(w_n197_0[0]),.din(w_dff_A_3DkbUKqV4_0),.clk(gclk));
	jdff dff_A_q4PeoTyl5_0(.dout(w_dff_A_3DkbUKqV4_0),.din(w_dff_A_q4PeoTyl5_0),.clk(gclk));
	jdff dff_A_32hI6N2n9_0(.dout(w_dff_A_q4PeoTyl5_0),.din(w_dff_A_32hI6N2n9_0),.clk(gclk));
	jdff dff_A_IYUO0ecr1_0(.dout(w_dff_A_32hI6N2n9_0),.din(w_dff_A_IYUO0ecr1_0),.clk(gclk));
	jdff dff_A_11nRX98N3_0(.dout(w_dff_A_IYUO0ecr1_0),.din(w_dff_A_11nRX98N3_0),.clk(gclk));
	jdff dff_A_T30xqLpp4_0(.dout(w_dff_A_11nRX98N3_0),.din(w_dff_A_T30xqLpp4_0),.clk(gclk));
	jdff dff_A_2gpDt1rw1_1(.dout(w_n193_0[1]),.din(w_dff_A_2gpDt1rw1_1),.clk(gclk));
	jdff dff_A_z4WWpocZ0_1(.dout(w_dff_A_2gpDt1rw1_1),.din(w_dff_A_z4WWpocZ0_1),.clk(gclk));
	jdff dff_A_BiEMJDwr2_1(.dout(w_dff_A_z4WWpocZ0_1),.din(w_dff_A_BiEMJDwr2_1),.clk(gclk));
	jdff dff_A_x3s1wrdr0_1(.dout(w_dff_A_BiEMJDwr2_1),.din(w_dff_A_x3s1wrdr0_1),.clk(gclk));
	jdff dff_A_CUXDsklJ4_1(.dout(w_dff_A_x3s1wrdr0_1),.din(w_dff_A_CUXDsklJ4_1),.clk(gclk));
	jdff dff_A_9Jbz5w6N9_1(.dout(w_dff_A_CUXDsklJ4_1),.din(w_dff_A_9Jbz5w6N9_1),.clk(gclk));
	jdff dff_A_s6t7iNYI6_1(.dout(w_dff_A_9Jbz5w6N9_1),.din(w_dff_A_s6t7iNYI6_1),.clk(gclk));
	jdff dff_B_4QZ46xG08_0(.din(n192),.dout(w_dff_B_4QZ46xG08_0),.clk(gclk));
	jdff dff_B_b6nSR68a2_0(.din(w_dff_B_4QZ46xG08_0),.dout(w_dff_B_b6nSR68a2_0),.clk(gclk));
	jdff dff_B_NJHj4LJQ3_0(.din(w_dff_B_b6nSR68a2_0),.dout(w_dff_B_NJHj4LJQ3_0),.clk(gclk));
	jdff dff_B_cylbLnVE1_0(.din(w_dff_B_NJHj4LJQ3_0),.dout(w_dff_B_cylbLnVE1_0),.clk(gclk));
	jdff dff_B_0xlbnkxf7_0(.din(w_dff_B_cylbLnVE1_0),.dout(w_dff_B_0xlbnkxf7_0),.clk(gclk));
	jdff dff_A_kkuwY2iN0_0(.dout(w_n191_0[0]),.din(w_dff_A_kkuwY2iN0_0),.clk(gclk));
	jdff dff_A_xEo5DSXc0_0(.dout(w_dff_A_kkuwY2iN0_0),.din(w_dff_A_xEo5DSXc0_0),.clk(gclk));
	jdff dff_A_JxBinVoZ4_0(.dout(w_dff_A_xEo5DSXc0_0),.din(w_dff_A_JxBinVoZ4_0),.clk(gclk));
	jdff dff_A_nUTgCvt80_0(.dout(w_dff_A_JxBinVoZ4_0),.din(w_dff_A_nUTgCvt80_0),.clk(gclk));
	jdff dff_A_r7iu4eT31_0(.dout(w_dff_A_nUTgCvt80_0),.din(w_dff_A_r7iu4eT31_0),.clk(gclk));
	jdff dff_A_PZtx4D5a9_0(.dout(w_dff_A_r7iu4eT31_0),.din(w_dff_A_PZtx4D5a9_0),.clk(gclk));
	jdff dff_A_D1zSyuGG8_0(.dout(w_dff_A_PZtx4D5a9_0),.din(w_dff_A_D1zSyuGG8_0),.clk(gclk));
	jdff dff_A_4WhcggbI7_0(.dout(w_dff_A_D1zSyuGG8_0),.din(w_dff_A_4WhcggbI7_0),.clk(gclk));
	jdff dff_A_6VDJmKIe8_0(.dout(w_dff_A_4WhcggbI7_0),.din(w_dff_A_6VDJmKIe8_0),.clk(gclk));
	jdff dff_A_AGZU92X91_0(.dout(w_dff_A_6VDJmKIe8_0),.din(w_dff_A_AGZU92X91_0),.clk(gclk));
	jdff dff_A_7EfEMMAw2_0(.dout(w_dff_A_AGZU92X91_0),.din(w_dff_A_7EfEMMAw2_0),.clk(gclk));
	jdff dff_A_gn9Dwxgk1_0(.dout(w_dff_A_7EfEMMAw2_0),.din(w_dff_A_gn9Dwxgk1_0),.clk(gclk));
	jdff dff_A_nbLpy6kM5_0(.dout(w_dff_A_gn9Dwxgk1_0),.din(w_dff_A_nbLpy6kM5_0),.clk(gclk));
	jdff dff_A_JYv7xi7H3_0(.dout(w_dff_A_nbLpy6kM5_0),.din(w_dff_A_JYv7xi7H3_0),.clk(gclk));
	jdff dff_A_Y4jSUqGe3_0(.dout(w_dff_A_JYv7xi7H3_0),.din(w_dff_A_Y4jSUqGe3_0),.clk(gclk));
	jdff dff_A_1xfANVUj8_0(.dout(w_dff_A_Y4jSUqGe3_0),.din(w_dff_A_1xfANVUj8_0),.clk(gclk));
	jdff dff_A_wYFRCQu26_0(.dout(w_dff_A_1xfANVUj8_0),.din(w_dff_A_wYFRCQu26_0),.clk(gclk));
	jdff dff_A_CHVy6Qct6_0(.dout(w_dff_A_wYFRCQu26_0),.din(w_dff_A_CHVy6Qct6_0),.clk(gclk));
	jdff dff_A_NztlICNx4_0(.dout(w_dff_A_CHVy6Qct6_0),.din(w_dff_A_NztlICNx4_0),.clk(gclk));
	jdff dff_A_K70pXfwm2_0(.dout(w_G53gat_0[0]),.din(w_dff_A_K70pXfwm2_0),.clk(gclk));
	jdff dff_A_rhgUzpww6_0(.dout(w_dff_A_K70pXfwm2_0),.din(w_dff_A_rhgUzpww6_0),.clk(gclk));
	jdff dff_A_lPudnZzQ4_0(.dout(w_dff_A_rhgUzpww6_0),.din(w_dff_A_lPudnZzQ4_0),.clk(gclk));
	jdff dff_A_Tqzg5ZiU4_0(.dout(w_dff_A_lPudnZzQ4_0),.din(w_dff_A_Tqzg5ZiU4_0),.clk(gclk));
	jdff dff_A_is7xcMgr9_0(.dout(w_dff_A_Tqzg5ZiU4_0),.din(w_dff_A_is7xcMgr9_0),.clk(gclk));
	jdff dff_A_ZSidA31H8_0(.dout(w_dff_A_is7xcMgr9_0),.din(w_dff_A_ZSidA31H8_0),.clk(gclk));
	jdff dff_A_AdleOg1T4_0(.dout(w_dff_A_ZSidA31H8_0),.din(w_dff_A_AdleOg1T4_0),.clk(gclk));
	jdff dff_A_2kr83mvm7_0(.dout(w_dff_A_AdleOg1T4_0),.din(w_dff_A_2kr83mvm7_0),.clk(gclk));
	jdff dff_A_7YB8gEZS0_0(.dout(w_dff_A_2kr83mvm7_0),.din(w_dff_A_7YB8gEZS0_0),.clk(gclk));
	jdff dff_A_72YPSi479_0(.dout(w_dff_A_7YB8gEZS0_0),.din(w_dff_A_72YPSi479_0),.clk(gclk));
	jdff dff_A_g7Y78fgg7_0(.dout(w_dff_A_72YPSi479_0),.din(w_dff_A_g7Y78fgg7_0),.clk(gclk));
	jdff dff_A_ijzhXmIl2_0(.dout(w_dff_A_g7Y78fgg7_0),.din(w_dff_A_ijzhXmIl2_0),.clk(gclk));
	jdff dff_A_5mq645bi0_0(.dout(w_dff_A_ijzhXmIl2_0),.din(w_dff_A_5mq645bi0_0),.clk(gclk));
	jdff dff_A_vOdb2YxJ8_0(.dout(w_dff_A_5mq645bi0_0),.din(w_dff_A_vOdb2YxJ8_0),.clk(gclk));
	jdff dff_A_Rp8YjN2A0_0(.dout(w_dff_A_vOdb2YxJ8_0),.din(w_dff_A_Rp8YjN2A0_0),.clk(gclk));
	jdff dff_A_wXz8MI1r6_0(.dout(w_dff_A_Rp8YjN2A0_0),.din(w_dff_A_wXz8MI1r6_0),.clk(gclk));
	jdff dff_A_iPjsRmrz4_0(.dout(w_dff_A_wXz8MI1r6_0),.din(w_dff_A_iPjsRmrz4_0),.clk(gclk));
	jdff dff_A_Qiowc9UD7_0(.dout(w_dff_A_iPjsRmrz4_0),.din(w_dff_A_Qiowc9UD7_0),.clk(gclk));
	jdff dff_A_eS2VW7jv4_0(.dout(w_dff_A_Qiowc9UD7_0),.din(w_dff_A_eS2VW7jv4_0),.clk(gclk));
	jdff dff_A_OYC4wMHD3_0(.dout(w_dff_A_eS2VW7jv4_0),.din(w_dff_A_OYC4wMHD3_0),.clk(gclk));
	jdff dff_A_rvv8PztO5_0(.dout(w_n184_0[0]),.din(w_dff_A_rvv8PztO5_0),.clk(gclk));
	jdff dff_A_39boRS979_0(.dout(w_dff_A_rvv8PztO5_0),.din(w_dff_A_39boRS979_0),.clk(gclk));
	jdff dff_A_NvpKZUwL4_0(.dout(w_dff_A_39boRS979_0),.din(w_dff_A_NvpKZUwL4_0),.clk(gclk));
	jdff dff_A_ySeg3elV5_0(.dout(w_dff_A_NvpKZUwL4_0),.din(w_dff_A_ySeg3elV5_0),.clk(gclk));
	jdff dff_A_CfgtonVu2_0(.dout(w_dff_A_ySeg3elV5_0),.din(w_dff_A_CfgtonVu2_0),.clk(gclk));
	jdff dff_A_ajlO7iq04_0(.dout(w_dff_A_CfgtonVu2_0),.din(w_dff_A_ajlO7iq04_0),.clk(gclk));
	jdff dff_B_TULCKkIv7_1(.din(n167),.dout(w_dff_B_TULCKkIv7_1),.clk(gclk));
	jdff dff_A_lOfZMnf54_0(.dout(w_n177_0[0]),.din(w_dff_A_lOfZMnf54_0),.clk(gclk));
	jdff dff_A_n6hXZ9SH3_0(.dout(w_dff_A_lOfZMnf54_0),.din(w_dff_A_n6hXZ9SH3_0),.clk(gclk));
	jdff dff_A_jUYZU3kF9_0(.dout(w_dff_A_n6hXZ9SH3_0),.din(w_dff_A_jUYZU3kF9_0),.clk(gclk));
	jdff dff_A_gevSWNzF0_0(.dout(w_dff_A_jUYZU3kF9_0),.din(w_dff_A_gevSWNzF0_0),.clk(gclk));
	jdff dff_A_6BGROkuE9_0(.dout(w_dff_A_gevSWNzF0_0),.din(w_dff_A_6BGROkuE9_0),.clk(gclk));
	jdff dff_A_eV97XeUj9_0(.dout(w_dff_A_6BGROkuE9_0),.din(w_dff_A_eV97XeUj9_0),.clk(gclk));
	jdff dff_A_Kf3ddpAR8_0(.dout(w_n174_0[0]),.din(w_dff_A_Kf3ddpAR8_0),.clk(gclk));
	jdff dff_A_AC3V1HOO4_0(.dout(w_dff_A_Kf3ddpAR8_0),.din(w_dff_A_AC3V1HOO4_0),.clk(gclk));
	jdff dff_A_WE7qvhvl3_0(.dout(w_dff_A_AC3V1HOO4_0),.din(w_dff_A_WE7qvhvl3_0),.clk(gclk));
	jdff dff_A_VMbfIxYJ9_0(.dout(w_dff_A_WE7qvhvl3_0),.din(w_dff_A_VMbfIxYJ9_0),.clk(gclk));
	jdff dff_A_Iyn24Ir93_0(.dout(w_dff_A_VMbfIxYJ9_0),.din(w_dff_A_Iyn24Ir93_0),.clk(gclk));
	jdff dff_A_1NHobVf29_0(.dout(w_dff_A_Iyn24Ir93_0),.din(w_dff_A_1NHobVf29_0),.clk(gclk));
	jdff dff_B_OOZQruHx0_1(.din(n172),.dout(w_dff_B_OOZQruHx0_1),.clk(gclk));
	jdff dff_B_c5c18Uis1_1(.din(w_dff_B_OOZQruHx0_1),.dout(w_dff_B_c5c18Uis1_1),.clk(gclk));
	jdff dff_B_PVqFOUhM9_1(.din(w_dff_B_c5c18Uis1_1),.dout(w_dff_B_PVqFOUhM9_1),.clk(gclk));
	jdff dff_B_sgkt7iPm9_1(.din(w_dff_B_PVqFOUhM9_1),.dout(w_dff_B_sgkt7iPm9_1),.clk(gclk));
	jdff dff_B_5SkpzC2A4_1(.din(w_dff_B_sgkt7iPm9_1),.dout(w_dff_B_5SkpzC2A4_1),.clk(gclk));
	jdff dff_B_vuzsV2FC6_1(.din(w_dff_B_5SkpzC2A4_1),.dout(w_dff_B_vuzsV2FC6_1),.clk(gclk));
	jdff dff_A_nC9RLLDY4_0(.dout(w_n170_0[0]),.din(w_dff_A_nC9RLLDY4_0),.clk(gclk));
	jdff dff_A_fSU0j8Yn2_0(.dout(w_dff_A_nC9RLLDY4_0),.din(w_dff_A_fSU0j8Yn2_0),.clk(gclk));
	jdff dff_A_5UjwFNuN8_0(.dout(w_dff_A_fSU0j8Yn2_0),.din(w_dff_A_5UjwFNuN8_0),.clk(gclk));
	jdff dff_A_I0B4DkU05_0(.dout(w_dff_A_5UjwFNuN8_0),.din(w_dff_A_I0B4DkU05_0),.clk(gclk));
	jdff dff_B_DacFIcBk5_2(.din(n170),.dout(w_dff_B_DacFIcBk5_2),.clk(gclk));
	jdff dff_B_i2Sflq2H1_0(.din(n169),.dout(w_dff_B_i2Sflq2H1_0),.clk(gclk));
	jdff dff_B_SlHUmUsE1_0(.din(w_dff_B_i2Sflq2H1_0),.dout(w_dff_B_SlHUmUsE1_0),.clk(gclk));
	jdff dff_B_nQ6YaW0S4_0(.din(w_dff_B_SlHUmUsE1_0),.dout(w_dff_B_nQ6YaW0S4_0),.clk(gclk));
	jdff dff_B_i8ozyrsk5_0(.din(w_dff_B_nQ6YaW0S4_0),.dout(w_dff_B_i8ozyrsk5_0),.clk(gclk));
	jdff dff_A_mIghtVWN7_0(.dout(w_n164_0[0]),.din(w_dff_A_mIghtVWN7_0),.clk(gclk));
	jdff dff_A_U6hHS9oy6_0(.dout(w_dff_A_mIghtVWN7_0),.din(w_dff_A_U6hHS9oy6_0),.clk(gclk));
	jdff dff_A_3A1so0WA4_0(.dout(w_dff_A_U6hHS9oy6_0),.din(w_dff_A_3A1so0WA4_0),.clk(gclk));
	jdff dff_A_M2mwOCZz0_0(.dout(w_dff_A_3A1so0WA4_0),.din(w_dff_A_M2mwOCZz0_0),.clk(gclk));
	jdff dff_A_2TjCq7Hh6_0(.dout(w_dff_A_M2mwOCZz0_0),.din(w_dff_A_2TjCq7Hh6_0),.clk(gclk));
	jdff dff_A_P8mWUwpS3_0(.dout(w_dff_A_2TjCq7Hh6_0),.din(w_dff_A_P8mWUwpS3_0),.clk(gclk));
	jdff dff_A_X4qN0ZtE2_0(.dout(w_n159_0[0]),.din(w_dff_A_X4qN0ZtE2_0),.clk(gclk));
	jdff dff_A_ZnHftyNV4_0(.dout(w_dff_A_X4qN0ZtE2_0),.din(w_dff_A_ZnHftyNV4_0),.clk(gclk));
	jdff dff_A_9cQavNd13_0(.dout(w_dff_A_ZnHftyNV4_0),.din(w_dff_A_9cQavNd13_0),.clk(gclk));
	jdff dff_A_pbaOLV8f9_0(.dout(w_dff_A_9cQavNd13_0),.din(w_dff_A_pbaOLV8f9_0),.clk(gclk));
	jdff dff_A_Ar5obENu8_0(.dout(w_dff_A_pbaOLV8f9_0),.din(w_dff_A_Ar5obENu8_0),.clk(gclk));
	jdff dff_A_3fWF9Vay3_0(.dout(w_dff_A_Ar5obENu8_0),.din(w_dff_A_3fWF9Vay3_0),.clk(gclk));
	jdff dff_A_X9fM55LS2_0(.dout(w_n156_0[0]),.din(w_dff_A_X9fM55LS2_0),.clk(gclk));
	jdff dff_A_5Q738wrw6_0(.dout(w_dff_A_X9fM55LS2_0),.din(w_dff_A_5Q738wrw6_0),.clk(gclk));
	jdff dff_A_DATfAEHS4_0(.dout(w_dff_A_5Q738wrw6_0),.din(w_dff_A_DATfAEHS4_0),.clk(gclk));
	jdff dff_A_gVjaJtsn2_0(.dout(w_dff_A_DATfAEHS4_0),.din(w_dff_A_gVjaJtsn2_0),.clk(gclk));
	jdff dff_A_bRsrjABE0_0(.dout(w_dff_A_gVjaJtsn2_0),.din(w_dff_A_bRsrjABE0_0),.clk(gclk));
	jdff dff_A_ZOGdPGs42_0(.dout(w_dff_A_bRsrjABE0_0),.din(w_dff_A_ZOGdPGs42_0),.clk(gclk));
	jdff dff_A_upZOs5PZ5_0(.dout(w_n154_0[0]),.din(w_dff_A_upZOs5PZ5_0),.clk(gclk));
	jdff dff_A_BdUgGSAh2_0(.dout(w_dff_A_upZOs5PZ5_0),.din(w_dff_A_BdUgGSAh2_0),.clk(gclk));
	jdff dff_A_Nc2x7Jwl2_0(.dout(w_dff_A_BdUgGSAh2_0),.din(w_dff_A_Nc2x7Jwl2_0),.clk(gclk));
	jdff dff_A_1mU1ZLEm8_0(.dout(w_dff_A_Nc2x7Jwl2_0),.din(w_dff_A_1mU1ZLEm8_0),.clk(gclk));
	jdff dff_A_nl7IyFXG9_0(.dout(w_dff_A_1mU1ZLEm8_0),.din(w_dff_A_nl7IyFXG9_0),.clk(gclk));
	jdff dff_B_ih3E6Wpi6_2(.din(n154),.dout(w_dff_B_ih3E6Wpi6_2),.clk(gclk));
	jdff dff_B_D617FD3g6_2(.din(w_dff_B_ih3E6Wpi6_2),.dout(w_dff_B_D617FD3g6_2),.clk(gclk));
	jdff dff_B_TAsBmQD71_2(.din(w_dff_B_D617FD3g6_2),.dout(w_dff_B_TAsBmQD71_2),.clk(gclk));
	jdff dff_B_m9OscV3G6_2(.din(w_dff_B_TAsBmQD71_2),.dout(w_dff_B_m9OscV3G6_2),.clk(gclk));
	jdff dff_B_0C65iaNx5_2(.din(w_dff_B_m9OscV3G6_2),.dout(w_dff_B_0C65iaNx5_2),.clk(gclk));
	jdff dff_B_f4x8NmUE9_2(.din(w_dff_B_0C65iaNx5_2),.dout(w_dff_B_f4x8NmUE9_2),.clk(gclk));
	jdff dff_B_6g7kN7jm8_2(.din(w_dff_B_f4x8NmUE9_2),.dout(w_dff_B_6g7kN7jm8_2),.clk(gclk));
	jdff dff_B_MybpwxhO4_2(.din(w_dff_B_6g7kN7jm8_2),.dout(w_dff_B_MybpwxhO4_2),.clk(gclk));
	jdff dff_B_Rv3whGh50_2(.din(w_dff_B_MybpwxhO4_2),.dout(w_dff_B_Rv3whGh50_2),.clk(gclk));
	jdff dff_B_ujhZzmE93_2(.din(w_dff_B_Rv3whGh50_2),.dout(w_dff_B_ujhZzmE93_2),.clk(gclk));
	jdff dff_B_p9htagI23_2(.din(w_dff_B_ujhZzmE93_2),.dout(w_dff_B_p9htagI23_2),.clk(gclk));
	jdff dff_B_7tnf8wmb0_2(.din(w_dff_B_p9htagI23_2),.dout(w_dff_B_7tnf8wmb0_2),.clk(gclk));
	jdff dff_B_IR8Bvya77_2(.din(w_dff_B_7tnf8wmb0_2),.dout(w_dff_B_IR8Bvya77_2),.clk(gclk));
	jdff dff_B_ynVHqGdP0_2(.din(w_dff_B_IR8Bvya77_2),.dout(w_dff_B_ynVHqGdP0_2),.clk(gclk));
	jdff dff_A_3OPq8lC90_0(.dout(w_G79gat_0[0]),.din(w_dff_A_3OPq8lC90_0),.clk(gclk));
	jdff dff_A_qLM8c9x33_0(.dout(w_dff_A_3OPq8lC90_0),.din(w_dff_A_qLM8c9x33_0),.clk(gclk));
	jdff dff_A_K8uVWCHg2_0(.dout(w_dff_A_qLM8c9x33_0),.din(w_dff_A_K8uVWCHg2_0),.clk(gclk));
	jdff dff_A_wQUjB8Sy9_0(.dout(w_dff_A_K8uVWCHg2_0),.din(w_dff_A_wQUjB8Sy9_0),.clk(gclk));
	jdff dff_A_dLf5Wvxq3_0(.dout(w_dff_A_wQUjB8Sy9_0),.din(w_dff_A_dLf5Wvxq3_0),.clk(gclk));
	jdff dff_A_3QiR7ewA2_0(.dout(w_dff_A_dLf5Wvxq3_0),.din(w_dff_A_3QiR7ewA2_0),.clk(gclk));
	jdff dff_A_iWa6xviI8_0(.dout(w_dff_A_3QiR7ewA2_0),.din(w_dff_A_iWa6xviI8_0),.clk(gclk));
	jdff dff_A_eklnG9MQ6_0(.dout(w_dff_A_iWa6xviI8_0),.din(w_dff_A_eklnG9MQ6_0),.clk(gclk));
	jdff dff_A_GBFYKOkz5_0(.dout(w_dff_A_eklnG9MQ6_0),.din(w_dff_A_GBFYKOkz5_0),.clk(gclk));
	jdff dff_A_c63E0tea8_0(.dout(w_dff_A_GBFYKOkz5_0),.din(w_dff_A_c63E0tea8_0),.clk(gclk));
	jdff dff_A_qMmAYXyr9_0(.dout(w_dff_A_c63E0tea8_0),.din(w_dff_A_qMmAYXyr9_0),.clk(gclk));
	jdff dff_A_qahQb5Qc7_0(.dout(w_dff_A_qMmAYXyr9_0),.din(w_dff_A_qahQb5Qc7_0),.clk(gclk));
	jdff dff_A_FT22x3K41_0(.dout(w_dff_A_qahQb5Qc7_0),.din(w_dff_A_FT22x3K41_0),.clk(gclk));
	jdff dff_A_FjkyvDqN9_0(.dout(w_dff_A_FT22x3K41_0),.din(w_dff_A_FjkyvDqN9_0),.clk(gclk));
	jdff dff_A_IcPR62ao3_0(.dout(w_dff_A_FjkyvDqN9_0),.din(w_dff_A_IcPR62ao3_0),.clk(gclk));
	jdff dff_A_dMFpHtVm4_1(.dout(w_n151_0[1]),.din(w_dff_A_dMFpHtVm4_1),.clk(gclk));
	jdff dff_A_7bWL3VEH3_1(.dout(w_dff_A_dMFpHtVm4_1),.din(w_dff_A_7bWL3VEH3_1),.clk(gclk));
	jdff dff_A_3vDhBz6t5_1(.dout(w_dff_A_7bWL3VEH3_1),.din(w_dff_A_3vDhBz6t5_1),.clk(gclk));
	jdff dff_A_d05E4w361_1(.dout(w_dff_A_3vDhBz6t5_1),.din(w_dff_A_d05E4w361_1),.clk(gclk));
	jdff dff_A_2wwBRVl54_1(.dout(w_dff_A_d05E4w361_1),.din(w_dff_A_2wwBRVl54_1),.clk(gclk));
	jdff dff_A_iswuUbvY4_1(.dout(w_dff_A_2wwBRVl54_1),.din(w_dff_A_iswuUbvY4_1),.clk(gclk));
	jdff dff_A_wSS7Uavd7_0(.dout(w_n150_0[0]),.din(w_dff_A_wSS7Uavd7_0),.clk(gclk));
	jdff dff_A_ahDzLQV77_0(.dout(w_dff_A_wSS7Uavd7_0),.din(w_dff_A_ahDzLQV77_0),.clk(gclk));
	jdff dff_A_tyBqzzah5_0(.dout(w_dff_A_ahDzLQV77_0),.din(w_dff_A_tyBqzzah5_0),.clk(gclk));
	jdff dff_A_lkFuCNfX4_0(.dout(w_dff_A_tyBqzzah5_0),.din(w_dff_A_lkFuCNfX4_0),.clk(gclk));
	jdff dff_A_YbFSinoe7_0(.dout(w_dff_A_lkFuCNfX4_0),.din(w_dff_A_YbFSinoe7_0),.clk(gclk));
	jdff dff_A_t3Hryi672_0(.dout(w_dff_A_YbFSinoe7_0),.din(w_dff_A_t3Hryi672_0),.clk(gclk));
	jdff dff_A_yj0eJcbk9_0(.dout(w_dff_A_t3Hryi672_0),.din(w_dff_A_yj0eJcbk9_0),.clk(gclk));
	jdff dff_A_iS7P584Y7_0(.dout(w_dff_A_yj0eJcbk9_0),.din(w_dff_A_iS7P584Y7_0),.clk(gclk));
	jdff dff_A_R5mgsJEh5_0(.dout(w_dff_A_iS7P584Y7_0),.din(w_dff_A_R5mgsJEh5_0),.clk(gclk));
	jdff dff_A_KNtmxcGp2_0(.dout(w_dff_A_R5mgsJEh5_0),.din(w_dff_A_KNtmxcGp2_0),.clk(gclk));
	jdff dff_A_FP4D0iMU9_0(.dout(w_dff_A_KNtmxcGp2_0),.din(w_dff_A_FP4D0iMU9_0),.clk(gclk));
	jdff dff_A_b787DLJQ7_0(.dout(w_dff_A_FP4D0iMU9_0),.din(w_dff_A_b787DLJQ7_0),.clk(gclk));
	jdff dff_B_3suSYngp4_2(.din(n150),.dout(w_dff_B_3suSYngp4_2),.clk(gclk));
	jdff dff_B_ryLnhs7O7_2(.din(w_dff_B_3suSYngp4_2),.dout(w_dff_B_ryLnhs7O7_2),.clk(gclk));
	jdff dff_B_nck2wWvV9_2(.din(w_dff_B_ryLnhs7O7_2),.dout(w_dff_B_nck2wWvV9_2),.clk(gclk));
	jdff dff_B_SgbJxtLR8_2(.din(w_dff_B_nck2wWvV9_2),.dout(w_dff_B_SgbJxtLR8_2),.clk(gclk));
	jdff dff_B_1bgoMqsc2_2(.din(w_dff_B_SgbJxtLR8_2),.dout(w_dff_B_1bgoMqsc2_2),.clk(gclk));
	jdff dff_B_4737DIKd2_2(.din(w_dff_B_1bgoMqsc2_2),.dout(w_dff_B_4737DIKd2_2),.clk(gclk));
	jdff dff_B_oJ0khUTh6_2(.din(w_dff_B_4737DIKd2_2),.dout(w_dff_B_oJ0khUTh6_2),.clk(gclk));
	jdff dff_A_CBhlU5Vi0_0(.dout(w_G66gat_0[0]),.din(w_dff_A_CBhlU5Vi0_0),.clk(gclk));
	jdff dff_A_Rhp8TIeZ8_0(.dout(w_dff_A_CBhlU5Vi0_0),.din(w_dff_A_Rhp8TIeZ8_0),.clk(gclk));
	jdff dff_A_hqIttyzW7_0(.dout(w_dff_A_Rhp8TIeZ8_0),.din(w_dff_A_hqIttyzW7_0),.clk(gclk));
	jdff dff_A_ggH5p7q20_0(.dout(w_dff_A_hqIttyzW7_0),.din(w_dff_A_ggH5p7q20_0),.clk(gclk));
	jdff dff_A_4LvNKKTI7_0(.dout(w_dff_A_ggH5p7q20_0),.din(w_dff_A_4LvNKKTI7_0),.clk(gclk));
	jdff dff_A_2Aj9k8949_0(.dout(w_dff_A_4LvNKKTI7_0),.din(w_dff_A_2Aj9k8949_0),.clk(gclk));
	jdff dff_A_WvQViioJ4_0(.dout(w_dff_A_2Aj9k8949_0),.din(w_dff_A_WvQViioJ4_0),.clk(gclk));
	jdff dff_A_36KIvm9k9_0(.dout(w_dff_A_WvQViioJ4_0),.din(w_dff_A_36KIvm9k9_0),.clk(gclk));
	jdff dff_A_rrQ8oGqq8_0(.dout(w_dff_A_36KIvm9k9_0),.din(w_dff_A_rrQ8oGqq8_0),.clk(gclk));
	jdff dff_A_grHjRU1c6_0(.dout(w_dff_A_rrQ8oGqq8_0),.din(w_dff_A_grHjRU1c6_0),.clk(gclk));
	jdff dff_A_38u79YLn2_0(.dout(w_dff_A_grHjRU1c6_0),.din(w_dff_A_38u79YLn2_0),.clk(gclk));
	jdff dff_A_Ip7mFw6K8_0(.dout(w_dff_A_38u79YLn2_0),.din(w_dff_A_Ip7mFw6K8_0),.clk(gclk));
	jdff dff_A_ylJ6p2Hj3_0(.dout(w_dff_A_Ip7mFw6K8_0),.din(w_dff_A_ylJ6p2Hj3_0),.clk(gclk));
	jdff dff_A_lpLg8iFg3_0(.dout(w_dff_A_ylJ6p2Hj3_0),.din(w_dff_A_lpLg8iFg3_0),.clk(gclk));
	jdff dff_A_tbpptluP1_0(.dout(w_dff_A_lpLg8iFg3_0),.din(w_dff_A_tbpptluP1_0),.clk(gclk));
	jdff dff_A_MxJo78O71_0(.dout(w_dff_A_tbpptluP1_0),.din(w_dff_A_MxJo78O71_0),.clk(gclk));
	jdff dff_A_LPShTF3E9_0(.dout(w_dff_A_MxJo78O71_0),.din(w_dff_A_LPShTF3E9_0),.clk(gclk));
	jdff dff_A_YLc1MDH15_0(.dout(w_dff_A_LPShTF3E9_0),.din(w_dff_A_YLc1MDH15_0),.clk(gclk));
	jdff dff_A_TfSFkQUk7_0(.dout(w_dff_A_YLc1MDH15_0),.din(w_dff_A_TfSFkQUk7_0),.clk(gclk));
	jdff dff_A_4L7SPVuI9_0(.dout(w_dff_A_TfSFkQUk7_0),.din(w_dff_A_4L7SPVuI9_0),.clk(gclk));
	jdff dff_A_qKQ1EjVd3_1(.dout(w_n146_0[1]),.din(w_dff_A_qKQ1EjVd3_1),.clk(gclk));
	jdff dff_A_CWr6yg7X2_1(.dout(w_dff_A_qKQ1EjVd3_1),.din(w_dff_A_CWr6yg7X2_1),.clk(gclk));
	jdff dff_A_OPhQx6q53_1(.dout(w_dff_A_CWr6yg7X2_1),.din(w_dff_A_OPhQx6q53_1),.clk(gclk));
	jdff dff_A_YDMdgSf06_1(.dout(w_dff_A_OPhQx6q53_1),.din(w_dff_A_YDMdgSf06_1),.clk(gclk));
	jdff dff_A_NHH8y1P76_0(.dout(w_n145_0[0]),.din(w_dff_A_NHH8y1P76_0),.clk(gclk));
	jdff dff_A_dy9ywEpf3_0(.dout(w_dff_A_NHH8y1P76_0),.din(w_dff_A_dy9ywEpf3_0),.clk(gclk));
	jdff dff_A_4Yn67P8E2_0(.dout(w_dff_A_dy9ywEpf3_0),.din(w_dff_A_4Yn67P8E2_0),.clk(gclk));
	jdff dff_A_36qhM1LE6_0(.dout(w_dff_A_4Yn67P8E2_0),.din(w_dff_A_36qhM1LE6_0),.clk(gclk));
	jdff dff_A_rqGOiAIo8_0(.dout(w_dff_A_36qhM1LE6_0),.din(w_dff_A_rqGOiAIo8_0),.clk(gclk));
	jdff dff_A_jggaCk2R5_0(.dout(w_dff_A_rqGOiAIo8_0),.din(w_dff_A_jggaCk2R5_0),.clk(gclk));
	jdff dff_A_TH3VM6Wq8_0(.dout(w_n142_0[0]),.din(w_dff_A_TH3VM6Wq8_0),.clk(gclk));
	jdff dff_B_L8xAIm631_1(.din(n112),.dout(w_dff_B_L8xAIm631_1),.clk(gclk));
	jdff dff_B_5HVIxTto7_1(.din(n116),.dout(w_dff_B_5HVIxTto7_1),.clk(gclk));
	jdff dff_A_KvN69eRv0_0(.dout(w_n132_0[0]),.din(w_dff_A_KvN69eRv0_0),.clk(gclk));
	jdff dff_A_8qC8Bxil9_0(.dout(w_dff_A_KvN69eRv0_0),.din(w_dff_A_8qC8Bxil9_0),.clk(gclk));
	jdff dff_A_Ahft7AOV4_0(.dout(w_dff_A_8qC8Bxil9_0),.din(w_dff_A_Ahft7AOV4_0),.clk(gclk));
	jdff dff_A_EvMmlDyf5_0(.dout(w_dff_A_Ahft7AOV4_0),.din(w_dff_A_EvMmlDyf5_0),.clk(gclk));
	jdff dff_A_0KBaRO998_0(.dout(w_dff_A_EvMmlDyf5_0),.din(w_dff_A_0KBaRO998_0),.clk(gclk));
	jdff dff_A_HxjKhfpm3_0(.dout(w_dff_A_0KBaRO998_0),.din(w_dff_A_HxjKhfpm3_0),.clk(gclk));
	jdff dff_A_FYfj79HQ6_0(.dout(w_n130_0[0]),.din(w_dff_A_FYfj79HQ6_0),.clk(gclk));
	jdff dff_A_nqUp2RTk9_0(.dout(w_dff_A_FYfj79HQ6_0),.din(w_dff_A_nqUp2RTk9_0),.clk(gclk));
	jdff dff_A_5TRk2knt2_0(.dout(w_dff_A_nqUp2RTk9_0),.din(w_dff_A_5TRk2knt2_0),.clk(gclk));
	jdff dff_A_55IHtMGb3_0(.dout(w_dff_A_5TRk2knt2_0),.din(w_dff_A_55IHtMGb3_0),.clk(gclk));
	jdff dff_A_ikW0gD047_0(.dout(w_dff_A_55IHtMGb3_0),.din(w_dff_A_ikW0gD047_0),.clk(gclk));
	jdff dff_A_rvw2qnGv6_1(.dout(w_n130_0[1]),.din(w_dff_A_rvw2qnGv6_1),.clk(gclk));
	jdff dff_A_LzYGizPC2_1(.dout(w_dff_A_rvw2qnGv6_1),.din(w_dff_A_LzYGizPC2_1),.clk(gclk));
	jdff dff_A_SrzJZZRR9_1(.dout(w_dff_A_LzYGizPC2_1),.din(w_dff_A_SrzJZZRR9_1),.clk(gclk));
	jdff dff_A_8EMDDm7r3_1(.dout(w_dff_A_SrzJZZRR9_1),.din(w_dff_A_8EMDDm7r3_1),.clk(gclk));
	jdff dff_A_Ss3t7B913_1(.dout(w_dff_A_8EMDDm7r3_1),.din(w_dff_A_Ss3t7B913_1),.clk(gclk));
	jdff dff_B_esKR7kkk1_3(.din(n130),.dout(w_dff_B_esKR7kkk1_3),.clk(gclk));
	jdff dff_B_yQY2moTH4_3(.din(w_dff_B_esKR7kkk1_3),.dout(w_dff_B_yQY2moTH4_3),.clk(gclk));
	jdff dff_B_oeXp4PmU3_3(.din(w_dff_B_yQY2moTH4_3),.dout(w_dff_B_oeXp4PmU3_3),.clk(gclk));
	jdff dff_B_ttlJSbP61_3(.din(w_dff_B_oeXp4PmU3_3),.dout(w_dff_B_ttlJSbP61_3),.clk(gclk));
	jdff dff_B_Qfl55UKq8_3(.din(w_dff_B_ttlJSbP61_3),.dout(w_dff_B_Qfl55UKq8_3),.clk(gclk));
	jdff dff_B_mKkf82ms6_3(.din(w_dff_B_Qfl55UKq8_3),.dout(w_dff_B_mKkf82ms6_3),.clk(gclk));
	jdff dff_B_duBsfNaE5_3(.din(w_dff_B_mKkf82ms6_3),.dout(w_dff_B_duBsfNaE5_3),.clk(gclk));
	jdff dff_A_hnpq7YPZ0_0(.dout(w_G21gat_1[0]),.din(w_dff_A_hnpq7YPZ0_0),.clk(gclk));
	jdff dff_A_6ZzR6NVO8_0(.dout(w_dff_A_hnpq7YPZ0_0),.din(w_dff_A_6ZzR6NVO8_0),.clk(gclk));
	jdff dff_A_IhUCNGIH8_0(.dout(w_dff_A_6ZzR6NVO8_0),.din(w_dff_A_IhUCNGIH8_0),.clk(gclk));
	jdff dff_A_yaCqGn8t2_0(.dout(w_dff_A_IhUCNGIH8_0),.din(w_dff_A_yaCqGn8t2_0),.clk(gclk));
	jdff dff_A_unDrCpin6_0(.dout(w_dff_A_yaCqGn8t2_0),.din(w_dff_A_unDrCpin6_0),.clk(gclk));
	jdff dff_A_alPvvsFh2_0(.dout(w_dff_A_unDrCpin6_0),.din(w_dff_A_alPvvsFh2_0),.clk(gclk));
	jdff dff_A_Mr5eIYlc5_0(.dout(w_dff_A_alPvvsFh2_0),.din(w_dff_A_Mr5eIYlc5_0),.clk(gclk));
	jdff dff_A_6wYury1T2_0(.dout(w_dff_A_Mr5eIYlc5_0),.din(w_dff_A_6wYury1T2_0),.clk(gclk));
	jdff dff_A_vz536jsF4_1(.dout(w_G21gat_0[1]),.din(w_dff_A_vz536jsF4_1),.clk(gclk));
	jdff dff_A_zOFjjEo51_1(.dout(w_dff_A_vz536jsF4_1),.din(w_dff_A_zOFjjEo51_1),.clk(gclk));
	jdff dff_A_OjvD6dLG8_1(.dout(w_dff_A_zOFjjEo51_1),.din(w_dff_A_OjvD6dLG8_1),.clk(gclk));
	jdff dff_A_JjBEHFzh0_1(.dout(w_dff_A_OjvD6dLG8_1),.din(w_dff_A_JjBEHFzh0_1),.clk(gclk));
	jdff dff_A_GIjglU9u6_1(.dout(w_dff_A_JjBEHFzh0_1),.din(w_dff_A_GIjglU9u6_1),.clk(gclk));
	jdff dff_A_elrsTPmC6_1(.dout(w_dff_A_GIjglU9u6_1),.din(w_dff_A_elrsTPmC6_1),.clk(gclk));
	jdff dff_A_gzX4iWzT6_1(.dout(w_dff_A_elrsTPmC6_1),.din(w_dff_A_gzX4iWzT6_1),.clk(gclk));
	jdff dff_A_wf3DvDfL8_1(.dout(w_dff_A_gzX4iWzT6_1),.din(w_dff_A_wf3DvDfL8_1),.clk(gclk));
	jdff dff_A_WHh6n79A7_1(.dout(w_dff_A_wf3DvDfL8_1),.din(w_dff_A_WHh6n79A7_1),.clk(gclk));
	jdff dff_A_LSGuI2nP5_1(.dout(w_dff_A_WHh6n79A7_1),.din(w_dff_A_LSGuI2nP5_1),.clk(gclk));
	jdff dff_A_MIwgaU5U1_1(.dout(w_dff_A_LSGuI2nP5_1),.din(w_dff_A_MIwgaU5U1_1),.clk(gclk));
	jdff dff_A_BmWdvScP5_1(.dout(w_dff_A_MIwgaU5U1_1),.din(w_dff_A_BmWdvScP5_1),.clk(gclk));
	jdff dff_A_ylkeI8A80_1(.dout(w_dff_A_BmWdvScP5_1),.din(w_dff_A_ylkeI8A80_1),.clk(gclk));
	jdff dff_A_P90YzDTl9_2(.dout(w_G21gat_0[2]),.din(w_dff_A_P90YzDTl9_2),.clk(gclk));
	jdff dff_A_kkPlUJ2S0_2(.dout(w_dff_A_P90YzDTl9_2),.din(w_dff_A_kkPlUJ2S0_2),.clk(gclk));
	jdff dff_A_boGCpCYk7_2(.dout(w_dff_A_kkPlUJ2S0_2),.din(w_dff_A_boGCpCYk7_2),.clk(gclk));
	jdff dff_A_r0km9SAv1_2(.dout(w_dff_A_boGCpCYk7_2),.din(w_dff_A_r0km9SAv1_2),.clk(gclk));
	jdff dff_A_cbe27X4j3_2(.dout(w_dff_A_r0km9SAv1_2),.din(w_dff_A_cbe27X4j3_2),.clk(gclk));
	jdff dff_A_FtHp9jB85_2(.dout(w_dff_A_cbe27X4j3_2),.din(w_dff_A_FtHp9jB85_2),.clk(gclk));
	jdff dff_A_1cc9wIDL4_2(.dout(w_dff_A_FtHp9jB85_2),.din(w_dff_A_1cc9wIDL4_2),.clk(gclk));
	jdff dff_A_2S56qNHh7_2(.dout(w_dff_A_1cc9wIDL4_2),.din(w_dff_A_2S56qNHh7_2),.clk(gclk));
	jdff dff_A_ngVAlWUj2_2(.dout(w_dff_A_2S56qNHh7_2),.din(w_dff_A_ngVAlWUj2_2),.clk(gclk));
	jdff dff_A_1LyjpzAE0_2(.dout(w_dff_A_ngVAlWUj2_2),.din(w_dff_A_1LyjpzAE0_2),.clk(gclk));
	jdff dff_A_8bhxMlF20_2(.dout(w_dff_A_1LyjpzAE0_2),.din(w_dff_A_8bhxMlF20_2),.clk(gclk));
	jdff dff_A_CgRXMc1o9_2(.dout(w_dff_A_8bhxMlF20_2),.din(w_dff_A_CgRXMc1o9_2),.clk(gclk));
	jdff dff_A_8CzVoGhG7_2(.dout(w_dff_A_CgRXMc1o9_2),.din(w_dff_A_8CzVoGhG7_2),.clk(gclk));
	jdff dff_A_pCSGokb38_0(.dout(w_n128_0[0]),.din(w_dff_A_pCSGokb38_0),.clk(gclk));
	jdff dff_A_IWZY9deA1_0(.dout(w_dff_A_pCSGokb38_0),.din(w_dff_A_IWZY9deA1_0),.clk(gclk));
	jdff dff_A_Qx3ogJgN7_0(.dout(w_dff_A_IWZY9deA1_0),.din(w_dff_A_Qx3ogJgN7_0),.clk(gclk));
	jdff dff_A_xCyHPCLS3_0(.dout(w_dff_A_Qx3ogJgN7_0),.din(w_dff_A_xCyHPCLS3_0),.clk(gclk));
	jdff dff_A_dRSkMPP55_0(.dout(w_dff_A_xCyHPCLS3_0),.din(w_dff_A_dRSkMPP55_0),.clk(gclk));
	jdff dff_A_nFqf8QzF1_0(.dout(w_dff_A_dRSkMPP55_0),.din(w_dff_A_nFqf8QzF1_0),.clk(gclk));
	jdff dff_A_2zuZ6jFB0_0(.dout(w_n126_0[0]),.din(w_dff_A_2zuZ6jFB0_0),.clk(gclk));
	jdff dff_A_D64y7Lok3_0(.dout(w_dff_A_2zuZ6jFB0_0),.din(w_dff_A_D64y7Lok3_0),.clk(gclk));
	jdff dff_A_nfY9ctfx9_0(.dout(w_dff_A_D64y7Lok3_0),.din(w_dff_A_nfY9ctfx9_0),.clk(gclk));
	jdff dff_A_6DMYWMBQ7_0(.dout(w_dff_A_nfY9ctfx9_0),.din(w_dff_A_6DMYWMBQ7_0),.clk(gclk));
	jdff dff_A_QLBicpOR7_0(.dout(w_dff_A_6DMYWMBQ7_0),.din(w_dff_A_QLBicpOR7_0),.clk(gclk));
	jdff dff_A_C7ESVwgH7_1(.dout(w_n126_0[1]),.din(w_dff_A_C7ESVwgH7_1),.clk(gclk));
	jdff dff_A_SNot2wgA3_1(.dout(w_dff_A_C7ESVwgH7_1),.din(w_dff_A_SNot2wgA3_1),.clk(gclk));
	jdff dff_A_p5ML6ha55_1(.dout(w_dff_A_SNot2wgA3_1),.din(w_dff_A_p5ML6ha55_1),.clk(gclk));
	jdff dff_A_sgt5feMI3_1(.dout(w_dff_A_p5ML6ha55_1),.din(w_dff_A_sgt5feMI3_1),.clk(gclk));
	jdff dff_A_u7RDWOiz3_1(.dout(w_dff_A_sgt5feMI3_1),.din(w_dff_A_u7RDWOiz3_1),.clk(gclk));
	jdff dff_B_7iFtbWKM7_3(.din(n126),.dout(w_dff_B_7iFtbWKM7_3),.clk(gclk));
	jdff dff_B_uckc6IQQ9_3(.din(w_dff_B_7iFtbWKM7_3),.dout(w_dff_B_uckc6IQQ9_3),.clk(gclk));
	jdff dff_B_GtsIZzQw2_3(.din(w_dff_B_uckc6IQQ9_3),.dout(w_dff_B_GtsIZzQw2_3),.clk(gclk));
	jdff dff_B_QL9zLZh95_3(.din(w_dff_B_GtsIZzQw2_3),.dout(w_dff_B_QL9zLZh95_3),.clk(gclk));
	jdff dff_B_C9hIiv3k6_3(.din(w_dff_B_QL9zLZh95_3),.dout(w_dff_B_C9hIiv3k6_3),.clk(gclk));
	jdff dff_B_DnfFyvX56_3(.din(w_dff_B_C9hIiv3k6_3),.dout(w_dff_B_DnfFyvX56_3),.clk(gclk));
	jdff dff_B_SWO0A4BS1_3(.din(w_dff_B_DnfFyvX56_3),.dout(w_dff_B_SWO0A4BS1_3),.clk(gclk));
	jdff dff_A_kcobK8Is2_0(.dout(w_G86gat_1[0]),.din(w_dff_A_kcobK8Is2_0),.clk(gclk));
	jdff dff_A_CQM9eZFe7_0(.dout(w_dff_A_kcobK8Is2_0),.din(w_dff_A_CQM9eZFe7_0),.clk(gclk));
	jdff dff_A_slPQWZ2C3_0(.dout(w_dff_A_CQM9eZFe7_0),.din(w_dff_A_slPQWZ2C3_0),.clk(gclk));
	jdff dff_A_TFALbzua9_0(.dout(w_dff_A_slPQWZ2C3_0),.din(w_dff_A_TFALbzua9_0),.clk(gclk));
	jdff dff_A_9EKSZZo06_0(.dout(w_dff_A_TFALbzua9_0),.din(w_dff_A_9EKSZZo06_0),.clk(gclk));
	jdff dff_A_cjXAEE6s3_0(.dout(w_dff_A_9EKSZZo06_0),.din(w_dff_A_cjXAEE6s3_0),.clk(gclk));
	jdff dff_A_BtYnkijl0_0(.dout(w_dff_A_cjXAEE6s3_0),.din(w_dff_A_BtYnkijl0_0),.clk(gclk));
	jdff dff_A_zpvm1eo74_0(.dout(w_dff_A_BtYnkijl0_0),.din(w_dff_A_zpvm1eo74_0),.clk(gclk));
	jdff dff_A_yvnGjsRs8_1(.dout(w_G86gat_0[1]),.din(w_dff_A_yvnGjsRs8_1),.clk(gclk));
	jdff dff_A_rw8qT8P43_1(.dout(w_dff_A_yvnGjsRs8_1),.din(w_dff_A_rw8qT8P43_1),.clk(gclk));
	jdff dff_A_jlDVpJ7x8_1(.dout(w_dff_A_rw8qT8P43_1),.din(w_dff_A_jlDVpJ7x8_1),.clk(gclk));
	jdff dff_A_bOKXQDzp5_1(.dout(w_dff_A_jlDVpJ7x8_1),.din(w_dff_A_bOKXQDzp5_1),.clk(gclk));
	jdff dff_A_ve1rEFdc6_1(.dout(w_dff_A_bOKXQDzp5_1),.din(w_dff_A_ve1rEFdc6_1),.clk(gclk));
	jdff dff_A_sVMokOZU3_1(.dout(w_dff_A_ve1rEFdc6_1),.din(w_dff_A_sVMokOZU3_1),.clk(gclk));
	jdff dff_A_KFc4OUjj6_1(.dout(w_dff_A_sVMokOZU3_1),.din(w_dff_A_KFc4OUjj6_1),.clk(gclk));
	jdff dff_A_GPzwGosk0_1(.dout(w_dff_A_KFc4OUjj6_1),.din(w_dff_A_GPzwGosk0_1),.clk(gclk));
	jdff dff_A_lRCmjHhC6_1(.dout(w_dff_A_GPzwGosk0_1),.din(w_dff_A_lRCmjHhC6_1),.clk(gclk));
	jdff dff_A_0xwpSxdc4_1(.dout(w_dff_A_lRCmjHhC6_1),.din(w_dff_A_0xwpSxdc4_1),.clk(gclk));
	jdff dff_A_4OjroygO6_1(.dout(w_dff_A_0xwpSxdc4_1),.din(w_dff_A_4OjroygO6_1),.clk(gclk));
	jdff dff_A_xsWauW9u4_1(.dout(w_dff_A_4OjroygO6_1),.din(w_dff_A_xsWauW9u4_1),.clk(gclk));
	jdff dff_A_3RY14p7Q2_1(.dout(w_dff_A_xsWauW9u4_1),.din(w_dff_A_3RY14p7Q2_1),.clk(gclk));
	jdff dff_A_ABVZFhL37_2(.dout(w_G86gat_0[2]),.din(w_dff_A_ABVZFhL37_2),.clk(gclk));
	jdff dff_A_zuVWxMWC9_2(.dout(w_dff_A_ABVZFhL37_2),.din(w_dff_A_zuVWxMWC9_2),.clk(gclk));
	jdff dff_A_WNcFqDLe9_2(.dout(w_dff_A_zuVWxMWC9_2),.din(w_dff_A_WNcFqDLe9_2),.clk(gclk));
	jdff dff_A_fzOGFt1a7_2(.dout(w_dff_A_WNcFqDLe9_2),.din(w_dff_A_fzOGFt1a7_2),.clk(gclk));
	jdff dff_A_ubA3NRgw2_2(.dout(w_dff_A_fzOGFt1a7_2),.din(w_dff_A_ubA3NRgw2_2),.clk(gclk));
	jdff dff_A_OOhARacv6_2(.dout(w_dff_A_ubA3NRgw2_2),.din(w_dff_A_OOhARacv6_2),.clk(gclk));
	jdff dff_A_hE7n0a4I7_2(.dout(w_dff_A_OOhARacv6_2),.din(w_dff_A_hE7n0a4I7_2),.clk(gclk));
	jdff dff_A_UoDmrJph5_2(.dout(w_dff_A_hE7n0a4I7_2),.din(w_dff_A_UoDmrJph5_2),.clk(gclk));
	jdff dff_A_zIohYmyg3_2(.dout(w_dff_A_UoDmrJph5_2),.din(w_dff_A_zIohYmyg3_2),.clk(gclk));
	jdff dff_A_Bq1laqnH5_2(.dout(w_dff_A_zIohYmyg3_2),.din(w_dff_A_Bq1laqnH5_2),.clk(gclk));
	jdff dff_A_RsgW4ij96_2(.dout(w_dff_A_Bq1laqnH5_2),.din(w_dff_A_RsgW4ij96_2),.clk(gclk));
	jdff dff_A_ktF3Za192_2(.dout(w_dff_A_RsgW4ij96_2),.din(w_dff_A_ktF3Za192_2),.clk(gclk));
	jdff dff_A_kTePh0YY1_2(.dout(w_dff_A_ktF3Za192_2),.din(w_dff_A_kTePh0YY1_2),.clk(gclk));
	jdff dff_B_rsRN4gi21_0(.din(n124),.dout(w_dff_B_rsRN4gi21_0),.clk(gclk));
	jdff dff_A_DD2EwS6E1_1(.dout(w_n123_0[1]),.din(w_dff_A_DD2EwS6E1_1),.clk(gclk));
	jdff dff_A_3mO9yJA19_1(.dout(w_dff_A_DD2EwS6E1_1),.din(w_dff_A_3mO9yJA19_1),.clk(gclk));
	jdff dff_A_GqZtSLYu0_1(.dout(w_dff_A_3mO9yJA19_1),.din(w_dff_A_GqZtSLYu0_1),.clk(gclk));
	jdff dff_A_LNLRBGh42_1(.dout(w_dff_A_GqZtSLYu0_1),.din(w_dff_A_LNLRBGh42_1),.clk(gclk));
	jdff dff_A_0GVK19w73_1(.dout(w_dff_A_LNLRBGh42_1),.din(w_dff_A_0GVK19w73_1),.clk(gclk));
	jdff dff_A_EUSJa4NQ3_0(.dout(w_G47gat_0[0]),.din(w_dff_A_EUSJa4NQ3_0),.clk(gclk));
	jdff dff_A_UzJrRbZe3_0(.dout(w_dff_A_EUSJa4NQ3_0),.din(w_dff_A_UzJrRbZe3_0),.clk(gclk));
	jdff dff_A_vFgpuMpX8_0(.dout(w_dff_A_UzJrRbZe3_0),.din(w_dff_A_vFgpuMpX8_0),.clk(gclk));
	jdff dff_A_jJt15PHk3_0(.dout(w_dff_A_vFgpuMpX8_0),.din(w_dff_A_jJt15PHk3_0),.clk(gclk));
	jdff dff_A_gObTqNUE4_0(.dout(w_dff_A_jJt15PHk3_0),.din(w_dff_A_gObTqNUE4_0),.clk(gclk));
	jdff dff_A_jE8scXq03_0(.dout(w_dff_A_gObTqNUE4_0),.din(w_dff_A_jE8scXq03_0),.clk(gclk));
	jdff dff_A_qyEOFRol2_0(.dout(w_dff_A_jE8scXq03_0),.din(w_dff_A_qyEOFRol2_0),.clk(gclk));
	jdff dff_A_RezMjxAs2_0(.dout(w_dff_A_qyEOFRol2_0),.din(w_dff_A_RezMjxAs2_0),.clk(gclk));
	jdff dff_A_s2sk7ri67_0(.dout(w_dff_A_RezMjxAs2_0),.din(w_dff_A_s2sk7ri67_0),.clk(gclk));
	jdff dff_A_0Hp699qs0_0(.dout(w_dff_A_s2sk7ri67_0),.din(w_dff_A_0Hp699qs0_0),.clk(gclk));
	jdff dff_A_4bkjgAZJ1_0(.dout(w_dff_A_0Hp699qs0_0),.din(w_dff_A_4bkjgAZJ1_0),.clk(gclk));
	jdff dff_A_cENlmcPz9_0(.dout(w_dff_A_4bkjgAZJ1_0),.din(w_dff_A_cENlmcPz9_0),.clk(gclk));
	jdff dff_A_7wffRQjy9_0(.dout(w_dff_A_cENlmcPz9_0),.din(w_dff_A_7wffRQjy9_0),.clk(gclk));
	jdff dff_B_Fv6m2CzD8_1(.din(n117),.dout(w_dff_B_Fv6m2CzD8_1),.clk(gclk));
	jdff dff_B_TmclbHEC8_1(.din(w_dff_B_Fv6m2CzD8_1),.dout(w_dff_B_TmclbHEC8_1),.clk(gclk));
	jdff dff_B_KBCDqDzO1_1(.din(w_dff_B_TmclbHEC8_1),.dout(w_dff_B_KBCDqDzO1_1),.clk(gclk));
	jdff dff_B_YhorwD8j4_1(.din(w_dff_B_KBCDqDzO1_1),.dout(w_dff_B_YhorwD8j4_1),.clk(gclk));
	jdff dff_B_wKH6W4uK7_1(.din(w_dff_B_YhorwD8j4_1),.dout(w_dff_B_wKH6W4uK7_1),.clk(gclk));
	jdff dff_B_aokus66T8_1(.din(w_dff_B_wKH6W4uK7_1),.dout(w_dff_B_aokus66T8_1),.clk(gclk));
	jdff dff_B_u6r39nYs8_1(.din(w_dff_B_aokus66T8_1),.dout(w_dff_B_u6r39nYs8_1),.clk(gclk));
	jdff dff_A_it2qwHqH0_0(.dout(w_G60gat_0[0]),.din(w_dff_A_it2qwHqH0_0),.clk(gclk));
	jdff dff_A_qwn3zPLH3_0(.dout(w_dff_A_it2qwHqH0_0),.din(w_dff_A_qwn3zPLH3_0),.clk(gclk));
	jdff dff_A_cyDwvHrD6_0(.dout(w_dff_A_qwn3zPLH3_0),.din(w_dff_A_cyDwvHrD6_0),.clk(gclk));
	jdff dff_A_wHUrBUHx2_0(.dout(w_dff_A_cyDwvHrD6_0),.din(w_dff_A_wHUrBUHx2_0),.clk(gclk));
	jdff dff_A_tm1iovNG2_0(.dout(w_dff_A_wHUrBUHx2_0),.din(w_dff_A_tm1iovNG2_0),.clk(gclk));
	jdff dff_A_fOcwSh3o6_0(.dout(w_dff_A_tm1iovNG2_0),.din(w_dff_A_fOcwSh3o6_0),.clk(gclk));
	jdff dff_A_ECDtJwif4_0(.dout(w_dff_A_fOcwSh3o6_0),.din(w_dff_A_ECDtJwif4_0),.clk(gclk));
	jdff dff_A_2GhpTHQo1_0(.dout(w_dff_A_ECDtJwif4_0),.din(w_dff_A_2GhpTHQo1_0),.clk(gclk));
	jdff dff_A_2S4R9faL7_0(.dout(w_dff_A_2GhpTHQo1_0),.din(w_dff_A_2S4R9faL7_0),.clk(gclk));
	jdff dff_A_ODmWjlRV5_0(.dout(w_dff_A_2S4R9faL7_0),.din(w_dff_A_ODmWjlRV5_0),.clk(gclk));
	jdff dff_A_rd3Fba8s6_0(.dout(w_dff_A_ODmWjlRV5_0),.din(w_dff_A_rd3Fba8s6_0),.clk(gclk));
	jdff dff_A_tko4XCxQ2_0(.dout(w_dff_A_rd3Fba8s6_0),.din(w_dff_A_tko4XCxQ2_0),.clk(gclk));
	jdff dff_A_tKksQxqR6_0(.dout(w_dff_A_tko4XCxQ2_0),.din(w_dff_A_tKksQxqR6_0),.clk(gclk));
	jdff dff_A_KEyb8s4Y9_1(.dout(w_G60gat_0[1]),.din(w_dff_A_KEyb8s4Y9_1),.clk(gclk));
	jdff dff_A_U5B2XVT57_1(.dout(w_dff_A_KEyb8s4Y9_1),.din(w_dff_A_U5B2XVT57_1),.clk(gclk));
	jdff dff_A_tgiBVSHu4_1(.dout(w_dff_A_U5B2XVT57_1),.din(w_dff_A_tgiBVSHu4_1),.clk(gclk));
	jdff dff_A_eucTybFG0_1(.dout(w_dff_A_tgiBVSHu4_1),.din(w_dff_A_eucTybFG0_1),.clk(gclk));
	jdff dff_A_dyrbwCaQ3_1(.dout(w_dff_A_eucTybFG0_1),.din(w_dff_A_dyrbwCaQ3_1),.clk(gclk));
	jdff dff_A_zPHajorB1_1(.dout(w_dff_A_dyrbwCaQ3_1),.din(w_dff_A_zPHajorB1_1),.clk(gclk));
	jdff dff_A_0r1rFZJN2_1(.dout(w_dff_A_zPHajorB1_1),.din(w_dff_A_0r1rFZJN2_1),.clk(gclk));
	jdff dff_A_gtyfAx5u2_1(.dout(w_dff_A_0r1rFZJN2_1),.din(w_dff_A_gtyfAx5u2_1),.clk(gclk));
	jdff dff_A_lyQsZuTS8_0(.dout(w_n115_0[0]),.din(w_dff_A_lyQsZuTS8_0),.clk(gclk));
	jdff dff_A_8PsZVu7s4_0(.dout(w_dff_A_lyQsZuTS8_0),.din(w_dff_A_8PsZVu7s4_0),.clk(gclk));
	jdff dff_A_4x2ufxxD8_0(.dout(w_n114_0[0]),.din(w_dff_A_4x2ufxxD8_0),.clk(gclk));
	jdff dff_A_5P6RYtYA6_0(.dout(w_dff_A_4x2ufxxD8_0),.din(w_dff_A_5P6RYtYA6_0),.clk(gclk));
	jdff dff_A_z7doHYr38_0(.dout(w_dff_A_5P6RYtYA6_0),.din(w_dff_A_z7doHYr38_0),.clk(gclk));
	jdff dff_A_bU20rqy65_0(.dout(w_dff_A_z7doHYr38_0),.din(w_dff_A_bU20rqy65_0),.clk(gclk));
	jdff dff_A_O709u4Bz7_0(.dout(w_dff_A_bU20rqy65_0),.din(w_dff_A_O709u4Bz7_0),.clk(gclk));
	jdff dff_A_2iAQPlyp8_0(.dout(w_dff_A_O709u4Bz7_0),.din(w_dff_A_2iAQPlyp8_0),.clk(gclk));
	jdff dff_A_hiYXJa653_0(.dout(w_G34gat_0[0]),.din(w_dff_A_hiYXJa653_0),.clk(gclk));
	jdff dff_A_ZkJX8wsO7_0(.dout(w_dff_A_hiYXJa653_0),.din(w_dff_A_ZkJX8wsO7_0),.clk(gclk));
	jdff dff_A_O1gGKJgq3_0(.dout(w_dff_A_ZkJX8wsO7_0),.din(w_dff_A_O1gGKJgq3_0),.clk(gclk));
	jdff dff_A_w1nJKGU09_0(.dout(w_dff_A_O1gGKJgq3_0),.din(w_dff_A_w1nJKGU09_0),.clk(gclk));
	jdff dff_A_GsPdezS24_0(.dout(w_dff_A_w1nJKGU09_0),.din(w_dff_A_GsPdezS24_0),.clk(gclk));
	jdff dff_A_EZTCzFBR7_0(.dout(w_dff_A_GsPdezS24_0),.din(w_dff_A_EZTCzFBR7_0),.clk(gclk));
	jdff dff_A_hAAFYBmp5_0(.dout(w_dff_A_EZTCzFBR7_0),.din(w_dff_A_hAAFYBmp5_0),.clk(gclk));
	jdff dff_A_kAASZgl22_0(.dout(w_dff_A_hAAFYBmp5_0),.din(w_dff_A_kAASZgl22_0),.clk(gclk));
	jdff dff_A_XCqU0mN41_0(.dout(w_dff_A_kAASZgl22_0),.din(w_dff_A_XCqU0mN41_0),.clk(gclk));
	jdff dff_A_ay6l1FQL0_0(.dout(w_dff_A_XCqU0mN41_0),.din(w_dff_A_ay6l1FQL0_0),.clk(gclk));
	jdff dff_A_doOqM7bH5_0(.dout(w_dff_A_ay6l1FQL0_0),.din(w_dff_A_doOqM7bH5_0),.clk(gclk));
	jdff dff_A_Ctzd03QN7_0(.dout(w_dff_A_doOqM7bH5_0),.din(w_dff_A_Ctzd03QN7_0),.clk(gclk));
	jdff dff_A_kTjO4ryG8_0(.dout(w_dff_A_Ctzd03QN7_0),.din(w_dff_A_kTjO4ryG8_0),.clk(gclk));
	jdff dff_A_2Esfz2Cc2_2(.dout(w_G34gat_0[2]),.din(w_dff_A_2Esfz2Cc2_2),.clk(gclk));
	jdff dff_A_kA7UKfZ70_2(.dout(w_dff_A_2Esfz2Cc2_2),.din(w_dff_A_kA7UKfZ70_2),.clk(gclk));
	jdff dff_A_FNMcSjCE6_2(.dout(w_dff_A_kA7UKfZ70_2),.din(w_dff_A_FNMcSjCE6_2),.clk(gclk));
	jdff dff_A_Sf7DTXvw4_2(.dout(w_dff_A_FNMcSjCE6_2),.din(w_dff_A_Sf7DTXvw4_2),.clk(gclk));
	jdff dff_A_IodsmCM40_2(.dout(w_dff_A_Sf7DTXvw4_2),.din(w_dff_A_IodsmCM40_2),.clk(gclk));
	jdff dff_A_OGXhtmPX5_2(.dout(w_dff_A_IodsmCM40_2),.din(w_dff_A_OGXhtmPX5_2),.clk(gclk));
	jdff dff_A_PJ5ac82i5_2(.dout(w_dff_A_OGXhtmPX5_2),.din(w_dff_A_PJ5ac82i5_2),.clk(gclk));
	jdff dff_A_HLRxu9hC8_2(.dout(w_dff_A_PJ5ac82i5_2),.din(w_dff_A_HLRxu9hC8_2),.clk(gclk));
	jdff dff_A_pdZLw88M9_0(.dout(w_n109_0[0]),.din(w_dff_A_pdZLw88M9_0),.clk(gclk));
	jdff dff_A_3T5QZSFe4_0(.dout(w_dff_A_pdZLw88M9_0),.din(w_dff_A_3T5QZSFe4_0),.clk(gclk));
	jdff dff_A_Ix1wpVIR0_0(.dout(w_dff_A_3T5QZSFe4_0),.din(w_dff_A_Ix1wpVIR0_0),.clk(gclk));
	jdff dff_A_QAVbQ8KG3_0(.dout(w_dff_A_Ix1wpVIR0_0),.din(w_dff_A_QAVbQ8KG3_0),.clk(gclk));
	jdff dff_A_ousPHLrB5_0(.dout(w_dff_A_QAVbQ8KG3_0),.din(w_dff_A_ousPHLrB5_0),.clk(gclk));
	jdff dff_A_riHUICMo6_0(.dout(w_dff_A_ousPHLrB5_0),.din(w_dff_A_riHUICMo6_0),.clk(gclk));
	jdff dff_A_1BCrSjlV2_0(.dout(w_n107_0[0]),.din(w_dff_A_1BCrSjlV2_0),.clk(gclk));
	jdff dff_A_ad8fcmtR1_0(.dout(w_dff_A_1BCrSjlV2_0),.din(w_dff_A_ad8fcmtR1_0),.clk(gclk));
	jdff dff_A_XH5Xx23o7_0(.dout(w_dff_A_ad8fcmtR1_0),.din(w_dff_A_XH5Xx23o7_0),.clk(gclk));
	jdff dff_A_MJcv7u0l3_0(.dout(w_dff_A_XH5Xx23o7_0),.din(w_dff_A_MJcv7u0l3_0),.clk(gclk));
	jdff dff_A_Klo8Z9nq0_0(.dout(w_dff_A_MJcv7u0l3_0),.din(w_dff_A_Klo8Z9nq0_0),.clk(gclk));
	jdff dff_B_vbNPuuRj4_2(.din(n107),.dout(w_dff_B_vbNPuuRj4_2),.clk(gclk));
	jdff dff_B_wXu0phGn4_2(.din(w_dff_B_vbNPuuRj4_2),.dout(w_dff_B_wXu0phGn4_2),.clk(gclk));
	jdff dff_B_TC71sZVX0_2(.din(w_dff_B_wXu0phGn4_2),.dout(w_dff_B_TC71sZVX0_2),.clk(gclk));
	jdff dff_B_riSjZN5b5_2(.din(w_dff_B_TC71sZVX0_2),.dout(w_dff_B_riSjZN5b5_2),.clk(gclk));
	jdff dff_B_yXinODag7_2(.din(w_dff_B_riSjZN5b5_2),.dout(w_dff_B_yXinODag7_2),.clk(gclk));
	jdff dff_B_Qo2yRTwU3_2(.din(w_dff_B_yXinODag7_2),.dout(w_dff_B_Qo2yRTwU3_2),.clk(gclk));
	jdff dff_B_Qpnbjv8i6_2(.din(w_dff_B_Qo2yRTwU3_2),.dout(w_dff_B_Qpnbjv8i6_2),.clk(gclk));
	jdff dff_A_1jLi4RYx1_0(.dout(w_G73gat_0[0]),.din(w_dff_A_1jLi4RYx1_0),.clk(gclk));
	jdff dff_A_hdwRdQAI2_0(.dout(w_dff_A_1jLi4RYx1_0),.din(w_dff_A_hdwRdQAI2_0),.clk(gclk));
	jdff dff_A_I0FAqYFk4_0(.dout(w_dff_A_hdwRdQAI2_0),.din(w_dff_A_I0FAqYFk4_0),.clk(gclk));
	jdff dff_A_RPQm22uG9_0(.dout(w_dff_A_I0FAqYFk4_0),.din(w_dff_A_RPQm22uG9_0),.clk(gclk));
	jdff dff_A_ToZX8LuQ5_0(.dout(w_dff_A_RPQm22uG9_0),.din(w_dff_A_ToZX8LuQ5_0),.clk(gclk));
	jdff dff_A_Eqvtuz0k7_0(.dout(w_dff_A_ToZX8LuQ5_0),.din(w_dff_A_Eqvtuz0k7_0),.clk(gclk));
	jdff dff_A_9Iq4itu71_0(.dout(w_dff_A_Eqvtuz0k7_0),.din(w_dff_A_9Iq4itu71_0),.clk(gclk));
	jdff dff_A_hgpJNaHG9_0(.dout(w_dff_A_9Iq4itu71_0),.din(w_dff_A_hgpJNaHG9_0),.clk(gclk));
	jdff dff_A_GEyPZXY59_0(.dout(w_dff_A_hgpJNaHG9_0),.din(w_dff_A_GEyPZXY59_0),.clk(gclk));
	jdff dff_A_85mXJdqJ6_0(.dout(w_dff_A_GEyPZXY59_0),.din(w_dff_A_85mXJdqJ6_0),.clk(gclk));
	jdff dff_A_XiE6s5Pe4_0(.dout(w_dff_A_85mXJdqJ6_0),.din(w_dff_A_XiE6s5Pe4_0),.clk(gclk));
	jdff dff_A_OxhLI8F16_0(.dout(w_dff_A_XiE6s5Pe4_0),.din(w_dff_A_OxhLI8F16_0),.clk(gclk));
	jdff dff_A_Uf4wyVZi1_0(.dout(w_dff_A_OxhLI8F16_0),.din(w_dff_A_Uf4wyVZi1_0),.clk(gclk));
	jdff dff_A_bmHSz2Tj0_1(.dout(w_G73gat_0[1]),.din(w_dff_A_bmHSz2Tj0_1),.clk(gclk));
	jdff dff_A_qlobzmpw6_1(.dout(w_dff_A_bmHSz2Tj0_1),.din(w_dff_A_qlobzmpw6_1),.clk(gclk));
	jdff dff_A_R441xY9b2_1(.dout(w_dff_A_qlobzmpw6_1),.din(w_dff_A_R441xY9b2_1),.clk(gclk));
	jdff dff_A_V0yOCIhw4_1(.dout(w_dff_A_R441xY9b2_1),.din(w_dff_A_V0yOCIhw4_1),.clk(gclk));
	jdff dff_A_gGJtaM9k0_1(.dout(w_dff_A_V0yOCIhw4_1),.din(w_dff_A_gGJtaM9k0_1),.clk(gclk));
	jdff dff_A_bRpoo7C77_1(.dout(w_dff_A_gGJtaM9k0_1),.din(w_dff_A_bRpoo7C77_1),.clk(gclk));
	jdff dff_A_0C47CxO73_1(.dout(w_dff_A_bRpoo7C77_1),.din(w_dff_A_0C47CxO73_1),.clk(gclk));
	jdff dff_A_LFlt7WTf2_1(.dout(w_dff_A_0C47CxO73_1),.din(w_dff_A_LFlt7WTf2_1),.clk(gclk));
	jdff dff_B_FIU4XNhX5_1(.din(n103),.dout(w_dff_B_FIU4XNhX5_1),.clk(gclk));
	jdff dff_B_E79sbgNT4_1(.din(w_dff_B_FIU4XNhX5_1),.dout(w_dff_B_E79sbgNT4_1),.clk(gclk));
	jdff dff_B_sox4Yx8h2_1(.din(w_dff_B_E79sbgNT4_1),.dout(w_dff_B_sox4Yx8h2_1),.clk(gclk));
	jdff dff_B_BH8cCgRW1_1(.din(w_dff_B_sox4Yx8h2_1),.dout(w_dff_B_BH8cCgRW1_1),.clk(gclk));
	jdff dff_B_1PvCAizf9_1(.din(w_dff_B_BH8cCgRW1_1),.dout(w_dff_B_1PvCAizf9_1),.clk(gclk));
	jdff dff_B_IY29OhhM2_1(.din(w_dff_B_1PvCAizf9_1),.dout(w_dff_B_IY29OhhM2_1),.clk(gclk));
	jdff dff_B_4aXRGgFB2_1(.din(w_dff_B_IY29OhhM2_1),.dout(w_dff_B_4aXRGgFB2_1),.clk(gclk));
	jdff dff_A_Bl0vePuy3_0(.dout(w_G99gat_0[0]),.din(w_dff_A_Bl0vePuy3_0),.clk(gclk));
	jdff dff_A_WPByknKX0_0(.dout(w_dff_A_Bl0vePuy3_0),.din(w_dff_A_WPByknKX0_0),.clk(gclk));
	jdff dff_A_psbqyxzE7_0(.dout(w_dff_A_WPByknKX0_0),.din(w_dff_A_psbqyxzE7_0),.clk(gclk));
	jdff dff_A_vAiuKXTl7_0(.dout(w_dff_A_psbqyxzE7_0),.din(w_dff_A_vAiuKXTl7_0),.clk(gclk));
	jdff dff_A_YDBVrOPt0_0(.dout(w_dff_A_vAiuKXTl7_0),.din(w_dff_A_YDBVrOPt0_0),.clk(gclk));
	jdff dff_A_KHOofYdl2_0(.dout(w_dff_A_YDBVrOPt0_0),.din(w_dff_A_KHOofYdl2_0),.clk(gclk));
	jdff dff_A_BlT9XUv15_0(.dout(w_dff_A_KHOofYdl2_0),.din(w_dff_A_BlT9XUv15_0),.clk(gclk));
	jdff dff_A_4MmouBb57_0(.dout(w_dff_A_BlT9XUv15_0),.din(w_dff_A_4MmouBb57_0),.clk(gclk));
	jdff dff_A_ryZQ9wY16_1(.dout(w_G99gat_0[1]),.din(w_dff_A_ryZQ9wY16_1),.clk(gclk));
	jdff dff_A_NzIrbV8u5_1(.dout(w_dff_A_ryZQ9wY16_1),.din(w_dff_A_NzIrbV8u5_1),.clk(gclk));
	jdff dff_A_NumHLs2G7_1(.dout(w_dff_A_NzIrbV8u5_1),.din(w_dff_A_NumHLs2G7_1),.clk(gclk));
	jdff dff_A_mZHBZK701_1(.dout(w_dff_A_NumHLs2G7_1),.din(w_dff_A_mZHBZK701_1),.clk(gclk));
	jdff dff_A_70pygJTa6_1(.dout(w_dff_A_mZHBZK701_1),.din(w_dff_A_70pygJTa6_1),.clk(gclk));
	jdff dff_A_PNlwz2hy0_1(.dout(w_dff_A_70pygJTa6_1),.din(w_dff_A_PNlwz2hy0_1),.clk(gclk));
	jdff dff_A_5DxUnceN5_1(.dout(w_dff_A_PNlwz2hy0_1),.din(w_dff_A_5DxUnceN5_1),.clk(gclk));
	jdff dff_A_u0Reuen91_1(.dout(w_dff_A_5DxUnceN5_1),.din(w_dff_A_u0Reuen91_1),.clk(gclk));
	jdff dff_A_3S0Noii19_1(.dout(w_dff_A_u0Reuen91_1),.din(w_dff_A_3S0Noii19_1),.clk(gclk));
	jdff dff_A_HOdmcer34_1(.dout(w_dff_A_3S0Noii19_1),.din(w_dff_A_HOdmcer34_1),.clk(gclk));
	jdff dff_A_Js6aPtXj6_1(.dout(w_dff_A_HOdmcer34_1),.din(w_dff_A_Js6aPtXj6_1),.clk(gclk));
	jdff dff_A_ixIbOInX5_1(.dout(w_dff_A_Js6aPtXj6_1),.din(w_dff_A_ixIbOInX5_1),.clk(gclk));
	jdff dff_A_3q3Udb6f2_1(.dout(w_dff_A_ixIbOInX5_1),.din(w_dff_A_3q3Udb6f2_1),.clk(gclk));
	jdff dff_A_3WhSAtBC6_0(.dout(w_n100_0[0]),.din(w_dff_A_3WhSAtBC6_0),.clk(gclk));
	jdff dff_A_C4yHK1bg7_0(.dout(w_dff_A_3WhSAtBC6_0),.din(w_dff_A_C4yHK1bg7_0),.clk(gclk));
	jdff dff_A_OHNi3BtC2_0(.dout(w_dff_A_C4yHK1bg7_0),.din(w_dff_A_OHNi3BtC2_0),.clk(gclk));
	jdff dff_A_tmvUf1fZ7_0(.dout(w_dff_A_OHNi3BtC2_0),.din(w_dff_A_tmvUf1fZ7_0),.clk(gclk));
	jdff dff_A_vry5MGvC5_0(.dout(w_dff_A_tmvUf1fZ7_0),.din(w_dff_A_vry5MGvC5_0),.clk(gclk));
	jdff dff_A_FycskBfx6_0(.dout(w_dff_A_vry5MGvC5_0),.din(w_dff_A_FycskBfx6_0),.clk(gclk));
	jdff dff_A_WYcYWevu1_0(.dout(w_n98_0[0]),.din(w_dff_A_WYcYWevu1_0),.clk(gclk));
	jdff dff_A_bNclPy5R3_0(.dout(w_dff_A_WYcYWevu1_0),.din(w_dff_A_bNclPy5R3_0),.clk(gclk));
	jdff dff_A_SBDThDsY3_0(.dout(w_dff_A_bNclPy5R3_0),.din(w_dff_A_SBDThDsY3_0),.clk(gclk));
	jdff dff_A_buxUTz049_0(.dout(w_dff_A_SBDThDsY3_0),.din(w_dff_A_buxUTz049_0),.clk(gclk));
	jdff dff_A_QQALszhd2_0(.dout(w_dff_A_buxUTz049_0),.din(w_dff_A_QQALszhd2_0),.clk(gclk));
	jdff dff_B_3SWlJP7U6_2(.din(n98),.dout(w_dff_B_3SWlJP7U6_2),.clk(gclk));
	jdff dff_B_H7EoF3O72_2(.din(w_dff_B_3SWlJP7U6_2),.dout(w_dff_B_H7EoF3O72_2),.clk(gclk));
	jdff dff_B_f6U0AA6u9_2(.din(w_dff_B_H7EoF3O72_2),.dout(w_dff_B_f6U0AA6u9_2),.clk(gclk));
	jdff dff_B_jiu8K6Mv4_2(.din(w_dff_B_f6U0AA6u9_2),.dout(w_dff_B_jiu8K6Mv4_2),.clk(gclk));
	jdff dff_B_h5wiugK65_2(.din(w_dff_B_jiu8K6Mv4_2),.dout(w_dff_B_h5wiugK65_2),.clk(gclk));
	jdff dff_B_0L1AhYIW6_2(.din(w_dff_B_h5wiugK65_2),.dout(w_dff_B_0L1AhYIW6_2),.clk(gclk));
	jdff dff_B_zzOnSQo75_2(.din(w_dff_B_0L1AhYIW6_2),.dout(w_dff_B_zzOnSQo75_2),.clk(gclk));
	jdff dff_A_pKoZdVtq3_0(.dout(w_G8gat_0[0]),.din(w_dff_A_pKoZdVtq3_0),.clk(gclk));
	jdff dff_A_LBmYrF4v2_0(.dout(w_dff_A_pKoZdVtq3_0),.din(w_dff_A_LBmYrF4v2_0),.clk(gclk));
	jdff dff_A_vkLkEUDb0_0(.dout(w_dff_A_LBmYrF4v2_0),.din(w_dff_A_vkLkEUDb0_0),.clk(gclk));
	jdff dff_A_8nGOXfmL3_0(.dout(w_dff_A_vkLkEUDb0_0),.din(w_dff_A_8nGOXfmL3_0),.clk(gclk));
	jdff dff_A_tckeineN2_0(.dout(w_dff_A_8nGOXfmL3_0),.din(w_dff_A_tckeineN2_0),.clk(gclk));
	jdff dff_A_V0OZ0ex87_0(.dout(w_dff_A_tckeineN2_0),.din(w_dff_A_V0OZ0ex87_0),.clk(gclk));
	jdff dff_A_RAQ7soBi6_0(.dout(w_dff_A_V0OZ0ex87_0),.din(w_dff_A_RAQ7soBi6_0),.clk(gclk));
	jdff dff_A_3gY0AY0h1_0(.dout(w_dff_A_RAQ7soBi6_0),.din(w_dff_A_3gY0AY0h1_0),.clk(gclk));
	jdff dff_A_stDXda203_0(.dout(w_dff_A_3gY0AY0h1_0),.din(w_dff_A_stDXda203_0),.clk(gclk));
	jdff dff_A_4wrPObSd0_0(.dout(w_dff_A_stDXda203_0),.din(w_dff_A_4wrPObSd0_0),.clk(gclk));
	jdff dff_A_inT0k7Z87_0(.dout(w_dff_A_4wrPObSd0_0),.din(w_dff_A_inT0k7Z87_0),.clk(gclk));
	jdff dff_A_5z3gmTeW9_0(.dout(w_dff_A_inT0k7Z87_0),.din(w_dff_A_5z3gmTeW9_0),.clk(gclk));
	jdff dff_A_BF8gCdAp4_0(.dout(w_dff_A_5z3gmTeW9_0),.din(w_dff_A_BF8gCdAp4_0),.clk(gclk));
	jdff dff_A_MGDYFj995_1(.dout(w_G8gat_0[1]),.din(w_dff_A_MGDYFj995_1),.clk(gclk));
	jdff dff_A_2T4XnEqm3_1(.dout(w_dff_A_MGDYFj995_1),.din(w_dff_A_2T4XnEqm3_1),.clk(gclk));
	jdff dff_A_Gm0vMFkY0_1(.dout(w_dff_A_2T4XnEqm3_1),.din(w_dff_A_Gm0vMFkY0_1),.clk(gclk));
	jdff dff_A_n64ETrL61_1(.dout(w_dff_A_Gm0vMFkY0_1),.din(w_dff_A_n64ETrL61_1),.clk(gclk));
	jdff dff_A_s1VW2A2j8_1(.dout(w_dff_A_n64ETrL61_1),.din(w_dff_A_s1VW2A2j8_1),.clk(gclk));
	jdff dff_A_mPsWAnai9_1(.dout(w_dff_A_s1VW2A2j8_1),.din(w_dff_A_mPsWAnai9_1),.clk(gclk));
	jdff dff_A_iXdroaPO2_1(.dout(w_dff_A_mPsWAnai9_1),.din(w_dff_A_iXdroaPO2_1),.clk(gclk));
	jdff dff_A_6l4mxBtJ8_1(.dout(w_dff_A_iXdroaPO2_1),.din(w_dff_A_6l4mxBtJ8_1),.clk(gclk));
	jdff dff_A_ZAq4GogY7_0(.dout(w_n96_0[0]),.din(w_dff_A_ZAq4GogY7_0),.clk(gclk));
	jdff dff_A_Zjd3FBVm9_0(.dout(w_dff_A_ZAq4GogY7_0),.din(w_dff_A_Zjd3FBVm9_0),.clk(gclk));
	jdff dff_A_hP8e5VEY4_0(.dout(w_dff_A_Zjd3FBVm9_0),.din(w_dff_A_hP8e5VEY4_0),.clk(gclk));
	jdff dff_A_E5jsua8o5_0(.dout(w_dff_A_hP8e5VEY4_0),.din(w_dff_A_E5jsua8o5_0),.clk(gclk));
	jdff dff_A_x77Iu3pY1_0(.dout(w_dff_A_E5jsua8o5_0),.din(w_dff_A_x77Iu3pY1_0),.clk(gclk));
	jdff dff_A_F1VAy6oj4_0(.dout(w_dff_A_x77Iu3pY1_0),.din(w_dff_A_F1VAy6oj4_0),.clk(gclk));
	jdff dff_B_1g27YgFr7_1(.din(n76),.dout(w_dff_B_1g27YgFr7_1),.clk(gclk));
	jdff dff_B_7jHgBMXL3_1(.din(n81),.dout(w_dff_B_7jHgBMXL3_1),.clk(gclk));
	jdff dff_A_YS5WvG4O8_0(.dout(w_n89_0[0]),.din(w_dff_A_YS5WvG4O8_0),.clk(gclk));
	jdff dff_A_RdscfmSd6_0(.dout(w_dff_A_YS5WvG4O8_0),.din(w_dff_A_RdscfmSd6_0),.clk(gclk));
	jdff dff_A_vs4Yte5a6_0(.dout(w_dff_A_RdscfmSd6_0),.din(w_dff_A_vs4Yte5a6_0),.clk(gclk));
	jdff dff_A_McmLrzke5_0(.dout(w_dff_A_vs4Yte5a6_0),.din(w_dff_A_McmLrzke5_0),.clk(gclk));
	jdff dff_A_TTdqR00b8_0(.dout(w_dff_A_McmLrzke5_0),.din(w_dff_A_TTdqR00b8_0),.clk(gclk));
	jdff dff_A_vcoSxdJH7_0(.dout(w_dff_A_TTdqR00b8_0),.din(w_dff_A_vcoSxdJH7_0),.clk(gclk));
	jdff dff_A_FNBBFI7k1_0(.dout(w_n84_0[0]),.din(w_dff_A_FNBBFI7k1_0),.clk(gclk));
	jdff dff_A_egyvezmP1_0(.dout(w_dff_A_FNBBFI7k1_0),.din(w_dff_A_egyvezmP1_0),.clk(gclk));
	jdff dff_A_KAqRUqc41_0(.dout(w_dff_A_egyvezmP1_0),.din(w_dff_A_KAqRUqc41_0),.clk(gclk));
	jdff dff_A_tNomMc159_0(.dout(w_dff_A_KAqRUqc41_0),.din(w_dff_A_tNomMc159_0),.clk(gclk));
	jdff dff_A_xxDRcru73_0(.dout(w_dff_A_tNomMc159_0),.din(w_dff_A_xxDRcru73_0),.clk(gclk));
	jdff dff_A_t6pyZeN27_0(.dout(w_dff_A_xxDRcru73_0),.din(w_dff_A_t6pyZeN27_0),.clk(gclk));
	jdff dff_A_0tDbL01y9_0(.dout(w_n82_0[0]),.din(w_dff_A_0tDbL01y9_0),.clk(gclk));
	jdff dff_A_QgsUMgbR2_0(.dout(w_dff_A_0tDbL01y9_0),.din(w_dff_A_QgsUMgbR2_0),.clk(gclk));
	jdff dff_A_zSvERz9r7_0(.dout(w_dff_A_QgsUMgbR2_0),.din(w_dff_A_zSvERz9r7_0),.clk(gclk));
	jdff dff_A_D8HQEZDm7_0(.dout(w_dff_A_zSvERz9r7_0),.din(w_dff_A_D8HQEZDm7_0),.clk(gclk));
	jdff dff_A_VUMppq5o2_0(.dout(w_dff_A_D8HQEZDm7_0),.din(w_dff_A_VUMppq5o2_0),.clk(gclk));
	jdff dff_A_PftCV0974_0(.dout(w_dff_A_VUMppq5o2_0),.din(w_dff_A_PftCV0974_0),.clk(gclk));
	jdff dff_A_H77QyUzX6_0(.dout(w_n79_0[0]),.din(w_dff_A_H77QyUzX6_0),.clk(gclk));
	jdff dff_A_ikqDVpKe9_0(.dout(w_dff_A_H77QyUzX6_0),.din(w_dff_A_ikqDVpKe9_0),.clk(gclk));
	jdff dff_A_6IvXc7H93_0(.dout(w_dff_A_ikqDVpKe9_0),.din(w_dff_A_6IvXc7H93_0),.clk(gclk));
	jdff dff_A_IEeZPfcm7_0(.dout(w_dff_A_6IvXc7H93_0),.din(w_dff_A_IEeZPfcm7_0),.clk(gclk));
	jdff dff_A_E3m0gHHM1_0(.dout(w_dff_A_IEeZPfcm7_0),.din(w_dff_A_E3m0gHHM1_0),.clk(gclk));
	jdff dff_A_0iX5VOvF3_0(.dout(w_dff_A_E3m0gHHM1_0),.din(w_dff_A_0iX5VOvF3_0),.clk(gclk));
	jdff dff_A_0KSjwQtd3_0(.dout(w_n78_0[0]),.din(w_dff_A_0KSjwQtd3_0),.clk(gclk));
	jdff dff_A_tJBtmbww6_0(.dout(w_dff_A_0KSjwQtd3_0),.din(w_dff_A_tJBtmbww6_0),.clk(gclk));
	jdff dff_A_KIGRHkPL2_0(.dout(w_dff_A_tJBtmbww6_0),.din(w_dff_A_KIGRHkPL2_0),.clk(gclk));
	jdff dff_A_3oa89vUu6_0(.dout(w_dff_A_KIGRHkPL2_0),.din(w_dff_A_3oa89vUu6_0),.clk(gclk));
	jdff dff_A_CAjglNfV7_0(.dout(w_n77_0[0]),.din(w_dff_A_CAjglNfV7_0),.clk(gclk));
	jdff dff_A_OU2Z0wSZ9_0(.dout(w_dff_A_CAjglNfV7_0),.din(w_dff_A_OU2Z0wSZ9_0),.clk(gclk));
	jdff dff_A_LbP9gmM75_0(.dout(w_dff_A_OU2Z0wSZ9_0),.din(w_dff_A_LbP9gmM75_0),.clk(gclk));
	jdff dff_A_qKygx8oj3_0(.dout(w_dff_A_LbP9gmM75_0),.din(w_dff_A_qKygx8oj3_0),.clk(gclk));
	jdff dff_A_H49QXB351_0(.dout(w_dff_A_qKygx8oj3_0),.din(w_dff_A_H49QXB351_0),.clk(gclk));
	jdff dff_A_DQdR1sTx9_0(.dout(w_dff_A_H49QXB351_0),.din(w_dff_A_DQdR1sTx9_0),.clk(gclk));
	jdff dff_A_0WKc5XU48_0(.dout(w_n73_0[0]),.din(w_dff_A_0WKc5XU48_0),.clk(gclk));
	jdff dff_A_1eDK6lYR9_0(.dout(w_dff_A_0WKc5XU48_0),.din(w_dff_A_1eDK6lYR9_0),.clk(gclk));
	jdff dff_A_b8Ik8HGI4_0(.dout(w_dff_A_1eDK6lYR9_0),.din(w_dff_A_b8Ik8HGI4_0),.clk(gclk));
	jdff dff_A_d4CkhFFo4_0(.dout(w_dff_A_b8Ik8HGI4_0),.din(w_dff_A_d4CkhFFo4_0),.clk(gclk));
	jdff dff_A_Km5hpih89_0(.dout(w_dff_A_d4CkhFFo4_0),.din(w_dff_A_Km5hpih89_0),.clk(gclk));
	jdff dff_A_p5hPemGS8_0(.dout(w_dff_A_Km5hpih89_0),.din(w_dff_A_p5hPemGS8_0),.clk(gclk));
	jdff dff_A_wgydJpYc2_0(.dout(w_n72_0[0]),.din(w_dff_A_wgydJpYc2_0),.clk(gclk));
	jdff dff_A_Fevppzgi7_0(.dout(w_dff_A_wgydJpYc2_0),.din(w_dff_A_Fevppzgi7_0),.clk(gclk));
	jdff dff_A_4rThsRKZ8_0(.dout(w_dff_A_Fevppzgi7_0),.din(w_dff_A_4rThsRKZ8_0),.clk(gclk));
	jdff dff_A_mjNe2c9q6_0(.dout(w_dff_A_4rThsRKZ8_0),.din(w_dff_A_mjNe2c9q6_0),.clk(gclk));
	jdff dff_A_UN8sB5N10_0(.dout(w_n71_0[0]),.din(w_dff_A_UN8sB5N10_0),.clk(gclk));
	jdff dff_A_cQUYckR48_0(.dout(w_dff_A_UN8sB5N10_0),.din(w_dff_A_cQUYckR48_0),.clk(gclk));
	jdff dff_A_vyhN0RL21_0(.dout(w_dff_A_cQUYckR48_0),.din(w_dff_A_vyhN0RL21_0),.clk(gclk));
	jdff dff_A_XmSAc9Y30_0(.dout(w_dff_A_vyhN0RL21_0),.din(w_dff_A_XmSAc9Y30_0),.clk(gclk));
	jdff dff_A_nPf3tF7K5_0(.dout(w_dff_A_XmSAc9Y30_0),.din(w_dff_A_nPf3tF7K5_0),.clk(gclk));
	jdff dff_A_im35mc7u0_0(.dout(w_dff_A_nPf3tF7K5_0),.din(w_dff_A_im35mc7u0_0),.clk(gclk));
	jdff dff_A_ibEiz88q1_0(.dout(w_n69_0[0]),.din(w_dff_A_ibEiz88q1_0),.clk(gclk));
	jdff dff_A_NQDn57kM7_0(.dout(w_dff_A_ibEiz88q1_0),.din(w_dff_A_NQDn57kM7_0),.clk(gclk));
	jdff dff_A_k8AqYqB49_0(.dout(w_dff_A_NQDn57kM7_0),.din(w_dff_A_k8AqYqB49_0),.clk(gclk));
	jdff dff_A_UEpzuz7S1_0(.dout(w_dff_A_k8AqYqB49_0),.din(w_dff_A_UEpzuz7S1_0),.clk(gclk));
	jdff dff_A_9tiFhrMz9_0(.dout(w_dff_A_UEpzuz7S1_0),.din(w_dff_A_9tiFhrMz9_0),.clk(gclk));
	jdff dff_B_N7AGX4IP8_2(.din(n69),.dout(w_dff_B_N7AGX4IP8_2),.clk(gclk));
	jdff dff_B_6G06KosA9_2(.din(w_dff_B_N7AGX4IP8_2),.dout(w_dff_B_6G06KosA9_2),.clk(gclk));
	jdff dff_B_KOAIJrsW4_2(.din(w_dff_B_6G06KosA9_2),.dout(w_dff_B_KOAIJrsW4_2),.clk(gclk));
	jdff dff_B_B4a7me5l3_2(.din(w_dff_B_KOAIJrsW4_2),.dout(w_dff_B_B4a7me5l3_2),.clk(gclk));
	jdff dff_B_fHVpo0DQ5_2(.din(w_dff_B_B4a7me5l3_2),.dout(w_dff_B_fHVpo0DQ5_2),.clk(gclk));
	jdff dff_B_YCdv7NHY3_2(.din(w_dff_B_fHVpo0DQ5_2),.dout(w_dff_B_YCdv7NHY3_2),.clk(gclk));
	jdff dff_B_R69DaiPJ4_2(.din(w_dff_B_YCdv7NHY3_2),.dout(w_dff_B_R69DaiPJ4_2),.clk(gclk));
	jdff dff_A_68eKiuOq4_0(.dout(w_G112gat_0[0]),.din(w_dff_A_68eKiuOq4_0),.clk(gclk));
	jdff dff_A_7s7x76Wm0_0(.dout(w_dff_A_68eKiuOq4_0),.din(w_dff_A_7s7x76Wm0_0),.clk(gclk));
	jdff dff_A_5VbRwkNE8_0(.dout(w_dff_A_7s7x76Wm0_0),.din(w_dff_A_5VbRwkNE8_0),.clk(gclk));
	jdff dff_A_DyW161X97_0(.dout(w_dff_A_5VbRwkNE8_0),.din(w_dff_A_DyW161X97_0),.clk(gclk));
	jdff dff_A_W2PdFSHR5_0(.dout(w_dff_A_DyW161X97_0),.din(w_dff_A_W2PdFSHR5_0),.clk(gclk));
	jdff dff_A_D6w4JkDp7_0(.dout(w_dff_A_W2PdFSHR5_0),.din(w_dff_A_D6w4JkDp7_0),.clk(gclk));
	jdff dff_A_8JH5ryuG1_0(.dout(w_dff_A_D6w4JkDp7_0),.din(w_dff_A_8JH5ryuG1_0),.clk(gclk));
	jdff dff_A_bNWg9gOY3_0(.dout(w_dff_A_8JH5ryuG1_0),.din(w_dff_A_bNWg9gOY3_0),.clk(gclk));
	jdff dff_A_5LwtncGv2_0(.dout(w_dff_A_bNWg9gOY3_0),.din(w_dff_A_5LwtncGv2_0),.clk(gclk));
	jdff dff_A_SY7nT9p57_0(.dout(w_dff_A_5LwtncGv2_0),.din(w_dff_A_SY7nT9p57_0),.clk(gclk));
	jdff dff_A_qDDjToK53_0(.dout(w_dff_A_SY7nT9p57_0),.din(w_dff_A_qDDjToK53_0),.clk(gclk));
	jdff dff_A_MEWjSqDL2_0(.dout(w_dff_A_qDDjToK53_0),.din(w_dff_A_MEWjSqDL2_0),.clk(gclk));
	jdff dff_A_y0ynk3B09_0(.dout(w_dff_A_MEWjSqDL2_0),.din(w_dff_A_y0ynk3B09_0),.clk(gclk));
	jdff dff_A_aPcuxAQt9_1(.dout(w_G112gat_0[1]),.din(w_dff_A_aPcuxAQt9_1),.clk(gclk));
	jdff dff_A_j4NiqdiA4_1(.dout(w_dff_A_aPcuxAQt9_1),.din(w_dff_A_j4NiqdiA4_1),.clk(gclk));
	jdff dff_A_ggz7T9v59_1(.dout(w_dff_A_j4NiqdiA4_1),.din(w_dff_A_ggz7T9v59_1),.clk(gclk));
	jdff dff_A_QceUSftn8_1(.dout(w_dff_A_ggz7T9v59_1),.din(w_dff_A_QceUSftn8_1),.clk(gclk));
	jdff dff_A_q5xRitIL5_1(.dout(w_dff_A_QceUSftn8_1),.din(w_dff_A_q5xRitIL5_1),.clk(gclk));
	jdff dff_A_tXyKoq2u0_1(.dout(w_dff_A_q5xRitIL5_1),.din(w_dff_A_tXyKoq2u0_1),.clk(gclk));
	jdff dff_A_PidPrwjK1_1(.dout(w_dff_A_tXyKoq2u0_1),.din(w_dff_A_PidPrwjK1_1),.clk(gclk));
	jdff dff_A_nAPqZLqT6_1(.dout(w_dff_A_PidPrwjK1_1),.din(w_dff_A_nAPqZLqT6_1),.clk(gclk));
	jdff dff_A_gJ6hF6OQ1_1(.dout(w_n139_0[1]),.din(w_dff_A_gJ6hF6OQ1_1),.clk(gclk));
	jdff dff_A_SqMnunAP0_1(.dout(w_dff_A_gJ6hF6OQ1_1),.din(w_dff_A_SqMnunAP0_1),.clk(gclk));
	jdff dff_A_x8GueNsS5_1(.dout(w_dff_A_SqMnunAP0_1),.din(w_dff_A_x8GueNsS5_1),.clk(gclk));
	jdff dff_A_69bqsicp0_1(.dout(w_dff_A_x8GueNsS5_1),.din(w_dff_A_69bqsicp0_1),.clk(gclk));
	jdff dff_A_VEwuRhUd5_1(.dout(w_dff_A_69bqsicp0_1),.din(w_dff_A_VEwuRhUd5_1),.clk(gclk));
	jdff dff_A_8uzRIjdi1_1(.dout(w_dff_A_VEwuRhUd5_1),.din(w_dff_A_8uzRIjdi1_1),.clk(gclk));
	jdff dff_B_psk07u3V0_1(.din(n50),.dout(w_dff_B_psk07u3V0_1),.clk(gclk));
	jdff dff_B_oqycvCM21_1(.din(n55),.dout(w_dff_B_oqycvCM21_1),.clk(gclk));
	jdff dff_A_MMSOLrkf9_0(.dout(w_G4gat_0[0]),.din(w_dff_A_MMSOLrkf9_0),.clk(gclk));
	jdff dff_A_EmbrQ3OK4_0(.dout(w_dff_A_MMSOLrkf9_0),.din(w_dff_A_EmbrQ3OK4_0),.clk(gclk));
	jdff dff_A_5EwA2DpY9_0(.dout(w_dff_A_EmbrQ3OK4_0),.din(w_dff_A_5EwA2DpY9_0),.clk(gclk));
	jdff dff_A_sSsn89L83_0(.dout(w_dff_A_5EwA2DpY9_0),.din(w_dff_A_sSsn89L83_0),.clk(gclk));
	jdff dff_A_5ABIk3ha6_0(.dout(w_dff_A_sSsn89L83_0),.din(w_dff_A_5ABIk3ha6_0),.clk(gclk));
	jdff dff_A_Rd3Iqsut7_0(.dout(w_dff_A_5ABIk3ha6_0),.din(w_dff_A_Rd3Iqsut7_0),.clk(gclk));
	jdff dff_A_B0KcFS5N3_0(.dout(w_dff_A_Rd3Iqsut7_0),.din(w_dff_A_B0KcFS5N3_0),.clk(gclk));
	jdff dff_A_OXR4KdRt3_2(.dout(w_G4gat_0[2]),.din(w_dff_A_OXR4KdRt3_2),.clk(gclk));
	jdff dff_A_HGZVjoyq2_0(.dout(w_n63_0[0]),.din(w_dff_A_HGZVjoyq2_0),.clk(gclk));
	jdff dff_A_y3JgxNnQ8_0(.dout(w_dff_A_HGZVjoyq2_0),.din(w_dff_A_y3JgxNnQ8_0),.clk(gclk));
	jdff dff_A_xSbHDy8M1_0(.dout(w_dff_A_y3JgxNnQ8_0),.din(w_dff_A_xSbHDy8M1_0),.clk(gclk));
	jdff dff_A_Zh6Zzmpx9_0(.dout(w_dff_A_xSbHDy8M1_0),.din(w_dff_A_Zh6Zzmpx9_0),.clk(gclk));
	jdff dff_A_GHmMaPQz1_0(.dout(w_dff_A_Zh6Zzmpx9_0),.din(w_dff_A_GHmMaPQz1_0),.clk(gclk));
	jdff dff_A_zxg6pJ4q5_0(.dout(w_G1gat_0[0]),.din(w_dff_A_zxg6pJ4q5_0),.clk(gclk));
	jdff dff_A_KlkLvP1s6_0(.dout(w_dff_A_zxg6pJ4q5_0),.din(w_dff_A_KlkLvP1s6_0),.clk(gclk));
	jdff dff_A_l6Ex0cdx4_0(.dout(w_dff_A_KlkLvP1s6_0),.din(w_dff_A_l6Ex0cdx4_0),.clk(gclk));
	jdff dff_A_wQCdnG0t0_0(.dout(w_dff_A_l6Ex0cdx4_0),.din(w_dff_A_wQCdnG0t0_0),.clk(gclk));
	jdff dff_A_unlN3uPJ9_0(.dout(w_dff_A_wQCdnG0t0_0),.din(w_dff_A_unlN3uPJ9_0),.clk(gclk));
	jdff dff_A_qMJdKDQo4_0(.dout(w_dff_A_unlN3uPJ9_0),.din(w_dff_A_qMJdKDQo4_0),.clk(gclk));
	jdff dff_A_A24A1gXq5_1(.dout(w_G1gat_0[1]),.din(w_dff_A_A24A1gXq5_1),.clk(gclk));
	jdff dff_A_poMtGWKM2_0(.dout(w_n61_0[0]),.din(w_dff_A_poMtGWKM2_0),.clk(gclk));
	jdff dff_A_BGrAfOEQ2_0(.dout(w_dff_A_poMtGWKM2_0),.din(w_dff_A_BGrAfOEQ2_0),.clk(gclk));
	jdff dff_A_KOnpoR7X3_0(.dout(w_dff_A_BGrAfOEQ2_0),.din(w_dff_A_KOnpoR7X3_0),.clk(gclk));
	jdff dff_A_xyIwAmPi0_0(.dout(w_dff_A_KOnpoR7X3_0),.din(w_dff_A_xyIwAmPi0_0),.clk(gclk));
	jdff dff_A_0ee1nJSj0_0(.dout(w_dff_A_xyIwAmPi0_0),.din(w_dff_A_0ee1nJSj0_0),.clk(gclk));
	jdff dff_A_mXeuhKAh9_0(.dout(w_G89gat_0[0]),.din(w_dff_A_mXeuhKAh9_0),.clk(gclk));
	jdff dff_A_WiEggLot0_0(.dout(w_dff_A_mXeuhKAh9_0),.din(w_dff_A_WiEggLot0_0),.clk(gclk));
	jdff dff_A_k2SMsEB40_0(.dout(w_dff_A_WiEggLot0_0),.din(w_dff_A_k2SMsEB40_0),.clk(gclk));
	jdff dff_A_Pdt8fVrR5_0(.dout(w_dff_A_k2SMsEB40_0),.din(w_dff_A_Pdt8fVrR5_0),.clk(gclk));
	jdff dff_A_Xslwsn9A7_0(.dout(w_dff_A_Pdt8fVrR5_0),.din(w_dff_A_Xslwsn9A7_0),.clk(gclk));
	jdff dff_A_VTHH7CAn5_0(.dout(w_dff_A_Xslwsn9A7_0),.din(w_dff_A_VTHH7CAn5_0),.clk(gclk));
	jdff dff_A_wx4vqfXc1_1(.dout(w_G89gat_0[1]),.din(w_dff_A_wx4vqfXc1_1),.clk(gclk));
	jdff dff_A_OtuWHIYh9_0(.dout(w_G56gat_0[0]),.din(w_dff_A_OtuWHIYh9_0),.clk(gclk));
	jdff dff_A_CQZXVABP2_0(.dout(w_dff_A_OtuWHIYh9_0),.din(w_dff_A_CQZXVABP2_0),.clk(gclk));
	jdff dff_A_t8svVLG17_0(.dout(w_dff_A_CQZXVABP2_0),.din(w_dff_A_t8svVLG17_0),.clk(gclk));
	jdff dff_A_4DJWQcyM2_0(.dout(w_dff_A_t8svVLG17_0),.din(w_dff_A_4DJWQcyM2_0),.clk(gclk));
	jdff dff_A_Gj9lJwna2_0(.dout(w_dff_A_4DJWQcyM2_0),.din(w_dff_A_Gj9lJwna2_0),.clk(gclk));
	jdff dff_A_fsi7MOdP6_0(.dout(w_dff_A_Gj9lJwna2_0),.din(w_dff_A_fsi7MOdP6_0),.clk(gclk));
	jdff dff_A_MpS27uXT9_0(.dout(w_dff_A_fsi7MOdP6_0),.din(w_dff_A_MpS27uXT9_0),.clk(gclk));
	jdff dff_A_LTw6E6Ql5_2(.dout(w_G56gat_0[2]),.din(w_dff_A_LTw6E6Ql5_2),.clk(gclk));
	jdff dff_A_b7HwALh75_0(.dout(w_n58_0[0]),.din(w_dff_A_b7HwALh75_0),.clk(gclk));
	jdff dff_A_tUTfemSi8_0(.dout(w_dff_A_b7HwALh75_0),.din(w_dff_A_tUTfemSi8_0),.clk(gclk));
	jdff dff_A_1qWtbnpy2_0(.dout(w_dff_A_tUTfemSi8_0),.din(w_dff_A_1qWtbnpy2_0),.clk(gclk));
	jdff dff_A_ZnTlYI2p8_0(.dout(w_dff_A_1qWtbnpy2_0),.din(w_dff_A_ZnTlYI2p8_0),.clk(gclk));
	jdff dff_A_bmwWrFaJ6_0(.dout(w_dff_A_ZnTlYI2p8_0),.din(w_dff_A_bmwWrFaJ6_0),.clk(gclk));
	jdff dff_A_SbywBC6r8_0(.dout(w_G50gat_0[0]),.din(w_dff_A_SbywBC6r8_0),.clk(gclk));
	jdff dff_A_2oG41Q1J2_0(.dout(w_dff_A_SbywBC6r8_0),.din(w_dff_A_2oG41Q1J2_0),.clk(gclk));
	jdff dff_A_368eFpuS7_0(.dout(w_dff_A_2oG41Q1J2_0),.din(w_dff_A_368eFpuS7_0),.clk(gclk));
	jdff dff_A_EeKppYKU2_0(.dout(w_dff_A_368eFpuS7_0),.din(w_dff_A_EeKppYKU2_0),.clk(gclk));
	jdff dff_A_e8Vraddr0_0(.dout(w_dff_A_EeKppYKU2_0),.din(w_dff_A_e8Vraddr0_0),.clk(gclk));
	jdff dff_A_XquBIlvv5_0(.dout(w_dff_A_e8Vraddr0_0),.din(w_dff_A_XquBIlvv5_0),.clk(gclk));
	jdff dff_A_o0bLKkPz9_1(.dout(w_G50gat_0[1]),.din(w_dff_A_o0bLKkPz9_1),.clk(gclk));
	jdff dff_A_sxEaZZfL4_0(.dout(w_G108gat_0[0]),.din(w_dff_A_sxEaZZfL4_0),.clk(gclk));
	jdff dff_A_3uv68hd12_0(.dout(w_dff_A_sxEaZZfL4_0),.din(w_dff_A_3uv68hd12_0),.clk(gclk));
	jdff dff_A_tMi8ojkN1_0(.dout(w_dff_A_3uv68hd12_0),.din(w_dff_A_tMi8ojkN1_0),.clk(gclk));
	jdff dff_A_gOAH3kGN4_0(.dout(w_dff_A_tMi8ojkN1_0),.din(w_dff_A_gOAH3kGN4_0),.clk(gclk));
	jdff dff_A_1NtzMFup5_0(.dout(w_dff_A_gOAH3kGN4_0),.din(w_dff_A_1NtzMFup5_0),.clk(gclk));
	jdff dff_A_saW5UnnJ7_0(.dout(w_dff_A_1NtzMFup5_0),.din(w_dff_A_saW5UnnJ7_0),.clk(gclk));
	jdff dff_A_Z5ttAmgn2_0(.dout(w_dff_A_saW5UnnJ7_0),.din(w_dff_A_Z5ttAmgn2_0),.clk(gclk));
	jdff dff_A_WgCxUncS6_2(.dout(w_G108gat_0[2]),.din(w_dff_A_WgCxUncS6_2),.clk(gclk));
	jdff dff_A_zpHSg7Vy4_0(.dout(w_n56_0[0]),.din(w_dff_A_zpHSg7Vy4_0),.clk(gclk));
	jdff dff_A_LL1rQsT87_0(.dout(w_dff_A_zpHSg7Vy4_0),.din(w_dff_A_LL1rQsT87_0),.clk(gclk));
	jdff dff_A_KVTmalWt2_0(.dout(w_dff_A_LL1rQsT87_0),.din(w_dff_A_KVTmalWt2_0),.clk(gclk));
	jdff dff_A_5OMAOq8G4_0(.dout(w_dff_A_KVTmalWt2_0),.din(w_dff_A_5OMAOq8G4_0),.clk(gclk));
	jdff dff_A_UoMNT9Qa5_0(.dout(w_dff_A_5OMAOq8G4_0),.din(w_dff_A_UoMNT9Qa5_0),.clk(gclk));
	jdff dff_A_C4ohPfNl4_0(.dout(w_G102gat_0[0]),.din(w_dff_A_C4ohPfNl4_0),.clk(gclk));
	jdff dff_A_iUHYDX1B0_0(.dout(w_dff_A_C4ohPfNl4_0),.din(w_dff_A_iUHYDX1B0_0),.clk(gclk));
	jdff dff_A_PWJzbRI75_0(.dout(w_dff_A_iUHYDX1B0_0),.din(w_dff_A_PWJzbRI75_0),.clk(gclk));
	jdff dff_A_2ulqc1dc6_0(.dout(w_dff_A_PWJzbRI75_0),.din(w_dff_A_2ulqc1dc6_0),.clk(gclk));
	jdff dff_A_KjHMfl831_0(.dout(w_dff_A_2ulqc1dc6_0),.din(w_dff_A_KjHMfl831_0),.clk(gclk));
	jdff dff_A_VjTQ0GMX3_0(.dout(w_dff_A_KjHMfl831_0),.din(w_dff_A_VjTQ0GMX3_0),.clk(gclk));
	jdff dff_A_uTzSJXu04_1(.dout(w_G102gat_0[1]),.din(w_dff_A_uTzSJXu04_1),.clk(gclk));
	jdff dff_A_fBEA9jxP0_0(.dout(w_G69gat_0[0]),.din(w_dff_A_fBEA9jxP0_0),.clk(gclk));
	jdff dff_A_OLfa3rfG0_0(.dout(w_dff_A_fBEA9jxP0_0),.din(w_dff_A_OLfa3rfG0_0),.clk(gclk));
	jdff dff_A_5EXQ7Kn36_0(.dout(w_dff_A_OLfa3rfG0_0),.din(w_dff_A_5EXQ7Kn36_0),.clk(gclk));
	jdff dff_A_zK5BxrtN3_0(.dout(w_dff_A_5EXQ7Kn36_0),.din(w_dff_A_zK5BxrtN3_0),.clk(gclk));
	jdff dff_A_isRDBUU88_0(.dout(w_dff_A_zK5BxrtN3_0),.din(w_dff_A_isRDBUU88_0),.clk(gclk));
	jdff dff_A_dvRx08Gc4_0(.dout(w_dff_A_isRDBUU88_0),.din(w_dff_A_dvRx08Gc4_0),.clk(gclk));
	jdff dff_A_Ge8B9hJt4_0(.dout(w_dff_A_dvRx08Gc4_0),.din(w_dff_A_Ge8B9hJt4_0),.clk(gclk));
	jdff dff_A_4g578riZ3_2(.dout(w_G69gat_0[2]),.din(w_dff_A_4g578riZ3_2),.clk(gclk));
	jdff dff_A_BWUVzlYy0_0(.dout(w_n53_0[0]),.din(w_dff_A_BWUVzlYy0_0),.clk(gclk));
	jdff dff_A_iqYffsIx4_0(.dout(w_dff_A_BWUVzlYy0_0),.din(w_dff_A_iqYffsIx4_0),.clk(gclk));
	jdff dff_A_7HGOLgLQ0_0(.dout(w_dff_A_iqYffsIx4_0),.din(w_dff_A_7HGOLgLQ0_0),.clk(gclk));
	jdff dff_A_8un81v9g3_0(.dout(w_dff_A_7HGOLgLQ0_0),.din(w_dff_A_8un81v9g3_0),.clk(gclk));
	jdff dff_A_QQxypFdR7_0(.dout(w_dff_A_8un81v9g3_0),.din(w_dff_A_QQxypFdR7_0),.clk(gclk));
	jdff dff_A_cOVi5QN32_0(.dout(w_G63gat_0[0]),.din(w_dff_A_cOVi5QN32_0),.clk(gclk));
	jdff dff_A_38LifaDN7_0(.dout(w_dff_A_cOVi5QN32_0),.din(w_dff_A_38LifaDN7_0),.clk(gclk));
	jdff dff_A_zy3GkgzL0_0(.dout(w_dff_A_38LifaDN7_0),.din(w_dff_A_zy3GkgzL0_0),.clk(gclk));
	jdff dff_A_VMN1DwnB5_0(.dout(w_dff_A_zy3GkgzL0_0),.din(w_dff_A_VMN1DwnB5_0),.clk(gclk));
	jdff dff_A_IO7KywT24_0(.dout(w_dff_A_VMN1DwnB5_0),.din(w_dff_A_IO7KywT24_0),.clk(gclk));
	jdff dff_A_HZbKt9s03_0(.dout(w_dff_A_IO7KywT24_0),.din(w_dff_A_HZbKt9s03_0),.clk(gclk));
	jdff dff_A_U0O983TN1_1(.dout(w_G63gat_0[1]),.din(w_dff_A_U0O983TN1_1),.clk(gclk));
	jdff dff_A_9XmdiHfa7_0(.dout(w_n52_0[0]),.din(w_dff_A_9XmdiHfa7_0),.clk(gclk));
	jdff dff_A_kxm4TQ1o1_0(.dout(w_dff_A_9XmdiHfa7_0),.din(w_dff_A_kxm4TQ1o1_0),.clk(gclk));
	jdff dff_A_9EIHA2mN8_0(.dout(w_dff_A_kxm4TQ1o1_0),.din(w_dff_A_9EIHA2mN8_0),.clk(gclk));
	jdff dff_A_3ykacEbC4_0(.dout(w_dff_A_9EIHA2mN8_0),.din(w_dff_A_3ykacEbC4_0),.clk(gclk));
	jdff dff_A_wAnMmerE8_1(.dout(w_G43gat_1[1]),.din(w_dff_A_wAnMmerE8_1),.clk(gclk));
	jdff dff_A_xghP78uJ2_1(.dout(w_G43gat_0[1]),.din(w_dff_A_xghP78uJ2_1),.clk(gclk));
	jdff dff_A_Pjmk4a686_2(.dout(w_G43gat_0[2]),.din(w_dff_A_Pjmk4a686_2),.clk(gclk));
	jdff dff_A_rMRatPpU3_0(.dout(w_G37gat_0[0]),.din(w_dff_A_rMRatPpU3_0),.clk(gclk));
	jdff dff_A_vKMgwbGJ8_0(.dout(w_dff_A_rMRatPpU3_0),.din(w_dff_A_vKMgwbGJ8_0),.clk(gclk));
	jdff dff_A_msD5FqKo8_0(.dout(w_dff_A_vKMgwbGJ8_0),.din(w_dff_A_msD5FqKo8_0),.clk(gclk));
	jdff dff_A_9KzMed2U8_0(.dout(w_dff_A_msD5FqKo8_0),.din(w_dff_A_9KzMed2U8_0),.clk(gclk));
	jdff dff_A_baAoJW3O6_0(.dout(w_dff_A_9KzMed2U8_0),.din(w_dff_A_baAoJW3O6_0),.clk(gclk));
	jdff dff_A_N4JjRjiX8_0(.dout(w_dff_A_baAoJW3O6_0),.din(w_dff_A_N4JjRjiX8_0),.clk(gclk));
	jdff dff_A_iK9sgUV75_1(.dout(w_G37gat_0[1]),.din(w_dff_A_iK9sgUV75_1),.clk(gclk));
	jdff dff_A_DbMQvbvi3_0(.dout(w_G17gat_0[0]),.din(w_dff_A_DbMQvbvi3_0),.clk(gclk));
	jdff dff_A_KSeK94Xh3_0(.dout(w_dff_A_DbMQvbvi3_0),.din(w_dff_A_KSeK94Xh3_0),.clk(gclk));
	jdff dff_A_RUCOTxEn2_0(.dout(w_dff_A_KSeK94Xh3_0),.din(w_dff_A_RUCOTxEn2_0),.clk(gclk));
	jdff dff_A_yjFjDUBe5_0(.dout(w_dff_A_RUCOTxEn2_0),.din(w_dff_A_yjFjDUBe5_0),.clk(gclk));
	jdff dff_A_nAqjQpYU9_0(.dout(w_dff_A_yjFjDUBe5_0),.din(w_dff_A_nAqjQpYU9_0),.clk(gclk));
	jdff dff_A_IAVnKPJE6_0(.dout(w_dff_A_nAqjQpYU9_0),.din(w_dff_A_IAVnKPJE6_0),.clk(gclk));
	jdff dff_A_xXeOIwou4_0(.dout(w_dff_A_IAVnKPJE6_0),.din(w_dff_A_xXeOIwou4_0),.clk(gclk));
	jdff dff_A_eny0RcZF5_2(.dout(w_G17gat_0[2]),.din(w_dff_A_eny0RcZF5_2),.clk(gclk));
	jdff dff_A_cjWThgh89_0(.dout(w_n47_0[0]),.din(w_dff_A_cjWThgh89_0),.clk(gclk));
	jdff dff_A_KRiWLSeP7_0(.dout(w_dff_A_cjWThgh89_0),.din(w_dff_A_KRiWLSeP7_0),.clk(gclk));
	jdff dff_A_thtnU7wY1_0(.dout(w_dff_A_KRiWLSeP7_0),.din(w_dff_A_thtnU7wY1_0),.clk(gclk));
	jdff dff_A_PSEeBRYd0_0(.dout(w_dff_A_thtnU7wY1_0),.din(w_dff_A_PSEeBRYd0_0),.clk(gclk));
	jdff dff_A_jrm4zwtG2_0(.dout(w_dff_A_PSEeBRYd0_0),.din(w_dff_A_jrm4zwtG2_0),.clk(gclk));
	jdff dff_A_n9yPRBbA0_0(.dout(w_G11gat_0[0]),.din(w_dff_A_n9yPRBbA0_0),.clk(gclk));
	jdff dff_A_YqfOQ8zT2_0(.dout(w_dff_A_n9yPRBbA0_0),.din(w_dff_A_YqfOQ8zT2_0),.clk(gclk));
	jdff dff_A_s83XpgJt9_0(.dout(w_dff_A_YqfOQ8zT2_0),.din(w_dff_A_s83XpgJt9_0),.clk(gclk));
	jdff dff_A_ZFI4vkSL7_0(.dout(w_dff_A_s83XpgJt9_0),.din(w_dff_A_ZFI4vkSL7_0),.clk(gclk));
	jdff dff_A_mtSJ8G1E7_0(.dout(w_dff_A_ZFI4vkSL7_0),.din(w_dff_A_mtSJ8G1E7_0),.clk(gclk));
	jdff dff_A_MQd5T3JC6_0(.dout(w_dff_A_mtSJ8G1E7_0),.din(w_dff_A_MQd5T3JC6_0),.clk(gclk));
	jdff dff_A_scHdCel47_1(.dout(w_G11gat_0[1]),.din(w_dff_A_scHdCel47_1),.clk(gclk));
	jdff dff_A_vq767C681_1(.dout(w_G30gat_0[1]),.din(w_dff_A_vq767C681_1),.clk(gclk));
	jdff dff_A_8fNpvyNO4_0(.dout(w_G24gat_0[0]),.din(w_dff_A_8fNpvyNO4_0),.clk(gclk));
	jdff dff_A_DMrYvpqC1_1(.dout(w_n44_0[1]),.din(w_dff_A_DMrYvpqC1_1),.clk(gclk));
	jdff dff_A_G8whc0Pr5_1(.dout(w_G82gat_0[1]),.din(w_dff_A_G8whc0Pr5_1),.clk(gclk));
	jdff dff_A_JHlZvLiu2_1(.dout(w_dff_A_G8whc0Pr5_1),.din(w_dff_A_JHlZvLiu2_1),.clk(gclk));
	jdff dff_A_y1wdbJ7V5_1(.dout(w_dff_A_JHlZvLiu2_1),.din(w_dff_A_y1wdbJ7V5_1),.clk(gclk));
	jdff dff_A_RTUJgqj54_1(.dout(w_dff_A_y1wdbJ7V5_1),.din(w_dff_A_RTUJgqj54_1),.clk(gclk));
	jdff dff_A_rZNTymzR4_1(.dout(w_dff_A_RTUJgqj54_1),.din(w_dff_A_rZNTymzR4_1),.clk(gclk));
	jdff dff_A_YrRtR3Ve0_1(.dout(w_dff_A_rZNTymzR4_1),.din(w_dff_A_YrRtR3Ve0_1),.clk(gclk));
	jdff dff_A_7hgsGo9G1_1(.dout(w_dff_A_YrRtR3Ve0_1),.din(w_dff_A_7hgsGo9G1_1),.clk(gclk));
	jdff dff_A_iYOw4pOk9_2(.dout(w_G82gat_0[2]),.din(w_dff_A_iYOw4pOk9_2),.clk(gclk));
	jdff dff_A_a5LUy0Jh0_0(.dout(w_n43_0[0]),.din(w_dff_A_a5LUy0Jh0_0),.clk(gclk));
	jdff dff_A_lmUF8aNa7_0(.dout(w_dff_A_a5LUy0Jh0_0),.din(w_dff_A_lmUF8aNa7_0),.clk(gclk));
	jdff dff_A_9aYZ00BV6_0(.dout(w_dff_A_lmUF8aNa7_0),.din(w_dff_A_9aYZ00BV6_0),.clk(gclk));
	jdff dff_A_58tyhiZ74_0(.dout(w_dff_A_9aYZ00BV6_0),.din(w_dff_A_58tyhiZ74_0),.clk(gclk));
	jdff dff_A_1S6iYLtK3_0(.dout(w_dff_A_58tyhiZ74_0),.din(w_dff_A_1S6iYLtK3_0),.clk(gclk));
	jdff dff_A_kmbyvGTf0_0(.dout(w_G76gat_0[0]),.din(w_dff_A_kmbyvGTf0_0),.clk(gclk));
	jdff dff_A_WsAkDPUO5_0(.dout(w_dff_A_kmbyvGTf0_0),.din(w_dff_A_WsAkDPUO5_0),.clk(gclk));
	jdff dff_A_JODcJSlN7_0(.dout(w_dff_A_WsAkDPUO5_0),.din(w_dff_A_JODcJSlN7_0),.clk(gclk));
	jdff dff_A_RgKDmBCP5_0(.dout(w_dff_A_JODcJSlN7_0),.din(w_dff_A_RgKDmBCP5_0),.clk(gclk));
	jdff dff_A_3N6aZG4V1_0(.dout(w_dff_A_RgKDmBCP5_0),.din(w_dff_A_3N6aZG4V1_0),.clk(gclk));
	jdff dff_A_Z8LXqTPZ1_0(.dout(w_dff_A_3N6aZG4V1_0),.din(w_dff_A_Z8LXqTPZ1_0),.clk(gclk));
	jdff dff_A_PUZJsGRG5_0(.dout(w_n87_0[0]),.din(w_dff_A_PUZJsGRG5_0),.clk(gclk));
	jdff dff_A_Vr9TnkqD2_0(.dout(w_dff_A_PUZJsGRG5_0),.din(w_dff_A_Vr9TnkqD2_0),.clk(gclk));
	jdff dff_A_jdyjcmOa7_0(.dout(w_dff_A_Vr9TnkqD2_0),.din(w_dff_A_jdyjcmOa7_0),.clk(gclk));
	jdff dff_A_E9ik2gEm3_0(.dout(w_dff_A_jdyjcmOa7_0),.din(w_dff_A_E9ik2gEm3_0),.clk(gclk));
	jdff dff_A_g0XFfzZl5_0(.dout(w_dff_A_E9ik2gEm3_0),.din(w_dff_A_g0XFfzZl5_0),.clk(gclk));
	jdff dff_A_st7JVpjz6_0(.dout(w_dff_A_g0XFfzZl5_0),.din(w_dff_A_st7JVpjz6_0),.clk(gclk));
	jdff dff_A_gp6QfW5O2_0(.dout(w_G95gat_0[0]),.din(w_dff_A_gp6QfW5O2_0),.clk(gclk));
	jdff dff_A_retoFnjf2_0(.dout(w_dff_A_gp6QfW5O2_0),.din(w_dff_A_retoFnjf2_0),.clk(gclk));
	jdff dff_A_pN3ggmc15_0(.dout(w_dff_A_retoFnjf2_0),.din(w_dff_A_pN3ggmc15_0),.clk(gclk));
	jdff dff_A_I6MPMl0M1_0(.dout(w_dff_A_pN3ggmc15_0),.din(w_dff_A_I6MPMl0M1_0),.clk(gclk));
	jdff dff_A_j00AEJWg8_0(.dout(w_dff_A_I6MPMl0M1_0),.din(w_dff_A_j00AEJWg8_0),.clk(gclk));
	jdff dff_A_nGIOe9D07_0(.dout(w_dff_A_j00AEJWg8_0),.din(w_dff_A_nGIOe9D07_0),.clk(gclk));
	jdff dff_A_F2J5LdON6_0(.dout(w_dff_A_nGIOe9D07_0),.din(w_dff_A_F2J5LdON6_0),.clk(gclk));
	jdff dff_A_AcISA6RU7_2(.dout(w_G95gat_0[2]),.din(w_dff_A_AcISA6RU7_2),.clk(gclk));
	jdff dff_A_tkBIfQCV9_1(.dout(w_G105gat_0[1]),.din(w_dff_A_tkBIfQCV9_1),.clk(gclk));
	jdff dff_A_YC0wFypt7_1(.dout(w_dff_A_tkBIfQCV9_1),.din(w_dff_A_YC0wFypt7_1),.clk(gclk));
	jdff dff_A_HMT7AyUD1_1(.dout(w_dff_A_YC0wFypt7_1),.din(w_dff_A_HMT7AyUD1_1),.clk(gclk));
	jdff dff_A_rIMszMo84_1(.dout(w_dff_A_HMT7AyUD1_1),.din(w_dff_A_rIMszMo84_1),.clk(gclk));
	jdff dff_A_B6clcUBo2_1(.dout(w_dff_A_rIMszMo84_1),.din(w_dff_A_B6clcUBo2_1),.clk(gclk));
	jdff dff_A_5HP8BIJ01_1(.dout(w_dff_A_B6clcUBo2_1),.din(w_dff_A_5HP8BIJ01_1),.clk(gclk));
	jdff dff_A_fDZDKLkV4_1(.dout(w_dff_A_5HP8BIJ01_1),.din(w_dff_A_fDZDKLkV4_1),.clk(gclk));
	jdff dff_A_y6qefsw96_1(.dout(w_dff_A_fDZDKLkV4_1),.din(w_dff_A_y6qefsw96_1),.clk(gclk));
	jdff dff_A_R2AnmVBV4_1(.dout(w_dff_A_y6qefsw96_1),.din(w_dff_A_R2AnmVBV4_1),.clk(gclk));
	jdff dff_A_lxZPLhBu6_1(.dout(w_dff_A_R2AnmVBV4_1),.din(w_dff_A_lxZPLhBu6_1),.clk(gclk));
	jdff dff_A_KdNP7kkJ2_1(.dout(w_dff_A_lxZPLhBu6_1),.din(w_dff_A_KdNP7kkJ2_1),.clk(gclk));
	jdff dff_A_0Re8soi95_1(.dout(w_dff_A_KdNP7kkJ2_1),.din(w_dff_A_0Re8soi95_1),.clk(gclk));
	jdff dff_A_2gHoIhD52_1(.dout(w_dff_A_0Re8soi95_1),.din(w_dff_A_2gHoIhD52_1),.clk(gclk));
	jdff dff_A_wxwzoTvF1_1(.dout(w_dff_A_2gHoIhD52_1),.din(w_dff_A_wxwzoTvF1_1),.clk(gclk));
	jdff dff_A_PYJI8UMC6_1(.dout(w_dff_A_wxwzoTvF1_1),.din(w_dff_A_PYJI8UMC6_1),.clk(gclk));
	jdff dff_A_MaxiYCp89_2(.dout(w_dff_A_4a1iUSTY4_0),.din(w_dff_A_MaxiYCp89_2),.clk(gclk));
	jdff dff_A_4a1iUSTY4_0(.dout(w_dff_A_RxCxpIGD6_0),.din(w_dff_A_4a1iUSTY4_0),.clk(gclk));
	jdff dff_A_RxCxpIGD6_0(.dout(w_dff_A_QWADezyW3_0),.din(w_dff_A_RxCxpIGD6_0),.clk(gclk));
	jdff dff_A_QWADezyW3_0(.dout(w_dff_A_uL6REXsy7_0),.din(w_dff_A_QWADezyW3_0),.clk(gclk));
	jdff dff_A_uL6REXsy7_0(.dout(w_dff_A_NAzGTNyg9_0),.din(w_dff_A_uL6REXsy7_0),.clk(gclk));
	jdff dff_A_NAzGTNyg9_0(.dout(w_dff_A_G2P8yfdL6_0),.din(w_dff_A_NAzGTNyg9_0),.clk(gclk));
	jdff dff_A_G2P8yfdL6_0(.dout(w_dff_A_auaaU9JO5_0),.din(w_dff_A_G2P8yfdL6_0),.clk(gclk));
	jdff dff_A_auaaU9JO5_0(.dout(w_dff_A_Z928laBU1_0),.din(w_dff_A_auaaU9JO5_0),.clk(gclk));
	jdff dff_A_Z928laBU1_0(.dout(w_dff_A_iTGutd682_0),.din(w_dff_A_Z928laBU1_0),.clk(gclk));
	jdff dff_A_iTGutd682_0(.dout(w_dff_A_h0b9DVmg1_0),.din(w_dff_A_iTGutd682_0),.clk(gclk));
	jdff dff_A_h0b9DVmg1_0(.dout(w_dff_A_7RCADPY52_0),.din(w_dff_A_h0b9DVmg1_0),.clk(gclk));
	jdff dff_A_7RCADPY52_0(.dout(w_dff_A_VWaVx4QM1_0),.din(w_dff_A_7RCADPY52_0),.clk(gclk));
	jdff dff_A_VWaVx4QM1_0(.dout(w_dff_A_51UUfiLp3_0),.din(w_dff_A_VWaVx4QM1_0),.clk(gclk));
	jdff dff_A_51UUfiLp3_0(.dout(w_dff_A_CKJaqjPo3_0),.din(w_dff_A_51UUfiLp3_0),.clk(gclk));
	jdff dff_A_CKJaqjPo3_0(.dout(w_dff_A_sgcmtF7V4_0),.din(w_dff_A_CKJaqjPo3_0),.clk(gclk));
	jdff dff_A_sgcmtF7V4_0(.dout(w_dff_A_okGHrDh63_0),.din(w_dff_A_sgcmtF7V4_0),.clk(gclk));
	jdff dff_A_okGHrDh63_0(.dout(w_dff_A_B9DHgZ8K7_0),.din(w_dff_A_okGHrDh63_0),.clk(gclk));
	jdff dff_A_B9DHgZ8K7_0(.dout(w_dff_A_cjO7Z7sD3_0),.din(w_dff_A_B9DHgZ8K7_0),.clk(gclk));
	jdff dff_A_cjO7Z7sD3_0(.dout(w_dff_A_GlggAXEA0_0),.din(w_dff_A_cjO7Z7sD3_0),.clk(gclk));
	jdff dff_A_GlggAXEA0_0(.dout(G223gat),.din(w_dff_A_GlggAXEA0_0),.clk(gclk));
	jdff dff_A_R3l9X8Gn8_1(.dout(w_dff_A_Gw6NYGQ52_0),.din(w_dff_A_R3l9X8Gn8_1),.clk(gclk));
	jdff dff_A_Gw6NYGQ52_0(.dout(w_dff_A_4ifcTakD8_0),.din(w_dff_A_Gw6NYGQ52_0),.clk(gclk));
	jdff dff_A_4ifcTakD8_0(.dout(w_dff_A_qQXOIv9C2_0),.din(w_dff_A_4ifcTakD8_0),.clk(gclk));
	jdff dff_A_qQXOIv9C2_0(.dout(w_dff_A_BWbWi0ka0_0),.din(w_dff_A_qQXOIv9C2_0),.clk(gclk));
	jdff dff_A_BWbWi0ka0_0(.dout(w_dff_A_w4Gaq2Dg0_0),.din(w_dff_A_BWbWi0ka0_0),.clk(gclk));
	jdff dff_A_w4Gaq2Dg0_0(.dout(w_dff_A_0k8GlC1P6_0),.din(w_dff_A_w4Gaq2Dg0_0),.clk(gclk));
	jdff dff_A_0k8GlC1P6_0(.dout(w_dff_A_QsnA1HsA9_0),.din(w_dff_A_0k8GlC1P6_0),.clk(gclk));
	jdff dff_A_QsnA1HsA9_0(.dout(w_dff_A_FJfEB19U4_0),.din(w_dff_A_QsnA1HsA9_0),.clk(gclk));
	jdff dff_A_FJfEB19U4_0(.dout(w_dff_A_CfF1bmPV9_0),.din(w_dff_A_FJfEB19U4_0),.clk(gclk));
	jdff dff_A_CfF1bmPV9_0(.dout(w_dff_A_4ZYY7OJs4_0),.din(w_dff_A_CfF1bmPV9_0),.clk(gclk));
	jdff dff_A_4ZYY7OJs4_0(.dout(w_dff_A_ALrhgiIh9_0),.din(w_dff_A_4ZYY7OJs4_0),.clk(gclk));
	jdff dff_A_ALrhgiIh9_0(.dout(w_dff_A_zl0zYyGv5_0),.din(w_dff_A_ALrhgiIh9_0),.clk(gclk));
	jdff dff_A_zl0zYyGv5_0(.dout(G329gat),.din(w_dff_A_zl0zYyGv5_0),.clk(gclk));
	jdff dff_A_cgYnHa567_1(.dout(w_dff_A_KJlCgD6r5_0),.din(w_dff_A_cgYnHa567_1),.clk(gclk));
	jdff dff_A_KJlCgD6r5_0(.dout(w_dff_A_FiOshWDZ9_0),.din(w_dff_A_KJlCgD6r5_0),.clk(gclk));
	jdff dff_A_FiOshWDZ9_0(.dout(w_dff_A_wAmORMbX5_0),.din(w_dff_A_FiOshWDZ9_0),.clk(gclk));
	jdff dff_A_wAmORMbX5_0(.dout(w_dff_A_ZswGhIHK6_0),.din(w_dff_A_wAmORMbX5_0),.clk(gclk));
	jdff dff_A_ZswGhIHK6_0(.dout(w_dff_A_vrpEtuVb5_0),.din(w_dff_A_ZswGhIHK6_0),.clk(gclk));
	jdff dff_A_vrpEtuVb5_0(.dout(G370gat),.din(w_dff_A_vrpEtuVb5_0),.clk(gclk));
	jdff dff_A_RCUy6P1j0_1(.dout(w_dff_A_9J82KA3Q7_0),.din(w_dff_A_RCUy6P1j0_1),.clk(gclk));
	jdff dff_A_9J82KA3Q7_0(.dout(G430gat),.din(w_dff_A_9J82KA3Q7_0),.clk(gclk));
endmodule

