/*

c499:
	jxor: 120
	jspl: 54
	jspl3: 64
	jnot: 8
	jcb: 2
	jdff: 405
	jand: 69

Summary:
	jxor: 120
	jspl: 54
	jspl3: 64
	jnot: 8
	jcb: 2
	jdff: 405
	jand: 69
*/

module c499(gclk, Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9, Gid10, Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19, Gid20, Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29, Gid30, Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr, God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10, God11, God12, God13, God14, God15, God16, God17, God18, God19, God20, God21, God22, God23, God24, God25, God26, God27, God28, God29, God30, God31);
	input gclk;
	input Gid0;
	input Gid1;
	input Gid2;
	input Gid3;
	input Gid4;
	input Gid5;
	input Gid6;
	input Gid7;
	input Gid8;
	input Gid9;
	input Gid10;
	input Gid11;
	input Gid12;
	input Gid13;
	input Gid14;
	input Gid15;
	input Gid16;
	input Gid17;
	input Gid18;
	input Gid19;
	input Gid20;
	input Gid21;
	input Gid22;
	input Gid23;
	input Gid24;
	input Gid25;
	input Gid26;
	input Gid27;
	input Gid28;
	input Gid29;
	input Gid30;
	input Gid31;
	input Gic0;
	input Gic1;
	input Gic2;
	input Gic3;
	input Gic4;
	input Gic5;
	input Gic6;
	input Gic7;
	input Gr;
	output God0;
	output God1;
	output God2;
	output God3;
	output God4;
	output God5;
	output God6;
	output God7;
	output God8;
	output God9;
	output God10;
	output God11;
	output God12;
	output God13;
	output God14;
	output God15;
	output God16;
	output God17;
	output God18;
	output God19;
	output God20;
	output God21;
	output God22;
	output God23;
	output God24;
	output God25;
	output God26;
	output God27;
	output God28;
	output God29;
	output God30;
	output God31;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n180;
	wire n182;
	wire n184;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n194;
	wire n196;
	wire n198;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n208;
	wire n210;
	wire n212;
	wire n214;
	wire n215;
	wire n217;
	wire n219;
	wire n221;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n236;
	wire n238;
	wire n240;
	wire n242;
	wire n243;
	wire n244;
	wire n246;
	wire n248;
	wire n250;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n257;
	wire n259;
	wire n261;
	wire n263;
	wire n264;
	wire n266;
	wire n268;
	wire n270;
	wire [2:0] w_Gid0_0;
	wire [2:0] w_Gid1_0;
	wire [2:0] w_Gid2_0;
	wire [2:0] w_Gid3_0;
	wire [2:0] w_Gid4_0;
	wire [2:0] w_Gid5_0;
	wire [2:0] w_Gid6_0;
	wire [2:0] w_Gid7_0;
	wire [2:0] w_Gid8_0;
	wire [2:0] w_Gid9_0;
	wire [2:0] w_Gid10_0;
	wire [2:0] w_Gid11_0;
	wire [2:0] w_Gid12_0;
	wire [2:0] w_Gid13_0;
	wire [2:0] w_Gid14_0;
	wire [2:0] w_Gid15_0;
	wire [2:0] w_Gid16_0;
	wire [2:0] w_Gid17_0;
	wire [2:0] w_Gid18_0;
	wire [2:0] w_Gid19_0;
	wire [2:0] w_Gid20_0;
	wire [2:0] w_Gid21_0;
	wire [2:0] w_Gid22_0;
	wire [2:0] w_Gid23_0;
	wire [2:0] w_Gid24_0;
	wire [2:0] w_Gid25_0;
	wire [2:0] w_Gid26_0;
	wire [2:0] w_Gid27_0;
	wire [2:0] w_Gid28_0;
	wire [2:0] w_Gid29_0;
	wire [2:0] w_Gid30_0;
	wire [2:0] w_Gid31_0;
	wire [2:0] w_Gr_0;
	wire [2:0] w_Gr_1;
	wire [2:0] w_Gr_2;
	wire [1:0] w_Gr_3;
	wire [1:0] w_n75_0;
	wire [1:0] w_n76_0;
	wire [1:0] w_n80_0;
	wire [1:0] w_n83_0;
	wire [1:0] w_n84_0;
	wire [2:0] w_n85_0;
	wire [2:0] w_n85_1;
	wire [1:0] w_n85_2;
	wire [1:0] w_n88_0;
	wire [1:0] w_n89_0;
	wire [1:0] w_n94_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n98_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n110_0;
	wire [2:0] w_n112_0;
	wire [2:0] w_n112_1;
	wire [2:0] w_n112_2;
	wire [1:0] w_n113_0;
	wire [1:0] w_n116_0;
	wire [1:0] w_n117_0;
	wire [2:0] w_n121_0;
	wire [2:0] w_n124_0;
	wire [1:0] w_n125_0;
	wire [2:0] w_n126_0;
	wire [2:0] w_n126_1;
	wire [1:0] w_n126_2;
	wire [1:0] w_n128_0;
	wire [1:0] w_n134_0;
	wire [1:0] w_n135_0;
	wire [1:0] w_n136_0;
	wire [1:0] w_n142_0;
	wire [1:0] w_n143_0;
	wire [2:0] w_n147_0;
	wire [2:0] w_n147_1;
	wire [1:0] w_n147_2;
	wire [2:0] w_n149_0;
	wire [2:0] w_n149_1;
	wire [1:0] w_n149_2;
	wire [1:0] w_n153_0;
	wire [1:0] w_n156_0;
	wire [2:0] w_n159_0;
	wire [2:0] w_n166_0;
	wire [2:0] w_n166_1;
	wire [2:0] w_n166_2;
	wire [1:0] w_n169_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n173_0;
	wire [1:0] w_n174_0;
	wire [1:0] w_n175_0;
	wire [2:0] w_n177_0;
	wire [1:0] w_n177_1;
	wire [2:0] w_n187_0;
	wire [2:0] w_n187_1;
	wire [1:0] w_n187_2;
	wire [1:0] w_n188_0;
	wire [1:0] w_n190_0;
	wire [2:0] w_n191_0;
	wire [1:0] w_n191_1;
	wire [1:0] w_n200_0;
	wire [2:0] w_n202_0;
	wire [2:0] w_n202_1;
	wire [1:0] w_n202_2;
	wire [1:0] w_n203_0;
	wire [2:0] w_n205_0;
	wire [1:0] w_n205_1;
	wire [2:0] w_n214_0;
	wire [1:0] w_n214_1;
	wire [1:0] w_n223_0;
	wire [1:0] w_n231_0;
	wire [1:0] w_n232_0;
	wire [2:0] w_n233_0;
	wire [1:0] w_n233_1;
	wire [1:0] w_n242_0;
	wire [2:0] w_n243_0;
	wire [1:0] w_n243_1;
	wire [1:0] w_n253_0;
	wire [2:0] w_n254_0;
	wire [1:0] w_n254_1;
	wire [2:0] w_n263_0;
	wire [1:0] w_n263_1;
	wire w_dff_A_xsHvLrT50_0;
	wire w_dff_B_A3cqmxTP5_2;
	wire w_dff_A_fHdPikeT7_1;
	wire w_dff_B_KtSH61WO6_2;
	wire w_dff_B_yyxcoOdw6_2;
	wire w_dff_A_CKBUldlp2_0;
	wire w_dff_A_7SxSECa31_0;
	wire w_dff_A_zSMxf2Hg5_0;
	wire w_dff_A_7V5asUu05_0;
	wire w_dff_A_tGSrHpHG2_0;
	wire w_dff_A_JNWAGWUt8_0;
	wire w_dff_A_9gAaidIj4_0;
	wire w_dff_A_kFFQf1lp7_0;
	wire w_dff_A_Uf1PxO8J5_0;
	wire w_dff_A_sxZdp59U5_0;
	wire w_dff_A_m2mR11So6_0;
	wire w_dff_A_xyTxYRt59_0;
	wire w_dff_A_V8stKZ9U4_0;
	wire w_dff_A_G9M1Bjrt0_0;
	wire w_dff_A_6MSWn3oX6_0;
	wire w_dff_A_e8wbs50M9_0;
	wire w_dff_B_b5epyP8x6_1;
	wire w_dff_B_hxqAOgCD5_1;
	wire w_dff_A_4IPXSKR66_0;
	wire w_dff_A_8MGPt5s03_0;
	wire w_dff_A_GjnX3kKg4_0;
	wire w_dff_A_NhYTO4iR6_0;
	wire w_dff_B_Rdj7wqLX1_2;
	wire w_dff_B_HItKXbww1_2;
	wire w_dff_B_gpYsGkyH9_2;
	wire w_dff_A_4a4Bc84i9_0;
	wire w_dff_A_CZswUChP3_0;
	wire w_dff_A_LvEISj5n0_0;
	wire w_dff_A_xrf3zG4d0_0;
	wire w_dff_B_ODVDWLU88_1;
	wire w_dff_B_HOwqrcPC7_1;
	wire w_dff_A_g0O7vAGz7_1;
	wire w_dff_A_Uas4QUmJ3_0;
	wire w_dff_A_AlCXvMgW0_0;
	wire w_dff_A_QeTBLKvK4_0;
	wire w_dff_A_W1E1wB682_0;
	wire w_dff_A_IvdKllUA9_0;
	wire w_dff_A_au9cLAnc1_2;
	wire w_dff_A_iYnrnaLZ9_2;
	wire w_dff_A_c8PAKLHG2_2;
	wire w_dff_A_2fp89xUw1_2;
	wire w_dff_A_I4pFocEd7_2;
	wire w_dff_A_w5AEq2sN0_0;
	wire w_dff_A_AcHISKVu4_0;
	wire w_dff_A_QY6P5fuv9_0;
	wire w_dff_A_MPzX67hC7_0;
	wire w_dff_A_VpyKfITQ2_0;
	wire w_dff_A_AY1ApXn43_0;
	wire w_dff_A_n7uOfbzP8_0;
	wire w_dff_A_irTlR0jg6_2;
	wire w_dff_A_ZshkRoN08_2;
	wire w_dff_A_p3hUBF6k6_2;
	wire w_dff_A_Rvo4aQ0m1_2;
	wire w_dff_A_0YxebjIB7_2;
	wire w_dff_B_b67s7T1b4_0;
	wire w_dff_A_RBghgPVD6_1;
	wire w_dff_A_kuX0xbhN0_0;
	wire w_dff_A_n1bXLGu77_0;
	wire w_dff_A_gFHqnZST6_0;
	wire w_dff_A_lTTVHCoY6_0;
	wire w_dff_A_HsFZPwNr8_0;
	wire w_dff_A_l09FAviz5_2;
	wire w_dff_A_vbRSpGdV3_2;
	wire w_dff_A_NioLwYLQ4_2;
	wire w_dff_A_558Tsuj70_2;
	wire w_dff_A_Fmw23bkx7_2;
	wire w_dff_A_IE9x3CTg7_0;
	wire w_dff_A_UnyKoXRX1_0;
	wire w_dff_A_VjxPrIe00_0;
	wire w_dff_A_m72EqgDs9_0;
	wire w_dff_A_1ZpFomE41_0;
	wire w_dff_A_gale4REy2_0;
	wire w_dff_A_1o9TibeK8_0;
	wire w_dff_A_tqXyFDpb1_0;
	wire w_dff_A_E95DKjEp2_0;
	wire w_dff_A_STeSXPb63_2;
	wire w_dff_A_JHBPrTm53_2;
	wire w_dff_A_NAlJo5TF6_2;
	wire w_dff_A_ClEVmivN9_2;
	wire w_dff_A_m2bEKbcd8_2;
	wire w_dff_B_5CFbhW9H9_0;
	wire w_dff_A_mBSGuVS72_0;
	wire w_dff_A_QdEEbRal4_0;
	wire w_dff_A_NLenSW1i8_0;
	wire w_dff_A_xLUXIChb1_0;
	wire w_dff_A_EYsURZ2f7_1;
	wire w_dff_A_JqDoPysW3_0;
	wire w_dff_A_Osgv8huM7_0;
	wire w_dff_A_EOr20ERz1_0;
	wire w_dff_A_k6MyJVur1_0;
	wire w_dff_A_qKHHdcJL0_0;
	wire w_dff_A_IFo2YrqA7_0;
	wire w_dff_A_paypljLX4_0;
	wire w_dff_A_X3DKZrh94_0;
	wire w_dff_A_pKEIzH8h8_0;
	wire w_dff_A_NQ7akYmb7_0;
	wire w_dff_A_yGMkx7uv1_0;
	wire w_dff_A_mmF43fjx4_0;
	wire w_dff_A_wKmK6h7u6_0;
	wire w_dff_A_4iHz0Oci6_0;
	wire w_dff_A_Cb4wNhcz0_0;
	wire w_dff_A_45CuhMzY4_0;
	wire w_dff_A_A0IBrAuK6_0;
	wire w_dff_A_p0jsRYB00_0;
	wire w_dff_A_MNhKk2F74_0;
	wire w_dff_A_7BOnHrtx5_0;
	wire w_dff_A_JGqyI7v55_0;
	wire w_dff_A_vsUBeMsF1_0;
	wire w_dff_A_QuA8xfCI1_0;
	wire w_dff_A_7U3Kpizm6_0;
	wire w_dff_A_uupUxC8h7_0;
	wire w_dff_A_qhHCfinI9_0;
	wire w_dff_A_zvgLAkvb8_0;
	wire w_dff_A_iGdvqOos6_0;
	wire w_dff_A_WZREt1t41_0;
	wire w_dff_A_12iKLGeb0_0;
	wire w_dff_A_PIwCzpr43_0;
	wire w_dff_A_fS6FLVyQ9_0;
	wire w_dff_A_ckgMQ0re1_0;
	wire w_dff_A_Ev5PtdyW4_0;
	wire w_dff_A_bPLUxzyp2_0;
	wire w_dff_A_kYblhX612_0;
	wire w_dff_A_rDiJ44VL5_1;
	wire w_dff_A_KfdWvmon5_0;
	wire w_dff_A_jynkVs1h9_0;
	wire w_dff_A_oMmIEPNC0_0;
	wire w_dff_A_saxYz4xk3_0;
	wire w_dff_A_7gtcvKQG4_0;
	wire w_dff_A_M1IXzDpf1_0;
	wire w_dff_A_MycwKLCo4_0;
	wire w_dff_A_uULW99Dd9_0;
	wire w_dff_A_6WBKOtYd4_0;
	wire w_dff_A_uYBDJQsx0_0;
	wire w_dff_A_17wcQfLi7_0;
	wire w_dff_A_MZLrsd2A0_0;
	wire w_dff_A_j8hRKf654_0;
	wire w_dff_A_Lvx1syXq2_0;
	wire w_dff_A_cMsqvbT91_0;
	wire w_dff_A_2LmZU9QV5_0;
	wire w_dff_A_bwssEJ8L3_0;
	wire w_dff_A_PJThdGI04_0;
	wire w_dff_A_OvIw5BR05_0;
	wire w_dff_A_TfB7wQkm3_0;
	wire w_dff_A_YJA1BUsx9_0;
	wire w_dff_A_2K0FPSDL4_0;
	wire w_dff_A_4jIbn53j8_0;
	wire w_dff_A_YGDNLoHi8_0;
	wire w_dff_A_zXNrUYCE9_0;
	wire w_dff_A_ijSwMVNU0_0;
	wire w_dff_A_93gcXRbU9_0;
	wire w_dff_A_hnchrOtX1_0;
	wire w_dff_A_9dIQSaS50_0;
	wire w_dff_A_fnQvHc5g1_0;
	wire w_dff_A_OQNCr2cb7_0;
	wire w_dff_A_dtDDVJN91_0;
	wire w_dff_A_f0DVnKwF7_0;
	wire w_dff_A_zi4CwLtO7_0;
	wire w_dff_A_NSwSjxau6_0;
	wire w_dff_A_7GamyOpk3_0;
	wire w_dff_B_e80MwPIa1_2;
	wire w_dff_B_2IKgjRfh7_2;
	wire w_dff_B_b6iKLfib8_2;
	wire w_dff_A_vckJMGo81_0;
	wire w_dff_A_WMI5uizx5_0;
	wire w_dff_A_y44YarSW0_0;
	wire w_dff_A_hWT5mOeY2_0;
	wire w_dff_A_l4byCqB86_0;
	wire w_dff_A_vRzVTpbT1_0;
	wire w_dff_A_q57cKHKq3_0;
	wire w_dff_A_j3IkkGoM5_0;
	wire w_dff_A_OxTmT3AS5_0;
	wire w_dff_A_5ZtQ9U0I5_0;
	wire w_dff_A_BjHxB8iY4_0;
	wire w_dff_A_kwwk4Y7Q9_0;
	wire w_dff_A_2oZjKsiF1_0;
	wire w_dff_A_LRvz497N3_0;
	wire w_dff_A_hGfYqPSD3_0;
	wire w_dff_A_ZiltNOEG8_0;
	wire w_dff_A_Y0ZhjNTM5_0;
	wire w_dff_A_FK4WOMqW0_0;
	wire w_dff_A_PfitI8gt2_0;
	wire w_dff_A_GGF5EFZ77_0;
	wire w_dff_A_WRyZI36C6_0;
	wire w_dff_A_M3ok0lhY9_0;
	wire w_dff_A_QrvOrU8h7_0;
	wire w_dff_A_LzkvNfCv8_0;
	wire w_dff_A_hr3MUg078_0;
	wire w_dff_A_5aET0P1v2_0;
	wire w_dff_A_nsfUXMgG0_0;
	wire w_dff_A_wEhcVPKc8_0;
	wire w_dff_A_GQcfvTwE3_0;
	wire w_dff_A_kwEauIa30_0;
	wire w_dff_A_xgfgeWQi3_0;
	wire w_dff_A_BYJ758UH1_0;
	wire w_dff_A_ueuhK2H97_0;
	wire w_dff_A_kZrjmoxk9_0;
	wire w_dff_A_uUiUz1DW2_0;
	wire w_dff_A_Ht497OWo8_0;
	wire w_dff_A_bZQMNXik2_0;
	wire w_dff_A_NFFpdhEI5_0;
	wire w_dff_A_RratTCgI9_0;
	wire w_dff_A_SqA8iIyR8_0;
	wire w_dff_A_XvLAby8w2_0;
	wire w_dff_A_IzZSqeq37_0;
	wire w_dff_A_PeIOuvWj4_0;
	wire w_dff_A_LAbieiDm0_0;
	wire w_dff_A_NTGyefKH4_0;
	wire w_dff_A_cxzokb8r0_0;
	wire w_dff_A_lJppg1qy9_0;
	wire w_dff_A_sptYYzdo1_0;
	wire w_dff_A_36yoWhlu0_0;
	wire w_dff_A_bMPtmkj41_0;
	wire w_dff_A_OdnjyUWN7_0;
	wire w_dff_A_ViKR0alW7_0;
	wire w_dff_A_OshFL5VS7_0;
	wire w_dff_A_21SCxWw11_0;
	wire w_dff_A_R5QegjHs6_0;
	wire w_dff_A_xcMew2LF5_0;
	wire w_dff_A_UZLJxiZ92_0;
	wire w_dff_A_yGtNHZTt5_0;
	wire w_dff_A_5Hmc8qTS5_0;
	wire w_dff_A_HSfLxjnM0_0;
	wire w_dff_A_WEFi1sWc6_0;
	wire w_dff_A_GncTWl2v3_0;
	wire w_dff_A_SpIEUzqS6_0;
	wire w_dff_A_RzSmkcoq7_0;
	wire w_dff_A_QtWbALBo5_0;
	wire w_dff_A_l7GTsDaa6_0;
	wire w_dff_A_Gg8XAR6R1_0;
	wire w_dff_A_QGGOFcGh8_0;
	wire w_dff_A_Ob80NA3b3_0;
	wire w_dff_A_8NJVnrL29_0;
	wire w_dff_A_Jzk2lz6J8_0;
	wire w_dff_A_ZLpKlT7Z7_0;
	wire w_dff_A_4OF9DJmF6_0;
	wire w_dff_A_CRAKeGGg2_0;
	wire w_dff_A_Wd6H7ox35_0;
	wire w_dff_A_4jr6RA0o0_0;
	wire w_dff_A_xLN5Qrlm2_0;
	wire w_dff_A_bP53vWSx8_0;
	wire w_dff_A_IloUHykN1_0;
	wire w_dff_A_moLtcGR57_0;
	wire w_dff_A_t7ggL07M9_0;
	wire w_dff_A_e0fZImGb1_0;
	wire w_dff_A_3QArWJJ35_0;
	wire w_dff_A_LMQccdJI8_0;
	wire w_dff_A_WV1roGcV3_0;
	wire w_dff_A_nfBAd0vj7_0;
	wire w_dff_A_lr4aCgXD3_0;
	wire w_dff_A_OCxnHt0k2_0;
	wire w_dff_A_Ev8pmVTN3_0;
	wire w_dff_A_hpAXw5dq3_0;
	wire w_dff_A_P9SqZ6Dj1_0;
	wire w_dff_A_C2Zl8j0U1_0;
	wire w_dff_A_CCABDGb92_0;
	wire w_dff_A_vWFFI2sx1_0;
	wire w_dff_A_bu5TOsZt2_0;
	wire w_dff_A_tteQgkbb5_0;
	wire w_dff_A_OQpiXoZq8_0;
	wire w_dff_A_yTlHa0bX0_0;
	wire w_dff_A_gPILNSDl6_0;
	wire w_dff_A_dTmzHv8y4_0;
	wire w_dff_A_f0UrF91r0_0;
	wire w_dff_A_rImIxOdU1_0;
	wire w_dff_A_DjH3obNe1_0;
	wire w_dff_A_CxycXzxt1_0;
	wire w_dff_A_ML2TD4h34_0;
	wire w_dff_A_PQ0Bq5HP4_0;
	wire w_dff_A_Bw250faj5_0;
	wire w_dff_A_Sl5E2Pss5_0;
	wire w_dff_A_xeROUAR32_0;
	wire w_dff_A_YOnF9Tbd0_0;
	wire w_dff_A_8bpDb2Qn9_0;
	wire w_dff_A_kHptG9EG0_0;
	wire w_dff_A_WRxhgMmC5_0;
	wire w_dff_A_DR6DxE9H1_0;
	wire w_dff_A_kLC6An7A8_0;
	wire w_dff_A_CNYpowAY2_0;
	wire w_dff_A_uuZuWW9G7_0;
	wire w_dff_A_ScXyqwmk5_0;
	wire w_dff_A_SMZUDPL52_0;
	wire w_dff_A_iJjnMfHd3_0;
	wire w_dff_A_Lke3J96z3_0;
	wire w_dff_A_fK9NmEFj1_0;
	wire w_dff_A_1Z8L5Wlo4_0;
	wire w_dff_A_qtPiHYIZ1_0;
	wire w_dff_A_GxhtbElV1_0;
	wire w_dff_A_4tSPT4ae0_0;
	wire w_dff_A_ShVlouA69_0;
	wire w_dff_A_HGrhehqR4_0;
	wire w_dff_A_yU5J5xKF7_0;
	wire w_dff_A_wW1QB6Ip8_0;
	wire w_dff_A_4eesJBAX1_0;
	wire w_dff_A_MvUKGEpP6_0;
	wire w_dff_A_CtIGVonJ4_0;
	wire w_dff_A_in8dp6GF0_0;
	wire w_dff_A_6GlIiAI46_0;
	wire w_dff_A_n2YyPnyt8_0;
	wire w_dff_A_8PAiNZnn2_0;
	wire w_dff_A_5ukHwWHE2_0;
	wire w_dff_A_fXFBxHfN8_0;
	wire w_dff_A_2xJHH95p7_0;
	wire w_dff_A_GW7inNXo9_0;
	wire w_dff_A_CIWDgkaH6_0;
	wire w_dff_A_EEZ76ch47_0;
	wire w_dff_A_XfsGqQgH9_0;
	wire w_dff_A_hP9CgISz6_0;
	wire w_dff_A_59J9n2YU4_0;
	wire w_dff_A_7Qkv7wzY2_0;
	wire w_dff_A_W47mm7Ai1_0;
	wire w_dff_A_dmj8I8wf4_0;
	wire w_dff_A_B7KuEblU4_0;
	wire w_dff_A_ZOKuz7Gy1_0;
	wire w_dff_A_6BDMHWkN3_0;
	wire w_dff_A_78wyfkzn7_0;
	wire w_dff_A_g81HgcgD1_0;
	wire w_dff_A_Uc3xER899_0;
	wire w_dff_A_f5HW29mj7_0;
	wire w_dff_A_9ho4Nn9t4_0;
	wire w_dff_A_WCTX8HK26_0;
	wire w_dff_A_fQt3MjJe2_0;
	wire w_dff_A_v9K8nSWP6_0;
	wire w_dff_A_qkUgSe8V2_0;
	wire w_dff_A_NwUPZEmv6_0;
	wire w_dff_A_vwV6qDiY0_0;
	wire w_dff_A_UePXeYo52_0;
	wire w_dff_A_90vmAjC44_0;
	wire w_dff_A_SV73FUkl9_0;
	wire w_dff_A_hoRlUHJb5_0;
	wire w_dff_A_XAjfJZzc0_0;
	wire w_dff_A_LvdBae3g4_0;
	wire w_dff_A_A0Gs43go1_0;
	wire w_dff_A_B0JUY8yP9_0;
	wire w_dff_A_URhjdKHN2_0;
	wire w_dff_A_LCjiDUSI8_0;
	wire w_dff_A_ANmPxrNb0_0;
	wire w_dff_A_NWEpgtfT4_0;
	wire w_dff_A_ZyKiFDdL6_0;
	wire w_dff_A_aElP0Gp81_0;
	wire w_dff_A_pHA9rxW93_0;
	wire w_dff_A_niuqIfuV8_0;
	wire w_dff_A_nKKuTyWB0_0;
	wire w_dff_A_S6Ku3KxG9_0;
	wire w_dff_A_iJEMv04R5_0;
	wire w_dff_A_BHGmYrIy3_0;
	wire w_dff_A_U7zZCN2Q6_0;
	wire w_dff_A_lJjb7aA84_0;
	wire w_dff_A_jvnZxQgd4_0;
	wire w_dff_A_13P3eB4r7_0;
	wire w_dff_A_NNrpbb4M1_0;
	wire w_dff_A_EH4UGlAo3_0;
	wire w_dff_A_4488NkMZ3_0;
	wire w_dff_A_MOmIMwaP9_0;
	wire w_dff_A_4wZLjRTf5_0;
	wire w_dff_A_64vW8LYs2_0;
	wire w_dff_A_T6SZeMnp1_0;
	wire w_dff_A_muIWvRze2_0;
	wire w_dff_A_es3LB2bb6_0;
	wire w_dff_A_O6iHzNyD7_0;
	wire w_dff_A_6ozCoOJb2_0;
	wire w_dff_A_Rv2ewegQ6_0;
	wire w_dff_A_OR6pGGhO9_0;
	wire w_dff_A_q9qdLaP40_0;
	wire w_dff_A_OLbfuIra7_0;
	wire w_dff_A_HIJJWWz61_0;
	wire w_dff_A_LT7ZlOYt8_0;
	wire w_dff_A_t6ipZzDX6_0;
	wire w_dff_A_DQCSUQqG6_0;
	wire w_dff_A_svqLrh3p5_0;
	wire w_dff_A_GkSNTNLK1_0;
	wire w_dff_A_smRNJj5V0_0;
	wire w_dff_A_g7AvD1lU2_0;
	wire w_dff_A_MXBC8gwc7_0;
	wire w_dff_A_XXgimxdL0_0;
	wire w_dff_A_BOD9uQUq4_0;
	wire w_dff_A_nkiiWIQD4_0;
	wire w_dff_A_y59Z0jRU0_0;
	wire w_dff_A_pFiZV1U81_0;
	wire w_dff_A_WBkR5y0F6_0;
	wire w_dff_A_D5KmenKw5_0;
	wire w_dff_A_GQ9VcaOp6_0;
	wire w_dff_A_p1WKOqjt3_0;
	wire w_dff_A_4lo1HaQU6_0;
	wire w_dff_A_6V26NkQY9_0;
	wire w_dff_A_tSQ47dtz9_0;
	wire w_dff_A_aebaVOIH5_0;
	wire w_dff_A_H2K6atbm7_0;
	wire w_dff_A_JLCdQGQ26_0;
	wire w_dff_A_vodje6d04_0;
	wire w_dff_A_PDVxLHao2_0;
	wire w_dff_A_73iZggXs5_0;
	wire w_dff_A_moRPC7wp3_0;
	wire w_dff_A_Mp2833Jr3_0;
	wire w_dff_A_TcFPoXcA1_0;
	wire w_dff_A_VIYnC5J50_0;
	wire w_dff_A_2Z9XcLd81_0;
	wire w_dff_A_odOsKShW0_0;
	wire w_dff_A_gAk31LJm6_0;
	wire w_dff_A_OMF8t8vb2_0;
	wire w_dff_A_QfoNNBsi3_0;
	jxor g000(.dina(w_Gid12_0[2]),.dinb(w_Gid8_0[2]),.dout(n73),.clk(gclk));
	jxor g001(.dina(w_Gid4_0[2]),.dinb(w_Gid0_0[2]),.dout(n74),.clk(gclk));
	jxor g002(.dina(n74),.dinb(n73),.dout(n75),.clk(gclk));
	jand g003(.dina(w_Gr_3[1]),.dinb(Gic0),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_n76_0[1]),.dinb(w_n75_0[1]),.dout(n77),.clk(gclk));
	jxor g005(.dina(w_Gid19_0[2]),.dinb(w_Gid18_0[2]),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_Gid17_0[2]),.dinb(w_Gid16_0[2]),.dout(n79),.clk(gclk));
	jxor g007(.dina(n79),.dinb(n78),.dout(n80),.clk(gclk));
	jxor g008(.dina(w_Gid23_0[2]),.dinb(w_Gid22_0[2]),.dout(n81),.clk(gclk));
	jxor g009(.dina(w_Gid21_0[2]),.dinb(w_Gid20_0[2]),.dout(n82),.clk(gclk));
	jxor g010(.dina(n82),.dinb(n81),.dout(n83),.clk(gclk));
	jxor g011(.dina(w_n83_0[1]),.dinb(w_n80_0[1]),.dout(n84),.clk(gclk));
	jxor g012(.dina(w_n84_0[1]),.dinb(n77),.dout(n85),.clk(gclk));
	jxor g013(.dina(w_Gid31_0[2]),.dinb(w_Gid27_0[2]),.dout(n86),.clk(gclk));
	jxor g014(.dina(w_Gid23_0[1]),.dinb(w_Gid19_0[1]),.dout(n87),.clk(gclk));
	jxor g015(.dina(n87),.dinb(n86),.dout(n88),.clk(gclk));
	jand g016(.dina(w_Gr_3[0]),.dinb(Gic7),.dout(n89),.clk(gclk));
	jnot g017(.din(w_n89_0[1]),.dout(n90),.clk(gclk));
	jxor g018(.dina(n90),.dinb(w_n88_0[1]),.dout(n91),.clk(gclk));
	jxor g019(.dina(w_Gid7_0[2]),.dinb(w_Gid6_0[2]),.dout(n92),.clk(gclk));
	jxor g020(.dina(w_Gid5_0[2]),.dinb(w_Gid4_0[1]),.dout(n93),.clk(gclk));
	jxor g021(.dina(n93),.dinb(n92),.dout(n94),.clk(gclk));
	jxor g022(.dina(w_Gid15_0[2]),.dinb(w_Gid14_0[2]),.dout(n95),.clk(gclk));
	jxor g023(.dina(w_Gid13_0[2]),.dinb(w_Gid12_0[1]),.dout(n96),.clk(gclk));
	jxor g024(.dina(n96),.dinb(n95),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_n97_0[1]),.dinb(w_n94_0[1]),.dout(n98),.clk(gclk));
	jxor g026(.dina(w_n98_0[1]),.dinb(n91),.dout(n99),.clk(gclk));
	jxor g027(.dina(w_Gid30_0[2]),.dinb(w_Gid26_0[2]),.dout(n100),.clk(gclk));
	jxor g028(.dina(w_Gid22_0[1]),.dinb(w_Gid18_0[1]),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n100),.dout(n102),.clk(gclk));
	jand g030(.dina(w_Gr_2[2]),.dinb(Gic6),.dout(n103),.clk(gclk));
	jxor g031(.dina(w_dff_B_b67s7T1b4_0),.dinb(n102),.dout(n104),.clk(gclk));
	jxor g032(.dina(w_Gid3_0[2]),.dinb(w_Gid2_0[2]),.dout(n105),.clk(gclk));
	jxor g033(.dina(w_Gid1_0[2]),.dinb(w_Gid0_0[1]),.dout(n106),.clk(gclk));
	jxor g034(.dina(n106),.dinb(n105),.dout(n107),.clk(gclk));
	jxor g035(.dina(w_Gid11_0[2]),.dinb(w_Gid10_0[2]),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_Gid9_0[2]),.dinb(w_Gid8_0[1]),.dout(n109),.clk(gclk));
	jxor g037(.dina(n109),.dinb(n108),.dout(n110),.clk(gclk));
	jxor g038(.dina(w_n110_0[1]),.dinb(w_n107_0[1]),.dout(n111),.clk(gclk));
	jxor g039(.dina(n111),.dinb(n104),.dout(n112),.clk(gclk));
	jand g040(.dina(w_n112_2[2]),.dinb(w_n99_0[1]),.dout(n113),.clk(gclk));
	jxor g041(.dina(w_Gid13_0[1]),.dinb(w_Gid9_0[1]),.dout(n114),.clk(gclk));
	jxor g042(.dina(w_Gid5_0[1]),.dinb(w_Gid1_0[1]),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(n114),.dout(n116),.clk(gclk));
	jand g044(.dina(w_Gr_2[1]),.dinb(Gic1),.dout(n117),.clk(gclk));
	jxor g045(.dina(w_n117_0[1]),.dinb(w_n116_0[1]),.dout(n118),.clk(gclk));
	jxor g046(.dina(w_Gid31_0[1]),.dinb(w_Gid30_0[1]),.dout(n119),.clk(gclk));
	jxor g047(.dina(w_Gid29_0[2]),.dinb(w_Gid28_0[2]),.dout(n120),.clk(gclk));
	jxor g048(.dina(n120),.dinb(n119),.dout(n121),.clk(gclk));
	jxor g049(.dina(w_Gid27_0[1]),.dinb(w_Gid26_0[1]),.dout(n122),.clk(gclk));
	jxor g050(.dina(w_Gid25_0[2]),.dinb(w_Gid24_0[2]),.dout(n123),.clk(gclk));
	jxor g051(.dina(n123),.dinb(n122),.dout(n124),.clk(gclk));
	jxor g052(.dina(w_n124_0[2]),.dinb(w_n121_0[2]),.dout(n125),.clk(gclk));
	jxor g053(.dina(w_n125_0[1]),.dinb(n118),.dout(n126),.clk(gclk));
	jxor g054(.dina(w_n126_2[1]),.dinb(w_n85_2[1]),.dout(n127),.clk(gclk));
	jand g055(.dina(w_Gr_2[0]),.dinb(Gic3),.dout(n128),.clk(gclk));
	jnot g056(.din(w_n128_0[1]),.dout(n129),.clk(gclk));
	jxor g057(.dina(n129),.dinb(w_n121_0[1]),.dout(n130),.clk(gclk));
	jxor g058(.dina(w_Gid15_0[1]),.dinb(w_Gid11_0[1]),.dout(n131),.clk(gclk));
	jxor g059(.dina(w_Gid7_0[1]),.dinb(w_Gid3_0[1]),.dout(n132),.clk(gclk));
	jxor g060(.dina(n132),.dinb(n131),.dout(n133),.clk(gclk));
	jxor g061(.dina(n133),.dinb(w_n83_0[0]),.dout(n134),.clk(gclk));
	jxor g062(.dina(w_n134_0[1]),.dinb(n130),.dout(n135),.clk(gclk));
	jand g063(.dina(w_Gr_1[2]),.dinb(Gic2),.dout(n136),.clk(gclk));
	jnot g064(.din(w_n136_0[1]),.dout(n137),.clk(gclk));
	jxor g065(.dina(n137),.dinb(w_n124_0[1]),.dout(n138),.clk(gclk));
	jxor g066(.dina(w_Gid14_0[1]),.dinb(w_Gid10_0[1]),.dout(n139),.clk(gclk));
	jxor g067(.dina(w_Gid6_0[1]),.dinb(w_Gid2_0[1]),.dout(n140),.clk(gclk));
	jxor g068(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g069(.dina(n141),.dinb(w_n80_0[0]),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_n142_0[1]),.dinb(n138),.dout(n143),.clk(gclk));
	jand g071(.dina(w_n143_0[1]),.dinb(w_n135_0[1]),.dout(n144),.clk(gclk));
	jand g072(.dina(n144),.dinb(n127),.dout(n145),.clk(gclk));
	jxor g073(.dina(w_n128_0[0]),.dinb(w_n121_0[0]),.dout(n146),.clk(gclk));
	jxor g074(.dina(w_n134_0[0]),.dinb(n146),.dout(n147),.clk(gclk));
	jxor g075(.dina(w_n136_0[0]),.dinb(w_n124_0[0]),.dout(n148),.clk(gclk));
	jxor g076(.dina(w_n142_0[0]),.dinb(n148),.dout(n149),.clk(gclk));
	jxor g077(.dina(w_n149_2[1]),.dinb(w_n147_2[1]),.dout(n150),.clk(gclk));
	jnot g078(.din(w_n76_0[0]),.dout(n151),.clk(gclk));
	jxor g079(.dina(n151),.dinb(w_n75_0[0]),.dout(n152),.clk(gclk));
	jxor g080(.dina(w_n84_0[0]),.dinb(n152),.dout(n153),.clk(gclk));
	jnot g081(.din(w_n117_0[0]),.dout(n154),.clk(gclk));
	jxor g082(.dina(n154),.dinb(w_n116_0[0]),.dout(n155),.clk(gclk));
	jxor g083(.dina(w_n125_0[0]),.dinb(n155),.dout(n156),.clk(gclk));
	jand g084(.dina(w_n156_0[1]),.dinb(w_n153_0[1]),.dout(n157),.clk(gclk));
	jand g085(.dina(n157),.dinb(n150),.dout(n158),.clk(gclk));
	jcb g086(.dina(n158),.dinb(n145),.dout(n159));
	jxor g087(.dina(w_Gid28_0[1]),.dinb(w_Gid24_0[1]),.dout(n160),.clk(gclk));
	jxor g088(.dina(w_Gid20_0[1]),.dinb(w_Gid16_0[1]),.dout(n161),.clk(gclk));
	jxor g089(.dina(n161),.dinb(n160),.dout(n162),.clk(gclk));
	jand g090(.dina(w_Gr_1[1]),.dinb(Gic4),.dout(n163),.clk(gclk));
	jxor g091(.dina(w_dff_B_5CFbhW9H9_0),.dinb(n162),.dout(n164),.clk(gclk));
	jxor g092(.dina(w_n107_0[0]),.dinb(w_n94_0[0]),.dout(n165),.clk(gclk));
	jxor g093(.dina(n165),.dinb(n164),.dout(n166),.clk(gclk));
	jxor g094(.dina(w_Gid29_0[1]),.dinb(w_Gid25_0[1]),.dout(n167),.clk(gclk));
	jxor g095(.dina(w_Gid21_0[1]),.dinb(w_Gid17_0[1]),.dout(n168),.clk(gclk));
	jxor g096(.dina(n168),.dinb(n167),.dout(n169),.clk(gclk));
	jand g097(.dina(w_Gr_1[0]),.dinb(Gic5),.dout(n170),.clk(gclk));
	jnot g098(.din(w_n170_0[1]),.dout(n171),.clk(gclk));
	jxor g099(.dina(n171),.dinb(w_n169_0[1]),.dout(n172),.clk(gclk));
	jxor g100(.dina(w_n110_0[0]),.dinb(w_n97_0[0]),.dout(n173),.clk(gclk));
	jxor g101(.dina(w_n173_0[1]),.dinb(n172),.dout(n174),.clk(gclk));
	jand g102(.dina(w_n174_0[1]),.dinb(w_n166_2[2]),.dout(n175),.clk(gclk));
	jand g103(.dina(w_n175_0[1]),.dinb(w_n159_0[2]),.dout(n176),.clk(gclk));
	jand g104(.dina(n176),.dinb(w_n113_0[1]),.dout(n177),.clk(gclk));
	jand g105(.dina(w_n177_1[1]),.dinb(w_n85_2[0]),.dout(n178),.clk(gclk));
	jxor g106(.dina(n178),.dinb(w_Gid0_0[0]),.dout(God0),.clk(gclk));
	jand g107(.dina(w_n177_1[0]),.dinb(w_n126_2[0]),.dout(n180),.clk(gclk));
	jxor g108(.dina(n180),.dinb(w_Gid1_0[0]),.dout(God1),.clk(gclk));
	jand g109(.dina(w_n177_0[2]),.dinb(w_n149_2[0]),.dout(n182),.clk(gclk));
	jxor g110(.dina(n182),.dinb(w_Gid2_0[0]),.dout(God2),.clk(gclk));
	jand g111(.dina(w_n177_0[1]),.dinb(w_n147_2[0]),.dout(n184),.clk(gclk));
	jxor g112(.dina(n184),.dinb(w_Gid3_0[0]),.dout(God3),.clk(gclk));
	jxor g113(.dina(w_n89_0[0]),.dinb(w_n88_0[0]),.dout(n186),.clk(gclk));
	jxor g114(.dina(w_n98_0[0]),.dinb(n186),.dout(n187),.clk(gclk));
	jnot g115(.din(w_n112_2[1]),.dout(n188),.clk(gclk));
	jand g116(.dina(w_n188_0[1]),.dinb(w_n187_2[1]),.dout(n189),.clk(gclk));
	jand g117(.dina(n189),.dinb(w_n159_0[1]),.dout(n190),.clk(gclk));
	jand g118(.dina(w_n190_0[1]),.dinb(w_n175_0[0]),.dout(n191),.clk(gclk));
	jand g119(.dina(w_n191_1[1]),.dinb(w_n85_1[2]),.dout(n192),.clk(gclk));
	jxor g120(.dina(n192),.dinb(w_Gid4_0[0]),.dout(God4),.clk(gclk));
	jand g121(.dina(w_n191_1[0]),.dinb(w_n126_1[2]),.dout(n194),.clk(gclk));
	jxor g122(.dina(n194),.dinb(w_Gid5_0[0]),.dout(God5),.clk(gclk));
	jand g123(.dina(w_n191_0[2]),.dinb(w_n149_1[2]),.dout(n196),.clk(gclk));
	jxor g124(.dina(n196),.dinb(w_Gid6_0[0]),.dout(God6),.clk(gclk));
	jand g125(.dina(w_n191_0[1]),.dinb(w_n147_1[2]),.dout(n198),.clk(gclk));
	jxor g126(.dina(n198),.dinb(w_Gid7_0[0]),.dout(God7),.clk(gclk));
	jnot g127(.din(w_n166_2[1]),.dout(n200),.clk(gclk));
	jxor g128(.dina(w_n170_0[0]),.dinb(w_n169_0[0]),.dout(n201),.clk(gclk));
	jxor g129(.dina(w_n173_0[0]),.dinb(n201),.dout(n202),.clk(gclk));
	jand g130(.dina(w_n202_2[1]),.dinb(w_n200_0[1]),.dout(n203),.clk(gclk));
	jand g131(.dina(w_n159_0[0]),.dinb(w_n113_0[0]),.dout(n204),.clk(gclk));
	jand g132(.dina(n204),.dinb(w_n203_0[1]),.dout(n205),.clk(gclk));
	jand g133(.dina(w_n205_1[1]),.dinb(w_n85_1[1]),.dout(n206),.clk(gclk));
	jxor g134(.dina(n206),.dinb(w_Gid8_0[0]),.dout(God8),.clk(gclk));
	jand g135(.dina(w_n205_1[0]),.dinb(w_n126_1[1]),.dout(n208),.clk(gclk));
	jxor g136(.dina(n208),.dinb(w_Gid9_0[0]),.dout(God9),.clk(gclk));
	jand g137(.dina(w_n205_0[2]),.dinb(w_n149_1[1]),.dout(n210),.clk(gclk));
	jxor g138(.dina(n210),.dinb(w_Gid10_0[0]),.dout(God10),.clk(gclk));
	jand g139(.dina(w_n205_0[1]),.dinb(w_n147_1[1]),.dout(n212),.clk(gclk));
	jxor g140(.dina(n212),.dinb(w_Gid11_0[0]),.dout(God11),.clk(gclk));
	jand g141(.dina(w_n203_0[0]),.dinb(w_n190_0[0]),.dout(n214),.clk(gclk));
	jand g142(.dina(w_n214_1[1]),.dinb(w_n85_1[0]),.dout(n215),.clk(gclk));
	jxor g143(.dina(n215),.dinb(w_Gid12_0[0]),.dout(God12),.clk(gclk));
	jand g144(.dina(w_n214_1[0]),.dinb(w_n126_1[0]),.dout(n217),.clk(gclk));
	jxor g145(.dina(n217),.dinb(w_Gid13_0[0]),.dout(God13),.clk(gclk));
	jand g146(.dina(w_n214_0[2]),.dinb(w_n149_1[0]),.dout(n219),.clk(gclk));
	jxor g147(.dina(n219),.dinb(w_Gid14_0[0]),.dout(God14),.clk(gclk));
	jand g148(.dina(w_n214_0[1]),.dinb(w_n147_1[0]),.dout(n221),.clk(gclk));
	jxor g149(.dina(n221),.dinb(w_Gid15_0[0]),.dout(God15),.clk(gclk));
	jand g150(.dina(w_n149_0[2]),.dinb(w_n135_0[0]),.dout(n223),.clk(gclk));
	jand g151(.dina(w_n156_0[0]),.dinb(w_n85_0[2]),.dout(n224),.clk(gclk));
	jxor g152(.dina(w_n112_2[0]),.dinb(w_n187_2[0]),.dout(n225),.clk(gclk));
	jand g153(.dina(n225),.dinb(w_n174_0[0]),.dout(n226),.clk(gclk));
	jand g154(.dina(n226),.dinb(w_n200_0[0]),.dout(n227),.clk(gclk));
	jxor g155(.dina(w_n202_2[0]),.dinb(w_n166_2[0]),.dout(n228),.clk(gclk));
	jand g156(.dina(n228),.dinb(w_n99_0[0]),.dout(n229),.clk(gclk));
	jand g157(.dina(n229),.dinb(w_n188_0[0]),.dout(n230),.clk(gclk));
	jcb g158(.dina(n230),.dinb(n227),.dout(n231));
	jand g159(.dina(w_n231_0[1]),.dinb(w_dff_B_hxqAOgCD5_1),.dout(n232),.clk(gclk));
	jand g160(.dina(w_n232_0[1]),.dinb(w_n223_0[1]),.dout(n233),.clk(gclk));
	jand g161(.dina(w_n233_1[1]),.dinb(w_n166_1[2]),.dout(n234),.clk(gclk));
	jxor g162(.dina(n234),.dinb(w_Gid16_0[0]),.dout(God16),.clk(gclk));
	jand g163(.dina(w_n233_1[0]),.dinb(w_n202_1[2]),.dout(n236),.clk(gclk));
	jxor g164(.dina(n236),.dinb(w_Gid17_0[0]),.dout(God17),.clk(gclk));
	jand g165(.dina(w_n233_0[2]),.dinb(w_n112_1[2]),.dout(n238),.clk(gclk));
	jxor g166(.dina(n238),.dinb(w_Gid18_0[0]),.dout(God18),.clk(gclk));
	jand g167(.dina(w_n233_0[1]),.dinb(w_n187_1[2]),.dout(n240),.clk(gclk));
	jxor g168(.dina(n240),.dinb(w_Gid19_0[0]),.dout(God19),.clk(gclk));
	jand g169(.dina(w_n143_0[0]),.dinb(w_n147_0[2]),.dout(n242),.clk(gclk));
	jand g170(.dina(w_n232_0[0]),.dinb(w_n242_0[1]),.dout(n243),.clk(gclk));
	jand g171(.dina(w_n243_1[1]),.dinb(w_n166_1[1]),.dout(n244),.clk(gclk));
	jxor g172(.dina(n244),.dinb(w_Gid20_0[0]),.dout(God20),.clk(gclk));
	jand g173(.dina(w_n243_1[0]),.dinb(w_n202_1[1]),.dout(n246),.clk(gclk));
	jxor g174(.dina(n246),.dinb(w_Gid21_0[0]),.dout(God21),.clk(gclk));
	jand g175(.dina(w_n243_0[2]),.dinb(w_n112_1[1]),.dout(n248),.clk(gclk));
	jxor g176(.dina(n248),.dinb(w_Gid22_0[0]),.dout(God22),.clk(gclk));
	jand g177(.dina(w_n243_0[1]),.dinb(w_n187_1[1]),.dout(n250),.clk(gclk));
	jxor g178(.dina(n250),.dinb(w_Gid23_0[0]),.dout(God23),.clk(gclk));
	jand g179(.dina(w_n126_0[2]),.dinb(w_n153_0[0]),.dout(n252),.clk(gclk));
	jand g180(.dina(w_n231_0[0]),.dinb(w_dff_B_HOwqrcPC7_1),.dout(n253),.clk(gclk));
	jand g181(.dina(w_n253_0[1]),.dinb(w_n223_0[0]),.dout(n254),.clk(gclk));
	jand g182(.dina(w_n254_1[1]),.dinb(w_n166_1[0]),.dout(n255),.clk(gclk));
	jxor g183(.dina(n255),.dinb(w_Gid24_0[0]),.dout(God24),.clk(gclk));
	jand g184(.dina(w_n254_1[0]),.dinb(w_n202_1[0]),.dout(n257),.clk(gclk));
	jxor g185(.dina(n257),.dinb(w_Gid25_0[0]),.dout(God25),.clk(gclk));
	jand g186(.dina(w_n254_0[2]),.dinb(w_n112_1[0]),.dout(n259),.clk(gclk));
	jxor g187(.dina(n259),.dinb(w_Gid26_0[0]),.dout(God26),.clk(gclk));
	jand g188(.dina(w_n254_0[1]),.dinb(w_n187_1[0]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_Gid27_0[0]),.dout(God27),.clk(gclk));
	jand g190(.dina(w_n253_0[0]),.dinb(w_n242_0[0]),.dout(n263),.clk(gclk));
	jand g191(.dina(w_n263_1[1]),.dinb(w_n166_0[2]),.dout(n264),.clk(gclk));
	jxor g192(.dina(n264),.dinb(w_Gid28_0[0]),.dout(God28),.clk(gclk));
	jand g193(.dina(w_n263_1[0]),.dinb(w_n202_0[2]),.dout(n266),.clk(gclk));
	jxor g194(.dina(n266),.dinb(w_Gid29_0[0]),.dout(God29),.clk(gclk));
	jand g195(.dina(w_n263_0[2]),.dinb(w_n112_0[2]),.dout(n268),.clk(gclk));
	jxor g196(.dina(n268),.dinb(w_Gid30_0[0]),.dout(God30),.clk(gclk));
	jand g197(.dina(w_n263_0[1]),.dinb(w_n187_0[2]),.dout(n270),.clk(gclk));
	jxor g198(.dina(n270),.dinb(w_Gid31_0[0]),.dout(God31),.clk(gclk));
	jspl3 jspl3_w_Gid0_0(.douta(w_dff_A_PJThdGI04_0),.doutb(w_Gid0_0[1]),.doutc(w_Gid0_0[2]),.din(Gid0));
	jspl3 jspl3_w_Gid1_0(.douta(w_dff_A_p0jsRYB00_0),.doutb(w_Gid1_0[1]),.doutc(w_Gid1_0[2]),.din(Gid1));
	jspl3 jspl3_w_Gid2_0(.douta(w_dff_A_FK4WOMqW0_0),.doutb(w_Gid2_0[1]),.doutc(w_Gid2_0[2]),.din(Gid2));
	jspl3 jspl3_w_Gid3_0(.douta(w_dff_A_fXFBxHfN8_0),.doutb(w_Gid3_0[1]),.doutc(w_Gid3_0[2]),.din(Gid3));
	jspl3 jspl3_w_Gid4_0(.douta(w_dff_A_6WBKOtYd4_0),.doutb(w_Gid4_0[1]),.doutc(w_Gid4_0[2]),.din(Gid4));
	jspl3 jspl3_w_Gid5_0(.douta(w_dff_A_pKEIzH8h8_0),.doutb(w_Gid5_0[1]),.doutc(w_Gid5_0[2]),.din(Gid5));
	jspl3 jspl3_w_Gid6_0(.douta(w_dff_A_OxTmT3AS5_0),.doutb(w_Gid6_0[1]),.doutc(w_Gid6_0[2]),.din(Gid6));
	jspl3 jspl3_w_Gid7_0(.douta(w_dff_A_wW1QB6Ip8_0),.doutb(w_Gid7_0[1]),.doutc(w_Gid7_0[2]),.din(Gid7));
	jspl3 jspl3_w_Gid8_0(.douta(w_dff_A_7GamyOpk3_0),.doutb(w_Gid8_0[1]),.doutc(w_Gid8_0[2]),.din(Gid8));
	jspl3 jspl3_w_Gid9_0(.douta(w_dff_A_kYblhX612_0),.doutb(w_Gid9_0[1]),.doutc(w_Gid9_0[2]),.din(Gid9));
	jspl3 jspl3_w_Gid10_0(.douta(w_dff_A_Ht497OWo8_0),.doutb(w_Gid10_0[1]),.doutc(w_Gid10_0[2]),.din(Gid10));
	jspl3 jspl3_w_Gid11_0(.douta(w_dff_A_9ho4Nn9t4_0),.doutb(w_Gid11_0[1]),.doutc(w_Gid11_0[2]),.din(Gid11));
	jspl3 jspl3_w_Gid12_0(.douta(w_dff_A_93gcXRbU9_0),.doutb(w_Gid12_0[1]),.doutc(w_Gid12_0[2]),.din(Gid12));
	jspl3 jspl3_w_Gid13_0(.douta(w_dff_A_zvgLAkvb8_0),.doutb(w_Gid13_0[1]),.doutc(w_Gid13_0[2]),.din(Gid13));
	jspl3 jspl3_w_Gid14_0(.douta(w_dff_A_nsfUXMgG0_0),.doutb(w_Gid14_0[1]),.doutc(w_Gid14_0[2]),.din(Gid14));
	jspl3 jspl3_w_Gid15_0(.douta(w_dff_A_W47mm7Ai1_0),.doutb(w_Gid15_0[1]),.doutc(w_Gid15_0[2]),.din(Gid15));
	jspl3 jspl3_w_Gid16_0(.douta(w_dff_A_xcMew2LF5_0),.doutb(w_Gid16_0[1]),.doutc(w_Gid16_0[2]),.din(Gid16));
	jspl3 jspl3_w_Gid17_0(.douta(w_dff_A_cxzokb8r0_0),.doutb(w_Gid17_0[1]),.doutc(w_Gid17_0[2]),.din(Gid17));
	jspl3 jspl3_w_Gid18_0(.douta(w_dff_A_4jr6RA0o0_0),.doutb(w_Gid18_0[1]),.doutc(w_Gid18_0[2]),.din(Gid18));
	jspl3 jspl3_w_Gid19_0(.douta(w_dff_A_l7GTsDaa6_0),.doutb(w_Gid19_0[1]),.doutc(w_Gid19_0[2]),.din(Gid19));
	jspl3 jspl3_w_Gid20_0(.douta(w_dff_A_aElP0Gp81_0),.doutb(w_Gid20_0[1]),.doutc(w_Gid20_0[2]),.din(Gid20));
	jspl3 jspl3_w_Gid21_0(.douta(w_dff_A_hoRlUHJb5_0),.doutb(w_Gid21_0[1]),.doutc(w_Gid21_0[2]),.din(Gid21));
	jspl3 jspl3_w_Gid22_0(.douta(w_dff_A_O6iHzNyD7_0),.doutb(w_Gid22_0[1]),.doutc(w_Gid22_0[2]),.din(Gid22));
	jspl3 jspl3_w_Gid23_0(.douta(w_dff_A_13P3eB4r7_0),.doutb(w_Gid23_0[1]),.doutc(w_Gid23_0[2]),.din(Gid23));
	jspl3 jspl3_w_Gid24_0(.douta(w_dff_A_OQpiXoZq8_0),.doutb(w_Gid24_0[1]),.doutc(w_Gid24_0[2]),.din(Gid24));
	jspl3 jspl3_w_Gid25_0(.douta(w_dff_A_lr4aCgXD3_0),.doutb(w_Gid25_0[1]),.doutc(w_Gid25_0[2]),.din(Gid25));
	jspl3 jspl3_w_Gid26_0(.douta(w_dff_A_uuZuWW9G7_0),.doutb(w_Gid26_0[1]),.doutc(w_Gid26_0[2]),.din(Gid26));
	jspl3 jspl3_w_Gid27_0(.douta(w_dff_A_Bw250faj5_0),.doutb(w_Gid27_0[1]),.doutc(w_Gid27_0[2]),.din(Gid27));
	jspl3 jspl3_w_Gid28_0(.douta(w_dff_A_D5KmenKw5_0),.doutb(w_Gid28_0[1]),.doutc(w_Gid28_0[2]),.din(Gid28));
	jspl3 jspl3_w_Gid29_0(.douta(w_dff_A_GkSNTNLK1_0),.doutb(w_Gid29_0[1]),.doutc(w_Gid29_0[2]),.din(Gid29));
	jspl3 jspl3_w_Gid30_0(.douta(w_dff_A_QfoNNBsi3_0),.doutb(w_Gid30_0[1]),.doutc(w_Gid30_0[2]),.din(Gid30));
	jspl3 jspl3_w_Gid31_0(.douta(w_dff_A_PDVxLHao2_0),.doutb(w_Gid31_0[1]),.doutc(w_Gid31_0[2]),.din(Gid31));
	jspl3 jspl3_w_Gr_0(.douta(w_Gr_0[0]),.doutb(w_Gr_0[1]),.doutc(w_Gr_0[2]),.din(Gr));
	jspl3 jspl3_w_Gr_1(.douta(w_Gr_1[0]),.doutb(w_Gr_1[1]),.doutc(w_Gr_1[2]),.din(w_Gr_0[0]));
	jspl3 jspl3_w_Gr_2(.douta(w_Gr_2[0]),.doutb(w_Gr_2[1]),.doutc(w_Gr_2[2]),.din(w_Gr_0[1]));
	jspl jspl_w_Gr_3(.douta(w_Gr_3[0]),.doutb(w_Gr_3[1]),.din(w_Gr_0[2]));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_dff_A_rDiJ44VL5_1),.din(n76));
	jspl jspl_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.din(n80));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_NhYTO4iR6_0),.doutb(w_n85_0[1]),.doutc(w_n85_0[2]),.din(n85));
	jspl3 jspl3_w_n85_1(.douta(w_n85_1[0]),.doutb(w_n85_1[1]),.doutc(w_n85_1[2]),.din(w_n85_0[0]));
	jspl jspl_w_n85_2(.douta(w_dff_A_e8wbs50M9_0),.doutb(w_n85_2[1]),.din(w_n85_0[1]));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n89_0(.douta(w_dff_A_IE9x3CTg7_0),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.din(n94));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n99_0(.douta(w_dff_A_w5AEq2sN0_0),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.din(n110));
	jspl3 jspl3_w_n112_0(.douta(w_dff_A_n7uOfbzP8_0),.doutb(w_n112_0[1]),.doutc(w_dff_A_0YxebjIB7_2),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_dff_A_fHdPikeT7_1),.din(w_dff_B_KtSH61WO6_2));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.din(n116));
	jspl jspl_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_EYsURZ2f7_1),.din(n117));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n124_0(.douta(w_n124_0[0]),.doutb(w_n124_0[1]),.doutc(w_n124_0[2]),.din(n124));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl3 jspl3_w_n126_0(.douta(w_dff_A_xLUXIChb1_0),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl3 jspl3_w_n126_1(.douta(w_n126_1[0]),.doutb(w_n126_1[1]),.doutc(w_n126_1[2]),.din(w_n126_0[0]));
	jspl jspl_w_n126_2(.douta(w_dff_A_xyTxYRt59_0),.doutb(w_n126_2[1]),.din(w_n126_0[1]));
	jspl jspl_w_n128_0(.douta(w_dff_A_6ozCoOJb2_0),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n134_0(.douta(w_n134_0[0]),.doutb(w_n134_0[1]),.din(n134));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.din(n135));
	jspl jspl_w_n136_0(.douta(w_dff_A_xLN5Qrlm2_0),.doutb(w_n136_0[1]),.din(n136));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl3 jspl3_w_n147_0(.douta(w_dff_A_Lke3J96z3_0),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl3 jspl3_w_n147_1(.douta(w_n147_1[0]),.doutb(w_n147_1[1]),.doutc(w_n147_1[2]),.din(w_n147_0[0]));
	jspl jspl_w_n147_2(.douta(w_dff_A_kFFQf1lp7_0),.doutb(w_n147_2[1]),.din(w_n147_0[1]));
	jspl3 jspl3_w_n149_0(.douta(w_dff_A_xrf3zG4d0_0),.doutb(w_n149_0[1]),.doutc(w_n149_0[2]),.din(n149));
	jspl3 jspl3_w_n149_1(.douta(w_n149_1[0]),.doutb(w_n149_1[1]),.doutc(w_n149_1[2]),.din(w_n149_0[0]));
	jspl jspl_w_n149_2(.douta(w_dff_A_7V5asUu05_0),.doutb(w_n149_2[1]),.din(w_n149_0[1]));
	jspl jspl_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.din(n153));
	jspl jspl_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.din(n156));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl3 jspl3_w_n166_0(.douta(w_dff_A_E95DKjEp2_0),.doutb(w_n166_0[1]),.doutc(w_dff_A_m2bEKbcd8_2),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.doutc(w_n166_1[2]),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_n166_2[2]),.din(w_n166_0[1]));
	jspl jspl_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_dff_A_VjxPrIe00_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.din(n173));
	jspl jspl_w_n174_0(.douta(w_dff_A_UnyKoXRX1_0),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_dff_A_xsHvLrT50_0),.doutb(w_n175_0[1]),.din(w_dff_B_A3cqmxTP5_2));
	jspl3 jspl3_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.doutc(w_n177_0[2]),.din(n177));
	jspl jspl_w_n177_1(.douta(w_n177_1[0]),.doutb(w_n177_1[1]),.din(w_n177_0[0]));
	jspl3 jspl3_w_n187_0(.douta(w_dff_A_HsFZPwNr8_0),.doutb(w_n187_0[1]),.doutc(w_dff_A_Fmw23bkx7_2),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_n187_1[0]),.doutb(w_n187_1[1]),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n187_2(.douta(w_n187_2[0]),.doutb(w_dff_A_RBghgPVD6_1),.din(w_n187_0[1]));
	jspl jspl_w_n188_0(.douta(w_dff_A_AcHISKVu4_0),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.din(n190));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n191_1(.douta(w_n191_1[0]),.doutb(w_n191_1[1]),.din(w_n191_0[0]));
	jspl jspl_w_n200_0(.douta(w_dff_A_m72EqgDs9_0),.doutb(w_n200_0[1]),.din(n200));
	jspl3 jspl3_w_n202_0(.douta(w_dff_A_IvdKllUA9_0),.doutb(w_n202_0[1]),.doutc(w_dff_A_I4pFocEd7_2),.din(n202));
	jspl3 jspl3_w_n202_1(.douta(w_n202_1[0]),.doutb(w_n202_1[1]),.doutc(w_n202_1[2]),.din(w_n202_0[0]));
	jspl jspl_w_n202_2(.douta(w_n202_2[0]),.doutb(w_dff_A_g0O7vAGz7_1),.din(w_n202_0[1]));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(w_dff_B_yyxcoOdw6_2));
	jspl3 jspl3_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.doutc(w_n205_0[2]),.din(n205));
	jspl jspl_w_n205_1(.douta(w_n205_1[0]),.doutb(w_n205_1[1]),.din(w_n205_0[0]));
	jspl3 jspl3_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.doutc(w_n214_0[2]),.din(n214));
	jspl jspl_w_n214_1(.douta(w_n214_1[0]),.doutb(w_n214_1[1]),.din(w_n214_0[0]));
	jspl jspl_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.din(w_dff_B_gpYsGkyH9_2));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.din(n231));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl jspl_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.din(w_n233_0[0]));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(w_dff_B_b6iKLfib8_2));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n243_1(.douta(w_n243_1[0]),.doutb(w_n243_1[1]),.din(w_n243_0[0]));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.din(n253));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl jspl_w_n254_1(.douta(w_n254_1[0]),.doutb(w_n254_1[1]),.din(w_n254_0[0]));
	jspl3 jspl3_w_n263_0(.douta(w_n263_0[0]),.doutb(w_n263_0[1]),.doutc(w_n263_0[2]),.din(n263));
	jspl jspl_w_n263_1(.douta(w_n263_1[0]),.doutb(w_n263_1[1]),.din(w_n263_0[0]));
	jdff dff_A_xsHvLrT50_0(.dout(w_n175_0[0]),.din(w_dff_A_xsHvLrT50_0),.clk(gclk));
	jdff dff_B_A3cqmxTP5_2(.din(n175),.dout(w_dff_B_A3cqmxTP5_2),.clk(gclk));
	jdff dff_A_fHdPikeT7_1(.dout(w_n113_0[1]),.din(w_dff_A_fHdPikeT7_1),.clk(gclk));
	jdff dff_B_KtSH61WO6_2(.din(n113),.dout(w_dff_B_KtSH61WO6_2),.clk(gclk));
	jdff dff_B_yyxcoOdw6_2(.din(n203),.dout(w_dff_B_yyxcoOdw6_2),.clk(gclk));
	jdff dff_A_CKBUldlp2_0(.dout(w_n149_2[0]),.din(w_dff_A_CKBUldlp2_0),.clk(gclk));
	jdff dff_A_7SxSECa31_0(.dout(w_dff_A_CKBUldlp2_0),.din(w_dff_A_7SxSECa31_0),.clk(gclk));
	jdff dff_A_zSMxf2Hg5_0(.dout(w_dff_A_7SxSECa31_0),.din(w_dff_A_zSMxf2Hg5_0),.clk(gclk));
	jdff dff_A_7V5asUu05_0(.dout(w_dff_A_zSMxf2Hg5_0),.din(w_dff_A_7V5asUu05_0),.clk(gclk));
	jdff dff_A_tGSrHpHG2_0(.dout(w_n147_2[0]),.din(w_dff_A_tGSrHpHG2_0),.clk(gclk));
	jdff dff_A_JNWAGWUt8_0(.dout(w_dff_A_tGSrHpHG2_0),.din(w_dff_A_JNWAGWUt8_0),.clk(gclk));
	jdff dff_A_9gAaidIj4_0(.dout(w_dff_A_JNWAGWUt8_0),.din(w_dff_A_9gAaidIj4_0),.clk(gclk));
	jdff dff_A_kFFQf1lp7_0(.dout(w_dff_A_9gAaidIj4_0),.din(w_dff_A_kFFQf1lp7_0),.clk(gclk));
	jdff dff_A_Uf1PxO8J5_0(.dout(w_n126_2[0]),.din(w_dff_A_Uf1PxO8J5_0),.clk(gclk));
	jdff dff_A_sxZdp59U5_0(.dout(w_dff_A_Uf1PxO8J5_0),.din(w_dff_A_sxZdp59U5_0),.clk(gclk));
	jdff dff_A_m2mR11So6_0(.dout(w_dff_A_sxZdp59U5_0),.din(w_dff_A_m2mR11So6_0),.clk(gclk));
	jdff dff_A_xyTxYRt59_0(.dout(w_dff_A_m2mR11So6_0),.din(w_dff_A_xyTxYRt59_0),.clk(gclk));
	jdff dff_A_V8stKZ9U4_0(.dout(w_n85_2[0]),.din(w_dff_A_V8stKZ9U4_0),.clk(gclk));
	jdff dff_A_G9M1Bjrt0_0(.dout(w_dff_A_V8stKZ9U4_0),.din(w_dff_A_G9M1Bjrt0_0),.clk(gclk));
	jdff dff_A_6MSWn3oX6_0(.dout(w_dff_A_G9M1Bjrt0_0),.din(w_dff_A_6MSWn3oX6_0),.clk(gclk));
	jdff dff_A_e8wbs50M9_0(.dout(w_dff_A_6MSWn3oX6_0),.din(w_dff_A_e8wbs50M9_0),.clk(gclk));
	jdff dff_B_b5epyP8x6_1(.din(n224),.dout(w_dff_B_b5epyP8x6_1),.clk(gclk));
	jdff dff_B_hxqAOgCD5_1(.din(w_dff_B_b5epyP8x6_1),.dout(w_dff_B_hxqAOgCD5_1),.clk(gclk));
	jdff dff_A_4IPXSKR66_0(.dout(w_n85_0[0]),.din(w_dff_A_4IPXSKR66_0),.clk(gclk));
	jdff dff_A_8MGPt5s03_0(.dout(w_dff_A_4IPXSKR66_0),.din(w_dff_A_8MGPt5s03_0),.clk(gclk));
	jdff dff_A_GjnX3kKg4_0(.dout(w_dff_A_8MGPt5s03_0),.din(w_dff_A_GjnX3kKg4_0),.clk(gclk));
	jdff dff_A_NhYTO4iR6_0(.dout(w_dff_A_GjnX3kKg4_0),.din(w_dff_A_NhYTO4iR6_0),.clk(gclk));
	jdff dff_B_Rdj7wqLX1_2(.din(n223),.dout(w_dff_B_Rdj7wqLX1_2),.clk(gclk));
	jdff dff_B_HItKXbww1_2(.din(w_dff_B_Rdj7wqLX1_2),.dout(w_dff_B_HItKXbww1_2),.clk(gclk));
	jdff dff_B_gpYsGkyH9_2(.din(w_dff_B_HItKXbww1_2),.dout(w_dff_B_gpYsGkyH9_2),.clk(gclk));
	jdff dff_A_4a4Bc84i9_0(.dout(w_n149_0[0]),.din(w_dff_A_4a4Bc84i9_0),.clk(gclk));
	jdff dff_A_CZswUChP3_0(.dout(w_dff_A_4a4Bc84i9_0),.din(w_dff_A_CZswUChP3_0),.clk(gclk));
	jdff dff_A_LvEISj5n0_0(.dout(w_dff_A_CZswUChP3_0),.din(w_dff_A_LvEISj5n0_0),.clk(gclk));
	jdff dff_A_xrf3zG4d0_0(.dout(w_dff_A_LvEISj5n0_0),.din(w_dff_A_xrf3zG4d0_0),.clk(gclk));
	jdff dff_B_ODVDWLU88_1(.din(n252),.dout(w_dff_B_ODVDWLU88_1),.clk(gclk));
	jdff dff_B_HOwqrcPC7_1(.din(w_dff_B_ODVDWLU88_1),.dout(w_dff_B_HOwqrcPC7_1),.clk(gclk));
	jdff dff_A_g0O7vAGz7_1(.dout(w_n202_2[1]),.din(w_dff_A_g0O7vAGz7_1),.clk(gclk));
	jdff dff_A_Uas4QUmJ3_0(.dout(w_n202_0[0]),.din(w_dff_A_Uas4QUmJ3_0),.clk(gclk));
	jdff dff_A_AlCXvMgW0_0(.dout(w_dff_A_Uas4QUmJ3_0),.din(w_dff_A_AlCXvMgW0_0),.clk(gclk));
	jdff dff_A_QeTBLKvK4_0(.dout(w_dff_A_AlCXvMgW0_0),.din(w_dff_A_QeTBLKvK4_0),.clk(gclk));
	jdff dff_A_W1E1wB682_0(.dout(w_dff_A_QeTBLKvK4_0),.din(w_dff_A_W1E1wB682_0),.clk(gclk));
	jdff dff_A_IvdKllUA9_0(.dout(w_dff_A_W1E1wB682_0),.din(w_dff_A_IvdKllUA9_0),.clk(gclk));
	jdff dff_A_au9cLAnc1_2(.dout(w_n202_0[2]),.din(w_dff_A_au9cLAnc1_2),.clk(gclk));
	jdff dff_A_iYnrnaLZ9_2(.dout(w_dff_A_au9cLAnc1_2),.din(w_dff_A_iYnrnaLZ9_2),.clk(gclk));
	jdff dff_A_c8PAKLHG2_2(.dout(w_dff_A_iYnrnaLZ9_2),.din(w_dff_A_c8PAKLHG2_2),.clk(gclk));
	jdff dff_A_2fp89xUw1_2(.dout(w_dff_A_c8PAKLHG2_2),.din(w_dff_A_2fp89xUw1_2),.clk(gclk));
	jdff dff_A_I4pFocEd7_2(.dout(w_dff_A_2fp89xUw1_2),.din(w_dff_A_I4pFocEd7_2),.clk(gclk));
	jdff dff_A_w5AEq2sN0_0(.dout(w_n99_0[0]),.din(w_dff_A_w5AEq2sN0_0),.clk(gclk));
	jdff dff_A_AcHISKVu4_0(.dout(w_n188_0[0]),.din(w_dff_A_AcHISKVu4_0),.clk(gclk));
	jdff dff_A_QY6P5fuv9_0(.dout(w_n112_0[0]),.din(w_dff_A_QY6P5fuv9_0),.clk(gclk));
	jdff dff_A_MPzX67hC7_0(.dout(w_dff_A_QY6P5fuv9_0),.din(w_dff_A_MPzX67hC7_0),.clk(gclk));
	jdff dff_A_VpyKfITQ2_0(.dout(w_dff_A_MPzX67hC7_0),.din(w_dff_A_VpyKfITQ2_0),.clk(gclk));
	jdff dff_A_AY1ApXn43_0(.dout(w_dff_A_VpyKfITQ2_0),.din(w_dff_A_AY1ApXn43_0),.clk(gclk));
	jdff dff_A_n7uOfbzP8_0(.dout(w_dff_A_AY1ApXn43_0),.din(w_dff_A_n7uOfbzP8_0),.clk(gclk));
	jdff dff_A_irTlR0jg6_2(.dout(w_n112_0[2]),.din(w_dff_A_irTlR0jg6_2),.clk(gclk));
	jdff dff_A_ZshkRoN08_2(.dout(w_dff_A_irTlR0jg6_2),.din(w_dff_A_ZshkRoN08_2),.clk(gclk));
	jdff dff_A_p3hUBF6k6_2(.dout(w_dff_A_ZshkRoN08_2),.din(w_dff_A_p3hUBF6k6_2),.clk(gclk));
	jdff dff_A_Rvo4aQ0m1_2(.dout(w_dff_A_p3hUBF6k6_2),.din(w_dff_A_Rvo4aQ0m1_2),.clk(gclk));
	jdff dff_A_0YxebjIB7_2(.dout(w_dff_A_Rvo4aQ0m1_2),.din(w_dff_A_0YxebjIB7_2),.clk(gclk));
	jdff dff_B_b67s7T1b4_0(.din(n103),.dout(w_dff_B_b67s7T1b4_0),.clk(gclk));
	jdff dff_A_RBghgPVD6_1(.dout(w_n187_2[1]),.din(w_dff_A_RBghgPVD6_1),.clk(gclk));
	jdff dff_A_kuX0xbhN0_0(.dout(w_n187_0[0]),.din(w_dff_A_kuX0xbhN0_0),.clk(gclk));
	jdff dff_A_n1bXLGu77_0(.dout(w_dff_A_kuX0xbhN0_0),.din(w_dff_A_n1bXLGu77_0),.clk(gclk));
	jdff dff_A_gFHqnZST6_0(.dout(w_dff_A_n1bXLGu77_0),.din(w_dff_A_gFHqnZST6_0),.clk(gclk));
	jdff dff_A_lTTVHCoY6_0(.dout(w_dff_A_gFHqnZST6_0),.din(w_dff_A_lTTVHCoY6_0),.clk(gclk));
	jdff dff_A_HsFZPwNr8_0(.dout(w_dff_A_lTTVHCoY6_0),.din(w_dff_A_HsFZPwNr8_0),.clk(gclk));
	jdff dff_A_l09FAviz5_2(.dout(w_n187_0[2]),.din(w_dff_A_l09FAviz5_2),.clk(gclk));
	jdff dff_A_vbRSpGdV3_2(.dout(w_dff_A_l09FAviz5_2),.din(w_dff_A_vbRSpGdV3_2),.clk(gclk));
	jdff dff_A_NioLwYLQ4_2(.dout(w_dff_A_vbRSpGdV3_2),.din(w_dff_A_NioLwYLQ4_2),.clk(gclk));
	jdff dff_A_558Tsuj70_2(.dout(w_dff_A_NioLwYLQ4_2),.din(w_dff_A_558Tsuj70_2),.clk(gclk));
	jdff dff_A_Fmw23bkx7_2(.dout(w_dff_A_558Tsuj70_2),.din(w_dff_A_Fmw23bkx7_2),.clk(gclk));
	jdff dff_A_IE9x3CTg7_0(.dout(w_n89_0[0]),.din(w_dff_A_IE9x3CTg7_0),.clk(gclk));
	jdff dff_A_UnyKoXRX1_0(.dout(w_n174_0[0]),.din(w_dff_A_UnyKoXRX1_0),.clk(gclk));
	jdff dff_A_VjxPrIe00_0(.dout(w_n170_0[0]),.din(w_dff_A_VjxPrIe00_0),.clk(gclk));
	jdff dff_A_m72EqgDs9_0(.dout(w_n200_0[0]),.din(w_dff_A_m72EqgDs9_0),.clk(gclk));
	jdff dff_A_1ZpFomE41_0(.dout(w_n166_0[0]),.din(w_dff_A_1ZpFomE41_0),.clk(gclk));
	jdff dff_A_gale4REy2_0(.dout(w_dff_A_1ZpFomE41_0),.din(w_dff_A_gale4REy2_0),.clk(gclk));
	jdff dff_A_1o9TibeK8_0(.dout(w_dff_A_gale4REy2_0),.din(w_dff_A_1o9TibeK8_0),.clk(gclk));
	jdff dff_A_tqXyFDpb1_0(.dout(w_dff_A_1o9TibeK8_0),.din(w_dff_A_tqXyFDpb1_0),.clk(gclk));
	jdff dff_A_E95DKjEp2_0(.dout(w_dff_A_tqXyFDpb1_0),.din(w_dff_A_E95DKjEp2_0),.clk(gclk));
	jdff dff_A_STeSXPb63_2(.dout(w_n166_0[2]),.din(w_dff_A_STeSXPb63_2),.clk(gclk));
	jdff dff_A_JHBPrTm53_2(.dout(w_dff_A_STeSXPb63_2),.din(w_dff_A_JHBPrTm53_2),.clk(gclk));
	jdff dff_A_NAlJo5TF6_2(.dout(w_dff_A_JHBPrTm53_2),.din(w_dff_A_NAlJo5TF6_2),.clk(gclk));
	jdff dff_A_ClEVmivN9_2(.dout(w_dff_A_NAlJo5TF6_2),.din(w_dff_A_ClEVmivN9_2),.clk(gclk));
	jdff dff_A_m2bEKbcd8_2(.dout(w_dff_A_ClEVmivN9_2),.din(w_dff_A_m2bEKbcd8_2),.clk(gclk));
	jdff dff_B_5CFbhW9H9_0(.din(n163),.dout(w_dff_B_5CFbhW9H9_0),.clk(gclk));
	jdff dff_A_mBSGuVS72_0(.dout(w_n126_0[0]),.din(w_dff_A_mBSGuVS72_0),.clk(gclk));
	jdff dff_A_QdEEbRal4_0(.dout(w_dff_A_mBSGuVS72_0),.din(w_dff_A_QdEEbRal4_0),.clk(gclk));
	jdff dff_A_NLenSW1i8_0(.dout(w_dff_A_QdEEbRal4_0),.din(w_dff_A_NLenSW1i8_0),.clk(gclk));
	jdff dff_A_xLUXIChb1_0(.dout(w_dff_A_NLenSW1i8_0),.din(w_dff_A_xLUXIChb1_0),.clk(gclk));
	jdff dff_A_EYsURZ2f7_1(.dout(w_n117_0[1]),.din(w_dff_A_EYsURZ2f7_1),.clk(gclk));
	jdff dff_A_JqDoPysW3_0(.dout(w_Gid5_0[0]),.din(w_dff_A_JqDoPysW3_0),.clk(gclk));
	jdff dff_A_Osgv8huM7_0(.dout(w_dff_A_JqDoPysW3_0),.din(w_dff_A_Osgv8huM7_0),.clk(gclk));
	jdff dff_A_EOr20ERz1_0(.dout(w_dff_A_Osgv8huM7_0),.din(w_dff_A_EOr20ERz1_0),.clk(gclk));
	jdff dff_A_k6MyJVur1_0(.dout(w_dff_A_EOr20ERz1_0),.din(w_dff_A_k6MyJVur1_0),.clk(gclk));
	jdff dff_A_qKHHdcJL0_0(.dout(w_dff_A_k6MyJVur1_0),.din(w_dff_A_qKHHdcJL0_0),.clk(gclk));
	jdff dff_A_IFo2YrqA7_0(.dout(w_dff_A_qKHHdcJL0_0),.din(w_dff_A_IFo2YrqA7_0),.clk(gclk));
	jdff dff_A_paypljLX4_0(.dout(w_dff_A_IFo2YrqA7_0),.din(w_dff_A_paypljLX4_0),.clk(gclk));
	jdff dff_A_X3DKZrh94_0(.dout(w_dff_A_paypljLX4_0),.din(w_dff_A_X3DKZrh94_0),.clk(gclk));
	jdff dff_A_pKEIzH8h8_0(.dout(w_dff_A_X3DKZrh94_0),.din(w_dff_A_pKEIzH8h8_0),.clk(gclk));
	jdff dff_A_NQ7akYmb7_0(.dout(w_Gid1_0[0]),.din(w_dff_A_NQ7akYmb7_0),.clk(gclk));
	jdff dff_A_yGMkx7uv1_0(.dout(w_dff_A_NQ7akYmb7_0),.din(w_dff_A_yGMkx7uv1_0),.clk(gclk));
	jdff dff_A_mmF43fjx4_0(.dout(w_dff_A_yGMkx7uv1_0),.din(w_dff_A_mmF43fjx4_0),.clk(gclk));
	jdff dff_A_wKmK6h7u6_0(.dout(w_dff_A_mmF43fjx4_0),.din(w_dff_A_wKmK6h7u6_0),.clk(gclk));
	jdff dff_A_4iHz0Oci6_0(.dout(w_dff_A_wKmK6h7u6_0),.din(w_dff_A_4iHz0Oci6_0),.clk(gclk));
	jdff dff_A_Cb4wNhcz0_0(.dout(w_dff_A_4iHz0Oci6_0),.din(w_dff_A_Cb4wNhcz0_0),.clk(gclk));
	jdff dff_A_45CuhMzY4_0(.dout(w_dff_A_Cb4wNhcz0_0),.din(w_dff_A_45CuhMzY4_0),.clk(gclk));
	jdff dff_A_A0IBrAuK6_0(.dout(w_dff_A_45CuhMzY4_0),.din(w_dff_A_A0IBrAuK6_0),.clk(gclk));
	jdff dff_A_p0jsRYB00_0(.dout(w_dff_A_A0IBrAuK6_0),.din(w_dff_A_p0jsRYB00_0),.clk(gclk));
	jdff dff_A_MNhKk2F74_0(.dout(w_Gid13_0[0]),.din(w_dff_A_MNhKk2F74_0),.clk(gclk));
	jdff dff_A_7BOnHrtx5_0(.dout(w_dff_A_MNhKk2F74_0),.din(w_dff_A_7BOnHrtx5_0),.clk(gclk));
	jdff dff_A_JGqyI7v55_0(.dout(w_dff_A_7BOnHrtx5_0),.din(w_dff_A_JGqyI7v55_0),.clk(gclk));
	jdff dff_A_vsUBeMsF1_0(.dout(w_dff_A_JGqyI7v55_0),.din(w_dff_A_vsUBeMsF1_0),.clk(gclk));
	jdff dff_A_QuA8xfCI1_0(.dout(w_dff_A_vsUBeMsF1_0),.din(w_dff_A_QuA8xfCI1_0),.clk(gclk));
	jdff dff_A_7U3Kpizm6_0(.dout(w_dff_A_QuA8xfCI1_0),.din(w_dff_A_7U3Kpizm6_0),.clk(gclk));
	jdff dff_A_uupUxC8h7_0(.dout(w_dff_A_7U3Kpizm6_0),.din(w_dff_A_uupUxC8h7_0),.clk(gclk));
	jdff dff_A_qhHCfinI9_0(.dout(w_dff_A_uupUxC8h7_0),.din(w_dff_A_qhHCfinI9_0),.clk(gclk));
	jdff dff_A_zvgLAkvb8_0(.dout(w_dff_A_qhHCfinI9_0),.din(w_dff_A_zvgLAkvb8_0),.clk(gclk));
	jdff dff_A_iGdvqOos6_0(.dout(w_Gid9_0[0]),.din(w_dff_A_iGdvqOos6_0),.clk(gclk));
	jdff dff_A_WZREt1t41_0(.dout(w_dff_A_iGdvqOos6_0),.din(w_dff_A_WZREt1t41_0),.clk(gclk));
	jdff dff_A_12iKLGeb0_0(.dout(w_dff_A_WZREt1t41_0),.din(w_dff_A_12iKLGeb0_0),.clk(gclk));
	jdff dff_A_PIwCzpr43_0(.dout(w_dff_A_12iKLGeb0_0),.din(w_dff_A_PIwCzpr43_0),.clk(gclk));
	jdff dff_A_fS6FLVyQ9_0(.dout(w_dff_A_PIwCzpr43_0),.din(w_dff_A_fS6FLVyQ9_0),.clk(gclk));
	jdff dff_A_ckgMQ0re1_0(.dout(w_dff_A_fS6FLVyQ9_0),.din(w_dff_A_ckgMQ0re1_0),.clk(gclk));
	jdff dff_A_Ev5PtdyW4_0(.dout(w_dff_A_ckgMQ0re1_0),.din(w_dff_A_Ev5PtdyW4_0),.clk(gclk));
	jdff dff_A_bPLUxzyp2_0(.dout(w_dff_A_Ev5PtdyW4_0),.din(w_dff_A_bPLUxzyp2_0),.clk(gclk));
	jdff dff_A_kYblhX612_0(.dout(w_dff_A_bPLUxzyp2_0),.din(w_dff_A_kYblhX612_0),.clk(gclk));
	jdff dff_A_rDiJ44VL5_1(.dout(w_n76_0[1]),.din(w_dff_A_rDiJ44VL5_1),.clk(gclk));
	jdff dff_A_KfdWvmon5_0(.dout(w_Gid4_0[0]),.din(w_dff_A_KfdWvmon5_0),.clk(gclk));
	jdff dff_A_jynkVs1h9_0(.dout(w_dff_A_KfdWvmon5_0),.din(w_dff_A_jynkVs1h9_0),.clk(gclk));
	jdff dff_A_oMmIEPNC0_0(.dout(w_dff_A_jynkVs1h9_0),.din(w_dff_A_oMmIEPNC0_0),.clk(gclk));
	jdff dff_A_saxYz4xk3_0(.dout(w_dff_A_oMmIEPNC0_0),.din(w_dff_A_saxYz4xk3_0),.clk(gclk));
	jdff dff_A_7gtcvKQG4_0(.dout(w_dff_A_saxYz4xk3_0),.din(w_dff_A_7gtcvKQG4_0),.clk(gclk));
	jdff dff_A_M1IXzDpf1_0(.dout(w_dff_A_7gtcvKQG4_0),.din(w_dff_A_M1IXzDpf1_0),.clk(gclk));
	jdff dff_A_MycwKLCo4_0(.dout(w_dff_A_M1IXzDpf1_0),.din(w_dff_A_MycwKLCo4_0),.clk(gclk));
	jdff dff_A_uULW99Dd9_0(.dout(w_dff_A_MycwKLCo4_0),.din(w_dff_A_uULW99Dd9_0),.clk(gclk));
	jdff dff_A_6WBKOtYd4_0(.dout(w_dff_A_uULW99Dd9_0),.din(w_dff_A_6WBKOtYd4_0),.clk(gclk));
	jdff dff_A_uYBDJQsx0_0(.dout(w_Gid0_0[0]),.din(w_dff_A_uYBDJQsx0_0),.clk(gclk));
	jdff dff_A_17wcQfLi7_0(.dout(w_dff_A_uYBDJQsx0_0),.din(w_dff_A_17wcQfLi7_0),.clk(gclk));
	jdff dff_A_MZLrsd2A0_0(.dout(w_dff_A_17wcQfLi7_0),.din(w_dff_A_MZLrsd2A0_0),.clk(gclk));
	jdff dff_A_j8hRKf654_0(.dout(w_dff_A_MZLrsd2A0_0),.din(w_dff_A_j8hRKf654_0),.clk(gclk));
	jdff dff_A_Lvx1syXq2_0(.dout(w_dff_A_j8hRKf654_0),.din(w_dff_A_Lvx1syXq2_0),.clk(gclk));
	jdff dff_A_cMsqvbT91_0(.dout(w_dff_A_Lvx1syXq2_0),.din(w_dff_A_cMsqvbT91_0),.clk(gclk));
	jdff dff_A_2LmZU9QV5_0(.dout(w_dff_A_cMsqvbT91_0),.din(w_dff_A_2LmZU9QV5_0),.clk(gclk));
	jdff dff_A_bwssEJ8L3_0(.dout(w_dff_A_2LmZU9QV5_0),.din(w_dff_A_bwssEJ8L3_0),.clk(gclk));
	jdff dff_A_PJThdGI04_0(.dout(w_dff_A_bwssEJ8L3_0),.din(w_dff_A_PJThdGI04_0),.clk(gclk));
	jdff dff_A_OvIw5BR05_0(.dout(w_Gid12_0[0]),.din(w_dff_A_OvIw5BR05_0),.clk(gclk));
	jdff dff_A_TfB7wQkm3_0(.dout(w_dff_A_OvIw5BR05_0),.din(w_dff_A_TfB7wQkm3_0),.clk(gclk));
	jdff dff_A_YJA1BUsx9_0(.dout(w_dff_A_TfB7wQkm3_0),.din(w_dff_A_YJA1BUsx9_0),.clk(gclk));
	jdff dff_A_2K0FPSDL4_0(.dout(w_dff_A_YJA1BUsx9_0),.din(w_dff_A_2K0FPSDL4_0),.clk(gclk));
	jdff dff_A_4jIbn53j8_0(.dout(w_dff_A_2K0FPSDL4_0),.din(w_dff_A_4jIbn53j8_0),.clk(gclk));
	jdff dff_A_YGDNLoHi8_0(.dout(w_dff_A_4jIbn53j8_0),.din(w_dff_A_YGDNLoHi8_0),.clk(gclk));
	jdff dff_A_zXNrUYCE9_0(.dout(w_dff_A_YGDNLoHi8_0),.din(w_dff_A_zXNrUYCE9_0),.clk(gclk));
	jdff dff_A_ijSwMVNU0_0(.dout(w_dff_A_zXNrUYCE9_0),.din(w_dff_A_ijSwMVNU0_0),.clk(gclk));
	jdff dff_A_93gcXRbU9_0(.dout(w_dff_A_ijSwMVNU0_0),.din(w_dff_A_93gcXRbU9_0),.clk(gclk));
	jdff dff_A_hnchrOtX1_0(.dout(w_Gid8_0[0]),.din(w_dff_A_hnchrOtX1_0),.clk(gclk));
	jdff dff_A_9dIQSaS50_0(.dout(w_dff_A_hnchrOtX1_0),.din(w_dff_A_9dIQSaS50_0),.clk(gclk));
	jdff dff_A_fnQvHc5g1_0(.dout(w_dff_A_9dIQSaS50_0),.din(w_dff_A_fnQvHc5g1_0),.clk(gclk));
	jdff dff_A_OQNCr2cb7_0(.dout(w_dff_A_fnQvHc5g1_0),.din(w_dff_A_OQNCr2cb7_0),.clk(gclk));
	jdff dff_A_dtDDVJN91_0(.dout(w_dff_A_OQNCr2cb7_0),.din(w_dff_A_dtDDVJN91_0),.clk(gclk));
	jdff dff_A_f0DVnKwF7_0(.dout(w_dff_A_dtDDVJN91_0),.din(w_dff_A_f0DVnKwF7_0),.clk(gclk));
	jdff dff_A_zi4CwLtO7_0(.dout(w_dff_A_f0DVnKwF7_0),.din(w_dff_A_zi4CwLtO7_0),.clk(gclk));
	jdff dff_A_NSwSjxau6_0(.dout(w_dff_A_zi4CwLtO7_0),.din(w_dff_A_NSwSjxau6_0),.clk(gclk));
	jdff dff_A_7GamyOpk3_0(.dout(w_dff_A_NSwSjxau6_0),.din(w_dff_A_7GamyOpk3_0),.clk(gclk));
	jdff dff_B_e80MwPIa1_2(.din(n242),.dout(w_dff_B_e80MwPIa1_2),.clk(gclk));
	jdff dff_B_2IKgjRfh7_2(.din(w_dff_B_e80MwPIa1_2),.dout(w_dff_B_2IKgjRfh7_2),.clk(gclk));
	jdff dff_B_b6iKLfib8_2(.din(w_dff_B_2IKgjRfh7_2),.dout(w_dff_B_b6iKLfib8_2),.clk(gclk));
	jdff dff_A_vckJMGo81_0(.dout(w_Gid6_0[0]),.din(w_dff_A_vckJMGo81_0),.clk(gclk));
	jdff dff_A_WMI5uizx5_0(.dout(w_dff_A_vckJMGo81_0),.din(w_dff_A_WMI5uizx5_0),.clk(gclk));
	jdff dff_A_y44YarSW0_0(.dout(w_dff_A_WMI5uizx5_0),.din(w_dff_A_y44YarSW0_0),.clk(gclk));
	jdff dff_A_hWT5mOeY2_0(.dout(w_dff_A_y44YarSW0_0),.din(w_dff_A_hWT5mOeY2_0),.clk(gclk));
	jdff dff_A_l4byCqB86_0(.dout(w_dff_A_hWT5mOeY2_0),.din(w_dff_A_l4byCqB86_0),.clk(gclk));
	jdff dff_A_vRzVTpbT1_0(.dout(w_dff_A_l4byCqB86_0),.din(w_dff_A_vRzVTpbT1_0),.clk(gclk));
	jdff dff_A_q57cKHKq3_0(.dout(w_dff_A_vRzVTpbT1_0),.din(w_dff_A_q57cKHKq3_0),.clk(gclk));
	jdff dff_A_j3IkkGoM5_0(.dout(w_dff_A_q57cKHKq3_0),.din(w_dff_A_j3IkkGoM5_0),.clk(gclk));
	jdff dff_A_OxTmT3AS5_0(.dout(w_dff_A_j3IkkGoM5_0),.din(w_dff_A_OxTmT3AS5_0),.clk(gclk));
	jdff dff_A_5ZtQ9U0I5_0(.dout(w_Gid2_0[0]),.din(w_dff_A_5ZtQ9U0I5_0),.clk(gclk));
	jdff dff_A_BjHxB8iY4_0(.dout(w_dff_A_5ZtQ9U0I5_0),.din(w_dff_A_BjHxB8iY4_0),.clk(gclk));
	jdff dff_A_kwwk4Y7Q9_0(.dout(w_dff_A_BjHxB8iY4_0),.din(w_dff_A_kwwk4Y7Q9_0),.clk(gclk));
	jdff dff_A_2oZjKsiF1_0(.dout(w_dff_A_kwwk4Y7Q9_0),.din(w_dff_A_2oZjKsiF1_0),.clk(gclk));
	jdff dff_A_LRvz497N3_0(.dout(w_dff_A_2oZjKsiF1_0),.din(w_dff_A_LRvz497N3_0),.clk(gclk));
	jdff dff_A_hGfYqPSD3_0(.dout(w_dff_A_LRvz497N3_0),.din(w_dff_A_hGfYqPSD3_0),.clk(gclk));
	jdff dff_A_ZiltNOEG8_0(.dout(w_dff_A_hGfYqPSD3_0),.din(w_dff_A_ZiltNOEG8_0),.clk(gclk));
	jdff dff_A_Y0ZhjNTM5_0(.dout(w_dff_A_ZiltNOEG8_0),.din(w_dff_A_Y0ZhjNTM5_0),.clk(gclk));
	jdff dff_A_FK4WOMqW0_0(.dout(w_dff_A_Y0ZhjNTM5_0),.din(w_dff_A_FK4WOMqW0_0),.clk(gclk));
	jdff dff_A_PfitI8gt2_0(.dout(w_Gid14_0[0]),.din(w_dff_A_PfitI8gt2_0),.clk(gclk));
	jdff dff_A_GGF5EFZ77_0(.dout(w_dff_A_PfitI8gt2_0),.din(w_dff_A_GGF5EFZ77_0),.clk(gclk));
	jdff dff_A_WRyZI36C6_0(.dout(w_dff_A_GGF5EFZ77_0),.din(w_dff_A_WRyZI36C6_0),.clk(gclk));
	jdff dff_A_M3ok0lhY9_0(.dout(w_dff_A_WRyZI36C6_0),.din(w_dff_A_M3ok0lhY9_0),.clk(gclk));
	jdff dff_A_QrvOrU8h7_0(.dout(w_dff_A_M3ok0lhY9_0),.din(w_dff_A_QrvOrU8h7_0),.clk(gclk));
	jdff dff_A_LzkvNfCv8_0(.dout(w_dff_A_QrvOrU8h7_0),.din(w_dff_A_LzkvNfCv8_0),.clk(gclk));
	jdff dff_A_hr3MUg078_0(.dout(w_dff_A_LzkvNfCv8_0),.din(w_dff_A_hr3MUg078_0),.clk(gclk));
	jdff dff_A_5aET0P1v2_0(.dout(w_dff_A_hr3MUg078_0),.din(w_dff_A_5aET0P1v2_0),.clk(gclk));
	jdff dff_A_nsfUXMgG0_0(.dout(w_dff_A_5aET0P1v2_0),.din(w_dff_A_nsfUXMgG0_0),.clk(gclk));
	jdff dff_A_wEhcVPKc8_0(.dout(w_Gid10_0[0]),.din(w_dff_A_wEhcVPKc8_0),.clk(gclk));
	jdff dff_A_GQcfvTwE3_0(.dout(w_dff_A_wEhcVPKc8_0),.din(w_dff_A_GQcfvTwE3_0),.clk(gclk));
	jdff dff_A_kwEauIa30_0(.dout(w_dff_A_GQcfvTwE3_0),.din(w_dff_A_kwEauIa30_0),.clk(gclk));
	jdff dff_A_xgfgeWQi3_0(.dout(w_dff_A_kwEauIa30_0),.din(w_dff_A_xgfgeWQi3_0),.clk(gclk));
	jdff dff_A_BYJ758UH1_0(.dout(w_dff_A_xgfgeWQi3_0),.din(w_dff_A_BYJ758UH1_0),.clk(gclk));
	jdff dff_A_ueuhK2H97_0(.dout(w_dff_A_BYJ758UH1_0),.din(w_dff_A_ueuhK2H97_0),.clk(gclk));
	jdff dff_A_kZrjmoxk9_0(.dout(w_dff_A_ueuhK2H97_0),.din(w_dff_A_kZrjmoxk9_0),.clk(gclk));
	jdff dff_A_uUiUz1DW2_0(.dout(w_dff_A_kZrjmoxk9_0),.din(w_dff_A_uUiUz1DW2_0),.clk(gclk));
	jdff dff_A_Ht497OWo8_0(.dout(w_dff_A_uUiUz1DW2_0),.din(w_dff_A_Ht497OWo8_0),.clk(gclk));
	jdff dff_A_bZQMNXik2_0(.dout(w_Gid17_0[0]),.din(w_dff_A_bZQMNXik2_0),.clk(gclk));
	jdff dff_A_NFFpdhEI5_0(.dout(w_dff_A_bZQMNXik2_0),.din(w_dff_A_NFFpdhEI5_0),.clk(gclk));
	jdff dff_A_RratTCgI9_0(.dout(w_dff_A_NFFpdhEI5_0),.din(w_dff_A_RratTCgI9_0),.clk(gclk));
	jdff dff_A_SqA8iIyR8_0(.dout(w_dff_A_RratTCgI9_0),.din(w_dff_A_SqA8iIyR8_0),.clk(gclk));
	jdff dff_A_XvLAby8w2_0(.dout(w_dff_A_SqA8iIyR8_0),.din(w_dff_A_XvLAby8w2_0),.clk(gclk));
	jdff dff_A_IzZSqeq37_0(.dout(w_dff_A_XvLAby8w2_0),.din(w_dff_A_IzZSqeq37_0),.clk(gclk));
	jdff dff_A_PeIOuvWj4_0(.dout(w_dff_A_IzZSqeq37_0),.din(w_dff_A_PeIOuvWj4_0),.clk(gclk));
	jdff dff_A_LAbieiDm0_0(.dout(w_dff_A_PeIOuvWj4_0),.din(w_dff_A_LAbieiDm0_0),.clk(gclk));
	jdff dff_A_NTGyefKH4_0(.dout(w_dff_A_LAbieiDm0_0),.din(w_dff_A_NTGyefKH4_0),.clk(gclk));
	jdff dff_A_cxzokb8r0_0(.dout(w_dff_A_NTGyefKH4_0),.din(w_dff_A_cxzokb8r0_0),.clk(gclk));
	jdff dff_A_lJppg1qy9_0(.dout(w_Gid16_0[0]),.din(w_dff_A_lJppg1qy9_0),.clk(gclk));
	jdff dff_A_sptYYzdo1_0(.dout(w_dff_A_lJppg1qy9_0),.din(w_dff_A_sptYYzdo1_0),.clk(gclk));
	jdff dff_A_36yoWhlu0_0(.dout(w_dff_A_sptYYzdo1_0),.din(w_dff_A_36yoWhlu0_0),.clk(gclk));
	jdff dff_A_bMPtmkj41_0(.dout(w_dff_A_36yoWhlu0_0),.din(w_dff_A_bMPtmkj41_0),.clk(gclk));
	jdff dff_A_OdnjyUWN7_0(.dout(w_dff_A_bMPtmkj41_0),.din(w_dff_A_OdnjyUWN7_0),.clk(gclk));
	jdff dff_A_ViKR0alW7_0(.dout(w_dff_A_OdnjyUWN7_0),.din(w_dff_A_ViKR0alW7_0),.clk(gclk));
	jdff dff_A_OshFL5VS7_0(.dout(w_dff_A_ViKR0alW7_0),.din(w_dff_A_OshFL5VS7_0),.clk(gclk));
	jdff dff_A_21SCxWw11_0(.dout(w_dff_A_OshFL5VS7_0),.din(w_dff_A_21SCxWw11_0),.clk(gclk));
	jdff dff_A_R5QegjHs6_0(.dout(w_dff_A_21SCxWw11_0),.din(w_dff_A_R5QegjHs6_0),.clk(gclk));
	jdff dff_A_xcMew2LF5_0(.dout(w_dff_A_R5QegjHs6_0),.din(w_dff_A_xcMew2LF5_0),.clk(gclk));
	jdff dff_A_UZLJxiZ92_0(.dout(w_Gid19_0[0]),.din(w_dff_A_UZLJxiZ92_0),.clk(gclk));
	jdff dff_A_yGtNHZTt5_0(.dout(w_dff_A_UZLJxiZ92_0),.din(w_dff_A_yGtNHZTt5_0),.clk(gclk));
	jdff dff_A_5Hmc8qTS5_0(.dout(w_dff_A_yGtNHZTt5_0),.din(w_dff_A_5Hmc8qTS5_0),.clk(gclk));
	jdff dff_A_HSfLxjnM0_0(.dout(w_dff_A_5Hmc8qTS5_0),.din(w_dff_A_HSfLxjnM0_0),.clk(gclk));
	jdff dff_A_WEFi1sWc6_0(.dout(w_dff_A_HSfLxjnM0_0),.din(w_dff_A_WEFi1sWc6_0),.clk(gclk));
	jdff dff_A_GncTWl2v3_0(.dout(w_dff_A_WEFi1sWc6_0),.din(w_dff_A_GncTWl2v3_0),.clk(gclk));
	jdff dff_A_SpIEUzqS6_0(.dout(w_dff_A_GncTWl2v3_0),.din(w_dff_A_SpIEUzqS6_0),.clk(gclk));
	jdff dff_A_RzSmkcoq7_0(.dout(w_dff_A_SpIEUzqS6_0),.din(w_dff_A_RzSmkcoq7_0),.clk(gclk));
	jdff dff_A_QtWbALBo5_0(.dout(w_dff_A_RzSmkcoq7_0),.din(w_dff_A_QtWbALBo5_0),.clk(gclk));
	jdff dff_A_l7GTsDaa6_0(.dout(w_dff_A_QtWbALBo5_0),.din(w_dff_A_l7GTsDaa6_0),.clk(gclk));
	jdff dff_A_Gg8XAR6R1_0(.dout(w_Gid18_0[0]),.din(w_dff_A_Gg8XAR6R1_0),.clk(gclk));
	jdff dff_A_QGGOFcGh8_0(.dout(w_dff_A_Gg8XAR6R1_0),.din(w_dff_A_QGGOFcGh8_0),.clk(gclk));
	jdff dff_A_Ob80NA3b3_0(.dout(w_dff_A_QGGOFcGh8_0),.din(w_dff_A_Ob80NA3b3_0),.clk(gclk));
	jdff dff_A_8NJVnrL29_0(.dout(w_dff_A_Ob80NA3b3_0),.din(w_dff_A_8NJVnrL29_0),.clk(gclk));
	jdff dff_A_Jzk2lz6J8_0(.dout(w_dff_A_8NJVnrL29_0),.din(w_dff_A_Jzk2lz6J8_0),.clk(gclk));
	jdff dff_A_ZLpKlT7Z7_0(.dout(w_dff_A_Jzk2lz6J8_0),.din(w_dff_A_ZLpKlT7Z7_0),.clk(gclk));
	jdff dff_A_4OF9DJmF6_0(.dout(w_dff_A_ZLpKlT7Z7_0),.din(w_dff_A_4OF9DJmF6_0),.clk(gclk));
	jdff dff_A_CRAKeGGg2_0(.dout(w_dff_A_4OF9DJmF6_0),.din(w_dff_A_CRAKeGGg2_0),.clk(gclk));
	jdff dff_A_Wd6H7ox35_0(.dout(w_dff_A_CRAKeGGg2_0),.din(w_dff_A_Wd6H7ox35_0),.clk(gclk));
	jdff dff_A_4jr6RA0o0_0(.dout(w_dff_A_Wd6H7ox35_0),.din(w_dff_A_4jr6RA0o0_0),.clk(gclk));
	jdff dff_A_xLN5Qrlm2_0(.dout(w_n136_0[0]),.din(w_dff_A_xLN5Qrlm2_0),.clk(gclk));
	jdff dff_A_bP53vWSx8_0(.dout(w_Gid25_0[0]),.din(w_dff_A_bP53vWSx8_0),.clk(gclk));
	jdff dff_A_IloUHykN1_0(.dout(w_dff_A_bP53vWSx8_0),.din(w_dff_A_IloUHykN1_0),.clk(gclk));
	jdff dff_A_moLtcGR57_0(.dout(w_dff_A_IloUHykN1_0),.din(w_dff_A_moLtcGR57_0),.clk(gclk));
	jdff dff_A_t7ggL07M9_0(.dout(w_dff_A_moLtcGR57_0),.din(w_dff_A_t7ggL07M9_0),.clk(gclk));
	jdff dff_A_e0fZImGb1_0(.dout(w_dff_A_t7ggL07M9_0),.din(w_dff_A_e0fZImGb1_0),.clk(gclk));
	jdff dff_A_3QArWJJ35_0(.dout(w_dff_A_e0fZImGb1_0),.din(w_dff_A_3QArWJJ35_0),.clk(gclk));
	jdff dff_A_LMQccdJI8_0(.dout(w_dff_A_3QArWJJ35_0),.din(w_dff_A_LMQccdJI8_0),.clk(gclk));
	jdff dff_A_WV1roGcV3_0(.dout(w_dff_A_LMQccdJI8_0),.din(w_dff_A_WV1roGcV3_0),.clk(gclk));
	jdff dff_A_nfBAd0vj7_0(.dout(w_dff_A_WV1roGcV3_0),.din(w_dff_A_nfBAd0vj7_0),.clk(gclk));
	jdff dff_A_lr4aCgXD3_0(.dout(w_dff_A_nfBAd0vj7_0),.din(w_dff_A_lr4aCgXD3_0),.clk(gclk));
	jdff dff_A_OCxnHt0k2_0(.dout(w_Gid24_0[0]),.din(w_dff_A_OCxnHt0k2_0),.clk(gclk));
	jdff dff_A_Ev8pmVTN3_0(.dout(w_dff_A_OCxnHt0k2_0),.din(w_dff_A_Ev8pmVTN3_0),.clk(gclk));
	jdff dff_A_hpAXw5dq3_0(.dout(w_dff_A_Ev8pmVTN3_0),.din(w_dff_A_hpAXw5dq3_0),.clk(gclk));
	jdff dff_A_P9SqZ6Dj1_0(.dout(w_dff_A_hpAXw5dq3_0),.din(w_dff_A_P9SqZ6Dj1_0),.clk(gclk));
	jdff dff_A_C2Zl8j0U1_0(.dout(w_dff_A_P9SqZ6Dj1_0),.din(w_dff_A_C2Zl8j0U1_0),.clk(gclk));
	jdff dff_A_CCABDGb92_0(.dout(w_dff_A_C2Zl8j0U1_0),.din(w_dff_A_CCABDGb92_0),.clk(gclk));
	jdff dff_A_vWFFI2sx1_0(.dout(w_dff_A_CCABDGb92_0),.din(w_dff_A_vWFFI2sx1_0),.clk(gclk));
	jdff dff_A_bu5TOsZt2_0(.dout(w_dff_A_vWFFI2sx1_0),.din(w_dff_A_bu5TOsZt2_0),.clk(gclk));
	jdff dff_A_tteQgkbb5_0(.dout(w_dff_A_bu5TOsZt2_0),.din(w_dff_A_tteQgkbb5_0),.clk(gclk));
	jdff dff_A_OQpiXoZq8_0(.dout(w_dff_A_tteQgkbb5_0),.din(w_dff_A_OQpiXoZq8_0),.clk(gclk));
	jdff dff_A_yTlHa0bX0_0(.dout(w_Gid27_0[0]),.din(w_dff_A_yTlHa0bX0_0),.clk(gclk));
	jdff dff_A_gPILNSDl6_0(.dout(w_dff_A_yTlHa0bX0_0),.din(w_dff_A_gPILNSDl6_0),.clk(gclk));
	jdff dff_A_dTmzHv8y4_0(.dout(w_dff_A_gPILNSDl6_0),.din(w_dff_A_dTmzHv8y4_0),.clk(gclk));
	jdff dff_A_f0UrF91r0_0(.dout(w_dff_A_dTmzHv8y4_0),.din(w_dff_A_f0UrF91r0_0),.clk(gclk));
	jdff dff_A_rImIxOdU1_0(.dout(w_dff_A_f0UrF91r0_0),.din(w_dff_A_rImIxOdU1_0),.clk(gclk));
	jdff dff_A_DjH3obNe1_0(.dout(w_dff_A_rImIxOdU1_0),.din(w_dff_A_DjH3obNe1_0),.clk(gclk));
	jdff dff_A_CxycXzxt1_0(.dout(w_dff_A_DjH3obNe1_0),.din(w_dff_A_CxycXzxt1_0),.clk(gclk));
	jdff dff_A_ML2TD4h34_0(.dout(w_dff_A_CxycXzxt1_0),.din(w_dff_A_ML2TD4h34_0),.clk(gclk));
	jdff dff_A_PQ0Bq5HP4_0(.dout(w_dff_A_ML2TD4h34_0),.din(w_dff_A_PQ0Bq5HP4_0),.clk(gclk));
	jdff dff_A_Bw250faj5_0(.dout(w_dff_A_PQ0Bq5HP4_0),.din(w_dff_A_Bw250faj5_0),.clk(gclk));
	jdff dff_A_Sl5E2Pss5_0(.dout(w_Gid26_0[0]),.din(w_dff_A_Sl5E2Pss5_0),.clk(gclk));
	jdff dff_A_xeROUAR32_0(.dout(w_dff_A_Sl5E2Pss5_0),.din(w_dff_A_xeROUAR32_0),.clk(gclk));
	jdff dff_A_YOnF9Tbd0_0(.dout(w_dff_A_xeROUAR32_0),.din(w_dff_A_YOnF9Tbd0_0),.clk(gclk));
	jdff dff_A_8bpDb2Qn9_0(.dout(w_dff_A_YOnF9Tbd0_0),.din(w_dff_A_8bpDb2Qn9_0),.clk(gclk));
	jdff dff_A_kHptG9EG0_0(.dout(w_dff_A_8bpDb2Qn9_0),.din(w_dff_A_kHptG9EG0_0),.clk(gclk));
	jdff dff_A_WRxhgMmC5_0(.dout(w_dff_A_kHptG9EG0_0),.din(w_dff_A_WRxhgMmC5_0),.clk(gclk));
	jdff dff_A_DR6DxE9H1_0(.dout(w_dff_A_WRxhgMmC5_0),.din(w_dff_A_DR6DxE9H1_0),.clk(gclk));
	jdff dff_A_kLC6An7A8_0(.dout(w_dff_A_DR6DxE9H1_0),.din(w_dff_A_kLC6An7A8_0),.clk(gclk));
	jdff dff_A_CNYpowAY2_0(.dout(w_dff_A_kLC6An7A8_0),.din(w_dff_A_CNYpowAY2_0),.clk(gclk));
	jdff dff_A_uuZuWW9G7_0(.dout(w_dff_A_CNYpowAY2_0),.din(w_dff_A_uuZuWW9G7_0),.clk(gclk));
	jdff dff_A_ScXyqwmk5_0(.dout(w_n147_0[0]),.din(w_dff_A_ScXyqwmk5_0),.clk(gclk));
	jdff dff_A_SMZUDPL52_0(.dout(w_dff_A_ScXyqwmk5_0),.din(w_dff_A_SMZUDPL52_0),.clk(gclk));
	jdff dff_A_iJjnMfHd3_0(.dout(w_dff_A_SMZUDPL52_0),.din(w_dff_A_iJjnMfHd3_0),.clk(gclk));
	jdff dff_A_Lke3J96z3_0(.dout(w_dff_A_iJjnMfHd3_0),.din(w_dff_A_Lke3J96z3_0),.clk(gclk));
	jdff dff_A_fK9NmEFj1_0(.dout(w_Gid7_0[0]),.din(w_dff_A_fK9NmEFj1_0),.clk(gclk));
	jdff dff_A_1Z8L5Wlo4_0(.dout(w_dff_A_fK9NmEFj1_0),.din(w_dff_A_1Z8L5Wlo4_0),.clk(gclk));
	jdff dff_A_qtPiHYIZ1_0(.dout(w_dff_A_1Z8L5Wlo4_0),.din(w_dff_A_qtPiHYIZ1_0),.clk(gclk));
	jdff dff_A_GxhtbElV1_0(.dout(w_dff_A_qtPiHYIZ1_0),.din(w_dff_A_GxhtbElV1_0),.clk(gclk));
	jdff dff_A_4tSPT4ae0_0(.dout(w_dff_A_GxhtbElV1_0),.din(w_dff_A_4tSPT4ae0_0),.clk(gclk));
	jdff dff_A_ShVlouA69_0(.dout(w_dff_A_4tSPT4ae0_0),.din(w_dff_A_ShVlouA69_0),.clk(gclk));
	jdff dff_A_HGrhehqR4_0(.dout(w_dff_A_ShVlouA69_0),.din(w_dff_A_HGrhehqR4_0),.clk(gclk));
	jdff dff_A_yU5J5xKF7_0(.dout(w_dff_A_HGrhehqR4_0),.din(w_dff_A_yU5J5xKF7_0),.clk(gclk));
	jdff dff_A_wW1QB6Ip8_0(.dout(w_dff_A_yU5J5xKF7_0),.din(w_dff_A_wW1QB6Ip8_0),.clk(gclk));
	jdff dff_A_4eesJBAX1_0(.dout(w_Gid3_0[0]),.din(w_dff_A_4eesJBAX1_0),.clk(gclk));
	jdff dff_A_MvUKGEpP6_0(.dout(w_dff_A_4eesJBAX1_0),.din(w_dff_A_MvUKGEpP6_0),.clk(gclk));
	jdff dff_A_CtIGVonJ4_0(.dout(w_dff_A_MvUKGEpP6_0),.din(w_dff_A_CtIGVonJ4_0),.clk(gclk));
	jdff dff_A_in8dp6GF0_0(.dout(w_dff_A_CtIGVonJ4_0),.din(w_dff_A_in8dp6GF0_0),.clk(gclk));
	jdff dff_A_6GlIiAI46_0(.dout(w_dff_A_in8dp6GF0_0),.din(w_dff_A_6GlIiAI46_0),.clk(gclk));
	jdff dff_A_n2YyPnyt8_0(.dout(w_dff_A_6GlIiAI46_0),.din(w_dff_A_n2YyPnyt8_0),.clk(gclk));
	jdff dff_A_8PAiNZnn2_0(.dout(w_dff_A_n2YyPnyt8_0),.din(w_dff_A_8PAiNZnn2_0),.clk(gclk));
	jdff dff_A_5ukHwWHE2_0(.dout(w_dff_A_8PAiNZnn2_0),.din(w_dff_A_5ukHwWHE2_0),.clk(gclk));
	jdff dff_A_fXFBxHfN8_0(.dout(w_dff_A_5ukHwWHE2_0),.din(w_dff_A_fXFBxHfN8_0),.clk(gclk));
	jdff dff_A_2xJHH95p7_0(.dout(w_Gid15_0[0]),.din(w_dff_A_2xJHH95p7_0),.clk(gclk));
	jdff dff_A_GW7inNXo9_0(.dout(w_dff_A_2xJHH95p7_0),.din(w_dff_A_GW7inNXo9_0),.clk(gclk));
	jdff dff_A_CIWDgkaH6_0(.dout(w_dff_A_GW7inNXo9_0),.din(w_dff_A_CIWDgkaH6_0),.clk(gclk));
	jdff dff_A_EEZ76ch47_0(.dout(w_dff_A_CIWDgkaH6_0),.din(w_dff_A_EEZ76ch47_0),.clk(gclk));
	jdff dff_A_XfsGqQgH9_0(.dout(w_dff_A_EEZ76ch47_0),.din(w_dff_A_XfsGqQgH9_0),.clk(gclk));
	jdff dff_A_hP9CgISz6_0(.dout(w_dff_A_XfsGqQgH9_0),.din(w_dff_A_hP9CgISz6_0),.clk(gclk));
	jdff dff_A_59J9n2YU4_0(.dout(w_dff_A_hP9CgISz6_0),.din(w_dff_A_59J9n2YU4_0),.clk(gclk));
	jdff dff_A_7Qkv7wzY2_0(.dout(w_dff_A_59J9n2YU4_0),.din(w_dff_A_7Qkv7wzY2_0),.clk(gclk));
	jdff dff_A_W47mm7Ai1_0(.dout(w_dff_A_7Qkv7wzY2_0),.din(w_dff_A_W47mm7Ai1_0),.clk(gclk));
	jdff dff_A_dmj8I8wf4_0(.dout(w_Gid11_0[0]),.din(w_dff_A_dmj8I8wf4_0),.clk(gclk));
	jdff dff_A_B7KuEblU4_0(.dout(w_dff_A_dmj8I8wf4_0),.din(w_dff_A_B7KuEblU4_0),.clk(gclk));
	jdff dff_A_ZOKuz7Gy1_0(.dout(w_dff_A_B7KuEblU4_0),.din(w_dff_A_ZOKuz7Gy1_0),.clk(gclk));
	jdff dff_A_6BDMHWkN3_0(.dout(w_dff_A_ZOKuz7Gy1_0),.din(w_dff_A_6BDMHWkN3_0),.clk(gclk));
	jdff dff_A_78wyfkzn7_0(.dout(w_dff_A_6BDMHWkN3_0),.din(w_dff_A_78wyfkzn7_0),.clk(gclk));
	jdff dff_A_g81HgcgD1_0(.dout(w_dff_A_78wyfkzn7_0),.din(w_dff_A_g81HgcgD1_0),.clk(gclk));
	jdff dff_A_Uc3xER899_0(.dout(w_dff_A_g81HgcgD1_0),.din(w_dff_A_Uc3xER899_0),.clk(gclk));
	jdff dff_A_f5HW29mj7_0(.dout(w_dff_A_Uc3xER899_0),.din(w_dff_A_f5HW29mj7_0),.clk(gclk));
	jdff dff_A_9ho4Nn9t4_0(.dout(w_dff_A_f5HW29mj7_0),.din(w_dff_A_9ho4Nn9t4_0),.clk(gclk));
	jdff dff_A_WCTX8HK26_0(.dout(w_Gid21_0[0]),.din(w_dff_A_WCTX8HK26_0),.clk(gclk));
	jdff dff_A_fQt3MjJe2_0(.dout(w_dff_A_WCTX8HK26_0),.din(w_dff_A_fQt3MjJe2_0),.clk(gclk));
	jdff dff_A_v9K8nSWP6_0(.dout(w_dff_A_fQt3MjJe2_0),.din(w_dff_A_v9K8nSWP6_0),.clk(gclk));
	jdff dff_A_qkUgSe8V2_0(.dout(w_dff_A_v9K8nSWP6_0),.din(w_dff_A_qkUgSe8V2_0),.clk(gclk));
	jdff dff_A_NwUPZEmv6_0(.dout(w_dff_A_qkUgSe8V2_0),.din(w_dff_A_NwUPZEmv6_0),.clk(gclk));
	jdff dff_A_vwV6qDiY0_0(.dout(w_dff_A_NwUPZEmv6_0),.din(w_dff_A_vwV6qDiY0_0),.clk(gclk));
	jdff dff_A_UePXeYo52_0(.dout(w_dff_A_vwV6qDiY0_0),.din(w_dff_A_UePXeYo52_0),.clk(gclk));
	jdff dff_A_90vmAjC44_0(.dout(w_dff_A_UePXeYo52_0),.din(w_dff_A_90vmAjC44_0),.clk(gclk));
	jdff dff_A_SV73FUkl9_0(.dout(w_dff_A_90vmAjC44_0),.din(w_dff_A_SV73FUkl9_0),.clk(gclk));
	jdff dff_A_hoRlUHJb5_0(.dout(w_dff_A_SV73FUkl9_0),.din(w_dff_A_hoRlUHJb5_0),.clk(gclk));
	jdff dff_A_XAjfJZzc0_0(.dout(w_Gid20_0[0]),.din(w_dff_A_XAjfJZzc0_0),.clk(gclk));
	jdff dff_A_LvdBae3g4_0(.dout(w_dff_A_XAjfJZzc0_0),.din(w_dff_A_LvdBae3g4_0),.clk(gclk));
	jdff dff_A_A0Gs43go1_0(.dout(w_dff_A_LvdBae3g4_0),.din(w_dff_A_A0Gs43go1_0),.clk(gclk));
	jdff dff_A_B0JUY8yP9_0(.dout(w_dff_A_A0Gs43go1_0),.din(w_dff_A_B0JUY8yP9_0),.clk(gclk));
	jdff dff_A_URhjdKHN2_0(.dout(w_dff_A_B0JUY8yP9_0),.din(w_dff_A_URhjdKHN2_0),.clk(gclk));
	jdff dff_A_LCjiDUSI8_0(.dout(w_dff_A_URhjdKHN2_0),.din(w_dff_A_LCjiDUSI8_0),.clk(gclk));
	jdff dff_A_ANmPxrNb0_0(.dout(w_dff_A_LCjiDUSI8_0),.din(w_dff_A_ANmPxrNb0_0),.clk(gclk));
	jdff dff_A_NWEpgtfT4_0(.dout(w_dff_A_ANmPxrNb0_0),.din(w_dff_A_NWEpgtfT4_0),.clk(gclk));
	jdff dff_A_ZyKiFDdL6_0(.dout(w_dff_A_NWEpgtfT4_0),.din(w_dff_A_ZyKiFDdL6_0),.clk(gclk));
	jdff dff_A_aElP0Gp81_0(.dout(w_dff_A_ZyKiFDdL6_0),.din(w_dff_A_aElP0Gp81_0),.clk(gclk));
	jdff dff_A_pHA9rxW93_0(.dout(w_Gid23_0[0]),.din(w_dff_A_pHA9rxW93_0),.clk(gclk));
	jdff dff_A_niuqIfuV8_0(.dout(w_dff_A_pHA9rxW93_0),.din(w_dff_A_niuqIfuV8_0),.clk(gclk));
	jdff dff_A_nKKuTyWB0_0(.dout(w_dff_A_niuqIfuV8_0),.din(w_dff_A_nKKuTyWB0_0),.clk(gclk));
	jdff dff_A_S6Ku3KxG9_0(.dout(w_dff_A_nKKuTyWB0_0),.din(w_dff_A_S6Ku3KxG9_0),.clk(gclk));
	jdff dff_A_iJEMv04R5_0(.dout(w_dff_A_S6Ku3KxG9_0),.din(w_dff_A_iJEMv04R5_0),.clk(gclk));
	jdff dff_A_BHGmYrIy3_0(.dout(w_dff_A_iJEMv04R5_0),.din(w_dff_A_BHGmYrIy3_0),.clk(gclk));
	jdff dff_A_U7zZCN2Q6_0(.dout(w_dff_A_BHGmYrIy3_0),.din(w_dff_A_U7zZCN2Q6_0),.clk(gclk));
	jdff dff_A_lJjb7aA84_0(.dout(w_dff_A_U7zZCN2Q6_0),.din(w_dff_A_lJjb7aA84_0),.clk(gclk));
	jdff dff_A_jvnZxQgd4_0(.dout(w_dff_A_lJjb7aA84_0),.din(w_dff_A_jvnZxQgd4_0),.clk(gclk));
	jdff dff_A_13P3eB4r7_0(.dout(w_dff_A_jvnZxQgd4_0),.din(w_dff_A_13P3eB4r7_0),.clk(gclk));
	jdff dff_A_NNrpbb4M1_0(.dout(w_Gid22_0[0]),.din(w_dff_A_NNrpbb4M1_0),.clk(gclk));
	jdff dff_A_EH4UGlAo3_0(.dout(w_dff_A_NNrpbb4M1_0),.din(w_dff_A_EH4UGlAo3_0),.clk(gclk));
	jdff dff_A_4488NkMZ3_0(.dout(w_dff_A_EH4UGlAo3_0),.din(w_dff_A_4488NkMZ3_0),.clk(gclk));
	jdff dff_A_MOmIMwaP9_0(.dout(w_dff_A_4488NkMZ3_0),.din(w_dff_A_MOmIMwaP9_0),.clk(gclk));
	jdff dff_A_4wZLjRTf5_0(.dout(w_dff_A_MOmIMwaP9_0),.din(w_dff_A_4wZLjRTf5_0),.clk(gclk));
	jdff dff_A_64vW8LYs2_0(.dout(w_dff_A_4wZLjRTf5_0),.din(w_dff_A_64vW8LYs2_0),.clk(gclk));
	jdff dff_A_T6SZeMnp1_0(.dout(w_dff_A_64vW8LYs2_0),.din(w_dff_A_T6SZeMnp1_0),.clk(gclk));
	jdff dff_A_muIWvRze2_0(.dout(w_dff_A_T6SZeMnp1_0),.din(w_dff_A_muIWvRze2_0),.clk(gclk));
	jdff dff_A_es3LB2bb6_0(.dout(w_dff_A_muIWvRze2_0),.din(w_dff_A_es3LB2bb6_0),.clk(gclk));
	jdff dff_A_O6iHzNyD7_0(.dout(w_dff_A_es3LB2bb6_0),.din(w_dff_A_O6iHzNyD7_0),.clk(gclk));
	jdff dff_A_6ozCoOJb2_0(.dout(w_n128_0[0]),.din(w_dff_A_6ozCoOJb2_0),.clk(gclk));
	jdff dff_A_Rv2ewegQ6_0(.dout(w_Gid29_0[0]),.din(w_dff_A_Rv2ewegQ6_0),.clk(gclk));
	jdff dff_A_OR6pGGhO9_0(.dout(w_dff_A_Rv2ewegQ6_0),.din(w_dff_A_OR6pGGhO9_0),.clk(gclk));
	jdff dff_A_q9qdLaP40_0(.dout(w_dff_A_OR6pGGhO9_0),.din(w_dff_A_q9qdLaP40_0),.clk(gclk));
	jdff dff_A_OLbfuIra7_0(.dout(w_dff_A_q9qdLaP40_0),.din(w_dff_A_OLbfuIra7_0),.clk(gclk));
	jdff dff_A_HIJJWWz61_0(.dout(w_dff_A_OLbfuIra7_0),.din(w_dff_A_HIJJWWz61_0),.clk(gclk));
	jdff dff_A_LT7ZlOYt8_0(.dout(w_dff_A_HIJJWWz61_0),.din(w_dff_A_LT7ZlOYt8_0),.clk(gclk));
	jdff dff_A_t6ipZzDX6_0(.dout(w_dff_A_LT7ZlOYt8_0),.din(w_dff_A_t6ipZzDX6_0),.clk(gclk));
	jdff dff_A_DQCSUQqG6_0(.dout(w_dff_A_t6ipZzDX6_0),.din(w_dff_A_DQCSUQqG6_0),.clk(gclk));
	jdff dff_A_svqLrh3p5_0(.dout(w_dff_A_DQCSUQqG6_0),.din(w_dff_A_svqLrh3p5_0),.clk(gclk));
	jdff dff_A_GkSNTNLK1_0(.dout(w_dff_A_svqLrh3p5_0),.din(w_dff_A_GkSNTNLK1_0),.clk(gclk));
	jdff dff_A_smRNJj5V0_0(.dout(w_Gid28_0[0]),.din(w_dff_A_smRNJj5V0_0),.clk(gclk));
	jdff dff_A_g7AvD1lU2_0(.dout(w_dff_A_smRNJj5V0_0),.din(w_dff_A_g7AvD1lU2_0),.clk(gclk));
	jdff dff_A_MXBC8gwc7_0(.dout(w_dff_A_g7AvD1lU2_0),.din(w_dff_A_MXBC8gwc7_0),.clk(gclk));
	jdff dff_A_XXgimxdL0_0(.dout(w_dff_A_MXBC8gwc7_0),.din(w_dff_A_XXgimxdL0_0),.clk(gclk));
	jdff dff_A_BOD9uQUq4_0(.dout(w_dff_A_XXgimxdL0_0),.din(w_dff_A_BOD9uQUq4_0),.clk(gclk));
	jdff dff_A_nkiiWIQD4_0(.dout(w_dff_A_BOD9uQUq4_0),.din(w_dff_A_nkiiWIQD4_0),.clk(gclk));
	jdff dff_A_y59Z0jRU0_0(.dout(w_dff_A_nkiiWIQD4_0),.din(w_dff_A_y59Z0jRU0_0),.clk(gclk));
	jdff dff_A_pFiZV1U81_0(.dout(w_dff_A_y59Z0jRU0_0),.din(w_dff_A_pFiZV1U81_0),.clk(gclk));
	jdff dff_A_WBkR5y0F6_0(.dout(w_dff_A_pFiZV1U81_0),.din(w_dff_A_WBkR5y0F6_0),.clk(gclk));
	jdff dff_A_D5KmenKw5_0(.dout(w_dff_A_WBkR5y0F6_0),.din(w_dff_A_D5KmenKw5_0),.clk(gclk));
	jdff dff_A_GQ9VcaOp6_0(.dout(w_Gid31_0[0]),.din(w_dff_A_GQ9VcaOp6_0),.clk(gclk));
	jdff dff_A_p1WKOqjt3_0(.dout(w_dff_A_GQ9VcaOp6_0),.din(w_dff_A_p1WKOqjt3_0),.clk(gclk));
	jdff dff_A_4lo1HaQU6_0(.dout(w_dff_A_p1WKOqjt3_0),.din(w_dff_A_4lo1HaQU6_0),.clk(gclk));
	jdff dff_A_6V26NkQY9_0(.dout(w_dff_A_4lo1HaQU6_0),.din(w_dff_A_6V26NkQY9_0),.clk(gclk));
	jdff dff_A_tSQ47dtz9_0(.dout(w_dff_A_6V26NkQY9_0),.din(w_dff_A_tSQ47dtz9_0),.clk(gclk));
	jdff dff_A_aebaVOIH5_0(.dout(w_dff_A_tSQ47dtz9_0),.din(w_dff_A_aebaVOIH5_0),.clk(gclk));
	jdff dff_A_H2K6atbm7_0(.dout(w_dff_A_aebaVOIH5_0),.din(w_dff_A_H2K6atbm7_0),.clk(gclk));
	jdff dff_A_JLCdQGQ26_0(.dout(w_dff_A_H2K6atbm7_0),.din(w_dff_A_JLCdQGQ26_0),.clk(gclk));
	jdff dff_A_vodje6d04_0(.dout(w_dff_A_JLCdQGQ26_0),.din(w_dff_A_vodje6d04_0),.clk(gclk));
	jdff dff_A_PDVxLHao2_0(.dout(w_dff_A_vodje6d04_0),.din(w_dff_A_PDVxLHao2_0),.clk(gclk));
	jdff dff_A_73iZggXs5_0(.dout(w_Gid30_0[0]),.din(w_dff_A_73iZggXs5_0),.clk(gclk));
	jdff dff_A_moRPC7wp3_0(.dout(w_dff_A_73iZggXs5_0),.din(w_dff_A_moRPC7wp3_0),.clk(gclk));
	jdff dff_A_Mp2833Jr3_0(.dout(w_dff_A_moRPC7wp3_0),.din(w_dff_A_Mp2833Jr3_0),.clk(gclk));
	jdff dff_A_TcFPoXcA1_0(.dout(w_dff_A_Mp2833Jr3_0),.din(w_dff_A_TcFPoXcA1_0),.clk(gclk));
	jdff dff_A_VIYnC5J50_0(.dout(w_dff_A_TcFPoXcA1_0),.din(w_dff_A_VIYnC5J50_0),.clk(gclk));
	jdff dff_A_2Z9XcLd81_0(.dout(w_dff_A_VIYnC5J50_0),.din(w_dff_A_2Z9XcLd81_0),.clk(gclk));
	jdff dff_A_odOsKShW0_0(.dout(w_dff_A_2Z9XcLd81_0),.din(w_dff_A_odOsKShW0_0),.clk(gclk));
	jdff dff_A_gAk31LJm6_0(.dout(w_dff_A_odOsKShW0_0),.din(w_dff_A_gAk31LJm6_0),.clk(gclk));
	jdff dff_A_OMF8t8vb2_0(.dout(w_dff_A_gAk31LJm6_0),.din(w_dff_A_OMF8t8vb2_0),.clk(gclk));
	jdff dff_A_QfoNNBsi3_0(.dout(w_dff_A_OMF8t8vb2_0),.din(w_dff_A_QfoNNBsi3_0),.clk(gclk));
endmodule

