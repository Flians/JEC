module rf_c499(Gic4, Gic2, Gid31, Gid30, Gid28, Gid10, Gic0, Gid8, Gid4, Gid2, Gic6, Gid14, Gid7, Gid15, Gid5, Gid1, Gid6, Gid11, Gic5, Gid9, Gic3, Gid25, Gid12, Gid0, Gr, Gic1, Gid13, Gid29, Gid16, Gid21, Gid17, Gid18, Gid22, Gid3, Gid19, Gic7, Gid23, Gid24, Gid26, Gid20, Gid27, God31, God30, God29, God9, God24, God10, God8, God16, God25, God19, God7, God11, God13, God6, God4, God17, God12, God23, God3, God2, God1, God0, God14, God15, God22, God20, God21, God5, God18, God26, God27, God28);
    input Gic4, Gic2, Gid31, Gid30, Gid28, Gid10, Gic0, Gid8, Gid4, Gid2, Gic6, Gid14, Gid7, Gid15, Gid5, Gid1, Gid6, Gid11, Gic5, Gid9, Gic3, Gid25, Gid12, Gid0, Gr, Gic1, Gid13, Gid29, Gid16, Gid21, Gid17, Gid18, Gid22, Gid3, Gid19, Gic7, Gid23, Gid24, Gid26, Gid20, Gid27;
    output God31, God30, God29, God9, God24, God10, God8, God16, God25, God19, God7, God11, God13, God6, God4, God17, God12, God23, God3, God2, God1, God0, God14, God15, God22, God20, God21, God5, God18, God26, God27, God28;
    wire n75;
    wire n78;
    wire n82;
    wire n86;
    wire n90;
    wire n94;
    wire n98;
    wire n102;
    wire n106;
    wire n110;
    wire n114;
    wire n118;
    wire n122;
    wire n126;
    wire n130;
    wire n133;
    wire n136;
    wire n140;
    wire n144;
    wire n148;
    wire n152;
    wire n156;
    wire n160;
    wire n164;
    wire n168;
    wire n172;
    wire n176;
    wire n180;
    wire n184;
    wire n188;
    wire n191;
    wire n195;
    wire n199;
    wire n203;
    wire n207;
    wire n211;
    wire n215;
    wire n219;
    wire n223;
    wire n227;
    wire n231;
    wire n235;
    wire n239;
    wire n243;
    wire n246;
    wire n250;
    wire n253;
    wire n257;
    wire n261;
    wire n265;
    wire n269;
    wire n273;
    wire n277;
    wire n281;
    wire n284;
    wire n287;
    wire n291;
    wire n295;
    wire n299;
    wire n303;
    wire n307;
    wire n311;
    wire n315;
    wire n319;
    wire n322;
    wire n326;
    wire n330;
    wire n334;
    wire n338;
    wire n342;
    wire n346;
    wire n350;
    wire n354;
    wire n358;
    wire n362;
    wire n366;
    wire n370;
    wire n374;
    wire n378;
    wire n381;
    wire n385;
    wire n389;
    wire n393;
    wire n397;
    wire n401;
    wire n405;
    wire n409;
    wire n412;
    wire n416;
    wire n420;
    wire n424;
    wire n428;
    wire n432;
    wire n436;
    wire n440;
    wire n444;
    wire n448;
    wire n452;
    wire n456;
    wire n460;
    wire n464;
    wire n468;
    wire n472;
    wire n476;
    wire n483;
    wire n487;
    wire n494;
    wire n498;
    wire n505;
    wire n509;
    wire n516;
    wire n520;
    wire n524;
    wire n528;
    wire n536;
    wire n544;
    wire n552;
    wire n559;
    wire n563;
    wire n567;
    wire n571;
    wire n575;
    wire n579;
    wire n583;
    wire n587;
    wire n591;
    wire n595;
    wire n599;
    wire n603;
    wire n607;
    wire n611;
    wire n615;
    wire n619;
    wire n623;
    wire n627;
    wire n631;
    wire n635;
    wire n639;
    wire n643;
    wire n647;
    wire n651;
    wire n655;
    wire n659;
    wire n663;
    wire n667;
    wire n671;
    wire n675;
    wire n679;
    wire n683;
    wire n687;
    wire n691;
    wire n699;
    wire n707;
    wire n715;
    wire n723;
    wire n727;
    wire n731;
    wire n735;
    wire n743;
    wire n751;
    wire n759;
    wire n767;
    wire n771;
    wire n775;
    wire n783;
    wire n791;
    wire n799;
    wire n807;
    wire n811;
    wire n819;
    wire n827;
    wire n835;
    wire n1216;
    wire n1218;
    wire n1221;
    wire n1224;
    wire n1227;
    wire n1230;
    wire n1233;
    wire n1236;
    wire n1239;
    wire n1242;
    wire n1245;
    wire n1248;
    wire n1251;
    wire n1254;
    wire n1257;
    wire n1260;
    wire n1263;
    wire n1266;
    wire n1269;
    wire n1272;
    wire n1275;
    wire n1278;
    wire n1281;
    wire n1284;
    wire n1287;
    wire n1290;
    wire n1293;
    wire n1296;
    wire n1299;
    wire n1302;
    wire n1305;
    wire n1308;
    wire n1311;
    wire n1314;
    wire n1317;
    wire n1320;
    wire n1323;
    wire n1327;
    wire n1330;
    wire n1332;
    wire n1335;
    wire n1338;
    wire n1341;
    wire n1344;
    wire n1347;
    wire n1350;
    wire n1353;
    wire n1356;
    wire n1359;
    wire n1362;
    wire n1365;
    wire n1368;
    wire n1371;
    wire n1375;
    wire n1377;
    wire n1380;
    wire n1383;
    wire n1386;
    wire n1389;
    wire n1392;
    wire n1395;
    wire n1398;
    wire n1401;
    wire n1404;
    wire n1407;
    wire n1410;
    wire n1413;
    wire n1416;
    wire n1419;
    wire n1422;
    wire n1425;
    wire n1428;
    wire n1431;
    wire n1434;
    wire n1437;
    wire n1440;
    wire n1443;
    wire n1446;
    wire n1449;
    wire n1452;
    wire n1455;
    wire n1458;
    wire n1461;
    wire n1464;
    wire n1467;
    wire n1470;
    wire n1473;
    wire n1477;
    wire n1479;
    wire n1482;
    wire n1485;
    wire n1488;
    wire n1491;
    wire n1494;
    wire n1497;
    wire n1500;
    wire n1503;
    wire n1506;
    wire n1509;
    wire n1512;
    wire n1515;
    wire n1518;
    wire n1521;
    wire n1524;
    wire n1527;
    wire n1530;
    wire n1533;
    wire n1536;
    wire n1539;
    wire n1542;
    wire n1545;
    wire n1548;
    wire n1551;
    wire n1554;
    wire n1557;
    wire n1560;
    wire n1563;
    wire n1566;
    wire n1569;
    wire n1572;
    wire n1575;
    wire n1578;
    wire n1581;
    wire n1584;
    wire n1587;
    wire n1590;
    wire n1593;
    wire n1596;
    wire n1599;
    wire n1602;
    wire n1605;
    wire n1608;
    wire n1611;
    wire n1614;
    wire n1618;
    wire n1621;
    wire n1623;
    wire n1626;
    wire n1629;
    wire n1632;
    wire n1635;
    wire n1638;
    wire n1641;
    wire n1644;
    wire n1647;
    wire n1650;
    wire n1653;
    wire n1656;
    wire n1659;
    wire n1662;
    wire n1665;
    wire n1668;
    wire n1671;
    wire n1674;
    wire n1677;
    wire n1680;
    wire n1683;
    wire n1686;
    wire n1689;
    wire n1692;
    wire n1695;
    wire n1698;
    wire n1701;
    wire n1704;
    wire n1707;
    wire n1710;
    wire n1713;
    wire n1716;
    wire n1719;
    wire n1722;
    wire n1725;
    wire n1728;
    wire n1731;
    wire n1734;
    wire n1737;
    wire n1740;
    wire n1743;
    wire n1746;
    wire n1749;
    wire n1752;
    wire n1755;
    wire n1758;
    wire n1761;
    wire n1764;
    wire n1767;
    wire n1770;
    wire n1773;
    wire n1776;
    wire n1779;
    wire n1782;
    wire n1785;
    wire n1788;
    wire n1791;
    wire n1794;
    wire n1797;
    wire n1800;
    wire n1803;
    wire n1806;
    wire n1809;
    wire n1812;
    wire n1815;
    wire n1818;
    wire n1821;
    wire n1824;
    wire n1827;
    wire n1830;
    wire n1833;
    wire n1836;
    wire n1839;
    wire n1842;
    wire n1845;
    wire n1848;
    wire n1851;
    wire n1854;
    wire n1857;
    wire n1860;
    wire n1863;
    wire n1866;
    wire n1869;
    wire n1872;
    wire n1875;
    wire n1878;
    wire n1881;
    wire n1884;
    wire n1887;
    wire n1890;
    wire n1893;
    wire n1896;
    wire n1899;
    wire n1902;
    wire n1905;
    wire n1908;
    wire n1911;
    wire n1914;
    wire n1917;
    wire n1920;
    wire n1923;
    wire n1926;
    wire n1929;
    wire n1932;
    wire n1935;
    wire n1938;
    wire n1941;
    wire n1944;
    wire n1947;
    wire n1950;
    wire n1953;
    wire n1956;
    wire n1959;
    wire n1962;
    wire n1965;
    wire n1968;
    wire n1971;
    wire n1974;
    wire n1977;
    wire n1980;
    wire n1983;
    wire n1986;
    wire n1989;
    wire n1992;
    wire n1995;
    wire n1998;
    wire n2001;
    wire n2004;
    wire n2007;
    wire n2010;
    wire n2013;
    wire n2016;
    wire n2019;
    wire n2022;
    wire n2025;
    wire n2028;
    wire n2031;
    wire n2034;
    wire n2037;
    wire n2040;
    wire n2043;
    wire n2046;
    wire n2049;
    wire n2052;
    wire n2055;
    wire n2058;
    wire n2061;
    wire n2064;
    wire n2067;
    wire n2070;
    wire n2073;
    wire n2076;
    wire n2079;
    wire n2082;
    wire n2085;
    wire n2088;
    wire n2091;
    wire n2094;
    wire n2097;
    wire n2100;
    wire n2103;
    wire n2106;
    wire n2109;
    wire n2112;
    wire n2115;
    wire n2118;
    wire n2121;
    wire n2124;
    wire n2127;
    wire n2130;
    wire n2133;
    wire n2136;
    wire n2139;
    wire n2142;
    wire n2145;
    wire n2148;
    wire n2151;
    wire n2154;
    wire n2157;
    wire n2160;
    wire n2163;
    wire n2166;
    wire n2169;
    wire n2172;
    wire n2175;
    wire n2178;
    wire n2181;
    wire n2184;
    wire n2187;
    wire n2190;
    wire n2193;
    wire n2196;
    wire n2199;
    wire n2202;
    wire n2205;
    wire n2208;
    wire n2211;
    wire n2214;
    wire n2217;
    wire n2220;
    wire n2223;
    wire n2226;
    wire n2229;
    wire n2232;
    wire n2235;
    wire n2238;
    wire n2241;
    wire n2244;
    wire n2247;
    wire n2250;
    wire n2253;
    wire n2256;
    wire n2259;
    wire n2262;
    wire n2265;
    wire n2268;
    wire n2271;
    wire n2274;
    wire n2277;
    wire n2280;
    wire n2283;
    wire n2286;
    wire n2289;
    wire n2292;
    wire n2295;
    wire n2298;
    wire n2301;
    wire n2304;
    wire n2307;
    wire n2310;
    wire n2313;
    wire n2316;
    wire n2319;
    wire n2322;
    wire n2325;
    wire n2328;
    wire n2331;
    wire n2334;
    wire n2337;
    wire n2340;
    wire n2343;
    wire n2346;
    wire n2349;
    wire n2352;
    wire n2355;
    wire n2358;
    wire n2361;
    wire n2364;
    wire n2367;
    wire n2370;
    wire n2373;
    wire n2376;
    wire n2379;
    wire n2382;
    wire n2385;
    wire n2388;
    wire n2391;
    wire n2394;
    wire n2397;
    wire n2400;
    wire n2403;
    wire n2406;
    wire n2409;
    wire n2412;
    wire n2415;
    wire n2418;
    wire n2421;
    wire n2424;
    wire n2427;
    wire n2430;
    wire n2433;
    wire n2436;
    wire n2439;
    wire n2442;
    wire n2445;
    wire n2448;
    wire n2451;
    wire n2454;
    wire n2457;
    wire n2460;
    wire n2463;
    wire n2466;
    wire n2469;
    wire n2472;
    wire n2475;
    wire n2478;
    wire n2481;
    wire n2484;
    wire n2487;
    wire n2490;
    wire n2493;
    jnot g000(.din(Gic0), .dout(n75));
    jnot g001(.din(Gr), .dout(n78));
    jor g002(.dinb(n75), .dina(n78), .dout(n82));
    jxor g003(.dinb(Gid16), .dina(Gid17), .dout(n86));
    jxor g004(.dinb(Gid18), .dina(Gid19), .dout(n90));
    jxor g005(.dinb(n86), .dina(n90), .dout(n94));
    jxor g006(.dinb(n82), .dina(n94), .dout(n98));
    jxor g007(.dinb(Gid0), .dina(Gid4), .dout(n102));
    jxor g008(.dinb(Gid8), .dina(Gid12), .dout(n106));
    jxor g009(.dinb(n102), .dina(n106), .dout(n110));
    jxor g010(.dinb(Gid20), .dina(Gid21), .dout(n114));
    jxor g011(.dinb(Gid22), .dina(Gid23), .dout(n118));
    jxor g012(.dinb(n114), .dina(n118), .dout(n122));
    jxor g013(.dinb(n110), .dina(n122), .dout(n126));
    jxor g014(.dinb(n98), .dina(n126), .dout(n130));
    jnot g015(.din(n130), .dout(n133));
    jnot g016(.din(Gic7), .dout(n136));
    jor g017(.dinb(n136), .dina(n78), .dout(n140));
    jxor g018(.dinb(Gid4), .dina(Gid5), .dout(n144));
    jxor g019(.dinb(Gid6), .dina(Gid7), .dout(n148));
    jxor g020(.dinb(n144), .dina(n148), .dout(n152));
    jxor g021(.dinb(n140), .dina(n152), .dout(n156));
    jxor g022(.dinb(Gid12), .dina(Gid13), .dout(n160));
    jxor g023(.dinb(Gid14), .dina(Gid15), .dout(n164));
    jxor g024(.dinb(n160), .dina(n164), .dout(n168));
    jxor g025(.dinb(Gid19), .dina(Gid23), .dout(n172));
    jxor g026(.dinb(Gid27), .dina(Gid31), .dout(n176));
    jxor g027(.dinb(n172), .dina(n176), .dout(n180));
    jxor g028(.dinb(n168), .dina(n180), .dout(n184));
    jxor g029(.dinb(n156), .dina(n184), .dout(n188));
    jnot g030(.din(Gic6), .dout(n191));
    jor g031(.dinb(n191), .dina(n78), .dout(n195));
    jxor g032(.dinb(Gid0), .dina(Gid1), .dout(n199));
    jxor g033(.dinb(Gid2), .dina(Gid3), .dout(n203));
    jxor g034(.dinb(n199), .dina(n203), .dout(n207));
    jxor g035(.dinb(n195), .dina(n207), .dout(n211));
    jxor g036(.dinb(Gid8), .dina(Gid9), .dout(n215));
    jxor g037(.dinb(Gid10), .dina(Gid11), .dout(n219));
    jxor g038(.dinb(n215), .dina(n219), .dout(n223));
    jxor g039(.dinb(Gid18), .dina(Gid22), .dout(n227));
    jxor g040(.dinb(Gid26), .dina(Gid30), .dout(n231));
    jxor g041(.dinb(n227), .dina(n231), .dout(n235));
    jxor g042(.dinb(n223), .dina(n235), .dout(n239));
    jxor g043(.dinb(n211), .dina(n239), .dout(n243));
    jnot g044(.din(n243), .dout(n246));
    jand g045(.dinb(n2145), .dina(n246), .dout(n250));
    jnot g046(.din(Gic4), .dout(n253));
    jor g047(.dinb(n253), .dina(n78), .dout(n257));
    jxor g048(.dinb(n152), .dina(n257), .dout(n261));
    jxor g049(.dinb(Gid16), .dina(Gid20), .dout(n265));
    jxor g050(.dinb(Gid24), .dina(Gid28), .dout(n269));
    jxor g051(.dinb(n265), .dina(n269), .dout(n273));
    jxor g052(.dinb(n207), .dina(n273), .dout(n277));
    jxor g053(.dinb(n261), .dina(n277), .dout(n281));
    jnot g054(.din(n281), .dout(n284));
    jnot g055(.din(Gic5), .dout(n287));
    jor g056(.dinb(n287), .dina(n78), .dout(n291));
    jxor g057(.dinb(n168), .dina(n291), .dout(n295));
    jxor g058(.dinb(Gid17), .dina(Gid21), .dout(n299));
    jxor g059(.dinb(Gid25), .dina(Gid29), .dout(n303));
    jxor g060(.dinb(n299), .dina(n303), .dout(n307));
    jxor g061(.dinb(n223), .dina(n307), .dout(n311));
    jxor g062(.dinb(n295), .dina(n311), .dout(n315));
    jand g063(.dinb(n284), .dina(n1446), .dout(n319));
    jnot g064(.din(Gic1), .dout(n322));
    jor g065(.dinb(n322), .dina(n78), .dout(n326));
    jxor g066(.dinb(Gid28), .dina(Gid29), .dout(n330));
    jxor g067(.dinb(Gid30), .dina(Gid31), .dout(n334));
    jxor g068(.dinb(n330), .dina(n334), .dout(n338));
    jxor g069(.dinb(n326), .dina(n338), .dout(n342));
    jxor g070(.dinb(Gid24), .dina(Gid25), .dout(n346));
    jxor g071(.dinb(Gid26), .dina(Gid27), .dout(n350));
    jxor g072(.dinb(n346), .dina(n350), .dout(n354));
    jxor g073(.dinb(Gid1), .dina(Gid5), .dout(n358));
    jxor g074(.dinb(Gid9), .dina(Gid13), .dout(n362));
    jxor g075(.dinb(n358), .dina(n362), .dout(n366));
    jxor g076(.dinb(n354), .dina(n366), .dout(n370));
    jxor g077(.dinb(n342), .dina(n370), .dout(n374));
    jxor g078(.dinb(n130), .dina(n374), .dout(n378));
    jnot g079(.din(Gic3), .dout(n381));
    jor g080(.dinb(n381), .dina(n78), .dout(n385));
    jxor g081(.dinb(n122), .dina(n385), .dout(n389));
    jxor g082(.dinb(Gid3), .dina(Gid7), .dout(n393));
    jxor g083(.dinb(Gid11), .dina(Gid15), .dout(n397));
    jxor g084(.dinb(n393), .dina(n397), .dout(n401));
    jxor g085(.dinb(n338), .dina(n401), .dout(n405));
    jxor g086(.dinb(n389), .dina(n405), .dout(n409));
    jnot g087(.din(Gic2), .dout(n412));
    jor g088(.dinb(n412), .dina(n78), .dout(n416));
    jxor g089(.dinb(n94), .dina(n416), .dout(n420));
    jxor g090(.dinb(Gid2), .dina(Gid6), .dout(n424));
    jxor g091(.dinb(Gid10), .dina(Gid14), .dout(n428));
    jxor g092(.dinb(n424), .dina(n428), .dout(n432));
    jxor g093(.dinb(n354), .dina(n432), .dout(n436));
    jxor g094(.dinb(n420), .dina(n436), .dout(n440));
    jand g095(.dinb(n409), .dina(n440), .dout(n444));
    jand g096(.dinb(n378), .dina(n444), .dout(n448));
    jxor g097(.dinb(n409), .dina(n440), .dout(n452));
    jand g098(.dinb(n130), .dina(n374), .dout(n456));
    jand g099(.dinb(n452), .dina(n456), .dout(n460));
    jor g100(.dinb(n448), .dina(n460), .dout(n464));
    jand g101(.dinb(n1216), .dina(n464), .dout(n468));
    jand g102(.dinb(n1236), .dina(n468), .dout(n472));
    jand g103(.dinb(n1221), .dina(n472), .dout(n476));
    jxor g104(.dinb(n2001), .dina(n476), .dout(God0));
    jnot g105(.din(n374), .dout(n483));
    jand g106(.dinb(n1227), .dina(n472), .dout(n487));
    jxor g107(.dinb(n1671), .dina(n487), .dout(God1));
    jnot g108(.din(n440), .dout(n494));
    jand g109(.dinb(n1233), .dina(n472), .dout(n498));
    jxor g110(.dinb(n1509), .dina(n498), .dout(God2));
    jnot g111(.din(n409), .dout(n505));
    jand g112(.dinb(n1245), .dina(n472), .dout(n509));
    jxor g113(.dinb(n1587), .dina(n509), .dout(God3));
    jnot g114(.din(n188), .dout(n516));
    jand g115(.dinb(n516), .dina(n1473), .dout(n520));
    jand g116(.dinb(n468), .dina(n1248), .dout(n524));
    jand g117(.dinb(n1218), .dina(n524), .dout(n528));
    jxor g118(.dinb(n2466), .dina(n528), .dout(God4));
    jand g119(.dinb(n1224), .dina(n524), .dout(n536));
    jxor g120(.dinb(n2436), .dina(n536), .dout(God5));
    jand g121(.dinb(n1230), .dina(n524), .dout(n544));
    jxor g122(.dinb(n2406), .dina(n544), .dout(God6));
    jand g123(.dinb(n1242), .dina(n524), .dout(n552));
    jxor g124(.dinb(n2376), .dina(n552), .dout(God7));
    jnot g125(.din(n315), .dout(n559));
    jand g126(.dinb(n1419), .dina(n559), .dout(n563));
    jand g127(.dinb(n250), .dina(n563), .dout(n567));
    jand g128(.dinb(n464), .dina(n567), .dout(n571));
    jand g129(.dinb(n1332), .dina(n571), .dout(n575));
    jxor g130(.dinb(n1974), .dina(n575), .dout(n579));
    jand g131(.dinb(n1623), .dina(n571), .dout(n583));
    jxor g132(.dinb(n1644), .dina(n583), .dout(n587));
    jand g133(.dinb(n1377), .dina(n571), .dout(n591));
    jxor g134(.dinb(n1482), .dina(n591), .dout(n595));
    jand g135(.dinb(n1539), .dina(n571), .dout(n599));
    jxor g136(.dinb(n1560), .dina(n599), .dout(n603));
    jand g137(.dinb(n520), .dina(n563), .dout(n607));
    jand g138(.dinb(n464), .dina(n607), .dout(n611));
    jand g139(.dinb(n1341), .dina(n611), .dout(n615));
    jxor g140(.dinb(n2349), .dina(n615), .dout(n619));
    jand g141(.dinb(n1632), .dina(n611), .dout(n623));
    jxor g142(.dinb(n2322), .dina(n623), .dout(n627));
    jand g143(.dinb(n1386), .dina(n611), .dout(n631));
    jxor g144(.dinb(n2295), .dina(n631), .dout(n635));
    jand g145(.dinb(n1548), .dina(n611), .dout(n639));
    jxor g146(.dinb(n2268), .dina(n639), .dout(n643));
    jand g147(.dinb(n133), .dina(n1641), .dout(n647));
    jand g148(.dinb(n1557), .dina(n494), .dout(n651));
    jxor g149(.dinb(n188), .dina(n243), .dout(n655));
    jand g150(.dinb(n281), .dina(n315), .dout(n659));
    jand g151(.dinb(n655), .dina(n659), .dout(n663));
    jxor g152(.dinb(n281), .dina(n315), .dout(n667));
    jand g153(.dinb(n188), .dina(n243), .dout(n671));
    jand g154(.dinb(n667), .dina(n671), .dout(n675));
    jor g155(.dinb(n663), .dina(n675), .dout(n679));
    jand g156(.dinb(n1375), .dina(n679), .dout(n683));
    jand g157(.dinb(n1330), .dina(n683), .dout(n687));
    jand g158(.dinb(n1266), .dina(n687), .dout(n691));
    jxor g159(.dinb(n2091), .dina(n691), .dout(God16));
    jand g160(.dinb(n1290), .dina(n687), .dout(n699));
    jxor g161(.dinb(n2061), .dina(n699), .dout(God17));
    jand g162(.dinb(n1314), .dina(n687), .dout(n707));
    jxor g163(.dinb(n2031), .dina(n707), .dout(God18));
    jand g164(.dinb(n1362), .dina(n687), .dout(n715));
    jxor g165(.dinb(n2238), .dina(n715), .dout(God19));
    jand g166(.dinb(n505), .dina(n1479), .dout(n723));
    jand g167(.dinb(n1477), .dina(n679), .dout(n727));
    jand g168(.dinb(n1330), .dina(n727), .dout(n731));
    jand g169(.dinb(n1254), .dina(n731), .dout(n735));
    jxor g170(.dinb(n1944), .dina(n735), .dout(God20));
    jand g171(.dinb(n1278), .dina(n731), .dout(n743));
    jxor g172(.dinb(n1914), .dina(n743), .dout(God21));
    jand g173(.dinb(n1302), .dina(n731), .dout(n751));
    jxor g174(.dinb(n1884), .dina(n751), .dout(God22));
    jand g175(.dinb(n1350), .dina(n731), .dout(n759));
    jxor g176(.dinb(n2208), .dina(n759), .dout(God23));
    jand g177(.dinb(n1881), .dina(n483), .dout(n767));
    jand g178(.dinb(n1621), .dina(n683), .dout(n771));
    jand g179(.dinb(n1407), .dina(n771), .dout(n775));
    jxor g180(.dinb(n1761), .dina(n775), .dout(God24));
    jand g181(.dinb(n1434), .dina(n771), .dout(n783));
    jxor g182(.dinb(n1731), .dina(n783), .dout(God25));
    jand g183(.dinb(n1461), .dina(n771), .dout(n791));
    jxor g184(.dinb(n1701), .dina(n791), .dout(God26));
    jand g185(.dinb(n2133), .dina(n771), .dout(n799));
    jxor g186(.dinb(n2178), .dina(n799), .dout(God27));
    jand g187(.dinb(n1621), .dina(n727), .dout(n807));
    jand g188(.dinb(n1395), .dina(n807), .dout(n811));
    jxor g189(.dinb(n1851), .dina(n811), .dout(God28));
    jand g190(.dinb(n1422), .dina(n807), .dout(n819));
    jxor g191(.dinb(n1821), .dina(n819), .dout(God29));
    jand g192(.dinb(n1449), .dina(n807), .dout(n827));
    jxor g193(.dinb(n1791), .dina(n827), .dout(God30));
    jand g194(.dinb(n2121), .dina(n807), .dout(n835));
    jxor g195(.dinb(n2148), .dina(n835), .dout(God31));
    jdff dff_A_0gFFnEVW4_2(.din(n643), .dout(God15));
    jdff dff_A_xwjecuNR3_2(.din(n635), .dout(God14));
    jdff dff_A_M993VYio7_2(.din(n627), .dout(God13));
    jdff dff_A_vUu1lEre9_2(.din(n619), .dout(God12));
    jdff dff_A_V82npY4S7_2(.din(n603), .dout(God11));
    jdff dff_A_BQoihez14_2(.din(n595), .dout(God10));
    jdff dff_A_phqVuheg8_2(.din(n587), .dout(God9));
    jdff dff_A_t28eNMZB9_2(.din(n579), .dout(God8));
    jdff dff_A_Q9QU7Bj22_0(.din(Gid4), .dout(n2493));
    jdff dff_A_u5U6dJIk9_0(.din(n2493), .dout(n2490));
    jdff dff_A_uewNRjes4_0(.din(n2490), .dout(n2487));
    jdff dff_A_uphu97sY5_0(.din(n2487), .dout(n2484));
    jdff dff_A_Bop2CZk01_0(.din(n2484), .dout(n2481));
    jdff dff_A_KSR6PYxZ3_0(.din(n2481), .dout(n2478));
    jdff dff_A_KLD5TaUO6_0(.din(n2478), .dout(n2475));
    jdff dff_A_tJ1TKZDb7_0(.din(n2475), .dout(n2472));
    jdff dff_A_rcKQSZOw1_0(.din(n2472), .dout(n2469));
    jdff dff_A_SJVqMlIB8_0(.din(n2469), .dout(n2466));
    jdff dff_A_FEjCAOOB9_0(.din(Gid5), .dout(n2463));
    jdff dff_A_nK0oOtDP6_0(.din(n2463), .dout(n2460));
    jdff dff_A_HM7LaCNQ1_0(.din(n2460), .dout(n2457));
    jdff dff_A_Os6jK8DZ6_0(.din(n2457), .dout(n2454));
    jdff dff_A_nC0QMXJo1_0(.din(n2454), .dout(n2451));
    jdff dff_A_lrYOVdYK3_0(.din(n2451), .dout(n2448));
    jdff dff_A_OJtApgAg7_0(.din(n2448), .dout(n2445));
    jdff dff_A_DAPceiDm1_0(.din(n2445), .dout(n2442));
    jdff dff_A_kJrN7nTn3_0(.din(n2442), .dout(n2439));
    jdff dff_A_UQFIFnTQ2_0(.din(n2439), .dout(n2436));
    jdff dff_A_uUCOQP0F4_0(.din(Gid6), .dout(n2433));
    jdff dff_A_YQ98d7MC7_0(.din(n2433), .dout(n2430));
    jdff dff_A_AWubdkLT4_0(.din(n2430), .dout(n2427));
    jdff dff_A_jNS75QVW0_0(.din(n2427), .dout(n2424));
    jdff dff_A_vP13EDxK5_0(.din(n2424), .dout(n2421));
    jdff dff_A_PoHwq2T92_0(.din(n2421), .dout(n2418));
    jdff dff_A_2RITnD434_0(.din(n2418), .dout(n2415));
    jdff dff_A_3GTPcaUq2_0(.din(n2415), .dout(n2412));
    jdff dff_A_iragpCK20_0(.din(n2412), .dout(n2409));
    jdff dff_A_zQgSfDyE2_0(.din(n2409), .dout(n2406));
    jdff dff_A_lscNnTKl6_0(.din(Gid7), .dout(n2403));
    jdff dff_A_elegr9Tb2_0(.din(n2403), .dout(n2400));
    jdff dff_A_5lMtpV8S1_0(.din(n2400), .dout(n2397));
    jdff dff_A_gi9z9JqQ7_0(.din(n2397), .dout(n2394));
    jdff dff_A_2Xk9XLIf5_0(.din(n2394), .dout(n2391));
    jdff dff_A_aT5wCdID9_0(.din(n2391), .dout(n2388));
    jdff dff_A_2gN5oCr33_0(.din(n2388), .dout(n2385));
    jdff dff_A_8EI5q0Y17_0(.din(n2385), .dout(n2382));
    jdff dff_A_5VyHml628_0(.din(n2382), .dout(n2379));
    jdff dff_A_7ujHyr9o1_0(.din(n2379), .dout(n2376));
    jdff dff_A_lvlshYzq9_0(.din(Gid12), .dout(n2373));
    jdff dff_A_k9L2HXLl0_0(.din(n2373), .dout(n2370));
    jdff dff_A_by4slmXY1_0(.din(n2370), .dout(n2367));
    jdff dff_A_m1sqM9th8_0(.din(n2367), .dout(n2364));
    jdff dff_A_ARGoS4l13_0(.din(n2364), .dout(n2361));
    jdff dff_A_R33jGjHD3_0(.din(n2361), .dout(n2358));
    jdff dff_A_K3Mrkb8M7_0(.din(n2358), .dout(n2355));
    jdff dff_A_qF1NASqO8_0(.din(n2355), .dout(n2352));
    jdff dff_A_bJrZfhqv3_0(.din(n2352), .dout(n2349));
    jdff dff_A_O2UE9IzC2_0(.din(Gid13), .dout(n2346));
    jdff dff_A_rMLrcsmc2_0(.din(n2346), .dout(n2343));
    jdff dff_A_eBfJ4Coj1_0(.din(n2343), .dout(n2340));
    jdff dff_A_ZlkRaivg2_0(.din(n2340), .dout(n2337));
    jdff dff_A_ZcpqnJ6x1_0(.din(n2337), .dout(n2334));
    jdff dff_A_6KtuZ0AG2_0(.din(n2334), .dout(n2331));
    jdff dff_A_mAXp9ONW6_0(.din(n2331), .dout(n2328));
    jdff dff_A_bprUAUkd5_0(.din(n2328), .dout(n2325));
    jdff dff_A_bTGgUHIj7_0(.din(n2325), .dout(n2322));
    jdff dff_A_nDFg7F1w9_0(.din(Gid14), .dout(n2319));
    jdff dff_A_xCy40D9R8_0(.din(n2319), .dout(n2316));
    jdff dff_A_hkZMM9wa3_0(.din(n2316), .dout(n2313));
    jdff dff_A_l1j6JX6B1_0(.din(n2313), .dout(n2310));
    jdff dff_A_jv9Hdcw18_0(.din(n2310), .dout(n2307));
    jdff dff_A_zdHGMoJ11_0(.din(n2307), .dout(n2304));
    jdff dff_A_dShX5IlL8_0(.din(n2304), .dout(n2301));
    jdff dff_A_Z1IMZcrX2_0(.din(n2301), .dout(n2298));
    jdff dff_A_OWcFprd26_0(.din(n2298), .dout(n2295));
    jdff dff_A_fQc3mC2M6_0(.din(Gid15), .dout(n2292));
    jdff dff_A_rnRe6E3z3_0(.din(n2292), .dout(n2289));
    jdff dff_A_d91xuzmG4_0(.din(n2289), .dout(n2286));
    jdff dff_A_KzL5nWyO5_0(.din(n2286), .dout(n2283));
    jdff dff_A_YGiECME14_0(.din(n2283), .dout(n2280));
    jdff dff_A_aIBlnj696_0(.din(n2280), .dout(n2277));
    jdff dff_A_YFxtvHIf0_0(.din(n2277), .dout(n2274));
    jdff dff_A_VcAUAAtf7_0(.din(n2274), .dout(n2271));
    jdff dff_A_CJbwMbIM4_0(.din(n2271), .dout(n2268));
    jdff dff_A_mL8s61KD1_0(.din(Gid19), .dout(n2265));
    jdff dff_A_wSARpwOI5_0(.din(n2265), .dout(n2262));
    jdff dff_A_TrVHqvel7_0(.din(n2262), .dout(n2259));
    jdff dff_A_BtdDMZw22_0(.din(n2259), .dout(n2256));
    jdff dff_A_BVYQKpOY1_0(.din(n2256), .dout(n2253));
    jdff dff_A_7YSPXMZk4_0(.din(n2253), .dout(n2250));
    jdff dff_A_nFSXwWmf8_0(.din(n2250), .dout(n2247));
    jdff dff_A_zMlzXqyE7_0(.din(n2247), .dout(n2244));
    jdff dff_A_7RLeG4eD5_0(.din(n2244), .dout(n2241));
    jdff dff_A_MU4e8yk37_0(.din(n2241), .dout(n2238));
    jdff dff_A_4HhG9E0g4_0(.din(Gid23), .dout(n2235));
    jdff dff_A_9ZY00dve4_0(.din(n2235), .dout(n2232));
    jdff dff_A_5ODI8vRM2_0(.din(n2232), .dout(n2229));
    jdff dff_A_jaRpQjHc8_0(.din(n2229), .dout(n2226));
    jdff dff_A_Ckzt9hw16_0(.din(n2226), .dout(n2223));
    jdff dff_A_LR1VdwX56_0(.din(n2223), .dout(n2220));
    jdff dff_A_EO95xqL32_0(.din(n2220), .dout(n2217));
    jdff dff_A_U0yyqX1C4_0(.din(n2217), .dout(n2214));
    jdff dff_B_Rte4w9es3_1(.din(n319), .dout(n1216));
    jdff dff_A_TdZSoHeu6_1(.din(n1332), .dout(n1218));
    jdff dff_A_6KPLnSfE3_2(.din(n1332), .dout(n1221));
    jdff dff_A_BhLGWC9X5_1(.din(n1623), .dout(n1224));
    jdff dff_A_B8CNvG0r6_2(.din(n1623), .dout(n1227));
    jdff dff_A_2yTkI1hH2_1(.din(n1377), .dout(n1230));
    jdff dff_A_q33zhwJ46_2(.din(n1377), .dout(n1233));
    jdff dff_A_2ABazkR04_1(.din(n1239), .dout(n1236));
    jdff dff_A_kyUciNE67_1(.din(n250), .dout(n1239));
    jdff dff_A_hLWWJtjJ9_1(.din(n1539), .dout(n1242));
    jdff dff_A_3aOtSkKJ2_2(.din(n1539), .dout(n1245));
    jdff dff_A_L1CkNsjZ1_1(.din(n1251), .dout(n1248));
    jdff dff_A_eQ2qaFeR9_1(.din(n520), .dout(n1251));
    jdff dff_A_sWanwmY18_0(.din(n1257), .dout(n1254));
    jdff dff_A_S66pMkgt8_0(.din(n1260), .dout(n1257));
    jdff dff_A_YLTzpJ3V6_0(.din(n1263), .dout(n1260));
    jdff dff_A_Sz4GEjpJ0_0(.din(n284), .dout(n1263));
    jdff dff_A_8oUWoO1h5_1(.din(n1269), .dout(n1266));
    jdff dff_A_Kh4rU1f75_1(.din(n1272), .dout(n1269));
    jdff dff_A_4Z5AXO532_1(.din(n1275), .dout(n1272));
    jdff dff_A_PFwnz67Q2_1(.din(n284), .dout(n1275));
    jdff dff_A_PPTg3Iav1_0(.din(n1281), .dout(n1278));
    jdff dff_A_7nI52sIH1_0(.din(n1284), .dout(n1281));
    jdff dff_A_rEKDNrAq3_0(.din(n1287), .dout(n1284));
    jdff dff_A_AfRShPpe1_0(.din(n559), .dout(n1287));
    jdff dff_A_eXdv9tdl2_1(.din(n1293), .dout(n1290));
    jdff dff_A_OZUH0gIg6_1(.din(n1296), .dout(n1293));
    jdff dff_A_2Ur3Tta55_1(.din(n1299), .dout(n1296));
    jdff dff_A_vi0FvzEj7_1(.din(n559), .dout(n1299));
    jdff dff_A_2uAaj9Bf0_0(.din(n1305), .dout(n1302));
    jdff dff_A_FuPINirv5_0(.din(n1308), .dout(n1305));
    jdff dff_A_PGUN6AGs3_0(.din(n1311), .dout(n1308));
    jdff dff_A_tPqZDPfm0_0(.din(n246), .dout(n1311));
    jdff dff_A_IDpmEh4b7_1(.din(n1317), .dout(n1314));
    jdff dff_A_WbBNiIxZ5_1(.din(n1320), .dout(n1317));
    jdff dff_A_kiW0wYSH5_1(.din(n1323), .dout(n1320));
    jdff dff_A_NS9FZHD09_1(.din(n246), .dout(n1323));
    jdff dff_B_HhewDILa3_2(.din(n647), .dout(n1327));
    jdff dff_B_0Hmst9Ao8_2(.din(n1327), .dout(n1330));
    jdff dff_A_2S3VPVf79_0(.din(n1335), .dout(n1332));
    jdff dff_A_vzCi34q87_0(.din(n1338), .dout(n1335));
    jdff dff_A_SCFHFwce0_0(.din(n133), .dout(n1338));
    jdff dff_A_fJv2Jp3o9_2(.din(n1344), .dout(n1341));
    jdff dff_A_C6xzG2D39_2(.din(n1347), .dout(n1344));
    jdff dff_A_prAwz9Vu2_2(.din(n133), .dout(n1347));
    jdff dff_A_7ixFlQiL8_0(.din(n1353), .dout(n1350));
    jdff dff_A_TwPnBrxg4_0(.din(n1356), .dout(n1353));
    jdff dff_A_TvcsOpbY5_0(.din(n1359), .dout(n1356));
    jdff dff_A_oAlwXBEk4_0(.din(n516), .dout(n1359));
    jdff dff_A_zHEqWZDn5_1(.din(n1365), .dout(n1362));
    jdff dff_A_3KxKLf872_1(.din(n1368), .dout(n1365));
    jdff dff_A_8DdwiIYg1_1(.din(n1371), .dout(n1368));
    jdff dff_A_vaeSNQw06_1(.din(n516), .dout(n1371));
    jdff dff_B_1lRPjpPb7_1(.din(n651), .dout(n1375));
    jdff dff_A_UYfCEhZU1_0(.din(n1380), .dout(n1377));
    jdff dff_A_Phz1k2l22_0(.din(n1383), .dout(n1380));
    jdff dff_A_RncceOAf9_0(.din(n494), .dout(n1383));
    jdff dff_A_P6FlqHA59_2(.din(n1389), .dout(n1386));
    jdff dff_A_dqAQLQcH0_2(.din(n1392), .dout(n1389));
    jdff dff_A_iJLQLhR73_2(.din(n494), .dout(n1392));
    jdff dff_A_epSb9qdl6_1(.din(n1398), .dout(n1395));
    jdff dff_A_jabU7rpU6_1(.din(n1401), .dout(n1398));
    jdff dff_A_LSR4ATTz1_1(.din(n1404), .dout(n1401));
    jdff dff_A_MWQtMVEZ6_1(.din(n284), .dout(n1404));
    jdff dff_A_AnxztkLF9_2(.din(n1410), .dout(n1407));
    jdff dff_A_1KQlsavk1_2(.din(n1413), .dout(n1410));
    jdff dff_A_V4ZTXYvZ3_2(.din(n1416), .dout(n1413));
    jdff dff_A_4o4B2lIS3_2(.din(n284), .dout(n1416));
    jdff dff_A_QtbBYnQl6_0(.din(n281), .dout(n1419));
    jdff dff_A_WWjFi0UX1_1(.din(n1425), .dout(n1422));
    jdff dff_A_IkUIFELm3_1(.din(n1428), .dout(n1425));
    jdff dff_A_7X4Ljqha9_1(.din(n1431), .dout(n1428));
    jdff dff_A_zffwGAEv4_1(.din(n559), .dout(n1431));
    jdff dff_A_KBaPVuYb3_2(.din(n1437), .dout(n1434));
    jdff dff_A_yj58tIyF3_2(.din(n1440), .dout(n1437));
    jdff dff_A_uYaAjGkO5_2(.din(n1443), .dout(n1440));
    jdff dff_A_Kw1437sK5_2(.din(n559), .dout(n1443));
    jdff dff_A_On7HNBGE5_1(.din(n315), .dout(n1446));
    jdff dff_A_CqwAOkyA1_1(.din(n1452), .dout(n1449));
    jdff dff_A_GXT2H5hE7_1(.din(n1455), .dout(n1452));
    jdff dff_A_droRYdtB6_1(.din(n1458), .dout(n1455));
    jdff dff_A_pG7nol8U6_1(.din(n246), .dout(n1458));
    jdff dff_A_OQYjVJfn6_2(.din(n1464), .dout(n1461));
    jdff dff_A_strRyCsJ7_2(.din(n1467), .dout(n1464));
    jdff dff_A_J7PpDoso4_2(.din(n1470), .dout(n1467));
    jdff dff_A_rWLW3Flm8_2(.din(n246), .dout(n1470));
    jdff dff_A_V9M7ah3w9_0(.din(n243), .dout(n1473));
    jdff dff_B_N7ictSn66_1(.din(n723), .dout(n1477));
    jdff dff_A_33RMobVg8_1(.din(n440), .dout(n1479));
    jdff dff_A_BnFN8U9V3_0(.din(n1485), .dout(n1482));
    jdff dff_A_MvTSmV1a7_0(.din(n1488), .dout(n1485));
    jdff dff_A_OGeO50AT2_0(.din(n1491), .dout(n1488));
    jdff dff_A_ekw8U2Yn3_0(.din(n1494), .dout(n1491));
    jdff dff_A_a9qtkZCR4_0(.din(n1497), .dout(n1494));
    jdff dff_A_14TJJhDQ2_0(.din(n1500), .dout(n1497));
    jdff dff_A_JfyyAggR3_0(.din(n1503), .dout(n1500));
    jdff dff_A_0Fj3mhkg6_0(.din(n1506), .dout(n1503));
    jdff dff_A_eNw4OvOL7_0(.din(Gid10), .dout(n1506));
    jdff dff_A_uzu088kf7_0(.din(n1512), .dout(n1509));
    jdff dff_A_1M6HnTol0_0(.din(n1515), .dout(n1512));
    jdff dff_A_KBZjQZSa4_0(.din(n1518), .dout(n1515));
    jdff dff_A_WApYmXMJ0_0(.din(n1521), .dout(n1518));
    jdff dff_A_seQvNnjn2_0(.din(n1524), .dout(n1521));
    jdff dff_A_4ntoCw6p3_0(.din(n1527), .dout(n1524));
    jdff dff_A_M5O6gD222_0(.din(n1530), .dout(n1527));
    jdff dff_A_5lRPa6kP6_0(.din(n1533), .dout(n1530));
    jdff dff_A_o0YPHncf4_0(.din(n1536), .dout(n1533));
    jdff dff_A_OKibUI7s5_0(.din(Gid2), .dout(n1536));
    jdff dff_A_bMlTEZej5_0(.din(n1542), .dout(n1539));
    jdff dff_A_fREsPi3E1_0(.din(n1545), .dout(n1542));
    jdff dff_A_t6RG7Zt14_0(.din(n505), .dout(n1545));
    jdff dff_A_Rjjfo0AW7_2(.din(n1551), .dout(n1548));
    jdff dff_A_GhWMT5938_2(.din(n1554), .dout(n1551));
    jdff dff_A_3XNOMt5T1_2(.din(n505), .dout(n1554));
    jdff dff_A_FO2hXmLY2_1(.din(n409), .dout(n1557));
    jdff dff_A_vPwUlBW37_0(.din(n1563), .dout(n1560));
    jdff dff_A_PhEFyMRB9_0(.din(n1566), .dout(n1563));
    jdff dff_A_OSux50RW4_0(.din(n1569), .dout(n1566));
    jdff dff_A_Y9B8Rzjy0_0(.din(n1572), .dout(n1569));
    jdff dff_A_0uwM0Kvi8_0(.din(n1575), .dout(n1572));
    jdff dff_A_4yXhrOGE4_0(.din(n1578), .dout(n1575));
    jdff dff_A_k6yO1LPW8_0(.din(n1581), .dout(n1578));
    jdff dff_A_zQ70HLrv4_0(.din(n1584), .dout(n1581));
    jdff dff_A_yRsTuwFj2_0(.din(Gid11), .dout(n1584));
    jdff dff_A_Tw6OxXSH2_0(.din(n1590), .dout(n1587));
    jdff dff_A_qXe8D67c3_0(.din(n1593), .dout(n1590));
    jdff dff_A_LxHPl93l3_0(.din(n1596), .dout(n1593));
    jdff dff_A_2BdazliQ7_0(.din(n1599), .dout(n1596));
    jdff dff_A_fUE2og6W6_0(.din(n1602), .dout(n1599));
    jdff dff_A_aaniOkpX3_0(.din(n1605), .dout(n1602));
    jdff dff_A_l7ObL10c7_0(.din(n1608), .dout(n1605));
    jdff dff_A_zSlgRA0O8_0(.din(n1611), .dout(n1608));
    jdff dff_A_7FGY6xaU5_0(.din(n1614), .dout(n1611));
    jdff dff_A_KHUXRvdL7_0(.din(Gid3), .dout(n1614));
    jdff dff_B_mWHhQsvF5_2(.din(n767), .dout(n1618));
    jdff dff_B_9twUOoy62_2(.din(n1618), .dout(n1621));
    jdff dff_A_G2E10bxz6_0(.din(n1626), .dout(n1623));
    jdff dff_A_GC0ibkMC1_0(.din(n1629), .dout(n1626));
    jdff dff_A_VNTPnrGY7_0(.din(n483), .dout(n1629));
    jdff dff_A_sFRoOlTJ8_2(.din(n1635), .dout(n1632));
    jdff dff_A_A391UrqM5_2(.din(n1638), .dout(n1635));
    jdff dff_A_dVt3nXuF0_2(.din(n483), .dout(n1638));
    jdff dff_A_gqixjLQh5_1(.din(n374), .dout(n1641));
    jdff dff_A_SWnw53He3_0(.din(n1647), .dout(n1644));
    jdff dff_A_CKzKrGB18_0(.din(n1650), .dout(n1647));
    jdff dff_A_AF4m5V6n6_0(.din(n1653), .dout(n1650));
    jdff dff_A_wAEQXdj32_0(.din(n1656), .dout(n1653));
    jdff dff_A_UYbbm1rk5_0(.din(n1659), .dout(n1656));
    jdff dff_A_JOiUTZgL4_0(.din(n1662), .dout(n1659));
    jdff dff_A_JhDOKjDH6_0(.din(n1665), .dout(n1662));
    jdff dff_A_4sLZQorV9_0(.din(n1668), .dout(n1665));
    jdff dff_A_5uodxngr2_0(.din(Gid9), .dout(n1668));
    jdff dff_A_aUldtjdY0_0(.din(n1674), .dout(n1671));
    jdff dff_A_wACvA3Qr6_0(.din(n1677), .dout(n1674));
    jdff dff_A_OogJDUR73_0(.din(n1680), .dout(n1677));
    jdff dff_A_pRblt9553_0(.din(n1683), .dout(n1680));
    jdff dff_A_toDSFF3U6_0(.din(n1686), .dout(n1683));
    jdff dff_A_fltqXaHr7_0(.din(n1689), .dout(n1686));
    jdff dff_A_Sl5llNbD9_0(.din(n1692), .dout(n1689));
    jdff dff_A_gAjXG29N7_0(.din(n1695), .dout(n1692));
    jdff dff_A_FwBczpJY7_0(.din(n1698), .dout(n1695));
    jdff dff_A_rzRBRAv01_0(.din(Gid1), .dout(n1698));
    jdff dff_A_IHN72d6R3_0(.din(n1704), .dout(n1701));
    jdff dff_A_UtLEqozy8_0(.din(n1707), .dout(n1704));
    jdff dff_A_MHie7kHn0_0(.din(n1710), .dout(n1707));
    jdff dff_A_0esC6ZKe8_0(.din(n1713), .dout(n1710));
    jdff dff_A_wDEpy8lL1_0(.din(n1716), .dout(n1713));
    jdff dff_A_Mv49l19D9_0(.din(n1719), .dout(n1716));
    jdff dff_A_zhybXctI1_0(.din(n1722), .dout(n1719));
    jdff dff_A_A3wFFSpk3_0(.din(n1725), .dout(n1722));
    jdff dff_A_47y8V22V9_0(.din(n1728), .dout(n1725));
    jdff dff_A_vLWxBEJx6_0(.din(Gid26), .dout(n1728));
    jdff dff_A_ZX4FFNas6_0(.din(n1734), .dout(n1731));
    jdff dff_A_Xfx9u2AJ8_0(.din(n1737), .dout(n1734));
    jdff dff_A_dBR6HYfx1_0(.din(n1740), .dout(n1737));
    jdff dff_A_r4ISNrTa8_0(.din(n1743), .dout(n1740));
    jdff dff_A_OZfdIsGw1_0(.din(n1746), .dout(n1743));
    jdff dff_A_pfjZ9vSC1_0(.din(n1749), .dout(n1746));
    jdff dff_A_0bVKRiT10_0(.din(n1752), .dout(n1749));
    jdff dff_A_rvc0P0ac6_0(.din(n1755), .dout(n1752));
    jdff dff_A_RbcBFmVd1_0(.din(n1758), .dout(n1755));
    jdff dff_A_9G3kIPMC3_0(.din(Gid25), .dout(n1758));
    jdff dff_A_gtE5ETZB7_0(.din(n1764), .dout(n1761));
    jdff dff_A_xLTxHeh53_0(.din(n1767), .dout(n1764));
    jdff dff_A_cWNTN2Kh0_0(.din(n1770), .dout(n1767));
    jdff dff_A_KtzlxNWX8_0(.din(n1773), .dout(n1770));
    jdff dff_A_IuTClk5m8_0(.din(n1776), .dout(n1773));
    jdff dff_A_DPQlQ9WG7_0(.din(n1779), .dout(n1776));
    jdff dff_A_qkpe5N1U3_0(.din(n1782), .dout(n1779));
    jdff dff_A_swttxSx32_0(.din(n1785), .dout(n1782));
    jdff dff_A_mwxQF4Gx8_0(.din(n1788), .dout(n1785));
    jdff dff_A_dd4JPFrE8_0(.din(Gid24), .dout(n1788));
    jdff dff_A_lbGUBpgO1_0(.din(n1794), .dout(n1791));
    jdff dff_A_JPYZM99P2_0(.din(n1797), .dout(n1794));
    jdff dff_A_f51ybZ9u9_0(.din(n1800), .dout(n1797));
    jdff dff_A_7NjTLA9B4_0(.din(n1803), .dout(n1800));
    jdff dff_A_cKPXaQXu4_0(.din(n1806), .dout(n1803));
    jdff dff_A_rjWFOxWc5_0(.din(n1809), .dout(n1806));
    jdff dff_A_cr50fjhn3_0(.din(n1812), .dout(n1809));
    jdff dff_A_JrKgJGNp3_0(.din(n1815), .dout(n1812));
    jdff dff_A_6mmsx3k63_0(.din(n1818), .dout(n1815));
    jdff dff_A_TZpTo5JX4_0(.din(Gid30), .dout(n1818));
    jdff dff_A_JX7wGKoY3_0(.din(n1824), .dout(n1821));
    jdff dff_A_if4ZQIqE3_0(.din(n1827), .dout(n1824));
    jdff dff_A_XOs7FRxQ7_0(.din(n1830), .dout(n1827));
    jdff dff_A_JQV1tsnl5_0(.din(n1833), .dout(n1830));
    jdff dff_A_mevcgLrD1_0(.din(n1836), .dout(n1833));
    jdff dff_A_SYHVpbdf0_0(.din(n1839), .dout(n1836));
    jdff dff_A_qdT5E7x65_0(.din(n1842), .dout(n1839));
    jdff dff_A_pDidJfOR4_0(.din(n1845), .dout(n1842));
    jdff dff_A_da3829Pt9_0(.din(n1848), .dout(n1845));
    jdff dff_A_a5AItAOo8_0(.din(Gid29), .dout(n1848));
    jdff dff_A_txPybEeQ9_0(.din(n1854), .dout(n1851));
    jdff dff_A_V05bALyb7_0(.din(n1857), .dout(n1854));
    jdff dff_A_ctYLBXow0_0(.din(n1860), .dout(n1857));
    jdff dff_A_0A1peUsx9_0(.din(n1863), .dout(n1860));
    jdff dff_A_BpPcuJPU4_0(.din(n1866), .dout(n1863));
    jdff dff_A_qmHKVTtT1_0(.din(n1869), .dout(n1866));
    jdff dff_A_5ygwasus8_0(.din(n1872), .dout(n1869));
    jdff dff_A_L2OxOXah8_0(.din(n1875), .dout(n1872));
    jdff dff_A_bJ6ShmnL5_0(.din(n1878), .dout(n1875));
    jdff dff_A_3oRQdi0j7_0(.din(Gid28), .dout(n1878));
    jdff dff_A_PyVA7EGn1_1(.din(n130), .dout(n1881));
    jdff dff_A_BtacOvqK5_0(.din(n1887), .dout(n1884));
    jdff dff_A_RJNDdF9y6_0(.din(n1890), .dout(n1887));
    jdff dff_A_fCZsKO7I5_0(.din(n1893), .dout(n1890));
    jdff dff_A_TZwdlQaY6_0(.din(n1896), .dout(n1893));
    jdff dff_A_WyjxEtHg9_0(.din(n1899), .dout(n1896));
    jdff dff_A_Vmn004ox3_0(.din(n1902), .dout(n1899));
    jdff dff_A_iGH9wmEz6_0(.din(n1905), .dout(n1902));
    jdff dff_A_yNHQbjuu0_0(.din(n1908), .dout(n1905));
    jdff dff_A_c20KbhyS3_0(.din(n1911), .dout(n1908));
    jdff dff_A_KunSXwVK0_0(.din(Gid22), .dout(n1911));
    jdff dff_A_lRp0t7UF0_0(.din(n1917), .dout(n1914));
    jdff dff_A_9M7aqyj65_0(.din(n1920), .dout(n1917));
    jdff dff_A_u7izM9Cn9_0(.din(n1923), .dout(n1920));
    jdff dff_A_frk0Qvs84_0(.din(n1926), .dout(n1923));
    jdff dff_A_u7TEIbvS7_0(.din(n1929), .dout(n1926));
    jdff dff_A_QvPMK6I32_0(.din(n1932), .dout(n1929));
    jdff dff_A_oEl98jT08_0(.din(n1935), .dout(n1932));
    jdff dff_A_6wx3TpP10_0(.din(n1938), .dout(n1935));
    jdff dff_A_xGDdqj0E7_0(.din(n1941), .dout(n1938));
    jdff dff_A_m2W6bpls3_0(.din(Gid21), .dout(n1941));
    jdff dff_A_Gi5xeoLN4_0(.din(n1947), .dout(n1944));
    jdff dff_A_TcDsCDqx4_0(.din(n1950), .dout(n1947));
    jdff dff_A_Ye7CRd2K2_0(.din(n1953), .dout(n1950));
    jdff dff_A_1LmDgkJP8_0(.din(n1956), .dout(n1953));
    jdff dff_A_G3H5DhMQ3_0(.din(n1959), .dout(n1956));
    jdff dff_A_vBoQbvAa6_0(.din(n1962), .dout(n1959));
    jdff dff_A_oL762PwQ9_0(.din(n1965), .dout(n1962));
    jdff dff_A_vb8dpYgl3_0(.din(n1968), .dout(n1965));
    jdff dff_A_a1BeJlsp6_0(.din(n1971), .dout(n1968));
    jdff dff_A_RyUKfDPN1_0(.din(Gid20), .dout(n1971));
    jdff dff_A_4KVCkl8i3_0(.din(n1977), .dout(n1974));
    jdff dff_A_nNjTufm59_0(.din(n1980), .dout(n1977));
    jdff dff_A_NrRiGeKo1_0(.din(n1983), .dout(n1980));
    jdff dff_A_ESfgqCBv0_0(.din(n1986), .dout(n1983));
    jdff dff_A_SeAbwVxP4_0(.din(n1989), .dout(n1986));
    jdff dff_A_mNR4Y6U18_0(.din(n1992), .dout(n1989));
    jdff dff_A_r0Ywc9aq7_0(.din(n1995), .dout(n1992));
    jdff dff_A_r4ktytZQ2_0(.din(n1998), .dout(n1995));
    jdff dff_A_AwHdmpig7_0(.din(Gid8), .dout(n1998));
    jdff dff_A_YjTEE3Pg0_0(.din(n2004), .dout(n2001));
    jdff dff_A_Cu7Fa5Za4_0(.din(n2007), .dout(n2004));
    jdff dff_A_fRTrJqm21_0(.din(n2010), .dout(n2007));
    jdff dff_A_6KK732pB3_0(.din(n2013), .dout(n2010));
    jdff dff_A_AyOpBqSA7_0(.din(n2016), .dout(n2013));
    jdff dff_A_0W79r3pP0_0(.din(n2019), .dout(n2016));
    jdff dff_A_bOAKxogg4_0(.din(n2022), .dout(n2019));
    jdff dff_A_jQVn1B2T5_0(.din(n2025), .dout(n2022));
    jdff dff_A_q7pJMTOM0_0(.din(n2028), .dout(n2025));
    jdff dff_A_BByNI0iY6_0(.din(Gid0), .dout(n2028));
    jdff dff_A_0o09eJDB8_0(.din(n2034), .dout(n2031));
    jdff dff_A_0k8BNKeL2_0(.din(n2037), .dout(n2034));
    jdff dff_A_lNJKa5Gs4_0(.din(n2040), .dout(n2037));
    jdff dff_A_vYRpx3jL0_0(.din(n2043), .dout(n2040));
    jdff dff_A_dkjIODqH8_0(.din(n2046), .dout(n2043));
    jdff dff_A_F2G7BfAI9_0(.din(n2049), .dout(n2046));
    jdff dff_A_1t5Wy7CZ1_0(.din(n2052), .dout(n2049));
    jdff dff_A_wP4Lbnov4_0(.din(n2055), .dout(n2052));
    jdff dff_A_qxzGUQ6h7_0(.din(n2058), .dout(n2055));
    jdff dff_A_vU1D6bgZ8_0(.din(Gid18), .dout(n2058));
    jdff dff_A_Hno60Ike5_0(.din(n2064), .dout(n2061));
    jdff dff_A_AWW1OFdr3_0(.din(n2067), .dout(n2064));
    jdff dff_A_Ch0EbdFD8_0(.din(n2070), .dout(n2067));
    jdff dff_A_ShDuunpI0_0(.din(n2073), .dout(n2070));
    jdff dff_A_UwjZBQ4v4_0(.din(n2076), .dout(n2073));
    jdff dff_A_QBKEX4JP5_0(.din(n2079), .dout(n2076));
    jdff dff_A_j3tkr4lD9_0(.din(n2082), .dout(n2079));
    jdff dff_A_Z6HM39KG5_0(.din(n2085), .dout(n2082));
    jdff dff_A_dp2cvq6m2_0(.din(n2088), .dout(n2085));
    jdff dff_A_WO8HeG3p8_0(.din(Gid17), .dout(n2088));
    jdff dff_A_sEaoKCku6_0(.din(n2094), .dout(n2091));
    jdff dff_A_66Z97chb2_0(.din(n2097), .dout(n2094));
    jdff dff_A_u3Ir0up57_0(.din(n2100), .dout(n2097));
    jdff dff_A_60mWSzSS8_0(.din(n2103), .dout(n2100));
    jdff dff_A_tRm41EB96_0(.din(n2106), .dout(n2103));
    jdff dff_A_8gw4dbGE5_0(.din(n2109), .dout(n2106));
    jdff dff_A_SLYlGsF47_0(.din(n2112), .dout(n2109));
    jdff dff_A_y9BVyr5U2_0(.din(n2115), .dout(n2112));
    jdff dff_A_uQRHRRbW1_0(.din(n2118), .dout(n2115));
    jdff dff_A_GsS2TZLX3_0(.din(Gid16), .dout(n2118));
    jdff dff_A_deQSb6i25_1(.din(n2124), .dout(n2121));
    jdff dff_A_oPlJmZpD1_1(.din(n2127), .dout(n2124));
    jdff dff_A_yDlRMZoa3_1(.din(n2130), .dout(n2127));
    jdff dff_A_cM2AZTWl7_1(.din(n516), .dout(n2130));
    jdff dff_A_0HSEoaew5_2(.din(n2136), .dout(n2133));
    jdff dff_A_9XG849Aw4_2(.din(n2139), .dout(n2136));
    jdff dff_A_fpj052yc5_2(.din(n2142), .dout(n2139));
    jdff dff_A_ZBKZozHu9_2(.din(n516), .dout(n2142));
    jdff dff_A_kssEyZ2b0_1(.din(n188), .dout(n2145));
    jdff dff_A_wigew52h3_0(.din(n2151), .dout(n2148));
    jdff dff_A_HDCfog407_0(.din(n2154), .dout(n2151));
    jdff dff_A_IjD9XFoy1_0(.din(n2157), .dout(n2154));
    jdff dff_A_g0G3o8nG5_0(.din(n2160), .dout(n2157));
    jdff dff_A_6CEhYrYR9_0(.din(n2163), .dout(n2160));
    jdff dff_A_tzStsJfK8_0(.din(n2166), .dout(n2163));
    jdff dff_A_iYlVlumC2_0(.din(n2169), .dout(n2166));
    jdff dff_A_peXKtfNH3_0(.din(n2172), .dout(n2169));
    jdff dff_A_kn0Hf9RC3_0(.din(n2175), .dout(n2172));
    jdff dff_A_UCk3kjV57_0(.din(Gid31), .dout(n2175));
    jdff dff_A_ypaPnnl45_0(.din(n2181), .dout(n2178));
    jdff dff_A_aK9jkWKe8_0(.din(n2184), .dout(n2181));
    jdff dff_A_i6mdCrtn4_0(.din(n2187), .dout(n2184));
    jdff dff_A_LkNOoy142_0(.din(n2190), .dout(n2187));
    jdff dff_A_dDxVUUBm9_0(.din(n2193), .dout(n2190));
    jdff dff_A_mzjkBW4y7_0(.din(n2196), .dout(n2193));
    jdff dff_A_2uqDLfHW2_0(.din(n2199), .dout(n2196));
    jdff dff_A_xa1uItNd7_0(.din(n2202), .dout(n2199));
    jdff dff_A_sqoJtCka8_0(.din(n2205), .dout(n2202));
    jdff dff_A_WJROMAW18_0(.din(Gid27), .dout(n2205));
    jdff dff_A_5CsYpWLa7_0(.din(n2211), .dout(n2208));
    jdff dff_A_fBQ3eCIP1_0(.din(n2214), .dout(n2211));
endmodule

