// Benchmark "top" written by ABC on Wed May 27 23:37:17 2020

module gf_multiplier ( 
    a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 , a8 ,
    a9 , a10 , a11 , a12 , a13 , a14 , a15 , a16 ,
    a17 , a18 , a19 , a20 , a21 , a22 , a23 , a24 ,
    a25 , a26 , a27 , a28 , a29 , a30 , a31 , a32 ,
    a33 , a34 , a35 , a36 , a37 , a38 , a39 , a40 ,
    a41 , a42 , a43 , a44 , a45 , a46 , a47 , a48 ,
    a49 , a50 , a51 , a52 , a53 , a54 , a55 , a56 ,
    a57 , a58 , a59 , a60 , a61 , a62 , a63 , b0 ,
    b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 , b9 ,
    b10 , b11 , b12 , b13 , b14 , b15 , b16 , b17 ,
    b18 , b19 , b20 , b21 , b22 , b23 , b24 , b25 ,
    b26 , b27 , b28 , b29 , b30 , b31 , b32 , b33 ,
    b34 , b35 , b36 , b37 , b38 , b39 , b40 , b41 ,
    b42 , b43 , b44 , b45 , b46 , b47 , b48 , b49 ,
    b50 , b51 , b52 , b53 , b54 , b55 , b56 , b57 ,
    b58 , b59 , b60 , b61 , b62 , b63 ,
    f0 , f1 , f2 , f3 , f4 , f5 , f6 , f7 , f8 ,
    f9 , f10 , f11 , f12 , f13 , f14 , f15 , f16 ,
    f17 , f18 , f19 , f20 , f21 , f22 , f23 , f24 ,
    f25 , f26 , f27 , f28 , f29 , f30 , f31 , f32 ,
    f33 , f34 , f35 , f36 , f37 , f38 , f39 , f40 ,
    f41 , f42 , f43 , f44 , f45 , f46 , f47 , f48 ,
    f49 , f50 , f51 , f52 , f53 , f54 , f55 , f56 ,
    f57 , f58 , f59 , f60 , f61 , f62 , f63 , f64 ,
    f65 , f66 , f67 , f68 , f69 , f70 , f71 , f72 ,
    f73 , f74 , f75 , f76 , f77 , f78 , f79 , f80 ,
    f81 , f82 , f83 , f84 , f85 , f86 , f87 , f88 ,
    f89 , f90 , f91 , f92 , f93 , f94 , f95 , f96 ,
    f97 , f98 , f99 , f100 , f101 , f102 , f103 ,
    f104 , f105 , f106 , f107 , f108 , f109 , f110 ,
    f111 , f112 , f113 , f114 , f115 , f116 , f117 ,
    f118 , f119 , f120 , f121 , f122 , f123 , f124 ,
    f125 , f126 , f127   );
  input  a0 , a1 , a2 , a3 , a4 , a5 , a6 , a7 ,
    a8 , a9 , a10 , a11 , a12 , a13 , a14 , a15 ,
    a16 , a17 , a18 , a19 , a20 , a21 , a22 , a23 ,
    a24 , a25 , a26 , a27 , a28 , a29 , a30 , a31 ,
    a32 , a33 , a34 , a35 , a36 , a37 , a38 , a39 ,
    a40 , a41 , a42 , a43 , a44 , a45 , a46 , a47 ,
    a48 , a49 , a50 , a51 , a52 , a53 , a54 , a55 ,
    a56 , a57 , a58 , a59 , a60 , a61 , a62 , a63 ,
    b0 , b1 , b2 , b3 , b4 , b5 , b6 , b7 , b8 ,
    b9 , b10 , b11 , b12 , b13 , b14 , b15 , b16 ,
    b17 , b18 , b19 , b20 , b21 , b22 , b23 , b24 ,
    b25 , b26 , b27 , b28 , b29 , b30 , b31 , b32 ,
    b33 , b34 , b35 , b36 , b37 , b38 , b39 , b40 ,
    b41 , b42 , b43 , b44 , b45 , b46 , b47 , b48 ,
    b49 , b50 , b51 , b52 , b53 , b54 , b55 , b56 ,
    b57 , b58 , b59 , b60 , b61 , b62 , b63 ;
  output f0 , f1 , f2 , f3 , f4 , f5 , f6 , f7 ,
    f8 , f9 , f10 , f11 , f12 , f13 , f14 , f15 ,
    f16 , f17 , f18 , f19 , f20 , f21 , f22 , f23 ,
    f24 , f25 , f26 , f27 , f28 , f29 , f30 , f31 ,
    f32 , f33 , f34 , f35 , f36 , f37 , f38 , f39 ,
    f40 , f41 , f42 , f43 , f44 , f45 , f46 , f47 ,
    f48 , f49 , f50 , f51 , f52 , f53 , f54 , f55 ,
    f56 , f57 , f58 , f59 , f60 , f61 , f62 , f63 ,
    f64 , f65 , f66 , f67 , f68 , f69 , f70 , f71 ,
    f72 , f73 , f74 , f75 , f76 , f77 , f78 , f79 ,
    f80 , f81 , f82 , f83 , f84 , f85 , f86 , f87 ,
    f88 , f89 , f90 , f91 , f92 , f93 , f94 , f95 ,
    f96 , f97 , f98 , f99 , f100 , f101 , f102 ,
    f103 , f104 , f105 , f106 , f107 , f108 , f109 ,
    f110 , f111 , f112 , f113 , f114 , f115 , f116 ,
    f117 , f118 , f119 , f120 , f121 , f122 , f123 ,
    f124 , f125 , f126 , f127 ;
  wire n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n348, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
    n380, n381, n382, n383, n384, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n478,
    n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
    n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
    n527, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n782, n783,
    n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
    n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
    n2423, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
    n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
    n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
    n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
    n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
    n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
    n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
    n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
    n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
    n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
    n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
    n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
    n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
    n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
    n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
    n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
    n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
    n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
    n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
    n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
    n4063, n4064, n4065, n4066, n4067, n4068, n4070, n4071, n4072, n4073,
    n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
    n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
    n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
    n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
    n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
    n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
    n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
    n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
    n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
    n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
    n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
    n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
    n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
    n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
    n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
    n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
    n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
    n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
    n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
    n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
    n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
    n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
    n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
    n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
    n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
    n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
    n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
    n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
    n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
    n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
    n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
    n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
    n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
    n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
    n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
    n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
    n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
    n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
    n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
    n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
    n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
    n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
    n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
    n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
    n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
    n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
    n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
    n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
    n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
    n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
    n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
    n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
    n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
    n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
    n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
    n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
    n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
    n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
    n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
    n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
    n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
    n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
    n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
    n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
    n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
    n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
    n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
    n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
    n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
    n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
    n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
    n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
    n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
    n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
    n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
    n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
    n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
    n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
    n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
    n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
    n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
    n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
    n6143, n6144, n6145, n6146, n6147, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
    n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
    n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
    n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
    n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
    n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
    n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
    n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
    n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
    n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
    n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
    n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
    n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
    n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
    n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
    n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
    n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
    n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
    n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
    n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
    n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
    n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
    n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
    n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
    n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
    n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
    n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
    n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
    n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
    n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
    n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
    n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7096, n7097,
    n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
    n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
    n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
    n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
    n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
    n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
    n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
    n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
    n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
    n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
    n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
    n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
    n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
    n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
    n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
    n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
    n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
    n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
    n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
    n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
    n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
    n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
    n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
    n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
    n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
    n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
    n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
    n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
    n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
    n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
    n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
    n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
    n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
    n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
    n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
    n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
    n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
    n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
    n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
    n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
    n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
    n7850, n7851, n7852, n7853, n7854, n7856, n7857, n7858, n7859, n7860,
    n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
    n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
    n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
    n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8121,
    n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
    n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
    n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
    n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
    n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
    n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
    n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
    n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
    n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
    n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
    n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
    n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
    n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
    n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
    n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
    n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
    n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
    n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
    n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
    n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
    n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
    n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
    n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
    n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
    n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
    n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
    n8382, n8383, n8384, n8385, n8386, n8388, n8389, n8390, n8391, n8392,
    n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
    n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
    n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
    n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
    n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
    n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
    n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
    n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
    n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
    n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
    n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
    n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
    n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
    n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
    n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
    n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
    n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
    n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
    n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
    n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
    n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
    n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
    n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
    n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
    n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
    n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
    n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
    n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
    n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
    n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
    n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
    n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
    n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
    n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
    n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
    n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
    n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
    n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
    n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
    n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
    n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
    n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
    n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
    n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
    n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
    n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
    n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
    n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
    n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
    n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
    n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9486,
    n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
    n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
    n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
    n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
    n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
    n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
    n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
    n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
    n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
    n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
    n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
    n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
    n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
    n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
    n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
    n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
    n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
    n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
    n9767, n9768, n9769, n9770, n9771, n9772, n9774, n9775, n9776, n9777,
    n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
    n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
    n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
    n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
    n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
    n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
    n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
    n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
    n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
    n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
    n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
    n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
    n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
    n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
    n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
    n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
    n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
    n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
    n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
    n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
    n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
    n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
    n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
    n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
    n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
    n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
    n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
    n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
    n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
    n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
    n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
    n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
    n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
    n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
    n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
    n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
    n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
    n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
    n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
    n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
    n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
    n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
    n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
    n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
    n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
    n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
    n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
    n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
    n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
    n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
    n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
    n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
    n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
    n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
    n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
    n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
    n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
    n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
    n10530, n10531, n10532, n10534, n10535, n10536, n10537, n10538, n10539,
    n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
    n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
    n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
    n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
    n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
    n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
    n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
    n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
    n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
    n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
    n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
    n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
    n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
    n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
    n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
    n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
    n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
    n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
    n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
    n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
    n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
    n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
    n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
    n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
    n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
    n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
    n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
    n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
    n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
    n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
    n10819, n10820, n10821, n10823, n10824, n10825, n10826, n10827, n10828,
    n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
    n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
    n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
    n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
    n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
    n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
    n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
    n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
    n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
    n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
    n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
    n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
    n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
    n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
    n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
    n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
    n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
    n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
    n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
    n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
    n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
    n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
    n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
    n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
    n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
    n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
    n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
    n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
    n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
    n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
    n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
    n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
    n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
    n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
    n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
    n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
    n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
    n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
    n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
    n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
    n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
    n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
    n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
    n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
    n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
    n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
    n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
    n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
    n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
    n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
    n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
    n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
    n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
    n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
    n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
    n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
    n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
    n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
    n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
    n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
    n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
    n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
    n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
    n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
    n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
    n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
    n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
    n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
    n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
    n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
    n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
    n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
    n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
    n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
    n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
    n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
    n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
    n11650, n11651, n11652, n11654, n11655, n11656, n11657, n11658, n11659,
    n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
    n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
    n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
    n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
    n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
    n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
    n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
    n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
    n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
    n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
    n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
    n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
    n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
    n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
    n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
    n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
    n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
    n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
    n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
    n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
    n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
    n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
    n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
    n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
    n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
    n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188, n12190, n12191, n12192,
    n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
    n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
    n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
    n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
    n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
    n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
    n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
    n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
    n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
    n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
    n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
    n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
    n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
    n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
    n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
    n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
    n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
    n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
    n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
    n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
    n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
    n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
    n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
    n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
    n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
    n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
    n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12454,
    n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
    n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
    n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
    n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
    n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
    n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
    n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
    n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
    n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
    n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
    n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
    n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
    n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
    n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
    n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
    n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
    n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
    n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
    n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
    n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
    n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
    n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
    n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
    n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
    n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
    n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
    n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
    n12707, n12708, n12709, n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
    n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
    n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
    n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
    n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
    n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
    n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
    n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
    n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
    n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
    n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
    n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
    n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
    n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
    n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
    n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
    n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
    n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
    n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
    n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
    n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
    n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
    n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
    n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
    n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
    n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
    n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
    n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
    n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
    n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
    n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
    n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
    n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
    n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13212, n13213,
    n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
    n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
    n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
    n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
    n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
    n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
    n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
    n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
    n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
    n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
    n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
    n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
    n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
    n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
    n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
    n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
    n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
    n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
    n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
    n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
    n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
    n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
    n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
    n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
    n13448, n13449, n13450, n13451, n13453, n13454, n13455, n13456, n13457,
    n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
    n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
    n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
    n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
    n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
    n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
    n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
    n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
    n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
    n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
    n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
    n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
    n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
    n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
    n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
    n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
    n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13691, n13692,
    n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
    n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
    n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
    n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
    n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
    n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
    n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
    n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
    n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
    n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
    n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
    n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
    n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
    n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
    n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
    n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
    n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
    n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
    n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
    n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
    n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
    n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
    n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
    n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
    n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
    n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
    n13927, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
    n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
    n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
    n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
    n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
    n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
    n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
    n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
    n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
    n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
    n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
    n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
    n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
    n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
    n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
    n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
    n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
    n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
    n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
    n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
    n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
    n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
    n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
    n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
    n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
    n14153, n14154, n14155, n14156, n14157, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
    n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
    n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
    n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
    n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
    n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
    n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
    n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
    n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
    n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
    n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
    n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
    n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14384, n14385, n14386, n14387, n14388,
    n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
    n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
    n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
    n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
    n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
    n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
    n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
    n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
    n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
    n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
    n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
    n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
    n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
    n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
    n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
    n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
    n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
    n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
    n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
    n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
    n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
    n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
    n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
    n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
    n14605, n14606, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
    n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
    n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
    n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
    n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
    n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
    n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
    n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
    n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
    n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
    n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
    n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
    n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
    n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
    n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
    n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
    n14822, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
    n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
    n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
    n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
    n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
    n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
    n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
    n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
    n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
    n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
    n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
    n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
    n15030, n15031, n15032, n15033, n15034, n15036, n15037, n15038, n15039,
    n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
    n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
    n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
    n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
    n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
    n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
    n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
    n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
    n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
    n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
    n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
    n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
    n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
    n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
    n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
    n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
    n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
    n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
    n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
    n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
    n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
    n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
    n15238, n15239, n15240, n15241, n15242, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
    n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
    n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
    n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
    n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
    n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
    n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
    n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
    n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
    n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
    n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
    n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
    n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
    n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
    n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
    n15446, n15447, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
    n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
    n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
    n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
    n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
    n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
    n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
    n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
    n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
    n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
    n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
    n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
    n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
    n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
    n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
    n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
    n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
    n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
    n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
    n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
    n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
    n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
    n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
    n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
    n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
    n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
    n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
    n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
    n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
    n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
    n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
    n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
    n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
    n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
    n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
    n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
    n15844, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
    n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
    n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
    n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
    n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
    n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
    n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
    n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
    n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
    n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
    n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
    n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
    n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
    n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
    n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
    n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
    n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
    n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
    n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
    n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
    n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
    n16034, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
    n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
    n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
    n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
    n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
    n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
    n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
    n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
    n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
    n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
    n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16220, n16222, n16223, n16224,
    n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
    n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
    n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
    n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
    n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
    n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
    n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
    n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
    n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
    n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
    n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
    n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
    n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
    n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
    n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
    n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
    n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
    n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
    n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
    n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
    n16405, n16406, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
    n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
    n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
    n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
    n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
    n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
    n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
    n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
    n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
    n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
    n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
    n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
    n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
    n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
    n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
    n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
    n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
    n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
    n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
    n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
    n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
    n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
    n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
    n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
    n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
    n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
    n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
    n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
    n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
    n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
    n16758, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
    n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
    n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
    n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
    n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
    n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
    n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
    n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
    n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
    n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
    n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
    n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
    n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
    n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
    n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
    n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
    n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
    n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
    n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
    n16930, n16931, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
    n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
    n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
    n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
    n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
    n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
    n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
    n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
    n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
    n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
    n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
    n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
    n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
    n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
    n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
    n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
    n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
    n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
    n17093, n17094, n17095, n17096, n17097, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
    n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
    n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
    n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
    n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
    n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
    n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
    n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
    n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
    n17256, n17257, n17258, n17259, n17261, n17262, n17263, n17264, n17265,
    n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
    n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
    n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
    n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
    n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
    n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
    n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
    n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
    n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
    n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
    n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
    n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
    n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
    n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
    n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
    n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
    n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
    n17419, n17420, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
    n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
    n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
    n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
    n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
    n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
    n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
    n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
    n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
    n17573, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
    n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
    n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
    n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
    n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
    n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
    n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
    n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
    n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
    n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
    n17718, n17719, n17720, n17721, n17722, n17724, n17725, n17726, n17727,
    n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
    n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
    n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
    n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
    n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
    n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
    n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
    n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
    n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
    n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
    n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
    n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
    n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
    n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
    n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
    n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17872,
    n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
    n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
    n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
    n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
    n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
    n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
    n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
    n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
    n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
    n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
    n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
    n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
    n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
    n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
    n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
    n18008, n18009, n18010, n18012, n18013, n18014, n18015, n18016, n18017,
    n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
    n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
    n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
    n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
    n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
    n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
    n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
    n18144, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
    n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
    n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
    n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
    n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
    n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
    n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
    n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
    n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
    n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
    n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
    n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
    n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
    n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
    n18271, n18272, n18273, n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
    n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
    n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
    n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
    n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
    n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
    n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
    n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
    n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
    n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
    n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
    n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
    n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
    n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
    n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
    n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
    n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
    n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
    n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
    n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
    n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
    n18516, n18517, n18518, n18519, n18520, n18522, n18523, n18524, n18525,
    n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
    n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
    n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
    n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
    n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
    n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
    n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
    n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
    n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
    n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
    n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
    n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
    n18634, n18635, n18636, n18638, n18639, n18640, n18641, n18642, n18643,
    n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
    n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
    n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
    n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
    n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
    n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
    n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18751, n18752,
    n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
    n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
    n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
    n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
    n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
    n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
    n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
    n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
    n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
    n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
    n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
    n18852, n18853, n18854, n18855, n18856, n18857, n18859, n18860, n18861,
    n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
    n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
    n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
    n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
    n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
    n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
    n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
    n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
    n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
    n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
    n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
    n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
    n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
    n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
    n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
    n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
    n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
    n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
    n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
    n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
    n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
    n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
    n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
    n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
    n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
    n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
    n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
    n19152, n19153, n19154, n19155, n19157, n19158, n19159, n19160, n19161,
    n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
    n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
    n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
    n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
    n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
    n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
    n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
    n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
    n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
    n19243, n19244, n19245, n19247, n19248, n19249, n19250, n19251, n19252,
    n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
    n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
    n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
    n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
    n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
    n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
    n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
    n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
    n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
    n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
    n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
    n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
    n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
    n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
    n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
    n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
    n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
    n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
    n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
    n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
    n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
    n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
    n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
    n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
    n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
    n19489, n19490, n19491, n19492, n19494, n19495, n19496, n19497, n19498,
    n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
    n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
    n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
    n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
    n19562, n19563, n19564, n19565, n19566, n19568, n19569, n19570, n19571,
    n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
    n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
    n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
    n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
    n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
    n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
    n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
    n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
    n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
    n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
    n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
    n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
    n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
    n19699, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
    n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
    n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
    n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
    n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
    n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
    n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19763,
    n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
    n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
    n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
    n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
    n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
    n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
    n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
    n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
    n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
    n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
    n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
    n19864, n19865, n19866, n19867, n19868, n19870, n19871, n19872, n19873,
    n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
    n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
    n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
    n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
    n19910, n19911, n19912, n19913, n19914, n19916, n19917, n19918, n19919,
    n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928,
    n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
    n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
    n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
    n19956, n19957, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
    n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
    n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
    n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992,
    n19993, n19994, n19995, n19996, n19998, n19999, n20000, n20001, n20002,
    n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
    n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
    n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20034, n20035, n20036, n20037, n20038, n20039,
    n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048,
    n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
    n20058, n20059, n20060, n20061, n20062, n20064, n20065, n20066, n20067,
    n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
    n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
    n20086, n20087, n20088, n20090, n20091, n20092, n20093, n20094, n20095,
    n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104,
    n20105, n20106, n20107, n20108, n20109, n20110, n20112, n20113, n20114,
    n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
    n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
    n20133, n20135, n20136, n20137, n20138, n20139, n20140, n20141;
  jand g00000(.dina(b0 ), .dinb(a0 ), .dout(f0 ));
  jxor g00001(.dina(a2 ), .dinb(a1 ), .dout(n257));
  jand g00002(.dina(n257), .dinb(a0 ), .dout(n258));
  jxor g00003(.dina(b1 ), .dinb(b0 ), .dout(n259));
  jand g00004(.dina(n259), .dinb(n258), .dout(n260));
  jnot g00005(.din(a0 ), .dout(n261));
  jand g00006(.dina(a1 ), .dinb(n261), .dout(n262));
  jand g00007(.dina(n262), .dinb(b0 ), .dout(n263));
  jor  g00008(.dina(n257), .dinb(n261), .dout(n264));
  jnot g00009(.din(n264), .dout(n265));
  jand g00010(.dina(n265), .dinb(b1 ), .dout(n266));
  jor  g00011(.dina(n266), .dinb(n263), .dout(n267));
  jor  g00012(.dina(n267), .dinb(n260), .dout(n268));
  jand g00013(.dina(f0 ), .dinb(a2 ), .dout(n269));
  jxor g00014(.dina(n269), .dinb(n268), .dout(f1 ));
  jnot g00015(.din(b0 ), .dout(n271));
  jand g00016(.dina(b1 ), .dinb(n271), .dout(n272));
  jxor g00017(.dina(n272), .dinb(b2 ), .dout(n273));
  jand g00018(.dina(n273), .dinb(n258), .dout(n274));
  jand g00019(.dina(n262), .dinb(b1 ), .dout(n275));
  jor  g00020(.dina(n275), .dinb(n274), .dout(n276));
  jand g00021(.dina(n265), .dinb(b2 ), .dout(n277));
  jnot g00022(.din(a2 ), .dout(n278));
  jor  g00023(.dina(n278), .dinb(a1 ), .dout(n279));
  jor  g00024(.dina(n279), .dinb(a0 ), .dout(n280));
  jnot g00025(.din(n280), .dout(n281));
  jand g00026(.dina(n281), .dinb(b0 ), .dout(n282));
  jor  g00027(.dina(n282), .dinb(n277), .dout(n283));
  jor  g00028(.dina(n283), .dinb(n276), .dout(n284));
  jor  g00029(.dina(f0 ), .dinb(n278), .dout(n285));
  jor  g00030(.dina(n285), .dinb(n268), .dout(n286));
  jand g00031(.dina(n286), .dinb(a2 ), .dout(n287));
  jxor g00032(.dina(n287), .dinb(n284), .dout(f2 ));
  jor  g00033(.dina(n286), .dinb(n284), .dout(n289));
  jxor g00034(.dina(a3 ), .dinb(a2 ), .dout(n290));
  jand g00035(.dina(n290), .dinb(b0 ), .dout(n291));
  jnot g00036(.din(n291), .dout(n292));
  jnot g00037(.din(b2 ), .dout(n293));
  jnot g00038(.din(n262), .dout(n294));
  jor  g00039(.dina(n294), .dinb(n293), .dout(n295));
  jnot g00040(.din(n258), .dout(n296));
  jxor g00041(.dina(b3 ), .dinb(b2 ), .dout(n297));
  jnot g00042(.din(n297), .dout(n298));
  jor  g00043(.dina(b2 ), .dinb(b0 ), .dout(n299));
  jand g00044(.dina(n299), .dinb(b1 ), .dout(n300));
  jxor g00045(.dina(n300), .dinb(n298), .dout(n301));
  jor  g00046(.dina(n301), .dinb(n296), .dout(n302));
  jnot g00047(.din(b3 ), .dout(n303));
  jor  g00048(.dina(n264), .dinb(n303), .dout(n304));
  jnot g00049(.din(b1 ), .dout(n305));
  jor  g00050(.dina(n280), .dinb(n305), .dout(n306));
  jand g00051(.dina(n306), .dinb(n304), .dout(n307));
  jand g00052(.dina(n307), .dinb(n302), .dout(n308));
  jand g00053(.dina(n308), .dinb(n295), .dout(n309));
  jxor g00054(.dina(n309), .dinb(n278), .dout(n310));
  jxor g00055(.dina(n310), .dinb(n292), .dout(n311));
  jxor g00056(.dina(n311), .dinb(n289), .dout(f3 ));
  jxor g00057(.dina(n309), .dinb(a2 ), .dout(n313));
  jor  g00058(.dina(n313), .dinb(n292), .dout(n314));
  jor  g00059(.dina(n311), .dinb(n289), .dout(n315));
  jand g00060(.dina(n315), .dinb(n314), .dout(n316));
  jxor g00061(.dina(a5 ), .dinb(a4 ), .dout(n317));
  jnot g00062(.din(n317), .dout(n318));
  jand g00063(.dina(n318), .dinb(n290), .dout(n319));
  jand g00064(.dina(n319), .dinb(b1 ), .dout(n320));
  jand g00065(.dina(n317), .dinb(n290), .dout(n321));
  jand g00066(.dina(n321), .dinb(n259), .dout(n322));
  jnot g00067(.din(n290), .dout(n323));
  jxor g00068(.dina(a4 ), .dinb(a3 ), .dout(n324));
  jand g00069(.dina(n324), .dinb(n323), .dout(n325));
  jand g00070(.dina(n325), .dinb(b0 ), .dout(n326));
  jor  g00071(.dina(n326), .dinb(n322), .dout(n327));
  jor  g00072(.dina(n327), .dinb(n320), .dout(n328));
  jnot g00073(.din(n328), .dout(n329));
  jand g00074(.dina(n291), .dinb(a5 ), .dout(n330));
  jxor g00075(.dina(n330), .dinb(n329), .dout(n331));
  jand g00076(.dina(b3 ), .dinb(b2 ), .dout(n332));
  jand g00077(.dina(n300), .dinb(n297), .dout(n333));
  jor  g00078(.dina(n333), .dinb(n332), .dout(n334));
  jxor g00079(.dina(b4 ), .dinb(b3 ), .dout(n335));
  jnot g00080(.din(n335), .dout(n336));
  jxor g00081(.dina(n336), .dinb(n334), .dout(n337));
  jor  g00082(.dina(n337), .dinb(n296), .dout(n338));
  jor  g00083(.dina(n294), .dinb(n303), .dout(n339));
  jnot g00084(.din(b4 ), .dout(n340));
  jor  g00085(.dina(n264), .dinb(n340), .dout(n341));
  jand g00086(.dina(n341), .dinb(n339), .dout(n342));
  jor  g00087(.dina(n280), .dinb(n293), .dout(n343));
  jand g00088(.dina(n343), .dinb(n342), .dout(n344));
  jand g00089(.dina(n344), .dinb(n338), .dout(n345));
  jxor g00090(.dina(n345), .dinb(a2 ), .dout(n346));
  jxor g00091(.dina(n346), .dinb(n331), .dout(n347));
  jnot g00092(.din(n347), .dout(n348));
  jxor g00093(.dina(n348), .dinb(n316), .dout(f4 ));
  jor  g00094(.dina(n346), .dinb(n331), .dout(n350));
  jor  g00095(.dina(n348), .dinb(n316), .dout(n351));
  jand g00096(.dina(n351), .dinb(n350), .dout(n352));
  jor  g00097(.dina(n324), .dinb(n290), .dout(n353));
  jor  g00098(.dina(n353), .dinb(n318), .dout(n354));
  jor  g00099(.dina(n354), .dinb(n271), .dout(n355));
  jand g00100(.dina(n319), .dinb(b2 ), .dout(n356));
  jnot g00101(.din(n356), .dout(n357));
  jand g00102(.dina(n357), .dinb(n355), .dout(n358));
  jand g00103(.dina(n321), .dinb(n273), .dout(n359));
  jand g00104(.dina(n325), .dinb(b1 ), .dout(n360));
  jor  g00105(.dina(n360), .dinb(n359), .dout(n361));
  jnot g00106(.din(n361), .dout(n362));
  jand g00107(.dina(n362), .dinb(n358), .dout(n363));
  jnot g00108(.din(a5 ), .dout(n364));
  jand g00109(.dina(n292), .dinb(a5 ), .dout(n365));
  jand g00110(.dina(n365), .dinb(n329), .dout(n366));
  jor  g00111(.dina(n366), .dinb(n364), .dout(n367));
  jxor g00112(.dina(n367), .dinb(n363), .dout(n368));
  jand g00113(.dina(b4 ), .dinb(b3 ), .dout(n369));
  jand g00114(.dina(n335), .dinb(n334), .dout(n370));
  jor  g00115(.dina(n370), .dinb(n369), .dout(n371));
  jxor g00116(.dina(b5 ), .dinb(b4 ), .dout(n372));
  jnot g00117(.din(n372), .dout(n373));
  jxor g00118(.dina(n373), .dinb(n371), .dout(n374));
  jor  g00119(.dina(n374), .dinb(n296), .dout(n375));
  jor  g00120(.dina(n294), .dinb(n340), .dout(n376));
  jnot g00121(.din(b5 ), .dout(n377));
  jor  g00122(.dina(n264), .dinb(n377), .dout(n378));
  jand g00123(.dina(n378), .dinb(n376), .dout(n379));
  jor  g00124(.dina(n280), .dinb(n303), .dout(n380));
  jand g00125(.dina(n380), .dinb(n379), .dout(n381));
  jand g00126(.dina(n381), .dinb(n375), .dout(n382));
  jxor g00127(.dina(n382), .dinb(a2 ), .dout(n383));
  jxor g00128(.dina(n383), .dinb(n368), .dout(n384));
  jxor g00129(.dina(n384), .dinb(n352), .dout(f5 ));
  jnot g00130(.din(n368), .dout(n386));
  jor  g00131(.dina(n383), .dinb(n386), .dout(n387));
  jor  g00132(.dina(n384), .dinb(n352), .dout(n388));
  jand g00133(.dina(n388), .dinb(n387), .dout(n389));
  jand g00134(.dina(n366), .dinb(n363), .dout(n390));
  jxor g00135(.dina(a6 ), .dinb(a5 ), .dout(n391));
  jand g00136(.dina(n391), .dinb(b0 ), .dout(n392));
  jxor g00137(.dina(n392), .dinb(n390), .dout(n393));
  jnot g00138(.din(n325), .dout(n394));
  jor  g00139(.dina(n394), .dinb(n293), .dout(n395));
  jor  g00140(.dina(n354), .dinb(n305), .dout(n396));
  jnot g00141(.din(n321), .dout(n397));
  jor  g00142(.dina(n397), .dinb(n301), .dout(n398));
  jnot g00143(.din(n319), .dout(n399));
  jor  g00144(.dina(n399), .dinb(n303), .dout(n400));
  jand g00145(.dina(n400), .dinb(n398), .dout(n401));
  jand g00146(.dina(n401), .dinb(n396), .dout(n402));
  jand g00147(.dina(n402), .dinb(n395), .dout(n403));
  jxor g00148(.dina(n403), .dinb(n364), .dout(n404));
  jxor g00149(.dina(n404), .dinb(n393), .dout(n405));
  jnot g00150(.din(n405), .dout(n406));
  jand g00151(.dina(b5 ), .dinb(b4 ), .dout(n407));
  jand g00152(.dina(n372), .dinb(n371), .dout(n408));
  jor  g00153(.dina(n408), .dinb(n407), .dout(n409));
  jxor g00154(.dina(b6 ), .dinb(b5 ), .dout(n410));
  jnot g00155(.din(n410), .dout(n411));
  jxor g00156(.dina(n411), .dinb(n409), .dout(n412));
  jor  g00157(.dina(n412), .dinb(n296), .dout(n413));
  jor  g00158(.dina(n280), .dinb(n340), .dout(n414));
  jnot g00159(.din(b6 ), .dout(n415));
  jor  g00160(.dina(n264), .dinb(n415), .dout(n416));
  jand g00161(.dina(n416), .dinb(n414), .dout(n417));
  jor  g00162(.dina(n294), .dinb(n377), .dout(n418));
  jand g00163(.dina(n418), .dinb(n417), .dout(n419));
  jand g00164(.dina(n419), .dinb(n413), .dout(n420));
  jxor g00165(.dina(n420), .dinb(a2 ), .dout(n421));
  jxor g00166(.dina(n421), .dinb(n406), .dout(n422));
  jnot g00167(.din(n422), .dout(n423));
  jxor g00168(.dina(n423), .dinb(n389), .dout(f6 ));
  jor  g00169(.dina(n421), .dinb(n406), .dout(n425));
  jor  g00170(.dina(n423), .dinb(n389), .dout(n426));
  jand g00171(.dina(n426), .dinb(n425), .dout(n427));
  jand g00172(.dina(n392), .dinb(n390), .dout(n428));
  jnot g00173(.din(n428), .dout(n429));
  jnot g00174(.din(n393), .dout(n430));
  jnot g00175(.din(n404), .dout(n431));
  jor  g00176(.dina(n431), .dinb(n430), .dout(n432));
  jand g00177(.dina(n432), .dinb(n429), .dout(n433));
  jxor g00178(.dina(a8 ), .dinb(a7 ), .dout(n434));
  jand g00179(.dina(n434), .dinb(n391), .dout(n435));
  jand g00180(.dina(n435), .dinb(n259), .dout(n436));
  jnot g00181(.din(n391), .dout(n437));
  jxor g00182(.dina(a7 ), .dinb(a6 ), .dout(n438));
  jand g00183(.dina(n438), .dinb(n437), .dout(n439));
  jand g00184(.dina(n439), .dinb(b0 ), .dout(n440));
  jnot g00185(.din(n434), .dout(n441));
  jand g00186(.dina(n441), .dinb(n391), .dout(n442));
  jand g00187(.dina(n442), .dinb(b1 ), .dout(n443));
  jor  g00188(.dina(n443), .dinb(n440), .dout(n444));
  jor  g00189(.dina(n444), .dinb(n436), .dout(n445));
  jnot g00190(.din(a8 ), .dout(n446));
  jnot g00191(.din(n392), .dout(n447));
  jor  g00192(.dina(n447), .dinb(n446), .dout(n448));
  jxor g00193(.dina(n448), .dinb(n445), .dout(n449));
  jor  g00194(.dina(n337), .dinb(n397), .dout(n450));
  jor  g00195(.dina(n399), .dinb(n340), .dout(n451));
  jor  g00196(.dina(n354), .dinb(n293), .dout(n452));
  jand g00197(.dina(n452), .dinb(n451), .dout(n453));
  jor  g00198(.dina(n394), .dinb(n303), .dout(n454));
  jand g00199(.dina(n454), .dinb(n453), .dout(n455));
  jand g00200(.dina(n455), .dinb(n450), .dout(n456));
  jxor g00201(.dina(n456), .dinb(a5 ), .dout(n457));
  jxor g00202(.dina(n457), .dinb(n449), .dout(n458));
  jnot g00203(.din(n458), .dout(n459));
  jxor g00204(.dina(n459), .dinb(n433), .dout(n460));
  jand g00205(.dina(b6 ), .dinb(b5 ), .dout(n461));
  jand g00206(.dina(n410), .dinb(n409), .dout(n462));
  jor  g00207(.dina(n462), .dinb(n461), .dout(n463));
  jxor g00208(.dina(b7 ), .dinb(b6 ), .dout(n464));
  jnot g00209(.din(n464), .dout(n465));
  jxor g00210(.dina(n465), .dinb(n463), .dout(n466));
  jor  g00211(.dina(n466), .dinb(n296), .dout(n467));
  jor  g00212(.dina(n294), .dinb(n415), .dout(n468));
  jnot g00213(.din(b7 ), .dout(n469));
  jor  g00214(.dina(n264), .dinb(n469), .dout(n470));
  jand g00215(.dina(n470), .dinb(n468), .dout(n471));
  jor  g00216(.dina(n280), .dinb(n377), .dout(n472));
  jand g00217(.dina(n472), .dinb(n471), .dout(n473));
  jand g00218(.dina(n473), .dinb(n467), .dout(n474));
  jxor g00219(.dina(n474), .dinb(a2 ), .dout(n475));
  jxor g00220(.dina(n475), .dinb(n460), .dout(n476));
  jxor g00221(.dina(n476), .dinb(n427), .dout(f7 ));
  jnot g00222(.din(n460), .dout(n478));
  jor  g00223(.dina(n475), .dinb(n478), .dout(n479));
  jor  g00224(.dina(n476), .dinb(n427), .dout(n480));
  jand g00225(.dina(n480), .dinb(n479), .dout(n481));
  jor  g00226(.dina(n457), .dinb(n449), .dout(n482));
  jor  g00227(.dina(n459), .dinb(n433), .dout(n483));
  jand g00228(.dina(n483), .dinb(n482), .dout(n484));
  jor  g00229(.dina(n438), .dinb(n391), .dout(n485));
  jor  g00230(.dina(n485), .dinb(n441), .dout(n486));
  jnot g00231(.din(n486), .dout(n487));
  jand g00232(.dina(n487), .dinb(b0 ), .dout(n488));
  jand g00233(.dina(n439), .dinb(b1 ), .dout(n489));
  jor  g00234(.dina(n489), .dinb(n488), .dout(n490));
  jand g00235(.dina(n435), .dinb(n273), .dout(n491));
  jand g00236(.dina(n442), .dinb(b2 ), .dout(n492));
  jor  g00237(.dina(n492), .dinb(n491), .dout(n493));
  jor  g00238(.dina(n493), .dinb(n490), .dout(n494));
  jnot g00239(.din(n445), .dout(n495));
  jand g00240(.dina(n447), .dinb(a8 ), .dout(n496));
  jand g00241(.dina(n496), .dinb(n495), .dout(n497));
  jnot g00242(.din(n497), .dout(n498));
  jand g00243(.dina(n498), .dinb(a8 ), .dout(n499));
  jxor g00244(.dina(n499), .dinb(n494), .dout(n500));
  jor  g00245(.dina(n374), .dinb(n397), .dout(n501));
  jor  g00246(.dina(n399), .dinb(n377), .dout(n502));
  jor  g00247(.dina(n354), .dinb(n303), .dout(n503));
  jand g00248(.dina(n503), .dinb(n502), .dout(n504));
  jor  g00249(.dina(n394), .dinb(n340), .dout(n505));
  jand g00250(.dina(n505), .dinb(n504), .dout(n506));
  jand g00251(.dina(n506), .dinb(n501), .dout(n507));
  jxor g00252(.dina(n507), .dinb(a5 ), .dout(n508));
  jxor g00253(.dina(n508), .dinb(n500), .dout(n509));
  jnot g00254(.din(n509), .dout(n510));
  jxor g00255(.dina(n510), .dinb(n484), .dout(n511));
  jand g00256(.dina(b7 ), .dinb(b6 ), .dout(n512));
  jand g00257(.dina(n464), .dinb(n463), .dout(n513));
  jor  g00258(.dina(n513), .dinb(n512), .dout(n514));
  jxor g00259(.dina(b8 ), .dinb(b7 ), .dout(n515));
  jnot g00260(.din(n515), .dout(n516));
  jxor g00261(.dina(n516), .dinb(n514), .dout(n517));
  jor  g00262(.dina(n517), .dinb(n296), .dout(n518));
  jnot g00263(.din(b8 ), .dout(n519));
  jor  g00264(.dina(n264), .dinb(n519), .dout(n520));
  jor  g00265(.dina(n294), .dinb(n469), .dout(n521));
  jor  g00266(.dina(n280), .dinb(n415), .dout(n522));
  jand g00267(.dina(n522), .dinb(n521), .dout(n523));
  jand g00268(.dina(n523), .dinb(n520), .dout(n524));
  jand g00269(.dina(n524), .dinb(n518), .dout(n525));
  jxor g00270(.dina(n525), .dinb(n278), .dout(n526));
  jxor g00271(.dina(n526), .dinb(n511), .dout(n527));
  jxor g00272(.dina(n527), .dinb(n481), .dout(f8 ));
  jnot g00273(.din(n526), .dout(n529));
  jor  g00274(.dina(n529), .dinb(n511), .dout(n530));
  jor  g00275(.dina(n527), .dinb(n481), .dout(n531));
  jand g00276(.dina(n531), .dinb(n530), .dout(n532));
  jnot g00277(.din(n500), .dout(n533));
  jor  g00278(.dina(n508), .dinb(n533), .dout(n534));
  jor  g00279(.dina(n509), .dinb(n484), .dout(n535));
  jand g00280(.dina(n535), .dinb(n534), .dout(n536));
  jor  g00281(.dina(n498), .dinb(n494), .dout(n537));
  jxor g00282(.dina(a9 ), .dinb(a8 ), .dout(n538));
  jand g00283(.dina(n538), .dinb(b0 ), .dout(n539));
  jnot g00284(.din(n539), .dout(n540));
  jxor g00285(.dina(n540), .dinb(n537), .dout(n541));
  jnot g00286(.din(n442), .dout(n542));
  jor  g00287(.dina(n542), .dinb(n303), .dout(n543));
  jnot g00288(.din(n435), .dout(n544));
  jor  g00289(.dina(n544), .dinb(n301), .dout(n545));
  jor  g00290(.dina(n486), .dinb(n305), .dout(n546));
  jnot g00291(.din(n439), .dout(n547));
  jor  g00292(.dina(n547), .dinb(n293), .dout(n548));
  jand g00293(.dina(n548), .dinb(n546), .dout(n549));
  jand g00294(.dina(n549), .dinb(n545), .dout(n550));
  jand g00295(.dina(n550), .dinb(n543), .dout(n551));
  jxor g00296(.dina(n551), .dinb(n446), .dout(n552));
  jxor g00297(.dina(n552), .dinb(n541), .dout(n553));
  jnot g00298(.din(n553), .dout(n554));
  jor  g00299(.dina(n412), .dinb(n397), .dout(n555));
  jor  g00300(.dina(n394), .dinb(n377), .dout(n556));
  jor  g00301(.dina(n354), .dinb(n340), .dout(n557));
  jand g00302(.dina(n557), .dinb(n556), .dout(n558));
  jor  g00303(.dina(n399), .dinb(n415), .dout(n559));
  jand g00304(.dina(n559), .dinb(n558), .dout(n560));
  jand g00305(.dina(n560), .dinb(n555), .dout(n561));
  jxor g00306(.dina(n561), .dinb(a5 ), .dout(n562));
  jxor g00307(.dina(n562), .dinb(n554), .dout(n563));
  jxor g00308(.dina(n563), .dinb(n536), .dout(n564));
  jand g00309(.dina(b8 ), .dinb(b7 ), .dout(n565));
  jand g00310(.dina(n515), .dinb(n514), .dout(n566));
  jor  g00311(.dina(n566), .dinb(n565), .dout(n567));
  jxor g00312(.dina(b9 ), .dinb(b8 ), .dout(n568));
  jnot g00313(.din(n568), .dout(n569));
  jxor g00314(.dina(n569), .dinb(n567), .dout(n570));
  jor  g00315(.dina(n570), .dinb(n296), .dout(n571));
  jnot g00316(.din(b9 ), .dout(n572));
  jor  g00317(.dina(n264), .dinb(n572), .dout(n573));
  jor  g00318(.dina(n294), .dinb(n519), .dout(n574));
  jor  g00319(.dina(n280), .dinb(n469), .dout(n575));
  jand g00320(.dina(n575), .dinb(n574), .dout(n576));
  jand g00321(.dina(n576), .dinb(n573), .dout(n577));
  jand g00322(.dina(n577), .dinb(n571), .dout(n578));
  jxor g00323(.dina(n578), .dinb(n278), .dout(n579));
  jxor g00324(.dina(n579), .dinb(n564), .dout(n580));
  jxor g00325(.dina(n580), .dinb(n532), .dout(f9 ));
  jnot g00326(.din(n579), .dout(n582));
  jor  g00327(.dina(n582), .dinb(n564), .dout(n583));
  jor  g00328(.dina(n580), .dinb(n532), .dout(n584));
  jand g00329(.dina(n584), .dinb(n583), .dout(n585));
  jor  g00330(.dina(n562), .dinb(n554), .dout(n586));
  jnot g00331(.din(n563), .dout(n587));
  jor  g00332(.dina(n587), .dinb(n536), .dout(n588));
  jand g00333(.dina(n588), .dinb(n586), .dout(n589));
  jnot g00334(.din(n537), .dout(n590));
  jand g00335(.dina(n539), .dinb(n590), .dout(n591));
  jand g00336(.dina(n552), .dinb(n541), .dout(n592));
  jor  g00337(.dina(n592), .dinb(n591), .dout(n593));
  jxor g00338(.dina(a11 ), .dinb(a10 ), .dout(n594));
  jand g00339(.dina(n594), .dinb(n538), .dout(n595));
  jand g00340(.dina(n595), .dinb(n259), .dout(n596));
  jnot g00341(.din(n538), .dout(n597));
  jxor g00342(.dina(a10 ), .dinb(a9 ), .dout(n598));
  jand g00343(.dina(n598), .dinb(n597), .dout(n599));
  jand g00344(.dina(n599), .dinb(b0 ), .dout(n600));
  jnot g00345(.din(n594), .dout(n601));
  jand g00346(.dina(n601), .dinb(n538), .dout(n602));
  jand g00347(.dina(n602), .dinb(b1 ), .dout(n603));
  jor  g00348(.dina(n603), .dinb(n600), .dout(n604));
  jor  g00349(.dina(n604), .dinb(n596), .dout(n605));
  jnot g00350(.din(a11 ), .dout(n606));
  jor  g00351(.dina(n540), .dinb(n606), .dout(n607));
  jxor g00352(.dina(n607), .dinb(n605), .dout(n608));
  jor  g00353(.dina(n544), .dinb(n337), .dout(n609));
  jor  g00354(.dina(n547), .dinb(n303), .dout(n610));
  jor  g00355(.dina(n486), .dinb(n293), .dout(n611));
  jand g00356(.dina(n611), .dinb(n610), .dout(n612));
  jor  g00357(.dina(n542), .dinb(n340), .dout(n613));
  jand g00358(.dina(n613), .dinb(n612), .dout(n614));
  jand g00359(.dina(n614), .dinb(n609), .dout(n615));
  jxor g00360(.dina(n615), .dinb(a8 ), .dout(n616));
  jxor g00361(.dina(n616), .dinb(n608), .dout(n617));
  jxor g00362(.dina(n617), .dinb(n593), .dout(n618));
  jnot g00363(.din(n618), .dout(n619));
  jor  g00364(.dina(n466), .dinb(n397), .dout(n620));
  jor  g00365(.dina(n394), .dinb(n415), .dout(n621));
  jor  g00366(.dina(n354), .dinb(n377), .dout(n622));
  jand g00367(.dina(n622), .dinb(n621), .dout(n623));
  jor  g00368(.dina(n399), .dinb(n469), .dout(n624));
  jand g00369(.dina(n624), .dinb(n623), .dout(n625));
  jand g00370(.dina(n625), .dinb(n620), .dout(n626));
  jxor g00371(.dina(n626), .dinb(a5 ), .dout(n627));
  jxor g00372(.dina(n627), .dinb(n619), .dout(n628));
  jxor g00373(.dina(n628), .dinb(n589), .dout(n629));
  jand g00374(.dina(b9 ), .dinb(b8 ), .dout(n630));
  jand g00375(.dina(n568), .dinb(n567), .dout(n631));
  jor  g00376(.dina(n631), .dinb(n630), .dout(n632));
  jxor g00377(.dina(b10 ), .dinb(b9 ), .dout(n633));
  jnot g00378(.din(n633), .dout(n634));
  jxor g00379(.dina(n634), .dinb(n632), .dout(n635));
  jor  g00380(.dina(n635), .dinb(n296), .dout(n636));
  jnot g00381(.din(b10 ), .dout(n637));
  jor  g00382(.dina(n264), .dinb(n637), .dout(n638));
  jor  g00383(.dina(n280), .dinb(n519), .dout(n639));
  jor  g00384(.dina(n294), .dinb(n572), .dout(n640));
  jand g00385(.dina(n640), .dinb(n639), .dout(n641));
  jand g00386(.dina(n641), .dinb(n638), .dout(n642));
  jand g00387(.dina(n642), .dinb(n636), .dout(n643));
  jxor g00388(.dina(n643), .dinb(n278), .dout(n644));
  jxor g00389(.dina(n644), .dinb(n629), .dout(n645));
  jxor g00390(.dina(n645), .dinb(n585), .dout(f10 ));
  jnot g00391(.din(n644), .dout(n647));
  jor  g00392(.dina(n647), .dinb(n629), .dout(n648));
  jor  g00393(.dina(n645), .dinb(n585), .dout(n649));
  jand g00394(.dina(n649), .dinb(n648), .dout(n650));
  jor  g00395(.dina(n627), .dinb(n619), .dout(n651));
  jnot g00396(.din(n628), .dout(n652));
  jor  g00397(.dina(n652), .dinb(n589), .dout(n653));
  jand g00398(.dina(n653), .dinb(n651), .dout(n654));
  jor  g00399(.dina(n616), .dinb(n608), .dout(n655));
  jand g00400(.dina(n617), .dinb(n593), .dout(n656));
  jnot g00401(.din(n656), .dout(n657));
  jand g00402(.dina(n657), .dinb(n655), .dout(n658));
  jor  g00403(.dina(n598), .dinb(n538), .dout(n659));
  jor  g00404(.dina(n659), .dinb(n601), .dout(n660));
  jnot g00405(.din(n660), .dout(n661));
  jand g00406(.dina(n661), .dinb(b0 ), .dout(n662));
  jand g00407(.dina(n602), .dinb(b2 ), .dout(n663));
  jor  g00408(.dina(n663), .dinb(n662), .dout(n664));
  jand g00409(.dina(n595), .dinb(n273), .dout(n665));
  jand g00410(.dina(n599), .dinb(b1 ), .dout(n666));
  jor  g00411(.dina(n666), .dinb(n665), .dout(n667));
  jor  g00412(.dina(n667), .dinb(n664), .dout(n668));
  jnot g00413(.din(n605), .dout(n669));
  jand g00414(.dina(n540), .dinb(a11 ), .dout(n670));
  jand g00415(.dina(n670), .dinb(n669), .dout(n671));
  jnot g00416(.din(n671), .dout(n672));
  jand g00417(.dina(n672), .dinb(a11 ), .dout(n673));
  jxor g00418(.dina(n673), .dinb(n668), .dout(n674));
  jnot g00419(.din(n674), .dout(n675));
  jor  g00420(.dina(n544), .dinb(n374), .dout(n676));
  jor  g00421(.dina(n547), .dinb(n340), .dout(n677));
  jor  g00422(.dina(n486), .dinb(n303), .dout(n678));
  jand g00423(.dina(n678), .dinb(n677), .dout(n679));
  jor  g00424(.dina(n542), .dinb(n377), .dout(n680));
  jand g00425(.dina(n680), .dinb(n679), .dout(n681));
  jand g00426(.dina(n681), .dinb(n676), .dout(n682));
  jxor g00427(.dina(n682), .dinb(a8 ), .dout(n683));
  jxor g00428(.dina(n683), .dinb(n675), .dout(n684));
  jnot g00429(.din(n684), .dout(n685));
  jxor g00430(.dina(n685), .dinb(n658), .dout(n686));
  jor  g00431(.dina(n517), .dinb(n397), .dout(n687));
  jor  g00432(.dina(n394), .dinb(n469), .dout(n688));
  jor  g00433(.dina(n399), .dinb(n519), .dout(n689));
  jor  g00434(.dina(n354), .dinb(n415), .dout(n690));
  jand g00435(.dina(n690), .dinb(n689), .dout(n691));
  jand g00436(.dina(n691), .dinb(n688), .dout(n692));
  jand g00437(.dina(n692), .dinb(n687), .dout(n693));
  jxor g00438(.dina(n693), .dinb(n364), .dout(n694));
  jxor g00439(.dina(n694), .dinb(n686), .dout(n695));
  jxor g00440(.dina(n695), .dinb(n654), .dout(n696));
  jand g00441(.dina(b10 ), .dinb(b9 ), .dout(n697));
  jand g00442(.dina(n633), .dinb(n632), .dout(n698));
  jor  g00443(.dina(n698), .dinb(n697), .dout(n699));
  jxor g00444(.dina(b11 ), .dinb(b10 ), .dout(n700));
  jnot g00445(.din(n700), .dout(n701));
  jxor g00446(.dina(n701), .dinb(n699), .dout(n702));
  jor  g00447(.dina(n702), .dinb(n296), .dout(n703));
  jnot g00448(.din(b11 ), .dout(n704));
  jor  g00449(.dina(n264), .dinb(n704), .dout(n705));
  jor  g00450(.dina(n294), .dinb(n637), .dout(n706));
  jor  g00451(.dina(n280), .dinb(n572), .dout(n707));
  jand g00452(.dina(n707), .dinb(n706), .dout(n708));
  jand g00453(.dina(n708), .dinb(n705), .dout(n709));
  jand g00454(.dina(n709), .dinb(n703), .dout(n710));
  jxor g00455(.dina(n710), .dinb(n278), .dout(n711));
  jxor g00456(.dina(n711), .dinb(n696), .dout(n712));
  jxor g00457(.dina(n712), .dinb(n650), .dout(f11 ));
  jnot g00458(.din(n711), .dout(n714));
  jor  g00459(.dina(n714), .dinb(n696), .dout(n715));
  jor  g00460(.dina(n712), .dinb(n650), .dout(n716));
  jand g00461(.dina(n716), .dinb(n715), .dout(n717));
  jor  g00462(.dina(n683), .dinb(n675), .dout(n718));
  jor  g00463(.dina(n685), .dinb(n658), .dout(n719));
  jand g00464(.dina(n719), .dinb(n718), .dout(n720));
  jor  g00465(.dina(n672), .dinb(n668), .dout(n721));
  jxor g00466(.dina(a12 ), .dinb(a11 ), .dout(n722));
  jand g00467(.dina(n722), .dinb(b0 ), .dout(n723));
  jnot g00468(.din(n723), .dout(n724));
  jxor g00469(.dina(n724), .dinb(n721), .dout(n725));
  jnot g00470(.din(n602), .dout(n726));
  jor  g00471(.dina(n726), .dinb(n303), .dout(n727));
  jnot g00472(.din(n595), .dout(n728));
  jor  g00473(.dina(n728), .dinb(n301), .dout(n729));
  jor  g00474(.dina(n660), .dinb(n305), .dout(n730));
  jnot g00475(.din(n599), .dout(n731));
  jor  g00476(.dina(n731), .dinb(n293), .dout(n732));
  jand g00477(.dina(n732), .dinb(n730), .dout(n733));
  jand g00478(.dina(n733), .dinb(n729), .dout(n734));
  jand g00479(.dina(n734), .dinb(n727), .dout(n735));
  jxor g00480(.dina(n735), .dinb(n606), .dout(n736));
  jxor g00481(.dina(n736), .dinb(n725), .dout(n737));
  jnot g00482(.din(n737), .dout(n738));
  jor  g00483(.dina(n544), .dinb(n412), .dout(n739));
  jor  g00484(.dina(n542), .dinb(n415), .dout(n740));
  jor  g00485(.dina(n486), .dinb(n340), .dout(n741));
  jand g00486(.dina(n741), .dinb(n740), .dout(n742));
  jor  g00487(.dina(n547), .dinb(n377), .dout(n743));
  jand g00488(.dina(n743), .dinb(n742), .dout(n744));
  jand g00489(.dina(n744), .dinb(n739), .dout(n745));
  jxor g00490(.dina(n745), .dinb(a8 ), .dout(n746));
  jxor g00491(.dina(n746), .dinb(n738), .dout(n747));
  jnot g00492(.din(n747), .dout(n748));
  jxor g00493(.dina(n748), .dinb(n720), .dout(n749));
  jor  g00494(.dina(n570), .dinb(n397), .dout(n750));
  jor  g00495(.dina(n354), .dinb(n469), .dout(n751));
  jor  g00496(.dina(n399), .dinb(n572), .dout(n752));
  jor  g00497(.dina(n394), .dinb(n519), .dout(n753));
  jand g00498(.dina(n753), .dinb(n752), .dout(n754));
  jand g00499(.dina(n754), .dinb(n751), .dout(n755));
  jand g00500(.dina(n755), .dinb(n750), .dout(n756));
  jxor g00501(.dina(n756), .dinb(n364), .dout(n757));
  jxor g00502(.dina(n757), .dinb(n749), .dout(n758));
  jand g00503(.dina(n694), .dinb(n686), .dout(n759));
  jnot g00504(.din(n759), .dout(n760));
  jnot g00505(.din(n695), .dout(n761));
  jor  g00506(.dina(n761), .dinb(n654), .dout(n762));
  jand g00507(.dina(n762), .dinb(n760), .dout(n763));
  jxor g00508(.dina(n763), .dinb(n758), .dout(n764));
  jand g00509(.dina(b11 ), .dinb(b10 ), .dout(n765));
  jand g00510(.dina(n700), .dinb(n699), .dout(n766));
  jor  g00511(.dina(n766), .dinb(n765), .dout(n767));
  jxor g00512(.dina(b12 ), .dinb(b11 ), .dout(n768));
  jnot g00513(.din(n768), .dout(n769));
  jxor g00514(.dina(n769), .dinb(n767), .dout(n770));
  jor  g00515(.dina(n770), .dinb(n296), .dout(n771));
  jnot g00516(.din(b12 ), .dout(n772));
  jor  g00517(.dina(n264), .dinb(n772), .dout(n773));
  jor  g00518(.dina(n294), .dinb(n704), .dout(n774));
  jor  g00519(.dina(n280), .dinb(n637), .dout(n775));
  jand g00520(.dina(n775), .dinb(n774), .dout(n776));
  jand g00521(.dina(n776), .dinb(n773), .dout(n777));
  jand g00522(.dina(n777), .dinb(n771), .dout(n778));
  jxor g00523(.dina(n778), .dinb(n278), .dout(n779));
  jxor g00524(.dina(n779), .dinb(n764), .dout(n780));
  jxor g00525(.dina(n780), .dinb(n717), .dout(f12 ));
  jnot g00526(.din(n779), .dout(n782));
  jor  g00527(.dina(n782), .dinb(n764), .dout(n783));
  jor  g00528(.dina(n780), .dinb(n717), .dout(n784));
  jand g00529(.dina(n784), .dinb(n783), .dout(n785));
  jand g00530(.dina(n757), .dinb(n749), .dout(n786));
  jnot g00531(.din(n786), .dout(n787));
  jnot g00532(.din(n758), .dout(n788));
  jor  g00533(.dina(n763), .dinb(n788), .dout(n789));
  jand g00534(.dina(n789), .dinb(n787), .dout(n790));
  jor  g00535(.dina(n746), .dinb(n738), .dout(n791));
  jor  g00536(.dina(n748), .dinb(n720), .dout(n792));
  jand g00537(.dina(n792), .dinb(n791), .dout(n793));
  jnot g00538(.din(n721), .dout(n794));
  jand g00539(.dina(n723), .dinb(n794), .dout(n795));
  jand g00540(.dina(n736), .dinb(n725), .dout(n796));
  jor  g00541(.dina(n796), .dinb(n795), .dout(n797));
  jxor g00542(.dina(a14 ), .dinb(a13 ), .dout(n798));
  jnot g00543(.din(n798), .dout(n799));
  jand g00544(.dina(n799), .dinb(n722), .dout(n800));
  jand g00545(.dina(n800), .dinb(b1 ), .dout(n801));
  jand g00546(.dina(n798), .dinb(n722), .dout(n802));
  jand g00547(.dina(n802), .dinb(n259), .dout(n803));
  jnot g00548(.din(n722), .dout(n804));
  jxor g00549(.dina(a13 ), .dinb(a12 ), .dout(n805));
  jand g00550(.dina(n805), .dinb(n804), .dout(n806));
  jand g00551(.dina(n806), .dinb(b0 ), .dout(n807));
  jor  g00552(.dina(n807), .dinb(n803), .dout(n808));
  jor  g00553(.dina(n808), .dinb(n801), .dout(n809));
  jnot g00554(.din(a14 ), .dout(n810));
  jor  g00555(.dina(n724), .dinb(n810), .dout(n811));
  jxor g00556(.dina(n811), .dinb(n809), .dout(n812));
  jor  g00557(.dina(n728), .dinb(n337), .dout(n813));
  jor  g00558(.dina(n731), .dinb(n303), .dout(n814));
  jor  g00559(.dina(n660), .dinb(n293), .dout(n815));
  jand g00560(.dina(n815), .dinb(n814), .dout(n816));
  jor  g00561(.dina(n726), .dinb(n340), .dout(n817));
  jand g00562(.dina(n817), .dinb(n816), .dout(n818));
  jand g00563(.dina(n818), .dinb(n813), .dout(n819));
  jxor g00564(.dina(n819), .dinb(a11 ), .dout(n820));
  jxor g00565(.dina(n820), .dinb(n812), .dout(n821));
  jxor g00566(.dina(n821), .dinb(n797), .dout(n822));
  jnot g00567(.din(n822), .dout(n823));
  jor  g00568(.dina(n466), .dinb(n544), .dout(n824));
  jor  g00569(.dina(n547), .dinb(n415), .dout(n825));
  jor  g00570(.dina(n486), .dinb(n377), .dout(n826));
  jand g00571(.dina(n826), .dinb(n825), .dout(n827));
  jor  g00572(.dina(n542), .dinb(n469), .dout(n828));
  jand g00573(.dina(n828), .dinb(n827), .dout(n829));
  jand g00574(.dina(n829), .dinb(n824), .dout(n830));
  jxor g00575(.dina(n830), .dinb(a8 ), .dout(n831));
  jxor g00576(.dina(n831), .dinb(n823), .dout(n832));
  jnot g00577(.din(n832), .dout(n833));
  jxor g00578(.dina(n833), .dinb(n793), .dout(n834));
  jor  g00579(.dina(n635), .dinb(n397), .dout(n835));
  jor  g00580(.dina(n354), .dinb(n519), .dout(n836));
  jor  g00581(.dina(n394), .dinb(n572), .dout(n837));
  jor  g00582(.dina(n399), .dinb(n637), .dout(n838));
  jand g00583(.dina(n838), .dinb(n837), .dout(n839));
  jand g00584(.dina(n839), .dinb(n836), .dout(n840));
  jand g00585(.dina(n840), .dinb(n835), .dout(n841));
  jxor g00586(.dina(n841), .dinb(n364), .dout(n842));
  jxor g00587(.dina(n842), .dinb(n834), .dout(n843));
  jxor g00588(.dina(n843), .dinb(n790), .dout(n844));
  jand g00589(.dina(b12 ), .dinb(b11 ), .dout(n845));
  jand g00590(.dina(n768), .dinb(n767), .dout(n846));
  jor  g00591(.dina(n846), .dinb(n845), .dout(n847));
  jxor g00592(.dina(b13 ), .dinb(b12 ), .dout(n848));
  jnot g00593(.din(n848), .dout(n849));
  jxor g00594(.dina(n849), .dinb(n847), .dout(n850));
  jor  g00595(.dina(n850), .dinb(n296), .dout(n851));
  jnot g00596(.din(b13 ), .dout(n852));
  jor  g00597(.dina(n264), .dinb(n852), .dout(n853));
  jor  g00598(.dina(n294), .dinb(n772), .dout(n854));
  jor  g00599(.dina(n280), .dinb(n704), .dout(n855));
  jand g00600(.dina(n855), .dinb(n854), .dout(n856));
  jand g00601(.dina(n856), .dinb(n853), .dout(n857));
  jand g00602(.dina(n857), .dinb(n851), .dout(n858));
  jxor g00603(.dina(n858), .dinb(n278), .dout(n859));
  jxor g00604(.dina(n859), .dinb(n844), .dout(n860));
  jxor g00605(.dina(n860), .dinb(n785), .dout(f13 ));
  jnot g00606(.din(n859), .dout(n862));
  jor  g00607(.dina(n862), .dinb(n844), .dout(n863));
  jor  g00608(.dina(n860), .dinb(n785), .dout(n864));
  jand g00609(.dina(n864), .dinb(n863), .dout(n865));
  jand g00610(.dina(n842), .dinb(n834), .dout(n866));
  jnot g00611(.din(n866), .dout(n867));
  jnot g00612(.din(n843), .dout(n868));
  jor  g00613(.dina(n868), .dinb(n790), .dout(n869));
  jand g00614(.dina(n869), .dinb(n867), .dout(n870));
  jor  g00615(.dina(n831), .dinb(n823), .dout(n871));
  jor  g00616(.dina(n833), .dinb(n793), .dout(n872));
  jand g00617(.dina(n872), .dinb(n871), .dout(n873));
  jor  g00618(.dina(n820), .dinb(n812), .dout(n874));
  jand g00619(.dina(n821), .dinb(n797), .dout(n875));
  jnot g00620(.din(n875), .dout(n876));
  jand g00621(.dina(n876), .dinb(n874), .dout(n877));
  jnot g00622(.din(n877), .dout(n878));
  jor  g00623(.dina(n805), .dinb(n722), .dout(n879));
  jor  g00624(.dina(n879), .dinb(n799), .dout(n880));
  jnot g00625(.din(n880), .dout(n881));
  jand g00626(.dina(n881), .dinb(b0 ), .dout(n882));
  jand g00627(.dina(n800), .dinb(b2 ), .dout(n883));
  jor  g00628(.dina(n883), .dinb(n882), .dout(n884));
  jand g00629(.dina(n802), .dinb(n273), .dout(n885));
  jand g00630(.dina(n806), .dinb(b1 ), .dout(n886));
  jor  g00631(.dina(n886), .dinb(n885), .dout(n887));
  jor  g00632(.dina(n887), .dinb(n884), .dout(n888));
  jnot g00633(.din(n809), .dout(n889));
  jand g00634(.dina(n724), .dinb(a14 ), .dout(n890));
  jand g00635(.dina(n890), .dinb(n889), .dout(n891));
  jnot g00636(.din(n891), .dout(n892));
  jand g00637(.dina(n892), .dinb(a14 ), .dout(n893));
  jxor g00638(.dina(n893), .dinb(n888), .dout(n894));
  jnot g00639(.din(n894), .dout(n895));
  jor  g00640(.dina(n728), .dinb(n374), .dout(n896));
  jor  g00641(.dina(n726), .dinb(n377), .dout(n897));
  jor  g00642(.dina(n660), .dinb(n303), .dout(n898));
  jand g00643(.dina(n898), .dinb(n897), .dout(n899));
  jor  g00644(.dina(n731), .dinb(n340), .dout(n900));
  jand g00645(.dina(n900), .dinb(n899), .dout(n901));
  jand g00646(.dina(n901), .dinb(n896), .dout(n902));
  jxor g00647(.dina(n902), .dinb(a11 ), .dout(n903));
  jxor g00648(.dina(n903), .dinb(n895), .dout(n904));
  jxor g00649(.dina(n904), .dinb(n878), .dout(n905));
  jor  g00650(.dina(n517), .dinb(n544), .dout(n906));
  jor  g00651(.dina(n542), .dinb(n519), .dout(n907));
  jor  g00652(.dina(n547), .dinb(n469), .dout(n908));
  jor  g00653(.dina(n486), .dinb(n415), .dout(n909));
  jand g00654(.dina(n909), .dinb(n908), .dout(n910));
  jand g00655(.dina(n910), .dinb(n907), .dout(n911));
  jand g00656(.dina(n911), .dinb(n906), .dout(n912));
  jxor g00657(.dina(n912), .dinb(n446), .dout(n913));
  jxor g00658(.dina(n913), .dinb(n905), .dout(n914));
  jnot g00659(.din(n914), .dout(n915));
  jxor g00660(.dina(n915), .dinb(n873), .dout(n916));
  jor  g00661(.dina(n702), .dinb(n397), .dout(n917));
  jor  g00662(.dina(n354), .dinb(n572), .dout(n918));
  jor  g00663(.dina(n399), .dinb(n704), .dout(n919));
  jor  g00664(.dina(n394), .dinb(n637), .dout(n920));
  jand g00665(.dina(n920), .dinb(n919), .dout(n921));
  jand g00666(.dina(n921), .dinb(n918), .dout(n922));
  jand g00667(.dina(n922), .dinb(n917), .dout(n923));
  jxor g00668(.dina(n923), .dinb(n364), .dout(n924));
  jxor g00669(.dina(n924), .dinb(n916), .dout(n925));
  jxor g00670(.dina(n925), .dinb(n870), .dout(n926));
  jand g00671(.dina(b13 ), .dinb(b12 ), .dout(n927));
  jand g00672(.dina(n848), .dinb(n847), .dout(n928));
  jor  g00673(.dina(n928), .dinb(n927), .dout(n929));
  jxor g00674(.dina(b14 ), .dinb(b13 ), .dout(n930));
  jnot g00675(.din(n930), .dout(n931));
  jxor g00676(.dina(n931), .dinb(n929), .dout(n932));
  jor  g00677(.dina(n932), .dinb(n296), .dout(n933));
  jnot g00678(.din(b14 ), .dout(n934));
  jor  g00679(.dina(n264), .dinb(n934), .dout(n935));
  jor  g00680(.dina(n294), .dinb(n852), .dout(n936));
  jor  g00681(.dina(n280), .dinb(n772), .dout(n937));
  jand g00682(.dina(n937), .dinb(n936), .dout(n938));
  jand g00683(.dina(n938), .dinb(n935), .dout(n939));
  jand g00684(.dina(n939), .dinb(n933), .dout(n940));
  jxor g00685(.dina(n940), .dinb(n278), .dout(n941));
  jxor g00686(.dina(n941), .dinb(n926), .dout(n942));
  jxor g00687(.dina(n942), .dinb(n865), .dout(f14 ));
  jnot g00688(.din(n941), .dout(n944));
  jor  g00689(.dina(n944), .dinb(n926), .dout(n945));
  jor  g00690(.dina(n942), .dinb(n865), .dout(n946));
  jand g00691(.dina(n946), .dinb(n945), .dout(n947));
  jand g00692(.dina(n924), .dinb(n916), .dout(n948));
  jnot g00693(.din(n948), .dout(n949));
  jnot g00694(.din(n925), .dout(n950));
  jor  g00695(.dina(n950), .dinb(n870), .dout(n951));
  jand g00696(.dina(n951), .dinb(n949), .dout(n952));
  jand g00697(.dina(n913), .dinb(n905), .dout(n953));
  jnot g00698(.din(n953), .dout(n954));
  jor  g00699(.dina(n915), .dinb(n873), .dout(n955));
  jand g00700(.dina(n955), .dinb(n954), .dout(n956));
  jor  g00701(.dina(n903), .dinb(n895), .dout(n957));
  jand g00702(.dina(n904), .dinb(n878), .dout(n958));
  jnot g00703(.din(n958), .dout(n959));
  jand g00704(.dina(n959), .dinb(n957), .dout(n960));
  jnot g00705(.din(n960), .dout(n961));
  jor  g00706(.dina(n892), .dinb(n888), .dout(n962));
  jxor g00707(.dina(a15 ), .dinb(a14 ), .dout(n963));
  jand g00708(.dina(n963), .dinb(b0 ), .dout(n964));
  jnot g00709(.din(n964), .dout(n965));
  jxor g00710(.dina(n965), .dinb(n962), .dout(n966));
  jnot g00711(.din(n806), .dout(n967));
  jor  g00712(.dina(n967), .dinb(n293), .dout(n968));
  jor  g00713(.dina(n880), .dinb(n305), .dout(n969));
  jnot g00714(.din(n802), .dout(n970));
  jor  g00715(.dina(n970), .dinb(n301), .dout(n971));
  jnot g00716(.din(n800), .dout(n972));
  jor  g00717(.dina(n972), .dinb(n303), .dout(n973));
  jand g00718(.dina(n973), .dinb(n971), .dout(n974));
  jand g00719(.dina(n974), .dinb(n969), .dout(n975));
  jand g00720(.dina(n975), .dinb(n968), .dout(n976));
  jxor g00721(.dina(n976), .dinb(n810), .dout(n977));
  jxor g00722(.dina(n977), .dinb(n966), .dout(n978));
  jnot g00723(.din(n978), .dout(n979));
  jor  g00724(.dina(n728), .dinb(n412), .dout(n980));
  jor  g00725(.dina(n726), .dinb(n415), .dout(n981));
  jor  g00726(.dina(n660), .dinb(n340), .dout(n982));
  jand g00727(.dina(n982), .dinb(n981), .dout(n983));
  jor  g00728(.dina(n731), .dinb(n377), .dout(n984));
  jand g00729(.dina(n984), .dinb(n983), .dout(n985));
  jand g00730(.dina(n985), .dinb(n980), .dout(n986));
  jxor g00731(.dina(n986), .dinb(a11 ), .dout(n987));
  jxor g00732(.dina(n987), .dinb(n979), .dout(n988));
  jxor g00733(.dina(n988), .dinb(n961), .dout(n989));
  jor  g00734(.dina(n570), .dinb(n544), .dout(n990));
  jor  g00735(.dina(n486), .dinb(n469), .dout(n991));
  jor  g00736(.dina(n542), .dinb(n572), .dout(n992));
  jor  g00737(.dina(n547), .dinb(n519), .dout(n993));
  jand g00738(.dina(n993), .dinb(n992), .dout(n994));
  jand g00739(.dina(n994), .dinb(n991), .dout(n995));
  jand g00740(.dina(n995), .dinb(n990), .dout(n996));
  jxor g00741(.dina(n996), .dinb(n446), .dout(n997));
  jxor g00742(.dina(n997), .dinb(n989), .dout(n998));
  jnot g00743(.din(n998), .dout(n999));
  jxor g00744(.dina(n999), .dinb(n956), .dout(n1000));
  jor  g00745(.dina(n770), .dinb(n397), .dout(n1001));
  jor  g00746(.dina(n354), .dinb(n637), .dout(n1002));
  jor  g00747(.dina(n394), .dinb(n704), .dout(n1003));
  jor  g00748(.dina(n399), .dinb(n772), .dout(n1004));
  jand g00749(.dina(n1004), .dinb(n1003), .dout(n1005));
  jand g00750(.dina(n1005), .dinb(n1002), .dout(n1006));
  jand g00751(.dina(n1006), .dinb(n1001), .dout(n1007));
  jxor g00752(.dina(n1007), .dinb(n364), .dout(n1008));
  jxor g00753(.dina(n1008), .dinb(n1000), .dout(n1009));
  jxor g00754(.dina(n1009), .dinb(n952), .dout(n1010));
  jand g00755(.dina(b14 ), .dinb(b13 ), .dout(n1011));
  jand g00756(.dina(n930), .dinb(n929), .dout(n1012));
  jor  g00757(.dina(n1012), .dinb(n1011), .dout(n1013));
  jxor g00758(.dina(b15 ), .dinb(b14 ), .dout(n1014));
  jnot g00759(.din(n1014), .dout(n1015));
  jxor g00760(.dina(n1015), .dinb(n1013), .dout(n1016));
  jor  g00761(.dina(n1016), .dinb(n296), .dout(n1017));
  jnot g00762(.din(b15 ), .dout(n1018));
  jor  g00763(.dina(n264), .dinb(n1018), .dout(n1019));
  jor  g00764(.dina(n294), .dinb(n934), .dout(n1020));
  jor  g00765(.dina(n280), .dinb(n852), .dout(n1021));
  jand g00766(.dina(n1021), .dinb(n1020), .dout(n1022));
  jand g00767(.dina(n1022), .dinb(n1019), .dout(n1023));
  jand g00768(.dina(n1023), .dinb(n1017), .dout(n1024));
  jxor g00769(.dina(n1024), .dinb(n278), .dout(n1025));
  jxor g00770(.dina(n1025), .dinb(n1010), .dout(n1026));
  jxor g00771(.dina(n1026), .dinb(n947), .dout(f15 ));
  jnot g00772(.din(n1025), .dout(n1028));
  jor  g00773(.dina(n1028), .dinb(n1010), .dout(n1029));
  jor  g00774(.dina(n1026), .dinb(n947), .dout(n1030));
  jand g00775(.dina(n1030), .dinb(n1029), .dout(n1031));
  jand g00776(.dina(n1008), .dinb(n1000), .dout(n1032));
  jnot g00777(.din(n1032), .dout(n1033));
  jnot g00778(.din(n1009), .dout(n1034));
  jor  g00779(.dina(n1034), .dinb(n952), .dout(n1035));
  jand g00780(.dina(n1035), .dinb(n1033), .dout(n1036));
  jand g00781(.dina(n997), .dinb(n989), .dout(n1037));
  jnot g00782(.din(n1037), .dout(n1038));
  jor  g00783(.dina(n999), .dinb(n956), .dout(n1039));
  jand g00784(.dina(n1039), .dinb(n1038), .dout(n1040));
  jor  g00785(.dina(n987), .dinb(n979), .dout(n1041));
  jand g00786(.dina(n988), .dinb(n961), .dout(n1042));
  jnot g00787(.din(n1042), .dout(n1043));
  jand g00788(.dina(n1043), .dinb(n1041), .dout(n1044));
  jnot g00789(.din(n962), .dout(n1045));
  jand g00790(.dina(n964), .dinb(n1045), .dout(n1046));
  jand g00791(.dina(n977), .dinb(n966), .dout(n1047));
  jor  g00792(.dina(n1047), .dinb(n1046), .dout(n1048));
  jxor g00793(.dina(a17 ), .dinb(a16 ), .dout(n1049));
  jnot g00794(.din(n1049), .dout(n1050));
  jand g00795(.dina(n1050), .dinb(n963), .dout(n1051));
  jand g00796(.dina(n1051), .dinb(b1 ), .dout(n1052));
  jand g00797(.dina(n1049), .dinb(n963), .dout(n1053));
  jand g00798(.dina(n1053), .dinb(n259), .dout(n1054));
  jnot g00799(.din(n963), .dout(n1055));
  jxor g00800(.dina(a16 ), .dinb(a15 ), .dout(n1056));
  jand g00801(.dina(n1056), .dinb(n1055), .dout(n1057));
  jand g00802(.dina(n1057), .dinb(b0 ), .dout(n1058));
  jor  g00803(.dina(n1058), .dinb(n1054), .dout(n1059));
  jor  g00804(.dina(n1059), .dinb(n1052), .dout(n1060));
  jnot g00805(.din(a17 ), .dout(n1061));
  jor  g00806(.dina(n965), .dinb(n1061), .dout(n1062));
  jxor g00807(.dina(n1062), .dinb(n1060), .dout(n1063));
  jor  g00808(.dina(n970), .dinb(n337), .dout(n1064));
  jor  g00809(.dina(n967), .dinb(n303), .dout(n1065));
  jor  g00810(.dina(n880), .dinb(n293), .dout(n1066));
  jand g00811(.dina(n1066), .dinb(n1065), .dout(n1067));
  jor  g00812(.dina(n972), .dinb(n340), .dout(n1068));
  jand g00813(.dina(n1068), .dinb(n1067), .dout(n1069));
  jand g00814(.dina(n1069), .dinb(n1064), .dout(n1070));
  jxor g00815(.dina(n1070), .dinb(a14 ), .dout(n1071));
  jxor g00816(.dina(n1071), .dinb(n1063), .dout(n1072));
  jxor g00817(.dina(n1072), .dinb(n1048), .dout(n1073));
  jnot g00818(.din(n1073), .dout(n1074));
  jor  g00819(.dina(n728), .dinb(n466), .dout(n1075));
  jor  g00820(.dina(n731), .dinb(n415), .dout(n1076));
  jor  g00821(.dina(n660), .dinb(n377), .dout(n1077));
  jand g00822(.dina(n1077), .dinb(n1076), .dout(n1078));
  jor  g00823(.dina(n726), .dinb(n469), .dout(n1079));
  jand g00824(.dina(n1079), .dinb(n1078), .dout(n1080));
  jand g00825(.dina(n1080), .dinb(n1075), .dout(n1081));
  jxor g00826(.dina(n1081), .dinb(a11 ), .dout(n1082));
  jxor g00827(.dina(n1082), .dinb(n1074), .dout(n1083));
  jnot g00828(.din(n1083), .dout(n1084));
  jxor g00829(.dina(n1084), .dinb(n1044), .dout(n1085));
  jor  g00830(.dina(n635), .dinb(n544), .dout(n1086));
  jor  g00831(.dina(n486), .dinb(n519), .dout(n1087));
  jor  g00832(.dina(n542), .dinb(n637), .dout(n1088));
  jor  g00833(.dina(n547), .dinb(n572), .dout(n1089));
  jand g00834(.dina(n1089), .dinb(n1088), .dout(n1090));
  jand g00835(.dina(n1090), .dinb(n1087), .dout(n1091));
  jand g00836(.dina(n1091), .dinb(n1086), .dout(n1092));
  jxor g00837(.dina(n1092), .dinb(n446), .dout(n1093));
  jxor g00838(.dina(n1093), .dinb(n1085), .dout(n1094));
  jxor g00839(.dina(n1094), .dinb(n1040), .dout(n1095));
  jor  g00840(.dina(n850), .dinb(n397), .dout(n1096));
  jor  g00841(.dina(n354), .dinb(n704), .dout(n1097));
  jor  g00842(.dina(n394), .dinb(n772), .dout(n1098));
  jor  g00843(.dina(n399), .dinb(n852), .dout(n1099));
  jand g00844(.dina(n1099), .dinb(n1098), .dout(n1100));
  jand g00845(.dina(n1100), .dinb(n1097), .dout(n1101));
  jand g00846(.dina(n1101), .dinb(n1096), .dout(n1102));
  jxor g00847(.dina(n1102), .dinb(n364), .dout(n1103));
  jxor g00848(.dina(n1103), .dinb(n1095), .dout(n1104));
  jnot g00849(.din(n1104), .dout(n1105));
  jxor g00850(.dina(n1105), .dinb(n1036), .dout(n1106));
  jand g00851(.dina(b15 ), .dinb(b14 ), .dout(n1107));
  jand g00852(.dina(n1014), .dinb(n1013), .dout(n1108));
  jor  g00853(.dina(n1108), .dinb(n1107), .dout(n1109));
  jxor g00854(.dina(b16 ), .dinb(b15 ), .dout(n1110));
  jnot g00855(.din(n1110), .dout(n1111));
  jxor g00856(.dina(n1111), .dinb(n1109), .dout(n1112));
  jor  g00857(.dina(n1112), .dinb(n296), .dout(n1113));
  jnot g00858(.din(b16 ), .dout(n1114));
  jor  g00859(.dina(n264), .dinb(n1114), .dout(n1115));
  jor  g00860(.dina(n294), .dinb(n1018), .dout(n1116));
  jor  g00861(.dina(n280), .dinb(n934), .dout(n1117));
  jand g00862(.dina(n1117), .dinb(n1116), .dout(n1118));
  jand g00863(.dina(n1118), .dinb(n1115), .dout(n1119));
  jand g00864(.dina(n1119), .dinb(n1113), .dout(n1120));
  jxor g00865(.dina(n1120), .dinb(n278), .dout(n1121));
  jxor g00866(.dina(n1121), .dinb(n1106), .dout(n1122));
  jxor g00867(.dina(n1122), .dinb(n1031), .dout(f16 ));
  jnot g00868(.din(n1121), .dout(n1124));
  jor  g00869(.dina(n1124), .dinb(n1106), .dout(n1125));
  jor  g00870(.dina(n1122), .dinb(n1031), .dout(n1126));
  jand g00871(.dina(n1126), .dinb(n1125), .dout(n1127));
  jnot g00872(.din(n1095), .dout(n1128));
  jand g00873(.dina(n1103), .dinb(n1128), .dout(n1129));
  jnot g00874(.din(n1129), .dout(n1130));
  jor  g00875(.dina(n1104), .dinb(n1036), .dout(n1131));
  jand g00876(.dina(n1131), .dinb(n1130), .dout(n1132));
  jand g00877(.dina(n1093), .dinb(n1085), .dout(n1133));
  jnot g00878(.din(n1040), .dout(n1134));
  jand g00879(.dina(n1094), .dinb(n1134), .dout(n1135));
  jor  g00880(.dina(n1135), .dinb(n1133), .dout(n1136));
  jor  g00881(.dina(n1082), .dinb(n1074), .dout(n1137));
  jor  g00882(.dina(n1084), .dinb(n1044), .dout(n1138));
  jand g00883(.dina(n1138), .dinb(n1137), .dout(n1139));
  jor  g00884(.dina(n1071), .dinb(n1063), .dout(n1140));
  jand g00885(.dina(n1072), .dinb(n1048), .dout(n1141));
  jnot g00886(.din(n1141), .dout(n1142));
  jand g00887(.dina(n1142), .dinb(n1140), .dout(n1143));
  jnot g00888(.din(n1143), .dout(n1144));
  jand g00889(.dina(n1057), .dinb(b1 ), .dout(n1145));
  jor  g00890(.dina(n1056), .dinb(n963), .dout(n1146));
  jor  g00891(.dina(n1146), .dinb(n1050), .dout(n1147));
  jnot g00892(.din(n1147), .dout(n1148));
  jand g00893(.dina(n1148), .dinb(b0 ), .dout(n1149));
  jand g00894(.dina(n1053), .dinb(n273), .dout(n1150));
  jand g00895(.dina(n1051), .dinb(b2 ), .dout(n1151));
  jor  g00896(.dina(n1151), .dinb(n1150), .dout(n1152));
  jor  g00897(.dina(n1152), .dinb(n1149), .dout(n1153));
  jor  g00898(.dina(n1153), .dinb(n1145), .dout(n1154));
  jnot g00899(.din(n1060), .dout(n1155));
  jand g00900(.dina(n965), .dinb(a17 ), .dout(n1156));
  jand g00901(.dina(n1156), .dinb(n1155), .dout(n1157));
  jnot g00902(.din(n1157), .dout(n1158));
  jand g00903(.dina(n1158), .dinb(a17 ), .dout(n1159));
  jxor g00904(.dina(n1159), .dinb(n1154), .dout(n1160));
  jnot g00905(.din(n1160), .dout(n1161));
  jor  g00906(.dina(n970), .dinb(n374), .dout(n1162));
  jor  g00907(.dina(n967), .dinb(n340), .dout(n1163));
  jor  g00908(.dina(n880), .dinb(n303), .dout(n1164));
  jand g00909(.dina(n1164), .dinb(n1163), .dout(n1165));
  jor  g00910(.dina(n972), .dinb(n377), .dout(n1166));
  jand g00911(.dina(n1166), .dinb(n1165), .dout(n1167));
  jand g00912(.dina(n1167), .dinb(n1162), .dout(n1168));
  jxor g00913(.dina(n1168), .dinb(a14 ), .dout(n1169));
  jxor g00914(.dina(n1169), .dinb(n1161), .dout(n1170));
  jxor g00915(.dina(n1170), .dinb(n1144), .dout(n1171));
  jnot g00916(.din(n1171), .dout(n1172));
  jor  g00917(.dina(n728), .dinb(n517), .dout(n1173));
  jor  g00918(.dina(n731), .dinb(n469), .dout(n1174));
  jor  g00919(.dina(n726), .dinb(n519), .dout(n1175));
  jor  g00920(.dina(n660), .dinb(n415), .dout(n1176));
  jand g00921(.dina(n1176), .dinb(n1175), .dout(n1177));
  jand g00922(.dina(n1177), .dinb(n1174), .dout(n1178));
  jand g00923(.dina(n1178), .dinb(n1173), .dout(n1179));
  jxor g00924(.dina(n1179), .dinb(a11 ), .dout(n1180));
  jxor g00925(.dina(n1180), .dinb(n1172), .dout(n1181));
  jnot g00926(.din(n1181), .dout(n1182));
  jxor g00927(.dina(n1182), .dinb(n1139), .dout(n1183));
  jor  g00928(.dina(n702), .dinb(n544), .dout(n1184));
  jor  g00929(.dina(n486), .dinb(n572), .dout(n1185));
  jor  g00930(.dina(n542), .dinb(n704), .dout(n1186));
  jor  g00931(.dina(n547), .dinb(n637), .dout(n1187));
  jand g00932(.dina(n1187), .dinb(n1186), .dout(n1188));
  jand g00933(.dina(n1188), .dinb(n1185), .dout(n1189));
  jand g00934(.dina(n1189), .dinb(n1184), .dout(n1190));
  jxor g00935(.dina(n1190), .dinb(n446), .dout(n1191));
  jxor g00936(.dina(n1191), .dinb(n1183), .dout(n1192));
  jxor g00937(.dina(n1192), .dinb(n1136), .dout(n1193));
  jor  g00938(.dina(n932), .dinb(n397), .dout(n1194));
  jor  g00939(.dina(n354), .dinb(n772), .dout(n1195));
  jor  g00940(.dina(n394), .dinb(n852), .dout(n1196));
  jor  g00941(.dina(n399), .dinb(n934), .dout(n1197));
  jand g00942(.dina(n1197), .dinb(n1196), .dout(n1198));
  jand g00943(.dina(n1198), .dinb(n1195), .dout(n1199));
  jand g00944(.dina(n1199), .dinb(n1194), .dout(n1200));
  jxor g00945(.dina(n1200), .dinb(n364), .dout(n1201));
  jxor g00946(.dina(n1201), .dinb(n1193), .dout(n1202));
  jxor g00947(.dina(n1202), .dinb(n1132), .dout(n1203));
  jand g00948(.dina(b16 ), .dinb(b15 ), .dout(n1204));
  jand g00949(.dina(n1110), .dinb(n1109), .dout(n1205));
  jor  g00950(.dina(n1205), .dinb(n1204), .dout(n1206));
  jxor g00951(.dina(b17 ), .dinb(b16 ), .dout(n1207));
  jnot g00952(.din(n1207), .dout(n1208));
  jxor g00953(.dina(n1208), .dinb(n1206), .dout(n1209));
  jor  g00954(.dina(n1209), .dinb(n296), .dout(n1210));
  jnot g00955(.din(b17 ), .dout(n1211));
  jor  g00956(.dina(n264), .dinb(n1211), .dout(n1212));
  jor  g00957(.dina(n294), .dinb(n1114), .dout(n1213));
  jor  g00958(.dina(n280), .dinb(n1018), .dout(n1214));
  jand g00959(.dina(n1214), .dinb(n1213), .dout(n1215));
  jand g00960(.dina(n1215), .dinb(n1212), .dout(n1216));
  jand g00961(.dina(n1216), .dinb(n1210), .dout(n1217));
  jxor g00962(.dina(n1217), .dinb(n278), .dout(n1218));
  jxor g00963(.dina(n1218), .dinb(n1203), .dout(n1219));
  jxor g00964(.dina(n1219), .dinb(n1127), .dout(f17 ));
  jnot g00965(.din(n1218), .dout(n1221));
  jor  g00966(.dina(n1221), .dinb(n1203), .dout(n1222));
  jor  g00967(.dina(n1219), .dinb(n1127), .dout(n1223));
  jand g00968(.dina(n1223), .dinb(n1222), .dout(n1224));
  jand g00969(.dina(n1201), .dinb(n1193), .dout(n1225));
  jnot g00970(.din(n1225), .dout(n1226));
  jnot g00971(.din(n1202), .dout(n1227));
  jor  g00972(.dina(n1227), .dinb(n1132), .dout(n1228));
  jand g00973(.dina(n1228), .dinb(n1226), .dout(n1229));
  jand g00974(.dina(n1191), .dinb(n1183), .dout(n1230));
  jand g00975(.dina(n1192), .dinb(n1136), .dout(n1231));
  jor  g00976(.dina(n1231), .dinb(n1230), .dout(n1232));
  jor  g00977(.dina(n1180), .dinb(n1172), .dout(n1233));
  jor  g00978(.dina(n1182), .dinb(n1139), .dout(n1234));
  jand g00979(.dina(n1234), .dinb(n1233), .dout(n1235));
  jor  g00980(.dina(n1169), .dinb(n1161), .dout(n1236));
  jand g00981(.dina(n1170), .dinb(n1144), .dout(n1237));
  jnot g00982(.din(n1237), .dout(n1238));
  jand g00983(.dina(n1238), .dinb(n1236), .dout(n1239));
  jnot g00984(.din(n1239), .dout(n1240));
  jor  g00985(.dina(n1158), .dinb(n1154), .dout(n1241));
  jxor g00986(.dina(a18 ), .dinb(a17 ), .dout(n1242));
  jand g00987(.dina(n1242), .dinb(b0 ), .dout(n1243));
  jnot g00988(.din(n1243), .dout(n1244));
  jxor g00989(.dina(n1244), .dinb(n1241), .dout(n1245));
  jnot g00990(.din(n1051), .dout(n1246));
  jor  g00991(.dina(n1246), .dinb(n303), .dout(n1247));
  jnot g00992(.din(n1053), .dout(n1248));
  jor  g00993(.dina(n1248), .dinb(n301), .dout(n1249));
  jor  g00994(.dina(n1147), .dinb(n305), .dout(n1250));
  jnot g00995(.din(n1057), .dout(n1251));
  jor  g00996(.dina(n1251), .dinb(n293), .dout(n1252));
  jand g00997(.dina(n1252), .dinb(n1250), .dout(n1253));
  jand g00998(.dina(n1253), .dinb(n1249), .dout(n1254));
  jand g00999(.dina(n1254), .dinb(n1247), .dout(n1255));
  jxor g01000(.dina(n1255), .dinb(n1061), .dout(n1256));
  jxor g01001(.dina(n1256), .dinb(n1245), .dout(n1257));
  jnot g01002(.din(n1257), .dout(n1258));
  jor  g01003(.dina(n970), .dinb(n412), .dout(n1259));
  jor  g01004(.dina(n972), .dinb(n415), .dout(n1260));
  jor  g01005(.dina(n880), .dinb(n340), .dout(n1261));
  jand g01006(.dina(n1261), .dinb(n1260), .dout(n1262));
  jor  g01007(.dina(n967), .dinb(n377), .dout(n1263));
  jand g01008(.dina(n1263), .dinb(n1262), .dout(n1264));
  jand g01009(.dina(n1264), .dinb(n1259), .dout(n1265));
  jxor g01010(.dina(n1265), .dinb(a14 ), .dout(n1266));
  jxor g01011(.dina(n1266), .dinb(n1258), .dout(n1267));
  jxor g01012(.dina(n1267), .dinb(n1240), .dout(n1268));
  jor  g01013(.dina(n728), .dinb(n570), .dout(n1269));
  jor  g01014(.dina(n660), .dinb(n469), .dout(n1270));
  jor  g01015(.dina(n731), .dinb(n519), .dout(n1271));
  jor  g01016(.dina(n726), .dinb(n572), .dout(n1272));
  jand g01017(.dina(n1272), .dinb(n1271), .dout(n1273));
  jand g01018(.dina(n1273), .dinb(n1270), .dout(n1274));
  jand g01019(.dina(n1274), .dinb(n1269), .dout(n1275));
  jxor g01020(.dina(n1275), .dinb(n606), .dout(n1276));
  jxor g01021(.dina(n1276), .dinb(n1268), .dout(n1277));
  jnot g01022(.din(n1277), .dout(n1278));
  jxor g01023(.dina(n1278), .dinb(n1235), .dout(n1279));
  jor  g01024(.dina(n770), .dinb(n544), .dout(n1280));
  jor  g01025(.dina(n486), .dinb(n637), .dout(n1281));
  jor  g01026(.dina(n547), .dinb(n704), .dout(n1282));
  jor  g01027(.dina(n542), .dinb(n772), .dout(n1283));
  jand g01028(.dina(n1283), .dinb(n1282), .dout(n1284));
  jand g01029(.dina(n1284), .dinb(n1281), .dout(n1285));
  jand g01030(.dina(n1285), .dinb(n1280), .dout(n1286));
  jxor g01031(.dina(n1286), .dinb(n446), .dout(n1287));
  jxor g01032(.dina(n1287), .dinb(n1279), .dout(n1288));
  jxor g01033(.dina(n1288), .dinb(n1232), .dout(n1289));
  jor  g01034(.dina(n1016), .dinb(n397), .dout(n1290));
  jor  g01035(.dina(n354), .dinb(n852), .dout(n1291));
  jor  g01036(.dina(n399), .dinb(n1018), .dout(n1292));
  jor  g01037(.dina(n394), .dinb(n934), .dout(n1293));
  jand g01038(.dina(n1293), .dinb(n1292), .dout(n1294));
  jand g01039(.dina(n1294), .dinb(n1291), .dout(n1295));
  jand g01040(.dina(n1295), .dinb(n1290), .dout(n1296));
  jxor g01041(.dina(n1296), .dinb(n364), .dout(n1297));
  jxor g01042(.dina(n1297), .dinb(n1289), .dout(n1298));
  jxor g01043(.dina(n1298), .dinb(n1229), .dout(n1299));
  jand g01044(.dina(b17 ), .dinb(b16 ), .dout(n1300));
  jand g01045(.dina(n1207), .dinb(n1206), .dout(n1301));
  jor  g01046(.dina(n1301), .dinb(n1300), .dout(n1302));
  jxor g01047(.dina(b18 ), .dinb(b17 ), .dout(n1303));
  jnot g01048(.din(n1303), .dout(n1304));
  jxor g01049(.dina(n1304), .dinb(n1302), .dout(n1305));
  jor  g01050(.dina(n1305), .dinb(n296), .dout(n1306));
  jnot g01051(.din(b18 ), .dout(n1307));
  jor  g01052(.dina(n264), .dinb(n1307), .dout(n1308));
  jor  g01053(.dina(n294), .dinb(n1211), .dout(n1309));
  jor  g01054(.dina(n280), .dinb(n1114), .dout(n1310));
  jand g01055(.dina(n1310), .dinb(n1309), .dout(n1311));
  jand g01056(.dina(n1311), .dinb(n1308), .dout(n1312));
  jand g01057(.dina(n1312), .dinb(n1306), .dout(n1313));
  jxor g01058(.dina(n1313), .dinb(n278), .dout(n1314));
  jxor g01059(.dina(n1314), .dinb(n1299), .dout(n1315));
  jxor g01060(.dina(n1315), .dinb(n1224), .dout(f18 ));
  jnot g01061(.din(n1314), .dout(n1317));
  jor  g01062(.dina(n1317), .dinb(n1299), .dout(n1318));
  jor  g01063(.dina(n1315), .dinb(n1224), .dout(n1319));
  jand g01064(.dina(n1319), .dinb(n1318), .dout(n1320));
  jand g01065(.dina(n1297), .dinb(n1289), .dout(n1321));
  jnot g01066(.din(n1321), .dout(n1322));
  jnot g01067(.din(n1298), .dout(n1323));
  jor  g01068(.dina(n1323), .dinb(n1229), .dout(n1324));
  jand g01069(.dina(n1324), .dinb(n1322), .dout(n1325));
  jand g01070(.dina(n1276), .dinb(n1268), .dout(n1326));
  jnot g01071(.din(n1326), .dout(n1327));
  jor  g01072(.dina(n1278), .dinb(n1235), .dout(n1328));
  jand g01073(.dina(n1328), .dinb(n1327), .dout(n1329));
  jor  g01074(.dina(n1266), .dinb(n1258), .dout(n1330));
  jand g01075(.dina(n1267), .dinb(n1240), .dout(n1331));
  jnot g01076(.din(n1331), .dout(n1332));
  jand g01077(.dina(n1332), .dinb(n1330), .dout(n1333));
  jnot g01078(.din(n1333), .dout(n1334));
  jnot g01079(.din(n1241), .dout(n1335));
  jand g01080(.dina(n1243), .dinb(n1335), .dout(n1336));
  jand g01081(.dina(n1256), .dinb(n1245), .dout(n1337));
  jor  g01082(.dina(n1337), .dinb(n1336), .dout(n1338));
  jxor g01083(.dina(a20 ), .dinb(a19 ), .dout(n1339));
  jand g01084(.dina(n1339), .dinb(n1242), .dout(n1340));
  jand g01085(.dina(n1340), .dinb(n259), .dout(n1341));
  jnot g01086(.din(n1242), .dout(n1342));
  jxor g01087(.dina(a19 ), .dinb(a18 ), .dout(n1343));
  jand g01088(.dina(n1343), .dinb(n1342), .dout(n1344));
  jand g01089(.dina(n1344), .dinb(b0 ), .dout(n1345));
  jnot g01090(.din(n1339), .dout(n1346));
  jand g01091(.dina(n1346), .dinb(n1242), .dout(n1347));
  jand g01092(.dina(n1347), .dinb(b1 ), .dout(n1348));
  jor  g01093(.dina(n1348), .dinb(n1345), .dout(n1349));
  jor  g01094(.dina(n1349), .dinb(n1341), .dout(n1350));
  jnot g01095(.din(a20 ), .dout(n1351));
  jor  g01096(.dina(n1244), .dinb(n1351), .dout(n1352));
  jxor g01097(.dina(n1352), .dinb(n1350), .dout(n1353));
  jor  g01098(.dina(n1248), .dinb(n337), .dout(n1354));
  jor  g01099(.dina(n1251), .dinb(n303), .dout(n1355));
  jor  g01100(.dina(n1147), .dinb(n293), .dout(n1356));
  jand g01101(.dina(n1356), .dinb(n1355), .dout(n1357));
  jor  g01102(.dina(n1246), .dinb(n340), .dout(n1358));
  jand g01103(.dina(n1358), .dinb(n1357), .dout(n1359));
  jand g01104(.dina(n1359), .dinb(n1354), .dout(n1360));
  jxor g01105(.dina(n1360), .dinb(a17 ), .dout(n1361));
  jxor g01106(.dina(n1361), .dinb(n1353), .dout(n1362));
  jxor g01107(.dina(n1362), .dinb(n1338), .dout(n1363));
  jnot g01108(.din(n1363), .dout(n1364));
  jor  g01109(.dina(n970), .dinb(n466), .dout(n1365));
  jor  g01110(.dina(n972), .dinb(n469), .dout(n1366));
  jor  g01111(.dina(n880), .dinb(n377), .dout(n1367));
  jand g01112(.dina(n1367), .dinb(n1366), .dout(n1368));
  jor  g01113(.dina(n967), .dinb(n415), .dout(n1369));
  jand g01114(.dina(n1369), .dinb(n1368), .dout(n1370));
  jand g01115(.dina(n1370), .dinb(n1365), .dout(n1371));
  jxor g01116(.dina(n1371), .dinb(a14 ), .dout(n1372));
  jxor g01117(.dina(n1372), .dinb(n1364), .dout(n1373));
  jxor g01118(.dina(n1373), .dinb(n1334), .dout(n1374));
  jor  g01119(.dina(n635), .dinb(n728), .dout(n1375));
  jor  g01120(.dina(n660), .dinb(n519), .dout(n1376));
  jor  g01121(.dina(n726), .dinb(n637), .dout(n1377));
  jor  g01122(.dina(n731), .dinb(n572), .dout(n1378));
  jand g01123(.dina(n1378), .dinb(n1377), .dout(n1379));
  jand g01124(.dina(n1379), .dinb(n1376), .dout(n1380));
  jand g01125(.dina(n1380), .dinb(n1375), .dout(n1381));
  jxor g01126(.dina(n1381), .dinb(n606), .dout(n1382));
  jxor g01127(.dina(n1382), .dinb(n1374), .dout(n1383));
  jnot g01128(.din(n1383), .dout(n1384));
  jxor g01129(.dina(n1384), .dinb(n1329), .dout(n1385));
  jor  g01130(.dina(n850), .dinb(n544), .dout(n1386));
  jor  g01131(.dina(n486), .dinb(n704), .dout(n1387));
  jor  g01132(.dina(n542), .dinb(n852), .dout(n1388));
  jor  g01133(.dina(n547), .dinb(n772), .dout(n1389));
  jand g01134(.dina(n1389), .dinb(n1388), .dout(n1390));
  jand g01135(.dina(n1390), .dinb(n1387), .dout(n1391));
  jand g01136(.dina(n1391), .dinb(n1386), .dout(n1392));
  jxor g01137(.dina(n1392), .dinb(n446), .dout(n1393));
  jxor g01138(.dina(n1393), .dinb(n1385), .dout(n1394));
  jand g01139(.dina(n1287), .dinb(n1279), .dout(n1395));
  jand g01140(.dina(n1288), .dinb(n1232), .dout(n1396));
  jor  g01141(.dina(n1396), .dinb(n1395), .dout(n1397));
  jxor g01142(.dina(n1397), .dinb(n1394), .dout(n1398));
  jor  g01143(.dina(n1112), .dinb(n397), .dout(n1399));
  jor  g01144(.dina(n354), .dinb(n934), .dout(n1400));
  jor  g01145(.dina(n394), .dinb(n1018), .dout(n1401));
  jor  g01146(.dina(n399), .dinb(n1114), .dout(n1402));
  jand g01147(.dina(n1402), .dinb(n1401), .dout(n1403));
  jand g01148(.dina(n1403), .dinb(n1400), .dout(n1404));
  jand g01149(.dina(n1404), .dinb(n1399), .dout(n1405));
  jxor g01150(.dina(n1405), .dinb(n364), .dout(n1406));
  jxor g01151(.dina(n1406), .dinb(n1398), .dout(n1407));
  jxor g01152(.dina(n1407), .dinb(n1325), .dout(n1408));
  jand g01153(.dina(b18 ), .dinb(b17 ), .dout(n1409));
  jand g01154(.dina(n1303), .dinb(n1302), .dout(n1410));
  jor  g01155(.dina(n1410), .dinb(n1409), .dout(n1411));
  jxor g01156(.dina(b19 ), .dinb(b18 ), .dout(n1412));
  jnot g01157(.din(n1412), .dout(n1413));
  jxor g01158(.dina(n1413), .dinb(n1411), .dout(n1414));
  jor  g01159(.dina(n1414), .dinb(n296), .dout(n1415));
  jnot g01160(.din(b19 ), .dout(n1416));
  jor  g01161(.dina(n264), .dinb(n1416), .dout(n1417));
  jor  g01162(.dina(n294), .dinb(n1307), .dout(n1418));
  jor  g01163(.dina(n280), .dinb(n1211), .dout(n1419));
  jand g01164(.dina(n1419), .dinb(n1418), .dout(n1420));
  jand g01165(.dina(n1420), .dinb(n1417), .dout(n1421));
  jand g01166(.dina(n1421), .dinb(n1415), .dout(n1422));
  jxor g01167(.dina(n1422), .dinb(n278), .dout(n1423));
  jxor g01168(.dina(n1423), .dinb(n1408), .dout(n1424));
  jxor g01169(.dina(n1424), .dinb(n1320), .dout(f19 ));
  jnot g01170(.din(n1423), .dout(n1426));
  jor  g01171(.dina(n1426), .dinb(n1408), .dout(n1427));
  jor  g01172(.dina(n1424), .dinb(n1320), .dout(n1428));
  jand g01173(.dina(n1428), .dinb(n1427), .dout(n1429));
  jand g01174(.dina(n1406), .dinb(n1398), .dout(n1430));
  jnot g01175(.din(n1430), .dout(n1431));
  jnot g01176(.din(n1407), .dout(n1432));
  jor  g01177(.dina(n1432), .dinb(n1325), .dout(n1433));
  jand g01178(.dina(n1433), .dinb(n1431), .dout(n1434));
  jand g01179(.dina(n1393), .dinb(n1385), .dout(n1435));
  jand g01180(.dina(n1397), .dinb(n1394), .dout(n1436));
  jor  g01181(.dina(n1436), .dinb(n1435), .dout(n1437));
  jand g01182(.dina(n1382), .dinb(n1374), .dout(n1438));
  jnot g01183(.din(n1438), .dout(n1439));
  jor  g01184(.dina(n1384), .dinb(n1329), .dout(n1440));
  jand g01185(.dina(n1440), .dinb(n1439), .dout(n1441));
  jor  g01186(.dina(n1372), .dinb(n1364), .dout(n1442));
  jand g01187(.dina(n1373), .dinb(n1334), .dout(n1443));
  jnot g01188(.din(n1443), .dout(n1444));
  jand g01189(.dina(n1444), .dinb(n1442), .dout(n1445));
  jnot g01190(.din(n1445), .dout(n1446));
  jor  g01191(.dina(n1361), .dinb(n1353), .dout(n1447));
  jand g01192(.dina(n1362), .dinb(n1338), .dout(n1448));
  jnot g01193(.din(n1448), .dout(n1449));
  jand g01194(.dina(n1449), .dinb(n1447), .dout(n1450));
  jnot g01195(.din(n1450), .dout(n1451));
  jor  g01196(.dina(n1343), .dinb(n1242), .dout(n1452));
  jor  g01197(.dina(n1452), .dinb(n1346), .dout(n1453));
  jnot g01198(.din(n1453), .dout(n1454));
  jand g01199(.dina(n1454), .dinb(b0 ), .dout(n1455));
  jand g01200(.dina(n1344), .dinb(b1 ), .dout(n1456));
  jor  g01201(.dina(n1456), .dinb(n1455), .dout(n1457));
  jand g01202(.dina(n1340), .dinb(n273), .dout(n1458));
  jand g01203(.dina(n1347), .dinb(b2 ), .dout(n1459));
  jor  g01204(.dina(n1459), .dinb(n1458), .dout(n1460));
  jor  g01205(.dina(n1460), .dinb(n1457), .dout(n1461));
  jnot g01206(.din(n1350), .dout(n1462));
  jand g01207(.dina(n1244), .dinb(a20 ), .dout(n1463));
  jand g01208(.dina(n1463), .dinb(n1462), .dout(n1464));
  jnot g01209(.din(n1464), .dout(n1465));
  jand g01210(.dina(n1465), .dinb(a20 ), .dout(n1466));
  jxor g01211(.dina(n1466), .dinb(n1461), .dout(n1467));
  jnot g01212(.din(n1467), .dout(n1468));
  jor  g01213(.dina(n1248), .dinb(n374), .dout(n1469));
  jor  g01214(.dina(n1251), .dinb(n340), .dout(n1470));
  jor  g01215(.dina(n1147), .dinb(n303), .dout(n1471));
  jand g01216(.dina(n1471), .dinb(n1470), .dout(n1472));
  jor  g01217(.dina(n1246), .dinb(n377), .dout(n1473));
  jand g01218(.dina(n1473), .dinb(n1472), .dout(n1474));
  jand g01219(.dina(n1474), .dinb(n1469), .dout(n1475));
  jxor g01220(.dina(n1475), .dinb(a17 ), .dout(n1476));
  jxor g01221(.dina(n1476), .dinb(n1468), .dout(n1477));
  jxor g01222(.dina(n1477), .dinb(n1451), .dout(n1478));
  jor  g01223(.dina(n970), .dinb(n517), .dout(n1479));
  jor  g01224(.dina(n967), .dinb(n469), .dout(n1480));
  jor  g01225(.dina(n972), .dinb(n519), .dout(n1481));
  jor  g01226(.dina(n880), .dinb(n415), .dout(n1482));
  jand g01227(.dina(n1482), .dinb(n1481), .dout(n1483));
  jand g01228(.dina(n1483), .dinb(n1480), .dout(n1484));
  jand g01229(.dina(n1484), .dinb(n1479), .dout(n1485));
  jxor g01230(.dina(n1485), .dinb(n810), .dout(n1486));
  jxor g01231(.dina(n1486), .dinb(n1478), .dout(n1487));
  jxor g01232(.dina(n1487), .dinb(n1446), .dout(n1488));
  jor  g01233(.dina(n702), .dinb(n728), .dout(n1489));
  jor  g01234(.dina(n660), .dinb(n572), .dout(n1490));
  jor  g01235(.dina(n726), .dinb(n704), .dout(n1491));
  jor  g01236(.dina(n731), .dinb(n637), .dout(n1492));
  jand g01237(.dina(n1492), .dinb(n1491), .dout(n1493));
  jand g01238(.dina(n1493), .dinb(n1490), .dout(n1494));
  jand g01239(.dina(n1494), .dinb(n1489), .dout(n1495));
  jxor g01240(.dina(n1495), .dinb(n606), .dout(n1496));
  jxor g01241(.dina(n1496), .dinb(n1488), .dout(n1497));
  jnot g01242(.din(n1497), .dout(n1498));
  jxor g01243(.dina(n1498), .dinb(n1441), .dout(n1499));
  jor  g01244(.dina(n932), .dinb(n544), .dout(n1500));
  jor  g01245(.dina(n486), .dinb(n772), .dout(n1501));
  jor  g01246(.dina(n547), .dinb(n852), .dout(n1502));
  jor  g01247(.dina(n542), .dinb(n934), .dout(n1503));
  jand g01248(.dina(n1503), .dinb(n1502), .dout(n1504));
  jand g01249(.dina(n1504), .dinb(n1501), .dout(n1505));
  jand g01250(.dina(n1505), .dinb(n1500), .dout(n1506));
  jxor g01251(.dina(n1506), .dinb(n446), .dout(n1507));
  jxor g01252(.dina(n1507), .dinb(n1499), .dout(n1508));
  jxor g01253(.dina(n1508), .dinb(n1437), .dout(n1509));
  jor  g01254(.dina(n1209), .dinb(n397), .dout(n1510));
  jor  g01255(.dina(n354), .dinb(n1018), .dout(n1511));
  jor  g01256(.dina(n399), .dinb(n1211), .dout(n1512));
  jor  g01257(.dina(n394), .dinb(n1114), .dout(n1513));
  jand g01258(.dina(n1513), .dinb(n1512), .dout(n1514));
  jand g01259(.dina(n1514), .dinb(n1511), .dout(n1515));
  jand g01260(.dina(n1515), .dinb(n1510), .dout(n1516));
  jxor g01261(.dina(n1516), .dinb(n364), .dout(n1517));
  jxor g01262(.dina(n1517), .dinb(n1509), .dout(n1518));
  jxor g01263(.dina(n1518), .dinb(n1434), .dout(n1519));
  jand g01264(.dina(b19 ), .dinb(b18 ), .dout(n1520));
  jand g01265(.dina(n1412), .dinb(n1411), .dout(n1521));
  jor  g01266(.dina(n1521), .dinb(n1520), .dout(n1522));
  jxor g01267(.dina(b20 ), .dinb(b19 ), .dout(n1523));
  jnot g01268(.din(n1523), .dout(n1524));
  jxor g01269(.dina(n1524), .dinb(n1522), .dout(n1525));
  jor  g01270(.dina(n1525), .dinb(n296), .dout(n1526));
  jnot g01271(.din(b20 ), .dout(n1527));
  jor  g01272(.dina(n264), .dinb(n1527), .dout(n1528));
  jor  g01273(.dina(n280), .dinb(n1307), .dout(n1529));
  jor  g01274(.dina(n294), .dinb(n1416), .dout(n1530));
  jand g01275(.dina(n1530), .dinb(n1529), .dout(n1531));
  jand g01276(.dina(n1531), .dinb(n1528), .dout(n1532));
  jand g01277(.dina(n1532), .dinb(n1526), .dout(n1533));
  jxor g01278(.dina(n1533), .dinb(n278), .dout(n1534));
  jxor g01279(.dina(n1534), .dinb(n1519), .dout(n1535));
  jxor g01280(.dina(n1535), .dinb(n1429), .dout(f20 ));
  jnot g01281(.din(n1534), .dout(n1537));
  jor  g01282(.dina(n1537), .dinb(n1519), .dout(n1538));
  jor  g01283(.dina(n1535), .dinb(n1429), .dout(n1539));
  jand g01284(.dina(n1539), .dinb(n1538), .dout(n1540));
  jand g01285(.dina(n1517), .dinb(n1509), .dout(n1541));
  jnot g01286(.din(n1541), .dout(n1542));
  jnot g01287(.din(n1518), .dout(n1543));
  jor  g01288(.dina(n1543), .dinb(n1434), .dout(n1544));
  jand g01289(.dina(n1544), .dinb(n1542), .dout(n1545));
  jand g01290(.dina(n1507), .dinb(n1499), .dout(n1546));
  jand g01291(.dina(n1508), .dinb(n1437), .dout(n1547));
  jor  g01292(.dina(n1547), .dinb(n1546), .dout(n1548));
  jand g01293(.dina(n1496), .dinb(n1488), .dout(n1549));
  jnot g01294(.din(n1549), .dout(n1550));
  jor  g01295(.dina(n1498), .dinb(n1441), .dout(n1551));
  jand g01296(.dina(n1551), .dinb(n1550), .dout(n1552));
  jand g01297(.dina(n1486), .dinb(n1478), .dout(n1553));
  jand g01298(.dina(n1487), .dinb(n1446), .dout(n1554));
  jor  g01299(.dina(n1554), .dinb(n1553), .dout(n1555));
  jor  g01300(.dina(n1476), .dinb(n1468), .dout(n1556));
  jand g01301(.dina(n1477), .dinb(n1451), .dout(n1557));
  jnot g01302(.din(n1557), .dout(n1558));
  jand g01303(.dina(n1558), .dinb(n1556), .dout(n1559));
  jnot g01304(.din(n1559), .dout(n1560));
  jor  g01305(.dina(n1465), .dinb(n1461), .dout(n1561));
  jxor g01306(.dina(a21 ), .dinb(a20 ), .dout(n1562));
  jand g01307(.dina(n1562), .dinb(b0 ), .dout(n1563));
  jnot g01308(.din(n1563), .dout(n1564));
  jxor g01309(.dina(n1564), .dinb(n1561), .dout(n1565));
  jnot g01310(.din(n1344), .dout(n1566));
  jor  g01311(.dina(n1566), .dinb(n293), .dout(n1567));
  jor  g01312(.dina(n1453), .dinb(n305), .dout(n1568));
  jnot g01313(.din(n1340), .dout(n1569));
  jor  g01314(.dina(n1569), .dinb(n301), .dout(n1570));
  jnot g01315(.din(n1347), .dout(n1571));
  jor  g01316(.dina(n1571), .dinb(n303), .dout(n1572));
  jand g01317(.dina(n1572), .dinb(n1570), .dout(n1573));
  jand g01318(.dina(n1573), .dinb(n1568), .dout(n1574));
  jand g01319(.dina(n1574), .dinb(n1567), .dout(n1575));
  jxor g01320(.dina(n1575), .dinb(n1351), .dout(n1576));
  jxor g01321(.dina(n1576), .dinb(n1565), .dout(n1577));
  jnot g01322(.din(n1577), .dout(n1578));
  jor  g01323(.dina(n1248), .dinb(n412), .dout(n1579));
  jor  g01324(.dina(n1251), .dinb(n377), .dout(n1580));
  jor  g01325(.dina(n1147), .dinb(n340), .dout(n1581));
  jand g01326(.dina(n1581), .dinb(n1580), .dout(n1582));
  jor  g01327(.dina(n1246), .dinb(n415), .dout(n1583));
  jand g01328(.dina(n1583), .dinb(n1582), .dout(n1584));
  jand g01329(.dina(n1584), .dinb(n1579), .dout(n1585));
  jxor g01330(.dina(n1585), .dinb(a17 ), .dout(n1586));
  jxor g01331(.dina(n1586), .dinb(n1578), .dout(n1587));
  jxor g01332(.dina(n1587), .dinb(n1560), .dout(n1588));
  jor  g01333(.dina(n970), .dinb(n570), .dout(n1589));
  jor  g01334(.dina(n880), .dinb(n469), .dout(n1590));
  jor  g01335(.dina(n967), .dinb(n519), .dout(n1591));
  jor  g01336(.dina(n972), .dinb(n572), .dout(n1592));
  jand g01337(.dina(n1592), .dinb(n1591), .dout(n1593));
  jand g01338(.dina(n1593), .dinb(n1590), .dout(n1594));
  jand g01339(.dina(n1594), .dinb(n1589), .dout(n1595));
  jxor g01340(.dina(n1595), .dinb(n810), .dout(n1596));
  jxor g01341(.dina(n1596), .dinb(n1588), .dout(n1597));
  jxor g01342(.dina(n1597), .dinb(n1555), .dout(n1598));
  jor  g01343(.dina(n770), .dinb(n728), .dout(n1599));
  jor  g01344(.dina(n660), .dinb(n637), .dout(n1600));
  jor  g01345(.dina(n726), .dinb(n772), .dout(n1601));
  jor  g01346(.dina(n731), .dinb(n704), .dout(n1602));
  jand g01347(.dina(n1602), .dinb(n1601), .dout(n1603));
  jand g01348(.dina(n1603), .dinb(n1600), .dout(n1604));
  jand g01349(.dina(n1604), .dinb(n1599), .dout(n1605));
  jxor g01350(.dina(n1605), .dinb(n606), .dout(n1606));
  jxor g01351(.dina(n1606), .dinb(n1598), .dout(n1607));
  jnot g01352(.din(n1607), .dout(n1608));
  jxor g01353(.dina(n1608), .dinb(n1552), .dout(n1609));
  jor  g01354(.dina(n1016), .dinb(n544), .dout(n1610));
  jor  g01355(.dina(n486), .dinb(n852), .dout(n1611));
  jor  g01356(.dina(n547), .dinb(n934), .dout(n1612));
  jor  g01357(.dina(n542), .dinb(n1018), .dout(n1613));
  jand g01358(.dina(n1613), .dinb(n1612), .dout(n1614));
  jand g01359(.dina(n1614), .dinb(n1611), .dout(n1615));
  jand g01360(.dina(n1615), .dinb(n1610), .dout(n1616));
  jxor g01361(.dina(n1616), .dinb(n446), .dout(n1617));
  jxor g01362(.dina(n1617), .dinb(n1609), .dout(n1618));
  jxor g01363(.dina(n1618), .dinb(n1548), .dout(n1619));
  jor  g01364(.dina(n1305), .dinb(n397), .dout(n1620));
  jor  g01365(.dina(n354), .dinb(n1114), .dout(n1621));
  jor  g01366(.dina(n394), .dinb(n1211), .dout(n1622));
  jor  g01367(.dina(n399), .dinb(n1307), .dout(n1623));
  jand g01368(.dina(n1623), .dinb(n1622), .dout(n1624));
  jand g01369(.dina(n1624), .dinb(n1621), .dout(n1625));
  jand g01370(.dina(n1625), .dinb(n1620), .dout(n1626));
  jxor g01371(.dina(n1626), .dinb(n364), .dout(n1627));
  jxor g01372(.dina(n1627), .dinb(n1619), .dout(n1628));
  jxor g01373(.dina(n1628), .dinb(n1545), .dout(n1629));
  jand g01374(.dina(b20 ), .dinb(b19 ), .dout(n1630));
  jand g01375(.dina(n1523), .dinb(n1522), .dout(n1631));
  jor  g01376(.dina(n1631), .dinb(n1630), .dout(n1632));
  jxor g01377(.dina(b21 ), .dinb(b20 ), .dout(n1633));
  jnot g01378(.din(n1633), .dout(n1634));
  jxor g01379(.dina(n1634), .dinb(n1632), .dout(n1635));
  jor  g01380(.dina(n1635), .dinb(n296), .dout(n1636));
  jnot g01381(.din(b21 ), .dout(n1637));
  jor  g01382(.dina(n264), .dinb(n1637), .dout(n1638));
  jor  g01383(.dina(n294), .dinb(n1527), .dout(n1639));
  jor  g01384(.dina(n280), .dinb(n1416), .dout(n1640));
  jand g01385(.dina(n1640), .dinb(n1639), .dout(n1641));
  jand g01386(.dina(n1641), .dinb(n1638), .dout(n1642));
  jand g01387(.dina(n1642), .dinb(n1636), .dout(n1643));
  jxor g01388(.dina(n1643), .dinb(n278), .dout(n1644));
  jxor g01389(.dina(n1644), .dinb(n1629), .dout(n1645));
  jxor g01390(.dina(n1645), .dinb(n1540), .dout(f21 ));
  jnot g01391(.din(n1644), .dout(n1647));
  jor  g01392(.dina(n1647), .dinb(n1629), .dout(n1648));
  jor  g01393(.dina(n1645), .dinb(n1540), .dout(n1649));
  jand g01394(.dina(n1649), .dinb(n1648), .dout(n1650));
  jand g01395(.dina(n1627), .dinb(n1619), .dout(n1651));
  jnot g01396(.din(n1651), .dout(n1652));
  jnot g01397(.din(n1628), .dout(n1653));
  jor  g01398(.dina(n1653), .dinb(n1545), .dout(n1654));
  jand g01399(.dina(n1654), .dinb(n1652), .dout(n1655));
  jand g01400(.dina(n1617), .dinb(n1609), .dout(n1656));
  jand g01401(.dina(n1618), .dinb(n1548), .dout(n1657));
  jor  g01402(.dina(n1657), .dinb(n1656), .dout(n1658));
  jand g01403(.dina(n1606), .dinb(n1598), .dout(n1659));
  jnot g01404(.din(n1659), .dout(n1660));
  jor  g01405(.dina(n1608), .dinb(n1552), .dout(n1661));
  jand g01406(.dina(n1661), .dinb(n1660), .dout(n1662));
  jand g01407(.dina(n1596), .dinb(n1588), .dout(n1663));
  jand g01408(.dina(n1597), .dinb(n1555), .dout(n1664));
  jor  g01409(.dina(n1664), .dinb(n1663), .dout(n1665));
  jor  g01410(.dina(n1586), .dinb(n1578), .dout(n1666));
  jand g01411(.dina(n1587), .dinb(n1560), .dout(n1667));
  jnot g01412(.din(n1667), .dout(n1668));
  jand g01413(.dina(n1668), .dinb(n1666), .dout(n1669));
  jnot g01414(.din(n1669), .dout(n1670));
  jnot g01415(.din(n1561), .dout(n1671));
  jand g01416(.dina(n1563), .dinb(n1671), .dout(n1672));
  jand g01417(.dina(n1576), .dinb(n1565), .dout(n1673));
  jor  g01418(.dina(n1673), .dinb(n1672), .dout(n1674));
  jxor g01419(.dina(a23 ), .dinb(a22 ), .dout(n1675));
  jand g01420(.dina(n1675), .dinb(n1562), .dout(n1676));
  jand g01421(.dina(n1676), .dinb(n259), .dout(n1677));
  jnot g01422(.din(n1562), .dout(n1678));
  jxor g01423(.dina(a22 ), .dinb(a21 ), .dout(n1679));
  jand g01424(.dina(n1679), .dinb(n1678), .dout(n1680));
  jand g01425(.dina(n1680), .dinb(b0 ), .dout(n1681));
  jnot g01426(.din(n1675), .dout(n1682));
  jand g01427(.dina(n1682), .dinb(n1562), .dout(n1683));
  jand g01428(.dina(n1683), .dinb(b1 ), .dout(n1684));
  jor  g01429(.dina(n1684), .dinb(n1681), .dout(n1685));
  jor  g01430(.dina(n1685), .dinb(n1677), .dout(n1686));
  jnot g01431(.din(a23 ), .dout(n1687));
  jor  g01432(.dina(n1564), .dinb(n1687), .dout(n1688));
  jxor g01433(.dina(n1688), .dinb(n1686), .dout(n1689));
  jor  g01434(.dina(n1569), .dinb(n337), .dout(n1690));
  jor  g01435(.dina(n1571), .dinb(n340), .dout(n1691));
  jor  g01436(.dina(n1453), .dinb(n293), .dout(n1692));
  jand g01437(.dina(n1692), .dinb(n1691), .dout(n1693));
  jor  g01438(.dina(n1566), .dinb(n303), .dout(n1694));
  jand g01439(.dina(n1694), .dinb(n1693), .dout(n1695));
  jand g01440(.dina(n1695), .dinb(n1690), .dout(n1696));
  jxor g01441(.dina(n1696), .dinb(a20 ), .dout(n1697));
  jxor g01442(.dina(n1697), .dinb(n1689), .dout(n1698));
  jxor g01443(.dina(n1698), .dinb(n1674), .dout(n1699));
  jnot g01444(.din(n1699), .dout(n1700));
  jor  g01445(.dina(n1248), .dinb(n466), .dout(n1701));
  jor  g01446(.dina(n1246), .dinb(n469), .dout(n1702));
  jor  g01447(.dina(n1147), .dinb(n377), .dout(n1703));
  jand g01448(.dina(n1703), .dinb(n1702), .dout(n1704));
  jor  g01449(.dina(n1251), .dinb(n415), .dout(n1705));
  jand g01450(.dina(n1705), .dinb(n1704), .dout(n1706));
  jand g01451(.dina(n1706), .dinb(n1701), .dout(n1707));
  jxor g01452(.dina(n1707), .dinb(a17 ), .dout(n1708));
  jxor g01453(.dina(n1708), .dinb(n1700), .dout(n1709));
  jxor g01454(.dina(n1709), .dinb(n1670), .dout(n1710));
  jor  g01455(.dina(n970), .dinb(n635), .dout(n1711));
  jor  g01456(.dina(n880), .dinb(n519), .dout(n1712));
  jor  g01457(.dina(n972), .dinb(n637), .dout(n1713));
  jor  g01458(.dina(n967), .dinb(n572), .dout(n1714));
  jand g01459(.dina(n1714), .dinb(n1713), .dout(n1715));
  jand g01460(.dina(n1715), .dinb(n1712), .dout(n1716));
  jand g01461(.dina(n1716), .dinb(n1711), .dout(n1717));
  jxor g01462(.dina(n1717), .dinb(n810), .dout(n1718));
  jxor g01463(.dina(n1718), .dinb(n1710), .dout(n1719));
  jxor g01464(.dina(n1719), .dinb(n1665), .dout(n1720));
  jor  g01465(.dina(n850), .dinb(n728), .dout(n1721));
  jor  g01466(.dina(n660), .dinb(n704), .dout(n1722));
  jor  g01467(.dina(n726), .dinb(n852), .dout(n1723));
  jor  g01468(.dina(n731), .dinb(n772), .dout(n1724));
  jand g01469(.dina(n1724), .dinb(n1723), .dout(n1725));
  jand g01470(.dina(n1725), .dinb(n1722), .dout(n1726));
  jand g01471(.dina(n1726), .dinb(n1721), .dout(n1727));
  jxor g01472(.dina(n1727), .dinb(n606), .dout(n1728));
  jxor g01473(.dina(n1728), .dinb(n1720), .dout(n1729));
  jnot g01474(.din(n1729), .dout(n1730));
  jxor g01475(.dina(n1730), .dinb(n1662), .dout(n1731));
  jor  g01476(.dina(n1112), .dinb(n544), .dout(n1732));
  jor  g01477(.dina(n486), .dinb(n934), .dout(n1733));
  jor  g01478(.dina(n547), .dinb(n1018), .dout(n1734));
  jor  g01479(.dina(n542), .dinb(n1114), .dout(n1735));
  jand g01480(.dina(n1735), .dinb(n1734), .dout(n1736));
  jand g01481(.dina(n1736), .dinb(n1733), .dout(n1737));
  jand g01482(.dina(n1737), .dinb(n1732), .dout(n1738));
  jxor g01483(.dina(n1738), .dinb(n446), .dout(n1739));
  jxor g01484(.dina(n1739), .dinb(n1731), .dout(n1740));
  jxor g01485(.dina(n1740), .dinb(n1658), .dout(n1741));
  jor  g01486(.dina(n1414), .dinb(n397), .dout(n1742));
  jor  g01487(.dina(n354), .dinb(n1211), .dout(n1743));
  jor  g01488(.dina(n394), .dinb(n1307), .dout(n1744));
  jor  g01489(.dina(n399), .dinb(n1416), .dout(n1745));
  jand g01490(.dina(n1745), .dinb(n1744), .dout(n1746));
  jand g01491(.dina(n1746), .dinb(n1743), .dout(n1747));
  jand g01492(.dina(n1747), .dinb(n1742), .dout(n1748));
  jxor g01493(.dina(n1748), .dinb(n364), .dout(n1749));
  jxor g01494(.dina(n1749), .dinb(n1741), .dout(n1750));
  jxor g01495(.dina(n1750), .dinb(n1655), .dout(n1751));
  jand g01496(.dina(b21 ), .dinb(b20 ), .dout(n1752));
  jand g01497(.dina(n1633), .dinb(n1632), .dout(n1753));
  jor  g01498(.dina(n1753), .dinb(n1752), .dout(n1754));
  jxor g01499(.dina(b22 ), .dinb(b21 ), .dout(n1755));
  jnot g01500(.din(n1755), .dout(n1756));
  jxor g01501(.dina(n1756), .dinb(n1754), .dout(n1757));
  jor  g01502(.dina(n1757), .dinb(n296), .dout(n1758));
  jnot g01503(.din(b22 ), .dout(n1759));
  jor  g01504(.dina(n264), .dinb(n1759), .dout(n1760));
  jor  g01505(.dina(n294), .dinb(n1637), .dout(n1761));
  jor  g01506(.dina(n280), .dinb(n1527), .dout(n1762));
  jand g01507(.dina(n1762), .dinb(n1761), .dout(n1763));
  jand g01508(.dina(n1763), .dinb(n1760), .dout(n1764));
  jand g01509(.dina(n1764), .dinb(n1758), .dout(n1765));
  jxor g01510(.dina(n1765), .dinb(n278), .dout(n1766));
  jxor g01511(.dina(n1766), .dinb(n1751), .dout(n1767));
  jxor g01512(.dina(n1767), .dinb(n1650), .dout(f22 ));
  jnot g01513(.din(n1766), .dout(n1769));
  jor  g01514(.dina(n1769), .dinb(n1751), .dout(n1770));
  jor  g01515(.dina(n1767), .dinb(n1650), .dout(n1771));
  jand g01516(.dina(n1771), .dinb(n1770), .dout(n1772));
  jand g01517(.dina(n1749), .dinb(n1741), .dout(n1773));
  jnot g01518(.din(n1773), .dout(n1774));
  jnot g01519(.din(n1750), .dout(n1775));
  jor  g01520(.dina(n1775), .dinb(n1655), .dout(n1776));
  jand g01521(.dina(n1776), .dinb(n1774), .dout(n1777));
  jand g01522(.dina(n1739), .dinb(n1731), .dout(n1778));
  jand g01523(.dina(n1740), .dinb(n1658), .dout(n1779));
  jor  g01524(.dina(n1779), .dinb(n1778), .dout(n1780));
  jand g01525(.dina(n1728), .dinb(n1720), .dout(n1781));
  jnot g01526(.din(n1781), .dout(n1782));
  jor  g01527(.dina(n1730), .dinb(n1662), .dout(n1783));
  jand g01528(.dina(n1783), .dinb(n1782), .dout(n1784));
  jand g01529(.dina(n1718), .dinb(n1710), .dout(n1785));
  jand g01530(.dina(n1719), .dinb(n1665), .dout(n1786));
  jor  g01531(.dina(n1786), .dinb(n1785), .dout(n1787));
  jor  g01532(.dina(n1708), .dinb(n1700), .dout(n1788));
  jand g01533(.dina(n1709), .dinb(n1670), .dout(n1789));
  jnot g01534(.din(n1789), .dout(n1790));
  jand g01535(.dina(n1790), .dinb(n1788), .dout(n1791));
  jnot g01536(.din(n1791), .dout(n1792));
  jor  g01537(.dina(n1248), .dinb(n517), .dout(n1793));
  jor  g01538(.dina(n1246), .dinb(n519), .dout(n1794));
  jor  g01539(.dina(n1251), .dinb(n469), .dout(n1795));
  jor  g01540(.dina(n1147), .dinb(n415), .dout(n1796));
  jand g01541(.dina(n1796), .dinb(n1795), .dout(n1797));
  jand g01542(.dina(n1797), .dinb(n1794), .dout(n1798));
  jand g01543(.dina(n1798), .dinb(n1793), .dout(n1799));
  jxor g01544(.dina(n1799), .dinb(n1061), .dout(n1800));
  jor  g01545(.dina(n1697), .dinb(n1689), .dout(n1801));
  jand g01546(.dina(n1698), .dinb(n1674), .dout(n1802));
  jnot g01547(.din(n1802), .dout(n1803));
  jand g01548(.dina(n1803), .dinb(n1801), .dout(n1804));
  jor  g01549(.dina(n1679), .dinb(n1562), .dout(n1805));
  jor  g01550(.dina(n1805), .dinb(n1682), .dout(n1806));
  jnot g01551(.din(n1806), .dout(n1807));
  jand g01552(.dina(n1807), .dinb(b0 ), .dout(n1808));
  jand g01553(.dina(n1680), .dinb(b1 ), .dout(n1809));
  jor  g01554(.dina(n1809), .dinb(n1808), .dout(n1810));
  jand g01555(.dina(n1676), .dinb(n273), .dout(n1811));
  jand g01556(.dina(n1683), .dinb(b2 ), .dout(n1812));
  jor  g01557(.dina(n1812), .dinb(n1811), .dout(n1813));
  jor  g01558(.dina(n1813), .dinb(n1810), .dout(n1814));
  jnot g01559(.din(n1686), .dout(n1815));
  jand g01560(.dina(n1564), .dinb(a23 ), .dout(n1816));
  jand g01561(.dina(n1816), .dinb(n1815), .dout(n1817));
  jnot g01562(.din(n1817), .dout(n1818));
  jand g01563(.dina(n1818), .dinb(a23 ), .dout(n1819));
  jxor g01564(.dina(n1819), .dinb(n1814), .dout(n1820));
  jor  g01565(.dina(n1569), .dinb(n374), .dout(n1821));
  jor  g01566(.dina(n1566), .dinb(n340), .dout(n1822));
  jor  g01567(.dina(n1453), .dinb(n303), .dout(n1823));
  jand g01568(.dina(n1823), .dinb(n1822), .dout(n1824));
  jor  g01569(.dina(n1571), .dinb(n377), .dout(n1825));
  jand g01570(.dina(n1825), .dinb(n1824), .dout(n1826));
  jand g01571(.dina(n1826), .dinb(n1821), .dout(n1827));
  jxor g01572(.dina(n1827), .dinb(a20 ), .dout(n1828));
  jxor g01573(.dina(n1828), .dinb(n1820), .dout(n1829));
  jxor g01574(.dina(n1829), .dinb(n1804), .dout(n1830));
  jxor g01575(.dina(n1830), .dinb(n1800), .dout(n1831));
  jxor g01576(.dina(n1831), .dinb(n1792), .dout(n1832));
  jor  g01577(.dina(n970), .dinb(n702), .dout(n1833));
  jor  g01578(.dina(n880), .dinb(n572), .dout(n1834));
  jor  g01579(.dina(n972), .dinb(n704), .dout(n1835));
  jor  g01580(.dina(n967), .dinb(n637), .dout(n1836));
  jand g01581(.dina(n1836), .dinb(n1835), .dout(n1837));
  jand g01582(.dina(n1837), .dinb(n1834), .dout(n1838));
  jand g01583(.dina(n1838), .dinb(n1833), .dout(n1839));
  jxor g01584(.dina(n1839), .dinb(n810), .dout(n1840));
  jxor g01585(.dina(n1840), .dinb(n1832), .dout(n1841));
  jxor g01586(.dina(n1841), .dinb(n1787), .dout(n1842));
  jor  g01587(.dina(n932), .dinb(n728), .dout(n1843));
  jor  g01588(.dina(n660), .dinb(n772), .dout(n1844));
  jor  g01589(.dina(n726), .dinb(n934), .dout(n1845));
  jor  g01590(.dina(n731), .dinb(n852), .dout(n1846));
  jand g01591(.dina(n1846), .dinb(n1845), .dout(n1847));
  jand g01592(.dina(n1847), .dinb(n1844), .dout(n1848));
  jand g01593(.dina(n1848), .dinb(n1843), .dout(n1849));
  jxor g01594(.dina(n1849), .dinb(n606), .dout(n1850));
  jxor g01595(.dina(n1850), .dinb(n1842), .dout(n1851));
  jnot g01596(.din(n1851), .dout(n1852));
  jxor g01597(.dina(n1852), .dinb(n1784), .dout(n1853));
  jor  g01598(.dina(n1209), .dinb(n544), .dout(n1854));
  jor  g01599(.dina(n486), .dinb(n1018), .dout(n1855));
  jor  g01600(.dina(n547), .dinb(n1114), .dout(n1856));
  jor  g01601(.dina(n542), .dinb(n1211), .dout(n1857));
  jand g01602(.dina(n1857), .dinb(n1856), .dout(n1858));
  jand g01603(.dina(n1858), .dinb(n1855), .dout(n1859));
  jand g01604(.dina(n1859), .dinb(n1854), .dout(n1860));
  jxor g01605(.dina(n1860), .dinb(n446), .dout(n1861));
  jxor g01606(.dina(n1861), .dinb(n1853), .dout(n1862));
  jxor g01607(.dina(n1862), .dinb(n1780), .dout(n1863));
  jor  g01608(.dina(n1525), .dinb(n397), .dout(n1864));
  jor  g01609(.dina(n354), .dinb(n1307), .dout(n1865));
  jor  g01610(.dina(n399), .dinb(n1527), .dout(n1866));
  jor  g01611(.dina(n394), .dinb(n1416), .dout(n1867));
  jand g01612(.dina(n1867), .dinb(n1866), .dout(n1868));
  jand g01613(.dina(n1868), .dinb(n1865), .dout(n1869));
  jand g01614(.dina(n1869), .dinb(n1864), .dout(n1870));
  jxor g01615(.dina(n1870), .dinb(n364), .dout(n1871));
  jxor g01616(.dina(n1871), .dinb(n1863), .dout(n1872));
  jxor g01617(.dina(n1872), .dinb(n1777), .dout(n1873));
  jand g01618(.dina(b22 ), .dinb(b21 ), .dout(n1874));
  jand g01619(.dina(n1755), .dinb(n1754), .dout(n1875));
  jor  g01620(.dina(n1875), .dinb(n1874), .dout(n1876));
  jxor g01621(.dina(b23 ), .dinb(b22 ), .dout(n1877));
  jnot g01622(.din(n1877), .dout(n1878));
  jxor g01623(.dina(n1878), .dinb(n1876), .dout(n1879));
  jor  g01624(.dina(n1879), .dinb(n296), .dout(n1880));
  jnot g01625(.din(b23 ), .dout(n1881));
  jor  g01626(.dina(n264), .dinb(n1881), .dout(n1882));
  jor  g01627(.dina(n294), .dinb(n1759), .dout(n1883));
  jor  g01628(.dina(n280), .dinb(n1637), .dout(n1884));
  jand g01629(.dina(n1884), .dinb(n1883), .dout(n1885));
  jand g01630(.dina(n1885), .dinb(n1882), .dout(n1886));
  jand g01631(.dina(n1886), .dinb(n1880), .dout(n1887));
  jxor g01632(.dina(n1887), .dinb(n278), .dout(n1888));
  jxor g01633(.dina(n1888), .dinb(n1873), .dout(n1889));
  jxor g01634(.dina(n1889), .dinb(n1772), .dout(f23 ));
  jnot g01635(.din(n1888), .dout(n1891));
  jor  g01636(.dina(n1891), .dinb(n1873), .dout(n1892));
  jor  g01637(.dina(n1889), .dinb(n1772), .dout(n1893));
  jand g01638(.dina(n1893), .dinb(n1892), .dout(n1894));
  jand g01639(.dina(n1871), .dinb(n1863), .dout(n1895));
  jnot g01640(.din(n1895), .dout(n1896));
  jnot g01641(.din(n1872), .dout(n1897));
  jor  g01642(.dina(n1897), .dinb(n1777), .dout(n1898));
  jand g01643(.dina(n1898), .dinb(n1896), .dout(n1899));
  jand g01644(.dina(n1861), .dinb(n1853), .dout(n1900));
  jand g01645(.dina(n1862), .dinb(n1780), .dout(n1901));
  jor  g01646(.dina(n1901), .dinb(n1900), .dout(n1902));
  jand g01647(.dina(n1850), .dinb(n1842), .dout(n1903));
  jnot g01648(.din(n1903), .dout(n1904));
  jor  g01649(.dina(n1852), .dinb(n1784), .dout(n1905));
  jand g01650(.dina(n1905), .dinb(n1904), .dout(n1906));
  jand g01651(.dina(n1840), .dinb(n1832), .dout(n1907));
  jand g01652(.dina(n1841), .dinb(n1787), .dout(n1908));
  jor  g01653(.dina(n1908), .dinb(n1907), .dout(n1909));
  jand g01654(.dina(n1830), .dinb(n1800), .dout(n1910));
  jand g01655(.dina(n1831), .dinb(n1792), .dout(n1911));
  jor  g01656(.dina(n1911), .dinb(n1910), .dout(n1912));
  jor  g01657(.dina(n1818), .dinb(n1814), .dout(n1913));
  jxor g01658(.dina(a24 ), .dinb(a23 ), .dout(n1914));
  jand g01659(.dina(n1914), .dinb(b0 ), .dout(n1915));
  jnot g01660(.din(n1915), .dout(n1916));
  jxor g01661(.dina(n1916), .dinb(n1913), .dout(n1917));
  jnot g01662(.din(n1680), .dout(n1918));
  jor  g01663(.dina(n1918), .dinb(n293), .dout(n1919));
  jor  g01664(.dina(n1806), .dinb(n305), .dout(n1920));
  jnot g01665(.din(n1676), .dout(n1921));
  jor  g01666(.dina(n1921), .dinb(n301), .dout(n1922));
  jnot g01667(.din(n1683), .dout(n1923));
  jor  g01668(.dina(n1923), .dinb(n303), .dout(n1924));
  jand g01669(.dina(n1924), .dinb(n1922), .dout(n1925));
  jand g01670(.dina(n1925), .dinb(n1920), .dout(n1926));
  jand g01671(.dina(n1926), .dinb(n1919), .dout(n1927));
  jxor g01672(.dina(n1927), .dinb(n1687), .dout(n1928));
  jxor g01673(.dina(n1928), .dinb(n1917), .dout(n1929));
  jnot g01674(.din(n1929), .dout(n1930));
  jor  g01675(.dina(n1569), .dinb(n412), .dout(n1931));
  jor  g01676(.dina(n1571), .dinb(n415), .dout(n1932));
  jor  g01677(.dina(n1453), .dinb(n340), .dout(n1933));
  jand g01678(.dina(n1933), .dinb(n1932), .dout(n1934));
  jor  g01679(.dina(n1566), .dinb(n377), .dout(n1935));
  jand g01680(.dina(n1935), .dinb(n1934), .dout(n1936));
  jand g01681(.dina(n1936), .dinb(n1931), .dout(n1937));
  jxor g01682(.dina(n1937), .dinb(a20 ), .dout(n1938));
  jxor g01683(.dina(n1938), .dinb(n1930), .dout(n1939));
  jnot g01684(.din(n1820), .dout(n1940));
  jand g01685(.dina(n1828), .dinb(n1940), .dout(n1941));
  jnot g01686(.din(n1941), .dout(n1942));
  jnot g01687(.din(n1804), .dout(n1943));
  jnot g01688(.din(n1828), .dout(n1944));
  jand g01689(.dina(n1944), .dinb(n1820), .dout(n1945));
  jor  g01690(.dina(n1945), .dinb(n1943), .dout(n1946));
  jand g01691(.dina(n1946), .dinb(n1942), .dout(n1947));
  jxor g01692(.dina(n1947), .dinb(n1939), .dout(n1948));
  jor  g01693(.dina(n1248), .dinb(n570), .dout(n1949));
  jor  g01694(.dina(n1147), .dinb(n469), .dout(n1950));
  jor  g01695(.dina(n1251), .dinb(n519), .dout(n1951));
  jor  g01696(.dina(n1246), .dinb(n572), .dout(n1952));
  jand g01697(.dina(n1952), .dinb(n1951), .dout(n1953));
  jand g01698(.dina(n1953), .dinb(n1950), .dout(n1954));
  jand g01699(.dina(n1954), .dinb(n1949), .dout(n1955));
  jxor g01700(.dina(n1955), .dinb(n1061), .dout(n1956));
  jxor g01701(.dina(n1956), .dinb(n1948), .dout(n1957));
  jxor g01702(.dina(n1957), .dinb(n1912), .dout(n1958));
  jor  g01703(.dina(n970), .dinb(n770), .dout(n1959));
  jor  g01704(.dina(n880), .dinb(n637), .dout(n1960));
  jor  g01705(.dina(n967), .dinb(n704), .dout(n1961));
  jor  g01706(.dina(n972), .dinb(n772), .dout(n1962));
  jand g01707(.dina(n1962), .dinb(n1961), .dout(n1963));
  jand g01708(.dina(n1963), .dinb(n1960), .dout(n1964));
  jand g01709(.dina(n1964), .dinb(n1959), .dout(n1965));
  jxor g01710(.dina(n1965), .dinb(n810), .dout(n1966));
  jxor g01711(.dina(n1966), .dinb(n1958), .dout(n1967));
  jxor g01712(.dina(n1967), .dinb(n1909), .dout(n1968));
  jor  g01713(.dina(n1016), .dinb(n728), .dout(n1969));
  jor  g01714(.dina(n660), .dinb(n852), .dout(n1970));
  jor  g01715(.dina(n731), .dinb(n934), .dout(n1971));
  jor  g01716(.dina(n726), .dinb(n1018), .dout(n1972));
  jand g01717(.dina(n1972), .dinb(n1971), .dout(n1973));
  jand g01718(.dina(n1973), .dinb(n1970), .dout(n1974));
  jand g01719(.dina(n1974), .dinb(n1969), .dout(n1975));
  jxor g01720(.dina(n1975), .dinb(n606), .dout(n1976));
  jxor g01721(.dina(n1976), .dinb(n1968), .dout(n1977));
  jnot g01722(.din(n1977), .dout(n1978));
  jxor g01723(.dina(n1978), .dinb(n1906), .dout(n1979));
  jor  g01724(.dina(n1305), .dinb(n544), .dout(n1980));
  jor  g01725(.dina(n486), .dinb(n1114), .dout(n1981));
  jor  g01726(.dina(n547), .dinb(n1211), .dout(n1982));
  jor  g01727(.dina(n542), .dinb(n1307), .dout(n1983));
  jand g01728(.dina(n1983), .dinb(n1982), .dout(n1984));
  jand g01729(.dina(n1984), .dinb(n1981), .dout(n1985));
  jand g01730(.dina(n1985), .dinb(n1980), .dout(n1986));
  jxor g01731(.dina(n1986), .dinb(n446), .dout(n1987));
  jxor g01732(.dina(n1987), .dinb(n1979), .dout(n1988));
  jxor g01733(.dina(n1988), .dinb(n1902), .dout(n1989));
  jor  g01734(.dina(n1635), .dinb(n397), .dout(n1990));
  jor  g01735(.dina(n354), .dinb(n1416), .dout(n1991));
  jor  g01736(.dina(n399), .dinb(n1637), .dout(n1992));
  jor  g01737(.dina(n394), .dinb(n1527), .dout(n1993));
  jand g01738(.dina(n1993), .dinb(n1992), .dout(n1994));
  jand g01739(.dina(n1994), .dinb(n1991), .dout(n1995));
  jand g01740(.dina(n1995), .dinb(n1990), .dout(n1996));
  jxor g01741(.dina(n1996), .dinb(n364), .dout(n1997));
  jxor g01742(.dina(n1997), .dinb(n1989), .dout(n1998));
  jxor g01743(.dina(n1998), .dinb(n1899), .dout(n1999));
  jand g01744(.dina(b23 ), .dinb(b22 ), .dout(n2000));
  jand g01745(.dina(n1877), .dinb(n1876), .dout(n2001));
  jor  g01746(.dina(n2001), .dinb(n2000), .dout(n2002));
  jxor g01747(.dina(b24 ), .dinb(b23 ), .dout(n2003));
  jnot g01748(.din(n2003), .dout(n2004));
  jxor g01749(.dina(n2004), .dinb(n2002), .dout(n2005));
  jor  g01750(.dina(n2005), .dinb(n296), .dout(n2006));
  jnot g01751(.din(b24 ), .dout(n2007));
  jor  g01752(.dina(n264), .dinb(n2007), .dout(n2008));
  jor  g01753(.dina(n294), .dinb(n1881), .dout(n2009));
  jor  g01754(.dina(n280), .dinb(n1759), .dout(n2010));
  jand g01755(.dina(n2010), .dinb(n2009), .dout(n2011));
  jand g01756(.dina(n2011), .dinb(n2008), .dout(n2012));
  jand g01757(.dina(n2012), .dinb(n2006), .dout(n2013));
  jxor g01758(.dina(n2013), .dinb(n278), .dout(n2014));
  jxor g01759(.dina(n2014), .dinb(n1999), .dout(n2015));
  jxor g01760(.dina(n2015), .dinb(n1894), .dout(f24 ));
  jnot g01761(.din(n2014), .dout(n2017));
  jor  g01762(.dina(n2017), .dinb(n1999), .dout(n2018));
  jor  g01763(.dina(n2015), .dinb(n1894), .dout(n2019));
  jand g01764(.dina(n2019), .dinb(n2018), .dout(n2020));
  jand g01765(.dina(n1997), .dinb(n1989), .dout(n2021));
  jnot g01766(.din(n2021), .dout(n2022));
  jnot g01767(.din(n1998), .dout(n2023));
  jor  g01768(.dina(n2023), .dinb(n1899), .dout(n2024));
  jand g01769(.dina(n2024), .dinb(n2022), .dout(n2025));
  jand g01770(.dina(n1987), .dinb(n1979), .dout(n2026));
  jand g01771(.dina(n1988), .dinb(n1902), .dout(n2027));
  jor  g01772(.dina(n2027), .dinb(n2026), .dout(n2028));
  jand g01773(.dina(n1976), .dinb(n1968), .dout(n2029));
  jnot g01774(.din(n2029), .dout(n2030));
  jor  g01775(.dina(n1978), .dinb(n1906), .dout(n2031));
  jand g01776(.dina(n2031), .dinb(n2030), .dout(n2032));
  jand g01777(.dina(n1956), .dinb(n1948), .dout(n2033));
  jand g01778(.dina(n1957), .dinb(n1912), .dout(n2034));
  jor  g01779(.dina(n2034), .dinb(n2033), .dout(n2035));
  jor  g01780(.dina(n1938), .dinb(n1930), .dout(n2036));
  jand g01781(.dina(n1947), .dinb(n1939), .dout(n2037));
  jnot g01782(.din(n2037), .dout(n2038));
  jand g01783(.dina(n2038), .dinb(n2036), .dout(n2039));
  jnot g01784(.din(n2039), .dout(n2040));
  jnot g01785(.din(n1913), .dout(n2041));
  jand g01786(.dina(n1915), .dinb(n2041), .dout(n2042));
  jand g01787(.dina(n1928), .dinb(n1917), .dout(n2043));
  jor  g01788(.dina(n2043), .dinb(n2042), .dout(n2044));
  jxor g01789(.dina(a26 ), .dinb(a25 ), .dout(n2045));
  jnot g01790(.din(n2045), .dout(n2046));
  jand g01791(.dina(n2046), .dinb(n1914), .dout(n2047));
  jand g01792(.dina(n2047), .dinb(b1 ), .dout(n2048));
  jand g01793(.dina(n2045), .dinb(n1914), .dout(n2049));
  jand g01794(.dina(n2049), .dinb(n259), .dout(n2050));
  jnot g01795(.din(n1914), .dout(n2051));
  jxor g01796(.dina(a25 ), .dinb(a24 ), .dout(n2052));
  jand g01797(.dina(n2052), .dinb(n2051), .dout(n2053));
  jand g01798(.dina(n2053), .dinb(b0 ), .dout(n2054));
  jor  g01799(.dina(n2054), .dinb(n2050), .dout(n2055));
  jor  g01800(.dina(n2055), .dinb(n2048), .dout(n2056));
  jnot g01801(.din(a26 ), .dout(n2057));
  jor  g01802(.dina(n1916), .dinb(n2057), .dout(n2058));
  jxor g01803(.dina(n2058), .dinb(n2056), .dout(n2059));
  jor  g01804(.dina(n1921), .dinb(n337), .dout(n2060));
  jor  g01805(.dina(n1923), .dinb(n340), .dout(n2061));
  jor  g01806(.dina(n1806), .dinb(n293), .dout(n2062));
  jand g01807(.dina(n2062), .dinb(n2061), .dout(n2063));
  jor  g01808(.dina(n1918), .dinb(n303), .dout(n2064));
  jand g01809(.dina(n2064), .dinb(n2063), .dout(n2065));
  jand g01810(.dina(n2065), .dinb(n2060), .dout(n2066));
  jxor g01811(.dina(n2066), .dinb(a23 ), .dout(n2067));
  jxor g01812(.dina(n2067), .dinb(n2059), .dout(n2068));
  jxor g01813(.dina(n2068), .dinb(n2044), .dout(n2069));
  jnot g01814(.din(n2069), .dout(n2070));
  jor  g01815(.dina(n1569), .dinb(n466), .dout(n2071));
  jor  g01816(.dina(n1566), .dinb(n415), .dout(n2072));
  jor  g01817(.dina(n1453), .dinb(n377), .dout(n2073));
  jand g01818(.dina(n2073), .dinb(n2072), .dout(n2074));
  jor  g01819(.dina(n1571), .dinb(n469), .dout(n2075));
  jand g01820(.dina(n2075), .dinb(n2074), .dout(n2076));
  jand g01821(.dina(n2076), .dinb(n2071), .dout(n2077));
  jxor g01822(.dina(n2077), .dinb(a20 ), .dout(n2078));
  jxor g01823(.dina(n2078), .dinb(n2070), .dout(n2079));
  jxor g01824(.dina(n2079), .dinb(n2040), .dout(n2080));
  jor  g01825(.dina(n1248), .dinb(n635), .dout(n2081));
  jor  g01826(.dina(n1147), .dinb(n519), .dout(n2082));
  jor  g01827(.dina(n1246), .dinb(n637), .dout(n2083));
  jor  g01828(.dina(n1251), .dinb(n572), .dout(n2084));
  jand g01829(.dina(n2084), .dinb(n2083), .dout(n2085));
  jand g01830(.dina(n2085), .dinb(n2082), .dout(n2086));
  jand g01831(.dina(n2086), .dinb(n2081), .dout(n2087));
  jxor g01832(.dina(n2087), .dinb(n1061), .dout(n2088));
  jxor g01833(.dina(n2088), .dinb(n2080), .dout(n2089));
  jxor g01834(.dina(n2089), .dinb(n2035), .dout(n2090));
  jor  g01835(.dina(n850), .dinb(n970), .dout(n2091));
  jor  g01836(.dina(n880), .dinb(n704), .dout(n2092));
  jor  g01837(.dina(n967), .dinb(n772), .dout(n2093));
  jor  g01838(.dina(n972), .dinb(n852), .dout(n2094));
  jand g01839(.dina(n2094), .dinb(n2093), .dout(n2095));
  jand g01840(.dina(n2095), .dinb(n2092), .dout(n2096));
  jand g01841(.dina(n2096), .dinb(n2091), .dout(n2097));
  jxor g01842(.dina(n2097), .dinb(n810), .dout(n2098));
  jxor g01843(.dina(n2098), .dinb(n2090), .dout(n2099));
  jand g01844(.dina(n1966), .dinb(n1958), .dout(n2100));
  jand g01845(.dina(n1967), .dinb(n1909), .dout(n2101));
  jor  g01846(.dina(n2101), .dinb(n2100), .dout(n2102));
  jxor g01847(.dina(n2102), .dinb(n2099), .dout(n2103));
  jor  g01848(.dina(n1112), .dinb(n728), .dout(n2104));
  jor  g01849(.dina(n660), .dinb(n934), .dout(n2105));
  jor  g01850(.dina(n726), .dinb(n1114), .dout(n2106));
  jor  g01851(.dina(n731), .dinb(n1018), .dout(n2107));
  jand g01852(.dina(n2107), .dinb(n2106), .dout(n2108));
  jand g01853(.dina(n2108), .dinb(n2105), .dout(n2109));
  jand g01854(.dina(n2109), .dinb(n2104), .dout(n2110));
  jxor g01855(.dina(n2110), .dinb(n606), .dout(n2111));
  jxor g01856(.dina(n2111), .dinb(n2103), .dout(n2112));
  jnot g01857(.din(n2112), .dout(n2113));
  jxor g01858(.dina(n2113), .dinb(n2032), .dout(n2114));
  jor  g01859(.dina(n1414), .dinb(n544), .dout(n2115));
  jor  g01860(.dina(n486), .dinb(n1211), .dout(n2116));
  jor  g01861(.dina(n547), .dinb(n1307), .dout(n2117));
  jor  g01862(.dina(n542), .dinb(n1416), .dout(n2118));
  jand g01863(.dina(n2118), .dinb(n2117), .dout(n2119));
  jand g01864(.dina(n2119), .dinb(n2116), .dout(n2120));
  jand g01865(.dina(n2120), .dinb(n2115), .dout(n2121));
  jxor g01866(.dina(n2121), .dinb(n446), .dout(n2122));
  jxor g01867(.dina(n2122), .dinb(n2114), .dout(n2123));
  jxor g01868(.dina(n2123), .dinb(n2028), .dout(n2124));
  jor  g01869(.dina(n1757), .dinb(n397), .dout(n2125));
  jor  g01870(.dina(n354), .dinb(n1527), .dout(n2126));
  jor  g01871(.dina(n399), .dinb(n1759), .dout(n2127));
  jor  g01872(.dina(n394), .dinb(n1637), .dout(n2128));
  jand g01873(.dina(n2128), .dinb(n2127), .dout(n2129));
  jand g01874(.dina(n2129), .dinb(n2126), .dout(n2130));
  jand g01875(.dina(n2130), .dinb(n2125), .dout(n2131));
  jxor g01876(.dina(n2131), .dinb(n364), .dout(n2132));
  jxor g01877(.dina(n2132), .dinb(n2124), .dout(n2133));
  jxor g01878(.dina(n2133), .dinb(n2025), .dout(n2134));
  jand g01879(.dina(b24 ), .dinb(b23 ), .dout(n2135));
  jand g01880(.dina(n2003), .dinb(n2002), .dout(n2136));
  jor  g01881(.dina(n2136), .dinb(n2135), .dout(n2137));
  jxor g01882(.dina(b25 ), .dinb(b24 ), .dout(n2138));
  jnot g01883(.din(n2138), .dout(n2139));
  jxor g01884(.dina(n2139), .dinb(n2137), .dout(n2140));
  jor  g01885(.dina(n2140), .dinb(n296), .dout(n2141));
  jnot g01886(.din(b25 ), .dout(n2142));
  jor  g01887(.dina(n264), .dinb(n2142), .dout(n2143));
  jor  g01888(.dina(n280), .dinb(n1881), .dout(n2144));
  jor  g01889(.dina(n294), .dinb(n2007), .dout(n2145));
  jand g01890(.dina(n2145), .dinb(n2144), .dout(n2146));
  jand g01891(.dina(n2146), .dinb(n2143), .dout(n2147));
  jand g01892(.dina(n2147), .dinb(n2141), .dout(n2148));
  jxor g01893(.dina(n2148), .dinb(n278), .dout(n2149));
  jxor g01894(.dina(n2149), .dinb(n2134), .dout(n2150));
  jxor g01895(.dina(n2150), .dinb(n2020), .dout(f25 ));
  jnot g01896(.din(n2149), .dout(n2152));
  jor  g01897(.dina(n2152), .dinb(n2134), .dout(n2153));
  jor  g01898(.dina(n2150), .dinb(n2020), .dout(n2154));
  jand g01899(.dina(n2154), .dinb(n2153), .dout(n2155));
  jand g01900(.dina(n2132), .dinb(n2124), .dout(n2156));
  jnot g01901(.din(n2156), .dout(n2157));
  jnot g01902(.din(n2133), .dout(n2158));
  jor  g01903(.dina(n2158), .dinb(n2025), .dout(n2159));
  jand g01904(.dina(n2159), .dinb(n2157), .dout(n2160));
  jand g01905(.dina(n2122), .dinb(n2114), .dout(n2161));
  jand g01906(.dina(n2123), .dinb(n2028), .dout(n2162));
  jor  g01907(.dina(n2162), .dinb(n2161), .dout(n2163));
  jand g01908(.dina(n2111), .dinb(n2103), .dout(n2164));
  jnot g01909(.din(n2164), .dout(n2165));
  jor  g01910(.dina(n2113), .dinb(n2032), .dout(n2166));
  jand g01911(.dina(n2166), .dinb(n2165), .dout(n2167));
  jand g01912(.dina(n2098), .dinb(n2090), .dout(n2168));
  jand g01913(.dina(n2102), .dinb(n2099), .dout(n2169));
  jor  g01914(.dina(n2169), .dinb(n2168), .dout(n2170));
  jand g01915(.dina(n2088), .dinb(n2080), .dout(n2171));
  jand g01916(.dina(n2089), .dinb(n2035), .dout(n2172));
  jor  g01917(.dina(n2172), .dinb(n2171), .dout(n2173));
  jor  g01918(.dina(n2078), .dinb(n2070), .dout(n2174));
  jand g01919(.dina(n2079), .dinb(n2040), .dout(n2175));
  jnot g01920(.din(n2175), .dout(n2176));
  jand g01921(.dina(n2176), .dinb(n2174), .dout(n2177));
  jnot g01922(.din(n2177), .dout(n2178));
  jor  g01923(.dina(n2067), .dinb(n2059), .dout(n2179));
  jand g01924(.dina(n2068), .dinb(n2044), .dout(n2180));
  jnot g01925(.din(n2180), .dout(n2181));
  jand g01926(.dina(n2181), .dinb(n2179), .dout(n2182));
  jnot g01927(.din(n2182), .dout(n2183));
  jand g01928(.dina(n2053), .dinb(b1 ), .dout(n2184));
  jor  g01929(.dina(n2052), .dinb(n1914), .dout(n2185));
  jor  g01930(.dina(n2185), .dinb(n2046), .dout(n2186));
  jnot g01931(.din(n2186), .dout(n2187));
  jand g01932(.dina(n2187), .dinb(b0 ), .dout(n2188));
  jand g01933(.dina(n2049), .dinb(n273), .dout(n2189));
  jand g01934(.dina(n2047), .dinb(b2 ), .dout(n2190));
  jor  g01935(.dina(n2190), .dinb(n2189), .dout(n2191));
  jor  g01936(.dina(n2191), .dinb(n2188), .dout(n2192));
  jor  g01937(.dina(n2192), .dinb(n2184), .dout(n2193));
  jnot g01938(.din(n2056), .dout(n2194));
  jand g01939(.dina(n1916), .dinb(a26 ), .dout(n2195));
  jand g01940(.dina(n2195), .dinb(n2194), .dout(n2196));
  jnot g01941(.din(n2196), .dout(n2197));
  jand g01942(.dina(n2197), .dinb(a26 ), .dout(n2198));
  jxor g01943(.dina(n2198), .dinb(n2193), .dout(n2199));
  jnot g01944(.din(n2199), .dout(n2200));
  jor  g01945(.dina(n1921), .dinb(n374), .dout(n2201));
  jor  g01946(.dina(n1923), .dinb(n377), .dout(n2202));
  jor  g01947(.dina(n1806), .dinb(n303), .dout(n2203));
  jand g01948(.dina(n2203), .dinb(n2202), .dout(n2204));
  jor  g01949(.dina(n1918), .dinb(n340), .dout(n2205));
  jand g01950(.dina(n2205), .dinb(n2204), .dout(n2206));
  jand g01951(.dina(n2206), .dinb(n2201), .dout(n2207));
  jxor g01952(.dina(n2207), .dinb(a23 ), .dout(n2208));
  jxor g01953(.dina(n2208), .dinb(n2200), .dout(n2209));
  jxor g01954(.dina(n2209), .dinb(n2183), .dout(n2210));
  jor  g01955(.dina(n1569), .dinb(n517), .dout(n2211));
  jor  g01956(.dina(n1571), .dinb(n519), .dout(n2212));
  jor  g01957(.dina(n1566), .dinb(n469), .dout(n2213));
  jor  g01958(.dina(n1453), .dinb(n415), .dout(n2214));
  jand g01959(.dina(n2214), .dinb(n2213), .dout(n2215));
  jand g01960(.dina(n2215), .dinb(n2212), .dout(n2216));
  jand g01961(.dina(n2216), .dinb(n2211), .dout(n2217));
  jxor g01962(.dina(n2217), .dinb(n1351), .dout(n2218));
  jxor g01963(.dina(n2218), .dinb(n2210), .dout(n2219));
  jxor g01964(.dina(n2219), .dinb(n2178), .dout(n2220));
  jor  g01965(.dina(n1248), .dinb(n702), .dout(n2221));
  jor  g01966(.dina(n1147), .dinb(n572), .dout(n2222));
  jor  g01967(.dina(n1251), .dinb(n637), .dout(n2223));
  jor  g01968(.dina(n1246), .dinb(n704), .dout(n2224));
  jand g01969(.dina(n2224), .dinb(n2223), .dout(n2225));
  jand g01970(.dina(n2225), .dinb(n2222), .dout(n2226));
  jand g01971(.dina(n2226), .dinb(n2221), .dout(n2227));
  jxor g01972(.dina(n2227), .dinb(n1061), .dout(n2228));
  jxor g01973(.dina(n2228), .dinb(n2220), .dout(n2229));
  jxor g01974(.dina(n2229), .dinb(n2173), .dout(n2230));
  jor  g01975(.dina(n932), .dinb(n970), .dout(n2231));
  jor  g01976(.dina(n880), .dinb(n772), .dout(n2232));
  jor  g01977(.dina(n967), .dinb(n852), .dout(n2233));
  jor  g01978(.dina(n972), .dinb(n934), .dout(n2234));
  jand g01979(.dina(n2234), .dinb(n2233), .dout(n2235));
  jand g01980(.dina(n2235), .dinb(n2232), .dout(n2236));
  jand g01981(.dina(n2236), .dinb(n2231), .dout(n2237));
  jxor g01982(.dina(n2237), .dinb(n810), .dout(n2238));
  jxor g01983(.dina(n2238), .dinb(n2230), .dout(n2239));
  jxor g01984(.dina(n2239), .dinb(n2170), .dout(n2240));
  jor  g01985(.dina(n1209), .dinb(n728), .dout(n2241));
  jor  g01986(.dina(n660), .dinb(n1018), .dout(n2242));
  jor  g01987(.dina(n726), .dinb(n1211), .dout(n2243));
  jor  g01988(.dina(n731), .dinb(n1114), .dout(n2244));
  jand g01989(.dina(n2244), .dinb(n2243), .dout(n2245));
  jand g01990(.dina(n2245), .dinb(n2242), .dout(n2246));
  jand g01991(.dina(n2246), .dinb(n2241), .dout(n2247));
  jxor g01992(.dina(n2247), .dinb(n606), .dout(n2248));
  jxor g01993(.dina(n2248), .dinb(n2240), .dout(n2249));
  jnot g01994(.din(n2249), .dout(n2250));
  jxor g01995(.dina(n2250), .dinb(n2167), .dout(n2251));
  jor  g01996(.dina(n1525), .dinb(n544), .dout(n2252));
  jor  g01997(.dina(n486), .dinb(n1307), .dout(n2253));
  jor  g01998(.dina(n547), .dinb(n1416), .dout(n2254));
  jor  g01999(.dina(n542), .dinb(n1527), .dout(n2255));
  jand g02000(.dina(n2255), .dinb(n2254), .dout(n2256));
  jand g02001(.dina(n2256), .dinb(n2253), .dout(n2257));
  jand g02002(.dina(n2257), .dinb(n2252), .dout(n2258));
  jxor g02003(.dina(n2258), .dinb(n446), .dout(n2259));
  jxor g02004(.dina(n2259), .dinb(n2251), .dout(n2260));
  jxor g02005(.dina(n2260), .dinb(n2163), .dout(n2261));
  jor  g02006(.dina(n1879), .dinb(n397), .dout(n2262));
  jor  g02007(.dina(n354), .dinb(n1637), .dout(n2263));
  jor  g02008(.dina(n394), .dinb(n1759), .dout(n2264));
  jor  g02009(.dina(n399), .dinb(n1881), .dout(n2265));
  jand g02010(.dina(n2265), .dinb(n2264), .dout(n2266));
  jand g02011(.dina(n2266), .dinb(n2263), .dout(n2267));
  jand g02012(.dina(n2267), .dinb(n2262), .dout(n2268));
  jxor g02013(.dina(n2268), .dinb(n364), .dout(n2269));
  jxor g02014(.dina(n2269), .dinb(n2261), .dout(n2270));
  jxor g02015(.dina(n2270), .dinb(n2160), .dout(n2271));
  jand g02016(.dina(b25 ), .dinb(b24 ), .dout(n2272));
  jand g02017(.dina(n2138), .dinb(n2137), .dout(n2273));
  jor  g02018(.dina(n2273), .dinb(n2272), .dout(n2274));
  jxor g02019(.dina(b26 ), .dinb(b25 ), .dout(n2275));
  jnot g02020(.din(n2275), .dout(n2276));
  jxor g02021(.dina(n2276), .dinb(n2274), .dout(n2277));
  jor  g02022(.dina(n2277), .dinb(n296), .dout(n2278));
  jnot g02023(.din(b26 ), .dout(n2279));
  jor  g02024(.dina(n264), .dinb(n2279), .dout(n2280));
  jor  g02025(.dina(n294), .dinb(n2142), .dout(n2281));
  jor  g02026(.dina(n280), .dinb(n2007), .dout(n2282));
  jand g02027(.dina(n2282), .dinb(n2281), .dout(n2283));
  jand g02028(.dina(n2283), .dinb(n2280), .dout(n2284));
  jand g02029(.dina(n2284), .dinb(n2278), .dout(n2285));
  jxor g02030(.dina(n2285), .dinb(n278), .dout(n2286));
  jxor g02031(.dina(n2286), .dinb(n2271), .dout(n2287));
  jxor g02032(.dina(n2287), .dinb(n2155), .dout(f26 ));
  jnot g02033(.din(n2286), .dout(n2289));
  jor  g02034(.dina(n2289), .dinb(n2271), .dout(n2290));
  jor  g02035(.dina(n2287), .dinb(n2155), .dout(n2291));
  jand g02036(.dina(n2291), .dinb(n2290), .dout(n2292));
  jand g02037(.dina(n2269), .dinb(n2261), .dout(n2293));
  jnot g02038(.din(n2293), .dout(n2294));
  jnot g02039(.din(n2270), .dout(n2295));
  jor  g02040(.dina(n2295), .dinb(n2160), .dout(n2296));
  jand g02041(.dina(n2296), .dinb(n2294), .dout(n2297));
  jand g02042(.dina(n2248), .dinb(n2240), .dout(n2298));
  jnot g02043(.din(n2298), .dout(n2299));
  jor  g02044(.dina(n2250), .dinb(n2167), .dout(n2300));
  jand g02045(.dina(n2300), .dinb(n2299), .dout(n2301));
  jand g02046(.dina(n2238), .dinb(n2230), .dout(n2302));
  jand g02047(.dina(n2239), .dinb(n2170), .dout(n2303));
  jor  g02048(.dina(n2303), .dinb(n2302), .dout(n2304));
  jand g02049(.dina(n2228), .dinb(n2220), .dout(n2305));
  jand g02050(.dina(n2229), .dinb(n2173), .dout(n2306));
  jor  g02051(.dina(n2306), .dinb(n2305), .dout(n2307));
  jand g02052(.dina(n2218), .dinb(n2210), .dout(n2308));
  jand g02053(.dina(n2219), .dinb(n2178), .dout(n2309));
  jor  g02054(.dina(n2309), .dinb(n2308), .dout(n2310));
  jor  g02055(.dina(n2208), .dinb(n2200), .dout(n2311));
  jand g02056(.dina(n2209), .dinb(n2183), .dout(n2312));
  jnot g02057(.din(n2312), .dout(n2313));
  jand g02058(.dina(n2313), .dinb(n2311), .dout(n2314));
  jnot g02059(.din(n2314), .dout(n2315));
  jor  g02060(.dina(n2197), .dinb(n2193), .dout(n2316));
  jxor g02061(.dina(a27 ), .dinb(a26 ), .dout(n2317));
  jand g02062(.dina(n2317), .dinb(b0 ), .dout(n2318));
  jnot g02063(.din(n2318), .dout(n2319));
  jxor g02064(.dina(n2319), .dinb(n2316), .dout(n2320));
  jnot g02065(.din(n2053), .dout(n2321));
  jor  g02066(.dina(n2321), .dinb(n293), .dout(n2322));
  jor  g02067(.dina(n2186), .dinb(n305), .dout(n2323));
  jnot g02068(.din(n2049), .dout(n2324));
  jor  g02069(.dina(n2324), .dinb(n301), .dout(n2325));
  jnot g02070(.din(n2047), .dout(n2326));
  jor  g02071(.dina(n2326), .dinb(n303), .dout(n2327));
  jand g02072(.dina(n2327), .dinb(n2325), .dout(n2328));
  jand g02073(.dina(n2328), .dinb(n2323), .dout(n2329));
  jand g02074(.dina(n2329), .dinb(n2322), .dout(n2330));
  jxor g02075(.dina(n2330), .dinb(n2057), .dout(n2331));
  jxor g02076(.dina(n2331), .dinb(n2320), .dout(n2332));
  jnot g02077(.din(n2332), .dout(n2333));
  jor  g02078(.dina(n1921), .dinb(n412), .dout(n2334));
  jor  g02079(.dina(n1918), .dinb(n377), .dout(n2335));
  jor  g02080(.dina(n1806), .dinb(n340), .dout(n2336));
  jand g02081(.dina(n2336), .dinb(n2335), .dout(n2337));
  jor  g02082(.dina(n1923), .dinb(n415), .dout(n2338));
  jand g02083(.dina(n2338), .dinb(n2337), .dout(n2339));
  jand g02084(.dina(n2339), .dinb(n2334), .dout(n2340));
  jxor g02085(.dina(n2340), .dinb(a23 ), .dout(n2341));
  jxor g02086(.dina(n2341), .dinb(n2333), .dout(n2342));
  jxor g02087(.dina(n2342), .dinb(n2315), .dout(n2343));
  jor  g02088(.dina(n1569), .dinb(n570), .dout(n2344));
  jor  g02089(.dina(n1453), .dinb(n469), .dout(n2345));
  jor  g02090(.dina(n1566), .dinb(n519), .dout(n2346));
  jor  g02091(.dina(n1571), .dinb(n572), .dout(n2347));
  jand g02092(.dina(n2347), .dinb(n2346), .dout(n2348));
  jand g02093(.dina(n2348), .dinb(n2345), .dout(n2349));
  jand g02094(.dina(n2349), .dinb(n2344), .dout(n2350));
  jxor g02095(.dina(n2350), .dinb(n1351), .dout(n2351));
  jxor g02096(.dina(n2351), .dinb(n2343), .dout(n2352));
  jxor g02097(.dina(n2352), .dinb(n2310), .dout(n2353));
  jor  g02098(.dina(n1248), .dinb(n770), .dout(n2354));
  jor  g02099(.dina(n1147), .dinb(n637), .dout(n2355));
  jor  g02100(.dina(n1251), .dinb(n704), .dout(n2356));
  jor  g02101(.dina(n1246), .dinb(n772), .dout(n2357));
  jand g02102(.dina(n2357), .dinb(n2356), .dout(n2358));
  jand g02103(.dina(n2358), .dinb(n2355), .dout(n2359));
  jand g02104(.dina(n2359), .dinb(n2354), .dout(n2360));
  jxor g02105(.dina(n2360), .dinb(n1061), .dout(n2361));
  jxor g02106(.dina(n2361), .dinb(n2353), .dout(n2362));
  jxor g02107(.dina(n2362), .dinb(n2307), .dout(n2363));
  jor  g02108(.dina(n1016), .dinb(n970), .dout(n2364));
  jor  g02109(.dina(n880), .dinb(n852), .dout(n2365));
  jor  g02110(.dina(n972), .dinb(n1018), .dout(n2366));
  jor  g02111(.dina(n967), .dinb(n934), .dout(n2367));
  jand g02112(.dina(n2367), .dinb(n2366), .dout(n2368));
  jand g02113(.dina(n2368), .dinb(n2365), .dout(n2369));
  jand g02114(.dina(n2369), .dinb(n2364), .dout(n2370));
  jxor g02115(.dina(n2370), .dinb(n810), .dout(n2371));
  jxor g02116(.dina(n2371), .dinb(n2363), .dout(n2372));
  jxor g02117(.dina(n2372), .dinb(n2304), .dout(n2373));
  jor  g02118(.dina(n1305), .dinb(n728), .dout(n2374));
  jor  g02119(.dina(n660), .dinb(n1114), .dout(n2375));
  jor  g02120(.dina(n726), .dinb(n1307), .dout(n2376));
  jor  g02121(.dina(n731), .dinb(n1211), .dout(n2377));
  jand g02122(.dina(n2377), .dinb(n2376), .dout(n2378));
  jand g02123(.dina(n2378), .dinb(n2375), .dout(n2379));
  jand g02124(.dina(n2379), .dinb(n2374), .dout(n2380));
  jxor g02125(.dina(n2380), .dinb(n606), .dout(n2381));
  jxor g02126(.dina(n2381), .dinb(n2373), .dout(n2382));
  jnot g02127(.din(n2382), .dout(n2383));
  jxor g02128(.dina(n2383), .dinb(n2301), .dout(n2384));
  jor  g02129(.dina(n1635), .dinb(n544), .dout(n2385));
  jor  g02130(.dina(n486), .dinb(n1416), .dout(n2386));
  jor  g02131(.dina(n547), .dinb(n1527), .dout(n2387));
  jor  g02132(.dina(n542), .dinb(n1637), .dout(n2388));
  jand g02133(.dina(n2388), .dinb(n2387), .dout(n2389));
  jand g02134(.dina(n2389), .dinb(n2386), .dout(n2390));
  jand g02135(.dina(n2390), .dinb(n2385), .dout(n2391));
  jxor g02136(.dina(n2391), .dinb(n446), .dout(n2392));
  jxor g02137(.dina(n2392), .dinb(n2384), .dout(n2393));
  jand g02138(.dina(n2259), .dinb(n2251), .dout(n2394));
  jand g02139(.dina(n2260), .dinb(n2163), .dout(n2395));
  jor  g02140(.dina(n2395), .dinb(n2394), .dout(n2396));
  jxor g02141(.dina(n2396), .dinb(n2393), .dout(n2397));
  jor  g02142(.dina(n2005), .dinb(n397), .dout(n2398));
  jor  g02143(.dina(n354), .dinb(n1759), .dout(n2399));
  jor  g02144(.dina(n394), .dinb(n1881), .dout(n2400));
  jor  g02145(.dina(n399), .dinb(n2007), .dout(n2401));
  jand g02146(.dina(n2401), .dinb(n2400), .dout(n2402));
  jand g02147(.dina(n2402), .dinb(n2399), .dout(n2403));
  jand g02148(.dina(n2403), .dinb(n2398), .dout(n2404));
  jxor g02149(.dina(n2404), .dinb(n364), .dout(n2405));
  jxor g02150(.dina(n2405), .dinb(n2397), .dout(n2406));
  jxor g02151(.dina(n2406), .dinb(n2297), .dout(n2407));
  jand g02152(.dina(b26 ), .dinb(b25 ), .dout(n2408));
  jand g02153(.dina(n2275), .dinb(n2274), .dout(n2409));
  jor  g02154(.dina(n2409), .dinb(n2408), .dout(n2410));
  jxor g02155(.dina(b27 ), .dinb(b26 ), .dout(n2411));
  jnot g02156(.din(n2411), .dout(n2412));
  jxor g02157(.dina(n2412), .dinb(n2410), .dout(n2413));
  jor  g02158(.dina(n2413), .dinb(n296), .dout(n2414));
  jnot g02159(.din(b27 ), .dout(n2415));
  jor  g02160(.dina(n264), .dinb(n2415), .dout(n2416));
  jor  g02161(.dina(n294), .dinb(n2279), .dout(n2417));
  jor  g02162(.dina(n280), .dinb(n2142), .dout(n2418));
  jand g02163(.dina(n2418), .dinb(n2417), .dout(n2419));
  jand g02164(.dina(n2419), .dinb(n2416), .dout(n2420));
  jand g02165(.dina(n2420), .dinb(n2414), .dout(n2421));
  jxor g02166(.dina(n2421), .dinb(n278), .dout(n2422));
  jxor g02167(.dina(n2422), .dinb(n2407), .dout(n2423));
  jxor g02168(.dina(n2423), .dinb(n2292), .dout(f27 ));
  jnot g02169(.din(n2422), .dout(n2425));
  jor  g02170(.dina(n2425), .dinb(n2407), .dout(n2426));
  jor  g02171(.dina(n2423), .dinb(n2292), .dout(n2427));
  jand g02172(.dina(n2427), .dinb(n2426), .dout(n2428));
  jand g02173(.dina(n2405), .dinb(n2397), .dout(n2429));
  jnot g02174(.din(n2429), .dout(n2430));
  jnot g02175(.din(n2406), .dout(n2431));
  jor  g02176(.dina(n2431), .dinb(n2297), .dout(n2432));
  jand g02177(.dina(n2432), .dinb(n2430), .dout(n2433));
  jand g02178(.dina(n2381), .dinb(n2373), .dout(n2434));
  jnot g02179(.din(n2434), .dout(n2435));
  jor  g02180(.dina(n2383), .dinb(n2301), .dout(n2436));
  jand g02181(.dina(n2436), .dinb(n2435), .dout(n2437));
  jand g02182(.dina(n2371), .dinb(n2363), .dout(n2438));
  jand g02183(.dina(n2372), .dinb(n2304), .dout(n2439));
  jor  g02184(.dina(n2439), .dinb(n2438), .dout(n2440));
  jand g02185(.dina(n2361), .dinb(n2353), .dout(n2441));
  jand g02186(.dina(n2362), .dinb(n2307), .dout(n2442));
  jor  g02187(.dina(n2442), .dinb(n2441), .dout(n2443));
  jand g02188(.dina(n2351), .dinb(n2343), .dout(n2444));
  jand g02189(.dina(n2352), .dinb(n2310), .dout(n2445));
  jor  g02190(.dina(n2445), .dinb(n2444), .dout(n2446));
  jor  g02191(.dina(n2341), .dinb(n2333), .dout(n2447));
  jand g02192(.dina(n2342), .dinb(n2315), .dout(n2448));
  jnot g02193(.din(n2448), .dout(n2449));
  jand g02194(.dina(n2449), .dinb(n2447), .dout(n2450));
  jnot g02195(.din(n2450), .dout(n2451));
  jnot g02196(.din(n2316), .dout(n2452));
  jand g02197(.dina(n2318), .dinb(n2452), .dout(n2453));
  jand g02198(.dina(n2331), .dinb(n2320), .dout(n2454));
  jor  g02199(.dina(n2454), .dinb(n2453), .dout(n2455));
  jxor g02200(.dina(a29 ), .dinb(a28 ), .dout(n2456));
  jnot g02201(.din(n2456), .dout(n2457));
  jand g02202(.dina(n2457), .dinb(n2317), .dout(n2458));
  jand g02203(.dina(n2458), .dinb(b1 ), .dout(n2459));
  jand g02204(.dina(n2456), .dinb(n2317), .dout(n2460));
  jand g02205(.dina(n2460), .dinb(n259), .dout(n2461));
  jnot g02206(.din(n2317), .dout(n2462));
  jxor g02207(.dina(a28 ), .dinb(a27 ), .dout(n2463));
  jand g02208(.dina(n2463), .dinb(n2462), .dout(n2464));
  jand g02209(.dina(n2464), .dinb(b0 ), .dout(n2465));
  jor  g02210(.dina(n2465), .dinb(n2461), .dout(n2466));
  jor  g02211(.dina(n2466), .dinb(n2459), .dout(n2467));
  jnot g02212(.din(a29 ), .dout(n2468));
  jor  g02213(.dina(n2319), .dinb(n2468), .dout(n2469));
  jxor g02214(.dina(n2469), .dinb(n2467), .dout(n2470));
  jor  g02215(.dina(n2324), .dinb(n337), .dout(n2471));
  jor  g02216(.dina(n2326), .dinb(n340), .dout(n2472));
  jor  g02217(.dina(n2186), .dinb(n293), .dout(n2473));
  jand g02218(.dina(n2473), .dinb(n2472), .dout(n2474));
  jor  g02219(.dina(n2321), .dinb(n303), .dout(n2475));
  jand g02220(.dina(n2475), .dinb(n2474), .dout(n2476));
  jand g02221(.dina(n2476), .dinb(n2471), .dout(n2477));
  jxor g02222(.dina(n2477), .dinb(a26 ), .dout(n2478));
  jxor g02223(.dina(n2478), .dinb(n2470), .dout(n2479));
  jxor g02224(.dina(n2479), .dinb(n2455), .dout(n2480));
  jnot g02225(.din(n2480), .dout(n2481));
  jor  g02226(.dina(n1921), .dinb(n466), .dout(n2482));
  jor  g02227(.dina(n1923), .dinb(n469), .dout(n2483));
  jor  g02228(.dina(n1806), .dinb(n377), .dout(n2484));
  jand g02229(.dina(n2484), .dinb(n2483), .dout(n2485));
  jor  g02230(.dina(n1918), .dinb(n415), .dout(n2486));
  jand g02231(.dina(n2486), .dinb(n2485), .dout(n2487));
  jand g02232(.dina(n2487), .dinb(n2482), .dout(n2488));
  jxor g02233(.dina(n2488), .dinb(a23 ), .dout(n2489));
  jxor g02234(.dina(n2489), .dinb(n2481), .dout(n2490));
  jxor g02235(.dina(n2490), .dinb(n2451), .dout(n2491));
  jor  g02236(.dina(n1569), .dinb(n635), .dout(n2492));
  jor  g02237(.dina(n1453), .dinb(n519), .dout(n2493));
  jor  g02238(.dina(n1566), .dinb(n572), .dout(n2494));
  jor  g02239(.dina(n1571), .dinb(n637), .dout(n2495));
  jand g02240(.dina(n2495), .dinb(n2494), .dout(n2496));
  jand g02241(.dina(n2496), .dinb(n2493), .dout(n2497));
  jand g02242(.dina(n2497), .dinb(n2492), .dout(n2498));
  jxor g02243(.dina(n2498), .dinb(n1351), .dout(n2499));
  jxor g02244(.dina(n2499), .dinb(n2491), .dout(n2500));
  jxor g02245(.dina(n2500), .dinb(n2446), .dout(n2501));
  jor  g02246(.dina(n1248), .dinb(n850), .dout(n2502));
  jor  g02247(.dina(n1147), .dinb(n704), .dout(n2503));
  jor  g02248(.dina(n1246), .dinb(n852), .dout(n2504));
  jor  g02249(.dina(n1251), .dinb(n772), .dout(n2505));
  jand g02250(.dina(n2505), .dinb(n2504), .dout(n2506));
  jand g02251(.dina(n2506), .dinb(n2503), .dout(n2507));
  jand g02252(.dina(n2507), .dinb(n2502), .dout(n2508));
  jxor g02253(.dina(n2508), .dinb(n1061), .dout(n2509));
  jxor g02254(.dina(n2509), .dinb(n2501), .dout(n2510));
  jxor g02255(.dina(n2510), .dinb(n2443), .dout(n2511));
  jor  g02256(.dina(n1112), .dinb(n970), .dout(n2512));
  jor  g02257(.dina(n880), .dinb(n934), .dout(n2513));
  jor  g02258(.dina(n972), .dinb(n1114), .dout(n2514));
  jor  g02259(.dina(n967), .dinb(n1018), .dout(n2515));
  jand g02260(.dina(n2515), .dinb(n2514), .dout(n2516));
  jand g02261(.dina(n2516), .dinb(n2513), .dout(n2517));
  jand g02262(.dina(n2517), .dinb(n2512), .dout(n2518));
  jxor g02263(.dina(n2518), .dinb(n810), .dout(n2519));
  jxor g02264(.dina(n2519), .dinb(n2511), .dout(n2520));
  jxor g02265(.dina(n2520), .dinb(n2440), .dout(n2521));
  jor  g02266(.dina(n1414), .dinb(n728), .dout(n2522));
  jor  g02267(.dina(n660), .dinb(n1211), .dout(n2523));
  jor  g02268(.dina(n731), .dinb(n1307), .dout(n2524));
  jor  g02269(.dina(n726), .dinb(n1416), .dout(n2525));
  jand g02270(.dina(n2525), .dinb(n2524), .dout(n2526));
  jand g02271(.dina(n2526), .dinb(n2523), .dout(n2527));
  jand g02272(.dina(n2527), .dinb(n2522), .dout(n2528));
  jxor g02273(.dina(n2528), .dinb(n606), .dout(n2529));
  jxor g02274(.dina(n2529), .dinb(n2521), .dout(n2530));
  jnot g02275(.din(n2530), .dout(n2531));
  jxor g02276(.dina(n2531), .dinb(n2437), .dout(n2532));
  jor  g02277(.dina(n1757), .dinb(n544), .dout(n2533));
  jor  g02278(.dina(n486), .dinb(n1527), .dout(n2534));
  jor  g02279(.dina(n542), .dinb(n1759), .dout(n2535));
  jor  g02280(.dina(n547), .dinb(n1637), .dout(n2536));
  jand g02281(.dina(n2536), .dinb(n2535), .dout(n2537));
  jand g02282(.dina(n2537), .dinb(n2534), .dout(n2538));
  jand g02283(.dina(n2538), .dinb(n2533), .dout(n2539));
  jxor g02284(.dina(n2539), .dinb(n446), .dout(n2540));
  jxor g02285(.dina(n2540), .dinb(n2532), .dout(n2541));
  jand g02286(.dina(n2392), .dinb(n2384), .dout(n2542));
  jand g02287(.dina(n2396), .dinb(n2393), .dout(n2543));
  jor  g02288(.dina(n2543), .dinb(n2542), .dout(n2544));
  jxor g02289(.dina(n2544), .dinb(n2541), .dout(n2545));
  jor  g02290(.dina(n2140), .dinb(n397), .dout(n2546));
  jor  g02291(.dina(n354), .dinb(n1881), .dout(n2547));
  jor  g02292(.dina(n394), .dinb(n2007), .dout(n2548));
  jor  g02293(.dina(n399), .dinb(n2142), .dout(n2549));
  jand g02294(.dina(n2549), .dinb(n2548), .dout(n2550));
  jand g02295(.dina(n2550), .dinb(n2547), .dout(n2551));
  jand g02296(.dina(n2551), .dinb(n2546), .dout(n2552));
  jxor g02297(.dina(n2552), .dinb(n364), .dout(n2553));
  jxor g02298(.dina(n2553), .dinb(n2545), .dout(n2554));
  jxor g02299(.dina(n2554), .dinb(n2433), .dout(n2555));
  jand g02300(.dina(b27 ), .dinb(b26 ), .dout(n2556));
  jand g02301(.dina(n2411), .dinb(n2410), .dout(n2557));
  jor  g02302(.dina(n2557), .dinb(n2556), .dout(n2558));
  jxor g02303(.dina(b28 ), .dinb(b27 ), .dout(n2559));
  jnot g02304(.din(n2559), .dout(n2560));
  jxor g02305(.dina(n2560), .dinb(n2558), .dout(n2561));
  jor  g02306(.dina(n2561), .dinb(n296), .dout(n2562));
  jnot g02307(.din(b28 ), .dout(n2563));
  jor  g02308(.dina(n264), .dinb(n2563), .dout(n2564));
  jor  g02309(.dina(n294), .dinb(n2415), .dout(n2565));
  jor  g02310(.dina(n280), .dinb(n2279), .dout(n2566));
  jand g02311(.dina(n2566), .dinb(n2565), .dout(n2567));
  jand g02312(.dina(n2567), .dinb(n2564), .dout(n2568));
  jand g02313(.dina(n2568), .dinb(n2562), .dout(n2569));
  jxor g02314(.dina(n2569), .dinb(n278), .dout(n2570));
  jxor g02315(.dina(n2570), .dinb(n2555), .dout(n2571));
  jxor g02316(.dina(n2571), .dinb(n2428), .dout(f28 ));
  jnot g02317(.din(n2570), .dout(n2573));
  jor  g02318(.dina(n2573), .dinb(n2555), .dout(n2574));
  jor  g02319(.dina(n2571), .dinb(n2428), .dout(n2575));
  jand g02320(.dina(n2575), .dinb(n2574), .dout(n2576));
  jand g02321(.dina(n2553), .dinb(n2545), .dout(n2577));
  jnot g02322(.din(n2577), .dout(n2578));
  jnot g02323(.din(n2554), .dout(n2579));
  jor  g02324(.dina(n2579), .dinb(n2433), .dout(n2580));
  jand g02325(.dina(n2580), .dinb(n2578), .dout(n2581));
  jand g02326(.dina(n2540), .dinb(n2532), .dout(n2582));
  jand g02327(.dina(n2544), .dinb(n2541), .dout(n2583));
  jor  g02328(.dina(n2583), .dinb(n2582), .dout(n2584));
  jand g02329(.dina(n2529), .dinb(n2521), .dout(n2585));
  jnot g02330(.din(n2585), .dout(n2586));
  jor  g02331(.dina(n2531), .dinb(n2437), .dout(n2587));
  jand g02332(.dina(n2587), .dinb(n2586), .dout(n2588));
  jand g02333(.dina(n2519), .dinb(n2511), .dout(n2589));
  jand g02334(.dina(n2520), .dinb(n2440), .dout(n2590));
  jor  g02335(.dina(n2590), .dinb(n2589), .dout(n2591));
  jand g02336(.dina(n2509), .dinb(n2501), .dout(n2592));
  jand g02337(.dina(n2510), .dinb(n2443), .dout(n2593));
  jor  g02338(.dina(n2593), .dinb(n2592), .dout(n2594));
  jand g02339(.dina(n2499), .dinb(n2491), .dout(n2595));
  jand g02340(.dina(n2500), .dinb(n2446), .dout(n2596));
  jor  g02341(.dina(n2596), .dinb(n2595), .dout(n2597));
  jor  g02342(.dina(n2489), .dinb(n2481), .dout(n2598));
  jand g02343(.dina(n2490), .dinb(n2451), .dout(n2599));
  jnot g02344(.din(n2599), .dout(n2600));
  jand g02345(.dina(n2600), .dinb(n2598), .dout(n2601));
  jnot g02346(.din(n2601), .dout(n2602));
  jor  g02347(.dina(n2478), .dinb(n2470), .dout(n2603));
  jand g02348(.dina(n2479), .dinb(n2455), .dout(n2604));
  jnot g02349(.din(n2604), .dout(n2605));
  jand g02350(.dina(n2605), .dinb(n2603), .dout(n2606));
  jnot g02351(.din(n2606), .dout(n2607));
  jor  g02352(.dina(n2463), .dinb(n2317), .dout(n2608));
  jor  g02353(.dina(n2608), .dinb(n2457), .dout(n2609));
  jnot g02354(.din(n2609), .dout(n2610));
  jand g02355(.dina(n2610), .dinb(b0 ), .dout(n2611));
  jand g02356(.dina(n2458), .dinb(b2 ), .dout(n2612));
  jor  g02357(.dina(n2612), .dinb(n2611), .dout(n2613));
  jand g02358(.dina(n2460), .dinb(n273), .dout(n2614));
  jand g02359(.dina(n2464), .dinb(b1 ), .dout(n2615));
  jor  g02360(.dina(n2615), .dinb(n2614), .dout(n2616));
  jor  g02361(.dina(n2616), .dinb(n2613), .dout(n2617));
  jnot g02362(.din(n2467), .dout(n2618));
  jand g02363(.dina(n2319), .dinb(a29 ), .dout(n2619));
  jand g02364(.dina(n2619), .dinb(n2618), .dout(n2620));
  jnot g02365(.din(n2620), .dout(n2621));
  jand g02366(.dina(n2621), .dinb(a29 ), .dout(n2622));
  jxor g02367(.dina(n2622), .dinb(n2617), .dout(n2623));
  jnot g02368(.din(n2623), .dout(n2624));
  jor  g02369(.dina(n2324), .dinb(n374), .dout(n2625));
  jor  g02370(.dina(n2326), .dinb(n377), .dout(n2626));
  jor  g02371(.dina(n2186), .dinb(n303), .dout(n2627));
  jand g02372(.dina(n2627), .dinb(n2626), .dout(n2628));
  jor  g02373(.dina(n2321), .dinb(n340), .dout(n2629));
  jand g02374(.dina(n2629), .dinb(n2628), .dout(n2630));
  jand g02375(.dina(n2630), .dinb(n2625), .dout(n2631));
  jxor g02376(.dina(n2631), .dinb(a26 ), .dout(n2632));
  jxor g02377(.dina(n2632), .dinb(n2624), .dout(n2633));
  jxor g02378(.dina(n2633), .dinb(n2607), .dout(n2634));
  jor  g02379(.dina(n1921), .dinb(n517), .dout(n2635));
  jor  g02380(.dina(n1918), .dinb(n469), .dout(n2636));
  jor  g02381(.dina(n1923), .dinb(n519), .dout(n2637));
  jor  g02382(.dina(n1806), .dinb(n415), .dout(n2638));
  jand g02383(.dina(n2638), .dinb(n2637), .dout(n2639));
  jand g02384(.dina(n2639), .dinb(n2636), .dout(n2640));
  jand g02385(.dina(n2640), .dinb(n2635), .dout(n2641));
  jxor g02386(.dina(n2641), .dinb(n1687), .dout(n2642));
  jxor g02387(.dina(n2642), .dinb(n2634), .dout(n2643));
  jxor g02388(.dina(n2643), .dinb(n2602), .dout(n2644));
  jor  g02389(.dina(n1569), .dinb(n702), .dout(n2645));
  jor  g02390(.dina(n1453), .dinb(n572), .dout(n2646));
  jor  g02391(.dina(n1566), .dinb(n637), .dout(n2647));
  jor  g02392(.dina(n1571), .dinb(n704), .dout(n2648));
  jand g02393(.dina(n2648), .dinb(n2647), .dout(n2649));
  jand g02394(.dina(n2649), .dinb(n2646), .dout(n2650));
  jand g02395(.dina(n2650), .dinb(n2645), .dout(n2651));
  jxor g02396(.dina(n2651), .dinb(n1351), .dout(n2652));
  jxor g02397(.dina(n2652), .dinb(n2644), .dout(n2653));
  jxor g02398(.dina(n2653), .dinb(n2597), .dout(n2654));
  jor  g02399(.dina(n1248), .dinb(n932), .dout(n2655));
  jor  g02400(.dina(n1147), .dinb(n772), .dout(n2656));
  jor  g02401(.dina(n1251), .dinb(n852), .dout(n2657));
  jor  g02402(.dina(n1246), .dinb(n934), .dout(n2658));
  jand g02403(.dina(n2658), .dinb(n2657), .dout(n2659));
  jand g02404(.dina(n2659), .dinb(n2656), .dout(n2660));
  jand g02405(.dina(n2660), .dinb(n2655), .dout(n2661));
  jxor g02406(.dina(n2661), .dinb(n1061), .dout(n2662));
  jxor g02407(.dina(n2662), .dinb(n2654), .dout(n2663));
  jxor g02408(.dina(n2663), .dinb(n2594), .dout(n2664));
  jor  g02409(.dina(n1209), .dinb(n970), .dout(n2665));
  jor  g02410(.dina(n880), .dinb(n1018), .dout(n2666));
  jor  g02411(.dina(n972), .dinb(n1211), .dout(n2667));
  jor  g02412(.dina(n967), .dinb(n1114), .dout(n2668));
  jand g02413(.dina(n2668), .dinb(n2667), .dout(n2669));
  jand g02414(.dina(n2669), .dinb(n2666), .dout(n2670));
  jand g02415(.dina(n2670), .dinb(n2665), .dout(n2671));
  jxor g02416(.dina(n2671), .dinb(n810), .dout(n2672));
  jxor g02417(.dina(n2672), .dinb(n2664), .dout(n2673));
  jxor g02418(.dina(n2673), .dinb(n2591), .dout(n2674));
  jor  g02419(.dina(n1525), .dinb(n728), .dout(n2675));
  jor  g02420(.dina(n660), .dinb(n1307), .dout(n2676));
  jor  g02421(.dina(n726), .dinb(n1527), .dout(n2677));
  jor  g02422(.dina(n731), .dinb(n1416), .dout(n2678));
  jand g02423(.dina(n2678), .dinb(n2677), .dout(n2679));
  jand g02424(.dina(n2679), .dinb(n2676), .dout(n2680));
  jand g02425(.dina(n2680), .dinb(n2675), .dout(n2681));
  jxor g02426(.dina(n2681), .dinb(n606), .dout(n2682));
  jxor g02427(.dina(n2682), .dinb(n2674), .dout(n2683));
  jnot g02428(.din(n2683), .dout(n2684));
  jxor g02429(.dina(n2684), .dinb(n2588), .dout(n2685));
  jor  g02430(.dina(n1879), .dinb(n544), .dout(n2686));
  jor  g02431(.dina(n486), .dinb(n1637), .dout(n2687));
  jor  g02432(.dina(n547), .dinb(n1759), .dout(n2688));
  jor  g02433(.dina(n542), .dinb(n1881), .dout(n2689));
  jand g02434(.dina(n2689), .dinb(n2688), .dout(n2690));
  jand g02435(.dina(n2690), .dinb(n2687), .dout(n2691));
  jand g02436(.dina(n2691), .dinb(n2686), .dout(n2692));
  jxor g02437(.dina(n2692), .dinb(n446), .dout(n2693));
  jxor g02438(.dina(n2693), .dinb(n2685), .dout(n2694));
  jxor g02439(.dina(n2694), .dinb(n2584), .dout(n2695));
  jor  g02440(.dina(n2277), .dinb(n397), .dout(n2696));
  jor  g02441(.dina(n354), .dinb(n2007), .dout(n2697));
  jor  g02442(.dina(n394), .dinb(n2142), .dout(n2698));
  jor  g02443(.dina(n399), .dinb(n2279), .dout(n2699));
  jand g02444(.dina(n2699), .dinb(n2698), .dout(n2700));
  jand g02445(.dina(n2700), .dinb(n2697), .dout(n2701));
  jand g02446(.dina(n2701), .dinb(n2696), .dout(n2702));
  jxor g02447(.dina(n2702), .dinb(n364), .dout(n2703));
  jxor g02448(.dina(n2703), .dinb(n2695), .dout(n2704));
  jxor g02449(.dina(n2704), .dinb(n2581), .dout(n2705));
  jand g02450(.dina(b28 ), .dinb(b27 ), .dout(n2706));
  jand g02451(.dina(n2559), .dinb(n2558), .dout(n2707));
  jor  g02452(.dina(n2707), .dinb(n2706), .dout(n2708));
  jxor g02453(.dina(b29 ), .dinb(b28 ), .dout(n2709));
  jnot g02454(.din(n2709), .dout(n2710));
  jxor g02455(.dina(n2710), .dinb(n2708), .dout(n2711));
  jor  g02456(.dina(n2711), .dinb(n296), .dout(n2712));
  jnot g02457(.din(b29 ), .dout(n2713));
  jor  g02458(.dina(n264), .dinb(n2713), .dout(n2714));
  jor  g02459(.dina(n294), .dinb(n2563), .dout(n2715));
  jor  g02460(.dina(n280), .dinb(n2415), .dout(n2716));
  jand g02461(.dina(n2716), .dinb(n2715), .dout(n2717));
  jand g02462(.dina(n2717), .dinb(n2714), .dout(n2718));
  jand g02463(.dina(n2718), .dinb(n2712), .dout(n2719));
  jxor g02464(.dina(n2719), .dinb(n278), .dout(n2720));
  jxor g02465(.dina(n2720), .dinb(n2705), .dout(n2721));
  jxor g02466(.dina(n2721), .dinb(n2576), .dout(f29 ));
  jnot g02467(.din(n2720), .dout(n2723));
  jor  g02468(.dina(n2723), .dinb(n2705), .dout(n2724));
  jor  g02469(.dina(n2721), .dinb(n2576), .dout(n2725));
  jand g02470(.dina(n2725), .dinb(n2724), .dout(n2726));
  jand g02471(.dina(n2703), .dinb(n2695), .dout(n2727));
  jnot g02472(.din(n2727), .dout(n2728));
  jnot g02473(.din(n2704), .dout(n2729));
  jor  g02474(.dina(n2729), .dinb(n2581), .dout(n2730));
  jand g02475(.dina(n2730), .dinb(n2728), .dout(n2731));
  jand g02476(.dina(n2693), .dinb(n2685), .dout(n2732));
  jand g02477(.dina(n2694), .dinb(n2584), .dout(n2733));
  jor  g02478(.dina(n2733), .dinb(n2732), .dout(n2734));
  jand g02479(.dina(n2682), .dinb(n2674), .dout(n2735));
  jnot g02480(.din(n2735), .dout(n2736));
  jor  g02481(.dina(n2684), .dinb(n2588), .dout(n2737));
  jand g02482(.dina(n2737), .dinb(n2736), .dout(n2738));
  jand g02483(.dina(n2672), .dinb(n2664), .dout(n2739));
  jand g02484(.dina(n2673), .dinb(n2591), .dout(n2740));
  jor  g02485(.dina(n2740), .dinb(n2739), .dout(n2741));
  jand g02486(.dina(n2662), .dinb(n2654), .dout(n2742));
  jand g02487(.dina(n2663), .dinb(n2594), .dout(n2743));
  jor  g02488(.dina(n2743), .dinb(n2742), .dout(n2744));
  jand g02489(.dina(n2652), .dinb(n2644), .dout(n2745));
  jand g02490(.dina(n2653), .dinb(n2597), .dout(n2746));
  jor  g02491(.dina(n2746), .dinb(n2745), .dout(n2747));
  jand g02492(.dina(n2642), .dinb(n2634), .dout(n2748));
  jand g02493(.dina(n2643), .dinb(n2602), .dout(n2749));
  jor  g02494(.dina(n2749), .dinb(n2748), .dout(n2750));
  jor  g02495(.dina(n2632), .dinb(n2624), .dout(n2751));
  jand g02496(.dina(n2633), .dinb(n2607), .dout(n2752));
  jnot g02497(.din(n2752), .dout(n2753));
  jand g02498(.dina(n2753), .dinb(n2751), .dout(n2754));
  jnot g02499(.din(n2754), .dout(n2755));
  jor  g02500(.dina(n2621), .dinb(n2617), .dout(n2756));
  jxor g02501(.dina(a30 ), .dinb(a29 ), .dout(n2757));
  jand g02502(.dina(n2757), .dinb(b0 ), .dout(n2758));
  jnot g02503(.din(n2758), .dout(n2759));
  jxor g02504(.dina(n2759), .dinb(n2756), .dout(n2760));
  jnot g02505(.din(n2458), .dout(n2761));
  jor  g02506(.dina(n2761), .dinb(n303), .dout(n2762));
  jor  g02507(.dina(n2609), .dinb(n305), .dout(n2763));
  jnot g02508(.din(n2460), .dout(n2764));
  jor  g02509(.dina(n2764), .dinb(n301), .dout(n2765));
  jnot g02510(.din(n2464), .dout(n2766));
  jor  g02511(.dina(n2766), .dinb(n293), .dout(n2767));
  jand g02512(.dina(n2767), .dinb(n2765), .dout(n2768));
  jand g02513(.dina(n2768), .dinb(n2763), .dout(n2769));
  jand g02514(.dina(n2769), .dinb(n2762), .dout(n2770));
  jxor g02515(.dina(n2770), .dinb(n2468), .dout(n2771));
  jxor g02516(.dina(n2771), .dinb(n2760), .dout(n2772));
  jnot g02517(.din(n2772), .dout(n2773));
  jor  g02518(.dina(n2324), .dinb(n412), .dout(n2774));
  jor  g02519(.dina(n2321), .dinb(n377), .dout(n2775));
  jor  g02520(.dina(n2186), .dinb(n340), .dout(n2776));
  jand g02521(.dina(n2776), .dinb(n2775), .dout(n2777));
  jor  g02522(.dina(n2326), .dinb(n415), .dout(n2778));
  jand g02523(.dina(n2778), .dinb(n2777), .dout(n2779));
  jand g02524(.dina(n2779), .dinb(n2774), .dout(n2780));
  jxor g02525(.dina(n2780), .dinb(a26 ), .dout(n2781));
  jxor g02526(.dina(n2781), .dinb(n2773), .dout(n2782));
  jxor g02527(.dina(n2782), .dinb(n2755), .dout(n2783));
  jor  g02528(.dina(n1921), .dinb(n570), .dout(n2784));
  jor  g02529(.dina(n1806), .dinb(n469), .dout(n2785));
  jor  g02530(.dina(n1918), .dinb(n519), .dout(n2786));
  jor  g02531(.dina(n1923), .dinb(n572), .dout(n2787));
  jand g02532(.dina(n2787), .dinb(n2786), .dout(n2788));
  jand g02533(.dina(n2788), .dinb(n2785), .dout(n2789));
  jand g02534(.dina(n2789), .dinb(n2784), .dout(n2790));
  jxor g02535(.dina(n2790), .dinb(n1687), .dout(n2791));
  jxor g02536(.dina(n2791), .dinb(n2783), .dout(n2792));
  jxor g02537(.dina(n2792), .dinb(n2750), .dout(n2793));
  jor  g02538(.dina(n1569), .dinb(n770), .dout(n2794));
  jor  g02539(.dina(n1453), .dinb(n637), .dout(n2795));
  jor  g02540(.dina(n1571), .dinb(n772), .dout(n2796));
  jor  g02541(.dina(n1566), .dinb(n704), .dout(n2797));
  jand g02542(.dina(n2797), .dinb(n2796), .dout(n2798));
  jand g02543(.dina(n2798), .dinb(n2795), .dout(n2799));
  jand g02544(.dina(n2799), .dinb(n2794), .dout(n2800));
  jxor g02545(.dina(n2800), .dinb(n1351), .dout(n2801));
  jxor g02546(.dina(n2801), .dinb(n2793), .dout(n2802));
  jxor g02547(.dina(n2802), .dinb(n2747), .dout(n2803));
  jor  g02548(.dina(n1248), .dinb(n1016), .dout(n2804));
  jor  g02549(.dina(n1147), .dinb(n852), .dout(n2805));
  jor  g02550(.dina(n1251), .dinb(n934), .dout(n2806));
  jor  g02551(.dina(n1246), .dinb(n1018), .dout(n2807));
  jand g02552(.dina(n2807), .dinb(n2806), .dout(n2808));
  jand g02553(.dina(n2808), .dinb(n2805), .dout(n2809));
  jand g02554(.dina(n2809), .dinb(n2804), .dout(n2810));
  jxor g02555(.dina(n2810), .dinb(n1061), .dout(n2811));
  jxor g02556(.dina(n2811), .dinb(n2803), .dout(n2812));
  jxor g02557(.dina(n2812), .dinb(n2744), .dout(n2813));
  jor  g02558(.dina(n1305), .dinb(n970), .dout(n2814));
  jor  g02559(.dina(n880), .dinb(n1114), .dout(n2815));
  jor  g02560(.dina(n967), .dinb(n1211), .dout(n2816));
  jor  g02561(.dina(n972), .dinb(n1307), .dout(n2817));
  jand g02562(.dina(n2817), .dinb(n2816), .dout(n2818));
  jand g02563(.dina(n2818), .dinb(n2815), .dout(n2819));
  jand g02564(.dina(n2819), .dinb(n2814), .dout(n2820));
  jxor g02565(.dina(n2820), .dinb(n810), .dout(n2821));
  jxor g02566(.dina(n2821), .dinb(n2813), .dout(n2822));
  jxor g02567(.dina(n2822), .dinb(n2741), .dout(n2823));
  jor  g02568(.dina(n1635), .dinb(n728), .dout(n2824));
  jor  g02569(.dina(n660), .dinb(n1416), .dout(n2825));
  jor  g02570(.dina(n731), .dinb(n1527), .dout(n2826));
  jor  g02571(.dina(n726), .dinb(n1637), .dout(n2827));
  jand g02572(.dina(n2827), .dinb(n2826), .dout(n2828));
  jand g02573(.dina(n2828), .dinb(n2825), .dout(n2829));
  jand g02574(.dina(n2829), .dinb(n2824), .dout(n2830));
  jxor g02575(.dina(n2830), .dinb(n606), .dout(n2831));
  jxor g02576(.dina(n2831), .dinb(n2823), .dout(n2832));
  jnot g02577(.din(n2832), .dout(n2833));
  jxor g02578(.dina(n2833), .dinb(n2738), .dout(n2834));
  jor  g02579(.dina(n2005), .dinb(n544), .dout(n2835));
  jor  g02580(.dina(n486), .dinb(n1759), .dout(n2836));
  jor  g02581(.dina(n542), .dinb(n2007), .dout(n2837));
  jor  g02582(.dina(n547), .dinb(n1881), .dout(n2838));
  jand g02583(.dina(n2838), .dinb(n2837), .dout(n2839));
  jand g02584(.dina(n2839), .dinb(n2836), .dout(n2840));
  jand g02585(.dina(n2840), .dinb(n2835), .dout(n2841));
  jxor g02586(.dina(n2841), .dinb(n446), .dout(n2842));
  jxor g02587(.dina(n2842), .dinb(n2834), .dout(n2843));
  jxor g02588(.dina(n2843), .dinb(n2734), .dout(n2844));
  jor  g02589(.dina(n2413), .dinb(n397), .dout(n2845));
  jor  g02590(.dina(n354), .dinb(n2142), .dout(n2846));
  jor  g02591(.dina(n394), .dinb(n2279), .dout(n2847));
  jor  g02592(.dina(n399), .dinb(n2415), .dout(n2848));
  jand g02593(.dina(n2848), .dinb(n2847), .dout(n2849));
  jand g02594(.dina(n2849), .dinb(n2846), .dout(n2850));
  jand g02595(.dina(n2850), .dinb(n2845), .dout(n2851));
  jxor g02596(.dina(n2851), .dinb(n364), .dout(n2852));
  jxor g02597(.dina(n2852), .dinb(n2844), .dout(n2853));
  jxor g02598(.dina(n2853), .dinb(n2731), .dout(n2854));
  jand g02599(.dina(b29 ), .dinb(b28 ), .dout(n2855));
  jand g02600(.dina(n2709), .dinb(n2708), .dout(n2856));
  jor  g02601(.dina(n2856), .dinb(n2855), .dout(n2857));
  jxor g02602(.dina(b30 ), .dinb(b29 ), .dout(n2858));
  jnot g02603(.din(n2858), .dout(n2859));
  jxor g02604(.dina(n2859), .dinb(n2857), .dout(n2860));
  jor  g02605(.dina(n2860), .dinb(n296), .dout(n2861));
  jnot g02606(.din(b30 ), .dout(n2862));
  jor  g02607(.dina(n264), .dinb(n2862), .dout(n2863));
  jor  g02608(.dina(n280), .dinb(n2563), .dout(n2864));
  jor  g02609(.dina(n294), .dinb(n2713), .dout(n2865));
  jand g02610(.dina(n2865), .dinb(n2864), .dout(n2866));
  jand g02611(.dina(n2866), .dinb(n2863), .dout(n2867));
  jand g02612(.dina(n2867), .dinb(n2861), .dout(n2868));
  jxor g02613(.dina(n2868), .dinb(n278), .dout(n2869));
  jxor g02614(.dina(n2869), .dinb(n2854), .dout(n2870));
  jxor g02615(.dina(n2870), .dinb(n2726), .dout(f30 ));
  jnot g02616(.din(n2869), .dout(n2872));
  jor  g02617(.dina(n2872), .dinb(n2854), .dout(n2873));
  jor  g02618(.dina(n2870), .dinb(n2726), .dout(n2874));
  jand g02619(.dina(n2874), .dinb(n2873), .dout(n2875));
  jand g02620(.dina(n2852), .dinb(n2844), .dout(n2876));
  jnot g02621(.din(n2876), .dout(n2877));
  jnot g02622(.din(n2853), .dout(n2878));
  jor  g02623(.dina(n2878), .dinb(n2731), .dout(n2879));
  jand g02624(.dina(n2879), .dinb(n2877), .dout(n2880));
  jand g02625(.dina(n2842), .dinb(n2834), .dout(n2881));
  jand g02626(.dina(n2843), .dinb(n2734), .dout(n2882));
  jor  g02627(.dina(n2882), .dinb(n2881), .dout(n2883));
  jand g02628(.dina(n2831), .dinb(n2823), .dout(n2884));
  jnot g02629(.din(n2884), .dout(n2885));
  jor  g02630(.dina(n2833), .dinb(n2738), .dout(n2886));
  jand g02631(.dina(n2886), .dinb(n2885), .dout(n2887));
  jand g02632(.dina(n2821), .dinb(n2813), .dout(n2888));
  jand g02633(.dina(n2822), .dinb(n2741), .dout(n2889));
  jor  g02634(.dina(n2889), .dinb(n2888), .dout(n2890));
  jand g02635(.dina(n2811), .dinb(n2803), .dout(n2891));
  jand g02636(.dina(n2812), .dinb(n2744), .dout(n2892));
  jor  g02637(.dina(n2892), .dinb(n2891), .dout(n2893));
  jand g02638(.dina(n2791), .dinb(n2783), .dout(n2894));
  jand g02639(.dina(n2792), .dinb(n2750), .dout(n2895));
  jor  g02640(.dina(n2895), .dinb(n2894), .dout(n2896));
  jor  g02641(.dina(n2781), .dinb(n2773), .dout(n2897));
  jand g02642(.dina(n2782), .dinb(n2755), .dout(n2898));
  jnot g02643(.din(n2898), .dout(n2899));
  jand g02644(.dina(n2899), .dinb(n2897), .dout(n2900));
  jnot g02645(.din(n2900), .dout(n2901));
  jnot g02646(.din(n2756), .dout(n2902));
  jand g02647(.dina(n2758), .dinb(n2902), .dout(n2903));
  jand g02648(.dina(n2771), .dinb(n2760), .dout(n2904));
  jor  g02649(.dina(n2904), .dinb(n2903), .dout(n2905));
  jxor g02650(.dina(a32 ), .dinb(a31 ), .dout(n2906));
  jand g02651(.dina(n2906), .dinb(n2757), .dout(n2907));
  jand g02652(.dina(n2907), .dinb(n259), .dout(n2908));
  jnot g02653(.din(n2757), .dout(n2909));
  jxor g02654(.dina(a31 ), .dinb(a30 ), .dout(n2910));
  jand g02655(.dina(n2910), .dinb(n2909), .dout(n2911));
  jand g02656(.dina(n2911), .dinb(b0 ), .dout(n2912));
  jnot g02657(.din(n2906), .dout(n2913));
  jand g02658(.dina(n2913), .dinb(n2757), .dout(n2914));
  jand g02659(.dina(n2914), .dinb(b1 ), .dout(n2915));
  jor  g02660(.dina(n2915), .dinb(n2912), .dout(n2916));
  jor  g02661(.dina(n2916), .dinb(n2908), .dout(n2917));
  jnot g02662(.din(a32 ), .dout(n2918));
  jor  g02663(.dina(n2759), .dinb(n2918), .dout(n2919));
  jxor g02664(.dina(n2919), .dinb(n2917), .dout(n2920));
  jor  g02665(.dina(n2764), .dinb(n337), .dout(n2921));
  jor  g02666(.dina(n2766), .dinb(n303), .dout(n2922));
  jor  g02667(.dina(n2609), .dinb(n293), .dout(n2923));
  jand g02668(.dina(n2923), .dinb(n2922), .dout(n2924));
  jor  g02669(.dina(n2761), .dinb(n340), .dout(n2925));
  jand g02670(.dina(n2925), .dinb(n2924), .dout(n2926));
  jand g02671(.dina(n2926), .dinb(n2921), .dout(n2927));
  jxor g02672(.dina(n2927), .dinb(a29 ), .dout(n2928));
  jxor g02673(.dina(n2928), .dinb(n2920), .dout(n2929));
  jxor g02674(.dina(n2929), .dinb(n2905), .dout(n2930));
  jnot g02675(.din(n2930), .dout(n2931));
  jor  g02676(.dina(n2324), .dinb(n466), .dout(n2932));
  jor  g02677(.dina(n2326), .dinb(n469), .dout(n2933));
  jor  g02678(.dina(n2186), .dinb(n377), .dout(n2934));
  jand g02679(.dina(n2934), .dinb(n2933), .dout(n2935));
  jor  g02680(.dina(n2321), .dinb(n415), .dout(n2936));
  jand g02681(.dina(n2936), .dinb(n2935), .dout(n2937));
  jand g02682(.dina(n2937), .dinb(n2932), .dout(n2938));
  jxor g02683(.dina(n2938), .dinb(a26 ), .dout(n2939));
  jxor g02684(.dina(n2939), .dinb(n2931), .dout(n2940));
  jxor g02685(.dina(n2940), .dinb(n2901), .dout(n2941));
  jor  g02686(.dina(n1921), .dinb(n635), .dout(n2942));
  jor  g02687(.dina(n1806), .dinb(n519), .dout(n2943));
  jor  g02688(.dina(n1918), .dinb(n572), .dout(n2944));
  jor  g02689(.dina(n1923), .dinb(n637), .dout(n2945));
  jand g02690(.dina(n2945), .dinb(n2944), .dout(n2946));
  jand g02691(.dina(n2946), .dinb(n2943), .dout(n2947));
  jand g02692(.dina(n2947), .dinb(n2942), .dout(n2948));
  jxor g02693(.dina(n2948), .dinb(n1687), .dout(n2949));
  jxor g02694(.dina(n2949), .dinb(n2941), .dout(n2950));
  jxor g02695(.dina(n2950), .dinb(n2896), .dout(n2951));
  jor  g02696(.dina(n1569), .dinb(n850), .dout(n2952));
  jor  g02697(.dina(n1453), .dinb(n704), .dout(n2953));
  jor  g02698(.dina(n1566), .dinb(n772), .dout(n2954));
  jor  g02699(.dina(n1571), .dinb(n852), .dout(n2955));
  jand g02700(.dina(n2955), .dinb(n2954), .dout(n2956));
  jand g02701(.dina(n2956), .dinb(n2953), .dout(n2957));
  jand g02702(.dina(n2957), .dinb(n2952), .dout(n2958));
  jxor g02703(.dina(n2958), .dinb(n1351), .dout(n2959));
  jxor g02704(.dina(n2959), .dinb(n2951), .dout(n2960));
  jand g02705(.dina(n2801), .dinb(n2793), .dout(n2961));
  jand g02706(.dina(n2802), .dinb(n2747), .dout(n2962));
  jor  g02707(.dina(n2962), .dinb(n2961), .dout(n2963));
  jxor g02708(.dina(n2963), .dinb(n2960), .dout(n2964));
  jor  g02709(.dina(n1112), .dinb(n1248), .dout(n2965));
  jor  g02710(.dina(n1147), .dinb(n934), .dout(n2966));
  jor  g02711(.dina(n1251), .dinb(n1018), .dout(n2967));
  jor  g02712(.dina(n1246), .dinb(n1114), .dout(n2968));
  jand g02713(.dina(n2968), .dinb(n2967), .dout(n2969));
  jand g02714(.dina(n2969), .dinb(n2966), .dout(n2970));
  jand g02715(.dina(n2970), .dinb(n2965), .dout(n2971));
  jxor g02716(.dina(n2971), .dinb(n1061), .dout(n2972));
  jxor g02717(.dina(n2972), .dinb(n2964), .dout(n2973));
  jxor g02718(.dina(n2973), .dinb(n2893), .dout(n2974));
  jor  g02719(.dina(n1414), .dinb(n970), .dout(n2975));
  jor  g02720(.dina(n880), .dinb(n1211), .dout(n2976));
  jor  g02721(.dina(n972), .dinb(n1416), .dout(n2977));
  jor  g02722(.dina(n967), .dinb(n1307), .dout(n2978));
  jand g02723(.dina(n2978), .dinb(n2977), .dout(n2979));
  jand g02724(.dina(n2979), .dinb(n2976), .dout(n2980));
  jand g02725(.dina(n2980), .dinb(n2975), .dout(n2981));
  jxor g02726(.dina(n2981), .dinb(n810), .dout(n2982));
  jxor g02727(.dina(n2982), .dinb(n2974), .dout(n2983));
  jxor g02728(.dina(n2983), .dinb(n2890), .dout(n2984));
  jor  g02729(.dina(n1757), .dinb(n728), .dout(n2985));
  jor  g02730(.dina(n660), .dinb(n1527), .dout(n2986));
  jor  g02731(.dina(n726), .dinb(n1759), .dout(n2987));
  jor  g02732(.dina(n731), .dinb(n1637), .dout(n2988));
  jand g02733(.dina(n2988), .dinb(n2987), .dout(n2989));
  jand g02734(.dina(n2989), .dinb(n2986), .dout(n2990));
  jand g02735(.dina(n2990), .dinb(n2985), .dout(n2991));
  jxor g02736(.dina(n2991), .dinb(n606), .dout(n2992));
  jxor g02737(.dina(n2992), .dinb(n2984), .dout(n2993));
  jnot g02738(.din(n2993), .dout(n2994));
  jxor g02739(.dina(n2994), .dinb(n2887), .dout(n2995));
  jor  g02740(.dina(n2140), .dinb(n544), .dout(n2996));
  jor  g02741(.dina(n486), .dinb(n1881), .dout(n2997));
  jor  g02742(.dina(n542), .dinb(n2142), .dout(n2998));
  jor  g02743(.dina(n547), .dinb(n2007), .dout(n2999));
  jand g02744(.dina(n2999), .dinb(n2998), .dout(n3000));
  jand g02745(.dina(n3000), .dinb(n2997), .dout(n3001));
  jand g02746(.dina(n3001), .dinb(n2996), .dout(n3002));
  jxor g02747(.dina(n3002), .dinb(n446), .dout(n3003));
  jxor g02748(.dina(n3003), .dinb(n2995), .dout(n3004));
  jxor g02749(.dina(n3004), .dinb(n2883), .dout(n3005));
  jor  g02750(.dina(n2561), .dinb(n397), .dout(n3006));
  jor  g02751(.dina(n354), .dinb(n2279), .dout(n3007));
  jor  g02752(.dina(n394), .dinb(n2415), .dout(n3008));
  jor  g02753(.dina(n399), .dinb(n2563), .dout(n3009));
  jand g02754(.dina(n3009), .dinb(n3008), .dout(n3010));
  jand g02755(.dina(n3010), .dinb(n3007), .dout(n3011));
  jand g02756(.dina(n3011), .dinb(n3006), .dout(n3012));
  jxor g02757(.dina(n3012), .dinb(n364), .dout(n3013));
  jxor g02758(.dina(n3013), .dinb(n3005), .dout(n3014));
  jxor g02759(.dina(n3014), .dinb(n2880), .dout(n3015));
  jand g02760(.dina(b30 ), .dinb(b29 ), .dout(n3016));
  jand g02761(.dina(n2858), .dinb(n2857), .dout(n3017));
  jor  g02762(.dina(n3017), .dinb(n3016), .dout(n3018));
  jxor g02763(.dina(b31 ), .dinb(b30 ), .dout(n3019));
  jnot g02764(.din(n3019), .dout(n3020));
  jxor g02765(.dina(n3020), .dinb(n3018), .dout(n3021));
  jor  g02766(.dina(n3021), .dinb(n296), .dout(n3022));
  jnot g02767(.din(b31 ), .dout(n3023));
  jor  g02768(.dina(n264), .dinb(n3023), .dout(n3024));
  jor  g02769(.dina(n294), .dinb(n2862), .dout(n3025));
  jor  g02770(.dina(n280), .dinb(n2713), .dout(n3026));
  jand g02771(.dina(n3026), .dinb(n3025), .dout(n3027));
  jand g02772(.dina(n3027), .dinb(n3024), .dout(n3028));
  jand g02773(.dina(n3028), .dinb(n3022), .dout(n3029));
  jxor g02774(.dina(n3029), .dinb(n278), .dout(n3030));
  jxor g02775(.dina(n3030), .dinb(n3015), .dout(n3031));
  jxor g02776(.dina(n3031), .dinb(n2875), .dout(f31 ));
  jnot g02777(.din(n3030), .dout(n3033));
  jor  g02778(.dina(n3033), .dinb(n3015), .dout(n3034));
  jor  g02779(.dina(n3031), .dinb(n2875), .dout(n3035));
  jand g02780(.dina(n3035), .dinb(n3034), .dout(n3036));
  jand g02781(.dina(n3013), .dinb(n3005), .dout(n3037));
  jnot g02782(.din(n3037), .dout(n3038));
  jnot g02783(.din(n3014), .dout(n3039));
  jor  g02784(.dina(n3039), .dinb(n2880), .dout(n3040));
  jand g02785(.dina(n3040), .dinb(n3038), .dout(n3041));
  jand g02786(.dina(n3003), .dinb(n2995), .dout(n3042));
  jand g02787(.dina(n3004), .dinb(n2883), .dout(n3043));
  jor  g02788(.dina(n3043), .dinb(n3042), .dout(n3044));
  jand g02789(.dina(n2992), .dinb(n2984), .dout(n3045));
  jnot g02790(.din(n3045), .dout(n3046));
  jor  g02791(.dina(n2994), .dinb(n2887), .dout(n3047));
  jand g02792(.dina(n3047), .dinb(n3046), .dout(n3048));
  jand g02793(.dina(n2982), .dinb(n2974), .dout(n3049));
  jand g02794(.dina(n2983), .dinb(n2890), .dout(n3050));
  jor  g02795(.dina(n3050), .dinb(n3049), .dout(n3051));
  jand g02796(.dina(n2972), .dinb(n2964), .dout(n3052));
  jand g02797(.dina(n2973), .dinb(n2893), .dout(n3053));
  jor  g02798(.dina(n3053), .dinb(n3052), .dout(n3054));
  jand g02799(.dina(n2959), .dinb(n2951), .dout(n3055));
  jand g02800(.dina(n2963), .dinb(n2960), .dout(n3056));
  jor  g02801(.dina(n3056), .dinb(n3055), .dout(n3057));
  jand g02802(.dina(n2949), .dinb(n2941), .dout(n3058));
  jand g02803(.dina(n2950), .dinb(n2896), .dout(n3059));
  jor  g02804(.dina(n3059), .dinb(n3058), .dout(n3060));
  jor  g02805(.dina(n2939), .dinb(n2931), .dout(n3061));
  jand g02806(.dina(n2940), .dinb(n2901), .dout(n3062));
  jnot g02807(.din(n3062), .dout(n3063));
  jand g02808(.dina(n3063), .dinb(n3061), .dout(n3064));
  jnot g02809(.din(n3064), .dout(n3065));
  jor  g02810(.dina(n2928), .dinb(n2920), .dout(n3066));
  jand g02811(.dina(n2929), .dinb(n2905), .dout(n3067));
  jnot g02812(.din(n3067), .dout(n3068));
  jand g02813(.dina(n3068), .dinb(n3066), .dout(n3069));
  jnot g02814(.din(n3069), .dout(n3070));
  jor  g02815(.dina(n2910), .dinb(n2757), .dout(n3071));
  jor  g02816(.dina(n3071), .dinb(n2913), .dout(n3072));
  jnot g02817(.din(n3072), .dout(n3073));
  jand g02818(.dina(n3073), .dinb(b0 ), .dout(n3074));
  jand g02819(.dina(n2911), .dinb(b1 ), .dout(n3075));
  jor  g02820(.dina(n3075), .dinb(n3074), .dout(n3076));
  jand g02821(.dina(n2907), .dinb(n273), .dout(n3077));
  jand g02822(.dina(n2914), .dinb(b2 ), .dout(n3078));
  jor  g02823(.dina(n3078), .dinb(n3077), .dout(n3079));
  jor  g02824(.dina(n3079), .dinb(n3076), .dout(n3080));
  jnot g02825(.din(n2917), .dout(n3081));
  jand g02826(.dina(n2759), .dinb(a32 ), .dout(n3082));
  jand g02827(.dina(n3082), .dinb(n3081), .dout(n3083));
  jnot g02828(.din(n3083), .dout(n3084));
  jand g02829(.dina(n3084), .dinb(a32 ), .dout(n3085));
  jxor g02830(.dina(n3085), .dinb(n3080), .dout(n3086));
  jnot g02831(.din(n3086), .dout(n3087));
  jor  g02832(.dina(n2764), .dinb(n374), .dout(n3088));
  jor  g02833(.dina(n2766), .dinb(n340), .dout(n3089));
  jor  g02834(.dina(n2609), .dinb(n303), .dout(n3090));
  jand g02835(.dina(n3090), .dinb(n3089), .dout(n3091));
  jor  g02836(.dina(n2761), .dinb(n377), .dout(n3092));
  jand g02837(.dina(n3092), .dinb(n3091), .dout(n3093));
  jand g02838(.dina(n3093), .dinb(n3088), .dout(n3094));
  jxor g02839(.dina(n3094), .dinb(a29 ), .dout(n3095));
  jxor g02840(.dina(n3095), .dinb(n3087), .dout(n3096));
  jxor g02841(.dina(n3096), .dinb(n3070), .dout(n3097));
  jor  g02842(.dina(n2324), .dinb(n517), .dout(n3098));
  jor  g02843(.dina(n2326), .dinb(n519), .dout(n3099));
  jor  g02844(.dina(n2321), .dinb(n469), .dout(n3100));
  jor  g02845(.dina(n2186), .dinb(n415), .dout(n3101));
  jand g02846(.dina(n3101), .dinb(n3100), .dout(n3102));
  jand g02847(.dina(n3102), .dinb(n3099), .dout(n3103));
  jand g02848(.dina(n3103), .dinb(n3098), .dout(n3104));
  jxor g02849(.dina(n3104), .dinb(n2057), .dout(n3105));
  jxor g02850(.dina(n3105), .dinb(n3097), .dout(n3106));
  jxor g02851(.dina(n3106), .dinb(n3065), .dout(n3107));
  jor  g02852(.dina(n1921), .dinb(n702), .dout(n3108));
  jor  g02853(.dina(n1806), .dinb(n572), .dout(n3109));
  jor  g02854(.dina(n1918), .dinb(n637), .dout(n3110));
  jor  g02855(.dina(n1923), .dinb(n704), .dout(n3111));
  jand g02856(.dina(n3111), .dinb(n3110), .dout(n3112));
  jand g02857(.dina(n3112), .dinb(n3109), .dout(n3113));
  jand g02858(.dina(n3113), .dinb(n3108), .dout(n3114));
  jxor g02859(.dina(n3114), .dinb(n1687), .dout(n3115));
  jxor g02860(.dina(n3115), .dinb(n3107), .dout(n3116));
  jxor g02861(.dina(n3116), .dinb(n3060), .dout(n3117));
  jor  g02862(.dina(n1569), .dinb(n932), .dout(n3118));
  jor  g02863(.dina(n1453), .dinb(n772), .dout(n3119));
  jor  g02864(.dina(n1566), .dinb(n852), .dout(n3120));
  jor  g02865(.dina(n1571), .dinb(n934), .dout(n3121));
  jand g02866(.dina(n3121), .dinb(n3120), .dout(n3122));
  jand g02867(.dina(n3122), .dinb(n3119), .dout(n3123));
  jand g02868(.dina(n3123), .dinb(n3118), .dout(n3124));
  jxor g02869(.dina(n3124), .dinb(n1351), .dout(n3125));
  jxor g02870(.dina(n3125), .dinb(n3117), .dout(n3126));
  jxor g02871(.dina(n3126), .dinb(n3057), .dout(n3127));
  jor  g02872(.dina(n1209), .dinb(n1248), .dout(n3128));
  jor  g02873(.dina(n1147), .dinb(n1018), .dout(n3129));
  jor  g02874(.dina(n1246), .dinb(n1211), .dout(n3130));
  jor  g02875(.dina(n1251), .dinb(n1114), .dout(n3131));
  jand g02876(.dina(n3131), .dinb(n3130), .dout(n3132));
  jand g02877(.dina(n3132), .dinb(n3129), .dout(n3133));
  jand g02878(.dina(n3133), .dinb(n3128), .dout(n3134));
  jxor g02879(.dina(n3134), .dinb(n1061), .dout(n3135));
  jxor g02880(.dina(n3135), .dinb(n3127), .dout(n3136));
  jxor g02881(.dina(n3136), .dinb(n3054), .dout(n3137));
  jor  g02882(.dina(n1525), .dinb(n970), .dout(n3138));
  jor  g02883(.dina(n880), .dinb(n1307), .dout(n3139));
  jor  g02884(.dina(n967), .dinb(n1416), .dout(n3140));
  jor  g02885(.dina(n972), .dinb(n1527), .dout(n3141));
  jand g02886(.dina(n3141), .dinb(n3140), .dout(n3142));
  jand g02887(.dina(n3142), .dinb(n3139), .dout(n3143));
  jand g02888(.dina(n3143), .dinb(n3138), .dout(n3144));
  jxor g02889(.dina(n3144), .dinb(n810), .dout(n3145));
  jxor g02890(.dina(n3145), .dinb(n3137), .dout(n3146));
  jxor g02891(.dina(n3146), .dinb(n3051), .dout(n3147));
  jor  g02892(.dina(n1879), .dinb(n728), .dout(n3148));
  jor  g02893(.dina(n660), .dinb(n1637), .dout(n3149));
  jor  g02894(.dina(n731), .dinb(n1759), .dout(n3150));
  jor  g02895(.dina(n726), .dinb(n1881), .dout(n3151));
  jand g02896(.dina(n3151), .dinb(n3150), .dout(n3152));
  jand g02897(.dina(n3152), .dinb(n3149), .dout(n3153));
  jand g02898(.dina(n3153), .dinb(n3148), .dout(n3154));
  jxor g02899(.dina(n3154), .dinb(n606), .dout(n3155));
  jxor g02900(.dina(n3155), .dinb(n3147), .dout(n3156));
  jnot g02901(.din(n3156), .dout(n3157));
  jxor g02902(.dina(n3157), .dinb(n3048), .dout(n3158));
  jor  g02903(.dina(n2277), .dinb(n544), .dout(n3159));
  jor  g02904(.dina(n486), .dinb(n2007), .dout(n3160));
  jor  g02905(.dina(n547), .dinb(n2142), .dout(n3161));
  jor  g02906(.dina(n542), .dinb(n2279), .dout(n3162));
  jand g02907(.dina(n3162), .dinb(n3161), .dout(n3163));
  jand g02908(.dina(n3163), .dinb(n3160), .dout(n3164));
  jand g02909(.dina(n3164), .dinb(n3159), .dout(n3165));
  jxor g02910(.dina(n3165), .dinb(n446), .dout(n3166));
  jxor g02911(.dina(n3166), .dinb(n3158), .dout(n3167));
  jxor g02912(.dina(n3167), .dinb(n3044), .dout(n3168));
  jor  g02913(.dina(n2711), .dinb(n397), .dout(n3169));
  jor  g02914(.dina(n354), .dinb(n2415), .dout(n3170));
  jor  g02915(.dina(n399), .dinb(n2713), .dout(n3171));
  jor  g02916(.dina(n394), .dinb(n2563), .dout(n3172));
  jand g02917(.dina(n3172), .dinb(n3171), .dout(n3173));
  jand g02918(.dina(n3173), .dinb(n3170), .dout(n3174));
  jand g02919(.dina(n3174), .dinb(n3169), .dout(n3175));
  jxor g02920(.dina(n3175), .dinb(n364), .dout(n3176));
  jxor g02921(.dina(n3176), .dinb(n3168), .dout(n3177));
  jxor g02922(.dina(n3177), .dinb(n3041), .dout(n3178));
  jand g02923(.dina(b31 ), .dinb(b30 ), .dout(n3179));
  jand g02924(.dina(n3019), .dinb(n3018), .dout(n3180));
  jor  g02925(.dina(n3180), .dinb(n3179), .dout(n3181));
  jxor g02926(.dina(b32 ), .dinb(b31 ), .dout(n3182));
  jnot g02927(.din(n3182), .dout(n3183));
  jxor g02928(.dina(n3183), .dinb(n3181), .dout(n3184));
  jor  g02929(.dina(n3184), .dinb(n296), .dout(n3185));
  jnot g02930(.din(b32 ), .dout(n3186));
  jor  g02931(.dina(n264), .dinb(n3186), .dout(n3187));
  jor  g02932(.dina(n280), .dinb(n2862), .dout(n3188));
  jor  g02933(.dina(n294), .dinb(n3023), .dout(n3189));
  jand g02934(.dina(n3189), .dinb(n3188), .dout(n3190));
  jand g02935(.dina(n3190), .dinb(n3187), .dout(n3191));
  jand g02936(.dina(n3191), .dinb(n3185), .dout(n3192));
  jxor g02937(.dina(n3192), .dinb(n278), .dout(n3193));
  jxor g02938(.dina(n3193), .dinb(n3178), .dout(n3194));
  jxor g02939(.dina(n3194), .dinb(n3036), .dout(f32 ));
  jnot g02940(.din(n3193), .dout(n3196));
  jor  g02941(.dina(n3196), .dinb(n3178), .dout(n3197));
  jor  g02942(.dina(n3194), .dinb(n3036), .dout(n3198));
  jand g02943(.dina(n3198), .dinb(n3197), .dout(n3199));
  jand g02944(.dina(n3176), .dinb(n3168), .dout(n3200));
  jnot g02945(.din(n3200), .dout(n3201));
  jnot g02946(.din(n3177), .dout(n3202));
  jor  g02947(.dina(n3202), .dinb(n3041), .dout(n3203));
  jand g02948(.dina(n3203), .dinb(n3201), .dout(n3204));
  jand g02949(.dina(n3166), .dinb(n3158), .dout(n3205));
  jand g02950(.dina(n3167), .dinb(n3044), .dout(n3206));
  jor  g02951(.dina(n3206), .dinb(n3205), .dout(n3207));
  jand g02952(.dina(n3155), .dinb(n3147), .dout(n3208));
  jnot g02953(.din(n3208), .dout(n3209));
  jor  g02954(.dina(n3157), .dinb(n3048), .dout(n3210));
  jand g02955(.dina(n3210), .dinb(n3209), .dout(n3211));
  jand g02956(.dina(n3145), .dinb(n3137), .dout(n3212));
  jand g02957(.dina(n3146), .dinb(n3051), .dout(n3213));
  jor  g02958(.dina(n3213), .dinb(n3212), .dout(n3214));
  jand g02959(.dina(n3135), .dinb(n3127), .dout(n3215));
  jand g02960(.dina(n3136), .dinb(n3054), .dout(n3216));
  jor  g02961(.dina(n3216), .dinb(n3215), .dout(n3217));
  jand g02962(.dina(n3125), .dinb(n3117), .dout(n3218));
  jand g02963(.dina(n3126), .dinb(n3057), .dout(n3219));
  jor  g02964(.dina(n3219), .dinb(n3218), .dout(n3220));
  jand g02965(.dina(n3115), .dinb(n3107), .dout(n3221));
  jand g02966(.dina(n3116), .dinb(n3060), .dout(n3222));
  jor  g02967(.dina(n3222), .dinb(n3221), .dout(n3223));
  jand g02968(.dina(n3105), .dinb(n3097), .dout(n3224));
  jand g02969(.dina(n3106), .dinb(n3065), .dout(n3225));
  jor  g02970(.dina(n3225), .dinb(n3224), .dout(n3226));
  jor  g02971(.dina(n3095), .dinb(n3087), .dout(n3227));
  jand g02972(.dina(n3096), .dinb(n3070), .dout(n3228));
  jnot g02973(.din(n3228), .dout(n3229));
  jand g02974(.dina(n3229), .dinb(n3227), .dout(n3230));
  jnot g02975(.din(n3230), .dout(n3231));
  jor  g02976(.dina(n3084), .dinb(n3080), .dout(n3232));
  jxor g02977(.dina(a33 ), .dinb(a32 ), .dout(n3233));
  jand g02978(.dina(n3233), .dinb(b0 ), .dout(n3234));
  jnot g02979(.din(n3234), .dout(n3235));
  jxor g02980(.dina(n3235), .dinb(n3232), .dout(n3236));
  jnot g02981(.din(n2914), .dout(n3237));
  jor  g02982(.dina(n3237), .dinb(n303), .dout(n3238));
  jnot g02983(.din(n2907), .dout(n3239));
  jor  g02984(.dina(n3239), .dinb(n301), .dout(n3240));
  jor  g02985(.dina(n3072), .dinb(n305), .dout(n3241));
  jnot g02986(.din(n2911), .dout(n3242));
  jor  g02987(.dina(n3242), .dinb(n293), .dout(n3243));
  jand g02988(.dina(n3243), .dinb(n3241), .dout(n3244));
  jand g02989(.dina(n3244), .dinb(n3240), .dout(n3245));
  jand g02990(.dina(n3245), .dinb(n3238), .dout(n3246));
  jxor g02991(.dina(n3246), .dinb(n2918), .dout(n3247));
  jxor g02992(.dina(n3247), .dinb(n3236), .dout(n3248));
  jnot g02993(.din(n3248), .dout(n3249));
  jor  g02994(.dina(n2764), .dinb(n412), .dout(n3250));
  jor  g02995(.dina(n2766), .dinb(n377), .dout(n3251));
  jor  g02996(.dina(n2609), .dinb(n340), .dout(n3252));
  jand g02997(.dina(n3252), .dinb(n3251), .dout(n3253));
  jor  g02998(.dina(n2761), .dinb(n415), .dout(n3254));
  jand g02999(.dina(n3254), .dinb(n3253), .dout(n3255));
  jand g03000(.dina(n3255), .dinb(n3250), .dout(n3256));
  jxor g03001(.dina(n3256), .dinb(a29 ), .dout(n3257));
  jxor g03002(.dina(n3257), .dinb(n3249), .dout(n3258));
  jxor g03003(.dina(n3258), .dinb(n3231), .dout(n3259));
  jor  g03004(.dina(n2324), .dinb(n570), .dout(n3260));
  jor  g03005(.dina(n2186), .dinb(n469), .dout(n3261));
  jor  g03006(.dina(n2326), .dinb(n572), .dout(n3262));
  jor  g03007(.dina(n2321), .dinb(n519), .dout(n3263));
  jand g03008(.dina(n3263), .dinb(n3262), .dout(n3264));
  jand g03009(.dina(n3264), .dinb(n3261), .dout(n3265));
  jand g03010(.dina(n3265), .dinb(n3260), .dout(n3266));
  jxor g03011(.dina(n3266), .dinb(n2057), .dout(n3267));
  jxor g03012(.dina(n3267), .dinb(n3259), .dout(n3268));
  jxor g03013(.dina(n3268), .dinb(n3226), .dout(n3269));
  jor  g03014(.dina(n1921), .dinb(n770), .dout(n3270));
  jor  g03015(.dina(n1806), .dinb(n637), .dout(n3271));
  jor  g03016(.dina(n1923), .dinb(n772), .dout(n3272));
  jor  g03017(.dina(n1918), .dinb(n704), .dout(n3273));
  jand g03018(.dina(n3273), .dinb(n3272), .dout(n3274));
  jand g03019(.dina(n3274), .dinb(n3271), .dout(n3275));
  jand g03020(.dina(n3275), .dinb(n3270), .dout(n3276));
  jxor g03021(.dina(n3276), .dinb(n1687), .dout(n3277));
  jxor g03022(.dina(n3277), .dinb(n3269), .dout(n3278));
  jxor g03023(.dina(n3278), .dinb(n3223), .dout(n3279));
  jor  g03024(.dina(n1569), .dinb(n1016), .dout(n3280));
  jor  g03025(.dina(n1453), .dinb(n852), .dout(n3281));
  jor  g03026(.dina(n1566), .dinb(n934), .dout(n3282));
  jor  g03027(.dina(n1571), .dinb(n1018), .dout(n3283));
  jand g03028(.dina(n3283), .dinb(n3282), .dout(n3284));
  jand g03029(.dina(n3284), .dinb(n3281), .dout(n3285));
  jand g03030(.dina(n3285), .dinb(n3280), .dout(n3286));
  jxor g03031(.dina(n3286), .dinb(n1351), .dout(n3287));
  jxor g03032(.dina(n3287), .dinb(n3279), .dout(n3288));
  jxor g03033(.dina(n3288), .dinb(n3220), .dout(n3289));
  jor  g03034(.dina(n1305), .dinb(n1248), .dout(n3290));
  jor  g03035(.dina(n1147), .dinb(n1114), .dout(n3291));
  jor  g03036(.dina(n1246), .dinb(n1307), .dout(n3292));
  jor  g03037(.dina(n1251), .dinb(n1211), .dout(n3293));
  jand g03038(.dina(n3293), .dinb(n3292), .dout(n3294));
  jand g03039(.dina(n3294), .dinb(n3291), .dout(n3295));
  jand g03040(.dina(n3295), .dinb(n3290), .dout(n3296));
  jxor g03041(.dina(n3296), .dinb(n1061), .dout(n3297));
  jxor g03042(.dina(n3297), .dinb(n3289), .dout(n3298));
  jxor g03043(.dina(n3298), .dinb(n3217), .dout(n3299));
  jor  g03044(.dina(n1635), .dinb(n970), .dout(n3300));
  jor  g03045(.dina(n880), .dinb(n1416), .dout(n3301));
  jor  g03046(.dina(n967), .dinb(n1527), .dout(n3302));
  jor  g03047(.dina(n972), .dinb(n1637), .dout(n3303));
  jand g03048(.dina(n3303), .dinb(n3302), .dout(n3304));
  jand g03049(.dina(n3304), .dinb(n3301), .dout(n3305));
  jand g03050(.dina(n3305), .dinb(n3300), .dout(n3306));
  jxor g03051(.dina(n3306), .dinb(n810), .dout(n3307));
  jxor g03052(.dina(n3307), .dinb(n3299), .dout(n3308));
  jxor g03053(.dina(n3308), .dinb(n3214), .dout(n3309));
  jor  g03054(.dina(n2005), .dinb(n728), .dout(n3310));
  jor  g03055(.dina(n660), .dinb(n1759), .dout(n3311));
  jor  g03056(.dina(n731), .dinb(n1881), .dout(n3312));
  jor  g03057(.dina(n726), .dinb(n2007), .dout(n3313));
  jand g03058(.dina(n3313), .dinb(n3312), .dout(n3314));
  jand g03059(.dina(n3314), .dinb(n3311), .dout(n3315));
  jand g03060(.dina(n3315), .dinb(n3310), .dout(n3316));
  jxor g03061(.dina(n3316), .dinb(n606), .dout(n3317));
  jxor g03062(.dina(n3317), .dinb(n3309), .dout(n3318));
  jnot g03063(.din(n3318), .dout(n3319));
  jxor g03064(.dina(n3319), .dinb(n3211), .dout(n3320));
  jor  g03065(.dina(n2413), .dinb(n544), .dout(n3321));
  jor  g03066(.dina(n486), .dinb(n2142), .dout(n3322));
  jor  g03067(.dina(n542), .dinb(n2415), .dout(n3323));
  jor  g03068(.dina(n547), .dinb(n2279), .dout(n3324));
  jand g03069(.dina(n3324), .dinb(n3323), .dout(n3325));
  jand g03070(.dina(n3325), .dinb(n3322), .dout(n3326));
  jand g03071(.dina(n3326), .dinb(n3321), .dout(n3327));
  jxor g03072(.dina(n3327), .dinb(n446), .dout(n3328));
  jxor g03073(.dina(n3328), .dinb(n3320), .dout(n3329));
  jxor g03074(.dina(n3329), .dinb(n3207), .dout(n3330));
  jor  g03075(.dina(n2860), .dinb(n397), .dout(n3331));
  jor  g03076(.dina(n354), .dinb(n2563), .dout(n3332));
  jor  g03077(.dina(n394), .dinb(n2713), .dout(n3333));
  jor  g03078(.dina(n399), .dinb(n2862), .dout(n3334));
  jand g03079(.dina(n3334), .dinb(n3333), .dout(n3335));
  jand g03080(.dina(n3335), .dinb(n3332), .dout(n3336));
  jand g03081(.dina(n3336), .dinb(n3331), .dout(n3337));
  jxor g03082(.dina(n3337), .dinb(n364), .dout(n3338));
  jxor g03083(.dina(n3338), .dinb(n3330), .dout(n3339));
  jxor g03084(.dina(n3339), .dinb(n3204), .dout(n3340));
  jand g03085(.dina(b32 ), .dinb(b31 ), .dout(n3341));
  jand g03086(.dina(n3182), .dinb(n3181), .dout(n3342));
  jor  g03087(.dina(n3342), .dinb(n3341), .dout(n3343));
  jxor g03088(.dina(b33 ), .dinb(b32 ), .dout(n3344));
  jnot g03089(.din(n3344), .dout(n3345));
  jxor g03090(.dina(n3345), .dinb(n3343), .dout(n3346));
  jor  g03091(.dina(n3346), .dinb(n296), .dout(n3347));
  jnot g03092(.din(b33 ), .dout(n3348));
  jor  g03093(.dina(n264), .dinb(n3348), .dout(n3349));
  jor  g03094(.dina(n280), .dinb(n3023), .dout(n3350));
  jor  g03095(.dina(n294), .dinb(n3186), .dout(n3351));
  jand g03096(.dina(n3351), .dinb(n3350), .dout(n3352));
  jand g03097(.dina(n3352), .dinb(n3349), .dout(n3353));
  jand g03098(.dina(n3353), .dinb(n3347), .dout(n3354));
  jxor g03099(.dina(n3354), .dinb(n278), .dout(n3355));
  jxor g03100(.dina(n3355), .dinb(n3340), .dout(n3356));
  jxor g03101(.dina(n3356), .dinb(n3199), .dout(f33 ));
  jnot g03102(.din(n3355), .dout(n3358));
  jor  g03103(.dina(n3358), .dinb(n3340), .dout(n3359));
  jor  g03104(.dina(n3356), .dinb(n3199), .dout(n3360));
  jand g03105(.dina(n3360), .dinb(n3359), .dout(n3361));
  jand g03106(.dina(n3338), .dinb(n3330), .dout(n3362));
  jnot g03107(.din(n3362), .dout(n3363));
  jnot g03108(.din(n3339), .dout(n3364));
  jor  g03109(.dina(n3364), .dinb(n3204), .dout(n3365));
  jand g03110(.dina(n3365), .dinb(n3363), .dout(n3366));
  jand g03111(.dina(n3328), .dinb(n3320), .dout(n3367));
  jand g03112(.dina(n3329), .dinb(n3207), .dout(n3368));
  jor  g03113(.dina(n3368), .dinb(n3367), .dout(n3369));
  jand g03114(.dina(n3317), .dinb(n3309), .dout(n3370));
  jnot g03115(.din(n3370), .dout(n3371));
  jor  g03116(.dina(n3319), .dinb(n3211), .dout(n3372));
  jand g03117(.dina(n3372), .dinb(n3371), .dout(n3373));
  jand g03118(.dina(n3307), .dinb(n3299), .dout(n3374));
  jand g03119(.dina(n3308), .dinb(n3214), .dout(n3375));
  jor  g03120(.dina(n3375), .dinb(n3374), .dout(n3376));
  jand g03121(.dina(n3297), .dinb(n3289), .dout(n3377));
  jand g03122(.dina(n3298), .dinb(n3217), .dout(n3378));
  jor  g03123(.dina(n3378), .dinb(n3377), .dout(n3379));
  jand g03124(.dina(n3287), .dinb(n3279), .dout(n3380));
  jand g03125(.dina(n3288), .dinb(n3220), .dout(n3381));
  jor  g03126(.dina(n3381), .dinb(n3380), .dout(n3382));
  jand g03127(.dina(n3277), .dinb(n3269), .dout(n3383));
  jand g03128(.dina(n3278), .dinb(n3223), .dout(n3384));
  jor  g03129(.dina(n3384), .dinb(n3383), .dout(n3385));
  jand g03130(.dina(n3267), .dinb(n3259), .dout(n3386));
  jand g03131(.dina(n3268), .dinb(n3226), .dout(n3387));
  jor  g03132(.dina(n3387), .dinb(n3386), .dout(n3388));
  jor  g03133(.dina(n3257), .dinb(n3249), .dout(n3389));
  jand g03134(.dina(n3258), .dinb(n3231), .dout(n3390));
  jnot g03135(.din(n3390), .dout(n3391));
  jand g03136(.dina(n3391), .dinb(n3389), .dout(n3392));
  jnot g03137(.din(n3392), .dout(n3393));
  jnot g03138(.din(n3232), .dout(n3394));
  jand g03139(.dina(n3234), .dinb(n3394), .dout(n3395));
  jand g03140(.dina(n3247), .dinb(n3236), .dout(n3396));
  jor  g03141(.dina(n3396), .dinb(n3395), .dout(n3397));
  jxor g03142(.dina(a35 ), .dinb(a34 ), .dout(n3398));
  jand g03143(.dina(n3398), .dinb(n3233), .dout(n3399));
  jand g03144(.dina(n3399), .dinb(n259), .dout(n3400));
  jnot g03145(.din(n3233), .dout(n3401));
  jxor g03146(.dina(a34 ), .dinb(a33 ), .dout(n3402));
  jand g03147(.dina(n3402), .dinb(n3401), .dout(n3403));
  jand g03148(.dina(n3403), .dinb(b0 ), .dout(n3404));
  jnot g03149(.din(n3398), .dout(n3405));
  jand g03150(.dina(n3405), .dinb(n3233), .dout(n3406));
  jand g03151(.dina(n3406), .dinb(b1 ), .dout(n3407));
  jor  g03152(.dina(n3407), .dinb(n3404), .dout(n3408));
  jor  g03153(.dina(n3408), .dinb(n3400), .dout(n3409));
  jnot g03154(.din(a35 ), .dout(n3410));
  jor  g03155(.dina(n3235), .dinb(n3410), .dout(n3411));
  jxor g03156(.dina(n3411), .dinb(n3409), .dout(n3412));
  jor  g03157(.dina(n3239), .dinb(n337), .dout(n3413));
  jor  g03158(.dina(n3237), .dinb(n340), .dout(n3414));
  jor  g03159(.dina(n3072), .dinb(n293), .dout(n3415));
  jand g03160(.dina(n3415), .dinb(n3414), .dout(n3416));
  jor  g03161(.dina(n3242), .dinb(n303), .dout(n3417));
  jand g03162(.dina(n3417), .dinb(n3416), .dout(n3418));
  jand g03163(.dina(n3418), .dinb(n3413), .dout(n3419));
  jxor g03164(.dina(n3419), .dinb(a32 ), .dout(n3420));
  jxor g03165(.dina(n3420), .dinb(n3412), .dout(n3421));
  jxor g03166(.dina(n3421), .dinb(n3397), .dout(n3422));
  jnot g03167(.din(n3422), .dout(n3423));
  jor  g03168(.dina(n2764), .dinb(n466), .dout(n3424));
  jor  g03169(.dina(n2766), .dinb(n415), .dout(n3425));
  jor  g03170(.dina(n2609), .dinb(n377), .dout(n3426));
  jand g03171(.dina(n3426), .dinb(n3425), .dout(n3427));
  jor  g03172(.dina(n2761), .dinb(n469), .dout(n3428));
  jand g03173(.dina(n3428), .dinb(n3427), .dout(n3429));
  jand g03174(.dina(n3429), .dinb(n3424), .dout(n3430));
  jxor g03175(.dina(n3430), .dinb(a29 ), .dout(n3431));
  jxor g03176(.dina(n3431), .dinb(n3423), .dout(n3432));
  jxor g03177(.dina(n3432), .dinb(n3393), .dout(n3433));
  jor  g03178(.dina(n2324), .dinb(n635), .dout(n3434));
  jor  g03179(.dina(n2186), .dinb(n519), .dout(n3435));
  jor  g03180(.dina(n2326), .dinb(n637), .dout(n3436));
  jor  g03181(.dina(n2321), .dinb(n572), .dout(n3437));
  jand g03182(.dina(n3437), .dinb(n3436), .dout(n3438));
  jand g03183(.dina(n3438), .dinb(n3435), .dout(n3439));
  jand g03184(.dina(n3439), .dinb(n3434), .dout(n3440));
  jxor g03185(.dina(n3440), .dinb(n2057), .dout(n3441));
  jxor g03186(.dina(n3441), .dinb(n3433), .dout(n3442));
  jxor g03187(.dina(n3442), .dinb(n3388), .dout(n3443));
  jor  g03188(.dina(n1921), .dinb(n850), .dout(n3444));
  jor  g03189(.dina(n1806), .dinb(n704), .dout(n3445));
  jor  g03190(.dina(n1923), .dinb(n852), .dout(n3446));
  jor  g03191(.dina(n1918), .dinb(n772), .dout(n3447));
  jand g03192(.dina(n3447), .dinb(n3446), .dout(n3448));
  jand g03193(.dina(n3448), .dinb(n3445), .dout(n3449));
  jand g03194(.dina(n3449), .dinb(n3444), .dout(n3450));
  jxor g03195(.dina(n3450), .dinb(n1687), .dout(n3451));
  jxor g03196(.dina(n3451), .dinb(n3443), .dout(n3452));
  jxor g03197(.dina(n3452), .dinb(n3385), .dout(n3453));
  jor  g03198(.dina(n1569), .dinb(n1112), .dout(n3454));
  jor  g03199(.dina(n1453), .dinb(n934), .dout(n3455));
  jor  g03200(.dina(n1566), .dinb(n1018), .dout(n3456));
  jor  g03201(.dina(n1571), .dinb(n1114), .dout(n3457));
  jand g03202(.dina(n3457), .dinb(n3456), .dout(n3458));
  jand g03203(.dina(n3458), .dinb(n3455), .dout(n3459));
  jand g03204(.dina(n3459), .dinb(n3454), .dout(n3460));
  jxor g03205(.dina(n3460), .dinb(n1351), .dout(n3461));
  jxor g03206(.dina(n3461), .dinb(n3453), .dout(n3462));
  jxor g03207(.dina(n3462), .dinb(n3382), .dout(n3463));
  jor  g03208(.dina(n1414), .dinb(n1248), .dout(n3464));
  jor  g03209(.dina(n1147), .dinb(n1211), .dout(n3465));
  jor  g03210(.dina(n1246), .dinb(n1416), .dout(n3466));
  jor  g03211(.dina(n1251), .dinb(n1307), .dout(n3467));
  jand g03212(.dina(n3467), .dinb(n3466), .dout(n3468));
  jand g03213(.dina(n3468), .dinb(n3465), .dout(n3469));
  jand g03214(.dina(n3469), .dinb(n3464), .dout(n3470));
  jxor g03215(.dina(n3470), .dinb(n1061), .dout(n3471));
  jxor g03216(.dina(n3471), .dinb(n3463), .dout(n3472));
  jxor g03217(.dina(n3472), .dinb(n3379), .dout(n3473));
  jor  g03218(.dina(n1757), .dinb(n970), .dout(n3474));
  jor  g03219(.dina(n880), .dinb(n1527), .dout(n3475));
  jor  g03220(.dina(n967), .dinb(n1637), .dout(n3476));
  jor  g03221(.dina(n972), .dinb(n1759), .dout(n3477));
  jand g03222(.dina(n3477), .dinb(n3476), .dout(n3478));
  jand g03223(.dina(n3478), .dinb(n3475), .dout(n3479));
  jand g03224(.dina(n3479), .dinb(n3474), .dout(n3480));
  jxor g03225(.dina(n3480), .dinb(n810), .dout(n3481));
  jxor g03226(.dina(n3481), .dinb(n3473), .dout(n3482));
  jxor g03227(.dina(n3482), .dinb(n3376), .dout(n3483));
  jor  g03228(.dina(n2140), .dinb(n728), .dout(n3484));
  jor  g03229(.dina(n660), .dinb(n1881), .dout(n3485));
  jor  g03230(.dina(n731), .dinb(n2007), .dout(n3486));
  jor  g03231(.dina(n726), .dinb(n2142), .dout(n3487));
  jand g03232(.dina(n3487), .dinb(n3486), .dout(n3488));
  jand g03233(.dina(n3488), .dinb(n3485), .dout(n3489));
  jand g03234(.dina(n3489), .dinb(n3484), .dout(n3490));
  jxor g03235(.dina(n3490), .dinb(n606), .dout(n3491));
  jxor g03236(.dina(n3491), .dinb(n3483), .dout(n3492));
  jnot g03237(.din(n3492), .dout(n3493));
  jxor g03238(.dina(n3493), .dinb(n3373), .dout(n3494));
  jor  g03239(.dina(n2561), .dinb(n544), .dout(n3495));
  jor  g03240(.dina(n486), .dinb(n2279), .dout(n3496));
  jor  g03241(.dina(n547), .dinb(n2415), .dout(n3497));
  jor  g03242(.dina(n542), .dinb(n2563), .dout(n3498));
  jand g03243(.dina(n3498), .dinb(n3497), .dout(n3499));
  jand g03244(.dina(n3499), .dinb(n3496), .dout(n3500));
  jand g03245(.dina(n3500), .dinb(n3495), .dout(n3501));
  jxor g03246(.dina(n3501), .dinb(n446), .dout(n3502));
  jxor g03247(.dina(n3502), .dinb(n3494), .dout(n3503));
  jxor g03248(.dina(n3503), .dinb(n3369), .dout(n3504));
  jor  g03249(.dina(n3021), .dinb(n397), .dout(n3505));
  jor  g03250(.dina(n354), .dinb(n2713), .dout(n3506));
  jor  g03251(.dina(n399), .dinb(n3023), .dout(n3507));
  jor  g03252(.dina(n394), .dinb(n2862), .dout(n3508));
  jand g03253(.dina(n3508), .dinb(n3507), .dout(n3509));
  jand g03254(.dina(n3509), .dinb(n3506), .dout(n3510));
  jand g03255(.dina(n3510), .dinb(n3505), .dout(n3511));
  jxor g03256(.dina(n3511), .dinb(n364), .dout(n3512));
  jxor g03257(.dina(n3512), .dinb(n3504), .dout(n3513));
  jxor g03258(.dina(n3513), .dinb(n3366), .dout(n3514));
  jand g03259(.dina(b33 ), .dinb(b32 ), .dout(n3515));
  jand g03260(.dina(n3344), .dinb(n3343), .dout(n3516));
  jor  g03261(.dina(n3516), .dinb(n3515), .dout(n3517));
  jxor g03262(.dina(b34 ), .dinb(b33 ), .dout(n3518));
  jnot g03263(.din(n3518), .dout(n3519));
  jxor g03264(.dina(n3519), .dinb(n3517), .dout(n3520));
  jor  g03265(.dina(n3520), .dinb(n296), .dout(n3521));
  jnot g03266(.din(b34 ), .dout(n3522));
  jor  g03267(.dina(n264), .dinb(n3522), .dout(n3523));
  jor  g03268(.dina(n280), .dinb(n3186), .dout(n3524));
  jor  g03269(.dina(n294), .dinb(n3348), .dout(n3525));
  jand g03270(.dina(n3525), .dinb(n3524), .dout(n3526));
  jand g03271(.dina(n3526), .dinb(n3523), .dout(n3527));
  jand g03272(.dina(n3527), .dinb(n3521), .dout(n3528));
  jxor g03273(.dina(n3528), .dinb(n278), .dout(n3529));
  jxor g03274(.dina(n3529), .dinb(n3514), .dout(n3530));
  jxor g03275(.dina(n3530), .dinb(n3361), .dout(f34 ));
  jnot g03276(.din(n3529), .dout(n3532));
  jor  g03277(.dina(n3532), .dinb(n3514), .dout(n3533));
  jor  g03278(.dina(n3530), .dinb(n3361), .dout(n3534));
  jand g03279(.dina(n3534), .dinb(n3533), .dout(n3535));
  jand g03280(.dina(n3512), .dinb(n3504), .dout(n3536));
  jnot g03281(.din(n3536), .dout(n3537));
  jnot g03282(.din(n3513), .dout(n3538));
  jor  g03283(.dina(n3538), .dinb(n3366), .dout(n3539));
  jand g03284(.dina(n3539), .dinb(n3537), .dout(n3540));
  jand g03285(.dina(n3502), .dinb(n3494), .dout(n3541));
  jand g03286(.dina(n3503), .dinb(n3369), .dout(n3542));
  jor  g03287(.dina(n3542), .dinb(n3541), .dout(n3543));
  jand g03288(.dina(n3491), .dinb(n3483), .dout(n3544));
  jnot g03289(.din(n3544), .dout(n3545));
  jor  g03290(.dina(n3493), .dinb(n3373), .dout(n3546));
  jand g03291(.dina(n3546), .dinb(n3545), .dout(n3547));
  jand g03292(.dina(n3481), .dinb(n3473), .dout(n3548));
  jand g03293(.dina(n3482), .dinb(n3376), .dout(n3549));
  jor  g03294(.dina(n3549), .dinb(n3548), .dout(n3550));
  jand g03295(.dina(n3471), .dinb(n3463), .dout(n3551));
  jand g03296(.dina(n3472), .dinb(n3379), .dout(n3552));
  jor  g03297(.dina(n3552), .dinb(n3551), .dout(n3553));
  jand g03298(.dina(n3461), .dinb(n3453), .dout(n3554));
  jand g03299(.dina(n3462), .dinb(n3382), .dout(n3555));
  jor  g03300(.dina(n3555), .dinb(n3554), .dout(n3556));
  jand g03301(.dina(n3451), .dinb(n3443), .dout(n3557));
  jand g03302(.dina(n3452), .dinb(n3385), .dout(n3558));
  jor  g03303(.dina(n3558), .dinb(n3557), .dout(n3559));
  jand g03304(.dina(n3441), .dinb(n3433), .dout(n3560));
  jand g03305(.dina(n3442), .dinb(n3388), .dout(n3561));
  jor  g03306(.dina(n3561), .dinb(n3560), .dout(n3562));
  jor  g03307(.dina(n3431), .dinb(n3423), .dout(n3563));
  jand g03308(.dina(n3432), .dinb(n3393), .dout(n3564));
  jnot g03309(.din(n3564), .dout(n3565));
  jand g03310(.dina(n3565), .dinb(n3563), .dout(n3566));
  jnot g03311(.din(n3566), .dout(n3567));
  jor  g03312(.dina(n3420), .dinb(n3412), .dout(n3568));
  jand g03313(.dina(n3421), .dinb(n3397), .dout(n3569));
  jnot g03314(.din(n3569), .dout(n3570));
  jand g03315(.dina(n3570), .dinb(n3568), .dout(n3571));
  jnot g03316(.din(n3571), .dout(n3572));
  jor  g03317(.dina(n3402), .dinb(n3233), .dout(n3573));
  jor  g03318(.dina(n3573), .dinb(n3405), .dout(n3574));
  jnot g03319(.din(n3574), .dout(n3575));
  jand g03320(.dina(n3575), .dinb(b0 ), .dout(n3576));
  jand g03321(.dina(n3406), .dinb(b2 ), .dout(n3577));
  jor  g03322(.dina(n3577), .dinb(n3576), .dout(n3578));
  jand g03323(.dina(n3399), .dinb(n273), .dout(n3579));
  jand g03324(.dina(n3403), .dinb(b1 ), .dout(n3580));
  jor  g03325(.dina(n3580), .dinb(n3579), .dout(n3581));
  jor  g03326(.dina(n3581), .dinb(n3578), .dout(n3582));
  jnot g03327(.din(n3409), .dout(n3583));
  jand g03328(.dina(n3235), .dinb(a35 ), .dout(n3584));
  jand g03329(.dina(n3584), .dinb(n3583), .dout(n3585));
  jnot g03330(.din(n3585), .dout(n3586));
  jand g03331(.dina(n3586), .dinb(a35 ), .dout(n3587));
  jxor g03332(.dina(n3587), .dinb(n3582), .dout(n3588));
  jnot g03333(.din(n3588), .dout(n3589));
  jor  g03334(.dina(n3239), .dinb(n374), .dout(n3590));
  jor  g03335(.dina(n3242), .dinb(n340), .dout(n3591));
  jor  g03336(.dina(n3072), .dinb(n303), .dout(n3592));
  jand g03337(.dina(n3592), .dinb(n3591), .dout(n3593));
  jor  g03338(.dina(n3237), .dinb(n377), .dout(n3594));
  jand g03339(.dina(n3594), .dinb(n3593), .dout(n3595));
  jand g03340(.dina(n3595), .dinb(n3590), .dout(n3596));
  jxor g03341(.dina(n3596), .dinb(a32 ), .dout(n3597));
  jxor g03342(.dina(n3597), .dinb(n3589), .dout(n3598));
  jxor g03343(.dina(n3598), .dinb(n3572), .dout(n3599));
  jor  g03344(.dina(n2764), .dinb(n517), .dout(n3600));
  jor  g03345(.dina(n2766), .dinb(n469), .dout(n3601));
  jor  g03346(.dina(n2761), .dinb(n519), .dout(n3602));
  jor  g03347(.dina(n2609), .dinb(n415), .dout(n3603));
  jand g03348(.dina(n3603), .dinb(n3602), .dout(n3604));
  jand g03349(.dina(n3604), .dinb(n3601), .dout(n3605));
  jand g03350(.dina(n3605), .dinb(n3600), .dout(n3606));
  jxor g03351(.dina(n3606), .dinb(n2468), .dout(n3607));
  jxor g03352(.dina(n3607), .dinb(n3599), .dout(n3608));
  jxor g03353(.dina(n3608), .dinb(n3567), .dout(n3609));
  jor  g03354(.dina(n2324), .dinb(n702), .dout(n3610));
  jor  g03355(.dina(n2186), .dinb(n572), .dout(n3611));
  jor  g03356(.dina(n2326), .dinb(n704), .dout(n3612));
  jor  g03357(.dina(n2321), .dinb(n637), .dout(n3613));
  jand g03358(.dina(n3613), .dinb(n3612), .dout(n3614));
  jand g03359(.dina(n3614), .dinb(n3611), .dout(n3615));
  jand g03360(.dina(n3615), .dinb(n3610), .dout(n3616));
  jxor g03361(.dina(n3616), .dinb(n2057), .dout(n3617));
  jxor g03362(.dina(n3617), .dinb(n3609), .dout(n3618));
  jxor g03363(.dina(n3618), .dinb(n3562), .dout(n3619));
  jor  g03364(.dina(n1921), .dinb(n932), .dout(n3620));
  jor  g03365(.dina(n1806), .dinb(n772), .dout(n3621));
  jor  g03366(.dina(n1918), .dinb(n852), .dout(n3622));
  jor  g03367(.dina(n1923), .dinb(n934), .dout(n3623));
  jand g03368(.dina(n3623), .dinb(n3622), .dout(n3624));
  jand g03369(.dina(n3624), .dinb(n3621), .dout(n3625));
  jand g03370(.dina(n3625), .dinb(n3620), .dout(n3626));
  jxor g03371(.dina(n3626), .dinb(n1687), .dout(n3627));
  jxor g03372(.dina(n3627), .dinb(n3619), .dout(n3628));
  jxor g03373(.dina(n3628), .dinb(n3559), .dout(n3629));
  jor  g03374(.dina(n1569), .dinb(n1209), .dout(n3630));
  jor  g03375(.dina(n1453), .dinb(n1018), .dout(n3631));
  jor  g03376(.dina(n1566), .dinb(n1114), .dout(n3632));
  jor  g03377(.dina(n1571), .dinb(n1211), .dout(n3633));
  jand g03378(.dina(n3633), .dinb(n3632), .dout(n3634));
  jand g03379(.dina(n3634), .dinb(n3631), .dout(n3635));
  jand g03380(.dina(n3635), .dinb(n3630), .dout(n3636));
  jxor g03381(.dina(n3636), .dinb(n1351), .dout(n3637));
  jxor g03382(.dina(n3637), .dinb(n3629), .dout(n3638));
  jxor g03383(.dina(n3638), .dinb(n3556), .dout(n3639));
  jor  g03384(.dina(n1525), .dinb(n1248), .dout(n3640));
  jor  g03385(.dina(n1147), .dinb(n1307), .dout(n3641));
  jor  g03386(.dina(n1246), .dinb(n1527), .dout(n3642));
  jor  g03387(.dina(n1251), .dinb(n1416), .dout(n3643));
  jand g03388(.dina(n3643), .dinb(n3642), .dout(n3644));
  jand g03389(.dina(n3644), .dinb(n3641), .dout(n3645));
  jand g03390(.dina(n3645), .dinb(n3640), .dout(n3646));
  jxor g03391(.dina(n3646), .dinb(n1061), .dout(n3647));
  jxor g03392(.dina(n3647), .dinb(n3639), .dout(n3648));
  jxor g03393(.dina(n3648), .dinb(n3553), .dout(n3649));
  jor  g03394(.dina(n1879), .dinb(n970), .dout(n3650));
  jor  g03395(.dina(n880), .dinb(n1637), .dout(n3651));
  jor  g03396(.dina(n967), .dinb(n1759), .dout(n3652));
  jor  g03397(.dina(n972), .dinb(n1881), .dout(n3653));
  jand g03398(.dina(n3653), .dinb(n3652), .dout(n3654));
  jand g03399(.dina(n3654), .dinb(n3651), .dout(n3655));
  jand g03400(.dina(n3655), .dinb(n3650), .dout(n3656));
  jxor g03401(.dina(n3656), .dinb(n810), .dout(n3657));
  jxor g03402(.dina(n3657), .dinb(n3649), .dout(n3658));
  jxor g03403(.dina(n3658), .dinb(n3550), .dout(n3659));
  jor  g03404(.dina(n2277), .dinb(n728), .dout(n3660));
  jor  g03405(.dina(n660), .dinb(n2007), .dout(n3661));
  jor  g03406(.dina(n726), .dinb(n2279), .dout(n3662));
  jor  g03407(.dina(n731), .dinb(n2142), .dout(n3663));
  jand g03408(.dina(n3663), .dinb(n3662), .dout(n3664));
  jand g03409(.dina(n3664), .dinb(n3661), .dout(n3665));
  jand g03410(.dina(n3665), .dinb(n3660), .dout(n3666));
  jxor g03411(.dina(n3666), .dinb(n606), .dout(n3667));
  jxor g03412(.dina(n3667), .dinb(n3659), .dout(n3668));
  jnot g03413(.din(n3668), .dout(n3669));
  jxor g03414(.dina(n3669), .dinb(n3547), .dout(n3670));
  jor  g03415(.dina(n2711), .dinb(n544), .dout(n3671));
  jor  g03416(.dina(n486), .dinb(n2415), .dout(n3672));
  jor  g03417(.dina(n547), .dinb(n2563), .dout(n3673));
  jor  g03418(.dina(n542), .dinb(n2713), .dout(n3674));
  jand g03419(.dina(n3674), .dinb(n3673), .dout(n3675));
  jand g03420(.dina(n3675), .dinb(n3672), .dout(n3676));
  jand g03421(.dina(n3676), .dinb(n3671), .dout(n3677));
  jxor g03422(.dina(n3677), .dinb(n446), .dout(n3678));
  jxor g03423(.dina(n3678), .dinb(n3670), .dout(n3679));
  jxor g03424(.dina(n3679), .dinb(n3543), .dout(n3680));
  jor  g03425(.dina(n3184), .dinb(n397), .dout(n3681));
  jor  g03426(.dina(n354), .dinb(n2862), .dout(n3682));
  jor  g03427(.dina(n394), .dinb(n3023), .dout(n3683));
  jor  g03428(.dina(n399), .dinb(n3186), .dout(n3684));
  jand g03429(.dina(n3684), .dinb(n3683), .dout(n3685));
  jand g03430(.dina(n3685), .dinb(n3682), .dout(n3686));
  jand g03431(.dina(n3686), .dinb(n3681), .dout(n3687));
  jxor g03432(.dina(n3687), .dinb(n364), .dout(n3688));
  jxor g03433(.dina(n3688), .dinb(n3680), .dout(n3689));
  jxor g03434(.dina(n3689), .dinb(n3540), .dout(n3690));
  jand g03435(.dina(b34 ), .dinb(b33 ), .dout(n3691));
  jand g03436(.dina(n3518), .dinb(n3517), .dout(n3692));
  jor  g03437(.dina(n3692), .dinb(n3691), .dout(n3693));
  jxor g03438(.dina(b35 ), .dinb(b34 ), .dout(n3694));
  jnot g03439(.din(n3694), .dout(n3695));
  jxor g03440(.dina(n3695), .dinb(n3693), .dout(n3696));
  jor  g03441(.dina(n3696), .dinb(n296), .dout(n3697));
  jnot g03442(.din(b35 ), .dout(n3698));
  jor  g03443(.dina(n264), .dinb(n3698), .dout(n3699));
  jor  g03444(.dina(n280), .dinb(n3348), .dout(n3700));
  jor  g03445(.dina(n294), .dinb(n3522), .dout(n3701));
  jand g03446(.dina(n3701), .dinb(n3700), .dout(n3702));
  jand g03447(.dina(n3702), .dinb(n3699), .dout(n3703));
  jand g03448(.dina(n3703), .dinb(n3697), .dout(n3704));
  jxor g03449(.dina(n3704), .dinb(n278), .dout(n3705));
  jxor g03450(.dina(n3705), .dinb(n3690), .dout(n3706));
  jxor g03451(.dina(n3706), .dinb(n3535), .dout(f35 ));
  jnot g03452(.din(n3705), .dout(n3708));
  jor  g03453(.dina(n3708), .dinb(n3690), .dout(n3709));
  jor  g03454(.dina(n3706), .dinb(n3535), .dout(n3710));
  jand g03455(.dina(n3710), .dinb(n3709), .dout(n3711));
  jand g03456(.dina(n3688), .dinb(n3680), .dout(n3712));
  jnot g03457(.din(n3712), .dout(n3713));
  jnot g03458(.din(n3689), .dout(n3714));
  jor  g03459(.dina(n3714), .dinb(n3540), .dout(n3715));
  jand g03460(.dina(n3715), .dinb(n3713), .dout(n3716));
  jand g03461(.dina(n3678), .dinb(n3670), .dout(n3717));
  jand g03462(.dina(n3679), .dinb(n3543), .dout(n3718));
  jor  g03463(.dina(n3718), .dinb(n3717), .dout(n3719));
  jand g03464(.dina(n3667), .dinb(n3659), .dout(n3720));
  jnot g03465(.din(n3720), .dout(n3721));
  jor  g03466(.dina(n3669), .dinb(n3547), .dout(n3722));
  jand g03467(.dina(n3722), .dinb(n3721), .dout(n3723));
  jand g03468(.dina(n3657), .dinb(n3649), .dout(n3724));
  jand g03469(.dina(n3658), .dinb(n3550), .dout(n3725));
  jor  g03470(.dina(n3725), .dinb(n3724), .dout(n3726));
  jand g03471(.dina(n3647), .dinb(n3639), .dout(n3727));
  jand g03472(.dina(n3648), .dinb(n3553), .dout(n3728));
  jor  g03473(.dina(n3728), .dinb(n3727), .dout(n3729));
  jand g03474(.dina(n3637), .dinb(n3629), .dout(n3730));
  jand g03475(.dina(n3638), .dinb(n3556), .dout(n3731));
  jor  g03476(.dina(n3731), .dinb(n3730), .dout(n3732));
  jand g03477(.dina(n3627), .dinb(n3619), .dout(n3733));
  jand g03478(.dina(n3628), .dinb(n3559), .dout(n3734));
  jor  g03479(.dina(n3734), .dinb(n3733), .dout(n3735));
  jand g03480(.dina(n3607), .dinb(n3599), .dout(n3736));
  jand g03481(.dina(n3608), .dinb(n3567), .dout(n3737));
  jor  g03482(.dina(n3737), .dinb(n3736), .dout(n3738));
  jor  g03483(.dina(n3597), .dinb(n3589), .dout(n3739));
  jand g03484(.dina(n3598), .dinb(n3572), .dout(n3740));
  jnot g03485(.din(n3740), .dout(n3741));
  jand g03486(.dina(n3741), .dinb(n3739), .dout(n3742));
  jnot g03487(.din(n3742), .dout(n3743));
  jor  g03488(.dina(n3586), .dinb(n3582), .dout(n3744));
  jxor g03489(.dina(a36 ), .dinb(a35 ), .dout(n3745));
  jand g03490(.dina(n3745), .dinb(b0 ), .dout(n3746));
  jnot g03491(.din(n3746), .dout(n3747));
  jxor g03492(.dina(n3747), .dinb(n3744), .dout(n3748));
  jnot g03493(.din(n3406), .dout(n3749));
  jor  g03494(.dina(n3749), .dinb(n303), .dout(n3750));
  jnot g03495(.din(n3399), .dout(n3751));
  jor  g03496(.dina(n3751), .dinb(n301), .dout(n3752));
  jor  g03497(.dina(n3574), .dinb(n305), .dout(n3753));
  jnot g03498(.din(n3403), .dout(n3754));
  jor  g03499(.dina(n3754), .dinb(n293), .dout(n3755));
  jand g03500(.dina(n3755), .dinb(n3753), .dout(n3756));
  jand g03501(.dina(n3756), .dinb(n3752), .dout(n3757));
  jand g03502(.dina(n3757), .dinb(n3750), .dout(n3758));
  jxor g03503(.dina(n3758), .dinb(n3410), .dout(n3759));
  jxor g03504(.dina(n3759), .dinb(n3748), .dout(n3760));
  jnot g03505(.din(n3760), .dout(n3761));
  jor  g03506(.dina(n3239), .dinb(n412), .dout(n3762));
  jor  g03507(.dina(n3237), .dinb(n415), .dout(n3763));
  jor  g03508(.dina(n3072), .dinb(n340), .dout(n3764));
  jand g03509(.dina(n3764), .dinb(n3763), .dout(n3765));
  jor  g03510(.dina(n3242), .dinb(n377), .dout(n3766));
  jand g03511(.dina(n3766), .dinb(n3765), .dout(n3767));
  jand g03512(.dina(n3767), .dinb(n3762), .dout(n3768));
  jxor g03513(.dina(n3768), .dinb(a32 ), .dout(n3769));
  jxor g03514(.dina(n3769), .dinb(n3761), .dout(n3770));
  jxor g03515(.dina(n3770), .dinb(n3743), .dout(n3771));
  jor  g03516(.dina(n2764), .dinb(n570), .dout(n3772));
  jor  g03517(.dina(n2609), .dinb(n469), .dout(n3773));
  jor  g03518(.dina(n2761), .dinb(n572), .dout(n3774));
  jor  g03519(.dina(n2766), .dinb(n519), .dout(n3775));
  jand g03520(.dina(n3775), .dinb(n3774), .dout(n3776));
  jand g03521(.dina(n3776), .dinb(n3773), .dout(n3777));
  jand g03522(.dina(n3777), .dinb(n3772), .dout(n3778));
  jxor g03523(.dina(n3778), .dinb(n2468), .dout(n3779));
  jxor g03524(.dina(n3779), .dinb(n3771), .dout(n3780));
  jxor g03525(.dina(n3780), .dinb(n3738), .dout(n3781));
  jor  g03526(.dina(n2324), .dinb(n770), .dout(n3782));
  jor  g03527(.dina(n2186), .dinb(n637), .dout(n3783));
  jor  g03528(.dina(n2326), .dinb(n772), .dout(n3784));
  jor  g03529(.dina(n2321), .dinb(n704), .dout(n3785));
  jand g03530(.dina(n3785), .dinb(n3784), .dout(n3786));
  jand g03531(.dina(n3786), .dinb(n3783), .dout(n3787));
  jand g03532(.dina(n3787), .dinb(n3782), .dout(n3788));
  jxor g03533(.dina(n3788), .dinb(n2057), .dout(n3789));
  jxor g03534(.dina(n3789), .dinb(n3781), .dout(n3790));
  jand g03535(.dina(n3617), .dinb(n3609), .dout(n3791));
  jand g03536(.dina(n3618), .dinb(n3562), .dout(n3792));
  jor  g03537(.dina(n3792), .dinb(n3791), .dout(n3793));
  jxor g03538(.dina(n3793), .dinb(n3790), .dout(n3794));
  jor  g03539(.dina(n1921), .dinb(n1016), .dout(n3795));
  jor  g03540(.dina(n1806), .dinb(n852), .dout(n3796));
  jor  g03541(.dina(n1918), .dinb(n934), .dout(n3797));
  jor  g03542(.dina(n1923), .dinb(n1018), .dout(n3798));
  jand g03543(.dina(n3798), .dinb(n3797), .dout(n3799));
  jand g03544(.dina(n3799), .dinb(n3796), .dout(n3800));
  jand g03545(.dina(n3800), .dinb(n3795), .dout(n3801));
  jxor g03546(.dina(n3801), .dinb(n1687), .dout(n3802));
  jxor g03547(.dina(n3802), .dinb(n3794), .dout(n3803));
  jxor g03548(.dina(n3803), .dinb(n3735), .dout(n3804));
  jor  g03549(.dina(n1569), .dinb(n1305), .dout(n3805));
  jor  g03550(.dina(n1453), .dinb(n1114), .dout(n3806));
  jor  g03551(.dina(n1571), .dinb(n1307), .dout(n3807));
  jor  g03552(.dina(n1566), .dinb(n1211), .dout(n3808));
  jand g03553(.dina(n3808), .dinb(n3807), .dout(n3809));
  jand g03554(.dina(n3809), .dinb(n3806), .dout(n3810));
  jand g03555(.dina(n3810), .dinb(n3805), .dout(n3811));
  jxor g03556(.dina(n3811), .dinb(n1351), .dout(n3812));
  jxor g03557(.dina(n3812), .dinb(n3804), .dout(n3813));
  jxor g03558(.dina(n3813), .dinb(n3732), .dout(n3814));
  jor  g03559(.dina(n1635), .dinb(n1248), .dout(n3815));
  jor  g03560(.dina(n1147), .dinb(n1416), .dout(n3816));
  jor  g03561(.dina(n1251), .dinb(n1527), .dout(n3817));
  jor  g03562(.dina(n1246), .dinb(n1637), .dout(n3818));
  jand g03563(.dina(n3818), .dinb(n3817), .dout(n3819));
  jand g03564(.dina(n3819), .dinb(n3816), .dout(n3820));
  jand g03565(.dina(n3820), .dinb(n3815), .dout(n3821));
  jxor g03566(.dina(n3821), .dinb(n1061), .dout(n3822));
  jxor g03567(.dina(n3822), .dinb(n3814), .dout(n3823));
  jxor g03568(.dina(n3823), .dinb(n3729), .dout(n3824));
  jor  g03569(.dina(n2005), .dinb(n970), .dout(n3825));
  jor  g03570(.dina(n880), .dinb(n1759), .dout(n3826));
  jor  g03571(.dina(n967), .dinb(n1881), .dout(n3827));
  jor  g03572(.dina(n972), .dinb(n2007), .dout(n3828));
  jand g03573(.dina(n3828), .dinb(n3827), .dout(n3829));
  jand g03574(.dina(n3829), .dinb(n3826), .dout(n3830));
  jand g03575(.dina(n3830), .dinb(n3825), .dout(n3831));
  jxor g03576(.dina(n3831), .dinb(n810), .dout(n3832));
  jxor g03577(.dina(n3832), .dinb(n3824), .dout(n3833));
  jxor g03578(.dina(n3833), .dinb(n3726), .dout(n3834));
  jor  g03579(.dina(n2413), .dinb(n728), .dout(n3835));
  jor  g03580(.dina(n660), .dinb(n2142), .dout(n3836));
  jor  g03581(.dina(n731), .dinb(n2279), .dout(n3837));
  jor  g03582(.dina(n726), .dinb(n2415), .dout(n3838));
  jand g03583(.dina(n3838), .dinb(n3837), .dout(n3839));
  jand g03584(.dina(n3839), .dinb(n3836), .dout(n3840));
  jand g03585(.dina(n3840), .dinb(n3835), .dout(n3841));
  jxor g03586(.dina(n3841), .dinb(n606), .dout(n3842));
  jxor g03587(.dina(n3842), .dinb(n3834), .dout(n3843));
  jnot g03588(.din(n3843), .dout(n3844));
  jxor g03589(.dina(n3844), .dinb(n3723), .dout(n3845));
  jor  g03590(.dina(n2860), .dinb(n544), .dout(n3846));
  jor  g03591(.dina(n486), .dinb(n2563), .dout(n3847));
  jor  g03592(.dina(n547), .dinb(n2713), .dout(n3848));
  jor  g03593(.dina(n542), .dinb(n2862), .dout(n3849));
  jand g03594(.dina(n3849), .dinb(n3848), .dout(n3850));
  jand g03595(.dina(n3850), .dinb(n3847), .dout(n3851));
  jand g03596(.dina(n3851), .dinb(n3846), .dout(n3852));
  jxor g03597(.dina(n3852), .dinb(n446), .dout(n3853));
  jxor g03598(.dina(n3853), .dinb(n3845), .dout(n3854));
  jxor g03599(.dina(n3854), .dinb(n3719), .dout(n3855));
  jor  g03600(.dina(n3346), .dinb(n397), .dout(n3856));
  jor  g03601(.dina(n354), .dinb(n3023), .dout(n3857));
  jor  g03602(.dina(n399), .dinb(n3348), .dout(n3858));
  jor  g03603(.dina(n394), .dinb(n3186), .dout(n3859));
  jand g03604(.dina(n3859), .dinb(n3858), .dout(n3860));
  jand g03605(.dina(n3860), .dinb(n3857), .dout(n3861));
  jand g03606(.dina(n3861), .dinb(n3856), .dout(n3862));
  jxor g03607(.dina(n3862), .dinb(n364), .dout(n3863));
  jxor g03608(.dina(n3863), .dinb(n3855), .dout(n3864));
  jxor g03609(.dina(n3864), .dinb(n3716), .dout(n3865));
  jand g03610(.dina(b35 ), .dinb(b34 ), .dout(n3866));
  jand g03611(.dina(n3694), .dinb(n3693), .dout(n3867));
  jor  g03612(.dina(n3867), .dinb(n3866), .dout(n3868));
  jxor g03613(.dina(b36 ), .dinb(b35 ), .dout(n3869));
  jnot g03614(.din(n3869), .dout(n3870));
  jxor g03615(.dina(n3870), .dinb(n3868), .dout(n3871));
  jor  g03616(.dina(n3871), .dinb(n296), .dout(n3872));
  jnot g03617(.din(b36 ), .dout(n3873));
  jor  g03618(.dina(n264), .dinb(n3873), .dout(n3874));
  jor  g03619(.dina(n280), .dinb(n3522), .dout(n3875));
  jor  g03620(.dina(n294), .dinb(n3698), .dout(n3876));
  jand g03621(.dina(n3876), .dinb(n3875), .dout(n3877));
  jand g03622(.dina(n3877), .dinb(n3874), .dout(n3878));
  jand g03623(.dina(n3878), .dinb(n3872), .dout(n3879));
  jxor g03624(.dina(n3879), .dinb(n278), .dout(n3880));
  jxor g03625(.dina(n3880), .dinb(n3865), .dout(n3881));
  jxor g03626(.dina(n3881), .dinb(n3711), .dout(f36 ));
  jnot g03627(.din(n3880), .dout(n3883));
  jor  g03628(.dina(n3883), .dinb(n3865), .dout(n3884));
  jor  g03629(.dina(n3881), .dinb(n3711), .dout(n3885));
  jand g03630(.dina(n3885), .dinb(n3884), .dout(n3886));
  jand g03631(.dina(n3863), .dinb(n3855), .dout(n3887));
  jnot g03632(.din(n3887), .dout(n3888));
  jnot g03633(.din(n3864), .dout(n3889));
  jor  g03634(.dina(n3889), .dinb(n3716), .dout(n3890));
  jand g03635(.dina(n3890), .dinb(n3888), .dout(n3891));
  jand g03636(.dina(n3853), .dinb(n3845), .dout(n3892));
  jand g03637(.dina(n3854), .dinb(n3719), .dout(n3893));
  jor  g03638(.dina(n3893), .dinb(n3892), .dout(n3894));
  jand g03639(.dina(n3842), .dinb(n3834), .dout(n3895));
  jnot g03640(.din(n3895), .dout(n3896));
  jor  g03641(.dina(n3844), .dinb(n3723), .dout(n3897));
  jand g03642(.dina(n3897), .dinb(n3896), .dout(n3898));
  jand g03643(.dina(n3832), .dinb(n3824), .dout(n3899));
  jand g03644(.dina(n3833), .dinb(n3726), .dout(n3900));
  jor  g03645(.dina(n3900), .dinb(n3899), .dout(n3901));
  jand g03646(.dina(n3822), .dinb(n3814), .dout(n3902));
  jand g03647(.dina(n3823), .dinb(n3729), .dout(n3903));
  jor  g03648(.dina(n3903), .dinb(n3902), .dout(n3904));
  jand g03649(.dina(n3812), .dinb(n3804), .dout(n3905));
  jand g03650(.dina(n3813), .dinb(n3732), .dout(n3906));
  jor  g03651(.dina(n3906), .dinb(n3905), .dout(n3907));
  jand g03652(.dina(n3802), .dinb(n3794), .dout(n3908));
  jand g03653(.dina(n3803), .dinb(n3735), .dout(n3909));
  jor  g03654(.dina(n3909), .dinb(n3908), .dout(n3910));
  jand g03655(.dina(n3789), .dinb(n3781), .dout(n3911));
  jand g03656(.dina(n3793), .dinb(n3790), .dout(n3912));
  jor  g03657(.dina(n3912), .dinb(n3911), .dout(n3913));
  jand g03658(.dina(n3779), .dinb(n3771), .dout(n3914));
  jand g03659(.dina(n3780), .dinb(n3738), .dout(n3915));
  jor  g03660(.dina(n3915), .dinb(n3914), .dout(n3916));
  jor  g03661(.dina(n3769), .dinb(n3761), .dout(n3917));
  jand g03662(.dina(n3770), .dinb(n3743), .dout(n3918));
  jnot g03663(.din(n3918), .dout(n3919));
  jand g03664(.dina(n3919), .dinb(n3917), .dout(n3920));
  jnot g03665(.din(n3920), .dout(n3921));
  jnot g03666(.din(n3744), .dout(n3922));
  jand g03667(.dina(n3746), .dinb(n3922), .dout(n3923));
  jand g03668(.dina(n3759), .dinb(n3748), .dout(n3924));
  jor  g03669(.dina(n3924), .dinb(n3923), .dout(n3925));
  jxor g03670(.dina(a38 ), .dinb(a37 ), .dout(n3926));
  jnot g03671(.din(n3926), .dout(n3927));
  jand g03672(.dina(n3927), .dinb(n3745), .dout(n3928));
  jand g03673(.dina(n3928), .dinb(b1 ), .dout(n3929));
  jand g03674(.dina(n3926), .dinb(n3745), .dout(n3930));
  jand g03675(.dina(n3930), .dinb(n259), .dout(n3931));
  jnot g03676(.din(n3745), .dout(n3932));
  jxor g03677(.dina(a37 ), .dinb(a36 ), .dout(n3933));
  jand g03678(.dina(n3933), .dinb(n3932), .dout(n3934));
  jand g03679(.dina(n3934), .dinb(b0 ), .dout(n3935));
  jor  g03680(.dina(n3935), .dinb(n3931), .dout(n3936));
  jor  g03681(.dina(n3936), .dinb(n3929), .dout(n3937));
  jnot g03682(.din(a38 ), .dout(n3938));
  jor  g03683(.dina(n3747), .dinb(n3938), .dout(n3939));
  jxor g03684(.dina(n3939), .dinb(n3937), .dout(n3940));
  jor  g03685(.dina(n3751), .dinb(n337), .dout(n3941));
  jor  g03686(.dina(n3754), .dinb(n303), .dout(n3942));
  jor  g03687(.dina(n3574), .dinb(n293), .dout(n3943));
  jand g03688(.dina(n3943), .dinb(n3942), .dout(n3944));
  jor  g03689(.dina(n3749), .dinb(n340), .dout(n3945));
  jand g03690(.dina(n3945), .dinb(n3944), .dout(n3946));
  jand g03691(.dina(n3946), .dinb(n3941), .dout(n3947));
  jxor g03692(.dina(n3947), .dinb(a35 ), .dout(n3948));
  jxor g03693(.dina(n3948), .dinb(n3940), .dout(n3949));
  jxor g03694(.dina(n3949), .dinb(n3925), .dout(n3950));
  jnot g03695(.din(n3950), .dout(n3951));
  jor  g03696(.dina(n3239), .dinb(n466), .dout(n3952));
  jor  g03697(.dina(n3242), .dinb(n415), .dout(n3953));
  jor  g03698(.dina(n3072), .dinb(n377), .dout(n3954));
  jand g03699(.dina(n3954), .dinb(n3953), .dout(n3955));
  jor  g03700(.dina(n3237), .dinb(n469), .dout(n3956));
  jand g03701(.dina(n3956), .dinb(n3955), .dout(n3957));
  jand g03702(.dina(n3957), .dinb(n3952), .dout(n3958));
  jxor g03703(.dina(n3958), .dinb(a32 ), .dout(n3959));
  jxor g03704(.dina(n3959), .dinb(n3951), .dout(n3960));
  jxor g03705(.dina(n3960), .dinb(n3921), .dout(n3961));
  jor  g03706(.dina(n2764), .dinb(n635), .dout(n3962));
  jor  g03707(.dina(n2609), .dinb(n519), .dout(n3963));
  jor  g03708(.dina(n2761), .dinb(n637), .dout(n3964));
  jor  g03709(.dina(n2766), .dinb(n572), .dout(n3965));
  jand g03710(.dina(n3965), .dinb(n3964), .dout(n3966));
  jand g03711(.dina(n3966), .dinb(n3963), .dout(n3967));
  jand g03712(.dina(n3967), .dinb(n3962), .dout(n3968));
  jxor g03713(.dina(n3968), .dinb(n2468), .dout(n3969));
  jxor g03714(.dina(n3969), .dinb(n3961), .dout(n3970));
  jxor g03715(.dina(n3970), .dinb(n3916), .dout(n3971));
  jor  g03716(.dina(n2324), .dinb(n850), .dout(n3972));
  jor  g03717(.dina(n2186), .dinb(n704), .dout(n3973));
  jor  g03718(.dina(n2321), .dinb(n772), .dout(n3974));
  jor  g03719(.dina(n2326), .dinb(n852), .dout(n3975));
  jand g03720(.dina(n3975), .dinb(n3974), .dout(n3976));
  jand g03721(.dina(n3976), .dinb(n3973), .dout(n3977));
  jand g03722(.dina(n3977), .dinb(n3972), .dout(n3978));
  jxor g03723(.dina(n3978), .dinb(n2057), .dout(n3979));
  jxor g03724(.dina(n3979), .dinb(n3971), .dout(n3980));
  jxor g03725(.dina(n3980), .dinb(n3913), .dout(n3981));
  jor  g03726(.dina(n1921), .dinb(n1112), .dout(n3982));
  jor  g03727(.dina(n1806), .dinb(n934), .dout(n3983));
  jor  g03728(.dina(n1918), .dinb(n1018), .dout(n3984));
  jor  g03729(.dina(n1923), .dinb(n1114), .dout(n3985));
  jand g03730(.dina(n3985), .dinb(n3984), .dout(n3986));
  jand g03731(.dina(n3986), .dinb(n3983), .dout(n3987));
  jand g03732(.dina(n3987), .dinb(n3982), .dout(n3988));
  jxor g03733(.dina(n3988), .dinb(n1687), .dout(n3989));
  jxor g03734(.dina(n3989), .dinb(n3981), .dout(n3990));
  jxor g03735(.dina(n3990), .dinb(n3910), .dout(n3991));
  jor  g03736(.dina(n1414), .dinb(n1569), .dout(n3992));
  jor  g03737(.dina(n1453), .dinb(n1211), .dout(n3993));
  jor  g03738(.dina(n1566), .dinb(n1307), .dout(n3994));
  jor  g03739(.dina(n1571), .dinb(n1416), .dout(n3995));
  jand g03740(.dina(n3995), .dinb(n3994), .dout(n3996));
  jand g03741(.dina(n3996), .dinb(n3993), .dout(n3997));
  jand g03742(.dina(n3997), .dinb(n3992), .dout(n3998));
  jxor g03743(.dina(n3998), .dinb(n1351), .dout(n3999));
  jxor g03744(.dina(n3999), .dinb(n3991), .dout(n4000));
  jxor g03745(.dina(n4000), .dinb(n3907), .dout(n4001));
  jor  g03746(.dina(n1757), .dinb(n1248), .dout(n4002));
  jor  g03747(.dina(n1147), .dinb(n1527), .dout(n4003));
  jor  g03748(.dina(n1251), .dinb(n1637), .dout(n4004));
  jor  g03749(.dina(n1246), .dinb(n1759), .dout(n4005));
  jand g03750(.dina(n4005), .dinb(n4004), .dout(n4006));
  jand g03751(.dina(n4006), .dinb(n4003), .dout(n4007));
  jand g03752(.dina(n4007), .dinb(n4002), .dout(n4008));
  jxor g03753(.dina(n4008), .dinb(n1061), .dout(n4009));
  jxor g03754(.dina(n4009), .dinb(n4001), .dout(n4010));
  jxor g03755(.dina(n4010), .dinb(n3904), .dout(n4011));
  jor  g03756(.dina(n2140), .dinb(n970), .dout(n4012));
  jor  g03757(.dina(n880), .dinb(n1881), .dout(n4013));
  jor  g03758(.dina(n967), .dinb(n2007), .dout(n4014));
  jor  g03759(.dina(n972), .dinb(n2142), .dout(n4015));
  jand g03760(.dina(n4015), .dinb(n4014), .dout(n4016));
  jand g03761(.dina(n4016), .dinb(n4013), .dout(n4017));
  jand g03762(.dina(n4017), .dinb(n4012), .dout(n4018));
  jxor g03763(.dina(n4018), .dinb(n810), .dout(n4019));
  jxor g03764(.dina(n4019), .dinb(n4011), .dout(n4020));
  jxor g03765(.dina(n4020), .dinb(n3901), .dout(n4021));
  jor  g03766(.dina(n2561), .dinb(n728), .dout(n4022));
  jor  g03767(.dina(n660), .dinb(n2279), .dout(n4023));
  jor  g03768(.dina(n726), .dinb(n2563), .dout(n4024));
  jor  g03769(.dina(n731), .dinb(n2415), .dout(n4025));
  jand g03770(.dina(n4025), .dinb(n4024), .dout(n4026));
  jand g03771(.dina(n4026), .dinb(n4023), .dout(n4027));
  jand g03772(.dina(n4027), .dinb(n4022), .dout(n4028));
  jxor g03773(.dina(n4028), .dinb(n606), .dout(n4029));
  jxor g03774(.dina(n4029), .dinb(n4021), .dout(n4030));
  jnot g03775(.din(n4030), .dout(n4031));
  jxor g03776(.dina(n4031), .dinb(n3898), .dout(n4032));
  jor  g03777(.dina(n3021), .dinb(n544), .dout(n4033));
  jor  g03778(.dina(n486), .dinb(n2713), .dout(n4034));
  jor  g03779(.dina(n547), .dinb(n2862), .dout(n4035));
  jor  g03780(.dina(n542), .dinb(n3023), .dout(n4036));
  jand g03781(.dina(n4036), .dinb(n4035), .dout(n4037));
  jand g03782(.dina(n4037), .dinb(n4034), .dout(n4038));
  jand g03783(.dina(n4038), .dinb(n4033), .dout(n4039));
  jxor g03784(.dina(n4039), .dinb(n446), .dout(n4040));
  jxor g03785(.dina(n4040), .dinb(n4032), .dout(n4041));
  jxor g03786(.dina(n4041), .dinb(n3894), .dout(n4042));
  jor  g03787(.dina(n3520), .dinb(n397), .dout(n4043));
  jor  g03788(.dina(n354), .dinb(n3186), .dout(n4044));
  jor  g03789(.dina(n399), .dinb(n3522), .dout(n4045));
  jor  g03790(.dina(n394), .dinb(n3348), .dout(n4046));
  jand g03791(.dina(n4046), .dinb(n4045), .dout(n4047));
  jand g03792(.dina(n4047), .dinb(n4044), .dout(n4048));
  jand g03793(.dina(n4048), .dinb(n4043), .dout(n4049));
  jxor g03794(.dina(n4049), .dinb(n364), .dout(n4050));
  jxor g03795(.dina(n4050), .dinb(n4042), .dout(n4051));
  jxor g03796(.dina(n4051), .dinb(n3891), .dout(n4052));
  jand g03797(.dina(b36 ), .dinb(b35 ), .dout(n4053));
  jand g03798(.dina(n3869), .dinb(n3868), .dout(n4054));
  jor  g03799(.dina(n4054), .dinb(n4053), .dout(n4055));
  jxor g03800(.dina(b37 ), .dinb(b36 ), .dout(n4056));
  jnot g03801(.din(n4056), .dout(n4057));
  jxor g03802(.dina(n4057), .dinb(n4055), .dout(n4058));
  jor  g03803(.dina(n4058), .dinb(n296), .dout(n4059));
  jnot g03804(.din(b37 ), .dout(n4060));
  jor  g03805(.dina(n264), .dinb(n4060), .dout(n4061));
  jor  g03806(.dina(n280), .dinb(n3698), .dout(n4062));
  jor  g03807(.dina(n294), .dinb(n3873), .dout(n4063));
  jand g03808(.dina(n4063), .dinb(n4062), .dout(n4064));
  jand g03809(.dina(n4064), .dinb(n4061), .dout(n4065));
  jand g03810(.dina(n4065), .dinb(n4059), .dout(n4066));
  jxor g03811(.dina(n4066), .dinb(n278), .dout(n4067));
  jxor g03812(.dina(n4067), .dinb(n4052), .dout(n4068));
  jxor g03813(.dina(n4068), .dinb(n3886), .dout(f37 ));
  jnot g03814(.din(n4067), .dout(n4070));
  jor  g03815(.dina(n4070), .dinb(n4052), .dout(n4071));
  jor  g03816(.dina(n4068), .dinb(n3886), .dout(n4072));
  jand g03817(.dina(n4072), .dinb(n4071), .dout(n4073));
  jand g03818(.dina(n4050), .dinb(n4042), .dout(n4074));
  jnot g03819(.din(n4074), .dout(n4075));
  jnot g03820(.din(n4051), .dout(n4076));
  jor  g03821(.dina(n4076), .dinb(n3891), .dout(n4077));
  jand g03822(.dina(n4077), .dinb(n4075), .dout(n4078));
  jand g03823(.dina(n4040), .dinb(n4032), .dout(n4079));
  jand g03824(.dina(n4041), .dinb(n3894), .dout(n4080));
  jor  g03825(.dina(n4080), .dinb(n4079), .dout(n4081));
  jand g03826(.dina(n4029), .dinb(n4021), .dout(n4082));
  jnot g03827(.din(n4082), .dout(n4083));
  jor  g03828(.dina(n4031), .dinb(n3898), .dout(n4084));
  jand g03829(.dina(n4084), .dinb(n4083), .dout(n4085));
  jand g03830(.dina(n4019), .dinb(n4011), .dout(n4086));
  jand g03831(.dina(n4020), .dinb(n3901), .dout(n4087));
  jor  g03832(.dina(n4087), .dinb(n4086), .dout(n4088));
  jand g03833(.dina(n4009), .dinb(n4001), .dout(n4089));
  jand g03834(.dina(n4010), .dinb(n3904), .dout(n4090));
  jor  g03835(.dina(n4090), .dinb(n4089), .dout(n4091));
  jand g03836(.dina(n3999), .dinb(n3991), .dout(n4092));
  jand g03837(.dina(n4000), .dinb(n3907), .dout(n4093));
  jor  g03838(.dina(n4093), .dinb(n4092), .dout(n4094));
  jand g03839(.dina(n3989), .dinb(n3981), .dout(n4095));
  jand g03840(.dina(n3990), .dinb(n3910), .dout(n4096));
  jor  g03841(.dina(n4096), .dinb(n4095), .dout(n4097));
  jand g03842(.dina(n3979), .dinb(n3971), .dout(n4098));
  jand g03843(.dina(n3980), .dinb(n3913), .dout(n4099));
  jor  g03844(.dina(n4099), .dinb(n4098), .dout(n4100));
  jand g03845(.dina(n3969), .dinb(n3961), .dout(n4101));
  jand g03846(.dina(n3970), .dinb(n3916), .dout(n4102));
  jor  g03847(.dina(n4102), .dinb(n4101), .dout(n4103));
  jor  g03848(.dina(n3959), .dinb(n3951), .dout(n4104));
  jand g03849(.dina(n3960), .dinb(n3921), .dout(n4105));
  jnot g03850(.din(n4105), .dout(n4106));
  jand g03851(.dina(n4106), .dinb(n4104), .dout(n4107));
  jnot g03852(.din(n4107), .dout(n4108));
  jor  g03853(.dina(n3948), .dinb(n3940), .dout(n4109));
  jand g03854(.dina(n3949), .dinb(n3925), .dout(n4110));
  jnot g03855(.din(n4110), .dout(n4111));
  jand g03856(.dina(n4111), .dinb(n4109), .dout(n4112));
  jnot g03857(.din(n4112), .dout(n4113));
  jand g03858(.dina(n3934), .dinb(b1 ), .dout(n4114));
  jor  g03859(.dina(n3933), .dinb(n3745), .dout(n4115));
  jor  g03860(.dina(n4115), .dinb(n3927), .dout(n4116));
  jnot g03861(.din(n4116), .dout(n4117));
  jand g03862(.dina(n4117), .dinb(b0 ), .dout(n4118));
  jand g03863(.dina(n3930), .dinb(n273), .dout(n4119));
  jand g03864(.dina(n3928), .dinb(b2 ), .dout(n4120));
  jor  g03865(.dina(n4120), .dinb(n4119), .dout(n4121));
  jor  g03866(.dina(n4121), .dinb(n4118), .dout(n4122));
  jor  g03867(.dina(n4122), .dinb(n4114), .dout(n4123));
  jnot g03868(.din(n3937), .dout(n4124));
  jand g03869(.dina(n3747), .dinb(a38 ), .dout(n4125));
  jand g03870(.dina(n4125), .dinb(n4124), .dout(n4126));
  jnot g03871(.din(n4126), .dout(n4127));
  jand g03872(.dina(n4127), .dinb(a38 ), .dout(n4128));
  jxor g03873(.dina(n4128), .dinb(n4123), .dout(n4129));
  jnot g03874(.din(n4129), .dout(n4130));
  jor  g03875(.dina(n3751), .dinb(n374), .dout(n4131));
  jor  g03876(.dina(n3754), .dinb(n340), .dout(n4132));
  jor  g03877(.dina(n3574), .dinb(n303), .dout(n4133));
  jand g03878(.dina(n4133), .dinb(n4132), .dout(n4134));
  jor  g03879(.dina(n3749), .dinb(n377), .dout(n4135));
  jand g03880(.dina(n4135), .dinb(n4134), .dout(n4136));
  jand g03881(.dina(n4136), .dinb(n4131), .dout(n4137));
  jxor g03882(.dina(n4137), .dinb(a35 ), .dout(n4138));
  jxor g03883(.dina(n4138), .dinb(n4130), .dout(n4139));
  jxor g03884(.dina(n4139), .dinb(n4113), .dout(n4140));
  jor  g03885(.dina(n3239), .dinb(n517), .dout(n4141));
  jor  g03886(.dina(n3237), .dinb(n519), .dout(n4142));
  jor  g03887(.dina(n3242), .dinb(n469), .dout(n4143));
  jor  g03888(.dina(n3072), .dinb(n415), .dout(n4144));
  jand g03889(.dina(n4144), .dinb(n4143), .dout(n4145));
  jand g03890(.dina(n4145), .dinb(n4142), .dout(n4146));
  jand g03891(.dina(n4146), .dinb(n4141), .dout(n4147));
  jxor g03892(.dina(n4147), .dinb(n2918), .dout(n4148));
  jxor g03893(.dina(n4148), .dinb(n4140), .dout(n4149));
  jxor g03894(.dina(n4149), .dinb(n4108), .dout(n4150));
  jor  g03895(.dina(n2764), .dinb(n702), .dout(n4151));
  jor  g03896(.dina(n2609), .dinb(n572), .dout(n4152));
  jor  g03897(.dina(n2761), .dinb(n704), .dout(n4153));
  jor  g03898(.dina(n2766), .dinb(n637), .dout(n4154));
  jand g03899(.dina(n4154), .dinb(n4153), .dout(n4155));
  jand g03900(.dina(n4155), .dinb(n4152), .dout(n4156));
  jand g03901(.dina(n4156), .dinb(n4151), .dout(n4157));
  jxor g03902(.dina(n4157), .dinb(n2468), .dout(n4158));
  jxor g03903(.dina(n4158), .dinb(n4150), .dout(n4159));
  jxor g03904(.dina(n4159), .dinb(n4103), .dout(n4160));
  jor  g03905(.dina(n2324), .dinb(n932), .dout(n4161));
  jor  g03906(.dina(n2186), .dinb(n772), .dout(n4162));
  jor  g03907(.dina(n2321), .dinb(n852), .dout(n4163));
  jor  g03908(.dina(n2326), .dinb(n934), .dout(n4164));
  jand g03909(.dina(n4164), .dinb(n4163), .dout(n4165));
  jand g03910(.dina(n4165), .dinb(n4162), .dout(n4166));
  jand g03911(.dina(n4166), .dinb(n4161), .dout(n4167));
  jxor g03912(.dina(n4167), .dinb(n2057), .dout(n4168));
  jxor g03913(.dina(n4168), .dinb(n4160), .dout(n4169));
  jxor g03914(.dina(n4169), .dinb(n4100), .dout(n4170));
  jor  g03915(.dina(n1921), .dinb(n1209), .dout(n4171));
  jor  g03916(.dina(n1806), .dinb(n1018), .dout(n4172));
  jor  g03917(.dina(n1923), .dinb(n1211), .dout(n4173));
  jor  g03918(.dina(n1918), .dinb(n1114), .dout(n4174));
  jand g03919(.dina(n4174), .dinb(n4173), .dout(n4175));
  jand g03920(.dina(n4175), .dinb(n4172), .dout(n4176));
  jand g03921(.dina(n4176), .dinb(n4171), .dout(n4177));
  jxor g03922(.dina(n4177), .dinb(n1687), .dout(n4178));
  jxor g03923(.dina(n4178), .dinb(n4170), .dout(n4179));
  jxor g03924(.dina(n4179), .dinb(n4097), .dout(n4180));
  jor  g03925(.dina(n1525), .dinb(n1569), .dout(n4181));
  jor  g03926(.dina(n1453), .dinb(n1307), .dout(n4182));
  jor  g03927(.dina(n1571), .dinb(n1527), .dout(n4183));
  jor  g03928(.dina(n1566), .dinb(n1416), .dout(n4184));
  jand g03929(.dina(n4184), .dinb(n4183), .dout(n4185));
  jand g03930(.dina(n4185), .dinb(n4182), .dout(n4186));
  jand g03931(.dina(n4186), .dinb(n4181), .dout(n4187));
  jxor g03932(.dina(n4187), .dinb(n1351), .dout(n4188));
  jxor g03933(.dina(n4188), .dinb(n4180), .dout(n4189));
  jxor g03934(.dina(n4189), .dinb(n4094), .dout(n4190));
  jor  g03935(.dina(n1879), .dinb(n1248), .dout(n4191));
  jor  g03936(.dina(n1147), .dinb(n1637), .dout(n4192));
  jor  g03937(.dina(n1246), .dinb(n1881), .dout(n4193));
  jor  g03938(.dina(n1251), .dinb(n1759), .dout(n4194));
  jand g03939(.dina(n4194), .dinb(n4193), .dout(n4195));
  jand g03940(.dina(n4195), .dinb(n4192), .dout(n4196));
  jand g03941(.dina(n4196), .dinb(n4191), .dout(n4197));
  jxor g03942(.dina(n4197), .dinb(n1061), .dout(n4198));
  jxor g03943(.dina(n4198), .dinb(n4190), .dout(n4199));
  jxor g03944(.dina(n4199), .dinb(n4091), .dout(n4200));
  jor  g03945(.dina(n2277), .dinb(n970), .dout(n4201));
  jor  g03946(.dina(n880), .dinb(n2007), .dout(n4202));
  jor  g03947(.dina(n967), .dinb(n2142), .dout(n4203));
  jor  g03948(.dina(n972), .dinb(n2279), .dout(n4204));
  jand g03949(.dina(n4204), .dinb(n4203), .dout(n4205));
  jand g03950(.dina(n4205), .dinb(n4202), .dout(n4206));
  jand g03951(.dina(n4206), .dinb(n4201), .dout(n4207));
  jxor g03952(.dina(n4207), .dinb(n810), .dout(n4208));
  jxor g03953(.dina(n4208), .dinb(n4200), .dout(n4209));
  jxor g03954(.dina(n4209), .dinb(n4088), .dout(n4210));
  jor  g03955(.dina(n2711), .dinb(n728), .dout(n4211));
  jor  g03956(.dina(n660), .dinb(n2415), .dout(n4212));
  jor  g03957(.dina(n731), .dinb(n2563), .dout(n4213));
  jor  g03958(.dina(n726), .dinb(n2713), .dout(n4214));
  jand g03959(.dina(n4214), .dinb(n4213), .dout(n4215));
  jand g03960(.dina(n4215), .dinb(n4212), .dout(n4216));
  jand g03961(.dina(n4216), .dinb(n4211), .dout(n4217));
  jxor g03962(.dina(n4217), .dinb(n606), .dout(n4218));
  jxor g03963(.dina(n4218), .dinb(n4210), .dout(n4219));
  jnot g03964(.din(n4219), .dout(n4220));
  jxor g03965(.dina(n4220), .dinb(n4085), .dout(n4221));
  jor  g03966(.dina(n3184), .dinb(n544), .dout(n4222));
  jor  g03967(.dina(n486), .dinb(n2862), .dout(n4223));
  jor  g03968(.dina(n547), .dinb(n3023), .dout(n4224));
  jor  g03969(.dina(n542), .dinb(n3186), .dout(n4225));
  jand g03970(.dina(n4225), .dinb(n4224), .dout(n4226));
  jand g03971(.dina(n4226), .dinb(n4223), .dout(n4227));
  jand g03972(.dina(n4227), .dinb(n4222), .dout(n4228));
  jxor g03973(.dina(n4228), .dinb(n446), .dout(n4229));
  jxor g03974(.dina(n4229), .dinb(n4221), .dout(n4230));
  jxor g03975(.dina(n4230), .dinb(n4081), .dout(n4231));
  jor  g03976(.dina(n3696), .dinb(n397), .dout(n4232));
  jor  g03977(.dina(n354), .dinb(n3348), .dout(n4233));
  jor  g03978(.dina(n399), .dinb(n3698), .dout(n4234));
  jor  g03979(.dina(n394), .dinb(n3522), .dout(n4235));
  jand g03980(.dina(n4235), .dinb(n4234), .dout(n4236));
  jand g03981(.dina(n4236), .dinb(n4233), .dout(n4237));
  jand g03982(.dina(n4237), .dinb(n4232), .dout(n4238));
  jxor g03983(.dina(n4238), .dinb(n364), .dout(n4239));
  jxor g03984(.dina(n4239), .dinb(n4231), .dout(n4240));
  jxor g03985(.dina(n4240), .dinb(n4078), .dout(n4241));
  jand g03986(.dina(b37 ), .dinb(b36 ), .dout(n4242));
  jand g03987(.dina(n4056), .dinb(n4055), .dout(n4243));
  jor  g03988(.dina(n4243), .dinb(n4242), .dout(n4244));
  jxor g03989(.dina(b38 ), .dinb(b37 ), .dout(n4245));
  jnot g03990(.din(n4245), .dout(n4246));
  jxor g03991(.dina(n4246), .dinb(n4244), .dout(n4247));
  jor  g03992(.dina(n4247), .dinb(n296), .dout(n4248));
  jnot g03993(.din(b38 ), .dout(n4249));
  jor  g03994(.dina(n264), .dinb(n4249), .dout(n4250));
  jor  g03995(.dina(n294), .dinb(n4060), .dout(n4251));
  jor  g03996(.dina(n280), .dinb(n3873), .dout(n4252));
  jand g03997(.dina(n4252), .dinb(n4251), .dout(n4253));
  jand g03998(.dina(n4253), .dinb(n4250), .dout(n4254));
  jand g03999(.dina(n4254), .dinb(n4248), .dout(n4255));
  jxor g04000(.dina(n4255), .dinb(n278), .dout(n4256));
  jxor g04001(.dina(n4256), .dinb(n4241), .dout(n4257));
  jxor g04002(.dina(n4257), .dinb(n4073), .dout(f38 ));
  jnot g04003(.din(n4256), .dout(n4259));
  jor  g04004(.dina(n4259), .dinb(n4241), .dout(n4260));
  jor  g04005(.dina(n4257), .dinb(n4073), .dout(n4261));
  jand g04006(.dina(n4261), .dinb(n4260), .dout(n4262));
  jand g04007(.dina(n4239), .dinb(n4231), .dout(n4263));
  jnot g04008(.din(n4263), .dout(n4264));
  jnot g04009(.din(n4240), .dout(n4265));
  jor  g04010(.dina(n4265), .dinb(n4078), .dout(n4266));
  jand g04011(.dina(n4266), .dinb(n4264), .dout(n4267));
  jand g04012(.dina(n4229), .dinb(n4221), .dout(n4268));
  jand g04013(.dina(n4230), .dinb(n4081), .dout(n4269));
  jor  g04014(.dina(n4269), .dinb(n4268), .dout(n4270));
  jand g04015(.dina(n4218), .dinb(n4210), .dout(n4271));
  jnot g04016(.din(n4271), .dout(n4272));
  jor  g04017(.dina(n4220), .dinb(n4085), .dout(n4273));
  jand g04018(.dina(n4273), .dinb(n4272), .dout(n4274));
  jand g04019(.dina(n4208), .dinb(n4200), .dout(n4275));
  jand g04020(.dina(n4209), .dinb(n4088), .dout(n4276));
  jor  g04021(.dina(n4276), .dinb(n4275), .dout(n4277));
  jand g04022(.dina(n4198), .dinb(n4190), .dout(n4278));
  jand g04023(.dina(n4199), .dinb(n4091), .dout(n4279));
  jor  g04024(.dina(n4279), .dinb(n4278), .dout(n4280));
  jand g04025(.dina(n4188), .dinb(n4180), .dout(n4281));
  jand g04026(.dina(n4189), .dinb(n4094), .dout(n4282));
  jor  g04027(.dina(n4282), .dinb(n4281), .dout(n4283));
  jand g04028(.dina(n4178), .dinb(n4170), .dout(n4284));
  jand g04029(.dina(n4179), .dinb(n4097), .dout(n4285));
  jor  g04030(.dina(n4285), .dinb(n4284), .dout(n4286));
  jand g04031(.dina(n4168), .dinb(n4160), .dout(n4287));
  jand g04032(.dina(n4169), .dinb(n4100), .dout(n4288));
  jor  g04033(.dina(n4288), .dinb(n4287), .dout(n4289));
  jand g04034(.dina(n4148), .dinb(n4140), .dout(n4290));
  jand g04035(.dina(n4149), .dinb(n4108), .dout(n4291));
  jor  g04036(.dina(n4291), .dinb(n4290), .dout(n4292));
  jor  g04037(.dina(n4138), .dinb(n4130), .dout(n4293));
  jand g04038(.dina(n4139), .dinb(n4113), .dout(n4294));
  jnot g04039(.din(n4294), .dout(n4295));
  jand g04040(.dina(n4295), .dinb(n4293), .dout(n4296));
  jnot g04041(.din(n4296), .dout(n4297));
  jor  g04042(.dina(n4127), .dinb(n4123), .dout(n4298));
  jxor g04043(.dina(a39 ), .dinb(a38 ), .dout(n4299));
  jand g04044(.dina(n4299), .dinb(b0 ), .dout(n4300));
  jnot g04045(.din(n4300), .dout(n4301));
  jxor g04046(.dina(n4301), .dinb(n4298), .dout(n4302));
  jnot g04047(.din(n3928), .dout(n4303));
  jor  g04048(.dina(n4303), .dinb(n303), .dout(n4304));
  jnot g04049(.din(n3930), .dout(n4305));
  jor  g04050(.dina(n4305), .dinb(n301), .dout(n4306));
  jor  g04051(.dina(n4116), .dinb(n305), .dout(n4307));
  jnot g04052(.din(n3934), .dout(n4308));
  jor  g04053(.dina(n4308), .dinb(n293), .dout(n4309));
  jand g04054(.dina(n4309), .dinb(n4307), .dout(n4310));
  jand g04055(.dina(n4310), .dinb(n4306), .dout(n4311));
  jand g04056(.dina(n4311), .dinb(n4304), .dout(n4312));
  jxor g04057(.dina(n4312), .dinb(n3938), .dout(n4313));
  jxor g04058(.dina(n4313), .dinb(n4302), .dout(n4314));
  jnot g04059(.din(n4314), .dout(n4315));
  jor  g04060(.dina(n3751), .dinb(n412), .dout(n4316));
  jor  g04061(.dina(n3749), .dinb(n415), .dout(n4317));
  jor  g04062(.dina(n3574), .dinb(n340), .dout(n4318));
  jand g04063(.dina(n4318), .dinb(n4317), .dout(n4319));
  jor  g04064(.dina(n3754), .dinb(n377), .dout(n4320));
  jand g04065(.dina(n4320), .dinb(n4319), .dout(n4321));
  jand g04066(.dina(n4321), .dinb(n4316), .dout(n4322));
  jxor g04067(.dina(n4322), .dinb(a35 ), .dout(n4323));
  jxor g04068(.dina(n4323), .dinb(n4315), .dout(n4324));
  jxor g04069(.dina(n4324), .dinb(n4297), .dout(n4325));
  jor  g04070(.dina(n3239), .dinb(n570), .dout(n4326));
  jor  g04071(.dina(n3072), .dinb(n469), .dout(n4327));
  jor  g04072(.dina(n3242), .dinb(n519), .dout(n4328));
  jor  g04073(.dina(n3237), .dinb(n572), .dout(n4329));
  jand g04074(.dina(n4329), .dinb(n4328), .dout(n4330));
  jand g04075(.dina(n4330), .dinb(n4327), .dout(n4331));
  jand g04076(.dina(n4331), .dinb(n4326), .dout(n4332));
  jxor g04077(.dina(n4332), .dinb(n2918), .dout(n4333));
  jxor g04078(.dina(n4333), .dinb(n4325), .dout(n4334));
  jxor g04079(.dina(n4334), .dinb(n4292), .dout(n4335));
  jor  g04080(.dina(n2764), .dinb(n770), .dout(n4336));
  jor  g04081(.dina(n2609), .dinb(n637), .dout(n4337));
  jor  g04082(.dina(n2761), .dinb(n772), .dout(n4338));
  jor  g04083(.dina(n2766), .dinb(n704), .dout(n4339));
  jand g04084(.dina(n4339), .dinb(n4338), .dout(n4340));
  jand g04085(.dina(n4340), .dinb(n4337), .dout(n4341));
  jand g04086(.dina(n4341), .dinb(n4336), .dout(n4342));
  jxor g04087(.dina(n4342), .dinb(n2468), .dout(n4343));
  jxor g04088(.dina(n4343), .dinb(n4335), .dout(n4344));
  jand g04089(.dina(n4158), .dinb(n4150), .dout(n4345));
  jand g04090(.dina(n4159), .dinb(n4103), .dout(n4346));
  jor  g04091(.dina(n4346), .dinb(n4345), .dout(n4347));
  jxor g04092(.dina(n4347), .dinb(n4344), .dout(n4348));
  jor  g04093(.dina(n2324), .dinb(n1016), .dout(n4349));
  jor  g04094(.dina(n2186), .dinb(n852), .dout(n4350));
  jor  g04095(.dina(n2321), .dinb(n934), .dout(n4351));
  jor  g04096(.dina(n2326), .dinb(n1018), .dout(n4352));
  jand g04097(.dina(n4352), .dinb(n4351), .dout(n4353));
  jand g04098(.dina(n4353), .dinb(n4350), .dout(n4354));
  jand g04099(.dina(n4354), .dinb(n4349), .dout(n4355));
  jxor g04100(.dina(n4355), .dinb(n2057), .dout(n4356));
  jxor g04101(.dina(n4356), .dinb(n4348), .dout(n4357));
  jxor g04102(.dina(n4357), .dinb(n4289), .dout(n4358));
  jor  g04103(.dina(n1921), .dinb(n1305), .dout(n4359));
  jor  g04104(.dina(n1806), .dinb(n1114), .dout(n4360));
  jor  g04105(.dina(n1918), .dinb(n1211), .dout(n4361));
  jor  g04106(.dina(n1923), .dinb(n1307), .dout(n4362));
  jand g04107(.dina(n4362), .dinb(n4361), .dout(n4363));
  jand g04108(.dina(n4363), .dinb(n4360), .dout(n4364));
  jand g04109(.dina(n4364), .dinb(n4359), .dout(n4365));
  jxor g04110(.dina(n4365), .dinb(n1687), .dout(n4366));
  jxor g04111(.dina(n4366), .dinb(n4358), .dout(n4367));
  jxor g04112(.dina(n4367), .dinb(n4286), .dout(n4368));
  jor  g04113(.dina(n1635), .dinb(n1569), .dout(n4369));
  jor  g04114(.dina(n1453), .dinb(n1416), .dout(n4370));
  jor  g04115(.dina(n1571), .dinb(n1637), .dout(n4371));
  jor  g04116(.dina(n1566), .dinb(n1527), .dout(n4372));
  jand g04117(.dina(n4372), .dinb(n4371), .dout(n4373));
  jand g04118(.dina(n4373), .dinb(n4370), .dout(n4374));
  jand g04119(.dina(n4374), .dinb(n4369), .dout(n4375));
  jxor g04120(.dina(n4375), .dinb(n1351), .dout(n4376));
  jxor g04121(.dina(n4376), .dinb(n4368), .dout(n4377));
  jxor g04122(.dina(n4377), .dinb(n4283), .dout(n4378));
  jor  g04123(.dina(n2005), .dinb(n1248), .dout(n4379));
  jor  g04124(.dina(n1147), .dinb(n1759), .dout(n4380));
  jor  g04125(.dina(n1251), .dinb(n1881), .dout(n4381));
  jor  g04126(.dina(n1246), .dinb(n2007), .dout(n4382));
  jand g04127(.dina(n4382), .dinb(n4381), .dout(n4383));
  jand g04128(.dina(n4383), .dinb(n4380), .dout(n4384));
  jand g04129(.dina(n4384), .dinb(n4379), .dout(n4385));
  jxor g04130(.dina(n4385), .dinb(n1061), .dout(n4386));
  jxor g04131(.dina(n4386), .dinb(n4378), .dout(n4387));
  jxor g04132(.dina(n4387), .dinb(n4280), .dout(n4388));
  jor  g04133(.dina(n2413), .dinb(n970), .dout(n4389));
  jor  g04134(.dina(n880), .dinb(n2142), .dout(n4390));
  jor  g04135(.dina(n967), .dinb(n2279), .dout(n4391));
  jor  g04136(.dina(n972), .dinb(n2415), .dout(n4392));
  jand g04137(.dina(n4392), .dinb(n4391), .dout(n4393));
  jand g04138(.dina(n4393), .dinb(n4390), .dout(n4394));
  jand g04139(.dina(n4394), .dinb(n4389), .dout(n4395));
  jxor g04140(.dina(n4395), .dinb(n810), .dout(n4396));
  jxor g04141(.dina(n4396), .dinb(n4388), .dout(n4397));
  jxor g04142(.dina(n4397), .dinb(n4277), .dout(n4398));
  jor  g04143(.dina(n2860), .dinb(n728), .dout(n4399));
  jor  g04144(.dina(n660), .dinb(n2563), .dout(n4400));
  jor  g04145(.dina(n726), .dinb(n2862), .dout(n4401));
  jor  g04146(.dina(n731), .dinb(n2713), .dout(n4402));
  jand g04147(.dina(n4402), .dinb(n4401), .dout(n4403));
  jand g04148(.dina(n4403), .dinb(n4400), .dout(n4404));
  jand g04149(.dina(n4404), .dinb(n4399), .dout(n4405));
  jxor g04150(.dina(n4405), .dinb(n606), .dout(n4406));
  jxor g04151(.dina(n4406), .dinb(n4398), .dout(n4407));
  jnot g04152(.din(n4407), .dout(n4408));
  jxor g04153(.dina(n4408), .dinb(n4274), .dout(n4409));
  jor  g04154(.dina(n3346), .dinb(n544), .dout(n4410));
  jor  g04155(.dina(n486), .dinb(n3023), .dout(n4411));
  jor  g04156(.dina(n542), .dinb(n3348), .dout(n4412));
  jor  g04157(.dina(n547), .dinb(n3186), .dout(n4413));
  jand g04158(.dina(n4413), .dinb(n4412), .dout(n4414));
  jand g04159(.dina(n4414), .dinb(n4411), .dout(n4415));
  jand g04160(.dina(n4415), .dinb(n4410), .dout(n4416));
  jxor g04161(.dina(n4416), .dinb(n446), .dout(n4417));
  jxor g04162(.dina(n4417), .dinb(n4409), .dout(n4418));
  jxor g04163(.dina(n4418), .dinb(n4270), .dout(n4419));
  jor  g04164(.dina(n3871), .dinb(n397), .dout(n4420));
  jor  g04165(.dina(n354), .dinb(n3522), .dout(n4421));
  jor  g04166(.dina(n394), .dinb(n3698), .dout(n4422));
  jor  g04167(.dina(n399), .dinb(n3873), .dout(n4423));
  jand g04168(.dina(n4423), .dinb(n4422), .dout(n4424));
  jand g04169(.dina(n4424), .dinb(n4421), .dout(n4425));
  jand g04170(.dina(n4425), .dinb(n4420), .dout(n4426));
  jxor g04171(.dina(n4426), .dinb(n364), .dout(n4427));
  jxor g04172(.dina(n4427), .dinb(n4419), .dout(n4428));
  jxor g04173(.dina(n4428), .dinb(n4267), .dout(n4429));
  jand g04174(.dina(b38 ), .dinb(b37 ), .dout(n4430));
  jand g04175(.dina(n4245), .dinb(n4244), .dout(n4431));
  jor  g04176(.dina(n4431), .dinb(n4430), .dout(n4432));
  jxor g04177(.dina(b39 ), .dinb(b38 ), .dout(n4433));
  jnot g04178(.din(n4433), .dout(n4434));
  jxor g04179(.dina(n4434), .dinb(n4432), .dout(n4435));
  jor  g04180(.dina(n4435), .dinb(n296), .dout(n4436));
  jnot g04181(.din(b39 ), .dout(n4437));
  jor  g04182(.dina(n264), .dinb(n4437), .dout(n4438));
  jor  g04183(.dina(n280), .dinb(n4060), .dout(n4439));
  jor  g04184(.dina(n294), .dinb(n4249), .dout(n4440));
  jand g04185(.dina(n4440), .dinb(n4439), .dout(n4441));
  jand g04186(.dina(n4441), .dinb(n4438), .dout(n4442));
  jand g04187(.dina(n4442), .dinb(n4436), .dout(n4443));
  jxor g04188(.dina(n4443), .dinb(n278), .dout(n4444));
  jxor g04189(.dina(n4444), .dinb(n4429), .dout(n4445));
  jxor g04190(.dina(n4445), .dinb(n4262), .dout(f39 ));
  jnot g04191(.din(n4444), .dout(n4447));
  jor  g04192(.dina(n4447), .dinb(n4429), .dout(n4448));
  jor  g04193(.dina(n4445), .dinb(n4262), .dout(n4449));
  jand g04194(.dina(n4449), .dinb(n4448), .dout(n4450));
  jand g04195(.dina(n4427), .dinb(n4419), .dout(n4451));
  jnot g04196(.din(n4451), .dout(n4452));
  jnot g04197(.din(n4428), .dout(n4453));
  jor  g04198(.dina(n4453), .dinb(n4267), .dout(n4454));
  jand g04199(.dina(n4454), .dinb(n4452), .dout(n4455));
  jand g04200(.dina(n4417), .dinb(n4409), .dout(n4456));
  jand g04201(.dina(n4418), .dinb(n4270), .dout(n4457));
  jor  g04202(.dina(n4457), .dinb(n4456), .dout(n4458));
  jand g04203(.dina(n4406), .dinb(n4398), .dout(n4459));
  jnot g04204(.din(n4459), .dout(n4460));
  jor  g04205(.dina(n4408), .dinb(n4274), .dout(n4461));
  jand g04206(.dina(n4461), .dinb(n4460), .dout(n4462));
  jand g04207(.dina(n4396), .dinb(n4388), .dout(n4463));
  jand g04208(.dina(n4397), .dinb(n4277), .dout(n4464));
  jor  g04209(.dina(n4464), .dinb(n4463), .dout(n4465));
  jand g04210(.dina(n4386), .dinb(n4378), .dout(n4466));
  jand g04211(.dina(n4387), .dinb(n4280), .dout(n4467));
  jor  g04212(.dina(n4467), .dinb(n4466), .dout(n4468));
  jand g04213(.dina(n4376), .dinb(n4368), .dout(n4469));
  jand g04214(.dina(n4377), .dinb(n4283), .dout(n4470));
  jor  g04215(.dina(n4470), .dinb(n4469), .dout(n4471));
  jand g04216(.dina(n4366), .dinb(n4358), .dout(n4472));
  jand g04217(.dina(n4367), .dinb(n4286), .dout(n4473));
  jor  g04218(.dina(n4473), .dinb(n4472), .dout(n4474));
  jand g04219(.dina(n4356), .dinb(n4348), .dout(n4475));
  jand g04220(.dina(n4357), .dinb(n4289), .dout(n4476));
  jor  g04221(.dina(n4476), .dinb(n4475), .dout(n4477));
  jand g04222(.dina(n4343), .dinb(n4335), .dout(n4478));
  jand g04223(.dina(n4347), .dinb(n4344), .dout(n4479));
  jor  g04224(.dina(n4479), .dinb(n4478), .dout(n4480));
  jand g04225(.dina(n4333), .dinb(n4325), .dout(n4481));
  jand g04226(.dina(n4334), .dinb(n4292), .dout(n4482));
  jor  g04227(.dina(n4482), .dinb(n4481), .dout(n4483));
  jor  g04228(.dina(n4323), .dinb(n4315), .dout(n4484));
  jand g04229(.dina(n4324), .dinb(n4297), .dout(n4485));
  jnot g04230(.din(n4485), .dout(n4486));
  jand g04231(.dina(n4486), .dinb(n4484), .dout(n4487));
  jnot g04232(.din(n4487), .dout(n4488));
  jnot g04233(.din(n4298), .dout(n4489));
  jand g04234(.dina(n4300), .dinb(n4489), .dout(n4490));
  jand g04235(.dina(n4313), .dinb(n4302), .dout(n4491));
  jor  g04236(.dina(n4491), .dinb(n4490), .dout(n4492));
  jxor g04237(.dina(a41 ), .dinb(a40 ), .dout(n4493));
  jand g04238(.dina(n4493), .dinb(n4299), .dout(n4494));
  jand g04239(.dina(n4494), .dinb(n259), .dout(n4495));
  jnot g04240(.din(n4299), .dout(n4496));
  jxor g04241(.dina(a40 ), .dinb(a39 ), .dout(n4497));
  jand g04242(.dina(n4497), .dinb(n4496), .dout(n4498));
  jand g04243(.dina(n4498), .dinb(b0 ), .dout(n4499));
  jnot g04244(.din(n4493), .dout(n4500));
  jand g04245(.dina(n4500), .dinb(n4299), .dout(n4501));
  jand g04246(.dina(n4501), .dinb(b1 ), .dout(n4502));
  jor  g04247(.dina(n4502), .dinb(n4499), .dout(n4503));
  jor  g04248(.dina(n4503), .dinb(n4495), .dout(n4504));
  jnot g04249(.din(a41 ), .dout(n4505));
  jor  g04250(.dina(n4301), .dinb(n4505), .dout(n4506));
  jxor g04251(.dina(n4506), .dinb(n4504), .dout(n4507));
  jor  g04252(.dina(n4305), .dinb(n337), .dout(n4508));
  jor  g04253(.dina(n4303), .dinb(n340), .dout(n4509));
  jor  g04254(.dina(n4116), .dinb(n293), .dout(n4510));
  jand g04255(.dina(n4510), .dinb(n4509), .dout(n4511));
  jor  g04256(.dina(n4308), .dinb(n303), .dout(n4512));
  jand g04257(.dina(n4512), .dinb(n4511), .dout(n4513));
  jand g04258(.dina(n4513), .dinb(n4508), .dout(n4514));
  jxor g04259(.dina(n4514), .dinb(a38 ), .dout(n4515));
  jxor g04260(.dina(n4515), .dinb(n4507), .dout(n4516));
  jxor g04261(.dina(n4516), .dinb(n4492), .dout(n4517));
  jnot g04262(.din(n4517), .dout(n4518));
  jor  g04263(.dina(n3751), .dinb(n466), .dout(n4519));
  jor  g04264(.dina(n3754), .dinb(n415), .dout(n4520));
  jor  g04265(.dina(n3574), .dinb(n377), .dout(n4521));
  jand g04266(.dina(n4521), .dinb(n4520), .dout(n4522));
  jor  g04267(.dina(n3749), .dinb(n469), .dout(n4523));
  jand g04268(.dina(n4523), .dinb(n4522), .dout(n4524));
  jand g04269(.dina(n4524), .dinb(n4519), .dout(n4525));
  jxor g04270(.dina(n4525), .dinb(a35 ), .dout(n4526));
  jxor g04271(.dina(n4526), .dinb(n4518), .dout(n4527));
  jxor g04272(.dina(n4527), .dinb(n4488), .dout(n4528));
  jor  g04273(.dina(n3239), .dinb(n635), .dout(n4529));
  jor  g04274(.dina(n3072), .dinb(n519), .dout(n4530));
  jor  g04275(.dina(n3237), .dinb(n637), .dout(n4531));
  jor  g04276(.dina(n3242), .dinb(n572), .dout(n4532));
  jand g04277(.dina(n4532), .dinb(n4531), .dout(n4533));
  jand g04278(.dina(n4533), .dinb(n4530), .dout(n4534));
  jand g04279(.dina(n4534), .dinb(n4529), .dout(n4535));
  jxor g04280(.dina(n4535), .dinb(n2918), .dout(n4536));
  jxor g04281(.dina(n4536), .dinb(n4528), .dout(n4537));
  jxor g04282(.dina(n4537), .dinb(n4483), .dout(n4538));
  jor  g04283(.dina(n2764), .dinb(n850), .dout(n4539));
  jor  g04284(.dina(n2609), .dinb(n704), .dout(n4540));
  jor  g04285(.dina(n2761), .dinb(n852), .dout(n4541));
  jor  g04286(.dina(n2766), .dinb(n772), .dout(n4542));
  jand g04287(.dina(n4542), .dinb(n4541), .dout(n4543));
  jand g04288(.dina(n4543), .dinb(n4540), .dout(n4544));
  jand g04289(.dina(n4544), .dinb(n4539), .dout(n4545));
  jxor g04290(.dina(n4545), .dinb(n2468), .dout(n4546));
  jxor g04291(.dina(n4546), .dinb(n4538), .dout(n4547));
  jxor g04292(.dina(n4547), .dinb(n4480), .dout(n4548));
  jor  g04293(.dina(n2324), .dinb(n1112), .dout(n4549));
  jor  g04294(.dina(n2186), .dinb(n934), .dout(n4550));
  jor  g04295(.dina(n2326), .dinb(n1114), .dout(n4551));
  jor  g04296(.dina(n2321), .dinb(n1018), .dout(n4552));
  jand g04297(.dina(n4552), .dinb(n4551), .dout(n4553));
  jand g04298(.dina(n4553), .dinb(n4550), .dout(n4554));
  jand g04299(.dina(n4554), .dinb(n4549), .dout(n4555));
  jxor g04300(.dina(n4555), .dinb(n2057), .dout(n4556));
  jxor g04301(.dina(n4556), .dinb(n4548), .dout(n4557));
  jxor g04302(.dina(n4557), .dinb(n4477), .dout(n4558));
  jor  g04303(.dina(n1921), .dinb(n1414), .dout(n4559));
  jor  g04304(.dina(n1806), .dinb(n1211), .dout(n4560));
  jor  g04305(.dina(n1918), .dinb(n1307), .dout(n4561));
  jor  g04306(.dina(n1923), .dinb(n1416), .dout(n4562));
  jand g04307(.dina(n4562), .dinb(n4561), .dout(n4563));
  jand g04308(.dina(n4563), .dinb(n4560), .dout(n4564));
  jand g04309(.dina(n4564), .dinb(n4559), .dout(n4565));
  jxor g04310(.dina(n4565), .dinb(n1687), .dout(n4566));
  jxor g04311(.dina(n4566), .dinb(n4558), .dout(n4567));
  jxor g04312(.dina(n4567), .dinb(n4474), .dout(n4568));
  jor  g04313(.dina(n1757), .dinb(n1569), .dout(n4569));
  jor  g04314(.dina(n1453), .dinb(n1527), .dout(n4570));
  jor  g04315(.dina(n1566), .dinb(n1637), .dout(n4571));
  jor  g04316(.dina(n1571), .dinb(n1759), .dout(n4572));
  jand g04317(.dina(n4572), .dinb(n4571), .dout(n4573));
  jand g04318(.dina(n4573), .dinb(n4570), .dout(n4574));
  jand g04319(.dina(n4574), .dinb(n4569), .dout(n4575));
  jxor g04320(.dina(n4575), .dinb(n1351), .dout(n4576));
  jxor g04321(.dina(n4576), .dinb(n4568), .dout(n4577));
  jxor g04322(.dina(n4577), .dinb(n4471), .dout(n4578));
  jor  g04323(.dina(n2140), .dinb(n1248), .dout(n4579));
  jor  g04324(.dina(n1147), .dinb(n1881), .dout(n4580));
  jor  g04325(.dina(n1246), .dinb(n2142), .dout(n4581));
  jor  g04326(.dina(n1251), .dinb(n2007), .dout(n4582));
  jand g04327(.dina(n4582), .dinb(n4581), .dout(n4583));
  jand g04328(.dina(n4583), .dinb(n4580), .dout(n4584));
  jand g04329(.dina(n4584), .dinb(n4579), .dout(n4585));
  jxor g04330(.dina(n4585), .dinb(n1061), .dout(n4586));
  jxor g04331(.dina(n4586), .dinb(n4578), .dout(n4587));
  jxor g04332(.dina(n4587), .dinb(n4468), .dout(n4588));
  jor  g04333(.dina(n2561), .dinb(n970), .dout(n4589));
  jor  g04334(.dina(n880), .dinb(n2279), .dout(n4590));
  jor  g04335(.dina(n972), .dinb(n2563), .dout(n4591));
  jor  g04336(.dina(n967), .dinb(n2415), .dout(n4592));
  jand g04337(.dina(n4592), .dinb(n4591), .dout(n4593));
  jand g04338(.dina(n4593), .dinb(n4590), .dout(n4594));
  jand g04339(.dina(n4594), .dinb(n4589), .dout(n4595));
  jxor g04340(.dina(n4595), .dinb(n810), .dout(n4596));
  jxor g04341(.dina(n4596), .dinb(n4588), .dout(n4597));
  jxor g04342(.dina(n4597), .dinb(n4465), .dout(n4598));
  jor  g04343(.dina(n3021), .dinb(n728), .dout(n4599));
  jor  g04344(.dina(n660), .dinb(n2713), .dout(n4600));
  jor  g04345(.dina(n731), .dinb(n2862), .dout(n4601));
  jor  g04346(.dina(n726), .dinb(n3023), .dout(n4602));
  jand g04347(.dina(n4602), .dinb(n4601), .dout(n4603));
  jand g04348(.dina(n4603), .dinb(n4600), .dout(n4604));
  jand g04349(.dina(n4604), .dinb(n4599), .dout(n4605));
  jxor g04350(.dina(n4605), .dinb(n606), .dout(n4606));
  jxor g04351(.dina(n4606), .dinb(n4598), .dout(n4607));
  jnot g04352(.din(n4607), .dout(n4608));
  jxor g04353(.dina(n4608), .dinb(n4462), .dout(n4609));
  jor  g04354(.dina(n3520), .dinb(n544), .dout(n4610));
  jor  g04355(.dina(n486), .dinb(n3186), .dout(n4611));
  jor  g04356(.dina(n547), .dinb(n3348), .dout(n4612));
  jor  g04357(.dina(n542), .dinb(n3522), .dout(n4613));
  jand g04358(.dina(n4613), .dinb(n4612), .dout(n4614));
  jand g04359(.dina(n4614), .dinb(n4611), .dout(n4615));
  jand g04360(.dina(n4615), .dinb(n4610), .dout(n4616));
  jxor g04361(.dina(n4616), .dinb(n446), .dout(n4617));
  jxor g04362(.dina(n4617), .dinb(n4609), .dout(n4618));
  jxor g04363(.dina(n4618), .dinb(n4458), .dout(n4619));
  jor  g04364(.dina(n4058), .dinb(n397), .dout(n4620));
  jor  g04365(.dina(n354), .dinb(n3698), .dout(n4621));
  jor  g04366(.dina(n394), .dinb(n3873), .dout(n4622));
  jor  g04367(.dina(n399), .dinb(n4060), .dout(n4623));
  jand g04368(.dina(n4623), .dinb(n4622), .dout(n4624));
  jand g04369(.dina(n4624), .dinb(n4621), .dout(n4625));
  jand g04370(.dina(n4625), .dinb(n4620), .dout(n4626));
  jxor g04371(.dina(n4626), .dinb(n364), .dout(n4627));
  jxor g04372(.dina(n4627), .dinb(n4619), .dout(n4628));
  jxor g04373(.dina(n4628), .dinb(n4455), .dout(n4629));
  jand g04374(.dina(b39 ), .dinb(b38 ), .dout(n4630));
  jand g04375(.dina(n4433), .dinb(n4432), .dout(n4631));
  jor  g04376(.dina(n4631), .dinb(n4630), .dout(n4632));
  jxor g04377(.dina(b40 ), .dinb(b39 ), .dout(n4633));
  jnot g04378(.din(n4633), .dout(n4634));
  jxor g04379(.dina(n4634), .dinb(n4632), .dout(n4635));
  jor  g04380(.dina(n4635), .dinb(n296), .dout(n4636));
  jnot g04381(.din(b40 ), .dout(n4637));
  jor  g04382(.dina(n264), .dinb(n4637), .dout(n4638));
  jor  g04383(.dina(n280), .dinb(n4249), .dout(n4639));
  jor  g04384(.dina(n294), .dinb(n4437), .dout(n4640));
  jand g04385(.dina(n4640), .dinb(n4639), .dout(n4641));
  jand g04386(.dina(n4641), .dinb(n4638), .dout(n4642));
  jand g04387(.dina(n4642), .dinb(n4636), .dout(n4643));
  jxor g04388(.dina(n4643), .dinb(n278), .dout(n4644));
  jxor g04389(.dina(n4644), .dinb(n4629), .dout(n4645));
  jxor g04390(.dina(n4645), .dinb(n4450), .dout(f40 ));
  jnot g04391(.din(n4644), .dout(n4647));
  jor  g04392(.dina(n4647), .dinb(n4629), .dout(n4648));
  jor  g04393(.dina(n4645), .dinb(n4450), .dout(n4649));
  jand g04394(.dina(n4649), .dinb(n4648), .dout(n4650));
  jand g04395(.dina(n4627), .dinb(n4619), .dout(n4651));
  jnot g04396(.din(n4651), .dout(n4652));
  jnot g04397(.din(n4628), .dout(n4653));
  jor  g04398(.dina(n4653), .dinb(n4455), .dout(n4654));
  jand g04399(.dina(n4654), .dinb(n4652), .dout(n4655));
  jand g04400(.dina(n4617), .dinb(n4609), .dout(n4656));
  jand g04401(.dina(n4618), .dinb(n4458), .dout(n4657));
  jor  g04402(.dina(n4657), .dinb(n4656), .dout(n4658));
  jand g04403(.dina(n4606), .dinb(n4598), .dout(n4659));
  jnot g04404(.din(n4659), .dout(n4660));
  jor  g04405(.dina(n4608), .dinb(n4462), .dout(n4661));
  jand g04406(.dina(n4661), .dinb(n4660), .dout(n4662));
  jand g04407(.dina(n4596), .dinb(n4588), .dout(n4663));
  jand g04408(.dina(n4597), .dinb(n4465), .dout(n4664));
  jor  g04409(.dina(n4664), .dinb(n4663), .dout(n4665));
  jand g04410(.dina(n4586), .dinb(n4578), .dout(n4666));
  jand g04411(.dina(n4587), .dinb(n4468), .dout(n4667));
  jor  g04412(.dina(n4667), .dinb(n4666), .dout(n4668));
  jand g04413(.dina(n4576), .dinb(n4568), .dout(n4669));
  jand g04414(.dina(n4577), .dinb(n4471), .dout(n4670));
  jor  g04415(.dina(n4670), .dinb(n4669), .dout(n4671));
  jand g04416(.dina(n4566), .dinb(n4558), .dout(n4672));
  jand g04417(.dina(n4567), .dinb(n4474), .dout(n4673));
  jor  g04418(.dina(n4673), .dinb(n4672), .dout(n4674));
  jand g04419(.dina(n4556), .dinb(n4548), .dout(n4675));
  jand g04420(.dina(n4557), .dinb(n4477), .dout(n4676));
  jor  g04421(.dina(n4676), .dinb(n4675), .dout(n4677));
  jand g04422(.dina(n4546), .dinb(n4538), .dout(n4678));
  jand g04423(.dina(n4547), .dinb(n4480), .dout(n4679));
  jor  g04424(.dina(n4679), .dinb(n4678), .dout(n4680));
  jand g04425(.dina(n4536), .dinb(n4528), .dout(n4681));
  jand g04426(.dina(n4537), .dinb(n4483), .dout(n4682));
  jor  g04427(.dina(n4682), .dinb(n4681), .dout(n4683));
  jor  g04428(.dina(n4526), .dinb(n4518), .dout(n4684));
  jand g04429(.dina(n4527), .dinb(n4488), .dout(n4685));
  jnot g04430(.din(n4685), .dout(n4686));
  jand g04431(.dina(n4686), .dinb(n4684), .dout(n4687));
  jnot g04432(.din(n4687), .dout(n4688));
  jor  g04433(.dina(n4515), .dinb(n4507), .dout(n4689));
  jand g04434(.dina(n4516), .dinb(n4492), .dout(n4690));
  jnot g04435(.din(n4690), .dout(n4691));
  jand g04436(.dina(n4691), .dinb(n4689), .dout(n4692));
  jnot g04437(.din(n4692), .dout(n4693));
  jand g04438(.dina(n4498), .dinb(b1 ), .dout(n4694));
  jor  g04439(.dina(n4497), .dinb(n4299), .dout(n4695));
  jor  g04440(.dina(n4695), .dinb(n4500), .dout(n4696));
  jnot g04441(.din(n4696), .dout(n4697));
  jand g04442(.dina(n4697), .dinb(b0 ), .dout(n4698));
  jand g04443(.dina(n4494), .dinb(n273), .dout(n4699));
  jand g04444(.dina(n4501), .dinb(b2 ), .dout(n4700));
  jor  g04445(.dina(n4700), .dinb(n4699), .dout(n4701));
  jor  g04446(.dina(n4701), .dinb(n4698), .dout(n4702));
  jor  g04447(.dina(n4702), .dinb(n4694), .dout(n4703));
  jnot g04448(.din(n4504), .dout(n4704));
  jand g04449(.dina(n4301), .dinb(a41 ), .dout(n4705));
  jand g04450(.dina(n4705), .dinb(n4704), .dout(n4706));
  jnot g04451(.din(n4706), .dout(n4707));
  jand g04452(.dina(n4707), .dinb(a41 ), .dout(n4708));
  jxor g04453(.dina(n4708), .dinb(n4703), .dout(n4709));
  jnot g04454(.din(n4709), .dout(n4710));
  jor  g04455(.dina(n4305), .dinb(n374), .dout(n4711));
  jor  g04456(.dina(n4303), .dinb(n377), .dout(n4712));
  jor  g04457(.dina(n4116), .dinb(n303), .dout(n4713));
  jand g04458(.dina(n4713), .dinb(n4712), .dout(n4714));
  jor  g04459(.dina(n4308), .dinb(n340), .dout(n4715));
  jand g04460(.dina(n4715), .dinb(n4714), .dout(n4716));
  jand g04461(.dina(n4716), .dinb(n4711), .dout(n4717));
  jxor g04462(.dina(n4717), .dinb(a38 ), .dout(n4718));
  jxor g04463(.dina(n4718), .dinb(n4710), .dout(n4719));
  jxor g04464(.dina(n4719), .dinb(n4693), .dout(n4720));
  jor  g04465(.dina(n3751), .dinb(n517), .dout(n4721));
  jor  g04466(.dina(n3754), .dinb(n469), .dout(n4722));
  jor  g04467(.dina(n3749), .dinb(n519), .dout(n4723));
  jor  g04468(.dina(n3574), .dinb(n415), .dout(n4724));
  jand g04469(.dina(n4724), .dinb(n4723), .dout(n4725));
  jand g04470(.dina(n4725), .dinb(n4722), .dout(n4726));
  jand g04471(.dina(n4726), .dinb(n4721), .dout(n4727));
  jxor g04472(.dina(n4727), .dinb(n3410), .dout(n4728));
  jxor g04473(.dina(n4728), .dinb(n4720), .dout(n4729));
  jxor g04474(.dina(n4729), .dinb(n4688), .dout(n4730));
  jor  g04475(.dina(n3239), .dinb(n702), .dout(n4731));
  jor  g04476(.dina(n3072), .dinb(n572), .dout(n4732));
  jor  g04477(.dina(n3237), .dinb(n704), .dout(n4733));
  jor  g04478(.dina(n3242), .dinb(n637), .dout(n4734));
  jand g04479(.dina(n4734), .dinb(n4733), .dout(n4735));
  jand g04480(.dina(n4735), .dinb(n4732), .dout(n4736));
  jand g04481(.dina(n4736), .dinb(n4731), .dout(n4737));
  jxor g04482(.dina(n4737), .dinb(n2918), .dout(n4738));
  jxor g04483(.dina(n4738), .dinb(n4730), .dout(n4739));
  jxor g04484(.dina(n4739), .dinb(n4683), .dout(n4740));
  jor  g04485(.dina(n2764), .dinb(n932), .dout(n4741));
  jor  g04486(.dina(n2609), .dinb(n772), .dout(n4742));
  jor  g04487(.dina(n2761), .dinb(n934), .dout(n4743));
  jor  g04488(.dina(n2766), .dinb(n852), .dout(n4744));
  jand g04489(.dina(n4744), .dinb(n4743), .dout(n4745));
  jand g04490(.dina(n4745), .dinb(n4742), .dout(n4746));
  jand g04491(.dina(n4746), .dinb(n4741), .dout(n4747));
  jxor g04492(.dina(n4747), .dinb(n2468), .dout(n4748));
  jxor g04493(.dina(n4748), .dinb(n4740), .dout(n4749));
  jxor g04494(.dina(n4749), .dinb(n4680), .dout(n4750));
  jor  g04495(.dina(n2324), .dinb(n1209), .dout(n4751));
  jor  g04496(.dina(n2186), .dinb(n1018), .dout(n4752));
  jor  g04497(.dina(n2321), .dinb(n1114), .dout(n4753));
  jor  g04498(.dina(n2326), .dinb(n1211), .dout(n4754));
  jand g04499(.dina(n4754), .dinb(n4753), .dout(n4755));
  jand g04500(.dina(n4755), .dinb(n4752), .dout(n4756));
  jand g04501(.dina(n4756), .dinb(n4751), .dout(n4757));
  jxor g04502(.dina(n4757), .dinb(n2057), .dout(n4758));
  jxor g04503(.dina(n4758), .dinb(n4750), .dout(n4759));
  jxor g04504(.dina(n4759), .dinb(n4677), .dout(n4760));
  jor  g04505(.dina(n1921), .dinb(n1525), .dout(n4761));
  jor  g04506(.dina(n1806), .dinb(n1307), .dout(n4762));
  jor  g04507(.dina(n1918), .dinb(n1416), .dout(n4763));
  jor  g04508(.dina(n1923), .dinb(n1527), .dout(n4764));
  jand g04509(.dina(n4764), .dinb(n4763), .dout(n4765));
  jand g04510(.dina(n4765), .dinb(n4762), .dout(n4766));
  jand g04511(.dina(n4766), .dinb(n4761), .dout(n4767));
  jxor g04512(.dina(n4767), .dinb(n1687), .dout(n4768));
  jxor g04513(.dina(n4768), .dinb(n4760), .dout(n4769));
  jxor g04514(.dina(n4769), .dinb(n4674), .dout(n4770));
  jor  g04515(.dina(n1879), .dinb(n1569), .dout(n4771));
  jor  g04516(.dina(n1453), .dinb(n1637), .dout(n4772));
  jor  g04517(.dina(n1571), .dinb(n1881), .dout(n4773));
  jor  g04518(.dina(n1566), .dinb(n1759), .dout(n4774));
  jand g04519(.dina(n4774), .dinb(n4773), .dout(n4775));
  jand g04520(.dina(n4775), .dinb(n4772), .dout(n4776));
  jand g04521(.dina(n4776), .dinb(n4771), .dout(n4777));
  jxor g04522(.dina(n4777), .dinb(n1351), .dout(n4778));
  jxor g04523(.dina(n4778), .dinb(n4770), .dout(n4779));
  jxor g04524(.dina(n4779), .dinb(n4671), .dout(n4780));
  jor  g04525(.dina(n2277), .dinb(n1248), .dout(n4781));
  jor  g04526(.dina(n1147), .dinb(n2007), .dout(n4782));
  jor  g04527(.dina(n1251), .dinb(n2142), .dout(n4783));
  jor  g04528(.dina(n1246), .dinb(n2279), .dout(n4784));
  jand g04529(.dina(n4784), .dinb(n4783), .dout(n4785));
  jand g04530(.dina(n4785), .dinb(n4782), .dout(n4786));
  jand g04531(.dina(n4786), .dinb(n4781), .dout(n4787));
  jxor g04532(.dina(n4787), .dinb(n1061), .dout(n4788));
  jxor g04533(.dina(n4788), .dinb(n4780), .dout(n4789));
  jxor g04534(.dina(n4789), .dinb(n4668), .dout(n4790));
  jor  g04535(.dina(n2711), .dinb(n970), .dout(n4791));
  jor  g04536(.dina(n880), .dinb(n2415), .dout(n4792));
  jor  g04537(.dina(n967), .dinb(n2563), .dout(n4793));
  jor  g04538(.dina(n972), .dinb(n2713), .dout(n4794));
  jand g04539(.dina(n4794), .dinb(n4793), .dout(n4795));
  jand g04540(.dina(n4795), .dinb(n4792), .dout(n4796));
  jand g04541(.dina(n4796), .dinb(n4791), .dout(n4797));
  jxor g04542(.dina(n4797), .dinb(n810), .dout(n4798));
  jxor g04543(.dina(n4798), .dinb(n4790), .dout(n4799));
  jxor g04544(.dina(n4799), .dinb(n4665), .dout(n4800));
  jor  g04545(.dina(n3184), .dinb(n728), .dout(n4801));
  jor  g04546(.dina(n660), .dinb(n2862), .dout(n4802));
  jor  g04547(.dina(n726), .dinb(n3186), .dout(n4803));
  jor  g04548(.dina(n731), .dinb(n3023), .dout(n4804));
  jand g04549(.dina(n4804), .dinb(n4803), .dout(n4805));
  jand g04550(.dina(n4805), .dinb(n4802), .dout(n4806));
  jand g04551(.dina(n4806), .dinb(n4801), .dout(n4807));
  jxor g04552(.dina(n4807), .dinb(n606), .dout(n4808));
  jxor g04553(.dina(n4808), .dinb(n4800), .dout(n4809));
  jnot g04554(.din(n4809), .dout(n4810));
  jxor g04555(.dina(n4810), .dinb(n4662), .dout(n4811));
  jor  g04556(.dina(n3696), .dinb(n544), .dout(n4812));
  jor  g04557(.dina(n486), .dinb(n3348), .dout(n4813));
  jor  g04558(.dina(n542), .dinb(n3698), .dout(n4814));
  jor  g04559(.dina(n547), .dinb(n3522), .dout(n4815));
  jand g04560(.dina(n4815), .dinb(n4814), .dout(n4816));
  jand g04561(.dina(n4816), .dinb(n4813), .dout(n4817));
  jand g04562(.dina(n4817), .dinb(n4812), .dout(n4818));
  jxor g04563(.dina(n4818), .dinb(n446), .dout(n4819));
  jxor g04564(.dina(n4819), .dinb(n4811), .dout(n4820));
  jxor g04565(.dina(n4820), .dinb(n4658), .dout(n4821));
  jor  g04566(.dina(n4247), .dinb(n397), .dout(n4822));
  jor  g04567(.dina(n354), .dinb(n3873), .dout(n4823));
  jor  g04568(.dina(n399), .dinb(n4249), .dout(n4824));
  jor  g04569(.dina(n394), .dinb(n4060), .dout(n4825));
  jand g04570(.dina(n4825), .dinb(n4824), .dout(n4826));
  jand g04571(.dina(n4826), .dinb(n4823), .dout(n4827));
  jand g04572(.dina(n4827), .dinb(n4822), .dout(n4828));
  jxor g04573(.dina(n4828), .dinb(n364), .dout(n4829));
  jxor g04574(.dina(n4829), .dinb(n4821), .dout(n4830));
  jxor g04575(.dina(n4830), .dinb(n4655), .dout(n4831));
  jand g04576(.dina(b40 ), .dinb(b39 ), .dout(n4832));
  jand g04577(.dina(n4633), .dinb(n4632), .dout(n4833));
  jor  g04578(.dina(n4833), .dinb(n4832), .dout(n4834));
  jxor g04579(.dina(b41 ), .dinb(b40 ), .dout(n4835));
  jnot g04580(.din(n4835), .dout(n4836));
  jxor g04581(.dina(n4836), .dinb(n4834), .dout(n4837));
  jor  g04582(.dina(n4837), .dinb(n296), .dout(n4838));
  jnot g04583(.din(b41 ), .dout(n4839));
  jor  g04584(.dina(n264), .dinb(n4839), .dout(n4840));
  jor  g04585(.dina(n294), .dinb(n4637), .dout(n4841));
  jor  g04586(.dina(n280), .dinb(n4437), .dout(n4842));
  jand g04587(.dina(n4842), .dinb(n4841), .dout(n4843));
  jand g04588(.dina(n4843), .dinb(n4840), .dout(n4844));
  jand g04589(.dina(n4844), .dinb(n4838), .dout(n4845));
  jxor g04590(.dina(n4845), .dinb(n278), .dout(n4846));
  jxor g04591(.dina(n4846), .dinb(n4831), .dout(n4847));
  jxor g04592(.dina(n4847), .dinb(n4650), .dout(f41 ));
  jnot g04593(.din(n4846), .dout(n4849));
  jor  g04594(.dina(n4849), .dinb(n4831), .dout(n4850));
  jor  g04595(.dina(n4847), .dinb(n4650), .dout(n4851));
  jand g04596(.dina(n4851), .dinb(n4850), .dout(n4852));
  jand g04597(.dina(n4829), .dinb(n4821), .dout(n4853));
  jnot g04598(.din(n4853), .dout(n4854));
  jnot g04599(.din(n4830), .dout(n4855));
  jor  g04600(.dina(n4855), .dinb(n4655), .dout(n4856));
  jand g04601(.dina(n4856), .dinb(n4854), .dout(n4857));
  jand g04602(.dina(n4819), .dinb(n4811), .dout(n4858));
  jand g04603(.dina(n4820), .dinb(n4658), .dout(n4859));
  jor  g04604(.dina(n4859), .dinb(n4858), .dout(n4860));
  jand g04605(.dina(n4808), .dinb(n4800), .dout(n4861));
  jnot g04606(.din(n4861), .dout(n4862));
  jor  g04607(.dina(n4810), .dinb(n4662), .dout(n4863));
  jand g04608(.dina(n4863), .dinb(n4862), .dout(n4864));
  jand g04609(.dina(n4798), .dinb(n4790), .dout(n4865));
  jand g04610(.dina(n4799), .dinb(n4665), .dout(n4866));
  jor  g04611(.dina(n4866), .dinb(n4865), .dout(n4867));
  jand g04612(.dina(n4788), .dinb(n4780), .dout(n4868));
  jand g04613(.dina(n4789), .dinb(n4668), .dout(n4869));
  jor  g04614(.dina(n4869), .dinb(n4868), .dout(n4870));
  jand g04615(.dina(n4778), .dinb(n4770), .dout(n4871));
  jand g04616(.dina(n4779), .dinb(n4671), .dout(n4872));
  jor  g04617(.dina(n4872), .dinb(n4871), .dout(n4873));
  jand g04618(.dina(n4768), .dinb(n4760), .dout(n4874));
  jand g04619(.dina(n4769), .dinb(n4674), .dout(n4875));
  jor  g04620(.dina(n4875), .dinb(n4874), .dout(n4876));
  jand g04621(.dina(n4758), .dinb(n4750), .dout(n4877));
  jand g04622(.dina(n4759), .dinb(n4677), .dout(n4878));
  jor  g04623(.dina(n4878), .dinb(n4877), .dout(n4879));
  jand g04624(.dina(n4748), .dinb(n4740), .dout(n4880));
  jand g04625(.dina(n4749), .dinb(n4680), .dout(n4881));
  jor  g04626(.dina(n4881), .dinb(n4880), .dout(n4882));
  jand g04627(.dina(n4738), .dinb(n4730), .dout(n4883));
  jand g04628(.dina(n4739), .dinb(n4683), .dout(n4884));
  jor  g04629(.dina(n4884), .dinb(n4883), .dout(n4885));
  jand g04630(.dina(n4728), .dinb(n4720), .dout(n4886));
  jand g04631(.dina(n4729), .dinb(n4688), .dout(n4887));
  jor  g04632(.dina(n4887), .dinb(n4886), .dout(n4888));
  jor  g04633(.dina(n4718), .dinb(n4710), .dout(n4889));
  jand g04634(.dina(n4719), .dinb(n4693), .dout(n4890));
  jnot g04635(.din(n4890), .dout(n4891));
  jand g04636(.dina(n4891), .dinb(n4889), .dout(n4892));
  jnot g04637(.din(n4892), .dout(n4893));
  jor  g04638(.dina(n4707), .dinb(n4703), .dout(n4894));
  jxor g04639(.dina(a42 ), .dinb(a41 ), .dout(n4895));
  jand g04640(.dina(n4895), .dinb(b0 ), .dout(n4896));
  jnot g04641(.din(n4896), .dout(n4897));
  jxor g04642(.dina(n4897), .dinb(n4894), .dout(n4898));
  jnot g04643(.din(n4501), .dout(n4899));
  jor  g04644(.dina(n4899), .dinb(n303), .dout(n4900));
  jor  g04645(.dina(n4696), .dinb(n305), .dout(n4901));
  jnot g04646(.din(n4494), .dout(n4902));
  jor  g04647(.dina(n4902), .dinb(n301), .dout(n4903));
  jnot g04648(.din(n4498), .dout(n4904));
  jor  g04649(.dina(n4904), .dinb(n293), .dout(n4905));
  jand g04650(.dina(n4905), .dinb(n4903), .dout(n4906));
  jand g04651(.dina(n4906), .dinb(n4901), .dout(n4907));
  jand g04652(.dina(n4907), .dinb(n4900), .dout(n4908));
  jxor g04653(.dina(n4908), .dinb(n4505), .dout(n4909));
  jxor g04654(.dina(n4909), .dinb(n4898), .dout(n4910));
  jnot g04655(.din(n4910), .dout(n4911));
  jor  g04656(.dina(n4305), .dinb(n412), .dout(n4912));
  jor  g04657(.dina(n4303), .dinb(n415), .dout(n4913));
  jor  g04658(.dina(n4116), .dinb(n340), .dout(n4914));
  jand g04659(.dina(n4914), .dinb(n4913), .dout(n4915));
  jor  g04660(.dina(n4308), .dinb(n377), .dout(n4916));
  jand g04661(.dina(n4916), .dinb(n4915), .dout(n4917));
  jand g04662(.dina(n4917), .dinb(n4912), .dout(n4918));
  jxor g04663(.dina(n4918), .dinb(a38 ), .dout(n4919));
  jxor g04664(.dina(n4919), .dinb(n4911), .dout(n4920));
  jxor g04665(.dina(n4920), .dinb(n4893), .dout(n4921));
  jor  g04666(.dina(n3751), .dinb(n570), .dout(n4922));
  jor  g04667(.dina(n3574), .dinb(n469), .dout(n4923));
  jor  g04668(.dina(n3749), .dinb(n572), .dout(n4924));
  jor  g04669(.dina(n3754), .dinb(n519), .dout(n4925));
  jand g04670(.dina(n4925), .dinb(n4924), .dout(n4926));
  jand g04671(.dina(n4926), .dinb(n4923), .dout(n4927));
  jand g04672(.dina(n4927), .dinb(n4922), .dout(n4928));
  jxor g04673(.dina(n4928), .dinb(n3410), .dout(n4929));
  jxor g04674(.dina(n4929), .dinb(n4921), .dout(n4930));
  jxor g04675(.dina(n4930), .dinb(n4888), .dout(n4931));
  jor  g04676(.dina(n3239), .dinb(n770), .dout(n4932));
  jor  g04677(.dina(n3072), .dinb(n637), .dout(n4933));
  jor  g04678(.dina(n3242), .dinb(n704), .dout(n4934));
  jor  g04679(.dina(n3237), .dinb(n772), .dout(n4935));
  jand g04680(.dina(n4935), .dinb(n4934), .dout(n4936));
  jand g04681(.dina(n4936), .dinb(n4933), .dout(n4937));
  jand g04682(.dina(n4937), .dinb(n4932), .dout(n4938));
  jxor g04683(.dina(n4938), .dinb(n2918), .dout(n4939));
  jxor g04684(.dina(n4939), .dinb(n4931), .dout(n4940));
  jxor g04685(.dina(n4940), .dinb(n4885), .dout(n4941));
  jor  g04686(.dina(n2764), .dinb(n1016), .dout(n4942));
  jor  g04687(.dina(n2609), .dinb(n852), .dout(n4943));
  jor  g04688(.dina(n2761), .dinb(n1018), .dout(n4944));
  jor  g04689(.dina(n2766), .dinb(n934), .dout(n4945));
  jand g04690(.dina(n4945), .dinb(n4944), .dout(n4946));
  jand g04691(.dina(n4946), .dinb(n4943), .dout(n4947));
  jand g04692(.dina(n4947), .dinb(n4942), .dout(n4948));
  jxor g04693(.dina(n4948), .dinb(n2468), .dout(n4949));
  jxor g04694(.dina(n4949), .dinb(n4941), .dout(n4950));
  jxor g04695(.dina(n4950), .dinb(n4882), .dout(n4951));
  jor  g04696(.dina(n2324), .dinb(n1305), .dout(n4952));
  jor  g04697(.dina(n2186), .dinb(n1114), .dout(n4953));
  jor  g04698(.dina(n2326), .dinb(n1307), .dout(n4954));
  jor  g04699(.dina(n2321), .dinb(n1211), .dout(n4955));
  jand g04700(.dina(n4955), .dinb(n4954), .dout(n4956));
  jand g04701(.dina(n4956), .dinb(n4953), .dout(n4957));
  jand g04702(.dina(n4957), .dinb(n4952), .dout(n4958));
  jxor g04703(.dina(n4958), .dinb(n2057), .dout(n4959));
  jxor g04704(.dina(n4959), .dinb(n4951), .dout(n4960));
  jxor g04705(.dina(n4960), .dinb(n4879), .dout(n4961));
  jor  g04706(.dina(n1921), .dinb(n1635), .dout(n4962));
  jor  g04707(.dina(n1806), .dinb(n1416), .dout(n4963));
  jor  g04708(.dina(n1918), .dinb(n1527), .dout(n4964));
  jor  g04709(.dina(n1923), .dinb(n1637), .dout(n4965));
  jand g04710(.dina(n4965), .dinb(n4964), .dout(n4966));
  jand g04711(.dina(n4966), .dinb(n4963), .dout(n4967));
  jand g04712(.dina(n4967), .dinb(n4962), .dout(n4968));
  jxor g04713(.dina(n4968), .dinb(n1687), .dout(n4969));
  jxor g04714(.dina(n4969), .dinb(n4961), .dout(n4970));
  jxor g04715(.dina(n4970), .dinb(n4876), .dout(n4971));
  jor  g04716(.dina(n2005), .dinb(n1569), .dout(n4972));
  jor  g04717(.dina(n1453), .dinb(n1759), .dout(n4973));
  jor  g04718(.dina(n1566), .dinb(n1881), .dout(n4974));
  jor  g04719(.dina(n1571), .dinb(n2007), .dout(n4975));
  jand g04720(.dina(n4975), .dinb(n4974), .dout(n4976));
  jand g04721(.dina(n4976), .dinb(n4973), .dout(n4977));
  jand g04722(.dina(n4977), .dinb(n4972), .dout(n4978));
  jxor g04723(.dina(n4978), .dinb(n1351), .dout(n4979));
  jxor g04724(.dina(n4979), .dinb(n4971), .dout(n4980));
  jxor g04725(.dina(n4980), .dinb(n4873), .dout(n4981));
  jor  g04726(.dina(n2413), .dinb(n1248), .dout(n4982));
  jor  g04727(.dina(n1147), .dinb(n2142), .dout(n4983));
  jor  g04728(.dina(n1251), .dinb(n2279), .dout(n4984));
  jor  g04729(.dina(n1246), .dinb(n2415), .dout(n4985));
  jand g04730(.dina(n4985), .dinb(n4984), .dout(n4986));
  jand g04731(.dina(n4986), .dinb(n4983), .dout(n4987));
  jand g04732(.dina(n4987), .dinb(n4982), .dout(n4988));
  jxor g04733(.dina(n4988), .dinb(n1061), .dout(n4989));
  jxor g04734(.dina(n4989), .dinb(n4981), .dout(n4990));
  jxor g04735(.dina(n4990), .dinb(n4870), .dout(n4991));
  jor  g04736(.dina(n2860), .dinb(n970), .dout(n4992));
  jor  g04737(.dina(n880), .dinb(n2563), .dout(n4993));
  jor  g04738(.dina(n967), .dinb(n2713), .dout(n4994));
  jor  g04739(.dina(n972), .dinb(n2862), .dout(n4995));
  jand g04740(.dina(n4995), .dinb(n4994), .dout(n4996));
  jand g04741(.dina(n4996), .dinb(n4993), .dout(n4997));
  jand g04742(.dina(n4997), .dinb(n4992), .dout(n4998));
  jxor g04743(.dina(n4998), .dinb(n810), .dout(n4999));
  jxor g04744(.dina(n4999), .dinb(n4991), .dout(n5000));
  jxor g04745(.dina(n5000), .dinb(n4867), .dout(n5001));
  jor  g04746(.dina(n3346), .dinb(n728), .dout(n5002));
  jor  g04747(.dina(n660), .dinb(n3023), .dout(n5003));
  jor  g04748(.dina(n726), .dinb(n3348), .dout(n5004));
  jor  g04749(.dina(n731), .dinb(n3186), .dout(n5005));
  jand g04750(.dina(n5005), .dinb(n5004), .dout(n5006));
  jand g04751(.dina(n5006), .dinb(n5003), .dout(n5007));
  jand g04752(.dina(n5007), .dinb(n5002), .dout(n5008));
  jxor g04753(.dina(n5008), .dinb(n606), .dout(n5009));
  jxor g04754(.dina(n5009), .dinb(n5001), .dout(n5010));
  jnot g04755(.din(n5010), .dout(n5011));
  jxor g04756(.dina(n5011), .dinb(n4864), .dout(n5012));
  jor  g04757(.dina(n3871), .dinb(n544), .dout(n5013));
  jor  g04758(.dina(n486), .dinb(n3522), .dout(n5014));
  jor  g04759(.dina(n542), .dinb(n3873), .dout(n5015));
  jor  g04760(.dina(n547), .dinb(n3698), .dout(n5016));
  jand g04761(.dina(n5016), .dinb(n5015), .dout(n5017));
  jand g04762(.dina(n5017), .dinb(n5014), .dout(n5018));
  jand g04763(.dina(n5018), .dinb(n5013), .dout(n5019));
  jxor g04764(.dina(n5019), .dinb(n446), .dout(n5020));
  jxor g04765(.dina(n5020), .dinb(n5012), .dout(n5021));
  jxor g04766(.dina(n5021), .dinb(n4860), .dout(n5022));
  jor  g04767(.dina(n4435), .dinb(n397), .dout(n5023));
  jor  g04768(.dina(n354), .dinb(n4060), .dout(n5024));
  jor  g04769(.dina(n399), .dinb(n4437), .dout(n5025));
  jor  g04770(.dina(n394), .dinb(n4249), .dout(n5026));
  jand g04771(.dina(n5026), .dinb(n5025), .dout(n5027));
  jand g04772(.dina(n5027), .dinb(n5024), .dout(n5028));
  jand g04773(.dina(n5028), .dinb(n5023), .dout(n5029));
  jxor g04774(.dina(n5029), .dinb(n364), .dout(n5030));
  jxor g04775(.dina(n5030), .dinb(n5022), .dout(n5031));
  jxor g04776(.dina(n5031), .dinb(n4857), .dout(n5032));
  jand g04777(.dina(b41 ), .dinb(b40 ), .dout(n5033));
  jand g04778(.dina(n4835), .dinb(n4834), .dout(n5034));
  jor  g04779(.dina(n5034), .dinb(n5033), .dout(n5035));
  jxor g04780(.dina(b42 ), .dinb(b41 ), .dout(n5036));
  jnot g04781(.din(n5036), .dout(n5037));
  jxor g04782(.dina(n5037), .dinb(n5035), .dout(n5038));
  jor  g04783(.dina(n5038), .dinb(n296), .dout(n5039));
  jnot g04784(.din(b42 ), .dout(n5040));
  jor  g04785(.dina(n264), .dinb(n5040), .dout(n5041));
  jor  g04786(.dina(n294), .dinb(n4839), .dout(n5042));
  jor  g04787(.dina(n280), .dinb(n4637), .dout(n5043));
  jand g04788(.dina(n5043), .dinb(n5042), .dout(n5044));
  jand g04789(.dina(n5044), .dinb(n5041), .dout(n5045));
  jand g04790(.dina(n5045), .dinb(n5039), .dout(n5046));
  jxor g04791(.dina(n5046), .dinb(n278), .dout(n5047));
  jxor g04792(.dina(n5047), .dinb(n5032), .dout(n5048));
  jxor g04793(.dina(n5048), .dinb(n4852), .dout(f42 ));
  jnot g04794(.din(n5047), .dout(n5050));
  jor  g04795(.dina(n5050), .dinb(n5032), .dout(n5051));
  jor  g04796(.dina(n5048), .dinb(n4852), .dout(n5052));
  jand g04797(.dina(n5052), .dinb(n5051), .dout(n5053));
  jand g04798(.dina(n5030), .dinb(n5022), .dout(n5054));
  jnot g04799(.din(n5054), .dout(n5055));
  jnot g04800(.din(n5031), .dout(n5056));
  jor  g04801(.dina(n5056), .dinb(n4857), .dout(n5057));
  jand g04802(.dina(n5057), .dinb(n5055), .dout(n5058));
  jand g04803(.dina(n5020), .dinb(n5012), .dout(n5059));
  jand g04804(.dina(n5021), .dinb(n4860), .dout(n5060));
  jor  g04805(.dina(n5060), .dinb(n5059), .dout(n5061));
  jand g04806(.dina(n5009), .dinb(n5001), .dout(n5062));
  jnot g04807(.din(n5062), .dout(n5063));
  jor  g04808(.dina(n5011), .dinb(n4864), .dout(n5064));
  jand g04809(.dina(n5064), .dinb(n5063), .dout(n5065));
  jand g04810(.dina(n4999), .dinb(n4991), .dout(n5066));
  jand g04811(.dina(n5000), .dinb(n4867), .dout(n5067));
  jor  g04812(.dina(n5067), .dinb(n5066), .dout(n5068));
  jand g04813(.dina(n4989), .dinb(n4981), .dout(n5069));
  jand g04814(.dina(n4990), .dinb(n4870), .dout(n5070));
  jor  g04815(.dina(n5070), .dinb(n5069), .dout(n5071));
  jand g04816(.dina(n4979), .dinb(n4971), .dout(n5072));
  jand g04817(.dina(n4980), .dinb(n4873), .dout(n5073));
  jor  g04818(.dina(n5073), .dinb(n5072), .dout(n5074));
  jand g04819(.dina(n4969), .dinb(n4961), .dout(n5075));
  jand g04820(.dina(n4970), .dinb(n4876), .dout(n5076));
  jor  g04821(.dina(n5076), .dinb(n5075), .dout(n5077));
  jand g04822(.dina(n4959), .dinb(n4951), .dout(n5078));
  jand g04823(.dina(n4960), .dinb(n4879), .dout(n5079));
  jor  g04824(.dina(n5079), .dinb(n5078), .dout(n5080));
  jand g04825(.dina(n4949), .dinb(n4941), .dout(n5081));
  jand g04826(.dina(n4950), .dinb(n4882), .dout(n5082));
  jor  g04827(.dina(n5082), .dinb(n5081), .dout(n5083));
  jand g04828(.dina(n4939), .dinb(n4931), .dout(n5084));
  jand g04829(.dina(n4940), .dinb(n4885), .dout(n5085));
  jor  g04830(.dina(n5085), .dinb(n5084), .dout(n5086));
  jand g04831(.dina(n4929), .dinb(n4921), .dout(n5087));
  jand g04832(.dina(n4930), .dinb(n4888), .dout(n5088));
  jor  g04833(.dina(n5088), .dinb(n5087), .dout(n5089));
  jor  g04834(.dina(n4919), .dinb(n4911), .dout(n5090));
  jand g04835(.dina(n4920), .dinb(n4893), .dout(n5091));
  jnot g04836(.din(n5091), .dout(n5092));
  jand g04837(.dina(n5092), .dinb(n5090), .dout(n5093));
  jnot g04838(.din(n5093), .dout(n5094));
  jnot g04839(.din(n4894), .dout(n5095));
  jand g04840(.dina(n4896), .dinb(n5095), .dout(n5096));
  jand g04841(.dina(n4909), .dinb(n4898), .dout(n5097));
  jor  g04842(.dina(n5097), .dinb(n5096), .dout(n5098));
  jxor g04843(.dina(a44 ), .dinb(a43 ), .dout(n5099));
  jand g04844(.dina(n5099), .dinb(n4895), .dout(n5100));
  jand g04845(.dina(n5100), .dinb(n259), .dout(n5101));
  jnot g04846(.din(n4895), .dout(n5102));
  jxor g04847(.dina(a43 ), .dinb(a42 ), .dout(n5103));
  jand g04848(.dina(n5103), .dinb(n5102), .dout(n5104));
  jand g04849(.dina(n5104), .dinb(b0 ), .dout(n5105));
  jnot g04850(.din(n5099), .dout(n5106));
  jand g04851(.dina(n5106), .dinb(n4895), .dout(n5107));
  jand g04852(.dina(n5107), .dinb(b1 ), .dout(n5108));
  jor  g04853(.dina(n5108), .dinb(n5105), .dout(n5109));
  jor  g04854(.dina(n5109), .dinb(n5101), .dout(n5110));
  jnot g04855(.din(a44 ), .dout(n5111));
  jor  g04856(.dina(n4897), .dinb(n5111), .dout(n5112));
  jxor g04857(.dina(n5112), .dinb(n5110), .dout(n5113));
  jor  g04858(.dina(n4902), .dinb(n337), .dout(n5114));
  jor  g04859(.dina(n4899), .dinb(n340), .dout(n5115));
  jor  g04860(.dina(n4696), .dinb(n293), .dout(n5116));
  jand g04861(.dina(n5116), .dinb(n5115), .dout(n5117));
  jor  g04862(.dina(n4904), .dinb(n303), .dout(n5118));
  jand g04863(.dina(n5118), .dinb(n5117), .dout(n5119));
  jand g04864(.dina(n5119), .dinb(n5114), .dout(n5120));
  jxor g04865(.dina(n5120), .dinb(a41 ), .dout(n5121));
  jxor g04866(.dina(n5121), .dinb(n5113), .dout(n5122));
  jxor g04867(.dina(n5122), .dinb(n5098), .dout(n5123));
  jnot g04868(.din(n5123), .dout(n5124));
  jor  g04869(.dina(n4305), .dinb(n466), .dout(n5125));
  jor  g04870(.dina(n4308), .dinb(n415), .dout(n5126));
  jor  g04871(.dina(n4116), .dinb(n377), .dout(n5127));
  jand g04872(.dina(n5127), .dinb(n5126), .dout(n5128));
  jor  g04873(.dina(n4303), .dinb(n469), .dout(n5129));
  jand g04874(.dina(n5129), .dinb(n5128), .dout(n5130));
  jand g04875(.dina(n5130), .dinb(n5125), .dout(n5131));
  jxor g04876(.dina(n5131), .dinb(a38 ), .dout(n5132));
  jxor g04877(.dina(n5132), .dinb(n5124), .dout(n5133));
  jxor g04878(.dina(n5133), .dinb(n5094), .dout(n5134));
  jor  g04879(.dina(n3751), .dinb(n635), .dout(n5135));
  jor  g04880(.dina(n3574), .dinb(n519), .dout(n5136));
  jor  g04881(.dina(n3749), .dinb(n637), .dout(n5137));
  jor  g04882(.dina(n3754), .dinb(n572), .dout(n5138));
  jand g04883(.dina(n5138), .dinb(n5137), .dout(n5139));
  jand g04884(.dina(n5139), .dinb(n5136), .dout(n5140));
  jand g04885(.dina(n5140), .dinb(n5135), .dout(n5141));
  jxor g04886(.dina(n5141), .dinb(n3410), .dout(n5142));
  jxor g04887(.dina(n5142), .dinb(n5134), .dout(n5143));
  jxor g04888(.dina(n5143), .dinb(n5089), .dout(n5144));
  jor  g04889(.dina(n3239), .dinb(n850), .dout(n5145));
  jor  g04890(.dina(n3072), .dinb(n704), .dout(n5146));
  jor  g04891(.dina(n3242), .dinb(n772), .dout(n5147));
  jor  g04892(.dina(n3237), .dinb(n852), .dout(n5148));
  jand g04893(.dina(n5148), .dinb(n5147), .dout(n5149));
  jand g04894(.dina(n5149), .dinb(n5146), .dout(n5150));
  jand g04895(.dina(n5150), .dinb(n5145), .dout(n5151));
  jxor g04896(.dina(n5151), .dinb(n2918), .dout(n5152));
  jxor g04897(.dina(n5152), .dinb(n5144), .dout(n5153));
  jxor g04898(.dina(n5153), .dinb(n5086), .dout(n5154));
  jor  g04899(.dina(n2764), .dinb(n1112), .dout(n5155));
  jor  g04900(.dina(n2609), .dinb(n934), .dout(n5156));
  jor  g04901(.dina(n2761), .dinb(n1114), .dout(n5157));
  jor  g04902(.dina(n2766), .dinb(n1018), .dout(n5158));
  jand g04903(.dina(n5158), .dinb(n5157), .dout(n5159));
  jand g04904(.dina(n5159), .dinb(n5156), .dout(n5160));
  jand g04905(.dina(n5160), .dinb(n5155), .dout(n5161));
  jxor g04906(.dina(n5161), .dinb(n2468), .dout(n5162));
  jxor g04907(.dina(n5162), .dinb(n5154), .dout(n5163));
  jxor g04908(.dina(n5163), .dinb(n5083), .dout(n5164));
  jor  g04909(.dina(n2324), .dinb(n1414), .dout(n5165));
  jor  g04910(.dina(n2186), .dinb(n1211), .dout(n5166));
  jor  g04911(.dina(n2321), .dinb(n1307), .dout(n5167));
  jor  g04912(.dina(n2326), .dinb(n1416), .dout(n5168));
  jand g04913(.dina(n5168), .dinb(n5167), .dout(n5169));
  jand g04914(.dina(n5169), .dinb(n5166), .dout(n5170));
  jand g04915(.dina(n5170), .dinb(n5165), .dout(n5171));
  jxor g04916(.dina(n5171), .dinb(n2057), .dout(n5172));
  jxor g04917(.dina(n5172), .dinb(n5164), .dout(n5173));
  jxor g04918(.dina(n5173), .dinb(n5080), .dout(n5174));
  jor  g04919(.dina(n1757), .dinb(n1921), .dout(n5175));
  jor  g04920(.dina(n1806), .dinb(n1527), .dout(n5176));
  jor  g04921(.dina(n1923), .dinb(n1759), .dout(n5177));
  jor  g04922(.dina(n1918), .dinb(n1637), .dout(n5178));
  jand g04923(.dina(n5178), .dinb(n5177), .dout(n5179));
  jand g04924(.dina(n5179), .dinb(n5176), .dout(n5180));
  jand g04925(.dina(n5180), .dinb(n5175), .dout(n5181));
  jxor g04926(.dina(n5181), .dinb(n1687), .dout(n5182));
  jxor g04927(.dina(n5182), .dinb(n5174), .dout(n5183));
  jxor g04928(.dina(n5183), .dinb(n5077), .dout(n5184));
  jor  g04929(.dina(n2140), .dinb(n1569), .dout(n5185));
  jor  g04930(.dina(n1453), .dinb(n1881), .dout(n5186));
  jor  g04931(.dina(n1566), .dinb(n2007), .dout(n5187));
  jor  g04932(.dina(n1571), .dinb(n2142), .dout(n5188));
  jand g04933(.dina(n5188), .dinb(n5187), .dout(n5189));
  jand g04934(.dina(n5189), .dinb(n5186), .dout(n5190));
  jand g04935(.dina(n5190), .dinb(n5185), .dout(n5191));
  jxor g04936(.dina(n5191), .dinb(n1351), .dout(n5192));
  jxor g04937(.dina(n5192), .dinb(n5184), .dout(n5193));
  jxor g04938(.dina(n5193), .dinb(n5074), .dout(n5194));
  jor  g04939(.dina(n2561), .dinb(n1248), .dout(n5195));
  jor  g04940(.dina(n1147), .dinb(n2279), .dout(n5196));
  jor  g04941(.dina(n1251), .dinb(n2415), .dout(n5197));
  jor  g04942(.dina(n1246), .dinb(n2563), .dout(n5198));
  jand g04943(.dina(n5198), .dinb(n5197), .dout(n5199));
  jand g04944(.dina(n5199), .dinb(n5196), .dout(n5200));
  jand g04945(.dina(n5200), .dinb(n5195), .dout(n5201));
  jxor g04946(.dina(n5201), .dinb(n1061), .dout(n5202));
  jxor g04947(.dina(n5202), .dinb(n5194), .dout(n5203));
  jxor g04948(.dina(n5203), .dinb(n5071), .dout(n5204));
  jor  g04949(.dina(n3021), .dinb(n970), .dout(n5205));
  jor  g04950(.dina(n880), .dinb(n2713), .dout(n5206));
  jor  g04951(.dina(n972), .dinb(n3023), .dout(n5207));
  jor  g04952(.dina(n967), .dinb(n2862), .dout(n5208));
  jand g04953(.dina(n5208), .dinb(n5207), .dout(n5209));
  jand g04954(.dina(n5209), .dinb(n5206), .dout(n5210));
  jand g04955(.dina(n5210), .dinb(n5205), .dout(n5211));
  jxor g04956(.dina(n5211), .dinb(n810), .dout(n5212));
  jxor g04957(.dina(n5212), .dinb(n5204), .dout(n5213));
  jxor g04958(.dina(n5213), .dinb(n5068), .dout(n5214));
  jor  g04959(.dina(n3520), .dinb(n728), .dout(n5215));
  jor  g04960(.dina(n660), .dinb(n3186), .dout(n5216));
  jor  g04961(.dina(n726), .dinb(n3522), .dout(n5217));
  jor  g04962(.dina(n731), .dinb(n3348), .dout(n5218));
  jand g04963(.dina(n5218), .dinb(n5217), .dout(n5219));
  jand g04964(.dina(n5219), .dinb(n5216), .dout(n5220));
  jand g04965(.dina(n5220), .dinb(n5215), .dout(n5221));
  jxor g04966(.dina(n5221), .dinb(n606), .dout(n5222));
  jxor g04967(.dina(n5222), .dinb(n5214), .dout(n5223));
  jnot g04968(.din(n5223), .dout(n5224));
  jxor g04969(.dina(n5224), .dinb(n5065), .dout(n5225));
  jor  g04970(.dina(n4058), .dinb(n544), .dout(n5226));
  jor  g04971(.dina(n486), .dinb(n3698), .dout(n5227));
  jor  g04972(.dina(n547), .dinb(n3873), .dout(n5228));
  jor  g04973(.dina(n542), .dinb(n4060), .dout(n5229));
  jand g04974(.dina(n5229), .dinb(n5228), .dout(n5230));
  jand g04975(.dina(n5230), .dinb(n5227), .dout(n5231));
  jand g04976(.dina(n5231), .dinb(n5226), .dout(n5232));
  jxor g04977(.dina(n5232), .dinb(n446), .dout(n5233));
  jxor g04978(.dina(n5233), .dinb(n5225), .dout(n5234));
  jxor g04979(.dina(n5234), .dinb(n5061), .dout(n5235));
  jor  g04980(.dina(n4635), .dinb(n397), .dout(n5236));
  jor  g04981(.dina(n354), .dinb(n4249), .dout(n5237));
  jor  g04982(.dina(n394), .dinb(n4437), .dout(n5238));
  jor  g04983(.dina(n399), .dinb(n4637), .dout(n5239));
  jand g04984(.dina(n5239), .dinb(n5238), .dout(n5240));
  jand g04985(.dina(n5240), .dinb(n5237), .dout(n5241));
  jand g04986(.dina(n5241), .dinb(n5236), .dout(n5242));
  jxor g04987(.dina(n5242), .dinb(n364), .dout(n5243));
  jxor g04988(.dina(n5243), .dinb(n5235), .dout(n5244));
  jxor g04989(.dina(n5244), .dinb(n5058), .dout(n5245));
  jand g04990(.dina(b42 ), .dinb(b41 ), .dout(n5246));
  jand g04991(.dina(n5036), .dinb(n5035), .dout(n5247));
  jor  g04992(.dina(n5247), .dinb(n5246), .dout(n5248));
  jxor g04993(.dina(b43 ), .dinb(b42 ), .dout(n5249));
  jnot g04994(.din(n5249), .dout(n5250));
  jxor g04995(.dina(n5250), .dinb(n5248), .dout(n5251));
  jor  g04996(.dina(n5251), .dinb(n296), .dout(n5252));
  jnot g04997(.din(b43 ), .dout(n5253));
  jor  g04998(.dina(n264), .dinb(n5253), .dout(n5254));
  jor  g04999(.dina(n294), .dinb(n5040), .dout(n5255));
  jor  g05000(.dina(n280), .dinb(n4839), .dout(n5256));
  jand g05001(.dina(n5256), .dinb(n5255), .dout(n5257));
  jand g05002(.dina(n5257), .dinb(n5254), .dout(n5258));
  jand g05003(.dina(n5258), .dinb(n5252), .dout(n5259));
  jxor g05004(.dina(n5259), .dinb(n278), .dout(n5260));
  jxor g05005(.dina(n5260), .dinb(n5245), .dout(n5261));
  jxor g05006(.dina(n5261), .dinb(n5053), .dout(f43 ));
  jnot g05007(.din(n5260), .dout(n5263));
  jor  g05008(.dina(n5263), .dinb(n5245), .dout(n5264));
  jor  g05009(.dina(n5261), .dinb(n5053), .dout(n5265));
  jand g05010(.dina(n5265), .dinb(n5264), .dout(n5266));
  jand g05011(.dina(n5243), .dinb(n5235), .dout(n5267));
  jnot g05012(.din(n5267), .dout(n5268));
  jnot g05013(.din(n5244), .dout(n5269));
  jor  g05014(.dina(n5269), .dinb(n5058), .dout(n5270));
  jand g05015(.dina(n5270), .dinb(n5268), .dout(n5271));
  jand g05016(.dina(n5233), .dinb(n5225), .dout(n5272));
  jand g05017(.dina(n5234), .dinb(n5061), .dout(n5273));
  jor  g05018(.dina(n5273), .dinb(n5272), .dout(n5274));
  jand g05019(.dina(n5222), .dinb(n5214), .dout(n5275));
  jnot g05020(.din(n5275), .dout(n5276));
  jor  g05021(.dina(n5224), .dinb(n5065), .dout(n5277));
  jand g05022(.dina(n5277), .dinb(n5276), .dout(n5278));
  jand g05023(.dina(n5212), .dinb(n5204), .dout(n5279));
  jand g05024(.dina(n5213), .dinb(n5068), .dout(n5280));
  jor  g05025(.dina(n5280), .dinb(n5279), .dout(n5281));
  jand g05026(.dina(n5202), .dinb(n5194), .dout(n5282));
  jand g05027(.dina(n5203), .dinb(n5071), .dout(n5283));
  jor  g05028(.dina(n5283), .dinb(n5282), .dout(n5284));
  jand g05029(.dina(n5192), .dinb(n5184), .dout(n5285));
  jand g05030(.dina(n5193), .dinb(n5074), .dout(n5286));
  jor  g05031(.dina(n5286), .dinb(n5285), .dout(n5287));
  jand g05032(.dina(n5182), .dinb(n5174), .dout(n5288));
  jand g05033(.dina(n5183), .dinb(n5077), .dout(n5289));
  jor  g05034(.dina(n5289), .dinb(n5288), .dout(n5290));
  jand g05035(.dina(n5172), .dinb(n5164), .dout(n5291));
  jand g05036(.dina(n5173), .dinb(n5080), .dout(n5292));
  jor  g05037(.dina(n5292), .dinb(n5291), .dout(n5293));
  jand g05038(.dina(n5162), .dinb(n5154), .dout(n5294));
  jand g05039(.dina(n5163), .dinb(n5083), .dout(n5295));
  jor  g05040(.dina(n5295), .dinb(n5294), .dout(n5296));
  jand g05041(.dina(n5152), .dinb(n5144), .dout(n5297));
  jand g05042(.dina(n5153), .dinb(n5086), .dout(n5298));
  jor  g05043(.dina(n5298), .dinb(n5297), .dout(n5299));
  jand g05044(.dina(n5142), .dinb(n5134), .dout(n5300));
  jand g05045(.dina(n5143), .dinb(n5089), .dout(n5301));
  jor  g05046(.dina(n5301), .dinb(n5300), .dout(n5302));
  jor  g05047(.dina(n5132), .dinb(n5124), .dout(n5303));
  jand g05048(.dina(n5133), .dinb(n5094), .dout(n5304));
  jnot g05049(.din(n5304), .dout(n5305));
  jand g05050(.dina(n5305), .dinb(n5303), .dout(n5306));
  jnot g05051(.din(n5306), .dout(n5307));
  jor  g05052(.dina(n5121), .dinb(n5113), .dout(n5308));
  jand g05053(.dina(n5122), .dinb(n5098), .dout(n5309));
  jnot g05054(.din(n5309), .dout(n5310));
  jand g05055(.dina(n5310), .dinb(n5308), .dout(n5311));
  jnot g05056(.din(n5311), .dout(n5312));
  jand g05057(.dina(n5104), .dinb(b1 ), .dout(n5313));
  jor  g05058(.dina(n5103), .dinb(n4895), .dout(n5314));
  jor  g05059(.dina(n5314), .dinb(n5106), .dout(n5315));
  jnot g05060(.din(n5315), .dout(n5316));
  jand g05061(.dina(n5316), .dinb(b0 ), .dout(n5317));
  jand g05062(.dina(n5100), .dinb(n273), .dout(n5318));
  jand g05063(.dina(n5107), .dinb(b2 ), .dout(n5319));
  jor  g05064(.dina(n5319), .dinb(n5318), .dout(n5320));
  jor  g05065(.dina(n5320), .dinb(n5317), .dout(n5321));
  jor  g05066(.dina(n5321), .dinb(n5313), .dout(n5322));
  jnot g05067(.din(n5110), .dout(n5323));
  jand g05068(.dina(n4897), .dinb(a44 ), .dout(n5324));
  jand g05069(.dina(n5324), .dinb(n5323), .dout(n5325));
  jnot g05070(.din(n5325), .dout(n5326));
  jand g05071(.dina(n5326), .dinb(a44 ), .dout(n5327));
  jxor g05072(.dina(n5327), .dinb(n5322), .dout(n5328));
  jnot g05073(.din(n5328), .dout(n5329));
  jor  g05074(.dina(n4902), .dinb(n374), .dout(n5330));
  jor  g05075(.dina(n4904), .dinb(n340), .dout(n5331));
  jor  g05076(.dina(n4696), .dinb(n303), .dout(n5332));
  jand g05077(.dina(n5332), .dinb(n5331), .dout(n5333));
  jor  g05078(.dina(n4899), .dinb(n377), .dout(n5334));
  jand g05079(.dina(n5334), .dinb(n5333), .dout(n5335));
  jand g05080(.dina(n5335), .dinb(n5330), .dout(n5336));
  jxor g05081(.dina(n5336), .dinb(a41 ), .dout(n5337));
  jxor g05082(.dina(n5337), .dinb(n5329), .dout(n5338));
  jxor g05083(.dina(n5338), .dinb(n5312), .dout(n5339));
  jnot g05084(.din(n5339), .dout(n5340));
  jor  g05085(.dina(n4305), .dinb(n517), .dout(n5341));
  jor  g05086(.dina(n4303), .dinb(n519), .dout(n5342));
  jor  g05087(.dina(n4308), .dinb(n469), .dout(n5343));
  jor  g05088(.dina(n4116), .dinb(n415), .dout(n5344));
  jand g05089(.dina(n5344), .dinb(n5343), .dout(n5345));
  jand g05090(.dina(n5345), .dinb(n5342), .dout(n5346));
  jand g05091(.dina(n5346), .dinb(n5341), .dout(n5347));
  jxor g05092(.dina(n5347), .dinb(a38 ), .dout(n5348));
  jxor g05093(.dina(n5348), .dinb(n5340), .dout(n5349));
  jxor g05094(.dina(n5349), .dinb(n5307), .dout(n5350));
  jor  g05095(.dina(n3751), .dinb(n702), .dout(n5351));
  jor  g05096(.dina(n3574), .dinb(n572), .dout(n5352));
  jor  g05097(.dina(n3749), .dinb(n704), .dout(n5353));
  jor  g05098(.dina(n3754), .dinb(n637), .dout(n5354));
  jand g05099(.dina(n5354), .dinb(n5353), .dout(n5355));
  jand g05100(.dina(n5355), .dinb(n5352), .dout(n5356));
  jand g05101(.dina(n5356), .dinb(n5351), .dout(n5357));
  jxor g05102(.dina(n5357), .dinb(n3410), .dout(n5358));
  jxor g05103(.dina(n5358), .dinb(n5350), .dout(n5359));
  jxor g05104(.dina(n5359), .dinb(n5302), .dout(n5360));
  jor  g05105(.dina(n3239), .dinb(n932), .dout(n5361));
  jor  g05106(.dina(n3072), .dinb(n772), .dout(n5362));
  jor  g05107(.dina(n3237), .dinb(n934), .dout(n5363));
  jor  g05108(.dina(n3242), .dinb(n852), .dout(n5364));
  jand g05109(.dina(n5364), .dinb(n5363), .dout(n5365));
  jand g05110(.dina(n5365), .dinb(n5362), .dout(n5366));
  jand g05111(.dina(n5366), .dinb(n5361), .dout(n5367));
  jxor g05112(.dina(n5367), .dinb(n2918), .dout(n5368));
  jxor g05113(.dina(n5368), .dinb(n5360), .dout(n5369));
  jxor g05114(.dina(n5369), .dinb(n5299), .dout(n5370));
  jor  g05115(.dina(n2764), .dinb(n1209), .dout(n5371));
  jor  g05116(.dina(n2609), .dinb(n1018), .dout(n5372));
  jor  g05117(.dina(n2761), .dinb(n1211), .dout(n5373));
  jor  g05118(.dina(n2766), .dinb(n1114), .dout(n5374));
  jand g05119(.dina(n5374), .dinb(n5373), .dout(n5375));
  jand g05120(.dina(n5375), .dinb(n5372), .dout(n5376));
  jand g05121(.dina(n5376), .dinb(n5371), .dout(n5377));
  jxor g05122(.dina(n5377), .dinb(n2468), .dout(n5378));
  jxor g05123(.dina(n5378), .dinb(n5370), .dout(n5379));
  jxor g05124(.dina(n5379), .dinb(n5296), .dout(n5380));
  jor  g05125(.dina(n2324), .dinb(n1525), .dout(n5381));
  jor  g05126(.dina(n2186), .dinb(n1307), .dout(n5382));
  jor  g05127(.dina(n2326), .dinb(n1527), .dout(n5383));
  jor  g05128(.dina(n2321), .dinb(n1416), .dout(n5384));
  jand g05129(.dina(n5384), .dinb(n5383), .dout(n5385));
  jand g05130(.dina(n5385), .dinb(n5382), .dout(n5386));
  jand g05131(.dina(n5386), .dinb(n5381), .dout(n5387));
  jxor g05132(.dina(n5387), .dinb(n2057), .dout(n5388));
  jxor g05133(.dina(n5388), .dinb(n5380), .dout(n5389));
  jxor g05134(.dina(n5389), .dinb(n5293), .dout(n5390));
  jor  g05135(.dina(n1879), .dinb(n1921), .dout(n5391));
  jor  g05136(.dina(n1806), .dinb(n1637), .dout(n5392));
  jor  g05137(.dina(n1923), .dinb(n1881), .dout(n5393));
  jor  g05138(.dina(n1918), .dinb(n1759), .dout(n5394));
  jand g05139(.dina(n5394), .dinb(n5393), .dout(n5395));
  jand g05140(.dina(n5395), .dinb(n5392), .dout(n5396));
  jand g05141(.dina(n5396), .dinb(n5391), .dout(n5397));
  jxor g05142(.dina(n5397), .dinb(n1687), .dout(n5398));
  jxor g05143(.dina(n5398), .dinb(n5390), .dout(n5399));
  jxor g05144(.dina(n5399), .dinb(n5290), .dout(n5400));
  jor  g05145(.dina(n2277), .dinb(n1569), .dout(n5401));
  jor  g05146(.dina(n1453), .dinb(n2007), .dout(n5402));
  jor  g05147(.dina(n1566), .dinb(n2142), .dout(n5403));
  jor  g05148(.dina(n1571), .dinb(n2279), .dout(n5404));
  jand g05149(.dina(n5404), .dinb(n5403), .dout(n5405));
  jand g05150(.dina(n5405), .dinb(n5402), .dout(n5406));
  jand g05151(.dina(n5406), .dinb(n5401), .dout(n5407));
  jxor g05152(.dina(n5407), .dinb(n1351), .dout(n5408));
  jxor g05153(.dina(n5408), .dinb(n5400), .dout(n5409));
  jxor g05154(.dina(n5409), .dinb(n5287), .dout(n5410));
  jor  g05155(.dina(n2711), .dinb(n1248), .dout(n5411));
  jor  g05156(.dina(n1147), .dinb(n2415), .dout(n5412));
  jor  g05157(.dina(n1251), .dinb(n2563), .dout(n5413));
  jor  g05158(.dina(n1246), .dinb(n2713), .dout(n5414));
  jand g05159(.dina(n5414), .dinb(n5413), .dout(n5415));
  jand g05160(.dina(n5415), .dinb(n5412), .dout(n5416));
  jand g05161(.dina(n5416), .dinb(n5411), .dout(n5417));
  jxor g05162(.dina(n5417), .dinb(n1061), .dout(n5418));
  jxor g05163(.dina(n5418), .dinb(n5410), .dout(n5419));
  jxor g05164(.dina(n5419), .dinb(n5284), .dout(n5420));
  jor  g05165(.dina(n3184), .dinb(n970), .dout(n5421));
  jor  g05166(.dina(n880), .dinb(n2862), .dout(n5422));
  jor  g05167(.dina(n967), .dinb(n3023), .dout(n5423));
  jor  g05168(.dina(n972), .dinb(n3186), .dout(n5424));
  jand g05169(.dina(n5424), .dinb(n5423), .dout(n5425));
  jand g05170(.dina(n5425), .dinb(n5422), .dout(n5426));
  jand g05171(.dina(n5426), .dinb(n5421), .dout(n5427));
  jxor g05172(.dina(n5427), .dinb(n810), .dout(n5428));
  jxor g05173(.dina(n5428), .dinb(n5420), .dout(n5429));
  jxor g05174(.dina(n5429), .dinb(n5281), .dout(n5430));
  jor  g05175(.dina(n3696), .dinb(n728), .dout(n5431));
  jor  g05176(.dina(n660), .dinb(n3348), .dout(n5432));
  jor  g05177(.dina(n726), .dinb(n3698), .dout(n5433));
  jor  g05178(.dina(n731), .dinb(n3522), .dout(n5434));
  jand g05179(.dina(n5434), .dinb(n5433), .dout(n5435));
  jand g05180(.dina(n5435), .dinb(n5432), .dout(n5436));
  jand g05181(.dina(n5436), .dinb(n5431), .dout(n5437));
  jxor g05182(.dina(n5437), .dinb(n606), .dout(n5438));
  jxor g05183(.dina(n5438), .dinb(n5430), .dout(n5439));
  jnot g05184(.din(n5439), .dout(n5440));
  jxor g05185(.dina(n5440), .dinb(n5278), .dout(n5441));
  jor  g05186(.dina(n4247), .dinb(n544), .dout(n5442));
  jor  g05187(.dina(n486), .dinb(n3873), .dout(n5443));
  jor  g05188(.dina(n547), .dinb(n4060), .dout(n5444));
  jor  g05189(.dina(n542), .dinb(n4249), .dout(n5445));
  jand g05190(.dina(n5445), .dinb(n5444), .dout(n5446));
  jand g05191(.dina(n5446), .dinb(n5443), .dout(n5447));
  jand g05192(.dina(n5447), .dinb(n5442), .dout(n5448));
  jxor g05193(.dina(n5448), .dinb(n446), .dout(n5449));
  jxor g05194(.dina(n5449), .dinb(n5441), .dout(n5450));
  jxor g05195(.dina(n5450), .dinb(n5274), .dout(n5451));
  jor  g05196(.dina(n4837), .dinb(n397), .dout(n5452));
  jor  g05197(.dina(n354), .dinb(n4437), .dout(n5453));
  jor  g05198(.dina(n394), .dinb(n4637), .dout(n5454));
  jor  g05199(.dina(n399), .dinb(n4839), .dout(n5455));
  jand g05200(.dina(n5455), .dinb(n5454), .dout(n5456));
  jand g05201(.dina(n5456), .dinb(n5453), .dout(n5457));
  jand g05202(.dina(n5457), .dinb(n5452), .dout(n5458));
  jxor g05203(.dina(n5458), .dinb(n364), .dout(n5459));
  jxor g05204(.dina(n5459), .dinb(n5451), .dout(n5460));
  jxor g05205(.dina(n5460), .dinb(n5271), .dout(n5461));
  jand g05206(.dina(b43 ), .dinb(b42 ), .dout(n5462));
  jand g05207(.dina(n5249), .dinb(n5248), .dout(n5463));
  jor  g05208(.dina(n5463), .dinb(n5462), .dout(n5464));
  jxor g05209(.dina(b44 ), .dinb(b43 ), .dout(n5465));
  jnot g05210(.din(n5465), .dout(n5466));
  jxor g05211(.dina(n5466), .dinb(n5464), .dout(n5467));
  jor  g05212(.dina(n5467), .dinb(n296), .dout(n5468));
  jnot g05213(.din(b44 ), .dout(n5469));
  jor  g05214(.dina(n264), .dinb(n5469), .dout(n5470));
  jor  g05215(.dina(n294), .dinb(n5253), .dout(n5471));
  jor  g05216(.dina(n280), .dinb(n5040), .dout(n5472));
  jand g05217(.dina(n5472), .dinb(n5471), .dout(n5473));
  jand g05218(.dina(n5473), .dinb(n5470), .dout(n5474));
  jand g05219(.dina(n5474), .dinb(n5468), .dout(n5475));
  jxor g05220(.dina(n5475), .dinb(n278), .dout(n5476));
  jxor g05221(.dina(n5476), .dinb(n5461), .dout(n5477));
  jxor g05222(.dina(n5477), .dinb(n5266), .dout(f44 ));
  jnot g05223(.din(n5476), .dout(n5479));
  jor  g05224(.dina(n5479), .dinb(n5461), .dout(n5480));
  jor  g05225(.dina(n5477), .dinb(n5266), .dout(n5481));
  jand g05226(.dina(n5481), .dinb(n5480), .dout(n5482));
  jand g05227(.dina(n5459), .dinb(n5451), .dout(n5483));
  jnot g05228(.din(n5483), .dout(n5484));
  jnot g05229(.din(n5460), .dout(n5485));
  jor  g05230(.dina(n5485), .dinb(n5271), .dout(n5486));
  jand g05231(.dina(n5486), .dinb(n5484), .dout(n5487));
  jand g05232(.dina(n5449), .dinb(n5441), .dout(n5488));
  jand g05233(.dina(n5450), .dinb(n5274), .dout(n5489));
  jor  g05234(.dina(n5489), .dinb(n5488), .dout(n5490));
  jand g05235(.dina(n5438), .dinb(n5430), .dout(n5491));
  jnot g05236(.din(n5491), .dout(n5492));
  jor  g05237(.dina(n5440), .dinb(n5278), .dout(n5493));
  jand g05238(.dina(n5493), .dinb(n5492), .dout(n5494));
  jand g05239(.dina(n5428), .dinb(n5420), .dout(n5495));
  jand g05240(.dina(n5429), .dinb(n5281), .dout(n5496));
  jor  g05241(.dina(n5496), .dinb(n5495), .dout(n5497));
  jand g05242(.dina(n5418), .dinb(n5410), .dout(n5498));
  jand g05243(.dina(n5419), .dinb(n5284), .dout(n5499));
  jor  g05244(.dina(n5499), .dinb(n5498), .dout(n5500));
  jand g05245(.dina(n5408), .dinb(n5400), .dout(n5501));
  jand g05246(.dina(n5409), .dinb(n5287), .dout(n5502));
  jor  g05247(.dina(n5502), .dinb(n5501), .dout(n5503));
  jand g05248(.dina(n5398), .dinb(n5390), .dout(n5504));
  jand g05249(.dina(n5399), .dinb(n5290), .dout(n5505));
  jor  g05250(.dina(n5505), .dinb(n5504), .dout(n5506));
  jand g05251(.dina(n5388), .dinb(n5380), .dout(n5507));
  jand g05252(.dina(n5389), .dinb(n5293), .dout(n5508));
  jor  g05253(.dina(n5508), .dinb(n5507), .dout(n5509));
  jand g05254(.dina(n5378), .dinb(n5370), .dout(n5510));
  jand g05255(.dina(n5379), .dinb(n5296), .dout(n5511));
  jor  g05256(.dina(n5511), .dinb(n5510), .dout(n5512));
  jand g05257(.dina(n5368), .dinb(n5360), .dout(n5513));
  jand g05258(.dina(n5369), .dinb(n5299), .dout(n5514));
  jor  g05259(.dina(n5514), .dinb(n5513), .dout(n5515));
  jand g05260(.dina(n5358), .dinb(n5350), .dout(n5516));
  jand g05261(.dina(n5359), .dinb(n5302), .dout(n5517));
  jor  g05262(.dina(n5517), .dinb(n5516), .dout(n5518));
  jor  g05263(.dina(n5348), .dinb(n5340), .dout(n5519));
  jand g05264(.dina(n5349), .dinb(n5307), .dout(n5520));
  jnot g05265(.din(n5520), .dout(n5521));
  jand g05266(.dina(n5521), .dinb(n5519), .dout(n5522));
  jnot g05267(.din(n5522), .dout(n5523));
  jor  g05268(.dina(n5337), .dinb(n5329), .dout(n5524));
  jand g05269(.dina(n5338), .dinb(n5312), .dout(n5525));
  jnot g05270(.din(n5525), .dout(n5526));
  jand g05271(.dina(n5526), .dinb(n5524), .dout(n5527));
  jnot g05272(.din(n5527), .dout(n5528));
  jor  g05273(.dina(n5326), .dinb(n5322), .dout(n5529));
  jxor g05274(.dina(a45 ), .dinb(a44 ), .dout(n5530));
  jand g05275(.dina(n5530), .dinb(b0 ), .dout(n5531));
  jnot g05276(.din(n5531), .dout(n5532));
  jxor g05277(.dina(n5532), .dinb(n5529), .dout(n5533));
  jnot g05278(.din(n5104), .dout(n5534));
  jor  g05279(.dina(n5534), .dinb(n293), .dout(n5535));
  jor  g05280(.dina(n5315), .dinb(n305), .dout(n5536));
  jnot g05281(.din(n5100), .dout(n5537));
  jor  g05282(.dina(n5537), .dinb(n301), .dout(n5538));
  jnot g05283(.din(n5107), .dout(n5539));
  jor  g05284(.dina(n5539), .dinb(n303), .dout(n5540));
  jand g05285(.dina(n5540), .dinb(n5538), .dout(n5541));
  jand g05286(.dina(n5541), .dinb(n5536), .dout(n5542));
  jand g05287(.dina(n5542), .dinb(n5535), .dout(n5543));
  jxor g05288(.dina(n5543), .dinb(n5111), .dout(n5544));
  jxor g05289(.dina(n5544), .dinb(n5533), .dout(n5545));
  jnot g05290(.din(n5545), .dout(n5546));
  jor  g05291(.dina(n4902), .dinb(n412), .dout(n5547));
  jor  g05292(.dina(n4899), .dinb(n415), .dout(n5548));
  jor  g05293(.dina(n4696), .dinb(n340), .dout(n5549));
  jand g05294(.dina(n5549), .dinb(n5548), .dout(n5550));
  jor  g05295(.dina(n4904), .dinb(n377), .dout(n5551));
  jand g05296(.dina(n5551), .dinb(n5550), .dout(n5552));
  jand g05297(.dina(n5552), .dinb(n5547), .dout(n5553));
  jxor g05298(.dina(n5553), .dinb(a41 ), .dout(n5554));
  jxor g05299(.dina(n5554), .dinb(n5546), .dout(n5555));
  jxor g05300(.dina(n5555), .dinb(n5528), .dout(n5556));
  jor  g05301(.dina(n4305), .dinb(n570), .dout(n5557));
  jor  g05302(.dina(n4116), .dinb(n469), .dout(n5558));
  jor  g05303(.dina(n4308), .dinb(n519), .dout(n5559));
  jor  g05304(.dina(n4303), .dinb(n572), .dout(n5560));
  jand g05305(.dina(n5560), .dinb(n5559), .dout(n5561));
  jand g05306(.dina(n5561), .dinb(n5558), .dout(n5562));
  jand g05307(.dina(n5562), .dinb(n5557), .dout(n5563));
  jxor g05308(.dina(n5563), .dinb(n3938), .dout(n5564));
  jxor g05309(.dina(n5564), .dinb(n5556), .dout(n5565));
  jxor g05310(.dina(n5565), .dinb(n5523), .dout(n5566));
  jor  g05311(.dina(n3751), .dinb(n770), .dout(n5567));
  jor  g05312(.dina(n3574), .dinb(n637), .dout(n5568));
  jor  g05313(.dina(n3749), .dinb(n772), .dout(n5569));
  jor  g05314(.dina(n3754), .dinb(n704), .dout(n5570));
  jand g05315(.dina(n5570), .dinb(n5569), .dout(n5571));
  jand g05316(.dina(n5571), .dinb(n5568), .dout(n5572));
  jand g05317(.dina(n5572), .dinb(n5567), .dout(n5573));
  jxor g05318(.dina(n5573), .dinb(n3410), .dout(n5574));
  jxor g05319(.dina(n5574), .dinb(n5566), .dout(n5575));
  jxor g05320(.dina(n5575), .dinb(n5518), .dout(n5576));
  jor  g05321(.dina(n3239), .dinb(n1016), .dout(n5577));
  jor  g05322(.dina(n3072), .dinb(n852), .dout(n5578));
  jor  g05323(.dina(n3237), .dinb(n1018), .dout(n5579));
  jor  g05324(.dina(n3242), .dinb(n934), .dout(n5580));
  jand g05325(.dina(n5580), .dinb(n5579), .dout(n5581));
  jand g05326(.dina(n5581), .dinb(n5578), .dout(n5582));
  jand g05327(.dina(n5582), .dinb(n5577), .dout(n5583));
  jxor g05328(.dina(n5583), .dinb(n2918), .dout(n5584));
  jxor g05329(.dina(n5584), .dinb(n5576), .dout(n5585));
  jxor g05330(.dina(n5585), .dinb(n5515), .dout(n5586));
  jor  g05331(.dina(n2764), .dinb(n1305), .dout(n5587));
  jor  g05332(.dina(n2609), .dinb(n1114), .dout(n5588));
  jor  g05333(.dina(n2761), .dinb(n1307), .dout(n5589));
  jor  g05334(.dina(n2766), .dinb(n1211), .dout(n5590));
  jand g05335(.dina(n5590), .dinb(n5589), .dout(n5591));
  jand g05336(.dina(n5591), .dinb(n5588), .dout(n5592));
  jand g05337(.dina(n5592), .dinb(n5587), .dout(n5593));
  jxor g05338(.dina(n5593), .dinb(n2468), .dout(n5594));
  jxor g05339(.dina(n5594), .dinb(n5586), .dout(n5595));
  jxor g05340(.dina(n5595), .dinb(n5512), .dout(n5596));
  jor  g05341(.dina(n2324), .dinb(n1635), .dout(n5597));
  jor  g05342(.dina(n2186), .dinb(n1416), .dout(n5598));
  jor  g05343(.dina(n2326), .dinb(n1637), .dout(n5599));
  jor  g05344(.dina(n2321), .dinb(n1527), .dout(n5600));
  jand g05345(.dina(n5600), .dinb(n5599), .dout(n5601));
  jand g05346(.dina(n5601), .dinb(n5598), .dout(n5602));
  jand g05347(.dina(n5602), .dinb(n5597), .dout(n5603));
  jxor g05348(.dina(n5603), .dinb(n2057), .dout(n5604));
  jxor g05349(.dina(n5604), .dinb(n5596), .dout(n5605));
  jxor g05350(.dina(n5605), .dinb(n5509), .dout(n5606));
  jor  g05351(.dina(n2005), .dinb(n1921), .dout(n5607));
  jor  g05352(.dina(n1806), .dinb(n1759), .dout(n5608));
  jor  g05353(.dina(n1923), .dinb(n2007), .dout(n5609));
  jor  g05354(.dina(n1918), .dinb(n1881), .dout(n5610));
  jand g05355(.dina(n5610), .dinb(n5609), .dout(n5611));
  jand g05356(.dina(n5611), .dinb(n5608), .dout(n5612));
  jand g05357(.dina(n5612), .dinb(n5607), .dout(n5613));
  jxor g05358(.dina(n5613), .dinb(n1687), .dout(n5614));
  jxor g05359(.dina(n5614), .dinb(n5606), .dout(n5615));
  jxor g05360(.dina(n5615), .dinb(n5506), .dout(n5616));
  jor  g05361(.dina(n2413), .dinb(n1569), .dout(n5617));
  jor  g05362(.dina(n1453), .dinb(n2142), .dout(n5618));
  jor  g05363(.dina(n1566), .dinb(n2279), .dout(n5619));
  jor  g05364(.dina(n1571), .dinb(n2415), .dout(n5620));
  jand g05365(.dina(n5620), .dinb(n5619), .dout(n5621));
  jand g05366(.dina(n5621), .dinb(n5618), .dout(n5622));
  jand g05367(.dina(n5622), .dinb(n5617), .dout(n5623));
  jxor g05368(.dina(n5623), .dinb(n1351), .dout(n5624));
  jxor g05369(.dina(n5624), .dinb(n5616), .dout(n5625));
  jxor g05370(.dina(n5625), .dinb(n5503), .dout(n5626));
  jor  g05371(.dina(n2860), .dinb(n1248), .dout(n5627));
  jor  g05372(.dina(n1147), .dinb(n2563), .dout(n5628));
  jor  g05373(.dina(n1246), .dinb(n2862), .dout(n5629));
  jor  g05374(.dina(n1251), .dinb(n2713), .dout(n5630));
  jand g05375(.dina(n5630), .dinb(n5629), .dout(n5631));
  jand g05376(.dina(n5631), .dinb(n5628), .dout(n5632));
  jand g05377(.dina(n5632), .dinb(n5627), .dout(n5633));
  jxor g05378(.dina(n5633), .dinb(n1061), .dout(n5634));
  jxor g05379(.dina(n5634), .dinb(n5626), .dout(n5635));
  jxor g05380(.dina(n5635), .dinb(n5500), .dout(n5636));
  jor  g05381(.dina(n3346), .dinb(n970), .dout(n5637));
  jor  g05382(.dina(n880), .dinb(n3023), .dout(n5638));
  jor  g05383(.dina(n967), .dinb(n3186), .dout(n5639));
  jor  g05384(.dina(n972), .dinb(n3348), .dout(n5640));
  jand g05385(.dina(n5640), .dinb(n5639), .dout(n5641));
  jand g05386(.dina(n5641), .dinb(n5638), .dout(n5642));
  jand g05387(.dina(n5642), .dinb(n5637), .dout(n5643));
  jxor g05388(.dina(n5643), .dinb(n810), .dout(n5644));
  jxor g05389(.dina(n5644), .dinb(n5636), .dout(n5645));
  jxor g05390(.dina(n5645), .dinb(n5497), .dout(n5646));
  jor  g05391(.dina(n3871), .dinb(n728), .dout(n5647));
  jor  g05392(.dina(n660), .dinb(n3522), .dout(n5648));
  jor  g05393(.dina(n726), .dinb(n3873), .dout(n5649));
  jor  g05394(.dina(n731), .dinb(n3698), .dout(n5650));
  jand g05395(.dina(n5650), .dinb(n5649), .dout(n5651));
  jand g05396(.dina(n5651), .dinb(n5648), .dout(n5652));
  jand g05397(.dina(n5652), .dinb(n5647), .dout(n5653));
  jxor g05398(.dina(n5653), .dinb(n606), .dout(n5654));
  jxor g05399(.dina(n5654), .dinb(n5646), .dout(n5655));
  jnot g05400(.din(n5655), .dout(n5656));
  jxor g05401(.dina(n5656), .dinb(n5494), .dout(n5657));
  jor  g05402(.dina(n4435), .dinb(n544), .dout(n5658));
  jor  g05403(.dina(n486), .dinb(n4060), .dout(n5659));
  jor  g05404(.dina(n547), .dinb(n4249), .dout(n5660));
  jor  g05405(.dina(n542), .dinb(n4437), .dout(n5661));
  jand g05406(.dina(n5661), .dinb(n5660), .dout(n5662));
  jand g05407(.dina(n5662), .dinb(n5659), .dout(n5663));
  jand g05408(.dina(n5663), .dinb(n5658), .dout(n5664));
  jxor g05409(.dina(n5664), .dinb(n446), .dout(n5665));
  jxor g05410(.dina(n5665), .dinb(n5657), .dout(n5666));
  jxor g05411(.dina(n5666), .dinb(n5490), .dout(n5667));
  jor  g05412(.dina(n5038), .dinb(n397), .dout(n5668));
  jor  g05413(.dina(n354), .dinb(n4637), .dout(n5669));
  jor  g05414(.dina(n394), .dinb(n4839), .dout(n5670));
  jor  g05415(.dina(n399), .dinb(n5040), .dout(n5671));
  jand g05416(.dina(n5671), .dinb(n5670), .dout(n5672));
  jand g05417(.dina(n5672), .dinb(n5669), .dout(n5673));
  jand g05418(.dina(n5673), .dinb(n5668), .dout(n5674));
  jxor g05419(.dina(n5674), .dinb(n364), .dout(n5675));
  jxor g05420(.dina(n5675), .dinb(n5667), .dout(n5676));
  jxor g05421(.dina(n5676), .dinb(n5487), .dout(n5677));
  jand g05422(.dina(b44 ), .dinb(b43 ), .dout(n5678));
  jand g05423(.dina(n5465), .dinb(n5464), .dout(n5679));
  jor  g05424(.dina(n5679), .dinb(n5678), .dout(n5680));
  jxor g05425(.dina(b45 ), .dinb(b44 ), .dout(n5681));
  jnot g05426(.din(n5681), .dout(n5682));
  jxor g05427(.dina(n5682), .dinb(n5680), .dout(n5683));
  jor  g05428(.dina(n5683), .dinb(n296), .dout(n5684));
  jnot g05429(.din(b45 ), .dout(n5685));
  jor  g05430(.dina(n264), .dinb(n5685), .dout(n5686));
  jor  g05431(.dina(n294), .dinb(n5469), .dout(n5687));
  jor  g05432(.dina(n280), .dinb(n5253), .dout(n5688));
  jand g05433(.dina(n5688), .dinb(n5687), .dout(n5689));
  jand g05434(.dina(n5689), .dinb(n5686), .dout(n5690));
  jand g05435(.dina(n5690), .dinb(n5684), .dout(n5691));
  jxor g05436(.dina(n5691), .dinb(n278), .dout(n5692));
  jxor g05437(.dina(n5692), .dinb(n5677), .dout(n5693));
  jxor g05438(.dina(n5693), .dinb(n5482), .dout(f45 ));
  jnot g05439(.din(n5692), .dout(n5695));
  jor  g05440(.dina(n5695), .dinb(n5677), .dout(n5696));
  jor  g05441(.dina(n5693), .dinb(n5482), .dout(n5697));
  jand g05442(.dina(n5697), .dinb(n5696), .dout(n5698));
  jand g05443(.dina(n5675), .dinb(n5667), .dout(n5699));
  jnot g05444(.din(n5699), .dout(n5700));
  jnot g05445(.din(n5676), .dout(n5701));
  jor  g05446(.dina(n5701), .dinb(n5487), .dout(n5702));
  jand g05447(.dina(n5702), .dinb(n5700), .dout(n5703));
  jand g05448(.dina(n5665), .dinb(n5657), .dout(n5704));
  jand g05449(.dina(n5666), .dinb(n5490), .dout(n5705));
  jor  g05450(.dina(n5705), .dinb(n5704), .dout(n5706));
  jand g05451(.dina(n5654), .dinb(n5646), .dout(n5707));
  jnot g05452(.din(n5707), .dout(n5708));
  jor  g05453(.dina(n5656), .dinb(n5494), .dout(n5709));
  jand g05454(.dina(n5709), .dinb(n5708), .dout(n5710));
  jand g05455(.dina(n5644), .dinb(n5636), .dout(n5711));
  jand g05456(.dina(n5645), .dinb(n5497), .dout(n5712));
  jor  g05457(.dina(n5712), .dinb(n5711), .dout(n5713));
  jand g05458(.dina(n5634), .dinb(n5626), .dout(n5714));
  jand g05459(.dina(n5635), .dinb(n5500), .dout(n5715));
  jor  g05460(.dina(n5715), .dinb(n5714), .dout(n5716));
  jand g05461(.dina(n5624), .dinb(n5616), .dout(n5717));
  jand g05462(.dina(n5625), .dinb(n5503), .dout(n5718));
  jor  g05463(.dina(n5718), .dinb(n5717), .dout(n5719));
  jand g05464(.dina(n5614), .dinb(n5606), .dout(n5720));
  jand g05465(.dina(n5615), .dinb(n5506), .dout(n5721));
  jor  g05466(.dina(n5721), .dinb(n5720), .dout(n5722));
  jand g05467(.dina(n5604), .dinb(n5596), .dout(n5723));
  jand g05468(.dina(n5605), .dinb(n5509), .dout(n5724));
  jor  g05469(.dina(n5724), .dinb(n5723), .dout(n5725));
  jand g05470(.dina(n5594), .dinb(n5586), .dout(n5726));
  jand g05471(.dina(n5595), .dinb(n5512), .dout(n5727));
  jor  g05472(.dina(n5727), .dinb(n5726), .dout(n5728));
  jand g05473(.dina(n5584), .dinb(n5576), .dout(n5729));
  jand g05474(.dina(n5585), .dinb(n5515), .dout(n5730));
  jor  g05475(.dina(n5730), .dinb(n5729), .dout(n5731));
  jand g05476(.dina(n5574), .dinb(n5566), .dout(n5732));
  jand g05477(.dina(n5575), .dinb(n5518), .dout(n5733));
  jor  g05478(.dina(n5733), .dinb(n5732), .dout(n5734));
  jand g05479(.dina(n5564), .dinb(n5556), .dout(n5735));
  jand g05480(.dina(n5565), .dinb(n5523), .dout(n5736));
  jor  g05481(.dina(n5736), .dinb(n5735), .dout(n5737));
  jor  g05482(.dina(n5554), .dinb(n5546), .dout(n5738));
  jand g05483(.dina(n5555), .dinb(n5528), .dout(n5739));
  jnot g05484(.din(n5739), .dout(n5740));
  jand g05485(.dina(n5740), .dinb(n5738), .dout(n5741));
  jnot g05486(.din(n5741), .dout(n5742));
  jnot g05487(.din(n5529), .dout(n5743));
  jand g05488(.dina(n5531), .dinb(n5743), .dout(n5744));
  jand g05489(.dina(n5544), .dinb(n5533), .dout(n5745));
  jor  g05490(.dina(n5745), .dinb(n5744), .dout(n5746));
  jxor g05491(.dina(a47 ), .dinb(a46 ), .dout(n5747));
  jand g05492(.dina(n5747), .dinb(n5530), .dout(n5748));
  jand g05493(.dina(n5748), .dinb(n259), .dout(n5749));
  jnot g05494(.din(n5530), .dout(n5750));
  jxor g05495(.dina(a46 ), .dinb(a45 ), .dout(n5751));
  jand g05496(.dina(n5751), .dinb(n5750), .dout(n5752));
  jand g05497(.dina(n5752), .dinb(b0 ), .dout(n5753));
  jnot g05498(.din(n5747), .dout(n5754));
  jand g05499(.dina(n5754), .dinb(n5530), .dout(n5755));
  jand g05500(.dina(n5755), .dinb(b1 ), .dout(n5756));
  jor  g05501(.dina(n5756), .dinb(n5753), .dout(n5757));
  jor  g05502(.dina(n5757), .dinb(n5749), .dout(n5758));
  jnot g05503(.din(a47 ), .dout(n5759));
  jor  g05504(.dina(n5532), .dinb(n5759), .dout(n5760));
  jxor g05505(.dina(n5760), .dinb(n5758), .dout(n5761));
  jor  g05506(.dina(n5537), .dinb(n337), .dout(n5762));
  jor  g05507(.dina(n5539), .dinb(n340), .dout(n5763));
  jor  g05508(.dina(n5315), .dinb(n293), .dout(n5764));
  jand g05509(.dina(n5764), .dinb(n5763), .dout(n5765));
  jor  g05510(.dina(n5534), .dinb(n303), .dout(n5766));
  jand g05511(.dina(n5766), .dinb(n5765), .dout(n5767));
  jand g05512(.dina(n5767), .dinb(n5762), .dout(n5768));
  jxor g05513(.dina(n5768), .dinb(a44 ), .dout(n5769));
  jxor g05514(.dina(n5769), .dinb(n5761), .dout(n5770));
  jxor g05515(.dina(n5770), .dinb(n5746), .dout(n5771));
  jnot g05516(.din(n5771), .dout(n5772));
  jor  g05517(.dina(n4902), .dinb(n466), .dout(n5773));
  jor  g05518(.dina(n4899), .dinb(n469), .dout(n5774));
  jor  g05519(.dina(n4696), .dinb(n377), .dout(n5775));
  jand g05520(.dina(n5775), .dinb(n5774), .dout(n5776));
  jor  g05521(.dina(n4904), .dinb(n415), .dout(n5777));
  jand g05522(.dina(n5777), .dinb(n5776), .dout(n5778));
  jand g05523(.dina(n5778), .dinb(n5773), .dout(n5779));
  jxor g05524(.dina(n5779), .dinb(a41 ), .dout(n5780));
  jxor g05525(.dina(n5780), .dinb(n5772), .dout(n5781));
  jxor g05526(.dina(n5781), .dinb(n5742), .dout(n5782));
  jor  g05527(.dina(n4305), .dinb(n635), .dout(n5783));
  jor  g05528(.dina(n4116), .dinb(n519), .dout(n5784));
  jor  g05529(.dina(n4303), .dinb(n637), .dout(n5785));
  jor  g05530(.dina(n4308), .dinb(n572), .dout(n5786));
  jand g05531(.dina(n5786), .dinb(n5785), .dout(n5787));
  jand g05532(.dina(n5787), .dinb(n5784), .dout(n5788));
  jand g05533(.dina(n5788), .dinb(n5783), .dout(n5789));
  jxor g05534(.dina(n5789), .dinb(n3938), .dout(n5790));
  jxor g05535(.dina(n5790), .dinb(n5782), .dout(n5791));
  jxor g05536(.dina(n5791), .dinb(n5737), .dout(n5792));
  jor  g05537(.dina(n3751), .dinb(n850), .dout(n5793));
  jor  g05538(.dina(n3574), .dinb(n704), .dout(n5794));
  jor  g05539(.dina(n3749), .dinb(n852), .dout(n5795));
  jor  g05540(.dina(n3754), .dinb(n772), .dout(n5796));
  jand g05541(.dina(n5796), .dinb(n5795), .dout(n5797));
  jand g05542(.dina(n5797), .dinb(n5794), .dout(n5798));
  jand g05543(.dina(n5798), .dinb(n5793), .dout(n5799));
  jxor g05544(.dina(n5799), .dinb(n3410), .dout(n5800));
  jxor g05545(.dina(n5800), .dinb(n5792), .dout(n5801));
  jxor g05546(.dina(n5801), .dinb(n5734), .dout(n5802));
  jor  g05547(.dina(n3239), .dinb(n1112), .dout(n5803));
  jor  g05548(.dina(n3072), .dinb(n934), .dout(n5804));
  jor  g05549(.dina(n3242), .dinb(n1018), .dout(n5805));
  jor  g05550(.dina(n3237), .dinb(n1114), .dout(n5806));
  jand g05551(.dina(n5806), .dinb(n5805), .dout(n5807));
  jand g05552(.dina(n5807), .dinb(n5804), .dout(n5808));
  jand g05553(.dina(n5808), .dinb(n5803), .dout(n5809));
  jxor g05554(.dina(n5809), .dinb(n2918), .dout(n5810));
  jxor g05555(.dina(n5810), .dinb(n5802), .dout(n5811));
  jxor g05556(.dina(n5811), .dinb(n5731), .dout(n5812));
  jor  g05557(.dina(n2764), .dinb(n1414), .dout(n5813));
  jor  g05558(.dina(n2609), .dinb(n1211), .dout(n5814));
  jor  g05559(.dina(n2761), .dinb(n1416), .dout(n5815));
  jor  g05560(.dina(n2766), .dinb(n1307), .dout(n5816));
  jand g05561(.dina(n5816), .dinb(n5815), .dout(n5817));
  jand g05562(.dina(n5817), .dinb(n5814), .dout(n5818));
  jand g05563(.dina(n5818), .dinb(n5813), .dout(n5819));
  jxor g05564(.dina(n5819), .dinb(n2468), .dout(n5820));
  jxor g05565(.dina(n5820), .dinb(n5812), .dout(n5821));
  jxor g05566(.dina(n5821), .dinb(n5728), .dout(n5822));
  jor  g05567(.dina(n2324), .dinb(n1757), .dout(n5823));
  jor  g05568(.dina(n2186), .dinb(n1527), .dout(n5824));
  jor  g05569(.dina(n2326), .dinb(n1759), .dout(n5825));
  jor  g05570(.dina(n2321), .dinb(n1637), .dout(n5826));
  jand g05571(.dina(n5826), .dinb(n5825), .dout(n5827));
  jand g05572(.dina(n5827), .dinb(n5824), .dout(n5828));
  jand g05573(.dina(n5828), .dinb(n5823), .dout(n5829));
  jxor g05574(.dina(n5829), .dinb(n2057), .dout(n5830));
  jxor g05575(.dina(n5830), .dinb(n5822), .dout(n5831));
  jxor g05576(.dina(n5831), .dinb(n5725), .dout(n5832));
  jor  g05577(.dina(n2140), .dinb(n1921), .dout(n5833));
  jor  g05578(.dina(n1806), .dinb(n1881), .dout(n5834));
  jor  g05579(.dina(n1923), .dinb(n2142), .dout(n5835));
  jor  g05580(.dina(n1918), .dinb(n2007), .dout(n5836));
  jand g05581(.dina(n5836), .dinb(n5835), .dout(n5837));
  jand g05582(.dina(n5837), .dinb(n5834), .dout(n5838));
  jand g05583(.dina(n5838), .dinb(n5833), .dout(n5839));
  jxor g05584(.dina(n5839), .dinb(n1687), .dout(n5840));
  jxor g05585(.dina(n5840), .dinb(n5832), .dout(n5841));
  jxor g05586(.dina(n5841), .dinb(n5722), .dout(n5842));
  jor  g05587(.dina(n2561), .dinb(n1569), .dout(n5843));
  jor  g05588(.dina(n1453), .dinb(n2279), .dout(n5844));
  jor  g05589(.dina(n1571), .dinb(n2563), .dout(n5845));
  jor  g05590(.dina(n1566), .dinb(n2415), .dout(n5846));
  jand g05591(.dina(n5846), .dinb(n5845), .dout(n5847));
  jand g05592(.dina(n5847), .dinb(n5844), .dout(n5848));
  jand g05593(.dina(n5848), .dinb(n5843), .dout(n5849));
  jxor g05594(.dina(n5849), .dinb(n1351), .dout(n5850));
  jxor g05595(.dina(n5850), .dinb(n5842), .dout(n5851));
  jxor g05596(.dina(n5851), .dinb(n5719), .dout(n5852));
  jor  g05597(.dina(n3021), .dinb(n1248), .dout(n5853));
  jor  g05598(.dina(n1147), .dinb(n2713), .dout(n5854));
  jor  g05599(.dina(n1246), .dinb(n3023), .dout(n5855));
  jor  g05600(.dina(n1251), .dinb(n2862), .dout(n5856));
  jand g05601(.dina(n5856), .dinb(n5855), .dout(n5857));
  jand g05602(.dina(n5857), .dinb(n5854), .dout(n5858));
  jand g05603(.dina(n5858), .dinb(n5853), .dout(n5859));
  jxor g05604(.dina(n5859), .dinb(n1061), .dout(n5860));
  jxor g05605(.dina(n5860), .dinb(n5852), .dout(n5861));
  jxor g05606(.dina(n5861), .dinb(n5716), .dout(n5862));
  jor  g05607(.dina(n3520), .dinb(n970), .dout(n5863));
  jor  g05608(.dina(n880), .dinb(n3186), .dout(n5864));
  jor  g05609(.dina(n967), .dinb(n3348), .dout(n5865));
  jor  g05610(.dina(n972), .dinb(n3522), .dout(n5866));
  jand g05611(.dina(n5866), .dinb(n5865), .dout(n5867));
  jand g05612(.dina(n5867), .dinb(n5864), .dout(n5868));
  jand g05613(.dina(n5868), .dinb(n5863), .dout(n5869));
  jxor g05614(.dina(n5869), .dinb(n810), .dout(n5870));
  jxor g05615(.dina(n5870), .dinb(n5862), .dout(n5871));
  jxor g05616(.dina(n5871), .dinb(n5713), .dout(n5872));
  jor  g05617(.dina(n4058), .dinb(n728), .dout(n5873));
  jor  g05618(.dina(n660), .dinb(n3698), .dout(n5874));
  jor  g05619(.dina(n731), .dinb(n3873), .dout(n5875));
  jor  g05620(.dina(n726), .dinb(n4060), .dout(n5876));
  jand g05621(.dina(n5876), .dinb(n5875), .dout(n5877));
  jand g05622(.dina(n5877), .dinb(n5874), .dout(n5878));
  jand g05623(.dina(n5878), .dinb(n5873), .dout(n5879));
  jxor g05624(.dina(n5879), .dinb(n606), .dout(n5880));
  jxor g05625(.dina(n5880), .dinb(n5872), .dout(n5881));
  jnot g05626(.din(n5881), .dout(n5882));
  jxor g05627(.dina(n5882), .dinb(n5710), .dout(n5883));
  jor  g05628(.dina(n4635), .dinb(n544), .dout(n5884));
  jor  g05629(.dina(n486), .dinb(n4249), .dout(n5885));
  jor  g05630(.dina(n542), .dinb(n4637), .dout(n5886));
  jor  g05631(.dina(n547), .dinb(n4437), .dout(n5887));
  jand g05632(.dina(n5887), .dinb(n5886), .dout(n5888));
  jand g05633(.dina(n5888), .dinb(n5885), .dout(n5889));
  jand g05634(.dina(n5889), .dinb(n5884), .dout(n5890));
  jxor g05635(.dina(n5890), .dinb(n446), .dout(n5891));
  jxor g05636(.dina(n5891), .dinb(n5883), .dout(n5892));
  jxor g05637(.dina(n5892), .dinb(n5706), .dout(n5893));
  jor  g05638(.dina(n5251), .dinb(n397), .dout(n5894));
  jor  g05639(.dina(n354), .dinb(n4839), .dout(n5895));
  jor  g05640(.dina(n399), .dinb(n5253), .dout(n5896));
  jor  g05641(.dina(n394), .dinb(n5040), .dout(n5897));
  jand g05642(.dina(n5897), .dinb(n5896), .dout(n5898));
  jand g05643(.dina(n5898), .dinb(n5895), .dout(n5899));
  jand g05644(.dina(n5899), .dinb(n5894), .dout(n5900));
  jxor g05645(.dina(n5900), .dinb(n364), .dout(n5901));
  jxor g05646(.dina(n5901), .dinb(n5893), .dout(n5902));
  jxor g05647(.dina(n5902), .dinb(n5703), .dout(n5903));
  jand g05648(.dina(b45 ), .dinb(b44 ), .dout(n5904));
  jand g05649(.dina(n5681), .dinb(n5680), .dout(n5905));
  jor  g05650(.dina(n5905), .dinb(n5904), .dout(n5906));
  jxor g05651(.dina(b46 ), .dinb(b45 ), .dout(n5907));
  jnot g05652(.din(n5907), .dout(n5908));
  jxor g05653(.dina(n5908), .dinb(n5906), .dout(n5909));
  jor  g05654(.dina(n5909), .dinb(n296), .dout(n5910));
  jnot g05655(.din(b46 ), .dout(n5911));
  jor  g05656(.dina(n264), .dinb(n5911), .dout(n5912));
  jor  g05657(.dina(n280), .dinb(n5469), .dout(n5913));
  jor  g05658(.dina(n294), .dinb(n5685), .dout(n5914));
  jand g05659(.dina(n5914), .dinb(n5913), .dout(n5915));
  jand g05660(.dina(n5915), .dinb(n5912), .dout(n5916));
  jand g05661(.dina(n5916), .dinb(n5910), .dout(n5917));
  jxor g05662(.dina(n5917), .dinb(n278), .dout(n5918));
  jxor g05663(.dina(n5918), .dinb(n5903), .dout(n5919));
  jxor g05664(.dina(n5919), .dinb(n5698), .dout(f46 ));
  jnot g05665(.din(n5918), .dout(n5921));
  jor  g05666(.dina(n5921), .dinb(n5903), .dout(n5922));
  jor  g05667(.dina(n5919), .dinb(n5698), .dout(n5923));
  jand g05668(.dina(n5923), .dinb(n5922), .dout(n5924));
  jand g05669(.dina(n5901), .dinb(n5893), .dout(n5925));
  jnot g05670(.din(n5925), .dout(n5926));
  jnot g05671(.din(n5902), .dout(n5927));
  jor  g05672(.dina(n5927), .dinb(n5703), .dout(n5928));
  jand g05673(.dina(n5928), .dinb(n5926), .dout(n5929));
  jand g05674(.dina(n5891), .dinb(n5883), .dout(n5930));
  jand g05675(.dina(n5892), .dinb(n5706), .dout(n5931));
  jor  g05676(.dina(n5931), .dinb(n5930), .dout(n5932));
  jand g05677(.dina(n5880), .dinb(n5872), .dout(n5933));
  jnot g05678(.din(n5933), .dout(n5934));
  jor  g05679(.dina(n5882), .dinb(n5710), .dout(n5935));
  jand g05680(.dina(n5935), .dinb(n5934), .dout(n5936));
  jand g05681(.dina(n5870), .dinb(n5862), .dout(n5937));
  jand g05682(.dina(n5871), .dinb(n5713), .dout(n5938));
  jor  g05683(.dina(n5938), .dinb(n5937), .dout(n5939));
  jand g05684(.dina(n5860), .dinb(n5852), .dout(n5940));
  jand g05685(.dina(n5861), .dinb(n5716), .dout(n5941));
  jor  g05686(.dina(n5941), .dinb(n5940), .dout(n5942));
  jand g05687(.dina(n5850), .dinb(n5842), .dout(n5943));
  jand g05688(.dina(n5851), .dinb(n5719), .dout(n5944));
  jor  g05689(.dina(n5944), .dinb(n5943), .dout(n5945));
  jand g05690(.dina(n5840), .dinb(n5832), .dout(n5946));
  jand g05691(.dina(n5841), .dinb(n5722), .dout(n5947));
  jor  g05692(.dina(n5947), .dinb(n5946), .dout(n5948));
  jand g05693(.dina(n5830), .dinb(n5822), .dout(n5949));
  jand g05694(.dina(n5831), .dinb(n5725), .dout(n5950));
  jor  g05695(.dina(n5950), .dinb(n5949), .dout(n5951));
  jand g05696(.dina(n5820), .dinb(n5812), .dout(n5952));
  jand g05697(.dina(n5821), .dinb(n5728), .dout(n5953));
  jor  g05698(.dina(n5953), .dinb(n5952), .dout(n5954));
  jand g05699(.dina(n5810), .dinb(n5802), .dout(n5955));
  jand g05700(.dina(n5811), .dinb(n5731), .dout(n5956));
  jor  g05701(.dina(n5956), .dinb(n5955), .dout(n5957));
  jand g05702(.dina(n5800), .dinb(n5792), .dout(n5958));
  jand g05703(.dina(n5801), .dinb(n5734), .dout(n5959));
  jor  g05704(.dina(n5959), .dinb(n5958), .dout(n5960));
  jand g05705(.dina(n5790), .dinb(n5782), .dout(n5961));
  jand g05706(.dina(n5791), .dinb(n5737), .dout(n5962));
  jor  g05707(.dina(n5962), .dinb(n5961), .dout(n5963));
  jor  g05708(.dina(n5780), .dinb(n5772), .dout(n5964));
  jand g05709(.dina(n5781), .dinb(n5742), .dout(n5965));
  jnot g05710(.din(n5965), .dout(n5966));
  jand g05711(.dina(n5966), .dinb(n5964), .dout(n5967));
  jnot g05712(.din(n5967), .dout(n5968));
  jor  g05713(.dina(n5769), .dinb(n5761), .dout(n5969));
  jand g05714(.dina(n5770), .dinb(n5746), .dout(n5970));
  jnot g05715(.din(n5970), .dout(n5971));
  jand g05716(.dina(n5971), .dinb(n5969), .dout(n5972));
  jnot g05717(.din(n5972), .dout(n5973));
  jor  g05718(.dina(n5751), .dinb(n5530), .dout(n5974));
  jor  g05719(.dina(n5974), .dinb(n5754), .dout(n5975));
  jnot g05720(.din(n5975), .dout(n5976));
  jand g05721(.dina(n5976), .dinb(b0 ), .dout(n5977));
  jand g05722(.dina(n5755), .dinb(b2 ), .dout(n5978));
  jor  g05723(.dina(n5978), .dinb(n5977), .dout(n5979));
  jand g05724(.dina(n5748), .dinb(n273), .dout(n5980));
  jand g05725(.dina(n5752), .dinb(b1 ), .dout(n5981));
  jor  g05726(.dina(n5981), .dinb(n5980), .dout(n5982));
  jor  g05727(.dina(n5982), .dinb(n5979), .dout(n5983));
  jnot g05728(.din(n5758), .dout(n5984));
  jand g05729(.dina(n5532), .dinb(a47 ), .dout(n5985));
  jand g05730(.dina(n5985), .dinb(n5984), .dout(n5986));
  jnot g05731(.din(n5986), .dout(n5987));
  jand g05732(.dina(n5987), .dinb(a47 ), .dout(n5988));
  jxor g05733(.dina(n5988), .dinb(n5983), .dout(n5989));
  jnot g05734(.din(n5989), .dout(n5990));
  jor  g05735(.dina(n5537), .dinb(n374), .dout(n5991));
  jor  g05736(.dina(n5534), .dinb(n340), .dout(n5992));
  jor  g05737(.dina(n5315), .dinb(n303), .dout(n5993));
  jand g05738(.dina(n5993), .dinb(n5992), .dout(n5994));
  jor  g05739(.dina(n5539), .dinb(n377), .dout(n5995));
  jand g05740(.dina(n5995), .dinb(n5994), .dout(n5996));
  jand g05741(.dina(n5996), .dinb(n5991), .dout(n5997));
  jxor g05742(.dina(n5997), .dinb(a44 ), .dout(n5998));
  jxor g05743(.dina(n5998), .dinb(n5990), .dout(n5999));
  jxor g05744(.dina(n5999), .dinb(n5973), .dout(n6000));
  jor  g05745(.dina(n4902), .dinb(n517), .dout(n6001));
  jor  g05746(.dina(n4904), .dinb(n469), .dout(n6002));
  jor  g05747(.dina(n4899), .dinb(n519), .dout(n6003));
  jor  g05748(.dina(n4696), .dinb(n415), .dout(n6004));
  jand g05749(.dina(n6004), .dinb(n6003), .dout(n6005));
  jand g05750(.dina(n6005), .dinb(n6002), .dout(n6006));
  jand g05751(.dina(n6006), .dinb(n6001), .dout(n6007));
  jxor g05752(.dina(n6007), .dinb(n4505), .dout(n6008));
  jxor g05753(.dina(n6008), .dinb(n6000), .dout(n6009));
  jxor g05754(.dina(n6009), .dinb(n5968), .dout(n6010));
  jor  g05755(.dina(n4305), .dinb(n702), .dout(n6011));
  jor  g05756(.dina(n4116), .dinb(n572), .dout(n6012));
  jor  g05757(.dina(n4308), .dinb(n637), .dout(n6013));
  jor  g05758(.dina(n4303), .dinb(n704), .dout(n6014));
  jand g05759(.dina(n6014), .dinb(n6013), .dout(n6015));
  jand g05760(.dina(n6015), .dinb(n6012), .dout(n6016));
  jand g05761(.dina(n6016), .dinb(n6011), .dout(n6017));
  jxor g05762(.dina(n6017), .dinb(n3938), .dout(n6018));
  jxor g05763(.dina(n6018), .dinb(n6010), .dout(n6019));
  jxor g05764(.dina(n6019), .dinb(n5963), .dout(n6020));
  jor  g05765(.dina(n3751), .dinb(n932), .dout(n6021));
  jor  g05766(.dina(n3574), .dinb(n772), .dout(n6022));
  jor  g05767(.dina(n3754), .dinb(n852), .dout(n6023));
  jor  g05768(.dina(n3749), .dinb(n934), .dout(n6024));
  jand g05769(.dina(n6024), .dinb(n6023), .dout(n6025));
  jand g05770(.dina(n6025), .dinb(n6022), .dout(n6026));
  jand g05771(.dina(n6026), .dinb(n6021), .dout(n6027));
  jxor g05772(.dina(n6027), .dinb(n3410), .dout(n6028));
  jxor g05773(.dina(n6028), .dinb(n6020), .dout(n6029));
  jxor g05774(.dina(n6029), .dinb(n5960), .dout(n6030));
  jor  g05775(.dina(n3239), .dinb(n1209), .dout(n6031));
  jor  g05776(.dina(n3072), .dinb(n1018), .dout(n6032));
  jor  g05777(.dina(n3237), .dinb(n1211), .dout(n6033));
  jor  g05778(.dina(n3242), .dinb(n1114), .dout(n6034));
  jand g05779(.dina(n6034), .dinb(n6033), .dout(n6035));
  jand g05780(.dina(n6035), .dinb(n6032), .dout(n6036));
  jand g05781(.dina(n6036), .dinb(n6031), .dout(n6037));
  jxor g05782(.dina(n6037), .dinb(n2918), .dout(n6038));
  jxor g05783(.dina(n6038), .dinb(n6030), .dout(n6039));
  jxor g05784(.dina(n6039), .dinb(n5957), .dout(n6040));
  jor  g05785(.dina(n2764), .dinb(n1525), .dout(n6041));
  jor  g05786(.dina(n2609), .dinb(n1307), .dout(n6042));
  jor  g05787(.dina(n2761), .dinb(n1527), .dout(n6043));
  jor  g05788(.dina(n2766), .dinb(n1416), .dout(n6044));
  jand g05789(.dina(n6044), .dinb(n6043), .dout(n6045));
  jand g05790(.dina(n6045), .dinb(n6042), .dout(n6046));
  jand g05791(.dina(n6046), .dinb(n6041), .dout(n6047));
  jxor g05792(.dina(n6047), .dinb(n2468), .dout(n6048));
  jxor g05793(.dina(n6048), .dinb(n6040), .dout(n6049));
  jxor g05794(.dina(n6049), .dinb(n5954), .dout(n6050));
  jor  g05795(.dina(n2324), .dinb(n1879), .dout(n6051));
  jor  g05796(.dina(n2186), .dinb(n1637), .dout(n6052));
  jor  g05797(.dina(n2326), .dinb(n1881), .dout(n6053));
  jor  g05798(.dina(n2321), .dinb(n1759), .dout(n6054));
  jand g05799(.dina(n6054), .dinb(n6053), .dout(n6055));
  jand g05800(.dina(n6055), .dinb(n6052), .dout(n6056));
  jand g05801(.dina(n6056), .dinb(n6051), .dout(n6057));
  jxor g05802(.dina(n6057), .dinb(n2057), .dout(n6058));
  jxor g05803(.dina(n6058), .dinb(n6050), .dout(n6059));
  jxor g05804(.dina(n6059), .dinb(n5951), .dout(n6060));
  jor  g05805(.dina(n2277), .dinb(n1921), .dout(n6061));
  jor  g05806(.dina(n1806), .dinb(n2007), .dout(n6062));
  jor  g05807(.dina(n1918), .dinb(n2142), .dout(n6063));
  jor  g05808(.dina(n1923), .dinb(n2279), .dout(n6064));
  jand g05809(.dina(n6064), .dinb(n6063), .dout(n6065));
  jand g05810(.dina(n6065), .dinb(n6062), .dout(n6066));
  jand g05811(.dina(n6066), .dinb(n6061), .dout(n6067));
  jxor g05812(.dina(n6067), .dinb(n1687), .dout(n6068));
  jxor g05813(.dina(n6068), .dinb(n6060), .dout(n6069));
  jxor g05814(.dina(n6069), .dinb(n5948), .dout(n6070));
  jor  g05815(.dina(n2711), .dinb(n1569), .dout(n6071));
  jor  g05816(.dina(n1453), .dinb(n2415), .dout(n6072));
  jor  g05817(.dina(n1566), .dinb(n2563), .dout(n6073));
  jor  g05818(.dina(n1571), .dinb(n2713), .dout(n6074));
  jand g05819(.dina(n6074), .dinb(n6073), .dout(n6075));
  jand g05820(.dina(n6075), .dinb(n6072), .dout(n6076));
  jand g05821(.dina(n6076), .dinb(n6071), .dout(n6077));
  jxor g05822(.dina(n6077), .dinb(n1351), .dout(n6078));
  jxor g05823(.dina(n6078), .dinb(n6070), .dout(n6079));
  jxor g05824(.dina(n6079), .dinb(n5945), .dout(n6080));
  jor  g05825(.dina(n3184), .dinb(n1248), .dout(n6081));
  jor  g05826(.dina(n1147), .dinb(n2862), .dout(n6082));
  jor  g05827(.dina(n1251), .dinb(n3023), .dout(n6083));
  jor  g05828(.dina(n1246), .dinb(n3186), .dout(n6084));
  jand g05829(.dina(n6084), .dinb(n6083), .dout(n6085));
  jand g05830(.dina(n6085), .dinb(n6082), .dout(n6086));
  jand g05831(.dina(n6086), .dinb(n6081), .dout(n6087));
  jxor g05832(.dina(n6087), .dinb(n1061), .dout(n6088));
  jxor g05833(.dina(n6088), .dinb(n6080), .dout(n6089));
  jxor g05834(.dina(n6089), .dinb(n5942), .dout(n6090));
  jor  g05835(.dina(n3696), .dinb(n970), .dout(n6091));
  jor  g05836(.dina(n880), .dinb(n3348), .dout(n6092));
  jor  g05837(.dina(n967), .dinb(n3522), .dout(n6093));
  jor  g05838(.dina(n972), .dinb(n3698), .dout(n6094));
  jand g05839(.dina(n6094), .dinb(n6093), .dout(n6095));
  jand g05840(.dina(n6095), .dinb(n6092), .dout(n6096));
  jand g05841(.dina(n6096), .dinb(n6091), .dout(n6097));
  jxor g05842(.dina(n6097), .dinb(n810), .dout(n6098));
  jxor g05843(.dina(n6098), .dinb(n6090), .dout(n6099));
  jxor g05844(.dina(n6099), .dinb(n5939), .dout(n6100));
  jor  g05845(.dina(n4247), .dinb(n728), .dout(n6101));
  jor  g05846(.dina(n660), .dinb(n3873), .dout(n6102));
  jor  g05847(.dina(n731), .dinb(n4060), .dout(n6103));
  jor  g05848(.dina(n726), .dinb(n4249), .dout(n6104));
  jand g05849(.dina(n6104), .dinb(n6103), .dout(n6105));
  jand g05850(.dina(n6105), .dinb(n6102), .dout(n6106));
  jand g05851(.dina(n6106), .dinb(n6101), .dout(n6107));
  jxor g05852(.dina(n6107), .dinb(n606), .dout(n6108));
  jxor g05853(.dina(n6108), .dinb(n6100), .dout(n6109));
  jnot g05854(.din(n6109), .dout(n6110));
  jxor g05855(.dina(n6110), .dinb(n5936), .dout(n6111));
  jor  g05856(.dina(n4837), .dinb(n544), .dout(n6112));
  jor  g05857(.dina(n486), .dinb(n4437), .dout(n6113));
  jor  g05858(.dina(n542), .dinb(n4839), .dout(n6114));
  jor  g05859(.dina(n547), .dinb(n4637), .dout(n6115));
  jand g05860(.dina(n6115), .dinb(n6114), .dout(n6116));
  jand g05861(.dina(n6116), .dinb(n6113), .dout(n6117));
  jand g05862(.dina(n6117), .dinb(n6112), .dout(n6118));
  jxor g05863(.dina(n6118), .dinb(n446), .dout(n6119));
  jxor g05864(.dina(n6119), .dinb(n6111), .dout(n6120));
  jxor g05865(.dina(n6120), .dinb(n5932), .dout(n6121));
  jor  g05866(.dina(n5467), .dinb(n397), .dout(n6122));
  jor  g05867(.dina(n354), .dinb(n5040), .dout(n6123));
  jor  g05868(.dina(n394), .dinb(n5253), .dout(n6124));
  jor  g05869(.dina(n399), .dinb(n5469), .dout(n6125));
  jand g05870(.dina(n6125), .dinb(n6124), .dout(n6126));
  jand g05871(.dina(n6126), .dinb(n6123), .dout(n6127));
  jand g05872(.dina(n6127), .dinb(n6122), .dout(n6128));
  jxor g05873(.dina(n6128), .dinb(n364), .dout(n6129));
  jxor g05874(.dina(n6129), .dinb(n6121), .dout(n6130));
  jxor g05875(.dina(n6130), .dinb(n5929), .dout(n6131));
  jand g05876(.dina(b46 ), .dinb(b45 ), .dout(n6132));
  jand g05877(.dina(n5907), .dinb(n5906), .dout(n6133));
  jor  g05878(.dina(n6133), .dinb(n6132), .dout(n6134));
  jxor g05879(.dina(b47 ), .dinb(b46 ), .dout(n6135));
  jnot g05880(.din(n6135), .dout(n6136));
  jxor g05881(.dina(n6136), .dinb(n6134), .dout(n6137));
  jor  g05882(.dina(n6137), .dinb(n296), .dout(n6138));
  jnot g05883(.din(b47 ), .dout(n6139));
  jor  g05884(.dina(n264), .dinb(n6139), .dout(n6140));
  jor  g05885(.dina(n294), .dinb(n5911), .dout(n6141));
  jor  g05886(.dina(n280), .dinb(n5685), .dout(n6142));
  jand g05887(.dina(n6142), .dinb(n6141), .dout(n6143));
  jand g05888(.dina(n6143), .dinb(n6140), .dout(n6144));
  jand g05889(.dina(n6144), .dinb(n6138), .dout(n6145));
  jxor g05890(.dina(n6145), .dinb(n278), .dout(n6146));
  jxor g05891(.dina(n6146), .dinb(n6131), .dout(n6147));
  jxor g05892(.dina(n6147), .dinb(n5924), .dout(f47 ));
  jnot g05893(.din(n6146), .dout(n6149));
  jor  g05894(.dina(n6149), .dinb(n6131), .dout(n6150));
  jor  g05895(.dina(n6147), .dinb(n5924), .dout(n6151));
  jand g05896(.dina(n6151), .dinb(n6150), .dout(n6152));
  jand g05897(.dina(n6129), .dinb(n6121), .dout(n6153));
  jnot g05898(.din(n6153), .dout(n6154));
  jnot g05899(.din(n6130), .dout(n6155));
  jor  g05900(.dina(n6155), .dinb(n5929), .dout(n6156));
  jand g05901(.dina(n6156), .dinb(n6154), .dout(n6157));
  jand g05902(.dina(n6119), .dinb(n6111), .dout(n6158));
  jand g05903(.dina(n6120), .dinb(n5932), .dout(n6159));
  jor  g05904(.dina(n6159), .dinb(n6158), .dout(n6160));
  jand g05905(.dina(n6108), .dinb(n6100), .dout(n6161));
  jnot g05906(.din(n6161), .dout(n6162));
  jor  g05907(.dina(n6110), .dinb(n5936), .dout(n6163));
  jand g05908(.dina(n6163), .dinb(n6162), .dout(n6164));
  jand g05909(.dina(n6098), .dinb(n6090), .dout(n6165));
  jand g05910(.dina(n6099), .dinb(n5939), .dout(n6166));
  jor  g05911(.dina(n6166), .dinb(n6165), .dout(n6167));
  jand g05912(.dina(n6088), .dinb(n6080), .dout(n6168));
  jand g05913(.dina(n6089), .dinb(n5942), .dout(n6169));
  jor  g05914(.dina(n6169), .dinb(n6168), .dout(n6170));
  jand g05915(.dina(n6078), .dinb(n6070), .dout(n6171));
  jand g05916(.dina(n6079), .dinb(n5945), .dout(n6172));
  jor  g05917(.dina(n6172), .dinb(n6171), .dout(n6173));
  jand g05918(.dina(n6068), .dinb(n6060), .dout(n6174));
  jand g05919(.dina(n6069), .dinb(n5948), .dout(n6175));
  jor  g05920(.dina(n6175), .dinb(n6174), .dout(n6176));
  jand g05921(.dina(n6058), .dinb(n6050), .dout(n6177));
  jand g05922(.dina(n6059), .dinb(n5951), .dout(n6178));
  jor  g05923(.dina(n6178), .dinb(n6177), .dout(n6179));
  jand g05924(.dina(n6048), .dinb(n6040), .dout(n6180));
  jand g05925(.dina(n6049), .dinb(n5954), .dout(n6181));
  jor  g05926(.dina(n6181), .dinb(n6180), .dout(n6182));
  jand g05927(.dina(n6038), .dinb(n6030), .dout(n6183));
  jand g05928(.dina(n6039), .dinb(n5957), .dout(n6184));
  jor  g05929(.dina(n6184), .dinb(n6183), .dout(n6185));
  jand g05930(.dina(n6028), .dinb(n6020), .dout(n6186));
  jand g05931(.dina(n6029), .dinb(n5960), .dout(n6187));
  jor  g05932(.dina(n6187), .dinb(n6186), .dout(n6188));
  jand g05933(.dina(n6018), .dinb(n6010), .dout(n6189));
  jand g05934(.dina(n6019), .dinb(n5963), .dout(n6190));
  jor  g05935(.dina(n6190), .dinb(n6189), .dout(n6191));
  jand g05936(.dina(n6008), .dinb(n6000), .dout(n6192));
  jand g05937(.dina(n6009), .dinb(n5968), .dout(n6193));
  jor  g05938(.dina(n6193), .dinb(n6192), .dout(n6194));
  jor  g05939(.dina(n5998), .dinb(n5990), .dout(n6195));
  jand g05940(.dina(n5999), .dinb(n5973), .dout(n6196));
  jnot g05941(.din(n6196), .dout(n6197));
  jand g05942(.dina(n6197), .dinb(n6195), .dout(n6198));
  jnot g05943(.din(n6198), .dout(n6199));
  jor  g05944(.dina(n5987), .dinb(n5983), .dout(n6200));
  jxor g05945(.dina(a48 ), .dinb(a47 ), .dout(n6201));
  jand g05946(.dina(n6201), .dinb(b0 ), .dout(n6202));
  jnot g05947(.din(n6202), .dout(n6203));
  jxor g05948(.dina(n6203), .dinb(n6200), .dout(n6204));
  jnot g05949(.din(n5755), .dout(n6205));
  jor  g05950(.dina(n6205), .dinb(n303), .dout(n6206));
  jnot g05951(.din(n5748), .dout(n6207));
  jor  g05952(.dina(n6207), .dinb(n301), .dout(n6208));
  jor  g05953(.dina(n5975), .dinb(n305), .dout(n6209));
  jnot g05954(.din(n5752), .dout(n6210));
  jor  g05955(.dina(n6210), .dinb(n293), .dout(n6211));
  jand g05956(.dina(n6211), .dinb(n6209), .dout(n6212));
  jand g05957(.dina(n6212), .dinb(n6208), .dout(n6213));
  jand g05958(.dina(n6213), .dinb(n6206), .dout(n6214));
  jxor g05959(.dina(n6214), .dinb(n5759), .dout(n6215));
  jxor g05960(.dina(n6215), .dinb(n6204), .dout(n6216));
  jnot g05961(.din(n6216), .dout(n6217));
  jor  g05962(.dina(n5537), .dinb(n412), .dout(n6218));
  jor  g05963(.dina(n5534), .dinb(n377), .dout(n6219));
  jor  g05964(.dina(n5315), .dinb(n340), .dout(n6220));
  jand g05965(.dina(n6220), .dinb(n6219), .dout(n6221));
  jor  g05966(.dina(n5539), .dinb(n415), .dout(n6222));
  jand g05967(.dina(n6222), .dinb(n6221), .dout(n6223));
  jand g05968(.dina(n6223), .dinb(n6218), .dout(n6224));
  jxor g05969(.dina(n6224), .dinb(a44 ), .dout(n6225));
  jxor g05970(.dina(n6225), .dinb(n6217), .dout(n6226));
  jxor g05971(.dina(n6226), .dinb(n6199), .dout(n6227));
  jor  g05972(.dina(n4902), .dinb(n570), .dout(n6228));
  jor  g05973(.dina(n4696), .dinb(n469), .dout(n6229));
  jor  g05974(.dina(n4899), .dinb(n572), .dout(n6230));
  jor  g05975(.dina(n4904), .dinb(n519), .dout(n6231));
  jand g05976(.dina(n6231), .dinb(n6230), .dout(n6232));
  jand g05977(.dina(n6232), .dinb(n6229), .dout(n6233));
  jand g05978(.dina(n6233), .dinb(n6228), .dout(n6234));
  jxor g05979(.dina(n6234), .dinb(n4505), .dout(n6235));
  jxor g05980(.dina(n6235), .dinb(n6227), .dout(n6236));
  jxor g05981(.dina(n6236), .dinb(n6194), .dout(n6237));
  jor  g05982(.dina(n4305), .dinb(n770), .dout(n6238));
  jor  g05983(.dina(n4116), .dinb(n637), .dout(n6239));
  jor  g05984(.dina(n4308), .dinb(n704), .dout(n6240));
  jor  g05985(.dina(n4303), .dinb(n772), .dout(n6241));
  jand g05986(.dina(n6241), .dinb(n6240), .dout(n6242));
  jand g05987(.dina(n6242), .dinb(n6239), .dout(n6243));
  jand g05988(.dina(n6243), .dinb(n6238), .dout(n6244));
  jxor g05989(.dina(n6244), .dinb(n3938), .dout(n6245));
  jxor g05990(.dina(n6245), .dinb(n6237), .dout(n6246));
  jxor g05991(.dina(n6246), .dinb(n6191), .dout(n6247));
  jor  g05992(.dina(n3751), .dinb(n1016), .dout(n6248));
  jor  g05993(.dina(n3574), .dinb(n852), .dout(n6249));
  jor  g05994(.dina(n3754), .dinb(n934), .dout(n6250));
  jor  g05995(.dina(n3749), .dinb(n1018), .dout(n6251));
  jand g05996(.dina(n6251), .dinb(n6250), .dout(n6252));
  jand g05997(.dina(n6252), .dinb(n6249), .dout(n6253));
  jand g05998(.dina(n6253), .dinb(n6248), .dout(n6254));
  jxor g05999(.dina(n6254), .dinb(n3410), .dout(n6255));
  jxor g06000(.dina(n6255), .dinb(n6247), .dout(n6256));
  jxor g06001(.dina(n6256), .dinb(n6188), .dout(n6257));
  jor  g06002(.dina(n3239), .dinb(n1305), .dout(n6258));
  jor  g06003(.dina(n3072), .dinb(n1114), .dout(n6259));
  jor  g06004(.dina(n3237), .dinb(n1307), .dout(n6260));
  jor  g06005(.dina(n3242), .dinb(n1211), .dout(n6261));
  jand g06006(.dina(n6261), .dinb(n6260), .dout(n6262));
  jand g06007(.dina(n6262), .dinb(n6259), .dout(n6263));
  jand g06008(.dina(n6263), .dinb(n6258), .dout(n6264));
  jxor g06009(.dina(n6264), .dinb(n2918), .dout(n6265));
  jxor g06010(.dina(n6265), .dinb(n6257), .dout(n6266));
  jxor g06011(.dina(n6266), .dinb(n6185), .dout(n6267));
  jor  g06012(.dina(n2764), .dinb(n1635), .dout(n6268));
  jor  g06013(.dina(n2609), .dinb(n1416), .dout(n6269));
  jor  g06014(.dina(n2761), .dinb(n1637), .dout(n6270));
  jor  g06015(.dina(n2766), .dinb(n1527), .dout(n6271));
  jand g06016(.dina(n6271), .dinb(n6270), .dout(n6272));
  jand g06017(.dina(n6272), .dinb(n6269), .dout(n6273));
  jand g06018(.dina(n6273), .dinb(n6268), .dout(n6274));
  jxor g06019(.dina(n6274), .dinb(n2468), .dout(n6275));
  jxor g06020(.dina(n6275), .dinb(n6267), .dout(n6276));
  jxor g06021(.dina(n6276), .dinb(n6182), .dout(n6277));
  jor  g06022(.dina(n2324), .dinb(n2005), .dout(n6278));
  jor  g06023(.dina(n2186), .dinb(n1759), .dout(n6279));
  jor  g06024(.dina(n2321), .dinb(n1881), .dout(n6280));
  jor  g06025(.dina(n2326), .dinb(n2007), .dout(n6281));
  jand g06026(.dina(n6281), .dinb(n6280), .dout(n6282));
  jand g06027(.dina(n6282), .dinb(n6279), .dout(n6283));
  jand g06028(.dina(n6283), .dinb(n6278), .dout(n6284));
  jxor g06029(.dina(n6284), .dinb(n2057), .dout(n6285));
  jxor g06030(.dina(n6285), .dinb(n6277), .dout(n6286));
  jxor g06031(.dina(n6286), .dinb(n6179), .dout(n6287));
  jor  g06032(.dina(n2413), .dinb(n1921), .dout(n6288));
  jor  g06033(.dina(n1806), .dinb(n2142), .dout(n6289));
  jor  g06034(.dina(n1918), .dinb(n2279), .dout(n6290));
  jor  g06035(.dina(n1923), .dinb(n2415), .dout(n6291));
  jand g06036(.dina(n6291), .dinb(n6290), .dout(n6292));
  jand g06037(.dina(n6292), .dinb(n6289), .dout(n6293));
  jand g06038(.dina(n6293), .dinb(n6288), .dout(n6294));
  jxor g06039(.dina(n6294), .dinb(n1687), .dout(n6295));
  jxor g06040(.dina(n6295), .dinb(n6287), .dout(n6296));
  jxor g06041(.dina(n6296), .dinb(n6176), .dout(n6297));
  jor  g06042(.dina(n2860), .dinb(n1569), .dout(n6298));
  jor  g06043(.dina(n1453), .dinb(n2563), .dout(n6299));
  jor  g06044(.dina(n1566), .dinb(n2713), .dout(n6300));
  jor  g06045(.dina(n1571), .dinb(n2862), .dout(n6301));
  jand g06046(.dina(n6301), .dinb(n6300), .dout(n6302));
  jand g06047(.dina(n6302), .dinb(n6299), .dout(n6303));
  jand g06048(.dina(n6303), .dinb(n6298), .dout(n6304));
  jxor g06049(.dina(n6304), .dinb(n1351), .dout(n6305));
  jxor g06050(.dina(n6305), .dinb(n6297), .dout(n6306));
  jxor g06051(.dina(n6306), .dinb(n6173), .dout(n6307));
  jor  g06052(.dina(n3346), .dinb(n1248), .dout(n6308));
  jor  g06053(.dina(n1147), .dinb(n3023), .dout(n6309));
  jor  g06054(.dina(n1251), .dinb(n3186), .dout(n6310));
  jor  g06055(.dina(n1246), .dinb(n3348), .dout(n6311));
  jand g06056(.dina(n6311), .dinb(n6310), .dout(n6312));
  jand g06057(.dina(n6312), .dinb(n6309), .dout(n6313));
  jand g06058(.dina(n6313), .dinb(n6308), .dout(n6314));
  jxor g06059(.dina(n6314), .dinb(n1061), .dout(n6315));
  jxor g06060(.dina(n6315), .dinb(n6307), .dout(n6316));
  jxor g06061(.dina(n6316), .dinb(n6170), .dout(n6317));
  jor  g06062(.dina(n3871), .dinb(n970), .dout(n6318));
  jor  g06063(.dina(n880), .dinb(n3522), .dout(n6319));
  jor  g06064(.dina(n972), .dinb(n3873), .dout(n6320));
  jor  g06065(.dina(n967), .dinb(n3698), .dout(n6321));
  jand g06066(.dina(n6321), .dinb(n6320), .dout(n6322));
  jand g06067(.dina(n6322), .dinb(n6319), .dout(n6323));
  jand g06068(.dina(n6323), .dinb(n6318), .dout(n6324));
  jxor g06069(.dina(n6324), .dinb(n810), .dout(n6325));
  jxor g06070(.dina(n6325), .dinb(n6317), .dout(n6326));
  jxor g06071(.dina(n6326), .dinb(n6167), .dout(n6327));
  jor  g06072(.dina(n4435), .dinb(n728), .dout(n6328));
  jor  g06073(.dina(n660), .dinb(n4060), .dout(n6329));
  jor  g06074(.dina(n731), .dinb(n4249), .dout(n6330));
  jor  g06075(.dina(n726), .dinb(n4437), .dout(n6331));
  jand g06076(.dina(n6331), .dinb(n6330), .dout(n6332));
  jand g06077(.dina(n6332), .dinb(n6329), .dout(n6333));
  jand g06078(.dina(n6333), .dinb(n6328), .dout(n6334));
  jxor g06079(.dina(n6334), .dinb(n606), .dout(n6335));
  jxor g06080(.dina(n6335), .dinb(n6327), .dout(n6336));
  jnot g06081(.din(n6336), .dout(n6337));
  jxor g06082(.dina(n6337), .dinb(n6164), .dout(n6338));
  jor  g06083(.dina(n5038), .dinb(n544), .dout(n6339));
  jor  g06084(.dina(n486), .dinb(n4637), .dout(n6340));
  jor  g06085(.dina(n542), .dinb(n5040), .dout(n6341));
  jor  g06086(.dina(n547), .dinb(n4839), .dout(n6342));
  jand g06087(.dina(n6342), .dinb(n6341), .dout(n6343));
  jand g06088(.dina(n6343), .dinb(n6340), .dout(n6344));
  jand g06089(.dina(n6344), .dinb(n6339), .dout(n6345));
  jxor g06090(.dina(n6345), .dinb(n446), .dout(n6346));
  jxor g06091(.dina(n6346), .dinb(n6338), .dout(n6347));
  jxor g06092(.dina(n6347), .dinb(n6160), .dout(n6348));
  jor  g06093(.dina(n5683), .dinb(n397), .dout(n6349));
  jor  g06094(.dina(n354), .dinb(n5253), .dout(n6350));
  jor  g06095(.dina(n394), .dinb(n5469), .dout(n6351));
  jor  g06096(.dina(n399), .dinb(n5685), .dout(n6352));
  jand g06097(.dina(n6352), .dinb(n6351), .dout(n6353));
  jand g06098(.dina(n6353), .dinb(n6350), .dout(n6354));
  jand g06099(.dina(n6354), .dinb(n6349), .dout(n6355));
  jxor g06100(.dina(n6355), .dinb(n364), .dout(n6356));
  jxor g06101(.dina(n6356), .dinb(n6348), .dout(n6357));
  jxor g06102(.dina(n6357), .dinb(n6157), .dout(n6358));
  jand g06103(.dina(b47 ), .dinb(b46 ), .dout(n6359));
  jand g06104(.dina(n6135), .dinb(n6134), .dout(n6360));
  jor  g06105(.dina(n6360), .dinb(n6359), .dout(n6361));
  jxor g06106(.dina(b48 ), .dinb(b47 ), .dout(n6362));
  jnot g06107(.din(n6362), .dout(n6363));
  jxor g06108(.dina(n6363), .dinb(n6361), .dout(n6364));
  jor  g06109(.dina(n6364), .dinb(n296), .dout(n6365));
  jnot g06110(.din(b48 ), .dout(n6366));
  jor  g06111(.dina(n264), .dinb(n6366), .dout(n6367));
  jor  g06112(.dina(n294), .dinb(n6139), .dout(n6368));
  jor  g06113(.dina(n280), .dinb(n5911), .dout(n6369));
  jand g06114(.dina(n6369), .dinb(n6368), .dout(n6370));
  jand g06115(.dina(n6370), .dinb(n6367), .dout(n6371));
  jand g06116(.dina(n6371), .dinb(n6365), .dout(n6372));
  jxor g06117(.dina(n6372), .dinb(n278), .dout(n6373));
  jxor g06118(.dina(n6373), .dinb(n6358), .dout(n6374));
  jxor g06119(.dina(n6374), .dinb(n6152), .dout(f48 ));
  jnot g06120(.din(n6373), .dout(n6376));
  jor  g06121(.dina(n6376), .dinb(n6358), .dout(n6377));
  jor  g06122(.dina(n6374), .dinb(n6152), .dout(n6378));
  jand g06123(.dina(n6378), .dinb(n6377), .dout(n6379));
  jand g06124(.dina(n6356), .dinb(n6348), .dout(n6380));
  jnot g06125(.din(n6380), .dout(n6381));
  jnot g06126(.din(n6357), .dout(n6382));
  jor  g06127(.dina(n6382), .dinb(n6157), .dout(n6383));
  jand g06128(.dina(n6383), .dinb(n6381), .dout(n6384));
  jand g06129(.dina(n6346), .dinb(n6338), .dout(n6385));
  jand g06130(.dina(n6347), .dinb(n6160), .dout(n6386));
  jor  g06131(.dina(n6386), .dinb(n6385), .dout(n6387));
  jand g06132(.dina(n6335), .dinb(n6327), .dout(n6388));
  jnot g06133(.din(n6388), .dout(n6389));
  jor  g06134(.dina(n6337), .dinb(n6164), .dout(n6390));
  jand g06135(.dina(n6390), .dinb(n6389), .dout(n6391));
  jand g06136(.dina(n6325), .dinb(n6317), .dout(n6392));
  jand g06137(.dina(n6326), .dinb(n6167), .dout(n6393));
  jor  g06138(.dina(n6393), .dinb(n6392), .dout(n6394));
  jand g06139(.dina(n6315), .dinb(n6307), .dout(n6395));
  jand g06140(.dina(n6316), .dinb(n6170), .dout(n6396));
  jor  g06141(.dina(n6396), .dinb(n6395), .dout(n6397));
  jand g06142(.dina(n6305), .dinb(n6297), .dout(n6398));
  jand g06143(.dina(n6306), .dinb(n6173), .dout(n6399));
  jor  g06144(.dina(n6399), .dinb(n6398), .dout(n6400));
  jand g06145(.dina(n6295), .dinb(n6287), .dout(n6401));
  jand g06146(.dina(n6296), .dinb(n6176), .dout(n6402));
  jor  g06147(.dina(n6402), .dinb(n6401), .dout(n6403));
  jand g06148(.dina(n6285), .dinb(n6277), .dout(n6404));
  jand g06149(.dina(n6286), .dinb(n6179), .dout(n6405));
  jor  g06150(.dina(n6405), .dinb(n6404), .dout(n6406));
  jand g06151(.dina(n6275), .dinb(n6267), .dout(n6407));
  jand g06152(.dina(n6276), .dinb(n6182), .dout(n6408));
  jor  g06153(.dina(n6408), .dinb(n6407), .dout(n6409));
  jand g06154(.dina(n6265), .dinb(n6257), .dout(n6410));
  jand g06155(.dina(n6266), .dinb(n6185), .dout(n6411));
  jor  g06156(.dina(n6411), .dinb(n6410), .dout(n6412));
  jand g06157(.dina(n6255), .dinb(n6247), .dout(n6413));
  jand g06158(.dina(n6256), .dinb(n6188), .dout(n6414));
  jor  g06159(.dina(n6414), .dinb(n6413), .dout(n6415));
  jand g06160(.dina(n6245), .dinb(n6237), .dout(n6416));
  jand g06161(.dina(n6246), .dinb(n6191), .dout(n6417));
  jor  g06162(.dina(n6417), .dinb(n6416), .dout(n6418));
  jand g06163(.dina(n6235), .dinb(n6227), .dout(n6419));
  jand g06164(.dina(n6236), .dinb(n6194), .dout(n6420));
  jor  g06165(.dina(n6420), .dinb(n6419), .dout(n6421));
  jor  g06166(.dina(n6225), .dinb(n6217), .dout(n6422));
  jand g06167(.dina(n6226), .dinb(n6199), .dout(n6423));
  jnot g06168(.din(n6423), .dout(n6424));
  jand g06169(.dina(n6424), .dinb(n6422), .dout(n6425));
  jnot g06170(.din(n6425), .dout(n6426));
  jnot g06171(.din(n6200), .dout(n6427));
  jand g06172(.dina(n6202), .dinb(n6427), .dout(n6428));
  jand g06173(.dina(n6215), .dinb(n6204), .dout(n6429));
  jor  g06174(.dina(n6429), .dinb(n6428), .dout(n6430));
  jxor g06175(.dina(a50 ), .dinb(a49 ), .dout(n6431));
  jnot g06176(.din(n6431), .dout(n6432));
  jand g06177(.dina(n6432), .dinb(n6201), .dout(n6433));
  jand g06178(.dina(n6433), .dinb(b1 ), .dout(n6434));
  jand g06179(.dina(n6431), .dinb(n6201), .dout(n6435));
  jand g06180(.dina(n6435), .dinb(n259), .dout(n6436));
  jnot g06181(.din(n6201), .dout(n6437));
  jxor g06182(.dina(a49 ), .dinb(a48 ), .dout(n6438));
  jand g06183(.dina(n6438), .dinb(n6437), .dout(n6439));
  jand g06184(.dina(n6439), .dinb(b0 ), .dout(n6440));
  jor  g06185(.dina(n6440), .dinb(n6436), .dout(n6441));
  jor  g06186(.dina(n6441), .dinb(n6434), .dout(n6442));
  jnot g06187(.din(a50 ), .dout(n6443));
  jor  g06188(.dina(n6203), .dinb(n6443), .dout(n6444));
  jxor g06189(.dina(n6444), .dinb(n6442), .dout(n6445));
  jor  g06190(.dina(n6207), .dinb(n337), .dout(n6446));
  jor  g06191(.dina(n6205), .dinb(n340), .dout(n6447));
  jor  g06192(.dina(n5975), .dinb(n293), .dout(n6448));
  jand g06193(.dina(n6448), .dinb(n6447), .dout(n6449));
  jor  g06194(.dina(n6210), .dinb(n303), .dout(n6450));
  jand g06195(.dina(n6450), .dinb(n6449), .dout(n6451));
  jand g06196(.dina(n6451), .dinb(n6446), .dout(n6452));
  jxor g06197(.dina(n6452), .dinb(a47 ), .dout(n6453));
  jxor g06198(.dina(n6453), .dinb(n6445), .dout(n6454));
  jxor g06199(.dina(n6454), .dinb(n6430), .dout(n6455));
  jnot g06200(.din(n6455), .dout(n6456));
  jor  g06201(.dina(n5537), .dinb(n466), .dout(n6457));
  jor  g06202(.dina(n5539), .dinb(n469), .dout(n6458));
  jor  g06203(.dina(n5315), .dinb(n377), .dout(n6459));
  jand g06204(.dina(n6459), .dinb(n6458), .dout(n6460));
  jor  g06205(.dina(n5534), .dinb(n415), .dout(n6461));
  jand g06206(.dina(n6461), .dinb(n6460), .dout(n6462));
  jand g06207(.dina(n6462), .dinb(n6457), .dout(n6463));
  jxor g06208(.dina(n6463), .dinb(a44 ), .dout(n6464));
  jxor g06209(.dina(n6464), .dinb(n6456), .dout(n6465));
  jxor g06210(.dina(n6465), .dinb(n6426), .dout(n6466));
  jor  g06211(.dina(n4902), .dinb(n635), .dout(n6467));
  jor  g06212(.dina(n4696), .dinb(n519), .dout(n6468));
  jor  g06213(.dina(n4899), .dinb(n637), .dout(n6469));
  jor  g06214(.dina(n4904), .dinb(n572), .dout(n6470));
  jand g06215(.dina(n6470), .dinb(n6469), .dout(n6471));
  jand g06216(.dina(n6471), .dinb(n6468), .dout(n6472));
  jand g06217(.dina(n6472), .dinb(n6467), .dout(n6473));
  jxor g06218(.dina(n6473), .dinb(n4505), .dout(n6474));
  jxor g06219(.dina(n6474), .dinb(n6466), .dout(n6475));
  jxor g06220(.dina(n6475), .dinb(n6421), .dout(n6476));
  jor  g06221(.dina(n4305), .dinb(n850), .dout(n6477));
  jor  g06222(.dina(n4116), .dinb(n704), .dout(n6478));
  jor  g06223(.dina(n4303), .dinb(n852), .dout(n6479));
  jor  g06224(.dina(n4308), .dinb(n772), .dout(n6480));
  jand g06225(.dina(n6480), .dinb(n6479), .dout(n6481));
  jand g06226(.dina(n6481), .dinb(n6478), .dout(n6482));
  jand g06227(.dina(n6482), .dinb(n6477), .dout(n6483));
  jxor g06228(.dina(n6483), .dinb(n3938), .dout(n6484));
  jxor g06229(.dina(n6484), .dinb(n6476), .dout(n6485));
  jxor g06230(.dina(n6485), .dinb(n6418), .dout(n6486));
  jor  g06231(.dina(n3751), .dinb(n1112), .dout(n6487));
  jor  g06232(.dina(n3574), .dinb(n934), .dout(n6488));
  jor  g06233(.dina(n3754), .dinb(n1018), .dout(n6489));
  jor  g06234(.dina(n3749), .dinb(n1114), .dout(n6490));
  jand g06235(.dina(n6490), .dinb(n6489), .dout(n6491));
  jand g06236(.dina(n6491), .dinb(n6488), .dout(n6492));
  jand g06237(.dina(n6492), .dinb(n6487), .dout(n6493));
  jxor g06238(.dina(n6493), .dinb(n3410), .dout(n6494));
  jxor g06239(.dina(n6494), .dinb(n6486), .dout(n6495));
  jxor g06240(.dina(n6495), .dinb(n6415), .dout(n6496));
  jor  g06241(.dina(n3239), .dinb(n1414), .dout(n6497));
  jor  g06242(.dina(n3072), .dinb(n1211), .dout(n6498));
  jor  g06243(.dina(n3237), .dinb(n1416), .dout(n6499));
  jor  g06244(.dina(n3242), .dinb(n1307), .dout(n6500));
  jand g06245(.dina(n6500), .dinb(n6499), .dout(n6501));
  jand g06246(.dina(n6501), .dinb(n6498), .dout(n6502));
  jand g06247(.dina(n6502), .dinb(n6497), .dout(n6503));
  jxor g06248(.dina(n6503), .dinb(n2918), .dout(n6504));
  jxor g06249(.dina(n6504), .dinb(n6496), .dout(n6505));
  jxor g06250(.dina(n6505), .dinb(n6412), .dout(n6506));
  jor  g06251(.dina(n2764), .dinb(n1757), .dout(n6507));
  jor  g06252(.dina(n2609), .dinb(n1527), .dout(n6508));
  jor  g06253(.dina(n2761), .dinb(n1759), .dout(n6509));
  jor  g06254(.dina(n2766), .dinb(n1637), .dout(n6510));
  jand g06255(.dina(n6510), .dinb(n6509), .dout(n6511));
  jand g06256(.dina(n6511), .dinb(n6508), .dout(n6512));
  jand g06257(.dina(n6512), .dinb(n6507), .dout(n6513));
  jxor g06258(.dina(n6513), .dinb(n2468), .dout(n6514));
  jxor g06259(.dina(n6514), .dinb(n6506), .dout(n6515));
  jxor g06260(.dina(n6515), .dinb(n6409), .dout(n6516));
  jor  g06261(.dina(n2140), .dinb(n2324), .dout(n6517));
  jor  g06262(.dina(n2186), .dinb(n1881), .dout(n6518));
  jor  g06263(.dina(n2321), .dinb(n2007), .dout(n6519));
  jor  g06264(.dina(n2326), .dinb(n2142), .dout(n6520));
  jand g06265(.dina(n6520), .dinb(n6519), .dout(n6521));
  jand g06266(.dina(n6521), .dinb(n6518), .dout(n6522));
  jand g06267(.dina(n6522), .dinb(n6517), .dout(n6523));
  jxor g06268(.dina(n6523), .dinb(n2057), .dout(n6524));
  jxor g06269(.dina(n6524), .dinb(n6516), .dout(n6525));
  jxor g06270(.dina(n6525), .dinb(n6406), .dout(n6526));
  jor  g06271(.dina(n2561), .dinb(n1921), .dout(n6527));
  jor  g06272(.dina(n1806), .dinb(n2279), .dout(n6528));
  jor  g06273(.dina(n1923), .dinb(n2563), .dout(n6529));
  jor  g06274(.dina(n1918), .dinb(n2415), .dout(n6530));
  jand g06275(.dina(n6530), .dinb(n6529), .dout(n6531));
  jand g06276(.dina(n6531), .dinb(n6528), .dout(n6532));
  jand g06277(.dina(n6532), .dinb(n6527), .dout(n6533));
  jxor g06278(.dina(n6533), .dinb(n1687), .dout(n6534));
  jxor g06279(.dina(n6534), .dinb(n6526), .dout(n6535));
  jxor g06280(.dina(n6535), .dinb(n6403), .dout(n6536));
  jor  g06281(.dina(n3021), .dinb(n1569), .dout(n6537));
  jor  g06282(.dina(n1453), .dinb(n2713), .dout(n6538));
  jor  g06283(.dina(n1566), .dinb(n2862), .dout(n6539));
  jor  g06284(.dina(n1571), .dinb(n3023), .dout(n6540));
  jand g06285(.dina(n6540), .dinb(n6539), .dout(n6541));
  jand g06286(.dina(n6541), .dinb(n6538), .dout(n6542));
  jand g06287(.dina(n6542), .dinb(n6537), .dout(n6543));
  jxor g06288(.dina(n6543), .dinb(n1351), .dout(n6544));
  jxor g06289(.dina(n6544), .dinb(n6536), .dout(n6545));
  jxor g06290(.dina(n6545), .dinb(n6400), .dout(n6546));
  jor  g06291(.dina(n3520), .dinb(n1248), .dout(n6547));
  jor  g06292(.dina(n1147), .dinb(n3186), .dout(n6548));
  jor  g06293(.dina(n1246), .dinb(n3522), .dout(n6549));
  jor  g06294(.dina(n1251), .dinb(n3348), .dout(n6550));
  jand g06295(.dina(n6550), .dinb(n6549), .dout(n6551));
  jand g06296(.dina(n6551), .dinb(n6548), .dout(n6552));
  jand g06297(.dina(n6552), .dinb(n6547), .dout(n6553));
  jxor g06298(.dina(n6553), .dinb(n1061), .dout(n6554));
  jxor g06299(.dina(n6554), .dinb(n6546), .dout(n6555));
  jxor g06300(.dina(n6555), .dinb(n6397), .dout(n6556));
  jor  g06301(.dina(n4058), .dinb(n970), .dout(n6557));
  jor  g06302(.dina(n880), .dinb(n3698), .dout(n6558));
  jor  g06303(.dina(n967), .dinb(n3873), .dout(n6559));
  jor  g06304(.dina(n972), .dinb(n4060), .dout(n6560));
  jand g06305(.dina(n6560), .dinb(n6559), .dout(n6561));
  jand g06306(.dina(n6561), .dinb(n6558), .dout(n6562));
  jand g06307(.dina(n6562), .dinb(n6557), .dout(n6563));
  jxor g06308(.dina(n6563), .dinb(n810), .dout(n6564));
  jxor g06309(.dina(n6564), .dinb(n6556), .dout(n6565));
  jxor g06310(.dina(n6565), .dinb(n6394), .dout(n6566));
  jor  g06311(.dina(n4635), .dinb(n728), .dout(n6567));
  jor  g06312(.dina(n660), .dinb(n4249), .dout(n6568));
  jor  g06313(.dina(n726), .dinb(n4637), .dout(n6569));
  jor  g06314(.dina(n731), .dinb(n4437), .dout(n6570));
  jand g06315(.dina(n6570), .dinb(n6569), .dout(n6571));
  jand g06316(.dina(n6571), .dinb(n6568), .dout(n6572));
  jand g06317(.dina(n6572), .dinb(n6567), .dout(n6573));
  jxor g06318(.dina(n6573), .dinb(n606), .dout(n6574));
  jxor g06319(.dina(n6574), .dinb(n6566), .dout(n6575));
  jnot g06320(.din(n6575), .dout(n6576));
  jxor g06321(.dina(n6576), .dinb(n6391), .dout(n6577));
  jor  g06322(.dina(n5251), .dinb(n544), .dout(n6578));
  jor  g06323(.dina(n486), .dinb(n4839), .dout(n6579));
  jor  g06324(.dina(n547), .dinb(n5040), .dout(n6580));
  jor  g06325(.dina(n542), .dinb(n5253), .dout(n6581));
  jand g06326(.dina(n6581), .dinb(n6580), .dout(n6582));
  jand g06327(.dina(n6582), .dinb(n6579), .dout(n6583));
  jand g06328(.dina(n6583), .dinb(n6578), .dout(n6584));
  jxor g06329(.dina(n6584), .dinb(n446), .dout(n6585));
  jxor g06330(.dina(n6585), .dinb(n6577), .dout(n6586));
  jxor g06331(.dina(n6586), .dinb(n6387), .dout(n6587));
  jor  g06332(.dina(n5909), .dinb(n397), .dout(n6588));
  jor  g06333(.dina(n354), .dinb(n5469), .dout(n6589));
  jor  g06334(.dina(n399), .dinb(n5911), .dout(n6590));
  jor  g06335(.dina(n394), .dinb(n5685), .dout(n6591));
  jand g06336(.dina(n6591), .dinb(n6590), .dout(n6592));
  jand g06337(.dina(n6592), .dinb(n6589), .dout(n6593));
  jand g06338(.dina(n6593), .dinb(n6588), .dout(n6594));
  jxor g06339(.dina(n6594), .dinb(n364), .dout(n6595));
  jxor g06340(.dina(n6595), .dinb(n6587), .dout(n6596));
  jxor g06341(.dina(n6596), .dinb(n6384), .dout(n6597));
  jand g06342(.dina(b48 ), .dinb(b47 ), .dout(n6598));
  jand g06343(.dina(n6362), .dinb(n6361), .dout(n6599));
  jor  g06344(.dina(n6599), .dinb(n6598), .dout(n6600));
  jxor g06345(.dina(b49 ), .dinb(b48 ), .dout(n6601));
  jnot g06346(.din(n6601), .dout(n6602));
  jxor g06347(.dina(n6602), .dinb(n6600), .dout(n6603));
  jor  g06348(.dina(n6603), .dinb(n296), .dout(n6604));
  jnot g06349(.din(b49 ), .dout(n6605));
  jor  g06350(.dina(n264), .dinb(n6605), .dout(n6606));
  jor  g06351(.dina(n280), .dinb(n6139), .dout(n6607));
  jor  g06352(.dina(n294), .dinb(n6366), .dout(n6608));
  jand g06353(.dina(n6608), .dinb(n6607), .dout(n6609));
  jand g06354(.dina(n6609), .dinb(n6606), .dout(n6610));
  jand g06355(.dina(n6610), .dinb(n6604), .dout(n6611));
  jxor g06356(.dina(n6611), .dinb(n278), .dout(n6612));
  jxor g06357(.dina(n6612), .dinb(n6597), .dout(n6613));
  jxor g06358(.dina(n6613), .dinb(n6379), .dout(f49 ));
  jnot g06359(.din(n6612), .dout(n6615));
  jor  g06360(.dina(n6615), .dinb(n6597), .dout(n6616));
  jor  g06361(.dina(n6613), .dinb(n6379), .dout(n6617));
  jand g06362(.dina(n6617), .dinb(n6616), .dout(n6618));
  jand g06363(.dina(n6595), .dinb(n6587), .dout(n6619));
  jnot g06364(.din(n6619), .dout(n6620));
  jnot g06365(.din(n6596), .dout(n6621));
  jor  g06366(.dina(n6621), .dinb(n6384), .dout(n6622));
  jand g06367(.dina(n6622), .dinb(n6620), .dout(n6623));
  jand g06368(.dina(n6585), .dinb(n6577), .dout(n6624));
  jand g06369(.dina(n6586), .dinb(n6387), .dout(n6625));
  jor  g06370(.dina(n6625), .dinb(n6624), .dout(n6626));
  jand g06371(.dina(n6574), .dinb(n6566), .dout(n6627));
  jnot g06372(.din(n6627), .dout(n6628));
  jor  g06373(.dina(n6576), .dinb(n6391), .dout(n6629));
  jand g06374(.dina(n6629), .dinb(n6628), .dout(n6630));
  jand g06375(.dina(n6564), .dinb(n6556), .dout(n6631));
  jand g06376(.dina(n6565), .dinb(n6394), .dout(n6632));
  jor  g06377(.dina(n6632), .dinb(n6631), .dout(n6633));
  jand g06378(.dina(n6554), .dinb(n6546), .dout(n6634));
  jand g06379(.dina(n6555), .dinb(n6397), .dout(n6635));
  jor  g06380(.dina(n6635), .dinb(n6634), .dout(n6636));
  jand g06381(.dina(n6544), .dinb(n6536), .dout(n6637));
  jand g06382(.dina(n6545), .dinb(n6400), .dout(n6638));
  jor  g06383(.dina(n6638), .dinb(n6637), .dout(n6639));
  jand g06384(.dina(n6534), .dinb(n6526), .dout(n6640));
  jand g06385(.dina(n6535), .dinb(n6403), .dout(n6641));
  jor  g06386(.dina(n6641), .dinb(n6640), .dout(n6642));
  jand g06387(.dina(n6524), .dinb(n6516), .dout(n6643));
  jand g06388(.dina(n6525), .dinb(n6406), .dout(n6644));
  jor  g06389(.dina(n6644), .dinb(n6643), .dout(n6645));
  jand g06390(.dina(n6514), .dinb(n6506), .dout(n6646));
  jand g06391(.dina(n6515), .dinb(n6409), .dout(n6647));
  jor  g06392(.dina(n6647), .dinb(n6646), .dout(n6648));
  jand g06393(.dina(n6504), .dinb(n6496), .dout(n6649));
  jand g06394(.dina(n6505), .dinb(n6412), .dout(n6650));
  jor  g06395(.dina(n6650), .dinb(n6649), .dout(n6651));
  jand g06396(.dina(n6494), .dinb(n6486), .dout(n6652));
  jand g06397(.dina(n6495), .dinb(n6415), .dout(n6653));
  jor  g06398(.dina(n6653), .dinb(n6652), .dout(n6654));
  jand g06399(.dina(n6484), .dinb(n6476), .dout(n6655));
  jand g06400(.dina(n6485), .dinb(n6418), .dout(n6656));
  jor  g06401(.dina(n6656), .dinb(n6655), .dout(n6657));
  jand g06402(.dina(n6474), .dinb(n6466), .dout(n6658));
  jand g06403(.dina(n6475), .dinb(n6421), .dout(n6659));
  jor  g06404(.dina(n6659), .dinb(n6658), .dout(n6660));
  jor  g06405(.dina(n6464), .dinb(n6456), .dout(n6661));
  jand g06406(.dina(n6465), .dinb(n6426), .dout(n6662));
  jnot g06407(.din(n6662), .dout(n6663));
  jand g06408(.dina(n6663), .dinb(n6661), .dout(n6664));
  jnot g06409(.din(n6664), .dout(n6665));
  jor  g06410(.dina(n6453), .dinb(n6445), .dout(n6666));
  jand g06411(.dina(n6454), .dinb(n6430), .dout(n6667));
  jnot g06412(.din(n6667), .dout(n6668));
  jand g06413(.dina(n6668), .dinb(n6666), .dout(n6669));
  jnot g06414(.din(n6669), .dout(n6670));
  jand g06415(.dina(n6439), .dinb(b1 ), .dout(n6671));
  jor  g06416(.dina(n6438), .dinb(n6201), .dout(n6672));
  jor  g06417(.dina(n6672), .dinb(n6432), .dout(n6673));
  jnot g06418(.din(n6673), .dout(n6674));
  jand g06419(.dina(n6674), .dinb(b0 ), .dout(n6675));
  jand g06420(.dina(n6435), .dinb(n273), .dout(n6676));
  jand g06421(.dina(n6433), .dinb(b2 ), .dout(n6677));
  jor  g06422(.dina(n6677), .dinb(n6676), .dout(n6678));
  jor  g06423(.dina(n6678), .dinb(n6675), .dout(n6679));
  jor  g06424(.dina(n6679), .dinb(n6671), .dout(n6680));
  jnot g06425(.din(n6442), .dout(n6681));
  jand g06426(.dina(n6203), .dinb(a50 ), .dout(n6682));
  jand g06427(.dina(n6682), .dinb(n6681), .dout(n6683));
  jnot g06428(.din(n6683), .dout(n6684));
  jand g06429(.dina(n6684), .dinb(a50 ), .dout(n6685));
  jxor g06430(.dina(n6685), .dinb(n6680), .dout(n6686));
  jnot g06431(.din(n6686), .dout(n6687));
  jor  g06432(.dina(n6207), .dinb(n374), .dout(n6688));
  jor  g06433(.dina(n6210), .dinb(n340), .dout(n6689));
  jor  g06434(.dina(n5975), .dinb(n303), .dout(n6690));
  jand g06435(.dina(n6690), .dinb(n6689), .dout(n6691));
  jor  g06436(.dina(n6205), .dinb(n377), .dout(n6692));
  jand g06437(.dina(n6692), .dinb(n6691), .dout(n6693));
  jand g06438(.dina(n6693), .dinb(n6688), .dout(n6694));
  jxor g06439(.dina(n6694), .dinb(a47 ), .dout(n6695));
  jxor g06440(.dina(n6695), .dinb(n6687), .dout(n6696));
  jxor g06441(.dina(n6696), .dinb(n6670), .dout(n6697));
  jor  g06442(.dina(n5537), .dinb(n517), .dout(n6698));
  jor  g06443(.dina(n5534), .dinb(n469), .dout(n6699));
  jor  g06444(.dina(n5539), .dinb(n519), .dout(n6700));
  jor  g06445(.dina(n5315), .dinb(n415), .dout(n6701));
  jand g06446(.dina(n6701), .dinb(n6700), .dout(n6702));
  jand g06447(.dina(n6702), .dinb(n6699), .dout(n6703));
  jand g06448(.dina(n6703), .dinb(n6698), .dout(n6704));
  jxor g06449(.dina(n6704), .dinb(n5111), .dout(n6705));
  jxor g06450(.dina(n6705), .dinb(n6697), .dout(n6706));
  jxor g06451(.dina(n6706), .dinb(n6665), .dout(n6707));
  jor  g06452(.dina(n4902), .dinb(n702), .dout(n6708));
  jor  g06453(.dina(n4696), .dinb(n572), .dout(n6709));
  jor  g06454(.dina(n4899), .dinb(n704), .dout(n6710));
  jor  g06455(.dina(n4904), .dinb(n637), .dout(n6711));
  jand g06456(.dina(n6711), .dinb(n6710), .dout(n6712));
  jand g06457(.dina(n6712), .dinb(n6709), .dout(n6713));
  jand g06458(.dina(n6713), .dinb(n6708), .dout(n6714));
  jxor g06459(.dina(n6714), .dinb(n4505), .dout(n6715));
  jxor g06460(.dina(n6715), .dinb(n6707), .dout(n6716));
  jxor g06461(.dina(n6716), .dinb(n6660), .dout(n6717));
  jor  g06462(.dina(n4305), .dinb(n932), .dout(n6718));
  jor  g06463(.dina(n4116), .dinb(n772), .dout(n6719));
  jor  g06464(.dina(n4308), .dinb(n852), .dout(n6720));
  jor  g06465(.dina(n4303), .dinb(n934), .dout(n6721));
  jand g06466(.dina(n6721), .dinb(n6720), .dout(n6722));
  jand g06467(.dina(n6722), .dinb(n6719), .dout(n6723));
  jand g06468(.dina(n6723), .dinb(n6718), .dout(n6724));
  jxor g06469(.dina(n6724), .dinb(n3938), .dout(n6725));
  jxor g06470(.dina(n6725), .dinb(n6717), .dout(n6726));
  jxor g06471(.dina(n6726), .dinb(n6657), .dout(n6727));
  jor  g06472(.dina(n3751), .dinb(n1209), .dout(n6728));
  jor  g06473(.dina(n3574), .dinb(n1018), .dout(n6729));
  jor  g06474(.dina(n3749), .dinb(n1211), .dout(n6730));
  jor  g06475(.dina(n3754), .dinb(n1114), .dout(n6731));
  jand g06476(.dina(n6731), .dinb(n6730), .dout(n6732));
  jand g06477(.dina(n6732), .dinb(n6729), .dout(n6733));
  jand g06478(.dina(n6733), .dinb(n6728), .dout(n6734));
  jxor g06479(.dina(n6734), .dinb(n3410), .dout(n6735));
  jxor g06480(.dina(n6735), .dinb(n6727), .dout(n6736));
  jxor g06481(.dina(n6736), .dinb(n6654), .dout(n6737));
  jor  g06482(.dina(n3239), .dinb(n1525), .dout(n6738));
  jor  g06483(.dina(n3072), .dinb(n1307), .dout(n6739));
  jor  g06484(.dina(n3242), .dinb(n1416), .dout(n6740));
  jor  g06485(.dina(n3237), .dinb(n1527), .dout(n6741));
  jand g06486(.dina(n6741), .dinb(n6740), .dout(n6742));
  jand g06487(.dina(n6742), .dinb(n6739), .dout(n6743));
  jand g06488(.dina(n6743), .dinb(n6738), .dout(n6744));
  jxor g06489(.dina(n6744), .dinb(n2918), .dout(n6745));
  jxor g06490(.dina(n6745), .dinb(n6737), .dout(n6746));
  jxor g06491(.dina(n6746), .dinb(n6651), .dout(n6747));
  jor  g06492(.dina(n2764), .dinb(n1879), .dout(n6748));
  jor  g06493(.dina(n2609), .dinb(n1637), .dout(n6749));
  jor  g06494(.dina(n2761), .dinb(n1881), .dout(n6750));
  jor  g06495(.dina(n2766), .dinb(n1759), .dout(n6751));
  jand g06496(.dina(n6751), .dinb(n6750), .dout(n6752));
  jand g06497(.dina(n6752), .dinb(n6749), .dout(n6753));
  jand g06498(.dina(n6753), .dinb(n6748), .dout(n6754));
  jxor g06499(.dina(n6754), .dinb(n2468), .dout(n6755));
  jxor g06500(.dina(n6755), .dinb(n6747), .dout(n6756));
  jxor g06501(.dina(n6756), .dinb(n6648), .dout(n6757));
  jor  g06502(.dina(n2277), .dinb(n2324), .dout(n6758));
  jor  g06503(.dina(n2186), .dinb(n2007), .dout(n6759));
  jor  g06504(.dina(n2326), .dinb(n2279), .dout(n6760));
  jor  g06505(.dina(n2321), .dinb(n2142), .dout(n6761));
  jand g06506(.dina(n6761), .dinb(n6760), .dout(n6762));
  jand g06507(.dina(n6762), .dinb(n6759), .dout(n6763));
  jand g06508(.dina(n6763), .dinb(n6758), .dout(n6764));
  jxor g06509(.dina(n6764), .dinb(n2057), .dout(n6765));
  jxor g06510(.dina(n6765), .dinb(n6757), .dout(n6766));
  jxor g06511(.dina(n6766), .dinb(n6645), .dout(n6767));
  jor  g06512(.dina(n2711), .dinb(n1921), .dout(n6768));
  jor  g06513(.dina(n1806), .dinb(n2415), .dout(n6769));
  jor  g06514(.dina(n1918), .dinb(n2563), .dout(n6770));
  jor  g06515(.dina(n1923), .dinb(n2713), .dout(n6771));
  jand g06516(.dina(n6771), .dinb(n6770), .dout(n6772));
  jand g06517(.dina(n6772), .dinb(n6769), .dout(n6773));
  jand g06518(.dina(n6773), .dinb(n6768), .dout(n6774));
  jxor g06519(.dina(n6774), .dinb(n1687), .dout(n6775));
  jxor g06520(.dina(n6775), .dinb(n6767), .dout(n6776));
  jxor g06521(.dina(n6776), .dinb(n6642), .dout(n6777));
  jor  g06522(.dina(n3184), .dinb(n1569), .dout(n6778));
  jor  g06523(.dina(n1453), .dinb(n2862), .dout(n6779));
  jor  g06524(.dina(n1566), .dinb(n3023), .dout(n6780));
  jor  g06525(.dina(n1571), .dinb(n3186), .dout(n6781));
  jand g06526(.dina(n6781), .dinb(n6780), .dout(n6782));
  jand g06527(.dina(n6782), .dinb(n6779), .dout(n6783));
  jand g06528(.dina(n6783), .dinb(n6778), .dout(n6784));
  jxor g06529(.dina(n6784), .dinb(n1351), .dout(n6785));
  jxor g06530(.dina(n6785), .dinb(n6777), .dout(n6786));
  jxor g06531(.dina(n6786), .dinb(n6639), .dout(n6787));
  jor  g06532(.dina(n3696), .dinb(n1248), .dout(n6788));
  jor  g06533(.dina(n1147), .dinb(n3348), .dout(n6789));
  jor  g06534(.dina(n1251), .dinb(n3522), .dout(n6790));
  jor  g06535(.dina(n1246), .dinb(n3698), .dout(n6791));
  jand g06536(.dina(n6791), .dinb(n6790), .dout(n6792));
  jand g06537(.dina(n6792), .dinb(n6789), .dout(n6793));
  jand g06538(.dina(n6793), .dinb(n6788), .dout(n6794));
  jxor g06539(.dina(n6794), .dinb(n1061), .dout(n6795));
  jxor g06540(.dina(n6795), .dinb(n6787), .dout(n6796));
  jxor g06541(.dina(n6796), .dinb(n6636), .dout(n6797));
  jor  g06542(.dina(n4247), .dinb(n970), .dout(n6798));
  jor  g06543(.dina(n880), .dinb(n3873), .dout(n6799));
  jor  g06544(.dina(n967), .dinb(n4060), .dout(n6800));
  jor  g06545(.dina(n972), .dinb(n4249), .dout(n6801));
  jand g06546(.dina(n6801), .dinb(n6800), .dout(n6802));
  jand g06547(.dina(n6802), .dinb(n6799), .dout(n6803));
  jand g06548(.dina(n6803), .dinb(n6798), .dout(n6804));
  jxor g06549(.dina(n6804), .dinb(n810), .dout(n6805));
  jxor g06550(.dina(n6805), .dinb(n6797), .dout(n6806));
  jxor g06551(.dina(n6806), .dinb(n6633), .dout(n6807));
  jor  g06552(.dina(n4837), .dinb(n728), .dout(n6808));
  jor  g06553(.dina(n660), .dinb(n4437), .dout(n6809));
  jor  g06554(.dina(n726), .dinb(n4839), .dout(n6810));
  jor  g06555(.dina(n731), .dinb(n4637), .dout(n6811));
  jand g06556(.dina(n6811), .dinb(n6810), .dout(n6812));
  jand g06557(.dina(n6812), .dinb(n6809), .dout(n6813));
  jand g06558(.dina(n6813), .dinb(n6808), .dout(n6814));
  jxor g06559(.dina(n6814), .dinb(n606), .dout(n6815));
  jxor g06560(.dina(n6815), .dinb(n6807), .dout(n6816));
  jnot g06561(.din(n6816), .dout(n6817));
  jxor g06562(.dina(n6817), .dinb(n6630), .dout(n6818));
  jor  g06563(.dina(n5467), .dinb(n544), .dout(n6819));
  jor  g06564(.dina(n486), .dinb(n5040), .dout(n6820));
  jor  g06565(.dina(n542), .dinb(n5469), .dout(n6821));
  jor  g06566(.dina(n547), .dinb(n5253), .dout(n6822));
  jand g06567(.dina(n6822), .dinb(n6821), .dout(n6823));
  jand g06568(.dina(n6823), .dinb(n6820), .dout(n6824));
  jand g06569(.dina(n6824), .dinb(n6819), .dout(n6825));
  jxor g06570(.dina(n6825), .dinb(n446), .dout(n6826));
  jxor g06571(.dina(n6826), .dinb(n6818), .dout(n6827));
  jxor g06572(.dina(n6827), .dinb(n6626), .dout(n6828));
  jor  g06573(.dina(n6137), .dinb(n397), .dout(n6829));
  jor  g06574(.dina(n354), .dinb(n5685), .dout(n6830));
  jor  g06575(.dina(n399), .dinb(n6139), .dout(n6831));
  jor  g06576(.dina(n394), .dinb(n5911), .dout(n6832));
  jand g06577(.dina(n6832), .dinb(n6831), .dout(n6833));
  jand g06578(.dina(n6833), .dinb(n6830), .dout(n6834));
  jand g06579(.dina(n6834), .dinb(n6829), .dout(n6835));
  jxor g06580(.dina(n6835), .dinb(n364), .dout(n6836));
  jxor g06581(.dina(n6836), .dinb(n6828), .dout(n6837));
  jxor g06582(.dina(n6837), .dinb(n6623), .dout(n6838));
  jand g06583(.dina(b49 ), .dinb(b48 ), .dout(n6839));
  jand g06584(.dina(n6601), .dinb(n6600), .dout(n6840));
  jor  g06585(.dina(n6840), .dinb(n6839), .dout(n6841));
  jxor g06586(.dina(b50 ), .dinb(b49 ), .dout(n6842));
  jnot g06587(.din(n6842), .dout(n6843));
  jxor g06588(.dina(n6843), .dinb(n6841), .dout(n6844));
  jor  g06589(.dina(n6844), .dinb(n296), .dout(n6845));
  jnot g06590(.din(b50 ), .dout(n6846));
  jor  g06591(.dina(n264), .dinb(n6846), .dout(n6847));
  jor  g06592(.dina(n294), .dinb(n6605), .dout(n6848));
  jor  g06593(.dina(n280), .dinb(n6366), .dout(n6849));
  jand g06594(.dina(n6849), .dinb(n6848), .dout(n6850));
  jand g06595(.dina(n6850), .dinb(n6847), .dout(n6851));
  jand g06596(.dina(n6851), .dinb(n6845), .dout(n6852));
  jxor g06597(.dina(n6852), .dinb(n278), .dout(n6853));
  jxor g06598(.dina(n6853), .dinb(n6838), .dout(n6854));
  jxor g06599(.dina(n6854), .dinb(n6618), .dout(f50 ));
  jnot g06600(.din(n6853), .dout(n6856));
  jor  g06601(.dina(n6856), .dinb(n6838), .dout(n6857));
  jor  g06602(.dina(n6854), .dinb(n6618), .dout(n6858));
  jand g06603(.dina(n6858), .dinb(n6857), .dout(n6859));
  jand g06604(.dina(n6836), .dinb(n6828), .dout(n6860));
  jnot g06605(.din(n6860), .dout(n6861));
  jnot g06606(.din(n6837), .dout(n6862));
  jor  g06607(.dina(n6862), .dinb(n6623), .dout(n6863));
  jand g06608(.dina(n6863), .dinb(n6861), .dout(n6864));
  jand g06609(.dina(n6826), .dinb(n6818), .dout(n6865));
  jand g06610(.dina(n6827), .dinb(n6626), .dout(n6866));
  jor  g06611(.dina(n6866), .dinb(n6865), .dout(n6867));
  jand g06612(.dina(n6805), .dinb(n6797), .dout(n6868));
  jand g06613(.dina(n6806), .dinb(n6633), .dout(n6869));
  jor  g06614(.dina(n6869), .dinb(n6868), .dout(n6870));
  jand g06615(.dina(n6795), .dinb(n6787), .dout(n6871));
  jand g06616(.dina(n6796), .dinb(n6636), .dout(n6872));
  jor  g06617(.dina(n6872), .dinb(n6871), .dout(n6873));
  jand g06618(.dina(n6785), .dinb(n6777), .dout(n6874));
  jand g06619(.dina(n6786), .dinb(n6639), .dout(n6875));
  jor  g06620(.dina(n6875), .dinb(n6874), .dout(n6876));
  jand g06621(.dina(n6775), .dinb(n6767), .dout(n6877));
  jand g06622(.dina(n6776), .dinb(n6642), .dout(n6878));
  jor  g06623(.dina(n6878), .dinb(n6877), .dout(n6879));
  jand g06624(.dina(n6765), .dinb(n6757), .dout(n6880));
  jand g06625(.dina(n6766), .dinb(n6645), .dout(n6881));
  jor  g06626(.dina(n6881), .dinb(n6880), .dout(n6882));
  jand g06627(.dina(n6755), .dinb(n6747), .dout(n6883));
  jand g06628(.dina(n6756), .dinb(n6648), .dout(n6884));
  jor  g06629(.dina(n6884), .dinb(n6883), .dout(n6885));
  jand g06630(.dina(n6745), .dinb(n6737), .dout(n6886));
  jand g06631(.dina(n6746), .dinb(n6651), .dout(n6887));
  jor  g06632(.dina(n6887), .dinb(n6886), .dout(n6888));
  jand g06633(.dina(n6735), .dinb(n6727), .dout(n6889));
  jand g06634(.dina(n6736), .dinb(n6654), .dout(n6890));
  jor  g06635(.dina(n6890), .dinb(n6889), .dout(n6891));
  jand g06636(.dina(n6725), .dinb(n6717), .dout(n6892));
  jand g06637(.dina(n6726), .dinb(n6657), .dout(n6893));
  jor  g06638(.dina(n6893), .dinb(n6892), .dout(n6894));
  jand g06639(.dina(n6715), .dinb(n6707), .dout(n6895));
  jand g06640(.dina(n6716), .dinb(n6660), .dout(n6896));
  jor  g06641(.dina(n6896), .dinb(n6895), .dout(n6897));
  jand g06642(.dina(n6705), .dinb(n6697), .dout(n6898));
  jand g06643(.dina(n6706), .dinb(n6665), .dout(n6899));
  jor  g06644(.dina(n6899), .dinb(n6898), .dout(n6900));
  jor  g06645(.dina(n6695), .dinb(n6687), .dout(n6901));
  jand g06646(.dina(n6696), .dinb(n6670), .dout(n6902));
  jnot g06647(.din(n6902), .dout(n6903));
  jand g06648(.dina(n6903), .dinb(n6901), .dout(n6904));
  jnot g06649(.din(n6904), .dout(n6905));
  jor  g06650(.dina(n6684), .dinb(n6680), .dout(n6906));
  jxor g06651(.dina(a51 ), .dinb(a50 ), .dout(n6907));
  jand g06652(.dina(n6907), .dinb(b0 ), .dout(n6908));
  jnot g06653(.din(n6908), .dout(n6909));
  jxor g06654(.dina(n6909), .dinb(n6906), .dout(n6910));
  jnot g06655(.din(n6439), .dout(n6911));
  jor  g06656(.dina(n6911), .dinb(n293), .dout(n6912));
  jor  g06657(.dina(n6673), .dinb(n305), .dout(n6913));
  jnot g06658(.din(n6435), .dout(n6914));
  jor  g06659(.dina(n6914), .dinb(n301), .dout(n6915));
  jnot g06660(.din(n6433), .dout(n6916));
  jor  g06661(.dina(n6916), .dinb(n303), .dout(n6917));
  jand g06662(.dina(n6917), .dinb(n6915), .dout(n6918));
  jand g06663(.dina(n6918), .dinb(n6913), .dout(n6919));
  jand g06664(.dina(n6919), .dinb(n6912), .dout(n6920));
  jxor g06665(.dina(n6920), .dinb(n6443), .dout(n6921));
  jxor g06666(.dina(n6921), .dinb(n6910), .dout(n6922));
  jnot g06667(.din(n6922), .dout(n6923));
  jor  g06668(.dina(n6207), .dinb(n412), .dout(n6924));
  jor  g06669(.dina(n6205), .dinb(n415), .dout(n6925));
  jor  g06670(.dina(n5975), .dinb(n340), .dout(n6926));
  jand g06671(.dina(n6926), .dinb(n6925), .dout(n6927));
  jor  g06672(.dina(n6210), .dinb(n377), .dout(n6928));
  jand g06673(.dina(n6928), .dinb(n6927), .dout(n6929));
  jand g06674(.dina(n6929), .dinb(n6924), .dout(n6930));
  jxor g06675(.dina(n6930), .dinb(a47 ), .dout(n6931));
  jxor g06676(.dina(n6931), .dinb(n6923), .dout(n6932));
  jxor g06677(.dina(n6932), .dinb(n6905), .dout(n6933));
  jor  g06678(.dina(n5537), .dinb(n570), .dout(n6934));
  jor  g06679(.dina(n5315), .dinb(n469), .dout(n6935));
  jor  g06680(.dina(n5534), .dinb(n519), .dout(n6936));
  jor  g06681(.dina(n5539), .dinb(n572), .dout(n6937));
  jand g06682(.dina(n6937), .dinb(n6936), .dout(n6938));
  jand g06683(.dina(n6938), .dinb(n6935), .dout(n6939));
  jand g06684(.dina(n6939), .dinb(n6934), .dout(n6940));
  jxor g06685(.dina(n6940), .dinb(n5111), .dout(n6941));
  jxor g06686(.dina(n6941), .dinb(n6933), .dout(n6942));
  jxor g06687(.dina(n6942), .dinb(n6900), .dout(n6943));
  jor  g06688(.dina(n4902), .dinb(n770), .dout(n6944));
  jor  g06689(.dina(n4696), .dinb(n637), .dout(n6945));
  jor  g06690(.dina(n4899), .dinb(n772), .dout(n6946));
  jor  g06691(.dina(n4904), .dinb(n704), .dout(n6947));
  jand g06692(.dina(n6947), .dinb(n6946), .dout(n6948));
  jand g06693(.dina(n6948), .dinb(n6945), .dout(n6949));
  jand g06694(.dina(n6949), .dinb(n6944), .dout(n6950));
  jxor g06695(.dina(n6950), .dinb(n4505), .dout(n6951));
  jxor g06696(.dina(n6951), .dinb(n6943), .dout(n6952));
  jxor g06697(.dina(n6952), .dinb(n6897), .dout(n6953));
  jor  g06698(.dina(n4305), .dinb(n1016), .dout(n6954));
  jor  g06699(.dina(n4116), .dinb(n852), .dout(n6955));
  jor  g06700(.dina(n4308), .dinb(n934), .dout(n6956));
  jor  g06701(.dina(n4303), .dinb(n1018), .dout(n6957));
  jand g06702(.dina(n6957), .dinb(n6956), .dout(n6958));
  jand g06703(.dina(n6958), .dinb(n6955), .dout(n6959));
  jand g06704(.dina(n6959), .dinb(n6954), .dout(n6960));
  jxor g06705(.dina(n6960), .dinb(n3938), .dout(n6961));
  jxor g06706(.dina(n6961), .dinb(n6953), .dout(n6962));
  jxor g06707(.dina(n6962), .dinb(n6894), .dout(n6963));
  jor  g06708(.dina(n3751), .dinb(n1305), .dout(n6964));
  jor  g06709(.dina(n3574), .dinb(n1114), .dout(n6965));
  jor  g06710(.dina(n3754), .dinb(n1211), .dout(n6966));
  jor  g06711(.dina(n3749), .dinb(n1307), .dout(n6967));
  jand g06712(.dina(n6967), .dinb(n6966), .dout(n6968));
  jand g06713(.dina(n6968), .dinb(n6965), .dout(n6969));
  jand g06714(.dina(n6969), .dinb(n6964), .dout(n6970));
  jxor g06715(.dina(n6970), .dinb(n3410), .dout(n6971));
  jxor g06716(.dina(n6971), .dinb(n6963), .dout(n6972));
  jxor g06717(.dina(n6972), .dinb(n6891), .dout(n6973));
  jor  g06718(.dina(n3239), .dinb(n1635), .dout(n6974));
  jor  g06719(.dina(n3072), .dinb(n1416), .dout(n6975));
  jor  g06720(.dina(n3242), .dinb(n1527), .dout(n6976));
  jor  g06721(.dina(n3237), .dinb(n1637), .dout(n6977));
  jand g06722(.dina(n6977), .dinb(n6976), .dout(n6978));
  jand g06723(.dina(n6978), .dinb(n6975), .dout(n6979));
  jand g06724(.dina(n6979), .dinb(n6974), .dout(n6980));
  jxor g06725(.dina(n6980), .dinb(n2918), .dout(n6981));
  jxor g06726(.dina(n6981), .dinb(n6973), .dout(n6982));
  jxor g06727(.dina(n6982), .dinb(n6888), .dout(n6983));
  jor  g06728(.dina(n2764), .dinb(n2005), .dout(n6984));
  jor  g06729(.dina(n2609), .dinb(n1759), .dout(n6985));
  jor  g06730(.dina(n2761), .dinb(n2007), .dout(n6986));
  jor  g06731(.dina(n2766), .dinb(n1881), .dout(n6987));
  jand g06732(.dina(n6987), .dinb(n6986), .dout(n6988));
  jand g06733(.dina(n6988), .dinb(n6985), .dout(n6989));
  jand g06734(.dina(n6989), .dinb(n6984), .dout(n6990));
  jxor g06735(.dina(n6990), .dinb(n2468), .dout(n6991));
  jxor g06736(.dina(n6991), .dinb(n6983), .dout(n6992));
  jxor g06737(.dina(n6992), .dinb(n6885), .dout(n6993));
  jor  g06738(.dina(n2413), .dinb(n2324), .dout(n6994));
  jor  g06739(.dina(n2186), .dinb(n2142), .dout(n6995));
  jor  g06740(.dina(n2326), .dinb(n2415), .dout(n6996));
  jor  g06741(.dina(n2321), .dinb(n2279), .dout(n6997));
  jand g06742(.dina(n6997), .dinb(n6996), .dout(n6998));
  jand g06743(.dina(n6998), .dinb(n6995), .dout(n6999));
  jand g06744(.dina(n6999), .dinb(n6994), .dout(n7000));
  jxor g06745(.dina(n7000), .dinb(n2057), .dout(n7001));
  jxor g06746(.dina(n7001), .dinb(n6993), .dout(n7002));
  jxor g06747(.dina(n7002), .dinb(n6882), .dout(n7003));
  jor  g06748(.dina(n2860), .dinb(n1921), .dout(n7004));
  jor  g06749(.dina(n1806), .dinb(n2563), .dout(n7005));
  jor  g06750(.dina(n1918), .dinb(n2713), .dout(n7006));
  jor  g06751(.dina(n1923), .dinb(n2862), .dout(n7007));
  jand g06752(.dina(n7007), .dinb(n7006), .dout(n7008));
  jand g06753(.dina(n7008), .dinb(n7005), .dout(n7009));
  jand g06754(.dina(n7009), .dinb(n7004), .dout(n7010));
  jxor g06755(.dina(n7010), .dinb(n1687), .dout(n7011));
  jxor g06756(.dina(n7011), .dinb(n7003), .dout(n7012));
  jxor g06757(.dina(n7012), .dinb(n6879), .dout(n7013));
  jor  g06758(.dina(n3346), .dinb(n1569), .dout(n7014));
  jor  g06759(.dina(n1453), .dinb(n3023), .dout(n7015));
  jor  g06760(.dina(n1566), .dinb(n3186), .dout(n7016));
  jor  g06761(.dina(n1571), .dinb(n3348), .dout(n7017));
  jand g06762(.dina(n7017), .dinb(n7016), .dout(n7018));
  jand g06763(.dina(n7018), .dinb(n7015), .dout(n7019));
  jand g06764(.dina(n7019), .dinb(n7014), .dout(n7020));
  jxor g06765(.dina(n7020), .dinb(n1351), .dout(n7021));
  jxor g06766(.dina(n7021), .dinb(n7013), .dout(n7022));
  jxor g06767(.dina(n7022), .dinb(n6876), .dout(n7023));
  jor  g06768(.dina(n3871), .dinb(n1248), .dout(n7024));
  jor  g06769(.dina(n1147), .dinb(n3522), .dout(n7025));
  jor  g06770(.dina(n1251), .dinb(n3698), .dout(n7026));
  jor  g06771(.dina(n1246), .dinb(n3873), .dout(n7027));
  jand g06772(.dina(n7027), .dinb(n7026), .dout(n7028));
  jand g06773(.dina(n7028), .dinb(n7025), .dout(n7029));
  jand g06774(.dina(n7029), .dinb(n7024), .dout(n7030));
  jxor g06775(.dina(n7030), .dinb(n1061), .dout(n7031));
  jxor g06776(.dina(n7031), .dinb(n7023), .dout(n7032));
  jxor g06777(.dina(n7032), .dinb(n6873), .dout(n7033));
  jor  g06778(.dina(n4435), .dinb(n970), .dout(n7034));
  jor  g06779(.dina(n880), .dinb(n4060), .dout(n7035));
  jor  g06780(.dina(n967), .dinb(n4249), .dout(n7036));
  jor  g06781(.dina(n972), .dinb(n4437), .dout(n7037));
  jand g06782(.dina(n7037), .dinb(n7036), .dout(n7038));
  jand g06783(.dina(n7038), .dinb(n7035), .dout(n7039));
  jand g06784(.dina(n7039), .dinb(n7034), .dout(n7040));
  jxor g06785(.dina(n7040), .dinb(n810), .dout(n7041));
  jxor g06786(.dina(n7041), .dinb(n7033), .dout(n7042));
  jxor g06787(.dina(n7042), .dinb(n6870), .dout(n7043));
  jor  g06788(.dina(n5038), .dinb(n728), .dout(n7044));
  jor  g06789(.dina(n660), .dinb(n4637), .dout(n7045));
  jor  g06790(.dina(n731), .dinb(n4839), .dout(n7046));
  jor  g06791(.dina(n726), .dinb(n5040), .dout(n7047));
  jand g06792(.dina(n7047), .dinb(n7046), .dout(n7048));
  jand g06793(.dina(n7048), .dinb(n7045), .dout(n7049));
  jand g06794(.dina(n7049), .dinb(n7044), .dout(n7050));
  jxor g06795(.dina(n7050), .dinb(n606), .dout(n7051));
  jxor g06796(.dina(n7051), .dinb(n7043), .dout(n7052));
  jnot g06797(.din(n7052), .dout(n7053));
  jand g06798(.dina(n6815), .dinb(n6807), .dout(n7054));
  jnot g06799(.din(n7054), .dout(n7055));
  jor  g06800(.dina(n6817), .dinb(n6630), .dout(n7056));
  jand g06801(.dina(n7056), .dinb(n7055), .dout(n7057));
  jxor g06802(.dina(n7057), .dinb(n7053), .dout(n7058));
  jor  g06803(.dina(n5683), .dinb(n544), .dout(n7059));
  jor  g06804(.dina(n486), .dinb(n5253), .dout(n7060));
  jor  g06805(.dina(n542), .dinb(n5685), .dout(n7061));
  jor  g06806(.dina(n547), .dinb(n5469), .dout(n7062));
  jand g06807(.dina(n7062), .dinb(n7061), .dout(n7063));
  jand g06808(.dina(n7063), .dinb(n7060), .dout(n7064));
  jand g06809(.dina(n7064), .dinb(n7059), .dout(n7065));
  jxor g06810(.dina(n7065), .dinb(n446), .dout(n7066));
  jxor g06811(.dina(n7066), .dinb(n7058), .dout(n7067));
  jxor g06812(.dina(n7067), .dinb(n6867), .dout(n7068));
  jor  g06813(.dina(n6364), .dinb(n397), .dout(n7069));
  jor  g06814(.dina(n354), .dinb(n5911), .dout(n7070));
  jor  g06815(.dina(n394), .dinb(n6139), .dout(n7071));
  jor  g06816(.dina(n399), .dinb(n6366), .dout(n7072));
  jand g06817(.dina(n7072), .dinb(n7071), .dout(n7073));
  jand g06818(.dina(n7073), .dinb(n7070), .dout(n7074));
  jand g06819(.dina(n7074), .dinb(n7069), .dout(n7075));
  jxor g06820(.dina(n7075), .dinb(n364), .dout(n7076));
  jxor g06821(.dina(n7076), .dinb(n7068), .dout(n7077));
  jxor g06822(.dina(n7077), .dinb(n6864), .dout(n7078));
  jand g06823(.dina(b50 ), .dinb(b49 ), .dout(n7079));
  jand g06824(.dina(n6842), .dinb(n6841), .dout(n7080));
  jor  g06825(.dina(n7080), .dinb(n7079), .dout(n7081));
  jxor g06826(.dina(b51 ), .dinb(b50 ), .dout(n7082));
  jnot g06827(.din(n7082), .dout(n7083));
  jxor g06828(.dina(n7083), .dinb(n7081), .dout(n7084));
  jor  g06829(.dina(n7084), .dinb(n296), .dout(n7085));
  jnot g06830(.din(b51 ), .dout(n7086));
  jor  g06831(.dina(n264), .dinb(n7086), .dout(n7087));
  jor  g06832(.dina(n280), .dinb(n6605), .dout(n7088));
  jor  g06833(.dina(n294), .dinb(n6846), .dout(n7089));
  jand g06834(.dina(n7089), .dinb(n7088), .dout(n7090));
  jand g06835(.dina(n7090), .dinb(n7087), .dout(n7091));
  jand g06836(.dina(n7091), .dinb(n7085), .dout(n7092));
  jxor g06837(.dina(n7092), .dinb(n278), .dout(n7093));
  jxor g06838(.dina(n7093), .dinb(n7078), .dout(n7094));
  jxor g06839(.dina(n7094), .dinb(n6859), .dout(f51 ));
  jnot g06840(.din(n7093), .dout(n7096));
  jor  g06841(.dina(n7096), .dinb(n7078), .dout(n7097));
  jor  g06842(.dina(n7094), .dinb(n6859), .dout(n7098));
  jand g06843(.dina(n7098), .dinb(n7097), .dout(n7099));
  jand g06844(.dina(n7076), .dinb(n7068), .dout(n7100));
  jnot g06845(.din(n7100), .dout(n7101));
  jnot g06846(.din(n7077), .dout(n7102));
  jor  g06847(.dina(n7102), .dinb(n6864), .dout(n7103));
  jand g06848(.dina(n7103), .dinb(n7101), .dout(n7104));
  jand g06849(.dina(n7066), .dinb(n7058), .dout(n7105));
  jand g06850(.dina(n7067), .dinb(n6867), .dout(n7106));
  jor  g06851(.dina(n7106), .dinb(n7105), .dout(n7107));
  jand g06852(.dina(n7051), .dinb(n7043), .dout(n7108));
  jnot g06853(.din(n7108), .dout(n7109));
  jor  g06854(.dina(n7057), .dinb(n7053), .dout(n7110));
  jand g06855(.dina(n7110), .dinb(n7109), .dout(n7111));
  jand g06856(.dina(n7041), .dinb(n7033), .dout(n7112));
  jand g06857(.dina(n7042), .dinb(n6870), .dout(n7113));
  jor  g06858(.dina(n7113), .dinb(n7112), .dout(n7114));
  jand g06859(.dina(n7031), .dinb(n7023), .dout(n7115));
  jand g06860(.dina(n7032), .dinb(n6873), .dout(n7116));
  jor  g06861(.dina(n7116), .dinb(n7115), .dout(n7117));
  jand g06862(.dina(n7021), .dinb(n7013), .dout(n7118));
  jand g06863(.dina(n7022), .dinb(n6876), .dout(n7119));
  jor  g06864(.dina(n7119), .dinb(n7118), .dout(n7120));
  jand g06865(.dina(n7011), .dinb(n7003), .dout(n7121));
  jand g06866(.dina(n7012), .dinb(n6879), .dout(n7122));
  jor  g06867(.dina(n7122), .dinb(n7121), .dout(n7123));
  jand g06868(.dina(n7001), .dinb(n6993), .dout(n7124));
  jand g06869(.dina(n7002), .dinb(n6882), .dout(n7125));
  jor  g06870(.dina(n7125), .dinb(n7124), .dout(n7126));
  jand g06871(.dina(n6991), .dinb(n6983), .dout(n7127));
  jand g06872(.dina(n6992), .dinb(n6885), .dout(n7128));
  jor  g06873(.dina(n7128), .dinb(n7127), .dout(n7129));
  jand g06874(.dina(n6981), .dinb(n6973), .dout(n7130));
  jand g06875(.dina(n6982), .dinb(n6888), .dout(n7131));
  jor  g06876(.dina(n7131), .dinb(n7130), .dout(n7132));
  jand g06877(.dina(n6971), .dinb(n6963), .dout(n7133));
  jand g06878(.dina(n6972), .dinb(n6891), .dout(n7134));
  jor  g06879(.dina(n7134), .dinb(n7133), .dout(n7135));
  jand g06880(.dina(n6961), .dinb(n6953), .dout(n7136));
  jand g06881(.dina(n6962), .dinb(n6894), .dout(n7137));
  jor  g06882(.dina(n7137), .dinb(n7136), .dout(n7138));
  jand g06883(.dina(n6951), .dinb(n6943), .dout(n7139));
  jand g06884(.dina(n6952), .dinb(n6897), .dout(n7140));
  jor  g06885(.dina(n7140), .dinb(n7139), .dout(n7141));
  jand g06886(.dina(n6941), .dinb(n6933), .dout(n7142));
  jand g06887(.dina(n6942), .dinb(n6900), .dout(n7143));
  jor  g06888(.dina(n7143), .dinb(n7142), .dout(n7144));
  jor  g06889(.dina(n6931), .dinb(n6923), .dout(n7145));
  jand g06890(.dina(n6932), .dinb(n6905), .dout(n7146));
  jnot g06891(.din(n7146), .dout(n7147));
  jand g06892(.dina(n7147), .dinb(n7145), .dout(n7148));
  jnot g06893(.din(n7148), .dout(n7149));
  jnot g06894(.din(n6906), .dout(n7150));
  jand g06895(.dina(n6908), .dinb(n7150), .dout(n7151));
  jand g06896(.dina(n6921), .dinb(n6910), .dout(n7152));
  jor  g06897(.dina(n7152), .dinb(n7151), .dout(n7153));
  jxor g06898(.dina(a53 ), .dinb(a52 ), .dout(n7154));
  jand g06899(.dina(n7154), .dinb(n6907), .dout(n7155));
  jand g06900(.dina(n7155), .dinb(n259), .dout(n7156));
  jnot g06901(.din(n6907), .dout(n7157));
  jxor g06902(.dina(a52 ), .dinb(a51 ), .dout(n7158));
  jand g06903(.dina(n7158), .dinb(n7157), .dout(n7159));
  jand g06904(.dina(n7159), .dinb(b0 ), .dout(n7160));
  jnot g06905(.din(n7154), .dout(n7161));
  jand g06906(.dina(n7161), .dinb(n6907), .dout(n7162));
  jand g06907(.dina(n7162), .dinb(b1 ), .dout(n7163));
  jor  g06908(.dina(n7163), .dinb(n7160), .dout(n7164));
  jor  g06909(.dina(n7164), .dinb(n7156), .dout(n7165));
  jnot g06910(.din(a53 ), .dout(n7166));
  jor  g06911(.dina(n6909), .dinb(n7166), .dout(n7167));
  jxor g06912(.dina(n7167), .dinb(n7165), .dout(n7168));
  jor  g06913(.dina(n6914), .dinb(n337), .dout(n7169));
  jor  g06914(.dina(n6916), .dinb(n340), .dout(n7170));
  jor  g06915(.dina(n6673), .dinb(n293), .dout(n7171));
  jand g06916(.dina(n7171), .dinb(n7170), .dout(n7172));
  jor  g06917(.dina(n6911), .dinb(n303), .dout(n7173));
  jand g06918(.dina(n7173), .dinb(n7172), .dout(n7174));
  jand g06919(.dina(n7174), .dinb(n7169), .dout(n7175));
  jxor g06920(.dina(n7175), .dinb(a50 ), .dout(n7176));
  jxor g06921(.dina(n7176), .dinb(n7168), .dout(n7177));
  jxor g06922(.dina(n7177), .dinb(n7153), .dout(n7178));
  jnot g06923(.din(n7178), .dout(n7179));
  jor  g06924(.dina(n6207), .dinb(n466), .dout(n7180));
  jor  g06925(.dina(n6205), .dinb(n469), .dout(n7181));
  jor  g06926(.dina(n5975), .dinb(n377), .dout(n7182));
  jand g06927(.dina(n7182), .dinb(n7181), .dout(n7183));
  jor  g06928(.dina(n6210), .dinb(n415), .dout(n7184));
  jand g06929(.dina(n7184), .dinb(n7183), .dout(n7185));
  jand g06930(.dina(n7185), .dinb(n7180), .dout(n7186));
  jxor g06931(.dina(n7186), .dinb(a47 ), .dout(n7187));
  jxor g06932(.dina(n7187), .dinb(n7179), .dout(n7188));
  jxor g06933(.dina(n7188), .dinb(n7149), .dout(n7189));
  jor  g06934(.dina(n5537), .dinb(n635), .dout(n7190));
  jor  g06935(.dina(n5315), .dinb(n519), .dout(n7191));
  jor  g06936(.dina(n5539), .dinb(n637), .dout(n7192));
  jor  g06937(.dina(n5534), .dinb(n572), .dout(n7193));
  jand g06938(.dina(n7193), .dinb(n7192), .dout(n7194));
  jand g06939(.dina(n7194), .dinb(n7191), .dout(n7195));
  jand g06940(.dina(n7195), .dinb(n7190), .dout(n7196));
  jxor g06941(.dina(n7196), .dinb(n5111), .dout(n7197));
  jxor g06942(.dina(n7197), .dinb(n7189), .dout(n7198));
  jxor g06943(.dina(n7198), .dinb(n7144), .dout(n7199));
  jor  g06944(.dina(n4902), .dinb(n850), .dout(n7200));
  jor  g06945(.dina(n4696), .dinb(n704), .dout(n7201));
  jor  g06946(.dina(n4904), .dinb(n772), .dout(n7202));
  jor  g06947(.dina(n4899), .dinb(n852), .dout(n7203));
  jand g06948(.dina(n7203), .dinb(n7202), .dout(n7204));
  jand g06949(.dina(n7204), .dinb(n7201), .dout(n7205));
  jand g06950(.dina(n7205), .dinb(n7200), .dout(n7206));
  jxor g06951(.dina(n7206), .dinb(n4505), .dout(n7207));
  jxor g06952(.dina(n7207), .dinb(n7199), .dout(n7208));
  jxor g06953(.dina(n7208), .dinb(n7141), .dout(n7209));
  jor  g06954(.dina(n4305), .dinb(n1112), .dout(n7210));
  jor  g06955(.dina(n4116), .dinb(n934), .dout(n7211));
  jor  g06956(.dina(n4308), .dinb(n1018), .dout(n7212));
  jor  g06957(.dina(n4303), .dinb(n1114), .dout(n7213));
  jand g06958(.dina(n7213), .dinb(n7212), .dout(n7214));
  jand g06959(.dina(n7214), .dinb(n7211), .dout(n7215));
  jand g06960(.dina(n7215), .dinb(n7210), .dout(n7216));
  jxor g06961(.dina(n7216), .dinb(n3938), .dout(n7217));
  jxor g06962(.dina(n7217), .dinb(n7209), .dout(n7218));
  jxor g06963(.dina(n7218), .dinb(n7138), .dout(n7219));
  jor  g06964(.dina(n3751), .dinb(n1414), .dout(n7220));
  jor  g06965(.dina(n3574), .dinb(n1211), .dout(n7221));
  jor  g06966(.dina(n3749), .dinb(n1416), .dout(n7222));
  jor  g06967(.dina(n3754), .dinb(n1307), .dout(n7223));
  jand g06968(.dina(n7223), .dinb(n7222), .dout(n7224));
  jand g06969(.dina(n7224), .dinb(n7221), .dout(n7225));
  jand g06970(.dina(n7225), .dinb(n7220), .dout(n7226));
  jxor g06971(.dina(n7226), .dinb(n3410), .dout(n7227));
  jxor g06972(.dina(n7227), .dinb(n7219), .dout(n7228));
  jxor g06973(.dina(n7228), .dinb(n7135), .dout(n7229));
  jor  g06974(.dina(n3239), .dinb(n1757), .dout(n7230));
  jor  g06975(.dina(n3072), .dinb(n1527), .dout(n7231));
  jor  g06976(.dina(n3237), .dinb(n1759), .dout(n7232));
  jor  g06977(.dina(n3242), .dinb(n1637), .dout(n7233));
  jand g06978(.dina(n7233), .dinb(n7232), .dout(n7234));
  jand g06979(.dina(n7234), .dinb(n7231), .dout(n7235));
  jand g06980(.dina(n7235), .dinb(n7230), .dout(n7236));
  jxor g06981(.dina(n7236), .dinb(n2918), .dout(n7237));
  jxor g06982(.dina(n7237), .dinb(n7229), .dout(n7238));
  jxor g06983(.dina(n7238), .dinb(n7132), .dout(n7239));
  jor  g06984(.dina(n2764), .dinb(n2140), .dout(n7240));
  jor  g06985(.dina(n2609), .dinb(n1881), .dout(n7241));
  jor  g06986(.dina(n2761), .dinb(n2142), .dout(n7242));
  jor  g06987(.dina(n2766), .dinb(n2007), .dout(n7243));
  jand g06988(.dina(n7243), .dinb(n7242), .dout(n7244));
  jand g06989(.dina(n7244), .dinb(n7241), .dout(n7245));
  jand g06990(.dina(n7245), .dinb(n7240), .dout(n7246));
  jxor g06991(.dina(n7246), .dinb(n2468), .dout(n7247));
  jxor g06992(.dina(n7247), .dinb(n7239), .dout(n7248));
  jxor g06993(.dina(n7248), .dinb(n7129), .dout(n7249));
  jor  g06994(.dina(n2561), .dinb(n2324), .dout(n7250));
  jor  g06995(.dina(n2186), .dinb(n2279), .dout(n7251));
  jor  g06996(.dina(n2326), .dinb(n2563), .dout(n7252));
  jor  g06997(.dina(n2321), .dinb(n2415), .dout(n7253));
  jand g06998(.dina(n7253), .dinb(n7252), .dout(n7254));
  jand g06999(.dina(n7254), .dinb(n7251), .dout(n7255));
  jand g07000(.dina(n7255), .dinb(n7250), .dout(n7256));
  jxor g07001(.dina(n7256), .dinb(n2057), .dout(n7257));
  jxor g07002(.dina(n7257), .dinb(n7249), .dout(n7258));
  jxor g07003(.dina(n7258), .dinb(n7126), .dout(n7259));
  jor  g07004(.dina(n3021), .dinb(n1921), .dout(n7260));
  jor  g07005(.dina(n1806), .dinb(n2713), .dout(n7261));
  jor  g07006(.dina(n1923), .dinb(n3023), .dout(n7262));
  jor  g07007(.dina(n1918), .dinb(n2862), .dout(n7263));
  jand g07008(.dina(n7263), .dinb(n7262), .dout(n7264));
  jand g07009(.dina(n7264), .dinb(n7261), .dout(n7265));
  jand g07010(.dina(n7265), .dinb(n7260), .dout(n7266));
  jxor g07011(.dina(n7266), .dinb(n1687), .dout(n7267));
  jxor g07012(.dina(n7267), .dinb(n7259), .dout(n7268));
  jxor g07013(.dina(n7268), .dinb(n7123), .dout(n7269));
  jor  g07014(.dina(n3520), .dinb(n1569), .dout(n7270));
  jor  g07015(.dina(n1453), .dinb(n3186), .dout(n7271));
  jor  g07016(.dina(n1566), .dinb(n3348), .dout(n7272));
  jor  g07017(.dina(n1571), .dinb(n3522), .dout(n7273));
  jand g07018(.dina(n7273), .dinb(n7272), .dout(n7274));
  jand g07019(.dina(n7274), .dinb(n7271), .dout(n7275));
  jand g07020(.dina(n7275), .dinb(n7270), .dout(n7276));
  jxor g07021(.dina(n7276), .dinb(n1351), .dout(n7277));
  jxor g07022(.dina(n7277), .dinb(n7269), .dout(n7278));
  jxor g07023(.dina(n7278), .dinb(n7120), .dout(n7279));
  jor  g07024(.dina(n4058), .dinb(n1248), .dout(n7280));
  jor  g07025(.dina(n1147), .dinb(n3698), .dout(n7281));
  jor  g07026(.dina(n1251), .dinb(n3873), .dout(n7282));
  jor  g07027(.dina(n1246), .dinb(n4060), .dout(n7283));
  jand g07028(.dina(n7283), .dinb(n7282), .dout(n7284));
  jand g07029(.dina(n7284), .dinb(n7281), .dout(n7285));
  jand g07030(.dina(n7285), .dinb(n7280), .dout(n7286));
  jxor g07031(.dina(n7286), .dinb(n1061), .dout(n7287));
  jxor g07032(.dina(n7287), .dinb(n7279), .dout(n7288));
  jxor g07033(.dina(n7288), .dinb(n7117), .dout(n7289));
  jor  g07034(.dina(n4635), .dinb(n970), .dout(n7290));
  jor  g07035(.dina(n880), .dinb(n4249), .dout(n7291));
  jor  g07036(.dina(n972), .dinb(n4637), .dout(n7292));
  jor  g07037(.dina(n967), .dinb(n4437), .dout(n7293));
  jand g07038(.dina(n7293), .dinb(n7292), .dout(n7294));
  jand g07039(.dina(n7294), .dinb(n7291), .dout(n7295));
  jand g07040(.dina(n7295), .dinb(n7290), .dout(n7296));
  jxor g07041(.dina(n7296), .dinb(n810), .dout(n7297));
  jxor g07042(.dina(n7297), .dinb(n7289), .dout(n7298));
  jxor g07043(.dina(n7298), .dinb(n7114), .dout(n7299));
  jor  g07044(.dina(n5251), .dinb(n728), .dout(n7300));
  jor  g07045(.dina(n660), .dinb(n4839), .dout(n7301));
  jor  g07046(.dina(n731), .dinb(n5040), .dout(n7302));
  jor  g07047(.dina(n726), .dinb(n5253), .dout(n7303));
  jand g07048(.dina(n7303), .dinb(n7302), .dout(n7304));
  jand g07049(.dina(n7304), .dinb(n7301), .dout(n7305));
  jand g07050(.dina(n7305), .dinb(n7300), .dout(n7306));
  jxor g07051(.dina(n7306), .dinb(n606), .dout(n7307));
  jxor g07052(.dina(n7307), .dinb(n7299), .dout(n7308));
  jnot g07053(.din(n7308), .dout(n7309));
  jxor g07054(.dina(n7309), .dinb(n7111), .dout(n7310));
  jor  g07055(.dina(n5909), .dinb(n544), .dout(n7311));
  jor  g07056(.dina(n486), .dinb(n5469), .dout(n7312));
  jor  g07057(.dina(n547), .dinb(n5685), .dout(n7313));
  jor  g07058(.dina(n542), .dinb(n5911), .dout(n7314));
  jand g07059(.dina(n7314), .dinb(n7313), .dout(n7315));
  jand g07060(.dina(n7315), .dinb(n7312), .dout(n7316));
  jand g07061(.dina(n7316), .dinb(n7311), .dout(n7317));
  jxor g07062(.dina(n7317), .dinb(n446), .dout(n7318));
  jxor g07063(.dina(n7318), .dinb(n7310), .dout(n7319));
  jxor g07064(.dina(n7319), .dinb(n7107), .dout(n7320));
  jor  g07065(.dina(n6603), .dinb(n397), .dout(n7321));
  jor  g07066(.dina(n354), .dinb(n6139), .dout(n7322));
  jor  g07067(.dina(n394), .dinb(n6366), .dout(n7323));
  jor  g07068(.dina(n399), .dinb(n6605), .dout(n7324));
  jand g07069(.dina(n7324), .dinb(n7323), .dout(n7325));
  jand g07070(.dina(n7325), .dinb(n7322), .dout(n7326));
  jand g07071(.dina(n7326), .dinb(n7321), .dout(n7327));
  jxor g07072(.dina(n7327), .dinb(n364), .dout(n7328));
  jxor g07073(.dina(n7328), .dinb(n7320), .dout(n7329));
  jxor g07074(.dina(n7329), .dinb(n7104), .dout(n7330));
  jand g07075(.dina(b51 ), .dinb(b50 ), .dout(n7331));
  jand g07076(.dina(n7082), .dinb(n7081), .dout(n7332));
  jor  g07077(.dina(n7332), .dinb(n7331), .dout(n7333));
  jxor g07078(.dina(b52 ), .dinb(b51 ), .dout(n7334));
  jnot g07079(.din(n7334), .dout(n7335));
  jxor g07080(.dina(n7335), .dinb(n7333), .dout(n7336));
  jor  g07081(.dina(n7336), .dinb(n296), .dout(n7337));
  jnot g07082(.din(b52 ), .dout(n7338));
  jor  g07083(.dina(n264), .dinb(n7338), .dout(n7339));
  jor  g07084(.dina(n294), .dinb(n7086), .dout(n7340));
  jor  g07085(.dina(n280), .dinb(n6846), .dout(n7341));
  jand g07086(.dina(n7341), .dinb(n7340), .dout(n7342));
  jand g07087(.dina(n7342), .dinb(n7339), .dout(n7343));
  jand g07088(.dina(n7343), .dinb(n7337), .dout(n7344));
  jxor g07089(.dina(n7344), .dinb(n278), .dout(n7345));
  jxor g07090(.dina(n7345), .dinb(n7330), .dout(n7346));
  jxor g07091(.dina(n7346), .dinb(n7099), .dout(f52 ));
  jnot g07092(.din(n7345), .dout(n7348));
  jor  g07093(.dina(n7348), .dinb(n7330), .dout(n7349));
  jor  g07094(.dina(n7346), .dinb(n7099), .dout(n7350));
  jand g07095(.dina(n7350), .dinb(n7349), .dout(n7351));
  jand g07096(.dina(n7328), .dinb(n7320), .dout(n7352));
  jnot g07097(.din(n7352), .dout(n7353));
  jnot g07098(.din(n7329), .dout(n7354));
  jor  g07099(.dina(n7354), .dinb(n7104), .dout(n7355));
  jand g07100(.dina(n7355), .dinb(n7353), .dout(n7356));
  jand g07101(.dina(n7318), .dinb(n7310), .dout(n7357));
  jand g07102(.dina(n7319), .dinb(n7107), .dout(n7358));
  jor  g07103(.dina(n7358), .dinb(n7357), .dout(n7359));
  jand g07104(.dina(n7307), .dinb(n7299), .dout(n7360));
  jnot g07105(.din(n7360), .dout(n7361));
  jor  g07106(.dina(n7309), .dinb(n7111), .dout(n7362));
  jand g07107(.dina(n7362), .dinb(n7361), .dout(n7363));
  jand g07108(.dina(n7297), .dinb(n7289), .dout(n7364));
  jand g07109(.dina(n7298), .dinb(n7114), .dout(n7365));
  jor  g07110(.dina(n7365), .dinb(n7364), .dout(n7366));
  jand g07111(.dina(n7287), .dinb(n7279), .dout(n7367));
  jand g07112(.dina(n7288), .dinb(n7117), .dout(n7368));
  jor  g07113(.dina(n7368), .dinb(n7367), .dout(n7369));
  jand g07114(.dina(n7277), .dinb(n7269), .dout(n7370));
  jand g07115(.dina(n7278), .dinb(n7120), .dout(n7371));
  jor  g07116(.dina(n7371), .dinb(n7370), .dout(n7372));
  jand g07117(.dina(n7267), .dinb(n7259), .dout(n7373));
  jand g07118(.dina(n7268), .dinb(n7123), .dout(n7374));
  jor  g07119(.dina(n7374), .dinb(n7373), .dout(n7375));
  jand g07120(.dina(n7257), .dinb(n7249), .dout(n7376));
  jand g07121(.dina(n7258), .dinb(n7126), .dout(n7377));
  jor  g07122(.dina(n7377), .dinb(n7376), .dout(n7378));
  jand g07123(.dina(n7247), .dinb(n7239), .dout(n7379));
  jand g07124(.dina(n7248), .dinb(n7129), .dout(n7380));
  jor  g07125(.dina(n7380), .dinb(n7379), .dout(n7381));
  jand g07126(.dina(n7237), .dinb(n7229), .dout(n7382));
  jand g07127(.dina(n7238), .dinb(n7132), .dout(n7383));
  jor  g07128(.dina(n7383), .dinb(n7382), .dout(n7384));
  jand g07129(.dina(n7227), .dinb(n7219), .dout(n7385));
  jand g07130(.dina(n7228), .dinb(n7135), .dout(n7386));
  jor  g07131(.dina(n7386), .dinb(n7385), .dout(n7387));
  jand g07132(.dina(n7217), .dinb(n7209), .dout(n7388));
  jand g07133(.dina(n7218), .dinb(n7138), .dout(n7389));
  jor  g07134(.dina(n7389), .dinb(n7388), .dout(n7390));
  jand g07135(.dina(n7207), .dinb(n7199), .dout(n7391));
  jand g07136(.dina(n7208), .dinb(n7141), .dout(n7392));
  jor  g07137(.dina(n7392), .dinb(n7391), .dout(n7393));
  jand g07138(.dina(n7197), .dinb(n7189), .dout(n7394));
  jand g07139(.dina(n7198), .dinb(n7144), .dout(n7395));
  jor  g07140(.dina(n7395), .dinb(n7394), .dout(n7396));
  jor  g07141(.dina(n7187), .dinb(n7179), .dout(n7397));
  jand g07142(.dina(n7188), .dinb(n7149), .dout(n7398));
  jnot g07143(.din(n7398), .dout(n7399));
  jand g07144(.dina(n7399), .dinb(n7397), .dout(n7400));
  jnot g07145(.din(n7400), .dout(n7401));
  jor  g07146(.dina(n6207), .dinb(n517), .dout(n7402));
  jor  g07147(.dina(n6205), .dinb(n519), .dout(n7403));
  jor  g07148(.dina(n6210), .dinb(n469), .dout(n7404));
  jor  g07149(.dina(n5975), .dinb(n415), .dout(n7405));
  jand g07150(.dina(n7405), .dinb(n7404), .dout(n7406));
  jand g07151(.dina(n7406), .dinb(n7403), .dout(n7407));
  jand g07152(.dina(n7407), .dinb(n7402), .dout(n7408));
  jxor g07153(.dina(n7408), .dinb(n5759), .dout(n7409));
  jor  g07154(.dina(n7176), .dinb(n7168), .dout(n7410));
  jand g07155(.dina(n7177), .dinb(n7153), .dout(n7411));
  jnot g07156(.din(n7411), .dout(n7412));
  jand g07157(.dina(n7412), .dinb(n7410), .dout(n7413));
  jor  g07158(.dina(n7158), .dinb(n6907), .dout(n7414));
  jor  g07159(.dina(n7414), .dinb(n7161), .dout(n7415));
  jnot g07160(.din(n7415), .dout(n7416));
  jand g07161(.dina(n7416), .dinb(b0 ), .dout(n7417));
  jand g07162(.dina(n7162), .dinb(b2 ), .dout(n7418));
  jor  g07163(.dina(n7418), .dinb(n7417), .dout(n7419));
  jand g07164(.dina(n7155), .dinb(n273), .dout(n7420));
  jand g07165(.dina(n7159), .dinb(b1 ), .dout(n7421));
  jor  g07166(.dina(n7421), .dinb(n7420), .dout(n7422));
  jor  g07167(.dina(n7422), .dinb(n7419), .dout(n7423));
  jnot g07168(.din(n7165), .dout(n7424));
  jand g07169(.dina(n6909), .dinb(a53 ), .dout(n7425));
  jand g07170(.dina(n7425), .dinb(n7424), .dout(n7426));
  jnot g07171(.din(n7426), .dout(n7427));
  jand g07172(.dina(n7427), .dinb(a53 ), .dout(n7428));
  jxor g07173(.dina(n7428), .dinb(n7423), .dout(n7429));
  jor  g07174(.dina(n6914), .dinb(n374), .dout(n7430));
  jor  g07175(.dina(n6911), .dinb(n340), .dout(n7431));
  jor  g07176(.dina(n6673), .dinb(n303), .dout(n7432));
  jand g07177(.dina(n7432), .dinb(n7431), .dout(n7433));
  jor  g07178(.dina(n6916), .dinb(n377), .dout(n7434));
  jand g07179(.dina(n7434), .dinb(n7433), .dout(n7435));
  jand g07180(.dina(n7435), .dinb(n7430), .dout(n7436));
  jxor g07181(.dina(n7436), .dinb(a50 ), .dout(n7437));
  jxor g07182(.dina(n7437), .dinb(n7429), .dout(n7438));
  jxor g07183(.dina(n7438), .dinb(n7413), .dout(n7439));
  jxor g07184(.dina(n7439), .dinb(n7409), .dout(n7440));
  jxor g07185(.dina(n7440), .dinb(n7401), .dout(n7441));
  jor  g07186(.dina(n5537), .dinb(n702), .dout(n7442));
  jor  g07187(.dina(n5315), .dinb(n572), .dout(n7443));
  jor  g07188(.dina(n5539), .dinb(n704), .dout(n7444));
  jor  g07189(.dina(n5534), .dinb(n637), .dout(n7445));
  jand g07190(.dina(n7445), .dinb(n7444), .dout(n7446));
  jand g07191(.dina(n7446), .dinb(n7443), .dout(n7447));
  jand g07192(.dina(n7447), .dinb(n7442), .dout(n7448));
  jxor g07193(.dina(n7448), .dinb(n5111), .dout(n7449));
  jxor g07194(.dina(n7449), .dinb(n7441), .dout(n7450));
  jxor g07195(.dina(n7450), .dinb(n7396), .dout(n7451));
  jor  g07196(.dina(n4902), .dinb(n932), .dout(n7452));
  jor  g07197(.dina(n4696), .dinb(n772), .dout(n7453));
  jor  g07198(.dina(n4899), .dinb(n934), .dout(n7454));
  jor  g07199(.dina(n4904), .dinb(n852), .dout(n7455));
  jand g07200(.dina(n7455), .dinb(n7454), .dout(n7456));
  jand g07201(.dina(n7456), .dinb(n7453), .dout(n7457));
  jand g07202(.dina(n7457), .dinb(n7452), .dout(n7458));
  jxor g07203(.dina(n7458), .dinb(n4505), .dout(n7459));
  jxor g07204(.dina(n7459), .dinb(n7451), .dout(n7460));
  jxor g07205(.dina(n7460), .dinb(n7393), .dout(n7461));
  jor  g07206(.dina(n4305), .dinb(n1209), .dout(n7462));
  jor  g07207(.dina(n4116), .dinb(n1018), .dout(n7463));
  jor  g07208(.dina(n4308), .dinb(n1114), .dout(n7464));
  jor  g07209(.dina(n4303), .dinb(n1211), .dout(n7465));
  jand g07210(.dina(n7465), .dinb(n7464), .dout(n7466));
  jand g07211(.dina(n7466), .dinb(n7463), .dout(n7467));
  jand g07212(.dina(n7467), .dinb(n7462), .dout(n7468));
  jxor g07213(.dina(n7468), .dinb(n3938), .dout(n7469));
  jxor g07214(.dina(n7469), .dinb(n7461), .dout(n7470));
  jxor g07215(.dina(n7470), .dinb(n7390), .dout(n7471));
  jor  g07216(.dina(n3751), .dinb(n1525), .dout(n7472));
  jor  g07217(.dina(n3574), .dinb(n1307), .dout(n7473));
  jor  g07218(.dina(n3749), .dinb(n1527), .dout(n7474));
  jor  g07219(.dina(n3754), .dinb(n1416), .dout(n7475));
  jand g07220(.dina(n7475), .dinb(n7474), .dout(n7476));
  jand g07221(.dina(n7476), .dinb(n7473), .dout(n7477));
  jand g07222(.dina(n7477), .dinb(n7472), .dout(n7478));
  jxor g07223(.dina(n7478), .dinb(n3410), .dout(n7479));
  jxor g07224(.dina(n7479), .dinb(n7471), .dout(n7480));
  jxor g07225(.dina(n7480), .dinb(n7387), .dout(n7481));
  jor  g07226(.dina(n3239), .dinb(n1879), .dout(n7482));
  jor  g07227(.dina(n3072), .dinb(n1637), .dout(n7483));
  jor  g07228(.dina(n3242), .dinb(n1759), .dout(n7484));
  jor  g07229(.dina(n3237), .dinb(n1881), .dout(n7485));
  jand g07230(.dina(n7485), .dinb(n7484), .dout(n7486));
  jand g07231(.dina(n7486), .dinb(n7483), .dout(n7487));
  jand g07232(.dina(n7487), .dinb(n7482), .dout(n7488));
  jxor g07233(.dina(n7488), .dinb(n2918), .dout(n7489));
  jxor g07234(.dina(n7489), .dinb(n7481), .dout(n7490));
  jxor g07235(.dina(n7490), .dinb(n7384), .dout(n7491));
  jor  g07236(.dina(n2764), .dinb(n2277), .dout(n7492));
  jor  g07237(.dina(n2609), .dinb(n2007), .dout(n7493));
  jor  g07238(.dina(n2761), .dinb(n2279), .dout(n7494));
  jor  g07239(.dina(n2766), .dinb(n2142), .dout(n7495));
  jand g07240(.dina(n7495), .dinb(n7494), .dout(n7496));
  jand g07241(.dina(n7496), .dinb(n7493), .dout(n7497));
  jand g07242(.dina(n7497), .dinb(n7492), .dout(n7498));
  jxor g07243(.dina(n7498), .dinb(n2468), .dout(n7499));
  jxor g07244(.dina(n7499), .dinb(n7491), .dout(n7500));
  jxor g07245(.dina(n7500), .dinb(n7381), .dout(n7501));
  jor  g07246(.dina(n2711), .dinb(n2324), .dout(n7502));
  jor  g07247(.dina(n2186), .dinb(n2415), .dout(n7503));
  jor  g07248(.dina(n2326), .dinb(n2713), .dout(n7504));
  jor  g07249(.dina(n2321), .dinb(n2563), .dout(n7505));
  jand g07250(.dina(n7505), .dinb(n7504), .dout(n7506));
  jand g07251(.dina(n7506), .dinb(n7503), .dout(n7507));
  jand g07252(.dina(n7507), .dinb(n7502), .dout(n7508));
  jxor g07253(.dina(n7508), .dinb(n2057), .dout(n7509));
  jxor g07254(.dina(n7509), .dinb(n7501), .dout(n7510));
  jxor g07255(.dina(n7510), .dinb(n7378), .dout(n7511));
  jor  g07256(.dina(n3184), .dinb(n1921), .dout(n7512));
  jor  g07257(.dina(n1806), .dinb(n2862), .dout(n7513));
  jor  g07258(.dina(n1923), .dinb(n3186), .dout(n7514));
  jor  g07259(.dina(n1918), .dinb(n3023), .dout(n7515));
  jand g07260(.dina(n7515), .dinb(n7514), .dout(n7516));
  jand g07261(.dina(n7516), .dinb(n7513), .dout(n7517));
  jand g07262(.dina(n7517), .dinb(n7512), .dout(n7518));
  jxor g07263(.dina(n7518), .dinb(n1687), .dout(n7519));
  jxor g07264(.dina(n7519), .dinb(n7511), .dout(n7520));
  jxor g07265(.dina(n7520), .dinb(n7375), .dout(n7521));
  jor  g07266(.dina(n3696), .dinb(n1569), .dout(n7522));
  jor  g07267(.dina(n1453), .dinb(n3348), .dout(n7523));
  jor  g07268(.dina(n1566), .dinb(n3522), .dout(n7524));
  jor  g07269(.dina(n1571), .dinb(n3698), .dout(n7525));
  jand g07270(.dina(n7525), .dinb(n7524), .dout(n7526));
  jand g07271(.dina(n7526), .dinb(n7523), .dout(n7527));
  jand g07272(.dina(n7527), .dinb(n7522), .dout(n7528));
  jxor g07273(.dina(n7528), .dinb(n1351), .dout(n7529));
  jxor g07274(.dina(n7529), .dinb(n7521), .dout(n7530));
  jxor g07275(.dina(n7530), .dinb(n7372), .dout(n7531));
  jor  g07276(.dina(n4247), .dinb(n1248), .dout(n7532));
  jor  g07277(.dina(n1147), .dinb(n3873), .dout(n7533));
  jor  g07278(.dina(n1246), .dinb(n4249), .dout(n7534));
  jor  g07279(.dina(n1251), .dinb(n4060), .dout(n7535));
  jand g07280(.dina(n7535), .dinb(n7534), .dout(n7536));
  jand g07281(.dina(n7536), .dinb(n7533), .dout(n7537));
  jand g07282(.dina(n7537), .dinb(n7532), .dout(n7538));
  jxor g07283(.dina(n7538), .dinb(n1061), .dout(n7539));
  jxor g07284(.dina(n7539), .dinb(n7531), .dout(n7540));
  jxor g07285(.dina(n7540), .dinb(n7369), .dout(n7541));
  jor  g07286(.dina(n4837), .dinb(n970), .dout(n7542));
  jor  g07287(.dina(n880), .dinb(n4437), .dout(n7543));
  jor  g07288(.dina(n967), .dinb(n4637), .dout(n7544));
  jor  g07289(.dina(n972), .dinb(n4839), .dout(n7545));
  jand g07290(.dina(n7545), .dinb(n7544), .dout(n7546));
  jand g07291(.dina(n7546), .dinb(n7543), .dout(n7547));
  jand g07292(.dina(n7547), .dinb(n7542), .dout(n7548));
  jxor g07293(.dina(n7548), .dinb(n810), .dout(n7549));
  jxor g07294(.dina(n7549), .dinb(n7541), .dout(n7550));
  jxor g07295(.dina(n7550), .dinb(n7366), .dout(n7551));
  jor  g07296(.dina(n5467), .dinb(n728), .dout(n7552));
  jor  g07297(.dina(n660), .dinb(n5040), .dout(n7553));
  jor  g07298(.dina(n726), .dinb(n5469), .dout(n7554));
  jor  g07299(.dina(n731), .dinb(n5253), .dout(n7555));
  jand g07300(.dina(n7555), .dinb(n7554), .dout(n7556));
  jand g07301(.dina(n7556), .dinb(n7553), .dout(n7557));
  jand g07302(.dina(n7557), .dinb(n7552), .dout(n7558));
  jxor g07303(.dina(n7558), .dinb(n606), .dout(n7559));
  jxor g07304(.dina(n7559), .dinb(n7551), .dout(n7560));
  jnot g07305(.din(n7560), .dout(n7561));
  jxor g07306(.dina(n7561), .dinb(n7363), .dout(n7562));
  jor  g07307(.dina(n6137), .dinb(n544), .dout(n7563));
  jor  g07308(.dina(n486), .dinb(n5685), .dout(n7564));
  jor  g07309(.dina(n547), .dinb(n5911), .dout(n7565));
  jor  g07310(.dina(n542), .dinb(n6139), .dout(n7566));
  jand g07311(.dina(n7566), .dinb(n7565), .dout(n7567));
  jand g07312(.dina(n7567), .dinb(n7564), .dout(n7568));
  jand g07313(.dina(n7568), .dinb(n7563), .dout(n7569));
  jxor g07314(.dina(n7569), .dinb(n446), .dout(n7570));
  jxor g07315(.dina(n7570), .dinb(n7562), .dout(n7571));
  jxor g07316(.dina(n7571), .dinb(n7359), .dout(n7572));
  jor  g07317(.dina(n6844), .dinb(n397), .dout(n7573));
  jor  g07318(.dina(n354), .dinb(n6366), .dout(n7574));
  jor  g07319(.dina(n394), .dinb(n6605), .dout(n7575));
  jor  g07320(.dina(n399), .dinb(n6846), .dout(n7576));
  jand g07321(.dina(n7576), .dinb(n7575), .dout(n7577));
  jand g07322(.dina(n7577), .dinb(n7574), .dout(n7578));
  jand g07323(.dina(n7578), .dinb(n7573), .dout(n7579));
  jxor g07324(.dina(n7579), .dinb(n364), .dout(n7580));
  jxor g07325(.dina(n7580), .dinb(n7572), .dout(n7581));
  jxor g07326(.dina(n7581), .dinb(n7356), .dout(n7582));
  jand g07327(.dina(b52 ), .dinb(b51 ), .dout(n7583));
  jand g07328(.dina(n7334), .dinb(n7333), .dout(n7584));
  jor  g07329(.dina(n7584), .dinb(n7583), .dout(n7585));
  jxor g07330(.dina(b53 ), .dinb(b52 ), .dout(n7586));
  jnot g07331(.din(n7586), .dout(n7587));
  jxor g07332(.dina(n7587), .dinb(n7585), .dout(n7588));
  jor  g07333(.dina(n7588), .dinb(n296), .dout(n7589));
  jnot g07334(.din(b53 ), .dout(n7590));
  jor  g07335(.dina(n264), .dinb(n7590), .dout(n7591));
  jor  g07336(.dina(n294), .dinb(n7338), .dout(n7592));
  jor  g07337(.dina(n280), .dinb(n7086), .dout(n7593));
  jand g07338(.dina(n7593), .dinb(n7592), .dout(n7594));
  jand g07339(.dina(n7594), .dinb(n7591), .dout(n7595));
  jand g07340(.dina(n7595), .dinb(n7589), .dout(n7596));
  jxor g07341(.dina(n7596), .dinb(n278), .dout(n7597));
  jxor g07342(.dina(n7597), .dinb(n7582), .dout(n7598));
  jxor g07343(.dina(n7598), .dinb(n7351), .dout(f53 ));
  jnot g07344(.din(n7597), .dout(n7600));
  jor  g07345(.dina(n7600), .dinb(n7582), .dout(n7601));
  jor  g07346(.dina(n7598), .dinb(n7351), .dout(n7602));
  jand g07347(.dina(n7602), .dinb(n7601), .dout(n7603));
  jand g07348(.dina(n7580), .dinb(n7572), .dout(n7604));
  jnot g07349(.din(n7604), .dout(n7605));
  jnot g07350(.din(n7581), .dout(n7606));
  jor  g07351(.dina(n7606), .dinb(n7356), .dout(n7607));
  jand g07352(.dina(n7607), .dinb(n7605), .dout(n7608));
  jand g07353(.dina(n7570), .dinb(n7562), .dout(n7609));
  jand g07354(.dina(n7571), .dinb(n7359), .dout(n7610));
  jor  g07355(.dina(n7610), .dinb(n7609), .dout(n7611));
  jand g07356(.dina(n7559), .dinb(n7551), .dout(n7612));
  jnot g07357(.din(n7612), .dout(n7613));
  jor  g07358(.dina(n7561), .dinb(n7363), .dout(n7614));
  jand g07359(.dina(n7614), .dinb(n7613), .dout(n7615));
  jand g07360(.dina(n7549), .dinb(n7541), .dout(n7616));
  jand g07361(.dina(n7550), .dinb(n7366), .dout(n7617));
  jor  g07362(.dina(n7617), .dinb(n7616), .dout(n7618));
  jand g07363(.dina(n7539), .dinb(n7531), .dout(n7619));
  jand g07364(.dina(n7540), .dinb(n7369), .dout(n7620));
  jor  g07365(.dina(n7620), .dinb(n7619), .dout(n7621));
  jand g07366(.dina(n7529), .dinb(n7521), .dout(n7622));
  jand g07367(.dina(n7530), .dinb(n7372), .dout(n7623));
  jor  g07368(.dina(n7623), .dinb(n7622), .dout(n7624));
  jand g07369(.dina(n7519), .dinb(n7511), .dout(n7625));
  jand g07370(.dina(n7520), .dinb(n7375), .dout(n7626));
  jor  g07371(.dina(n7626), .dinb(n7625), .dout(n7627));
  jand g07372(.dina(n7509), .dinb(n7501), .dout(n7628));
  jand g07373(.dina(n7510), .dinb(n7378), .dout(n7629));
  jor  g07374(.dina(n7629), .dinb(n7628), .dout(n7630));
  jand g07375(.dina(n7499), .dinb(n7491), .dout(n7631));
  jand g07376(.dina(n7500), .dinb(n7381), .dout(n7632));
  jor  g07377(.dina(n7632), .dinb(n7631), .dout(n7633));
  jand g07378(.dina(n7489), .dinb(n7481), .dout(n7634));
  jand g07379(.dina(n7490), .dinb(n7384), .dout(n7635));
  jor  g07380(.dina(n7635), .dinb(n7634), .dout(n7636));
  jand g07381(.dina(n7479), .dinb(n7471), .dout(n7637));
  jand g07382(.dina(n7480), .dinb(n7387), .dout(n7638));
  jor  g07383(.dina(n7638), .dinb(n7637), .dout(n7639));
  jand g07384(.dina(n7469), .dinb(n7461), .dout(n7640));
  jand g07385(.dina(n7470), .dinb(n7390), .dout(n7641));
  jor  g07386(.dina(n7641), .dinb(n7640), .dout(n7642));
  jand g07387(.dina(n7459), .dinb(n7451), .dout(n7643));
  jand g07388(.dina(n7460), .dinb(n7393), .dout(n7644));
  jor  g07389(.dina(n7644), .dinb(n7643), .dout(n7645));
  jand g07390(.dina(n7449), .dinb(n7441), .dout(n7646));
  jand g07391(.dina(n7450), .dinb(n7396), .dout(n7647));
  jor  g07392(.dina(n7647), .dinb(n7646), .dout(n7648));
  jand g07393(.dina(n7439), .dinb(n7409), .dout(n7649));
  jand g07394(.dina(n7440), .dinb(n7401), .dout(n7650));
  jor  g07395(.dina(n7650), .dinb(n7649), .dout(n7651));
  jor  g07396(.dina(n7427), .dinb(n7423), .dout(n7652));
  jxor g07397(.dina(a54 ), .dinb(a53 ), .dout(n7653));
  jand g07398(.dina(n7653), .dinb(b0 ), .dout(n7654));
  jnot g07399(.din(n7654), .dout(n7655));
  jxor g07400(.dina(n7655), .dinb(n7652), .dout(n7656));
  jnot g07401(.din(n7159), .dout(n7657));
  jor  g07402(.dina(n7657), .dinb(n293), .dout(n7658));
  jor  g07403(.dina(n7415), .dinb(n305), .dout(n7659));
  jnot g07404(.din(n7155), .dout(n7660));
  jor  g07405(.dina(n7660), .dinb(n301), .dout(n7661));
  jnot g07406(.din(n7162), .dout(n7662));
  jor  g07407(.dina(n7662), .dinb(n303), .dout(n7663));
  jand g07408(.dina(n7663), .dinb(n7661), .dout(n7664));
  jand g07409(.dina(n7664), .dinb(n7659), .dout(n7665));
  jand g07410(.dina(n7665), .dinb(n7658), .dout(n7666));
  jxor g07411(.dina(n7666), .dinb(n7166), .dout(n7667));
  jxor g07412(.dina(n7667), .dinb(n7656), .dout(n7668));
  jnot g07413(.din(n7668), .dout(n7669));
  jor  g07414(.dina(n6914), .dinb(n412), .dout(n7670));
  jor  g07415(.dina(n6916), .dinb(n415), .dout(n7671));
  jor  g07416(.dina(n6673), .dinb(n340), .dout(n7672));
  jand g07417(.dina(n7672), .dinb(n7671), .dout(n7673));
  jor  g07418(.dina(n6911), .dinb(n377), .dout(n7674));
  jand g07419(.dina(n7674), .dinb(n7673), .dout(n7675));
  jand g07420(.dina(n7675), .dinb(n7670), .dout(n7676));
  jxor g07421(.dina(n7676), .dinb(a50 ), .dout(n7677));
  jxor g07422(.dina(n7677), .dinb(n7669), .dout(n7678));
  jnot g07423(.din(n7429), .dout(n7679));
  jand g07424(.dina(n7437), .dinb(n7679), .dout(n7680));
  jnot g07425(.din(n7680), .dout(n7681));
  jnot g07426(.din(n7413), .dout(n7682));
  jnot g07427(.din(n7437), .dout(n7683));
  jand g07428(.dina(n7683), .dinb(n7429), .dout(n7684));
  jor  g07429(.dina(n7684), .dinb(n7682), .dout(n7685));
  jand g07430(.dina(n7685), .dinb(n7681), .dout(n7686));
  jxor g07431(.dina(n7686), .dinb(n7678), .dout(n7687));
  jor  g07432(.dina(n6207), .dinb(n570), .dout(n7688));
  jor  g07433(.dina(n5975), .dinb(n469), .dout(n7689));
  jor  g07434(.dina(n6205), .dinb(n572), .dout(n7690));
  jor  g07435(.dina(n6210), .dinb(n519), .dout(n7691));
  jand g07436(.dina(n7691), .dinb(n7690), .dout(n7692));
  jand g07437(.dina(n7692), .dinb(n7689), .dout(n7693));
  jand g07438(.dina(n7693), .dinb(n7688), .dout(n7694));
  jxor g07439(.dina(n7694), .dinb(n5759), .dout(n7695));
  jxor g07440(.dina(n7695), .dinb(n7687), .dout(n7696));
  jxor g07441(.dina(n7696), .dinb(n7651), .dout(n7697));
  jor  g07442(.dina(n5537), .dinb(n770), .dout(n7698));
  jor  g07443(.dina(n5315), .dinb(n637), .dout(n7699));
  jor  g07444(.dina(n5534), .dinb(n704), .dout(n7700));
  jor  g07445(.dina(n5539), .dinb(n772), .dout(n7701));
  jand g07446(.dina(n7701), .dinb(n7700), .dout(n7702));
  jand g07447(.dina(n7702), .dinb(n7699), .dout(n7703));
  jand g07448(.dina(n7703), .dinb(n7698), .dout(n7704));
  jxor g07449(.dina(n7704), .dinb(n5111), .dout(n7705));
  jxor g07450(.dina(n7705), .dinb(n7697), .dout(n7706));
  jxor g07451(.dina(n7706), .dinb(n7648), .dout(n7707));
  jor  g07452(.dina(n4902), .dinb(n1016), .dout(n7708));
  jor  g07453(.dina(n4696), .dinb(n852), .dout(n7709));
  jor  g07454(.dina(n4899), .dinb(n1018), .dout(n7710));
  jor  g07455(.dina(n4904), .dinb(n934), .dout(n7711));
  jand g07456(.dina(n7711), .dinb(n7710), .dout(n7712));
  jand g07457(.dina(n7712), .dinb(n7709), .dout(n7713));
  jand g07458(.dina(n7713), .dinb(n7708), .dout(n7714));
  jxor g07459(.dina(n7714), .dinb(n4505), .dout(n7715));
  jxor g07460(.dina(n7715), .dinb(n7707), .dout(n7716));
  jxor g07461(.dina(n7716), .dinb(n7645), .dout(n7717));
  jor  g07462(.dina(n4305), .dinb(n1305), .dout(n7718));
  jor  g07463(.dina(n4116), .dinb(n1114), .dout(n7719));
  jor  g07464(.dina(n4303), .dinb(n1307), .dout(n7720));
  jor  g07465(.dina(n4308), .dinb(n1211), .dout(n7721));
  jand g07466(.dina(n7721), .dinb(n7720), .dout(n7722));
  jand g07467(.dina(n7722), .dinb(n7719), .dout(n7723));
  jand g07468(.dina(n7723), .dinb(n7718), .dout(n7724));
  jxor g07469(.dina(n7724), .dinb(n3938), .dout(n7725));
  jxor g07470(.dina(n7725), .dinb(n7717), .dout(n7726));
  jxor g07471(.dina(n7726), .dinb(n7642), .dout(n7727));
  jor  g07472(.dina(n3751), .dinb(n1635), .dout(n7728));
  jor  g07473(.dina(n3574), .dinb(n1416), .dout(n7729));
  jor  g07474(.dina(n3754), .dinb(n1527), .dout(n7730));
  jor  g07475(.dina(n3749), .dinb(n1637), .dout(n7731));
  jand g07476(.dina(n7731), .dinb(n7730), .dout(n7732));
  jand g07477(.dina(n7732), .dinb(n7729), .dout(n7733));
  jand g07478(.dina(n7733), .dinb(n7728), .dout(n7734));
  jxor g07479(.dina(n7734), .dinb(n3410), .dout(n7735));
  jxor g07480(.dina(n7735), .dinb(n7727), .dout(n7736));
  jxor g07481(.dina(n7736), .dinb(n7639), .dout(n7737));
  jor  g07482(.dina(n3239), .dinb(n2005), .dout(n7738));
  jor  g07483(.dina(n3072), .dinb(n1759), .dout(n7739));
  jor  g07484(.dina(n3237), .dinb(n2007), .dout(n7740));
  jor  g07485(.dina(n3242), .dinb(n1881), .dout(n7741));
  jand g07486(.dina(n7741), .dinb(n7740), .dout(n7742));
  jand g07487(.dina(n7742), .dinb(n7739), .dout(n7743));
  jand g07488(.dina(n7743), .dinb(n7738), .dout(n7744));
  jxor g07489(.dina(n7744), .dinb(n2918), .dout(n7745));
  jxor g07490(.dina(n7745), .dinb(n7737), .dout(n7746));
  jxor g07491(.dina(n7746), .dinb(n7636), .dout(n7747));
  jor  g07492(.dina(n2764), .dinb(n2413), .dout(n7748));
  jor  g07493(.dina(n2609), .dinb(n2142), .dout(n7749));
  jor  g07494(.dina(n2761), .dinb(n2415), .dout(n7750));
  jor  g07495(.dina(n2766), .dinb(n2279), .dout(n7751));
  jand g07496(.dina(n7751), .dinb(n7750), .dout(n7752));
  jand g07497(.dina(n7752), .dinb(n7749), .dout(n7753));
  jand g07498(.dina(n7753), .dinb(n7748), .dout(n7754));
  jxor g07499(.dina(n7754), .dinb(n2468), .dout(n7755));
  jxor g07500(.dina(n7755), .dinb(n7747), .dout(n7756));
  jxor g07501(.dina(n7756), .dinb(n7633), .dout(n7757));
  jor  g07502(.dina(n2860), .dinb(n2324), .dout(n7758));
  jor  g07503(.dina(n2186), .dinb(n2563), .dout(n7759));
  jor  g07504(.dina(n2321), .dinb(n2713), .dout(n7760));
  jor  g07505(.dina(n2326), .dinb(n2862), .dout(n7761));
  jand g07506(.dina(n7761), .dinb(n7760), .dout(n7762));
  jand g07507(.dina(n7762), .dinb(n7759), .dout(n7763));
  jand g07508(.dina(n7763), .dinb(n7758), .dout(n7764));
  jxor g07509(.dina(n7764), .dinb(n2057), .dout(n7765));
  jxor g07510(.dina(n7765), .dinb(n7757), .dout(n7766));
  jxor g07511(.dina(n7766), .dinb(n7630), .dout(n7767));
  jor  g07512(.dina(n3346), .dinb(n1921), .dout(n7768));
  jor  g07513(.dina(n1806), .dinb(n3023), .dout(n7769));
  jor  g07514(.dina(n1923), .dinb(n3348), .dout(n7770));
  jor  g07515(.dina(n1918), .dinb(n3186), .dout(n7771));
  jand g07516(.dina(n7771), .dinb(n7770), .dout(n7772));
  jand g07517(.dina(n7772), .dinb(n7769), .dout(n7773));
  jand g07518(.dina(n7773), .dinb(n7768), .dout(n7774));
  jxor g07519(.dina(n7774), .dinb(n1687), .dout(n7775));
  jxor g07520(.dina(n7775), .dinb(n7767), .dout(n7776));
  jxor g07521(.dina(n7776), .dinb(n7627), .dout(n7777));
  jor  g07522(.dina(n3871), .dinb(n1569), .dout(n7778));
  jor  g07523(.dina(n1453), .dinb(n3522), .dout(n7779));
  jor  g07524(.dina(n1566), .dinb(n3698), .dout(n7780));
  jor  g07525(.dina(n1571), .dinb(n3873), .dout(n7781));
  jand g07526(.dina(n7781), .dinb(n7780), .dout(n7782));
  jand g07527(.dina(n7782), .dinb(n7779), .dout(n7783));
  jand g07528(.dina(n7783), .dinb(n7778), .dout(n7784));
  jxor g07529(.dina(n7784), .dinb(n1351), .dout(n7785));
  jxor g07530(.dina(n7785), .dinb(n7777), .dout(n7786));
  jxor g07531(.dina(n7786), .dinb(n7624), .dout(n7787));
  jor  g07532(.dina(n4435), .dinb(n1248), .dout(n7788));
  jor  g07533(.dina(n1147), .dinb(n4060), .dout(n7789));
  jor  g07534(.dina(n1251), .dinb(n4249), .dout(n7790));
  jor  g07535(.dina(n1246), .dinb(n4437), .dout(n7791));
  jand g07536(.dina(n7791), .dinb(n7790), .dout(n7792));
  jand g07537(.dina(n7792), .dinb(n7789), .dout(n7793));
  jand g07538(.dina(n7793), .dinb(n7788), .dout(n7794));
  jxor g07539(.dina(n7794), .dinb(n1061), .dout(n7795));
  jxor g07540(.dina(n7795), .dinb(n7787), .dout(n7796));
  jxor g07541(.dina(n7796), .dinb(n7621), .dout(n7797));
  jor  g07542(.dina(n5038), .dinb(n970), .dout(n7798));
  jor  g07543(.dina(n880), .dinb(n4637), .dout(n7799));
  jor  g07544(.dina(n967), .dinb(n4839), .dout(n7800));
  jor  g07545(.dina(n972), .dinb(n5040), .dout(n7801));
  jand g07546(.dina(n7801), .dinb(n7800), .dout(n7802));
  jand g07547(.dina(n7802), .dinb(n7799), .dout(n7803));
  jand g07548(.dina(n7803), .dinb(n7798), .dout(n7804));
  jxor g07549(.dina(n7804), .dinb(n810), .dout(n7805));
  jxor g07550(.dina(n7805), .dinb(n7797), .dout(n7806));
  jxor g07551(.dina(n7806), .dinb(n7618), .dout(n7807));
  jor  g07552(.dina(n5683), .dinb(n728), .dout(n7808));
  jor  g07553(.dina(n660), .dinb(n5253), .dout(n7809));
  jor  g07554(.dina(n726), .dinb(n5685), .dout(n7810));
  jor  g07555(.dina(n731), .dinb(n5469), .dout(n7811));
  jand g07556(.dina(n7811), .dinb(n7810), .dout(n7812));
  jand g07557(.dina(n7812), .dinb(n7809), .dout(n7813));
  jand g07558(.dina(n7813), .dinb(n7808), .dout(n7814));
  jxor g07559(.dina(n7814), .dinb(n606), .dout(n7815));
  jxor g07560(.dina(n7815), .dinb(n7807), .dout(n7816));
  jnot g07561(.din(n7816), .dout(n7817));
  jxor g07562(.dina(n7817), .dinb(n7615), .dout(n7818));
  jor  g07563(.dina(n6364), .dinb(n544), .dout(n7819));
  jor  g07564(.dina(n486), .dinb(n5911), .dout(n7820));
  jor  g07565(.dina(n547), .dinb(n6139), .dout(n7821));
  jor  g07566(.dina(n542), .dinb(n6366), .dout(n7822));
  jand g07567(.dina(n7822), .dinb(n7821), .dout(n7823));
  jand g07568(.dina(n7823), .dinb(n7820), .dout(n7824));
  jand g07569(.dina(n7824), .dinb(n7819), .dout(n7825));
  jxor g07570(.dina(n7825), .dinb(n446), .dout(n7826));
  jxor g07571(.dina(n7826), .dinb(n7818), .dout(n7827));
  jxor g07572(.dina(n7827), .dinb(n7611), .dout(n7828));
  jor  g07573(.dina(n7084), .dinb(n397), .dout(n7829));
  jor  g07574(.dina(n354), .dinb(n6605), .dout(n7830));
  jor  g07575(.dina(n394), .dinb(n6846), .dout(n7831));
  jor  g07576(.dina(n399), .dinb(n7086), .dout(n7832));
  jand g07577(.dina(n7832), .dinb(n7831), .dout(n7833));
  jand g07578(.dina(n7833), .dinb(n7830), .dout(n7834));
  jand g07579(.dina(n7834), .dinb(n7829), .dout(n7835));
  jxor g07580(.dina(n7835), .dinb(n364), .dout(n7836));
  jxor g07581(.dina(n7836), .dinb(n7828), .dout(n7837));
  jxor g07582(.dina(n7837), .dinb(n7608), .dout(n7838));
  jand g07583(.dina(b53 ), .dinb(b52 ), .dout(n7839));
  jand g07584(.dina(n7586), .dinb(n7585), .dout(n7840));
  jor  g07585(.dina(n7840), .dinb(n7839), .dout(n7841));
  jxor g07586(.dina(b54 ), .dinb(b53 ), .dout(n7842));
  jnot g07587(.din(n7842), .dout(n7843));
  jxor g07588(.dina(n7843), .dinb(n7841), .dout(n7844));
  jor  g07589(.dina(n7844), .dinb(n296), .dout(n7845));
  jnot g07590(.din(b54 ), .dout(n7846));
  jor  g07591(.dina(n264), .dinb(n7846), .dout(n7847));
  jor  g07592(.dina(n280), .dinb(n7338), .dout(n7848));
  jor  g07593(.dina(n294), .dinb(n7590), .dout(n7849));
  jand g07594(.dina(n7849), .dinb(n7848), .dout(n7850));
  jand g07595(.dina(n7850), .dinb(n7847), .dout(n7851));
  jand g07596(.dina(n7851), .dinb(n7845), .dout(n7852));
  jxor g07597(.dina(n7852), .dinb(n278), .dout(n7853));
  jxor g07598(.dina(n7853), .dinb(n7838), .dout(n7854));
  jxor g07599(.dina(n7854), .dinb(n7603), .dout(f54 ));
  jnot g07600(.din(n7853), .dout(n7856));
  jor  g07601(.dina(n7856), .dinb(n7838), .dout(n7857));
  jor  g07602(.dina(n7854), .dinb(n7603), .dout(n7858));
  jand g07603(.dina(n7858), .dinb(n7857), .dout(n7859));
  jand g07604(.dina(n7836), .dinb(n7828), .dout(n7860));
  jnot g07605(.din(n7860), .dout(n7861));
  jnot g07606(.din(n7837), .dout(n7862));
  jor  g07607(.dina(n7862), .dinb(n7608), .dout(n7863));
  jand g07608(.dina(n7863), .dinb(n7861), .dout(n7864));
  jand g07609(.dina(n7826), .dinb(n7818), .dout(n7865));
  jand g07610(.dina(n7827), .dinb(n7611), .dout(n7866));
  jor  g07611(.dina(n7866), .dinb(n7865), .dout(n7867));
  jand g07612(.dina(n7815), .dinb(n7807), .dout(n7868));
  jnot g07613(.din(n7868), .dout(n7869));
  jor  g07614(.dina(n7817), .dinb(n7615), .dout(n7870));
  jand g07615(.dina(n7870), .dinb(n7869), .dout(n7871));
  jand g07616(.dina(n7805), .dinb(n7797), .dout(n7872));
  jand g07617(.dina(n7806), .dinb(n7618), .dout(n7873));
  jor  g07618(.dina(n7873), .dinb(n7872), .dout(n7874));
  jand g07619(.dina(n7795), .dinb(n7787), .dout(n7875));
  jand g07620(.dina(n7796), .dinb(n7621), .dout(n7876));
  jor  g07621(.dina(n7876), .dinb(n7875), .dout(n7877));
  jand g07622(.dina(n7785), .dinb(n7777), .dout(n7878));
  jand g07623(.dina(n7786), .dinb(n7624), .dout(n7879));
  jor  g07624(.dina(n7879), .dinb(n7878), .dout(n7880));
  jand g07625(.dina(n7775), .dinb(n7767), .dout(n7881));
  jand g07626(.dina(n7776), .dinb(n7627), .dout(n7882));
  jor  g07627(.dina(n7882), .dinb(n7881), .dout(n7883));
  jand g07628(.dina(n7765), .dinb(n7757), .dout(n7884));
  jand g07629(.dina(n7766), .dinb(n7630), .dout(n7885));
  jor  g07630(.dina(n7885), .dinb(n7884), .dout(n7886));
  jand g07631(.dina(n7755), .dinb(n7747), .dout(n7887));
  jand g07632(.dina(n7756), .dinb(n7633), .dout(n7888));
  jor  g07633(.dina(n7888), .dinb(n7887), .dout(n7889));
  jand g07634(.dina(n7745), .dinb(n7737), .dout(n7890));
  jand g07635(.dina(n7746), .dinb(n7636), .dout(n7891));
  jor  g07636(.dina(n7891), .dinb(n7890), .dout(n7892));
  jand g07637(.dina(n7735), .dinb(n7727), .dout(n7893));
  jand g07638(.dina(n7736), .dinb(n7639), .dout(n7894));
  jor  g07639(.dina(n7894), .dinb(n7893), .dout(n7895));
  jand g07640(.dina(n7725), .dinb(n7717), .dout(n7896));
  jand g07641(.dina(n7726), .dinb(n7642), .dout(n7897));
  jor  g07642(.dina(n7897), .dinb(n7896), .dout(n7898));
  jand g07643(.dina(n7715), .dinb(n7707), .dout(n7899));
  jand g07644(.dina(n7716), .dinb(n7645), .dout(n7900));
  jor  g07645(.dina(n7900), .dinb(n7899), .dout(n7901));
  jand g07646(.dina(n7705), .dinb(n7697), .dout(n7902));
  jand g07647(.dina(n7706), .dinb(n7648), .dout(n7903));
  jor  g07648(.dina(n7903), .dinb(n7902), .dout(n7904));
  jand g07649(.dina(n7695), .dinb(n7687), .dout(n7905));
  jand g07650(.dina(n7696), .dinb(n7651), .dout(n7906));
  jor  g07651(.dina(n7906), .dinb(n7905), .dout(n7907));
  jor  g07652(.dina(n7677), .dinb(n7669), .dout(n7908));
  jand g07653(.dina(n7686), .dinb(n7678), .dout(n7909));
  jnot g07654(.din(n7909), .dout(n7910));
  jand g07655(.dina(n7910), .dinb(n7908), .dout(n7911));
  jnot g07656(.din(n7911), .dout(n7912));
  jnot g07657(.din(n7652), .dout(n7913));
  jand g07658(.dina(n7654), .dinb(n7913), .dout(n7914));
  jand g07659(.dina(n7667), .dinb(n7656), .dout(n7915));
  jor  g07660(.dina(n7915), .dinb(n7914), .dout(n7916));
  jxor g07661(.dina(a56 ), .dinb(a55 ), .dout(n7917));
  jand g07662(.dina(n7917), .dinb(n7653), .dout(n7918));
  jand g07663(.dina(n7918), .dinb(n259), .dout(n7919));
  jnot g07664(.din(n7653), .dout(n7920));
  jxor g07665(.dina(a55 ), .dinb(a54 ), .dout(n7921));
  jand g07666(.dina(n7921), .dinb(n7920), .dout(n7922));
  jand g07667(.dina(n7922), .dinb(b0 ), .dout(n7923));
  jnot g07668(.din(n7917), .dout(n7924));
  jand g07669(.dina(n7924), .dinb(n7653), .dout(n7925));
  jand g07670(.dina(n7925), .dinb(b1 ), .dout(n7926));
  jor  g07671(.dina(n7926), .dinb(n7923), .dout(n7927));
  jor  g07672(.dina(n7927), .dinb(n7919), .dout(n7928));
  jnot g07673(.din(a56 ), .dout(n7929));
  jor  g07674(.dina(n7655), .dinb(n7929), .dout(n7930));
  jxor g07675(.dina(n7930), .dinb(n7928), .dout(n7931));
  jor  g07676(.dina(n7660), .dinb(n337), .dout(n7932));
  jor  g07677(.dina(n7662), .dinb(n340), .dout(n7933));
  jor  g07678(.dina(n7415), .dinb(n293), .dout(n7934));
  jand g07679(.dina(n7934), .dinb(n7933), .dout(n7935));
  jor  g07680(.dina(n7657), .dinb(n303), .dout(n7936));
  jand g07681(.dina(n7936), .dinb(n7935), .dout(n7937));
  jand g07682(.dina(n7937), .dinb(n7932), .dout(n7938));
  jxor g07683(.dina(n7938), .dinb(a53 ), .dout(n7939));
  jxor g07684(.dina(n7939), .dinb(n7931), .dout(n7940));
  jxor g07685(.dina(n7940), .dinb(n7916), .dout(n7941));
  jnot g07686(.din(n7941), .dout(n7942));
  jor  g07687(.dina(n6914), .dinb(n466), .dout(n7943));
  jor  g07688(.dina(n6916), .dinb(n469), .dout(n7944));
  jor  g07689(.dina(n6673), .dinb(n377), .dout(n7945));
  jand g07690(.dina(n7945), .dinb(n7944), .dout(n7946));
  jor  g07691(.dina(n6911), .dinb(n415), .dout(n7947));
  jand g07692(.dina(n7947), .dinb(n7946), .dout(n7948));
  jand g07693(.dina(n7948), .dinb(n7943), .dout(n7949));
  jxor g07694(.dina(n7949), .dinb(a50 ), .dout(n7950));
  jxor g07695(.dina(n7950), .dinb(n7942), .dout(n7951));
  jxor g07696(.dina(n7951), .dinb(n7912), .dout(n7952));
  jor  g07697(.dina(n6207), .dinb(n635), .dout(n7953));
  jor  g07698(.dina(n5975), .dinb(n519), .dout(n7954));
  jor  g07699(.dina(n6205), .dinb(n637), .dout(n7955));
  jor  g07700(.dina(n6210), .dinb(n572), .dout(n7956));
  jand g07701(.dina(n7956), .dinb(n7955), .dout(n7957));
  jand g07702(.dina(n7957), .dinb(n7954), .dout(n7958));
  jand g07703(.dina(n7958), .dinb(n7953), .dout(n7959));
  jxor g07704(.dina(n7959), .dinb(n5759), .dout(n7960));
  jxor g07705(.dina(n7960), .dinb(n7952), .dout(n7961));
  jxor g07706(.dina(n7961), .dinb(n7907), .dout(n7962));
  jor  g07707(.dina(n5537), .dinb(n850), .dout(n7963));
  jor  g07708(.dina(n5315), .dinb(n704), .dout(n7964));
  jor  g07709(.dina(n5539), .dinb(n852), .dout(n7965));
  jor  g07710(.dina(n5534), .dinb(n772), .dout(n7966));
  jand g07711(.dina(n7966), .dinb(n7965), .dout(n7967));
  jand g07712(.dina(n7967), .dinb(n7964), .dout(n7968));
  jand g07713(.dina(n7968), .dinb(n7963), .dout(n7969));
  jxor g07714(.dina(n7969), .dinb(n5111), .dout(n7970));
  jxor g07715(.dina(n7970), .dinb(n7962), .dout(n7971));
  jxor g07716(.dina(n7971), .dinb(n7904), .dout(n7972));
  jor  g07717(.dina(n4902), .dinb(n1112), .dout(n7973));
  jor  g07718(.dina(n4696), .dinb(n934), .dout(n7974));
  jor  g07719(.dina(n4899), .dinb(n1114), .dout(n7975));
  jor  g07720(.dina(n4904), .dinb(n1018), .dout(n7976));
  jand g07721(.dina(n7976), .dinb(n7975), .dout(n7977));
  jand g07722(.dina(n7977), .dinb(n7974), .dout(n7978));
  jand g07723(.dina(n7978), .dinb(n7973), .dout(n7979));
  jxor g07724(.dina(n7979), .dinb(n4505), .dout(n7980));
  jxor g07725(.dina(n7980), .dinb(n7972), .dout(n7981));
  jxor g07726(.dina(n7981), .dinb(n7901), .dout(n7982));
  jor  g07727(.dina(n4305), .dinb(n1414), .dout(n7983));
  jor  g07728(.dina(n4116), .dinb(n1211), .dout(n7984));
  jor  g07729(.dina(n4308), .dinb(n1307), .dout(n7985));
  jor  g07730(.dina(n4303), .dinb(n1416), .dout(n7986));
  jand g07731(.dina(n7986), .dinb(n7985), .dout(n7987));
  jand g07732(.dina(n7987), .dinb(n7984), .dout(n7988));
  jand g07733(.dina(n7988), .dinb(n7983), .dout(n7989));
  jxor g07734(.dina(n7989), .dinb(n3938), .dout(n7990));
  jxor g07735(.dina(n7990), .dinb(n7982), .dout(n7991));
  jxor g07736(.dina(n7991), .dinb(n7898), .dout(n7992));
  jor  g07737(.dina(n3751), .dinb(n1757), .dout(n7993));
  jor  g07738(.dina(n3574), .dinb(n1527), .dout(n7994));
  jor  g07739(.dina(n3754), .dinb(n1637), .dout(n7995));
  jor  g07740(.dina(n3749), .dinb(n1759), .dout(n7996));
  jand g07741(.dina(n7996), .dinb(n7995), .dout(n7997));
  jand g07742(.dina(n7997), .dinb(n7994), .dout(n7998));
  jand g07743(.dina(n7998), .dinb(n7993), .dout(n7999));
  jxor g07744(.dina(n7999), .dinb(n3410), .dout(n8000));
  jxor g07745(.dina(n8000), .dinb(n7992), .dout(n8001));
  jxor g07746(.dina(n8001), .dinb(n7895), .dout(n8002));
  jor  g07747(.dina(n3239), .dinb(n2140), .dout(n8003));
  jor  g07748(.dina(n3072), .dinb(n1881), .dout(n8004));
  jor  g07749(.dina(n3237), .dinb(n2142), .dout(n8005));
  jor  g07750(.dina(n3242), .dinb(n2007), .dout(n8006));
  jand g07751(.dina(n8006), .dinb(n8005), .dout(n8007));
  jand g07752(.dina(n8007), .dinb(n8004), .dout(n8008));
  jand g07753(.dina(n8008), .dinb(n8003), .dout(n8009));
  jxor g07754(.dina(n8009), .dinb(n2918), .dout(n8010));
  jxor g07755(.dina(n8010), .dinb(n8002), .dout(n8011));
  jxor g07756(.dina(n8011), .dinb(n7892), .dout(n8012));
  jor  g07757(.dina(n2561), .dinb(n2764), .dout(n8013));
  jor  g07758(.dina(n2609), .dinb(n2279), .dout(n8014));
  jor  g07759(.dina(n2761), .dinb(n2563), .dout(n8015));
  jor  g07760(.dina(n2766), .dinb(n2415), .dout(n8016));
  jand g07761(.dina(n8016), .dinb(n8015), .dout(n8017));
  jand g07762(.dina(n8017), .dinb(n8014), .dout(n8018));
  jand g07763(.dina(n8018), .dinb(n8013), .dout(n8019));
  jxor g07764(.dina(n8019), .dinb(n2468), .dout(n8020));
  jxor g07765(.dina(n8020), .dinb(n8012), .dout(n8021));
  jxor g07766(.dina(n8021), .dinb(n7889), .dout(n8022));
  jor  g07767(.dina(n3021), .dinb(n2324), .dout(n8023));
  jor  g07768(.dina(n2186), .dinb(n2713), .dout(n8024));
  jor  g07769(.dina(n2321), .dinb(n2862), .dout(n8025));
  jor  g07770(.dina(n2326), .dinb(n3023), .dout(n8026));
  jand g07771(.dina(n8026), .dinb(n8025), .dout(n8027));
  jand g07772(.dina(n8027), .dinb(n8024), .dout(n8028));
  jand g07773(.dina(n8028), .dinb(n8023), .dout(n8029));
  jxor g07774(.dina(n8029), .dinb(n2057), .dout(n8030));
  jxor g07775(.dina(n8030), .dinb(n8022), .dout(n8031));
  jxor g07776(.dina(n8031), .dinb(n7886), .dout(n8032));
  jor  g07777(.dina(n3520), .dinb(n1921), .dout(n8033));
  jor  g07778(.dina(n1806), .dinb(n3186), .dout(n8034));
  jor  g07779(.dina(n1923), .dinb(n3522), .dout(n8035));
  jor  g07780(.dina(n1918), .dinb(n3348), .dout(n8036));
  jand g07781(.dina(n8036), .dinb(n8035), .dout(n8037));
  jand g07782(.dina(n8037), .dinb(n8034), .dout(n8038));
  jand g07783(.dina(n8038), .dinb(n8033), .dout(n8039));
  jxor g07784(.dina(n8039), .dinb(n1687), .dout(n8040));
  jxor g07785(.dina(n8040), .dinb(n8032), .dout(n8041));
  jxor g07786(.dina(n8041), .dinb(n7883), .dout(n8042));
  jor  g07787(.dina(n4058), .dinb(n1569), .dout(n8043));
  jor  g07788(.dina(n1453), .dinb(n3698), .dout(n8044));
  jor  g07789(.dina(n1566), .dinb(n3873), .dout(n8045));
  jor  g07790(.dina(n1571), .dinb(n4060), .dout(n8046));
  jand g07791(.dina(n8046), .dinb(n8045), .dout(n8047));
  jand g07792(.dina(n8047), .dinb(n8044), .dout(n8048));
  jand g07793(.dina(n8048), .dinb(n8043), .dout(n8049));
  jxor g07794(.dina(n8049), .dinb(n1351), .dout(n8050));
  jxor g07795(.dina(n8050), .dinb(n8042), .dout(n8051));
  jxor g07796(.dina(n8051), .dinb(n7880), .dout(n8052));
  jor  g07797(.dina(n4635), .dinb(n1248), .dout(n8053));
  jor  g07798(.dina(n1147), .dinb(n4249), .dout(n8054));
  jor  g07799(.dina(n1246), .dinb(n4637), .dout(n8055));
  jor  g07800(.dina(n1251), .dinb(n4437), .dout(n8056));
  jand g07801(.dina(n8056), .dinb(n8055), .dout(n8057));
  jand g07802(.dina(n8057), .dinb(n8054), .dout(n8058));
  jand g07803(.dina(n8058), .dinb(n8053), .dout(n8059));
  jxor g07804(.dina(n8059), .dinb(n1061), .dout(n8060));
  jxor g07805(.dina(n8060), .dinb(n8052), .dout(n8061));
  jxor g07806(.dina(n8061), .dinb(n7877), .dout(n8062));
  jor  g07807(.dina(n5251), .dinb(n970), .dout(n8063));
  jor  g07808(.dina(n880), .dinb(n4839), .dout(n8064));
  jor  g07809(.dina(n967), .dinb(n5040), .dout(n8065));
  jor  g07810(.dina(n972), .dinb(n5253), .dout(n8066));
  jand g07811(.dina(n8066), .dinb(n8065), .dout(n8067));
  jand g07812(.dina(n8067), .dinb(n8064), .dout(n8068));
  jand g07813(.dina(n8068), .dinb(n8063), .dout(n8069));
  jxor g07814(.dina(n8069), .dinb(n810), .dout(n8070));
  jxor g07815(.dina(n8070), .dinb(n8062), .dout(n8071));
  jxor g07816(.dina(n8071), .dinb(n7874), .dout(n8072));
  jor  g07817(.dina(n5909), .dinb(n728), .dout(n8073));
  jor  g07818(.dina(n660), .dinb(n5469), .dout(n8074));
  jor  g07819(.dina(n731), .dinb(n5685), .dout(n8075));
  jor  g07820(.dina(n726), .dinb(n5911), .dout(n8076));
  jand g07821(.dina(n8076), .dinb(n8075), .dout(n8077));
  jand g07822(.dina(n8077), .dinb(n8074), .dout(n8078));
  jand g07823(.dina(n8078), .dinb(n8073), .dout(n8079));
  jxor g07824(.dina(n8079), .dinb(n606), .dout(n8080));
  jxor g07825(.dina(n8080), .dinb(n8072), .dout(n8081));
  jnot g07826(.din(n8081), .dout(n8082));
  jxor g07827(.dina(n8082), .dinb(n7871), .dout(n8083));
  jor  g07828(.dina(n6603), .dinb(n544), .dout(n8084));
  jor  g07829(.dina(n486), .dinb(n6139), .dout(n8085));
  jor  g07830(.dina(n547), .dinb(n6366), .dout(n8086));
  jor  g07831(.dina(n542), .dinb(n6605), .dout(n8087));
  jand g07832(.dina(n8087), .dinb(n8086), .dout(n8088));
  jand g07833(.dina(n8088), .dinb(n8085), .dout(n8089));
  jand g07834(.dina(n8089), .dinb(n8084), .dout(n8090));
  jxor g07835(.dina(n8090), .dinb(n446), .dout(n8091));
  jxor g07836(.dina(n8091), .dinb(n8083), .dout(n8092));
  jxor g07837(.dina(n8092), .dinb(n7867), .dout(n8093));
  jor  g07838(.dina(n7336), .dinb(n397), .dout(n8094));
  jor  g07839(.dina(n354), .dinb(n6846), .dout(n8095));
  jor  g07840(.dina(n399), .dinb(n7338), .dout(n8096));
  jor  g07841(.dina(n394), .dinb(n7086), .dout(n8097));
  jand g07842(.dina(n8097), .dinb(n8096), .dout(n8098));
  jand g07843(.dina(n8098), .dinb(n8095), .dout(n8099));
  jand g07844(.dina(n8099), .dinb(n8094), .dout(n8100));
  jxor g07845(.dina(n8100), .dinb(n364), .dout(n8101));
  jxor g07846(.dina(n8101), .dinb(n8093), .dout(n8102));
  jxor g07847(.dina(n8102), .dinb(n7864), .dout(n8103));
  jand g07848(.dina(b54 ), .dinb(b53 ), .dout(n8104));
  jand g07849(.dina(n7842), .dinb(n7841), .dout(n8105));
  jor  g07850(.dina(n8105), .dinb(n8104), .dout(n8106));
  jxor g07851(.dina(b55 ), .dinb(b54 ), .dout(n8107));
  jnot g07852(.din(n8107), .dout(n8108));
  jxor g07853(.dina(n8108), .dinb(n8106), .dout(n8109));
  jor  g07854(.dina(n8109), .dinb(n296), .dout(n8110));
  jnot g07855(.din(b55 ), .dout(n8111));
  jor  g07856(.dina(n264), .dinb(n8111), .dout(n8112));
  jor  g07857(.dina(n280), .dinb(n7590), .dout(n8113));
  jor  g07858(.dina(n294), .dinb(n7846), .dout(n8114));
  jand g07859(.dina(n8114), .dinb(n8113), .dout(n8115));
  jand g07860(.dina(n8115), .dinb(n8112), .dout(n8116));
  jand g07861(.dina(n8116), .dinb(n8110), .dout(n8117));
  jxor g07862(.dina(n8117), .dinb(n278), .dout(n8118));
  jxor g07863(.dina(n8118), .dinb(n8103), .dout(n8119));
  jxor g07864(.dina(n8119), .dinb(n7859), .dout(f55 ));
  jnot g07865(.din(n8118), .dout(n8121));
  jor  g07866(.dina(n8121), .dinb(n8103), .dout(n8122));
  jor  g07867(.dina(n8119), .dinb(n7859), .dout(n8123));
  jand g07868(.dina(n8123), .dinb(n8122), .dout(n8124));
  jand g07869(.dina(n8101), .dinb(n8093), .dout(n8125));
  jnot g07870(.din(n8125), .dout(n8126));
  jnot g07871(.din(n8102), .dout(n8127));
  jor  g07872(.dina(n8127), .dinb(n7864), .dout(n8128));
  jand g07873(.dina(n8128), .dinb(n8126), .dout(n8129));
  jand g07874(.dina(n8091), .dinb(n8083), .dout(n8130));
  jand g07875(.dina(n8092), .dinb(n7867), .dout(n8131));
  jor  g07876(.dina(n8131), .dinb(n8130), .dout(n8132));
  jand g07877(.dina(n8080), .dinb(n8072), .dout(n8133));
  jnot g07878(.din(n8133), .dout(n8134));
  jor  g07879(.dina(n8082), .dinb(n7871), .dout(n8135));
  jand g07880(.dina(n8135), .dinb(n8134), .dout(n8136));
  jand g07881(.dina(n8070), .dinb(n8062), .dout(n8137));
  jand g07882(.dina(n8071), .dinb(n7874), .dout(n8138));
  jor  g07883(.dina(n8138), .dinb(n8137), .dout(n8139));
  jand g07884(.dina(n8060), .dinb(n8052), .dout(n8140));
  jand g07885(.dina(n8061), .dinb(n7877), .dout(n8141));
  jor  g07886(.dina(n8141), .dinb(n8140), .dout(n8142));
  jand g07887(.dina(n8050), .dinb(n8042), .dout(n8143));
  jand g07888(.dina(n8051), .dinb(n7880), .dout(n8144));
  jor  g07889(.dina(n8144), .dinb(n8143), .dout(n8145));
  jand g07890(.dina(n8040), .dinb(n8032), .dout(n8146));
  jand g07891(.dina(n8041), .dinb(n7883), .dout(n8147));
  jor  g07892(.dina(n8147), .dinb(n8146), .dout(n8148));
  jand g07893(.dina(n8030), .dinb(n8022), .dout(n8149));
  jand g07894(.dina(n8031), .dinb(n7886), .dout(n8150));
  jor  g07895(.dina(n8150), .dinb(n8149), .dout(n8151));
  jand g07896(.dina(n8020), .dinb(n8012), .dout(n8152));
  jand g07897(.dina(n8021), .dinb(n7889), .dout(n8153));
  jor  g07898(.dina(n8153), .dinb(n8152), .dout(n8154));
  jand g07899(.dina(n8010), .dinb(n8002), .dout(n8155));
  jand g07900(.dina(n8011), .dinb(n7892), .dout(n8156));
  jor  g07901(.dina(n8156), .dinb(n8155), .dout(n8157));
  jand g07902(.dina(n8000), .dinb(n7992), .dout(n8158));
  jand g07903(.dina(n8001), .dinb(n7895), .dout(n8159));
  jor  g07904(.dina(n8159), .dinb(n8158), .dout(n8160));
  jand g07905(.dina(n7990), .dinb(n7982), .dout(n8161));
  jand g07906(.dina(n7991), .dinb(n7898), .dout(n8162));
  jor  g07907(.dina(n8162), .dinb(n8161), .dout(n8163));
  jand g07908(.dina(n7980), .dinb(n7972), .dout(n8164));
  jand g07909(.dina(n7981), .dinb(n7901), .dout(n8165));
  jor  g07910(.dina(n8165), .dinb(n8164), .dout(n8166));
  jand g07911(.dina(n7970), .dinb(n7962), .dout(n8167));
  jand g07912(.dina(n7971), .dinb(n7904), .dout(n8168));
  jor  g07913(.dina(n8168), .dinb(n8167), .dout(n8169));
  jand g07914(.dina(n7960), .dinb(n7952), .dout(n8170));
  jand g07915(.dina(n7961), .dinb(n7907), .dout(n8171));
  jor  g07916(.dina(n8171), .dinb(n8170), .dout(n8172));
  jor  g07917(.dina(n7950), .dinb(n7942), .dout(n8173));
  jand g07918(.dina(n7951), .dinb(n7912), .dout(n8174));
  jnot g07919(.din(n8174), .dout(n8175));
  jand g07920(.dina(n8175), .dinb(n8173), .dout(n8176));
  jnot g07921(.din(n8176), .dout(n8177));
  jor  g07922(.dina(n7939), .dinb(n7931), .dout(n8178));
  jand g07923(.dina(n7940), .dinb(n7916), .dout(n8179));
  jnot g07924(.din(n8179), .dout(n8180));
  jand g07925(.dina(n8180), .dinb(n8178), .dout(n8181));
  jnot g07926(.din(n8181), .dout(n8182));
  jand g07927(.dina(n7922), .dinb(b1 ), .dout(n8183));
  jor  g07928(.dina(n7921), .dinb(n7653), .dout(n8184));
  jor  g07929(.dina(n8184), .dinb(n7924), .dout(n8185));
  jnot g07930(.din(n8185), .dout(n8186));
  jand g07931(.dina(n8186), .dinb(b0 ), .dout(n8187));
  jand g07932(.dina(n7918), .dinb(n273), .dout(n8188));
  jand g07933(.dina(n7925), .dinb(b2 ), .dout(n8189));
  jor  g07934(.dina(n8189), .dinb(n8188), .dout(n8190));
  jor  g07935(.dina(n8190), .dinb(n8187), .dout(n8191));
  jor  g07936(.dina(n8191), .dinb(n8183), .dout(n8192));
  jnot g07937(.din(n7928), .dout(n8193));
  jand g07938(.dina(n7655), .dinb(a56 ), .dout(n8194));
  jand g07939(.dina(n8194), .dinb(n8193), .dout(n8195));
  jnot g07940(.din(n8195), .dout(n8196));
  jand g07941(.dina(n8196), .dinb(a56 ), .dout(n8197));
  jxor g07942(.dina(n8197), .dinb(n8192), .dout(n8198));
  jnot g07943(.din(n8198), .dout(n8199));
  jor  g07944(.dina(n7660), .dinb(n374), .dout(n8200));
  jor  g07945(.dina(n7662), .dinb(n377), .dout(n8201));
  jor  g07946(.dina(n7415), .dinb(n303), .dout(n8202));
  jand g07947(.dina(n8202), .dinb(n8201), .dout(n8203));
  jor  g07948(.dina(n7657), .dinb(n340), .dout(n8204));
  jand g07949(.dina(n8204), .dinb(n8203), .dout(n8205));
  jand g07950(.dina(n8205), .dinb(n8200), .dout(n8206));
  jxor g07951(.dina(n8206), .dinb(a53 ), .dout(n8207));
  jxor g07952(.dina(n8207), .dinb(n8199), .dout(n8208));
  jxor g07953(.dina(n8208), .dinb(n8182), .dout(n8209));
  jor  g07954(.dina(n6914), .dinb(n517), .dout(n8210));
  jor  g07955(.dina(n6916), .dinb(n519), .dout(n8211));
  jor  g07956(.dina(n6911), .dinb(n469), .dout(n8212));
  jor  g07957(.dina(n6673), .dinb(n415), .dout(n8213));
  jand g07958(.dina(n8213), .dinb(n8212), .dout(n8214));
  jand g07959(.dina(n8214), .dinb(n8211), .dout(n8215));
  jand g07960(.dina(n8215), .dinb(n8210), .dout(n8216));
  jxor g07961(.dina(n8216), .dinb(n6443), .dout(n8217));
  jxor g07962(.dina(n8217), .dinb(n8209), .dout(n8218));
  jxor g07963(.dina(n8218), .dinb(n8177), .dout(n8219));
  jor  g07964(.dina(n6207), .dinb(n702), .dout(n8220));
  jor  g07965(.dina(n5975), .dinb(n572), .dout(n8221));
  jor  g07966(.dina(n6205), .dinb(n704), .dout(n8222));
  jor  g07967(.dina(n6210), .dinb(n637), .dout(n8223));
  jand g07968(.dina(n8223), .dinb(n8222), .dout(n8224));
  jand g07969(.dina(n8224), .dinb(n8221), .dout(n8225));
  jand g07970(.dina(n8225), .dinb(n8220), .dout(n8226));
  jxor g07971(.dina(n8226), .dinb(n5759), .dout(n8227));
  jxor g07972(.dina(n8227), .dinb(n8219), .dout(n8228));
  jxor g07973(.dina(n8228), .dinb(n8172), .dout(n8229));
  jor  g07974(.dina(n5537), .dinb(n932), .dout(n8230));
  jor  g07975(.dina(n5315), .dinb(n772), .dout(n8231));
  jor  g07976(.dina(n5539), .dinb(n934), .dout(n8232));
  jor  g07977(.dina(n5534), .dinb(n852), .dout(n8233));
  jand g07978(.dina(n8233), .dinb(n8232), .dout(n8234));
  jand g07979(.dina(n8234), .dinb(n8231), .dout(n8235));
  jand g07980(.dina(n8235), .dinb(n8230), .dout(n8236));
  jxor g07981(.dina(n8236), .dinb(n5111), .dout(n8237));
  jxor g07982(.dina(n8237), .dinb(n8229), .dout(n8238));
  jxor g07983(.dina(n8238), .dinb(n8169), .dout(n8239));
  jor  g07984(.dina(n4902), .dinb(n1209), .dout(n8240));
  jor  g07985(.dina(n4696), .dinb(n1018), .dout(n8241));
  jor  g07986(.dina(n4904), .dinb(n1114), .dout(n8242));
  jor  g07987(.dina(n4899), .dinb(n1211), .dout(n8243));
  jand g07988(.dina(n8243), .dinb(n8242), .dout(n8244));
  jand g07989(.dina(n8244), .dinb(n8241), .dout(n8245));
  jand g07990(.dina(n8245), .dinb(n8240), .dout(n8246));
  jxor g07991(.dina(n8246), .dinb(n4505), .dout(n8247));
  jxor g07992(.dina(n8247), .dinb(n8239), .dout(n8248));
  jxor g07993(.dina(n8248), .dinb(n8166), .dout(n8249));
  jor  g07994(.dina(n4305), .dinb(n1525), .dout(n8250));
  jor  g07995(.dina(n4116), .dinb(n1307), .dout(n8251));
  jor  g07996(.dina(n4303), .dinb(n1527), .dout(n8252));
  jor  g07997(.dina(n4308), .dinb(n1416), .dout(n8253));
  jand g07998(.dina(n8253), .dinb(n8252), .dout(n8254));
  jand g07999(.dina(n8254), .dinb(n8251), .dout(n8255));
  jand g08000(.dina(n8255), .dinb(n8250), .dout(n8256));
  jxor g08001(.dina(n8256), .dinb(n3938), .dout(n8257));
  jxor g08002(.dina(n8257), .dinb(n8249), .dout(n8258));
  jxor g08003(.dina(n8258), .dinb(n8163), .dout(n8259));
  jor  g08004(.dina(n3751), .dinb(n1879), .dout(n8260));
  jor  g08005(.dina(n3574), .dinb(n1637), .dout(n8261));
  jor  g08006(.dina(n3749), .dinb(n1881), .dout(n8262));
  jor  g08007(.dina(n3754), .dinb(n1759), .dout(n8263));
  jand g08008(.dina(n8263), .dinb(n8262), .dout(n8264));
  jand g08009(.dina(n8264), .dinb(n8261), .dout(n8265));
  jand g08010(.dina(n8265), .dinb(n8260), .dout(n8266));
  jxor g08011(.dina(n8266), .dinb(n3410), .dout(n8267));
  jxor g08012(.dina(n8267), .dinb(n8259), .dout(n8268));
  jxor g08013(.dina(n8268), .dinb(n8160), .dout(n8269));
  jor  g08014(.dina(n3239), .dinb(n2277), .dout(n8270));
  jor  g08015(.dina(n3072), .dinb(n2007), .dout(n8271));
  jor  g08016(.dina(n3242), .dinb(n2142), .dout(n8272));
  jor  g08017(.dina(n3237), .dinb(n2279), .dout(n8273));
  jand g08018(.dina(n8273), .dinb(n8272), .dout(n8274));
  jand g08019(.dina(n8274), .dinb(n8271), .dout(n8275));
  jand g08020(.dina(n8275), .dinb(n8270), .dout(n8276));
  jxor g08021(.dina(n8276), .dinb(n2918), .dout(n8277));
  jxor g08022(.dina(n8277), .dinb(n8269), .dout(n8278));
  jxor g08023(.dina(n8278), .dinb(n8157), .dout(n8279));
  jor  g08024(.dina(n2711), .dinb(n2764), .dout(n8280));
  jor  g08025(.dina(n2609), .dinb(n2415), .dout(n8281));
  jor  g08026(.dina(n2761), .dinb(n2713), .dout(n8282));
  jor  g08027(.dina(n2766), .dinb(n2563), .dout(n8283));
  jand g08028(.dina(n8283), .dinb(n8282), .dout(n8284));
  jand g08029(.dina(n8284), .dinb(n8281), .dout(n8285));
  jand g08030(.dina(n8285), .dinb(n8280), .dout(n8286));
  jxor g08031(.dina(n8286), .dinb(n2468), .dout(n8287));
  jxor g08032(.dina(n8287), .dinb(n8279), .dout(n8288));
  jxor g08033(.dina(n8288), .dinb(n8154), .dout(n8289));
  jor  g08034(.dina(n3184), .dinb(n2324), .dout(n8290));
  jor  g08035(.dina(n2186), .dinb(n2862), .dout(n8291));
  jor  g08036(.dina(n2321), .dinb(n3023), .dout(n8292));
  jor  g08037(.dina(n2326), .dinb(n3186), .dout(n8293));
  jand g08038(.dina(n8293), .dinb(n8292), .dout(n8294));
  jand g08039(.dina(n8294), .dinb(n8291), .dout(n8295));
  jand g08040(.dina(n8295), .dinb(n8290), .dout(n8296));
  jxor g08041(.dina(n8296), .dinb(n2057), .dout(n8297));
  jxor g08042(.dina(n8297), .dinb(n8289), .dout(n8298));
  jxor g08043(.dina(n8298), .dinb(n8151), .dout(n8299));
  jor  g08044(.dina(n3696), .dinb(n1921), .dout(n8300));
  jor  g08045(.dina(n1806), .dinb(n3348), .dout(n8301));
  jor  g08046(.dina(n1918), .dinb(n3522), .dout(n8302));
  jor  g08047(.dina(n1923), .dinb(n3698), .dout(n8303));
  jand g08048(.dina(n8303), .dinb(n8302), .dout(n8304));
  jand g08049(.dina(n8304), .dinb(n8301), .dout(n8305));
  jand g08050(.dina(n8305), .dinb(n8300), .dout(n8306));
  jxor g08051(.dina(n8306), .dinb(n1687), .dout(n8307));
  jxor g08052(.dina(n8307), .dinb(n8299), .dout(n8308));
  jxor g08053(.dina(n8308), .dinb(n8148), .dout(n8309));
  jor  g08054(.dina(n4247), .dinb(n1569), .dout(n8310));
  jor  g08055(.dina(n1453), .dinb(n3873), .dout(n8311));
  jor  g08056(.dina(n1566), .dinb(n4060), .dout(n8312));
  jor  g08057(.dina(n1571), .dinb(n4249), .dout(n8313));
  jand g08058(.dina(n8313), .dinb(n8312), .dout(n8314));
  jand g08059(.dina(n8314), .dinb(n8311), .dout(n8315));
  jand g08060(.dina(n8315), .dinb(n8310), .dout(n8316));
  jxor g08061(.dina(n8316), .dinb(n1351), .dout(n8317));
  jxor g08062(.dina(n8317), .dinb(n8309), .dout(n8318));
  jxor g08063(.dina(n8318), .dinb(n8145), .dout(n8319));
  jor  g08064(.dina(n4837), .dinb(n1248), .dout(n8320));
  jor  g08065(.dina(n1147), .dinb(n4437), .dout(n8321));
  jor  g08066(.dina(n1246), .dinb(n4839), .dout(n8322));
  jor  g08067(.dina(n1251), .dinb(n4637), .dout(n8323));
  jand g08068(.dina(n8323), .dinb(n8322), .dout(n8324));
  jand g08069(.dina(n8324), .dinb(n8321), .dout(n8325));
  jand g08070(.dina(n8325), .dinb(n8320), .dout(n8326));
  jxor g08071(.dina(n8326), .dinb(n1061), .dout(n8327));
  jxor g08072(.dina(n8327), .dinb(n8319), .dout(n8328));
  jxor g08073(.dina(n8328), .dinb(n8142), .dout(n8329));
  jor  g08074(.dina(n5467), .dinb(n970), .dout(n8330));
  jor  g08075(.dina(n880), .dinb(n5040), .dout(n8331));
  jor  g08076(.dina(n967), .dinb(n5253), .dout(n8332));
  jor  g08077(.dina(n972), .dinb(n5469), .dout(n8333));
  jand g08078(.dina(n8333), .dinb(n8332), .dout(n8334));
  jand g08079(.dina(n8334), .dinb(n8331), .dout(n8335));
  jand g08080(.dina(n8335), .dinb(n8330), .dout(n8336));
  jxor g08081(.dina(n8336), .dinb(n810), .dout(n8337));
  jxor g08082(.dina(n8337), .dinb(n8329), .dout(n8338));
  jxor g08083(.dina(n8338), .dinb(n8139), .dout(n8339));
  jor  g08084(.dina(n6137), .dinb(n728), .dout(n8340));
  jor  g08085(.dina(n660), .dinb(n5685), .dout(n8341));
  jor  g08086(.dina(n731), .dinb(n5911), .dout(n8342));
  jor  g08087(.dina(n726), .dinb(n6139), .dout(n8343));
  jand g08088(.dina(n8343), .dinb(n8342), .dout(n8344));
  jand g08089(.dina(n8344), .dinb(n8341), .dout(n8345));
  jand g08090(.dina(n8345), .dinb(n8340), .dout(n8346));
  jxor g08091(.dina(n8346), .dinb(n606), .dout(n8347));
  jxor g08092(.dina(n8347), .dinb(n8339), .dout(n8348));
  jxor g08093(.dina(n8348), .dinb(n8136), .dout(n8349));
  jor  g08094(.dina(n6844), .dinb(n544), .dout(n8350));
  jor  g08095(.dina(n486), .dinb(n6366), .dout(n8351));
  jor  g08096(.dina(n547), .dinb(n6605), .dout(n8352));
  jor  g08097(.dina(n542), .dinb(n6846), .dout(n8353));
  jand g08098(.dina(n8353), .dinb(n8352), .dout(n8354));
  jand g08099(.dina(n8354), .dinb(n8351), .dout(n8355));
  jand g08100(.dina(n8355), .dinb(n8350), .dout(n8356));
  jxor g08101(.dina(n8356), .dinb(n446), .dout(n8357));
  jxor g08102(.dina(n8357), .dinb(n8349), .dout(n8358));
  jnot g08103(.din(n8358), .dout(n8359));
  jxor g08104(.dina(n8359), .dinb(n8132), .dout(n8360));
  jor  g08105(.dina(n7588), .dinb(n397), .dout(n8361));
  jor  g08106(.dina(n354), .dinb(n7086), .dout(n8362));
  jor  g08107(.dina(n399), .dinb(n7590), .dout(n8363));
  jor  g08108(.dina(n394), .dinb(n7338), .dout(n8364));
  jand g08109(.dina(n8364), .dinb(n8363), .dout(n8365));
  jand g08110(.dina(n8365), .dinb(n8362), .dout(n8366));
  jand g08111(.dina(n8366), .dinb(n8361), .dout(n8367));
  jxor g08112(.dina(n8367), .dinb(n364), .dout(n8368));
  jxor g08113(.dina(n8368), .dinb(n8360), .dout(n8369));
  jxor g08114(.dina(n8369), .dinb(n8129), .dout(n8370));
  jand g08115(.dina(b55 ), .dinb(b54 ), .dout(n8371));
  jand g08116(.dina(n8107), .dinb(n8106), .dout(n8372));
  jor  g08117(.dina(n8372), .dinb(n8371), .dout(n8373));
  jxor g08118(.dina(b56 ), .dinb(b55 ), .dout(n8374));
  jnot g08119(.din(n8374), .dout(n8375));
  jxor g08120(.dina(n8375), .dinb(n8373), .dout(n8376));
  jor  g08121(.dina(n8376), .dinb(n296), .dout(n8377));
  jnot g08122(.din(b56 ), .dout(n8378));
  jor  g08123(.dina(n264), .dinb(n8378), .dout(n8379));
  jor  g08124(.dina(n280), .dinb(n7846), .dout(n8380));
  jor  g08125(.dina(n294), .dinb(n8111), .dout(n8381));
  jand g08126(.dina(n8381), .dinb(n8380), .dout(n8382));
  jand g08127(.dina(n8382), .dinb(n8379), .dout(n8383));
  jand g08128(.dina(n8383), .dinb(n8377), .dout(n8384));
  jxor g08129(.dina(n8384), .dinb(n278), .dout(n8385));
  jxor g08130(.dina(n8385), .dinb(n8370), .dout(n8386));
  jxor g08131(.dina(n8386), .dinb(n8124), .dout(f56 ));
  jnot g08132(.din(n8385), .dout(n8388));
  jor  g08133(.dina(n8388), .dinb(n8370), .dout(n8389));
  jor  g08134(.dina(n8386), .dinb(n8124), .dout(n8390));
  jand g08135(.dina(n8390), .dinb(n8389), .dout(n8391));
  jand g08136(.dina(n8368), .dinb(n8360), .dout(n8392));
  jnot g08137(.din(n8392), .dout(n8393));
  jnot g08138(.din(n8369), .dout(n8394));
  jor  g08139(.dina(n8394), .dinb(n8129), .dout(n8395));
  jand g08140(.dina(n8395), .dinb(n8393), .dout(n8396));
  jnot g08141(.din(n8349), .dout(n8397));
  jand g08142(.dina(n8357), .dinb(n8397), .dout(n8398));
  jand g08143(.dina(n8359), .dinb(n8132), .dout(n8399));
  jor  g08144(.dina(n8399), .dinb(n8398), .dout(n8400));
  jand g08145(.dina(n8347), .dinb(n8339), .dout(n8401));
  jnot g08146(.din(n8136), .dout(n8402));
  jand g08147(.dina(n8348), .dinb(n8402), .dout(n8403));
  jor  g08148(.dina(n8403), .dinb(n8401), .dout(n8404));
  jand g08149(.dina(n8337), .dinb(n8329), .dout(n8405));
  jand g08150(.dina(n8338), .dinb(n8139), .dout(n8406));
  jor  g08151(.dina(n8406), .dinb(n8405), .dout(n8407));
  jand g08152(.dina(n8327), .dinb(n8319), .dout(n8408));
  jand g08153(.dina(n8328), .dinb(n8142), .dout(n8409));
  jor  g08154(.dina(n8409), .dinb(n8408), .dout(n8410));
  jand g08155(.dina(n8317), .dinb(n8309), .dout(n8411));
  jand g08156(.dina(n8318), .dinb(n8145), .dout(n8412));
  jor  g08157(.dina(n8412), .dinb(n8411), .dout(n8413));
  jand g08158(.dina(n8307), .dinb(n8299), .dout(n8414));
  jand g08159(.dina(n8308), .dinb(n8148), .dout(n8415));
  jor  g08160(.dina(n8415), .dinb(n8414), .dout(n8416));
  jand g08161(.dina(n8297), .dinb(n8289), .dout(n8417));
  jand g08162(.dina(n8298), .dinb(n8151), .dout(n8418));
  jor  g08163(.dina(n8418), .dinb(n8417), .dout(n8419));
  jand g08164(.dina(n8287), .dinb(n8279), .dout(n8420));
  jand g08165(.dina(n8288), .dinb(n8154), .dout(n8421));
  jor  g08166(.dina(n8421), .dinb(n8420), .dout(n8422));
  jand g08167(.dina(n8277), .dinb(n8269), .dout(n8423));
  jand g08168(.dina(n8278), .dinb(n8157), .dout(n8424));
  jor  g08169(.dina(n8424), .dinb(n8423), .dout(n8425));
  jand g08170(.dina(n8267), .dinb(n8259), .dout(n8426));
  jand g08171(.dina(n8268), .dinb(n8160), .dout(n8427));
  jor  g08172(.dina(n8427), .dinb(n8426), .dout(n8428));
  jand g08173(.dina(n8257), .dinb(n8249), .dout(n8429));
  jand g08174(.dina(n8258), .dinb(n8163), .dout(n8430));
  jor  g08175(.dina(n8430), .dinb(n8429), .dout(n8431));
  jand g08176(.dina(n8247), .dinb(n8239), .dout(n8432));
  jand g08177(.dina(n8248), .dinb(n8166), .dout(n8433));
  jor  g08178(.dina(n8433), .dinb(n8432), .dout(n8434));
  jand g08179(.dina(n8237), .dinb(n8229), .dout(n8435));
  jand g08180(.dina(n8238), .dinb(n8169), .dout(n8436));
  jor  g08181(.dina(n8436), .dinb(n8435), .dout(n8437));
  jand g08182(.dina(n8227), .dinb(n8219), .dout(n8438));
  jand g08183(.dina(n8228), .dinb(n8172), .dout(n8439));
  jor  g08184(.dina(n8439), .dinb(n8438), .dout(n8440));
  jand g08185(.dina(n8217), .dinb(n8209), .dout(n8441));
  jand g08186(.dina(n8218), .dinb(n8177), .dout(n8442));
  jor  g08187(.dina(n8442), .dinb(n8441), .dout(n8443));
  jor  g08188(.dina(n8207), .dinb(n8199), .dout(n8444));
  jand g08189(.dina(n8208), .dinb(n8182), .dout(n8445));
  jnot g08190(.din(n8445), .dout(n8446));
  jand g08191(.dina(n8446), .dinb(n8444), .dout(n8447));
  jnot g08192(.din(n8447), .dout(n8448));
  jor  g08193(.dina(n8196), .dinb(n8192), .dout(n8449));
  jxor g08194(.dina(a57 ), .dinb(a56 ), .dout(n8450));
  jand g08195(.dina(n8450), .dinb(b0 ), .dout(n8451));
  jnot g08196(.din(n8451), .dout(n8452));
  jxor g08197(.dina(n8452), .dinb(n8449), .dout(n8453));
  jnot g08198(.din(n7925), .dout(n8454));
  jor  g08199(.dina(n8454), .dinb(n303), .dout(n8455));
  jor  g08200(.dina(n8185), .dinb(n305), .dout(n8456));
  jnot g08201(.din(n7918), .dout(n8457));
  jor  g08202(.dina(n8457), .dinb(n301), .dout(n8458));
  jnot g08203(.din(n7922), .dout(n8459));
  jor  g08204(.dina(n8459), .dinb(n293), .dout(n8460));
  jand g08205(.dina(n8460), .dinb(n8458), .dout(n8461));
  jand g08206(.dina(n8461), .dinb(n8456), .dout(n8462));
  jand g08207(.dina(n8462), .dinb(n8455), .dout(n8463));
  jxor g08208(.dina(n8463), .dinb(n7929), .dout(n8464));
  jxor g08209(.dina(n8464), .dinb(n8453), .dout(n8465));
  jnot g08210(.din(n8465), .dout(n8466));
  jor  g08211(.dina(n7660), .dinb(n412), .dout(n8467));
  jor  g08212(.dina(n7662), .dinb(n415), .dout(n8468));
  jor  g08213(.dina(n7415), .dinb(n340), .dout(n8469));
  jand g08214(.dina(n8469), .dinb(n8468), .dout(n8470));
  jor  g08215(.dina(n7657), .dinb(n377), .dout(n8471));
  jand g08216(.dina(n8471), .dinb(n8470), .dout(n8472));
  jand g08217(.dina(n8472), .dinb(n8467), .dout(n8473));
  jxor g08218(.dina(n8473), .dinb(a53 ), .dout(n8474));
  jxor g08219(.dina(n8474), .dinb(n8466), .dout(n8475));
  jxor g08220(.dina(n8475), .dinb(n8448), .dout(n8476));
  jor  g08221(.dina(n6914), .dinb(n570), .dout(n8477));
  jor  g08222(.dina(n6673), .dinb(n469), .dout(n8478));
  jor  g08223(.dina(n6911), .dinb(n519), .dout(n8479));
  jor  g08224(.dina(n6916), .dinb(n572), .dout(n8480));
  jand g08225(.dina(n8480), .dinb(n8479), .dout(n8481));
  jand g08226(.dina(n8481), .dinb(n8478), .dout(n8482));
  jand g08227(.dina(n8482), .dinb(n8477), .dout(n8483));
  jxor g08228(.dina(n8483), .dinb(n6443), .dout(n8484));
  jxor g08229(.dina(n8484), .dinb(n8476), .dout(n8485));
  jxor g08230(.dina(n8485), .dinb(n8443), .dout(n8486));
  jor  g08231(.dina(n6207), .dinb(n770), .dout(n8487));
  jor  g08232(.dina(n5975), .dinb(n637), .dout(n8488));
  jor  g08233(.dina(n6210), .dinb(n704), .dout(n8489));
  jor  g08234(.dina(n6205), .dinb(n772), .dout(n8490));
  jand g08235(.dina(n8490), .dinb(n8489), .dout(n8491));
  jand g08236(.dina(n8491), .dinb(n8488), .dout(n8492));
  jand g08237(.dina(n8492), .dinb(n8487), .dout(n8493));
  jxor g08238(.dina(n8493), .dinb(n5759), .dout(n8494));
  jxor g08239(.dina(n8494), .dinb(n8486), .dout(n8495));
  jxor g08240(.dina(n8495), .dinb(n8440), .dout(n8496));
  jor  g08241(.dina(n5537), .dinb(n1016), .dout(n8497));
  jor  g08242(.dina(n5315), .dinb(n852), .dout(n8498));
  jor  g08243(.dina(n5534), .dinb(n934), .dout(n8499));
  jor  g08244(.dina(n5539), .dinb(n1018), .dout(n8500));
  jand g08245(.dina(n8500), .dinb(n8499), .dout(n8501));
  jand g08246(.dina(n8501), .dinb(n8498), .dout(n8502));
  jand g08247(.dina(n8502), .dinb(n8497), .dout(n8503));
  jxor g08248(.dina(n8503), .dinb(n5111), .dout(n8504));
  jxor g08249(.dina(n8504), .dinb(n8496), .dout(n8505));
  jxor g08250(.dina(n8505), .dinb(n8437), .dout(n8506));
  jor  g08251(.dina(n4902), .dinb(n1305), .dout(n8507));
  jor  g08252(.dina(n4696), .dinb(n1114), .dout(n8508));
  jor  g08253(.dina(n4904), .dinb(n1211), .dout(n8509));
  jor  g08254(.dina(n4899), .dinb(n1307), .dout(n8510));
  jand g08255(.dina(n8510), .dinb(n8509), .dout(n8511));
  jand g08256(.dina(n8511), .dinb(n8508), .dout(n8512));
  jand g08257(.dina(n8512), .dinb(n8507), .dout(n8513));
  jxor g08258(.dina(n8513), .dinb(n4505), .dout(n8514));
  jxor g08259(.dina(n8514), .dinb(n8506), .dout(n8515));
  jxor g08260(.dina(n8515), .dinb(n8434), .dout(n8516));
  jor  g08261(.dina(n4305), .dinb(n1635), .dout(n8517));
  jor  g08262(.dina(n4116), .dinb(n1416), .dout(n8518));
  jor  g08263(.dina(n4303), .dinb(n1637), .dout(n8519));
  jor  g08264(.dina(n4308), .dinb(n1527), .dout(n8520));
  jand g08265(.dina(n8520), .dinb(n8519), .dout(n8521));
  jand g08266(.dina(n8521), .dinb(n8518), .dout(n8522));
  jand g08267(.dina(n8522), .dinb(n8517), .dout(n8523));
  jxor g08268(.dina(n8523), .dinb(n3938), .dout(n8524));
  jxor g08269(.dina(n8524), .dinb(n8516), .dout(n8525));
  jxor g08270(.dina(n8525), .dinb(n8431), .dout(n8526));
  jor  g08271(.dina(n3751), .dinb(n2005), .dout(n8527));
  jor  g08272(.dina(n3574), .dinb(n1759), .dout(n8528));
  jor  g08273(.dina(n3754), .dinb(n1881), .dout(n8529));
  jor  g08274(.dina(n3749), .dinb(n2007), .dout(n8530));
  jand g08275(.dina(n8530), .dinb(n8529), .dout(n8531));
  jand g08276(.dina(n8531), .dinb(n8528), .dout(n8532));
  jand g08277(.dina(n8532), .dinb(n8527), .dout(n8533));
  jxor g08278(.dina(n8533), .dinb(n3410), .dout(n8534));
  jxor g08279(.dina(n8534), .dinb(n8526), .dout(n8535));
  jxor g08280(.dina(n8535), .dinb(n8428), .dout(n8536));
  jor  g08281(.dina(n3239), .dinb(n2413), .dout(n8537));
  jor  g08282(.dina(n3072), .dinb(n2142), .dout(n8538));
  jor  g08283(.dina(n3242), .dinb(n2279), .dout(n8539));
  jor  g08284(.dina(n3237), .dinb(n2415), .dout(n8540));
  jand g08285(.dina(n8540), .dinb(n8539), .dout(n8541));
  jand g08286(.dina(n8541), .dinb(n8538), .dout(n8542));
  jand g08287(.dina(n8542), .dinb(n8537), .dout(n8543));
  jxor g08288(.dina(n8543), .dinb(n2918), .dout(n8544));
  jxor g08289(.dina(n8544), .dinb(n8536), .dout(n8545));
  jxor g08290(.dina(n8545), .dinb(n8425), .dout(n8546));
  jor  g08291(.dina(n2860), .dinb(n2764), .dout(n8547));
  jor  g08292(.dina(n2609), .dinb(n2563), .dout(n8548));
  jor  g08293(.dina(n2761), .dinb(n2862), .dout(n8549));
  jor  g08294(.dina(n2766), .dinb(n2713), .dout(n8550));
  jand g08295(.dina(n8550), .dinb(n8549), .dout(n8551));
  jand g08296(.dina(n8551), .dinb(n8548), .dout(n8552));
  jand g08297(.dina(n8552), .dinb(n8547), .dout(n8553));
  jxor g08298(.dina(n8553), .dinb(n2468), .dout(n8554));
  jxor g08299(.dina(n8554), .dinb(n8546), .dout(n8555));
  jxor g08300(.dina(n8555), .dinb(n8422), .dout(n8556));
  jor  g08301(.dina(n3346), .dinb(n2324), .dout(n8557));
  jor  g08302(.dina(n2186), .dinb(n3023), .dout(n8558));
  jor  g08303(.dina(n2321), .dinb(n3186), .dout(n8559));
  jor  g08304(.dina(n2326), .dinb(n3348), .dout(n8560));
  jand g08305(.dina(n8560), .dinb(n8559), .dout(n8561));
  jand g08306(.dina(n8561), .dinb(n8558), .dout(n8562));
  jand g08307(.dina(n8562), .dinb(n8557), .dout(n8563));
  jxor g08308(.dina(n8563), .dinb(n2057), .dout(n8564));
  jxor g08309(.dina(n8564), .dinb(n8556), .dout(n8565));
  jxor g08310(.dina(n8565), .dinb(n8419), .dout(n8566));
  jor  g08311(.dina(n3871), .dinb(n1921), .dout(n8567));
  jor  g08312(.dina(n1806), .dinb(n3522), .dout(n8568));
  jor  g08313(.dina(n1918), .dinb(n3698), .dout(n8569));
  jor  g08314(.dina(n1923), .dinb(n3873), .dout(n8570));
  jand g08315(.dina(n8570), .dinb(n8569), .dout(n8571));
  jand g08316(.dina(n8571), .dinb(n8568), .dout(n8572));
  jand g08317(.dina(n8572), .dinb(n8567), .dout(n8573));
  jxor g08318(.dina(n8573), .dinb(n1687), .dout(n8574));
  jxor g08319(.dina(n8574), .dinb(n8566), .dout(n8575));
  jxor g08320(.dina(n8575), .dinb(n8416), .dout(n8576));
  jor  g08321(.dina(n4435), .dinb(n1569), .dout(n8577));
  jor  g08322(.dina(n1453), .dinb(n4060), .dout(n8578));
  jor  g08323(.dina(n1566), .dinb(n4249), .dout(n8579));
  jor  g08324(.dina(n1571), .dinb(n4437), .dout(n8580));
  jand g08325(.dina(n8580), .dinb(n8579), .dout(n8581));
  jand g08326(.dina(n8581), .dinb(n8578), .dout(n8582));
  jand g08327(.dina(n8582), .dinb(n8577), .dout(n8583));
  jxor g08328(.dina(n8583), .dinb(n1351), .dout(n8584));
  jxor g08329(.dina(n8584), .dinb(n8576), .dout(n8585));
  jxor g08330(.dina(n8585), .dinb(n8413), .dout(n8586));
  jor  g08331(.dina(n5038), .dinb(n1248), .dout(n8587));
  jor  g08332(.dina(n1147), .dinb(n4637), .dout(n8588));
  jor  g08333(.dina(n1246), .dinb(n5040), .dout(n8589));
  jor  g08334(.dina(n1251), .dinb(n4839), .dout(n8590));
  jand g08335(.dina(n8590), .dinb(n8589), .dout(n8591));
  jand g08336(.dina(n8591), .dinb(n8588), .dout(n8592));
  jand g08337(.dina(n8592), .dinb(n8587), .dout(n8593));
  jxor g08338(.dina(n8593), .dinb(n1061), .dout(n8594));
  jxor g08339(.dina(n8594), .dinb(n8586), .dout(n8595));
  jxor g08340(.dina(n8595), .dinb(n8410), .dout(n8596));
  jor  g08341(.dina(n5683), .dinb(n970), .dout(n8597));
  jor  g08342(.dina(n880), .dinb(n5253), .dout(n8598));
  jor  g08343(.dina(n967), .dinb(n5469), .dout(n8599));
  jor  g08344(.dina(n972), .dinb(n5685), .dout(n8600));
  jand g08345(.dina(n8600), .dinb(n8599), .dout(n8601));
  jand g08346(.dina(n8601), .dinb(n8598), .dout(n8602));
  jand g08347(.dina(n8602), .dinb(n8597), .dout(n8603));
  jxor g08348(.dina(n8603), .dinb(n810), .dout(n8604));
  jxor g08349(.dina(n8604), .dinb(n8596), .dout(n8605));
  jxor g08350(.dina(n8605), .dinb(n8407), .dout(n8606));
  jor  g08351(.dina(n6364), .dinb(n728), .dout(n8607));
  jor  g08352(.dina(n660), .dinb(n5911), .dout(n8608));
  jor  g08353(.dina(n726), .dinb(n6366), .dout(n8609));
  jor  g08354(.dina(n731), .dinb(n6139), .dout(n8610));
  jand g08355(.dina(n8610), .dinb(n8609), .dout(n8611));
  jand g08356(.dina(n8611), .dinb(n8608), .dout(n8612));
  jand g08357(.dina(n8612), .dinb(n8607), .dout(n8613));
  jxor g08358(.dina(n8613), .dinb(n606), .dout(n8614));
  jxor g08359(.dina(n8614), .dinb(n8606), .dout(n8615));
  jxor g08360(.dina(n8615), .dinb(n8404), .dout(n8616));
  jor  g08361(.dina(n7084), .dinb(n544), .dout(n8617));
  jor  g08362(.dina(n486), .dinb(n6605), .dout(n8618));
  jor  g08363(.dina(n547), .dinb(n6846), .dout(n8619));
  jor  g08364(.dina(n542), .dinb(n7086), .dout(n8620));
  jand g08365(.dina(n8620), .dinb(n8619), .dout(n8621));
  jand g08366(.dina(n8621), .dinb(n8618), .dout(n8622));
  jand g08367(.dina(n8622), .dinb(n8617), .dout(n8623));
  jxor g08368(.dina(n8623), .dinb(n446), .dout(n8624));
  jxor g08369(.dina(n8624), .dinb(n8616), .dout(n8625));
  jxor g08370(.dina(n8625), .dinb(n8400), .dout(n8626));
  jor  g08371(.dina(n7844), .dinb(n397), .dout(n8627));
  jor  g08372(.dina(n354), .dinb(n7338), .dout(n8628));
  jor  g08373(.dina(n399), .dinb(n7846), .dout(n8629));
  jor  g08374(.dina(n394), .dinb(n7590), .dout(n8630));
  jand g08375(.dina(n8630), .dinb(n8629), .dout(n8631));
  jand g08376(.dina(n8631), .dinb(n8628), .dout(n8632));
  jand g08377(.dina(n8632), .dinb(n8627), .dout(n8633));
  jxor g08378(.dina(n8633), .dinb(n364), .dout(n8634));
  jxor g08379(.dina(n8634), .dinb(n8626), .dout(n8635));
  jxor g08380(.dina(n8635), .dinb(n8396), .dout(n8636));
  jand g08381(.dina(b56 ), .dinb(b55 ), .dout(n8637));
  jand g08382(.dina(n8374), .dinb(n8373), .dout(n8638));
  jor  g08383(.dina(n8638), .dinb(n8637), .dout(n8639));
  jxor g08384(.dina(b57 ), .dinb(b56 ), .dout(n8640));
  jnot g08385(.din(n8640), .dout(n8641));
  jxor g08386(.dina(n8641), .dinb(n8639), .dout(n8642));
  jor  g08387(.dina(n8642), .dinb(n296), .dout(n8643));
  jnot g08388(.din(b57 ), .dout(n8644));
  jor  g08389(.dina(n264), .dinb(n8644), .dout(n8645));
  jor  g08390(.dina(n280), .dinb(n8111), .dout(n8646));
  jor  g08391(.dina(n294), .dinb(n8378), .dout(n8647));
  jand g08392(.dina(n8647), .dinb(n8646), .dout(n8648));
  jand g08393(.dina(n8648), .dinb(n8645), .dout(n8649));
  jand g08394(.dina(n8649), .dinb(n8643), .dout(n8650));
  jxor g08395(.dina(n8650), .dinb(n278), .dout(n8651));
  jxor g08396(.dina(n8651), .dinb(n8636), .dout(n8652));
  jxor g08397(.dina(n8652), .dinb(n8391), .dout(f57 ));
  jnot g08398(.din(n8651), .dout(n8654));
  jor  g08399(.dina(n8654), .dinb(n8636), .dout(n8655));
  jor  g08400(.dina(n8652), .dinb(n8391), .dout(n8656));
  jand g08401(.dina(n8656), .dinb(n8655), .dout(n8657));
  jand g08402(.dina(n8634), .dinb(n8626), .dout(n8658));
  jnot g08403(.din(n8658), .dout(n8659));
  jnot g08404(.din(n8635), .dout(n8660));
  jor  g08405(.dina(n8660), .dinb(n8396), .dout(n8661));
  jand g08406(.dina(n8661), .dinb(n8659), .dout(n8662));
  jand g08407(.dina(n8624), .dinb(n8616), .dout(n8663));
  jand g08408(.dina(n8625), .dinb(n8400), .dout(n8664));
  jor  g08409(.dina(n8664), .dinb(n8663), .dout(n8665));
  jand g08410(.dina(n8614), .dinb(n8606), .dout(n8666));
  jand g08411(.dina(n8615), .dinb(n8404), .dout(n8667));
  jor  g08412(.dina(n8667), .dinb(n8666), .dout(n8668));
  jand g08413(.dina(n8604), .dinb(n8596), .dout(n8669));
  jand g08414(.dina(n8605), .dinb(n8407), .dout(n8670));
  jor  g08415(.dina(n8670), .dinb(n8669), .dout(n8671));
  jand g08416(.dina(n8594), .dinb(n8586), .dout(n8672));
  jand g08417(.dina(n8595), .dinb(n8410), .dout(n8673));
  jor  g08418(.dina(n8673), .dinb(n8672), .dout(n8674));
  jand g08419(.dina(n8584), .dinb(n8576), .dout(n8675));
  jand g08420(.dina(n8585), .dinb(n8413), .dout(n8676));
  jor  g08421(.dina(n8676), .dinb(n8675), .dout(n8677));
  jand g08422(.dina(n8574), .dinb(n8566), .dout(n8678));
  jand g08423(.dina(n8575), .dinb(n8416), .dout(n8679));
  jor  g08424(.dina(n8679), .dinb(n8678), .dout(n8680));
  jand g08425(.dina(n8564), .dinb(n8556), .dout(n8681));
  jand g08426(.dina(n8565), .dinb(n8419), .dout(n8682));
  jor  g08427(.dina(n8682), .dinb(n8681), .dout(n8683));
  jand g08428(.dina(n8554), .dinb(n8546), .dout(n8684));
  jand g08429(.dina(n8555), .dinb(n8422), .dout(n8685));
  jor  g08430(.dina(n8685), .dinb(n8684), .dout(n8686));
  jand g08431(.dina(n8544), .dinb(n8536), .dout(n8687));
  jand g08432(.dina(n8545), .dinb(n8425), .dout(n8688));
  jor  g08433(.dina(n8688), .dinb(n8687), .dout(n8689));
  jand g08434(.dina(n8534), .dinb(n8526), .dout(n8690));
  jand g08435(.dina(n8535), .dinb(n8428), .dout(n8691));
  jor  g08436(.dina(n8691), .dinb(n8690), .dout(n8692));
  jand g08437(.dina(n8524), .dinb(n8516), .dout(n8693));
  jand g08438(.dina(n8525), .dinb(n8431), .dout(n8694));
  jor  g08439(.dina(n8694), .dinb(n8693), .dout(n8695));
  jand g08440(.dina(n8514), .dinb(n8506), .dout(n8696));
  jand g08441(.dina(n8515), .dinb(n8434), .dout(n8697));
  jor  g08442(.dina(n8697), .dinb(n8696), .dout(n8698));
  jand g08443(.dina(n8504), .dinb(n8496), .dout(n8699));
  jand g08444(.dina(n8505), .dinb(n8437), .dout(n8700));
  jor  g08445(.dina(n8700), .dinb(n8699), .dout(n8701));
  jand g08446(.dina(n8494), .dinb(n8486), .dout(n8702));
  jand g08447(.dina(n8495), .dinb(n8440), .dout(n8703));
  jor  g08448(.dina(n8703), .dinb(n8702), .dout(n8704));
  jand g08449(.dina(n8484), .dinb(n8476), .dout(n8705));
  jand g08450(.dina(n8485), .dinb(n8443), .dout(n8706));
  jor  g08451(.dina(n8706), .dinb(n8705), .dout(n8707));
  jor  g08452(.dina(n8474), .dinb(n8466), .dout(n8708));
  jand g08453(.dina(n8475), .dinb(n8448), .dout(n8709));
  jnot g08454(.din(n8709), .dout(n8710));
  jand g08455(.dina(n8710), .dinb(n8708), .dout(n8711));
  jnot g08456(.din(n8711), .dout(n8712));
  jnot g08457(.din(n8449), .dout(n8713));
  jand g08458(.dina(n8451), .dinb(n8713), .dout(n8714));
  jand g08459(.dina(n8464), .dinb(n8453), .dout(n8715));
  jor  g08460(.dina(n8715), .dinb(n8714), .dout(n8716));
  jxor g08461(.dina(a59 ), .dinb(a58 ), .dout(n8717));
  jand g08462(.dina(n8717), .dinb(n8450), .dout(n8718));
  jand g08463(.dina(n8718), .dinb(n259), .dout(n8719));
  jnot g08464(.din(n8450), .dout(n8720));
  jxor g08465(.dina(a58 ), .dinb(a57 ), .dout(n8721));
  jand g08466(.dina(n8721), .dinb(n8720), .dout(n8722));
  jand g08467(.dina(n8722), .dinb(b0 ), .dout(n8723));
  jnot g08468(.din(n8717), .dout(n8724));
  jand g08469(.dina(n8724), .dinb(n8450), .dout(n8725));
  jand g08470(.dina(n8725), .dinb(b1 ), .dout(n8726));
  jor  g08471(.dina(n8726), .dinb(n8723), .dout(n8727));
  jor  g08472(.dina(n8727), .dinb(n8719), .dout(n8728));
  jnot g08473(.din(a59 ), .dout(n8729));
  jor  g08474(.dina(n8452), .dinb(n8729), .dout(n8730));
  jxor g08475(.dina(n8730), .dinb(n8728), .dout(n8731));
  jor  g08476(.dina(n8457), .dinb(n337), .dout(n8732));
  jor  g08477(.dina(n8459), .dinb(n303), .dout(n8733));
  jor  g08478(.dina(n8185), .dinb(n293), .dout(n8734));
  jand g08479(.dina(n8734), .dinb(n8733), .dout(n8735));
  jor  g08480(.dina(n8454), .dinb(n340), .dout(n8736));
  jand g08481(.dina(n8736), .dinb(n8735), .dout(n8737));
  jand g08482(.dina(n8737), .dinb(n8732), .dout(n8738));
  jxor g08483(.dina(n8738), .dinb(a56 ), .dout(n8739));
  jxor g08484(.dina(n8739), .dinb(n8731), .dout(n8740));
  jxor g08485(.dina(n8740), .dinb(n8716), .dout(n8741));
  jnot g08486(.din(n8741), .dout(n8742));
  jor  g08487(.dina(n7660), .dinb(n466), .dout(n8743));
  jor  g08488(.dina(n7662), .dinb(n469), .dout(n8744));
  jor  g08489(.dina(n7415), .dinb(n377), .dout(n8745));
  jand g08490(.dina(n8745), .dinb(n8744), .dout(n8746));
  jor  g08491(.dina(n7657), .dinb(n415), .dout(n8747));
  jand g08492(.dina(n8747), .dinb(n8746), .dout(n8748));
  jand g08493(.dina(n8748), .dinb(n8743), .dout(n8749));
  jxor g08494(.dina(n8749), .dinb(a53 ), .dout(n8750));
  jxor g08495(.dina(n8750), .dinb(n8742), .dout(n8751));
  jxor g08496(.dina(n8751), .dinb(n8712), .dout(n8752));
  jor  g08497(.dina(n6914), .dinb(n635), .dout(n8753));
  jor  g08498(.dina(n6673), .dinb(n519), .dout(n8754));
  jor  g08499(.dina(n6911), .dinb(n572), .dout(n8755));
  jor  g08500(.dina(n6916), .dinb(n637), .dout(n8756));
  jand g08501(.dina(n8756), .dinb(n8755), .dout(n8757));
  jand g08502(.dina(n8757), .dinb(n8754), .dout(n8758));
  jand g08503(.dina(n8758), .dinb(n8753), .dout(n8759));
  jxor g08504(.dina(n8759), .dinb(n6443), .dout(n8760));
  jxor g08505(.dina(n8760), .dinb(n8752), .dout(n8761));
  jxor g08506(.dina(n8761), .dinb(n8707), .dout(n8762));
  jor  g08507(.dina(n6207), .dinb(n850), .dout(n8763));
  jor  g08508(.dina(n5975), .dinb(n704), .dout(n8764));
  jor  g08509(.dina(n6210), .dinb(n772), .dout(n8765));
  jor  g08510(.dina(n6205), .dinb(n852), .dout(n8766));
  jand g08511(.dina(n8766), .dinb(n8765), .dout(n8767));
  jand g08512(.dina(n8767), .dinb(n8764), .dout(n8768));
  jand g08513(.dina(n8768), .dinb(n8763), .dout(n8769));
  jxor g08514(.dina(n8769), .dinb(n5759), .dout(n8770));
  jxor g08515(.dina(n8770), .dinb(n8762), .dout(n8771));
  jxor g08516(.dina(n8771), .dinb(n8704), .dout(n8772));
  jor  g08517(.dina(n5537), .dinb(n1112), .dout(n8773));
  jor  g08518(.dina(n5315), .dinb(n934), .dout(n8774));
  jor  g08519(.dina(n5539), .dinb(n1114), .dout(n8775));
  jor  g08520(.dina(n5534), .dinb(n1018), .dout(n8776));
  jand g08521(.dina(n8776), .dinb(n8775), .dout(n8777));
  jand g08522(.dina(n8777), .dinb(n8774), .dout(n8778));
  jand g08523(.dina(n8778), .dinb(n8773), .dout(n8779));
  jxor g08524(.dina(n8779), .dinb(n5111), .dout(n8780));
  jxor g08525(.dina(n8780), .dinb(n8772), .dout(n8781));
  jxor g08526(.dina(n8781), .dinb(n8701), .dout(n8782));
  jor  g08527(.dina(n4902), .dinb(n1414), .dout(n8783));
  jor  g08528(.dina(n4696), .dinb(n1211), .dout(n8784));
  jor  g08529(.dina(n4899), .dinb(n1416), .dout(n8785));
  jor  g08530(.dina(n4904), .dinb(n1307), .dout(n8786));
  jand g08531(.dina(n8786), .dinb(n8785), .dout(n8787));
  jand g08532(.dina(n8787), .dinb(n8784), .dout(n8788));
  jand g08533(.dina(n8788), .dinb(n8783), .dout(n8789));
  jxor g08534(.dina(n8789), .dinb(n4505), .dout(n8790));
  jxor g08535(.dina(n8790), .dinb(n8782), .dout(n8791));
  jxor g08536(.dina(n8791), .dinb(n8698), .dout(n8792));
  jor  g08537(.dina(n4305), .dinb(n1757), .dout(n8793));
  jor  g08538(.dina(n4116), .dinb(n1527), .dout(n8794));
  jor  g08539(.dina(n4308), .dinb(n1637), .dout(n8795));
  jor  g08540(.dina(n4303), .dinb(n1759), .dout(n8796));
  jand g08541(.dina(n8796), .dinb(n8795), .dout(n8797));
  jand g08542(.dina(n8797), .dinb(n8794), .dout(n8798));
  jand g08543(.dina(n8798), .dinb(n8793), .dout(n8799));
  jxor g08544(.dina(n8799), .dinb(n3938), .dout(n8800));
  jxor g08545(.dina(n8800), .dinb(n8792), .dout(n8801));
  jxor g08546(.dina(n8801), .dinb(n8695), .dout(n8802));
  jor  g08547(.dina(n3751), .dinb(n2140), .dout(n8803));
  jor  g08548(.dina(n3574), .dinb(n1881), .dout(n8804));
  jor  g08549(.dina(n3754), .dinb(n2007), .dout(n8805));
  jor  g08550(.dina(n3749), .dinb(n2142), .dout(n8806));
  jand g08551(.dina(n8806), .dinb(n8805), .dout(n8807));
  jand g08552(.dina(n8807), .dinb(n8804), .dout(n8808));
  jand g08553(.dina(n8808), .dinb(n8803), .dout(n8809));
  jxor g08554(.dina(n8809), .dinb(n3410), .dout(n8810));
  jxor g08555(.dina(n8810), .dinb(n8802), .dout(n8811));
  jxor g08556(.dina(n8811), .dinb(n8692), .dout(n8812));
  jor  g08557(.dina(n3239), .dinb(n2561), .dout(n8813));
  jor  g08558(.dina(n3072), .dinb(n2279), .dout(n8814));
  jor  g08559(.dina(n3237), .dinb(n2563), .dout(n8815));
  jor  g08560(.dina(n3242), .dinb(n2415), .dout(n8816));
  jand g08561(.dina(n8816), .dinb(n8815), .dout(n8817));
  jand g08562(.dina(n8817), .dinb(n8814), .dout(n8818));
  jand g08563(.dina(n8818), .dinb(n8813), .dout(n8819));
  jxor g08564(.dina(n8819), .dinb(n2918), .dout(n8820));
  jxor g08565(.dina(n8820), .dinb(n8812), .dout(n8821));
  jxor g08566(.dina(n8821), .dinb(n8689), .dout(n8822));
  jor  g08567(.dina(n3021), .dinb(n2764), .dout(n8823));
  jor  g08568(.dina(n2609), .dinb(n2713), .dout(n8824));
  jor  g08569(.dina(n2761), .dinb(n3023), .dout(n8825));
  jor  g08570(.dina(n2766), .dinb(n2862), .dout(n8826));
  jand g08571(.dina(n8826), .dinb(n8825), .dout(n8827));
  jand g08572(.dina(n8827), .dinb(n8824), .dout(n8828));
  jand g08573(.dina(n8828), .dinb(n8823), .dout(n8829));
  jxor g08574(.dina(n8829), .dinb(n2468), .dout(n8830));
  jxor g08575(.dina(n8830), .dinb(n8822), .dout(n8831));
  jxor g08576(.dina(n8831), .dinb(n8686), .dout(n8832));
  jor  g08577(.dina(n3520), .dinb(n2324), .dout(n8833));
  jor  g08578(.dina(n2186), .dinb(n3186), .dout(n8834));
  jor  g08579(.dina(n2321), .dinb(n3348), .dout(n8835));
  jor  g08580(.dina(n2326), .dinb(n3522), .dout(n8836));
  jand g08581(.dina(n8836), .dinb(n8835), .dout(n8837));
  jand g08582(.dina(n8837), .dinb(n8834), .dout(n8838));
  jand g08583(.dina(n8838), .dinb(n8833), .dout(n8839));
  jxor g08584(.dina(n8839), .dinb(n2057), .dout(n8840));
  jxor g08585(.dina(n8840), .dinb(n8832), .dout(n8841));
  jxor g08586(.dina(n8841), .dinb(n8683), .dout(n8842));
  jor  g08587(.dina(n4058), .dinb(n1921), .dout(n8843));
  jor  g08588(.dina(n1806), .dinb(n3698), .dout(n8844));
  jor  g08589(.dina(n1923), .dinb(n4060), .dout(n8845));
  jor  g08590(.dina(n1918), .dinb(n3873), .dout(n8846));
  jand g08591(.dina(n8846), .dinb(n8845), .dout(n8847));
  jand g08592(.dina(n8847), .dinb(n8844), .dout(n8848));
  jand g08593(.dina(n8848), .dinb(n8843), .dout(n8849));
  jxor g08594(.dina(n8849), .dinb(n1687), .dout(n8850));
  jxor g08595(.dina(n8850), .dinb(n8842), .dout(n8851));
  jxor g08596(.dina(n8851), .dinb(n8680), .dout(n8852));
  jor  g08597(.dina(n4635), .dinb(n1569), .dout(n8853));
  jor  g08598(.dina(n1453), .dinb(n4249), .dout(n8854));
  jor  g08599(.dina(n1566), .dinb(n4437), .dout(n8855));
  jor  g08600(.dina(n1571), .dinb(n4637), .dout(n8856));
  jand g08601(.dina(n8856), .dinb(n8855), .dout(n8857));
  jand g08602(.dina(n8857), .dinb(n8854), .dout(n8858));
  jand g08603(.dina(n8858), .dinb(n8853), .dout(n8859));
  jxor g08604(.dina(n8859), .dinb(n1351), .dout(n8860));
  jxor g08605(.dina(n8860), .dinb(n8852), .dout(n8861));
  jxor g08606(.dina(n8861), .dinb(n8677), .dout(n8862));
  jor  g08607(.dina(n5251), .dinb(n1248), .dout(n8863));
  jor  g08608(.dina(n1147), .dinb(n4839), .dout(n8864));
  jor  g08609(.dina(n1246), .dinb(n5253), .dout(n8865));
  jor  g08610(.dina(n1251), .dinb(n5040), .dout(n8866));
  jand g08611(.dina(n8866), .dinb(n8865), .dout(n8867));
  jand g08612(.dina(n8867), .dinb(n8864), .dout(n8868));
  jand g08613(.dina(n8868), .dinb(n8863), .dout(n8869));
  jxor g08614(.dina(n8869), .dinb(n1061), .dout(n8870));
  jxor g08615(.dina(n8870), .dinb(n8862), .dout(n8871));
  jxor g08616(.dina(n8871), .dinb(n8674), .dout(n8872));
  jor  g08617(.dina(n5909), .dinb(n970), .dout(n8873));
  jor  g08618(.dina(n880), .dinb(n5469), .dout(n8874));
  jor  g08619(.dina(n972), .dinb(n5911), .dout(n8875));
  jor  g08620(.dina(n967), .dinb(n5685), .dout(n8876));
  jand g08621(.dina(n8876), .dinb(n8875), .dout(n8877));
  jand g08622(.dina(n8877), .dinb(n8874), .dout(n8878));
  jand g08623(.dina(n8878), .dinb(n8873), .dout(n8879));
  jxor g08624(.dina(n8879), .dinb(n810), .dout(n8880));
  jxor g08625(.dina(n8880), .dinb(n8872), .dout(n8881));
  jxor g08626(.dina(n8881), .dinb(n8671), .dout(n8882));
  jor  g08627(.dina(n6603), .dinb(n728), .dout(n8883));
  jor  g08628(.dina(n660), .dinb(n6139), .dout(n8884));
  jor  g08629(.dina(n731), .dinb(n6366), .dout(n8885));
  jor  g08630(.dina(n726), .dinb(n6605), .dout(n8886));
  jand g08631(.dina(n8886), .dinb(n8885), .dout(n8887));
  jand g08632(.dina(n8887), .dinb(n8884), .dout(n8888));
  jand g08633(.dina(n8888), .dinb(n8883), .dout(n8889));
  jxor g08634(.dina(n8889), .dinb(n606), .dout(n8890));
  jxor g08635(.dina(n8890), .dinb(n8882), .dout(n8891));
  jxor g08636(.dina(n8891), .dinb(n8668), .dout(n8892));
  jor  g08637(.dina(n7336), .dinb(n544), .dout(n8893));
  jor  g08638(.dina(n486), .dinb(n6846), .dout(n8894));
  jor  g08639(.dina(n547), .dinb(n7086), .dout(n8895));
  jor  g08640(.dina(n542), .dinb(n7338), .dout(n8896));
  jand g08641(.dina(n8896), .dinb(n8895), .dout(n8897));
  jand g08642(.dina(n8897), .dinb(n8894), .dout(n8898));
  jand g08643(.dina(n8898), .dinb(n8893), .dout(n8899));
  jxor g08644(.dina(n8899), .dinb(n446), .dout(n8900));
  jxor g08645(.dina(n8900), .dinb(n8892), .dout(n8901));
  jxor g08646(.dina(n8901), .dinb(n8665), .dout(n8902));
  jor  g08647(.dina(n8109), .dinb(n397), .dout(n8903));
  jor  g08648(.dina(n354), .dinb(n7590), .dout(n8904));
  jor  g08649(.dina(n394), .dinb(n7846), .dout(n8905));
  jor  g08650(.dina(n399), .dinb(n8111), .dout(n8906));
  jand g08651(.dina(n8906), .dinb(n8905), .dout(n8907));
  jand g08652(.dina(n8907), .dinb(n8904), .dout(n8908));
  jand g08653(.dina(n8908), .dinb(n8903), .dout(n8909));
  jxor g08654(.dina(n8909), .dinb(n364), .dout(n8910));
  jxor g08655(.dina(n8910), .dinb(n8902), .dout(n8911));
  jxor g08656(.dina(n8911), .dinb(n8662), .dout(n8912));
  jand g08657(.dina(b57 ), .dinb(b56 ), .dout(n8913));
  jand g08658(.dina(n8640), .dinb(n8639), .dout(n8914));
  jor  g08659(.dina(n8914), .dinb(n8913), .dout(n8915));
  jxor g08660(.dina(b58 ), .dinb(b57 ), .dout(n8916));
  jnot g08661(.din(n8916), .dout(n8917));
  jxor g08662(.dina(n8917), .dinb(n8915), .dout(n8918));
  jor  g08663(.dina(n8918), .dinb(n296), .dout(n8919));
  jnot g08664(.din(b58 ), .dout(n8920));
  jor  g08665(.dina(n264), .dinb(n8920), .dout(n8921));
  jor  g08666(.dina(n294), .dinb(n8644), .dout(n8922));
  jor  g08667(.dina(n280), .dinb(n8378), .dout(n8923));
  jand g08668(.dina(n8923), .dinb(n8922), .dout(n8924));
  jand g08669(.dina(n8924), .dinb(n8921), .dout(n8925));
  jand g08670(.dina(n8925), .dinb(n8919), .dout(n8926));
  jxor g08671(.dina(n8926), .dinb(n278), .dout(n8927));
  jxor g08672(.dina(n8927), .dinb(n8912), .dout(n8928));
  jxor g08673(.dina(n8928), .dinb(n8657), .dout(f58 ));
  jnot g08674(.din(n8927), .dout(n8930));
  jor  g08675(.dina(n8930), .dinb(n8912), .dout(n8931));
  jor  g08676(.dina(n8928), .dinb(n8657), .dout(n8932));
  jand g08677(.dina(n8932), .dinb(n8931), .dout(n8933));
  jand g08678(.dina(n8910), .dinb(n8902), .dout(n8934));
  jnot g08679(.din(n8934), .dout(n8935));
  jnot g08680(.din(n8911), .dout(n8936));
  jor  g08681(.dina(n8936), .dinb(n8662), .dout(n8937));
  jand g08682(.dina(n8937), .dinb(n8935), .dout(n8938));
  jand g08683(.dina(n8900), .dinb(n8892), .dout(n8939));
  jand g08684(.dina(n8901), .dinb(n8665), .dout(n8940));
  jor  g08685(.dina(n8940), .dinb(n8939), .dout(n8941));
  jand g08686(.dina(n8890), .dinb(n8882), .dout(n8942));
  jand g08687(.dina(n8891), .dinb(n8668), .dout(n8943));
  jor  g08688(.dina(n8943), .dinb(n8942), .dout(n8944));
  jand g08689(.dina(n8880), .dinb(n8872), .dout(n8945));
  jand g08690(.dina(n8881), .dinb(n8671), .dout(n8946));
  jor  g08691(.dina(n8946), .dinb(n8945), .dout(n8947));
  jand g08692(.dina(n8870), .dinb(n8862), .dout(n8948));
  jand g08693(.dina(n8871), .dinb(n8674), .dout(n8949));
  jor  g08694(.dina(n8949), .dinb(n8948), .dout(n8950));
  jand g08695(.dina(n8860), .dinb(n8852), .dout(n8951));
  jand g08696(.dina(n8861), .dinb(n8677), .dout(n8952));
  jor  g08697(.dina(n8952), .dinb(n8951), .dout(n8953));
  jand g08698(.dina(n8850), .dinb(n8842), .dout(n8954));
  jand g08699(.dina(n8851), .dinb(n8680), .dout(n8955));
  jor  g08700(.dina(n8955), .dinb(n8954), .dout(n8956));
  jand g08701(.dina(n8840), .dinb(n8832), .dout(n8957));
  jand g08702(.dina(n8841), .dinb(n8683), .dout(n8958));
  jor  g08703(.dina(n8958), .dinb(n8957), .dout(n8959));
  jand g08704(.dina(n8830), .dinb(n8822), .dout(n8960));
  jand g08705(.dina(n8831), .dinb(n8686), .dout(n8961));
  jor  g08706(.dina(n8961), .dinb(n8960), .dout(n8962));
  jand g08707(.dina(n8820), .dinb(n8812), .dout(n8963));
  jand g08708(.dina(n8821), .dinb(n8689), .dout(n8964));
  jor  g08709(.dina(n8964), .dinb(n8963), .dout(n8965));
  jand g08710(.dina(n8810), .dinb(n8802), .dout(n8966));
  jand g08711(.dina(n8811), .dinb(n8692), .dout(n8967));
  jor  g08712(.dina(n8967), .dinb(n8966), .dout(n8968));
  jand g08713(.dina(n8800), .dinb(n8792), .dout(n8969));
  jand g08714(.dina(n8801), .dinb(n8695), .dout(n8970));
  jor  g08715(.dina(n8970), .dinb(n8969), .dout(n8971));
  jand g08716(.dina(n8790), .dinb(n8782), .dout(n8972));
  jand g08717(.dina(n8791), .dinb(n8698), .dout(n8973));
  jor  g08718(.dina(n8973), .dinb(n8972), .dout(n8974));
  jand g08719(.dina(n8780), .dinb(n8772), .dout(n8975));
  jand g08720(.dina(n8781), .dinb(n8701), .dout(n8976));
  jor  g08721(.dina(n8976), .dinb(n8975), .dout(n8977));
  jand g08722(.dina(n8770), .dinb(n8762), .dout(n8978));
  jand g08723(.dina(n8771), .dinb(n8704), .dout(n8979));
  jor  g08724(.dina(n8979), .dinb(n8978), .dout(n8980));
  jand g08725(.dina(n8760), .dinb(n8752), .dout(n8981));
  jand g08726(.dina(n8761), .dinb(n8707), .dout(n8982));
  jor  g08727(.dina(n8982), .dinb(n8981), .dout(n8983));
  jor  g08728(.dina(n8750), .dinb(n8742), .dout(n8984));
  jand g08729(.dina(n8751), .dinb(n8712), .dout(n8985));
  jnot g08730(.din(n8985), .dout(n8986));
  jand g08731(.dina(n8986), .dinb(n8984), .dout(n8987));
  jnot g08732(.din(n8987), .dout(n8988));
  jor  g08733(.dina(n7660), .dinb(n517), .dout(n8989));
  jor  g08734(.dina(n7657), .dinb(n469), .dout(n8990));
  jor  g08735(.dina(n7662), .dinb(n519), .dout(n8991));
  jor  g08736(.dina(n7415), .dinb(n415), .dout(n8992));
  jand g08737(.dina(n8992), .dinb(n8991), .dout(n8993));
  jand g08738(.dina(n8993), .dinb(n8990), .dout(n8994));
  jand g08739(.dina(n8994), .dinb(n8989), .dout(n8995));
  jxor g08740(.dina(n8995), .dinb(n7166), .dout(n8996));
  jor  g08741(.dina(n8739), .dinb(n8731), .dout(n8997));
  jand g08742(.dina(n8740), .dinb(n8716), .dout(n8998));
  jnot g08743(.din(n8998), .dout(n8999));
  jand g08744(.dina(n8999), .dinb(n8997), .dout(n9000));
  jand g08745(.dina(n8722), .dinb(b1 ), .dout(n9001));
  jor  g08746(.dina(n8721), .dinb(n8450), .dout(n9002));
  jor  g08747(.dina(n9002), .dinb(n8724), .dout(n9003));
  jnot g08748(.din(n9003), .dout(n9004));
  jand g08749(.dina(n9004), .dinb(b0 ), .dout(n9005));
  jand g08750(.dina(n8718), .dinb(n273), .dout(n9006));
  jand g08751(.dina(n8725), .dinb(b2 ), .dout(n9007));
  jor  g08752(.dina(n9007), .dinb(n9006), .dout(n9008));
  jor  g08753(.dina(n9008), .dinb(n9005), .dout(n9009));
  jor  g08754(.dina(n9009), .dinb(n9001), .dout(n9010));
  jnot g08755(.din(n8728), .dout(n9011));
  jand g08756(.dina(n8452), .dinb(a59 ), .dout(n9012));
  jand g08757(.dina(n9012), .dinb(n9011), .dout(n9013));
  jnot g08758(.din(n9013), .dout(n9014));
  jand g08759(.dina(n9014), .dinb(a59 ), .dout(n9015));
  jxor g08760(.dina(n9015), .dinb(n9010), .dout(n9016));
  jor  g08761(.dina(n8457), .dinb(n374), .dout(n9017));
  jor  g08762(.dina(n8454), .dinb(n377), .dout(n9018));
  jor  g08763(.dina(n8185), .dinb(n303), .dout(n9019));
  jand g08764(.dina(n9019), .dinb(n9018), .dout(n9020));
  jor  g08765(.dina(n8459), .dinb(n340), .dout(n9021));
  jand g08766(.dina(n9021), .dinb(n9020), .dout(n9022));
  jand g08767(.dina(n9022), .dinb(n9017), .dout(n9023));
  jxor g08768(.dina(n9023), .dinb(a56 ), .dout(n9024));
  jxor g08769(.dina(n9024), .dinb(n9016), .dout(n9025));
  jxor g08770(.dina(n9025), .dinb(n9000), .dout(n9026));
  jxor g08771(.dina(n9026), .dinb(n8996), .dout(n9027));
  jxor g08772(.dina(n9027), .dinb(n8988), .dout(n9028));
  jor  g08773(.dina(n6914), .dinb(n702), .dout(n9029));
  jor  g08774(.dina(n6673), .dinb(n572), .dout(n9030));
  jor  g08775(.dina(n6916), .dinb(n704), .dout(n9031));
  jor  g08776(.dina(n6911), .dinb(n637), .dout(n9032));
  jand g08777(.dina(n9032), .dinb(n9031), .dout(n9033));
  jand g08778(.dina(n9033), .dinb(n9030), .dout(n9034));
  jand g08779(.dina(n9034), .dinb(n9029), .dout(n9035));
  jxor g08780(.dina(n9035), .dinb(n6443), .dout(n9036));
  jxor g08781(.dina(n9036), .dinb(n9028), .dout(n9037));
  jxor g08782(.dina(n9037), .dinb(n8983), .dout(n9038));
  jor  g08783(.dina(n6207), .dinb(n932), .dout(n9039));
  jor  g08784(.dina(n5975), .dinb(n772), .dout(n9040));
  jor  g08785(.dina(n6210), .dinb(n852), .dout(n9041));
  jor  g08786(.dina(n6205), .dinb(n934), .dout(n9042));
  jand g08787(.dina(n9042), .dinb(n9041), .dout(n9043));
  jand g08788(.dina(n9043), .dinb(n9040), .dout(n9044));
  jand g08789(.dina(n9044), .dinb(n9039), .dout(n9045));
  jxor g08790(.dina(n9045), .dinb(n5759), .dout(n9046));
  jxor g08791(.dina(n9046), .dinb(n9038), .dout(n9047));
  jxor g08792(.dina(n9047), .dinb(n8980), .dout(n9048));
  jor  g08793(.dina(n5537), .dinb(n1209), .dout(n9049));
  jor  g08794(.dina(n5315), .dinb(n1018), .dout(n9050));
  jor  g08795(.dina(n5539), .dinb(n1211), .dout(n9051));
  jor  g08796(.dina(n5534), .dinb(n1114), .dout(n9052));
  jand g08797(.dina(n9052), .dinb(n9051), .dout(n9053));
  jand g08798(.dina(n9053), .dinb(n9050), .dout(n9054));
  jand g08799(.dina(n9054), .dinb(n9049), .dout(n9055));
  jxor g08800(.dina(n9055), .dinb(n5111), .dout(n9056));
  jxor g08801(.dina(n9056), .dinb(n9048), .dout(n9057));
  jxor g08802(.dina(n9057), .dinb(n8977), .dout(n9058));
  jor  g08803(.dina(n4902), .dinb(n1525), .dout(n9059));
  jor  g08804(.dina(n4696), .dinb(n1307), .dout(n9060));
  jor  g08805(.dina(n4899), .dinb(n1527), .dout(n9061));
  jor  g08806(.dina(n4904), .dinb(n1416), .dout(n9062));
  jand g08807(.dina(n9062), .dinb(n9061), .dout(n9063));
  jand g08808(.dina(n9063), .dinb(n9060), .dout(n9064));
  jand g08809(.dina(n9064), .dinb(n9059), .dout(n9065));
  jxor g08810(.dina(n9065), .dinb(n4505), .dout(n9066));
  jxor g08811(.dina(n9066), .dinb(n9058), .dout(n9067));
  jxor g08812(.dina(n9067), .dinb(n8974), .dout(n9068));
  jor  g08813(.dina(n4305), .dinb(n1879), .dout(n9069));
  jor  g08814(.dina(n4116), .dinb(n1637), .dout(n9070));
  jor  g08815(.dina(n4308), .dinb(n1759), .dout(n9071));
  jor  g08816(.dina(n4303), .dinb(n1881), .dout(n9072));
  jand g08817(.dina(n9072), .dinb(n9071), .dout(n9073));
  jand g08818(.dina(n9073), .dinb(n9070), .dout(n9074));
  jand g08819(.dina(n9074), .dinb(n9069), .dout(n9075));
  jxor g08820(.dina(n9075), .dinb(n3938), .dout(n9076));
  jxor g08821(.dina(n9076), .dinb(n9068), .dout(n9077));
  jxor g08822(.dina(n9077), .dinb(n8971), .dout(n9078));
  jor  g08823(.dina(n3751), .dinb(n2277), .dout(n9079));
  jor  g08824(.dina(n3574), .dinb(n2007), .dout(n9080));
  jor  g08825(.dina(n3754), .dinb(n2142), .dout(n9081));
  jor  g08826(.dina(n3749), .dinb(n2279), .dout(n9082));
  jand g08827(.dina(n9082), .dinb(n9081), .dout(n9083));
  jand g08828(.dina(n9083), .dinb(n9080), .dout(n9084));
  jand g08829(.dina(n9084), .dinb(n9079), .dout(n9085));
  jxor g08830(.dina(n9085), .dinb(n3410), .dout(n9086));
  jxor g08831(.dina(n9086), .dinb(n9078), .dout(n9087));
  jxor g08832(.dina(n9087), .dinb(n8968), .dout(n9088));
  jor  g08833(.dina(n3239), .dinb(n2711), .dout(n9089));
  jor  g08834(.dina(n3072), .dinb(n2415), .dout(n9090));
  jor  g08835(.dina(n3242), .dinb(n2563), .dout(n9091));
  jor  g08836(.dina(n3237), .dinb(n2713), .dout(n9092));
  jand g08837(.dina(n9092), .dinb(n9091), .dout(n9093));
  jand g08838(.dina(n9093), .dinb(n9090), .dout(n9094));
  jand g08839(.dina(n9094), .dinb(n9089), .dout(n9095));
  jxor g08840(.dina(n9095), .dinb(n2918), .dout(n9096));
  jxor g08841(.dina(n9096), .dinb(n9088), .dout(n9097));
  jxor g08842(.dina(n9097), .dinb(n8965), .dout(n9098));
  jor  g08843(.dina(n3184), .dinb(n2764), .dout(n9099));
  jor  g08844(.dina(n2609), .dinb(n2862), .dout(n9100));
  jor  g08845(.dina(n2761), .dinb(n3186), .dout(n9101));
  jor  g08846(.dina(n2766), .dinb(n3023), .dout(n9102));
  jand g08847(.dina(n9102), .dinb(n9101), .dout(n9103));
  jand g08848(.dina(n9103), .dinb(n9100), .dout(n9104));
  jand g08849(.dina(n9104), .dinb(n9099), .dout(n9105));
  jxor g08850(.dina(n9105), .dinb(n2468), .dout(n9106));
  jxor g08851(.dina(n9106), .dinb(n9098), .dout(n9107));
  jxor g08852(.dina(n9107), .dinb(n8962), .dout(n9108));
  jor  g08853(.dina(n3696), .dinb(n2324), .dout(n9109));
  jor  g08854(.dina(n2186), .dinb(n3348), .dout(n9110));
  jor  g08855(.dina(n2321), .dinb(n3522), .dout(n9111));
  jor  g08856(.dina(n2326), .dinb(n3698), .dout(n9112));
  jand g08857(.dina(n9112), .dinb(n9111), .dout(n9113));
  jand g08858(.dina(n9113), .dinb(n9110), .dout(n9114));
  jand g08859(.dina(n9114), .dinb(n9109), .dout(n9115));
  jxor g08860(.dina(n9115), .dinb(n2057), .dout(n9116));
  jxor g08861(.dina(n9116), .dinb(n9108), .dout(n9117));
  jxor g08862(.dina(n9117), .dinb(n8959), .dout(n9118));
  jor  g08863(.dina(n4247), .dinb(n1921), .dout(n9119));
  jor  g08864(.dina(n1806), .dinb(n3873), .dout(n9120));
  jor  g08865(.dina(n1918), .dinb(n4060), .dout(n9121));
  jor  g08866(.dina(n1923), .dinb(n4249), .dout(n9122));
  jand g08867(.dina(n9122), .dinb(n9121), .dout(n9123));
  jand g08868(.dina(n9123), .dinb(n9120), .dout(n9124));
  jand g08869(.dina(n9124), .dinb(n9119), .dout(n9125));
  jxor g08870(.dina(n9125), .dinb(n1687), .dout(n9126));
  jxor g08871(.dina(n9126), .dinb(n9118), .dout(n9127));
  jxor g08872(.dina(n9127), .dinb(n8956), .dout(n9128));
  jor  g08873(.dina(n4837), .dinb(n1569), .dout(n9129));
  jor  g08874(.dina(n1453), .dinb(n4437), .dout(n9130));
  jor  g08875(.dina(n1566), .dinb(n4637), .dout(n9131));
  jor  g08876(.dina(n1571), .dinb(n4839), .dout(n9132));
  jand g08877(.dina(n9132), .dinb(n9131), .dout(n9133));
  jand g08878(.dina(n9133), .dinb(n9130), .dout(n9134));
  jand g08879(.dina(n9134), .dinb(n9129), .dout(n9135));
  jxor g08880(.dina(n9135), .dinb(n1351), .dout(n9136));
  jxor g08881(.dina(n9136), .dinb(n9128), .dout(n9137));
  jxor g08882(.dina(n9137), .dinb(n8953), .dout(n9138));
  jor  g08883(.dina(n5467), .dinb(n1248), .dout(n9139));
  jor  g08884(.dina(n1147), .dinb(n5040), .dout(n9140));
  jor  g08885(.dina(n1251), .dinb(n5253), .dout(n9141));
  jor  g08886(.dina(n1246), .dinb(n5469), .dout(n9142));
  jand g08887(.dina(n9142), .dinb(n9141), .dout(n9143));
  jand g08888(.dina(n9143), .dinb(n9140), .dout(n9144));
  jand g08889(.dina(n9144), .dinb(n9139), .dout(n9145));
  jxor g08890(.dina(n9145), .dinb(n1061), .dout(n9146));
  jxor g08891(.dina(n9146), .dinb(n9138), .dout(n9147));
  jxor g08892(.dina(n9147), .dinb(n8950), .dout(n9148));
  jor  g08893(.dina(n6137), .dinb(n970), .dout(n9149));
  jor  g08894(.dina(n880), .dinb(n5685), .dout(n9150));
  jor  g08895(.dina(n972), .dinb(n6139), .dout(n9151));
  jor  g08896(.dina(n967), .dinb(n5911), .dout(n9152));
  jand g08897(.dina(n9152), .dinb(n9151), .dout(n9153));
  jand g08898(.dina(n9153), .dinb(n9150), .dout(n9154));
  jand g08899(.dina(n9154), .dinb(n9149), .dout(n9155));
  jxor g08900(.dina(n9155), .dinb(n810), .dout(n9156));
  jxor g08901(.dina(n9156), .dinb(n9148), .dout(n9157));
  jxor g08902(.dina(n9157), .dinb(n8947), .dout(n9158));
  jor  g08903(.dina(n6844), .dinb(n728), .dout(n9159));
  jor  g08904(.dina(n660), .dinb(n6366), .dout(n9160));
  jor  g08905(.dina(n726), .dinb(n6846), .dout(n9161));
  jor  g08906(.dina(n731), .dinb(n6605), .dout(n9162));
  jand g08907(.dina(n9162), .dinb(n9161), .dout(n9163));
  jand g08908(.dina(n9163), .dinb(n9160), .dout(n9164));
  jand g08909(.dina(n9164), .dinb(n9159), .dout(n9165));
  jxor g08910(.dina(n9165), .dinb(n606), .dout(n9166));
  jxor g08911(.dina(n9166), .dinb(n9158), .dout(n9167));
  jxor g08912(.dina(n9167), .dinb(n8944), .dout(n9168));
  jor  g08913(.dina(n7588), .dinb(n544), .dout(n9169));
  jor  g08914(.dina(n486), .dinb(n7086), .dout(n9170));
  jor  g08915(.dina(n547), .dinb(n7338), .dout(n9171));
  jor  g08916(.dina(n542), .dinb(n7590), .dout(n9172));
  jand g08917(.dina(n9172), .dinb(n9171), .dout(n9173));
  jand g08918(.dina(n9173), .dinb(n9170), .dout(n9174));
  jand g08919(.dina(n9174), .dinb(n9169), .dout(n9175));
  jxor g08920(.dina(n9175), .dinb(n446), .dout(n9176));
  jxor g08921(.dina(n9176), .dinb(n9168), .dout(n9177));
  jxor g08922(.dina(n9177), .dinb(n8941), .dout(n9178));
  jor  g08923(.dina(n8376), .dinb(n397), .dout(n9179));
  jor  g08924(.dina(n354), .dinb(n7846), .dout(n9180));
  jor  g08925(.dina(n394), .dinb(n8111), .dout(n9181));
  jor  g08926(.dina(n399), .dinb(n8378), .dout(n9182));
  jand g08927(.dina(n9182), .dinb(n9181), .dout(n9183));
  jand g08928(.dina(n9183), .dinb(n9180), .dout(n9184));
  jand g08929(.dina(n9184), .dinb(n9179), .dout(n9185));
  jxor g08930(.dina(n9185), .dinb(n364), .dout(n9186));
  jxor g08931(.dina(n9186), .dinb(n9178), .dout(n9187));
  jand g08932(.dina(b58 ), .dinb(b57 ), .dout(n9188));
  jand g08933(.dina(n8916), .dinb(n8915), .dout(n9189));
  jor  g08934(.dina(n9189), .dinb(n9188), .dout(n9190));
  jxor g08935(.dina(b59 ), .dinb(b58 ), .dout(n9191));
  jnot g08936(.din(n9191), .dout(n9192));
  jxor g08937(.dina(n9192), .dinb(n9190), .dout(n9193));
  jor  g08938(.dina(n9193), .dinb(n296), .dout(n9194));
  jnot g08939(.din(b59 ), .dout(n9195));
  jor  g08940(.dina(n264), .dinb(n9195), .dout(n9196));
  jor  g08941(.dina(n294), .dinb(n8920), .dout(n9197));
  jor  g08942(.dina(n280), .dinb(n8644), .dout(n9198));
  jand g08943(.dina(n9198), .dinb(n9197), .dout(n9199));
  jand g08944(.dina(n9199), .dinb(n9196), .dout(n9200));
  jand g08945(.dina(n9200), .dinb(n9194), .dout(n9201));
  jxor g08946(.dina(n9201), .dinb(n278), .dout(n9202));
  jxor g08947(.dina(n9202), .dinb(n9187), .dout(n9203));
  jxor g08948(.dina(n9203), .dinb(n8938), .dout(n9204));
  jxor g08949(.dina(n9204), .dinb(n8933), .dout(f59 ));
  jnot g08950(.din(n8938), .dout(n9206));
  jand g08951(.dina(n9203), .dinb(n9206), .dout(n9207));
  jnot g08952(.din(n9207), .dout(n9208));
  jor  g08953(.dina(n9204), .dinb(n8933), .dout(n9209));
  jand g08954(.dina(n9209), .dinb(n9208), .dout(n9210));
  jand g08955(.dina(n9186), .dinb(n9178), .dout(n9211));
  jand g08956(.dina(n9202), .dinb(n9187), .dout(n9212));
  jor  g08957(.dina(n9212), .dinb(n9211), .dout(n9213));
  jnot g08958(.din(n9213), .dout(n9214));
  jand g08959(.dina(n9176), .dinb(n9168), .dout(n9215));
  jand g08960(.dina(n9177), .dinb(n8941), .dout(n9216));
  jor  g08961(.dina(n9216), .dinb(n9215), .dout(n9217));
  jand g08962(.dina(n9166), .dinb(n9158), .dout(n9218));
  jand g08963(.dina(n9167), .dinb(n8944), .dout(n9219));
  jor  g08964(.dina(n9219), .dinb(n9218), .dout(n9220));
  jand g08965(.dina(n9156), .dinb(n9148), .dout(n9221));
  jand g08966(.dina(n9157), .dinb(n8947), .dout(n9222));
  jor  g08967(.dina(n9222), .dinb(n9221), .dout(n9223));
  jand g08968(.dina(n9146), .dinb(n9138), .dout(n9224));
  jand g08969(.dina(n9147), .dinb(n8950), .dout(n9225));
  jor  g08970(.dina(n9225), .dinb(n9224), .dout(n9226));
  jand g08971(.dina(n9136), .dinb(n9128), .dout(n9227));
  jand g08972(.dina(n9137), .dinb(n8953), .dout(n9228));
  jor  g08973(.dina(n9228), .dinb(n9227), .dout(n9229));
  jand g08974(.dina(n9126), .dinb(n9118), .dout(n9230));
  jand g08975(.dina(n9127), .dinb(n8956), .dout(n9231));
  jor  g08976(.dina(n9231), .dinb(n9230), .dout(n9232));
  jand g08977(.dina(n9116), .dinb(n9108), .dout(n9233));
  jand g08978(.dina(n9117), .dinb(n8959), .dout(n9234));
  jor  g08979(.dina(n9234), .dinb(n9233), .dout(n9235));
  jand g08980(.dina(n9106), .dinb(n9098), .dout(n9236));
  jand g08981(.dina(n9107), .dinb(n8962), .dout(n9237));
  jor  g08982(.dina(n9237), .dinb(n9236), .dout(n9238));
  jand g08983(.dina(n9096), .dinb(n9088), .dout(n9239));
  jand g08984(.dina(n9097), .dinb(n8965), .dout(n9240));
  jor  g08985(.dina(n9240), .dinb(n9239), .dout(n9241));
  jand g08986(.dina(n9086), .dinb(n9078), .dout(n9242));
  jand g08987(.dina(n9087), .dinb(n8968), .dout(n9243));
  jor  g08988(.dina(n9243), .dinb(n9242), .dout(n9244));
  jand g08989(.dina(n9076), .dinb(n9068), .dout(n9245));
  jand g08990(.dina(n9077), .dinb(n8971), .dout(n9246));
  jor  g08991(.dina(n9246), .dinb(n9245), .dout(n9247));
  jand g08992(.dina(n9066), .dinb(n9058), .dout(n9248));
  jand g08993(.dina(n9067), .dinb(n8974), .dout(n9249));
  jor  g08994(.dina(n9249), .dinb(n9248), .dout(n9250));
  jand g08995(.dina(n9056), .dinb(n9048), .dout(n9251));
  jand g08996(.dina(n9057), .dinb(n8977), .dout(n9252));
  jor  g08997(.dina(n9252), .dinb(n9251), .dout(n9253));
  jand g08998(.dina(n9046), .dinb(n9038), .dout(n9254));
  jand g08999(.dina(n9047), .dinb(n8980), .dout(n9255));
  jor  g09000(.dina(n9255), .dinb(n9254), .dout(n9256));
  jand g09001(.dina(n9036), .dinb(n9028), .dout(n9257));
  jand g09002(.dina(n9037), .dinb(n8983), .dout(n9258));
  jor  g09003(.dina(n9258), .dinb(n9257), .dout(n9259));
  jand g09004(.dina(n9026), .dinb(n8996), .dout(n9260));
  jand g09005(.dina(n9027), .dinb(n8988), .dout(n9261));
  jor  g09006(.dina(n9261), .dinb(n9260), .dout(n9262));
  jor  g09007(.dina(n9014), .dinb(n9010), .dout(n9263));
  jxor g09008(.dina(a60 ), .dinb(a59 ), .dout(n9264));
  jand g09009(.dina(n9264), .dinb(b0 ), .dout(n9265));
  jnot g09010(.din(n9265), .dout(n9266));
  jxor g09011(.dina(n9266), .dinb(n9263), .dout(n9267));
  jnot g09012(.din(n8725), .dout(n9268));
  jor  g09013(.dina(n9268), .dinb(n303), .dout(n9269));
  jor  g09014(.dina(n9003), .dinb(n305), .dout(n9270));
  jnot g09015(.din(n8718), .dout(n9271));
  jor  g09016(.dina(n9271), .dinb(n301), .dout(n9272));
  jnot g09017(.din(n8722), .dout(n9273));
  jor  g09018(.dina(n9273), .dinb(n293), .dout(n9274));
  jand g09019(.dina(n9274), .dinb(n9272), .dout(n9275));
  jand g09020(.dina(n9275), .dinb(n9270), .dout(n9276));
  jand g09021(.dina(n9276), .dinb(n9269), .dout(n9277));
  jxor g09022(.dina(n9277), .dinb(n8729), .dout(n9278));
  jxor g09023(.dina(n9278), .dinb(n9267), .dout(n9279));
  jnot g09024(.din(n9279), .dout(n9280));
  jor  g09025(.dina(n8457), .dinb(n412), .dout(n9281));
  jor  g09026(.dina(n8454), .dinb(n415), .dout(n9282));
  jor  g09027(.dina(n8185), .dinb(n340), .dout(n9283));
  jand g09028(.dina(n9283), .dinb(n9282), .dout(n9284));
  jor  g09029(.dina(n8459), .dinb(n377), .dout(n9285));
  jand g09030(.dina(n9285), .dinb(n9284), .dout(n9286));
  jand g09031(.dina(n9286), .dinb(n9281), .dout(n9287));
  jxor g09032(.dina(n9287), .dinb(a56 ), .dout(n9288));
  jxor g09033(.dina(n9288), .dinb(n9280), .dout(n9289));
  jnot g09034(.din(n9016), .dout(n9290));
  jand g09035(.dina(n9024), .dinb(n9290), .dout(n9291));
  jnot g09036(.din(n9291), .dout(n9292));
  jnot g09037(.din(n9000), .dout(n9293));
  jnot g09038(.din(n9024), .dout(n9294));
  jand g09039(.dina(n9294), .dinb(n9016), .dout(n9295));
  jor  g09040(.dina(n9295), .dinb(n9293), .dout(n9296));
  jand g09041(.dina(n9296), .dinb(n9292), .dout(n9297));
  jxor g09042(.dina(n9297), .dinb(n9289), .dout(n9298));
  jor  g09043(.dina(n7660), .dinb(n570), .dout(n9299));
  jor  g09044(.dina(n7415), .dinb(n469), .dout(n9300));
  jor  g09045(.dina(n7657), .dinb(n519), .dout(n9301));
  jor  g09046(.dina(n7662), .dinb(n572), .dout(n9302));
  jand g09047(.dina(n9302), .dinb(n9301), .dout(n9303));
  jand g09048(.dina(n9303), .dinb(n9300), .dout(n9304));
  jand g09049(.dina(n9304), .dinb(n9299), .dout(n9305));
  jxor g09050(.dina(n9305), .dinb(n7166), .dout(n9306));
  jxor g09051(.dina(n9306), .dinb(n9298), .dout(n9307));
  jxor g09052(.dina(n9307), .dinb(n9262), .dout(n9308));
  jor  g09053(.dina(n6914), .dinb(n770), .dout(n9309));
  jor  g09054(.dina(n6673), .dinb(n637), .dout(n9310));
  jor  g09055(.dina(n6916), .dinb(n772), .dout(n9311));
  jor  g09056(.dina(n6911), .dinb(n704), .dout(n9312));
  jand g09057(.dina(n9312), .dinb(n9311), .dout(n9313));
  jand g09058(.dina(n9313), .dinb(n9310), .dout(n9314));
  jand g09059(.dina(n9314), .dinb(n9309), .dout(n9315));
  jxor g09060(.dina(n9315), .dinb(n6443), .dout(n9316));
  jxor g09061(.dina(n9316), .dinb(n9308), .dout(n9317));
  jxor g09062(.dina(n9317), .dinb(n9259), .dout(n9318));
  jor  g09063(.dina(n6207), .dinb(n1016), .dout(n9319));
  jor  g09064(.dina(n5975), .dinb(n852), .dout(n9320));
  jor  g09065(.dina(n6205), .dinb(n1018), .dout(n9321));
  jor  g09066(.dina(n6210), .dinb(n934), .dout(n9322));
  jand g09067(.dina(n9322), .dinb(n9321), .dout(n9323));
  jand g09068(.dina(n9323), .dinb(n9320), .dout(n9324));
  jand g09069(.dina(n9324), .dinb(n9319), .dout(n9325));
  jxor g09070(.dina(n9325), .dinb(n5759), .dout(n9326));
  jxor g09071(.dina(n9326), .dinb(n9318), .dout(n9327));
  jxor g09072(.dina(n9327), .dinb(n9256), .dout(n9328));
  jor  g09073(.dina(n5537), .dinb(n1305), .dout(n9329));
  jor  g09074(.dina(n5315), .dinb(n1114), .dout(n9330));
  jor  g09075(.dina(n5534), .dinb(n1211), .dout(n9331));
  jor  g09076(.dina(n5539), .dinb(n1307), .dout(n9332));
  jand g09077(.dina(n9332), .dinb(n9331), .dout(n9333));
  jand g09078(.dina(n9333), .dinb(n9330), .dout(n9334));
  jand g09079(.dina(n9334), .dinb(n9329), .dout(n9335));
  jxor g09080(.dina(n9335), .dinb(n5111), .dout(n9336));
  jxor g09081(.dina(n9336), .dinb(n9328), .dout(n9337));
  jxor g09082(.dina(n9337), .dinb(n9253), .dout(n9338));
  jor  g09083(.dina(n4902), .dinb(n1635), .dout(n9339));
  jor  g09084(.dina(n4696), .dinb(n1416), .dout(n9340));
  jor  g09085(.dina(n4904), .dinb(n1527), .dout(n9341));
  jor  g09086(.dina(n4899), .dinb(n1637), .dout(n9342));
  jand g09087(.dina(n9342), .dinb(n9341), .dout(n9343));
  jand g09088(.dina(n9343), .dinb(n9340), .dout(n9344));
  jand g09089(.dina(n9344), .dinb(n9339), .dout(n9345));
  jxor g09090(.dina(n9345), .dinb(n4505), .dout(n9346));
  jxor g09091(.dina(n9346), .dinb(n9338), .dout(n9347));
  jxor g09092(.dina(n9347), .dinb(n9250), .dout(n9348));
  jor  g09093(.dina(n4305), .dinb(n2005), .dout(n9349));
  jor  g09094(.dina(n4116), .dinb(n1759), .dout(n9350));
  jor  g09095(.dina(n4308), .dinb(n1881), .dout(n9351));
  jor  g09096(.dina(n4303), .dinb(n2007), .dout(n9352));
  jand g09097(.dina(n9352), .dinb(n9351), .dout(n9353));
  jand g09098(.dina(n9353), .dinb(n9350), .dout(n9354));
  jand g09099(.dina(n9354), .dinb(n9349), .dout(n9355));
  jxor g09100(.dina(n9355), .dinb(n3938), .dout(n9356));
  jxor g09101(.dina(n9356), .dinb(n9348), .dout(n9357));
  jxor g09102(.dina(n9357), .dinb(n9247), .dout(n9358));
  jor  g09103(.dina(n3751), .dinb(n2413), .dout(n9359));
  jor  g09104(.dina(n3574), .dinb(n2142), .dout(n9360));
  jor  g09105(.dina(n3754), .dinb(n2279), .dout(n9361));
  jor  g09106(.dina(n3749), .dinb(n2415), .dout(n9362));
  jand g09107(.dina(n9362), .dinb(n9361), .dout(n9363));
  jand g09108(.dina(n9363), .dinb(n9360), .dout(n9364));
  jand g09109(.dina(n9364), .dinb(n9359), .dout(n9365));
  jxor g09110(.dina(n9365), .dinb(n3410), .dout(n9366));
  jxor g09111(.dina(n9366), .dinb(n9358), .dout(n9367));
  jxor g09112(.dina(n9367), .dinb(n9244), .dout(n9368));
  jor  g09113(.dina(n3239), .dinb(n2860), .dout(n9369));
  jor  g09114(.dina(n3072), .dinb(n2563), .dout(n9370));
  jor  g09115(.dina(n3242), .dinb(n2713), .dout(n9371));
  jor  g09116(.dina(n3237), .dinb(n2862), .dout(n9372));
  jand g09117(.dina(n9372), .dinb(n9371), .dout(n9373));
  jand g09118(.dina(n9373), .dinb(n9370), .dout(n9374));
  jand g09119(.dina(n9374), .dinb(n9369), .dout(n9375));
  jxor g09120(.dina(n9375), .dinb(n2918), .dout(n9376));
  jxor g09121(.dina(n9376), .dinb(n9368), .dout(n9377));
  jxor g09122(.dina(n9377), .dinb(n9241), .dout(n9378));
  jor  g09123(.dina(n3346), .dinb(n2764), .dout(n9379));
  jor  g09124(.dina(n2609), .dinb(n3023), .dout(n9380));
  jor  g09125(.dina(n2761), .dinb(n3348), .dout(n9381));
  jor  g09126(.dina(n2766), .dinb(n3186), .dout(n9382));
  jand g09127(.dina(n9382), .dinb(n9381), .dout(n9383));
  jand g09128(.dina(n9383), .dinb(n9380), .dout(n9384));
  jand g09129(.dina(n9384), .dinb(n9379), .dout(n9385));
  jxor g09130(.dina(n9385), .dinb(n2468), .dout(n9386));
  jxor g09131(.dina(n9386), .dinb(n9378), .dout(n9387));
  jxor g09132(.dina(n9387), .dinb(n9238), .dout(n9388));
  jor  g09133(.dina(n3871), .dinb(n2324), .dout(n9389));
  jor  g09134(.dina(n2186), .dinb(n3522), .dout(n9390));
  jor  g09135(.dina(n2326), .dinb(n3873), .dout(n9391));
  jor  g09136(.dina(n2321), .dinb(n3698), .dout(n9392));
  jand g09137(.dina(n9392), .dinb(n9391), .dout(n9393));
  jand g09138(.dina(n9393), .dinb(n9390), .dout(n9394));
  jand g09139(.dina(n9394), .dinb(n9389), .dout(n9395));
  jxor g09140(.dina(n9395), .dinb(n2057), .dout(n9396));
  jxor g09141(.dina(n9396), .dinb(n9388), .dout(n9397));
  jxor g09142(.dina(n9397), .dinb(n9235), .dout(n9398));
  jor  g09143(.dina(n4435), .dinb(n1921), .dout(n9399));
  jor  g09144(.dina(n1806), .dinb(n4060), .dout(n9400));
  jor  g09145(.dina(n1918), .dinb(n4249), .dout(n9401));
  jor  g09146(.dina(n1923), .dinb(n4437), .dout(n9402));
  jand g09147(.dina(n9402), .dinb(n9401), .dout(n9403));
  jand g09148(.dina(n9403), .dinb(n9400), .dout(n9404));
  jand g09149(.dina(n9404), .dinb(n9399), .dout(n9405));
  jxor g09150(.dina(n9405), .dinb(n1687), .dout(n9406));
  jxor g09151(.dina(n9406), .dinb(n9398), .dout(n9407));
  jxor g09152(.dina(n9407), .dinb(n9232), .dout(n9408));
  jor  g09153(.dina(n5038), .dinb(n1569), .dout(n9409));
  jor  g09154(.dina(n1453), .dinb(n4637), .dout(n9410));
  jor  g09155(.dina(n1566), .dinb(n4839), .dout(n9411));
  jor  g09156(.dina(n1571), .dinb(n5040), .dout(n9412));
  jand g09157(.dina(n9412), .dinb(n9411), .dout(n9413));
  jand g09158(.dina(n9413), .dinb(n9410), .dout(n9414));
  jand g09159(.dina(n9414), .dinb(n9409), .dout(n9415));
  jxor g09160(.dina(n9415), .dinb(n1351), .dout(n9416));
  jxor g09161(.dina(n9416), .dinb(n9408), .dout(n9417));
  jxor g09162(.dina(n9417), .dinb(n9229), .dout(n9418));
  jor  g09163(.dina(n5683), .dinb(n1248), .dout(n9419));
  jor  g09164(.dina(n1147), .dinb(n5253), .dout(n9420));
  jor  g09165(.dina(n1251), .dinb(n5469), .dout(n9421));
  jor  g09166(.dina(n1246), .dinb(n5685), .dout(n9422));
  jand g09167(.dina(n9422), .dinb(n9421), .dout(n9423));
  jand g09168(.dina(n9423), .dinb(n9420), .dout(n9424));
  jand g09169(.dina(n9424), .dinb(n9419), .dout(n9425));
  jxor g09170(.dina(n9425), .dinb(n1061), .dout(n9426));
  jxor g09171(.dina(n9426), .dinb(n9418), .dout(n9427));
  jxor g09172(.dina(n9427), .dinb(n9226), .dout(n9428));
  jor  g09173(.dina(n6364), .dinb(n970), .dout(n9429));
  jor  g09174(.dina(n880), .dinb(n5911), .dout(n9430));
  jor  g09175(.dina(n972), .dinb(n6366), .dout(n9431));
  jor  g09176(.dina(n967), .dinb(n6139), .dout(n9432));
  jand g09177(.dina(n9432), .dinb(n9431), .dout(n9433));
  jand g09178(.dina(n9433), .dinb(n9430), .dout(n9434));
  jand g09179(.dina(n9434), .dinb(n9429), .dout(n9435));
  jxor g09180(.dina(n9435), .dinb(n810), .dout(n9436));
  jxor g09181(.dina(n9436), .dinb(n9428), .dout(n9437));
  jxor g09182(.dina(n9437), .dinb(n9223), .dout(n9438));
  jor  g09183(.dina(n7084), .dinb(n728), .dout(n9439));
  jor  g09184(.dina(n660), .dinb(n6605), .dout(n9440));
  jor  g09185(.dina(n731), .dinb(n6846), .dout(n9441));
  jor  g09186(.dina(n726), .dinb(n7086), .dout(n9442));
  jand g09187(.dina(n9442), .dinb(n9441), .dout(n9443));
  jand g09188(.dina(n9443), .dinb(n9440), .dout(n9444));
  jand g09189(.dina(n9444), .dinb(n9439), .dout(n9445));
  jxor g09190(.dina(n9445), .dinb(n606), .dout(n9446));
  jxor g09191(.dina(n9446), .dinb(n9438), .dout(n9447));
  jxor g09192(.dina(n9447), .dinb(n9220), .dout(n9448));
  jor  g09193(.dina(n7844), .dinb(n544), .dout(n9449));
  jor  g09194(.dina(n486), .dinb(n7338), .dout(n9450));
  jor  g09195(.dina(n547), .dinb(n7590), .dout(n9451));
  jor  g09196(.dina(n542), .dinb(n7846), .dout(n9452));
  jand g09197(.dina(n9452), .dinb(n9451), .dout(n9453));
  jand g09198(.dina(n9453), .dinb(n9450), .dout(n9454));
  jand g09199(.dina(n9454), .dinb(n9449), .dout(n9455));
  jxor g09200(.dina(n9455), .dinb(n446), .dout(n9456));
  jxor g09201(.dina(n9456), .dinb(n9448), .dout(n9457));
  jxor g09202(.dina(n9457), .dinb(n9217), .dout(n9458));
  jor  g09203(.dina(n8642), .dinb(n397), .dout(n9459));
  jor  g09204(.dina(n354), .dinb(n8111), .dout(n9460));
  jor  g09205(.dina(n399), .dinb(n8644), .dout(n9461));
  jor  g09206(.dina(n394), .dinb(n8378), .dout(n9462));
  jand g09207(.dina(n9462), .dinb(n9461), .dout(n9463));
  jand g09208(.dina(n9463), .dinb(n9460), .dout(n9464));
  jand g09209(.dina(n9464), .dinb(n9459), .dout(n9465));
  jxor g09210(.dina(n9465), .dinb(n364), .dout(n9466));
  jxor g09211(.dina(n9466), .dinb(n9458), .dout(n9467));
  jand g09212(.dina(b59 ), .dinb(b58 ), .dout(n9468));
  jand g09213(.dina(n9191), .dinb(n9190), .dout(n9469));
  jor  g09214(.dina(n9469), .dinb(n9468), .dout(n9470));
  jxor g09215(.dina(b60 ), .dinb(b59 ), .dout(n9471));
  jnot g09216(.din(n9471), .dout(n9472));
  jxor g09217(.dina(n9472), .dinb(n9470), .dout(n9473));
  jor  g09218(.dina(n9473), .dinb(n296), .dout(n9474));
  jnot g09219(.din(b60 ), .dout(n9475));
  jor  g09220(.dina(n264), .dinb(n9475), .dout(n9476));
  jor  g09221(.dina(n280), .dinb(n8920), .dout(n9477));
  jor  g09222(.dina(n294), .dinb(n9195), .dout(n9478));
  jand g09223(.dina(n9478), .dinb(n9477), .dout(n9479));
  jand g09224(.dina(n9479), .dinb(n9476), .dout(n9480));
  jand g09225(.dina(n9480), .dinb(n9474), .dout(n9481));
  jxor g09226(.dina(n9481), .dinb(n278), .dout(n9482));
  jxor g09227(.dina(n9482), .dinb(n9467), .dout(n9483));
  jxor g09228(.dina(n9483), .dinb(n9214), .dout(n9484));
  jxor g09229(.dina(n9484), .dinb(n9210), .dout(f60 ));
  jand g09230(.dina(n9466), .dinb(n9458), .dout(n9486));
  jand g09231(.dina(n9482), .dinb(n9467), .dout(n9487));
  jor  g09232(.dina(n9487), .dinb(n9486), .dout(n9488));
  jnot g09233(.din(n9488), .dout(n9489));
  jand g09234(.dina(n9456), .dinb(n9448), .dout(n9490));
  jand g09235(.dina(n9457), .dinb(n9217), .dout(n9491));
  jor  g09236(.dina(n9491), .dinb(n9490), .dout(n9492));
  jand g09237(.dina(n9446), .dinb(n9438), .dout(n9493));
  jand g09238(.dina(n9447), .dinb(n9220), .dout(n9494));
  jor  g09239(.dina(n9494), .dinb(n9493), .dout(n9495));
  jand g09240(.dina(n9436), .dinb(n9428), .dout(n9496));
  jand g09241(.dina(n9437), .dinb(n9223), .dout(n9497));
  jor  g09242(.dina(n9497), .dinb(n9496), .dout(n9498));
  jand g09243(.dina(n9426), .dinb(n9418), .dout(n9499));
  jand g09244(.dina(n9427), .dinb(n9226), .dout(n9500));
  jor  g09245(.dina(n9500), .dinb(n9499), .dout(n9501));
  jand g09246(.dina(n9416), .dinb(n9408), .dout(n9502));
  jand g09247(.dina(n9417), .dinb(n9229), .dout(n9503));
  jor  g09248(.dina(n9503), .dinb(n9502), .dout(n9504));
  jand g09249(.dina(n9406), .dinb(n9398), .dout(n9505));
  jand g09250(.dina(n9407), .dinb(n9232), .dout(n9506));
  jor  g09251(.dina(n9506), .dinb(n9505), .dout(n9507));
  jand g09252(.dina(n9396), .dinb(n9388), .dout(n9508));
  jand g09253(.dina(n9397), .dinb(n9235), .dout(n9509));
  jor  g09254(.dina(n9509), .dinb(n9508), .dout(n9510));
  jand g09255(.dina(n9386), .dinb(n9378), .dout(n9511));
  jand g09256(.dina(n9387), .dinb(n9238), .dout(n9512));
  jor  g09257(.dina(n9512), .dinb(n9511), .dout(n9513));
  jand g09258(.dina(n9376), .dinb(n9368), .dout(n9514));
  jand g09259(.dina(n9377), .dinb(n9241), .dout(n9515));
  jor  g09260(.dina(n9515), .dinb(n9514), .dout(n9516));
  jand g09261(.dina(n9366), .dinb(n9358), .dout(n9517));
  jand g09262(.dina(n9367), .dinb(n9244), .dout(n9518));
  jor  g09263(.dina(n9518), .dinb(n9517), .dout(n9519));
  jand g09264(.dina(n9356), .dinb(n9348), .dout(n9520));
  jand g09265(.dina(n9357), .dinb(n9247), .dout(n9521));
  jor  g09266(.dina(n9521), .dinb(n9520), .dout(n9522));
  jand g09267(.dina(n9346), .dinb(n9338), .dout(n9523));
  jand g09268(.dina(n9347), .dinb(n9250), .dout(n9524));
  jor  g09269(.dina(n9524), .dinb(n9523), .dout(n9525));
  jand g09270(.dina(n9336), .dinb(n9328), .dout(n9526));
  jand g09271(.dina(n9337), .dinb(n9253), .dout(n9527));
  jor  g09272(.dina(n9527), .dinb(n9526), .dout(n9528));
  jand g09273(.dina(n9326), .dinb(n9318), .dout(n9529));
  jand g09274(.dina(n9327), .dinb(n9256), .dout(n9530));
  jor  g09275(.dina(n9530), .dinb(n9529), .dout(n9531));
  jand g09276(.dina(n9316), .dinb(n9308), .dout(n9532));
  jand g09277(.dina(n9317), .dinb(n9259), .dout(n9533));
  jor  g09278(.dina(n9533), .dinb(n9532), .dout(n9534));
  jand g09279(.dina(n9306), .dinb(n9298), .dout(n9535));
  jand g09280(.dina(n9307), .dinb(n9262), .dout(n9536));
  jor  g09281(.dina(n9536), .dinb(n9535), .dout(n9537));
  jor  g09282(.dina(n9288), .dinb(n9280), .dout(n9538));
  jand g09283(.dina(n9297), .dinb(n9289), .dout(n9539));
  jnot g09284(.din(n9539), .dout(n9540));
  jand g09285(.dina(n9540), .dinb(n9538), .dout(n9541));
  jnot g09286(.din(n9541), .dout(n9542));
  jnot g09287(.din(n9263), .dout(n9543));
  jand g09288(.dina(n9265), .dinb(n9543), .dout(n9544));
  jand g09289(.dina(n9278), .dinb(n9267), .dout(n9545));
  jor  g09290(.dina(n9545), .dinb(n9544), .dout(n9546));
  jxor g09291(.dina(a62 ), .dinb(a61 ), .dout(n9547));
  jand g09292(.dina(n9547), .dinb(n9264), .dout(n9548));
  jand g09293(.dina(n9548), .dinb(n259), .dout(n9549));
  jnot g09294(.din(n9264), .dout(n9550));
  jxor g09295(.dina(a61 ), .dinb(a60 ), .dout(n9551));
  jand g09296(.dina(n9551), .dinb(n9550), .dout(n9552));
  jand g09297(.dina(n9552), .dinb(b0 ), .dout(n9553));
  jnot g09298(.din(n9547), .dout(n9554));
  jand g09299(.dina(n9554), .dinb(n9264), .dout(n9555));
  jand g09300(.dina(n9555), .dinb(b1 ), .dout(n9556));
  jor  g09301(.dina(n9556), .dinb(n9553), .dout(n9557));
  jor  g09302(.dina(n9557), .dinb(n9549), .dout(n9558));
  jnot g09303(.din(a62 ), .dout(n9559));
  jor  g09304(.dina(n9266), .dinb(n9559), .dout(n9560));
  jxor g09305(.dina(n9560), .dinb(n9558), .dout(n9561));
  jor  g09306(.dina(n9271), .dinb(n337), .dout(n9562));
  jor  g09307(.dina(n9268), .dinb(n340), .dout(n9563));
  jor  g09308(.dina(n9003), .dinb(n293), .dout(n9564));
  jand g09309(.dina(n9564), .dinb(n9563), .dout(n9565));
  jor  g09310(.dina(n9273), .dinb(n303), .dout(n9566));
  jand g09311(.dina(n9566), .dinb(n9565), .dout(n9567));
  jand g09312(.dina(n9567), .dinb(n9562), .dout(n9568));
  jxor g09313(.dina(n9568), .dinb(a59 ), .dout(n9569));
  jxor g09314(.dina(n9569), .dinb(n9561), .dout(n9570));
  jxor g09315(.dina(n9570), .dinb(n9546), .dout(n9571));
  jnot g09316(.din(n9571), .dout(n9572));
  jor  g09317(.dina(n8457), .dinb(n466), .dout(n9573));
  jor  g09318(.dina(n8454), .dinb(n469), .dout(n9574));
  jor  g09319(.dina(n8185), .dinb(n377), .dout(n9575));
  jand g09320(.dina(n9575), .dinb(n9574), .dout(n9576));
  jor  g09321(.dina(n8459), .dinb(n415), .dout(n9577));
  jand g09322(.dina(n9577), .dinb(n9576), .dout(n9578));
  jand g09323(.dina(n9578), .dinb(n9573), .dout(n9579));
  jxor g09324(.dina(n9579), .dinb(a56 ), .dout(n9580));
  jxor g09325(.dina(n9580), .dinb(n9572), .dout(n9581));
  jxor g09326(.dina(n9581), .dinb(n9542), .dout(n9582));
  jor  g09327(.dina(n7660), .dinb(n635), .dout(n9583));
  jor  g09328(.dina(n7415), .dinb(n519), .dout(n9584));
  jor  g09329(.dina(n7657), .dinb(n572), .dout(n9585));
  jor  g09330(.dina(n7662), .dinb(n637), .dout(n9586));
  jand g09331(.dina(n9586), .dinb(n9585), .dout(n9587));
  jand g09332(.dina(n9587), .dinb(n9584), .dout(n9588));
  jand g09333(.dina(n9588), .dinb(n9583), .dout(n9589));
  jxor g09334(.dina(n9589), .dinb(n7166), .dout(n9590));
  jxor g09335(.dina(n9590), .dinb(n9582), .dout(n9591));
  jxor g09336(.dina(n9591), .dinb(n9537), .dout(n9592));
  jor  g09337(.dina(n6914), .dinb(n850), .dout(n9593));
  jor  g09338(.dina(n6673), .dinb(n704), .dout(n9594));
  jor  g09339(.dina(n6911), .dinb(n772), .dout(n9595));
  jor  g09340(.dina(n6916), .dinb(n852), .dout(n9596));
  jand g09341(.dina(n9596), .dinb(n9595), .dout(n9597));
  jand g09342(.dina(n9597), .dinb(n9594), .dout(n9598));
  jand g09343(.dina(n9598), .dinb(n9593), .dout(n9599));
  jxor g09344(.dina(n9599), .dinb(n6443), .dout(n9600));
  jxor g09345(.dina(n9600), .dinb(n9592), .dout(n9601));
  jxor g09346(.dina(n9601), .dinb(n9534), .dout(n9602));
  jor  g09347(.dina(n6207), .dinb(n1112), .dout(n9603));
  jor  g09348(.dina(n5975), .dinb(n934), .dout(n9604));
  jor  g09349(.dina(n6205), .dinb(n1114), .dout(n9605));
  jor  g09350(.dina(n6210), .dinb(n1018), .dout(n9606));
  jand g09351(.dina(n9606), .dinb(n9605), .dout(n9607));
  jand g09352(.dina(n9607), .dinb(n9604), .dout(n9608));
  jand g09353(.dina(n9608), .dinb(n9603), .dout(n9609));
  jxor g09354(.dina(n9609), .dinb(n5759), .dout(n9610));
  jxor g09355(.dina(n9610), .dinb(n9602), .dout(n9611));
  jxor g09356(.dina(n9611), .dinb(n9531), .dout(n9612));
  jor  g09357(.dina(n5537), .dinb(n1414), .dout(n9613));
  jor  g09358(.dina(n5315), .dinb(n1211), .dout(n9614));
  jor  g09359(.dina(n5539), .dinb(n1416), .dout(n9615));
  jor  g09360(.dina(n5534), .dinb(n1307), .dout(n9616));
  jand g09361(.dina(n9616), .dinb(n9615), .dout(n9617));
  jand g09362(.dina(n9617), .dinb(n9614), .dout(n9618));
  jand g09363(.dina(n9618), .dinb(n9613), .dout(n9619));
  jxor g09364(.dina(n9619), .dinb(n5111), .dout(n9620));
  jxor g09365(.dina(n9620), .dinb(n9612), .dout(n9621));
  jxor g09366(.dina(n9621), .dinb(n9528), .dout(n9622));
  jor  g09367(.dina(n4902), .dinb(n1757), .dout(n9623));
  jor  g09368(.dina(n4696), .dinb(n1527), .dout(n9624));
  jor  g09369(.dina(n4904), .dinb(n1637), .dout(n9625));
  jor  g09370(.dina(n4899), .dinb(n1759), .dout(n9626));
  jand g09371(.dina(n9626), .dinb(n9625), .dout(n9627));
  jand g09372(.dina(n9627), .dinb(n9624), .dout(n9628));
  jand g09373(.dina(n9628), .dinb(n9623), .dout(n9629));
  jxor g09374(.dina(n9629), .dinb(n4505), .dout(n9630));
  jxor g09375(.dina(n9630), .dinb(n9622), .dout(n9631));
  jxor g09376(.dina(n9631), .dinb(n9525), .dout(n9632));
  jor  g09377(.dina(n4305), .dinb(n2140), .dout(n9633));
  jor  g09378(.dina(n4116), .dinb(n1881), .dout(n9634));
  jor  g09379(.dina(n4308), .dinb(n2007), .dout(n9635));
  jor  g09380(.dina(n4303), .dinb(n2142), .dout(n9636));
  jand g09381(.dina(n9636), .dinb(n9635), .dout(n9637));
  jand g09382(.dina(n9637), .dinb(n9634), .dout(n9638));
  jand g09383(.dina(n9638), .dinb(n9633), .dout(n9639));
  jxor g09384(.dina(n9639), .dinb(n3938), .dout(n9640));
  jxor g09385(.dina(n9640), .dinb(n9632), .dout(n9641));
  jxor g09386(.dina(n9641), .dinb(n9522), .dout(n9642));
  jor  g09387(.dina(n3751), .dinb(n2561), .dout(n9643));
  jor  g09388(.dina(n3574), .dinb(n2279), .dout(n9644));
  jor  g09389(.dina(n3754), .dinb(n2415), .dout(n9645));
  jor  g09390(.dina(n3749), .dinb(n2563), .dout(n9646));
  jand g09391(.dina(n9646), .dinb(n9645), .dout(n9647));
  jand g09392(.dina(n9647), .dinb(n9644), .dout(n9648));
  jand g09393(.dina(n9648), .dinb(n9643), .dout(n9649));
  jxor g09394(.dina(n9649), .dinb(n3410), .dout(n9650));
  jxor g09395(.dina(n9650), .dinb(n9642), .dout(n9651));
  jxor g09396(.dina(n9651), .dinb(n9519), .dout(n9652));
  jor  g09397(.dina(n3021), .dinb(n3239), .dout(n9653));
  jor  g09398(.dina(n3072), .dinb(n2713), .dout(n9654));
  jor  g09399(.dina(n3242), .dinb(n2862), .dout(n9655));
  jor  g09400(.dina(n3237), .dinb(n3023), .dout(n9656));
  jand g09401(.dina(n9656), .dinb(n9655), .dout(n9657));
  jand g09402(.dina(n9657), .dinb(n9654), .dout(n9658));
  jand g09403(.dina(n9658), .dinb(n9653), .dout(n9659));
  jxor g09404(.dina(n9659), .dinb(n2918), .dout(n9660));
  jxor g09405(.dina(n9660), .dinb(n9652), .dout(n9661));
  jxor g09406(.dina(n9661), .dinb(n9516), .dout(n9662));
  jor  g09407(.dina(n3520), .dinb(n2764), .dout(n9663));
  jor  g09408(.dina(n2609), .dinb(n3186), .dout(n9664));
  jor  g09409(.dina(n2761), .dinb(n3522), .dout(n9665));
  jor  g09410(.dina(n2766), .dinb(n3348), .dout(n9666));
  jand g09411(.dina(n9666), .dinb(n9665), .dout(n9667));
  jand g09412(.dina(n9667), .dinb(n9664), .dout(n9668));
  jand g09413(.dina(n9668), .dinb(n9663), .dout(n9669));
  jxor g09414(.dina(n9669), .dinb(n2468), .dout(n9670));
  jxor g09415(.dina(n9670), .dinb(n9662), .dout(n9671));
  jxor g09416(.dina(n9671), .dinb(n9513), .dout(n9672));
  jor  g09417(.dina(n4058), .dinb(n2324), .dout(n9673));
  jor  g09418(.dina(n2186), .dinb(n3698), .dout(n9674));
  jor  g09419(.dina(n2321), .dinb(n3873), .dout(n9675));
  jor  g09420(.dina(n2326), .dinb(n4060), .dout(n9676));
  jand g09421(.dina(n9676), .dinb(n9675), .dout(n9677));
  jand g09422(.dina(n9677), .dinb(n9674), .dout(n9678));
  jand g09423(.dina(n9678), .dinb(n9673), .dout(n9679));
  jxor g09424(.dina(n9679), .dinb(n2057), .dout(n9680));
  jxor g09425(.dina(n9680), .dinb(n9672), .dout(n9681));
  jxor g09426(.dina(n9681), .dinb(n9510), .dout(n9682));
  jor  g09427(.dina(n4635), .dinb(n1921), .dout(n9683));
  jor  g09428(.dina(n1806), .dinb(n4249), .dout(n9684));
  jor  g09429(.dina(n1923), .dinb(n4637), .dout(n9685));
  jor  g09430(.dina(n1918), .dinb(n4437), .dout(n9686));
  jand g09431(.dina(n9686), .dinb(n9685), .dout(n9687));
  jand g09432(.dina(n9687), .dinb(n9684), .dout(n9688));
  jand g09433(.dina(n9688), .dinb(n9683), .dout(n9689));
  jxor g09434(.dina(n9689), .dinb(n1687), .dout(n9690));
  jxor g09435(.dina(n9690), .dinb(n9682), .dout(n9691));
  jxor g09436(.dina(n9691), .dinb(n9507), .dout(n9692));
  jor  g09437(.dina(n5251), .dinb(n1569), .dout(n9693));
  jor  g09438(.dina(n1453), .dinb(n4839), .dout(n9694));
  jor  g09439(.dina(n1566), .dinb(n5040), .dout(n9695));
  jor  g09440(.dina(n1571), .dinb(n5253), .dout(n9696));
  jand g09441(.dina(n9696), .dinb(n9695), .dout(n9697));
  jand g09442(.dina(n9697), .dinb(n9694), .dout(n9698));
  jand g09443(.dina(n9698), .dinb(n9693), .dout(n9699));
  jxor g09444(.dina(n9699), .dinb(n1351), .dout(n9700));
  jxor g09445(.dina(n9700), .dinb(n9692), .dout(n9701));
  jxor g09446(.dina(n9701), .dinb(n9504), .dout(n9702));
  jor  g09447(.dina(n5909), .dinb(n1248), .dout(n9703));
  jor  g09448(.dina(n1147), .dinb(n5469), .dout(n9704));
  jor  g09449(.dina(n1251), .dinb(n5685), .dout(n9705));
  jor  g09450(.dina(n1246), .dinb(n5911), .dout(n9706));
  jand g09451(.dina(n9706), .dinb(n9705), .dout(n9707));
  jand g09452(.dina(n9707), .dinb(n9704), .dout(n9708));
  jand g09453(.dina(n9708), .dinb(n9703), .dout(n9709));
  jxor g09454(.dina(n9709), .dinb(n1061), .dout(n9710));
  jxor g09455(.dina(n9710), .dinb(n9702), .dout(n9711));
  jxor g09456(.dina(n9711), .dinb(n9501), .dout(n9712));
  jor  g09457(.dina(n6603), .dinb(n970), .dout(n9713));
  jor  g09458(.dina(n880), .dinb(n6139), .dout(n9714));
  jor  g09459(.dina(n967), .dinb(n6366), .dout(n9715));
  jor  g09460(.dina(n972), .dinb(n6605), .dout(n9716));
  jand g09461(.dina(n9716), .dinb(n9715), .dout(n9717));
  jand g09462(.dina(n9717), .dinb(n9714), .dout(n9718));
  jand g09463(.dina(n9718), .dinb(n9713), .dout(n9719));
  jxor g09464(.dina(n9719), .dinb(n810), .dout(n9720));
  jxor g09465(.dina(n9720), .dinb(n9712), .dout(n9721));
  jxor g09466(.dina(n9721), .dinb(n9498), .dout(n9722));
  jor  g09467(.dina(n7336), .dinb(n728), .dout(n9723));
  jor  g09468(.dina(n660), .dinb(n6846), .dout(n9724));
  jor  g09469(.dina(n726), .dinb(n7338), .dout(n9725));
  jor  g09470(.dina(n731), .dinb(n7086), .dout(n9726));
  jand g09471(.dina(n9726), .dinb(n9725), .dout(n9727));
  jand g09472(.dina(n9727), .dinb(n9724), .dout(n9728));
  jand g09473(.dina(n9728), .dinb(n9723), .dout(n9729));
  jxor g09474(.dina(n9729), .dinb(n606), .dout(n9730));
  jxor g09475(.dina(n9730), .dinb(n9722), .dout(n9731));
  jxor g09476(.dina(n9731), .dinb(n9495), .dout(n9732));
  jor  g09477(.dina(n8109), .dinb(n544), .dout(n9733));
  jor  g09478(.dina(n486), .dinb(n7590), .dout(n9734));
  jor  g09479(.dina(n547), .dinb(n7846), .dout(n9735));
  jor  g09480(.dina(n542), .dinb(n8111), .dout(n9736));
  jand g09481(.dina(n9736), .dinb(n9735), .dout(n9737));
  jand g09482(.dina(n9737), .dinb(n9734), .dout(n9738));
  jand g09483(.dina(n9738), .dinb(n9733), .dout(n9739));
  jxor g09484(.dina(n9739), .dinb(n446), .dout(n9740));
  jxor g09485(.dina(n9740), .dinb(n9732), .dout(n9741));
  jxor g09486(.dina(n9741), .dinb(n9492), .dout(n9742));
  jor  g09487(.dina(n8918), .dinb(n397), .dout(n9743));
  jor  g09488(.dina(n354), .dinb(n8378), .dout(n9744));
  jor  g09489(.dina(n394), .dinb(n8644), .dout(n9745));
  jor  g09490(.dina(n399), .dinb(n8920), .dout(n9746));
  jand g09491(.dina(n9746), .dinb(n9745), .dout(n9747));
  jand g09492(.dina(n9747), .dinb(n9744), .dout(n9748));
  jand g09493(.dina(n9748), .dinb(n9743), .dout(n9749));
  jxor g09494(.dina(n9749), .dinb(n364), .dout(n9750));
  jxor g09495(.dina(n9750), .dinb(n9742), .dout(n9751));
  jand g09496(.dina(b60 ), .dinb(b59 ), .dout(n9752));
  jand g09497(.dina(n9471), .dinb(n9470), .dout(n9753));
  jor  g09498(.dina(n9753), .dinb(n9752), .dout(n9754));
  jxor g09499(.dina(b61 ), .dinb(b60 ), .dout(n9755));
  jnot g09500(.din(n9755), .dout(n9756));
  jxor g09501(.dina(n9756), .dinb(n9754), .dout(n9757));
  jor  g09502(.dina(n9757), .dinb(n296), .dout(n9758));
  jnot g09503(.din(b61 ), .dout(n9759));
  jor  g09504(.dina(n264), .dinb(n9759), .dout(n9760));
  jor  g09505(.dina(n294), .dinb(n9475), .dout(n9761));
  jor  g09506(.dina(n280), .dinb(n9195), .dout(n9762));
  jand g09507(.dina(n9762), .dinb(n9761), .dout(n9763));
  jand g09508(.dina(n9763), .dinb(n9760), .dout(n9764));
  jand g09509(.dina(n9764), .dinb(n9758), .dout(n9765));
  jxor g09510(.dina(n9765), .dinb(n278), .dout(n9766));
  jxor g09511(.dina(n9766), .dinb(n9751), .dout(n9767));
  jxor g09512(.dina(n9767), .dinb(n9489), .dout(n9768));
  jand g09513(.dina(n9483), .dinb(n9213), .dout(n9769));
  jnot g09514(.din(n9769), .dout(n9770));
  jor  g09515(.dina(n9484), .dinb(n9210), .dout(n9771));
  jand g09516(.dina(n9771), .dinb(n9770), .dout(n9772));
  jxor g09517(.dina(n9772), .dinb(n9768), .dout(f61 ));
  jand g09518(.dina(n9767), .dinb(n9488), .dout(n9774));
  jnot g09519(.din(n9774), .dout(n9775));
  jor  g09520(.dina(n9772), .dinb(n9768), .dout(n9776));
  jand g09521(.dina(n9776), .dinb(n9775), .dout(n9777));
  jand g09522(.dina(n9750), .dinb(n9742), .dout(n9778));
  jand g09523(.dina(n9766), .dinb(n9751), .dout(n9779));
  jor  g09524(.dina(n9779), .dinb(n9778), .dout(n9780));
  jnot g09525(.din(n9780), .dout(n9781));
  jand g09526(.dina(n9740), .dinb(n9732), .dout(n9782));
  jand g09527(.dina(n9741), .dinb(n9492), .dout(n9783));
  jor  g09528(.dina(n9783), .dinb(n9782), .dout(n9784));
  jand g09529(.dina(n9730), .dinb(n9722), .dout(n9785));
  jand g09530(.dina(n9731), .dinb(n9495), .dout(n9786));
  jor  g09531(.dina(n9786), .dinb(n9785), .dout(n9787));
  jand g09532(.dina(n9720), .dinb(n9712), .dout(n9788));
  jand g09533(.dina(n9721), .dinb(n9498), .dout(n9789));
  jor  g09534(.dina(n9789), .dinb(n9788), .dout(n9790));
  jand g09535(.dina(n9710), .dinb(n9702), .dout(n9791));
  jand g09536(.dina(n9711), .dinb(n9501), .dout(n9792));
  jor  g09537(.dina(n9792), .dinb(n9791), .dout(n9793));
  jand g09538(.dina(n9700), .dinb(n9692), .dout(n9794));
  jand g09539(.dina(n9701), .dinb(n9504), .dout(n9795));
  jor  g09540(.dina(n9795), .dinb(n9794), .dout(n9796));
  jand g09541(.dina(n9690), .dinb(n9682), .dout(n9797));
  jand g09542(.dina(n9691), .dinb(n9507), .dout(n9798));
  jor  g09543(.dina(n9798), .dinb(n9797), .dout(n9799));
  jand g09544(.dina(n9680), .dinb(n9672), .dout(n9800));
  jand g09545(.dina(n9681), .dinb(n9510), .dout(n9801));
  jor  g09546(.dina(n9801), .dinb(n9800), .dout(n9802));
  jand g09547(.dina(n9670), .dinb(n9662), .dout(n9803));
  jand g09548(.dina(n9671), .dinb(n9513), .dout(n9804));
  jor  g09549(.dina(n9804), .dinb(n9803), .dout(n9805));
  jand g09550(.dina(n9660), .dinb(n9652), .dout(n9806));
  jand g09551(.dina(n9661), .dinb(n9516), .dout(n9807));
  jor  g09552(.dina(n9807), .dinb(n9806), .dout(n9808));
  jand g09553(.dina(n9650), .dinb(n9642), .dout(n9809));
  jand g09554(.dina(n9651), .dinb(n9519), .dout(n9810));
  jor  g09555(.dina(n9810), .dinb(n9809), .dout(n9811));
  jand g09556(.dina(n9640), .dinb(n9632), .dout(n9812));
  jand g09557(.dina(n9641), .dinb(n9522), .dout(n9813));
  jor  g09558(.dina(n9813), .dinb(n9812), .dout(n9814));
  jand g09559(.dina(n9630), .dinb(n9622), .dout(n9815));
  jand g09560(.dina(n9631), .dinb(n9525), .dout(n9816));
  jor  g09561(.dina(n9816), .dinb(n9815), .dout(n9817));
  jand g09562(.dina(n9620), .dinb(n9612), .dout(n9818));
  jand g09563(.dina(n9621), .dinb(n9528), .dout(n9819));
  jor  g09564(.dina(n9819), .dinb(n9818), .dout(n9820));
  jand g09565(.dina(n9610), .dinb(n9602), .dout(n9821));
  jand g09566(.dina(n9611), .dinb(n9531), .dout(n9822));
  jor  g09567(.dina(n9822), .dinb(n9821), .dout(n9823));
  jand g09568(.dina(n9600), .dinb(n9592), .dout(n9824));
  jand g09569(.dina(n9601), .dinb(n9534), .dout(n9825));
  jor  g09570(.dina(n9825), .dinb(n9824), .dout(n9826));
  jand g09571(.dina(n9590), .dinb(n9582), .dout(n9827));
  jand g09572(.dina(n9591), .dinb(n9537), .dout(n9828));
  jor  g09573(.dina(n9828), .dinb(n9827), .dout(n9829));
  jor  g09574(.dina(n9580), .dinb(n9572), .dout(n9830));
  jand g09575(.dina(n9581), .dinb(n9542), .dout(n9831));
  jnot g09576(.din(n9831), .dout(n9832));
  jand g09577(.dina(n9832), .dinb(n9830), .dout(n9833));
  jnot g09578(.din(n9833), .dout(n9834));
  jor  g09579(.dina(n8457), .dinb(n517), .dout(n9835));
  jor  g09580(.dina(n8454), .dinb(n519), .dout(n9836));
  jor  g09581(.dina(n8459), .dinb(n469), .dout(n9837));
  jor  g09582(.dina(n8185), .dinb(n415), .dout(n9838));
  jand g09583(.dina(n9838), .dinb(n9837), .dout(n9839));
  jand g09584(.dina(n9839), .dinb(n9836), .dout(n9840));
  jand g09585(.dina(n9840), .dinb(n9835), .dout(n9841));
  jxor g09586(.dina(n9841), .dinb(n7929), .dout(n9842));
  jor  g09587(.dina(n9569), .dinb(n9561), .dout(n9843));
  jand g09588(.dina(n9570), .dinb(n9546), .dout(n9844));
  jnot g09589(.din(n9844), .dout(n9845));
  jand g09590(.dina(n9845), .dinb(n9843), .dout(n9846));
  jand g09591(.dina(n9552), .dinb(b1 ), .dout(n9847));
  jor  g09592(.dina(n9551), .dinb(n9264), .dout(n9848));
  jor  g09593(.dina(n9848), .dinb(n9554), .dout(n9849));
  jnot g09594(.din(n9849), .dout(n9850));
  jand g09595(.dina(n9850), .dinb(b0 ), .dout(n9851));
  jand g09596(.dina(n9548), .dinb(n273), .dout(n9852));
  jand g09597(.dina(n9555), .dinb(b2 ), .dout(n9853));
  jor  g09598(.dina(n9853), .dinb(n9852), .dout(n9854));
  jor  g09599(.dina(n9854), .dinb(n9851), .dout(n9855));
  jor  g09600(.dina(n9855), .dinb(n9847), .dout(n9856));
  jnot g09601(.din(n9558), .dout(n9857));
  jand g09602(.dina(n9266), .dinb(a62 ), .dout(n9858));
  jand g09603(.dina(n9858), .dinb(n9857), .dout(n9859));
  jnot g09604(.din(n9859), .dout(n9860));
  jand g09605(.dina(n9860), .dinb(a62 ), .dout(n9861));
  jxor g09606(.dina(n9861), .dinb(n9856), .dout(n9862));
  jor  g09607(.dina(n9271), .dinb(n374), .dout(n9863));
  jor  g09608(.dina(n9268), .dinb(n377), .dout(n9864));
  jor  g09609(.dina(n9003), .dinb(n303), .dout(n9865));
  jand g09610(.dina(n9865), .dinb(n9864), .dout(n9866));
  jor  g09611(.dina(n9273), .dinb(n340), .dout(n9867));
  jand g09612(.dina(n9867), .dinb(n9866), .dout(n9868));
  jand g09613(.dina(n9868), .dinb(n9863), .dout(n9869));
  jxor g09614(.dina(n9869), .dinb(a59 ), .dout(n9870));
  jxor g09615(.dina(n9870), .dinb(n9862), .dout(n9871));
  jxor g09616(.dina(n9871), .dinb(n9846), .dout(n9872));
  jxor g09617(.dina(n9872), .dinb(n9842), .dout(n9873));
  jxor g09618(.dina(n9873), .dinb(n9834), .dout(n9874));
  jor  g09619(.dina(n7660), .dinb(n702), .dout(n9875));
  jor  g09620(.dina(n7415), .dinb(n572), .dout(n9876));
  jor  g09621(.dina(n7657), .dinb(n637), .dout(n9877));
  jor  g09622(.dina(n7662), .dinb(n704), .dout(n9878));
  jand g09623(.dina(n9878), .dinb(n9877), .dout(n9879));
  jand g09624(.dina(n9879), .dinb(n9876), .dout(n9880));
  jand g09625(.dina(n9880), .dinb(n9875), .dout(n9881));
  jxor g09626(.dina(n9881), .dinb(n7166), .dout(n9882));
  jxor g09627(.dina(n9882), .dinb(n9874), .dout(n9883));
  jxor g09628(.dina(n9883), .dinb(n9829), .dout(n9884));
  jor  g09629(.dina(n6914), .dinb(n932), .dout(n9885));
  jor  g09630(.dina(n6673), .dinb(n772), .dout(n9886));
  jor  g09631(.dina(n6911), .dinb(n852), .dout(n9887));
  jor  g09632(.dina(n6916), .dinb(n934), .dout(n9888));
  jand g09633(.dina(n9888), .dinb(n9887), .dout(n9889));
  jand g09634(.dina(n9889), .dinb(n9886), .dout(n9890));
  jand g09635(.dina(n9890), .dinb(n9885), .dout(n9891));
  jxor g09636(.dina(n9891), .dinb(n6443), .dout(n9892));
  jxor g09637(.dina(n9892), .dinb(n9884), .dout(n9893));
  jxor g09638(.dina(n9893), .dinb(n9826), .dout(n9894));
  jor  g09639(.dina(n6207), .dinb(n1209), .dout(n9895));
  jor  g09640(.dina(n5975), .dinb(n1018), .dout(n9896));
  jor  g09641(.dina(n6205), .dinb(n1211), .dout(n9897));
  jor  g09642(.dina(n6210), .dinb(n1114), .dout(n9898));
  jand g09643(.dina(n9898), .dinb(n9897), .dout(n9899));
  jand g09644(.dina(n9899), .dinb(n9896), .dout(n9900));
  jand g09645(.dina(n9900), .dinb(n9895), .dout(n9901));
  jxor g09646(.dina(n9901), .dinb(n5759), .dout(n9902));
  jxor g09647(.dina(n9902), .dinb(n9894), .dout(n9903));
  jxor g09648(.dina(n9903), .dinb(n9823), .dout(n9904));
  jor  g09649(.dina(n5537), .dinb(n1525), .dout(n9905));
  jor  g09650(.dina(n5315), .dinb(n1307), .dout(n9906));
  jor  g09651(.dina(n5539), .dinb(n1527), .dout(n9907));
  jor  g09652(.dina(n5534), .dinb(n1416), .dout(n9908));
  jand g09653(.dina(n9908), .dinb(n9907), .dout(n9909));
  jand g09654(.dina(n9909), .dinb(n9906), .dout(n9910));
  jand g09655(.dina(n9910), .dinb(n9905), .dout(n9911));
  jxor g09656(.dina(n9911), .dinb(n5111), .dout(n9912));
  jxor g09657(.dina(n9912), .dinb(n9904), .dout(n9913));
  jxor g09658(.dina(n9913), .dinb(n9820), .dout(n9914));
  jor  g09659(.dina(n4902), .dinb(n1879), .dout(n9915));
  jor  g09660(.dina(n4696), .dinb(n1637), .dout(n9916));
  jor  g09661(.dina(n4904), .dinb(n1759), .dout(n9917));
  jor  g09662(.dina(n4899), .dinb(n1881), .dout(n9918));
  jand g09663(.dina(n9918), .dinb(n9917), .dout(n9919));
  jand g09664(.dina(n9919), .dinb(n9916), .dout(n9920));
  jand g09665(.dina(n9920), .dinb(n9915), .dout(n9921));
  jxor g09666(.dina(n9921), .dinb(n4505), .dout(n9922));
  jxor g09667(.dina(n9922), .dinb(n9914), .dout(n9923));
  jxor g09668(.dina(n9923), .dinb(n9817), .dout(n9924));
  jor  g09669(.dina(n4305), .dinb(n2277), .dout(n9925));
  jor  g09670(.dina(n4116), .dinb(n2007), .dout(n9926));
  jor  g09671(.dina(n4308), .dinb(n2142), .dout(n9927));
  jor  g09672(.dina(n4303), .dinb(n2279), .dout(n9928));
  jand g09673(.dina(n9928), .dinb(n9927), .dout(n9929));
  jand g09674(.dina(n9929), .dinb(n9926), .dout(n9930));
  jand g09675(.dina(n9930), .dinb(n9925), .dout(n9931));
  jxor g09676(.dina(n9931), .dinb(n3938), .dout(n9932));
  jxor g09677(.dina(n9932), .dinb(n9924), .dout(n9933));
  jxor g09678(.dina(n9933), .dinb(n9814), .dout(n9934));
  jor  g09679(.dina(n3751), .dinb(n2711), .dout(n9935));
  jor  g09680(.dina(n3574), .dinb(n2415), .dout(n9936));
  jor  g09681(.dina(n3754), .dinb(n2563), .dout(n9937));
  jor  g09682(.dina(n3749), .dinb(n2713), .dout(n9938));
  jand g09683(.dina(n9938), .dinb(n9937), .dout(n9939));
  jand g09684(.dina(n9939), .dinb(n9936), .dout(n9940));
  jand g09685(.dina(n9940), .dinb(n9935), .dout(n9941));
  jxor g09686(.dina(n9941), .dinb(n3410), .dout(n9942));
  jxor g09687(.dina(n9942), .dinb(n9934), .dout(n9943));
  jxor g09688(.dina(n9943), .dinb(n9811), .dout(n9944));
  jor  g09689(.dina(n3184), .dinb(n3239), .dout(n9945));
  jor  g09690(.dina(n3072), .dinb(n2862), .dout(n9946));
  jor  g09691(.dina(n3242), .dinb(n3023), .dout(n9947));
  jor  g09692(.dina(n3237), .dinb(n3186), .dout(n9948));
  jand g09693(.dina(n9948), .dinb(n9947), .dout(n9949));
  jand g09694(.dina(n9949), .dinb(n9946), .dout(n9950));
  jand g09695(.dina(n9950), .dinb(n9945), .dout(n9951));
  jxor g09696(.dina(n9951), .dinb(n2918), .dout(n9952));
  jxor g09697(.dina(n9952), .dinb(n9944), .dout(n9953));
  jxor g09698(.dina(n9953), .dinb(n9808), .dout(n9954));
  jor  g09699(.dina(n3696), .dinb(n2764), .dout(n9955));
  jor  g09700(.dina(n2609), .dinb(n3348), .dout(n9956));
  jor  g09701(.dina(n2761), .dinb(n3698), .dout(n9957));
  jor  g09702(.dina(n2766), .dinb(n3522), .dout(n9958));
  jand g09703(.dina(n9958), .dinb(n9957), .dout(n9959));
  jand g09704(.dina(n9959), .dinb(n9956), .dout(n9960));
  jand g09705(.dina(n9960), .dinb(n9955), .dout(n9961));
  jxor g09706(.dina(n9961), .dinb(n2468), .dout(n9962));
  jxor g09707(.dina(n9962), .dinb(n9954), .dout(n9963));
  jxor g09708(.dina(n9963), .dinb(n9805), .dout(n9964));
  jor  g09709(.dina(n4247), .dinb(n2324), .dout(n9965));
  jor  g09710(.dina(n2186), .dinb(n3873), .dout(n9966));
  jor  g09711(.dina(n2321), .dinb(n4060), .dout(n9967));
  jor  g09712(.dina(n2326), .dinb(n4249), .dout(n9968));
  jand g09713(.dina(n9968), .dinb(n9967), .dout(n9969));
  jand g09714(.dina(n9969), .dinb(n9966), .dout(n9970));
  jand g09715(.dina(n9970), .dinb(n9965), .dout(n9971));
  jxor g09716(.dina(n9971), .dinb(n2057), .dout(n9972));
  jxor g09717(.dina(n9972), .dinb(n9964), .dout(n9973));
  jxor g09718(.dina(n9973), .dinb(n9802), .dout(n9974));
  jor  g09719(.dina(n4837), .dinb(n1921), .dout(n9975));
  jor  g09720(.dina(n1806), .dinb(n4437), .dout(n9976));
  jor  g09721(.dina(n1918), .dinb(n4637), .dout(n9977));
  jor  g09722(.dina(n1923), .dinb(n4839), .dout(n9978));
  jand g09723(.dina(n9978), .dinb(n9977), .dout(n9979));
  jand g09724(.dina(n9979), .dinb(n9976), .dout(n9980));
  jand g09725(.dina(n9980), .dinb(n9975), .dout(n9981));
  jxor g09726(.dina(n9981), .dinb(n1687), .dout(n9982));
  jxor g09727(.dina(n9982), .dinb(n9974), .dout(n9983));
  jxor g09728(.dina(n9983), .dinb(n9799), .dout(n9984));
  jor  g09729(.dina(n5467), .dinb(n1569), .dout(n9985));
  jor  g09730(.dina(n1453), .dinb(n5040), .dout(n9986));
  jor  g09731(.dina(n1571), .dinb(n5469), .dout(n9987));
  jor  g09732(.dina(n1566), .dinb(n5253), .dout(n9988));
  jand g09733(.dina(n9988), .dinb(n9987), .dout(n9989));
  jand g09734(.dina(n9989), .dinb(n9986), .dout(n9990));
  jand g09735(.dina(n9990), .dinb(n9985), .dout(n9991));
  jxor g09736(.dina(n9991), .dinb(n1351), .dout(n9992));
  jxor g09737(.dina(n9992), .dinb(n9984), .dout(n9993));
  jxor g09738(.dina(n9993), .dinb(n9796), .dout(n9994));
  jor  g09739(.dina(n6137), .dinb(n1248), .dout(n9995));
  jor  g09740(.dina(n1147), .dinb(n5685), .dout(n9996));
  jor  g09741(.dina(n1251), .dinb(n5911), .dout(n9997));
  jor  g09742(.dina(n1246), .dinb(n6139), .dout(n9998));
  jand g09743(.dina(n9998), .dinb(n9997), .dout(n9999));
  jand g09744(.dina(n9999), .dinb(n9996), .dout(n10000));
  jand g09745(.dina(n10000), .dinb(n9995), .dout(n10001));
  jxor g09746(.dina(n10001), .dinb(n1061), .dout(n10002));
  jxor g09747(.dina(n10002), .dinb(n9994), .dout(n10003));
  jxor g09748(.dina(n10003), .dinb(n9793), .dout(n10004));
  jor  g09749(.dina(n6844), .dinb(n970), .dout(n10005));
  jor  g09750(.dina(n880), .dinb(n6366), .dout(n10006));
  jor  g09751(.dina(n967), .dinb(n6605), .dout(n10007));
  jor  g09752(.dina(n972), .dinb(n6846), .dout(n10008));
  jand g09753(.dina(n10008), .dinb(n10007), .dout(n10009));
  jand g09754(.dina(n10009), .dinb(n10006), .dout(n10010));
  jand g09755(.dina(n10010), .dinb(n10005), .dout(n10011));
  jxor g09756(.dina(n10011), .dinb(n810), .dout(n10012));
  jxor g09757(.dina(n10012), .dinb(n10004), .dout(n10013));
  jxor g09758(.dina(n10013), .dinb(n9790), .dout(n10014));
  jor  g09759(.dina(n7588), .dinb(n728), .dout(n10015));
  jor  g09760(.dina(n660), .dinb(n7086), .dout(n10016));
  jor  g09761(.dina(n731), .dinb(n7338), .dout(n10017));
  jor  g09762(.dina(n726), .dinb(n7590), .dout(n10018));
  jand g09763(.dina(n10018), .dinb(n10017), .dout(n10019));
  jand g09764(.dina(n10019), .dinb(n10016), .dout(n10020));
  jand g09765(.dina(n10020), .dinb(n10015), .dout(n10021));
  jxor g09766(.dina(n10021), .dinb(n606), .dout(n10022));
  jxor g09767(.dina(n10022), .dinb(n10014), .dout(n10023));
  jxor g09768(.dina(n10023), .dinb(n9787), .dout(n10024));
  jor  g09769(.dina(n8376), .dinb(n544), .dout(n10025));
  jor  g09770(.dina(n486), .dinb(n7846), .dout(n10026));
  jor  g09771(.dina(n547), .dinb(n8111), .dout(n10027));
  jor  g09772(.dina(n542), .dinb(n8378), .dout(n10028));
  jand g09773(.dina(n10028), .dinb(n10027), .dout(n10029));
  jand g09774(.dina(n10029), .dinb(n10026), .dout(n10030));
  jand g09775(.dina(n10030), .dinb(n10025), .dout(n10031));
  jxor g09776(.dina(n10031), .dinb(n446), .dout(n10032));
  jxor g09777(.dina(n10032), .dinb(n10024), .dout(n10033));
  jor  g09778(.dina(n9193), .dinb(n397), .dout(n10034));
  jor  g09779(.dina(n354), .dinb(n8644), .dout(n10035));
  jor  g09780(.dina(n394), .dinb(n8920), .dout(n10036));
  jor  g09781(.dina(n399), .dinb(n9195), .dout(n10037));
  jand g09782(.dina(n10037), .dinb(n10036), .dout(n10038));
  jand g09783(.dina(n10038), .dinb(n10035), .dout(n10039));
  jand g09784(.dina(n10039), .dinb(n10034), .dout(n10040));
  jxor g09785(.dina(n10040), .dinb(n364), .dout(n10041));
  jxor g09786(.dina(n10041), .dinb(n10033), .dout(n10042));
  jxor g09787(.dina(n10042), .dinb(n9784), .dout(n10043));
  jand g09788(.dina(b61 ), .dinb(b60 ), .dout(n10044));
  jand g09789(.dina(n9755), .dinb(n9754), .dout(n10045));
  jor  g09790(.dina(n10045), .dinb(n10044), .dout(n10046));
  jxor g09791(.dina(b62 ), .dinb(b61 ), .dout(n10047));
  jnot g09792(.din(n10047), .dout(n10048));
  jxor g09793(.dina(n10048), .dinb(n10046), .dout(n10049));
  jor  g09794(.dina(n10049), .dinb(n296), .dout(n10050));
  jnot g09795(.din(b62 ), .dout(n10051));
  jor  g09796(.dina(n264), .dinb(n10051), .dout(n10052));
  jor  g09797(.dina(n280), .dinb(n9475), .dout(n10053));
  jor  g09798(.dina(n294), .dinb(n9759), .dout(n10054));
  jand g09799(.dina(n10054), .dinb(n10053), .dout(n10055));
  jand g09800(.dina(n10055), .dinb(n10052), .dout(n10056));
  jand g09801(.dina(n10056), .dinb(n10050), .dout(n10057));
  jxor g09802(.dina(n10057), .dinb(n278), .dout(n10058));
  jxor g09803(.dina(n10058), .dinb(n10043), .dout(n10059));
  jxor g09804(.dina(n10059), .dinb(n9781), .dout(n10060));
  jxor g09805(.dina(n10060), .dinb(n9777), .dout(f62 ));
  jand g09806(.dina(n10059), .dinb(n9780), .dout(n10062));
  jnot g09807(.din(n10062), .dout(n10063));
  jor  g09808(.dina(n10060), .dinb(n9777), .dout(n10064));
  jand g09809(.dina(n10064), .dinb(n10063), .dout(n10065));
  jand g09810(.dina(n10042), .dinb(n9784), .dout(n10066));
  jand g09811(.dina(n10058), .dinb(n10043), .dout(n10067));
  jor  g09812(.dina(n10067), .dinb(n10066), .dout(n10068));
  jnot g09813(.din(n10068), .dout(n10069));
  jand g09814(.dina(n10032), .dinb(n10024), .dout(n10070));
  jand g09815(.dina(n10041), .dinb(n10033), .dout(n10071));
  jor  g09816(.dina(n10071), .dinb(n10070), .dout(n10072));
  jand g09817(.dina(n10022), .dinb(n10014), .dout(n10073));
  jand g09818(.dina(n10023), .dinb(n9787), .dout(n10074));
  jor  g09819(.dina(n10074), .dinb(n10073), .dout(n10075));
  jand g09820(.dina(n10012), .dinb(n10004), .dout(n10076));
  jand g09821(.dina(n10013), .dinb(n9790), .dout(n10077));
  jor  g09822(.dina(n10077), .dinb(n10076), .dout(n10078));
  jand g09823(.dina(n10002), .dinb(n9994), .dout(n10079));
  jand g09824(.dina(n10003), .dinb(n9793), .dout(n10080));
  jor  g09825(.dina(n10080), .dinb(n10079), .dout(n10081));
  jand g09826(.dina(n9992), .dinb(n9984), .dout(n10082));
  jand g09827(.dina(n9993), .dinb(n9796), .dout(n10083));
  jor  g09828(.dina(n10083), .dinb(n10082), .dout(n10084));
  jand g09829(.dina(n9982), .dinb(n9974), .dout(n10085));
  jand g09830(.dina(n9983), .dinb(n9799), .dout(n10086));
  jor  g09831(.dina(n10086), .dinb(n10085), .dout(n10087));
  jand g09832(.dina(n9972), .dinb(n9964), .dout(n10088));
  jand g09833(.dina(n9973), .dinb(n9802), .dout(n10089));
  jor  g09834(.dina(n10089), .dinb(n10088), .dout(n10090));
  jand g09835(.dina(n9962), .dinb(n9954), .dout(n10091));
  jand g09836(.dina(n9963), .dinb(n9805), .dout(n10092));
  jor  g09837(.dina(n10092), .dinb(n10091), .dout(n10093));
  jand g09838(.dina(n9952), .dinb(n9944), .dout(n10094));
  jand g09839(.dina(n9953), .dinb(n9808), .dout(n10095));
  jor  g09840(.dina(n10095), .dinb(n10094), .dout(n10096));
  jand g09841(.dina(n9932), .dinb(n9924), .dout(n10097));
  jand g09842(.dina(n9933), .dinb(n9814), .dout(n10098));
  jor  g09843(.dina(n10098), .dinb(n10097), .dout(n10099));
  jand g09844(.dina(n9922), .dinb(n9914), .dout(n10100));
  jand g09845(.dina(n9923), .dinb(n9817), .dout(n10101));
  jor  g09846(.dina(n10101), .dinb(n10100), .dout(n10102));
  jand g09847(.dina(n9912), .dinb(n9904), .dout(n10103));
  jand g09848(.dina(n9913), .dinb(n9820), .dout(n10104));
  jor  g09849(.dina(n10104), .dinb(n10103), .dout(n10105));
  jand g09850(.dina(n9902), .dinb(n9894), .dout(n10106));
  jand g09851(.dina(n9903), .dinb(n9823), .dout(n10107));
  jor  g09852(.dina(n10107), .dinb(n10106), .dout(n10108));
  jand g09853(.dina(n9892), .dinb(n9884), .dout(n10109));
  jand g09854(.dina(n9893), .dinb(n9826), .dout(n10110));
  jor  g09855(.dina(n10110), .dinb(n10109), .dout(n10111));
  jand g09856(.dina(n9882), .dinb(n9874), .dout(n10112));
  jand g09857(.dina(n9883), .dinb(n9829), .dout(n10113));
  jor  g09858(.dina(n10113), .dinb(n10112), .dout(n10114));
  jand g09859(.dina(n9872), .dinb(n9842), .dout(n10115));
  jand g09860(.dina(n9873), .dinb(n9834), .dout(n10116));
  jor  g09861(.dina(n10116), .dinb(n10115), .dout(n10117));
  jnot g09862(.din(n9870), .dout(n10118));
  jand g09863(.dina(n10118), .dinb(n9862), .dout(n10119));
  jnot g09864(.din(n10119), .dout(n10120));
  jnot g09865(.din(n9862), .dout(n10121));
  jand g09866(.dina(n9870), .dinb(n10121), .dout(n10122));
  jor  g09867(.dina(n10122), .dinb(n9846), .dout(n10123));
  jand g09868(.dina(n10123), .dinb(n10120), .dout(n10124));
  jnot g09869(.din(n10124), .dout(n10125));
  jor  g09870(.dina(n9860), .dinb(n9856), .dout(n10126));
  jnot g09871(.din(n10126), .dout(n10127));
  jxor g09872(.dina(a63 ), .dinb(n9559), .dout(n10128));
  jnot g09873(.din(n10128), .dout(n10129));
  jand g09874(.dina(n10129), .dinb(b0 ), .dout(n10130));
  jxor g09875(.dina(n10130), .dinb(n10127), .dout(n10131));
  jnot g09876(.din(n9555), .dout(n10132));
  jor  g09877(.dina(n10132), .dinb(n303), .dout(n10133));
  jnot g09878(.din(n9548), .dout(n10134));
  jor  g09879(.dina(n10134), .dinb(n301), .dout(n10135));
  jor  g09880(.dina(n9849), .dinb(n305), .dout(n10136));
  jnot g09881(.din(n9552), .dout(n10137));
  jor  g09882(.dina(n10137), .dinb(n293), .dout(n10138));
  jand g09883(.dina(n10138), .dinb(n10136), .dout(n10139));
  jand g09884(.dina(n10139), .dinb(n10135), .dout(n10140));
  jand g09885(.dina(n10140), .dinb(n10133), .dout(n10141));
  jxor g09886(.dina(n10141), .dinb(n9559), .dout(n10142));
  jxor g09887(.dina(n10142), .dinb(n10131), .dout(n10143));
  jnot g09888(.din(n10143), .dout(n10144));
  jor  g09889(.dina(n9271), .dinb(n412), .dout(n10145));
  jor  g09890(.dina(n9273), .dinb(n377), .dout(n10146));
  jor  g09891(.dina(n9003), .dinb(n340), .dout(n10147));
  jand g09892(.dina(n10147), .dinb(n10146), .dout(n10148));
  jor  g09893(.dina(n9268), .dinb(n415), .dout(n10149));
  jand g09894(.dina(n10149), .dinb(n10148), .dout(n10150));
  jand g09895(.dina(n10150), .dinb(n10145), .dout(n10151));
  jxor g09896(.dina(n10151), .dinb(a59 ), .dout(n10152));
  jxor g09897(.dina(n10152), .dinb(n10144), .dout(n10153));
  jxor g09898(.dina(n10153), .dinb(n10125), .dout(n10154));
  jor  g09899(.dina(n8457), .dinb(n570), .dout(n10155));
  jor  g09900(.dina(n8185), .dinb(n469), .dout(n10156));
  jor  g09901(.dina(n8454), .dinb(n572), .dout(n10157));
  jor  g09902(.dina(n8459), .dinb(n519), .dout(n10158));
  jand g09903(.dina(n10158), .dinb(n10157), .dout(n10159));
  jand g09904(.dina(n10159), .dinb(n10156), .dout(n10160));
  jand g09905(.dina(n10160), .dinb(n10155), .dout(n10161));
  jxor g09906(.dina(n10161), .dinb(n7929), .dout(n10162));
  jxor g09907(.dina(n10162), .dinb(n10154), .dout(n10163));
  jxor g09908(.dina(n10163), .dinb(n10117), .dout(n10164));
  jor  g09909(.dina(n7660), .dinb(n770), .dout(n10165));
  jor  g09910(.dina(n7415), .dinb(n637), .dout(n10166));
  jor  g09911(.dina(n7657), .dinb(n704), .dout(n10167));
  jor  g09912(.dina(n7662), .dinb(n772), .dout(n10168));
  jand g09913(.dina(n10168), .dinb(n10167), .dout(n10169));
  jand g09914(.dina(n10169), .dinb(n10166), .dout(n10170));
  jand g09915(.dina(n10170), .dinb(n10165), .dout(n10171));
  jxor g09916(.dina(n10171), .dinb(n7166), .dout(n10172));
  jxor g09917(.dina(n10172), .dinb(n10164), .dout(n10173));
  jxor g09918(.dina(n10173), .dinb(n10114), .dout(n10174));
  jor  g09919(.dina(n6914), .dinb(n1016), .dout(n10175));
  jor  g09920(.dina(n6673), .dinb(n852), .dout(n10176));
  jor  g09921(.dina(n6911), .dinb(n934), .dout(n10177));
  jor  g09922(.dina(n6916), .dinb(n1018), .dout(n10178));
  jand g09923(.dina(n10178), .dinb(n10177), .dout(n10179));
  jand g09924(.dina(n10179), .dinb(n10176), .dout(n10180));
  jand g09925(.dina(n10180), .dinb(n10175), .dout(n10181));
  jxor g09926(.dina(n10181), .dinb(n6443), .dout(n10182));
  jxor g09927(.dina(n10182), .dinb(n10174), .dout(n10183));
  jxor g09928(.dina(n10183), .dinb(n10111), .dout(n10184));
  jor  g09929(.dina(n6207), .dinb(n1305), .dout(n10185));
  jor  g09930(.dina(n5975), .dinb(n1114), .dout(n10186));
  jor  g09931(.dina(n6210), .dinb(n1211), .dout(n10187));
  jor  g09932(.dina(n6205), .dinb(n1307), .dout(n10188));
  jand g09933(.dina(n10188), .dinb(n10187), .dout(n10189));
  jand g09934(.dina(n10189), .dinb(n10186), .dout(n10190));
  jand g09935(.dina(n10190), .dinb(n10185), .dout(n10191));
  jxor g09936(.dina(n10191), .dinb(n5759), .dout(n10192));
  jxor g09937(.dina(n10192), .dinb(n10184), .dout(n10193));
  jxor g09938(.dina(n10193), .dinb(n10108), .dout(n10194));
  jor  g09939(.dina(n5537), .dinb(n1635), .dout(n10195));
  jor  g09940(.dina(n5315), .dinb(n1416), .dout(n10196));
  jor  g09941(.dina(n5534), .dinb(n1527), .dout(n10197));
  jor  g09942(.dina(n5539), .dinb(n1637), .dout(n10198));
  jand g09943(.dina(n10198), .dinb(n10197), .dout(n10199));
  jand g09944(.dina(n10199), .dinb(n10196), .dout(n10200));
  jand g09945(.dina(n10200), .dinb(n10195), .dout(n10201));
  jxor g09946(.dina(n10201), .dinb(n5111), .dout(n10202));
  jxor g09947(.dina(n10202), .dinb(n10194), .dout(n10203));
  jxor g09948(.dina(n10203), .dinb(n10105), .dout(n10204));
  jor  g09949(.dina(n4902), .dinb(n2005), .dout(n10205));
  jor  g09950(.dina(n4696), .dinb(n1759), .dout(n10206));
  jor  g09951(.dina(n4904), .dinb(n1881), .dout(n10207));
  jor  g09952(.dina(n4899), .dinb(n2007), .dout(n10208));
  jand g09953(.dina(n10208), .dinb(n10207), .dout(n10209));
  jand g09954(.dina(n10209), .dinb(n10206), .dout(n10210));
  jand g09955(.dina(n10210), .dinb(n10205), .dout(n10211));
  jxor g09956(.dina(n10211), .dinb(n4505), .dout(n10212));
  jxor g09957(.dina(n10212), .dinb(n10204), .dout(n10213));
  jxor g09958(.dina(n10213), .dinb(n10102), .dout(n10214));
  jor  g09959(.dina(n4305), .dinb(n2413), .dout(n10215));
  jor  g09960(.dina(n4116), .dinb(n2142), .dout(n10216));
  jor  g09961(.dina(n4308), .dinb(n2279), .dout(n10217));
  jor  g09962(.dina(n4303), .dinb(n2415), .dout(n10218));
  jand g09963(.dina(n10218), .dinb(n10217), .dout(n10219));
  jand g09964(.dina(n10219), .dinb(n10216), .dout(n10220));
  jand g09965(.dina(n10220), .dinb(n10215), .dout(n10221));
  jxor g09966(.dina(n10221), .dinb(n3938), .dout(n10222));
  jxor g09967(.dina(n10222), .dinb(n10214), .dout(n10223));
  jxor g09968(.dina(n10223), .dinb(n10099), .dout(n10224));
  jor  g09969(.dina(n3751), .dinb(n2860), .dout(n10225));
  jor  g09970(.dina(n3574), .dinb(n2563), .dout(n10226));
  jor  g09971(.dina(n3754), .dinb(n2713), .dout(n10227));
  jor  g09972(.dina(n3749), .dinb(n2862), .dout(n10228));
  jand g09973(.dina(n10228), .dinb(n10227), .dout(n10229));
  jand g09974(.dina(n10229), .dinb(n10226), .dout(n10230));
  jand g09975(.dina(n10230), .dinb(n10225), .dout(n10231));
  jxor g09976(.dina(n10231), .dinb(n3410), .dout(n10232));
  jxor g09977(.dina(n10232), .dinb(n10224), .dout(n10233));
  jand g09978(.dina(n9942), .dinb(n9934), .dout(n10234));
  jand g09979(.dina(n9943), .dinb(n9811), .dout(n10235));
  jor  g09980(.dina(n10235), .dinb(n10234), .dout(n10236));
  jxor g09981(.dina(n10236), .dinb(n10233), .dout(n10237));
  jor  g09982(.dina(n3346), .dinb(n3239), .dout(n10238));
  jor  g09983(.dina(n3072), .dinb(n3023), .dout(n10239));
  jor  g09984(.dina(n3237), .dinb(n3348), .dout(n10240));
  jor  g09985(.dina(n3242), .dinb(n3186), .dout(n10241));
  jand g09986(.dina(n10241), .dinb(n10240), .dout(n10242));
  jand g09987(.dina(n10242), .dinb(n10239), .dout(n10243));
  jand g09988(.dina(n10243), .dinb(n10238), .dout(n10244));
  jxor g09989(.dina(n10244), .dinb(n2918), .dout(n10245));
  jxor g09990(.dina(n10245), .dinb(n10237), .dout(n10246));
  jxor g09991(.dina(n10246), .dinb(n10096), .dout(n10247));
  jor  g09992(.dina(n3871), .dinb(n2764), .dout(n10248));
  jor  g09993(.dina(n2609), .dinb(n3522), .dout(n10249));
  jor  g09994(.dina(n2761), .dinb(n3873), .dout(n10250));
  jor  g09995(.dina(n2766), .dinb(n3698), .dout(n10251));
  jand g09996(.dina(n10251), .dinb(n10250), .dout(n10252));
  jand g09997(.dina(n10252), .dinb(n10249), .dout(n10253));
  jand g09998(.dina(n10253), .dinb(n10248), .dout(n10254));
  jxor g09999(.dina(n10254), .dinb(n2468), .dout(n10255));
  jxor g10000(.dina(n10255), .dinb(n10247), .dout(n10256));
  jxor g10001(.dina(n10256), .dinb(n10093), .dout(n10257));
  jor  g10002(.dina(n4435), .dinb(n2324), .dout(n10258));
  jor  g10003(.dina(n2186), .dinb(n4060), .dout(n10259));
  jor  g10004(.dina(n2321), .dinb(n4249), .dout(n10260));
  jor  g10005(.dina(n2326), .dinb(n4437), .dout(n10261));
  jand g10006(.dina(n10261), .dinb(n10260), .dout(n10262));
  jand g10007(.dina(n10262), .dinb(n10259), .dout(n10263));
  jand g10008(.dina(n10263), .dinb(n10258), .dout(n10264));
  jxor g10009(.dina(n10264), .dinb(n2057), .dout(n10265));
  jxor g10010(.dina(n10265), .dinb(n10257), .dout(n10266));
  jxor g10011(.dina(n10266), .dinb(n10090), .dout(n10267));
  jor  g10012(.dina(n5038), .dinb(n1921), .dout(n10268));
  jor  g10013(.dina(n1806), .dinb(n4637), .dout(n10269));
  jor  g10014(.dina(n1923), .dinb(n5040), .dout(n10270));
  jor  g10015(.dina(n1918), .dinb(n4839), .dout(n10271));
  jand g10016(.dina(n10271), .dinb(n10270), .dout(n10272));
  jand g10017(.dina(n10272), .dinb(n10269), .dout(n10273));
  jand g10018(.dina(n10273), .dinb(n10268), .dout(n10274));
  jxor g10019(.dina(n10274), .dinb(n1687), .dout(n10275));
  jxor g10020(.dina(n10275), .dinb(n10267), .dout(n10276));
  jxor g10021(.dina(n10276), .dinb(n10087), .dout(n10277));
  jor  g10022(.dina(n5683), .dinb(n1569), .dout(n10278));
  jor  g10023(.dina(n1453), .dinb(n5253), .dout(n10279));
  jor  g10024(.dina(n1566), .dinb(n5469), .dout(n10280));
  jor  g10025(.dina(n1571), .dinb(n5685), .dout(n10281));
  jand g10026(.dina(n10281), .dinb(n10280), .dout(n10282));
  jand g10027(.dina(n10282), .dinb(n10279), .dout(n10283));
  jand g10028(.dina(n10283), .dinb(n10278), .dout(n10284));
  jxor g10029(.dina(n10284), .dinb(n1351), .dout(n10285));
  jxor g10030(.dina(n10285), .dinb(n10277), .dout(n10286));
  jxor g10031(.dina(n10286), .dinb(n10084), .dout(n10287));
  jor  g10032(.dina(n6364), .dinb(n1248), .dout(n10288));
  jor  g10033(.dina(n1147), .dinb(n5911), .dout(n10289));
  jor  g10034(.dina(n1246), .dinb(n6366), .dout(n10290));
  jor  g10035(.dina(n1251), .dinb(n6139), .dout(n10291));
  jand g10036(.dina(n10291), .dinb(n10290), .dout(n10292));
  jand g10037(.dina(n10292), .dinb(n10289), .dout(n10293));
  jand g10038(.dina(n10293), .dinb(n10288), .dout(n10294));
  jxor g10039(.dina(n10294), .dinb(n1061), .dout(n10295));
  jxor g10040(.dina(n10295), .dinb(n10287), .dout(n10296));
  jxor g10041(.dina(n10296), .dinb(n10081), .dout(n10297));
  jor  g10042(.dina(n7084), .dinb(n970), .dout(n10298));
  jor  g10043(.dina(n880), .dinb(n6605), .dout(n10299));
  jor  g10044(.dina(n967), .dinb(n6846), .dout(n10300));
  jor  g10045(.dina(n972), .dinb(n7086), .dout(n10301));
  jand g10046(.dina(n10301), .dinb(n10300), .dout(n10302));
  jand g10047(.dina(n10302), .dinb(n10299), .dout(n10303));
  jand g10048(.dina(n10303), .dinb(n10298), .dout(n10304));
  jxor g10049(.dina(n10304), .dinb(n810), .dout(n10305));
  jxor g10050(.dina(n10305), .dinb(n10297), .dout(n10306));
  jxor g10051(.dina(n10306), .dinb(n10078), .dout(n10307));
  jor  g10052(.dina(n7844), .dinb(n728), .dout(n10308));
  jor  g10053(.dina(n660), .dinb(n7338), .dout(n10309));
  jor  g10054(.dina(n731), .dinb(n7590), .dout(n10310));
  jor  g10055(.dina(n726), .dinb(n7846), .dout(n10311));
  jand g10056(.dina(n10311), .dinb(n10310), .dout(n10312));
  jand g10057(.dina(n10312), .dinb(n10309), .dout(n10313));
  jand g10058(.dina(n10313), .dinb(n10308), .dout(n10314));
  jxor g10059(.dina(n10314), .dinb(n606), .dout(n10315));
  jxor g10060(.dina(n10315), .dinb(n10307), .dout(n10316));
  jxor g10061(.dina(n10316), .dinb(n10075), .dout(n10317));
  jor  g10062(.dina(n8642), .dinb(n544), .dout(n10318));
  jor  g10063(.dina(n486), .dinb(n8111), .dout(n10319));
  jor  g10064(.dina(n542), .dinb(n8644), .dout(n10320));
  jor  g10065(.dina(n547), .dinb(n8378), .dout(n10321));
  jand g10066(.dina(n10321), .dinb(n10320), .dout(n10322));
  jand g10067(.dina(n10322), .dinb(n10319), .dout(n10323));
  jand g10068(.dina(n10323), .dinb(n10318), .dout(n10324));
  jxor g10069(.dina(n10324), .dinb(n446), .dout(n10325));
  jxor g10070(.dina(n10325), .dinb(n10317), .dout(n10326));
  jor  g10071(.dina(n9473), .dinb(n397), .dout(n10327));
  jor  g10072(.dina(n354), .dinb(n8920), .dout(n10328));
  jor  g10073(.dina(n399), .dinb(n9475), .dout(n10329));
  jor  g10074(.dina(n394), .dinb(n9195), .dout(n10330));
  jand g10075(.dina(n10330), .dinb(n10329), .dout(n10331));
  jand g10076(.dina(n10331), .dinb(n10328), .dout(n10332));
  jand g10077(.dina(n10332), .dinb(n10327), .dout(n10333));
  jxor g10078(.dina(n10333), .dinb(n364), .dout(n10334));
  jxor g10079(.dina(n10334), .dinb(n10326), .dout(n10335));
  jxor g10080(.dina(n10335), .dinb(n10072), .dout(n10336));
  jand g10081(.dina(b62 ), .dinb(b61 ), .dout(n10337));
  jnot g10082(.din(n10337), .dout(n10338));
  jnot g10083(.din(n10044), .dout(n10339));
  jnot g10084(.din(n9752), .dout(n10340));
  jnot g10085(.din(n9468), .dout(n10341));
  jnot g10086(.din(n9188), .dout(n10342));
  jnot g10087(.din(n8913), .dout(n10343));
  jnot g10088(.din(n8637), .dout(n10344));
  jnot g10089(.din(n8371), .dout(n10345));
  jnot g10090(.din(n8104), .dout(n10346));
  jnot g10091(.din(n7839), .dout(n10347));
  jnot g10092(.din(n7583), .dout(n10348));
  jnot g10093(.din(n7331), .dout(n10349));
  jnot g10094(.din(n7079), .dout(n10350));
  jnot g10095(.din(n6839), .dout(n10351));
  jnot g10096(.din(n6598), .dout(n10352));
  jnot g10097(.din(n6359), .dout(n10353));
  jnot g10098(.din(n6132), .dout(n10354));
  jnot g10099(.din(n5904), .dout(n10355));
  jnot g10100(.din(n5678), .dout(n10356));
  jnot g10101(.din(n5462), .dout(n10357));
  jnot g10102(.din(n5246), .dout(n10358));
  jnot g10103(.din(n5033), .dout(n10359));
  jnot g10104(.din(n4832), .dout(n10360));
  jnot g10105(.din(n4630), .dout(n10361));
  jnot g10106(.din(n4430), .dout(n10362));
  jnot g10107(.din(n4242), .dout(n10363));
  jnot g10108(.din(n4053), .dout(n10364));
  jnot g10109(.din(n3866), .dout(n10365));
  jnot g10110(.din(n3691), .dout(n10366));
  jnot g10111(.din(n3515), .dout(n10367));
  jnot g10112(.din(n3341), .dout(n10368));
  jnot g10113(.din(n3179), .dout(n10369));
  jnot g10114(.din(n3016), .dout(n10370));
  jnot g10115(.din(n2855), .dout(n10371));
  jnot g10116(.din(n2706), .dout(n10372));
  jnot g10117(.din(n2556), .dout(n10373));
  jnot g10118(.din(n2408), .dout(n10374));
  jnot g10119(.din(n2272), .dout(n10375));
  jnot g10120(.din(n2135), .dout(n10376));
  jnot g10121(.din(n2000), .dout(n10377));
  jnot g10122(.din(n1874), .dout(n10378));
  jnot g10123(.din(n1752), .dout(n10379));
  jnot g10124(.din(n1630), .dout(n10380));
  jnot g10125(.din(n1520), .dout(n10381));
  jnot g10126(.din(n1409), .dout(n10382));
  jnot g10127(.din(n1300), .dout(n10383));
  jnot g10128(.din(n1204), .dout(n10384));
  jnot g10129(.din(n1107), .dout(n10385));
  jnot g10130(.din(n1011), .dout(n10386));
  jnot g10131(.din(n927), .dout(n10387));
  jnot g10132(.din(n845), .dout(n10388));
  jnot g10133(.din(n765), .dout(n10389));
  jnot g10134(.din(n697), .dout(n10390));
  jnot g10135(.din(n630), .dout(n10391));
  jnot g10136(.din(n565), .dout(n10392));
  jnot g10137(.din(n512), .dout(n10393));
  jnot g10138(.din(n461), .dout(n10394));
  jnot g10139(.din(n407), .dout(n10395));
  jnot g10140(.din(n369), .dout(n10396));
  jnot g10141(.din(n332), .dout(n10397));
  jand g10142(.dina(n293), .dinb(n271), .dout(n10398));
  jor  g10143(.dina(n10398), .dinb(n305), .dout(n10399));
  jor  g10144(.dina(n10399), .dinb(n298), .dout(n10400));
  jand g10145(.dina(n10400), .dinb(n10397), .dout(n10401));
  jor  g10146(.dina(n336), .dinb(n10401), .dout(n10402));
  jand g10147(.dina(n10402), .dinb(n10396), .dout(n10403));
  jor  g10148(.dina(n373), .dinb(n10403), .dout(n10404));
  jand g10149(.dina(n10404), .dinb(n10395), .dout(n10405));
  jor  g10150(.dina(n411), .dinb(n10405), .dout(n10406));
  jand g10151(.dina(n10406), .dinb(n10394), .dout(n10407));
  jor  g10152(.dina(n465), .dinb(n10407), .dout(n10408));
  jand g10153(.dina(n10408), .dinb(n10393), .dout(n10409));
  jor  g10154(.dina(n516), .dinb(n10409), .dout(n10410));
  jand g10155(.dina(n10410), .dinb(n10392), .dout(n10411));
  jor  g10156(.dina(n569), .dinb(n10411), .dout(n10412));
  jand g10157(.dina(n10412), .dinb(n10391), .dout(n10413));
  jor  g10158(.dina(n634), .dinb(n10413), .dout(n10414));
  jand g10159(.dina(n10414), .dinb(n10390), .dout(n10415));
  jor  g10160(.dina(n701), .dinb(n10415), .dout(n10416));
  jand g10161(.dina(n10416), .dinb(n10389), .dout(n10417));
  jor  g10162(.dina(n769), .dinb(n10417), .dout(n10418));
  jand g10163(.dina(n10418), .dinb(n10388), .dout(n10419));
  jor  g10164(.dina(n849), .dinb(n10419), .dout(n10420));
  jand g10165(.dina(n10420), .dinb(n10387), .dout(n10421));
  jor  g10166(.dina(n931), .dinb(n10421), .dout(n10422));
  jand g10167(.dina(n10422), .dinb(n10386), .dout(n10423));
  jor  g10168(.dina(n1015), .dinb(n10423), .dout(n10424));
  jand g10169(.dina(n10424), .dinb(n10385), .dout(n10425));
  jor  g10170(.dina(n1111), .dinb(n10425), .dout(n10426));
  jand g10171(.dina(n10426), .dinb(n10384), .dout(n10427));
  jor  g10172(.dina(n1208), .dinb(n10427), .dout(n10428));
  jand g10173(.dina(n10428), .dinb(n10383), .dout(n10429));
  jor  g10174(.dina(n1304), .dinb(n10429), .dout(n10430));
  jand g10175(.dina(n10430), .dinb(n10382), .dout(n10431));
  jor  g10176(.dina(n1413), .dinb(n10431), .dout(n10432));
  jand g10177(.dina(n10432), .dinb(n10381), .dout(n10433));
  jor  g10178(.dina(n1524), .dinb(n10433), .dout(n10434));
  jand g10179(.dina(n10434), .dinb(n10380), .dout(n10435));
  jor  g10180(.dina(n1634), .dinb(n10435), .dout(n10436));
  jand g10181(.dina(n10436), .dinb(n10379), .dout(n10437));
  jor  g10182(.dina(n1756), .dinb(n10437), .dout(n10438));
  jand g10183(.dina(n10438), .dinb(n10378), .dout(n10439));
  jor  g10184(.dina(n1878), .dinb(n10439), .dout(n10440));
  jand g10185(.dina(n10440), .dinb(n10377), .dout(n10441));
  jor  g10186(.dina(n2004), .dinb(n10441), .dout(n10442));
  jand g10187(.dina(n10442), .dinb(n10376), .dout(n10443));
  jor  g10188(.dina(n2139), .dinb(n10443), .dout(n10444));
  jand g10189(.dina(n10444), .dinb(n10375), .dout(n10445));
  jor  g10190(.dina(n2276), .dinb(n10445), .dout(n10446));
  jand g10191(.dina(n10446), .dinb(n10374), .dout(n10447));
  jor  g10192(.dina(n2412), .dinb(n10447), .dout(n10448));
  jand g10193(.dina(n10448), .dinb(n10373), .dout(n10449));
  jor  g10194(.dina(n2560), .dinb(n10449), .dout(n10450));
  jand g10195(.dina(n10450), .dinb(n10372), .dout(n10451));
  jor  g10196(.dina(n2710), .dinb(n10451), .dout(n10452));
  jand g10197(.dina(n10452), .dinb(n10371), .dout(n10453));
  jor  g10198(.dina(n2859), .dinb(n10453), .dout(n10454));
  jand g10199(.dina(n10454), .dinb(n10370), .dout(n10455));
  jor  g10200(.dina(n3020), .dinb(n10455), .dout(n10456));
  jand g10201(.dina(n10456), .dinb(n10369), .dout(n10457));
  jor  g10202(.dina(n3183), .dinb(n10457), .dout(n10458));
  jand g10203(.dina(n10458), .dinb(n10368), .dout(n10459));
  jor  g10204(.dina(n3345), .dinb(n10459), .dout(n10460));
  jand g10205(.dina(n10460), .dinb(n10367), .dout(n10461));
  jor  g10206(.dina(n3519), .dinb(n10461), .dout(n10462));
  jand g10207(.dina(n10462), .dinb(n10366), .dout(n10463));
  jor  g10208(.dina(n3695), .dinb(n10463), .dout(n10464));
  jand g10209(.dina(n10464), .dinb(n10365), .dout(n10465));
  jor  g10210(.dina(n3870), .dinb(n10465), .dout(n10466));
  jand g10211(.dina(n10466), .dinb(n10364), .dout(n10467));
  jor  g10212(.dina(n4057), .dinb(n10467), .dout(n10468));
  jand g10213(.dina(n10468), .dinb(n10363), .dout(n10469));
  jor  g10214(.dina(n4246), .dinb(n10469), .dout(n10470));
  jand g10215(.dina(n10470), .dinb(n10362), .dout(n10471));
  jor  g10216(.dina(n4434), .dinb(n10471), .dout(n10472));
  jand g10217(.dina(n10472), .dinb(n10361), .dout(n10473));
  jor  g10218(.dina(n4634), .dinb(n10473), .dout(n10474));
  jand g10219(.dina(n10474), .dinb(n10360), .dout(n10475));
  jor  g10220(.dina(n4836), .dinb(n10475), .dout(n10476));
  jand g10221(.dina(n10476), .dinb(n10359), .dout(n10477));
  jor  g10222(.dina(n5037), .dinb(n10477), .dout(n10478));
  jand g10223(.dina(n10478), .dinb(n10358), .dout(n10479));
  jor  g10224(.dina(n5250), .dinb(n10479), .dout(n10480));
  jand g10225(.dina(n10480), .dinb(n10357), .dout(n10481));
  jor  g10226(.dina(n5466), .dinb(n10481), .dout(n10482));
  jand g10227(.dina(n10482), .dinb(n10356), .dout(n10483));
  jor  g10228(.dina(n5682), .dinb(n10483), .dout(n10484));
  jand g10229(.dina(n10484), .dinb(n10355), .dout(n10485));
  jor  g10230(.dina(n5908), .dinb(n10485), .dout(n10486));
  jand g10231(.dina(n10486), .dinb(n10354), .dout(n10487));
  jor  g10232(.dina(n6136), .dinb(n10487), .dout(n10488));
  jand g10233(.dina(n10488), .dinb(n10353), .dout(n10489));
  jor  g10234(.dina(n6363), .dinb(n10489), .dout(n10490));
  jand g10235(.dina(n10490), .dinb(n10352), .dout(n10491));
  jor  g10236(.dina(n6602), .dinb(n10491), .dout(n10492));
  jand g10237(.dina(n10492), .dinb(n10351), .dout(n10493));
  jor  g10238(.dina(n6843), .dinb(n10493), .dout(n10494));
  jand g10239(.dina(n10494), .dinb(n10350), .dout(n10495));
  jor  g10240(.dina(n7083), .dinb(n10495), .dout(n10496));
  jand g10241(.dina(n10496), .dinb(n10349), .dout(n10497));
  jor  g10242(.dina(n7335), .dinb(n10497), .dout(n10498));
  jand g10243(.dina(n10498), .dinb(n10348), .dout(n10499));
  jor  g10244(.dina(n7587), .dinb(n10499), .dout(n10500));
  jand g10245(.dina(n10500), .dinb(n10347), .dout(n10501));
  jor  g10246(.dina(n7843), .dinb(n10501), .dout(n10502));
  jand g10247(.dina(n10502), .dinb(n10346), .dout(n10503));
  jor  g10248(.dina(n8108), .dinb(n10503), .dout(n10504));
  jand g10249(.dina(n10504), .dinb(n10345), .dout(n10505));
  jor  g10250(.dina(n8375), .dinb(n10505), .dout(n10506));
  jand g10251(.dina(n10506), .dinb(n10344), .dout(n10507));
  jor  g10252(.dina(n8641), .dinb(n10507), .dout(n10508));
  jand g10253(.dina(n10508), .dinb(n10343), .dout(n10509));
  jor  g10254(.dina(n8917), .dinb(n10509), .dout(n10510));
  jand g10255(.dina(n10510), .dinb(n10342), .dout(n10511));
  jor  g10256(.dina(n9192), .dinb(n10511), .dout(n10512));
  jand g10257(.dina(n10512), .dinb(n10341), .dout(n10513));
  jor  g10258(.dina(n9472), .dinb(n10513), .dout(n10514));
  jand g10259(.dina(n10514), .dinb(n10340), .dout(n10515));
  jor  g10260(.dina(n9756), .dinb(n10515), .dout(n10516));
  jand g10261(.dina(n10516), .dinb(n10339), .dout(n10517));
  jor  g10262(.dina(n10048), .dinb(n10517), .dout(n10518));
  jand g10263(.dina(n10518), .dinb(n10338), .dout(n10519));
  jxor g10264(.dina(b63 ), .dinb(b62 ), .dout(n10520));
  jxor g10265(.dina(n10520), .dinb(n10519), .dout(n10521));
  jor  g10266(.dina(n10521), .dinb(n296), .dout(n10522));
  jnot g10267(.din(b63 ), .dout(n10523));
  jor  g10268(.dina(n264), .dinb(n10523), .dout(n10524));
  jor  g10269(.dina(n294), .dinb(n10051), .dout(n10525));
  jor  g10270(.dina(n280), .dinb(n9759), .dout(n10526));
  jand g10271(.dina(n10526), .dinb(n10525), .dout(n10527));
  jand g10272(.dina(n10527), .dinb(n10524), .dout(n10528));
  jand g10273(.dina(n10528), .dinb(n10522), .dout(n10529));
  jxor g10274(.dina(n10529), .dinb(n278), .dout(n10530));
  jxor g10275(.dina(n10530), .dinb(n10336), .dout(n10531));
  jxor g10276(.dina(n10531), .dinb(n10069), .dout(n10532));
  jxor g10277(.dina(n10532), .dinb(n10065), .dout(f63 ));
  jnot g10278(.din(n10336), .dout(n10534));
  jxor g10279(.dina(n10530), .dinb(n10534), .dout(n10535));
  jor  g10280(.dina(n10535), .dinb(n10069), .dout(n10536));
  jor  g10281(.dina(n10532), .dinb(n10065), .dout(n10537));
  jand g10282(.dina(n10537), .dinb(n10536), .dout(n10538));
  jand g10283(.dina(n10335), .dinb(n10072), .dout(n10539));
  jnot g10284(.din(n10539), .dout(n10540));
  jxor g10285(.dina(n10529), .dinb(a2 ), .dout(n10541));
  jor  g10286(.dina(n10541), .dinb(n10534), .dout(n10542));
  jand g10287(.dina(n10542), .dinb(n10540), .dout(n10543));
  jand g10288(.dina(n10325), .dinb(n10317), .dout(n10544));
  jand g10289(.dina(n10334), .dinb(n10326), .dout(n10545));
  jor  g10290(.dina(n10545), .dinb(n10544), .dout(n10546));
  jand g10291(.dina(n10315), .dinb(n10307), .dout(n10547));
  jand g10292(.dina(n10316), .dinb(n10075), .dout(n10548));
  jor  g10293(.dina(n10548), .dinb(n10547), .dout(n10549));
  jand g10294(.dina(n10305), .dinb(n10297), .dout(n10550));
  jand g10295(.dina(n10306), .dinb(n10078), .dout(n10551));
  jor  g10296(.dina(n10551), .dinb(n10550), .dout(n10552));
  jand g10297(.dina(n10295), .dinb(n10287), .dout(n10553));
  jand g10298(.dina(n10296), .dinb(n10081), .dout(n10554));
  jor  g10299(.dina(n10554), .dinb(n10553), .dout(n10555));
  jand g10300(.dina(n10285), .dinb(n10277), .dout(n10556));
  jand g10301(.dina(n10286), .dinb(n10084), .dout(n10557));
  jor  g10302(.dina(n10557), .dinb(n10556), .dout(n10558));
  jand g10303(.dina(n10275), .dinb(n10267), .dout(n10559));
  jand g10304(.dina(n10276), .dinb(n10087), .dout(n10560));
  jor  g10305(.dina(n10560), .dinb(n10559), .dout(n10561));
  jand g10306(.dina(n10265), .dinb(n10257), .dout(n10562));
  jand g10307(.dina(n10266), .dinb(n10090), .dout(n10563));
  jor  g10308(.dina(n10563), .dinb(n10562), .dout(n10564));
  jand g10309(.dina(n10255), .dinb(n10247), .dout(n10565));
  jand g10310(.dina(n10256), .dinb(n10093), .dout(n10566));
  jor  g10311(.dina(n10566), .dinb(n10565), .dout(n10567));
  jand g10312(.dina(n10245), .dinb(n10237), .dout(n10568));
  jand g10313(.dina(n10246), .dinb(n10096), .dout(n10569));
  jor  g10314(.dina(n10569), .dinb(n10568), .dout(n10570));
  jand g10315(.dina(n10222), .dinb(n10214), .dout(n10571));
  jand g10316(.dina(n10223), .dinb(n10099), .dout(n10572));
  jor  g10317(.dina(n10572), .dinb(n10571), .dout(n10573));
  jand g10318(.dina(n10212), .dinb(n10204), .dout(n10574));
  jand g10319(.dina(n10213), .dinb(n10102), .dout(n10575));
  jor  g10320(.dina(n10575), .dinb(n10574), .dout(n10576));
  jand g10321(.dina(n10202), .dinb(n10194), .dout(n10577));
  jand g10322(.dina(n10203), .dinb(n10105), .dout(n10578));
  jor  g10323(.dina(n10578), .dinb(n10577), .dout(n10579));
  jand g10324(.dina(n10182), .dinb(n10174), .dout(n10580));
  jand g10325(.dina(n10183), .dinb(n10111), .dout(n10581));
  jor  g10326(.dina(n10581), .dinb(n10580), .dout(n10582));
  jand g10327(.dina(n10162), .dinb(n10154), .dout(n10583));
  jand g10328(.dina(n10163), .dinb(n10117), .dout(n10584));
  jor  g10329(.dina(n10584), .dinb(n10583), .dout(n10585));
  jor  g10330(.dina(n10152), .dinb(n10144), .dout(n10586));
  jand g10331(.dina(n10153), .dinb(n10125), .dout(n10587));
  jnot g10332(.din(n10587), .dout(n10588));
  jand g10333(.dina(n10588), .dinb(n10586), .dout(n10589));
  jnot g10334(.din(n10589), .dout(n10590));
  jand g10335(.dina(n10130), .dinb(n10127), .dout(n10591));
  jand g10336(.dina(n10142), .dinb(n10131), .dout(n10592));
  jor  g10337(.dina(n10592), .dinb(n10591), .dout(n10593));
  jand g10338(.dina(a63 ), .dinb(a62 ), .dout(n10594));
  jand g10339(.dina(n10594), .dinb(b0 ), .dout(n10595));
  jand g10340(.dina(n10129), .dinb(b1 ), .dout(n10596));
  jor  g10341(.dina(n10596), .dinb(n10595), .dout(n10597));
  jnot g10342(.din(n10597), .dout(n10598));
  jor  g10343(.dina(n10134), .dinb(n337), .dout(n10599));
  jor  g10344(.dina(n10137), .dinb(n303), .dout(n10600));
  jor  g10345(.dina(n9849), .dinb(n293), .dout(n10601));
  jand g10346(.dina(n10601), .dinb(n10600), .dout(n10602));
  jor  g10347(.dina(n10132), .dinb(n340), .dout(n10603));
  jand g10348(.dina(n10603), .dinb(n10602), .dout(n10604));
  jand g10349(.dina(n10604), .dinb(n10599), .dout(n10605));
  jxor g10350(.dina(n10605), .dinb(a62 ), .dout(n10606));
  jxor g10351(.dina(n10606), .dinb(n10598), .dout(n10607));
  jxor g10352(.dina(n10607), .dinb(n10593), .dout(n10608));
  jnot g10353(.din(n10608), .dout(n10609));
  jor  g10354(.dina(n9271), .dinb(n466), .dout(n10610));
  jor  g10355(.dina(n9268), .dinb(n469), .dout(n10611));
  jor  g10356(.dina(n9003), .dinb(n377), .dout(n10612));
  jand g10357(.dina(n10612), .dinb(n10611), .dout(n10613));
  jor  g10358(.dina(n9273), .dinb(n415), .dout(n10614));
  jand g10359(.dina(n10614), .dinb(n10613), .dout(n10615));
  jand g10360(.dina(n10615), .dinb(n10610), .dout(n10616));
  jxor g10361(.dina(n10616), .dinb(a59 ), .dout(n10617));
  jxor g10362(.dina(n10617), .dinb(n10609), .dout(n10618));
  jxor g10363(.dina(n10618), .dinb(n10590), .dout(n10619));
  jor  g10364(.dina(n8457), .dinb(n635), .dout(n10620));
  jor  g10365(.dina(n8185), .dinb(n519), .dout(n10621));
  jor  g10366(.dina(n8459), .dinb(n572), .dout(n10622));
  jor  g10367(.dina(n8454), .dinb(n637), .dout(n10623));
  jand g10368(.dina(n10623), .dinb(n10622), .dout(n10624));
  jand g10369(.dina(n10624), .dinb(n10621), .dout(n10625));
  jand g10370(.dina(n10625), .dinb(n10620), .dout(n10626));
  jxor g10371(.dina(n10626), .dinb(n7929), .dout(n10627));
  jxor g10372(.dina(n10627), .dinb(n10619), .dout(n10628));
  jxor g10373(.dina(n10628), .dinb(n10585), .dout(n10629));
  jor  g10374(.dina(n7660), .dinb(n850), .dout(n10630));
  jor  g10375(.dina(n7415), .dinb(n704), .dout(n10631));
  jor  g10376(.dina(n7662), .dinb(n852), .dout(n10632));
  jor  g10377(.dina(n7657), .dinb(n772), .dout(n10633));
  jand g10378(.dina(n10633), .dinb(n10632), .dout(n10634));
  jand g10379(.dina(n10634), .dinb(n10631), .dout(n10635));
  jand g10380(.dina(n10635), .dinb(n10630), .dout(n10636));
  jxor g10381(.dina(n10636), .dinb(n7166), .dout(n10637));
  jxor g10382(.dina(n10637), .dinb(n10629), .dout(n10638));
  jand g10383(.dina(n10172), .dinb(n10164), .dout(n10639));
  jand g10384(.dina(n10173), .dinb(n10114), .dout(n10640));
  jor  g10385(.dina(n10640), .dinb(n10639), .dout(n10641));
  jxor g10386(.dina(n10641), .dinb(n10638), .dout(n10642));
  jor  g10387(.dina(n6914), .dinb(n1112), .dout(n10643));
  jor  g10388(.dina(n6673), .dinb(n934), .dout(n10644));
  jor  g10389(.dina(n6911), .dinb(n1018), .dout(n10645));
  jor  g10390(.dina(n6916), .dinb(n1114), .dout(n10646));
  jand g10391(.dina(n10646), .dinb(n10645), .dout(n10647));
  jand g10392(.dina(n10647), .dinb(n10644), .dout(n10648));
  jand g10393(.dina(n10648), .dinb(n10643), .dout(n10649));
  jxor g10394(.dina(n10649), .dinb(n6443), .dout(n10650));
  jxor g10395(.dina(n10650), .dinb(n10642), .dout(n10651));
  jxor g10396(.dina(n10651), .dinb(n10582), .dout(n10652));
  jor  g10397(.dina(n6207), .dinb(n1414), .dout(n10653));
  jor  g10398(.dina(n5975), .dinb(n1211), .dout(n10654));
  jor  g10399(.dina(n6210), .dinb(n1307), .dout(n10655));
  jor  g10400(.dina(n6205), .dinb(n1416), .dout(n10656));
  jand g10401(.dina(n10656), .dinb(n10655), .dout(n10657));
  jand g10402(.dina(n10657), .dinb(n10654), .dout(n10658));
  jand g10403(.dina(n10658), .dinb(n10653), .dout(n10659));
  jxor g10404(.dina(n10659), .dinb(n5759), .dout(n10660));
  jxor g10405(.dina(n10660), .dinb(n10652), .dout(n10661));
  jand g10406(.dina(n10192), .dinb(n10184), .dout(n10662));
  jand g10407(.dina(n10193), .dinb(n10108), .dout(n10663));
  jor  g10408(.dina(n10663), .dinb(n10662), .dout(n10664));
  jxor g10409(.dina(n10664), .dinb(n10661), .dout(n10665));
  jor  g10410(.dina(n5537), .dinb(n1757), .dout(n10666));
  jor  g10411(.dina(n5315), .dinb(n1527), .dout(n10667));
  jor  g10412(.dina(n5534), .dinb(n1637), .dout(n10668));
  jor  g10413(.dina(n5539), .dinb(n1759), .dout(n10669));
  jand g10414(.dina(n10669), .dinb(n10668), .dout(n10670));
  jand g10415(.dina(n10670), .dinb(n10667), .dout(n10671));
  jand g10416(.dina(n10671), .dinb(n10666), .dout(n10672));
  jxor g10417(.dina(n10672), .dinb(n5111), .dout(n10673));
  jxor g10418(.dina(n10673), .dinb(n10665), .dout(n10674));
  jxor g10419(.dina(n10674), .dinb(n10579), .dout(n10675));
  jor  g10420(.dina(n4902), .dinb(n2140), .dout(n10676));
  jor  g10421(.dina(n4696), .dinb(n1881), .dout(n10677));
  jor  g10422(.dina(n4899), .dinb(n2142), .dout(n10678));
  jor  g10423(.dina(n4904), .dinb(n2007), .dout(n10679));
  jand g10424(.dina(n10679), .dinb(n10678), .dout(n10680));
  jand g10425(.dina(n10680), .dinb(n10677), .dout(n10681));
  jand g10426(.dina(n10681), .dinb(n10676), .dout(n10682));
  jxor g10427(.dina(n10682), .dinb(n4505), .dout(n10683));
  jxor g10428(.dina(n10683), .dinb(n10675), .dout(n10684));
  jxor g10429(.dina(n10684), .dinb(n10576), .dout(n10685));
  jor  g10430(.dina(n4305), .dinb(n2561), .dout(n10686));
  jor  g10431(.dina(n4116), .dinb(n2279), .dout(n10687));
  jor  g10432(.dina(n4308), .dinb(n2415), .dout(n10688));
  jor  g10433(.dina(n4303), .dinb(n2563), .dout(n10689));
  jand g10434(.dina(n10689), .dinb(n10688), .dout(n10690));
  jand g10435(.dina(n10690), .dinb(n10687), .dout(n10691));
  jand g10436(.dina(n10691), .dinb(n10686), .dout(n10692));
  jxor g10437(.dina(n10692), .dinb(n3938), .dout(n10693));
  jxor g10438(.dina(n10693), .dinb(n10685), .dout(n10694));
  jxor g10439(.dina(n10694), .dinb(n10573), .dout(n10695));
  jor  g10440(.dina(n3751), .dinb(n3021), .dout(n10696));
  jor  g10441(.dina(n3574), .dinb(n2713), .dout(n10697));
  jor  g10442(.dina(n3754), .dinb(n2862), .dout(n10698));
  jor  g10443(.dina(n3749), .dinb(n3023), .dout(n10699));
  jand g10444(.dina(n10699), .dinb(n10698), .dout(n10700));
  jand g10445(.dina(n10700), .dinb(n10697), .dout(n10701));
  jand g10446(.dina(n10701), .dinb(n10696), .dout(n10702));
  jxor g10447(.dina(n10702), .dinb(n3410), .dout(n10703));
  jxor g10448(.dina(n10703), .dinb(n10695), .dout(n10704));
  jand g10449(.dina(n10232), .dinb(n10224), .dout(n10705));
  jand g10450(.dina(n10236), .dinb(n10233), .dout(n10706));
  jor  g10451(.dina(n10706), .dinb(n10705), .dout(n10707));
  jxor g10452(.dina(n10707), .dinb(n10704), .dout(n10708));
  jor  g10453(.dina(n3520), .dinb(n3239), .dout(n10709));
  jor  g10454(.dina(n3072), .dinb(n3186), .dout(n10710));
  jor  g10455(.dina(n3237), .dinb(n3522), .dout(n10711));
  jor  g10456(.dina(n3242), .dinb(n3348), .dout(n10712));
  jand g10457(.dina(n10712), .dinb(n10711), .dout(n10713));
  jand g10458(.dina(n10713), .dinb(n10710), .dout(n10714));
  jand g10459(.dina(n10714), .dinb(n10709), .dout(n10715));
  jxor g10460(.dina(n10715), .dinb(n2918), .dout(n10716));
  jxor g10461(.dina(n10716), .dinb(n10708), .dout(n10717));
  jxor g10462(.dina(n10717), .dinb(n10570), .dout(n10718));
  jor  g10463(.dina(n4058), .dinb(n2764), .dout(n10719));
  jor  g10464(.dina(n2609), .dinb(n3698), .dout(n10720));
  jor  g10465(.dina(n2761), .dinb(n4060), .dout(n10721));
  jor  g10466(.dina(n2766), .dinb(n3873), .dout(n10722));
  jand g10467(.dina(n10722), .dinb(n10721), .dout(n10723));
  jand g10468(.dina(n10723), .dinb(n10720), .dout(n10724));
  jand g10469(.dina(n10724), .dinb(n10719), .dout(n10725));
  jxor g10470(.dina(n10725), .dinb(n2468), .dout(n10726));
  jxor g10471(.dina(n10726), .dinb(n10718), .dout(n10727));
  jxor g10472(.dina(n10727), .dinb(n10567), .dout(n10728));
  jor  g10473(.dina(n4635), .dinb(n2324), .dout(n10729));
  jor  g10474(.dina(n2186), .dinb(n4249), .dout(n10730));
  jor  g10475(.dina(n2326), .dinb(n4637), .dout(n10731));
  jor  g10476(.dina(n2321), .dinb(n4437), .dout(n10732));
  jand g10477(.dina(n10732), .dinb(n10731), .dout(n10733));
  jand g10478(.dina(n10733), .dinb(n10730), .dout(n10734));
  jand g10479(.dina(n10734), .dinb(n10729), .dout(n10735));
  jxor g10480(.dina(n10735), .dinb(n2057), .dout(n10736));
  jxor g10481(.dina(n10736), .dinb(n10728), .dout(n10737));
  jxor g10482(.dina(n10737), .dinb(n10564), .dout(n10738));
  jor  g10483(.dina(n5251), .dinb(n1921), .dout(n10739));
  jor  g10484(.dina(n1806), .dinb(n4839), .dout(n10740));
  jor  g10485(.dina(n1918), .dinb(n5040), .dout(n10741));
  jor  g10486(.dina(n1923), .dinb(n5253), .dout(n10742));
  jand g10487(.dina(n10742), .dinb(n10741), .dout(n10743));
  jand g10488(.dina(n10743), .dinb(n10740), .dout(n10744));
  jand g10489(.dina(n10744), .dinb(n10739), .dout(n10745));
  jxor g10490(.dina(n10745), .dinb(n1687), .dout(n10746));
  jxor g10491(.dina(n10746), .dinb(n10738), .dout(n10747));
  jxor g10492(.dina(n10747), .dinb(n10561), .dout(n10748));
  jor  g10493(.dina(n5909), .dinb(n1569), .dout(n10749));
  jor  g10494(.dina(n1453), .dinb(n5469), .dout(n10750));
  jor  g10495(.dina(n1566), .dinb(n5685), .dout(n10751));
  jor  g10496(.dina(n1571), .dinb(n5911), .dout(n10752));
  jand g10497(.dina(n10752), .dinb(n10751), .dout(n10753));
  jand g10498(.dina(n10753), .dinb(n10750), .dout(n10754));
  jand g10499(.dina(n10754), .dinb(n10749), .dout(n10755));
  jxor g10500(.dina(n10755), .dinb(n1351), .dout(n10756));
  jxor g10501(.dina(n10756), .dinb(n10748), .dout(n10757));
  jxor g10502(.dina(n10757), .dinb(n10558), .dout(n10758));
  jor  g10503(.dina(n6603), .dinb(n1248), .dout(n10759));
  jor  g10504(.dina(n1147), .dinb(n6139), .dout(n10760));
  jor  g10505(.dina(n1251), .dinb(n6366), .dout(n10761));
  jor  g10506(.dina(n1246), .dinb(n6605), .dout(n10762));
  jand g10507(.dina(n10762), .dinb(n10761), .dout(n10763));
  jand g10508(.dina(n10763), .dinb(n10760), .dout(n10764));
  jand g10509(.dina(n10764), .dinb(n10759), .dout(n10765));
  jxor g10510(.dina(n10765), .dinb(n1061), .dout(n10766));
  jxor g10511(.dina(n10766), .dinb(n10758), .dout(n10767));
  jxor g10512(.dina(n10767), .dinb(n10555), .dout(n10768));
  jor  g10513(.dina(n7336), .dinb(n970), .dout(n10769));
  jor  g10514(.dina(n880), .dinb(n6846), .dout(n10770));
  jor  g10515(.dina(n972), .dinb(n7338), .dout(n10771));
  jor  g10516(.dina(n967), .dinb(n7086), .dout(n10772));
  jand g10517(.dina(n10772), .dinb(n10771), .dout(n10773));
  jand g10518(.dina(n10773), .dinb(n10770), .dout(n10774));
  jand g10519(.dina(n10774), .dinb(n10769), .dout(n10775));
  jxor g10520(.dina(n10775), .dinb(n810), .dout(n10776));
  jxor g10521(.dina(n10776), .dinb(n10768), .dout(n10777));
  jxor g10522(.dina(n10777), .dinb(n10552), .dout(n10778));
  jor  g10523(.dina(n8109), .dinb(n728), .dout(n10779));
  jor  g10524(.dina(n660), .dinb(n7590), .dout(n10780));
  jor  g10525(.dina(n731), .dinb(n7846), .dout(n10781));
  jor  g10526(.dina(n726), .dinb(n8111), .dout(n10782));
  jand g10527(.dina(n10782), .dinb(n10781), .dout(n10783));
  jand g10528(.dina(n10783), .dinb(n10780), .dout(n10784));
  jand g10529(.dina(n10784), .dinb(n10779), .dout(n10785));
  jxor g10530(.dina(n10785), .dinb(n606), .dout(n10786));
  jxor g10531(.dina(n10786), .dinb(n10778), .dout(n10787));
  jxor g10532(.dina(n10787), .dinb(n10549), .dout(n10788));
  jor  g10533(.dina(n8918), .dinb(n544), .dout(n10789));
  jor  g10534(.dina(n486), .dinb(n8378), .dout(n10790));
  jor  g10535(.dina(n547), .dinb(n8644), .dout(n10791));
  jor  g10536(.dina(n542), .dinb(n8920), .dout(n10792));
  jand g10537(.dina(n10792), .dinb(n10791), .dout(n10793));
  jand g10538(.dina(n10793), .dinb(n10790), .dout(n10794));
  jand g10539(.dina(n10794), .dinb(n10789), .dout(n10795));
  jxor g10540(.dina(n10795), .dinb(n446), .dout(n10796));
  jxor g10541(.dina(n10796), .dinb(n10788), .dout(n10797));
  jor  g10542(.dina(n9757), .dinb(n397), .dout(n10798));
  jor  g10543(.dina(n354), .dinb(n9195), .dout(n10799));
  jor  g10544(.dina(n394), .dinb(n9475), .dout(n10800));
  jor  g10545(.dina(n399), .dinb(n9759), .dout(n10801));
  jand g10546(.dina(n10801), .dinb(n10800), .dout(n10802));
  jand g10547(.dina(n10802), .dinb(n10799), .dout(n10803));
  jand g10548(.dina(n10803), .dinb(n10798), .dout(n10804));
  jxor g10549(.dina(n10804), .dinb(n364), .dout(n10805));
  jxor g10550(.dina(n10805), .dinb(n10797), .dout(n10806));
  jxor g10551(.dina(n10806), .dinb(n10546), .dout(n10807));
  jor  g10552(.dina(b63 ), .dinb(n10051), .dout(n10808));
  jor  g10553(.dina(n10808), .dinb(n10519), .dout(n10809));
  jand g10554(.dina(n10047), .dinb(n10046), .dout(n10810));
  jor  g10555(.dina(n10810), .dinb(b62 ), .dout(n10811));
  jor  g10556(.dina(n10811), .dinb(n10523), .dout(n10812));
  jand g10557(.dina(n10812), .dinb(n10809), .dout(n10813));
  jor  g10558(.dina(n10813), .dinb(n296), .dout(n10814));
  jor  g10559(.dina(n280), .dinb(n10051), .dout(n10815));
  jor  g10560(.dina(n294), .dinb(n10523), .dout(n10816));
  jand g10561(.dina(n10816), .dinb(n10815), .dout(n10817));
  jand g10562(.dina(n10817), .dinb(n10814), .dout(n10818));
  jxor g10563(.dina(n10818), .dinb(n278), .dout(n10819));
  jxor g10564(.dina(n10819), .dinb(n10807), .dout(n10820));
  jxor g10565(.dina(n10820), .dinb(n10543), .dout(n10821));
  jxor g10566(.dina(n10821), .dinb(n10538), .dout(f64 ));
  jand g10567(.dina(n10806), .dinb(n10546), .dout(n10823));
  jnot g10568(.din(n10823), .dout(n10824));
  jnot g10569(.din(n10807), .dout(n10825));
  jnot g10570(.din(n10819), .dout(n10826));
  jor  g10571(.dina(n10826), .dinb(n10825), .dout(n10827));
  jand g10572(.dina(n10827), .dinb(n10824), .dout(n10828));
  jand g10573(.dina(n10796), .dinb(n10788), .dout(n10829));
  jand g10574(.dina(n10805), .dinb(n10797), .dout(n10830));
  jor  g10575(.dina(n10830), .dinb(n10829), .dout(n10831));
  jand g10576(.dina(n10811), .dinb(b63 ), .dout(n10832));
  jand g10577(.dina(n10832), .dinb(n258), .dout(n10833));
  jnot g10578(.din(n10833), .dout(n10834));
  jor  g10579(.dina(n10834), .dinb(a2 ), .dout(n10835));
  jand g10580(.dina(n281), .dinb(b63 ), .dout(n10836));
  jor  g10581(.dina(n10836), .dinb(n278), .dout(n10837));
  jor  g10582(.dina(n10837), .dinb(n10833), .dout(n10838));
  jand g10583(.dina(n10838), .dinb(n10835), .dout(n10839));
  jxor g10584(.dina(n10839), .dinb(n10831), .dout(n10840));
  jand g10585(.dina(n10786), .dinb(n10778), .dout(n10841));
  jand g10586(.dina(n10787), .dinb(n10549), .dout(n10842));
  jor  g10587(.dina(n10842), .dinb(n10841), .dout(n10843));
  jand g10588(.dina(n10776), .dinb(n10768), .dout(n10844));
  jand g10589(.dina(n10777), .dinb(n10552), .dout(n10845));
  jor  g10590(.dina(n10845), .dinb(n10844), .dout(n10846));
  jand g10591(.dina(n10766), .dinb(n10758), .dout(n10847));
  jand g10592(.dina(n10767), .dinb(n10555), .dout(n10848));
  jor  g10593(.dina(n10848), .dinb(n10847), .dout(n10849));
  jand g10594(.dina(n10756), .dinb(n10748), .dout(n10850));
  jand g10595(.dina(n10757), .dinb(n10558), .dout(n10851));
  jor  g10596(.dina(n10851), .dinb(n10850), .dout(n10852));
  jand g10597(.dina(n10746), .dinb(n10738), .dout(n10853));
  jand g10598(.dina(n10747), .dinb(n10561), .dout(n10854));
  jor  g10599(.dina(n10854), .dinb(n10853), .dout(n10855));
  jand g10600(.dina(n10736), .dinb(n10728), .dout(n10856));
  jand g10601(.dina(n10737), .dinb(n10564), .dout(n10857));
  jor  g10602(.dina(n10857), .dinb(n10856), .dout(n10858));
  jand g10603(.dina(n10726), .dinb(n10718), .dout(n10859));
  jand g10604(.dina(n10727), .dinb(n10567), .dout(n10860));
  jor  g10605(.dina(n10860), .dinb(n10859), .dout(n10861));
  jand g10606(.dina(n10716), .dinb(n10708), .dout(n10862));
  jand g10607(.dina(n10717), .dinb(n10570), .dout(n10863));
  jor  g10608(.dina(n10863), .dinb(n10862), .dout(n10864));
  jand g10609(.dina(n10703), .dinb(n10695), .dout(n10865));
  jand g10610(.dina(n10707), .dinb(n10704), .dout(n10866));
  jor  g10611(.dina(n10866), .dinb(n10865), .dout(n10867));
  jand g10612(.dina(n10693), .dinb(n10685), .dout(n10868));
  jand g10613(.dina(n10694), .dinb(n10573), .dout(n10869));
  jor  g10614(.dina(n10869), .dinb(n10868), .dout(n10870));
  jand g10615(.dina(n10683), .dinb(n10675), .dout(n10871));
  jand g10616(.dina(n10684), .dinb(n10576), .dout(n10872));
  jor  g10617(.dina(n10872), .dinb(n10871), .dout(n10873));
  jand g10618(.dina(n10673), .dinb(n10665), .dout(n10874));
  jand g10619(.dina(n10674), .dinb(n10579), .dout(n10875));
  jor  g10620(.dina(n10875), .dinb(n10874), .dout(n10876));
  jand g10621(.dina(n10660), .dinb(n10652), .dout(n10877));
  jand g10622(.dina(n10664), .dinb(n10661), .dout(n10878));
  jor  g10623(.dina(n10878), .dinb(n10877), .dout(n10879));
  jand g10624(.dina(n10650), .dinb(n10642), .dout(n10880));
  jand g10625(.dina(n10651), .dinb(n10582), .dout(n10881));
  jor  g10626(.dina(n10881), .dinb(n10880), .dout(n10882));
  jand g10627(.dina(n10637), .dinb(n10629), .dout(n10883));
  jand g10628(.dina(n10641), .dinb(n10638), .dout(n10884));
  jor  g10629(.dina(n10884), .dinb(n10883), .dout(n10885));
  jand g10630(.dina(n10627), .dinb(n10619), .dout(n10886));
  jand g10631(.dina(n10628), .dinb(n10585), .dout(n10887));
  jor  g10632(.dina(n10887), .dinb(n10886), .dout(n10888));
  jor  g10633(.dina(n10617), .dinb(n10609), .dout(n10889));
  jand g10634(.dina(n10618), .dinb(n10590), .dout(n10890));
  jnot g10635(.din(n10890), .dout(n10891));
  jand g10636(.dina(n10891), .dinb(n10889), .dout(n10892));
  jnot g10637(.din(n10892), .dout(n10893));
  jor  g10638(.dina(n10606), .dinb(n10598), .dout(n10894));
  jand g10639(.dina(n10607), .dinb(n10593), .dout(n10895));
  jnot g10640(.din(n10895), .dout(n10896));
  jand g10641(.dina(n10896), .dinb(n10894), .dout(n10897));
  jnot g10642(.din(n10897), .dout(n10898));
  jand g10643(.dina(n10594), .dinb(b1 ), .dout(n10899));
  jand g10644(.dina(n10129), .dinb(b2 ), .dout(n10900));
  jor  g10645(.dina(n10900), .dinb(n10899), .dout(n10901));
  jnot g10646(.din(n10901), .dout(n10902));
  jor  g10647(.dina(n10134), .dinb(n374), .dout(n10903));
  jor  g10648(.dina(n10132), .dinb(n377), .dout(n10904));
  jor  g10649(.dina(n9849), .dinb(n303), .dout(n10905));
  jand g10650(.dina(n10905), .dinb(n10904), .dout(n10906));
  jor  g10651(.dina(n10137), .dinb(n340), .dout(n10907));
  jand g10652(.dina(n10907), .dinb(n10906), .dout(n10908));
  jand g10653(.dina(n10908), .dinb(n10903), .dout(n10909));
  jxor g10654(.dina(n10909), .dinb(a62 ), .dout(n10910));
  jxor g10655(.dina(n10910), .dinb(n10902), .dout(n10911));
  jxor g10656(.dina(n10911), .dinb(n10898), .dout(n10912));
  jor  g10657(.dina(n9271), .dinb(n517), .dout(n10913));
  jor  g10658(.dina(n9273), .dinb(n469), .dout(n10914));
  jor  g10659(.dina(n9268), .dinb(n519), .dout(n10915));
  jor  g10660(.dina(n9003), .dinb(n415), .dout(n10916));
  jand g10661(.dina(n10916), .dinb(n10915), .dout(n10917));
  jand g10662(.dina(n10917), .dinb(n10914), .dout(n10918));
  jand g10663(.dina(n10918), .dinb(n10913), .dout(n10919));
  jxor g10664(.dina(n10919), .dinb(n8729), .dout(n10920));
  jxor g10665(.dina(n10920), .dinb(n10912), .dout(n10921));
  jxor g10666(.dina(n10921), .dinb(n10893), .dout(n10922));
  jor  g10667(.dina(n8457), .dinb(n702), .dout(n10923));
  jor  g10668(.dina(n8185), .dinb(n572), .dout(n10924));
  jor  g10669(.dina(n8454), .dinb(n704), .dout(n10925));
  jor  g10670(.dina(n8459), .dinb(n637), .dout(n10926));
  jand g10671(.dina(n10926), .dinb(n10925), .dout(n10927));
  jand g10672(.dina(n10927), .dinb(n10924), .dout(n10928));
  jand g10673(.dina(n10928), .dinb(n10923), .dout(n10929));
  jxor g10674(.dina(n10929), .dinb(n7929), .dout(n10930));
  jxor g10675(.dina(n10930), .dinb(n10922), .dout(n10931));
  jxor g10676(.dina(n10931), .dinb(n10888), .dout(n10932));
  jor  g10677(.dina(n7660), .dinb(n932), .dout(n10933));
  jor  g10678(.dina(n7415), .dinb(n772), .dout(n10934));
  jor  g10679(.dina(n7662), .dinb(n934), .dout(n10935));
  jor  g10680(.dina(n7657), .dinb(n852), .dout(n10936));
  jand g10681(.dina(n10936), .dinb(n10935), .dout(n10937));
  jand g10682(.dina(n10937), .dinb(n10934), .dout(n10938));
  jand g10683(.dina(n10938), .dinb(n10933), .dout(n10939));
  jxor g10684(.dina(n10939), .dinb(n7166), .dout(n10940));
  jxor g10685(.dina(n10940), .dinb(n10932), .dout(n10941));
  jxor g10686(.dina(n10941), .dinb(n10885), .dout(n10942));
  jor  g10687(.dina(n6914), .dinb(n1209), .dout(n10943));
  jor  g10688(.dina(n6673), .dinb(n1018), .dout(n10944));
  jor  g10689(.dina(n6916), .dinb(n1211), .dout(n10945));
  jor  g10690(.dina(n6911), .dinb(n1114), .dout(n10946));
  jand g10691(.dina(n10946), .dinb(n10945), .dout(n10947));
  jand g10692(.dina(n10947), .dinb(n10944), .dout(n10948));
  jand g10693(.dina(n10948), .dinb(n10943), .dout(n10949));
  jxor g10694(.dina(n10949), .dinb(n6443), .dout(n10950));
  jxor g10695(.dina(n10950), .dinb(n10942), .dout(n10951));
  jxor g10696(.dina(n10951), .dinb(n10882), .dout(n10952));
  jor  g10697(.dina(n6207), .dinb(n1525), .dout(n10953));
  jor  g10698(.dina(n5975), .dinb(n1307), .dout(n10954));
  jor  g10699(.dina(n6210), .dinb(n1416), .dout(n10955));
  jor  g10700(.dina(n6205), .dinb(n1527), .dout(n10956));
  jand g10701(.dina(n10956), .dinb(n10955), .dout(n10957));
  jand g10702(.dina(n10957), .dinb(n10954), .dout(n10958));
  jand g10703(.dina(n10958), .dinb(n10953), .dout(n10959));
  jxor g10704(.dina(n10959), .dinb(n5759), .dout(n10960));
  jxor g10705(.dina(n10960), .dinb(n10952), .dout(n10961));
  jxor g10706(.dina(n10961), .dinb(n10879), .dout(n10962));
  jor  g10707(.dina(n5537), .dinb(n1879), .dout(n10963));
  jor  g10708(.dina(n5315), .dinb(n1637), .dout(n10964));
  jor  g10709(.dina(n5534), .dinb(n1759), .dout(n10965));
  jor  g10710(.dina(n5539), .dinb(n1881), .dout(n10966));
  jand g10711(.dina(n10966), .dinb(n10965), .dout(n10967));
  jand g10712(.dina(n10967), .dinb(n10964), .dout(n10968));
  jand g10713(.dina(n10968), .dinb(n10963), .dout(n10969));
  jxor g10714(.dina(n10969), .dinb(n5111), .dout(n10970));
  jxor g10715(.dina(n10970), .dinb(n10962), .dout(n10971));
  jxor g10716(.dina(n10971), .dinb(n10876), .dout(n10972));
  jor  g10717(.dina(n4902), .dinb(n2277), .dout(n10973));
  jor  g10718(.dina(n4696), .dinb(n2007), .dout(n10974));
  jor  g10719(.dina(n4904), .dinb(n2142), .dout(n10975));
  jor  g10720(.dina(n4899), .dinb(n2279), .dout(n10976));
  jand g10721(.dina(n10976), .dinb(n10975), .dout(n10977));
  jand g10722(.dina(n10977), .dinb(n10974), .dout(n10978));
  jand g10723(.dina(n10978), .dinb(n10973), .dout(n10979));
  jxor g10724(.dina(n10979), .dinb(n4505), .dout(n10980));
  jxor g10725(.dina(n10980), .dinb(n10972), .dout(n10981));
  jxor g10726(.dina(n10981), .dinb(n10873), .dout(n10982));
  jor  g10727(.dina(n4305), .dinb(n2711), .dout(n10983));
  jor  g10728(.dina(n4116), .dinb(n2415), .dout(n10984));
  jor  g10729(.dina(n4303), .dinb(n2713), .dout(n10985));
  jor  g10730(.dina(n4308), .dinb(n2563), .dout(n10986));
  jand g10731(.dina(n10986), .dinb(n10985), .dout(n10987));
  jand g10732(.dina(n10987), .dinb(n10984), .dout(n10988));
  jand g10733(.dina(n10988), .dinb(n10983), .dout(n10989));
  jxor g10734(.dina(n10989), .dinb(n3938), .dout(n10990));
  jxor g10735(.dina(n10990), .dinb(n10982), .dout(n10991));
  jxor g10736(.dina(n10991), .dinb(n10870), .dout(n10992));
  jor  g10737(.dina(n3751), .dinb(n3184), .dout(n10993));
  jor  g10738(.dina(n3574), .dinb(n2862), .dout(n10994));
  jor  g10739(.dina(n3754), .dinb(n3023), .dout(n10995));
  jor  g10740(.dina(n3749), .dinb(n3186), .dout(n10996));
  jand g10741(.dina(n10996), .dinb(n10995), .dout(n10997));
  jand g10742(.dina(n10997), .dinb(n10994), .dout(n10998));
  jand g10743(.dina(n10998), .dinb(n10993), .dout(n10999));
  jxor g10744(.dina(n10999), .dinb(n3410), .dout(n11000));
  jxor g10745(.dina(n11000), .dinb(n10992), .dout(n11001));
  jxor g10746(.dina(n11001), .dinb(n10867), .dout(n11002));
  jor  g10747(.dina(n3696), .dinb(n3239), .dout(n11003));
  jor  g10748(.dina(n3072), .dinb(n3348), .dout(n11004));
  jor  g10749(.dina(n3242), .dinb(n3522), .dout(n11005));
  jor  g10750(.dina(n3237), .dinb(n3698), .dout(n11006));
  jand g10751(.dina(n11006), .dinb(n11005), .dout(n11007));
  jand g10752(.dina(n11007), .dinb(n11004), .dout(n11008));
  jand g10753(.dina(n11008), .dinb(n11003), .dout(n11009));
  jxor g10754(.dina(n11009), .dinb(n2918), .dout(n11010));
  jxor g10755(.dina(n11010), .dinb(n11002), .dout(n11011));
  jxor g10756(.dina(n11011), .dinb(n10864), .dout(n11012));
  jor  g10757(.dina(n4247), .dinb(n2764), .dout(n11013));
  jor  g10758(.dina(n2609), .dinb(n3873), .dout(n11014));
  jor  g10759(.dina(n2761), .dinb(n4249), .dout(n11015));
  jor  g10760(.dina(n2766), .dinb(n4060), .dout(n11016));
  jand g10761(.dina(n11016), .dinb(n11015), .dout(n11017));
  jand g10762(.dina(n11017), .dinb(n11014), .dout(n11018));
  jand g10763(.dina(n11018), .dinb(n11013), .dout(n11019));
  jxor g10764(.dina(n11019), .dinb(n2468), .dout(n11020));
  jxor g10765(.dina(n11020), .dinb(n11012), .dout(n11021));
  jxor g10766(.dina(n11021), .dinb(n10861), .dout(n11022));
  jor  g10767(.dina(n4837), .dinb(n2324), .dout(n11023));
  jor  g10768(.dina(n2186), .dinb(n4437), .dout(n11024));
  jor  g10769(.dina(n2326), .dinb(n4839), .dout(n11025));
  jor  g10770(.dina(n2321), .dinb(n4637), .dout(n11026));
  jand g10771(.dina(n11026), .dinb(n11025), .dout(n11027));
  jand g10772(.dina(n11027), .dinb(n11024), .dout(n11028));
  jand g10773(.dina(n11028), .dinb(n11023), .dout(n11029));
  jxor g10774(.dina(n11029), .dinb(n2057), .dout(n11030));
  jxor g10775(.dina(n11030), .dinb(n11022), .dout(n11031));
  jxor g10776(.dina(n11031), .dinb(n10858), .dout(n11032));
  jor  g10777(.dina(n5467), .dinb(n1921), .dout(n11033));
  jor  g10778(.dina(n1806), .dinb(n5040), .dout(n11034));
  jor  g10779(.dina(n1923), .dinb(n5469), .dout(n11035));
  jor  g10780(.dina(n1918), .dinb(n5253), .dout(n11036));
  jand g10781(.dina(n11036), .dinb(n11035), .dout(n11037));
  jand g10782(.dina(n11037), .dinb(n11034), .dout(n11038));
  jand g10783(.dina(n11038), .dinb(n11033), .dout(n11039));
  jxor g10784(.dina(n11039), .dinb(n1687), .dout(n11040));
  jxor g10785(.dina(n11040), .dinb(n11032), .dout(n11041));
  jxor g10786(.dina(n11041), .dinb(n10855), .dout(n11042));
  jor  g10787(.dina(n6137), .dinb(n1569), .dout(n11043));
  jor  g10788(.dina(n1453), .dinb(n5685), .dout(n11044));
  jor  g10789(.dina(n1566), .dinb(n5911), .dout(n11045));
  jor  g10790(.dina(n1571), .dinb(n6139), .dout(n11046));
  jand g10791(.dina(n11046), .dinb(n11045), .dout(n11047));
  jand g10792(.dina(n11047), .dinb(n11044), .dout(n11048));
  jand g10793(.dina(n11048), .dinb(n11043), .dout(n11049));
  jxor g10794(.dina(n11049), .dinb(n1351), .dout(n11050));
  jxor g10795(.dina(n11050), .dinb(n11042), .dout(n11051));
  jxor g10796(.dina(n11051), .dinb(n10852), .dout(n11052));
  jor  g10797(.dina(n6844), .dinb(n1248), .dout(n11053));
  jor  g10798(.dina(n1147), .dinb(n6366), .dout(n11054));
  jor  g10799(.dina(n1246), .dinb(n6846), .dout(n11055));
  jor  g10800(.dina(n1251), .dinb(n6605), .dout(n11056));
  jand g10801(.dina(n11056), .dinb(n11055), .dout(n11057));
  jand g10802(.dina(n11057), .dinb(n11054), .dout(n11058));
  jand g10803(.dina(n11058), .dinb(n11053), .dout(n11059));
  jxor g10804(.dina(n11059), .dinb(n1061), .dout(n11060));
  jxor g10805(.dina(n11060), .dinb(n11052), .dout(n11061));
  jxor g10806(.dina(n11061), .dinb(n10849), .dout(n11062));
  jor  g10807(.dina(n7588), .dinb(n970), .dout(n11063));
  jor  g10808(.dina(n880), .dinb(n7086), .dout(n11064));
  jor  g10809(.dina(n972), .dinb(n7590), .dout(n11065));
  jor  g10810(.dina(n967), .dinb(n7338), .dout(n11066));
  jand g10811(.dina(n11066), .dinb(n11065), .dout(n11067));
  jand g10812(.dina(n11067), .dinb(n11064), .dout(n11068));
  jand g10813(.dina(n11068), .dinb(n11063), .dout(n11069));
  jxor g10814(.dina(n11069), .dinb(n810), .dout(n11070));
  jxor g10815(.dina(n11070), .dinb(n11062), .dout(n11071));
  jxor g10816(.dina(n11071), .dinb(n10846), .dout(n11072));
  jor  g10817(.dina(n8376), .dinb(n728), .dout(n11073));
  jor  g10818(.dina(n660), .dinb(n7846), .dout(n11074));
  jor  g10819(.dina(n731), .dinb(n8111), .dout(n11075));
  jor  g10820(.dina(n726), .dinb(n8378), .dout(n11076));
  jand g10821(.dina(n11076), .dinb(n11075), .dout(n11077));
  jand g10822(.dina(n11077), .dinb(n11074), .dout(n11078));
  jand g10823(.dina(n11078), .dinb(n11073), .dout(n11079));
  jxor g10824(.dina(n11079), .dinb(n606), .dout(n11080));
  jxor g10825(.dina(n11080), .dinb(n11072), .dout(n11081));
  jor  g10826(.dina(n9193), .dinb(n544), .dout(n11082));
  jor  g10827(.dina(n486), .dinb(n8644), .dout(n11083));
  jor  g10828(.dina(n547), .dinb(n8920), .dout(n11084));
  jor  g10829(.dina(n542), .dinb(n9195), .dout(n11085));
  jand g10830(.dina(n11085), .dinb(n11084), .dout(n11086));
  jand g10831(.dina(n11086), .dinb(n11083), .dout(n11087));
  jand g10832(.dina(n11087), .dinb(n11082), .dout(n11088));
  jxor g10833(.dina(n11088), .dinb(n446), .dout(n11089));
  jxor g10834(.dina(n11089), .dinb(n11081), .dout(n11090));
  jxor g10835(.dina(n11090), .dinb(n10843), .dout(n11091));
  jor  g10836(.dina(n10049), .dinb(n397), .dout(n11092));
  jor  g10837(.dina(n354), .dinb(n9475), .dout(n11093));
  jor  g10838(.dina(n394), .dinb(n9759), .dout(n11094));
  jor  g10839(.dina(n399), .dinb(n10051), .dout(n11095));
  jand g10840(.dina(n11095), .dinb(n11094), .dout(n11096));
  jand g10841(.dina(n11096), .dinb(n11093), .dout(n11097));
  jand g10842(.dina(n11097), .dinb(n11092), .dout(n11098));
  jxor g10843(.dina(n11098), .dinb(n364), .dout(n11099));
  jxor g10844(.dina(n11099), .dinb(n11091), .dout(n11100));
  jnot g10845(.din(n11100), .dout(n11101));
  jxor g10846(.dina(n11101), .dinb(n10840), .dout(n11102));
  jxor g10847(.dina(n11102), .dinb(n10828), .dout(n11103));
  jnot g10848(.din(n10820), .dout(n11104));
  jor  g10849(.dina(n11104), .dinb(n10543), .dout(n11105));
  jor  g10850(.dina(n10821), .dinb(n10538), .dout(n11106));
  jand g10851(.dina(n11106), .dinb(n11105), .dout(n11107));
  jxor g10852(.dina(n11107), .dinb(n11103), .dout(f65 ));
  jnot g10853(.din(n10831), .dout(n11109));
  jor  g10854(.dina(n10839), .dinb(n11109), .dout(n11110));
  jor  g10855(.dina(n11101), .dinb(n10840), .dout(n11111));
  jand g10856(.dina(n11111), .dinb(n11110), .dout(n11112));
  jand g10857(.dina(n11090), .dinb(n10843), .dout(n11113));
  jand g10858(.dina(n11099), .dinb(n11091), .dout(n11114));
  jor  g10859(.dina(n11114), .dinb(n11113), .dout(n11115));
  jor  g10860(.dina(n10521), .dinb(n397), .dout(n11116));
  jor  g10861(.dina(n354), .dinb(n9759), .dout(n11117));
  jor  g10862(.dina(n394), .dinb(n10051), .dout(n11118));
  jor  g10863(.dina(n399), .dinb(n10523), .dout(n11119));
  jand g10864(.dina(n11119), .dinb(n11118), .dout(n11120));
  jand g10865(.dina(n11120), .dinb(n11117), .dout(n11121));
  jand g10866(.dina(n11121), .dinb(n11116), .dout(n11122));
  jxor g10867(.dina(n11122), .dinb(n364), .dout(n11123));
  jxor g10868(.dina(n11123), .dinb(n11115), .dout(n11124));
  jand g10869(.dina(n11070), .dinb(n11062), .dout(n11125));
  jand g10870(.dina(n11071), .dinb(n10846), .dout(n11126));
  jor  g10871(.dina(n11126), .dinb(n11125), .dout(n11127));
  jor  g10872(.dina(n8642), .dinb(n728), .dout(n11128));
  jor  g10873(.dina(n660), .dinb(n8111), .dout(n11129));
  jor  g10874(.dina(n731), .dinb(n8378), .dout(n11130));
  jor  g10875(.dina(n726), .dinb(n8644), .dout(n11131));
  jand g10876(.dina(n11131), .dinb(n11130), .dout(n11132));
  jand g10877(.dina(n11132), .dinb(n11129), .dout(n11133));
  jand g10878(.dina(n11133), .dinb(n11128), .dout(n11134));
  jxor g10879(.dina(n11134), .dinb(n606), .dout(n11135));
  jxor g10880(.dina(n11135), .dinb(n11127), .dout(n11136));
  jand g10881(.dina(n11050), .dinb(n11042), .dout(n11137));
  jand g10882(.dina(n11051), .dinb(n10852), .dout(n11138));
  jor  g10883(.dina(n11138), .dinb(n11137), .dout(n11139));
  jor  g10884(.dina(n7084), .dinb(n1248), .dout(n11140));
  jor  g10885(.dina(n1147), .dinb(n6605), .dout(n11141));
  jor  g10886(.dina(n1246), .dinb(n7086), .dout(n11142));
  jor  g10887(.dina(n1251), .dinb(n6846), .dout(n11143));
  jand g10888(.dina(n11143), .dinb(n11142), .dout(n11144));
  jand g10889(.dina(n11144), .dinb(n11141), .dout(n11145));
  jand g10890(.dina(n11145), .dinb(n11140), .dout(n11146));
  jxor g10891(.dina(n11146), .dinb(n1061), .dout(n11147));
  jxor g10892(.dina(n11147), .dinb(n11139), .dout(n11148));
  jand g10893(.dina(n11040), .dinb(n11032), .dout(n11149));
  jand g10894(.dina(n11041), .dinb(n10855), .dout(n11150));
  jor  g10895(.dina(n11150), .dinb(n11149), .dout(n11151));
  jor  g10896(.dina(n6364), .dinb(n1569), .dout(n11152));
  jor  g10897(.dina(n1453), .dinb(n5911), .dout(n11153));
  jor  g10898(.dina(n1566), .dinb(n6139), .dout(n11154));
  jor  g10899(.dina(n1571), .dinb(n6366), .dout(n11155));
  jand g10900(.dina(n11155), .dinb(n11154), .dout(n11156));
  jand g10901(.dina(n11156), .dinb(n11153), .dout(n11157));
  jand g10902(.dina(n11157), .dinb(n11152), .dout(n11158));
  jxor g10903(.dina(n11158), .dinb(n1351), .dout(n11159));
  jxor g10904(.dina(n11159), .dinb(n11151), .dout(n11160));
  jand g10905(.dina(n11030), .dinb(n11022), .dout(n11161));
  jand g10906(.dina(n11031), .dinb(n10858), .dout(n11162));
  jor  g10907(.dina(n11162), .dinb(n11161), .dout(n11163));
  jor  g10908(.dina(n5683), .dinb(n1921), .dout(n11164));
  jor  g10909(.dina(n1806), .dinb(n5253), .dout(n11165));
  jor  g10910(.dina(n1918), .dinb(n5469), .dout(n11166));
  jor  g10911(.dina(n1923), .dinb(n5685), .dout(n11167));
  jand g10912(.dina(n11167), .dinb(n11166), .dout(n11168));
  jand g10913(.dina(n11168), .dinb(n11165), .dout(n11169));
  jand g10914(.dina(n11169), .dinb(n11164), .dout(n11170));
  jxor g10915(.dina(n11170), .dinb(n1687), .dout(n11171));
  jxor g10916(.dina(n11171), .dinb(n11163), .dout(n11172));
  jand g10917(.dina(n11020), .dinb(n11012), .dout(n11173));
  jand g10918(.dina(n11021), .dinb(n10861), .dout(n11174));
  jor  g10919(.dina(n11174), .dinb(n11173), .dout(n11175));
  jor  g10920(.dina(n5038), .dinb(n2324), .dout(n11176));
  jor  g10921(.dina(n2186), .dinb(n4637), .dout(n11177));
  jor  g10922(.dina(n2321), .dinb(n4839), .dout(n11178));
  jor  g10923(.dina(n2326), .dinb(n5040), .dout(n11179));
  jand g10924(.dina(n11179), .dinb(n11178), .dout(n11180));
  jand g10925(.dina(n11180), .dinb(n11177), .dout(n11181));
  jand g10926(.dina(n11181), .dinb(n11176), .dout(n11182));
  jxor g10927(.dina(n11182), .dinb(n2057), .dout(n11183));
  jxor g10928(.dina(n11183), .dinb(n11175), .dout(n11184));
  jand g10929(.dina(n11010), .dinb(n11002), .dout(n11185));
  jand g10930(.dina(n11011), .dinb(n10864), .dout(n11186));
  jor  g10931(.dina(n11186), .dinb(n11185), .dout(n11187));
  jor  g10932(.dina(n4435), .dinb(n2764), .dout(n11188));
  jor  g10933(.dina(n2609), .dinb(n4060), .dout(n11189));
  jor  g10934(.dina(n2761), .dinb(n4437), .dout(n11190));
  jor  g10935(.dina(n2766), .dinb(n4249), .dout(n11191));
  jand g10936(.dina(n11191), .dinb(n11190), .dout(n11192));
  jand g10937(.dina(n11192), .dinb(n11189), .dout(n11193));
  jand g10938(.dina(n11193), .dinb(n11188), .dout(n11194));
  jxor g10939(.dina(n11194), .dinb(n2468), .dout(n11195));
  jxor g10940(.dina(n11195), .dinb(n11187), .dout(n11196));
  jand g10941(.dina(n10980), .dinb(n10972), .dout(n11197));
  jand g10942(.dina(n10981), .dinb(n10873), .dout(n11198));
  jor  g10943(.dina(n11198), .dinb(n11197), .dout(n11199));
  jand g10944(.dina(n10970), .dinb(n10962), .dout(n11200));
  jand g10945(.dina(n10971), .dinb(n10876), .dout(n11201));
  jor  g10946(.dina(n11201), .dinb(n11200), .dout(n11202));
  jand g10947(.dina(n10950), .dinb(n10942), .dout(n11203));
  jand g10948(.dina(n10951), .dinb(n10882), .dout(n11204));
  jor  g10949(.dina(n11204), .dinb(n11203), .dout(n11205));
  jand g10950(.dina(n10940), .dinb(n10932), .dout(n11206));
  jand g10951(.dina(n10941), .dinb(n10885), .dout(n11207));
  jor  g10952(.dina(n11207), .dinb(n11206), .dout(n11208));
  jand g10953(.dina(n10930), .dinb(n10922), .dout(n11209));
  jand g10954(.dina(n10931), .dinb(n10888), .dout(n11210));
  jor  g10955(.dina(n11210), .dinb(n11209), .dout(n11211));
  jand g10956(.dina(n10920), .dinb(n10912), .dout(n11212));
  jand g10957(.dina(n10921), .dinb(n10893), .dout(n11213));
  jor  g10958(.dina(n11213), .dinb(n11212), .dout(n11214));
  jor  g10959(.dina(n10910), .dinb(n10902), .dout(n11215));
  jand g10960(.dina(n10911), .dinb(n10898), .dout(n11216));
  jnot g10961(.din(n11216), .dout(n11217));
  jand g10962(.dina(n11217), .dinb(n11215), .dout(n11218));
  jnot g10963(.din(n11218), .dout(n11219));
  jand g10964(.dina(n10594), .dinb(b2 ), .dout(n11220));
  jand g10965(.dina(n10129), .dinb(b3 ), .dout(n11221));
  jor  g10966(.dina(n11221), .dinb(n11220), .dout(n11222));
  jxor g10967(.dina(n11222), .dinb(a2 ), .dout(n11223));
  jnot g10968(.din(n11223), .dout(n11224));
  jor  g10969(.dina(n10134), .dinb(n412), .dout(n11225));
  jor  g10970(.dina(n10132), .dinb(n415), .dout(n11226));
  jor  g10971(.dina(n9849), .dinb(n340), .dout(n11227));
  jand g10972(.dina(n11227), .dinb(n11226), .dout(n11228));
  jor  g10973(.dina(n10137), .dinb(n377), .dout(n11229));
  jand g10974(.dina(n11229), .dinb(n11228), .dout(n11230));
  jand g10975(.dina(n11230), .dinb(n11225), .dout(n11231));
  jxor g10976(.dina(n11231), .dinb(a62 ), .dout(n11232));
  jxor g10977(.dina(n11232), .dinb(n11224), .dout(n11233));
  jxor g10978(.dina(n11233), .dinb(n11219), .dout(n11234));
  jor  g10979(.dina(n9271), .dinb(n570), .dout(n11235));
  jor  g10980(.dina(n9003), .dinb(n469), .dout(n11236));
  jor  g10981(.dina(n9273), .dinb(n519), .dout(n11237));
  jor  g10982(.dina(n9268), .dinb(n572), .dout(n11238));
  jand g10983(.dina(n11238), .dinb(n11237), .dout(n11239));
  jand g10984(.dina(n11239), .dinb(n11236), .dout(n11240));
  jand g10985(.dina(n11240), .dinb(n11235), .dout(n11241));
  jxor g10986(.dina(n11241), .dinb(n8729), .dout(n11242));
  jxor g10987(.dina(n11242), .dinb(n11234), .dout(n11243));
  jxor g10988(.dina(n11243), .dinb(n11214), .dout(n11244));
  jor  g10989(.dina(n8457), .dinb(n770), .dout(n11245));
  jor  g10990(.dina(n8185), .dinb(n637), .dout(n11246));
  jor  g10991(.dina(n8459), .dinb(n704), .dout(n11247));
  jor  g10992(.dina(n8454), .dinb(n772), .dout(n11248));
  jand g10993(.dina(n11248), .dinb(n11247), .dout(n11249));
  jand g10994(.dina(n11249), .dinb(n11246), .dout(n11250));
  jand g10995(.dina(n11250), .dinb(n11245), .dout(n11251));
  jxor g10996(.dina(n11251), .dinb(n7929), .dout(n11252));
  jxor g10997(.dina(n11252), .dinb(n11244), .dout(n11253));
  jxor g10998(.dina(n11253), .dinb(n11211), .dout(n11254));
  jor  g10999(.dina(n7660), .dinb(n1016), .dout(n11255));
  jor  g11000(.dina(n7415), .dinb(n852), .dout(n11256));
  jor  g11001(.dina(n7657), .dinb(n934), .dout(n11257));
  jor  g11002(.dina(n7662), .dinb(n1018), .dout(n11258));
  jand g11003(.dina(n11258), .dinb(n11257), .dout(n11259));
  jand g11004(.dina(n11259), .dinb(n11256), .dout(n11260));
  jand g11005(.dina(n11260), .dinb(n11255), .dout(n11261));
  jxor g11006(.dina(n11261), .dinb(n7166), .dout(n11262));
  jxor g11007(.dina(n11262), .dinb(n11254), .dout(n11263));
  jxor g11008(.dina(n11263), .dinb(n11208), .dout(n11264));
  jor  g11009(.dina(n6914), .dinb(n1305), .dout(n11265));
  jor  g11010(.dina(n6673), .dinb(n1114), .dout(n11266));
  jor  g11011(.dina(n6911), .dinb(n1211), .dout(n11267));
  jor  g11012(.dina(n6916), .dinb(n1307), .dout(n11268));
  jand g11013(.dina(n11268), .dinb(n11267), .dout(n11269));
  jand g11014(.dina(n11269), .dinb(n11266), .dout(n11270));
  jand g11015(.dina(n11270), .dinb(n11265), .dout(n11271));
  jxor g11016(.dina(n11271), .dinb(n6443), .dout(n11272));
  jxor g11017(.dina(n11272), .dinb(n11264), .dout(n11273));
  jxor g11018(.dina(n11273), .dinb(n11205), .dout(n11274));
  jor  g11019(.dina(n6207), .dinb(n1635), .dout(n11275));
  jor  g11020(.dina(n5975), .dinb(n1416), .dout(n11276));
  jor  g11021(.dina(n6210), .dinb(n1527), .dout(n11277));
  jor  g11022(.dina(n6205), .dinb(n1637), .dout(n11278));
  jand g11023(.dina(n11278), .dinb(n11277), .dout(n11279));
  jand g11024(.dina(n11279), .dinb(n11276), .dout(n11280));
  jand g11025(.dina(n11280), .dinb(n11275), .dout(n11281));
  jxor g11026(.dina(n11281), .dinb(n5759), .dout(n11282));
  jxor g11027(.dina(n11282), .dinb(n11274), .dout(n11283));
  jand g11028(.dina(n10960), .dinb(n10952), .dout(n11284));
  jand g11029(.dina(n10961), .dinb(n10879), .dout(n11285));
  jor  g11030(.dina(n11285), .dinb(n11284), .dout(n11286));
  jxor g11031(.dina(n11286), .dinb(n11283), .dout(n11287));
  jor  g11032(.dina(n5537), .dinb(n2005), .dout(n11288));
  jor  g11033(.dina(n5315), .dinb(n1759), .dout(n11289));
  jor  g11034(.dina(n5534), .dinb(n1881), .dout(n11290));
  jor  g11035(.dina(n5539), .dinb(n2007), .dout(n11291));
  jand g11036(.dina(n11291), .dinb(n11290), .dout(n11292));
  jand g11037(.dina(n11292), .dinb(n11289), .dout(n11293));
  jand g11038(.dina(n11293), .dinb(n11288), .dout(n11294));
  jxor g11039(.dina(n11294), .dinb(n5111), .dout(n11295));
  jxor g11040(.dina(n11295), .dinb(n11287), .dout(n11296));
  jxor g11041(.dina(n11296), .dinb(n11202), .dout(n11297));
  jor  g11042(.dina(n4902), .dinb(n2413), .dout(n11298));
  jor  g11043(.dina(n4696), .dinb(n2142), .dout(n11299));
  jor  g11044(.dina(n4899), .dinb(n2415), .dout(n11300));
  jor  g11045(.dina(n4904), .dinb(n2279), .dout(n11301));
  jand g11046(.dina(n11301), .dinb(n11300), .dout(n11302));
  jand g11047(.dina(n11302), .dinb(n11299), .dout(n11303));
  jand g11048(.dina(n11303), .dinb(n11298), .dout(n11304));
  jxor g11049(.dina(n11304), .dinb(n4505), .dout(n11305));
  jxor g11050(.dina(n11305), .dinb(n11297), .dout(n11306));
  jxor g11051(.dina(n11306), .dinb(n11199), .dout(n11307));
  jor  g11052(.dina(n4305), .dinb(n2860), .dout(n11308));
  jor  g11053(.dina(n4116), .dinb(n2563), .dout(n11309));
  jor  g11054(.dina(n4308), .dinb(n2713), .dout(n11310));
  jor  g11055(.dina(n4303), .dinb(n2862), .dout(n11311));
  jand g11056(.dina(n11311), .dinb(n11310), .dout(n11312));
  jand g11057(.dina(n11312), .dinb(n11309), .dout(n11313));
  jand g11058(.dina(n11313), .dinb(n11308), .dout(n11314));
  jxor g11059(.dina(n11314), .dinb(n3938), .dout(n11315));
  jxor g11060(.dina(n11315), .dinb(n11307), .dout(n11316));
  jand g11061(.dina(n10990), .dinb(n10982), .dout(n11317));
  jand g11062(.dina(n10991), .dinb(n10870), .dout(n11318));
  jor  g11063(.dina(n11318), .dinb(n11317), .dout(n11319));
  jxor g11064(.dina(n11319), .dinb(n11316), .dout(n11320));
  jor  g11065(.dina(n3751), .dinb(n3346), .dout(n11321));
  jor  g11066(.dina(n3574), .dinb(n3023), .dout(n11322));
  jor  g11067(.dina(n3754), .dinb(n3186), .dout(n11323));
  jor  g11068(.dina(n3749), .dinb(n3348), .dout(n11324));
  jand g11069(.dina(n11324), .dinb(n11323), .dout(n11325));
  jand g11070(.dina(n11325), .dinb(n11322), .dout(n11326));
  jand g11071(.dina(n11326), .dinb(n11321), .dout(n11327));
  jxor g11072(.dina(n11327), .dinb(n3410), .dout(n11328));
  jxor g11073(.dina(n11328), .dinb(n11320), .dout(n11329));
  jand g11074(.dina(n11000), .dinb(n10992), .dout(n11330));
  jand g11075(.dina(n11001), .dinb(n10867), .dout(n11331));
  jor  g11076(.dina(n11331), .dinb(n11330), .dout(n11332));
  jor  g11077(.dina(n3871), .dinb(n3239), .dout(n11333));
  jor  g11078(.dina(n3072), .dinb(n3522), .dout(n11334));
  jor  g11079(.dina(n3242), .dinb(n3698), .dout(n11335));
  jor  g11080(.dina(n3237), .dinb(n3873), .dout(n11336));
  jand g11081(.dina(n11336), .dinb(n11335), .dout(n11337));
  jand g11082(.dina(n11337), .dinb(n11334), .dout(n11338));
  jand g11083(.dina(n11338), .dinb(n11333), .dout(n11339));
  jxor g11084(.dina(n11339), .dinb(n2918), .dout(n11340));
  jxor g11085(.dina(n11340), .dinb(n11332), .dout(n11341));
  jxor g11086(.dina(n11341), .dinb(n11329), .dout(n11342));
  jxor g11087(.dina(n11342), .dinb(n11196), .dout(n11343));
  jxor g11088(.dina(n11343), .dinb(n11184), .dout(n11344));
  jxor g11089(.dina(n11344), .dinb(n11172), .dout(n11345));
  jxor g11090(.dina(n11345), .dinb(n11160), .dout(n11346));
  jxor g11091(.dina(n11346), .dinb(n11148), .dout(n11347));
  jand g11092(.dina(n11060), .dinb(n11052), .dout(n11348));
  jand g11093(.dina(n11061), .dinb(n10849), .dout(n11349));
  jor  g11094(.dina(n11349), .dinb(n11348), .dout(n11350));
  jor  g11095(.dina(n7844), .dinb(n970), .dout(n11351));
  jor  g11096(.dina(n880), .dinb(n7338), .dout(n11352));
  jor  g11097(.dina(n967), .dinb(n7590), .dout(n11353));
  jor  g11098(.dina(n972), .dinb(n7846), .dout(n11354));
  jand g11099(.dina(n11354), .dinb(n11353), .dout(n11355));
  jand g11100(.dina(n11355), .dinb(n11352), .dout(n11356));
  jand g11101(.dina(n11356), .dinb(n11351), .dout(n11357));
  jxor g11102(.dina(n11357), .dinb(n810), .dout(n11358));
  jxor g11103(.dina(n11358), .dinb(n11350), .dout(n11359));
  jxor g11104(.dina(n11359), .dinb(n11347), .dout(n11360));
  jxor g11105(.dina(n11360), .dinb(n11136), .dout(n11361));
  jand g11106(.dina(n11080), .dinb(n11072), .dout(n11362));
  jand g11107(.dina(n11089), .dinb(n11081), .dout(n11363));
  jor  g11108(.dina(n11363), .dinb(n11362), .dout(n11364));
  jor  g11109(.dina(n9473), .dinb(n544), .dout(n11365));
  jor  g11110(.dina(n486), .dinb(n8920), .dout(n11366));
  jor  g11111(.dina(n542), .dinb(n9475), .dout(n11367));
  jor  g11112(.dina(n547), .dinb(n9195), .dout(n11368));
  jand g11113(.dina(n11368), .dinb(n11367), .dout(n11369));
  jand g11114(.dina(n11369), .dinb(n11366), .dout(n11370));
  jand g11115(.dina(n11370), .dinb(n11365), .dout(n11371));
  jxor g11116(.dina(n11371), .dinb(n446), .dout(n11372));
  jxor g11117(.dina(n11372), .dinb(n11364), .dout(n11373));
  jxor g11118(.dina(n11373), .dinb(n11361), .dout(n11374));
  jxor g11119(.dina(n11374), .dinb(n11124), .dout(n11375));
  jxor g11120(.dina(n11375), .dinb(n11112), .dout(n11376));
  jnot g11121(.din(n11102), .dout(n11377));
  jor  g11122(.dina(n11377), .dinb(n10828), .dout(n11378));
  jor  g11123(.dina(n11107), .dinb(n11103), .dout(n11379));
  jand g11124(.dina(n11379), .dinb(n11378), .dout(n11380));
  jxor g11125(.dina(n11380), .dinb(n11376), .dout(f66 ));
  jnot g11126(.din(n11375), .dout(n11382));
  jor  g11127(.dina(n11382), .dinb(n11112), .dout(n11383));
  jor  g11128(.dina(n11380), .dinb(n11376), .dout(n11384));
  jand g11129(.dina(n11384), .dinb(n11383), .dout(n11385));
  jand g11130(.dina(n11123), .dinb(n11115), .dout(n11386));
  jand g11131(.dina(n11374), .dinb(n11124), .dout(n11387));
  jor  g11132(.dina(n11387), .dinb(n11386), .dout(n11388));
  jand g11133(.dina(n11147), .dinb(n11139), .dout(n11389));
  jand g11134(.dina(n11346), .dinb(n11148), .dout(n11390));
  jor  g11135(.dina(n11390), .dinb(n11389), .dout(n11391));
  jor  g11136(.dina(n8109), .dinb(n970), .dout(n11392));
  jor  g11137(.dina(n880), .dinb(n7590), .dout(n11393));
  jor  g11138(.dina(n967), .dinb(n7846), .dout(n11394));
  jor  g11139(.dina(n972), .dinb(n8111), .dout(n11395));
  jand g11140(.dina(n11395), .dinb(n11394), .dout(n11396));
  jand g11141(.dina(n11396), .dinb(n11393), .dout(n11397));
  jand g11142(.dina(n11397), .dinb(n11392), .dout(n11398));
  jxor g11143(.dina(n11398), .dinb(n810), .dout(n11399));
  jxor g11144(.dina(n11399), .dinb(n11391), .dout(n11400));
  jand g11145(.dina(n11171), .dinb(n11163), .dout(n11401));
  jand g11146(.dina(n11344), .dinb(n11172), .dout(n11402));
  jor  g11147(.dina(n11402), .dinb(n11401), .dout(n11403));
  jor  g11148(.dina(n6603), .dinb(n1569), .dout(n11404));
  jor  g11149(.dina(n1453), .dinb(n6139), .dout(n11405));
  jor  g11150(.dina(n1566), .dinb(n6366), .dout(n11406));
  jor  g11151(.dina(n1571), .dinb(n6605), .dout(n11407));
  jand g11152(.dina(n11407), .dinb(n11406), .dout(n11408));
  jand g11153(.dina(n11408), .dinb(n11405), .dout(n11409));
  jand g11154(.dina(n11409), .dinb(n11404), .dout(n11410));
  jxor g11155(.dina(n11410), .dinb(n1351), .dout(n11411));
  jxor g11156(.dina(n11411), .dinb(n11403), .dout(n11412));
  jand g11157(.dina(n11195), .dinb(n11187), .dout(n11413));
  jand g11158(.dina(n11342), .dinb(n11196), .dout(n11414));
  jor  g11159(.dina(n11414), .dinb(n11413), .dout(n11415));
  jor  g11160(.dina(n5251), .dinb(n2324), .dout(n11416));
  jor  g11161(.dina(n2186), .dinb(n4839), .dout(n11417));
  jor  g11162(.dina(n2321), .dinb(n5040), .dout(n11418));
  jor  g11163(.dina(n2326), .dinb(n5253), .dout(n11419));
  jand g11164(.dina(n11419), .dinb(n11418), .dout(n11420));
  jand g11165(.dina(n11420), .dinb(n11417), .dout(n11421));
  jand g11166(.dina(n11421), .dinb(n11416), .dout(n11422));
  jxor g11167(.dina(n11422), .dinb(n2057), .dout(n11423));
  jxor g11168(.dina(n11423), .dinb(n11415), .dout(n11424));
  jand g11169(.dina(n11319), .dinb(n11316), .dout(n11425));
  jand g11170(.dina(n11328), .dinb(n11320), .dout(n11426));
  jor  g11171(.dina(n11426), .dinb(n11425), .dout(n11427));
  jor  g11172(.dina(n4058), .dinb(n3239), .dout(n11428));
  jor  g11173(.dina(n3072), .dinb(n3698), .dout(n11429));
  jor  g11174(.dina(n3237), .dinb(n4060), .dout(n11430));
  jor  g11175(.dina(n3242), .dinb(n3873), .dout(n11431));
  jand g11176(.dina(n11431), .dinb(n11430), .dout(n11432));
  jand g11177(.dina(n11432), .dinb(n11429), .dout(n11433));
  jand g11178(.dina(n11433), .dinb(n11428), .dout(n11434));
  jxor g11179(.dina(n11434), .dinb(n2918), .dout(n11435));
  jxor g11180(.dina(n11435), .dinb(n11427), .dout(n11436));
  jand g11181(.dina(n11306), .dinb(n11199), .dout(n11437));
  jand g11182(.dina(n11315), .dinb(n11307), .dout(n11438));
  jor  g11183(.dina(n11438), .dinb(n11437), .dout(n11439));
  jand g11184(.dina(n11296), .dinb(n11202), .dout(n11440));
  jand g11185(.dina(n11305), .dinb(n11297), .dout(n11441));
  jor  g11186(.dina(n11441), .dinb(n11440), .dout(n11442));
  jand g11187(.dina(n11286), .dinb(n11283), .dout(n11443));
  jand g11188(.dina(n11295), .dinb(n11287), .dout(n11444));
  jor  g11189(.dina(n11444), .dinb(n11443), .dout(n11445));
  jand g11190(.dina(n11273), .dinb(n11205), .dout(n11446));
  jand g11191(.dina(n11282), .dinb(n11274), .dout(n11447));
  jor  g11192(.dina(n11447), .dinb(n11446), .dout(n11448));
  jand g11193(.dina(n11263), .dinb(n11208), .dout(n11449));
  jand g11194(.dina(n11272), .dinb(n11264), .dout(n11450));
  jor  g11195(.dina(n11450), .dinb(n11449), .dout(n11451));
  jand g11196(.dina(n11253), .dinb(n11211), .dout(n11452));
  jand g11197(.dina(n11262), .dinb(n11254), .dout(n11453));
  jor  g11198(.dina(n11453), .dinb(n11452), .dout(n11454));
  jand g11199(.dina(n11233), .dinb(n11219), .dout(n11455));
  jand g11200(.dina(n11242), .dinb(n11234), .dout(n11456));
  jor  g11201(.dina(n11456), .dinb(n11455), .dout(n11457));
  jand g11202(.dina(n11222), .dinb(a2 ), .dout(n11458));
  jnot g11203(.din(n11458), .dout(n11459));
  jor  g11204(.dina(n11232), .dinb(n11224), .dout(n11460));
  jand g11205(.dina(n11460), .dinb(n11459), .dout(n11461));
  jnot g11206(.din(n11461), .dout(n11462));
  jand g11207(.dina(n10594), .dinb(b3 ), .dout(n11463));
  jand g11208(.dina(n10129), .dinb(b4 ), .dout(n11464));
  jor  g11209(.dina(n11464), .dinb(n11463), .dout(n11465));
  jxor g11210(.dina(n11465), .dinb(a2 ), .dout(n11466));
  jnot g11211(.din(n11466), .dout(n11467));
  jor  g11212(.dina(n10134), .dinb(n466), .dout(n11468));
  jor  g11213(.dina(n10132), .dinb(n469), .dout(n11469));
  jor  g11214(.dina(n9849), .dinb(n377), .dout(n11470));
  jand g11215(.dina(n11470), .dinb(n11469), .dout(n11471));
  jor  g11216(.dina(n10137), .dinb(n415), .dout(n11472));
  jand g11217(.dina(n11472), .dinb(n11471), .dout(n11473));
  jand g11218(.dina(n11473), .dinb(n11468), .dout(n11474));
  jxor g11219(.dina(n11474), .dinb(a62 ), .dout(n11475));
  jxor g11220(.dina(n11475), .dinb(n11467), .dout(n11476));
  jxor g11221(.dina(n11476), .dinb(n11462), .dout(n11477));
  jor  g11222(.dina(n9271), .dinb(n635), .dout(n11478));
  jor  g11223(.dina(n9003), .dinb(n519), .dout(n11479));
  jor  g11224(.dina(n9268), .dinb(n637), .dout(n11480));
  jor  g11225(.dina(n9273), .dinb(n572), .dout(n11481));
  jand g11226(.dina(n11481), .dinb(n11480), .dout(n11482));
  jand g11227(.dina(n11482), .dinb(n11479), .dout(n11483));
  jand g11228(.dina(n11483), .dinb(n11478), .dout(n11484));
  jxor g11229(.dina(n11484), .dinb(n8729), .dout(n11485));
  jxor g11230(.dina(n11485), .dinb(n11477), .dout(n11486));
  jxor g11231(.dina(n11486), .dinb(n11457), .dout(n11487));
  jor  g11232(.dina(n8457), .dinb(n850), .dout(n11488));
  jor  g11233(.dina(n8185), .dinb(n704), .dout(n11489));
  jor  g11234(.dina(n8459), .dinb(n772), .dout(n11490));
  jor  g11235(.dina(n8454), .dinb(n852), .dout(n11491));
  jand g11236(.dina(n11491), .dinb(n11490), .dout(n11492));
  jand g11237(.dina(n11492), .dinb(n11489), .dout(n11493));
  jand g11238(.dina(n11493), .dinb(n11488), .dout(n11494));
  jxor g11239(.dina(n11494), .dinb(n7929), .dout(n11495));
  jxor g11240(.dina(n11495), .dinb(n11487), .dout(n11496));
  jand g11241(.dina(n11243), .dinb(n11214), .dout(n11497));
  jand g11242(.dina(n11252), .dinb(n11244), .dout(n11498));
  jor  g11243(.dina(n11498), .dinb(n11497), .dout(n11499));
  jxor g11244(.dina(n11499), .dinb(n11496), .dout(n11500));
  jor  g11245(.dina(n7660), .dinb(n1112), .dout(n11501));
  jor  g11246(.dina(n7415), .dinb(n934), .dout(n11502));
  jor  g11247(.dina(n7657), .dinb(n1018), .dout(n11503));
  jor  g11248(.dina(n7662), .dinb(n1114), .dout(n11504));
  jand g11249(.dina(n11504), .dinb(n11503), .dout(n11505));
  jand g11250(.dina(n11505), .dinb(n11502), .dout(n11506));
  jand g11251(.dina(n11506), .dinb(n11501), .dout(n11507));
  jxor g11252(.dina(n11507), .dinb(n7166), .dout(n11508));
  jxor g11253(.dina(n11508), .dinb(n11500), .dout(n11509));
  jxor g11254(.dina(n11509), .dinb(n11454), .dout(n11510));
  jor  g11255(.dina(n6914), .dinb(n1414), .dout(n11511));
  jor  g11256(.dina(n6673), .dinb(n1211), .dout(n11512));
  jor  g11257(.dina(n6916), .dinb(n1416), .dout(n11513));
  jor  g11258(.dina(n6911), .dinb(n1307), .dout(n11514));
  jand g11259(.dina(n11514), .dinb(n11513), .dout(n11515));
  jand g11260(.dina(n11515), .dinb(n11512), .dout(n11516));
  jand g11261(.dina(n11516), .dinb(n11511), .dout(n11517));
  jxor g11262(.dina(n11517), .dinb(n6443), .dout(n11518));
  jxor g11263(.dina(n11518), .dinb(n11510), .dout(n11519));
  jxor g11264(.dina(n11519), .dinb(n11451), .dout(n11520));
  jor  g11265(.dina(n6207), .dinb(n1757), .dout(n11521));
  jor  g11266(.dina(n5975), .dinb(n1527), .dout(n11522));
  jor  g11267(.dina(n6210), .dinb(n1637), .dout(n11523));
  jor  g11268(.dina(n6205), .dinb(n1759), .dout(n11524));
  jand g11269(.dina(n11524), .dinb(n11523), .dout(n11525));
  jand g11270(.dina(n11525), .dinb(n11522), .dout(n11526));
  jand g11271(.dina(n11526), .dinb(n11521), .dout(n11527));
  jxor g11272(.dina(n11527), .dinb(n5759), .dout(n11528));
  jxor g11273(.dina(n11528), .dinb(n11520), .dout(n11529));
  jxor g11274(.dina(n11529), .dinb(n11448), .dout(n11530));
  jor  g11275(.dina(n5537), .dinb(n2140), .dout(n11531));
  jor  g11276(.dina(n5315), .dinb(n1881), .dout(n11532));
  jor  g11277(.dina(n5539), .dinb(n2142), .dout(n11533));
  jor  g11278(.dina(n5534), .dinb(n2007), .dout(n11534));
  jand g11279(.dina(n11534), .dinb(n11533), .dout(n11535));
  jand g11280(.dina(n11535), .dinb(n11532), .dout(n11536));
  jand g11281(.dina(n11536), .dinb(n11531), .dout(n11537));
  jxor g11282(.dina(n11537), .dinb(n5111), .dout(n11538));
  jxor g11283(.dina(n11538), .dinb(n11530), .dout(n11539));
  jxor g11284(.dina(n11539), .dinb(n11445), .dout(n11540));
  jor  g11285(.dina(n4902), .dinb(n2561), .dout(n11541));
  jor  g11286(.dina(n4696), .dinb(n2279), .dout(n11542));
  jor  g11287(.dina(n4899), .dinb(n2563), .dout(n11543));
  jor  g11288(.dina(n4904), .dinb(n2415), .dout(n11544));
  jand g11289(.dina(n11544), .dinb(n11543), .dout(n11545));
  jand g11290(.dina(n11545), .dinb(n11542), .dout(n11546));
  jand g11291(.dina(n11546), .dinb(n11541), .dout(n11547));
  jxor g11292(.dina(n11547), .dinb(n4505), .dout(n11548));
  jxor g11293(.dina(n11548), .dinb(n11540), .dout(n11549));
  jxor g11294(.dina(n11549), .dinb(n11442), .dout(n11550));
  jor  g11295(.dina(n4305), .dinb(n3021), .dout(n11551));
  jor  g11296(.dina(n4116), .dinb(n2713), .dout(n11552));
  jor  g11297(.dina(n4308), .dinb(n2862), .dout(n11553));
  jor  g11298(.dina(n4303), .dinb(n3023), .dout(n11554));
  jand g11299(.dina(n11554), .dinb(n11553), .dout(n11555));
  jand g11300(.dina(n11555), .dinb(n11552), .dout(n11556));
  jand g11301(.dina(n11556), .dinb(n11551), .dout(n11557));
  jxor g11302(.dina(n11557), .dinb(n3938), .dout(n11558));
  jxor g11303(.dina(n11558), .dinb(n11550), .dout(n11559));
  jxor g11304(.dina(n11559), .dinb(n11439), .dout(n11560));
  jor  g11305(.dina(n3520), .dinb(n3751), .dout(n11561));
  jor  g11306(.dina(n3574), .dinb(n3186), .dout(n11562));
  jor  g11307(.dina(n3749), .dinb(n3522), .dout(n11563));
  jor  g11308(.dina(n3754), .dinb(n3348), .dout(n11564));
  jand g11309(.dina(n11564), .dinb(n11563), .dout(n11565));
  jand g11310(.dina(n11565), .dinb(n11562), .dout(n11566));
  jand g11311(.dina(n11566), .dinb(n11561), .dout(n11567));
  jxor g11312(.dina(n11567), .dinb(n3410), .dout(n11568));
  jxor g11313(.dina(n11568), .dinb(n11560), .dout(n11569));
  jxor g11314(.dina(n11569), .dinb(n11436), .dout(n11570));
  jand g11315(.dina(n11340), .dinb(n11332), .dout(n11571));
  jand g11316(.dina(n11341), .dinb(n11329), .dout(n11572));
  jor  g11317(.dina(n11572), .dinb(n11571), .dout(n11573));
  jor  g11318(.dina(n4635), .dinb(n2764), .dout(n11574));
  jor  g11319(.dina(n2609), .dinb(n4249), .dout(n11575));
  jor  g11320(.dina(n2761), .dinb(n4637), .dout(n11576));
  jor  g11321(.dina(n2766), .dinb(n4437), .dout(n11577));
  jand g11322(.dina(n11577), .dinb(n11576), .dout(n11578));
  jand g11323(.dina(n11578), .dinb(n11575), .dout(n11579));
  jand g11324(.dina(n11579), .dinb(n11574), .dout(n11580));
  jxor g11325(.dina(n11580), .dinb(n2468), .dout(n11581));
  jxor g11326(.dina(n11581), .dinb(n11573), .dout(n11582));
  jxor g11327(.dina(n11582), .dinb(n11570), .dout(n11583));
  jxor g11328(.dina(n11583), .dinb(n11424), .dout(n11584));
  jand g11329(.dina(n11183), .dinb(n11175), .dout(n11585));
  jand g11330(.dina(n11343), .dinb(n11184), .dout(n11586));
  jor  g11331(.dina(n11586), .dinb(n11585), .dout(n11587));
  jor  g11332(.dina(n5909), .dinb(n1921), .dout(n11588));
  jor  g11333(.dina(n1806), .dinb(n5469), .dout(n11589));
  jor  g11334(.dina(n1918), .dinb(n5685), .dout(n11590));
  jor  g11335(.dina(n1923), .dinb(n5911), .dout(n11591));
  jand g11336(.dina(n11591), .dinb(n11590), .dout(n11592));
  jand g11337(.dina(n11592), .dinb(n11589), .dout(n11593));
  jand g11338(.dina(n11593), .dinb(n11588), .dout(n11594));
  jxor g11339(.dina(n11594), .dinb(n1687), .dout(n11595));
  jxor g11340(.dina(n11595), .dinb(n11587), .dout(n11596));
  jxor g11341(.dina(n11596), .dinb(n11584), .dout(n11597));
  jxor g11342(.dina(n11597), .dinb(n11412), .dout(n11598));
  jand g11343(.dina(n11159), .dinb(n11151), .dout(n11599));
  jand g11344(.dina(n11345), .dinb(n11160), .dout(n11600));
  jor  g11345(.dina(n11600), .dinb(n11599), .dout(n11601));
  jor  g11346(.dina(n7336), .dinb(n1248), .dout(n11602));
  jor  g11347(.dina(n1147), .dinb(n6846), .dout(n11603));
  jor  g11348(.dina(n1246), .dinb(n7338), .dout(n11604));
  jor  g11349(.dina(n1251), .dinb(n7086), .dout(n11605));
  jand g11350(.dina(n11605), .dinb(n11604), .dout(n11606));
  jand g11351(.dina(n11606), .dinb(n11603), .dout(n11607));
  jand g11352(.dina(n11607), .dinb(n11602), .dout(n11608));
  jxor g11353(.dina(n11608), .dinb(n1061), .dout(n11609));
  jxor g11354(.dina(n11609), .dinb(n11601), .dout(n11610));
  jxor g11355(.dina(n11610), .dinb(n11598), .dout(n11611));
  jxor g11356(.dina(n11611), .dinb(n11400), .dout(n11612));
  jand g11357(.dina(n11358), .dinb(n11350), .dout(n11613));
  jand g11358(.dina(n11359), .dinb(n11347), .dout(n11614));
  jor  g11359(.dina(n11614), .dinb(n11613), .dout(n11615));
  jor  g11360(.dina(n8918), .dinb(n728), .dout(n11616));
  jor  g11361(.dina(n660), .dinb(n8378), .dout(n11617));
  jor  g11362(.dina(n726), .dinb(n8920), .dout(n11618));
  jor  g11363(.dina(n731), .dinb(n8644), .dout(n11619));
  jand g11364(.dina(n11619), .dinb(n11618), .dout(n11620));
  jand g11365(.dina(n11620), .dinb(n11617), .dout(n11621));
  jand g11366(.dina(n11621), .dinb(n11616), .dout(n11622));
  jxor g11367(.dina(n11622), .dinb(n606), .dout(n11623));
  jxor g11368(.dina(n11623), .dinb(n11615), .dout(n11624));
  jxor g11369(.dina(n11624), .dinb(n11612), .dout(n11625));
  jand g11370(.dina(n11135), .dinb(n11127), .dout(n11626));
  jand g11371(.dina(n11360), .dinb(n11136), .dout(n11627));
  jor  g11372(.dina(n11627), .dinb(n11626), .dout(n11628));
  jor  g11373(.dina(n9757), .dinb(n544), .dout(n11629));
  jor  g11374(.dina(n486), .dinb(n9195), .dout(n11630));
  jor  g11375(.dina(n547), .dinb(n9475), .dout(n11631));
  jor  g11376(.dina(n542), .dinb(n9759), .dout(n11632));
  jand g11377(.dina(n11632), .dinb(n11631), .dout(n11633));
  jand g11378(.dina(n11633), .dinb(n11630), .dout(n11634));
  jand g11379(.dina(n11634), .dinb(n11629), .dout(n11635));
  jxor g11380(.dina(n11635), .dinb(n446), .dout(n11636));
  jxor g11381(.dina(n11636), .dinb(n11628), .dout(n11637));
  jxor g11382(.dina(n11637), .dinb(n11625), .dout(n11638));
  jand g11383(.dina(n11372), .dinb(n11364), .dout(n11639));
  jand g11384(.dina(n11373), .dinb(n11361), .dout(n11640));
  jor  g11385(.dina(n11640), .dinb(n11639), .dout(n11641));
  jnot g11386(.din(n11641), .dout(n11642));
  jor  g11387(.dina(n10813), .dinb(n397), .dout(n11643));
  jor  g11388(.dina(n354), .dinb(n10051), .dout(n11644));
  jor  g11389(.dina(n394), .dinb(n10523), .dout(n11645));
  jand g11390(.dina(n11645), .dinb(n11644), .dout(n11646));
  jand g11391(.dina(n11646), .dinb(n11643), .dout(n11647));
  jxor g11392(.dina(n11647), .dinb(a5 ), .dout(n11648));
  jxor g11393(.dina(n11648), .dinb(n11642), .dout(n11649));
  jxor g11394(.dina(n11649), .dinb(n11638), .dout(n11650));
  jxor g11395(.dina(n11650), .dinb(n11388), .dout(n11651));
  jnot g11396(.din(n11651), .dout(n11652));
  jxor g11397(.dina(n11652), .dinb(n11385), .dout(f67 ));
  jand g11398(.dina(n11650), .dinb(n11388), .dout(n11654));
  jnot g11399(.din(n11654), .dout(n11655));
  jor  g11400(.dina(n11652), .dinb(n11385), .dout(n11656));
  jand g11401(.dina(n11656), .dinb(n11655), .dout(n11657));
  jor  g11402(.dina(n11648), .dinb(n11642), .dout(n11658));
  jand g11403(.dina(n11649), .dinb(n11638), .dout(n11659));
  jnot g11404(.din(n11659), .dout(n11660));
  jand g11405(.dina(n11660), .dinb(n11658), .dout(n11661));
  jnot g11406(.din(n11661), .dout(n11662));
  jand g11407(.dina(n11399), .dinb(n11391), .dout(n11663));
  jand g11408(.dina(n11611), .dinb(n11400), .dout(n11664));
  jor  g11409(.dina(n11664), .dinb(n11663), .dout(n11665));
  jor  g11410(.dina(n9193), .dinb(n728), .dout(n11666));
  jor  g11411(.dina(n660), .dinb(n8644), .dout(n11667));
  jor  g11412(.dina(n731), .dinb(n8920), .dout(n11668));
  jor  g11413(.dina(n726), .dinb(n9195), .dout(n11669));
  jand g11414(.dina(n11669), .dinb(n11668), .dout(n11670));
  jand g11415(.dina(n11670), .dinb(n11667), .dout(n11671));
  jand g11416(.dina(n11671), .dinb(n11666), .dout(n11672));
  jxor g11417(.dina(n11672), .dinb(n606), .dout(n11673));
  jxor g11418(.dina(n11673), .dinb(n11665), .dout(n11674));
  jand g11419(.dina(n11411), .dinb(n11403), .dout(n11675));
  jand g11420(.dina(n11597), .dinb(n11412), .dout(n11676));
  jor  g11421(.dina(n11676), .dinb(n11675), .dout(n11677));
  jor  g11422(.dina(n7588), .dinb(n1248), .dout(n11678));
  jor  g11423(.dina(n1147), .dinb(n7086), .dout(n11679));
  jor  g11424(.dina(n1251), .dinb(n7338), .dout(n11680));
  jor  g11425(.dina(n1246), .dinb(n7590), .dout(n11681));
  jand g11426(.dina(n11681), .dinb(n11680), .dout(n11682));
  jand g11427(.dina(n11682), .dinb(n11679), .dout(n11683));
  jand g11428(.dina(n11683), .dinb(n11678), .dout(n11684));
  jxor g11429(.dina(n11684), .dinb(n1061), .dout(n11685));
  jxor g11430(.dina(n11685), .dinb(n11677), .dout(n11686));
  jand g11431(.dina(n11423), .dinb(n11415), .dout(n11687));
  jand g11432(.dina(n11583), .dinb(n11424), .dout(n11688));
  jor  g11433(.dina(n11688), .dinb(n11687), .dout(n11689));
  jor  g11434(.dina(n6137), .dinb(n1921), .dout(n11690));
  jor  g11435(.dina(n1806), .dinb(n5685), .dout(n11691));
  jor  g11436(.dina(n1918), .dinb(n5911), .dout(n11692));
  jor  g11437(.dina(n1923), .dinb(n6139), .dout(n11693));
  jand g11438(.dina(n11693), .dinb(n11692), .dout(n11694));
  jand g11439(.dina(n11694), .dinb(n11691), .dout(n11695));
  jand g11440(.dina(n11695), .dinb(n11690), .dout(n11696));
  jxor g11441(.dina(n11696), .dinb(n1687), .dout(n11697));
  jxor g11442(.dina(n11697), .dinb(n11689), .dout(n11698));
  jand g11443(.dina(n11435), .dinb(n11427), .dout(n11699));
  jand g11444(.dina(n11569), .dinb(n11436), .dout(n11700));
  jor  g11445(.dina(n11700), .dinb(n11699), .dout(n11701));
  jor  g11446(.dina(n4837), .dinb(n2764), .dout(n11702));
  jor  g11447(.dina(n2609), .dinb(n4437), .dout(n11703));
  jor  g11448(.dina(n2761), .dinb(n4839), .dout(n11704));
  jor  g11449(.dina(n2766), .dinb(n4637), .dout(n11705));
  jand g11450(.dina(n11705), .dinb(n11704), .dout(n11706));
  jand g11451(.dina(n11706), .dinb(n11703), .dout(n11707));
  jand g11452(.dina(n11707), .dinb(n11702), .dout(n11708));
  jxor g11453(.dina(n11708), .dinb(n2468), .dout(n11709));
  jxor g11454(.dina(n11709), .dinb(n11701), .dout(n11710));
  jand g11455(.dina(n11559), .dinb(n11439), .dout(n11711));
  jand g11456(.dina(n11568), .dinb(n11560), .dout(n11712));
  jor  g11457(.dina(n11712), .dinb(n11711), .dout(n11713));
  jor  g11458(.dina(n4247), .dinb(n3239), .dout(n11714));
  jor  g11459(.dina(n3072), .dinb(n3873), .dout(n11715));
  jor  g11460(.dina(n3242), .dinb(n4060), .dout(n11716));
  jor  g11461(.dina(n3237), .dinb(n4249), .dout(n11717));
  jand g11462(.dina(n11717), .dinb(n11716), .dout(n11718));
  jand g11463(.dina(n11718), .dinb(n11715), .dout(n11719));
  jand g11464(.dina(n11719), .dinb(n11714), .dout(n11720));
  jxor g11465(.dina(n11720), .dinb(n2918), .dout(n11721));
  jxor g11466(.dina(n11721), .dinb(n11713), .dout(n11722));
  jand g11467(.dina(n11539), .dinb(n11445), .dout(n11723));
  jand g11468(.dina(n11548), .dinb(n11540), .dout(n11724));
  jor  g11469(.dina(n11724), .dinb(n11723), .dout(n11725));
  jand g11470(.dina(n11529), .dinb(n11448), .dout(n11726));
  jand g11471(.dina(n11538), .dinb(n11530), .dout(n11727));
  jor  g11472(.dina(n11727), .dinb(n11726), .dout(n11728));
  jand g11473(.dina(n11519), .dinb(n11451), .dout(n11729));
  jand g11474(.dina(n11528), .dinb(n11520), .dout(n11730));
  jor  g11475(.dina(n11730), .dinb(n11729), .dout(n11731));
  jand g11476(.dina(n11499), .dinb(n11496), .dout(n11732));
  jand g11477(.dina(n11508), .dinb(n11500), .dout(n11733));
  jor  g11478(.dina(n11733), .dinb(n11732), .dout(n11734));
  jand g11479(.dina(n11486), .dinb(n11457), .dout(n11735));
  jand g11480(.dina(n11495), .dinb(n11487), .dout(n11736));
  jor  g11481(.dina(n11736), .dinb(n11735), .dout(n11737));
  jand g11482(.dina(n11465), .dinb(a2 ), .dout(n11738));
  jnot g11483(.din(n11738), .dout(n11739));
  jor  g11484(.dina(n11475), .dinb(n11467), .dout(n11740));
  jand g11485(.dina(n11740), .dinb(n11739), .dout(n11741));
  jnot g11486(.din(n11741), .dout(n11742));
  jand g11487(.dina(n10594), .dinb(b4 ), .dout(n11743));
  jand g11488(.dina(n10129), .dinb(b5 ), .dout(n11744));
  jor  g11489(.dina(n11744), .dinb(n11743), .dout(n11745));
  jxor g11490(.dina(n11745), .dinb(a2 ), .dout(n11746));
  jor  g11491(.dina(n10134), .dinb(n517), .dout(n11747));
  jor  g11492(.dina(n10137), .dinb(n469), .dout(n11748));
  jor  g11493(.dina(n10132), .dinb(n519), .dout(n11749));
  jor  g11494(.dina(n9849), .dinb(n415), .dout(n11750));
  jand g11495(.dina(n11750), .dinb(n11749), .dout(n11751));
  jand g11496(.dina(n11751), .dinb(n11748), .dout(n11752));
  jand g11497(.dina(n11752), .dinb(n11747), .dout(n11753));
  jxor g11498(.dina(n11753), .dinb(n9559), .dout(n11754));
  jxor g11499(.dina(n11754), .dinb(n11746), .dout(n11755));
  jxor g11500(.dina(n11755), .dinb(n11742), .dout(n11756));
  jor  g11501(.dina(n9271), .dinb(n702), .dout(n11757));
  jor  g11502(.dina(n9003), .dinb(n572), .dout(n11758));
  jor  g11503(.dina(n9273), .dinb(n637), .dout(n11759));
  jor  g11504(.dina(n9268), .dinb(n704), .dout(n11760));
  jand g11505(.dina(n11760), .dinb(n11759), .dout(n11761));
  jand g11506(.dina(n11761), .dinb(n11758), .dout(n11762));
  jand g11507(.dina(n11762), .dinb(n11757), .dout(n11763));
  jxor g11508(.dina(n11763), .dinb(n8729), .dout(n11764));
  jxor g11509(.dina(n11764), .dinb(n11756), .dout(n11765));
  jand g11510(.dina(n11476), .dinb(n11462), .dout(n11766));
  jand g11511(.dina(n11485), .dinb(n11477), .dout(n11767));
  jor  g11512(.dina(n11767), .dinb(n11766), .dout(n11768));
  jxor g11513(.dina(n11768), .dinb(n11765), .dout(n11769));
  jor  g11514(.dina(n8457), .dinb(n932), .dout(n11770));
  jor  g11515(.dina(n8185), .dinb(n772), .dout(n11771));
  jor  g11516(.dina(n8459), .dinb(n852), .dout(n11772));
  jor  g11517(.dina(n8454), .dinb(n934), .dout(n11773));
  jand g11518(.dina(n11773), .dinb(n11772), .dout(n11774));
  jand g11519(.dina(n11774), .dinb(n11771), .dout(n11775));
  jand g11520(.dina(n11775), .dinb(n11770), .dout(n11776));
  jxor g11521(.dina(n11776), .dinb(n7929), .dout(n11777));
  jxor g11522(.dina(n11777), .dinb(n11769), .dout(n11778));
  jxor g11523(.dina(n11778), .dinb(n11737), .dout(n11779));
  jor  g11524(.dina(n7660), .dinb(n1209), .dout(n11780));
  jor  g11525(.dina(n7415), .dinb(n1018), .dout(n11781));
  jor  g11526(.dina(n7662), .dinb(n1211), .dout(n11782));
  jor  g11527(.dina(n7657), .dinb(n1114), .dout(n11783));
  jand g11528(.dina(n11783), .dinb(n11782), .dout(n11784));
  jand g11529(.dina(n11784), .dinb(n11781), .dout(n11785));
  jand g11530(.dina(n11785), .dinb(n11780), .dout(n11786));
  jxor g11531(.dina(n11786), .dinb(n7166), .dout(n11787));
  jxor g11532(.dina(n11787), .dinb(n11779), .dout(n11788));
  jxor g11533(.dina(n11788), .dinb(n11734), .dout(n11789));
  jor  g11534(.dina(n6914), .dinb(n1525), .dout(n11790));
  jor  g11535(.dina(n6673), .dinb(n1307), .dout(n11791));
  jor  g11536(.dina(n6916), .dinb(n1527), .dout(n11792));
  jor  g11537(.dina(n6911), .dinb(n1416), .dout(n11793));
  jand g11538(.dina(n11793), .dinb(n11792), .dout(n11794));
  jand g11539(.dina(n11794), .dinb(n11791), .dout(n11795));
  jand g11540(.dina(n11795), .dinb(n11790), .dout(n11796));
  jxor g11541(.dina(n11796), .dinb(n6443), .dout(n11797));
  jxor g11542(.dina(n11797), .dinb(n11789), .dout(n11798));
  jand g11543(.dina(n11509), .dinb(n11454), .dout(n11799));
  jand g11544(.dina(n11518), .dinb(n11510), .dout(n11800));
  jor  g11545(.dina(n11800), .dinb(n11799), .dout(n11801));
  jxor g11546(.dina(n11801), .dinb(n11798), .dout(n11802));
  jor  g11547(.dina(n6207), .dinb(n1879), .dout(n11803));
  jor  g11548(.dina(n5975), .dinb(n1637), .dout(n11804));
  jor  g11549(.dina(n6205), .dinb(n1881), .dout(n11805));
  jor  g11550(.dina(n6210), .dinb(n1759), .dout(n11806));
  jand g11551(.dina(n11806), .dinb(n11805), .dout(n11807));
  jand g11552(.dina(n11807), .dinb(n11804), .dout(n11808));
  jand g11553(.dina(n11808), .dinb(n11803), .dout(n11809));
  jxor g11554(.dina(n11809), .dinb(n5759), .dout(n11810));
  jxor g11555(.dina(n11810), .dinb(n11802), .dout(n11811));
  jxor g11556(.dina(n11811), .dinb(n11731), .dout(n11812));
  jor  g11557(.dina(n5537), .dinb(n2277), .dout(n11813));
  jor  g11558(.dina(n5315), .dinb(n2007), .dout(n11814));
  jor  g11559(.dina(n5539), .dinb(n2279), .dout(n11815));
  jor  g11560(.dina(n5534), .dinb(n2142), .dout(n11816));
  jand g11561(.dina(n11816), .dinb(n11815), .dout(n11817));
  jand g11562(.dina(n11817), .dinb(n11814), .dout(n11818));
  jand g11563(.dina(n11818), .dinb(n11813), .dout(n11819));
  jxor g11564(.dina(n11819), .dinb(n5111), .dout(n11820));
  jxor g11565(.dina(n11820), .dinb(n11812), .dout(n11821));
  jxor g11566(.dina(n11821), .dinb(n11728), .dout(n11822));
  jor  g11567(.dina(n4902), .dinb(n2711), .dout(n11823));
  jor  g11568(.dina(n4696), .dinb(n2415), .dout(n11824));
  jor  g11569(.dina(n4899), .dinb(n2713), .dout(n11825));
  jor  g11570(.dina(n4904), .dinb(n2563), .dout(n11826));
  jand g11571(.dina(n11826), .dinb(n11825), .dout(n11827));
  jand g11572(.dina(n11827), .dinb(n11824), .dout(n11828));
  jand g11573(.dina(n11828), .dinb(n11823), .dout(n11829));
  jxor g11574(.dina(n11829), .dinb(n4505), .dout(n11830));
  jxor g11575(.dina(n11830), .dinb(n11822), .dout(n11831));
  jxor g11576(.dina(n11831), .dinb(n11725), .dout(n11832));
  jor  g11577(.dina(n4305), .dinb(n3184), .dout(n11833));
  jor  g11578(.dina(n4116), .dinb(n2862), .dout(n11834));
  jor  g11579(.dina(n4308), .dinb(n3023), .dout(n11835));
  jor  g11580(.dina(n4303), .dinb(n3186), .dout(n11836));
  jand g11581(.dina(n11836), .dinb(n11835), .dout(n11837));
  jand g11582(.dina(n11837), .dinb(n11834), .dout(n11838));
  jand g11583(.dina(n11838), .dinb(n11833), .dout(n11839));
  jxor g11584(.dina(n11839), .dinb(n3938), .dout(n11840));
  jxor g11585(.dina(n11840), .dinb(n11832), .dout(n11841));
  jand g11586(.dina(n11549), .dinb(n11442), .dout(n11842));
  jand g11587(.dina(n11558), .dinb(n11550), .dout(n11843));
  jor  g11588(.dina(n11843), .dinb(n11842), .dout(n11844));
  jxor g11589(.dina(n11844), .dinb(n11841), .dout(n11845));
  jor  g11590(.dina(n3696), .dinb(n3751), .dout(n11846));
  jor  g11591(.dina(n3574), .dinb(n3348), .dout(n11847));
  jor  g11592(.dina(n3754), .dinb(n3522), .dout(n11848));
  jor  g11593(.dina(n3749), .dinb(n3698), .dout(n11849));
  jand g11594(.dina(n11849), .dinb(n11848), .dout(n11850));
  jand g11595(.dina(n11850), .dinb(n11847), .dout(n11851));
  jand g11596(.dina(n11851), .dinb(n11846), .dout(n11852));
  jxor g11597(.dina(n11852), .dinb(n3410), .dout(n11853));
  jxor g11598(.dina(n11853), .dinb(n11845), .dout(n11854));
  jxor g11599(.dina(n11854), .dinb(n11722), .dout(n11855));
  jxor g11600(.dina(n11855), .dinb(n11710), .dout(n11856));
  jand g11601(.dina(n11581), .dinb(n11573), .dout(n11857));
  jand g11602(.dina(n11582), .dinb(n11570), .dout(n11858));
  jor  g11603(.dina(n11858), .dinb(n11857), .dout(n11859));
  jor  g11604(.dina(n5467), .dinb(n2324), .dout(n11860));
  jor  g11605(.dina(n2186), .dinb(n5040), .dout(n11861));
  jor  g11606(.dina(n2321), .dinb(n5253), .dout(n11862));
  jor  g11607(.dina(n2326), .dinb(n5469), .dout(n11863));
  jand g11608(.dina(n11863), .dinb(n11862), .dout(n11864));
  jand g11609(.dina(n11864), .dinb(n11861), .dout(n11865));
  jand g11610(.dina(n11865), .dinb(n11860), .dout(n11866));
  jxor g11611(.dina(n11866), .dinb(n2057), .dout(n11867));
  jxor g11612(.dina(n11867), .dinb(n11859), .dout(n11868));
  jxor g11613(.dina(n11868), .dinb(n11856), .dout(n11869));
  jxor g11614(.dina(n11869), .dinb(n11698), .dout(n11870));
  jand g11615(.dina(n11595), .dinb(n11587), .dout(n11871));
  jand g11616(.dina(n11596), .dinb(n11584), .dout(n11872));
  jor  g11617(.dina(n11872), .dinb(n11871), .dout(n11873));
  jor  g11618(.dina(n6844), .dinb(n1569), .dout(n11874));
  jor  g11619(.dina(n1453), .dinb(n6366), .dout(n11875));
  jor  g11620(.dina(n1566), .dinb(n6605), .dout(n11876));
  jor  g11621(.dina(n1571), .dinb(n6846), .dout(n11877));
  jand g11622(.dina(n11877), .dinb(n11876), .dout(n11878));
  jand g11623(.dina(n11878), .dinb(n11875), .dout(n11879));
  jand g11624(.dina(n11879), .dinb(n11874), .dout(n11880));
  jxor g11625(.dina(n11880), .dinb(n1351), .dout(n11881));
  jxor g11626(.dina(n11881), .dinb(n11873), .dout(n11882));
  jxor g11627(.dina(n11882), .dinb(n11870), .dout(n11883));
  jxor g11628(.dina(n11883), .dinb(n11686), .dout(n11884));
  jand g11629(.dina(n11609), .dinb(n11601), .dout(n11885));
  jand g11630(.dina(n11610), .dinb(n11598), .dout(n11886));
  jor  g11631(.dina(n11886), .dinb(n11885), .dout(n11887));
  jor  g11632(.dina(n8376), .dinb(n970), .dout(n11888));
  jor  g11633(.dina(n880), .dinb(n7846), .dout(n11889));
  jor  g11634(.dina(n972), .dinb(n8378), .dout(n11890));
  jor  g11635(.dina(n967), .dinb(n8111), .dout(n11891));
  jand g11636(.dina(n11891), .dinb(n11890), .dout(n11892));
  jand g11637(.dina(n11892), .dinb(n11889), .dout(n11893));
  jand g11638(.dina(n11893), .dinb(n11888), .dout(n11894));
  jxor g11639(.dina(n11894), .dinb(n810), .dout(n11895));
  jxor g11640(.dina(n11895), .dinb(n11887), .dout(n11896));
  jxor g11641(.dina(n11896), .dinb(n11884), .dout(n11897));
  jxor g11642(.dina(n11897), .dinb(n11674), .dout(n11898));
  jand g11643(.dina(n11623), .dinb(n11615), .dout(n11899));
  jand g11644(.dina(n11624), .dinb(n11612), .dout(n11900));
  jor  g11645(.dina(n11900), .dinb(n11899), .dout(n11901));
  jor  g11646(.dina(n10049), .dinb(n544), .dout(n11902));
  jor  g11647(.dina(n486), .dinb(n9475), .dout(n11903));
  jor  g11648(.dina(n547), .dinb(n9759), .dout(n11904));
  jor  g11649(.dina(n542), .dinb(n10051), .dout(n11905));
  jand g11650(.dina(n11905), .dinb(n11904), .dout(n11906));
  jand g11651(.dina(n11906), .dinb(n11903), .dout(n11907));
  jand g11652(.dina(n11907), .dinb(n11902), .dout(n11908));
  jxor g11653(.dina(n11908), .dinb(n446), .dout(n11909));
  jxor g11654(.dina(n11909), .dinb(n11901), .dout(n11910));
  jxor g11655(.dina(n11910), .dinb(n11898), .dout(n11911));
  jand g11656(.dina(n11636), .dinb(n11628), .dout(n11912));
  jand g11657(.dina(n11637), .dinb(n11625), .dout(n11913));
  jor  g11658(.dina(n11913), .dinb(n11912), .dout(n11914));
  jnot g11659(.din(n11914), .dout(n11915));
  jnot g11660(.din(n354), .dout(n11916));
  jand g11661(.dina(n11916), .dinb(b63 ), .dout(n11917));
  jand g11662(.dina(n10832), .dinb(n321), .dout(n11918));
  jor  g11663(.dina(n11918), .dinb(n11917), .dout(n11919));
  jxor g11664(.dina(n11919), .dinb(n364), .dout(n11920));
  jxor g11665(.dina(n11920), .dinb(n11915), .dout(n11921));
  jxor g11666(.dina(n11921), .dinb(n11911), .dout(n11922));
  jxor g11667(.dina(n11922), .dinb(n11662), .dout(n11923));
  jnot g11668(.din(n11923), .dout(n11924));
  jxor g11669(.dina(n11924), .dinb(n11657), .dout(f68 ));
  jand g11670(.dina(n11922), .dinb(n11662), .dout(n11926));
  jnot g11671(.din(n11926), .dout(n11927));
  jor  g11672(.dina(n11924), .dinb(n11657), .dout(n11928));
  jand g11673(.dina(n11928), .dinb(n11927), .dout(n11929));
  jor  g11674(.dina(n11920), .dinb(n11915), .dout(n11930));
  jand g11675(.dina(n11921), .dinb(n11911), .dout(n11931));
  jnot g11676(.din(n11931), .dout(n11932));
  jand g11677(.dina(n11932), .dinb(n11930), .dout(n11933));
  jnot g11678(.din(n11933), .dout(n11934));
  jand g11679(.dina(n11909), .dinb(n11901), .dout(n11935));
  jand g11680(.dina(n11910), .dinb(n11898), .dout(n11936));
  jor  g11681(.dina(n11936), .dinb(n11935), .dout(n11937));
  jor  g11682(.dina(n10521), .dinb(n544), .dout(n11938));
  jor  g11683(.dina(n486), .dinb(n9759), .dout(n11939));
  jor  g11684(.dina(n547), .dinb(n10051), .dout(n11940));
  jor  g11685(.dina(n542), .dinb(n10523), .dout(n11941));
  jand g11686(.dina(n11941), .dinb(n11940), .dout(n11942));
  jand g11687(.dina(n11942), .dinb(n11939), .dout(n11943));
  jand g11688(.dina(n11943), .dinb(n11938), .dout(n11944));
  jxor g11689(.dina(n11944), .dinb(n446), .dout(n11945));
  jxor g11690(.dina(n11945), .dinb(n11937), .dout(n11946));
  jand g11691(.dina(n11673), .dinb(n11665), .dout(n11947));
  jand g11692(.dina(n11897), .dinb(n11674), .dout(n11948));
  jor  g11693(.dina(n11948), .dinb(n11947), .dout(n11949));
  jor  g11694(.dina(n9473), .dinb(n728), .dout(n11950));
  jor  g11695(.dina(n660), .dinb(n8920), .dout(n11951));
  jor  g11696(.dina(n726), .dinb(n9475), .dout(n11952));
  jor  g11697(.dina(n731), .dinb(n9195), .dout(n11953));
  jand g11698(.dina(n11953), .dinb(n11952), .dout(n11954));
  jand g11699(.dina(n11954), .dinb(n11951), .dout(n11955));
  jand g11700(.dina(n11955), .dinb(n11950), .dout(n11956));
  jxor g11701(.dina(n11956), .dinb(n606), .dout(n11957));
  jxor g11702(.dina(n11957), .dinb(n11949), .dout(n11958));
  jand g11703(.dina(n11895), .dinb(n11887), .dout(n11959));
  jand g11704(.dina(n11896), .dinb(n11884), .dout(n11960));
  jor  g11705(.dina(n11960), .dinb(n11959), .dout(n11961));
  jor  g11706(.dina(n8642), .dinb(n970), .dout(n11962));
  jor  g11707(.dina(n880), .dinb(n8111), .dout(n11963));
  jor  g11708(.dina(n972), .dinb(n8644), .dout(n11964));
  jor  g11709(.dina(n967), .dinb(n8378), .dout(n11965));
  jand g11710(.dina(n11965), .dinb(n11964), .dout(n11966));
  jand g11711(.dina(n11966), .dinb(n11963), .dout(n11967));
  jand g11712(.dina(n11967), .dinb(n11962), .dout(n11968));
  jxor g11713(.dina(n11968), .dinb(n810), .dout(n11969));
  jxor g11714(.dina(n11969), .dinb(n11961), .dout(n11970));
  jand g11715(.dina(n11685), .dinb(n11677), .dout(n11971));
  jand g11716(.dina(n11883), .dinb(n11686), .dout(n11972));
  jor  g11717(.dina(n11972), .dinb(n11971), .dout(n11973));
  jor  g11718(.dina(n7844), .dinb(n1248), .dout(n11974));
  jor  g11719(.dina(n1147), .dinb(n7338), .dout(n11975));
  jor  g11720(.dina(n1251), .dinb(n7590), .dout(n11976));
  jor  g11721(.dina(n1246), .dinb(n7846), .dout(n11977));
  jand g11722(.dina(n11977), .dinb(n11976), .dout(n11978));
  jand g11723(.dina(n11978), .dinb(n11975), .dout(n11979));
  jand g11724(.dina(n11979), .dinb(n11974), .dout(n11980));
  jxor g11725(.dina(n11980), .dinb(n1061), .dout(n11981));
  jxor g11726(.dina(n11981), .dinb(n11973), .dout(n11982));
  jand g11727(.dina(n11881), .dinb(n11873), .dout(n11983));
  jand g11728(.dina(n11882), .dinb(n11870), .dout(n11984));
  jor  g11729(.dina(n11984), .dinb(n11983), .dout(n11985));
  jor  g11730(.dina(n7084), .dinb(n1569), .dout(n11986));
  jor  g11731(.dina(n1453), .dinb(n6605), .dout(n11987));
  jor  g11732(.dina(n1566), .dinb(n6846), .dout(n11988));
  jor  g11733(.dina(n1571), .dinb(n7086), .dout(n11989));
  jand g11734(.dina(n11989), .dinb(n11988), .dout(n11990));
  jand g11735(.dina(n11990), .dinb(n11987), .dout(n11991));
  jand g11736(.dina(n11991), .dinb(n11986), .dout(n11992));
  jxor g11737(.dina(n11992), .dinb(n1351), .dout(n11993));
  jxor g11738(.dina(n11993), .dinb(n11985), .dout(n11994));
  jand g11739(.dina(n11697), .dinb(n11689), .dout(n11995));
  jand g11740(.dina(n11869), .dinb(n11698), .dout(n11996));
  jor  g11741(.dina(n11996), .dinb(n11995), .dout(n11997));
  jor  g11742(.dina(n6364), .dinb(n1921), .dout(n11998));
  jor  g11743(.dina(n1806), .dinb(n5911), .dout(n11999));
  jor  g11744(.dina(n1923), .dinb(n6366), .dout(n12000));
  jor  g11745(.dina(n1918), .dinb(n6139), .dout(n12001));
  jand g11746(.dina(n12001), .dinb(n12000), .dout(n12002));
  jand g11747(.dina(n12002), .dinb(n11999), .dout(n12003));
  jand g11748(.dina(n12003), .dinb(n11998), .dout(n12004));
  jxor g11749(.dina(n12004), .dinb(n1687), .dout(n12005));
  jxor g11750(.dina(n12005), .dinb(n11997), .dout(n12006));
  jand g11751(.dina(n11709), .dinb(n11701), .dout(n12007));
  jand g11752(.dina(n11855), .dinb(n11710), .dout(n12008));
  jor  g11753(.dina(n12008), .dinb(n12007), .dout(n12009));
  jor  g11754(.dina(n5038), .dinb(n2764), .dout(n12010));
  jor  g11755(.dina(n2609), .dinb(n4637), .dout(n12011));
  jor  g11756(.dina(n2761), .dinb(n5040), .dout(n12012));
  jor  g11757(.dina(n2766), .dinb(n4839), .dout(n12013));
  jand g11758(.dina(n12013), .dinb(n12012), .dout(n12014));
  jand g11759(.dina(n12014), .dinb(n12011), .dout(n12015));
  jand g11760(.dina(n12015), .dinb(n12010), .dout(n12016));
  jxor g11761(.dina(n12016), .dinb(n2468), .dout(n12017));
  jxor g11762(.dina(n12017), .dinb(n12009), .dout(n12018));
  jand g11763(.dina(n11844), .dinb(n11841), .dout(n12019));
  jand g11764(.dina(n11853), .dinb(n11845), .dout(n12020));
  jor  g11765(.dina(n12020), .dinb(n12019), .dout(n12021));
  jand g11766(.dina(n11831), .dinb(n11725), .dout(n12022));
  jand g11767(.dina(n11840), .dinb(n11832), .dout(n12023));
  jor  g11768(.dina(n12023), .dinb(n12022), .dout(n12024));
  jand g11769(.dina(n11821), .dinb(n11728), .dout(n12025));
  jand g11770(.dina(n11830), .dinb(n11822), .dout(n12026));
  jor  g11771(.dina(n12026), .dinb(n12025), .dout(n12027));
  jand g11772(.dina(n11811), .dinb(n11731), .dout(n12028));
  jand g11773(.dina(n11820), .dinb(n11812), .dout(n12029));
  jor  g11774(.dina(n12029), .dinb(n12028), .dout(n12030));
  jand g11775(.dina(n11801), .dinb(n11798), .dout(n12031));
  jand g11776(.dina(n11810), .dinb(n11802), .dout(n12032));
  jor  g11777(.dina(n12032), .dinb(n12031), .dout(n12033));
  jand g11778(.dina(n11788), .dinb(n11734), .dout(n12034));
  jand g11779(.dina(n11797), .dinb(n11789), .dout(n12035));
  jor  g11780(.dina(n12035), .dinb(n12034), .dout(n12036));
  jand g11781(.dina(n11778), .dinb(n11737), .dout(n12037));
  jand g11782(.dina(n11787), .dinb(n11779), .dout(n12038));
  jor  g11783(.dina(n12038), .dinb(n12037), .dout(n12039));
  jand g11784(.dina(n11768), .dinb(n11765), .dout(n12040));
  jand g11785(.dina(n11777), .dinb(n11769), .dout(n12041));
  jor  g11786(.dina(n12041), .dinb(n12040), .dout(n12042));
  jand g11787(.dina(n11755), .dinb(n11742), .dout(n12043));
  jand g11788(.dina(n11764), .dinb(n11756), .dout(n12044));
  jor  g11789(.dina(n12044), .dinb(n12043), .dout(n12045));
  jand g11790(.dina(n11745), .dinb(a2 ), .dout(n12046));
  jand g11791(.dina(n11754), .dinb(n11746), .dout(n12047));
  jor  g11792(.dina(n12047), .dinb(n12046), .dout(n12048));
  jand g11793(.dina(n10594), .dinb(b5 ), .dout(n12049));
  jand g11794(.dina(n10129), .dinb(b6 ), .dout(n12050));
  jor  g11795(.dina(n12050), .dinb(n12049), .dout(n12051));
  jxor g11796(.dina(a5 ), .dinb(a2 ), .dout(n12052));
  jxor g11797(.dina(n12052), .dinb(n12051), .dout(n12053));
  jxor g11798(.dina(n12053), .dinb(n12048), .dout(n12054));
  jor  g11799(.dina(n10134), .dinb(n570), .dout(n12055));
  jor  g11800(.dina(n9849), .dinb(n469), .dout(n12056));
  jor  g11801(.dina(n10137), .dinb(n519), .dout(n12057));
  jor  g11802(.dina(n10132), .dinb(n572), .dout(n12058));
  jand g11803(.dina(n12058), .dinb(n12057), .dout(n12059));
  jand g11804(.dina(n12059), .dinb(n12056), .dout(n12060));
  jand g11805(.dina(n12060), .dinb(n12055), .dout(n12061));
  jxor g11806(.dina(n12061), .dinb(n9559), .dout(n12062));
  jxor g11807(.dina(n12062), .dinb(n12054), .dout(n12063));
  jor  g11808(.dina(n9271), .dinb(n770), .dout(n12064));
  jor  g11809(.dina(n9003), .dinb(n637), .dout(n12065));
  jor  g11810(.dina(n9268), .dinb(n772), .dout(n12066));
  jor  g11811(.dina(n9273), .dinb(n704), .dout(n12067));
  jand g11812(.dina(n12067), .dinb(n12066), .dout(n12068));
  jand g11813(.dina(n12068), .dinb(n12065), .dout(n12069));
  jand g11814(.dina(n12069), .dinb(n12064), .dout(n12070));
  jxor g11815(.dina(n12070), .dinb(n8729), .dout(n12071));
  jxor g11816(.dina(n12071), .dinb(n12063), .dout(n12072));
  jxor g11817(.dina(n12072), .dinb(n12045), .dout(n12073));
  jor  g11818(.dina(n8457), .dinb(n1016), .dout(n12074));
  jor  g11819(.dina(n8185), .dinb(n852), .dout(n12075));
  jor  g11820(.dina(n8459), .dinb(n934), .dout(n12076));
  jor  g11821(.dina(n8454), .dinb(n1018), .dout(n12077));
  jand g11822(.dina(n12077), .dinb(n12076), .dout(n12078));
  jand g11823(.dina(n12078), .dinb(n12075), .dout(n12079));
  jand g11824(.dina(n12079), .dinb(n12074), .dout(n12080));
  jxor g11825(.dina(n12080), .dinb(n7929), .dout(n12081));
  jxor g11826(.dina(n12081), .dinb(n12073), .dout(n12082));
  jxor g11827(.dina(n12082), .dinb(n12042), .dout(n12083));
  jor  g11828(.dina(n7660), .dinb(n1305), .dout(n12084));
  jor  g11829(.dina(n7415), .dinb(n1114), .dout(n12085));
  jor  g11830(.dina(n7657), .dinb(n1211), .dout(n12086));
  jor  g11831(.dina(n7662), .dinb(n1307), .dout(n12087));
  jand g11832(.dina(n12087), .dinb(n12086), .dout(n12088));
  jand g11833(.dina(n12088), .dinb(n12085), .dout(n12089));
  jand g11834(.dina(n12089), .dinb(n12084), .dout(n12090));
  jxor g11835(.dina(n12090), .dinb(n7166), .dout(n12091));
  jxor g11836(.dina(n12091), .dinb(n12083), .dout(n12092));
  jxor g11837(.dina(n12092), .dinb(n12039), .dout(n12093));
  jor  g11838(.dina(n6914), .dinb(n1635), .dout(n12094));
  jor  g11839(.dina(n6673), .dinb(n1416), .dout(n12095));
  jor  g11840(.dina(n6911), .dinb(n1527), .dout(n12096));
  jor  g11841(.dina(n6916), .dinb(n1637), .dout(n12097));
  jand g11842(.dina(n12097), .dinb(n12096), .dout(n12098));
  jand g11843(.dina(n12098), .dinb(n12095), .dout(n12099));
  jand g11844(.dina(n12099), .dinb(n12094), .dout(n12100));
  jxor g11845(.dina(n12100), .dinb(n6443), .dout(n12101));
  jxor g11846(.dina(n12101), .dinb(n12093), .dout(n12102));
  jxor g11847(.dina(n12102), .dinb(n12036), .dout(n12103));
  jor  g11848(.dina(n6207), .dinb(n2005), .dout(n12104));
  jor  g11849(.dina(n5975), .dinb(n1759), .dout(n12105));
  jor  g11850(.dina(n6205), .dinb(n2007), .dout(n12106));
  jor  g11851(.dina(n6210), .dinb(n1881), .dout(n12107));
  jand g11852(.dina(n12107), .dinb(n12106), .dout(n12108));
  jand g11853(.dina(n12108), .dinb(n12105), .dout(n12109));
  jand g11854(.dina(n12109), .dinb(n12104), .dout(n12110));
  jxor g11855(.dina(n12110), .dinb(n5759), .dout(n12111));
  jxor g11856(.dina(n12111), .dinb(n12103), .dout(n12112));
  jxor g11857(.dina(n12112), .dinb(n12033), .dout(n12113));
  jor  g11858(.dina(n5537), .dinb(n2413), .dout(n12114));
  jor  g11859(.dina(n5315), .dinb(n2142), .dout(n12115));
  jor  g11860(.dina(n5534), .dinb(n2279), .dout(n12116));
  jor  g11861(.dina(n5539), .dinb(n2415), .dout(n12117));
  jand g11862(.dina(n12117), .dinb(n12116), .dout(n12118));
  jand g11863(.dina(n12118), .dinb(n12115), .dout(n12119));
  jand g11864(.dina(n12119), .dinb(n12114), .dout(n12120));
  jxor g11865(.dina(n12120), .dinb(n5111), .dout(n12121));
  jxor g11866(.dina(n12121), .dinb(n12113), .dout(n12122));
  jxor g11867(.dina(n12122), .dinb(n12030), .dout(n12123));
  jor  g11868(.dina(n4902), .dinb(n2860), .dout(n12124));
  jor  g11869(.dina(n4696), .dinb(n2563), .dout(n12125));
  jor  g11870(.dina(n4904), .dinb(n2713), .dout(n12126));
  jor  g11871(.dina(n4899), .dinb(n2862), .dout(n12127));
  jand g11872(.dina(n12127), .dinb(n12126), .dout(n12128));
  jand g11873(.dina(n12128), .dinb(n12125), .dout(n12129));
  jand g11874(.dina(n12129), .dinb(n12124), .dout(n12130));
  jxor g11875(.dina(n12130), .dinb(n4505), .dout(n12131));
  jxor g11876(.dina(n12131), .dinb(n12123), .dout(n12132));
  jxor g11877(.dina(n12132), .dinb(n12027), .dout(n12133));
  jor  g11878(.dina(n4305), .dinb(n3346), .dout(n12134));
  jor  g11879(.dina(n4116), .dinb(n3023), .dout(n12135));
  jor  g11880(.dina(n4308), .dinb(n3186), .dout(n12136));
  jor  g11881(.dina(n4303), .dinb(n3348), .dout(n12137));
  jand g11882(.dina(n12137), .dinb(n12136), .dout(n12138));
  jand g11883(.dina(n12138), .dinb(n12135), .dout(n12139));
  jand g11884(.dina(n12139), .dinb(n12134), .dout(n12140));
  jxor g11885(.dina(n12140), .dinb(n3938), .dout(n12141));
  jxor g11886(.dina(n12141), .dinb(n12133), .dout(n12142));
  jxor g11887(.dina(n12142), .dinb(n12024), .dout(n12143));
  jor  g11888(.dina(n3871), .dinb(n3751), .dout(n12144));
  jor  g11889(.dina(n3574), .dinb(n3522), .dout(n12145));
  jor  g11890(.dina(n3749), .dinb(n3873), .dout(n12146));
  jor  g11891(.dina(n3754), .dinb(n3698), .dout(n12147));
  jand g11892(.dina(n12147), .dinb(n12146), .dout(n12148));
  jand g11893(.dina(n12148), .dinb(n12145), .dout(n12149));
  jand g11894(.dina(n12149), .dinb(n12144), .dout(n12150));
  jxor g11895(.dina(n12150), .dinb(n3410), .dout(n12151));
  jxor g11896(.dina(n12151), .dinb(n12143), .dout(n12152));
  jxor g11897(.dina(n12152), .dinb(n12021), .dout(n12153));
  jand g11898(.dina(n11721), .dinb(n11713), .dout(n12154));
  jand g11899(.dina(n11854), .dinb(n11722), .dout(n12155));
  jor  g11900(.dina(n12155), .dinb(n12154), .dout(n12156));
  jor  g11901(.dina(n4435), .dinb(n3239), .dout(n12157));
  jor  g11902(.dina(n3072), .dinb(n4060), .dout(n12158));
  jor  g11903(.dina(n3242), .dinb(n4249), .dout(n12159));
  jor  g11904(.dina(n3237), .dinb(n4437), .dout(n12160));
  jand g11905(.dina(n12160), .dinb(n12159), .dout(n12161));
  jand g11906(.dina(n12161), .dinb(n12158), .dout(n12162));
  jand g11907(.dina(n12162), .dinb(n12157), .dout(n12163));
  jxor g11908(.dina(n12163), .dinb(n2918), .dout(n12164));
  jxor g11909(.dina(n12164), .dinb(n12156), .dout(n12165));
  jxor g11910(.dina(n12165), .dinb(n12153), .dout(n12166));
  jxor g11911(.dina(n12166), .dinb(n12018), .dout(n12167));
  jand g11912(.dina(n11867), .dinb(n11859), .dout(n12168));
  jand g11913(.dina(n11868), .dinb(n11856), .dout(n12169));
  jor  g11914(.dina(n12169), .dinb(n12168), .dout(n12170));
  jor  g11915(.dina(n5683), .dinb(n2324), .dout(n12171));
  jor  g11916(.dina(n2186), .dinb(n5253), .dout(n12172));
  jor  g11917(.dina(n2321), .dinb(n5469), .dout(n12173));
  jor  g11918(.dina(n2326), .dinb(n5685), .dout(n12174));
  jand g11919(.dina(n12174), .dinb(n12173), .dout(n12175));
  jand g11920(.dina(n12175), .dinb(n12172), .dout(n12176));
  jand g11921(.dina(n12176), .dinb(n12171), .dout(n12177));
  jxor g11922(.dina(n12177), .dinb(n2057), .dout(n12178));
  jxor g11923(.dina(n12178), .dinb(n12170), .dout(n12179));
  jxor g11924(.dina(n12179), .dinb(n12167), .dout(n12180));
  jxor g11925(.dina(n12180), .dinb(n12006), .dout(n12181));
  jxor g11926(.dina(n12181), .dinb(n11994), .dout(n12182));
  jxor g11927(.dina(n12182), .dinb(n11982), .dout(n12183));
  jxor g11928(.dina(n12183), .dinb(n11970), .dout(n12184));
  jxor g11929(.dina(n12184), .dinb(n11958), .dout(n12185));
  jxor g11930(.dina(n12185), .dinb(n11946), .dout(n12186));
  jxor g11931(.dina(n12186), .dinb(n11934), .dout(n12187));
  jnot g11932(.din(n12187), .dout(n12188));
  jxor g11933(.dina(n12188), .dinb(n11929), .dout(f69 ));
  jand g11934(.dina(n12186), .dinb(n11934), .dout(n12190));
  jnot g11935(.din(n12190), .dout(n12191));
  jor  g11936(.dina(n12188), .dinb(n11929), .dout(n12192));
  jand g11937(.dina(n12192), .dinb(n12191), .dout(n12193));
  jand g11938(.dina(n11945), .dinb(n11937), .dout(n12194));
  jand g11939(.dina(n12185), .dinb(n11946), .dout(n12195));
  jor  g11940(.dina(n12195), .dinb(n12194), .dout(n12196));
  jand g11941(.dina(n11957), .dinb(n11949), .dout(n12197));
  jand g11942(.dina(n12184), .dinb(n11958), .dout(n12198));
  jor  g11943(.dina(n12198), .dinb(n12197), .dout(n12199));
  jnot g11944(.din(n12199), .dout(n12200));
  jor  g11945(.dina(n10813), .dinb(n544), .dout(n12201));
  jor  g11946(.dina(n486), .dinb(n10051), .dout(n12202));
  jor  g11947(.dina(n547), .dinb(n10523), .dout(n12203));
  jand g11948(.dina(n12203), .dinb(n12202), .dout(n12204));
  jand g11949(.dina(n12204), .dinb(n12201), .dout(n12205));
  jxor g11950(.dina(n12205), .dinb(a8 ), .dout(n12206));
  jxor g11951(.dina(n12206), .dinb(n12200), .dout(n12207));
  jand g11952(.dina(n11969), .dinb(n11961), .dout(n12208));
  jand g11953(.dina(n12183), .dinb(n11970), .dout(n12209));
  jor  g11954(.dina(n12209), .dinb(n12208), .dout(n12210));
  jor  g11955(.dina(n9757), .dinb(n728), .dout(n12211));
  jor  g11956(.dina(n660), .dinb(n9195), .dout(n12212));
  jor  g11957(.dina(n731), .dinb(n9475), .dout(n12213));
  jor  g11958(.dina(n726), .dinb(n9759), .dout(n12214));
  jand g11959(.dina(n12214), .dinb(n12213), .dout(n12215));
  jand g11960(.dina(n12215), .dinb(n12212), .dout(n12216));
  jand g11961(.dina(n12216), .dinb(n12211), .dout(n12217));
  jxor g11962(.dina(n12217), .dinb(n606), .dout(n12218));
  jxor g11963(.dina(n12218), .dinb(n12210), .dout(n12219));
  jand g11964(.dina(n11981), .dinb(n11973), .dout(n12220));
  jand g11965(.dina(n12182), .dinb(n11982), .dout(n12221));
  jor  g11966(.dina(n12221), .dinb(n12220), .dout(n12222));
  jor  g11967(.dina(n8918), .dinb(n970), .dout(n12223));
  jor  g11968(.dina(n880), .dinb(n8378), .dout(n12224));
  jor  g11969(.dina(n972), .dinb(n8920), .dout(n12225));
  jor  g11970(.dina(n967), .dinb(n8644), .dout(n12226));
  jand g11971(.dina(n12226), .dinb(n12225), .dout(n12227));
  jand g11972(.dina(n12227), .dinb(n12224), .dout(n12228));
  jand g11973(.dina(n12228), .dinb(n12223), .dout(n12229));
  jxor g11974(.dina(n12229), .dinb(n810), .dout(n12230));
  jxor g11975(.dina(n12230), .dinb(n12222), .dout(n12231));
  jand g11976(.dina(n11993), .dinb(n11985), .dout(n12232));
  jand g11977(.dina(n12181), .dinb(n11994), .dout(n12233));
  jor  g11978(.dina(n12233), .dinb(n12232), .dout(n12234));
  jor  g11979(.dina(n8109), .dinb(n1248), .dout(n12235));
  jor  g11980(.dina(n1147), .dinb(n7590), .dout(n12236));
  jor  g11981(.dina(n1246), .dinb(n8111), .dout(n12237));
  jor  g11982(.dina(n1251), .dinb(n7846), .dout(n12238));
  jand g11983(.dina(n12238), .dinb(n12237), .dout(n12239));
  jand g11984(.dina(n12239), .dinb(n12236), .dout(n12240));
  jand g11985(.dina(n12240), .dinb(n12235), .dout(n12241));
  jxor g11986(.dina(n12241), .dinb(n1061), .dout(n12242));
  jxor g11987(.dina(n12242), .dinb(n12234), .dout(n12243));
  jand g11988(.dina(n12005), .dinb(n11997), .dout(n12244));
  jand g11989(.dina(n12180), .dinb(n12006), .dout(n12245));
  jor  g11990(.dina(n12245), .dinb(n12244), .dout(n12246));
  jor  g11991(.dina(n7336), .dinb(n1569), .dout(n12247));
  jor  g11992(.dina(n1453), .dinb(n6846), .dout(n12248));
  jor  g11993(.dina(n1571), .dinb(n7338), .dout(n12249));
  jor  g11994(.dina(n1566), .dinb(n7086), .dout(n12250));
  jand g11995(.dina(n12250), .dinb(n12249), .dout(n12251));
  jand g11996(.dina(n12251), .dinb(n12248), .dout(n12252));
  jand g11997(.dina(n12252), .dinb(n12247), .dout(n12253));
  jxor g11998(.dina(n12253), .dinb(n1351), .dout(n12254));
  jxor g11999(.dina(n12254), .dinb(n12246), .dout(n12255));
  jand g12000(.dina(n12017), .dinb(n12009), .dout(n12256));
  jand g12001(.dina(n12166), .dinb(n12018), .dout(n12257));
  jor  g12002(.dina(n12257), .dinb(n12256), .dout(n12258));
  jor  g12003(.dina(n5909), .dinb(n2324), .dout(n12259));
  jor  g12004(.dina(n2186), .dinb(n5469), .dout(n12260));
  jor  g12005(.dina(n2326), .dinb(n5911), .dout(n12261));
  jor  g12006(.dina(n2321), .dinb(n5685), .dout(n12262));
  jand g12007(.dina(n12262), .dinb(n12261), .dout(n12263));
  jand g12008(.dina(n12263), .dinb(n12260), .dout(n12264));
  jand g12009(.dina(n12264), .dinb(n12259), .dout(n12265));
  jxor g12010(.dina(n12265), .dinb(n2057), .dout(n12266));
  jxor g12011(.dina(n12266), .dinb(n12258), .dout(n12267));
  jand g12012(.dina(n12164), .dinb(n12156), .dout(n12268));
  jand g12013(.dina(n12165), .dinb(n12153), .dout(n12269));
  jor  g12014(.dina(n12269), .dinb(n12268), .dout(n12270));
  jor  g12015(.dina(n5251), .dinb(n2764), .dout(n12271));
  jor  g12016(.dina(n2609), .dinb(n4839), .dout(n12272));
  jor  g12017(.dina(n2761), .dinb(n5253), .dout(n12273));
  jor  g12018(.dina(n2766), .dinb(n5040), .dout(n12274));
  jand g12019(.dina(n12274), .dinb(n12273), .dout(n12275));
  jand g12020(.dina(n12275), .dinb(n12272), .dout(n12276));
  jand g12021(.dina(n12276), .dinb(n12271), .dout(n12277));
  jxor g12022(.dina(n12277), .dinb(n2468), .dout(n12278));
  jxor g12023(.dina(n12278), .dinb(n12270), .dout(n12279));
  jand g12024(.dina(n12151), .dinb(n12143), .dout(n12280));
  jand g12025(.dina(n12152), .dinb(n12021), .dout(n12281));
  jor  g12026(.dina(n12281), .dinb(n12280), .dout(n12282));
  jor  g12027(.dina(n4635), .dinb(n3239), .dout(n12283));
  jor  g12028(.dina(n3072), .dinb(n4249), .dout(n12284));
  jor  g12029(.dina(n3237), .dinb(n4637), .dout(n12285));
  jor  g12030(.dina(n3242), .dinb(n4437), .dout(n12286));
  jand g12031(.dina(n12286), .dinb(n12285), .dout(n12287));
  jand g12032(.dina(n12287), .dinb(n12284), .dout(n12288));
  jand g12033(.dina(n12288), .dinb(n12283), .dout(n12289));
  jxor g12034(.dina(n12289), .dinb(n2918), .dout(n12290));
  jxor g12035(.dina(n12290), .dinb(n12282), .dout(n12291));
  jand g12036(.dina(n12141), .dinb(n12133), .dout(n12292));
  jand g12037(.dina(n12142), .dinb(n12024), .dout(n12293));
  jor  g12038(.dina(n12293), .dinb(n12292), .dout(n12294));
  jand g12039(.dina(n12121), .dinb(n12113), .dout(n12295));
  jand g12040(.dina(n12122), .dinb(n12030), .dout(n12296));
  jor  g12041(.dina(n12296), .dinb(n12295), .dout(n12297));
  jand g12042(.dina(n12111), .dinb(n12103), .dout(n12298));
  jand g12043(.dina(n12112), .dinb(n12033), .dout(n12299));
  jor  g12044(.dina(n12299), .dinb(n12298), .dout(n12300));
  jand g12045(.dina(n12101), .dinb(n12093), .dout(n12301));
  jand g12046(.dina(n12102), .dinb(n12036), .dout(n12302));
  jor  g12047(.dina(n12302), .dinb(n12301), .dout(n12303));
  jand g12048(.dina(n12091), .dinb(n12083), .dout(n12304));
  jand g12049(.dina(n12092), .dinb(n12039), .dout(n12305));
  jor  g12050(.dina(n12305), .dinb(n12304), .dout(n12306));
  jand g12051(.dina(n12081), .dinb(n12073), .dout(n12307));
  jand g12052(.dina(n12082), .dinb(n12042), .dout(n12308));
  jor  g12053(.dina(n12308), .dinb(n12307), .dout(n12309));
  jand g12054(.dina(n12071), .dinb(n12063), .dout(n12310));
  jand g12055(.dina(n12072), .dinb(n12045), .dout(n12311));
  jor  g12056(.dina(n12311), .dinb(n12310), .dout(n12312));
  jand g12057(.dina(n12053), .dinb(n12048), .dout(n12313));
  jand g12058(.dina(n12062), .dinb(n12054), .dout(n12314));
  jor  g12059(.dina(n12314), .dinb(n12313), .dout(n12315));
  jand g12060(.dina(n364), .dinb(n278), .dout(n12316));
  jand g12061(.dina(n12052), .dinb(n12051), .dout(n12317));
  jor  g12062(.dina(n12317), .dinb(n12316), .dout(n12318));
  jand g12063(.dina(n10594), .dinb(b6 ), .dout(n12319));
  jand g12064(.dina(n10129), .dinb(b7 ), .dout(n12320));
  jor  g12065(.dina(n12320), .dinb(n12319), .dout(n12321));
  jnot g12066(.din(n12321), .dout(n12322));
  jxor g12067(.dina(n12322), .dinb(n12318), .dout(n12323));
  jor  g12068(.dina(n10134), .dinb(n635), .dout(n12324));
  jor  g12069(.dina(n9849), .dinb(n519), .dout(n12325));
  jor  g12070(.dina(n10137), .dinb(n572), .dout(n12326));
  jor  g12071(.dina(n10132), .dinb(n637), .dout(n12327));
  jand g12072(.dina(n12327), .dinb(n12326), .dout(n12328));
  jand g12073(.dina(n12328), .dinb(n12325), .dout(n12329));
  jand g12074(.dina(n12329), .dinb(n12324), .dout(n12330));
  jxor g12075(.dina(n12330), .dinb(n9559), .dout(n12331));
  jxor g12076(.dina(n12331), .dinb(n12323), .dout(n12332));
  jxor g12077(.dina(n12332), .dinb(n12315), .dout(n12333));
  jor  g12078(.dina(n9271), .dinb(n850), .dout(n12334));
  jor  g12079(.dina(n9003), .dinb(n704), .dout(n12335));
  jor  g12080(.dina(n9268), .dinb(n852), .dout(n12336));
  jor  g12081(.dina(n9273), .dinb(n772), .dout(n12337));
  jand g12082(.dina(n12337), .dinb(n12336), .dout(n12338));
  jand g12083(.dina(n12338), .dinb(n12335), .dout(n12339));
  jand g12084(.dina(n12339), .dinb(n12334), .dout(n12340));
  jxor g12085(.dina(n12340), .dinb(n8729), .dout(n12341));
  jxor g12086(.dina(n12341), .dinb(n12333), .dout(n12342));
  jxor g12087(.dina(n12342), .dinb(n12312), .dout(n12343));
  jor  g12088(.dina(n8457), .dinb(n1112), .dout(n12344));
  jor  g12089(.dina(n8185), .dinb(n934), .dout(n12345));
  jor  g12090(.dina(n8459), .dinb(n1018), .dout(n12346));
  jor  g12091(.dina(n8454), .dinb(n1114), .dout(n12347));
  jand g12092(.dina(n12347), .dinb(n12346), .dout(n12348));
  jand g12093(.dina(n12348), .dinb(n12345), .dout(n12349));
  jand g12094(.dina(n12349), .dinb(n12344), .dout(n12350));
  jxor g12095(.dina(n12350), .dinb(n7929), .dout(n12351));
  jxor g12096(.dina(n12351), .dinb(n12343), .dout(n12352));
  jxor g12097(.dina(n12352), .dinb(n12309), .dout(n12353));
  jor  g12098(.dina(n7660), .dinb(n1414), .dout(n12354));
  jor  g12099(.dina(n7415), .dinb(n1211), .dout(n12355));
  jor  g12100(.dina(n7657), .dinb(n1307), .dout(n12356));
  jor  g12101(.dina(n7662), .dinb(n1416), .dout(n12357));
  jand g12102(.dina(n12357), .dinb(n12356), .dout(n12358));
  jand g12103(.dina(n12358), .dinb(n12355), .dout(n12359));
  jand g12104(.dina(n12359), .dinb(n12354), .dout(n12360));
  jxor g12105(.dina(n12360), .dinb(n7166), .dout(n12361));
  jxor g12106(.dina(n12361), .dinb(n12353), .dout(n12362));
  jxor g12107(.dina(n12362), .dinb(n12306), .dout(n12363));
  jor  g12108(.dina(n6914), .dinb(n1757), .dout(n12364));
  jor  g12109(.dina(n6673), .dinb(n1527), .dout(n12365));
  jor  g12110(.dina(n6911), .dinb(n1637), .dout(n12366));
  jor  g12111(.dina(n6916), .dinb(n1759), .dout(n12367));
  jand g12112(.dina(n12367), .dinb(n12366), .dout(n12368));
  jand g12113(.dina(n12368), .dinb(n12365), .dout(n12369));
  jand g12114(.dina(n12369), .dinb(n12364), .dout(n12370));
  jxor g12115(.dina(n12370), .dinb(n6443), .dout(n12371));
  jxor g12116(.dina(n12371), .dinb(n12363), .dout(n12372));
  jxor g12117(.dina(n12372), .dinb(n12303), .dout(n12373));
  jor  g12118(.dina(n6207), .dinb(n2140), .dout(n12374));
  jor  g12119(.dina(n5975), .dinb(n1881), .dout(n12375));
  jor  g12120(.dina(n6205), .dinb(n2142), .dout(n12376));
  jor  g12121(.dina(n6210), .dinb(n2007), .dout(n12377));
  jand g12122(.dina(n12377), .dinb(n12376), .dout(n12378));
  jand g12123(.dina(n12378), .dinb(n12375), .dout(n12379));
  jand g12124(.dina(n12379), .dinb(n12374), .dout(n12380));
  jxor g12125(.dina(n12380), .dinb(n5759), .dout(n12381));
  jxor g12126(.dina(n12381), .dinb(n12373), .dout(n12382));
  jxor g12127(.dina(n12382), .dinb(n12300), .dout(n12383));
  jor  g12128(.dina(n5537), .dinb(n2561), .dout(n12384));
  jor  g12129(.dina(n5315), .dinb(n2279), .dout(n12385));
  jor  g12130(.dina(n5539), .dinb(n2563), .dout(n12386));
  jor  g12131(.dina(n5534), .dinb(n2415), .dout(n12387));
  jand g12132(.dina(n12387), .dinb(n12386), .dout(n12388));
  jand g12133(.dina(n12388), .dinb(n12385), .dout(n12389));
  jand g12134(.dina(n12389), .dinb(n12384), .dout(n12390));
  jxor g12135(.dina(n12390), .dinb(n5111), .dout(n12391));
  jxor g12136(.dina(n12391), .dinb(n12383), .dout(n12392));
  jxor g12137(.dina(n12392), .dinb(n12297), .dout(n12393));
  jor  g12138(.dina(n4902), .dinb(n3021), .dout(n12394));
  jor  g12139(.dina(n4696), .dinb(n2713), .dout(n12395));
  jor  g12140(.dina(n4899), .dinb(n3023), .dout(n12396));
  jor  g12141(.dina(n4904), .dinb(n2862), .dout(n12397));
  jand g12142(.dina(n12397), .dinb(n12396), .dout(n12398));
  jand g12143(.dina(n12398), .dinb(n12395), .dout(n12399));
  jand g12144(.dina(n12399), .dinb(n12394), .dout(n12400));
  jxor g12145(.dina(n12400), .dinb(n4505), .dout(n12401));
  jxor g12146(.dina(n12401), .dinb(n12393), .dout(n12402));
  jnot g12147(.din(n12123), .dout(n12403));
  jnot g12148(.din(n12131), .dout(n12404));
  jand g12149(.dina(n12404), .dinb(n12403), .dout(n12405));
  jnot g12150(.din(n12405), .dout(n12406));
  jand g12151(.dina(n12131), .dinb(n12123), .dout(n12407));
  jor  g12152(.dina(n12407), .dinb(n12027), .dout(n12408));
  jand g12153(.dina(n12408), .dinb(n12406), .dout(n12409));
  jxor g12154(.dina(n12409), .dinb(n12402), .dout(n12410));
  jor  g12155(.dina(n4305), .dinb(n3520), .dout(n12411));
  jor  g12156(.dina(n4116), .dinb(n3186), .dout(n12412));
  jor  g12157(.dina(n4303), .dinb(n3522), .dout(n12413));
  jor  g12158(.dina(n4308), .dinb(n3348), .dout(n12414));
  jand g12159(.dina(n12414), .dinb(n12413), .dout(n12415));
  jand g12160(.dina(n12415), .dinb(n12412), .dout(n12416));
  jand g12161(.dina(n12416), .dinb(n12411), .dout(n12417));
  jxor g12162(.dina(n12417), .dinb(n3938), .dout(n12418));
  jxor g12163(.dina(n12418), .dinb(n12410), .dout(n12419));
  jxor g12164(.dina(n12419), .dinb(n12294), .dout(n12420));
  jor  g12165(.dina(n4058), .dinb(n3751), .dout(n12421));
  jor  g12166(.dina(n3574), .dinb(n3698), .dout(n12422));
  jor  g12167(.dina(n3749), .dinb(n4060), .dout(n12423));
  jor  g12168(.dina(n3754), .dinb(n3873), .dout(n12424));
  jand g12169(.dina(n12424), .dinb(n12423), .dout(n12425));
  jand g12170(.dina(n12425), .dinb(n12422), .dout(n12426));
  jand g12171(.dina(n12426), .dinb(n12421), .dout(n12427));
  jxor g12172(.dina(n12427), .dinb(n3410), .dout(n12428));
  jxor g12173(.dina(n12428), .dinb(n12420), .dout(n12429));
  jxor g12174(.dina(n12429), .dinb(n12291), .dout(n12430));
  jxor g12175(.dina(n12430), .dinb(n12279), .dout(n12431));
  jxor g12176(.dina(n12431), .dinb(n12267), .dout(n12432));
  jand g12177(.dina(n12178), .dinb(n12170), .dout(n12433));
  jand g12178(.dina(n12179), .dinb(n12167), .dout(n12434));
  jor  g12179(.dina(n12434), .dinb(n12433), .dout(n12435));
  jor  g12180(.dina(n6603), .dinb(n1921), .dout(n12436));
  jor  g12181(.dina(n1806), .dinb(n6139), .dout(n12437));
  jor  g12182(.dina(n1918), .dinb(n6366), .dout(n12438));
  jor  g12183(.dina(n1923), .dinb(n6605), .dout(n12439));
  jand g12184(.dina(n12439), .dinb(n12438), .dout(n12440));
  jand g12185(.dina(n12440), .dinb(n12437), .dout(n12441));
  jand g12186(.dina(n12441), .dinb(n12436), .dout(n12442));
  jxor g12187(.dina(n12442), .dinb(n1687), .dout(n12443));
  jxor g12188(.dina(n12443), .dinb(n12435), .dout(n12444));
  jxor g12189(.dina(n12444), .dinb(n12432), .dout(n12445));
  jxor g12190(.dina(n12445), .dinb(n12255), .dout(n12446));
  jxor g12191(.dina(n12446), .dinb(n12243), .dout(n12447));
  jxor g12192(.dina(n12447), .dinb(n12231), .dout(n12448));
  jxor g12193(.dina(n12448), .dinb(n12219), .dout(n12449));
  jxor g12194(.dina(n12449), .dinb(n12207), .dout(n12450));
  jxor g12195(.dina(n12450), .dinb(n12196), .dout(n12451));
  jnot g12196(.din(n12451), .dout(n12452));
  jxor g12197(.dina(n12452), .dinb(n12193), .dout(f70 ));
  jand g12198(.dina(n12450), .dinb(n12196), .dout(n12454));
  jnot g12199(.din(n12454), .dout(n12455));
  jor  g12200(.dina(n12452), .dinb(n12193), .dout(n12456));
  jand g12201(.dina(n12456), .dinb(n12455), .dout(n12457));
  jor  g12202(.dina(n12206), .dinb(n12200), .dout(n12458));
  jand g12203(.dina(n12449), .dinb(n12207), .dout(n12459));
  jnot g12204(.din(n12459), .dout(n12460));
  jand g12205(.dina(n12460), .dinb(n12458), .dout(n12461));
  jnot g12206(.din(n12461), .dout(n12462));
  jand g12207(.dina(n12254), .dinb(n12246), .dout(n12463));
  jand g12208(.dina(n12445), .dinb(n12255), .dout(n12464));
  jor  g12209(.dina(n12464), .dinb(n12463), .dout(n12465));
  jor  g12210(.dina(n8376), .dinb(n1248), .dout(n12466));
  jor  g12211(.dina(n1147), .dinb(n7846), .dout(n12467));
  jor  g12212(.dina(n1251), .dinb(n8111), .dout(n12468));
  jor  g12213(.dina(n1246), .dinb(n8378), .dout(n12469));
  jand g12214(.dina(n12469), .dinb(n12468), .dout(n12470));
  jand g12215(.dina(n12470), .dinb(n12467), .dout(n12471));
  jand g12216(.dina(n12471), .dinb(n12466), .dout(n12472));
  jxor g12217(.dina(n12472), .dinb(n1061), .dout(n12473));
  jxor g12218(.dina(n12473), .dinb(n12465), .dout(n12474));
  jand g12219(.dina(n12266), .dinb(n12258), .dout(n12475));
  jand g12220(.dina(n12431), .dinb(n12267), .dout(n12476));
  jor  g12221(.dina(n12476), .dinb(n12475), .dout(n12477));
  jor  g12222(.dina(n6844), .dinb(n1921), .dout(n12478));
  jor  g12223(.dina(n1806), .dinb(n6366), .dout(n12479));
  jor  g12224(.dina(n1918), .dinb(n6605), .dout(n12480));
  jor  g12225(.dina(n1923), .dinb(n6846), .dout(n12481));
  jand g12226(.dina(n12481), .dinb(n12480), .dout(n12482));
  jand g12227(.dina(n12482), .dinb(n12479), .dout(n12483));
  jand g12228(.dina(n12483), .dinb(n12478), .dout(n12484));
  jxor g12229(.dina(n12484), .dinb(n1687), .dout(n12485));
  jxor g12230(.dina(n12485), .dinb(n12477), .dout(n12486));
  jand g12231(.dina(n12290), .dinb(n12282), .dout(n12487));
  jand g12232(.dina(n12429), .dinb(n12291), .dout(n12488));
  jor  g12233(.dina(n12488), .dinb(n12487), .dout(n12489));
  jor  g12234(.dina(n5467), .dinb(n2764), .dout(n12490));
  jor  g12235(.dina(n2609), .dinb(n5040), .dout(n12491));
  jor  g12236(.dina(n2761), .dinb(n5469), .dout(n12492));
  jor  g12237(.dina(n2766), .dinb(n5253), .dout(n12493));
  jand g12238(.dina(n12493), .dinb(n12492), .dout(n12494));
  jand g12239(.dina(n12494), .dinb(n12491), .dout(n12495));
  jand g12240(.dina(n12495), .dinb(n12490), .dout(n12496));
  jxor g12241(.dina(n12496), .dinb(n2468), .dout(n12497));
  jxor g12242(.dina(n12497), .dinb(n12489), .dout(n12498));
  jand g12243(.dina(n12419), .dinb(n12294), .dout(n12499));
  jand g12244(.dina(n12428), .dinb(n12420), .dout(n12500));
  jor  g12245(.dina(n12500), .dinb(n12499), .dout(n12501));
  jor  g12246(.dina(n4837), .dinb(n3239), .dout(n12502));
  jor  g12247(.dina(n3072), .dinb(n4437), .dout(n12503));
  jor  g12248(.dina(n3237), .dinb(n4839), .dout(n12504));
  jor  g12249(.dina(n3242), .dinb(n4637), .dout(n12505));
  jand g12250(.dina(n12505), .dinb(n12504), .dout(n12506));
  jand g12251(.dina(n12506), .dinb(n12503), .dout(n12507));
  jand g12252(.dina(n12507), .dinb(n12502), .dout(n12508));
  jxor g12253(.dina(n12508), .dinb(n2918), .dout(n12509));
  jxor g12254(.dina(n12509), .dinb(n12501), .dout(n12510));
  jand g12255(.dina(n12409), .dinb(n12402), .dout(n12511));
  jand g12256(.dina(n12418), .dinb(n12410), .dout(n12512));
  jor  g12257(.dina(n12512), .dinb(n12511), .dout(n12513));
  jand g12258(.dina(n12382), .dinb(n12300), .dout(n12514));
  jand g12259(.dina(n12391), .dinb(n12383), .dout(n12515));
  jor  g12260(.dina(n12515), .dinb(n12514), .dout(n12516));
  jand g12261(.dina(n12372), .dinb(n12303), .dout(n12517));
  jand g12262(.dina(n12381), .dinb(n12373), .dout(n12518));
  jor  g12263(.dina(n12518), .dinb(n12517), .dout(n12519));
  jand g12264(.dina(n12362), .dinb(n12306), .dout(n12520));
  jand g12265(.dina(n12371), .dinb(n12363), .dout(n12521));
  jor  g12266(.dina(n12521), .dinb(n12520), .dout(n12522));
  jand g12267(.dina(n12352), .dinb(n12309), .dout(n12523));
  jand g12268(.dina(n12361), .dinb(n12353), .dout(n12524));
  jor  g12269(.dina(n12524), .dinb(n12523), .dout(n12525));
  jand g12270(.dina(n12342), .dinb(n12312), .dout(n12526));
  jand g12271(.dina(n12351), .dinb(n12343), .dout(n12527));
  jor  g12272(.dina(n12527), .dinb(n12526), .dout(n12528));
  jand g12273(.dina(n12332), .dinb(n12315), .dout(n12529));
  jand g12274(.dina(n12341), .dinb(n12333), .dout(n12530));
  jor  g12275(.dina(n12530), .dinb(n12529), .dout(n12531));
  jand g12276(.dina(n12322), .dinb(n12318), .dout(n12532));
  jand g12277(.dina(n12331), .dinb(n12323), .dout(n12533));
  jor  g12278(.dina(n12533), .dinb(n12532), .dout(n12534));
  jand g12279(.dina(n10594), .dinb(b7 ), .dout(n12535));
  jand g12280(.dina(n10129), .dinb(b8 ), .dout(n12536));
  jor  g12281(.dina(n12536), .dinb(n12535), .dout(n12537));
  jnot g12282(.din(n12537), .dout(n12538));
  jxor g12283(.dina(n12538), .dinb(n12321), .dout(n12539));
  jxor g12284(.dina(n12539), .dinb(n12534), .dout(n12540));
  jor  g12285(.dina(n10134), .dinb(n702), .dout(n12541));
  jor  g12286(.dina(n9849), .dinb(n572), .dout(n12542));
  jor  g12287(.dina(n10132), .dinb(n704), .dout(n12543));
  jor  g12288(.dina(n10137), .dinb(n637), .dout(n12544));
  jand g12289(.dina(n12544), .dinb(n12543), .dout(n12545));
  jand g12290(.dina(n12545), .dinb(n12542), .dout(n12546));
  jand g12291(.dina(n12546), .dinb(n12541), .dout(n12547));
  jxor g12292(.dina(n12547), .dinb(n9559), .dout(n12548));
  jxor g12293(.dina(n12548), .dinb(n12540), .dout(n12549));
  jor  g12294(.dina(n9271), .dinb(n932), .dout(n12550));
  jor  g12295(.dina(n9003), .dinb(n772), .dout(n12551));
  jor  g12296(.dina(n9268), .dinb(n934), .dout(n12552));
  jor  g12297(.dina(n9273), .dinb(n852), .dout(n12553));
  jand g12298(.dina(n12553), .dinb(n12552), .dout(n12554));
  jand g12299(.dina(n12554), .dinb(n12551), .dout(n12555));
  jand g12300(.dina(n12555), .dinb(n12550), .dout(n12556));
  jxor g12301(.dina(n12556), .dinb(n8729), .dout(n12557));
  jxor g12302(.dina(n12557), .dinb(n12549), .dout(n12558));
  jxor g12303(.dina(n12558), .dinb(n12531), .dout(n12559));
  jor  g12304(.dina(n8457), .dinb(n1209), .dout(n12560));
  jor  g12305(.dina(n8185), .dinb(n1018), .dout(n12561));
  jor  g12306(.dina(n8459), .dinb(n1114), .dout(n12562));
  jor  g12307(.dina(n8454), .dinb(n1211), .dout(n12563));
  jand g12308(.dina(n12563), .dinb(n12562), .dout(n12564));
  jand g12309(.dina(n12564), .dinb(n12561), .dout(n12565));
  jand g12310(.dina(n12565), .dinb(n12560), .dout(n12566));
  jxor g12311(.dina(n12566), .dinb(n7929), .dout(n12567));
  jxor g12312(.dina(n12567), .dinb(n12559), .dout(n12568));
  jxor g12313(.dina(n12568), .dinb(n12528), .dout(n12569));
  jor  g12314(.dina(n7660), .dinb(n1525), .dout(n12570));
  jor  g12315(.dina(n7415), .dinb(n1307), .dout(n12571));
  jor  g12316(.dina(n7662), .dinb(n1527), .dout(n12572));
  jor  g12317(.dina(n7657), .dinb(n1416), .dout(n12573));
  jand g12318(.dina(n12573), .dinb(n12572), .dout(n12574));
  jand g12319(.dina(n12574), .dinb(n12571), .dout(n12575));
  jand g12320(.dina(n12575), .dinb(n12570), .dout(n12576));
  jxor g12321(.dina(n12576), .dinb(n7166), .dout(n12577));
  jxor g12322(.dina(n12577), .dinb(n12569), .dout(n12578));
  jxor g12323(.dina(n12578), .dinb(n12525), .dout(n12579));
  jor  g12324(.dina(n6914), .dinb(n1879), .dout(n12580));
  jor  g12325(.dina(n6673), .dinb(n1637), .dout(n12581));
  jor  g12326(.dina(n6916), .dinb(n1881), .dout(n12582));
  jor  g12327(.dina(n6911), .dinb(n1759), .dout(n12583));
  jand g12328(.dina(n12583), .dinb(n12582), .dout(n12584));
  jand g12329(.dina(n12584), .dinb(n12581), .dout(n12585));
  jand g12330(.dina(n12585), .dinb(n12580), .dout(n12586));
  jxor g12331(.dina(n12586), .dinb(n6443), .dout(n12587));
  jxor g12332(.dina(n12587), .dinb(n12579), .dout(n12588));
  jxor g12333(.dina(n12588), .dinb(n12522), .dout(n12589));
  jor  g12334(.dina(n6207), .dinb(n2277), .dout(n12590));
  jor  g12335(.dina(n5975), .dinb(n2007), .dout(n12591));
  jor  g12336(.dina(n6210), .dinb(n2142), .dout(n12592));
  jor  g12337(.dina(n6205), .dinb(n2279), .dout(n12593));
  jand g12338(.dina(n12593), .dinb(n12592), .dout(n12594));
  jand g12339(.dina(n12594), .dinb(n12591), .dout(n12595));
  jand g12340(.dina(n12595), .dinb(n12590), .dout(n12596));
  jxor g12341(.dina(n12596), .dinb(n5759), .dout(n12597));
  jxor g12342(.dina(n12597), .dinb(n12589), .dout(n12598));
  jxor g12343(.dina(n12598), .dinb(n12519), .dout(n12599));
  jor  g12344(.dina(n5537), .dinb(n2711), .dout(n12600));
  jor  g12345(.dina(n5315), .dinb(n2415), .dout(n12601));
  jor  g12346(.dina(n5539), .dinb(n2713), .dout(n12602));
  jor  g12347(.dina(n5534), .dinb(n2563), .dout(n12603));
  jand g12348(.dina(n12603), .dinb(n12602), .dout(n12604));
  jand g12349(.dina(n12604), .dinb(n12601), .dout(n12605));
  jand g12350(.dina(n12605), .dinb(n12600), .dout(n12606));
  jxor g12351(.dina(n12606), .dinb(n5111), .dout(n12607));
  jxor g12352(.dina(n12607), .dinb(n12599), .dout(n12608));
  jxor g12353(.dina(n12608), .dinb(n12516), .dout(n12609));
  jor  g12354(.dina(n4902), .dinb(n3184), .dout(n12610));
  jor  g12355(.dina(n4696), .dinb(n2862), .dout(n12611));
  jor  g12356(.dina(n4904), .dinb(n3023), .dout(n12612));
  jor  g12357(.dina(n4899), .dinb(n3186), .dout(n12613));
  jand g12358(.dina(n12613), .dinb(n12612), .dout(n12614));
  jand g12359(.dina(n12614), .dinb(n12611), .dout(n12615));
  jand g12360(.dina(n12615), .dinb(n12610), .dout(n12616));
  jxor g12361(.dina(n12616), .dinb(n4505), .dout(n12617));
  jxor g12362(.dina(n12617), .dinb(n12609), .dout(n12618));
  jand g12363(.dina(n12392), .dinb(n12297), .dout(n12619));
  jand g12364(.dina(n12401), .dinb(n12393), .dout(n12620));
  jor  g12365(.dina(n12620), .dinb(n12619), .dout(n12621));
  jxor g12366(.dina(n12621), .dinb(n12618), .dout(n12622));
  jor  g12367(.dina(n4305), .dinb(n3696), .dout(n12623));
  jor  g12368(.dina(n4116), .dinb(n3348), .dout(n12624));
  jor  g12369(.dina(n4303), .dinb(n3698), .dout(n12625));
  jor  g12370(.dina(n4308), .dinb(n3522), .dout(n12626));
  jand g12371(.dina(n12626), .dinb(n12625), .dout(n12627));
  jand g12372(.dina(n12627), .dinb(n12624), .dout(n12628));
  jand g12373(.dina(n12628), .dinb(n12623), .dout(n12629));
  jxor g12374(.dina(n12629), .dinb(n3938), .dout(n12630));
  jxor g12375(.dina(n12630), .dinb(n12622), .dout(n12631));
  jxor g12376(.dina(n12631), .dinb(n12513), .dout(n12632));
  jor  g12377(.dina(n4247), .dinb(n3751), .dout(n12633));
  jor  g12378(.dina(n3574), .dinb(n3873), .dout(n12634));
  jor  g12379(.dina(n3754), .dinb(n4060), .dout(n12635));
  jor  g12380(.dina(n3749), .dinb(n4249), .dout(n12636));
  jand g12381(.dina(n12636), .dinb(n12635), .dout(n12637));
  jand g12382(.dina(n12637), .dinb(n12634), .dout(n12638));
  jand g12383(.dina(n12638), .dinb(n12633), .dout(n12639));
  jxor g12384(.dina(n12639), .dinb(n3410), .dout(n12640));
  jxor g12385(.dina(n12640), .dinb(n12632), .dout(n12641));
  jxor g12386(.dina(n12641), .dinb(n12510), .dout(n12642));
  jxor g12387(.dina(n12642), .dinb(n12498), .dout(n12643));
  jand g12388(.dina(n12278), .dinb(n12270), .dout(n12644));
  jand g12389(.dina(n12430), .dinb(n12279), .dout(n12645));
  jor  g12390(.dina(n12645), .dinb(n12644), .dout(n12646));
  jor  g12391(.dina(n6137), .dinb(n2324), .dout(n12647));
  jor  g12392(.dina(n2186), .dinb(n5685), .dout(n12648));
  jor  g12393(.dina(n2321), .dinb(n5911), .dout(n12649));
  jor  g12394(.dina(n2326), .dinb(n6139), .dout(n12650));
  jand g12395(.dina(n12650), .dinb(n12649), .dout(n12651));
  jand g12396(.dina(n12651), .dinb(n12648), .dout(n12652));
  jand g12397(.dina(n12652), .dinb(n12647), .dout(n12653));
  jxor g12398(.dina(n12653), .dinb(n2057), .dout(n12654));
  jxor g12399(.dina(n12654), .dinb(n12646), .dout(n12655));
  jxor g12400(.dina(n12655), .dinb(n12643), .dout(n12656));
  jxor g12401(.dina(n12656), .dinb(n12486), .dout(n12657));
  jand g12402(.dina(n12443), .dinb(n12435), .dout(n12658));
  jand g12403(.dina(n12444), .dinb(n12432), .dout(n12659));
  jor  g12404(.dina(n12659), .dinb(n12658), .dout(n12660));
  jor  g12405(.dina(n7588), .dinb(n1569), .dout(n12661));
  jor  g12406(.dina(n1453), .dinb(n7086), .dout(n12662));
  jor  g12407(.dina(n1571), .dinb(n7590), .dout(n12663));
  jor  g12408(.dina(n1566), .dinb(n7338), .dout(n12664));
  jand g12409(.dina(n12664), .dinb(n12663), .dout(n12665));
  jand g12410(.dina(n12665), .dinb(n12662), .dout(n12666));
  jand g12411(.dina(n12666), .dinb(n12661), .dout(n12667));
  jxor g12412(.dina(n12667), .dinb(n1351), .dout(n12668));
  jxor g12413(.dina(n12668), .dinb(n12660), .dout(n12669));
  jxor g12414(.dina(n12669), .dinb(n12657), .dout(n12670));
  jxor g12415(.dina(n12670), .dinb(n12474), .dout(n12671));
  jand g12416(.dina(n12242), .dinb(n12234), .dout(n12672));
  jand g12417(.dina(n12446), .dinb(n12243), .dout(n12673));
  jor  g12418(.dina(n12673), .dinb(n12672), .dout(n12674));
  jor  g12419(.dina(n9193), .dinb(n970), .dout(n12675));
  jor  g12420(.dina(n880), .dinb(n8644), .dout(n12676));
  jor  g12421(.dina(n967), .dinb(n8920), .dout(n12677));
  jor  g12422(.dina(n972), .dinb(n9195), .dout(n12678));
  jand g12423(.dina(n12678), .dinb(n12677), .dout(n12679));
  jand g12424(.dina(n12679), .dinb(n12676), .dout(n12680));
  jand g12425(.dina(n12680), .dinb(n12675), .dout(n12681));
  jxor g12426(.dina(n12681), .dinb(n810), .dout(n12682));
  jxor g12427(.dina(n12682), .dinb(n12674), .dout(n12683));
  jxor g12428(.dina(n12683), .dinb(n12671), .dout(n12684));
  jand g12429(.dina(n12230), .dinb(n12222), .dout(n12685));
  jand g12430(.dina(n12447), .dinb(n12231), .dout(n12686));
  jor  g12431(.dina(n12686), .dinb(n12685), .dout(n12687));
  jor  g12432(.dina(n10049), .dinb(n728), .dout(n12688));
  jor  g12433(.dina(n660), .dinb(n9475), .dout(n12689));
  jor  g12434(.dina(n731), .dinb(n9759), .dout(n12690));
  jor  g12435(.dina(n726), .dinb(n10051), .dout(n12691));
  jand g12436(.dina(n12691), .dinb(n12690), .dout(n12692));
  jand g12437(.dina(n12692), .dinb(n12689), .dout(n12693));
  jand g12438(.dina(n12693), .dinb(n12688), .dout(n12694));
  jxor g12439(.dina(n12694), .dinb(n606), .dout(n12695));
  jxor g12440(.dina(n12695), .dinb(n12687), .dout(n12696));
  jxor g12441(.dina(n12696), .dinb(n12684), .dout(n12697));
  jand g12442(.dina(n12218), .dinb(n12210), .dout(n12698));
  jand g12443(.dina(n12448), .dinb(n12219), .dout(n12699));
  jor  g12444(.dina(n12699), .dinb(n12698), .dout(n12700));
  jnot g12445(.din(n12700), .dout(n12701));
  jand g12446(.dina(n487), .dinb(b63 ), .dout(n12702));
  jand g12447(.dina(n10832), .dinb(n435), .dout(n12703));
  jor  g12448(.dina(n12703), .dinb(n12702), .dout(n12704));
  jxor g12449(.dina(n12704), .dinb(n446), .dout(n12705));
  jxor g12450(.dina(n12705), .dinb(n12701), .dout(n12706));
  jxor g12451(.dina(n12706), .dinb(n12697), .dout(n12707));
  jxor g12452(.dina(n12707), .dinb(n12462), .dout(n12708));
  jnot g12453(.din(n12708), .dout(n12709));
  jxor g12454(.dina(n12709), .dinb(n12457), .dout(f71 ));
  jand g12455(.dina(n12707), .dinb(n12462), .dout(n12711));
  jnot g12456(.din(n12711), .dout(n12712));
  jor  g12457(.dina(n12709), .dinb(n12457), .dout(n12713));
  jand g12458(.dina(n12713), .dinb(n12712), .dout(n12714));
  jor  g12459(.dina(n12705), .dinb(n12701), .dout(n12715));
  jand g12460(.dina(n12706), .dinb(n12697), .dout(n12716));
  jnot g12461(.din(n12716), .dout(n12717));
  jand g12462(.dina(n12717), .dinb(n12715), .dout(n12718));
  jnot g12463(.din(n12718), .dout(n12719));
  jand g12464(.dina(n12695), .dinb(n12687), .dout(n12720));
  jand g12465(.dina(n12696), .dinb(n12684), .dout(n12721));
  jor  g12466(.dina(n12721), .dinb(n12720), .dout(n12722));
  jor  g12467(.dina(n10521), .dinb(n728), .dout(n12723));
  jor  g12468(.dina(n660), .dinb(n9759), .dout(n12724));
  jor  g12469(.dina(n726), .dinb(n10523), .dout(n12725));
  jor  g12470(.dina(n731), .dinb(n10051), .dout(n12726));
  jand g12471(.dina(n12726), .dinb(n12725), .dout(n12727));
  jand g12472(.dina(n12727), .dinb(n12724), .dout(n12728));
  jand g12473(.dina(n12728), .dinb(n12723), .dout(n12729));
  jxor g12474(.dina(n12729), .dinb(n606), .dout(n12730));
  jxor g12475(.dina(n12730), .dinb(n12722), .dout(n12731));
  jand g12476(.dina(n12682), .dinb(n12674), .dout(n12732));
  jand g12477(.dina(n12683), .dinb(n12671), .dout(n12733));
  jor  g12478(.dina(n12733), .dinb(n12732), .dout(n12734));
  jor  g12479(.dina(n9473), .dinb(n970), .dout(n12735));
  jor  g12480(.dina(n880), .dinb(n8920), .dout(n12736));
  jor  g12481(.dina(n972), .dinb(n9475), .dout(n12737));
  jor  g12482(.dina(n967), .dinb(n9195), .dout(n12738));
  jand g12483(.dina(n12738), .dinb(n12737), .dout(n12739));
  jand g12484(.dina(n12739), .dinb(n12736), .dout(n12740));
  jand g12485(.dina(n12740), .dinb(n12735), .dout(n12741));
  jxor g12486(.dina(n12741), .dinb(n810), .dout(n12742));
  jxor g12487(.dina(n12742), .dinb(n12734), .dout(n12743));
  jand g12488(.dina(n12473), .dinb(n12465), .dout(n12744));
  jand g12489(.dina(n12670), .dinb(n12474), .dout(n12745));
  jor  g12490(.dina(n12745), .dinb(n12744), .dout(n12746));
  jor  g12491(.dina(n8642), .dinb(n1248), .dout(n12747));
  jor  g12492(.dina(n1147), .dinb(n8111), .dout(n12748));
  jor  g12493(.dina(n1251), .dinb(n8378), .dout(n12749));
  jor  g12494(.dina(n1246), .dinb(n8644), .dout(n12750));
  jand g12495(.dina(n12750), .dinb(n12749), .dout(n12751));
  jand g12496(.dina(n12751), .dinb(n12748), .dout(n12752));
  jand g12497(.dina(n12752), .dinb(n12747), .dout(n12753));
  jxor g12498(.dina(n12753), .dinb(n1061), .dout(n12754));
  jxor g12499(.dina(n12754), .dinb(n12746), .dout(n12755));
  jand g12500(.dina(n12485), .dinb(n12477), .dout(n12756));
  jand g12501(.dina(n12656), .dinb(n12486), .dout(n12757));
  jor  g12502(.dina(n12757), .dinb(n12756), .dout(n12758));
  jor  g12503(.dina(n7084), .dinb(n1921), .dout(n12759));
  jor  g12504(.dina(n1806), .dinb(n6605), .dout(n12760));
  jor  g12505(.dina(n1918), .dinb(n6846), .dout(n12761));
  jor  g12506(.dina(n1923), .dinb(n7086), .dout(n12762));
  jand g12507(.dina(n12762), .dinb(n12761), .dout(n12763));
  jand g12508(.dina(n12763), .dinb(n12760), .dout(n12764));
  jand g12509(.dina(n12764), .dinb(n12759), .dout(n12765));
  jxor g12510(.dina(n12765), .dinb(n1687), .dout(n12766));
  jxor g12511(.dina(n12766), .dinb(n12758), .dout(n12767));
  jand g12512(.dina(n12654), .dinb(n12646), .dout(n12768));
  jand g12513(.dina(n12655), .dinb(n12643), .dout(n12769));
  jor  g12514(.dina(n12769), .dinb(n12768), .dout(n12770));
  jor  g12515(.dina(n6364), .dinb(n2324), .dout(n12771));
  jor  g12516(.dina(n2186), .dinb(n5911), .dout(n12772));
  jor  g12517(.dina(n2321), .dinb(n6139), .dout(n12773));
  jor  g12518(.dina(n2326), .dinb(n6366), .dout(n12774));
  jand g12519(.dina(n12774), .dinb(n12773), .dout(n12775));
  jand g12520(.dina(n12775), .dinb(n12772), .dout(n12776));
  jand g12521(.dina(n12776), .dinb(n12771), .dout(n12777));
  jxor g12522(.dina(n12777), .dinb(n2057), .dout(n12778));
  jxor g12523(.dina(n12778), .dinb(n12770), .dout(n12779));
  jand g12524(.dina(n12509), .dinb(n12501), .dout(n12780));
  jand g12525(.dina(n12641), .dinb(n12510), .dout(n12781));
  jor  g12526(.dina(n12781), .dinb(n12780), .dout(n12782));
  jor  g12527(.dina(n5038), .dinb(n3239), .dout(n12783));
  jor  g12528(.dina(n3072), .dinb(n4637), .dout(n12784));
  jor  g12529(.dina(n3242), .dinb(n4839), .dout(n12785));
  jor  g12530(.dina(n3237), .dinb(n5040), .dout(n12786));
  jand g12531(.dina(n12786), .dinb(n12785), .dout(n12787));
  jand g12532(.dina(n12787), .dinb(n12784), .dout(n12788));
  jand g12533(.dina(n12788), .dinb(n12783), .dout(n12789));
  jxor g12534(.dina(n12789), .dinb(n2918), .dout(n12790));
  jxor g12535(.dina(n12790), .dinb(n12782), .dout(n12791));
  jand g12536(.dina(n12631), .dinb(n12513), .dout(n12792));
  jand g12537(.dina(n12640), .dinb(n12632), .dout(n12793));
  jor  g12538(.dina(n12793), .dinb(n12792), .dout(n12794));
  jand g12539(.dina(n12621), .dinb(n12618), .dout(n12795));
  jand g12540(.dina(n12630), .dinb(n12622), .dout(n12796));
  jor  g12541(.dina(n12796), .dinb(n12795), .dout(n12797));
  jand g12542(.dina(n12608), .dinb(n12516), .dout(n12798));
  jand g12543(.dina(n12617), .dinb(n12609), .dout(n12799));
  jor  g12544(.dina(n12799), .dinb(n12798), .dout(n12800));
  jor  g12545(.dina(n4902), .dinb(n3346), .dout(n12801));
  jor  g12546(.dina(n4696), .dinb(n3023), .dout(n12802));
  jor  g12547(.dina(n4899), .dinb(n3348), .dout(n12803));
  jor  g12548(.dina(n4904), .dinb(n3186), .dout(n12804));
  jand g12549(.dina(n12804), .dinb(n12803), .dout(n12805));
  jand g12550(.dina(n12805), .dinb(n12802), .dout(n12806));
  jand g12551(.dina(n12806), .dinb(n12801), .dout(n12807));
  jxor g12552(.dina(n12807), .dinb(n4505), .dout(n12808));
  jand g12553(.dina(n12598), .dinb(n12519), .dout(n12809));
  jand g12554(.dina(n12607), .dinb(n12599), .dout(n12810));
  jor  g12555(.dina(n12810), .dinb(n12809), .dout(n12811));
  jand g12556(.dina(n12588), .dinb(n12522), .dout(n12812));
  jand g12557(.dina(n12597), .dinb(n12589), .dout(n12813));
  jor  g12558(.dina(n12813), .dinb(n12812), .dout(n12814));
  jand g12559(.dina(n12578), .dinb(n12525), .dout(n12815));
  jand g12560(.dina(n12587), .dinb(n12579), .dout(n12816));
  jor  g12561(.dina(n12816), .dinb(n12815), .dout(n12817));
  jand g12562(.dina(n12568), .dinb(n12528), .dout(n12818));
  jand g12563(.dina(n12577), .dinb(n12569), .dout(n12819));
  jor  g12564(.dina(n12819), .dinb(n12818), .dout(n12820));
  jand g12565(.dina(n12558), .dinb(n12531), .dout(n12821));
  jand g12566(.dina(n12567), .dinb(n12559), .dout(n12822));
  jor  g12567(.dina(n12822), .dinb(n12821), .dout(n12823));
  jand g12568(.dina(n12548), .dinb(n12540), .dout(n12824));
  jand g12569(.dina(n12557), .dinb(n12549), .dout(n12825));
  jor  g12570(.dina(n12825), .dinb(n12824), .dout(n12826));
  jand g12571(.dina(n12538), .dinb(n12321), .dout(n12827));
  jand g12572(.dina(n12539), .dinb(n12534), .dout(n12828));
  jor  g12573(.dina(n12828), .dinb(n12827), .dout(n12829));
  jand g12574(.dina(n10594), .dinb(b8 ), .dout(n12830));
  jand g12575(.dina(n10129), .dinb(b9 ), .dout(n12831));
  jor  g12576(.dina(n12831), .dinb(n12830), .dout(n12832));
  jxor g12577(.dina(n12537), .dinb(n446), .dout(n12833));
  jxor g12578(.dina(n12833), .dinb(n12832), .dout(n12834));
  jxor g12579(.dina(n12834), .dinb(n12829), .dout(n12835));
  jor  g12580(.dina(n10134), .dinb(n770), .dout(n12836));
  jor  g12581(.dina(n9849), .dinb(n637), .dout(n12837));
  jor  g12582(.dina(n10137), .dinb(n704), .dout(n12838));
  jor  g12583(.dina(n10132), .dinb(n772), .dout(n12839));
  jand g12584(.dina(n12839), .dinb(n12838), .dout(n12840));
  jand g12585(.dina(n12840), .dinb(n12837), .dout(n12841));
  jand g12586(.dina(n12841), .dinb(n12836), .dout(n12842));
  jxor g12587(.dina(n12842), .dinb(n9559), .dout(n12843));
  jxor g12588(.dina(n12843), .dinb(n12835), .dout(n12844));
  jor  g12589(.dina(n9271), .dinb(n1016), .dout(n12845));
  jor  g12590(.dina(n9003), .dinb(n852), .dout(n12846));
  jor  g12591(.dina(n9268), .dinb(n1018), .dout(n12847));
  jor  g12592(.dina(n9273), .dinb(n934), .dout(n12848));
  jand g12593(.dina(n12848), .dinb(n12847), .dout(n12849));
  jand g12594(.dina(n12849), .dinb(n12846), .dout(n12850));
  jand g12595(.dina(n12850), .dinb(n12845), .dout(n12851));
  jxor g12596(.dina(n12851), .dinb(n8729), .dout(n12852));
  jxor g12597(.dina(n12852), .dinb(n12844), .dout(n12853));
  jxor g12598(.dina(n12853), .dinb(n12826), .dout(n12854));
  jor  g12599(.dina(n8457), .dinb(n1305), .dout(n12855));
  jor  g12600(.dina(n8185), .dinb(n1114), .dout(n12856));
  jor  g12601(.dina(n8454), .dinb(n1307), .dout(n12857));
  jor  g12602(.dina(n8459), .dinb(n1211), .dout(n12858));
  jand g12603(.dina(n12858), .dinb(n12857), .dout(n12859));
  jand g12604(.dina(n12859), .dinb(n12856), .dout(n12860));
  jand g12605(.dina(n12860), .dinb(n12855), .dout(n12861));
  jxor g12606(.dina(n12861), .dinb(n7929), .dout(n12862));
  jxor g12607(.dina(n12862), .dinb(n12854), .dout(n12863));
  jxor g12608(.dina(n12863), .dinb(n12823), .dout(n12864));
  jor  g12609(.dina(n7660), .dinb(n1635), .dout(n12865));
  jor  g12610(.dina(n7415), .dinb(n1416), .dout(n12866));
  jor  g12611(.dina(n7662), .dinb(n1637), .dout(n12867));
  jor  g12612(.dina(n7657), .dinb(n1527), .dout(n12868));
  jand g12613(.dina(n12868), .dinb(n12867), .dout(n12869));
  jand g12614(.dina(n12869), .dinb(n12866), .dout(n12870));
  jand g12615(.dina(n12870), .dinb(n12865), .dout(n12871));
  jxor g12616(.dina(n12871), .dinb(n7166), .dout(n12872));
  jxor g12617(.dina(n12872), .dinb(n12864), .dout(n12873));
  jxor g12618(.dina(n12873), .dinb(n12820), .dout(n12874));
  jor  g12619(.dina(n6914), .dinb(n2005), .dout(n12875));
  jor  g12620(.dina(n6673), .dinb(n1759), .dout(n12876));
  jor  g12621(.dina(n6911), .dinb(n1881), .dout(n12877));
  jor  g12622(.dina(n6916), .dinb(n2007), .dout(n12878));
  jand g12623(.dina(n12878), .dinb(n12877), .dout(n12879));
  jand g12624(.dina(n12879), .dinb(n12876), .dout(n12880));
  jand g12625(.dina(n12880), .dinb(n12875), .dout(n12881));
  jxor g12626(.dina(n12881), .dinb(n6443), .dout(n12882));
  jxor g12627(.dina(n12882), .dinb(n12874), .dout(n12883));
  jxor g12628(.dina(n12883), .dinb(n12817), .dout(n12884));
  jor  g12629(.dina(n6207), .dinb(n2413), .dout(n12885));
  jor  g12630(.dina(n5975), .dinb(n2142), .dout(n12886));
  jor  g12631(.dina(n6205), .dinb(n2415), .dout(n12887));
  jor  g12632(.dina(n6210), .dinb(n2279), .dout(n12888));
  jand g12633(.dina(n12888), .dinb(n12887), .dout(n12889));
  jand g12634(.dina(n12889), .dinb(n12886), .dout(n12890));
  jand g12635(.dina(n12890), .dinb(n12885), .dout(n12891));
  jxor g12636(.dina(n12891), .dinb(n5759), .dout(n12892));
  jxor g12637(.dina(n12892), .dinb(n12884), .dout(n12893));
  jxor g12638(.dina(n12893), .dinb(n12814), .dout(n12894));
  jor  g12639(.dina(n5537), .dinb(n2860), .dout(n12895));
  jor  g12640(.dina(n5315), .dinb(n2563), .dout(n12896));
  jor  g12641(.dina(n5534), .dinb(n2713), .dout(n12897));
  jor  g12642(.dina(n5539), .dinb(n2862), .dout(n12898));
  jand g12643(.dina(n12898), .dinb(n12897), .dout(n12899));
  jand g12644(.dina(n12899), .dinb(n12896), .dout(n12900));
  jand g12645(.dina(n12900), .dinb(n12895), .dout(n12901));
  jxor g12646(.dina(n12901), .dinb(n5111), .dout(n12902));
  jxor g12647(.dina(n12902), .dinb(n12894), .dout(n12903));
  jxor g12648(.dina(n12903), .dinb(n12811), .dout(n12904));
  jxor g12649(.dina(n12904), .dinb(n12808), .dout(n12905));
  jxor g12650(.dina(n12905), .dinb(n12800), .dout(n12906));
  jor  g12651(.dina(n4305), .dinb(n3871), .dout(n12907));
  jor  g12652(.dina(n4116), .dinb(n3522), .dout(n12908));
  jor  g12653(.dina(n4308), .dinb(n3698), .dout(n12909));
  jor  g12654(.dina(n4303), .dinb(n3873), .dout(n12910));
  jand g12655(.dina(n12910), .dinb(n12909), .dout(n12911));
  jand g12656(.dina(n12911), .dinb(n12908), .dout(n12912));
  jand g12657(.dina(n12912), .dinb(n12907), .dout(n12913));
  jxor g12658(.dina(n12913), .dinb(n3938), .dout(n12914));
  jxor g12659(.dina(n12914), .dinb(n12906), .dout(n12915));
  jxor g12660(.dina(n12915), .dinb(n12797), .dout(n12916));
  jor  g12661(.dina(n4435), .dinb(n3751), .dout(n12917));
  jor  g12662(.dina(n3574), .dinb(n4060), .dout(n12918));
  jor  g12663(.dina(n3754), .dinb(n4249), .dout(n12919));
  jor  g12664(.dina(n3749), .dinb(n4437), .dout(n12920));
  jand g12665(.dina(n12920), .dinb(n12919), .dout(n12921));
  jand g12666(.dina(n12921), .dinb(n12918), .dout(n12922));
  jand g12667(.dina(n12922), .dinb(n12917), .dout(n12923));
  jxor g12668(.dina(n12923), .dinb(n3410), .dout(n12924));
  jxor g12669(.dina(n12924), .dinb(n12916), .dout(n12925));
  jxor g12670(.dina(n12925), .dinb(n12794), .dout(n12926));
  jxor g12671(.dina(n12926), .dinb(n12791), .dout(n12927));
  jand g12672(.dina(n12497), .dinb(n12489), .dout(n12928));
  jand g12673(.dina(n12642), .dinb(n12498), .dout(n12929));
  jor  g12674(.dina(n12929), .dinb(n12928), .dout(n12930));
  jor  g12675(.dina(n5683), .dinb(n2764), .dout(n12931));
  jor  g12676(.dina(n2609), .dinb(n5253), .dout(n12932));
  jor  g12677(.dina(n2761), .dinb(n5685), .dout(n12933));
  jor  g12678(.dina(n2766), .dinb(n5469), .dout(n12934));
  jand g12679(.dina(n12934), .dinb(n12933), .dout(n12935));
  jand g12680(.dina(n12935), .dinb(n12932), .dout(n12936));
  jand g12681(.dina(n12936), .dinb(n12931), .dout(n12937));
  jxor g12682(.dina(n12937), .dinb(n2468), .dout(n12938));
  jxor g12683(.dina(n12938), .dinb(n12930), .dout(n12939));
  jxor g12684(.dina(n12939), .dinb(n12927), .dout(n12940));
  jxor g12685(.dina(n12940), .dinb(n12779), .dout(n12941));
  jxor g12686(.dina(n12941), .dinb(n12767), .dout(n12942));
  jand g12687(.dina(n12668), .dinb(n12660), .dout(n12943));
  jand g12688(.dina(n12669), .dinb(n12657), .dout(n12944));
  jor  g12689(.dina(n12944), .dinb(n12943), .dout(n12945));
  jor  g12690(.dina(n7844), .dinb(n1569), .dout(n12946));
  jor  g12691(.dina(n1453), .dinb(n7338), .dout(n12947));
  jor  g12692(.dina(n1566), .dinb(n7590), .dout(n12948));
  jor  g12693(.dina(n1571), .dinb(n7846), .dout(n12949));
  jand g12694(.dina(n12949), .dinb(n12948), .dout(n12950));
  jand g12695(.dina(n12950), .dinb(n12947), .dout(n12951));
  jand g12696(.dina(n12951), .dinb(n12946), .dout(n12952));
  jxor g12697(.dina(n12952), .dinb(n1351), .dout(n12953));
  jxor g12698(.dina(n12953), .dinb(n12945), .dout(n12954));
  jxor g12699(.dina(n12954), .dinb(n12942), .dout(n12955));
  jxor g12700(.dina(n12955), .dinb(n12755), .dout(n12956));
  jxor g12701(.dina(n12956), .dinb(n12743), .dout(n12957));
  jxor g12702(.dina(n12957), .dinb(n12731), .dout(n12958));
  jxor g12703(.dina(n12958), .dinb(n12719), .dout(n12959));
  jnot g12704(.din(n12959), .dout(n12960));
  jxor g12705(.dina(n12960), .dinb(n12714), .dout(f72 ));
  jand g12706(.dina(n12958), .dinb(n12719), .dout(n12962));
  jnot g12707(.din(n12962), .dout(n12963));
  jor  g12708(.dina(n12960), .dinb(n12714), .dout(n12964));
  jand g12709(.dina(n12964), .dinb(n12963), .dout(n12965));
  jand g12710(.dina(n12730), .dinb(n12722), .dout(n12966));
  jand g12711(.dina(n12957), .dinb(n12731), .dout(n12967));
  jor  g12712(.dina(n12967), .dinb(n12966), .dout(n12968));
  jand g12713(.dina(n12754), .dinb(n12746), .dout(n12969));
  jand g12714(.dina(n12955), .dinb(n12755), .dout(n12970));
  jor  g12715(.dina(n12970), .dinb(n12969), .dout(n12971));
  jor  g12716(.dina(n9757), .dinb(n970), .dout(n12972));
  jor  g12717(.dina(n880), .dinb(n9195), .dout(n12973));
  jor  g12718(.dina(n967), .dinb(n9475), .dout(n12974));
  jor  g12719(.dina(n972), .dinb(n9759), .dout(n12975));
  jand g12720(.dina(n12975), .dinb(n12974), .dout(n12976));
  jand g12721(.dina(n12976), .dinb(n12973), .dout(n12977));
  jand g12722(.dina(n12977), .dinb(n12972), .dout(n12978));
  jxor g12723(.dina(n12978), .dinb(n810), .dout(n12979));
  jxor g12724(.dina(n12979), .dinb(n12971), .dout(n12980));
  jand g12725(.dina(n12766), .dinb(n12758), .dout(n12981));
  jand g12726(.dina(n12941), .dinb(n12767), .dout(n12982));
  jor  g12727(.dina(n12982), .dinb(n12981), .dout(n12983));
  jor  g12728(.dina(n8109), .dinb(n1569), .dout(n12984));
  jor  g12729(.dina(n1453), .dinb(n7590), .dout(n12985));
  jor  g12730(.dina(n1571), .dinb(n8111), .dout(n12986));
  jor  g12731(.dina(n1566), .dinb(n7846), .dout(n12987));
  jand g12732(.dina(n12987), .dinb(n12986), .dout(n12988));
  jand g12733(.dina(n12988), .dinb(n12985), .dout(n12989));
  jand g12734(.dina(n12989), .dinb(n12984), .dout(n12990));
  jxor g12735(.dina(n12990), .dinb(n1351), .dout(n12991));
  jxor g12736(.dina(n12991), .dinb(n12983), .dout(n12992));
  jand g12737(.dina(n12778), .dinb(n12770), .dout(n12993));
  jand g12738(.dina(n12940), .dinb(n12779), .dout(n12994));
  jor  g12739(.dina(n12994), .dinb(n12993), .dout(n12995));
  jor  g12740(.dina(n7336), .dinb(n1921), .dout(n12996));
  jor  g12741(.dina(n1806), .dinb(n6846), .dout(n12997));
  jor  g12742(.dina(n1923), .dinb(n7338), .dout(n12998));
  jor  g12743(.dina(n1918), .dinb(n7086), .dout(n12999));
  jand g12744(.dina(n12999), .dinb(n12998), .dout(n13000));
  jand g12745(.dina(n13000), .dinb(n12997), .dout(n13001));
  jand g12746(.dina(n13001), .dinb(n12996), .dout(n13002));
  jxor g12747(.dina(n13002), .dinb(n1687), .dout(n13003));
  jxor g12748(.dina(n13003), .dinb(n12995), .dout(n13004));
  jand g12749(.dina(n12938), .dinb(n12930), .dout(n13005));
  jand g12750(.dina(n12939), .dinb(n12927), .dout(n13006));
  jor  g12751(.dina(n13006), .dinb(n13005), .dout(n13007));
  jor  g12752(.dina(n6603), .dinb(n2324), .dout(n13008));
  jor  g12753(.dina(n2186), .dinb(n6139), .dout(n13009));
  jor  g12754(.dina(n2326), .dinb(n6605), .dout(n13010));
  jor  g12755(.dina(n2321), .dinb(n6366), .dout(n13011));
  jand g12756(.dina(n13011), .dinb(n13010), .dout(n13012));
  jand g12757(.dina(n13012), .dinb(n13009), .dout(n13013));
  jand g12758(.dina(n13013), .dinb(n13008), .dout(n13014));
  jxor g12759(.dina(n13014), .dinb(n2057), .dout(n13015));
  jxor g12760(.dina(n13015), .dinb(n13007), .dout(n13016));
  jand g12761(.dina(n12924), .dinb(n12916), .dout(n13017));
  jand g12762(.dina(n12925), .dinb(n12794), .dout(n13018));
  jor  g12763(.dina(n13018), .dinb(n13017), .dout(n13019));
  jor  g12764(.dina(n5251), .dinb(n3239), .dout(n13020));
  jor  g12765(.dina(n3072), .dinb(n4839), .dout(n13021));
  jor  g12766(.dina(n3242), .dinb(n5040), .dout(n13022));
  jor  g12767(.dina(n3237), .dinb(n5253), .dout(n13023));
  jand g12768(.dina(n13023), .dinb(n13022), .dout(n13024));
  jand g12769(.dina(n13024), .dinb(n13021), .dout(n13025));
  jand g12770(.dina(n13025), .dinb(n13020), .dout(n13026));
  jxor g12771(.dina(n13026), .dinb(n2918), .dout(n13027));
  jxor g12772(.dina(n13027), .dinb(n13019), .dout(n13028));
  jand g12773(.dina(n12914), .dinb(n12906), .dout(n13029));
  jand g12774(.dina(n12915), .dinb(n12797), .dout(n13030));
  jor  g12775(.dina(n13030), .dinb(n13029), .dout(n13031));
  jand g12776(.dina(n12904), .dinb(n12808), .dout(n13032));
  jand g12777(.dina(n12905), .dinb(n12800), .dout(n13033));
  jor  g12778(.dina(n13033), .dinb(n13032), .dout(n13034));
  jand g12779(.dina(n12892), .dinb(n12884), .dout(n13035));
  jand g12780(.dina(n12893), .dinb(n12814), .dout(n13036));
  jor  g12781(.dina(n13036), .dinb(n13035), .dout(n13037));
  jand g12782(.dina(n12882), .dinb(n12874), .dout(n13038));
  jand g12783(.dina(n12883), .dinb(n12817), .dout(n13039));
  jor  g12784(.dina(n13039), .dinb(n13038), .dout(n13040));
  jand g12785(.dina(n12872), .dinb(n12864), .dout(n13041));
  jand g12786(.dina(n12873), .dinb(n12820), .dout(n13042));
  jor  g12787(.dina(n13042), .dinb(n13041), .dout(n13043));
  jand g12788(.dina(n12862), .dinb(n12854), .dout(n13044));
  jand g12789(.dina(n12863), .dinb(n12823), .dout(n13045));
  jor  g12790(.dina(n13045), .dinb(n13044), .dout(n13046));
  jand g12791(.dina(n12852), .dinb(n12844), .dout(n13047));
  jand g12792(.dina(n12853), .dinb(n12826), .dout(n13048));
  jor  g12793(.dina(n13048), .dinb(n13047), .dout(n13049));
  jand g12794(.dina(n12834), .dinb(n12829), .dout(n13050));
  jand g12795(.dina(n12843), .dinb(n12835), .dout(n13051));
  jor  g12796(.dina(n13051), .dinb(n13050), .dout(n13052));
  jand g12797(.dina(n10594), .dinb(b9 ), .dout(n13053));
  jand g12798(.dina(n10129), .dinb(b10 ), .dout(n13054));
  jor  g12799(.dina(n13054), .dinb(n13053), .dout(n13055));
  jnot g12800(.din(n13055), .dout(n13056));
  jand g12801(.dina(n12537), .dinb(n446), .dout(n13057));
  jand g12802(.dina(n12833), .dinb(n12832), .dout(n13058));
  jor  g12803(.dina(n13058), .dinb(n13057), .dout(n13059));
  jxor g12804(.dina(n13059), .dinb(n13056), .dout(n13060));
  jor  g12805(.dina(n10134), .dinb(n850), .dout(n13061));
  jor  g12806(.dina(n9849), .dinb(n704), .dout(n13062));
  jor  g12807(.dina(n10137), .dinb(n772), .dout(n13063));
  jor  g12808(.dina(n10132), .dinb(n852), .dout(n13064));
  jand g12809(.dina(n13064), .dinb(n13063), .dout(n13065));
  jand g12810(.dina(n13065), .dinb(n13062), .dout(n13066));
  jand g12811(.dina(n13066), .dinb(n13061), .dout(n13067));
  jxor g12812(.dina(n13067), .dinb(n9559), .dout(n13068));
  jxor g12813(.dina(n13068), .dinb(n13060), .dout(n13069));
  jxor g12814(.dina(n13069), .dinb(n13052), .dout(n13070));
  jor  g12815(.dina(n9271), .dinb(n1112), .dout(n13071));
  jor  g12816(.dina(n9003), .dinb(n934), .dout(n13072));
  jor  g12817(.dina(n9268), .dinb(n1114), .dout(n13073));
  jor  g12818(.dina(n9273), .dinb(n1018), .dout(n13074));
  jand g12819(.dina(n13074), .dinb(n13073), .dout(n13075));
  jand g12820(.dina(n13075), .dinb(n13072), .dout(n13076));
  jand g12821(.dina(n13076), .dinb(n13071), .dout(n13077));
  jxor g12822(.dina(n13077), .dinb(n8729), .dout(n13078));
  jxor g12823(.dina(n13078), .dinb(n13070), .dout(n13079));
  jxor g12824(.dina(n13079), .dinb(n13049), .dout(n13080));
  jor  g12825(.dina(n8457), .dinb(n1414), .dout(n13081));
  jor  g12826(.dina(n8185), .dinb(n1211), .dout(n13082));
  jor  g12827(.dina(n8454), .dinb(n1416), .dout(n13083));
  jor  g12828(.dina(n8459), .dinb(n1307), .dout(n13084));
  jand g12829(.dina(n13084), .dinb(n13083), .dout(n13085));
  jand g12830(.dina(n13085), .dinb(n13082), .dout(n13086));
  jand g12831(.dina(n13086), .dinb(n13081), .dout(n13087));
  jxor g12832(.dina(n13087), .dinb(n7929), .dout(n13088));
  jxor g12833(.dina(n13088), .dinb(n13080), .dout(n13089));
  jxor g12834(.dina(n13089), .dinb(n13046), .dout(n13090));
  jor  g12835(.dina(n7660), .dinb(n1757), .dout(n13091));
  jor  g12836(.dina(n7415), .dinb(n1527), .dout(n13092));
  jor  g12837(.dina(n7662), .dinb(n1759), .dout(n13093));
  jor  g12838(.dina(n7657), .dinb(n1637), .dout(n13094));
  jand g12839(.dina(n13094), .dinb(n13093), .dout(n13095));
  jand g12840(.dina(n13095), .dinb(n13092), .dout(n13096));
  jand g12841(.dina(n13096), .dinb(n13091), .dout(n13097));
  jxor g12842(.dina(n13097), .dinb(n7166), .dout(n13098));
  jxor g12843(.dina(n13098), .dinb(n13090), .dout(n13099));
  jxor g12844(.dina(n13099), .dinb(n13043), .dout(n13100));
  jor  g12845(.dina(n6914), .dinb(n2140), .dout(n13101));
  jor  g12846(.dina(n6673), .dinb(n1881), .dout(n13102));
  jor  g12847(.dina(n6916), .dinb(n2142), .dout(n13103));
  jor  g12848(.dina(n6911), .dinb(n2007), .dout(n13104));
  jand g12849(.dina(n13104), .dinb(n13103), .dout(n13105));
  jand g12850(.dina(n13105), .dinb(n13102), .dout(n13106));
  jand g12851(.dina(n13106), .dinb(n13101), .dout(n13107));
  jxor g12852(.dina(n13107), .dinb(n6443), .dout(n13108));
  jxor g12853(.dina(n13108), .dinb(n13100), .dout(n13109));
  jxor g12854(.dina(n13109), .dinb(n13040), .dout(n13110));
  jor  g12855(.dina(n6207), .dinb(n2561), .dout(n13111));
  jor  g12856(.dina(n5975), .dinb(n2279), .dout(n13112));
  jor  g12857(.dina(n6210), .dinb(n2415), .dout(n13113));
  jor  g12858(.dina(n6205), .dinb(n2563), .dout(n13114));
  jand g12859(.dina(n13114), .dinb(n13113), .dout(n13115));
  jand g12860(.dina(n13115), .dinb(n13112), .dout(n13116));
  jand g12861(.dina(n13116), .dinb(n13111), .dout(n13117));
  jxor g12862(.dina(n13117), .dinb(n5759), .dout(n13118));
  jxor g12863(.dina(n13118), .dinb(n13110), .dout(n13119));
  jxor g12864(.dina(n13119), .dinb(n13037), .dout(n13120));
  jor  g12865(.dina(n5537), .dinb(n3021), .dout(n13121));
  jor  g12866(.dina(n5315), .dinb(n2713), .dout(n13122));
  jor  g12867(.dina(n5539), .dinb(n3023), .dout(n13123));
  jor  g12868(.dina(n5534), .dinb(n2862), .dout(n13124));
  jand g12869(.dina(n13124), .dinb(n13123), .dout(n13125));
  jand g12870(.dina(n13125), .dinb(n13122), .dout(n13126));
  jand g12871(.dina(n13126), .dinb(n13121), .dout(n13127));
  jxor g12872(.dina(n13127), .dinb(n5111), .dout(n13128));
  jxor g12873(.dina(n13128), .dinb(n13120), .dout(n13129));
  jnot g12874(.din(n12894), .dout(n13130));
  jnot g12875(.din(n12902), .dout(n13131));
  jand g12876(.dina(n13131), .dinb(n13130), .dout(n13132));
  jnot g12877(.din(n13132), .dout(n13133));
  jand g12878(.dina(n12902), .dinb(n12894), .dout(n13134));
  jor  g12879(.dina(n13134), .dinb(n12811), .dout(n13135));
  jand g12880(.dina(n13135), .dinb(n13133), .dout(n13136));
  jxor g12881(.dina(n13136), .dinb(n13129), .dout(n13137));
  jor  g12882(.dina(n4902), .dinb(n3520), .dout(n13138));
  jor  g12883(.dina(n4696), .dinb(n3186), .dout(n13139));
  jor  g12884(.dina(n4899), .dinb(n3522), .dout(n13140));
  jor  g12885(.dina(n4904), .dinb(n3348), .dout(n13141));
  jand g12886(.dina(n13141), .dinb(n13140), .dout(n13142));
  jand g12887(.dina(n13142), .dinb(n13139), .dout(n13143));
  jand g12888(.dina(n13143), .dinb(n13138), .dout(n13144));
  jxor g12889(.dina(n13144), .dinb(n4505), .dout(n13145));
  jxor g12890(.dina(n13145), .dinb(n13137), .dout(n13146));
  jxor g12891(.dina(n13146), .dinb(n13034), .dout(n13147));
  jor  g12892(.dina(n4058), .dinb(n4305), .dout(n13148));
  jor  g12893(.dina(n4116), .dinb(n3698), .dout(n13149));
  jor  g12894(.dina(n4308), .dinb(n3873), .dout(n13150));
  jor  g12895(.dina(n4303), .dinb(n4060), .dout(n13151));
  jand g12896(.dina(n13151), .dinb(n13150), .dout(n13152));
  jand g12897(.dina(n13152), .dinb(n13149), .dout(n13153));
  jand g12898(.dina(n13153), .dinb(n13148), .dout(n13154));
  jxor g12899(.dina(n13154), .dinb(n3938), .dout(n13155));
  jxor g12900(.dina(n13155), .dinb(n13147), .dout(n13156));
  jxor g12901(.dina(n13156), .dinb(n13031), .dout(n13157));
  jor  g12902(.dina(n4635), .dinb(n3751), .dout(n13158));
  jor  g12903(.dina(n3574), .dinb(n4249), .dout(n13159));
  jor  g12904(.dina(n3749), .dinb(n4637), .dout(n13160));
  jor  g12905(.dina(n3754), .dinb(n4437), .dout(n13161));
  jand g12906(.dina(n13161), .dinb(n13160), .dout(n13162));
  jand g12907(.dina(n13162), .dinb(n13159), .dout(n13163));
  jand g12908(.dina(n13163), .dinb(n13158), .dout(n13164));
  jxor g12909(.dina(n13164), .dinb(n3410), .dout(n13165));
  jxor g12910(.dina(n13165), .dinb(n13157), .dout(n13166));
  jxor g12911(.dina(n13166), .dinb(n13028), .dout(n13167));
  jand g12912(.dina(n12790), .dinb(n12782), .dout(n13168));
  jand g12913(.dina(n12926), .dinb(n12791), .dout(n13169));
  jor  g12914(.dina(n13169), .dinb(n13168), .dout(n13170));
  jor  g12915(.dina(n5909), .dinb(n2764), .dout(n13171));
  jor  g12916(.dina(n2609), .dinb(n5469), .dout(n13172));
  jor  g12917(.dina(n2761), .dinb(n5911), .dout(n13173));
  jor  g12918(.dina(n2766), .dinb(n5685), .dout(n13174));
  jand g12919(.dina(n13174), .dinb(n13173), .dout(n13175));
  jand g12920(.dina(n13175), .dinb(n13172), .dout(n13176));
  jand g12921(.dina(n13176), .dinb(n13171), .dout(n13177));
  jxor g12922(.dina(n13177), .dinb(n2468), .dout(n13178));
  jxor g12923(.dina(n13178), .dinb(n13170), .dout(n13179));
  jxor g12924(.dina(n13179), .dinb(n13167), .dout(n13180));
  jxor g12925(.dina(n13180), .dinb(n13016), .dout(n13181));
  jxor g12926(.dina(n13181), .dinb(n13004), .dout(n13182));
  jxor g12927(.dina(n13182), .dinb(n12992), .dout(n13183));
  jand g12928(.dina(n12953), .dinb(n12945), .dout(n13184));
  jand g12929(.dina(n12954), .dinb(n12942), .dout(n13185));
  jor  g12930(.dina(n13185), .dinb(n13184), .dout(n13186));
  jor  g12931(.dina(n8918), .dinb(n1248), .dout(n13187));
  jor  g12932(.dina(n1147), .dinb(n8378), .dout(n13188));
  jor  g12933(.dina(n1251), .dinb(n8644), .dout(n13189));
  jor  g12934(.dina(n1246), .dinb(n8920), .dout(n13190));
  jand g12935(.dina(n13190), .dinb(n13189), .dout(n13191));
  jand g12936(.dina(n13191), .dinb(n13188), .dout(n13192));
  jand g12937(.dina(n13192), .dinb(n13187), .dout(n13193));
  jxor g12938(.dina(n13193), .dinb(n1061), .dout(n13194));
  jxor g12939(.dina(n13194), .dinb(n13186), .dout(n13195));
  jxor g12940(.dina(n13195), .dinb(n13183), .dout(n13196));
  jxor g12941(.dina(n13196), .dinb(n12980), .dout(n13197));
  jand g12942(.dina(n12742), .dinb(n12734), .dout(n13198));
  jand g12943(.dina(n12956), .dinb(n12743), .dout(n13199));
  jor  g12944(.dina(n13199), .dinb(n13198), .dout(n13200));
  jor  g12945(.dina(n10813), .dinb(n728), .dout(n13201));
  jor  g12946(.dina(n660), .dinb(n10051), .dout(n13202));
  jor  g12947(.dina(n731), .dinb(n10523), .dout(n13203));
  jand g12948(.dina(n13203), .dinb(n13202), .dout(n13204));
  jand g12949(.dina(n13204), .dinb(n13201), .dout(n13205));
  jxor g12950(.dina(n13205), .dinb(n606), .dout(n13206));
  jxor g12951(.dina(n13206), .dinb(n13200), .dout(n13207));
  jxor g12952(.dina(n13207), .dinb(n13197), .dout(n13208));
  jxor g12953(.dina(n13208), .dinb(n12968), .dout(n13209));
  jnot g12954(.din(n13209), .dout(n13210));
  jxor g12955(.dina(n13210), .dinb(n12965), .dout(f73 ));
  jand g12956(.dina(n13208), .dinb(n12968), .dout(n13212));
  jnot g12957(.din(n13212), .dout(n13213));
  jor  g12958(.dina(n13210), .dinb(n12965), .dout(n13214));
  jand g12959(.dina(n13214), .dinb(n13213), .dout(n13215));
  jand g12960(.dina(n13206), .dinb(n13200), .dout(n13216));
  jand g12961(.dina(n13207), .dinb(n13197), .dout(n13217));
  jor  g12962(.dina(n13217), .dinb(n13216), .dout(n13218));
  jand g12963(.dina(n12979), .dinb(n12971), .dout(n13219));
  jand g12964(.dina(n13196), .dinb(n12980), .dout(n13220));
  jor  g12965(.dina(n13220), .dinb(n13219), .dout(n13221));
  jnot g12966(.din(n13221), .dout(n13222));
  jand g12967(.dina(n661), .dinb(b63 ), .dout(n13223));
  jand g12968(.dina(n10832), .dinb(n595), .dout(n13224));
  jor  g12969(.dina(n13224), .dinb(n13223), .dout(n13225));
  jxor g12970(.dina(n13225), .dinb(n606), .dout(n13226));
  jxor g12971(.dina(n13226), .dinb(n13222), .dout(n13227));
  jand g12972(.dina(n13194), .dinb(n13186), .dout(n13228));
  jand g12973(.dina(n13195), .dinb(n13183), .dout(n13229));
  jor  g12974(.dina(n13229), .dinb(n13228), .dout(n13230));
  jor  g12975(.dina(n10049), .dinb(n970), .dout(n13231));
  jor  g12976(.dina(n880), .dinb(n9475), .dout(n13232));
  jor  g12977(.dina(n967), .dinb(n9759), .dout(n13233));
  jor  g12978(.dina(n972), .dinb(n10051), .dout(n13234));
  jand g12979(.dina(n13234), .dinb(n13233), .dout(n13235));
  jand g12980(.dina(n13235), .dinb(n13232), .dout(n13236));
  jand g12981(.dina(n13236), .dinb(n13231), .dout(n13237));
  jxor g12982(.dina(n13237), .dinb(n810), .dout(n13238));
  jxor g12983(.dina(n13238), .dinb(n13230), .dout(n13239));
  jand g12984(.dina(n12991), .dinb(n12983), .dout(n13240));
  jand g12985(.dina(n13182), .dinb(n12992), .dout(n13241));
  jor  g12986(.dina(n13241), .dinb(n13240), .dout(n13242));
  jor  g12987(.dina(n9193), .dinb(n1248), .dout(n13243));
  jor  g12988(.dina(n1147), .dinb(n8644), .dout(n13244));
  jor  g12989(.dina(n1251), .dinb(n8920), .dout(n13245));
  jor  g12990(.dina(n1246), .dinb(n9195), .dout(n13246));
  jand g12991(.dina(n13246), .dinb(n13245), .dout(n13247));
  jand g12992(.dina(n13247), .dinb(n13244), .dout(n13248));
  jand g12993(.dina(n13248), .dinb(n13243), .dout(n13249));
  jxor g12994(.dina(n13249), .dinb(n1061), .dout(n13250));
  jxor g12995(.dina(n13250), .dinb(n13242), .dout(n13251));
  jand g12996(.dina(n13003), .dinb(n12995), .dout(n13252));
  jand g12997(.dina(n13181), .dinb(n13004), .dout(n13253));
  jor  g12998(.dina(n13253), .dinb(n13252), .dout(n13254));
  jor  g12999(.dina(n8376), .dinb(n1569), .dout(n13255));
  jor  g13000(.dina(n1453), .dinb(n7846), .dout(n13256));
  jor  g13001(.dina(n1566), .dinb(n8111), .dout(n13257));
  jor  g13002(.dina(n1571), .dinb(n8378), .dout(n13258));
  jand g13003(.dina(n13258), .dinb(n13257), .dout(n13259));
  jand g13004(.dina(n13259), .dinb(n13256), .dout(n13260));
  jand g13005(.dina(n13260), .dinb(n13255), .dout(n13261));
  jxor g13006(.dina(n13261), .dinb(n1351), .dout(n13262));
  jxor g13007(.dina(n13262), .dinb(n13254), .dout(n13263));
  jand g13008(.dina(n13178), .dinb(n13170), .dout(n13264));
  jand g13009(.dina(n13179), .dinb(n13167), .dout(n13265));
  jor  g13010(.dina(n13265), .dinb(n13264), .dout(n13266));
  jor  g13011(.dina(n6844), .dinb(n2324), .dout(n13267));
  jor  g13012(.dina(n2186), .dinb(n6366), .dout(n13268));
  jor  g13013(.dina(n2321), .dinb(n6605), .dout(n13269));
  jor  g13014(.dina(n2326), .dinb(n6846), .dout(n13270));
  jand g13015(.dina(n13270), .dinb(n13269), .dout(n13271));
  jand g13016(.dina(n13271), .dinb(n13268), .dout(n13272));
  jand g13017(.dina(n13272), .dinb(n13267), .dout(n13273));
  jxor g13018(.dina(n13273), .dinb(n2057), .dout(n13274));
  jxor g13019(.dina(n13274), .dinb(n13266), .dout(n13275));
  jand g13020(.dina(n13027), .dinb(n13019), .dout(n13276));
  jand g13021(.dina(n13166), .dinb(n13028), .dout(n13277));
  jor  g13022(.dina(n13277), .dinb(n13276), .dout(n13278));
  jor  g13023(.dina(n6137), .dinb(n2764), .dout(n13279));
  jor  g13024(.dina(n2609), .dinb(n5685), .dout(n13280));
  jor  g13025(.dina(n2761), .dinb(n6139), .dout(n13281));
  jor  g13026(.dina(n2766), .dinb(n5911), .dout(n13282));
  jand g13027(.dina(n13282), .dinb(n13281), .dout(n13283));
  jand g13028(.dina(n13283), .dinb(n13280), .dout(n13284));
  jand g13029(.dina(n13284), .dinb(n13279), .dout(n13285));
  jxor g13030(.dina(n13285), .dinb(n2468), .dout(n13286));
  jxor g13031(.dina(n13286), .dinb(n13278), .dout(n13287));
  jand g13032(.dina(n13156), .dinb(n13031), .dout(n13288));
  jand g13033(.dina(n13165), .dinb(n13157), .dout(n13289));
  jor  g13034(.dina(n13289), .dinb(n13288), .dout(n13290));
  jor  g13035(.dina(n5467), .dinb(n3239), .dout(n13291));
  jor  g13036(.dina(n3072), .dinb(n5040), .dout(n13292));
  jor  g13037(.dina(n3242), .dinb(n5253), .dout(n13293));
  jor  g13038(.dina(n3237), .dinb(n5469), .dout(n13294));
  jand g13039(.dina(n13294), .dinb(n13293), .dout(n13295));
  jand g13040(.dina(n13295), .dinb(n13292), .dout(n13296));
  jand g13041(.dina(n13296), .dinb(n13291), .dout(n13297));
  jxor g13042(.dina(n13297), .dinb(n2918), .dout(n13298));
  jxor g13043(.dina(n13298), .dinb(n13290), .dout(n13299));
  jand g13044(.dina(n13146), .dinb(n13034), .dout(n13300));
  jand g13045(.dina(n13155), .dinb(n13147), .dout(n13301));
  jor  g13046(.dina(n13301), .dinb(n13300), .dout(n13302));
  jand g13047(.dina(n13136), .dinb(n13129), .dout(n13303));
  jand g13048(.dina(n13145), .dinb(n13137), .dout(n13304));
  jor  g13049(.dina(n13304), .dinb(n13303), .dout(n13305));
  jand g13050(.dina(n13109), .dinb(n13040), .dout(n13306));
  jand g13051(.dina(n13118), .dinb(n13110), .dout(n13307));
  jor  g13052(.dina(n13307), .dinb(n13306), .dout(n13308));
  jand g13053(.dina(n13099), .dinb(n13043), .dout(n13309));
  jand g13054(.dina(n13108), .dinb(n13100), .dout(n13310));
  jor  g13055(.dina(n13310), .dinb(n13309), .dout(n13311));
  jand g13056(.dina(n13089), .dinb(n13046), .dout(n13312));
  jand g13057(.dina(n13098), .dinb(n13090), .dout(n13313));
  jor  g13058(.dina(n13313), .dinb(n13312), .dout(n13314));
  jand g13059(.dina(n13079), .dinb(n13049), .dout(n13315));
  jand g13060(.dina(n13088), .dinb(n13080), .dout(n13316));
  jor  g13061(.dina(n13316), .dinb(n13315), .dout(n13317));
  jand g13062(.dina(n13069), .dinb(n13052), .dout(n13318));
  jand g13063(.dina(n13078), .dinb(n13070), .dout(n13319));
  jor  g13064(.dina(n13319), .dinb(n13318), .dout(n13320));
  jand g13065(.dina(n13059), .dinb(n13056), .dout(n13321));
  jand g13066(.dina(n13068), .dinb(n13060), .dout(n13322));
  jor  g13067(.dina(n13322), .dinb(n13321), .dout(n13323));
  jand g13068(.dina(n10594), .dinb(b10 ), .dout(n13324));
  jand g13069(.dina(n10129), .dinb(b11 ), .dout(n13325));
  jor  g13070(.dina(n13325), .dinb(n13324), .dout(n13326));
  jxor g13071(.dina(n13326), .dinb(n13056), .dout(n13327));
  jxor g13072(.dina(n13327), .dinb(n13323), .dout(n13328));
  jor  g13073(.dina(n10134), .dinb(n932), .dout(n13329));
  jor  g13074(.dina(n9849), .dinb(n772), .dout(n13330));
  jor  g13075(.dina(n10132), .dinb(n934), .dout(n13331));
  jor  g13076(.dina(n10137), .dinb(n852), .dout(n13332));
  jand g13077(.dina(n13332), .dinb(n13331), .dout(n13333));
  jand g13078(.dina(n13333), .dinb(n13330), .dout(n13334));
  jand g13079(.dina(n13334), .dinb(n13329), .dout(n13335));
  jxor g13080(.dina(n13335), .dinb(n9559), .dout(n13336));
  jxor g13081(.dina(n13336), .dinb(n13328), .dout(n13337));
  jor  g13082(.dina(n9271), .dinb(n1209), .dout(n13338));
  jor  g13083(.dina(n9003), .dinb(n1018), .dout(n13339));
  jor  g13084(.dina(n9273), .dinb(n1114), .dout(n13340));
  jor  g13085(.dina(n9268), .dinb(n1211), .dout(n13341));
  jand g13086(.dina(n13341), .dinb(n13340), .dout(n13342));
  jand g13087(.dina(n13342), .dinb(n13339), .dout(n13343));
  jand g13088(.dina(n13343), .dinb(n13338), .dout(n13344));
  jxor g13089(.dina(n13344), .dinb(n8729), .dout(n13345));
  jxor g13090(.dina(n13345), .dinb(n13337), .dout(n13346));
  jxor g13091(.dina(n13346), .dinb(n13320), .dout(n13347));
  jor  g13092(.dina(n8457), .dinb(n1525), .dout(n13348));
  jor  g13093(.dina(n8185), .dinb(n1307), .dout(n13349));
  jor  g13094(.dina(n8459), .dinb(n1416), .dout(n13350));
  jor  g13095(.dina(n8454), .dinb(n1527), .dout(n13351));
  jand g13096(.dina(n13351), .dinb(n13350), .dout(n13352));
  jand g13097(.dina(n13352), .dinb(n13349), .dout(n13353));
  jand g13098(.dina(n13353), .dinb(n13348), .dout(n13354));
  jxor g13099(.dina(n13354), .dinb(n7929), .dout(n13355));
  jxor g13100(.dina(n13355), .dinb(n13347), .dout(n13356));
  jxor g13101(.dina(n13356), .dinb(n13317), .dout(n13357));
  jor  g13102(.dina(n7660), .dinb(n1879), .dout(n13358));
  jor  g13103(.dina(n7415), .dinb(n1637), .dout(n13359));
  jor  g13104(.dina(n7662), .dinb(n1881), .dout(n13360));
  jor  g13105(.dina(n7657), .dinb(n1759), .dout(n13361));
  jand g13106(.dina(n13361), .dinb(n13360), .dout(n13362));
  jand g13107(.dina(n13362), .dinb(n13359), .dout(n13363));
  jand g13108(.dina(n13363), .dinb(n13358), .dout(n13364));
  jxor g13109(.dina(n13364), .dinb(n7166), .dout(n13365));
  jxor g13110(.dina(n13365), .dinb(n13357), .dout(n13366));
  jxor g13111(.dina(n13366), .dinb(n13314), .dout(n13367));
  jor  g13112(.dina(n6914), .dinb(n2277), .dout(n13368));
  jor  g13113(.dina(n6673), .dinb(n2007), .dout(n13369));
  jor  g13114(.dina(n6916), .dinb(n2279), .dout(n13370));
  jor  g13115(.dina(n6911), .dinb(n2142), .dout(n13371));
  jand g13116(.dina(n13371), .dinb(n13370), .dout(n13372));
  jand g13117(.dina(n13372), .dinb(n13369), .dout(n13373));
  jand g13118(.dina(n13373), .dinb(n13368), .dout(n13374));
  jxor g13119(.dina(n13374), .dinb(n6443), .dout(n13375));
  jxor g13120(.dina(n13375), .dinb(n13367), .dout(n13376));
  jxor g13121(.dina(n13376), .dinb(n13311), .dout(n13377));
  jor  g13122(.dina(n6207), .dinb(n2711), .dout(n13378));
  jor  g13123(.dina(n5975), .dinb(n2415), .dout(n13379));
  jor  g13124(.dina(n6210), .dinb(n2563), .dout(n13380));
  jor  g13125(.dina(n6205), .dinb(n2713), .dout(n13381));
  jand g13126(.dina(n13381), .dinb(n13380), .dout(n13382));
  jand g13127(.dina(n13382), .dinb(n13379), .dout(n13383));
  jand g13128(.dina(n13383), .dinb(n13378), .dout(n13384));
  jxor g13129(.dina(n13384), .dinb(n5759), .dout(n13385));
  jxor g13130(.dina(n13385), .dinb(n13377), .dout(n13386));
  jxor g13131(.dina(n13386), .dinb(n13308), .dout(n13387));
  jor  g13132(.dina(n5537), .dinb(n3184), .dout(n13388));
  jor  g13133(.dina(n5315), .dinb(n2862), .dout(n13389));
  jor  g13134(.dina(n5539), .dinb(n3186), .dout(n13390));
  jor  g13135(.dina(n5534), .dinb(n3023), .dout(n13391));
  jand g13136(.dina(n13391), .dinb(n13390), .dout(n13392));
  jand g13137(.dina(n13392), .dinb(n13389), .dout(n13393));
  jand g13138(.dina(n13393), .dinb(n13388), .dout(n13394));
  jxor g13139(.dina(n13394), .dinb(n5111), .dout(n13395));
  jxor g13140(.dina(n13395), .dinb(n13387), .dout(n13396));
  jand g13141(.dina(n13119), .dinb(n13037), .dout(n13397));
  jand g13142(.dina(n13128), .dinb(n13120), .dout(n13398));
  jor  g13143(.dina(n13398), .dinb(n13397), .dout(n13399));
  jxor g13144(.dina(n13399), .dinb(n13396), .dout(n13400));
  jor  g13145(.dina(n4902), .dinb(n3696), .dout(n13401));
  jor  g13146(.dina(n4696), .dinb(n3348), .dout(n13402));
  jor  g13147(.dina(n4904), .dinb(n3522), .dout(n13403));
  jor  g13148(.dina(n4899), .dinb(n3698), .dout(n13404));
  jand g13149(.dina(n13404), .dinb(n13403), .dout(n13405));
  jand g13150(.dina(n13405), .dinb(n13402), .dout(n13406));
  jand g13151(.dina(n13406), .dinb(n13401), .dout(n13407));
  jxor g13152(.dina(n13407), .dinb(n4505), .dout(n13408));
  jxor g13153(.dina(n13408), .dinb(n13400), .dout(n13409));
  jxor g13154(.dina(n13409), .dinb(n13305), .dout(n13410));
  jor  g13155(.dina(n4247), .dinb(n4305), .dout(n13411));
  jor  g13156(.dina(n4116), .dinb(n3873), .dout(n13412));
  jor  g13157(.dina(n4308), .dinb(n4060), .dout(n13413));
  jor  g13158(.dina(n4303), .dinb(n4249), .dout(n13414));
  jand g13159(.dina(n13414), .dinb(n13413), .dout(n13415));
  jand g13160(.dina(n13415), .dinb(n13412), .dout(n13416));
  jand g13161(.dina(n13416), .dinb(n13411), .dout(n13417));
  jxor g13162(.dina(n13417), .dinb(n3938), .dout(n13418));
  jxor g13163(.dina(n13418), .dinb(n13410), .dout(n13419));
  jxor g13164(.dina(n13419), .dinb(n13302), .dout(n13420));
  jor  g13165(.dina(n4837), .dinb(n3751), .dout(n13421));
  jor  g13166(.dina(n3574), .dinb(n4437), .dout(n13422));
  jor  g13167(.dina(n3754), .dinb(n4637), .dout(n13423));
  jor  g13168(.dina(n3749), .dinb(n4839), .dout(n13424));
  jand g13169(.dina(n13424), .dinb(n13423), .dout(n13425));
  jand g13170(.dina(n13425), .dinb(n13422), .dout(n13426));
  jand g13171(.dina(n13426), .dinb(n13421), .dout(n13427));
  jxor g13172(.dina(n13427), .dinb(n3410), .dout(n13428));
  jxor g13173(.dina(n13428), .dinb(n13420), .dout(n13429));
  jxor g13174(.dina(n13429), .dinb(n13299), .dout(n13430));
  jxor g13175(.dina(n13430), .dinb(n13287), .dout(n13431));
  jxor g13176(.dina(n13431), .dinb(n13275), .dout(n13432));
  jand g13177(.dina(n13015), .dinb(n13007), .dout(n13433));
  jand g13178(.dina(n13180), .dinb(n13016), .dout(n13434));
  jor  g13179(.dina(n13434), .dinb(n13433), .dout(n13435));
  jor  g13180(.dina(n7588), .dinb(n1921), .dout(n13436));
  jor  g13181(.dina(n1806), .dinb(n7086), .dout(n13437));
  jor  g13182(.dina(n1923), .dinb(n7590), .dout(n13438));
  jor  g13183(.dina(n1918), .dinb(n7338), .dout(n13439));
  jand g13184(.dina(n13439), .dinb(n13438), .dout(n13440));
  jand g13185(.dina(n13440), .dinb(n13437), .dout(n13441));
  jand g13186(.dina(n13441), .dinb(n13436), .dout(n13442));
  jxor g13187(.dina(n13442), .dinb(n1687), .dout(n13443));
  jxor g13188(.dina(n13443), .dinb(n13435), .dout(n13444));
  jxor g13189(.dina(n13444), .dinb(n13432), .dout(n13445));
  jxor g13190(.dina(n13445), .dinb(n13263), .dout(n13446));
  jxor g13191(.dina(n13446), .dinb(n13251), .dout(n13447));
  jxor g13192(.dina(n13447), .dinb(n13239), .dout(n13448));
  jxor g13193(.dina(n13448), .dinb(n13227), .dout(n13449));
  jxor g13194(.dina(n13449), .dinb(n13218), .dout(n13450));
  jnot g13195(.din(n13450), .dout(n13451));
  jxor g13196(.dina(n13451), .dinb(n13215), .dout(f74 ));
  jand g13197(.dina(n13449), .dinb(n13218), .dout(n13453));
  jnot g13198(.din(n13453), .dout(n13454));
  jor  g13199(.dina(n13451), .dinb(n13215), .dout(n13455));
  jand g13200(.dina(n13455), .dinb(n13454), .dout(n13456));
  jor  g13201(.dina(n13226), .dinb(n13222), .dout(n13457));
  jand g13202(.dina(n13448), .dinb(n13227), .dout(n13458));
  jnot g13203(.din(n13458), .dout(n13459));
  jand g13204(.dina(n13459), .dinb(n13457), .dout(n13460));
  jnot g13205(.din(n13460), .dout(n13461));
  jand g13206(.dina(n13238), .dinb(n13230), .dout(n13462));
  jand g13207(.dina(n13447), .dinb(n13239), .dout(n13463));
  jor  g13208(.dina(n13463), .dinb(n13462), .dout(n13464));
  jor  g13209(.dina(n10521), .dinb(n970), .dout(n13465));
  jor  g13210(.dina(n880), .dinb(n9759), .dout(n13466));
  jor  g13211(.dina(n967), .dinb(n10051), .dout(n13467));
  jor  g13212(.dina(n972), .dinb(n10523), .dout(n13468));
  jand g13213(.dina(n13468), .dinb(n13467), .dout(n13469));
  jand g13214(.dina(n13469), .dinb(n13466), .dout(n13470));
  jand g13215(.dina(n13470), .dinb(n13465), .dout(n13471));
  jxor g13216(.dina(n13471), .dinb(n810), .dout(n13472));
  jxor g13217(.dina(n13472), .dinb(n13464), .dout(n13473));
  jand g13218(.dina(n13250), .dinb(n13242), .dout(n13474));
  jand g13219(.dina(n13446), .dinb(n13251), .dout(n13475));
  jor  g13220(.dina(n13475), .dinb(n13474), .dout(n13476));
  jor  g13221(.dina(n9473), .dinb(n1248), .dout(n13477));
  jor  g13222(.dina(n1147), .dinb(n8920), .dout(n13478));
  jor  g13223(.dina(n1251), .dinb(n9195), .dout(n13479));
  jor  g13224(.dina(n1246), .dinb(n9475), .dout(n13480));
  jand g13225(.dina(n13480), .dinb(n13479), .dout(n13481));
  jand g13226(.dina(n13481), .dinb(n13478), .dout(n13482));
  jand g13227(.dina(n13482), .dinb(n13477), .dout(n13483));
  jxor g13228(.dina(n13483), .dinb(n1061), .dout(n13484));
  jxor g13229(.dina(n13484), .dinb(n13476), .dout(n13485));
  jand g13230(.dina(n13262), .dinb(n13254), .dout(n13486));
  jand g13231(.dina(n13445), .dinb(n13263), .dout(n13487));
  jor  g13232(.dina(n13487), .dinb(n13486), .dout(n13488));
  jor  g13233(.dina(n8642), .dinb(n1569), .dout(n13489));
  jor  g13234(.dina(n1453), .dinb(n8111), .dout(n13490));
  jor  g13235(.dina(n1566), .dinb(n8378), .dout(n13491));
  jor  g13236(.dina(n1571), .dinb(n8644), .dout(n13492));
  jand g13237(.dina(n13492), .dinb(n13491), .dout(n13493));
  jand g13238(.dina(n13493), .dinb(n13490), .dout(n13494));
  jand g13239(.dina(n13494), .dinb(n13489), .dout(n13495));
  jxor g13240(.dina(n13495), .dinb(n1351), .dout(n13496));
  jxor g13241(.dina(n13496), .dinb(n13488), .dout(n13497));
  jand g13242(.dina(n13274), .dinb(n13266), .dout(n13498));
  jand g13243(.dina(n13431), .dinb(n13275), .dout(n13499));
  jor  g13244(.dina(n13499), .dinb(n13498), .dout(n13500));
  jor  g13245(.dina(n7084), .dinb(n2324), .dout(n13501));
  jor  g13246(.dina(n2186), .dinb(n6605), .dout(n13502));
  jor  g13247(.dina(n2321), .dinb(n6846), .dout(n13503));
  jor  g13248(.dina(n2326), .dinb(n7086), .dout(n13504));
  jand g13249(.dina(n13504), .dinb(n13503), .dout(n13505));
  jand g13250(.dina(n13505), .dinb(n13502), .dout(n13506));
  jand g13251(.dina(n13506), .dinb(n13501), .dout(n13507));
  jxor g13252(.dina(n13507), .dinb(n2057), .dout(n13508));
  jxor g13253(.dina(n13508), .dinb(n13500), .dout(n13509));
  jand g13254(.dina(n13286), .dinb(n13278), .dout(n13510));
  jand g13255(.dina(n13430), .dinb(n13287), .dout(n13511));
  jor  g13256(.dina(n13511), .dinb(n13510), .dout(n13512));
  jor  g13257(.dina(n6364), .dinb(n2764), .dout(n13513));
  jor  g13258(.dina(n2609), .dinb(n5911), .dout(n13514));
  jor  g13259(.dina(n2761), .dinb(n6366), .dout(n13515));
  jor  g13260(.dina(n2766), .dinb(n6139), .dout(n13516));
  jand g13261(.dina(n13516), .dinb(n13515), .dout(n13517));
  jand g13262(.dina(n13517), .dinb(n13514), .dout(n13518));
  jand g13263(.dina(n13518), .dinb(n13513), .dout(n13519));
  jxor g13264(.dina(n13519), .dinb(n2468), .dout(n13520));
  jxor g13265(.dina(n13520), .dinb(n13512), .dout(n13521));
  jand g13266(.dina(n13419), .dinb(n13302), .dout(n13522));
  jand g13267(.dina(n13428), .dinb(n13420), .dout(n13523));
  jor  g13268(.dina(n13523), .dinb(n13522), .dout(n13524));
  jand g13269(.dina(n13409), .dinb(n13305), .dout(n13525));
  jand g13270(.dina(n13418), .dinb(n13410), .dout(n13526));
  jor  g13271(.dina(n13526), .dinb(n13525), .dout(n13527));
  jand g13272(.dina(n13399), .dinb(n13396), .dout(n13528));
  jand g13273(.dina(n13408), .dinb(n13400), .dout(n13529));
  jor  g13274(.dina(n13529), .dinb(n13528), .dout(n13530));
  jand g13275(.dina(n13386), .dinb(n13308), .dout(n13531));
  jand g13276(.dina(n13395), .dinb(n13387), .dout(n13532));
  jor  g13277(.dina(n13532), .dinb(n13531), .dout(n13533));
  jand g13278(.dina(n13376), .dinb(n13311), .dout(n13534));
  jand g13279(.dina(n13385), .dinb(n13377), .dout(n13535));
  jor  g13280(.dina(n13535), .dinb(n13534), .dout(n13536));
  jand g13281(.dina(n13366), .dinb(n13314), .dout(n13537));
  jand g13282(.dina(n13375), .dinb(n13367), .dout(n13538));
  jor  g13283(.dina(n13538), .dinb(n13537), .dout(n13539));
  jand g13284(.dina(n13356), .dinb(n13317), .dout(n13540));
  jand g13285(.dina(n13365), .dinb(n13357), .dout(n13541));
  jor  g13286(.dina(n13541), .dinb(n13540), .dout(n13542));
  jand g13287(.dina(n13346), .dinb(n13320), .dout(n13543));
  jand g13288(.dina(n13355), .dinb(n13347), .dout(n13544));
  jor  g13289(.dina(n13544), .dinb(n13543), .dout(n13545));
  jand g13290(.dina(n13336), .dinb(n13328), .dout(n13546));
  jand g13291(.dina(n13345), .dinb(n13337), .dout(n13547));
  jor  g13292(.dina(n13547), .dinb(n13546), .dout(n13548));
  jand g13293(.dina(n13326), .dinb(n13056), .dout(n13549));
  jand g13294(.dina(n13327), .dinb(n13323), .dout(n13550));
  jor  g13295(.dina(n13550), .dinb(n13549), .dout(n13551));
  jand g13296(.dina(n10594), .dinb(b11 ), .dout(n13552));
  jand g13297(.dina(n10129), .dinb(b12 ), .dout(n13553));
  jor  g13298(.dina(n13553), .dinb(n13552), .dout(n13554));
  jxor g13299(.dina(n13055), .dinb(n606), .dout(n13555));
  jxor g13300(.dina(n13555), .dinb(n13554), .dout(n13556));
  jor  g13301(.dina(n10134), .dinb(n1016), .dout(n13557));
  jor  g13302(.dina(n9849), .dinb(n852), .dout(n13558));
  jor  g13303(.dina(n10137), .dinb(n934), .dout(n13559));
  jor  g13304(.dina(n10132), .dinb(n1018), .dout(n13560));
  jand g13305(.dina(n13560), .dinb(n13559), .dout(n13561));
  jand g13306(.dina(n13561), .dinb(n13558), .dout(n13562));
  jand g13307(.dina(n13562), .dinb(n13557), .dout(n13563));
  jxor g13308(.dina(n13563), .dinb(n9559), .dout(n13564));
  jxor g13309(.dina(n13564), .dinb(n13556), .dout(n13565));
  jxor g13310(.dina(n13565), .dinb(n13551), .dout(n13566));
  jor  g13311(.dina(n9271), .dinb(n1305), .dout(n13567));
  jor  g13312(.dina(n9003), .dinb(n1114), .dout(n13568));
  jor  g13313(.dina(n9268), .dinb(n1307), .dout(n13569));
  jor  g13314(.dina(n9273), .dinb(n1211), .dout(n13570));
  jand g13315(.dina(n13570), .dinb(n13569), .dout(n13571));
  jand g13316(.dina(n13571), .dinb(n13568), .dout(n13572));
  jand g13317(.dina(n13572), .dinb(n13567), .dout(n13573));
  jxor g13318(.dina(n13573), .dinb(n8729), .dout(n13574));
  jxor g13319(.dina(n13574), .dinb(n13566), .dout(n13575));
  jxor g13320(.dina(n13575), .dinb(n13548), .dout(n13576));
  jor  g13321(.dina(n8457), .dinb(n1635), .dout(n13577));
  jor  g13322(.dina(n8185), .dinb(n1416), .dout(n13578));
  jor  g13323(.dina(n8459), .dinb(n1527), .dout(n13579));
  jor  g13324(.dina(n8454), .dinb(n1637), .dout(n13580));
  jand g13325(.dina(n13580), .dinb(n13579), .dout(n13581));
  jand g13326(.dina(n13581), .dinb(n13578), .dout(n13582));
  jand g13327(.dina(n13582), .dinb(n13577), .dout(n13583));
  jxor g13328(.dina(n13583), .dinb(n7929), .dout(n13584));
  jxor g13329(.dina(n13584), .dinb(n13576), .dout(n13585));
  jxor g13330(.dina(n13585), .dinb(n13545), .dout(n13586));
  jor  g13331(.dina(n7660), .dinb(n2005), .dout(n13587));
  jor  g13332(.dina(n7415), .dinb(n1759), .dout(n13588));
  jor  g13333(.dina(n7657), .dinb(n1881), .dout(n13589));
  jor  g13334(.dina(n7662), .dinb(n2007), .dout(n13590));
  jand g13335(.dina(n13590), .dinb(n13589), .dout(n13591));
  jand g13336(.dina(n13591), .dinb(n13588), .dout(n13592));
  jand g13337(.dina(n13592), .dinb(n13587), .dout(n13593));
  jxor g13338(.dina(n13593), .dinb(n7166), .dout(n13594));
  jxor g13339(.dina(n13594), .dinb(n13586), .dout(n13595));
  jxor g13340(.dina(n13595), .dinb(n13542), .dout(n13596));
  jor  g13341(.dina(n6914), .dinb(n2413), .dout(n13597));
  jor  g13342(.dina(n6673), .dinb(n2142), .dout(n13598));
  jor  g13343(.dina(n6916), .dinb(n2415), .dout(n13599));
  jor  g13344(.dina(n6911), .dinb(n2279), .dout(n13600));
  jand g13345(.dina(n13600), .dinb(n13599), .dout(n13601));
  jand g13346(.dina(n13601), .dinb(n13598), .dout(n13602));
  jand g13347(.dina(n13602), .dinb(n13597), .dout(n13603));
  jxor g13348(.dina(n13603), .dinb(n6443), .dout(n13604));
  jxor g13349(.dina(n13604), .dinb(n13596), .dout(n13605));
  jxor g13350(.dina(n13605), .dinb(n13539), .dout(n13606));
  jor  g13351(.dina(n6207), .dinb(n2860), .dout(n13607));
  jor  g13352(.dina(n5975), .dinb(n2563), .dout(n13608));
  jor  g13353(.dina(n6210), .dinb(n2713), .dout(n13609));
  jor  g13354(.dina(n6205), .dinb(n2862), .dout(n13610));
  jand g13355(.dina(n13610), .dinb(n13609), .dout(n13611));
  jand g13356(.dina(n13611), .dinb(n13608), .dout(n13612));
  jand g13357(.dina(n13612), .dinb(n13607), .dout(n13613));
  jxor g13358(.dina(n13613), .dinb(n5759), .dout(n13614));
  jxor g13359(.dina(n13614), .dinb(n13606), .dout(n13615));
  jxor g13360(.dina(n13615), .dinb(n13536), .dout(n13616));
  jor  g13361(.dina(n5537), .dinb(n3346), .dout(n13617));
  jor  g13362(.dina(n5315), .dinb(n3023), .dout(n13618));
  jor  g13363(.dina(n5534), .dinb(n3186), .dout(n13619));
  jor  g13364(.dina(n5539), .dinb(n3348), .dout(n13620));
  jand g13365(.dina(n13620), .dinb(n13619), .dout(n13621));
  jand g13366(.dina(n13621), .dinb(n13618), .dout(n13622));
  jand g13367(.dina(n13622), .dinb(n13617), .dout(n13623));
  jxor g13368(.dina(n13623), .dinb(n5111), .dout(n13624));
  jxor g13369(.dina(n13624), .dinb(n13616), .dout(n13625));
  jxor g13370(.dina(n13625), .dinb(n13533), .dout(n13626));
  jor  g13371(.dina(n4902), .dinb(n3871), .dout(n13627));
  jor  g13372(.dina(n4696), .dinb(n3522), .dout(n13628));
  jor  g13373(.dina(n4904), .dinb(n3698), .dout(n13629));
  jor  g13374(.dina(n4899), .dinb(n3873), .dout(n13630));
  jand g13375(.dina(n13630), .dinb(n13629), .dout(n13631));
  jand g13376(.dina(n13631), .dinb(n13628), .dout(n13632));
  jand g13377(.dina(n13632), .dinb(n13627), .dout(n13633));
  jxor g13378(.dina(n13633), .dinb(n4505), .dout(n13634));
  jxor g13379(.dina(n13634), .dinb(n13626), .dout(n13635));
  jxor g13380(.dina(n13635), .dinb(n13530), .dout(n13636));
  jor  g13381(.dina(n4435), .dinb(n4305), .dout(n13637));
  jor  g13382(.dina(n4116), .dinb(n4060), .dout(n13638));
  jor  g13383(.dina(n4303), .dinb(n4437), .dout(n13639));
  jor  g13384(.dina(n4308), .dinb(n4249), .dout(n13640));
  jand g13385(.dina(n13640), .dinb(n13639), .dout(n13641));
  jand g13386(.dina(n13641), .dinb(n13638), .dout(n13642));
  jand g13387(.dina(n13642), .dinb(n13637), .dout(n13643));
  jxor g13388(.dina(n13643), .dinb(n3938), .dout(n13644));
  jxor g13389(.dina(n13644), .dinb(n13636), .dout(n13645));
  jxor g13390(.dina(n13645), .dinb(n13527), .dout(n13646));
  jor  g13391(.dina(n5038), .dinb(n3751), .dout(n13647));
  jor  g13392(.dina(n3574), .dinb(n4637), .dout(n13648));
  jor  g13393(.dina(n3754), .dinb(n4839), .dout(n13649));
  jor  g13394(.dina(n3749), .dinb(n5040), .dout(n13650));
  jand g13395(.dina(n13650), .dinb(n13649), .dout(n13651));
  jand g13396(.dina(n13651), .dinb(n13648), .dout(n13652));
  jand g13397(.dina(n13652), .dinb(n13647), .dout(n13653));
  jxor g13398(.dina(n13653), .dinb(n3410), .dout(n13654));
  jxor g13399(.dina(n13654), .dinb(n13646), .dout(n13655));
  jxor g13400(.dina(n13655), .dinb(n13524), .dout(n13656));
  jand g13401(.dina(n13298), .dinb(n13290), .dout(n13657));
  jand g13402(.dina(n13429), .dinb(n13299), .dout(n13658));
  jor  g13403(.dina(n13658), .dinb(n13657), .dout(n13659));
  jor  g13404(.dina(n5683), .dinb(n3239), .dout(n13660));
  jor  g13405(.dina(n3072), .dinb(n5253), .dout(n13661));
  jor  g13406(.dina(n3242), .dinb(n5469), .dout(n13662));
  jor  g13407(.dina(n3237), .dinb(n5685), .dout(n13663));
  jand g13408(.dina(n13663), .dinb(n13662), .dout(n13664));
  jand g13409(.dina(n13664), .dinb(n13661), .dout(n13665));
  jand g13410(.dina(n13665), .dinb(n13660), .dout(n13666));
  jxor g13411(.dina(n13666), .dinb(n2918), .dout(n13667));
  jxor g13412(.dina(n13667), .dinb(n13659), .dout(n13668));
  jxor g13413(.dina(n13668), .dinb(n13656), .dout(n13669));
  jxor g13414(.dina(n13669), .dinb(n13521), .dout(n13670));
  jxor g13415(.dina(n13670), .dinb(n13509), .dout(n13671));
  jand g13416(.dina(n13443), .dinb(n13435), .dout(n13672));
  jand g13417(.dina(n13444), .dinb(n13432), .dout(n13673));
  jor  g13418(.dina(n13673), .dinb(n13672), .dout(n13674));
  jor  g13419(.dina(n7844), .dinb(n1921), .dout(n13675));
  jor  g13420(.dina(n1806), .dinb(n7338), .dout(n13676));
  jor  g13421(.dina(n1918), .dinb(n7590), .dout(n13677));
  jor  g13422(.dina(n1923), .dinb(n7846), .dout(n13678));
  jand g13423(.dina(n13678), .dinb(n13677), .dout(n13679));
  jand g13424(.dina(n13679), .dinb(n13676), .dout(n13680));
  jand g13425(.dina(n13680), .dinb(n13675), .dout(n13681));
  jxor g13426(.dina(n13681), .dinb(n1687), .dout(n13682));
  jxor g13427(.dina(n13682), .dinb(n13674), .dout(n13683));
  jxor g13428(.dina(n13683), .dinb(n13671), .dout(n13684));
  jxor g13429(.dina(n13684), .dinb(n13497), .dout(n13685));
  jxor g13430(.dina(n13685), .dinb(n13485), .dout(n13686));
  jxor g13431(.dina(n13686), .dinb(n13473), .dout(n13687));
  jxor g13432(.dina(n13687), .dinb(n13461), .dout(n13688));
  jnot g13433(.din(n13688), .dout(n13689));
  jxor g13434(.dina(n13689), .dinb(n13456), .dout(f75 ));
  jand g13435(.dina(n13687), .dinb(n13461), .dout(n13691));
  jnot g13436(.din(n13691), .dout(n13692));
  jor  g13437(.dina(n13689), .dinb(n13456), .dout(n13693));
  jand g13438(.dina(n13693), .dinb(n13692), .dout(n13694));
  jand g13439(.dina(n13472), .dinb(n13464), .dout(n13695));
  jand g13440(.dina(n13686), .dinb(n13473), .dout(n13696));
  jor  g13441(.dina(n13696), .dinb(n13695), .dout(n13697));
  jand g13442(.dina(n13508), .dinb(n13500), .dout(n13698));
  jand g13443(.dina(n13670), .dinb(n13509), .dout(n13699));
  jor  g13444(.dina(n13699), .dinb(n13698), .dout(n13700));
  jor  g13445(.dina(n8109), .dinb(n1921), .dout(n13701));
  jor  g13446(.dina(n1806), .dinb(n7590), .dout(n13702));
  jor  g13447(.dina(n1918), .dinb(n7846), .dout(n13703));
  jor  g13448(.dina(n1923), .dinb(n8111), .dout(n13704));
  jand g13449(.dina(n13704), .dinb(n13703), .dout(n13705));
  jand g13450(.dina(n13705), .dinb(n13702), .dout(n13706));
  jand g13451(.dina(n13706), .dinb(n13701), .dout(n13707));
  jxor g13452(.dina(n13707), .dinb(n1687), .dout(n13708));
  jxor g13453(.dina(n13708), .dinb(n13700), .dout(n13709));
  jand g13454(.dina(n13520), .dinb(n13512), .dout(n13710));
  jand g13455(.dina(n13669), .dinb(n13521), .dout(n13711));
  jor  g13456(.dina(n13711), .dinb(n13710), .dout(n13712));
  jor  g13457(.dina(n7336), .dinb(n2324), .dout(n13713));
  jor  g13458(.dina(n2186), .dinb(n6846), .dout(n13714));
  jor  g13459(.dina(n2326), .dinb(n7338), .dout(n13715));
  jor  g13460(.dina(n2321), .dinb(n7086), .dout(n13716));
  jand g13461(.dina(n13716), .dinb(n13715), .dout(n13717));
  jand g13462(.dina(n13717), .dinb(n13714), .dout(n13718));
  jand g13463(.dina(n13718), .dinb(n13713), .dout(n13719));
  jxor g13464(.dina(n13719), .dinb(n2057), .dout(n13720));
  jxor g13465(.dina(n13720), .dinb(n13712), .dout(n13721));
  jand g13466(.dina(n13667), .dinb(n13659), .dout(n13722));
  jand g13467(.dina(n13668), .dinb(n13656), .dout(n13723));
  jor  g13468(.dina(n13723), .dinb(n13722), .dout(n13724));
  jor  g13469(.dina(n6603), .dinb(n2764), .dout(n13725));
  jor  g13470(.dina(n2609), .dinb(n6139), .dout(n13726));
  jor  g13471(.dina(n2761), .dinb(n6605), .dout(n13727));
  jor  g13472(.dina(n2766), .dinb(n6366), .dout(n13728));
  jand g13473(.dina(n13728), .dinb(n13727), .dout(n13729));
  jand g13474(.dina(n13729), .dinb(n13726), .dout(n13730));
  jand g13475(.dina(n13730), .dinb(n13725), .dout(n13731));
  jxor g13476(.dina(n13731), .dinb(n2468), .dout(n13732));
  jxor g13477(.dina(n13732), .dinb(n13724), .dout(n13733));
  jand g13478(.dina(n13644), .dinb(n13636), .dout(n13734));
  jand g13479(.dina(n13645), .dinb(n13527), .dout(n13735));
  jor  g13480(.dina(n13735), .dinb(n13734), .dout(n13736));
  jand g13481(.dina(n13634), .dinb(n13626), .dout(n13737));
  jand g13482(.dina(n13635), .dinb(n13530), .dout(n13738));
  jor  g13483(.dina(n13738), .dinb(n13737), .dout(n13739));
  jand g13484(.dina(n13624), .dinb(n13616), .dout(n13740));
  jand g13485(.dina(n13625), .dinb(n13533), .dout(n13741));
  jor  g13486(.dina(n13741), .dinb(n13740), .dout(n13742));
  jand g13487(.dina(n13604), .dinb(n13596), .dout(n13743));
  jand g13488(.dina(n13605), .dinb(n13539), .dout(n13744));
  jor  g13489(.dina(n13744), .dinb(n13743), .dout(n13745));
  jand g13490(.dina(n13594), .dinb(n13586), .dout(n13746));
  jand g13491(.dina(n13595), .dinb(n13542), .dout(n13747));
  jor  g13492(.dina(n13747), .dinb(n13746), .dout(n13748));
  jand g13493(.dina(n13584), .dinb(n13576), .dout(n13749));
  jand g13494(.dina(n13585), .dinb(n13545), .dout(n13750));
  jor  g13495(.dina(n13750), .dinb(n13749), .dout(n13751));
  jand g13496(.dina(n13574), .dinb(n13566), .dout(n13752));
  jand g13497(.dina(n13575), .dinb(n13548), .dout(n13753));
  jor  g13498(.dina(n13753), .dinb(n13752), .dout(n13754));
  jand g13499(.dina(n13564), .dinb(n13556), .dout(n13755));
  jand g13500(.dina(n13565), .dinb(n13551), .dout(n13756));
  jor  g13501(.dina(n13756), .dinb(n13755), .dout(n13757));
  jand g13502(.dina(n10594), .dinb(b12 ), .dout(n13758));
  jand g13503(.dina(n10129), .dinb(b13 ), .dout(n13759));
  jor  g13504(.dina(n13759), .dinb(n13758), .dout(n13760));
  jnot g13505(.din(n13760), .dout(n13761));
  jand g13506(.dina(n13055), .dinb(n606), .dout(n13762));
  jand g13507(.dina(n13555), .dinb(n13554), .dout(n13763));
  jor  g13508(.dina(n13763), .dinb(n13762), .dout(n13764));
  jxor g13509(.dina(n13764), .dinb(n13761), .dout(n13765));
  jor  g13510(.dina(n10134), .dinb(n1112), .dout(n13766));
  jor  g13511(.dina(n9849), .dinb(n934), .dout(n13767));
  jor  g13512(.dina(n10132), .dinb(n1114), .dout(n13768));
  jor  g13513(.dina(n10137), .dinb(n1018), .dout(n13769));
  jand g13514(.dina(n13769), .dinb(n13768), .dout(n13770));
  jand g13515(.dina(n13770), .dinb(n13767), .dout(n13771));
  jand g13516(.dina(n13771), .dinb(n13766), .dout(n13772));
  jxor g13517(.dina(n13772), .dinb(n9559), .dout(n13773));
  jxor g13518(.dina(n13773), .dinb(n13765), .dout(n13774));
  jxor g13519(.dina(n13774), .dinb(n13757), .dout(n13775));
  jor  g13520(.dina(n9271), .dinb(n1414), .dout(n13776));
  jor  g13521(.dina(n9003), .dinb(n1211), .dout(n13777));
  jor  g13522(.dina(n9273), .dinb(n1307), .dout(n13778));
  jor  g13523(.dina(n9268), .dinb(n1416), .dout(n13779));
  jand g13524(.dina(n13779), .dinb(n13778), .dout(n13780));
  jand g13525(.dina(n13780), .dinb(n13777), .dout(n13781));
  jand g13526(.dina(n13781), .dinb(n13776), .dout(n13782));
  jxor g13527(.dina(n13782), .dinb(n8729), .dout(n13783));
  jxor g13528(.dina(n13783), .dinb(n13775), .dout(n13784));
  jxor g13529(.dina(n13784), .dinb(n13754), .dout(n13785));
  jor  g13530(.dina(n8457), .dinb(n1757), .dout(n13786));
  jor  g13531(.dina(n8185), .dinb(n1527), .dout(n13787));
  jor  g13532(.dina(n8459), .dinb(n1637), .dout(n13788));
  jor  g13533(.dina(n8454), .dinb(n1759), .dout(n13789));
  jand g13534(.dina(n13789), .dinb(n13788), .dout(n13790));
  jand g13535(.dina(n13790), .dinb(n13787), .dout(n13791));
  jand g13536(.dina(n13791), .dinb(n13786), .dout(n13792));
  jxor g13537(.dina(n13792), .dinb(n7929), .dout(n13793));
  jxor g13538(.dina(n13793), .dinb(n13785), .dout(n13794));
  jxor g13539(.dina(n13794), .dinb(n13751), .dout(n13795));
  jor  g13540(.dina(n7660), .dinb(n2140), .dout(n13796));
  jor  g13541(.dina(n7415), .dinb(n1881), .dout(n13797));
  jor  g13542(.dina(n7662), .dinb(n2142), .dout(n13798));
  jor  g13543(.dina(n7657), .dinb(n2007), .dout(n13799));
  jand g13544(.dina(n13799), .dinb(n13798), .dout(n13800));
  jand g13545(.dina(n13800), .dinb(n13797), .dout(n13801));
  jand g13546(.dina(n13801), .dinb(n13796), .dout(n13802));
  jxor g13547(.dina(n13802), .dinb(n7166), .dout(n13803));
  jxor g13548(.dina(n13803), .dinb(n13795), .dout(n13804));
  jxor g13549(.dina(n13804), .dinb(n13748), .dout(n13805));
  jor  g13550(.dina(n6914), .dinb(n2561), .dout(n13806));
  jor  g13551(.dina(n6673), .dinb(n2279), .dout(n13807));
  jor  g13552(.dina(n6911), .dinb(n2415), .dout(n13808));
  jor  g13553(.dina(n6916), .dinb(n2563), .dout(n13809));
  jand g13554(.dina(n13809), .dinb(n13808), .dout(n13810));
  jand g13555(.dina(n13810), .dinb(n13807), .dout(n13811));
  jand g13556(.dina(n13811), .dinb(n13806), .dout(n13812));
  jxor g13557(.dina(n13812), .dinb(n6443), .dout(n13813));
  jxor g13558(.dina(n13813), .dinb(n13805), .dout(n13814));
  jxor g13559(.dina(n13814), .dinb(n13745), .dout(n13815));
  jor  g13560(.dina(n6207), .dinb(n3021), .dout(n13816));
  jor  g13561(.dina(n5975), .dinb(n2713), .dout(n13817));
  jor  g13562(.dina(n6210), .dinb(n2862), .dout(n13818));
  jor  g13563(.dina(n6205), .dinb(n3023), .dout(n13819));
  jand g13564(.dina(n13819), .dinb(n13818), .dout(n13820));
  jand g13565(.dina(n13820), .dinb(n13817), .dout(n13821));
  jand g13566(.dina(n13821), .dinb(n13816), .dout(n13822));
  jxor g13567(.dina(n13822), .dinb(n5759), .dout(n13823));
  jxor g13568(.dina(n13823), .dinb(n13815), .dout(n13824));
  jnot g13569(.din(n13606), .dout(n13825));
  jnot g13570(.din(n13614), .dout(n13826));
  jand g13571(.dina(n13826), .dinb(n13825), .dout(n13827));
  jnot g13572(.din(n13827), .dout(n13828));
  jand g13573(.dina(n13614), .dinb(n13606), .dout(n13829));
  jor  g13574(.dina(n13829), .dinb(n13536), .dout(n13830));
  jand g13575(.dina(n13830), .dinb(n13828), .dout(n13831));
  jxor g13576(.dina(n13831), .dinb(n13824), .dout(n13832));
  jor  g13577(.dina(n5537), .dinb(n3520), .dout(n13833));
  jor  g13578(.dina(n5315), .dinb(n3186), .dout(n13834));
  jor  g13579(.dina(n5534), .dinb(n3348), .dout(n13835));
  jor  g13580(.dina(n5539), .dinb(n3522), .dout(n13836));
  jand g13581(.dina(n13836), .dinb(n13835), .dout(n13837));
  jand g13582(.dina(n13837), .dinb(n13834), .dout(n13838));
  jand g13583(.dina(n13838), .dinb(n13833), .dout(n13839));
  jxor g13584(.dina(n13839), .dinb(n5111), .dout(n13840));
  jxor g13585(.dina(n13840), .dinb(n13832), .dout(n13841));
  jxor g13586(.dina(n13841), .dinb(n13742), .dout(n13842));
  jor  g13587(.dina(n4902), .dinb(n4058), .dout(n13843));
  jor  g13588(.dina(n4696), .dinb(n3698), .dout(n13844));
  jor  g13589(.dina(n4899), .dinb(n4060), .dout(n13845));
  jor  g13590(.dina(n4904), .dinb(n3873), .dout(n13846));
  jand g13591(.dina(n13846), .dinb(n13845), .dout(n13847));
  jand g13592(.dina(n13847), .dinb(n13844), .dout(n13848));
  jand g13593(.dina(n13848), .dinb(n13843), .dout(n13849));
  jxor g13594(.dina(n13849), .dinb(n4505), .dout(n13850));
  jxor g13595(.dina(n13850), .dinb(n13842), .dout(n13851));
  jxor g13596(.dina(n13851), .dinb(n13739), .dout(n13852));
  jor  g13597(.dina(n4635), .dinb(n4305), .dout(n13853));
  jor  g13598(.dina(n4116), .dinb(n4249), .dout(n13854));
  jor  g13599(.dina(n4303), .dinb(n4637), .dout(n13855));
  jor  g13600(.dina(n4308), .dinb(n4437), .dout(n13856));
  jand g13601(.dina(n13856), .dinb(n13855), .dout(n13857));
  jand g13602(.dina(n13857), .dinb(n13854), .dout(n13858));
  jand g13603(.dina(n13858), .dinb(n13853), .dout(n13859));
  jxor g13604(.dina(n13859), .dinb(n3938), .dout(n13860));
  jxor g13605(.dina(n13860), .dinb(n13852), .dout(n13861));
  jxor g13606(.dina(n13861), .dinb(n13736), .dout(n13862));
  jor  g13607(.dina(n5251), .dinb(n3751), .dout(n13863));
  jor  g13608(.dina(n3574), .dinb(n4839), .dout(n13864));
  jor  g13609(.dina(n3754), .dinb(n5040), .dout(n13865));
  jor  g13610(.dina(n3749), .dinb(n5253), .dout(n13866));
  jand g13611(.dina(n13866), .dinb(n13865), .dout(n13867));
  jand g13612(.dina(n13867), .dinb(n13864), .dout(n13868));
  jand g13613(.dina(n13868), .dinb(n13863), .dout(n13869));
  jxor g13614(.dina(n13869), .dinb(n3410), .dout(n13870));
  jxor g13615(.dina(n13870), .dinb(n13862), .dout(n13871));
  jand g13616(.dina(n13654), .dinb(n13646), .dout(n13872));
  jand g13617(.dina(n13655), .dinb(n13524), .dout(n13873));
  jor  g13618(.dina(n13873), .dinb(n13872), .dout(n13874));
  jor  g13619(.dina(n5909), .dinb(n3239), .dout(n13875));
  jor  g13620(.dina(n3072), .dinb(n5469), .dout(n13876));
  jor  g13621(.dina(n3242), .dinb(n5685), .dout(n13877));
  jor  g13622(.dina(n3237), .dinb(n5911), .dout(n13878));
  jand g13623(.dina(n13878), .dinb(n13877), .dout(n13879));
  jand g13624(.dina(n13879), .dinb(n13876), .dout(n13880));
  jand g13625(.dina(n13880), .dinb(n13875), .dout(n13881));
  jxor g13626(.dina(n13881), .dinb(n2918), .dout(n13882));
  jxor g13627(.dina(n13882), .dinb(n13874), .dout(n13883));
  jxor g13628(.dina(n13883), .dinb(n13871), .dout(n13884));
  jxor g13629(.dina(n13884), .dinb(n13733), .dout(n13885));
  jxor g13630(.dina(n13885), .dinb(n13721), .dout(n13886));
  jxor g13631(.dina(n13886), .dinb(n13709), .dout(n13887));
  jand g13632(.dina(n13682), .dinb(n13674), .dout(n13888));
  jand g13633(.dina(n13683), .dinb(n13671), .dout(n13889));
  jor  g13634(.dina(n13889), .dinb(n13888), .dout(n13890));
  jor  g13635(.dina(n8918), .dinb(n1569), .dout(n13891));
  jor  g13636(.dina(n1453), .dinb(n8378), .dout(n13892));
  jor  g13637(.dina(n1566), .dinb(n8644), .dout(n13893));
  jor  g13638(.dina(n1571), .dinb(n8920), .dout(n13894));
  jand g13639(.dina(n13894), .dinb(n13893), .dout(n13895));
  jand g13640(.dina(n13895), .dinb(n13892), .dout(n13896));
  jand g13641(.dina(n13896), .dinb(n13891), .dout(n13897));
  jxor g13642(.dina(n13897), .dinb(n1351), .dout(n13898));
  jxor g13643(.dina(n13898), .dinb(n13890), .dout(n13899));
  jxor g13644(.dina(n13899), .dinb(n13887), .dout(n13900));
  jand g13645(.dina(n13496), .dinb(n13488), .dout(n13901));
  jand g13646(.dina(n13684), .dinb(n13497), .dout(n13902));
  jor  g13647(.dina(n13902), .dinb(n13901), .dout(n13903));
  jor  g13648(.dina(n9757), .dinb(n1248), .dout(n13904));
  jor  g13649(.dina(n1147), .dinb(n9195), .dout(n13905));
  jor  g13650(.dina(n1251), .dinb(n9475), .dout(n13906));
  jor  g13651(.dina(n1246), .dinb(n9759), .dout(n13907));
  jand g13652(.dina(n13907), .dinb(n13906), .dout(n13908));
  jand g13653(.dina(n13908), .dinb(n13905), .dout(n13909));
  jand g13654(.dina(n13909), .dinb(n13904), .dout(n13910));
  jxor g13655(.dina(n13910), .dinb(n1061), .dout(n13911));
  jxor g13656(.dina(n13911), .dinb(n13903), .dout(n13912));
  jxor g13657(.dina(n13912), .dinb(n13900), .dout(n13913));
  jand g13658(.dina(n13484), .dinb(n13476), .dout(n13914));
  jand g13659(.dina(n13685), .dinb(n13485), .dout(n13915));
  jor  g13660(.dina(n13915), .dinb(n13914), .dout(n13916));
  jnot g13661(.din(n13916), .dout(n13917));
  jor  g13662(.dina(n967), .dinb(n10523), .dout(n13918));
  jor  g13663(.dina(n10813), .dinb(n970), .dout(n13919));
  jor  g13664(.dina(n880), .dinb(n10051), .dout(n13920));
  jand g13665(.dina(n13920), .dinb(n13919), .dout(n13921));
  jand g13666(.dina(n13921), .dinb(n13918), .dout(n13922));
  jxor g13667(.dina(n13922), .dinb(a14 ), .dout(n13923));
  jxor g13668(.dina(n13923), .dinb(n13917), .dout(n13924));
  jxor g13669(.dina(n13924), .dinb(n13913), .dout(n13925));
  jxor g13670(.dina(n13925), .dinb(n13697), .dout(n13926));
  jnot g13671(.din(n13926), .dout(n13927));
  jxor g13672(.dina(n13927), .dinb(n13694), .dout(f76 ));
  jand g13673(.dina(n13925), .dinb(n13697), .dout(n13929));
  jnot g13674(.din(n13929), .dout(n13930));
  jor  g13675(.dina(n13927), .dinb(n13694), .dout(n13931));
  jand g13676(.dina(n13931), .dinb(n13930), .dout(n13932));
  jor  g13677(.dina(n13923), .dinb(n13917), .dout(n13933));
  jand g13678(.dina(n13924), .dinb(n13913), .dout(n13934));
  jnot g13679(.din(n13934), .dout(n13935));
  jand g13680(.dina(n13935), .dinb(n13933), .dout(n13936));
  jnot g13681(.din(n13936), .dout(n13937));
  jand g13682(.dina(n13708), .dinb(n13700), .dout(n13938));
  jand g13683(.dina(n13886), .dinb(n13709), .dout(n13939));
  jor  g13684(.dina(n13939), .dinb(n13938), .dout(n13940));
  jor  g13685(.dina(n9193), .dinb(n1569), .dout(n13941));
  jor  g13686(.dina(n1453), .dinb(n8644), .dout(n13942));
  jor  g13687(.dina(n1566), .dinb(n8920), .dout(n13943));
  jor  g13688(.dina(n1571), .dinb(n9195), .dout(n13944));
  jand g13689(.dina(n13944), .dinb(n13943), .dout(n13945));
  jand g13690(.dina(n13945), .dinb(n13942), .dout(n13946));
  jand g13691(.dina(n13946), .dinb(n13941), .dout(n13947));
  jxor g13692(.dina(n13947), .dinb(n1351), .dout(n13948));
  jxor g13693(.dina(n13948), .dinb(n13940), .dout(n13949));
  jand g13694(.dina(n13720), .dinb(n13712), .dout(n13950));
  jand g13695(.dina(n13885), .dinb(n13721), .dout(n13951));
  jor  g13696(.dina(n13951), .dinb(n13950), .dout(n13952));
  jor  g13697(.dina(n8376), .dinb(n1921), .dout(n13953));
  jor  g13698(.dina(n1806), .dinb(n7846), .dout(n13954));
  jor  g13699(.dina(n1923), .dinb(n8378), .dout(n13955));
  jor  g13700(.dina(n1918), .dinb(n8111), .dout(n13956));
  jand g13701(.dina(n13956), .dinb(n13955), .dout(n13957));
  jand g13702(.dina(n13957), .dinb(n13954), .dout(n13958));
  jand g13703(.dina(n13958), .dinb(n13953), .dout(n13959));
  jxor g13704(.dina(n13959), .dinb(n1687), .dout(n13960));
  jxor g13705(.dina(n13960), .dinb(n13952), .dout(n13961));
  jand g13706(.dina(n13732), .dinb(n13724), .dout(n13962));
  jand g13707(.dina(n13884), .dinb(n13733), .dout(n13963));
  jor  g13708(.dina(n13963), .dinb(n13962), .dout(n13964));
  jor  g13709(.dina(n7588), .dinb(n2324), .dout(n13965));
  jor  g13710(.dina(n2186), .dinb(n7086), .dout(n13966));
  jor  g13711(.dina(n2326), .dinb(n7590), .dout(n13967));
  jor  g13712(.dina(n2321), .dinb(n7338), .dout(n13968));
  jand g13713(.dina(n13968), .dinb(n13967), .dout(n13969));
  jand g13714(.dina(n13969), .dinb(n13966), .dout(n13970));
  jand g13715(.dina(n13970), .dinb(n13965), .dout(n13971));
  jxor g13716(.dina(n13971), .dinb(n2057), .dout(n13972));
  jxor g13717(.dina(n13972), .dinb(n13964), .dout(n13973));
  jand g13718(.dina(n13882), .dinb(n13874), .dout(n13974));
  jand g13719(.dina(n13883), .dinb(n13871), .dout(n13975));
  jor  g13720(.dina(n13975), .dinb(n13974), .dout(n13976));
  jor  g13721(.dina(n6844), .dinb(n2764), .dout(n13977));
  jor  g13722(.dina(n2609), .dinb(n6366), .dout(n13978));
  jor  g13723(.dina(n2761), .dinb(n6846), .dout(n13979));
  jor  g13724(.dina(n2766), .dinb(n6605), .dout(n13980));
  jand g13725(.dina(n13980), .dinb(n13979), .dout(n13981));
  jand g13726(.dina(n13981), .dinb(n13978), .dout(n13982));
  jand g13727(.dina(n13982), .dinb(n13977), .dout(n13983));
  jxor g13728(.dina(n13983), .dinb(n2468), .dout(n13984));
  jxor g13729(.dina(n13984), .dinb(n13976), .dout(n13985));
  jand g13730(.dina(n13861), .dinb(n13736), .dout(n13986));
  jand g13731(.dina(n13870), .dinb(n13862), .dout(n13987));
  jor  g13732(.dina(n13987), .dinb(n13986), .dout(n13988));
  jor  g13733(.dina(n6137), .dinb(n3239), .dout(n13989));
  jor  g13734(.dina(n3072), .dinb(n5685), .dout(n13990));
  jor  g13735(.dina(n3242), .dinb(n5911), .dout(n13991));
  jor  g13736(.dina(n3237), .dinb(n6139), .dout(n13992));
  jand g13737(.dina(n13992), .dinb(n13991), .dout(n13993));
  jand g13738(.dina(n13993), .dinb(n13990), .dout(n13994));
  jand g13739(.dina(n13994), .dinb(n13989), .dout(n13995));
  jxor g13740(.dina(n13995), .dinb(n2918), .dout(n13996));
  jxor g13741(.dina(n13996), .dinb(n13988), .dout(n13997));
  jand g13742(.dina(n13851), .dinb(n13739), .dout(n13998));
  jand g13743(.dina(n13860), .dinb(n13852), .dout(n13999));
  jor  g13744(.dina(n13999), .dinb(n13998), .dout(n14000));
  jand g13745(.dina(n13841), .dinb(n13742), .dout(n14001));
  jand g13746(.dina(n13850), .dinb(n13842), .dout(n14002));
  jor  g13747(.dina(n14002), .dinb(n14001), .dout(n14003));
  jand g13748(.dina(n13831), .dinb(n13824), .dout(n14004));
  jand g13749(.dina(n13840), .dinb(n13832), .dout(n14005));
  jor  g13750(.dina(n14005), .dinb(n14004), .dout(n14006));
  jand g13751(.dina(n13814), .dinb(n13745), .dout(n14007));
  jand g13752(.dina(n13823), .dinb(n13815), .dout(n14008));
  jor  g13753(.dina(n14008), .dinb(n14007), .dout(n14009));
  jand g13754(.dina(n13804), .dinb(n13748), .dout(n14010));
  jand g13755(.dina(n13813), .dinb(n13805), .dout(n14011));
  jor  g13756(.dina(n14011), .dinb(n14010), .dout(n14012));
  jand g13757(.dina(n13794), .dinb(n13751), .dout(n14013));
  jand g13758(.dina(n13803), .dinb(n13795), .dout(n14014));
  jor  g13759(.dina(n14014), .dinb(n14013), .dout(n14015));
  jand g13760(.dina(n13784), .dinb(n13754), .dout(n14016));
  jand g13761(.dina(n13793), .dinb(n13785), .dout(n14017));
  jor  g13762(.dina(n14017), .dinb(n14016), .dout(n14018));
  jand g13763(.dina(n13774), .dinb(n13757), .dout(n14019));
  jand g13764(.dina(n13783), .dinb(n13775), .dout(n14020));
  jor  g13765(.dina(n14020), .dinb(n14019), .dout(n14021));
  jand g13766(.dina(n13764), .dinb(n13761), .dout(n14022));
  jand g13767(.dina(n13773), .dinb(n13765), .dout(n14023));
  jor  g13768(.dina(n14023), .dinb(n14022), .dout(n14024));
  jand g13769(.dina(n10594), .dinb(b13 ), .dout(n14025));
  jand g13770(.dina(n10129), .dinb(b14 ), .dout(n14026));
  jor  g13771(.dina(n14026), .dinb(n14025), .dout(n14027));
  jxor g13772(.dina(n14027), .dinb(n13761), .dout(n14028));
  jor  g13773(.dina(n10134), .dinb(n1209), .dout(n14029));
  jor  g13774(.dina(n9849), .dinb(n1018), .dout(n14030));
  jor  g13775(.dina(n10137), .dinb(n1114), .dout(n14031));
  jor  g13776(.dina(n10132), .dinb(n1211), .dout(n14032));
  jand g13777(.dina(n14032), .dinb(n14031), .dout(n14033));
  jand g13778(.dina(n14033), .dinb(n14030), .dout(n14034));
  jand g13779(.dina(n14034), .dinb(n14029), .dout(n14035));
  jxor g13780(.dina(n14035), .dinb(n9559), .dout(n14036));
  jxor g13781(.dina(n14036), .dinb(n14028), .dout(n14037));
  jxor g13782(.dina(n14037), .dinb(n14024), .dout(n14038));
  jor  g13783(.dina(n9271), .dinb(n1525), .dout(n14039));
  jor  g13784(.dina(n9003), .dinb(n1307), .dout(n14040));
  jor  g13785(.dina(n9273), .dinb(n1416), .dout(n14041));
  jor  g13786(.dina(n9268), .dinb(n1527), .dout(n14042));
  jand g13787(.dina(n14042), .dinb(n14041), .dout(n14043));
  jand g13788(.dina(n14043), .dinb(n14040), .dout(n14044));
  jand g13789(.dina(n14044), .dinb(n14039), .dout(n14045));
  jxor g13790(.dina(n14045), .dinb(n8729), .dout(n14046));
  jxor g13791(.dina(n14046), .dinb(n14038), .dout(n14047));
  jxor g13792(.dina(n14047), .dinb(n14021), .dout(n14048));
  jor  g13793(.dina(n8457), .dinb(n1879), .dout(n14049));
  jor  g13794(.dina(n8185), .dinb(n1637), .dout(n14050));
  jor  g13795(.dina(n8454), .dinb(n1881), .dout(n14051));
  jor  g13796(.dina(n8459), .dinb(n1759), .dout(n14052));
  jand g13797(.dina(n14052), .dinb(n14051), .dout(n14053));
  jand g13798(.dina(n14053), .dinb(n14050), .dout(n14054));
  jand g13799(.dina(n14054), .dinb(n14049), .dout(n14055));
  jxor g13800(.dina(n14055), .dinb(n7929), .dout(n14056));
  jxor g13801(.dina(n14056), .dinb(n14048), .dout(n14057));
  jxor g13802(.dina(n14057), .dinb(n14018), .dout(n14058));
  jor  g13803(.dina(n7660), .dinb(n2277), .dout(n14059));
  jor  g13804(.dina(n7415), .dinb(n2007), .dout(n14060));
  jor  g13805(.dina(n7662), .dinb(n2279), .dout(n14061));
  jor  g13806(.dina(n7657), .dinb(n2142), .dout(n14062));
  jand g13807(.dina(n14062), .dinb(n14061), .dout(n14063));
  jand g13808(.dina(n14063), .dinb(n14060), .dout(n14064));
  jand g13809(.dina(n14064), .dinb(n14059), .dout(n14065));
  jxor g13810(.dina(n14065), .dinb(n7166), .dout(n14066));
  jxor g13811(.dina(n14066), .dinb(n14058), .dout(n14067));
  jxor g13812(.dina(n14067), .dinb(n14015), .dout(n14068));
  jor  g13813(.dina(n6914), .dinb(n2711), .dout(n14069));
  jor  g13814(.dina(n6673), .dinb(n2415), .dout(n14070));
  jor  g13815(.dina(n6916), .dinb(n2713), .dout(n14071));
  jor  g13816(.dina(n6911), .dinb(n2563), .dout(n14072));
  jand g13817(.dina(n14072), .dinb(n14071), .dout(n14073));
  jand g13818(.dina(n14073), .dinb(n14070), .dout(n14074));
  jand g13819(.dina(n14074), .dinb(n14069), .dout(n14075));
  jxor g13820(.dina(n14075), .dinb(n6443), .dout(n14076));
  jxor g13821(.dina(n14076), .dinb(n14068), .dout(n14077));
  jxor g13822(.dina(n14077), .dinb(n14012), .dout(n14078));
  jor  g13823(.dina(n6207), .dinb(n3184), .dout(n14079));
  jor  g13824(.dina(n5975), .dinb(n2862), .dout(n14080));
  jor  g13825(.dina(n6210), .dinb(n3023), .dout(n14081));
  jor  g13826(.dina(n6205), .dinb(n3186), .dout(n14082));
  jand g13827(.dina(n14082), .dinb(n14081), .dout(n14083));
  jand g13828(.dina(n14083), .dinb(n14080), .dout(n14084));
  jand g13829(.dina(n14084), .dinb(n14079), .dout(n14085));
  jxor g13830(.dina(n14085), .dinb(n5759), .dout(n14086));
  jxor g13831(.dina(n14086), .dinb(n14078), .dout(n14087));
  jxor g13832(.dina(n14087), .dinb(n14009), .dout(n14088));
  jor  g13833(.dina(n5537), .dinb(n3696), .dout(n14089));
  jor  g13834(.dina(n5315), .dinb(n3348), .dout(n14090));
  jor  g13835(.dina(n5539), .dinb(n3698), .dout(n14091));
  jor  g13836(.dina(n5534), .dinb(n3522), .dout(n14092));
  jand g13837(.dina(n14092), .dinb(n14091), .dout(n14093));
  jand g13838(.dina(n14093), .dinb(n14090), .dout(n14094));
  jand g13839(.dina(n14094), .dinb(n14089), .dout(n14095));
  jxor g13840(.dina(n14095), .dinb(n5111), .dout(n14096));
  jxor g13841(.dina(n14096), .dinb(n14088), .dout(n14097));
  jxor g13842(.dina(n14097), .dinb(n14006), .dout(n14098));
  jor  g13843(.dina(n4902), .dinb(n4247), .dout(n14099));
  jor  g13844(.dina(n4696), .dinb(n3873), .dout(n14100));
  jor  g13845(.dina(n4904), .dinb(n4060), .dout(n14101));
  jor  g13846(.dina(n4899), .dinb(n4249), .dout(n14102));
  jand g13847(.dina(n14102), .dinb(n14101), .dout(n14103));
  jand g13848(.dina(n14103), .dinb(n14100), .dout(n14104));
  jand g13849(.dina(n14104), .dinb(n14099), .dout(n14105));
  jxor g13850(.dina(n14105), .dinb(n4505), .dout(n14106));
  jxor g13851(.dina(n14106), .dinb(n14098), .dout(n14107));
  jxor g13852(.dina(n14107), .dinb(n14003), .dout(n14108));
  jor  g13853(.dina(n4837), .dinb(n4305), .dout(n14109));
  jor  g13854(.dina(n4116), .dinb(n4437), .dout(n14110));
  jor  g13855(.dina(n4303), .dinb(n4839), .dout(n14111));
  jor  g13856(.dina(n4308), .dinb(n4637), .dout(n14112));
  jand g13857(.dina(n14112), .dinb(n14111), .dout(n14113));
  jand g13858(.dina(n14113), .dinb(n14110), .dout(n14114));
  jand g13859(.dina(n14114), .dinb(n14109), .dout(n14115));
  jxor g13860(.dina(n14115), .dinb(n3938), .dout(n14116));
  jxor g13861(.dina(n14116), .dinb(n14108), .dout(n14117));
  jxor g13862(.dina(n14117), .dinb(n14000), .dout(n14118));
  jor  g13863(.dina(n5467), .dinb(n3751), .dout(n14119));
  jor  g13864(.dina(n3574), .dinb(n5040), .dout(n14120));
  jor  g13865(.dina(n3754), .dinb(n5253), .dout(n14121));
  jor  g13866(.dina(n3749), .dinb(n5469), .dout(n14122));
  jand g13867(.dina(n14122), .dinb(n14121), .dout(n14123));
  jand g13868(.dina(n14123), .dinb(n14120), .dout(n14124));
  jand g13869(.dina(n14124), .dinb(n14119), .dout(n14125));
  jxor g13870(.dina(n14125), .dinb(n3410), .dout(n14126));
  jxor g13871(.dina(n14126), .dinb(n14118), .dout(n14127));
  jxor g13872(.dina(n14127), .dinb(n13997), .dout(n14128));
  jxor g13873(.dina(n14128), .dinb(n13985), .dout(n14129));
  jxor g13874(.dina(n14129), .dinb(n13973), .dout(n14130));
  jxor g13875(.dina(n14130), .dinb(n13961), .dout(n14131));
  jxor g13876(.dina(n14131), .dinb(n13949), .dout(n14132));
  jand g13877(.dina(n13898), .dinb(n13890), .dout(n14133));
  jand g13878(.dina(n13899), .dinb(n13887), .dout(n14134));
  jor  g13879(.dina(n14134), .dinb(n14133), .dout(n14135));
  jor  g13880(.dina(n10049), .dinb(n1248), .dout(n14136));
  jor  g13881(.dina(n1147), .dinb(n9475), .dout(n14137));
  jor  g13882(.dina(n1251), .dinb(n9759), .dout(n14138));
  jor  g13883(.dina(n1246), .dinb(n10051), .dout(n14139));
  jand g13884(.dina(n14139), .dinb(n14138), .dout(n14140));
  jand g13885(.dina(n14140), .dinb(n14137), .dout(n14141));
  jand g13886(.dina(n14141), .dinb(n14136), .dout(n14142));
  jxor g13887(.dina(n14142), .dinb(n1061), .dout(n14143));
  jxor g13888(.dina(n14143), .dinb(n14135), .dout(n14144));
  jxor g13889(.dina(n14144), .dinb(n14132), .dout(n14145));
  jand g13890(.dina(n13911), .dinb(n13903), .dout(n14146));
  jand g13891(.dina(n13912), .dinb(n13900), .dout(n14147));
  jor  g13892(.dina(n14147), .dinb(n14146), .dout(n14148));
  jnot g13893(.din(n14148), .dout(n14149));
  jand g13894(.dina(n881), .dinb(b63 ), .dout(n14150));
  jand g13895(.dina(n10832), .dinb(n802), .dout(n14151));
  jor  g13896(.dina(n14151), .dinb(n14150), .dout(n14152));
  jxor g13897(.dina(n14152), .dinb(n810), .dout(n14153));
  jxor g13898(.dina(n14153), .dinb(n14149), .dout(n14154));
  jxor g13899(.dina(n14154), .dinb(n14145), .dout(n14155));
  jxor g13900(.dina(n14155), .dinb(n13937), .dout(n14156));
  jnot g13901(.din(n14156), .dout(n14157));
  jxor g13902(.dina(n14157), .dinb(n13932), .dout(f77 ));
  jor  g13903(.dina(n14153), .dinb(n14149), .dout(n14159));
  jand g13904(.dina(n14154), .dinb(n14145), .dout(n14160));
  jnot g13905(.din(n14160), .dout(n14161));
  jand g13906(.dina(n14161), .dinb(n14159), .dout(n14162));
  jnot g13907(.din(n14162), .dout(n14163));
  jand g13908(.dina(n13948), .dinb(n13940), .dout(n14164));
  jand g13909(.dina(n14131), .dinb(n13949), .dout(n14165));
  jor  g13910(.dina(n14165), .dinb(n14164), .dout(n14166));
  jor  g13911(.dina(n9473), .dinb(n1569), .dout(n14167));
  jor  g13912(.dina(n1453), .dinb(n8920), .dout(n14168));
  jor  g13913(.dina(n1566), .dinb(n9195), .dout(n14169));
  jor  g13914(.dina(n1571), .dinb(n9475), .dout(n14170));
  jand g13915(.dina(n14170), .dinb(n14169), .dout(n14171));
  jand g13916(.dina(n14171), .dinb(n14168), .dout(n14172));
  jand g13917(.dina(n14172), .dinb(n14167), .dout(n14173));
  jxor g13918(.dina(n14173), .dinb(n1351), .dout(n14174));
  jxor g13919(.dina(n14174), .dinb(n14166), .dout(n14175));
  jand g13920(.dina(n13960), .dinb(n13952), .dout(n14176));
  jand g13921(.dina(n14130), .dinb(n13961), .dout(n14177));
  jor  g13922(.dina(n14177), .dinb(n14176), .dout(n14178));
  jor  g13923(.dina(n8642), .dinb(n1921), .dout(n14179));
  jor  g13924(.dina(n1806), .dinb(n8111), .dout(n14180));
  jor  g13925(.dina(n1923), .dinb(n8644), .dout(n14181));
  jor  g13926(.dina(n1918), .dinb(n8378), .dout(n14182));
  jand g13927(.dina(n14182), .dinb(n14181), .dout(n14183));
  jand g13928(.dina(n14183), .dinb(n14180), .dout(n14184));
  jand g13929(.dina(n14184), .dinb(n14179), .dout(n14185));
  jxor g13930(.dina(n14185), .dinb(n1687), .dout(n14186));
  jxor g13931(.dina(n14186), .dinb(n14178), .dout(n14187));
  jand g13932(.dina(n13972), .dinb(n13964), .dout(n14188));
  jand g13933(.dina(n14129), .dinb(n13973), .dout(n14189));
  jor  g13934(.dina(n14189), .dinb(n14188), .dout(n14190));
  jor  g13935(.dina(n7844), .dinb(n2324), .dout(n14191));
  jor  g13936(.dina(n2186), .dinb(n7338), .dout(n14192));
  jor  g13937(.dina(n2326), .dinb(n7846), .dout(n14193));
  jor  g13938(.dina(n2321), .dinb(n7590), .dout(n14194));
  jand g13939(.dina(n14194), .dinb(n14193), .dout(n14195));
  jand g13940(.dina(n14195), .dinb(n14192), .dout(n14196));
  jand g13941(.dina(n14196), .dinb(n14191), .dout(n14197));
  jxor g13942(.dina(n14197), .dinb(n2057), .dout(n14198));
  jxor g13943(.dina(n14198), .dinb(n14190), .dout(n14199));
  jand g13944(.dina(n13984), .dinb(n13976), .dout(n14200));
  jand g13945(.dina(n14128), .dinb(n13985), .dout(n14201));
  jor  g13946(.dina(n14201), .dinb(n14200), .dout(n14202));
  jor  g13947(.dina(n7084), .dinb(n2764), .dout(n14203));
  jor  g13948(.dina(n2609), .dinb(n6605), .dout(n14204));
  jor  g13949(.dina(n2761), .dinb(n7086), .dout(n14205));
  jor  g13950(.dina(n2766), .dinb(n6846), .dout(n14206));
  jand g13951(.dina(n14206), .dinb(n14205), .dout(n14207));
  jand g13952(.dina(n14207), .dinb(n14204), .dout(n14208));
  jand g13953(.dina(n14208), .dinb(n14203), .dout(n14209));
  jxor g13954(.dina(n14209), .dinb(n2468), .dout(n14210));
  jxor g13955(.dina(n14210), .dinb(n14202), .dout(n14211));
  jand g13956(.dina(n14117), .dinb(n14000), .dout(n14212));
  jand g13957(.dina(n14126), .dinb(n14118), .dout(n14213));
  jor  g13958(.dina(n14213), .dinb(n14212), .dout(n14214));
  jand g13959(.dina(n14107), .dinb(n14003), .dout(n14215));
  jand g13960(.dina(n14116), .dinb(n14108), .dout(n14216));
  jor  g13961(.dina(n14216), .dinb(n14215), .dout(n14217));
  jand g13962(.dina(n14097), .dinb(n14006), .dout(n14218));
  jand g13963(.dina(n14106), .dinb(n14098), .dout(n14219));
  jor  g13964(.dina(n14219), .dinb(n14218), .dout(n14220));
  jand g13965(.dina(n14087), .dinb(n14009), .dout(n14221));
  jand g13966(.dina(n14096), .dinb(n14088), .dout(n14222));
  jor  g13967(.dina(n14222), .dinb(n14221), .dout(n14223));
  jand g13968(.dina(n14077), .dinb(n14012), .dout(n14224));
  jand g13969(.dina(n14086), .dinb(n14078), .dout(n14225));
  jor  g13970(.dina(n14225), .dinb(n14224), .dout(n14226));
  jand g13971(.dina(n14067), .dinb(n14015), .dout(n14227));
  jand g13972(.dina(n14076), .dinb(n14068), .dout(n14228));
  jor  g13973(.dina(n14228), .dinb(n14227), .dout(n14229));
  jand g13974(.dina(n14057), .dinb(n14018), .dout(n14230));
  jand g13975(.dina(n14066), .dinb(n14058), .dout(n14231));
  jor  g13976(.dina(n14231), .dinb(n14230), .dout(n14232));
  jand g13977(.dina(n14047), .dinb(n14021), .dout(n14233));
  jand g13978(.dina(n14056), .dinb(n14048), .dout(n14234));
  jor  g13979(.dina(n14234), .dinb(n14233), .dout(n14235));
  jand g13980(.dina(n14037), .dinb(n14024), .dout(n14236));
  jand g13981(.dina(n14046), .dinb(n14038), .dout(n14237));
  jor  g13982(.dina(n14237), .dinb(n14236), .dout(n14238));
  jand g13983(.dina(n14027), .dinb(n13761), .dout(n14239));
  jand g13984(.dina(n14036), .dinb(n14028), .dout(n14240));
  jor  g13985(.dina(n14240), .dinb(n14239), .dout(n14241));
  jand g13986(.dina(n10594), .dinb(b14 ), .dout(n14242));
  jand g13987(.dina(n10129), .dinb(b15 ), .dout(n14243));
  jor  g13988(.dina(n14243), .dinb(n14242), .dout(n14244));
  jxor g13989(.dina(n14244), .dinb(n810), .dout(n14245));
  jxor g13990(.dina(n14245), .dinb(n13760), .dout(n14246));
  jor  g13991(.dina(n10134), .dinb(n1305), .dout(n14247));
  jor  g13992(.dina(n9849), .dinb(n1114), .dout(n14248));
  jor  g13993(.dina(n10137), .dinb(n1211), .dout(n14249));
  jor  g13994(.dina(n10132), .dinb(n1307), .dout(n14250));
  jand g13995(.dina(n14250), .dinb(n14249), .dout(n14251));
  jand g13996(.dina(n14251), .dinb(n14248), .dout(n14252));
  jand g13997(.dina(n14252), .dinb(n14247), .dout(n14253));
  jxor g13998(.dina(n14253), .dinb(n9559), .dout(n14254));
  jxor g13999(.dina(n14254), .dinb(n14246), .dout(n14255));
  jxor g14000(.dina(n14255), .dinb(n14241), .dout(n14256));
  jor  g14001(.dina(n9271), .dinb(n1635), .dout(n14257));
  jor  g14002(.dina(n9003), .dinb(n1416), .dout(n14258));
  jor  g14003(.dina(n9268), .dinb(n1637), .dout(n14259));
  jor  g14004(.dina(n9273), .dinb(n1527), .dout(n14260));
  jand g14005(.dina(n14260), .dinb(n14259), .dout(n14261));
  jand g14006(.dina(n14261), .dinb(n14258), .dout(n14262));
  jand g14007(.dina(n14262), .dinb(n14257), .dout(n14263));
  jxor g14008(.dina(n14263), .dinb(n8729), .dout(n14264));
  jxor g14009(.dina(n14264), .dinb(n14256), .dout(n14265));
  jxor g14010(.dina(n14265), .dinb(n14238), .dout(n14266));
  jor  g14011(.dina(n8457), .dinb(n2005), .dout(n14267));
  jor  g14012(.dina(n8185), .dinb(n1759), .dout(n14268));
  jor  g14013(.dina(n8454), .dinb(n2007), .dout(n14269));
  jor  g14014(.dina(n8459), .dinb(n1881), .dout(n14270));
  jand g14015(.dina(n14270), .dinb(n14269), .dout(n14271));
  jand g14016(.dina(n14271), .dinb(n14268), .dout(n14272));
  jand g14017(.dina(n14272), .dinb(n14267), .dout(n14273));
  jxor g14018(.dina(n14273), .dinb(n7929), .dout(n14274));
  jxor g14019(.dina(n14274), .dinb(n14266), .dout(n14275));
  jxor g14020(.dina(n14275), .dinb(n14235), .dout(n14276));
  jor  g14021(.dina(n7660), .dinb(n2413), .dout(n14277));
  jor  g14022(.dina(n7415), .dinb(n2142), .dout(n14278));
  jor  g14023(.dina(n7662), .dinb(n2415), .dout(n14279));
  jor  g14024(.dina(n7657), .dinb(n2279), .dout(n14280));
  jand g14025(.dina(n14280), .dinb(n14279), .dout(n14281));
  jand g14026(.dina(n14281), .dinb(n14278), .dout(n14282));
  jand g14027(.dina(n14282), .dinb(n14277), .dout(n14283));
  jxor g14028(.dina(n14283), .dinb(n7166), .dout(n14284));
  jxor g14029(.dina(n14284), .dinb(n14276), .dout(n14285));
  jxor g14030(.dina(n14285), .dinb(n14232), .dout(n14286));
  jor  g14031(.dina(n6914), .dinb(n2860), .dout(n14287));
  jor  g14032(.dina(n6673), .dinb(n2563), .dout(n14288));
  jor  g14033(.dina(n6911), .dinb(n2713), .dout(n14289));
  jor  g14034(.dina(n6916), .dinb(n2862), .dout(n14290));
  jand g14035(.dina(n14290), .dinb(n14289), .dout(n14291));
  jand g14036(.dina(n14291), .dinb(n14288), .dout(n14292));
  jand g14037(.dina(n14292), .dinb(n14287), .dout(n14293));
  jxor g14038(.dina(n14293), .dinb(n6443), .dout(n14294));
  jxor g14039(.dina(n14294), .dinb(n14286), .dout(n14295));
  jxor g14040(.dina(n14295), .dinb(n14229), .dout(n14296));
  jor  g14041(.dina(n6207), .dinb(n3346), .dout(n14297));
  jor  g14042(.dina(n5975), .dinb(n3023), .dout(n14298));
  jor  g14043(.dina(n6205), .dinb(n3348), .dout(n14299));
  jor  g14044(.dina(n6210), .dinb(n3186), .dout(n14300));
  jand g14045(.dina(n14300), .dinb(n14299), .dout(n14301));
  jand g14046(.dina(n14301), .dinb(n14298), .dout(n14302));
  jand g14047(.dina(n14302), .dinb(n14297), .dout(n14303));
  jxor g14048(.dina(n14303), .dinb(n5759), .dout(n14304));
  jxor g14049(.dina(n14304), .dinb(n14296), .dout(n14305));
  jxor g14050(.dina(n14305), .dinb(n14226), .dout(n14306));
  jor  g14051(.dina(n5537), .dinb(n3871), .dout(n14307));
  jor  g14052(.dina(n5315), .dinb(n3522), .dout(n14308));
  jor  g14053(.dina(n5539), .dinb(n3873), .dout(n14309));
  jor  g14054(.dina(n5534), .dinb(n3698), .dout(n14310));
  jand g14055(.dina(n14310), .dinb(n14309), .dout(n14311));
  jand g14056(.dina(n14311), .dinb(n14308), .dout(n14312));
  jand g14057(.dina(n14312), .dinb(n14307), .dout(n14313));
  jxor g14058(.dina(n14313), .dinb(n5111), .dout(n14314));
  jxor g14059(.dina(n14314), .dinb(n14306), .dout(n14315));
  jxor g14060(.dina(n14315), .dinb(n14223), .dout(n14316));
  jor  g14061(.dina(n4902), .dinb(n4435), .dout(n14317));
  jor  g14062(.dina(n4696), .dinb(n4060), .dout(n14318));
  jor  g14063(.dina(n4899), .dinb(n4437), .dout(n14319));
  jor  g14064(.dina(n4904), .dinb(n4249), .dout(n14320));
  jand g14065(.dina(n14320), .dinb(n14319), .dout(n14321));
  jand g14066(.dina(n14321), .dinb(n14318), .dout(n14322));
  jand g14067(.dina(n14322), .dinb(n14317), .dout(n14323));
  jxor g14068(.dina(n14323), .dinb(n4505), .dout(n14324));
  jxor g14069(.dina(n14324), .dinb(n14316), .dout(n14325));
  jxor g14070(.dina(n14325), .dinb(n14220), .dout(n14326));
  jor  g14071(.dina(n5038), .dinb(n4305), .dout(n14327));
  jor  g14072(.dina(n4116), .dinb(n4637), .dout(n14328));
  jor  g14073(.dina(n4308), .dinb(n4839), .dout(n14329));
  jor  g14074(.dina(n4303), .dinb(n5040), .dout(n14330));
  jand g14075(.dina(n14330), .dinb(n14329), .dout(n14331));
  jand g14076(.dina(n14331), .dinb(n14328), .dout(n14332));
  jand g14077(.dina(n14332), .dinb(n14327), .dout(n14333));
  jxor g14078(.dina(n14333), .dinb(n3938), .dout(n14334));
  jxor g14079(.dina(n14334), .dinb(n14326), .dout(n14335));
  jxor g14080(.dina(n14335), .dinb(n14217), .dout(n14336));
  jor  g14081(.dina(n5683), .dinb(n3751), .dout(n14337));
  jor  g14082(.dina(n3574), .dinb(n5253), .dout(n14338));
  jor  g14083(.dina(n3754), .dinb(n5469), .dout(n14339));
  jor  g14084(.dina(n3749), .dinb(n5685), .dout(n14340));
  jand g14085(.dina(n14340), .dinb(n14339), .dout(n14341));
  jand g14086(.dina(n14341), .dinb(n14338), .dout(n14342));
  jand g14087(.dina(n14342), .dinb(n14337), .dout(n14343));
  jxor g14088(.dina(n14343), .dinb(n3410), .dout(n14344));
  jxor g14089(.dina(n14344), .dinb(n14336), .dout(n14345));
  jxor g14090(.dina(n14345), .dinb(n14214), .dout(n14346));
  jand g14091(.dina(n13996), .dinb(n13988), .dout(n14347));
  jand g14092(.dina(n14127), .dinb(n13997), .dout(n14348));
  jor  g14093(.dina(n14348), .dinb(n14347), .dout(n14349));
  jor  g14094(.dina(n6364), .dinb(n3239), .dout(n14350));
  jor  g14095(.dina(n3072), .dinb(n5911), .dout(n14351));
  jor  g14096(.dina(n3242), .dinb(n6139), .dout(n14352));
  jor  g14097(.dina(n3237), .dinb(n6366), .dout(n14353));
  jand g14098(.dina(n14353), .dinb(n14352), .dout(n14354));
  jand g14099(.dina(n14354), .dinb(n14351), .dout(n14355));
  jand g14100(.dina(n14355), .dinb(n14350), .dout(n14356));
  jxor g14101(.dina(n14356), .dinb(n2918), .dout(n14357));
  jxor g14102(.dina(n14357), .dinb(n14349), .dout(n14358));
  jxor g14103(.dina(n14358), .dinb(n14346), .dout(n14359));
  jxor g14104(.dina(n14359), .dinb(n14211), .dout(n14360));
  jxor g14105(.dina(n14360), .dinb(n14199), .dout(n14361));
  jxor g14106(.dina(n14361), .dinb(n14187), .dout(n14362));
  jxor g14107(.dina(n14362), .dinb(n14175), .dout(n14363));
  jand g14108(.dina(n14143), .dinb(n14135), .dout(n14364));
  jand g14109(.dina(n14144), .dinb(n14132), .dout(n14365));
  jor  g14110(.dina(n14365), .dinb(n14364), .dout(n14366));
  jor  g14111(.dina(n10521), .dinb(n1248), .dout(n14367));
  jor  g14112(.dina(n1147), .dinb(n9759), .dout(n14368));
  jor  g14113(.dina(n1246), .dinb(n10523), .dout(n14369));
  jor  g14114(.dina(n1251), .dinb(n10051), .dout(n14370));
  jand g14115(.dina(n14370), .dinb(n14369), .dout(n14371));
  jand g14116(.dina(n14371), .dinb(n14368), .dout(n14372));
  jand g14117(.dina(n14372), .dinb(n14367), .dout(n14373));
  jxor g14118(.dina(n14373), .dinb(n1061), .dout(n14374));
  jxor g14119(.dina(n14374), .dinb(n14366), .dout(n14375));
  jxor g14120(.dina(n14375), .dinb(n14363), .dout(n14376));
  jxor g14121(.dina(n14376), .dinb(n14163), .dout(n14377));
  jnot g14122(.din(n14377), .dout(n14378));
  jand g14123(.dina(n14155), .dinb(n13937), .dout(n14379));
  jnot g14124(.din(n14379), .dout(n14380));
  jor  g14125(.dina(n14157), .dinb(n13932), .dout(n14381));
  jand g14126(.dina(n14381), .dinb(n14380), .dout(n14382));
  jxor g14127(.dina(n14382), .dinb(n14378), .dout(f78 ));
  jand g14128(.dina(n14374), .dinb(n14366), .dout(n14384));
  jand g14129(.dina(n14375), .dinb(n14363), .dout(n14385));
  jor  g14130(.dina(n14385), .dinb(n14384), .dout(n14386));
  jand g14131(.dina(n14174), .dinb(n14166), .dout(n14387));
  jand g14132(.dina(n14362), .dinb(n14175), .dout(n14388));
  jor  g14133(.dina(n14388), .dinb(n14387), .dout(n14389));
  jor  g14134(.dina(n10813), .dinb(n1248), .dout(n14390));
  jor  g14135(.dina(n1147), .dinb(n10051), .dout(n14391));
  jor  g14136(.dina(n1251), .dinb(n10523), .dout(n14392));
  jand g14137(.dina(n14392), .dinb(n14391), .dout(n14393));
  jand g14138(.dina(n14393), .dinb(n14390), .dout(n14394));
  jxor g14139(.dina(n14394), .dinb(n1061), .dout(n14395));
  jxor g14140(.dina(n14395), .dinb(n14389), .dout(n14396));
  jand g14141(.dina(n14186), .dinb(n14178), .dout(n14397));
  jand g14142(.dina(n14361), .dinb(n14187), .dout(n14398));
  jor  g14143(.dina(n14398), .dinb(n14397), .dout(n14399));
  jor  g14144(.dina(n9757), .dinb(n1569), .dout(n14400));
  jor  g14145(.dina(n1453), .dinb(n9195), .dout(n14401));
  jor  g14146(.dina(n1566), .dinb(n9475), .dout(n14402));
  jor  g14147(.dina(n1571), .dinb(n9759), .dout(n14403));
  jand g14148(.dina(n14403), .dinb(n14402), .dout(n14404));
  jand g14149(.dina(n14404), .dinb(n14401), .dout(n14405));
  jand g14150(.dina(n14405), .dinb(n14400), .dout(n14406));
  jxor g14151(.dina(n14406), .dinb(n1351), .dout(n14407));
  jxor g14152(.dina(n14407), .dinb(n14399), .dout(n14408));
  jand g14153(.dina(n14198), .dinb(n14190), .dout(n14409));
  jand g14154(.dina(n14360), .dinb(n14199), .dout(n14410));
  jor  g14155(.dina(n14410), .dinb(n14409), .dout(n14411));
  jor  g14156(.dina(n8918), .dinb(n1921), .dout(n14412));
  jor  g14157(.dina(n1806), .dinb(n8378), .dout(n14413));
  jor  g14158(.dina(n1918), .dinb(n8644), .dout(n14414));
  jor  g14159(.dina(n1923), .dinb(n8920), .dout(n14415));
  jand g14160(.dina(n14415), .dinb(n14414), .dout(n14416));
  jand g14161(.dina(n14416), .dinb(n14413), .dout(n14417));
  jand g14162(.dina(n14417), .dinb(n14412), .dout(n14418));
  jxor g14163(.dina(n14418), .dinb(n1687), .dout(n14419));
  jxor g14164(.dina(n14419), .dinb(n14411), .dout(n14420));
  jand g14165(.dina(n14210), .dinb(n14202), .dout(n14421));
  jand g14166(.dina(n14359), .dinb(n14211), .dout(n14422));
  jor  g14167(.dina(n14422), .dinb(n14421), .dout(n14423));
  jor  g14168(.dina(n8109), .dinb(n2324), .dout(n14424));
  jor  g14169(.dina(n2186), .dinb(n7590), .dout(n14425));
  jor  g14170(.dina(n2321), .dinb(n7846), .dout(n14426));
  jor  g14171(.dina(n2326), .dinb(n8111), .dout(n14427));
  jand g14172(.dina(n14427), .dinb(n14426), .dout(n14428));
  jand g14173(.dina(n14428), .dinb(n14425), .dout(n14429));
  jand g14174(.dina(n14429), .dinb(n14424), .dout(n14430));
  jxor g14175(.dina(n14430), .dinb(n2057), .dout(n14431));
  jxor g14176(.dina(n14431), .dinb(n14423), .dout(n14432));
  jand g14177(.dina(n14357), .dinb(n14349), .dout(n14433));
  jand g14178(.dina(n14358), .dinb(n14346), .dout(n14434));
  jor  g14179(.dina(n14434), .dinb(n14433), .dout(n14435));
  jor  g14180(.dina(n7336), .dinb(n2764), .dout(n14436));
  jor  g14181(.dina(n2609), .dinb(n6846), .dout(n14437));
  jor  g14182(.dina(n2761), .dinb(n7338), .dout(n14438));
  jor  g14183(.dina(n2766), .dinb(n7086), .dout(n14439));
  jand g14184(.dina(n14439), .dinb(n14438), .dout(n14440));
  jand g14185(.dina(n14440), .dinb(n14437), .dout(n14441));
  jand g14186(.dina(n14441), .dinb(n14436), .dout(n14442));
  jxor g14187(.dina(n14442), .dinb(n2468), .dout(n14443));
  jxor g14188(.dina(n14443), .dinb(n14435), .dout(n14444));
  jand g14189(.dina(n14344), .dinb(n14336), .dout(n14445));
  jand g14190(.dina(n14345), .dinb(n14214), .dout(n14446));
  jor  g14191(.dina(n14446), .dinb(n14445), .dout(n14447));
  jor  g14192(.dina(n6603), .dinb(n3239), .dout(n14448));
  jor  g14193(.dina(n3072), .dinb(n6139), .dout(n14449));
  jor  g14194(.dina(n3237), .dinb(n6605), .dout(n14450));
  jor  g14195(.dina(n3242), .dinb(n6366), .dout(n14451));
  jand g14196(.dina(n14451), .dinb(n14450), .dout(n14452));
  jand g14197(.dina(n14452), .dinb(n14449), .dout(n14453));
  jand g14198(.dina(n14453), .dinb(n14448), .dout(n14454));
  jxor g14199(.dina(n14454), .dinb(n2918), .dout(n14455));
  jxor g14200(.dina(n14455), .dinb(n14447), .dout(n14456));
  jand g14201(.dina(n14334), .dinb(n14326), .dout(n14457));
  jand g14202(.dina(n14335), .dinb(n14217), .dout(n14458));
  jor  g14203(.dina(n14458), .dinb(n14457), .dout(n14459));
  jand g14204(.dina(n14324), .dinb(n14316), .dout(n14460));
  jand g14205(.dina(n14325), .dinb(n14220), .dout(n14461));
  jor  g14206(.dina(n14461), .dinb(n14460), .dout(n14462));
  jand g14207(.dina(n14314), .dinb(n14306), .dout(n14463));
  jand g14208(.dina(n14315), .dinb(n14223), .dout(n14464));
  jor  g14209(.dina(n14464), .dinb(n14463), .dout(n14465));
  jand g14210(.dina(n14304), .dinb(n14296), .dout(n14466));
  jand g14211(.dina(n14305), .dinb(n14226), .dout(n14467));
  jor  g14212(.dina(n14467), .dinb(n14466), .dout(n14468));
  jand g14213(.dina(n14294), .dinb(n14286), .dout(n14469));
  jand g14214(.dina(n14295), .dinb(n14229), .dout(n14470));
  jor  g14215(.dina(n14470), .dinb(n14469), .dout(n14471));
  jand g14216(.dina(n14264), .dinb(n14256), .dout(n14472));
  jand g14217(.dina(n14265), .dinb(n14238), .dout(n14473));
  jor  g14218(.dina(n14473), .dinb(n14472), .dout(n14474));
  jand g14219(.dina(n14254), .dinb(n14246), .dout(n14475));
  jand g14220(.dina(n14255), .dinb(n14241), .dout(n14476));
  jor  g14221(.dina(n14476), .dinb(n14475), .dout(n14477));
  jand g14222(.dina(n10594), .dinb(b15 ), .dout(n14478));
  jand g14223(.dina(n10129), .dinb(b16 ), .dout(n14479));
  jor  g14224(.dina(n14479), .dinb(n14478), .dout(n14480));
  jnot g14225(.din(n14480), .dout(n14481));
  jand g14226(.dina(n14244), .dinb(n810), .dout(n14482));
  jand g14227(.dina(n14245), .dinb(n13760), .dout(n14483));
  jor  g14228(.dina(n14483), .dinb(n14482), .dout(n14484));
  jxor g14229(.dina(n14484), .dinb(n14481), .dout(n14485));
  jor  g14230(.dina(n10134), .dinb(n1414), .dout(n14486));
  jor  g14231(.dina(n9849), .dinb(n1211), .dout(n14487));
  jor  g14232(.dina(n10137), .dinb(n1307), .dout(n14488));
  jor  g14233(.dina(n10132), .dinb(n1416), .dout(n14489));
  jand g14234(.dina(n14489), .dinb(n14488), .dout(n14490));
  jand g14235(.dina(n14490), .dinb(n14487), .dout(n14491));
  jand g14236(.dina(n14491), .dinb(n14486), .dout(n14492));
  jxor g14237(.dina(n14492), .dinb(n9559), .dout(n14493));
  jxor g14238(.dina(n14493), .dinb(n14485), .dout(n14494));
  jxor g14239(.dina(n14494), .dinb(n14477), .dout(n14495));
  jor  g14240(.dina(n9271), .dinb(n1757), .dout(n14496));
  jor  g14241(.dina(n9003), .dinb(n1527), .dout(n14497));
  jor  g14242(.dina(n9273), .dinb(n1637), .dout(n14498));
  jor  g14243(.dina(n9268), .dinb(n1759), .dout(n14499));
  jand g14244(.dina(n14499), .dinb(n14498), .dout(n14500));
  jand g14245(.dina(n14500), .dinb(n14497), .dout(n14501));
  jand g14246(.dina(n14501), .dinb(n14496), .dout(n14502));
  jxor g14247(.dina(n14502), .dinb(n8729), .dout(n14503));
  jxor g14248(.dina(n14503), .dinb(n14495), .dout(n14504));
  jxor g14249(.dina(n14504), .dinb(n14474), .dout(n14505));
  jor  g14250(.dina(n8457), .dinb(n2140), .dout(n14506));
  jor  g14251(.dina(n8185), .dinb(n1881), .dout(n14507));
  jor  g14252(.dina(n8454), .dinb(n2142), .dout(n14508));
  jor  g14253(.dina(n8459), .dinb(n2007), .dout(n14509));
  jand g14254(.dina(n14509), .dinb(n14508), .dout(n14510));
  jand g14255(.dina(n14510), .dinb(n14507), .dout(n14511));
  jand g14256(.dina(n14511), .dinb(n14506), .dout(n14512));
  jxor g14257(.dina(n14512), .dinb(n7929), .dout(n14513));
  jxor g14258(.dina(n14513), .dinb(n14505), .dout(n14514));
  jnot g14259(.din(n14266), .dout(n14515));
  jnot g14260(.din(n14274), .dout(n14516));
  jand g14261(.dina(n14516), .dinb(n14515), .dout(n14517));
  jnot g14262(.din(n14517), .dout(n14518));
  jand g14263(.dina(n14274), .dinb(n14266), .dout(n14519));
  jor  g14264(.dina(n14519), .dinb(n14235), .dout(n14520));
  jand g14265(.dina(n14520), .dinb(n14518), .dout(n14521));
  jxor g14266(.dina(n14521), .dinb(n14514), .dout(n14522));
  jor  g14267(.dina(n7660), .dinb(n2561), .dout(n14523));
  jor  g14268(.dina(n7415), .dinb(n2279), .dout(n14524));
  jor  g14269(.dina(n7657), .dinb(n2415), .dout(n14525));
  jor  g14270(.dina(n7662), .dinb(n2563), .dout(n14526));
  jand g14271(.dina(n14526), .dinb(n14525), .dout(n14527));
  jand g14272(.dina(n14527), .dinb(n14524), .dout(n14528));
  jand g14273(.dina(n14528), .dinb(n14523), .dout(n14529));
  jxor g14274(.dina(n14529), .dinb(n7166), .dout(n14530));
  jxor g14275(.dina(n14530), .dinb(n14522), .dout(n14531));
  jand g14276(.dina(n14284), .dinb(n14276), .dout(n14532));
  jand g14277(.dina(n14285), .dinb(n14232), .dout(n14533));
  jor  g14278(.dina(n14533), .dinb(n14532), .dout(n14534));
  jxor g14279(.dina(n14534), .dinb(n14531), .dout(n14535));
  jor  g14280(.dina(n6914), .dinb(n3021), .dout(n14536));
  jor  g14281(.dina(n6673), .dinb(n2713), .dout(n14537));
  jor  g14282(.dina(n6916), .dinb(n3023), .dout(n14538));
  jor  g14283(.dina(n6911), .dinb(n2862), .dout(n14539));
  jand g14284(.dina(n14539), .dinb(n14538), .dout(n14540));
  jand g14285(.dina(n14540), .dinb(n14537), .dout(n14541));
  jand g14286(.dina(n14541), .dinb(n14536), .dout(n14542));
  jxor g14287(.dina(n14542), .dinb(n6443), .dout(n14543));
  jxor g14288(.dina(n14543), .dinb(n14535), .dout(n14544));
  jxor g14289(.dina(n14544), .dinb(n14471), .dout(n14545));
  jor  g14290(.dina(n6207), .dinb(n3520), .dout(n14546));
  jor  g14291(.dina(n5975), .dinb(n3186), .dout(n14547));
  jor  g14292(.dina(n6210), .dinb(n3348), .dout(n14548));
  jor  g14293(.dina(n6205), .dinb(n3522), .dout(n14549));
  jand g14294(.dina(n14549), .dinb(n14548), .dout(n14550));
  jand g14295(.dina(n14550), .dinb(n14547), .dout(n14551));
  jand g14296(.dina(n14551), .dinb(n14546), .dout(n14552));
  jxor g14297(.dina(n14552), .dinb(n5759), .dout(n14553));
  jxor g14298(.dina(n14553), .dinb(n14545), .dout(n14554));
  jxor g14299(.dina(n14554), .dinb(n14468), .dout(n14555));
  jor  g14300(.dina(n5537), .dinb(n4058), .dout(n14556));
  jor  g14301(.dina(n5315), .dinb(n3698), .dout(n14557));
  jor  g14302(.dina(n5539), .dinb(n4060), .dout(n14558));
  jor  g14303(.dina(n5534), .dinb(n3873), .dout(n14559));
  jand g14304(.dina(n14559), .dinb(n14558), .dout(n14560));
  jand g14305(.dina(n14560), .dinb(n14557), .dout(n14561));
  jand g14306(.dina(n14561), .dinb(n14556), .dout(n14562));
  jxor g14307(.dina(n14562), .dinb(n5111), .dout(n14563));
  jxor g14308(.dina(n14563), .dinb(n14555), .dout(n14564));
  jxor g14309(.dina(n14564), .dinb(n14465), .dout(n14565));
  jor  g14310(.dina(n4635), .dinb(n4902), .dout(n14566));
  jor  g14311(.dina(n4696), .dinb(n4249), .dout(n14567));
  jor  g14312(.dina(n4904), .dinb(n4437), .dout(n14568));
  jor  g14313(.dina(n4899), .dinb(n4637), .dout(n14569));
  jand g14314(.dina(n14569), .dinb(n14568), .dout(n14570));
  jand g14315(.dina(n14570), .dinb(n14567), .dout(n14571));
  jand g14316(.dina(n14571), .dinb(n14566), .dout(n14572));
  jxor g14317(.dina(n14572), .dinb(n4505), .dout(n14573));
  jxor g14318(.dina(n14573), .dinb(n14565), .dout(n14574));
  jxor g14319(.dina(n14574), .dinb(n14462), .dout(n14575));
  jor  g14320(.dina(n5251), .dinb(n4305), .dout(n14576));
  jor  g14321(.dina(n4116), .dinb(n4839), .dout(n14577));
  jor  g14322(.dina(n4308), .dinb(n5040), .dout(n14578));
  jor  g14323(.dina(n4303), .dinb(n5253), .dout(n14579));
  jand g14324(.dina(n14579), .dinb(n14578), .dout(n14580));
  jand g14325(.dina(n14580), .dinb(n14577), .dout(n14581));
  jand g14326(.dina(n14581), .dinb(n14576), .dout(n14582));
  jxor g14327(.dina(n14582), .dinb(n3938), .dout(n14583));
  jxor g14328(.dina(n14583), .dinb(n14575), .dout(n14584));
  jxor g14329(.dina(n14584), .dinb(n14459), .dout(n14585));
  jor  g14330(.dina(n5909), .dinb(n3751), .dout(n14586));
  jor  g14331(.dina(n3574), .dinb(n5469), .dout(n14587));
  jor  g14332(.dina(n3754), .dinb(n5685), .dout(n14588));
  jor  g14333(.dina(n3749), .dinb(n5911), .dout(n14589));
  jand g14334(.dina(n14589), .dinb(n14588), .dout(n14590));
  jand g14335(.dina(n14590), .dinb(n14587), .dout(n14591));
  jand g14336(.dina(n14591), .dinb(n14586), .dout(n14592));
  jxor g14337(.dina(n14592), .dinb(n3410), .dout(n14593));
  jxor g14338(.dina(n14593), .dinb(n14585), .dout(n14594));
  jxor g14339(.dina(n14594), .dinb(n14456), .dout(n14595));
  jxor g14340(.dina(n14595), .dinb(n14444), .dout(n14596));
  jxor g14341(.dina(n14596), .dinb(n14432), .dout(n14597));
  jxor g14342(.dina(n14597), .dinb(n14420), .dout(n14598));
  jxor g14343(.dina(n14598), .dinb(n14408), .dout(n14599));
  jxor g14344(.dina(n14599), .dinb(n14396), .dout(n14600));
  jxor g14345(.dina(n14600), .dinb(n14386), .dout(n14601));
  jnot g14346(.din(n14601), .dout(n14602));
  jand g14347(.dina(n14376), .dinb(n14163), .dout(n14603));
  jnot g14348(.din(n14603), .dout(n14604));
  jor  g14349(.dina(n14382), .dinb(n14378), .dout(n14605));
  jand g14350(.dina(n14605), .dinb(n14604), .dout(n14606));
  jxor g14351(.dina(n14606), .dinb(n14602), .dout(f79 ));
  jand g14352(.dina(n14600), .dinb(n14386), .dout(n14608));
  jnot g14353(.din(n14608), .dout(n14609));
  jor  g14354(.dina(n14606), .dinb(n14602), .dout(n14610));
  jand g14355(.dina(n14610), .dinb(n14609), .dout(n14611));
  jand g14356(.dina(n14395), .dinb(n14389), .dout(n14612));
  jand g14357(.dina(n14599), .dinb(n14396), .dout(n14613));
  jor  g14358(.dina(n14613), .dinb(n14612), .dout(n14614));
  jand g14359(.dina(n14419), .dinb(n14411), .dout(n14615));
  jand g14360(.dina(n14597), .dinb(n14420), .dout(n14616));
  jor  g14361(.dina(n14616), .dinb(n14615), .dout(n14617));
  jor  g14362(.dina(n10049), .dinb(n1569), .dout(n14618));
  jor  g14363(.dina(n1453), .dinb(n9475), .dout(n14619));
  jor  g14364(.dina(n1571), .dinb(n10051), .dout(n14620));
  jor  g14365(.dina(n1566), .dinb(n9759), .dout(n14621));
  jand g14366(.dina(n14621), .dinb(n14620), .dout(n14622));
  jand g14367(.dina(n14622), .dinb(n14619), .dout(n14623));
  jand g14368(.dina(n14623), .dinb(n14618), .dout(n14624));
  jxor g14369(.dina(n14624), .dinb(n1351), .dout(n14625));
  jxor g14370(.dina(n14625), .dinb(n14617), .dout(n14626));
  jand g14371(.dina(n14443), .dinb(n14435), .dout(n14627));
  jand g14372(.dina(n14595), .dinb(n14444), .dout(n14628));
  jor  g14373(.dina(n14628), .dinb(n14627), .dout(n14629));
  jor  g14374(.dina(n8376), .dinb(n2324), .dout(n14630));
  jor  g14375(.dina(n2186), .dinb(n7846), .dout(n14631));
  jor  g14376(.dina(n2321), .dinb(n8111), .dout(n14632));
  jor  g14377(.dina(n2326), .dinb(n8378), .dout(n14633));
  jand g14378(.dina(n14633), .dinb(n14632), .dout(n14634));
  jand g14379(.dina(n14634), .dinb(n14631), .dout(n14635));
  jand g14380(.dina(n14635), .dinb(n14630), .dout(n14636));
  jxor g14381(.dina(n14636), .dinb(n2057), .dout(n14637));
  jxor g14382(.dina(n14637), .dinb(n14629), .dout(n14638));
  jand g14383(.dina(n14455), .dinb(n14447), .dout(n14639));
  jand g14384(.dina(n14594), .dinb(n14456), .dout(n14640));
  jor  g14385(.dina(n14640), .dinb(n14639), .dout(n14641));
  jor  g14386(.dina(n7588), .dinb(n2764), .dout(n14642));
  jor  g14387(.dina(n2609), .dinb(n7086), .dout(n14643));
  jor  g14388(.dina(n2761), .dinb(n7590), .dout(n14644));
  jor  g14389(.dina(n2766), .dinb(n7338), .dout(n14645));
  jand g14390(.dina(n14645), .dinb(n14644), .dout(n14646));
  jand g14391(.dina(n14646), .dinb(n14643), .dout(n14647));
  jand g14392(.dina(n14647), .dinb(n14642), .dout(n14648));
  jxor g14393(.dina(n14648), .dinb(n2468), .dout(n14649));
  jxor g14394(.dina(n14649), .dinb(n14641), .dout(n14650));
  jand g14395(.dina(n14584), .dinb(n14459), .dout(n14651));
  jand g14396(.dina(n14593), .dinb(n14585), .dout(n14652));
  jor  g14397(.dina(n14652), .dinb(n14651), .dout(n14653));
  jor  g14398(.dina(n6844), .dinb(n3239), .dout(n14654));
  jor  g14399(.dina(n3072), .dinb(n6366), .dout(n14655));
  jor  g14400(.dina(n3237), .dinb(n6846), .dout(n14656));
  jor  g14401(.dina(n3242), .dinb(n6605), .dout(n14657));
  jand g14402(.dina(n14657), .dinb(n14656), .dout(n14658));
  jand g14403(.dina(n14658), .dinb(n14655), .dout(n14659));
  jand g14404(.dina(n14659), .dinb(n14654), .dout(n14660));
  jxor g14405(.dina(n14660), .dinb(n2918), .dout(n14661));
  jxor g14406(.dina(n14661), .dinb(n14653), .dout(n14662));
  jand g14407(.dina(n14574), .dinb(n14462), .dout(n14663));
  jand g14408(.dina(n14583), .dinb(n14575), .dout(n14664));
  jor  g14409(.dina(n14664), .dinb(n14663), .dout(n14665));
  jand g14410(.dina(n14564), .dinb(n14465), .dout(n14666));
  jand g14411(.dina(n14573), .dinb(n14565), .dout(n14667));
  jor  g14412(.dina(n14667), .dinb(n14666), .dout(n14668));
  jand g14413(.dina(n14554), .dinb(n14468), .dout(n14669));
  jand g14414(.dina(n14563), .dinb(n14555), .dout(n14670));
  jor  g14415(.dina(n14670), .dinb(n14669), .dout(n14671));
  jand g14416(.dina(n14544), .dinb(n14471), .dout(n14672));
  jand g14417(.dina(n14553), .dinb(n14545), .dout(n14673));
  jor  g14418(.dina(n14673), .dinb(n14672), .dout(n14674));
  jand g14419(.dina(n14534), .dinb(n14531), .dout(n14675));
  jand g14420(.dina(n14543), .dinb(n14535), .dout(n14676));
  jor  g14421(.dina(n14676), .dinb(n14675), .dout(n14677));
  jand g14422(.dina(n14521), .dinb(n14514), .dout(n14678));
  jand g14423(.dina(n14530), .dinb(n14522), .dout(n14679));
  jor  g14424(.dina(n14679), .dinb(n14678), .dout(n14680));
  jand g14425(.dina(n14504), .dinb(n14474), .dout(n14681));
  jand g14426(.dina(n14513), .dinb(n14505), .dout(n14682));
  jor  g14427(.dina(n14682), .dinb(n14681), .dout(n14683));
  jand g14428(.dina(n14494), .dinb(n14477), .dout(n14684));
  jand g14429(.dina(n14503), .dinb(n14495), .dout(n14685));
  jor  g14430(.dina(n14685), .dinb(n14684), .dout(n14686));
  jand g14431(.dina(n14484), .dinb(n14481), .dout(n14687));
  jand g14432(.dina(n14493), .dinb(n14485), .dout(n14688));
  jor  g14433(.dina(n14688), .dinb(n14687), .dout(n14689));
  jand g14434(.dina(n10594), .dinb(b16 ), .dout(n14690));
  jand g14435(.dina(n10129), .dinb(b17 ), .dout(n14691));
  jor  g14436(.dina(n14691), .dinb(n14690), .dout(n14692));
  jnot g14437(.din(n14692), .dout(n14693));
  jxor g14438(.dina(n14693), .dinb(n14480), .dout(n14694));
  jor  g14439(.dina(n10134), .dinb(n1525), .dout(n14695));
  jor  g14440(.dina(n9849), .dinb(n1307), .dout(n14696));
  jor  g14441(.dina(n10137), .dinb(n1416), .dout(n14697));
  jor  g14442(.dina(n10132), .dinb(n1527), .dout(n14698));
  jand g14443(.dina(n14698), .dinb(n14697), .dout(n14699));
  jand g14444(.dina(n14699), .dinb(n14696), .dout(n14700));
  jand g14445(.dina(n14700), .dinb(n14695), .dout(n14701));
  jxor g14446(.dina(n14701), .dinb(n9559), .dout(n14702));
  jxor g14447(.dina(n14702), .dinb(n14694), .dout(n14703));
  jxor g14448(.dina(n14703), .dinb(n14689), .dout(n14704));
  jor  g14449(.dina(n9271), .dinb(n1879), .dout(n14705));
  jor  g14450(.dina(n9003), .dinb(n1637), .dout(n14706));
  jor  g14451(.dina(n9273), .dinb(n1759), .dout(n14707));
  jor  g14452(.dina(n9268), .dinb(n1881), .dout(n14708));
  jand g14453(.dina(n14708), .dinb(n14707), .dout(n14709));
  jand g14454(.dina(n14709), .dinb(n14706), .dout(n14710));
  jand g14455(.dina(n14710), .dinb(n14705), .dout(n14711));
  jxor g14456(.dina(n14711), .dinb(n8729), .dout(n14712));
  jxor g14457(.dina(n14712), .dinb(n14704), .dout(n14713));
  jxor g14458(.dina(n14713), .dinb(n14686), .dout(n14714));
  jor  g14459(.dina(n8457), .dinb(n2277), .dout(n14715));
  jor  g14460(.dina(n8185), .dinb(n2007), .dout(n14716));
  jor  g14461(.dina(n8454), .dinb(n2279), .dout(n14717));
  jor  g14462(.dina(n8459), .dinb(n2142), .dout(n14718));
  jand g14463(.dina(n14718), .dinb(n14717), .dout(n14719));
  jand g14464(.dina(n14719), .dinb(n14716), .dout(n14720));
  jand g14465(.dina(n14720), .dinb(n14715), .dout(n14721));
  jxor g14466(.dina(n14721), .dinb(n7929), .dout(n14722));
  jxor g14467(.dina(n14722), .dinb(n14714), .dout(n14723));
  jxor g14468(.dina(n14723), .dinb(n14683), .dout(n14724));
  jor  g14469(.dina(n7660), .dinb(n2711), .dout(n14725));
  jor  g14470(.dina(n7415), .dinb(n2415), .dout(n14726));
  jor  g14471(.dina(n7662), .dinb(n2713), .dout(n14727));
  jor  g14472(.dina(n7657), .dinb(n2563), .dout(n14728));
  jand g14473(.dina(n14728), .dinb(n14727), .dout(n14729));
  jand g14474(.dina(n14729), .dinb(n14726), .dout(n14730));
  jand g14475(.dina(n14730), .dinb(n14725), .dout(n14731));
  jxor g14476(.dina(n14731), .dinb(n7166), .dout(n14732));
  jxor g14477(.dina(n14732), .dinb(n14724), .dout(n14733));
  jxor g14478(.dina(n14733), .dinb(n14680), .dout(n14734));
  jor  g14479(.dina(n6914), .dinb(n3184), .dout(n14735));
  jor  g14480(.dina(n6673), .dinb(n2862), .dout(n14736));
  jor  g14481(.dina(n6911), .dinb(n3023), .dout(n14737));
  jor  g14482(.dina(n6916), .dinb(n3186), .dout(n14738));
  jand g14483(.dina(n14738), .dinb(n14737), .dout(n14739));
  jand g14484(.dina(n14739), .dinb(n14736), .dout(n14740));
  jand g14485(.dina(n14740), .dinb(n14735), .dout(n14741));
  jxor g14486(.dina(n14741), .dinb(n6443), .dout(n14742));
  jxor g14487(.dina(n14742), .dinb(n14734), .dout(n14743));
  jxor g14488(.dina(n14743), .dinb(n14677), .dout(n14744));
  jor  g14489(.dina(n6207), .dinb(n3696), .dout(n14745));
  jor  g14490(.dina(n5975), .dinb(n3348), .dout(n14746));
  jor  g14491(.dina(n6205), .dinb(n3698), .dout(n14747));
  jor  g14492(.dina(n6210), .dinb(n3522), .dout(n14748));
  jand g14493(.dina(n14748), .dinb(n14747), .dout(n14749));
  jand g14494(.dina(n14749), .dinb(n14746), .dout(n14750));
  jand g14495(.dina(n14750), .dinb(n14745), .dout(n14751));
  jxor g14496(.dina(n14751), .dinb(n5759), .dout(n14752));
  jxor g14497(.dina(n14752), .dinb(n14744), .dout(n14753));
  jxor g14498(.dina(n14753), .dinb(n14674), .dout(n14754));
  jor  g14499(.dina(n5537), .dinb(n4247), .dout(n14755));
  jor  g14500(.dina(n5315), .dinb(n3873), .dout(n14756));
  jor  g14501(.dina(n5539), .dinb(n4249), .dout(n14757));
  jor  g14502(.dina(n5534), .dinb(n4060), .dout(n14758));
  jand g14503(.dina(n14758), .dinb(n14757), .dout(n14759));
  jand g14504(.dina(n14759), .dinb(n14756), .dout(n14760));
  jand g14505(.dina(n14760), .dinb(n14755), .dout(n14761));
  jxor g14506(.dina(n14761), .dinb(n5111), .dout(n14762));
  jxor g14507(.dina(n14762), .dinb(n14754), .dout(n14763));
  jxor g14508(.dina(n14763), .dinb(n14671), .dout(n14764));
  jor  g14509(.dina(n4837), .dinb(n4902), .dout(n14765));
  jor  g14510(.dina(n4696), .dinb(n4437), .dout(n14766));
  jor  g14511(.dina(n4899), .dinb(n4839), .dout(n14767));
  jor  g14512(.dina(n4904), .dinb(n4637), .dout(n14768));
  jand g14513(.dina(n14768), .dinb(n14767), .dout(n14769));
  jand g14514(.dina(n14769), .dinb(n14766), .dout(n14770));
  jand g14515(.dina(n14770), .dinb(n14765), .dout(n14771));
  jxor g14516(.dina(n14771), .dinb(n4505), .dout(n14772));
  jxor g14517(.dina(n14772), .dinb(n14764), .dout(n14773));
  jxor g14518(.dina(n14773), .dinb(n14668), .dout(n14774));
  jor  g14519(.dina(n5467), .dinb(n4305), .dout(n14775));
  jor  g14520(.dina(n4116), .dinb(n5040), .dout(n14776));
  jor  g14521(.dina(n4308), .dinb(n5253), .dout(n14777));
  jor  g14522(.dina(n4303), .dinb(n5469), .dout(n14778));
  jand g14523(.dina(n14778), .dinb(n14777), .dout(n14779));
  jand g14524(.dina(n14779), .dinb(n14776), .dout(n14780));
  jand g14525(.dina(n14780), .dinb(n14775), .dout(n14781));
  jxor g14526(.dina(n14781), .dinb(n3938), .dout(n14782));
  jxor g14527(.dina(n14782), .dinb(n14774), .dout(n14783));
  jxor g14528(.dina(n14783), .dinb(n14665), .dout(n14784));
  jor  g14529(.dina(n6137), .dinb(n3751), .dout(n14785));
  jor  g14530(.dina(n3574), .dinb(n5685), .dout(n14786));
  jor  g14531(.dina(n3754), .dinb(n5911), .dout(n14787));
  jor  g14532(.dina(n3749), .dinb(n6139), .dout(n14788));
  jand g14533(.dina(n14788), .dinb(n14787), .dout(n14789));
  jand g14534(.dina(n14789), .dinb(n14786), .dout(n14790));
  jand g14535(.dina(n14790), .dinb(n14785), .dout(n14791));
  jxor g14536(.dina(n14791), .dinb(n3410), .dout(n14792));
  jxor g14537(.dina(n14792), .dinb(n14784), .dout(n14793));
  jxor g14538(.dina(n14793), .dinb(n14662), .dout(n14794));
  jxor g14539(.dina(n14794), .dinb(n14650), .dout(n14795));
  jxor g14540(.dina(n14795), .dinb(n14638), .dout(n14796));
  jand g14541(.dina(n14431), .dinb(n14423), .dout(n14797));
  jand g14542(.dina(n14596), .dinb(n14432), .dout(n14798));
  jor  g14543(.dina(n14798), .dinb(n14797), .dout(n14799));
  jor  g14544(.dina(n9193), .dinb(n1921), .dout(n14800));
  jor  g14545(.dina(n1806), .dinb(n8644), .dout(n14801));
  jor  g14546(.dina(n1918), .dinb(n8920), .dout(n14802));
  jor  g14547(.dina(n1923), .dinb(n9195), .dout(n14803));
  jand g14548(.dina(n14803), .dinb(n14802), .dout(n14804));
  jand g14549(.dina(n14804), .dinb(n14801), .dout(n14805));
  jand g14550(.dina(n14805), .dinb(n14800), .dout(n14806));
  jxor g14551(.dina(n14806), .dinb(n1687), .dout(n14807));
  jxor g14552(.dina(n14807), .dinb(n14799), .dout(n14808));
  jxor g14553(.dina(n14808), .dinb(n14796), .dout(n14809));
  jxor g14554(.dina(n14809), .dinb(n14626), .dout(n14810));
  jand g14555(.dina(n14407), .dinb(n14399), .dout(n14811));
  jand g14556(.dina(n14598), .dinb(n14408), .dout(n14812));
  jor  g14557(.dina(n14812), .dinb(n14811), .dout(n14813));
  jnot g14558(.din(n14813), .dout(n14814));
  jand g14559(.dina(n1148), .dinb(b63 ), .dout(n14815));
  jand g14560(.dina(n10832), .dinb(n1053), .dout(n14816));
  jor  g14561(.dina(n14816), .dinb(n14815), .dout(n14817));
  jxor g14562(.dina(n14817), .dinb(n1061), .dout(n14818));
  jxor g14563(.dina(n14818), .dinb(n14814), .dout(n14819));
  jxor g14564(.dina(n14819), .dinb(n14810), .dout(n14820));
  jxor g14565(.dina(n14820), .dinb(n14614), .dout(n14821));
  jnot g14566(.din(n14821), .dout(n14822));
  jxor g14567(.dina(n14822), .dinb(n14611), .dout(f80 ));
  jand g14568(.dina(n14820), .dinb(n14614), .dout(n14824));
  jnot g14569(.din(n14824), .dout(n14825));
  jor  g14570(.dina(n14822), .dinb(n14611), .dout(n14826));
  jand g14571(.dina(n14826), .dinb(n14825), .dout(n14827));
  jor  g14572(.dina(n14818), .dinb(n14814), .dout(n14828));
  jand g14573(.dina(n14819), .dinb(n14810), .dout(n14829));
  jnot g14574(.din(n14829), .dout(n14830));
  jand g14575(.dina(n14830), .dinb(n14828), .dout(n14831));
  jnot g14576(.din(n14831), .dout(n14832));
  jand g14577(.dina(n14625), .dinb(n14617), .dout(n14833));
  jand g14578(.dina(n14809), .dinb(n14626), .dout(n14834));
  jor  g14579(.dina(n14834), .dinb(n14833), .dout(n14835));
  jor  g14580(.dina(n10521), .dinb(n1569), .dout(n14836));
  jor  g14581(.dina(n1453), .dinb(n9759), .dout(n14837));
  jor  g14582(.dina(n1566), .dinb(n10051), .dout(n14838));
  jor  g14583(.dina(n1571), .dinb(n10523), .dout(n14839));
  jand g14584(.dina(n14839), .dinb(n14838), .dout(n14840));
  jand g14585(.dina(n14840), .dinb(n14837), .dout(n14841));
  jand g14586(.dina(n14841), .dinb(n14836), .dout(n14842));
  jxor g14587(.dina(n14842), .dinb(n1351), .dout(n14843));
  jxor g14588(.dina(n14843), .dinb(n14835), .dout(n14844));
  jand g14589(.dina(n14807), .dinb(n14799), .dout(n14845));
  jand g14590(.dina(n14808), .dinb(n14796), .dout(n14846));
  jor  g14591(.dina(n14846), .dinb(n14845), .dout(n14847));
  jor  g14592(.dina(n9473), .dinb(n1921), .dout(n14848));
  jor  g14593(.dina(n1806), .dinb(n8920), .dout(n14849));
  jor  g14594(.dina(n1923), .dinb(n9475), .dout(n14850));
  jor  g14595(.dina(n1918), .dinb(n9195), .dout(n14851));
  jand g14596(.dina(n14851), .dinb(n14850), .dout(n14852));
  jand g14597(.dina(n14852), .dinb(n14849), .dout(n14853));
  jand g14598(.dina(n14853), .dinb(n14848), .dout(n14854));
  jxor g14599(.dina(n14854), .dinb(n1687), .dout(n14855));
  jxor g14600(.dina(n14855), .dinb(n14847), .dout(n14856));
  jand g14601(.dina(n14637), .dinb(n14629), .dout(n14857));
  jand g14602(.dina(n14795), .dinb(n14638), .dout(n14858));
  jor  g14603(.dina(n14858), .dinb(n14857), .dout(n14859));
  jor  g14604(.dina(n8642), .dinb(n2324), .dout(n14860));
  jor  g14605(.dina(n2186), .dinb(n8111), .dout(n14861));
  jor  g14606(.dina(n2321), .dinb(n8378), .dout(n14862));
  jor  g14607(.dina(n2326), .dinb(n8644), .dout(n14863));
  jand g14608(.dina(n14863), .dinb(n14862), .dout(n14864));
  jand g14609(.dina(n14864), .dinb(n14861), .dout(n14865));
  jand g14610(.dina(n14865), .dinb(n14860), .dout(n14866));
  jxor g14611(.dina(n14866), .dinb(n2057), .dout(n14867));
  jxor g14612(.dina(n14867), .dinb(n14859), .dout(n14868));
  jand g14613(.dina(n14649), .dinb(n14641), .dout(n14869));
  jand g14614(.dina(n14794), .dinb(n14650), .dout(n14870));
  jor  g14615(.dina(n14870), .dinb(n14869), .dout(n14871));
  jor  g14616(.dina(n7844), .dinb(n2764), .dout(n14872));
  jor  g14617(.dina(n2609), .dinb(n7338), .dout(n14873));
  jor  g14618(.dina(n2761), .dinb(n7846), .dout(n14874));
  jor  g14619(.dina(n2766), .dinb(n7590), .dout(n14875));
  jand g14620(.dina(n14875), .dinb(n14874), .dout(n14876));
  jand g14621(.dina(n14876), .dinb(n14873), .dout(n14877));
  jand g14622(.dina(n14877), .dinb(n14872), .dout(n14878));
  jxor g14623(.dina(n14878), .dinb(n2468), .dout(n14879));
  jxor g14624(.dina(n14879), .dinb(n14871), .dout(n14880));
  jand g14625(.dina(n14783), .dinb(n14665), .dout(n14881));
  jand g14626(.dina(n14792), .dinb(n14784), .dout(n14882));
  jor  g14627(.dina(n14882), .dinb(n14881), .dout(n14883));
  jand g14628(.dina(n14773), .dinb(n14668), .dout(n14884));
  jand g14629(.dina(n14782), .dinb(n14774), .dout(n14885));
  jor  g14630(.dina(n14885), .dinb(n14884), .dout(n14886));
  jand g14631(.dina(n14763), .dinb(n14671), .dout(n14887));
  jand g14632(.dina(n14772), .dinb(n14764), .dout(n14888));
  jor  g14633(.dina(n14888), .dinb(n14887), .dout(n14889));
  jand g14634(.dina(n14753), .dinb(n14674), .dout(n14890));
  jand g14635(.dina(n14762), .dinb(n14754), .dout(n14891));
  jor  g14636(.dina(n14891), .dinb(n14890), .dout(n14892));
  jand g14637(.dina(n14743), .dinb(n14677), .dout(n14893));
  jand g14638(.dina(n14752), .dinb(n14744), .dout(n14894));
  jor  g14639(.dina(n14894), .dinb(n14893), .dout(n14895));
  jand g14640(.dina(n14723), .dinb(n14683), .dout(n14896));
  jand g14641(.dina(n14732), .dinb(n14724), .dout(n14897));
  jor  g14642(.dina(n14897), .dinb(n14896), .dout(n14898));
  jand g14643(.dina(n14713), .dinb(n14686), .dout(n14899));
  jand g14644(.dina(n14722), .dinb(n14714), .dout(n14900));
  jor  g14645(.dina(n14900), .dinb(n14899), .dout(n14901));
  jand g14646(.dina(n14703), .dinb(n14689), .dout(n14902));
  jand g14647(.dina(n14712), .dinb(n14704), .dout(n14903));
  jor  g14648(.dina(n14903), .dinb(n14902), .dout(n14904));
  jand g14649(.dina(n14693), .dinb(n14480), .dout(n14905));
  jand g14650(.dina(n14702), .dinb(n14694), .dout(n14906));
  jor  g14651(.dina(n14906), .dinb(n14905), .dout(n14907));
  jand g14652(.dina(n10594), .dinb(b17 ), .dout(n14908));
  jand g14653(.dina(n10129), .dinb(b18 ), .dout(n14909));
  jor  g14654(.dina(n14909), .dinb(n14908), .dout(n14910));
  jxor g14655(.dina(n14910), .dinb(n1061), .dout(n14911));
  jxor g14656(.dina(n14911), .dinb(n14692), .dout(n14912));
  jor  g14657(.dina(n10134), .dinb(n1635), .dout(n14913));
  jor  g14658(.dina(n9849), .dinb(n1416), .dout(n14914));
  jor  g14659(.dina(n10132), .dinb(n1637), .dout(n14915));
  jor  g14660(.dina(n10137), .dinb(n1527), .dout(n14916));
  jand g14661(.dina(n14916), .dinb(n14915), .dout(n14917));
  jand g14662(.dina(n14917), .dinb(n14914), .dout(n14918));
  jand g14663(.dina(n14918), .dinb(n14913), .dout(n14919));
  jxor g14664(.dina(n14919), .dinb(n9559), .dout(n14920));
  jxor g14665(.dina(n14920), .dinb(n14912), .dout(n14921));
  jxor g14666(.dina(n14921), .dinb(n14907), .dout(n14922));
  jor  g14667(.dina(n9271), .dinb(n2005), .dout(n14923));
  jor  g14668(.dina(n9003), .dinb(n1759), .dout(n14924));
  jor  g14669(.dina(n9268), .dinb(n2007), .dout(n14925));
  jor  g14670(.dina(n9273), .dinb(n1881), .dout(n14926));
  jand g14671(.dina(n14926), .dinb(n14925), .dout(n14927));
  jand g14672(.dina(n14927), .dinb(n14924), .dout(n14928));
  jand g14673(.dina(n14928), .dinb(n14923), .dout(n14929));
  jxor g14674(.dina(n14929), .dinb(n8729), .dout(n14930));
  jxor g14675(.dina(n14930), .dinb(n14922), .dout(n14931));
  jxor g14676(.dina(n14931), .dinb(n14904), .dout(n14932));
  jor  g14677(.dina(n8457), .dinb(n2413), .dout(n14933));
  jor  g14678(.dina(n8185), .dinb(n2142), .dout(n14934));
  jor  g14679(.dina(n8459), .dinb(n2279), .dout(n14935));
  jor  g14680(.dina(n8454), .dinb(n2415), .dout(n14936));
  jand g14681(.dina(n14936), .dinb(n14935), .dout(n14937));
  jand g14682(.dina(n14937), .dinb(n14934), .dout(n14938));
  jand g14683(.dina(n14938), .dinb(n14933), .dout(n14939));
  jxor g14684(.dina(n14939), .dinb(n7929), .dout(n14940));
  jxor g14685(.dina(n14940), .dinb(n14932), .dout(n14941));
  jxor g14686(.dina(n14941), .dinb(n14901), .dout(n14942));
  jor  g14687(.dina(n7660), .dinb(n2860), .dout(n14943));
  jor  g14688(.dina(n7415), .dinb(n2563), .dout(n14944));
  jor  g14689(.dina(n7657), .dinb(n2713), .dout(n14945));
  jor  g14690(.dina(n7662), .dinb(n2862), .dout(n14946));
  jand g14691(.dina(n14946), .dinb(n14945), .dout(n14947));
  jand g14692(.dina(n14947), .dinb(n14944), .dout(n14948));
  jand g14693(.dina(n14948), .dinb(n14943), .dout(n14949));
  jxor g14694(.dina(n14949), .dinb(n7166), .dout(n14950));
  jxor g14695(.dina(n14950), .dinb(n14942), .dout(n14951));
  jxor g14696(.dina(n14951), .dinb(n14898), .dout(n14952));
  jand g14697(.dina(n14733), .dinb(n14680), .dout(n14953));
  jand g14698(.dina(n14742), .dinb(n14734), .dout(n14954));
  jor  g14699(.dina(n14954), .dinb(n14953), .dout(n14955));
  jor  g14700(.dina(n6914), .dinb(n3346), .dout(n14956));
  jor  g14701(.dina(n6673), .dinb(n3023), .dout(n14957));
  jor  g14702(.dina(n6916), .dinb(n3348), .dout(n14958));
  jor  g14703(.dina(n6911), .dinb(n3186), .dout(n14959));
  jand g14704(.dina(n14959), .dinb(n14958), .dout(n14960));
  jand g14705(.dina(n14960), .dinb(n14957), .dout(n14961));
  jand g14706(.dina(n14961), .dinb(n14956), .dout(n14962));
  jxor g14707(.dina(n14962), .dinb(n6443), .dout(n14963));
  jxor g14708(.dina(n14963), .dinb(n14955), .dout(n14964));
  jxor g14709(.dina(n14964), .dinb(n14952), .dout(n14965));
  jor  g14710(.dina(n6207), .dinb(n3871), .dout(n14966));
  jor  g14711(.dina(n5975), .dinb(n3522), .dout(n14967));
  jor  g14712(.dina(n6205), .dinb(n3873), .dout(n14968));
  jor  g14713(.dina(n6210), .dinb(n3698), .dout(n14969));
  jand g14714(.dina(n14969), .dinb(n14968), .dout(n14970));
  jand g14715(.dina(n14970), .dinb(n14967), .dout(n14971));
  jand g14716(.dina(n14971), .dinb(n14966), .dout(n14972));
  jxor g14717(.dina(n14972), .dinb(n5759), .dout(n14973));
  jxor g14718(.dina(n14973), .dinb(n14965), .dout(n14974));
  jxor g14719(.dina(n14974), .dinb(n14895), .dout(n14975));
  jor  g14720(.dina(n5537), .dinb(n4435), .dout(n14976));
  jor  g14721(.dina(n5315), .dinb(n4060), .dout(n14977));
  jor  g14722(.dina(n5534), .dinb(n4249), .dout(n14978));
  jor  g14723(.dina(n5539), .dinb(n4437), .dout(n14979));
  jand g14724(.dina(n14979), .dinb(n14978), .dout(n14980));
  jand g14725(.dina(n14980), .dinb(n14977), .dout(n14981));
  jand g14726(.dina(n14981), .dinb(n14976), .dout(n14982));
  jxor g14727(.dina(n14982), .dinb(n5111), .dout(n14983));
  jxor g14728(.dina(n14983), .dinb(n14975), .dout(n14984));
  jxor g14729(.dina(n14984), .dinb(n14892), .dout(n14985));
  jor  g14730(.dina(n5038), .dinb(n4902), .dout(n14986));
  jor  g14731(.dina(n4696), .dinb(n4637), .dout(n14987));
  jor  g14732(.dina(n4899), .dinb(n5040), .dout(n14988));
  jor  g14733(.dina(n4904), .dinb(n4839), .dout(n14989));
  jand g14734(.dina(n14989), .dinb(n14988), .dout(n14990));
  jand g14735(.dina(n14990), .dinb(n14987), .dout(n14991));
  jand g14736(.dina(n14991), .dinb(n14986), .dout(n14992));
  jxor g14737(.dina(n14992), .dinb(n4505), .dout(n14993));
  jxor g14738(.dina(n14993), .dinb(n14985), .dout(n14994));
  jxor g14739(.dina(n14994), .dinb(n14889), .dout(n14995));
  jor  g14740(.dina(n5683), .dinb(n4305), .dout(n14996));
  jor  g14741(.dina(n4116), .dinb(n5253), .dout(n14997));
  jor  g14742(.dina(n4303), .dinb(n5685), .dout(n14998));
  jor  g14743(.dina(n4308), .dinb(n5469), .dout(n14999));
  jand g14744(.dina(n14999), .dinb(n14998), .dout(n15000));
  jand g14745(.dina(n15000), .dinb(n14997), .dout(n15001));
  jand g14746(.dina(n15001), .dinb(n14996), .dout(n15002));
  jxor g14747(.dina(n15002), .dinb(n3938), .dout(n15003));
  jxor g14748(.dina(n15003), .dinb(n14995), .dout(n15004));
  jxor g14749(.dina(n15004), .dinb(n14886), .dout(n15005));
  jor  g14750(.dina(n6364), .dinb(n3751), .dout(n15006));
  jor  g14751(.dina(n3574), .dinb(n5911), .dout(n15007));
  jor  g14752(.dina(n3749), .dinb(n6366), .dout(n15008));
  jor  g14753(.dina(n3754), .dinb(n6139), .dout(n15009));
  jand g14754(.dina(n15009), .dinb(n15008), .dout(n15010));
  jand g14755(.dina(n15010), .dinb(n15007), .dout(n15011));
  jand g14756(.dina(n15011), .dinb(n15006), .dout(n15012));
  jxor g14757(.dina(n15012), .dinb(n3410), .dout(n15013));
  jxor g14758(.dina(n15013), .dinb(n15005), .dout(n15014));
  jxor g14759(.dina(n15014), .dinb(n14883), .dout(n15015));
  jand g14760(.dina(n14661), .dinb(n14653), .dout(n15016));
  jand g14761(.dina(n14793), .dinb(n14662), .dout(n15017));
  jor  g14762(.dina(n15017), .dinb(n15016), .dout(n15018));
  jor  g14763(.dina(n7084), .dinb(n3239), .dout(n15019));
  jor  g14764(.dina(n3072), .dinb(n6605), .dout(n15020));
  jor  g14765(.dina(n3237), .dinb(n7086), .dout(n15021));
  jor  g14766(.dina(n3242), .dinb(n6846), .dout(n15022));
  jand g14767(.dina(n15022), .dinb(n15021), .dout(n15023));
  jand g14768(.dina(n15023), .dinb(n15020), .dout(n15024));
  jand g14769(.dina(n15024), .dinb(n15019), .dout(n15025));
  jxor g14770(.dina(n15025), .dinb(n2918), .dout(n15026));
  jxor g14771(.dina(n15026), .dinb(n15018), .dout(n15027));
  jxor g14772(.dina(n15027), .dinb(n15015), .dout(n15028));
  jxor g14773(.dina(n15028), .dinb(n14880), .dout(n15029));
  jxor g14774(.dina(n15029), .dinb(n14868), .dout(n15030));
  jxor g14775(.dina(n15030), .dinb(n14856), .dout(n15031));
  jxor g14776(.dina(n15031), .dinb(n14844), .dout(n15032));
  jxor g14777(.dina(n15032), .dinb(n14832), .dout(n15033));
  jnot g14778(.din(n15033), .dout(n15034));
  jxor g14779(.dina(n15034), .dinb(n14827), .dout(f81 ));
  jand g14780(.dina(n15032), .dinb(n14832), .dout(n15036));
  jnot g14781(.din(n15036), .dout(n15037));
  jor  g14782(.dina(n15034), .dinb(n14827), .dout(n15038));
  jand g14783(.dina(n15038), .dinb(n15037), .dout(n15039));
  jand g14784(.dina(n14843), .dinb(n14835), .dout(n15040));
  jand g14785(.dina(n15031), .dinb(n14844), .dout(n15041));
  jor  g14786(.dina(n15041), .dinb(n15040), .dout(n15042));
  jand g14787(.dina(n14867), .dinb(n14859), .dout(n15043));
  jand g14788(.dina(n15029), .dinb(n14868), .dout(n15044));
  jor  g14789(.dina(n15044), .dinb(n15043), .dout(n15045));
  jor  g14790(.dina(n9757), .dinb(n1921), .dout(n15046));
  jor  g14791(.dina(n1806), .dinb(n9195), .dout(n15047));
  jor  g14792(.dina(n1918), .dinb(n9475), .dout(n15048));
  jor  g14793(.dina(n1923), .dinb(n9759), .dout(n15049));
  jand g14794(.dina(n15049), .dinb(n15048), .dout(n15050));
  jand g14795(.dina(n15050), .dinb(n15047), .dout(n15051));
  jand g14796(.dina(n15051), .dinb(n15046), .dout(n15052));
  jxor g14797(.dina(n15052), .dinb(n1687), .dout(n15053));
  jxor g14798(.dina(n15053), .dinb(n15045), .dout(n15054));
  jand g14799(.dina(n14879), .dinb(n14871), .dout(n15055));
  jand g14800(.dina(n15028), .dinb(n14880), .dout(n15056));
  jor  g14801(.dina(n15056), .dinb(n15055), .dout(n15057));
  jor  g14802(.dina(n8918), .dinb(n2324), .dout(n15058));
  jor  g14803(.dina(n2186), .dinb(n8378), .dout(n15059));
  jor  g14804(.dina(n2326), .dinb(n8920), .dout(n15060));
  jor  g14805(.dina(n2321), .dinb(n8644), .dout(n15061));
  jand g14806(.dina(n15061), .dinb(n15060), .dout(n15062));
  jand g14807(.dina(n15062), .dinb(n15059), .dout(n15063));
  jand g14808(.dina(n15063), .dinb(n15058), .dout(n15064));
  jxor g14809(.dina(n15064), .dinb(n2057), .dout(n15065));
  jxor g14810(.dina(n15065), .dinb(n15057), .dout(n15066));
  jand g14811(.dina(n15026), .dinb(n15018), .dout(n15067));
  jand g14812(.dina(n15027), .dinb(n15015), .dout(n15068));
  jor  g14813(.dina(n15068), .dinb(n15067), .dout(n15069));
  jor  g14814(.dina(n8109), .dinb(n2764), .dout(n15070));
  jor  g14815(.dina(n2609), .dinb(n7590), .dout(n15071));
  jor  g14816(.dina(n2761), .dinb(n8111), .dout(n15072));
  jor  g14817(.dina(n2766), .dinb(n7846), .dout(n15073));
  jand g14818(.dina(n15073), .dinb(n15072), .dout(n15074));
  jand g14819(.dina(n15074), .dinb(n15071), .dout(n15075));
  jand g14820(.dina(n15075), .dinb(n15070), .dout(n15076));
  jxor g14821(.dina(n15076), .dinb(n2468), .dout(n15077));
  jxor g14822(.dina(n15077), .dinb(n15069), .dout(n15078));
  jand g14823(.dina(n15013), .dinb(n15005), .dout(n15079));
  jand g14824(.dina(n15014), .dinb(n14883), .dout(n15080));
  jor  g14825(.dina(n15080), .dinb(n15079), .dout(n15081));
  jor  g14826(.dina(n7336), .dinb(n3239), .dout(n15082));
  jor  g14827(.dina(n3072), .dinb(n6846), .dout(n15083));
  jor  g14828(.dina(n3242), .dinb(n7086), .dout(n15084));
  jor  g14829(.dina(n3237), .dinb(n7338), .dout(n15085));
  jand g14830(.dina(n15085), .dinb(n15084), .dout(n15086));
  jand g14831(.dina(n15086), .dinb(n15083), .dout(n15087));
  jand g14832(.dina(n15087), .dinb(n15082), .dout(n15088));
  jxor g14833(.dina(n15088), .dinb(n2918), .dout(n15089));
  jxor g14834(.dina(n15089), .dinb(n15081), .dout(n15090));
  jand g14835(.dina(n15003), .dinb(n14995), .dout(n15091));
  jand g14836(.dina(n15004), .dinb(n14886), .dout(n15092));
  jor  g14837(.dina(n15092), .dinb(n15091), .dout(n15093));
  jand g14838(.dina(n14993), .dinb(n14985), .dout(n15094));
  jand g14839(.dina(n14994), .dinb(n14889), .dout(n15095));
  jor  g14840(.dina(n15095), .dinb(n15094), .dout(n15096));
  jand g14841(.dina(n14983), .dinb(n14975), .dout(n15097));
  jand g14842(.dina(n14984), .dinb(n14892), .dout(n15098));
  jor  g14843(.dina(n15098), .dinb(n15097), .dout(n15099));
  jand g14844(.dina(n14973), .dinb(n14965), .dout(n15100));
  jand g14845(.dina(n14974), .dinb(n14895), .dout(n15101));
  jor  g14846(.dina(n15101), .dinb(n15100), .dout(n15102));
  jand g14847(.dina(n14963), .dinb(n14955), .dout(n15103));
  jand g14848(.dina(n14964), .dinb(n14952), .dout(n15104));
  jor  g14849(.dina(n15104), .dinb(n15103), .dout(n15105));
  jand g14850(.dina(n14950), .dinb(n14942), .dout(n15106));
  jand g14851(.dina(n14951), .dinb(n14898), .dout(n15107));
  jor  g14852(.dina(n15107), .dinb(n15106), .dout(n15108));
  jand g14853(.dina(n14930), .dinb(n14922), .dout(n15109));
  jand g14854(.dina(n14931), .dinb(n14904), .dout(n15110));
  jor  g14855(.dina(n15110), .dinb(n15109), .dout(n15111));
  jand g14856(.dina(n10594), .dinb(b18 ), .dout(n15112));
  jand g14857(.dina(n10129), .dinb(b19 ), .dout(n15113));
  jor  g14858(.dina(n15113), .dinb(n15112), .dout(n15114));
  jnot g14859(.din(n15114), .dout(n15115));
  jand g14860(.dina(n14910), .dinb(n1061), .dout(n15116));
  jand g14861(.dina(n14911), .dinb(n14692), .dout(n15117));
  jor  g14862(.dina(n15117), .dinb(n15116), .dout(n15118));
  jxor g14863(.dina(n15118), .dinb(n15115), .dout(n15119));
  jor  g14864(.dina(n10134), .dinb(n1757), .dout(n15120));
  jor  g14865(.dina(n9849), .dinb(n1527), .dout(n15121));
  jor  g14866(.dina(n10132), .dinb(n1759), .dout(n15122));
  jor  g14867(.dina(n10137), .dinb(n1637), .dout(n15123));
  jand g14868(.dina(n15123), .dinb(n15122), .dout(n15124));
  jand g14869(.dina(n15124), .dinb(n15121), .dout(n15125));
  jand g14870(.dina(n15125), .dinb(n15120), .dout(n15126));
  jxor g14871(.dina(n15126), .dinb(n9559), .dout(n15127));
  jxor g14872(.dina(n15127), .dinb(n15119), .dout(n15128));
  jand g14873(.dina(n14920), .dinb(n14912), .dout(n15129));
  jand g14874(.dina(n14921), .dinb(n14907), .dout(n15130));
  jor  g14875(.dina(n15130), .dinb(n15129), .dout(n15131));
  jxor g14876(.dina(n15131), .dinb(n15128), .dout(n15132));
  jor  g14877(.dina(n9271), .dinb(n2140), .dout(n15133));
  jor  g14878(.dina(n9003), .dinb(n1881), .dout(n15134));
  jor  g14879(.dina(n9273), .dinb(n2007), .dout(n15135));
  jor  g14880(.dina(n9268), .dinb(n2142), .dout(n15136));
  jand g14881(.dina(n15136), .dinb(n15135), .dout(n15137));
  jand g14882(.dina(n15137), .dinb(n15134), .dout(n15138));
  jand g14883(.dina(n15138), .dinb(n15133), .dout(n15139));
  jxor g14884(.dina(n15139), .dinb(n8729), .dout(n15140));
  jxor g14885(.dina(n15140), .dinb(n15132), .dout(n15141));
  jxor g14886(.dina(n15141), .dinb(n15111), .dout(n15142));
  jor  g14887(.dina(n8457), .dinb(n2561), .dout(n15143));
  jor  g14888(.dina(n8185), .dinb(n2279), .dout(n15144));
  jor  g14889(.dina(n8459), .dinb(n2415), .dout(n15145));
  jor  g14890(.dina(n8454), .dinb(n2563), .dout(n15146));
  jand g14891(.dina(n15146), .dinb(n15145), .dout(n15147));
  jand g14892(.dina(n15147), .dinb(n15144), .dout(n15148));
  jand g14893(.dina(n15148), .dinb(n15143), .dout(n15149));
  jxor g14894(.dina(n15149), .dinb(n7929), .dout(n15150));
  jxor g14895(.dina(n15150), .dinb(n15142), .dout(n15151));
  jand g14896(.dina(n14940), .dinb(n14932), .dout(n15152));
  jand g14897(.dina(n14941), .dinb(n14901), .dout(n15153));
  jor  g14898(.dina(n15153), .dinb(n15152), .dout(n15154));
  jxor g14899(.dina(n15154), .dinb(n15151), .dout(n15155));
  jor  g14900(.dina(n7660), .dinb(n3021), .dout(n15156));
  jor  g14901(.dina(n7415), .dinb(n2713), .dout(n15157));
  jor  g14902(.dina(n7657), .dinb(n2862), .dout(n15158));
  jor  g14903(.dina(n7662), .dinb(n3023), .dout(n15159));
  jand g14904(.dina(n15159), .dinb(n15158), .dout(n15160));
  jand g14905(.dina(n15160), .dinb(n15157), .dout(n15161));
  jand g14906(.dina(n15161), .dinb(n15156), .dout(n15162));
  jxor g14907(.dina(n15162), .dinb(n7166), .dout(n15163));
  jxor g14908(.dina(n15163), .dinb(n15155), .dout(n15164));
  jxor g14909(.dina(n15164), .dinb(n15108), .dout(n15165));
  jor  g14910(.dina(n6914), .dinb(n3520), .dout(n15166));
  jor  g14911(.dina(n6673), .dinb(n3186), .dout(n15167));
  jor  g14912(.dina(n6911), .dinb(n3348), .dout(n15168));
  jor  g14913(.dina(n6916), .dinb(n3522), .dout(n15169));
  jand g14914(.dina(n15169), .dinb(n15168), .dout(n15170));
  jand g14915(.dina(n15170), .dinb(n15167), .dout(n15171));
  jand g14916(.dina(n15171), .dinb(n15166), .dout(n15172));
  jxor g14917(.dina(n15172), .dinb(n6443), .dout(n15173));
  jxor g14918(.dina(n15173), .dinb(n15165), .dout(n15174));
  jxor g14919(.dina(n15174), .dinb(n15105), .dout(n15175));
  jor  g14920(.dina(n6207), .dinb(n4058), .dout(n15176));
  jor  g14921(.dina(n5975), .dinb(n3698), .dout(n15177));
  jor  g14922(.dina(n6210), .dinb(n3873), .dout(n15178));
  jor  g14923(.dina(n6205), .dinb(n4060), .dout(n15179));
  jand g14924(.dina(n15179), .dinb(n15178), .dout(n15180));
  jand g14925(.dina(n15180), .dinb(n15177), .dout(n15181));
  jand g14926(.dina(n15181), .dinb(n15176), .dout(n15182));
  jxor g14927(.dina(n15182), .dinb(n5759), .dout(n15183));
  jxor g14928(.dina(n15183), .dinb(n15175), .dout(n15184));
  jxor g14929(.dina(n15184), .dinb(n15102), .dout(n15185));
  jor  g14930(.dina(n5537), .dinb(n4635), .dout(n15186));
  jor  g14931(.dina(n5315), .dinb(n4249), .dout(n15187));
  jor  g14932(.dina(n5539), .dinb(n4637), .dout(n15188));
  jor  g14933(.dina(n5534), .dinb(n4437), .dout(n15189));
  jand g14934(.dina(n15189), .dinb(n15188), .dout(n15190));
  jand g14935(.dina(n15190), .dinb(n15187), .dout(n15191));
  jand g14936(.dina(n15191), .dinb(n15186), .dout(n15192));
  jxor g14937(.dina(n15192), .dinb(n5111), .dout(n15193));
  jxor g14938(.dina(n15193), .dinb(n15185), .dout(n15194));
  jxor g14939(.dina(n15194), .dinb(n15099), .dout(n15195));
  jor  g14940(.dina(n5251), .dinb(n4902), .dout(n15196));
  jor  g14941(.dina(n4696), .dinb(n4839), .dout(n15197));
  jor  g14942(.dina(n4899), .dinb(n5253), .dout(n15198));
  jor  g14943(.dina(n4904), .dinb(n5040), .dout(n15199));
  jand g14944(.dina(n15199), .dinb(n15198), .dout(n15200));
  jand g14945(.dina(n15200), .dinb(n15197), .dout(n15201));
  jand g14946(.dina(n15201), .dinb(n15196), .dout(n15202));
  jxor g14947(.dina(n15202), .dinb(n4505), .dout(n15203));
  jxor g14948(.dina(n15203), .dinb(n15195), .dout(n15204));
  jxor g14949(.dina(n15204), .dinb(n15096), .dout(n15205));
  jor  g14950(.dina(n5909), .dinb(n4305), .dout(n15206));
  jor  g14951(.dina(n4116), .dinb(n5469), .dout(n15207));
  jor  g14952(.dina(n4303), .dinb(n5911), .dout(n15208));
  jor  g14953(.dina(n4308), .dinb(n5685), .dout(n15209));
  jand g14954(.dina(n15209), .dinb(n15208), .dout(n15210));
  jand g14955(.dina(n15210), .dinb(n15207), .dout(n15211));
  jand g14956(.dina(n15211), .dinb(n15206), .dout(n15212));
  jxor g14957(.dina(n15212), .dinb(n3938), .dout(n15213));
  jxor g14958(.dina(n15213), .dinb(n15205), .dout(n15214));
  jxor g14959(.dina(n15214), .dinb(n15093), .dout(n15215));
  jor  g14960(.dina(n6603), .dinb(n3751), .dout(n15216));
  jor  g14961(.dina(n3574), .dinb(n6139), .dout(n15217));
  jor  g14962(.dina(n3754), .dinb(n6366), .dout(n15218));
  jor  g14963(.dina(n3749), .dinb(n6605), .dout(n15219));
  jand g14964(.dina(n15219), .dinb(n15218), .dout(n15220));
  jand g14965(.dina(n15220), .dinb(n15217), .dout(n15221));
  jand g14966(.dina(n15221), .dinb(n15216), .dout(n15222));
  jxor g14967(.dina(n15222), .dinb(n3410), .dout(n15223));
  jxor g14968(.dina(n15223), .dinb(n15215), .dout(n15224));
  jxor g14969(.dina(n15224), .dinb(n15090), .dout(n15225));
  jxor g14970(.dina(n15225), .dinb(n15078), .dout(n15226));
  jxor g14971(.dina(n15226), .dinb(n15066), .dout(n15227));
  jxor g14972(.dina(n15227), .dinb(n15054), .dout(n15228));
  jand g14973(.dina(n14855), .dinb(n14847), .dout(n15229));
  jand g14974(.dina(n15030), .dinb(n14856), .dout(n15230));
  jor  g14975(.dina(n15230), .dinb(n15229), .dout(n15231));
  jnot g14976(.din(n15231), .dout(n15232));
  jor  g14977(.dina(n10813), .dinb(n1569), .dout(n15233));
  jor  g14978(.dina(n1453), .dinb(n10051), .dout(n15234));
  jor  g14979(.dina(n1566), .dinb(n10523), .dout(n15235));
  jand g14980(.dina(n15235), .dinb(n15234), .dout(n15236));
  jand g14981(.dina(n15236), .dinb(n15233), .dout(n15237));
  jxor g14982(.dina(n15237), .dinb(a20 ), .dout(n15238));
  jxor g14983(.dina(n15238), .dinb(n15232), .dout(n15239));
  jxor g14984(.dina(n15239), .dinb(n15228), .dout(n15240));
  jxor g14985(.dina(n15240), .dinb(n15042), .dout(n15241));
  jnot g14986(.din(n15241), .dout(n15242));
  jxor g14987(.dina(n15242), .dinb(n15039), .dout(f82 ));
  jand g14988(.dina(n15240), .dinb(n15042), .dout(n15244));
  jnot g14989(.din(n15244), .dout(n15245));
  jor  g14990(.dina(n15242), .dinb(n15039), .dout(n15246));
  jand g14991(.dina(n15246), .dinb(n15245), .dout(n15247));
  jor  g14992(.dina(n15238), .dinb(n15232), .dout(n15248));
  jand g14993(.dina(n15239), .dinb(n15228), .dout(n15249));
  jnot g14994(.din(n15249), .dout(n15250));
  jand g14995(.dina(n15250), .dinb(n15248), .dout(n15251));
  jnot g14996(.din(n15251), .dout(n15252));
  jand g14997(.dina(n15053), .dinb(n15045), .dout(n15253));
  jand g14998(.dina(n15227), .dinb(n15054), .dout(n15254));
  jor  g14999(.dina(n15254), .dinb(n15253), .dout(n15255));
  jnot g15000(.din(n15255), .dout(n15256));
  jand g15001(.dina(n1454), .dinb(b63 ), .dout(n15257));
  jand g15002(.dina(n10832), .dinb(n1340), .dout(n15258));
  jor  g15003(.dina(n15258), .dinb(n15257), .dout(n15259));
  jxor g15004(.dina(n15259), .dinb(n1351), .dout(n15260));
  jxor g15005(.dina(n15260), .dinb(n15256), .dout(n15261));
  jand g15006(.dina(n15065), .dinb(n15057), .dout(n15262));
  jand g15007(.dina(n15226), .dinb(n15066), .dout(n15263));
  jor  g15008(.dina(n15263), .dinb(n15262), .dout(n15264));
  jor  g15009(.dina(n10049), .dinb(n1921), .dout(n15265));
  jor  g15010(.dina(n1806), .dinb(n9475), .dout(n15266));
  jor  g15011(.dina(n1923), .dinb(n10051), .dout(n15267));
  jor  g15012(.dina(n1918), .dinb(n9759), .dout(n15268));
  jand g15013(.dina(n15268), .dinb(n15267), .dout(n15269));
  jand g15014(.dina(n15269), .dinb(n15266), .dout(n15270));
  jand g15015(.dina(n15270), .dinb(n15265), .dout(n15271));
  jxor g15016(.dina(n15271), .dinb(n1687), .dout(n15272));
  jxor g15017(.dina(n15272), .dinb(n15264), .dout(n15273));
  jand g15018(.dina(n15077), .dinb(n15069), .dout(n15274));
  jand g15019(.dina(n15225), .dinb(n15078), .dout(n15275));
  jor  g15020(.dina(n15275), .dinb(n15274), .dout(n15276));
  jor  g15021(.dina(n9193), .dinb(n2324), .dout(n15277));
  jor  g15022(.dina(n2186), .dinb(n8644), .dout(n15278));
  jor  g15023(.dina(n2326), .dinb(n9195), .dout(n15279));
  jor  g15024(.dina(n2321), .dinb(n8920), .dout(n15280));
  jand g15025(.dina(n15280), .dinb(n15279), .dout(n15281));
  jand g15026(.dina(n15281), .dinb(n15278), .dout(n15282));
  jand g15027(.dina(n15282), .dinb(n15277), .dout(n15283));
  jxor g15028(.dina(n15283), .dinb(n2057), .dout(n15284));
  jxor g15029(.dina(n15284), .dinb(n15276), .dout(n15285));
  jand g15030(.dina(n15089), .dinb(n15081), .dout(n15286));
  jand g15031(.dina(n15224), .dinb(n15090), .dout(n15287));
  jor  g15032(.dina(n15287), .dinb(n15286), .dout(n15288));
  jor  g15033(.dina(n8376), .dinb(n2764), .dout(n15289));
  jor  g15034(.dina(n2609), .dinb(n7846), .dout(n15290));
  jor  g15035(.dina(n2761), .dinb(n8378), .dout(n15291));
  jor  g15036(.dina(n2766), .dinb(n8111), .dout(n15292));
  jand g15037(.dina(n15292), .dinb(n15291), .dout(n15293));
  jand g15038(.dina(n15293), .dinb(n15290), .dout(n15294));
  jand g15039(.dina(n15294), .dinb(n15289), .dout(n15295));
  jxor g15040(.dina(n15295), .dinb(n2468), .dout(n15296));
  jxor g15041(.dina(n15296), .dinb(n15288), .dout(n15297));
  jand g15042(.dina(n15214), .dinb(n15093), .dout(n15298));
  jand g15043(.dina(n15223), .dinb(n15215), .dout(n15299));
  jor  g15044(.dina(n15299), .dinb(n15298), .dout(n15300));
  jor  g15045(.dina(n7588), .dinb(n3239), .dout(n15301));
  jor  g15046(.dina(n3072), .dinb(n7086), .dout(n15302));
  jor  g15047(.dina(n3242), .dinb(n7338), .dout(n15303));
  jor  g15048(.dina(n3237), .dinb(n7590), .dout(n15304));
  jand g15049(.dina(n15304), .dinb(n15303), .dout(n15305));
  jand g15050(.dina(n15305), .dinb(n15302), .dout(n15306));
  jand g15051(.dina(n15306), .dinb(n15301), .dout(n15307));
  jxor g15052(.dina(n15307), .dinb(n2918), .dout(n15308));
  jxor g15053(.dina(n15308), .dinb(n15300), .dout(n15309));
  jand g15054(.dina(n15204), .dinb(n15096), .dout(n15310));
  jand g15055(.dina(n15213), .dinb(n15205), .dout(n15311));
  jor  g15056(.dina(n15311), .dinb(n15310), .dout(n15312));
  jand g15057(.dina(n15194), .dinb(n15099), .dout(n15313));
  jand g15058(.dina(n15203), .dinb(n15195), .dout(n15314));
  jor  g15059(.dina(n15314), .dinb(n15313), .dout(n15315));
  jand g15060(.dina(n15184), .dinb(n15102), .dout(n15316));
  jand g15061(.dina(n15193), .dinb(n15185), .dout(n15317));
  jor  g15062(.dina(n15317), .dinb(n15316), .dout(n15318));
  jand g15063(.dina(n15174), .dinb(n15105), .dout(n15319));
  jand g15064(.dina(n15183), .dinb(n15175), .dout(n15320));
  jor  g15065(.dina(n15320), .dinb(n15319), .dout(n15321));
  jand g15066(.dina(n15164), .dinb(n15108), .dout(n15322));
  jand g15067(.dina(n15173), .dinb(n15165), .dout(n15323));
  jor  g15068(.dina(n15323), .dinb(n15322), .dout(n15324));
  jand g15069(.dina(n15154), .dinb(n15151), .dout(n15325));
  jand g15070(.dina(n15163), .dinb(n15155), .dout(n15326));
  jor  g15071(.dina(n15326), .dinb(n15325), .dout(n15327));
  jand g15072(.dina(n15141), .dinb(n15111), .dout(n15328));
  jand g15073(.dina(n15150), .dinb(n15142), .dout(n15329));
  jor  g15074(.dina(n15329), .dinb(n15328), .dout(n15330));
  jand g15075(.dina(n15131), .dinb(n15128), .dout(n15331));
  jand g15076(.dina(n15140), .dinb(n15132), .dout(n15332));
  jor  g15077(.dina(n15332), .dinb(n15331), .dout(n15333));
  jand g15078(.dina(n15118), .dinb(n15115), .dout(n15334));
  jand g15079(.dina(n15127), .dinb(n15119), .dout(n15335));
  jor  g15080(.dina(n15335), .dinb(n15334), .dout(n15336));
  jand g15081(.dina(n10594), .dinb(b19 ), .dout(n15337));
  jand g15082(.dina(n10129), .dinb(b20 ), .dout(n15338));
  jor  g15083(.dina(n15338), .dinb(n15337), .dout(n15339));
  jnot g15084(.din(n15339), .dout(n15340));
  jxor g15085(.dina(n15340), .dinb(n15114), .dout(n15341));
  jor  g15086(.dina(n10134), .dinb(n1879), .dout(n15342));
  jor  g15087(.dina(n9849), .dinb(n1637), .dout(n15343));
  jor  g15088(.dina(n10137), .dinb(n1759), .dout(n15344));
  jor  g15089(.dina(n10132), .dinb(n1881), .dout(n15345));
  jand g15090(.dina(n15345), .dinb(n15344), .dout(n15346));
  jand g15091(.dina(n15346), .dinb(n15343), .dout(n15347));
  jand g15092(.dina(n15347), .dinb(n15342), .dout(n15348));
  jxor g15093(.dina(n15348), .dinb(n9559), .dout(n15349));
  jxor g15094(.dina(n15349), .dinb(n15341), .dout(n15350));
  jxor g15095(.dina(n15350), .dinb(n15336), .dout(n15351));
  jor  g15096(.dina(n9271), .dinb(n2277), .dout(n15352));
  jor  g15097(.dina(n9003), .dinb(n2007), .dout(n15353));
  jor  g15098(.dina(n9268), .dinb(n2279), .dout(n15354));
  jor  g15099(.dina(n9273), .dinb(n2142), .dout(n15355));
  jand g15100(.dina(n15355), .dinb(n15354), .dout(n15356));
  jand g15101(.dina(n15356), .dinb(n15353), .dout(n15357));
  jand g15102(.dina(n15357), .dinb(n15352), .dout(n15358));
  jxor g15103(.dina(n15358), .dinb(n8729), .dout(n15359));
  jxor g15104(.dina(n15359), .dinb(n15351), .dout(n15360));
  jxor g15105(.dina(n15360), .dinb(n15333), .dout(n15361));
  jor  g15106(.dina(n8457), .dinb(n2711), .dout(n15362));
  jor  g15107(.dina(n8185), .dinb(n2415), .dout(n15363));
  jor  g15108(.dina(n8459), .dinb(n2563), .dout(n15364));
  jor  g15109(.dina(n8454), .dinb(n2713), .dout(n15365));
  jand g15110(.dina(n15365), .dinb(n15364), .dout(n15366));
  jand g15111(.dina(n15366), .dinb(n15363), .dout(n15367));
  jand g15112(.dina(n15367), .dinb(n15362), .dout(n15368));
  jxor g15113(.dina(n15368), .dinb(n7929), .dout(n15369));
  jxor g15114(.dina(n15369), .dinb(n15361), .dout(n15370));
  jxor g15115(.dina(n15370), .dinb(n15330), .dout(n15371));
  jor  g15116(.dina(n7660), .dinb(n3184), .dout(n15372));
  jor  g15117(.dina(n7415), .dinb(n2862), .dout(n15373));
  jor  g15118(.dina(n7662), .dinb(n3186), .dout(n15374));
  jor  g15119(.dina(n7657), .dinb(n3023), .dout(n15375));
  jand g15120(.dina(n15375), .dinb(n15374), .dout(n15376));
  jand g15121(.dina(n15376), .dinb(n15373), .dout(n15377));
  jand g15122(.dina(n15377), .dinb(n15372), .dout(n15378));
  jxor g15123(.dina(n15378), .dinb(n7166), .dout(n15379));
  jxor g15124(.dina(n15379), .dinb(n15371), .dout(n15380));
  jxor g15125(.dina(n15380), .dinb(n15327), .dout(n15381));
  jor  g15126(.dina(n6914), .dinb(n3696), .dout(n15382));
  jor  g15127(.dina(n6673), .dinb(n3348), .dout(n15383));
  jor  g15128(.dina(n6916), .dinb(n3698), .dout(n15384));
  jor  g15129(.dina(n6911), .dinb(n3522), .dout(n15385));
  jand g15130(.dina(n15385), .dinb(n15384), .dout(n15386));
  jand g15131(.dina(n15386), .dinb(n15383), .dout(n15387));
  jand g15132(.dina(n15387), .dinb(n15382), .dout(n15388));
  jxor g15133(.dina(n15388), .dinb(n6443), .dout(n15389));
  jxor g15134(.dina(n15389), .dinb(n15381), .dout(n15390));
  jxor g15135(.dina(n15390), .dinb(n15324), .dout(n15391));
  jor  g15136(.dina(n6207), .dinb(n4247), .dout(n15392));
  jor  g15137(.dina(n5975), .dinb(n3873), .dout(n15393));
  jor  g15138(.dina(n6210), .dinb(n4060), .dout(n15394));
  jor  g15139(.dina(n6205), .dinb(n4249), .dout(n15395));
  jand g15140(.dina(n15395), .dinb(n15394), .dout(n15396));
  jand g15141(.dina(n15396), .dinb(n15393), .dout(n15397));
  jand g15142(.dina(n15397), .dinb(n15392), .dout(n15398));
  jxor g15143(.dina(n15398), .dinb(n5759), .dout(n15399));
  jxor g15144(.dina(n15399), .dinb(n15391), .dout(n15400));
  jxor g15145(.dina(n15400), .dinb(n15321), .dout(n15401));
  jor  g15146(.dina(n5537), .dinb(n4837), .dout(n15402));
  jor  g15147(.dina(n5315), .dinb(n4437), .dout(n15403));
  jor  g15148(.dina(n5534), .dinb(n4637), .dout(n15404));
  jor  g15149(.dina(n5539), .dinb(n4839), .dout(n15405));
  jand g15150(.dina(n15405), .dinb(n15404), .dout(n15406));
  jand g15151(.dina(n15406), .dinb(n15403), .dout(n15407));
  jand g15152(.dina(n15407), .dinb(n15402), .dout(n15408));
  jxor g15153(.dina(n15408), .dinb(n5111), .dout(n15409));
  jxor g15154(.dina(n15409), .dinb(n15401), .dout(n15410));
  jxor g15155(.dina(n15410), .dinb(n15318), .dout(n15411));
  jor  g15156(.dina(n5467), .dinb(n4902), .dout(n15412));
  jor  g15157(.dina(n4696), .dinb(n5040), .dout(n15413));
  jor  g15158(.dina(n4899), .dinb(n5469), .dout(n15414));
  jor  g15159(.dina(n4904), .dinb(n5253), .dout(n15415));
  jand g15160(.dina(n15415), .dinb(n15414), .dout(n15416));
  jand g15161(.dina(n15416), .dinb(n15413), .dout(n15417));
  jand g15162(.dina(n15417), .dinb(n15412), .dout(n15418));
  jxor g15163(.dina(n15418), .dinb(n4505), .dout(n15419));
  jxor g15164(.dina(n15419), .dinb(n15411), .dout(n15420));
  jxor g15165(.dina(n15420), .dinb(n15315), .dout(n15421));
  jor  g15166(.dina(n6137), .dinb(n4305), .dout(n15422));
  jor  g15167(.dina(n4116), .dinb(n5685), .dout(n15423));
  jor  g15168(.dina(n4308), .dinb(n5911), .dout(n15424));
  jor  g15169(.dina(n4303), .dinb(n6139), .dout(n15425));
  jand g15170(.dina(n15425), .dinb(n15424), .dout(n15426));
  jand g15171(.dina(n15426), .dinb(n15423), .dout(n15427));
  jand g15172(.dina(n15427), .dinb(n15422), .dout(n15428));
  jxor g15173(.dina(n15428), .dinb(n3938), .dout(n15429));
  jxor g15174(.dina(n15429), .dinb(n15421), .dout(n15430));
  jxor g15175(.dina(n15430), .dinb(n15312), .dout(n15431));
  jor  g15176(.dina(n6844), .dinb(n3751), .dout(n15432));
  jor  g15177(.dina(n3574), .dinb(n6366), .dout(n15433));
  jor  g15178(.dina(n3754), .dinb(n6605), .dout(n15434));
  jor  g15179(.dina(n3749), .dinb(n6846), .dout(n15435));
  jand g15180(.dina(n15435), .dinb(n15434), .dout(n15436));
  jand g15181(.dina(n15436), .dinb(n15433), .dout(n15437));
  jand g15182(.dina(n15437), .dinb(n15432), .dout(n15438));
  jxor g15183(.dina(n15438), .dinb(n3410), .dout(n15439));
  jxor g15184(.dina(n15439), .dinb(n15431), .dout(n15440));
  jxor g15185(.dina(n15440), .dinb(n15309), .dout(n15441));
  jxor g15186(.dina(n15441), .dinb(n15297), .dout(n15442));
  jxor g15187(.dina(n15442), .dinb(n15285), .dout(n15443));
  jxor g15188(.dina(n15443), .dinb(n15273), .dout(n15444));
  jxor g15189(.dina(n15444), .dinb(n15261), .dout(n15445));
  jxor g15190(.dina(n15445), .dinb(n15252), .dout(n15446));
  jnot g15191(.din(n15446), .dout(n15447));
  jxor g15192(.dina(n15447), .dinb(n15247), .dout(f83 ));
  jor  g15193(.dina(n15260), .dinb(n15256), .dout(n15449));
  jand g15194(.dina(n15444), .dinb(n15261), .dout(n15450));
  jnot g15195(.din(n15450), .dout(n15451));
  jand g15196(.dina(n15451), .dinb(n15449), .dout(n15452));
  jnot g15197(.din(n15452), .dout(n15453));
  jand g15198(.dina(n15272), .dinb(n15264), .dout(n15454));
  jand g15199(.dina(n15443), .dinb(n15273), .dout(n15455));
  jor  g15200(.dina(n15455), .dinb(n15454), .dout(n15456));
  jor  g15201(.dina(n10521), .dinb(n1921), .dout(n15457));
  jor  g15202(.dina(n1806), .dinb(n9759), .dout(n15458));
  jor  g15203(.dina(n1918), .dinb(n10051), .dout(n15459));
  jor  g15204(.dina(n1923), .dinb(n10523), .dout(n15460));
  jand g15205(.dina(n15460), .dinb(n15459), .dout(n15461));
  jand g15206(.dina(n15461), .dinb(n15458), .dout(n15462));
  jand g15207(.dina(n15462), .dinb(n15457), .dout(n15463));
  jxor g15208(.dina(n15463), .dinb(n1687), .dout(n15464));
  jxor g15209(.dina(n15464), .dinb(n15456), .dout(n15465));
  jand g15210(.dina(n15284), .dinb(n15276), .dout(n15466));
  jand g15211(.dina(n15442), .dinb(n15285), .dout(n15467));
  jor  g15212(.dina(n15467), .dinb(n15466), .dout(n15468));
  jor  g15213(.dina(n9473), .dinb(n2324), .dout(n15469));
  jor  g15214(.dina(n2186), .dinb(n8920), .dout(n15470));
  jor  g15215(.dina(n2326), .dinb(n9475), .dout(n15471));
  jor  g15216(.dina(n2321), .dinb(n9195), .dout(n15472));
  jand g15217(.dina(n15472), .dinb(n15471), .dout(n15473));
  jand g15218(.dina(n15473), .dinb(n15470), .dout(n15474));
  jand g15219(.dina(n15474), .dinb(n15469), .dout(n15475));
  jxor g15220(.dina(n15475), .dinb(n2057), .dout(n15476));
  jxor g15221(.dina(n15476), .dinb(n15468), .dout(n15477));
  jand g15222(.dina(n15296), .dinb(n15288), .dout(n15478));
  jand g15223(.dina(n15441), .dinb(n15297), .dout(n15479));
  jor  g15224(.dina(n15479), .dinb(n15478), .dout(n15480));
  jor  g15225(.dina(n8642), .dinb(n2764), .dout(n15481));
  jor  g15226(.dina(n2609), .dinb(n8111), .dout(n15482));
  jor  g15227(.dina(n2761), .dinb(n8644), .dout(n15483));
  jor  g15228(.dina(n2766), .dinb(n8378), .dout(n15484));
  jand g15229(.dina(n15484), .dinb(n15483), .dout(n15485));
  jand g15230(.dina(n15485), .dinb(n15482), .dout(n15486));
  jand g15231(.dina(n15486), .dinb(n15481), .dout(n15487));
  jxor g15232(.dina(n15487), .dinb(n2468), .dout(n15488));
  jxor g15233(.dina(n15488), .dinb(n15480), .dout(n15489));
  jand g15234(.dina(n15308), .dinb(n15300), .dout(n15490));
  jand g15235(.dina(n15440), .dinb(n15309), .dout(n15491));
  jor  g15236(.dina(n15491), .dinb(n15490), .dout(n15492));
  jor  g15237(.dina(n7844), .dinb(n3239), .dout(n15493));
  jor  g15238(.dina(n3072), .dinb(n7338), .dout(n15494));
  jor  g15239(.dina(n3242), .dinb(n7590), .dout(n15495));
  jor  g15240(.dina(n3237), .dinb(n7846), .dout(n15496));
  jand g15241(.dina(n15496), .dinb(n15495), .dout(n15497));
  jand g15242(.dina(n15497), .dinb(n15494), .dout(n15498));
  jand g15243(.dina(n15498), .dinb(n15493), .dout(n15499));
  jxor g15244(.dina(n15499), .dinb(n2918), .dout(n15500));
  jxor g15245(.dina(n15500), .dinb(n15492), .dout(n15501));
  jand g15246(.dina(n15430), .dinb(n15312), .dout(n15502));
  jand g15247(.dina(n15439), .dinb(n15431), .dout(n15503));
  jor  g15248(.dina(n15503), .dinb(n15502), .dout(n15504));
  jand g15249(.dina(n15420), .dinb(n15315), .dout(n15505));
  jand g15250(.dina(n15429), .dinb(n15421), .dout(n15506));
  jor  g15251(.dina(n15506), .dinb(n15505), .dout(n15507));
  jand g15252(.dina(n15410), .dinb(n15318), .dout(n15508));
  jand g15253(.dina(n15419), .dinb(n15411), .dout(n15509));
  jor  g15254(.dina(n15509), .dinb(n15508), .dout(n15510));
  jand g15255(.dina(n15400), .dinb(n15321), .dout(n15511));
  jand g15256(.dina(n15409), .dinb(n15401), .dout(n15512));
  jor  g15257(.dina(n15512), .dinb(n15511), .dout(n15513));
  jand g15258(.dina(n15390), .dinb(n15324), .dout(n15514));
  jand g15259(.dina(n15399), .dinb(n15391), .dout(n15515));
  jor  g15260(.dina(n15515), .dinb(n15514), .dout(n15516));
  jand g15261(.dina(n15380), .dinb(n15327), .dout(n15517));
  jand g15262(.dina(n15389), .dinb(n15381), .dout(n15518));
  jor  g15263(.dina(n15518), .dinb(n15517), .dout(n15519));
  jand g15264(.dina(n15360), .dinb(n15333), .dout(n15520));
  jand g15265(.dina(n15369), .dinb(n15361), .dout(n15521));
  jor  g15266(.dina(n15521), .dinb(n15520), .dout(n15522));
  jand g15267(.dina(n15350), .dinb(n15336), .dout(n15523));
  jand g15268(.dina(n15359), .dinb(n15351), .dout(n15524));
  jor  g15269(.dina(n15524), .dinb(n15523), .dout(n15525));
  jand g15270(.dina(n15340), .dinb(n15114), .dout(n15526));
  jand g15271(.dina(n15349), .dinb(n15341), .dout(n15527));
  jor  g15272(.dina(n15527), .dinb(n15526), .dout(n15528));
  jand g15273(.dina(n10594), .dinb(b20 ), .dout(n15529));
  jand g15274(.dina(n10129), .dinb(b21 ), .dout(n15530));
  jor  g15275(.dina(n15530), .dinb(n15529), .dout(n15531));
  jxor g15276(.dina(n15531), .dinb(n1351), .dout(n15532));
  jxor g15277(.dina(n15532), .dinb(n15339), .dout(n15533));
  jor  g15278(.dina(n10134), .dinb(n2005), .dout(n15534));
  jor  g15279(.dina(n9849), .dinb(n1759), .dout(n15535));
  jor  g15280(.dina(n10137), .dinb(n1881), .dout(n15536));
  jor  g15281(.dina(n10132), .dinb(n2007), .dout(n15537));
  jand g15282(.dina(n15537), .dinb(n15536), .dout(n15538));
  jand g15283(.dina(n15538), .dinb(n15535), .dout(n15539));
  jand g15284(.dina(n15539), .dinb(n15534), .dout(n15540));
  jxor g15285(.dina(n15540), .dinb(n9559), .dout(n15541));
  jxor g15286(.dina(n15541), .dinb(n15533), .dout(n15542));
  jxor g15287(.dina(n15542), .dinb(n15528), .dout(n15543));
  jor  g15288(.dina(n9271), .dinb(n2413), .dout(n15544));
  jor  g15289(.dina(n9003), .dinb(n2142), .dout(n15545));
  jor  g15290(.dina(n9273), .dinb(n2279), .dout(n15546));
  jor  g15291(.dina(n9268), .dinb(n2415), .dout(n15547));
  jand g15292(.dina(n15547), .dinb(n15546), .dout(n15548));
  jand g15293(.dina(n15548), .dinb(n15545), .dout(n15549));
  jand g15294(.dina(n15549), .dinb(n15544), .dout(n15550));
  jxor g15295(.dina(n15550), .dinb(n8729), .dout(n15551));
  jxor g15296(.dina(n15551), .dinb(n15543), .dout(n15552));
  jxor g15297(.dina(n15552), .dinb(n15525), .dout(n15553));
  jor  g15298(.dina(n8457), .dinb(n2860), .dout(n15554));
  jor  g15299(.dina(n8185), .dinb(n2563), .dout(n15555));
  jor  g15300(.dina(n8454), .dinb(n2862), .dout(n15556));
  jor  g15301(.dina(n8459), .dinb(n2713), .dout(n15557));
  jand g15302(.dina(n15557), .dinb(n15556), .dout(n15558));
  jand g15303(.dina(n15558), .dinb(n15555), .dout(n15559));
  jand g15304(.dina(n15559), .dinb(n15554), .dout(n15560));
  jxor g15305(.dina(n15560), .dinb(n7929), .dout(n15561));
  jxor g15306(.dina(n15561), .dinb(n15553), .dout(n15562));
  jxor g15307(.dina(n15562), .dinb(n15522), .dout(n15563));
  jand g15308(.dina(n15370), .dinb(n15330), .dout(n15564));
  jand g15309(.dina(n15379), .dinb(n15371), .dout(n15565));
  jor  g15310(.dina(n15565), .dinb(n15564), .dout(n15566));
  jor  g15311(.dina(n7660), .dinb(n3346), .dout(n15567));
  jor  g15312(.dina(n7415), .dinb(n3023), .dout(n15568));
  jor  g15313(.dina(n7662), .dinb(n3348), .dout(n15569));
  jor  g15314(.dina(n7657), .dinb(n3186), .dout(n15570));
  jand g15315(.dina(n15570), .dinb(n15569), .dout(n15571));
  jand g15316(.dina(n15571), .dinb(n15568), .dout(n15572));
  jand g15317(.dina(n15572), .dinb(n15567), .dout(n15573));
  jxor g15318(.dina(n15573), .dinb(n7166), .dout(n15574));
  jxor g15319(.dina(n15574), .dinb(n15566), .dout(n15575));
  jxor g15320(.dina(n15575), .dinb(n15563), .dout(n15576));
  jor  g15321(.dina(n6914), .dinb(n3871), .dout(n15577));
  jor  g15322(.dina(n6673), .dinb(n3522), .dout(n15578));
  jor  g15323(.dina(n6916), .dinb(n3873), .dout(n15579));
  jor  g15324(.dina(n6911), .dinb(n3698), .dout(n15580));
  jand g15325(.dina(n15580), .dinb(n15579), .dout(n15581));
  jand g15326(.dina(n15581), .dinb(n15578), .dout(n15582));
  jand g15327(.dina(n15582), .dinb(n15577), .dout(n15583));
  jxor g15328(.dina(n15583), .dinb(n6443), .dout(n15584));
  jxor g15329(.dina(n15584), .dinb(n15576), .dout(n15585));
  jxor g15330(.dina(n15585), .dinb(n15519), .dout(n15586));
  jor  g15331(.dina(n6207), .dinb(n4435), .dout(n15587));
  jor  g15332(.dina(n5975), .dinb(n4060), .dout(n15588));
  jor  g15333(.dina(n6205), .dinb(n4437), .dout(n15589));
  jor  g15334(.dina(n6210), .dinb(n4249), .dout(n15590));
  jand g15335(.dina(n15590), .dinb(n15589), .dout(n15591));
  jand g15336(.dina(n15591), .dinb(n15588), .dout(n15592));
  jand g15337(.dina(n15592), .dinb(n15587), .dout(n15593));
  jxor g15338(.dina(n15593), .dinb(n5759), .dout(n15594));
  jxor g15339(.dina(n15594), .dinb(n15586), .dout(n15595));
  jxor g15340(.dina(n15595), .dinb(n15516), .dout(n15596));
  jor  g15341(.dina(n5537), .dinb(n5038), .dout(n15597));
  jor  g15342(.dina(n5315), .dinb(n4637), .dout(n15598));
  jor  g15343(.dina(n5534), .dinb(n4839), .dout(n15599));
  jor  g15344(.dina(n5539), .dinb(n5040), .dout(n15600));
  jand g15345(.dina(n15600), .dinb(n15599), .dout(n15601));
  jand g15346(.dina(n15601), .dinb(n15598), .dout(n15602));
  jand g15347(.dina(n15602), .dinb(n15597), .dout(n15603));
  jxor g15348(.dina(n15603), .dinb(n5111), .dout(n15604));
  jxor g15349(.dina(n15604), .dinb(n15596), .dout(n15605));
  jxor g15350(.dina(n15605), .dinb(n15513), .dout(n15606));
  jor  g15351(.dina(n5683), .dinb(n4902), .dout(n15607));
  jor  g15352(.dina(n4696), .dinb(n5253), .dout(n15608));
  jor  g15353(.dina(n4904), .dinb(n5469), .dout(n15609));
  jor  g15354(.dina(n4899), .dinb(n5685), .dout(n15610));
  jand g15355(.dina(n15610), .dinb(n15609), .dout(n15611));
  jand g15356(.dina(n15611), .dinb(n15608), .dout(n15612));
  jand g15357(.dina(n15612), .dinb(n15607), .dout(n15613));
  jxor g15358(.dina(n15613), .dinb(n4505), .dout(n15614));
  jxor g15359(.dina(n15614), .dinb(n15606), .dout(n15615));
  jxor g15360(.dina(n15615), .dinb(n15510), .dout(n15616));
  jor  g15361(.dina(n6364), .dinb(n4305), .dout(n15617));
  jor  g15362(.dina(n4116), .dinb(n5911), .dout(n15618));
  jor  g15363(.dina(n4308), .dinb(n6139), .dout(n15619));
  jor  g15364(.dina(n4303), .dinb(n6366), .dout(n15620));
  jand g15365(.dina(n15620), .dinb(n15619), .dout(n15621));
  jand g15366(.dina(n15621), .dinb(n15618), .dout(n15622));
  jand g15367(.dina(n15622), .dinb(n15617), .dout(n15623));
  jxor g15368(.dina(n15623), .dinb(n3938), .dout(n15624));
  jxor g15369(.dina(n15624), .dinb(n15616), .dout(n15625));
  jxor g15370(.dina(n15625), .dinb(n15507), .dout(n15626));
  jor  g15371(.dina(n7084), .dinb(n3751), .dout(n15627));
  jor  g15372(.dina(n3574), .dinb(n6605), .dout(n15628));
  jor  g15373(.dina(n3749), .dinb(n7086), .dout(n15629));
  jor  g15374(.dina(n3754), .dinb(n6846), .dout(n15630));
  jand g15375(.dina(n15630), .dinb(n15629), .dout(n15631));
  jand g15376(.dina(n15631), .dinb(n15628), .dout(n15632));
  jand g15377(.dina(n15632), .dinb(n15627), .dout(n15633));
  jxor g15378(.dina(n15633), .dinb(n3410), .dout(n15634));
  jxor g15379(.dina(n15634), .dinb(n15626), .dout(n15635));
  jxor g15380(.dina(n15635), .dinb(n15504), .dout(n15636));
  jxor g15381(.dina(n15636), .dinb(n15501), .dout(n15637));
  jxor g15382(.dina(n15637), .dinb(n15489), .dout(n15638));
  jxor g15383(.dina(n15638), .dinb(n15477), .dout(n15639));
  jxor g15384(.dina(n15639), .dinb(n15465), .dout(n15640));
  jxor g15385(.dina(n15640), .dinb(n15453), .dout(n15641));
  jnot g15386(.din(n15641), .dout(n15642));
  jand g15387(.dina(n15445), .dinb(n15252), .dout(n15643));
  jnot g15388(.din(n15643), .dout(n15644));
  jor  g15389(.dina(n15447), .dinb(n15247), .dout(n15645));
  jand g15390(.dina(n15645), .dinb(n15644), .dout(n15646));
  jxor g15391(.dina(n15646), .dinb(n15642), .dout(f84 ));
  jand g15392(.dina(n15464), .dinb(n15456), .dout(n15648));
  jand g15393(.dina(n15639), .dinb(n15465), .dout(n15649));
  jor  g15394(.dina(n15649), .dinb(n15648), .dout(n15650));
  jand g15395(.dina(n15476), .dinb(n15468), .dout(n15651));
  jand g15396(.dina(n15638), .dinb(n15477), .dout(n15652));
  jor  g15397(.dina(n15652), .dinb(n15651), .dout(n15653));
  jor  g15398(.dina(n10813), .dinb(n1921), .dout(n15654));
  jor  g15399(.dina(n1806), .dinb(n10051), .dout(n15655));
  jor  g15400(.dina(n1918), .dinb(n10523), .dout(n15656));
  jand g15401(.dina(n15656), .dinb(n15655), .dout(n15657));
  jand g15402(.dina(n15657), .dinb(n15654), .dout(n15658));
  jxor g15403(.dina(n15658), .dinb(n1687), .dout(n15659));
  jxor g15404(.dina(n15659), .dinb(n15653), .dout(n15660));
  jand g15405(.dina(n15488), .dinb(n15480), .dout(n15661));
  jand g15406(.dina(n15637), .dinb(n15489), .dout(n15662));
  jor  g15407(.dina(n15662), .dinb(n15661), .dout(n15663));
  jor  g15408(.dina(n9757), .dinb(n2324), .dout(n15664));
  jor  g15409(.dina(n2186), .dinb(n9195), .dout(n15665));
  jor  g15410(.dina(n2321), .dinb(n9475), .dout(n15666));
  jor  g15411(.dina(n2326), .dinb(n9759), .dout(n15667));
  jand g15412(.dina(n15667), .dinb(n15666), .dout(n15668));
  jand g15413(.dina(n15668), .dinb(n15665), .dout(n15669));
  jand g15414(.dina(n15669), .dinb(n15664), .dout(n15670));
  jxor g15415(.dina(n15670), .dinb(n2057), .dout(n15671));
  jxor g15416(.dina(n15671), .dinb(n15663), .dout(n15672));
  jand g15417(.dina(n15500), .dinb(n15492), .dout(n15673));
  jand g15418(.dina(n15636), .dinb(n15501), .dout(n15674));
  jor  g15419(.dina(n15674), .dinb(n15673), .dout(n15675));
  jor  g15420(.dina(n8918), .dinb(n2764), .dout(n15676));
  jor  g15421(.dina(n2609), .dinb(n8378), .dout(n15677));
  jor  g15422(.dina(n2761), .dinb(n8920), .dout(n15678));
  jor  g15423(.dina(n2766), .dinb(n8644), .dout(n15679));
  jand g15424(.dina(n15679), .dinb(n15678), .dout(n15680));
  jand g15425(.dina(n15680), .dinb(n15677), .dout(n15681));
  jand g15426(.dina(n15681), .dinb(n15676), .dout(n15682));
  jxor g15427(.dina(n15682), .dinb(n2468), .dout(n15683));
  jxor g15428(.dina(n15683), .dinb(n15675), .dout(n15684));
  jand g15429(.dina(n15624), .dinb(n15616), .dout(n15685));
  jand g15430(.dina(n15625), .dinb(n15507), .dout(n15686));
  jor  g15431(.dina(n15686), .dinb(n15685), .dout(n15687));
  jand g15432(.dina(n15614), .dinb(n15606), .dout(n15688));
  jand g15433(.dina(n15615), .dinb(n15510), .dout(n15689));
  jor  g15434(.dina(n15689), .dinb(n15688), .dout(n15690));
  jand g15435(.dina(n15604), .dinb(n15596), .dout(n15691));
  jand g15436(.dina(n15605), .dinb(n15513), .dout(n15692));
  jor  g15437(.dina(n15692), .dinb(n15691), .dout(n15693));
  jand g15438(.dina(n15594), .dinb(n15586), .dout(n15694));
  jand g15439(.dina(n15595), .dinb(n15516), .dout(n15695));
  jor  g15440(.dina(n15695), .dinb(n15694), .dout(n15696));
  jand g15441(.dina(n15584), .dinb(n15576), .dout(n15697));
  jand g15442(.dina(n15585), .dinb(n15519), .dout(n15698));
  jor  g15443(.dina(n15698), .dinb(n15697), .dout(n15699));
  jand g15444(.dina(n15574), .dinb(n15566), .dout(n15700));
  jand g15445(.dina(n15575), .dinb(n15563), .dout(n15701));
  jor  g15446(.dina(n15701), .dinb(n15700), .dout(n15702));
  jand g15447(.dina(n15561), .dinb(n15553), .dout(n15703));
  jand g15448(.dina(n15562), .dinb(n15522), .dout(n15704));
  jor  g15449(.dina(n15704), .dinb(n15703), .dout(n15705));
  jand g15450(.dina(n15551), .dinb(n15543), .dout(n15706));
  jand g15451(.dina(n15552), .dinb(n15525), .dout(n15707));
  jor  g15452(.dina(n15707), .dinb(n15706), .dout(n15708));
  jand g15453(.dina(n15541), .dinb(n15533), .dout(n15709));
  jand g15454(.dina(n15542), .dinb(n15528), .dout(n15710));
  jor  g15455(.dina(n15710), .dinb(n15709), .dout(n15711));
  jand g15456(.dina(n10594), .dinb(b21 ), .dout(n15712));
  jand g15457(.dina(n10129), .dinb(b22 ), .dout(n15713));
  jor  g15458(.dina(n15713), .dinb(n15712), .dout(n15714));
  jnot g15459(.din(n15714), .dout(n15715));
  jand g15460(.dina(n15531), .dinb(n1351), .dout(n15716));
  jand g15461(.dina(n15532), .dinb(n15339), .dout(n15717));
  jor  g15462(.dina(n15717), .dinb(n15716), .dout(n15718));
  jxor g15463(.dina(n15718), .dinb(n15715), .dout(n15719));
  jor  g15464(.dina(n10134), .dinb(n2140), .dout(n15720));
  jor  g15465(.dina(n9849), .dinb(n1881), .dout(n15721));
  jor  g15466(.dina(n10137), .dinb(n2007), .dout(n15722));
  jor  g15467(.dina(n10132), .dinb(n2142), .dout(n15723));
  jand g15468(.dina(n15723), .dinb(n15722), .dout(n15724));
  jand g15469(.dina(n15724), .dinb(n15721), .dout(n15725));
  jand g15470(.dina(n15725), .dinb(n15720), .dout(n15726));
  jxor g15471(.dina(n15726), .dinb(n9559), .dout(n15727));
  jxor g15472(.dina(n15727), .dinb(n15719), .dout(n15728));
  jxor g15473(.dina(n15728), .dinb(n15711), .dout(n15729));
  jor  g15474(.dina(n9271), .dinb(n2561), .dout(n15730));
  jor  g15475(.dina(n9003), .dinb(n2279), .dout(n15731));
  jor  g15476(.dina(n9268), .dinb(n2563), .dout(n15732));
  jor  g15477(.dina(n9273), .dinb(n2415), .dout(n15733));
  jand g15478(.dina(n15733), .dinb(n15732), .dout(n15734));
  jand g15479(.dina(n15734), .dinb(n15731), .dout(n15735));
  jand g15480(.dina(n15735), .dinb(n15730), .dout(n15736));
  jxor g15481(.dina(n15736), .dinb(n8729), .dout(n15737));
  jxor g15482(.dina(n15737), .dinb(n15729), .dout(n15738));
  jxor g15483(.dina(n15738), .dinb(n15708), .dout(n15739));
  jor  g15484(.dina(n8457), .dinb(n3021), .dout(n15740));
  jor  g15485(.dina(n8185), .dinb(n2713), .dout(n15741));
  jor  g15486(.dina(n8454), .dinb(n3023), .dout(n15742));
  jor  g15487(.dina(n8459), .dinb(n2862), .dout(n15743));
  jand g15488(.dina(n15743), .dinb(n15742), .dout(n15744));
  jand g15489(.dina(n15744), .dinb(n15741), .dout(n15745));
  jand g15490(.dina(n15745), .dinb(n15740), .dout(n15746));
  jxor g15491(.dina(n15746), .dinb(n7929), .dout(n15747));
  jxor g15492(.dina(n15747), .dinb(n15739), .dout(n15748));
  jxor g15493(.dina(n15748), .dinb(n15705), .dout(n15749));
  jor  g15494(.dina(n7660), .dinb(n3520), .dout(n15750));
  jor  g15495(.dina(n7415), .dinb(n3186), .dout(n15751));
  jor  g15496(.dina(n7657), .dinb(n3348), .dout(n15752));
  jor  g15497(.dina(n7662), .dinb(n3522), .dout(n15753));
  jand g15498(.dina(n15753), .dinb(n15752), .dout(n15754));
  jand g15499(.dina(n15754), .dinb(n15751), .dout(n15755));
  jand g15500(.dina(n15755), .dinb(n15750), .dout(n15756));
  jxor g15501(.dina(n15756), .dinb(n7166), .dout(n15757));
  jxor g15502(.dina(n15757), .dinb(n15749), .dout(n15758));
  jxor g15503(.dina(n15758), .dinb(n15702), .dout(n15759));
  jor  g15504(.dina(n6914), .dinb(n4058), .dout(n15760));
  jor  g15505(.dina(n6673), .dinb(n3698), .dout(n15761));
  jor  g15506(.dina(n6911), .dinb(n3873), .dout(n15762));
  jor  g15507(.dina(n6916), .dinb(n4060), .dout(n15763));
  jand g15508(.dina(n15763), .dinb(n15762), .dout(n15764));
  jand g15509(.dina(n15764), .dinb(n15761), .dout(n15765));
  jand g15510(.dina(n15765), .dinb(n15760), .dout(n15766));
  jxor g15511(.dina(n15766), .dinb(n6443), .dout(n15767));
  jxor g15512(.dina(n15767), .dinb(n15759), .dout(n15768));
  jxor g15513(.dina(n15768), .dinb(n15699), .dout(n15769));
  jor  g15514(.dina(n6207), .dinb(n4635), .dout(n15770));
  jor  g15515(.dina(n5975), .dinb(n4249), .dout(n15771));
  jor  g15516(.dina(n6205), .dinb(n4637), .dout(n15772));
  jor  g15517(.dina(n6210), .dinb(n4437), .dout(n15773));
  jand g15518(.dina(n15773), .dinb(n15772), .dout(n15774));
  jand g15519(.dina(n15774), .dinb(n15771), .dout(n15775));
  jand g15520(.dina(n15775), .dinb(n15770), .dout(n15776));
  jxor g15521(.dina(n15776), .dinb(n5759), .dout(n15777));
  jxor g15522(.dina(n15777), .dinb(n15769), .dout(n15778));
  jxor g15523(.dina(n15778), .dinb(n15696), .dout(n15779));
  jor  g15524(.dina(n5251), .dinb(n5537), .dout(n15780));
  jor  g15525(.dina(n5315), .dinb(n4839), .dout(n15781));
  jor  g15526(.dina(n5539), .dinb(n5253), .dout(n15782));
  jor  g15527(.dina(n5534), .dinb(n5040), .dout(n15783));
  jand g15528(.dina(n15783), .dinb(n15782), .dout(n15784));
  jand g15529(.dina(n15784), .dinb(n15781), .dout(n15785));
  jand g15530(.dina(n15785), .dinb(n15780), .dout(n15786));
  jxor g15531(.dina(n15786), .dinb(n5111), .dout(n15787));
  jxor g15532(.dina(n15787), .dinb(n15779), .dout(n15788));
  jxor g15533(.dina(n15788), .dinb(n15693), .dout(n15789));
  jor  g15534(.dina(n5909), .dinb(n4902), .dout(n15790));
  jor  g15535(.dina(n4696), .dinb(n5469), .dout(n15791));
  jor  g15536(.dina(n4904), .dinb(n5685), .dout(n15792));
  jor  g15537(.dina(n4899), .dinb(n5911), .dout(n15793));
  jand g15538(.dina(n15793), .dinb(n15792), .dout(n15794));
  jand g15539(.dina(n15794), .dinb(n15791), .dout(n15795));
  jand g15540(.dina(n15795), .dinb(n15790), .dout(n15796));
  jxor g15541(.dina(n15796), .dinb(n4505), .dout(n15797));
  jxor g15542(.dina(n15797), .dinb(n15789), .dout(n15798));
  jxor g15543(.dina(n15798), .dinb(n15690), .dout(n15799));
  jor  g15544(.dina(n6603), .dinb(n4305), .dout(n15800));
  jor  g15545(.dina(n4116), .dinb(n6139), .dout(n15801));
  jor  g15546(.dina(n4303), .dinb(n6605), .dout(n15802));
  jor  g15547(.dina(n4308), .dinb(n6366), .dout(n15803));
  jand g15548(.dina(n15803), .dinb(n15802), .dout(n15804));
  jand g15549(.dina(n15804), .dinb(n15801), .dout(n15805));
  jand g15550(.dina(n15805), .dinb(n15800), .dout(n15806));
  jxor g15551(.dina(n15806), .dinb(n3938), .dout(n15807));
  jxor g15552(.dina(n15807), .dinb(n15799), .dout(n15808));
  jxor g15553(.dina(n15808), .dinb(n15687), .dout(n15809));
  jor  g15554(.dina(n7336), .dinb(n3751), .dout(n15810));
  jor  g15555(.dina(n3574), .dinb(n6846), .dout(n15811));
  jor  g15556(.dina(n3754), .dinb(n7086), .dout(n15812));
  jor  g15557(.dina(n3749), .dinb(n7338), .dout(n15813));
  jand g15558(.dina(n15813), .dinb(n15812), .dout(n15814));
  jand g15559(.dina(n15814), .dinb(n15811), .dout(n15815));
  jand g15560(.dina(n15815), .dinb(n15810), .dout(n15816));
  jxor g15561(.dina(n15816), .dinb(n3410), .dout(n15817));
  jxor g15562(.dina(n15817), .dinb(n15809), .dout(n15818));
  jor  g15563(.dina(n8109), .dinb(n3239), .dout(n15819));
  jor  g15564(.dina(n3072), .dinb(n7590), .dout(n15820));
  jor  g15565(.dina(n3242), .dinb(n7846), .dout(n15821));
  jor  g15566(.dina(n3237), .dinb(n8111), .dout(n15822));
  jand g15567(.dina(n15822), .dinb(n15821), .dout(n15823));
  jand g15568(.dina(n15823), .dinb(n15820), .dout(n15824));
  jand g15569(.dina(n15824), .dinb(n15819), .dout(n15825));
  jxor g15570(.dina(n15825), .dinb(n2918), .dout(n15826));
  jnot g15571(.din(n15626), .dout(n15827));
  jnot g15572(.din(n15634), .dout(n15828));
  jand g15573(.dina(n15828), .dinb(n15827), .dout(n15829));
  jnot g15574(.din(n15829), .dout(n15830));
  jand g15575(.dina(n15634), .dinb(n15626), .dout(n15831));
  jor  g15576(.dina(n15831), .dinb(n15504), .dout(n15832));
  jand g15577(.dina(n15832), .dinb(n15830), .dout(n15833));
  jxor g15578(.dina(n15833), .dinb(n15826), .dout(n15834));
  jxor g15579(.dina(n15834), .dinb(n15818), .dout(n15835));
  jxor g15580(.dina(n15835), .dinb(n15684), .dout(n15836));
  jxor g15581(.dina(n15836), .dinb(n15672), .dout(n15837));
  jxor g15582(.dina(n15837), .dinb(n15660), .dout(n15838));
  jxor g15583(.dina(n15838), .dinb(n15650), .dout(n15839));
  jnot g15584(.din(n15839), .dout(n15840));
  jand g15585(.dina(n15640), .dinb(n15453), .dout(n15841));
  jnot g15586(.din(n15841), .dout(n15842));
  jor  g15587(.dina(n15646), .dinb(n15642), .dout(n15843));
  jand g15588(.dina(n15843), .dinb(n15842), .dout(n15844));
  jxor g15589(.dina(n15844), .dinb(n15840), .dout(f85 ));
  jand g15590(.dina(n15838), .dinb(n15650), .dout(n15846));
  jnot g15591(.din(n15846), .dout(n15847));
  jor  g15592(.dina(n15844), .dinb(n15840), .dout(n15848));
  jand g15593(.dina(n15848), .dinb(n15847), .dout(n15849));
  jand g15594(.dina(n15659), .dinb(n15653), .dout(n15850));
  jand g15595(.dina(n15837), .dinb(n15660), .dout(n15851));
  jor  g15596(.dina(n15851), .dinb(n15850), .dout(n15852));
  jand g15597(.dina(n15671), .dinb(n15663), .dout(n15853));
  jand g15598(.dina(n15836), .dinb(n15672), .dout(n15854));
  jor  g15599(.dina(n15854), .dinb(n15853), .dout(n15855));
  jnot g15600(.din(n15855), .dout(n15856));
  jand g15601(.dina(n1807), .dinb(b63 ), .dout(n15857));
  jand g15602(.dina(n10832), .dinb(n1676), .dout(n15858));
  jor  g15603(.dina(n15858), .dinb(n15857), .dout(n15859));
  jxor g15604(.dina(n15859), .dinb(n1687), .dout(n15860));
  jxor g15605(.dina(n15860), .dinb(n15856), .dout(n15861));
  jand g15606(.dina(n15683), .dinb(n15675), .dout(n15862));
  jand g15607(.dina(n15835), .dinb(n15684), .dout(n15863));
  jor  g15608(.dina(n15863), .dinb(n15862), .dout(n15864));
  jor  g15609(.dina(n10049), .dinb(n2324), .dout(n15865));
  jor  g15610(.dina(n2186), .dinb(n9475), .dout(n15866));
  jor  g15611(.dina(n2321), .dinb(n9759), .dout(n15867));
  jor  g15612(.dina(n2326), .dinb(n10051), .dout(n15868));
  jand g15613(.dina(n15868), .dinb(n15867), .dout(n15869));
  jand g15614(.dina(n15869), .dinb(n15866), .dout(n15870));
  jand g15615(.dina(n15870), .dinb(n15865), .dout(n15871));
  jxor g15616(.dina(n15871), .dinb(n2057), .dout(n15872));
  jxor g15617(.dina(n15872), .dinb(n15864), .dout(n15873));
  jand g15618(.dina(n15808), .dinb(n15687), .dout(n15874));
  jand g15619(.dina(n15817), .dinb(n15809), .dout(n15875));
  jor  g15620(.dina(n15875), .dinb(n15874), .dout(n15876));
  jor  g15621(.dina(n8376), .dinb(n3239), .dout(n15877));
  jor  g15622(.dina(n3072), .dinb(n7846), .dout(n15878));
  jor  g15623(.dina(n3237), .dinb(n8378), .dout(n15879));
  jor  g15624(.dina(n3242), .dinb(n8111), .dout(n15880));
  jand g15625(.dina(n15880), .dinb(n15879), .dout(n15881));
  jand g15626(.dina(n15881), .dinb(n15878), .dout(n15882));
  jand g15627(.dina(n15882), .dinb(n15877), .dout(n15883));
  jxor g15628(.dina(n15883), .dinb(n2918), .dout(n15884));
  jxor g15629(.dina(n15884), .dinb(n15876), .dout(n15885));
  jand g15630(.dina(n15798), .dinb(n15690), .dout(n15886));
  jand g15631(.dina(n15807), .dinb(n15799), .dout(n15887));
  jor  g15632(.dina(n15887), .dinb(n15886), .dout(n15888));
  jand g15633(.dina(n15788), .dinb(n15693), .dout(n15889));
  jand g15634(.dina(n15797), .dinb(n15789), .dout(n15890));
  jor  g15635(.dina(n15890), .dinb(n15889), .dout(n15891));
  jand g15636(.dina(n15778), .dinb(n15696), .dout(n15892));
  jand g15637(.dina(n15787), .dinb(n15779), .dout(n15893));
  jor  g15638(.dina(n15893), .dinb(n15892), .dout(n15894));
  jand g15639(.dina(n15768), .dinb(n15699), .dout(n15895));
  jand g15640(.dina(n15777), .dinb(n15769), .dout(n15896));
  jor  g15641(.dina(n15896), .dinb(n15895), .dout(n15897));
  jand g15642(.dina(n15758), .dinb(n15702), .dout(n15898));
  jand g15643(.dina(n15767), .dinb(n15759), .dout(n15899));
  jor  g15644(.dina(n15899), .dinb(n15898), .dout(n15900));
  jand g15645(.dina(n15748), .dinb(n15705), .dout(n15901));
  jand g15646(.dina(n15757), .dinb(n15749), .dout(n15902));
  jor  g15647(.dina(n15902), .dinb(n15901), .dout(n15903));
  jand g15648(.dina(n15738), .dinb(n15708), .dout(n15904));
  jand g15649(.dina(n15747), .dinb(n15739), .dout(n15905));
  jor  g15650(.dina(n15905), .dinb(n15904), .dout(n15906));
  jand g15651(.dina(n15728), .dinb(n15711), .dout(n15907));
  jand g15652(.dina(n15737), .dinb(n15729), .dout(n15908));
  jor  g15653(.dina(n15908), .dinb(n15907), .dout(n15909));
  jand g15654(.dina(n15718), .dinb(n15715), .dout(n15910));
  jand g15655(.dina(n15727), .dinb(n15719), .dout(n15911));
  jor  g15656(.dina(n15911), .dinb(n15910), .dout(n15912));
  jand g15657(.dina(n10594), .dinb(b22 ), .dout(n15913));
  jand g15658(.dina(n10129), .dinb(b23 ), .dout(n15914));
  jor  g15659(.dina(n15914), .dinb(n15913), .dout(n15915));
  jnot g15660(.din(n15915), .dout(n15916));
  jxor g15661(.dina(n15916), .dinb(n15714), .dout(n15917));
  jor  g15662(.dina(n10134), .dinb(n2277), .dout(n15918));
  jor  g15663(.dina(n9849), .dinb(n2007), .dout(n15919));
  jor  g15664(.dina(n10137), .dinb(n2142), .dout(n15920));
  jor  g15665(.dina(n10132), .dinb(n2279), .dout(n15921));
  jand g15666(.dina(n15921), .dinb(n15920), .dout(n15922));
  jand g15667(.dina(n15922), .dinb(n15919), .dout(n15923));
  jand g15668(.dina(n15923), .dinb(n15918), .dout(n15924));
  jxor g15669(.dina(n15924), .dinb(n9559), .dout(n15925));
  jxor g15670(.dina(n15925), .dinb(n15917), .dout(n15926));
  jxor g15671(.dina(n15926), .dinb(n15912), .dout(n15927));
  jor  g15672(.dina(n9271), .dinb(n2711), .dout(n15928));
  jor  g15673(.dina(n9003), .dinb(n2415), .dout(n15929));
  jor  g15674(.dina(n9268), .dinb(n2713), .dout(n15930));
  jor  g15675(.dina(n9273), .dinb(n2563), .dout(n15931));
  jand g15676(.dina(n15931), .dinb(n15930), .dout(n15932));
  jand g15677(.dina(n15932), .dinb(n15929), .dout(n15933));
  jand g15678(.dina(n15933), .dinb(n15928), .dout(n15934));
  jxor g15679(.dina(n15934), .dinb(n8729), .dout(n15935));
  jxor g15680(.dina(n15935), .dinb(n15927), .dout(n15936));
  jxor g15681(.dina(n15936), .dinb(n15909), .dout(n15937));
  jor  g15682(.dina(n8457), .dinb(n3184), .dout(n15938));
  jor  g15683(.dina(n8185), .dinb(n2862), .dout(n15939));
  jor  g15684(.dina(n8459), .dinb(n3023), .dout(n15940));
  jor  g15685(.dina(n8454), .dinb(n3186), .dout(n15941));
  jand g15686(.dina(n15941), .dinb(n15940), .dout(n15942));
  jand g15687(.dina(n15942), .dinb(n15939), .dout(n15943));
  jand g15688(.dina(n15943), .dinb(n15938), .dout(n15944));
  jxor g15689(.dina(n15944), .dinb(n7929), .dout(n15945));
  jxor g15690(.dina(n15945), .dinb(n15937), .dout(n15946));
  jxor g15691(.dina(n15946), .dinb(n15906), .dout(n15947));
  jor  g15692(.dina(n7660), .dinb(n3696), .dout(n15948));
  jor  g15693(.dina(n7415), .dinb(n3348), .dout(n15949));
  jor  g15694(.dina(n7657), .dinb(n3522), .dout(n15950));
  jor  g15695(.dina(n7662), .dinb(n3698), .dout(n15951));
  jand g15696(.dina(n15951), .dinb(n15950), .dout(n15952));
  jand g15697(.dina(n15952), .dinb(n15949), .dout(n15953));
  jand g15698(.dina(n15953), .dinb(n15948), .dout(n15954));
  jxor g15699(.dina(n15954), .dinb(n7166), .dout(n15955));
  jxor g15700(.dina(n15955), .dinb(n15947), .dout(n15956));
  jxor g15701(.dina(n15956), .dinb(n15903), .dout(n15957));
  jor  g15702(.dina(n6914), .dinb(n4247), .dout(n15958));
  jor  g15703(.dina(n6673), .dinb(n3873), .dout(n15959));
  jor  g15704(.dina(n6911), .dinb(n4060), .dout(n15960));
  jor  g15705(.dina(n6916), .dinb(n4249), .dout(n15961));
  jand g15706(.dina(n15961), .dinb(n15960), .dout(n15962));
  jand g15707(.dina(n15962), .dinb(n15959), .dout(n15963));
  jand g15708(.dina(n15963), .dinb(n15958), .dout(n15964));
  jxor g15709(.dina(n15964), .dinb(n6443), .dout(n15965));
  jxor g15710(.dina(n15965), .dinb(n15957), .dout(n15966));
  jxor g15711(.dina(n15966), .dinb(n15900), .dout(n15967));
  jor  g15712(.dina(n6207), .dinb(n4837), .dout(n15968));
  jor  g15713(.dina(n5975), .dinb(n4437), .dout(n15969));
  jor  g15714(.dina(n6210), .dinb(n4637), .dout(n15970));
  jor  g15715(.dina(n6205), .dinb(n4839), .dout(n15971));
  jand g15716(.dina(n15971), .dinb(n15970), .dout(n15972));
  jand g15717(.dina(n15972), .dinb(n15969), .dout(n15973));
  jand g15718(.dina(n15973), .dinb(n15968), .dout(n15974));
  jxor g15719(.dina(n15974), .dinb(n5759), .dout(n15975));
  jxor g15720(.dina(n15975), .dinb(n15967), .dout(n15976));
  jxor g15721(.dina(n15976), .dinb(n15897), .dout(n15977));
  jor  g15722(.dina(n5467), .dinb(n5537), .dout(n15978));
  jor  g15723(.dina(n5315), .dinb(n5040), .dout(n15979));
  jor  g15724(.dina(n5539), .dinb(n5469), .dout(n15980));
  jor  g15725(.dina(n5534), .dinb(n5253), .dout(n15981));
  jand g15726(.dina(n15981), .dinb(n15980), .dout(n15982));
  jand g15727(.dina(n15982), .dinb(n15979), .dout(n15983));
  jand g15728(.dina(n15983), .dinb(n15978), .dout(n15984));
  jxor g15729(.dina(n15984), .dinb(n5111), .dout(n15985));
  jxor g15730(.dina(n15985), .dinb(n15977), .dout(n15986));
  jxor g15731(.dina(n15986), .dinb(n15894), .dout(n15987));
  jor  g15732(.dina(n6137), .dinb(n4902), .dout(n15988));
  jor  g15733(.dina(n4696), .dinb(n5685), .dout(n15989));
  jor  g15734(.dina(n4904), .dinb(n5911), .dout(n15990));
  jor  g15735(.dina(n4899), .dinb(n6139), .dout(n15991));
  jand g15736(.dina(n15991), .dinb(n15990), .dout(n15992));
  jand g15737(.dina(n15992), .dinb(n15989), .dout(n15993));
  jand g15738(.dina(n15993), .dinb(n15988), .dout(n15994));
  jxor g15739(.dina(n15994), .dinb(n4505), .dout(n15995));
  jxor g15740(.dina(n15995), .dinb(n15987), .dout(n15996));
  jxor g15741(.dina(n15996), .dinb(n15891), .dout(n15997));
  jor  g15742(.dina(n6844), .dinb(n4305), .dout(n15998));
  jor  g15743(.dina(n4116), .dinb(n6366), .dout(n15999));
  jor  g15744(.dina(n4303), .dinb(n6846), .dout(n16000));
  jor  g15745(.dina(n4308), .dinb(n6605), .dout(n16001));
  jand g15746(.dina(n16001), .dinb(n16000), .dout(n16002));
  jand g15747(.dina(n16002), .dinb(n15999), .dout(n16003));
  jand g15748(.dina(n16003), .dinb(n15998), .dout(n16004));
  jxor g15749(.dina(n16004), .dinb(n3938), .dout(n16005));
  jxor g15750(.dina(n16005), .dinb(n15997), .dout(n16006));
  jxor g15751(.dina(n16006), .dinb(n15888), .dout(n16007));
  jor  g15752(.dina(n7588), .dinb(n3751), .dout(n16008));
  jor  g15753(.dina(n3574), .dinb(n7086), .dout(n16009));
  jor  g15754(.dina(n3749), .dinb(n7590), .dout(n16010));
  jor  g15755(.dina(n3754), .dinb(n7338), .dout(n16011));
  jand g15756(.dina(n16011), .dinb(n16010), .dout(n16012));
  jand g15757(.dina(n16012), .dinb(n16009), .dout(n16013));
  jand g15758(.dina(n16013), .dinb(n16008), .dout(n16014));
  jxor g15759(.dina(n16014), .dinb(n3410), .dout(n16015));
  jxor g15760(.dina(n16015), .dinb(n16007), .dout(n16016));
  jxor g15761(.dina(n16016), .dinb(n15885), .dout(n16017));
  jand g15762(.dina(n15833), .dinb(n15826), .dout(n16018));
  jand g15763(.dina(n15834), .dinb(n15818), .dout(n16019));
  jor  g15764(.dina(n16019), .dinb(n16018), .dout(n16020));
  jor  g15765(.dina(n9193), .dinb(n2764), .dout(n16021));
  jor  g15766(.dina(n2609), .dinb(n8644), .dout(n16022));
  jor  g15767(.dina(n2761), .dinb(n9195), .dout(n16023));
  jor  g15768(.dina(n2766), .dinb(n8920), .dout(n16024));
  jand g15769(.dina(n16024), .dinb(n16023), .dout(n16025));
  jand g15770(.dina(n16025), .dinb(n16022), .dout(n16026));
  jand g15771(.dina(n16026), .dinb(n16021), .dout(n16027));
  jxor g15772(.dina(n16027), .dinb(n2468), .dout(n16028));
  jxor g15773(.dina(n16028), .dinb(n16020), .dout(n16029));
  jxor g15774(.dina(n16029), .dinb(n16017), .dout(n16030));
  jxor g15775(.dina(n16030), .dinb(n15873), .dout(n16031));
  jxor g15776(.dina(n16031), .dinb(n15861), .dout(n16032));
  jxor g15777(.dina(n16032), .dinb(n15852), .dout(n16033));
  jnot g15778(.din(n16033), .dout(n16034));
  jxor g15779(.dina(n16034), .dinb(n15849), .dout(f86 ));
  jand g15780(.dina(n16032), .dinb(n15852), .dout(n16036));
  jnot g15781(.din(n16036), .dout(n16037));
  jor  g15782(.dina(n16034), .dinb(n15849), .dout(n16038));
  jand g15783(.dina(n16038), .dinb(n16037), .dout(n16039));
  jor  g15784(.dina(n15860), .dinb(n15856), .dout(n16040));
  jand g15785(.dina(n16031), .dinb(n15861), .dout(n16041));
  jnot g15786(.din(n16041), .dout(n16042));
  jand g15787(.dina(n16042), .dinb(n16040), .dout(n16043));
  jnot g15788(.din(n16043), .dout(n16044));
  jand g15789(.dina(n15872), .dinb(n15864), .dout(n16045));
  jand g15790(.dina(n16030), .dinb(n15873), .dout(n16046));
  jor  g15791(.dina(n16046), .dinb(n16045), .dout(n16047));
  jor  g15792(.dina(n10521), .dinb(n2324), .dout(n16048));
  jor  g15793(.dina(n2186), .dinb(n9759), .dout(n16049));
  jor  g15794(.dina(n2321), .dinb(n10051), .dout(n16050));
  jor  g15795(.dina(n2326), .dinb(n10523), .dout(n16051));
  jand g15796(.dina(n16051), .dinb(n16050), .dout(n16052));
  jand g15797(.dina(n16052), .dinb(n16049), .dout(n16053));
  jand g15798(.dina(n16053), .dinb(n16048), .dout(n16054));
  jxor g15799(.dina(n16054), .dinb(n2057), .dout(n16055));
  jxor g15800(.dina(n16055), .dinb(n16047), .dout(n16056));
  jand g15801(.dina(n16028), .dinb(n16020), .dout(n16057));
  jand g15802(.dina(n16029), .dinb(n16017), .dout(n16058));
  jor  g15803(.dina(n16058), .dinb(n16057), .dout(n16059));
  jor  g15804(.dina(n9473), .dinb(n2764), .dout(n16060));
  jor  g15805(.dina(n2609), .dinb(n8920), .dout(n16061));
  jor  g15806(.dina(n2761), .dinb(n9475), .dout(n16062));
  jor  g15807(.dina(n2766), .dinb(n9195), .dout(n16063));
  jand g15808(.dina(n16063), .dinb(n16062), .dout(n16064));
  jand g15809(.dina(n16064), .dinb(n16061), .dout(n16065));
  jand g15810(.dina(n16065), .dinb(n16060), .dout(n16066));
  jxor g15811(.dina(n16066), .dinb(n2468), .dout(n16067));
  jxor g15812(.dina(n16067), .dinb(n16059), .dout(n16068));
  jand g15813(.dina(n15884), .dinb(n15876), .dout(n16069));
  jand g15814(.dina(n16016), .dinb(n15885), .dout(n16070));
  jor  g15815(.dina(n16070), .dinb(n16069), .dout(n16071));
  jor  g15816(.dina(n8642), .dinb(n3239), .dout(n16072));
  jor  g15817(.dina(n3072), .dinb(n8111), .dout(n16073));
  jor  g15818(.dina(n3237), .dinb(n8644), .dout(n16074));
  jor  g15819(.dina(n3242), .dinb(n8378), .dout(n16075));
  jand g15820(.dina(n16075), .dinb(n16074), .dout(n16076));
  jand g15821(.dina(n16076), .dinb(n16073), .dout(n16077));
  jand g15822(.dina(n16077), .dinb(n16072), .dout(n16078));
  jxor g15823(.dina(n16078), .dinb(n2918), .dout(n16079));
  jxor g15824(.dina(n16079), .dinb(n16071), .dout(n16080));
  jand g15825(.dina(n16006), .dinb(n15888), .dout(n16081));
  jand g15826(.dina(n16015), .dinb(n16007), .dout(n16082));
  jor  g15827(.dina(n16082), .dinb(n16081), .dout(n16083));
  jand g15828(.dina(n15996), .dinb(n15891), .dout(n16084));
  jand g15829(.dina(n16005), .dinb(n15997), .dout(n16085));
  jor  g15830(.dina(n16085), .dinb(n16084), .dout(n16086));
  jand g15831(.dina(n15986), .dinb(n15894), .dout(n16087));
  jand g15832(.dina(n15995), .dinb(n15987), .dout(n16088));
  jor  g15833(.dina(n16088), .dinb(n16087), .dout(n16089));
  jand g15834(.dina(n15976), .dinb(n15897), .dout(n16090));
  jand g15835(.dina(n15985), .dinb(n15977), .dout(n16091));
  jor  g15836(.dina(n16091), .dinb(n16090), .dout(n16092));
  jand g15837(.dina(n15966), .dinb(n15900), .dout(n16093));
  jand g15838(.dina(n15975), .dinb(n15967), .dout(n16094));
  jor  g15839(.dina(n16094), .dinb(n16093), .dout(n16095));
  jand g15840(.dina(n15956), .dinb(n15903), .dout(n16096));
  jand g15841(.dina(n15965), .dinb(n15957), .dout(n16097));
  jor  g15842(.dina(n16097), .dinb(n16096), .dout(n16098));
  jand g15843(.dina(n15946), .dinb(n15906), .dout(n16099));
  jand g15844(.dina(n15955), .dinb(n15947), .dout(n16100));
  jor  g15845(.dina(n16100), .dinb(n16099), .dout(n16101));
  jand g15846(.dina(n15926), .dinb(n15912), .dout(n16102));
  jand g15847(.dina(n15935), .dinb(n15927), .dout(n16103));
  jor  g15848(.dina(n16103), .dinb(n16102), .dout(n16104));
  jand g15849(.dina(n15916), .dinb(n15714), .dout(n16105));
  jand g15850(.dina(n15925), .dinb(n15917), .dout(n16106));
  jor  g15851(.dina(n16106), .dinb(n16105), .dout(n16107));
  jand g15852(.dina(n10594), .dinb(b23 ), .dout(n16108));
  jand g15853(.dina(n10129), .dinb(b24 ), .dout(n16109));
  jor  g15854(.dina(n16109), .dinb(n16108), .dout(n16110));
  jxor g15855(.dina(n16110), .dinb(n1687), .dout(n16111));
  jxor g15856(.dina(n16111), .dinb(n15915), .dout(n16112));
  jor  g15857(.dina(n10134), .dinb(n2413), .dout(n16113));
  jor  g15858(.dina(n9849), .dinb(n2142), .dout(n16114));
  jor  g15859(.dina(n10137), .dinb(n2279), .dout(n16115));
  jor  g15860(.dina(n10132), .dinb(n2415), .dout(n16116));
  jand g15861(.dina(n16116), .dinb(n16115), .dout(n16117));
  jand g15862(.dina(n16117), .dinb(n16114), .dout(n16118));
  jand g15863(.dina(n16118), .dinb(n16113), .dout(n16119));
  jxor g15864(.dina(n16119), .dinb(n9559), .dout(n16120));
  jxor g15865(.dina(n16120), .dinb(n16112), .dout(n16121));
  jxor g15866(.dina(n16121), .dinb(n16107), .dout(n16122));
  jor  g15867(.dina(n9271), .dinb(n2860), .dout(n16123));
  jor  g15868(.dina(n9003), .dinb(n2563), .dout(n16124));
  jor  g15869(.dina(n9268), .dinb(n2862), .dout(n16125));
  jor  g15870(.dina(n9273), .dinb(n2713), .dout(n16126));
  jand g15871(.dina(n16126), .dinb(n16125), .dout(n16127));
  jand g15872(.dina(n16127), .dinb(n16124), .dout(n16128));
  jand g15873(.dina(n16128), .dinb(n16123), .dout(n16129));
  jxor g15874(.dina(n16129), .dinb(n8729), .dout(n16130));
  jxor g15875(.dina(n16130), .dinb(n16122), .dout(n16131));
  jxor g15876(.dina(n16131), .dinb(n16104), .dout(n16132));
  jand g15877(.dina(n15936), .dinb(n15909), .dout(n16133));
  jand g15878(.dina(n15945), .dinb(n15937), .dout(n16134));
  jor  g15879(.dina(n16134), .dinb(n16133), .dout(n16135));
  jor  g15880(.dina(n8457), .dinb(n3346), .dout(n16136));
  jor  g15881(.dina(n8185), .dinb(n3023), .dout(n16137));
  jor  g15882(.dina(n8459), .dinb(n3186), .dout(n16138));
  jor  g15883(.dina(n8454), .dinb(n3348), .dout(n16139));
  jand g15884(.dina(n16139), .dinb(n16138), .dout(n16140));
  jand g15885(.dina(n16140), .dinb(n16137), .dout(n16141));
  jand g15886(.dina(n16141), .dinb(n16136), .dout(n16142));
  jxor g15887(.dina(n16142), .dinb(n7929), .dout(n16143));
  jxor g15888(.dina(n16143), .dinb(n16135), .dout(n16144));
  jxor g15889(.dina(n16144), .dinb(n16132), .dout(n16145));
  jor  g15890(.dina(n7660), .dinb(n3871), .dout(n16146));
  jor  g15891(.dina(n7415), .dinb(n3522), .dout(n16147));
  jor  g15892(.dina(n7657), .dinb(n3698), .dout(n16148));
  jor  g15893(.dina(n7662), .dinb(n3873), .dout(n16149));
  jand g15894(.dina(n16149), .dinb(n16148), .dout(n16150));
  jand g15895(.dina(n16150), .dinb(n16147), .dout(n16151));
  jand g15896(.dina(n16151), .dinb(n16146), .dout(n16152));
  jxor g15897(.dina(n16152), .dinb(n7166), .dout(n16153));
  jxor g15898(.dina(n16153), .dinb(n16145), .dout(n16154));
  jxor g15899(.dina(n16154), .dinb(n16101), .dout(n16155));
  jor  g15900(.dina(n6914), .dinb(n4435), .dout(n16156));
  jor  g15901(.dina(n6673), .dinb(n4060), .dout(n16157));
  jor  g15902(.dina(n6911), .dinb(n4249), .dout(n16158));
  jor  g15903(.dina(n6916), .dinb(n4437), .dout(n16159));
  jand g15904(.dina(n16159), .dinb(n16158), .dout(n16160));
  jand g15905(.dina(n16160), .dinb(n16157), .dout(n16161));
  jand g15906(.dina(n16161), .dinb(n16156), .dout(n16162));
  jxor g15907(.dina(n16162), .dinb(n6443), .dout(n16163));
  jxor g15908(.dina(n16163), .dinb(n16155), .dout(n16164));
  jxor g15909(.dina(n16164), .dinb(n16098), .dout(n16165));
  jor  g15910(.dina(n6207), .dinb(n5038), .dout(n16166));
  jor  g15911(.dina(n5975), .dinb(n4637), .dout(n16167));
  jor  g15912(.dina(n6210), .dinb(n4839), .dout(n16168));
  jor  g15913(.dina(n6205), .dinb(n5040), .dout(n16169));
  jand g15914(.dina(n16169), .dinb(n16168), .dout(n16170));
  jand g15915(.dina(n16170), .dinb(n16167), .dout(n16171));
  jand g15916(.dina(n16171), .dinb(n16166), .dout(n16172));
  jxor g15917(.dina(n16172), .dinb(n5759), .dout(n16173));
  jxor g15918(.dina(n16173), .dinb(n16165), .dout(n16174));
  jxor g15919(.dina(n16174), .dinb(n16095), .dout(n16175));
  jor  g15920(.dina(n5683), .dinb(n5537), .dout(n16176));
  jor  g15921(.dina(n5315), .dinb(n5253), .dout(n16177));
  jor  g15922(.dina(n5539), .dinb(n5685), .dout(n16178));
  jor  g15923(.dina(n5534), .dinb(n5469), .dout(n16179));
  jand g15924(.dina(n16179), .dinb(n16178), .dout(n16180));
  jand g15925(.dina(n16180), .dinb(n16177), .dout(n16181));
  jand g15926(.dina(n16181), .dinb(n16176), .dout(n16182));
  jxor g15927(.dina(n16182), .dinb(n5111), .dout(n16183));
  jxor g15928(.dina(n16183), .dinb(n16175), .dout(n16184));
  jxor g15929(.dina(n16184), .dinb(n16092), .dout(n16185));
  jor  g15930(.dina(n6364), .dinb(n4902), .dout(n16186));
  jor  g15931(.dina(n4696), .dinb(n5911), .dout(n16187));
  jor  g15932(.dina(n4899), .dinb(n6366), .dout(n16188));
  jor  g15933(.dina(n4904), .dinb(n6139), .dout(n16189));
  jand g15934(.dina(n16189), .dinb(n16188), .dout(n16190));
  jand g15935(.dina(n16190), .dinb(n16187), .dout(n16191));
  jand g15936(.dina(n16191), .dinb(n16186), .dout(n16192));
  jxor g15937(.dina(n16192), .dinb(n4505), .dout(n16193));
  jxor g15938(.dina(n16193), .dinb(n16185), .dout(n16194));
  jxor g15939(.dina(n16194), .dinb(n16089), .dout(n16195));
  jor  g15940(.dina(n7084), .dinb(n4305), .dout(n16196));
  jor  g15941(.dina(n4116), .dinb(n6605), .dout(n16197));
  jor  g15942(.dina(n4308), .dinb(n6846), .dout(n16198));
  jor  g15943(.dina(n4303), .dinb(n7086), .dout(n16199));
  jand g15944(.dina(n16199), .dinb(n16198), .dout(n16200));
  jand g15945(.dina(n16200), .dinb(n16197), .dout(n16201));
  jand g15946(.dina(n16201), .dinb(n16196), .dout(n16202));
  jxor g15947(.dina(n16202), .dinb(n3938), .dout(n16203));
  jxor g15948(.dina(n16203), .dinb(n16195), .dout(n16204));
  jxor g15949(.dina(n16204), .dinb(n16086), .dout(n16205));
  jor  g15950(.dina(n7844), .dinb(n3751), .dout(n16206));
  jor  g15951(.dina(n3574), .dinb(n7338), .dout(n16207));
  jor  g15952(.dina(n3749), .dinb(n7846), .dout(n16208));
  jor  g15953(.dina(n3754), .dinb(n7590), .dout(n16209));
  jand g15954(.dina(n16209), .dinb(n16208), .dout(n16210));
  jand g15955(.dina(n16210), .dinb(n16207), .dout(n16211));
  jand g15956(.dina(n16211), .dinb(n16206), .dout(n16212));
  jxor g15957(.dina(n16212), .dinb(n3410), .dout(n16213));
  jxor g15958(.dina(n16213), .dinb(n16205), .dout(n16214));
  jxor g15959(.dina(n16214), .dinb(n16083), .dout(n16215));
  jxor g15960(.dina(n16215), .dinb(n16080), .dout(n16216));
  jxor g15961(.dina(n16216), .dinb(n16068), .dout(n16217));
  jxor g15962(.dina(n16217), .dinb(n16056), .dout(n16218));
  jxor g15963(.dina(n16218), .dinb(n16044), .dout(n16219));
  jnot g15964(.din(n16219), .dout(n16220));
  jxor g15965(.dina(n16220), .dinb(n16039), .dout(f87 ));
  jand g15966(.dina(n16218), .dinb(n16044), .dout(n16222));
  jnot g15967(.din(n16222), .dout(n16223));
  jor  g15968(.dina(n16220), .dinb(n16039), .dout(n16224));
  jand g15969(.dina(n16224), .dinb(n16223), .dout(n16225));
  jand g15970(.dina(n16055), .dinb(n16047), .dout(n16226));
  jand g15971(.dina(n16217), .dinb(n16056), .dout(n16227));
  jor  g15972(.dina(n16227), .dinb(n16226), .dout(n16228));
  jand g15973(.dina(n16213), .dinb(n16205), .dout(n16229));
  jand g15974(.dina(n16214), .dinb(n16083), .dout(n16230));
  jor  g15975(.dina(n16230), .dinb(n16229), .dout(n16231));
  jor  g15976(.dina(n8918), .dinb(n3239), .dout(n16232));
  jor  g15977(.dina(n3072), .dinb(n8378), .dout(n16233));
  jor  g15978(.dina(n3242), .dinb(n8644), .dout(n16234));
  jor  g15979(.dina(n3237), .dinb(n8920), .dout(n16235));
  jand g15980(.dina(n16235), .dinb(n16234), .dout(n16236));
  jand g15981(.dina(n16236), .dinb(n16233), .dout(n16237));
  jand g15982(.dina(n16237), .dinb(n16232), .dout(n16238));
  jxor g15983(.dina(n16238), .dinb(n2918), .dout(n16239));
  jxor g15984(.dina(n16239), .dinb(n16231), .dout(n16240));
  jand g15985(.dina(n16193), .dinb(n16185), .dout(n16241));
  jand g15986(.dina(n16194), .dinb(n16089), .dout(n16242));
  jor  g15987(.dina(n16242), .dinb(n16241), .dout(n16243));
  jand g15988(.dina(n16183), .dinb(n16175), .dout(n16244));
  jand g15989(.dina(n16184), .dinb(n16092), .dout(n16245));
  jor  g15990(.dina(n16245), .dinb(n16244), .dout(n16246));
  jand g15991(.dina(n16173), .dinb(n16165), .dout(n16247));
  jand g15992(.dina(n16174), .dinb(n16095), .dout(n16248));
  jor  g15993(.dina(n16248), .dinb(n16247), .dout(n16249));
  jand g15994(.dina(n16163), .dinb(n16155), .dout(n16250));
  jand g15995(.dina(n16164), .dinb(n16098), .dout(n16251));
  jor  g15996(.dina(n16251), .dinb(n16250), .dout(n16252));
  jand g15997(.dina(n16153), .dinb(n16145), .dout(n16253));
  jand g15998(.dina(n16154), .dinb(n16101), .dout(n16254));
  jor  g15999(.dina(n16254), .dinb(n16253), .dout(n16255));
  jand g16000(.dina(n16143), .dinb(n16135), .dout(n16256));
  jand g16001(.dina(n16144), .dinb(n16132), .dout(n16257));
  jor  g16002(.dina(n16257), .dinb(n16256), .dout(n16258));
  jand g16003(.dina(n16130), .dinb(n16122), .dout(n16259));
  jand g16004(.dina(n16131), .dinb(n16104), .dout(n16260));
  jor  g16005(.dina(n16260), .dinb(n16259), .dout(n16261));
  jand g16006(.dina(n16120), .dinb(n16112), .dout(n16262));
  jand g16007(.dina(n16121), .dinb(n16107), .dout(n16263));
  jor  g16008(.dina(n16263), .dinb(n16262), .dout(n16264));
  jand g16009(.dina(n10594), .dinb(b24 ), .dout(n16265));
  jand g16010(.dina(n10129), .dinb(b25 ), .dout(n16266));
  jor  g16011(.dina(n16266), .dinb(n16265), .dout(n16267));
  jnot g16012(.din(n16267), .dout(n16268));
  jand g16013(.dina(n16110), .dinb(n1687), .dout(n16269));
  jand g16014(.dina(n16111), .dinb(n15915), .dout(n16270));
  jor  g16015(.dina(n16270), .dinb(n16269), .dout(n16271));
  jxor g16016(.dina(n16271), .dinb(n16268), .dout(n16272));
  jor  g16017(.dina(n10134), .dinb(n2561), .dout(n16273));
  jor  g16018(.dina(n9849), .dinb(n2279), .dout(n16274));
  jor  g16019(.dina(n10137), .dinb(n2415), .dout(n16275));
  jor  g16020(.dina(n10132), .dinb(n2563), .dout(n16276));
  jand g16021(.dina(n16276), .dinb(n16275), .dout(n16277));
  jand g16022(.dina(n16277), .dinb(n16274), .dout(n16278));
  jand g16023(.dina(n16278), .dinb(n16273), .dout(n16279));
  jxor g16024(.dina(n16279), .dinb(n9559), .dout(n16280));
  jxor g16025(.dina(n16280), .dinb(n16272), .dout(n16281));
  jxor g16026(.dina(n16281), .dinb(n16264), .dout(n16282));
  jor  g16027(.dina(n9271), .dinb(n3021), .dout(n16283));
  jor  g16028(.dina(n9003), .dinb(n2713), .dout(n16284));
  jor  g16029(.dina(n9273), .dinb(n2862), .dout(n16285));
  jor  g16030(.dina(n9268), .dinb(n3023), .dout(n16286));
  jand g16031(.dina(n16286), .dinb(n16285), .dout(n16287));
  jand g16032(.dina(n16287), .dinb(n16284), .dout(n16288));
  jand g16033(.dina(n16288), .dinb(n16283), .dout(n16289));
  jxor g16034(.dina(n16289), .dinb(n8729), .dout(n16290));
  jxor g16035(.dina(n16290), .dinb(n16282), .dout(n16291));
  jxor g16036(.dina(n16291), .dinb(n16261), .dout(n16292));
  jor  g16037(.dina(n8457), .dinb(n3520), .dout(n16293));
  jor  g16038(.dina(n8185), .dinb(n3186), .dout(n16294));
  jor  g16039(.dina(n8454), .dinb(n3522), .dout(n16295));
  jor  g16040(.dina(n8459), .dinb(n3348), .dout(n16296));
  jand g16041(.dina(n16296), .dinb(n16295), .dout(n16297));
  jand g16042(.dina(n16297), .dinb(n16294), .dout(n16298));
  jand g16043(.dina(n16298), .dinb(n16293), .dout(n16299));
  jxor g16044(.dina(n16299), .dinb(n7929), .dout(n16300));
  jxor g16045(.dina(n16300), .dinb(n16292), .dout(n16301));
  jxor g16046(.dina(n16301), .dinb(n16258), .dout(n16302));
  jor  g16047(.dina(n7660), .dinb(n4058), .dout(n16303));
  jor  g16048(.dina(n7415), .dinb(n3698), .dout(n16304));
  jor  g16049(.dina(n7662), .dinb(n4060), .dout(n16305));
  jor  g16050(.dina(n7657), .dinb(n3873), .dout(n16306));
  jand g16051(.dina(n16306), .dinb(n16305), .dout(n16307));
  jand g16052(.dina(n16307), .dinb(n16304), .dout(n16308));
  jand g16053(.dina(n16308), .dinb(n16303), .dout(n16309));
  jxor g16054(.dina(n16309), .dinb(n7166), .dout(n16310));
  jxor g16055(.dina(n16310), .dinb(n16302), .dout(n16311));
  jxor g16056(.dina(n16311), .dinb(n16255), .dout(n16312));
  jor  g16057(.dina(n6914), .dinb(n4635), .dout(n16313));
  jor  g16058(.dina(n6673), .dinb(n4249), .dout(n16314));
  jor  g16059(.dina(n6911), .dinb(n4437), .dout(n16315));
  jor  g16060(.dina(n6916), .dinb(n4637), .dout(n16316));
  jand g16061(.dina(n16316), .dinb(n16315), .dout(n16317));
  jand g16062(.dina(n16317), .dinb(n16314), .dout(n16318));
  jand g16063(.dina(n16318), .dinb(n16313), .dout(n16319));
  jxor g16064(.dina(n16319), .dinb(n6443), .dout(n16320));
  jxor g16065(.dina(n16320), .dinb(n16312), .dout(n16321));
  jxor g16066(.dina(n16321), .dinb(n16252), .dout(n16322));
  jor  g16067(.dina(n6207), .dinb(n5251), .dout(n16323));
  jor  g16068(.dina(n5975), .dinb(n4839), .dout(n16324));
  jor  g16069(.dina(n6205), .dinb(n5253), .dout(n16325));
  jor  g16070(.dina(n6210), .dinb(n5040), .dout(n16326));
  jand g16071(.dina(n16326), .dinb(n16325), .dout(n16327));
  jand g16072(.dina(n16327), .dinb(n16324), .dout(n16328));
  jand g16073(.dina(n16328), .dinb(n16323), .dout(n16329));
  jxor g16074(.dina(n16329), .dinb(n5759), .dout(n16330));
  jxor g16075(.dina(n16330), .dinb(n16322), .dout(n16331));
  jxor g16076(.dina(n16331), .dinb(n16249), .dout(n16332));
  jor  g16077(.dina(n5909), .dinb(n5537), .dout(n16333));
  jor  g16078(.dina(n5315), .dinb(n5469), .dout(n16334));
  jor  g16079(.dina(n5539), .dinb(n5911), .dout(n16335));
  jor  g16080(.dina(n5534), .dinb(n5685), .dout(n16336));
  jand g16081(.dina(n16336), .dinb(n16335), .dout(n16337));
  jand g16082(.dina(n16337), .dinb(n16334), .dout(n16338));
  jand g16083(.dina(n16338), .dinb(n16333), .dout(n16339));
  jxor g16084(.dina(n16339), .dinb(n5111), .dout(n16340));
  jxor g16085(.dina(n16340), .dinb(n16332), .dout(n16341));
  jxor g16086(.dina(n16341), .dinb(n16246), .dout(n16342));
  jor  g16087(.dina(n6603), .dinb(n4902), .dout(n16343));
  jor  g16088(.dina(n4696), .dinb(n6139), .dout(n16344));
  jor  g16089(.dina(n4899), .dinb(n6605), .dout(n16345));
  jor  g16090(.dina(n4904), .dinb(n6366), .dout(n16346));
  jand g16091(.dina(n16346), .dinb(n16345), .dout(n16347));
  jand g16092(.dina(n16347), .dinb(n16344), .dout(n16348));
  jand g16093(.dina(n16348), .dinb(n16343), .dout(n16349));
  jxor g16094(.dina(n16349), .dinb(n4505), .dout(n16350));
  jxor g16095(.dina(n16350), .dinb(n16342), .dout(n16351));
  jxor g16096(.dina(n16351), .dinb(n16243), .dout(n16352));
  jor  g16097(.dina(n7336), .dinb(n4305), .dout(n16353));
  jor  g16098(.dina(n4116), .dinb(n6846), .dout(n16354));
  jor  g16099(.dina(n4308), .dinb(n7086), .dout(n16355));
  jor  g16100(.dina(n4303), .dinb(n7338), .dout(n16356));
  jand g16101(.dina(n16356), .dinb(n16355), .dout(n16357));
  jand g16102(.dina(n16357), .dinb(n16354), .dout(n16358));
  jand g16103(.dina(n16358), .dinb(n16353), .dout(n16359));
  jxor g16104(.dina(n16359), .dinb(n3938), .dout(n16360));
  jxor g16105(.dina(n16360), .dinb(n16352), .dout(n16361));
  jnot g16106(.din(n16195), .dout(n16362));
  jnot g16107(.din(n16203), .dout(n16363));
  jand g16108(.dina(n16363), .dinb(n16362), .dout(n16364));
  jnot g16109(.din(n16364), .dout(n16365));
  jand g16110(.dina(n16203), .dinb(n16195), .dout(n16366));
  jor  g16111(.dina(n16366), .dinb(n16086), .dout(n16367));
  jand g16112(.dina(n16367), .dinb(n16365), .dout(n16368));
  jxor g16113(.dina(n16368), .dinb(n16361), .dout(n16369));
  jor  g16114(.dina(n8109), .dinb(n3751), .dout(n16370));
  jor  g16115(.dina(n3574), .dinb(n7590), .dout(n16371));
  jor  g16116(.dina(n3754), .dinb(n7846), .dout(n16372));
  jor  g16117(.dina(n3749), .dinb(n8111), .dout(n16373));
  jand g16118(.dina(n16373), .dinb(n16372), .dout(n16374));
  jand g16119(.dina(n16374), .dinb(n16371), .dout(n16375));
  jand g16120(.dina(n16375), .dinb(n16370), .dout(n16376));
  jxor g16121(.dina(n16376), .dinb(n3410), .dout(n16377));
  jxor g16122(.dina(n16377), .dinb(n16369), .dout(n16378));
  jxor g16123(.dina(n16378), .dinb(n16240), .dout(n16379));
  jand g16124(.dina(n16079), .dinb(n16071), .dout(n16380));
  jand g16125(.dina(n16215), .dinb(n16080), .dout(n16381));
  jor  g16126(.dina(n16381), .dinb(n16380), .dout(n16382));
  jor  g16127(.dina(n9757), .dinb(n2764), .dout(n16383));
  jor  g16128(.dina(n2609), .dinb(n9195), .dout(n16384));
  jor  g16129(.dina(n2761), .dinb(n9759), .dout(n16385));
  jor  g16130(.dina(n2766), .dinb(n9475), .dout(n16386));
  jand g16131(.dina(n16386), .dinb(n16385), .dout(n16387));
  jand g16132(.dina(n16387), .dinb(n16384), .dout(n16388));
  jand g16133(.dina(n16388), .dinb(n16383), .dout(n16389));
  jxor g16134(.dina(n16389), .dinb(n2468), .dout(n16390));
  jxor g16135(.dina(n16390), .dinb(n16382), .dout(n16391));
  jxor g16136(.dina(n16391), .dinb(n16379), .dout(n16392));
  jand g16137(.dina(n16067), .dinb(n16059), .dout(n16393));
  jand g16138(.dina(n16216), .dinb(n16068), .dout(n16394));
  jor  g16139(.dina(n16394), .dinb(n16393), .dout(n16395));
  jnot g16140(.din(n16395), .dout(n16396));
  jor  g16141(.dina(n10813), .dinb(n2324), .dout(n16397));
  jor  g16142(.dina(n2186), .dinb(n10051), .dout(n16398));
  jor  g16143(.dina(n2321), .dinb(n10523), .dout(n16399));
  jand g16144(.dina(n16399), .dinb(n16398), .dout(n16400));
  jand g16145(.dina(n16400), .dinb(n16397), .dout(n16401));
  jxor g16146(.dina(n16401), .dinb(a26 ), .dout(n16402));
  jxor g16147(.dina(n16402), .dinb(n16396), .dout(n16403));
  jxor g16148(.dina(n16403), .dinb(n16392), .dout(n16404));
  jxor g16149(.dina(n16404), .dinb(n16228), .dout(n16405));
  jnot g16150(.din(n16405), .dout(n16406));
  jxor g16151(.dina(n16406), .dinb(n16225), .dout(f88 ));
  jand g16152(.dina(n16404), .dinb(n16228), .dout(n16408));
  jnot g16153(.din(n16408), .dout(n16409));
  jor  g16154(.dina(n16406), .dinb(n16225), .dout(n16410));
  jand g16155(.dina(n16410), .dinb(n16409), .dout(n16411));
  jor  g16156(.dina(n16402), .dinb(n16396), .dout(n16412));
  jand g16157(.dina(n16403), .dinb(n16392), .dout(n16413));
  jnot g16158(.din(n16413), .dout(n16414));
  jand g16159(.dina(n16414), .dinb(n16412), .dout(n16415));
  jnot g16160(.din(n16415), .dout(n16416));
  jand g16161(.dina(n16239), .dinb(n16231), .dout(n16417));
  jand g16162(.dina(n16378), .dinb(n16240), .dout(n16418));
  jor  g16163(.dina(n16418), .dinb(n16417), .dout(n16419));
  jor  g16164(.dina(n10049), .dinb(n2764), .dout(n16420));
  jor  g16165(.dina(n2609), .dinb(n9475), .dout(n16421));
  jor  g16166(.dina(n2761), .dinb(n10051), .dout(n16422));
  jor  g16167(.dina(n2766), .dinb(n9759), .dout(n16423));
  jand g16168(.dina(n16423), .dinb(n16422), .dout(n16424));
  jand g16169(.dina(n16424), .dinb(n16421), .dout(n16425));
  jand g16170(.dina(n16425), .dinb(n16420), .dout(n16426));
  jxor g16171(.dina(n16426), .dinb(n2468), .dout(n16427));
  jxor g16172(.dina(n16427), .dinb(n16419), .dout(n16428));
  jand g16173(.dina(n16368), .dinb(n16361), .dout(n16429));
  jand g16174(.dina(n16377), .dinb(n16369), .dout(n16430));
  jor  g16175(.dina(n16430), .dinb(n16429), .dout(n16431));
  jor  g16176(.dina(n9193), .dinb(n3239), .dout(n16432));
  jor  g16177(.dina(n3072), .dinb(n8644), .dout(n16433));
  jor  g16178(.dina(n3242), .dinb(n8920), .dout(n16434));
  jor  g16179(.dina(n3237), .dinb(n9195), .dout(n16435));
  jand g16180(.dina(n16435), .dinb(n16434), .dout(n16436));
  jand g16181(.dina(n16436), .dinb(n16433), .dout(n16437));
  jand g16182(.dina(n16437), .dinb(n16432), .dout(n16438));
  jxor g16183(.dina(n16438), .dinb(n2918), .dout(n16439));
  jxor g16184(.dina(n16439), .dinb(n16431), .dout(n16440));
  jand g16185(.dina(n16351), .dinb(n16243), .dout(n16441));
  jand g16186(.dina(n16360), .dinb(n16352), .dout(n16442));
  jor  g16187(.dina(n16442), .dinb(n16441), .dout(n16443));
  jand g16188(.dina(n16341), .dinb(n16246), .dout(n16444));
  jand g16189(.dina(n16350), .dinb(n16342), .dout(n16445));
  jor  g16190(.dina(n16445), .dinb(n16444), .dout(n16446));
  jand g16191(.dina(n16331), .dinb(n16249), .dout(n16447));
  jand g16192(.dina(n16340), .dinb(n16332), .dout(n16448));
  jor  g16193(.dina(n16448), .dinb(n16447), .dout(n16449));
  jand g16194(.dina(n16321), .dinb(n16252), .dout(n16450));
  jand g16195(.dina(n16330), .dinb(n16322), .dout(n16451));
  jor  g16196(.dina(n16451), .dinb(n16450), .dout(n16452));
  jand g16197(.dina(n16311), .dinb(n16255), .dout(n16453));
  jand g16198(.dina(n16320), .dinb(n16312), .dout(n16454));
  jor  g16199(.dina(n16454), .dinb(n16453), .dout(n16455));
  jand g16200(.dina(n16301), .dinb(n16258), .dout(n16456));
  jand g16201(.dina(n16310), .dinb(n16302), .dout(n16457));
  jor  g16202(.dina(n16457), .dinb(n16456), .dout(n16458));
  jand g16203(.dina(n16291), .dinb(n16261), .dout(n16459));
  jand g16204(.dina(n16300), .dinb(n16292), .dout(n16460));
  jor  g16205(.dina(n16460), .dinb(n16459), .dout(n16461));
  jand g16206(.dina(n16281), .dinb(n16264), .dout(n16462));
  jand g16207(.dina(n16290), .dinb(n16282), .dout(n16463));
  jor  g16208(.dina(n16463), .dinb(n16462), .dout(n16464));
  jand g16209(.dina(n16271), .dinb(n16268), .dout(n16465));
  jand g16210(.dina(n16280), .dinb(n16272), .dout(n16466));
  jor  g16211(.dina(n16466), .dinb(n16465), .dout(n16467));
  jand g16212(.dina(n10594), .dinb(b25 ), .dout(n16468));
  jand g16213(.dina(n10129), .dinb(b26 ), .dout(n16469));
  jor  g16214(.dina(n16469), .dinb(n16468), .dout(n16470));
  jnot g16215(.din(n16470), .dout(n16471));
  jxor g16216(.dina(n16471), .dinb(n16267), .dout(n16472));
  jor  g16217(.dina(n10134), .dinb(n2711), .dout(n16473));
  jor  g16218(.dina(n9849), .dinb(n2415), .dout(n16474));
  jor  g16219(.dina(n10137), .dinb(n2563), .dout(n16475));
  jor  g16220(.dina(n10132), .dinb(n2713), .dout(n16476));
  jand g16221(.dina(n16476), .dinb(n16475), .dout(n16477));
  jand g16222(.dina(n16477), .dinb(n16474), .dout(n16478));
  jand g16223(.dina(n16478), .dinb(n16473), .dout(n16479));
  jxor g16224(.dina(n16479), .dinb(n9559), .dout(n16480));
  jxor g16225(.dina(n16480), .dinb(n16472), .dout(n16481));
  jxor g16226(.dina(n16481), .dinb(n16467), .dout(n16482));
  jor  g16227(.dina(n9271), .dinb(n3184), .dout(n16483));
  jor  g16228(.dina(n9003), .dinb(n2862), .dout(n16484));
  jor  g16229(.dina(n9273), .dinb(n3023), .dout(n16485));
  jor  g16230(.dina(n9268), .dinb(n3186), .dout(n16486));
  jand g16231(.dina(n16486), .dinb(n16485), .dout(n16487));
  jand g16232(.dina(n16487), .dinb(n16484), .dout(n16488));
  jand g16233(.dina(n16488), .dinb(n16483), .dout(n16489));
  jxor g16234(.dina(n16489), .dinb(n8729), .dout(n16490));
  jxor g16235(.dina(n16490), .dinb(n16482), .dout(n16491));
  jxor g16236(.dina(n16491), .dinb(n16464), .dout(n16492));
  jor  g16237(.dina(n8457), .dinb(n3696), .dout(n16493));
  jor  g16238(.dina(n8185), .dinb(n3348), .dout(n16494));
  jor  g16239(.dina(n8454), .dinb(n3698), .dout(n16495));
  jor  g16240(.dina(n8459), .dinb(n3522), .dout(n16496));
  jand g16241(.dina(n16496), .dinb(n16495), .dout(n16497));
  jand g16242(.dina(n16497), .dinb(n16494), .dout(n16498));
  jand g16243(.dina(n16498), .dinb(n16493), .dout(n16499));
  jxor g16244(.dina(n16499), .dinb(n7929), .dout(n16500));
  jxor g16245(.dina(n16500), .dinb(n16492), .dout(n16501));
  jxor g16246(.dina(n16501), .dinb(n16461), .dout(n16502));
  jor  g16247(.dina(n7660), .dinb(n4247), .dout(n16503));
  jor  g16248(.dina(n7415), .dinb(n3873), .dout(n16504));
  jor  g16249(.dina(n7657), .dinb(n4060), .dout(n16505));
  jor  g16250(.dina(n7662), .dinb(n4249), .dout(n16506));
  jand g16251(.dina(n16506), .dinb(n16505), .dout(n16507));
  jand g16252(.dina(n16507), .dinb(n16504), .dout(n16508));
  jand g16253(.dina(n16508), .dinb(n16503), .dout(n16509));
  jxor g16254(.dina(n16509), .dinb(n7166), .dout(n16510));
  jxor g16255(.dina(n16510), .dinb(n16502), .dout(n16511));
  jxor g16256(.dina(n16511), .dinb(n16458), .dout(n16512));
  jor  g16257(.dina(n6914), .dinb(n4837), .dout(n16513));
  jor  g16258(.dina(n6673), .dinb(n4437), .dout(n16514));
  jor  g16259(.dina(n6911), .dinb(n4637), .dout(n16515));
  jor  g16260(.dina(n6916), .dinb(n4839), .dout(n16516));
  jand g16261(.dina(n16516), .dinb(n16515), .dout(n16517));
  jand g16262(.dina(n16517), .dinb(n16514), .dout(n16518));
  jand g16263(.dina(n16518), .dinb(n16513), .dout(n16519));
  jxor g16264(.dina(n16519), .dinb(n6443), .dout(n16520));
  jxor g16265(.dina(n16520), .dinb(n16512), .dout(n16521));
  jxor g16266(.dina(n16521), .dinb(n16455), .dout(n16522));
  jor  g16267(.dina(n6207), .dinb(n5467), .dout(n16523));
  jor  g16268(.dina(n5975), .dinb(n5040), .dout(n16524));
  jor  g16269(.dina(n6210), .dinb(n5253), .dout(n16525));
  jor  g16270(.dina(n6205), .dinb(n5469), .dout(n16526));
  jand g16271(.dina(n16526), .dinb(n16525), .dout(n16527));
  jand g16272(.dina(n16527), .dinb(n16524), .dout(n16528));
  jand g16273(.dina(n16528), .dinb(n16523), .dout(n16529));
  jxor g16274(.dina(n16529), .dinb(n5759), .dout(n16530));
  jxor g16275(.dina(n16530), .dinb(n16522), .dout(n16531));
  jxor g16276(.dina(n16531), .dinb(n16452), .dout(n16532));
  jor  g16277(.dina(n6137), .dinb(n5537), .dout(n16533));
  jor  g16278(.dina(n5315), .dinb(n5685), .dout(n16534));
  jor  g16279(.dina(n5534), .dinb(n5911), .dout(n16535));
  jor  g16280(.dina(n5539), .dinb(n6139), .dout(n16536));
  jand g16281(.dina(n16536), .dinb(n16535), .dout(n16537));
  jand g16282(.dina(n16537), .dinb(n16534), .dout(n16538));
  jand g16283(.dina(n16538), .dinb(n16533), .dout(n16539));
  jxor g16284(.dina(n16539), .dinb(n5111), .dout(n16540));
  jxor g16285(.dina(n16540), .dinb(n16532), .dout(n16541));
  jxor g16286(.dina(n16541), .dinb(n16449), .dout(n16542));
  jor  g16287(.dina(n6844), .dinb(n4902), .dout(n16543));
  jor  g16288(.dina(n4696), .dinb(n6366), .dout(n16544));
  jor  g16289(.dina(n4899), .dinb(n6846), .dout(n16545));
  jor  g16290(.dina(n4904), .dinb(n6605), .dout(n16546));
  jand g16291(.dina(n16546), .dinb(n16545), .dout(n16547));
  jand g16292(.dina(n16547), .dinb(n16544), .dout(n16548));
  jand g16293(.dina(n16548), .dinb(n16543), .dout(n16549));
  jxor g16294(.dina(n16549), .dinb(n4505), .dout(n16550));
  jxor g16295(.dina(n16550), .dinb(n16542), .dout(n16551));
  jxor g16296(.dina(n16551), .dinb(n16446), .dout(n16552));
  jor  g16297(.dina(n7588), .dinb(n4305), .dout(n16553));
  jor  g16298(.dina(n4116), .dinb(n7086), .dout(n16554));
  jor  g16299(.dina(n4308), .dinb(n7338), .dout(n16555));
  jor  g16300(.dina(n4303), .dinb(n7590), .dout(n16556));
  jand g16301(.dina(n16556), .dinb(n16555), .dout(n16557));
  jand g16302(.dina(n16557), .dinb(n16554), .dout(n16558));
  jand g16303(.dina(n16558), .dinb(n16553), .dout(n16559));
  jxor g16304(.dina(n16559), .dinb(n3938), .dout(n16560));
  jxor g16305(.dina(n16560), .dinb(n16552), .dout(n16561));
  jxor g16306(.dina(n16561), .dinb(n16443), .dout(n16562));
  jor  g16307(.dina(n8376), .dinb(n3751), .dout(n16563));
  jor  g16308(.dina(n3574), .dinb(n7846), .dout(n16564));
  jor  g16309(.dina(n3754), .dinb(n8111), .dout(n16565));
  jor  g16310(.dina(n3749), .dinb(n8378), .dout(n16566));
  jand g16311(.dina(n16566), .dinb(n16565), .dout(n16567));
  jand g16312(.dina(n16567), .dinb(n16564), .dout(n16568));
  jand g16313(.dina(n16568), .dinb(n16563), .dout(n16569));
  jxor g16314(.dina(n16569), .dinb(n3410), .dout(n16570));
  jxor g16315(.dina(n16570), .dinb(n16562), .dout(n16571));
  jxor g16316(.dina(n16571), .dinb(n16440), .dout(n16572));
  jxor g16317(.dina(n16572), .dinb(n16428), .dout(n16573));
  jand g16318(.dina(n16390), .dinb(n16382), .dout(n16574));
  jand g16319(.dina(n16391), .dinb(n16379), .dout(n16575));
  jor  g16320(.dina(n16575), .dinb(n16574), .dout(n16576));
  jnot g16321(.din(n16576), .dout(n16577));
  jand g16322(.dina(n2187), .dinb(b63 ), .dout(n16578));
  jand g16323(.dina(n10832), .dinb(n2049), .dout(n16579));
  jor  g16324(.dina(n16579), .dinb(n16578), .dout(n16580));
  jxor g16325(.dina(n16580), .dinb(n2057), .dout(n16581));
  jxor g16326(.dina(n16581), .dinb(n16577), .dout(n16582));
  jxor g16327(.dina(n16582), .dinb(n16573), .dout(n16583));
  jxor g16328(.dina(n16583), .dinb(n16416), .dout(n16584));
  jnot g16329(.din(n16584), .dout(n16585));
  jxor g16330(.dina(n16585), .dinb(n16411), .dout(f89 ));
  jor  g16331(.dina(n16581), .dinb(n16577), .dout(n16587));
  jand g16332(.dina(n16582), .dinb(n16573), .dout(n16588));
  jnot g16333(.din(n16588), .dout(n16589));
  jand g16334(.dina(n16589), .dinb(n16587), .dout(n16590));
  jnot g16335(.din(n16590), .dout(n16591));
  jand g16336(.dina(n16427), .dinb(n16419), .dout(n16592));
  jand g16337(.dina(n16572), .dinb(n16428), .dout(n16593));
  jor  g16338(.dina(n16593), .dinb(n16592), .dout(n16594));
  jor  g16339(.dina(n10521), .dinb(n2764), .dout(n16595));
  jor  g16340(.dina(n2609), .dinb(n9759), .dout(n16596));
  jor  g16341(.dina(n2761), .dinb(n10523), .dout(n16597));
  jor  g16342(.dina(n2766), .dinb(n10051), .dout(n16598));
  jand g16343(.dina(n16598), .dinb(n16597), .dout(n16599));
  jand g16344(.dina(n16599), .dinb(n16596), .dout(n16600));
  jand g16345(.dina(n16600), .dinb(n16595), .dout(n16601));
  jxor g16346(.dina(n16601), .dinb(n2468), .dout(n16602));
  jxor g16347(.dina(n16602), .dinb(n16594), .dout(n16603));
  jand g16348(.dina(n16561), .dinb(n16443), .dout(n16604));
  jand g16349(.dina(n16570), .dinb(n16562), .dout(n16605));
  jor  g16350(.dina(n16605), .dinb(n16604), .dout(n16606));
  jand g16351(.dina(n16551), .dinb(n16446), .dout(n16607));
  jand g16352(.dina(n16560), .dinb(n16552), .dout(n16608));
  jor  g16353(.dina(n16608), .dinb(n16607), .dout(n16609));
  jand g16354(.dina(n16541), .dinb(n16449), .dout(n16610));
  jand g16355(.dina(n16550), .dinb(n16542), .dout(n16611));
  jor  g16356(.dina(n16611), .dinb(n16610), .dout(n16612));
  jand g16357(.dina(n16531), .dinb(n16452), .dout(n16613));
  jand g16358(.dina(n16540), .dinb(n16532), .dout(n16614));
  jor  g16359(.dina(n16614), .dinb(n16613), .dout(n16615));
  jand g16360(.dina(n16521), .dinb(n16455), .dout(n16616));
  jand g16361(.dina(n16530), .dinb(n16522), .dout(n16617));
  jor  g16362(.dina(n16617), .dinb(n16616), .dout(n16618));
  jand g16363(.dina(n16511), .dinb(n16458), .dout(n16619));
  jand g16364(.dina(n16520), .dinb(n16512), .dout(n16620));
  jor  g16365(.dina(n16620), .dinb(n16619), .dout(n16621));
  jand g16366(.dina(n16501), .dinb(n16461), .dout(n16622));
  jand g16367(.dina(n16510), .dinb(n16502), .dout(n16623));
  jor  g16368(.dina(n16623), .dinb(n16622), .dout(n16624));
  jand g16369(.dina(n16491), .dinb(n16464), .dout(n16625));
  jand g16370(.dina(n16500), .dinb(n16492), .dout(n16626));
  jor  g16371(.dina(n16626), .dinb(n16625), .dout(n16627));
  jand g16372(.dina(n16481), .dinb(n16467), .dout(n16628));
  jand g16373(.dina(n16490), .dinb(n16482), .dout(n16629));
  jor  g16374(.dina(n16629), .dinb(n16628), .dout(n16630));
  jor  g16375(.dina(n9271), .dinb(n3346), .dout(n16631));
  jor  g16376(.dina(n9003), .dinb(n3023), .dout(n16632));
  jor  g16377(.dina(n9268), .dinb(n3348), .dout(n16633));
  jor  g16378(.dina(n9273), .dinb(n3186), .dout(n16634));
  jand g16379(.dina(n16634), .dinb(n16633), .dout(n16635));
  jand g16380(.dina(n16635), .dinb(n16632), .dout(n16636));
  jand g16381(.dina(n16636), .dinb(n16631), .dout(n16637));
  jxor g16382(.dina(n16637), .dinb(n8729), .dout(n16638));
  jxor g16383(.dina(n16638), .dinb(n16630), .dout(n16639));
  jand g16384(.dina(n16471), .dinb(n16267), .dout(n16640));
  jand g16385(.dina(n16480), .dinb(n16472), .dout(n16641));
  jor  g16386(.dina(n16641), .dinb(n16640), .dout(n16642));
  jand g16387(.dina(n10594), .dinb(b26 ), .dout(n16643));
  jand g16388(.dina(n10129), .dinb(b27 ), .dout(n16644));
  jor  g16389(.dina(n16644), .dinb(n16643), .dout(n16645));
  jxor g16390(.dina(n16645), .dinb(n2057), .dout(n16646));
  jxor g16391(.dina(n16646), .dinb(n16470), .dout(n16647));
  jxor g16392(.dina(n16647), .dinb(n16642), .dout(n16648));
  jor  g16393(.dina(n10134), .dinb(n2860), .dout(n16649));
  jor  g16394(.dina(n9849), .dinb(n2563), .dout(n16650));
  jor  g16395(.dina(n10132), .dinb(n2862), .dout(n16651));
  jor  g16396(.dina(n10137), .dinb(n2713), .dout(n16652));
  jand g16397(.dina(n16652), .dinb(n16651), .dout(n16653));
  jand g16398(.dina(n16653), .dinb(n16650), .dout(n16654));
  jand g16399(.dina(n16654), .dinb(n16649), .dout(n16655));
  jxor g16400(.dina(n16655), .dinb(n9559), .dout(n16656));
  jxor g16401(.dina(n16656), .dinb(n16648), .dout(n16657));
  jxor g16402(.dina(n16657), .dinb(n16639), .dout(n16658));
  jor  g16403(.dina(n8457), .dinb(n3871), .dout(n16659));
  jor  g16404(.dina(n8185), .dinb(n3522), .dout(n16660));
  jor  g16405(.dina(n8454), .dinb(n3873), .dout(n16661));
  jor  g16406(.dina(n8459), .dinb(n3698), .dout(n16662));
  jand g16407(.dina(n16662), .dinb(n16661), .dout(n16663));
  jand g16408(.dina(n16663), .dinb(n16660), .dout(n16664));
  jand g16409(.dina(n16664), .dinb(n16659), .dout(n16665));
  jxor g16410(.dina(n16665), .dinb(n7929), .dout(n16666));
  jxor g16411(.dina(n16666), .dinb(n16658), .dout(n16667));
  jxor g16412(.dina(n16667), .dinb(n16627), .dout(n16668));
  jor  g16413(.dina(n7660), .dinb(n4435), .dout(n16669));
  jor  g16414(.dina(n7415), .dinb(n4060), .dout(n16670));
  jor  g16415(.dina(n7657), .dinb(n4249), .dout(n16671));
  jor  g16416(.dina(n7662), .dinb(n4437), .dout(n16672));
  jand g16417(.dina(n16672), .dinb(n16671), .dout(n16673));
  jand g16418(.dina(n16673), .dinb(n16670), .dout(n16674));
  jand g16419(.dina(n16674), .dinb(n16669), .dout(n16675));
  jxor g16420(.dina(n16675), .dinb(n7166), .dout(n16676));
  jxor g16421(.dina(n16676), .dinb(n16668), .dout(n16677));
  jxor g16422(.dina(n16677), .dinb(n16624), .dout(n16678));
  jor  g16423(.dina(n6914), .dinb(n5038), .dout(n16679));
  jor  g16424(.dina(n6673), .dinb(n4637), .dout(n16680));
  jor  g16425(.dina(n6911), .dinb(n4839), .dout(n16681));
  jor  g16426(.dina(n6916), .dinb(n5040), .dout(n16682));
  jand g16427(.dina(n16682), .dinb(n16681), .dout(n16683));
  jand g16428(.dina(n16683), .dinb(n16680), .dout(n16684));
  jand g16429(.dina(n16684), .dinb(n16679), .dout(n16685));
  jxor g16430(.dina(n16685), .dinb(n6443), .dout(n16686));
  jxor g16431(.dina(n16686), .dinb(n16678), .dout(n16687));
  jxor g16432(.dina(n16687), .dinb(n16621), .dout(n16688));
  jor  g16433(.dina(n6207), .dinb(n5683), .dout(n16689));
  jor  g16434(.dina(n5975), .dinb(n5253), .dout(n16690));
  jor  g16435(.dina(n6205), .dinb(n5685), .dout(n16691));
  jor  g16436(.dina(n6210), .dinb(n5469), .dout(n16692));
  jand g16437(.dina(n16692), .dinb(n16691), .dout(n16693));
  jand g16438(.dina(n16693), .dinb(n16690), .dout(n16694));
  jand g16439(.dina(n16694), .dinb(n16689), .dout(n16695));
  jxor g16440(.dina(n16695), .dinb(n5759), .dout(n16696));
  jxor g16441(.dina(n16696), .dinb(n16688), .dout(n16697));
  jxor g16442(.dina(n16697), .dinb(n16618), .dout(n16698));
  jor  g16443(.dina(n6364), .dinb(n5537), .dout(n16699));
  jor  g16444(.dina(n5315), .dinb(n5911), .dout(n16700));
  jor  g16445(.dina(n5534), .dinb(n6139), .dout(n16701));
  jor  g16446(.dina(n5539), .dinb(n6366), .dout(n16702));
  jand g16447(.dina(n16702), .dinb(n16701), .dout(n16703));
  jand g16448(.dina(n16703), .dinb(n16700), .dout(n16704));
  jand g16449(.dina(n16704), .dinb(n16699), .dout(n16705));
  jxor g16450(.dina(n16705), .dinb(n5111), .dout(n16706));
  jxor g16451(.dina(n16706), .dinb(n16698), .dout(n16707));
  jxor g16452(.dina(n16707), .dinb(n16615), .dout(n16708));
  jor  g16453(.dina(n7084), .dinb(n4902), .dout(n16709));
  jor  g16454(.dina(n4696), .dinb(n6605), .dout(n16710));
  jor  g16455(.dina(n4904), .dinb(n6846), .dout(n16711));
  jor  g16456(.dina(n4899), .dinb(n7086), .dout(n16712));
  jand g16457(.dina(n16712), .dinb(n16711), .dout(n16713));
  jand g16458(.dina(n16713), .dinb(n16710), .dout(n16714));
  jand g16459(.dina(n16714), .dinb(n16709), .dout(n16715));
  jxor g16460(.dina(n16715), .dinb(n4505), .dout(n16716));
  jxor g16461(.dina(n16716), .dinb(n16708), .dout(n16717));
  jxor g16462(.dina(n16717), .dinb(n16612), .dout(n16718));
  jor  g16463(.dina(n7844), .dinb(n4305), .dout(n16719));
  jor  g16464(.dina(n4116), .dinb(n7338), .dout(n16720));
  jor  g16465(.dina(n4308), .dinb(n7590), .dout(n16721));
  jor  g16466(.dina(n4303), .dinb(n7846), .dout(n16722));
  jand g16467(.dina(n16722), .dinb(n16721), .dout(n16723));
  jand g16468(.dina(n16723), .dinb(n16720), .dout(n16724));
  jand g16469(.dina(n16724), .dinb(n16719), .dout(n16725));
  jxor g16470(.dina(n16725), .dinb(n3938), .dout(n16726));
  jxor g16471(.dina(n16726), .dinb(n16718), .dout(n16727));
  jxor g16472(.dina(n16727), .dinb(n16609), .dout(n16728));
  jor  g16473(.dina(n8642), .dinb(n3751), .dout(n16729));
  jor  g16474(.dina(n3574), .dinb(n8111), .dout(n16730));
  jor  g16475(.dina(n3754), .dinb(n8378), .dout(n16731));
  jor  g16476(.dina(n3749), .dinb(n8644), .dout(n16732));
  jand g16477(.dina(n16732), .dinb(n16731), .dout(n16733));
  jand g16478(.dina(n16733), .dinb(n16730), .dout(n16734));
  jand g16479(.dina(n16734), .dinb(n16729), .dout(n16735));
  jxor g16480(.dina(n16735), .dinb(n3410), .dout(n16736));
  jxor g16481(.dina(n16736), .dinb(n16728), .dout(n16737));
  jxor g16482(.dina(n16737), .dinb(n16606), .dout(n16738));
  jand g16483(.dina(n16439), .dinb(n16431), .dout(n16739));
  jand g16484(.dina(n16571), .dinb(n16440), .dout(n16740));
  jor  g16485(.dina(n16740), .dinb(n16739), .dout(n16741));
  jor  g16486(.dina(n9473), .dinb(n3239), .dout(n16742));
  jor  g16487(.dina(n3072), .dinb(n8920), .dout(n16743));
  jor  g16488(.dina(n3237), .dinb(n9475), .dout(n16744));
  jor  g16489(.dina(n3242), .dinb(n9195), .dout(n16745));
  jand g16490(.dina(n16745), .dinb(n16744), .dout(n16746));
  jand g16491(.dina(n16746), .dinb(n16743), .dout(n16747));
  jand g16492(.dina(n16747), .dinb(n16742), .dout(n16748));
  jxor g16493(.dina(n16748), .dinb(n2918), .dout(n16749));
  jxor g16494(.dina(n16749), .dinb(n16741), .dout(n16750));
  jxor g16495(.dina(n16750), .dinb(n16738), .dout(n16751));
  jxor g16496(.dina(n16751), .dinb(n16603), .dout(n16752));
  jxor g16497(.dina(n16752), .dinb(n16591), .dout(n16753));
  jnot g16498(.din(n16753), .dout(n16754));
  jand g16499(.dina(n16583), .dinb(n16416), .dout(n16755));
  jnot g16500(.din(n16755), .dout(n16756));
  jor  g16501(.dina(n16585), .dinb(n16411), .dout(n16757));
  jand g16502(.dina(n16757), .dinb(n16756), .dout(n16758));
  jxor g16503(.dina(n16758), .dinb(n16754), .dout(f90 ));
  jand g16504(.dina(n16602), .dinb(n16594), .dout(n16760));
  jand g16505(.dina(n16751), .dinb(n16603), .dout(n16761));
  jor  g16506(.dina(n16761), .dinb(n16760), .dout(n16762));
  jand g16507(.dina(n16749), .dinb(n16741), .dout(n16763));
  jand g16508(.dina(n16750), .dinb(n16738), .dout(n16764));
  jor  g16509(.dina(n16764), .dinb(n16763), .dout(n16765));
  jnot g16510(.din(n16765), .dout(n16766));
  jor  g16511(.dina(n10813), .dinb(n2764), .dout(n16767));
  jor  g16512(.dina(n2609), .dinb(n10051), .dout(n16768));
  jor  g16513(.dina(n2766), .dinb(n10523), .dout(n16769));
  jand g16514(.dina(n16769), .dinb(n16768), .dout(n16770));
  jand g16515(.dina(n16770), .dinb(n16767), .dout(n16771));
  jxor g16516(.dina(n16771), .dinb(a29 ), .dout(n16772));
  jxor g16517(.dina(n16772), .dinb(n16766), .dout(n16773));
  jand g16518(.dina(n16736), .dinb(n16728), .dout(n16774));
  jand g16519(.dina(n16737), .dinb(n16606), .dout(n16775));
  jor  g16520(.dina(n16775), .dinb(n16774), .dout(n16776));
  jor  g16521(.dina(n9757), .dinb(n3239), .dout(n16777));
  jor  g16522(.dina(n3072), .dinb(n9195), .dout(n16778));
  jor  g16523(.dina(n3242), .dinb(n9475), .dout(n16779));
  jor  g16524(.dina(n3237), .dinb(n9759), .dout(n16780));
  jand g16525(.dina(n16780), .dinb(n16779), .dout(n16781));
  jand g16526(.dina(n16781), .dinb(n16778), .dout(n16782));
  jand g16527(.dina(n16782), .dinb(n16777), .dout(n16783));
  jxor g16528(.dina(n16783), .dinb(n2918), .dout(n16784));
  jxor g16529(.dina(n16784), .dinb(n16776), .dout(n16785));
  jand g16530(.dina(n16726), .dinb(n16718), .dout(n16786));
  jand g16531(.dina(n16727), .dinb(n16609), .dout(n16787));
  jor  g16532(.dina(n16787), .dinb(n16786), .dout(n16788));
  jand g16533(.dina(n16706), .dinb(n16698), .dout(n16789));
  jand g16534(.dina(n16707), .dinb(n16615), .dout(n16790));
  jor  g16535(.dina(n16790), .dinb(n16789), .dout(n16791));
  jand g16536(.dina(n16696), .dinb(n16688), .dout(n16792));
  jand g16537(.dina(n16697), .dinb(n16618), .dout(n16793));
  jor  g16538(.dina(n16793), .dinb(n16792), .dout(n16794));
  jand g16539(.dina(n16686), .dinb(n16678), .dout(n16795));
  jand g16540(.dina(n16687), .dinb(n16621), .dout(n16796));
  jor  g16541(.dina(n16796), .dinb(n16795), .dout(n16797));
  jand g16542(.dina(n16676), .dinb(n16668), .dout(n16798));
  jand g16543(.dina(n16677), .dinb(n16624), .dout(n16799));
  jor  g16544(.dina(n16799), .dinb(n16798), .dout(n16800));
  jand g16545(.dina(n16666), .dinb(n16658), .dout(n16801));
  jand g16546(.dina(n16667), .dinb(n16627), .dout(n16802));
  jor  g16547(.dina(n16802), .dinb(n16801), .dout(n16803));
  jand g16548(.dina(n16638), .dinb(n16630), .dout(n16804));
  jand g16549(.dina(n16657), .dinb(n16639), .dout(n16805));
  jor  g16550(.dina(n16805), .dinb(n16804), .dout(n16806));
  jand g16551(.dina(n10594), .dinb(b27 ), .dout(n16807));
  jand g16552(.dina(n10129), .dinb(b28 ), .dout(n16808));
  jor  g16553(.dina(n16808), .dinb(n16807), .dout(n16809));
  jnot g16554(.din(n16809), .dout(n16810));
  jand g16555(.dina(n16645), .dinb(n2057), .dout(n16811));
  jand g16556(.dina(n16646), .dinb(n16470), .dout(n16812));
  jor  g16557(.dina(n16812), .dinb(n16811), .dout(n16813));
  jxor g16558(.dina(n16813), .dinb(n16810), .dout(n16814));
  jor  g16559(.dina(n10134), .dinb(n3021), .dout(n16815));
  jor  g16560(.dina(n9849), .dinb(n2713), .dout(n16816));
  jor  g16561(.dina(n10132), .dinb(n3023), .dout(n16817));
  jor  g16562(.dina(n10137), .dinb(n2862), .dout(n16818));
  jand g16563(.dina(n16818), .dinb(n16817), .dout(n16819));
  jand g16564(.dina(n16819), .dinb(n16816), .dout(n16820));
  jand g16565(.dina(n16820), .dinb(n16815), .dout(n16821));
  jxor g16566(.dina(n16821), .dinb(n9559), .dout(n16822));
  jxor g16567(.dina(n16822), .dinb(n16814), .dout(n16823));
  jand g16568(.dina(n16647), .dinb(n16642), .dout(n16824));
  jand g16569(.dina(n16656), .dinb(n16648), .dout(n16825));
  jor  g16570(.dina(n16825), .dinb(n16824), .dout(n16826));
  jxor g16571(.dina(n16826), .dinb(n16823), .dout(n16827));
  jor  g16572(.dina(n9271), .dinb(n3520), .dout(n16828));
  jor  g16573(.dina(n9003), .dinb(n3186), .dout(n16829));
  jor  g16574(.dina(n9273), .dinb(n3348), .dout(n16830));
  jor  g16575(.dina(n9268), .dinb(n3522), .dout(n16831));
  jand g16576(.dina(n16831), .dinb(n16830), .dout(n16832));
  jand g16577(.dina(n16832), .dinb(n16829), .dout(n16833));
  jand g16578(.dina(n16833), .dinb(n16828), .dout(n16834));
  jxor g16579(.dina(n16834), .dinb(n8729), .dout(n16835));
  jxor g16580(.dina(n16835), .dinb(n16827), .dout(n16836));
  jxor g16581(.dina(n16836), .dinb(n16806), .dout(n16837));
  jor  g16582(.dina(n8457), .dinb(n4058), .dout(n16838));
  jor  g16583(.dina(n8185), .dinb(n3698), .dout(n16839));
  jor  g16584(.dina(n8459), .dinb(n3873), .dout(n16840));
  jor  g16585(.dina(n8454), .dinb(n4060), .dout(n16841));
  jand g16586(.dina(n16841), .dinb(n16840), .dout(n16842));
  jand g16587(.dina(n16842), .dinb(n16839), .dout(n16843));
  jand g16588(.dina(n16843), .dinb(n16838), .dout(n16844));
  jxor g16589(.dina(n16844), .dinb(n7929), .dout(n16845));
  jxor g16590(.dina(n16845), .dinb(n16837), .dout(n16846));
  jxor g16591(.dina(n16846), .dinb(n16803), .dout(n16847));
  jor  g16592(.dina(n7660), .dinb(n4635), .dout(n16848));
  jor  g16593(.dina(n7415), .dinb(n4249), .dout(n16849));
  jor  g16594(.dina(n7657), .dinb(n4437), .dout(n16850));
  jor  g16595(.dina(n7662), .dinb(n4637), .dout(n16851));
  jand g16596(.dina(n16851), .dinb(n16850), .dout(n16852));
  jand g16597(.dina(n16852), .dinb(n16849), .dout(n16853));
  jand g16598(.dina(n16853), .dinb(n16848), .dout(n16854));
  jxor g16599(.dina(n16854), .dinb(n7166), .dout(n16855));
  jxor g16600(.dina(n16855), .dinb(n16847), .dout(n16856));
  jxor g16601(.dina(n16856), .dinb(n16800), .dout(n16857));
  jor  g16602(.dina(n6914), .dinb(n5251), .dout(n16858));
  jor  g16603(.dina(n6673), .dinb(n4839), .dout(n16859));
  jor  g16604(.dina(n6911), .dinb(n5040), .dout(n16860));
  jor  g16605(.dina(n6916), .dinb(n5253), .dout(n16861));
  jand g16606(.dina(n16861), .dinb(n16860), .dout(n16862));
  jand g16607(.dina(n16862), .dinb(n16859), .dout(n16863));
  jand g16608(.dina(n16863), .dinb(n16858), .dout(n16864));
  jxor g16609(.dina(n16864), .dinb(n6443), .dout(n16865));
  jxor g16610(.dina(n16865), .dinb(n16857), .dout(n16866));
  jxor g16611(.dina(n16866), .dinb(n16797), .dout(n16867));
  jor  g16612(.dina(n5909), .dinb(n6207), .dout(n16868));
  jor  g16613(.dina(n5975), .dinb(n5469), .dout(n16869));
  jor  g16614(.dina(n6210), .dinb(n5685), .dout(n16870));
  jor  g16615(.dina(n6205), .dinb(n5911), .dout(n16871));
  jand g16616(.dina(n16871), .dinb(n16870), .dout(n16872));
  jand g16617(.dina(n16872), .dinb(n16869), .dout(n16873));
  jand g16618(.dina(n16873), .dinb(n16868), .dout(n16874));
  jxor g16619(.dina(n16874), .dinb(n5759), .dout(n16875));
  jxor g16620(.dina(n16875), .dinb(n16867), .dout(n16876));
  jxor g16621(.dina(n16876), .dinb(n16794), .dout(n16877));
  jor  g16622(.dina(n6603), .dinb(n5537), .dout(n16878));
  jor  g16623(.dina(n5315), .dinb(n6139), .dout(n16879));
  jor  g16624(.dina(n5539), .dinb(n6605), .dout(n16880));
  jor  g16625(.dina(n5534), .dinb(n6366), .dout(n16881));
  jand g16626(.dina(n16881), .dinb(n16880), .dout(n16882));
  jand g16627(.dina(n16882), .dinb(n16879), .dout(n16883));
  jand g16628(.dina(n16883), .dinb(n16878), .dout(n16884));
  jxor g16629(.dina(n16884), .dinb(n5111), .dout(n16885));
  jxor g16630(.dina(n16885), .dinb(n16877), .dout(n16886));
  jxor g16631(.dina(n16886), .dinb(n16791), .dout(n16887));
  jor  g16632(.dina(n7336), .dinb(n4902), .dout(n16888));
  jor  g16633(.dina(n4696), .dinb(n6846), .dout(n16889));
  jor  g16634(.dina(n4899), .dinb(n7338), .dout(n16890));
  jor  g16635(.dina(n4904), .dinb(n7086), .dout(n16891));
  jand g16636(.dina(n16891), .dinb(n16890), .dout(n16892));
  jand g16637(.dina(n16892), .dinb(n16889), .dout(n16893));
  jand g16638(.dina(n16893), .dinb(n16888), .dout(n16894));
  jxor g16639(.dina(n16894), .dinb(n4505), .dout(n16895));
  jxor g16640(.dina(n16895), .dinb(n16887), .dout(n16896));
  jnot g16641(.din(n16708), .dout(n16897));
  jnot g16642(.din(n16716), .dout(n16898));
  jand g16643(.dina(n16898), .dinb(n16897), .dout(n16899));
  jnot g16644(.din(n16899), .dout(n16900));
  jand g16645(.dina(n16716), .dinb(n16708), .dout(n16901));
  jor  g16646(.dina(n16901), .dinb(n16612), .dout(n16902));
  jand g16647(.dina(n16902), .dinb(n16900), .dout(n16903));
  jxor g16648(.dina(n16903), .dinb(n16896), .dout(n16904));
  jor  g16649(.dina(n8109), .dinb(n4305), .dout(n16905));
  jor  g16650(.dina(n4116), .dinb(n7590), .dout(n16906));
  jor  g16651(.dina(n4303), .dinb(n8111), .dout(n16907));
  jor  g16652(.dina(n4308), .dinb(n7846), .dout(n16908));
  jand g16653(.dina(n16908), .dinb(n16907), .dout(n16909));
  jand g16654(.dina(n16909), .dinb(n16906), .dout(n16910));
  jand g16655(.dina(n16910), .dinb(n16905), .dout(n16911));
  jxor g16656(.dina(n16911), .dinb(n3938), .dout(n16912));
  jxor g16657(.dina(n16912), .dinb(n16904), .dout(n16913));
  jxor g16658(.dina(n16913), .dinb(n16788), .dout(n16914));
  jor  g16659(.dina(n8918), .dinb(n3751), .dout(n16915));
  jor  g16660(.dina(n3574), .dinb(n8378), .dout(n16916));
  jor  g16661(.dina(n3754), .dinb(n8644), .dout(n16917));
  jor  g16662(.dina(n3749), .dinb(n8920), .dout(n16918));
  jand g16663(.dina(n16918), .dinb(n16917), .dout(n16919));
  jand g16664(.dina(n16919), .dinb(n16916), .dout(n16920));
  jand g16665(.dina(n16920), .dinb(n16915), .dout(n16921));
  jxor g16666(.dina(n16921), .dinb(n3410), .dout(n16922));
  jxor g16667(.dina(n16922), .dinb(n16914), .dout(n16923));
  jxor g16668(.dina(n16923), .dinb(n16785), .dout(n16924));
  jxor g16669(.dina(n16924), .dinb(n16773), .dout(n16925));
  jxor g16670(.dina(n16925), .dinb(n16762), .dout(n16926));
  jnot g16671(.din(n16926), .dout(n16927));
  jand g16672(.dina(n16752), .dinb(n16591), .dout(n16928));
  jnot g16673(.din(n16928), .dout(n16929));
  jor  g16674(.dina(n16758), .dinb(n16754), .dout(n16930));
  jand g16675(.dina(n16930), .dinb(n16929), .dout(n16931));
  jxor g16676(.dina(n16931), .dinb(n16927), .dout(f91 ));
  jand g16677(.dina(n16925), .dinb(n16762), .dout(n16933));
  jnot g16678(.din(n16933), .dout(n16934));
  jor  g16679(.dina(n16931), .dinb(n16927), .dout(n16935));
  jand g16680(.dina(n16935), .dinb(n16934), .dout(n16936));
  jor  g16681(.dina(n16772), .dinb(n16766), .dout(n16937));
  jand g16682(.dina(n16924), .dinb(n16773), .dout(n16938));
  jnot g16683(.din(n16938), .dout(n16939));
  jand g16684(.dina(n16939), .dinb(n16937), .dout(n16940));
  jnot g16685(.din(n16940), .dout(n16941));
  jand g16686(.dina(n16913), .dinb(n16788), .dout(n16942));
  jand g16687(.dina(n16922), .dinb(n16914), .dout(n16943));
  jor  g16688(.dina(n16943), .dinb(n16942), .dout(n16944));
  jor  g16689(.dina(n10049), .dinb(n3239), .dout(n16945));
  jor  g16690(.dina(n3072), .dinb(n9475), .dout(n16946));
  jor  g16691(.dina(n3237), .dinb(n10051), .dout(n16947));
  jor  g16692(.dina(n3242), .dinb(n9759), .dout(n16948));
  jand g16693(.dina(n16948), .dinb(n16947), .dout(n16949));
  jand g16694(.dina(n16949), .dinb(n16946), .dout(n16950));
  jand g16695(.dina(n16950), .dinb(n16945), .dout(n16951));
  jxor g16696(.dina(n16951), .dinb(n2918), .dout(n16952));
  jxor g16697(.dina(n16952), .dinb(n16944), .dout(n16953));
  jand g16698(.dina(n16903), .dinb(n16896), .dout(n16954));
  jand g16699(.dina(n16912), .dinb(n16904), .dout(n16955));
  jor  g16700(.dina(n16955), .dinb(n16954), .dout(n16956));
  jand g16701(.dina(n16886), .dinb(n16791), .dout(n16957));
  jand g16702(.dina(n16895), .dinb(n16887), .dout(n16958));
  jor  g16703(.dina(n16958), .dinb(n16957), .dout(n16959));
  jand g16704(.dina(n16876), .dinb(n16794), .dout(n16960));
  jand g16705(.dina(n16885), .dinb(n16877), .dout(n16961));
  jor  g16706(.dina(n16961), .dinb(n16960), .dout(n16962));
  jand g16707(.dina(n16866), .dinb(n16797), .dout(n16963));
  jand g16708(.dina(n16875), .dinb(n16867), .dout(n16964));
  jor  g16709(.dina(n16964), .dinb(n16963), .dout(n16965));
  jand g16710(.dina(n16856), .dinb(n16800), .dout(n16966));
  jand g16711(.dina(n16865), .dinb(n16857), .dout(n16967));
  jor  g16712(.dina(n16967), .dinb(n16966), .dout(n16968));
  jand g16713(.dina(n16846), .dinb(n16803), .dout(n16969));
  jand g16714(.dina(n16855), .dinb(n16847), .dout(n16970));
  jor  g16715(.dina(n16970), .dinb(n16969), .dout(n16971));
  jand g16716(.dina(n16836), .dinb(n16806), .dout(n16972));
  jand g16717(.dina(n16845), .dinb(n16837), .dout(n16973));
  jor  g16718(.dina(n16973), .dinb(n16972), .dout(n16974));
  jand g16719(.dina(n16826), .dinb(n16823), .dout(n16975));
  jand g16720(.dina(n16835), .dinb(n16827), .dout(n16976));
  jor  g16721(.dina(n16976), .dinb(n16975), .dout(n16977));
  jand g16722(.dina(n16813), .dinb(n16810), .dout(n16978));
  jand g16723(.dina(n16822), .dinb(n16814), .dout(n16979));
  jor  g16724(.dina(n16979), .dinb(n16978), .dout(n16980));
  jand g16725(.dina(n10594), .dinb(b28 ), .dout(n16981));
  jand g16726(.dina(n10129), .dinb(b29 ), .dout(n16982));
  jor  g16727(.dina(n16982), .dinb(n16981), .dout(n16983));
  jnot g16728(.din(n16983), .dout(n16984));
  jxor g16729(.dina(n16984), .dinb(n16809), .dout(n16985));
  jxor g16730(.dina(n16985), .dinb(n16980), .dout(n16986));
  jor  g16731(.dina(n10134), .dinb(n3184), .dout(n16987));
  jor  g16732(.dina(n9849), .dinb(n2862), .dout(n16988));
  jor  g16733(.dina(n10132), .dinb(n3186), .dout(n16989));
  jor  g16734(.dina(n10137), .dinb(n3023), .dout(n16990));
  jand g16735(.dina(n16990), .dinb(n16989), .dout(n16991));
  jand g16736(.dina(n16991), .dinb(n16988), .dout(n16992));
  jand g16737(.dina(n16992), .dinb(n16987), .dout(n16993));
  jxor g16738(.dina(n16993), .dinb(n9559), .dout(n16994));
  jxor g16739(.dina(n16994), .dinb(n16986), .dout(n16995));
  jor  g16740(.dina(n9271), .dinb(n3696), .dout(n16996));
  jor  g16741(.dina(n9003), .dinb(n3348), .dout(n16997));
  jor  g16742(.dina(n9273), .dinb(n3522), .dout(n16998));
  jor  g16743(.dina(n9268), .dinb(n3698), .dout(n16999));
  jand g16744(.dina(n16999), .dinb(n16998), .dout(n17000));
  jand g16745(.dina(n17000), .dinb(n16997), .dout(n17001));
  jand g16746(.dina(n17001), .dinb(n16996), .dout(n17002));
  jxor g16747(.dina(n17002), .dinb(n8729), .dout(n17003));
  jxor g16748(.dina(n17003), .dinb(n16995), .dout(n17004));
  jxor g16749(.dina(n17004), .dinb(n16977), .dout(n17005));
  jor  g16750(.dina(n8457), .dinb(n4247), .dout(n17006));
  jor  g16751(.dina(n8185), .dinb(n3873), .dout(n17007));
  jor  g16752(.dina(n8454), .dinb(n4249), .dout(n17008));
  jor  g16753(.dina(n8459), .dinb(n4060), .dout(n17009));
  jand g16754(.dina(n17009), .dinb(n17008), .dout(n17010));
  jand g16755(.dina(n17010), .dinb(n17007), .dout(n17011));
  jand g16756(.dina(n17011), .dinb(n17006), .dout(n17012));
  jxor g16757(.dina(n17012), .dinb(n7929), .dout(n17013));
  jxor g16758(.dina(n17013), .dinb(n17005), .dout(n17014));
  jxor g16759(.dina(n17014), .dinb(n16974), .dout(n17015));
  jor  g16760(.dina(n7660), .dinb(n4837), .dout(n17016));
  jor  g16761(.dina(n7415), .dinb(n4437), .dout(n17017));
  jor  g16762(.dina(n7657), .dinb(n4637), .dout(n17018));
  jor  g16763(.dina(n7662), .dinb(n4839), .dout(n17019));
  jand g16764(.dina(n17019), .dinb(n17018), .dout(n17020));
  jand g16765(.dina(n17020), .dinb(n17017), .dout(n17021));
  jand g16766(.dina(n17021), .dinb(n17016), .dout(n17022));
  jxor g16767(.dina(n17022), .dinb(n7166), .dout(n17023));
  jxor g16768(.dina(n17023), .dinb(n17015), .dout(n17024));
  jxor g16769(.dina(n17024), .dinb(n16971), .dout(n17025));
  jor  g16770(.dina(n6914), .dinb(n5467), .dout(n17026));
  jor  g16771(.dina(n6673), .dinb(n5040), .dout(n17027));
  jor  g16772(.dina(n6916), .dinb(n5469), .dout(n17028));
  jor  g16773(.dina(n6911), .dinb(n5253), .dout(n17029));
  jand g16774(.dina(n17029), .dinb(n17028), .dout(n17030));
  jand g16775(.dina(n17030), .dinb(n17027), .dout(n17031));
  jand g16776(.dina(n17031), .dinb(n17026), .dout(n17032));
  jxor g16777(.dina(n17032), .dinb(n6443), .dout(n17033));
  jxor g16778(.dina(n17033), .dinb(n17025), .dout(n17034));
  jxor g16779(.dina(n17034), .dinb(n16968), .dout(n17035));
  jor  g16780(.dina(n6137), .dinb(n6207), .dout(n17036));
  jor  g16781(.dina(n5975), .dinb(n5685), .dout(n17037));
  jor  g16782(.dina(n6210), .dinb(n5911), .dout(n17038));
  jor  g16783(.dina(n6205), .dinb(n6139), .dout(n17039));
  jand g16784(.dina(n17039), .dinb(n17038), .dout(n17040));
  jand g16785(.dina(n17040), .dinb(n17037), .dout(n17041));
  jand g16786(.dina(n17041), .dinb(n17036), .dout(n17042));
  jxor g16787(.dina(n17042), .dinb(n5759), .dout(n17043));
  jxor g16788(.dina(n17043), .dinb(n17035), .dout(n17044));
  jxor g16789(.dina(n17044), .dinb(n16965), .dout(n17045));
  jor  g16790(.dina(n6844), .dinb(n5537), .dout(n17046));
  jor  g16791(.dina(n5315), .dinb(n6366), .dout(n17047));
  jor  g16792(.dina(n5534), .dinb(n6605), .dout(n17048));
  jor  g16793(.dina(n5539), .dinb(n6846), .dout(n17049));
  jand g16794(.dina(n17049), .dinb(n17048), .dout(n17050));
  jand g16795(.dina(n17050), .dinb(n17047), .dout(n17051));
  jand g16796(.dina(n17051), .dinb(n17046), .dout(n17052));
  jxor g16797(.dina(n17052), .dinb(n5111), .dout(n17053));
  jxor g16798(.dina(n17053), .dinb(n17045), .dout(n17054));
  jxor g16799(.dina(n17054), .dinb(n16962), .dout(n17055));
  jor  g16800(.dina(n7588), .dinb(n4902), .dout(n17056));
  jor  g16801(.dina(n4696), .dinb(n7086), .dout(n17057));
  jor  g16802(.dina(n4904), .dinb(n7338), .dout(n17058));
  jor  g16803(.dina(n4899), .dinb(n7590), .dout(n17059));
  jand g16804(.dina(n17059), .dinb(n17058), .dout(n17060));
  jand g16805(.dina(n17060), .dinb(n17057), .dout(n17061));
  jand g16806(.dina(n17061), .dinb(n17056), .dout(n17062));
  jxor g16807(.dina(n17062), .dinb(n4505), .dout(n17063));
  jxor g16808(.dina(n17063), .dinb(n17055), .dout(n17064));
  jxor g16809(.dina(n17064), .dinb(n16959), .dout(n17065));
  jor  g16810(.dina(n8376), .dinb(n4305), .dout(n17066));
  jor  g16811(.dina(n4116), .dinb(n7846), .dout(n17067));
  jor  g16812(.dina(n4303), .dinb(n8378), .dout(n17068));
  jor  g16813(.dina(n4308), .dinb(n8111), .dout(n17069));
  jand g16814(.dina(n17069), .dinb(n17068), .dout(n17070));
  jand g16815(.dina(n17070), .dinb(n17067), .dout(n17071));
  jand g16816(.dina(n17071), .dinb(n17066), .dout(n17072));
  jxor g16817(.dina(n17072), .dinb(n3938), .dout(n17073));
  jxor g16818(.dina(n17073), .dinb(n17065), .dout(n17074));
  jxor g16819(.dina(n17074), .dinb(n16956), .dout(n17075));
  jor  g16820(.dina(n9193), .dinb(n3751), .dout(n17076));
  jor  g16821(.dina(n3574), .dinb(n8644), .dout(n17077));
  jor  g16822(.dina(n3754), .dinb(n8920), .dout(n17078));
  jor  g16823(.dina(n3749), .dinb(n9195), .dout(n17079));
  jand g16824(.dina(n17079), .dinb(n17078), .dout(n17080));
  jand g16825(.dina(n17080), .dinb(n17077), .dout(n17081));
  jand g16826(.dina(n17081), .dinb(n17076), .dout(n17082));
  jxor g16827(.dina(n17082), .dinb(n3410), .dout(n17083));
  jxor g16828(.dina(n17083), .dinb(n17075), .dout(n17084));
  jxor g16829(.dina(n17084), .dinb(n16953), .dout(n17085));
  jand g16830(.dina(n16784), .dinb(n16776), .dout(n17086));
  jand g16831(.dina(n16923), .dinb(n16785), .dout(n17087));
  jor  g16832(.dina(n17087), .dinb(n17086), .dout(n17088));
  jnot g16833(.din(n17088), .dout(n17089));
  jand g16834(.dina(n2610), .dinb(b63 ), .dout(n17090));
  jand g16835(.dina(n10832), .dinb(n2460), .dout(n17091));
  jor  g16836(.dina(n17091), .dinb(n17090), .dout(n17092));
  jxor g16837(.dina(n17092), .dinb(n2468), .dout(n17093));
  jxor g16838(.dina(n17093), .dinb(n17089), .dout(n17094));
  jxor g16839(.dina(n17094), .dinb(n17085), .dout(n17095));
  jxor g16840(.dina(n17095), .dinb(n16941), .dout(n17096));
  jnot g16841(.din(n17096), .dout(n17097));
  jxor g16842(.dina(n17097), .dinb(n16936), .dout(f92 ));
  jand g16843(.dina(n17095), .dinb(n16941), .dout(n17099));
  jnot g16844(.din(n17099), .dout(n17100));
  jor  g16845(.dina(n17097), .dinb(n16936), .dout(n17101));
  jand g16846(.dina(n17101), .dinb(n17100), .dout(n17102));
  jor  g16847(.dina(n17093), .dinb(n17089), .dout(n17103));
  jand g16848(.dina(n17094), .dinb(n17085), .dout(n17104));
  jnot g16849(.din(n17104), .dout(n17105));
  jand g16850(.dina(n17105), .dinb(n17103), .dout(n17106));
  jnot g16851(.din(n17106), .dout(n17107));
  jand g16852(.dina(n17074), .dinb(n16956), .dout(n17108));
  jand g16853(.dina(n17083), .dinb(n17075), .dout(n17109));
  jor  g16854(.dina(n17109), .dinb(n17108), .dout(n17110));
  jand g16855(.dina(n17064), .dinb(n16959), .dout(n17111));
  jand g16856(.dina(n17073), .dinb(n17065), .dout(n17112));
  jor  g16857(.dina(n17112), .dinb(n17111), .dout(n17113));
  jand g16858(.dina(n17054), .dinb(n16962), .dout(n17114));
  jand g16859(.dina(n17063), .dinb(n17055), .dout(n17115));
  jor  g16860(.dina(n17115), .dinb(n17114), .dout(n17116));
  jor  g16861(.dina(n7844), .dinb(n4902), .dout(n17117));
  jor  g16862(.dina(n4696), .dinb(n7338), .dout(n17118));
  jor  g16863(.dina(n4899), .dinb(n7846), .dout(n17119));
  jor  g16864(.dina(n4904), .dinb(n7590), .dout(n17120));
  jand g16865(.dina(n17120), .dinb(n17119), .dout(n17121));
  jand g16866(.dina(n17121), .dinb(n17118), .dout(n17122));
  jand g16867(.dina(n17122), .dinb(n17117), .dout(n17123));
  jxor g16868(.dina(n17123), .dinb(n4505), .dout(n17124));
  jnot g16869(.din(n17124), .dout(n17125));
  jand g16870(.dina(n17044), .dinb(n16965), .dout(n17126));
  jand g16871(.dina(n17053), .dinb(n17045), .dout(n17127));
  jor  g16872(.dina(n17127), .dinb(n17126), .dout(n17128));
  jand g16873(.dina(n17034), .dinb(n16968), .dout(n17129));
  jand g16874(.dina(n17043), .dinb(n17035), .dout(n17130));
  jor  g16875(.dina(n17130), .dinb(n17129), .dout(n17131));
  jand g16876(.dina(n17024), .dinb(n16971), .dout(n17132));
  jand g16877(.dina(n17033), .dinb(n17025), .dout(n17133));
  jor  g16878(.dina(n17133), .dinb(n17132), .dout(n17134));
  jand g16879(.dina(n17014), .dinb(n16974), .dout(n17135));
  jand g16880(.dina(n17023), .dinb(n17015), .dout(n17136));
  jor  g16881(.dina(n17136), .dinb(n17135), .dout(n17137));
  jand g16882(.dina(n17004), .dinb(n16977), .dout(n17138));
  jand g16883(.dina(n17013), .dinb(n17005), .dout(n17139));
  jor  g16884(.dina(n17139), .dinb(n17138), .dout(n17140));
  jand g16885(.dina(n16994), .dinb(n16986), .dout(n17141));
  jand g16886(.dina(n17003), .dinb(n16995), .dout(n17142));
  jor  g16887(.dina(n17142), .dinb(n17141), .dout(n17143));
  jand g16888(.dina(n16984), .dinb(n16809), .dout(n17144));
  jand g16889(.dina(n16985), .dinb(n16980), .dout(n17145));
  jor  g16890(.dina(n17145), .dinb(n17144), .dout(n17146));
  jand g16891(.dina(n10594), .dinb(b29 ), .dout(n17147));
  jand g16892(.dina(n10129), .dinb(b30 ), .dout(n17148));
  jor  g16893(.dina(n17148), .dinb(n17147), .dout(n17149));
  jxor g16894(.dina(n17149), .dinb(n2468), .dout(n17150));
  jxor g16895(.dina(n17150), .dinb(n16983), .dout(n17151));
  jxor g16896(.dina(n17151), .dinb(n17146), .dout(n17152));
  jor  g16897(.dina(n10134), .dinb(n3346), .dout(n17153));
  jor  g16898(.dina(n9849), .dinb(n3023), .dout(n17154));
  jor  g16899(.dina(n10137), .dinb(n3186), .dout(n17155));
  jor  g16900(.dina(n10132), .dinb(n3348), .dout(n17156));
  jand g16901(.dina(n17156), .dinb(n17155), .dout(n17157));
  jand g16902(.dina(n17157), .dinb(n17154), .dout(n17158));
  jand g16903(.dina(n17158), .dinb(n17153), .dout(n17159));
  jxor g16904(.dina(n17159), .dinb(n9559), .dout(n17160));
  jxor g16905(.dina(n17160), .dinb(n17152), .dout(n17161));
  jor  g16906(.dina(n9271), .dinb(n3871), .dout(n17162));
  jor  g16907(.dina(n9003), .dinb(n3522), .dout(n17163));
  jor  g16908(.dina(n9273), .dinb(n3698), .dout(n17164));
  jor  g16909(.dina(n9268), .dinb(n3873), .dout(n17165));
  jand g16910(.dina(n17165), .dinb(n17164), .dout(n17166));
  jand g16911(.dina(n17166), .dinb(n17163), .dout(n17167));
  jand g16912(.dina(n17167), .dinb(n17162), .dout(n17168));
  jxor g16913(.dina(n17168), .dinb(n8729), .dout(n17169));
  jxor g16914(.dina(n17169), .dinb(n17161), .dout(n17170));
  jxor g16915(.dina(n17170), .dinb(n17143), .dout(n17171));
  jor  g16916(.dina(n8457), .dinb(n4435), .dout(n17172));
  jor  g16917(.dina(n8185), .dinb(n4060), .dout(n17173));
  jor  g16918(.dina(n8459), .dinb(n4249), .dout(n17174));
  jor  g16919(.dina(n8454), .dinb(n4437), .dout(n17175));
  jand g16920(.dina(n17175), .dinb(n17174), .dout(n17176));
  jand g16921(.dina(n17176), .dinb(n17173), .dout(n17177));
  jand g16922(.dina(n17177), .dinb(n17172), .dout(n17178));
  jxor g16923(.dina(n17178), .dinb(n7929), .dout(n17179));
  jxor g16924(.dina(n17179), .dinb(n17171), .dout(n17180));
  jxor g16925(.dina(n17180), .dinb(n17140), .dout(n17181));
  jor  g16926(.dina(n7660), .dinb(n5038), .dout(n17182));
  jor  g16927(.dina(n7415), .dinb(n4637), .dout(n17183));
  jor  g16928(.dina(n7657), .dinb(n4839), .dout(n17184));
  jor  g16929(.dina(n7662), .dinb(n5040), .dout(n17185));
  jand g16930(.dina(n17185), .dinb(n17184), .dout(n17186));
  jand g16931(.dina(n17186), .dinb(n17183), .dout(n17187));
  jand g16932(.dina(n17187), .dinb(n17182), .dout(n17188));
  jxor g16933(.dina(n17188), .dinb(n7166), .dout(n17189));
  jxor g16934(.dina(n17189), .dinb(n17181), .dout(n17190));
  jxor g16935(.dina(n17190), .dinb(n17137), .dout(n17191));
  jor  g16936(.dina(n6914), .dinb(n5683), .dout(n17192));
  jor  g16937(.dina(n6673), .dinb(n5253), .dout(n17193));
  jor  g16938(.dina(n6916), .dinb(n5685), .dout(n17194));
  jor  g16939(.dina(n6911), .dinb(n5469), .dout(n17195));
  jand g16940(.dina(n17195), .dinb(n17194), .dout(n17196));
  jand g16941(.dina(n17196), .dinb(n17193), .dout(n17197));
  jand g16942(.dina(n17197), .dinb(n17192), .dout(n17198));
  jxor g16943(.dina(n17198), .dinb(n6443), .dout(n17199));
  jxor g16944(.dina(n17199), .dinb(n17191), .dout(n17200));
  jxor g16945(.dina(n17200), .dinb(n17134), .dout(n17201));
  jor  g16946(.dina(n6364), .dinb(n6207), .dout(n17202));
  jor  g16947(.dina(n5975), .dinb(n5911), .dout(n17203));
  jor  g16948(.dina(n6205), .dinb(n6366), .dout(n17204));
  jor  g16949(.dina(n6210), .dinb(n6139), .dout(n17205));
  jand g16950(.dina(n17205), .dinb(n17204), .dout(n17206));
  jand g16951(.dina(n17206), .dinb(n17203), .dout(n17207));
  jand g16952(.dina(n17207), .dinb(n17202), .dout(n17208));
  jxor g16953(.dina(n17208), .dinb(n5759), .dout(n17209));
  jxor g16954(.dina(n17209), .dinb(n17201), .dout(n17210));
  jxor g16955(.dina(n17210), .dinb(n17131), .dout(n17211));
  jnot g16956(.din(n17211), .dout(n17212));
  jor  g16957(.dina(n7084), .dinb(n5537), .dout(n17213));
  jor  g16958(.dina(n5315), .dinb(n6605), .dout(n17214));
  jor  g16959(.dina(n5534), .dinb(n6846), .dout(n17215));
  jor  g16960(.dina(n5539), .dinb(n7086), .dout(n17216));
  jand g16961(.dina(n17216), .dinb(n17215), .dout(n17217));
  jand g16962(.dina(n17217), .dinb(n17214), .dout(n17218));
  jand g16963(.dina(n17218), .dinb(n17213), .dout(n17219));
  jxor g16964(.dina(n17219), .dinb(n5111), .dout(n17220));
  jxor g16965(.dina(n17220), .dinb(n17212), .dout(n17221));
  jxor g16966(.dina(n17221), .dinb(n17128), .dout(n17222));
  jxor g16967(.dina(n17222), .dinb(n17125), .dout(n17223));
  jxor g16968(.dina(n17223), .dinb(n17116), .dout(n17224));
  jor  g16969(.dina(n8642), .dinb(n4305), .dout(n17225));
  jor  g16970(.dina(n4116), .dinb(n8111), .dout(n17226));
  jor  g16971(.dina(n4308), .dinb(n8378), .dout(n17227));
  jor  g16972(.dina(n4303), .dinb(n8644), .dout(n17228));
  jand g16973(.dina(n17228), .dinb(n17227), .dout(n17229));
  jand g16974(.dina(n17229), .dinb(n17226), .dout(n17230));
  jand g16975(.dina(n17230), .dinb(n17225), .dout(n17231));
  jxor g16976(.dina(n17231), .dinb(n3938), .dout(n17232));
  jxor g16977(.dina(n17232), .dinb(n17224), .dout(n17233));
  jxor g16978(.dina(n17233), .dinb(n17113), .dout(n17234));
  jor  g16979(.dina(n9473), .dinb(n3751), .dout(n17235));
  jor  g16980(.dina(n3574), .dinb(n8920), .dout(n17236));
  jor  g16981(.dina(n3754), .dinb(n9195), .dout(n17237));
  jor  g16982(.dina(n3749), .dinb(n9475), .dout(n17238));
  jand g16983(.dina(n17238), .dinb(n17237), .dout(n17239));
  jand g16984(.dina(n17239), .dinb(n17236), .dout(n17240));
  jand g16985(.dina(n17240), .dinb(n17235), .dout(n17241));
  jxor g16986(.dina(n17241), .dinb(n3410), .dout(n17242));
  jxor g16987(.dina(n17242), .dinb(n17234), .dout(n17243));
  jxor g16988(.dina(n17243), .dinb(n17110), .dout(n17244));
  jand g16989(.dina(n16952), .dinb(n16944), .dout(n17245));
  jand g16990(.dina(n17084), .dinb(n16953), .dout(n17246));
  jor  g16991(.dina(n17246), .dinb(n17245), .dout(n17247));
  jor  g16992(.dina(n10521), .dinb(n3239), .dout(n17248));
  jor  g16993(.dina(n3072), .dinb(n9759), .dout(n17249));
  jor  g16994(.dina(n3242), .dinb(n10051), .dout(n17250));
  jor  g16995(.dina(n3237), .dinb(n10523), .dout(n17251));
  jand g16996(.dina(n17251), .dinb(n17250), .dout(n17252));
  jand g16997(.dina(n17252), .dinb(n17249), .dout(n17253));
  jand g16998(.dina(n17253), .dinb(n17248), .dout(n17254));
  jxor g16999(.dina(n17254), .dinb(n2918), .dout(n17255));
  jxor g17000(.dina(n17255), .dinb(n17247), .dout(n17256));
  jxor g17001(.dina(n17256), .dinb(n17244), .dout(n17257));
  jxor g17002(.dina(n17257), .dinb(n17107), .dout(n17258));
  jnot g17003(.din(n17258), .dout(n17259));
  jxor g17004(.dina(n17259), .dinb(n17102), .dout(f93 ));
  jand g17005(.dina(n17257), .dinb(n17107), .dout(n17261));
  jnot g17006(.din(n17261), .dout(n17262));
  jor  g17007(.dina(n17259), .dinb(n17102), .dout(n17263));
  jand g17008(.dina(n17263), .dinb(n17262), .dout(n17264));
  jand g17009(.dina(n17255), .dinb(n17247), .dout(n17265));
  jand g17010(.dina(n17256), .dinb(n17244), .dout(n17266));
  jor  g17011(.dina(n17266), .dinb(n17265), .dout(n17267));
  jand g17012(.dina(n17242), .dinb(n17234), .dout(n17268));
  jand g17013(.dina(n17243), .dinb(n17110), .dout(n17269));
  jor  g17014(.dina(n17269), .dinb(n17268), .dout(n17270));
  jnot g17015(.din(n17270), .dout(n17271));
  jor  g17016(.dina(n10813), .dinb(n3239), .dout(n17272));
  jor  g17017(.dina(n3072), .dinb(n10051), .dout(n17273));
  jor  g17018(.dina(n3242), .dinb(n10523), .dout(n17274));
  jand g17019(.dina(n17274), .dinb(n17273), .dout(n17275));
  jand g17020(.dina(n17275), .dinb(n17272), .dout(n17276));
  jxor g17021(.dina(n17276), .dinb(a32 ), .dout(n17277));
  jxor g17022(.dina(n17277), .dinb(n17271), .dout(n17278));
  jand g17023(.dina(n17232), .dinb(n17224), .dout(n17279));
  jand g17024(.dina(n17233), .dinb(n17113), .dout(n17280));
  jor  g17025(.dina(n17280), .dinb(n17279), .dout(n17281));
  jor  g17026(.dina(n17222), .dinb(n17125), .dout(n17282));
  jand g17027(.dina(n17223), .dinb(n17116), .dout(n17283));
  jnot g17028(.din(n17283), .dout(n17284));
  jand g17029(.dina(n17284), .dinb(n17282), .dout(n17285));
  jnot g17030(.din(n17285), .dout(n17286));
  jand g17031(.dina(n17209), .dinb(n17201), .dout(n17287));
  jand g17032(.dina(n17210), .dinb(n17131), .dout(n17288));
  jor  g17033(.dina(n17288), .dinb(n17287), .dout(n17289));
  jand g17034(.dina(n17199), .dinb(n17191), .dout(n17290));
  jand g17035(.dina(n17200), .dinb(n17134), .dout(n17291));
  jor  g17036(.dina(n17291), .dinb(n17290), .dout(n17292));
  jand g17037(.dina(n17189), .dinb(n17181), .dout(n17293));
  jand g17038(.dina(n17190), .dinb(n17137), .dout(n17294));
  jor  g17039(.dina(n17294), .dinb(n17293), .dout(n17295));
  jand g17040(.dina(n17179), .dinb(n17171), .dout(n17296));
  jand g17041(.dina(n17180), .dinb(n17140), .dout(n17297));
  jor  g17042(.dina(n17297), .dinb(n17296), .dout(n17298));
  jand g17043(.dina(n17169), .dinb(n17161), .dout(n17299));
  jand g17044(.dina(n17170), .dinb(n17143), .dout(n17300));
  jor  g17045(.dina(n17300), .dinb(n17299), .dout(n17301));
  jand g17046(.dina(n17151), .dinb(n17146), .dout(n17302));
  jand g17047(.dina(n17160), .dinb(n17152), .dout(n17303));
  jor  g17048(.dina(n17303), .dinb(n17302), .dout(n17304));
  jand g17049(.dina(n10594), .dinb(b30 ), .dout(n17305));
  jand g17050(.dina(n10129), .dinb(b31 ), .dout(n17306));
  jor  g17051(.dina(n17306), .dinb(n17305), .dout(n17307));
  jnot g17052(.din(n17307), .dout(n17308));
  jand g17053(.dina(n17149), .dinb(n2468), .dout(n17309));
  jand g17054(.dina(n17150), .dinb(n16983), .dout(n17310));
  jor  g17055(.dina(n17310), .dinb(n17309), .dout(n17311));
  jxor g17056(.dina(n17311), .dinb(n17308), .dout(n17312));
  jor  g17057(.dina(n10134), .dinb(n3520), .dout(n17313));
  jor  g17058(.dina(n9849), .dinb(n3186), .dout(n17314));
  jor  g17059(.dina(n10137), .dinb(n3348), .dout(n17315));
  jor  g17060(.dina(n10132), .dinb(n3522), .dout(n17316));
  jand g17061(.dina(n17316), .dinb(n17315), .dout(n17317));
  jand g17062(.dina(n17317), .dinb(n17314), .dout(n17318));
  jand g17063(.dina(n17318), .dinb(n17313), .dout(n17319));
  jxor g17064(.dina(n17319), .dinb(n9559), .dout(n17320));
  jxor g17065(.dina(n17320), .dinb(n17312), .dout(n17321));
  jxor g17066(.dina(n17321), .dinb(n17304), .dout(n17322));
  jor  g17067(.dina(n9271), .dinb(n4058), .dout(n17323));
  jor  g17068(.dina(n9003), .dinb(n3698), .dout(n17324));
  jor  g17069(.dina(n9268), .dinb(n4060), .dout(n17325));
  jor  g17070(.dina(n9273), .dinb(n3873), .dout(n17326));
  jand g17071(.dina(n17326), .dinb(n17325), .dout(n17327));
  jand g17072(.dina(n17327), .dinb(n17324), .dout(n17328));
  jand g17073(.dina(n17328), .dinb(n17323), .dout(n17329));
  jxor g17074(.dina(n17329), .dinb(n8729), .dout(n17330));
  jxor g17075(.dina(n17330), .dinb(n17322), .dout(n17331));
  jxor g17076(.dina(n17331), .dinb(n17301), .dout(n17332));
  jor  g17077(.dina(n8457), .dinb(n4635), .dout(n17333));
  jor  g17078(.dina(n8185), .dinb(n4249), .dout(n17334));
  jor  g17079(.dina(n8459), .dinb(n4437), .dout(n17335));
  jor  g17080(.dina(n8454), .dinb(n4637), .dout(n17336));
  jand g17081(.dina(n17336), .dinb(n17335), .dout(n17337));
  jand g17082(.dina(n17337), .dinb(n17334), .dout(n17338));
  jand g17083(.dina(n17338), .dinb(n17333), .dout(n17339));
  jxor g17084(.dina(n17339), .dinb(n7929), .dout(n17340));
  jxor g17085(.dina(n17340), .dinb(n17332), .dout(n17341));
  jxor g17086(.dina(n17341), .dinb(n17298), .dout(n17342));
  jor  g17087(.dina(n7660), .dinb(n5251), .dout(n17343));
  jor  g17088(.dina(n7415), .dinb(n4839), .dout(n17344));
  jor  g17089(.dina(n7662), .dinb(n5253), .dout(n17345));
  jor  g17090(.dina(n7657), .dinb(n5040), .dout(n17346));
  jand g17091(.dina(n17346), .dinb(n17345), .dout(n17347));
  jand g17092(.dina(n17347), .dinb(n17344), .dout(n17348));
  jand g17093(.dina(n17348), .dinb(n17343), .dout(n17349));
  jxor g17094(.dina(n17349), .dinb(n7166), .dout(n17350));
  jxor g17095(.dina(n17350), .dinb(n17342), .dout(n17351));
  jxor g17096(.dina(n17351), .dinb(n17295), .dout(n17352));
  jor  g17097(.dina(n6914), .dinb(n5909), .dout(n17353));
  jor  g17098(.dina(n6673), .dinb(n5469), .dout(n17354));
  jor  g17099(.dina(n6911), .dinb(n5685), .dout(n17355));
  jor  g17100(.dina(n6916), .dinb(n5911), .dout(n17356));
  jand g17101(.dina(n17356), .dinb(n17355), .dout(n17357));
  jand g17102(.dina(n17357), .dinb(n17354), .dout(n17358));
  jand g17103(.dina(n17358), .dinb(n17353), .dout(n17359));
  jxor g17104(.dina(n17359), .dinb(n6443), .dout(n17360));
  jxor g17105(.dina(n17360), .dinb(n17352), .dout(n17361));
  jxor g17106(.dina(n17361), .dinb(n17292), .dout(n17362));
  jor  g17107(.dina(n6603), .dinb(n6207), .dout(n17363));
  jor  g17108(.dina(n5975), .dinb(n6139), .dout(n17364));
  jor  g17109(.dina(n6205), .dinb(n6605), .dout(n17365));
  jor  g17110(.dina(n6210), .dinb(n6366), .dout(n17366));
  jand g17111(.dina(n17366), .dinb(n17365), .dout(n17367));
  jand g17112(.dina(n17367), .dinb(n17364), .dout(n17368));
  jand g17113(.dina(n17368), .dinb(n17363), .dout(n17369));
  jxor g17114(.dina(n17369), .dinb(n5759), .dout(n17370));
  jxor g17115(.dina(n17370), .dinb(n17362), .dout(n17371));
  jxor g17116(.dina(n17371), .dinb(n17289), .dout(n17372));
  jor  g17117(.dina(n7336), .dinb(n5537), .dout(n17373));
  jor  g17118(.dina(n5315), .dinb(n6846), .dout(n17374));
  jor  g17119(.dina(n5534), .dinb(n7086), .dout(n17375));
  jor  g17120(.dina(n5539), .dinb(n7338), .dout(n17376));
  jand g17121(.dina(n17376), .dinb(n17375), .dout(n17377));
  jand g17122(.dina(n17377), .dinb(n17374), .dout(n17378));
  jand g17123(.dina(n17378), .dinb(n17373), .dout(n17379));
  jxor g17124(.dina(n17379), .dinb(n5111), .dout(n17380));
  jxor g17125(.dina(n17380), .dinb(n17372), .dout(n17381));
  jnot g17126(.din(n17220), .dout(n17382));
  jand g17127(.dina(n17382), .dinb(n17212), .dout(n17383));
  jnot g17128(.din(n17383), .dout(n17384));
  jand g17129(.dina(n17220), .dinb(n17211), .dout(n17385));
  jor  g17130(.dina(n17385), .dinb(n17128), .dout(n17386));
  jand g17131(.dina(n17386), .dinb(n17384), .dout(n17387));
  jxor g17132(.dina(n17387), .dinb(n17381), .dout(n17388));
  jor  g17133(.dina(n8109), .dinb(n4902), .dout(n17389));
  jor  g17134(.dina(n4696), .dinb(n7590), .dout(n17390));
  jor  g17135(.dina(n4904), .dinb(n7846), .dout(n17391));
  jor  g17136(.dina(n4899), .dinb(n8111), .dout(n17392));
  jand g17137(.dina(n17392), .dinb(n17391), .dout(n17393));
  jand g17138(.dina(n17393), .dinb(n17390), .dout(n17394));
  jand g17139(.dina(n17394), .dinb(n17389), .dout(n17395));
  jxor g17140(.dina(n17395), .dinb(n4505), .dout(n17396));
  jxor g17141(.dina(n17396), .dinb(n17388), .dout(n17397));
  jxor g17142(.dina(n17397), .dinb(n17286), .dout(n17398));
  jor  g17143(.dina(n8918), .dinb(n4305), .dout(n17399));
  jor  g17144(.dina(n4116), .dinb(n8378), .dout(n17400));
  jor  g17145(.dina(n4308), .dinb(n8644), .dout(n17401));
  jor  g17146(.dina(n4303), .dinb(n8920), .dout(n17402));
  jand g17147(.dina(n17402), .dinb(n17401), .dout(n17403));
  jand g17148(.dina(n17403), .dinb(n17400), .dout(n17404));
  jand g17149(.dina(n17404), .dinb(n17399), .dout(n17405));
  jxor g17150(.dina(n17405), .dinb(n3938), .dout(n17406));
  jxor g17151(.dina(n17406), .dinb(n17398), .dout(n17407));
  jxor g17152(.dina(n17407), .dinb(n17281), .dout(n17408));
  jor  g17153(.dina(n9757), .dinb(n3751), .dout(n17409));
  jor  g17154(.dina(n3574), .dinb(n9195), .dout(n17410));
  jor  g17155(.dina(n3754), .dinb(n9475), .dout(n17411));
  jor  g17156(.dina(n3749), .dinb(n9759), .dout(n17412));
  jand g17157(.dina(n17412), .dinb(n17411), .dout(n17413));
  jand g17158(.dina(n17413), .dinb(n17410), .dout(n17414));
  jand g17159(.dina(n17414), .dinb(n17409), .dout(n17415));
  jxor g17160(.dina(n17415), .dinb(n3410), .dout(n17416));
  jxor g17161(.dina(n17416), .dinb(n17408), .dout(n17417));
  jxor g17162(.dina(n17417), .dinb(n17278), .dout(n17418));
  jxor g17163(.dina(n17418), .dinb(n17267), .dout(n17419));
  jnot g17164(.din(n17419), .dout(n17420));
  jxor g17165(.dina(n17420), .dinb(n17264), .dout(f94 ));
  jand g17166(.dina(n17418), .dinb(n17267), .dout(n17422));
  jnot g17167(.din(n17422), .dout(n17423));
  jor  g17168(.dina(n17420), .dinb(n17264), .dout(n17424));
  jand g17169(.dina(n17424), .dinb(n17423), .dout(n17425));
  jor  g17170(.dina(n17277), .dinb(n17271), .dout(n17426));
  jand g17171(.dina(n17417), .dinb(n17278), .dout(n17427));
  jnot g17172(.din(n17427), .dout(n17428));
  jand g17173(.dina(n17428), .dinb(n17426), .dout(n17429));
  jnot g17174(.din(n17429), .dout(n17430));
  jand g17175(.dina(n17407), .dinb(n17281), .dout(n17431));
  jand g17176(.dina(n17416), .dinb(n17408), .dout(n17432));
  jor  g17177(.dina(n17432), .dinb(n17431), .dout(n17433));
  jnot g17178(.din(n17433), .dout(n17434));
  jand g17179(.dina(n3073), .dinb(b63 ), .dout(n17435));
  jand g17180(.dina(n10832), .dinb(n2907), .dout(n17436));
  jor  g17181(.dina(n17436), .dinb(n17435), .dout(n17437));
  jxor g17182(.dina(n17437), .dinb(n2918), .dout(n17438));
  jxor g17183(.dina(n17438), .dinb(n17434), .dout(n17439));
  jand g17184(.dina(n17397), .dinb(n17286), .dout(n17440));
  jand g17185(.dina(n17406), .dinb(n17398), .dout(n17441));
  jor  g17186(.dina(n17441), .dinb(n17440), .dout(n17442));
  jand g17187(.dina(n17387), .dinb(n17381), .dout(n17443));
  jand g17188(.dina(n17396), .dinb(n17388), .dout(n17444));
  jor  g17189(.dina(n17444), .dinb(n17443), .dout(n17445));
  jand g17190(.dina(n17371), .dinb(n17289), .dout(n17446));
  jand g17191(.dina(n17380), .dinb(n17372), .dout(n17447));
  jor  g17192(.dina(n17447), .dinb(n17446), .dout(n17448));
  jand g17193(.dina(n17361), .dinb(n17292), .dout(n17449));
  jand g17194(.dina(n17370), .dinb(n17362), .dout(n17450));
  jor  g17195(.dina(n17450), .dinb(n17449), .dout(n17451));
  jand g17196(.dina(n17351), .dinb(n17295), .dout(n17452));
  jand g17197(.dina(n17360), .dinb(n17352), .dout(n17453));
  jor  g17198(.dina(n17453), .dinb(n17452), .dout(n17454));
  jand g17199(.dina(n17341), .dinb(n17298), .dout(n17455));
  jand g17200(.dina(n17350), .dinb(n17342), .dout(n17456));
  jor  g17201(.dina(n17456), .dinb(n17455), .dout(n17457));
  jand g17202(.dina(n17331), .dinb(n17301), .dout(n17458));
  jand g17203(.dina(n17340), .dinb(n17332), .dout(n17459));
  jor  g17204(.dina(n17459), .dinb(n17458), .dout(n17460));
  jand g17205(.dina(n17321), .dinb(n17304), .dout(n17461));
  jand g17206(.dina(n17330), .dinb(n17322), .dout(n17462));
  jor  g17207(.dina(n17462), .dinb(n17461), .dout(n17463));
  jand g17208(.dina(n17311), .dinb(n17308), .dout(n17464));
  jand g17209(.dina(n17320), .dinb(n17312), .dout(n17465));
  jor  g17210(.dina(n17465), .dinb(n17464), .dout(n17466));
  jand g17211(.dina(n10594), .dinb(b31 ), .dout(n17467));
  jand g17212(.dina(n10129), .dinb(b32 ), .dout(n17468));
  jor  g17213(.dina(n17468), .dinb(n17467), .dout(n17469));
  jnot g17214(.din(n17469), .dout(n17470));
  jxor g17215(.dina(n17470), .dinb(n17307), .dout(n17471));
  jxor g17216(.dina(n17471), .dinb(n17466), .dout(n17472));
  jor  g17217(.dina(n10134), .dinb(n3696), .dout(n17473));
  jor  g17218(.dina(n9849), .dinb(n3348), .dout(n17474));
  jor  g17219(.dina(n10137), .dinb(n3522), .dout(n17475));
  jor  g17220(.dina(n10132), .dinb(n3698), .dout(n17476));
  jand g17221(.dina(n17476), .dinb(n17475), .dout(n17477));
  jand g17222(.dina(n17477), .dinb(n17474), .dout(n17478));
  jand g17223(.dina(n17478), .dinb(n17473), .dout(n17479));
  jxor g17224(.dina(n17479), .dinb(n9559), .dout(n17480));
  jxor g17225(.dina(n17480), .dinb(n17472), .dout(n17481));
  jor  g17226(.dina(n9271), .dinb(n4247), .dout(n17482));
  jor  g17227(.dina(n9003), .dinb(n3873), .dout(n17483));
  jor  g17228(.dina(n9273), .dinb(n4060), .dout(n17484));
  jor  g17229(.dina(n9268), .dinb(n4249), .dout(n17485));
  jand g17230(.dina(n17485), .dinb(n17484), .dout(n17486));
  jand g17231(.dina(n17486), .dinb(n17483), .dout(n17487));
  jand g17232(.dina(n17487), .dinb(n17482), .dout(n17488));
  jxor g17233(.dina(n17488), .dinb(n8729), .dout(n17489));
  jxor g17234(.dina(n17489), .dinb(n17481), .dout(n17490));
  jxor g17235(.dina(n17490), .dinb(n17463), .dout(n17491));
  jor  g17236(.dina(n8457), .dinb(n4837), .dout(n17492));
  jor  g17237(.dina(n8185), .dinb(n4437), .dout(n17493));
  jor  g17238(.dina(n8454), .dinb(n4839), .dout(n17494));
  jor  g17239(.dina(n8459), .dinb(n4637), .dout(n17495));
  jand g17240(.dina(n17495), .dinb(n17494), .dout(n17496));
  jand g17241(.dina(n17496), .dinb(n17493), .dout(n17497));
  jand g17242(.dina(n17497), .dinb(n17492), .dout(n17498));
  jxor g17243(.dina(n17498), .dinb(n7929), .dout(n17499));
  jxor g17244(.dina(n17499), .dinb(n17491), .dout(n17500));
  jxor g17245(.dina(n17500), .dinb(n17460), .dout(n17501));
  jor  g17246(.dina(n7660), .dinb(n5467), .dout(n17502));
  jor  g17247(.dina(n7415), .dinb(n5040), .dout(n17503));
  jor  g17248(.dina(n7657), .dinb(n5253), .dout(n17504));
  jor  g17249(.dina(n7662), .dinb(n5469), .dout(n17505));
  jand g17250(.dina(n17505), .dinb(n17504), .dout(n17506));
  jand g17251(.dina(n17506), .dinb(n17503), .dout(n17507));
  jand g17252(.dina(n17507), .dinb(n17502), .dout(n17508));
  jxor g17253(.dina(n17508), .dinb(n7166), .dout(n17509));
  jxor g17254(.dina(n17509), .dinb(n17501), .dout(n17510));
  jxor g17255(.dina(n17510), .dinb(n17457), .dout(n17511));
  jor  g17256(.dina(n6914), .dinb(n6137), .dout(n17512));
  jor  g17257(.dina(n6673), .dinb(n5685), .dout(n17513));
  jor  g17258(.dina(n6911), .dinb(n5911), .dout(n17514));
  jor  g17259(.dina(n6916), .dinb(n6139), .dout(n17515));
  jand g17260(.dina(n17515), .dinb(n17514), .dout(n17516));
  jand g17261(.dina(n17516), .dinb(n17513), .dout(n17517));
  jand g17262(.dina(n17517), .dinb(n17512), .dout(n17518));
  jxor g17263(.dina(n17518), .dinb(n6443), .dout(n17519));
  jxor g17264(.dina(n17519), .dinb(n17511), .dout(n17520));
  jxor g17265(.dina(n17520), .dinb(n17454), .dout(n17521));
  jor  g17266(.dina(n6844), .dinb(n6207), .dout(n17522));
  jor  g17267(.dina(n5975), .dinb(n6366), .dout(n17523));
  jor  g17268(.dina(n6210), .dinb(n6605), .dout(n17524));
  jor  g17269(.dina(n6205), .dinb(n6846), .dout(n17525));
  jand g17270(.dina(n17525), .dinb(n17524), .dout(n17526));
  jand g17271(.dina(n17526), .dinb(n17523), .dout(n17527));
  jand g17272(.dina(n17527), .dinb(n17522), .dout(n17528));
  jxor g17273(.dina(n17528), .dinb(n5759), .dout(n17529));
  jxor g17274(.dina(n17529), .dinb(n17521), .dout(n17530));
  jxor g17275(.dina(n17530), .dinb(n17451), .dout(n17531));
  jor  g17276(.dina(n7588), .dinb(n5537), .dout(n17532));
  jor  g17277(.dina(n5315), .dinb(n7086), .dout(n17533));
  jor  g17278(.dina(n5534), .dinb(n7338), .dout(n17534));
  jor  g17279(.dina(n5539), .dinb(n7590), .dout(n17535));
  jand g17280(.dina(n17535), .dinb(n17534), .dout(n17536));
  jand g17281(.dina(n17536), .dinb(n17533), .dout(n17537));
  jand g17282(.dina(n17537), .dinb(n17532), .dout(n17538));
  jxor g17283(.dina(n17538), .dinb(n5111), .dout(n17539));
  jxor g17284(.dina(n17539), .dinb(n17531), .dout(n17540));
  jxor g17285(.dina(n17540), .dinb(n17448), .dout(n17541));
  jor  g17286(.dina(n8376), .dinb(n4902), .dout(n17542));
  jor  g17287(.dina(n4696), .dinb(n7846), .dout(n17543));
  jor  g17288(.dina(n4904), .dinb(n8111), .dout(n17544));
  jor  g17289(.dina(n4899), .dinb(n8378), .dout(n17545));
  jand g17290(.dina(n17545), .dinb(n17544), .dout(n17546));
  jand g17291(.dina(n17546), .dinb(n17543), .dout(n17547));
  jand g17292(.dina(n17547), .dinb(n17542), .dout(n17548));
  jxor g17293(.dina(n17548), .dinb(n4505), .dout(n17549));
  jxor g17294(.dina(n17549), .dinb(n17541), .dout(n17550));
  jxor g17295(.dina(n17550), .dinb(n17445), .dout(n17551));
  jor  g17296(.dina(n9193), .dinb(n4305), .dout(n17552));
  jor  g17297(.dina(n4116), .dinb(n8644), .dout(n17553));
  jor  g17298(.dina(n4308), .dinb(n8920), .dout(n17554));
  jor  g17299(.dina(n4303), .dinb(n9195), .dout(n17555));
  jand g17300(.dina(n17555), .dinb(n17554), .dout(n17556));
  jand g17301(.dina(n17556), .dinb(n17553), .dout(n17557));
  jand g17302(.dina(n17557), .dinb(n17552), .dout(n17558));
  jxor g17303(.dina(n17558), .dinb(n3938), .dout(n17559));
  jxor g17304(.dina(n17559), .dinb(n17551), .dout(n17560));
  jxor g17305(.dina(n17560), .dinb(n17442), .dout(n17561));
  jor  g17306(.dina(n10049), .dinb(n3751), .dout(n17562));
  jor  g17307(.dina(n3574), .dinb(n9475), .dout(n17563));
  jor  g17308(.dina(n3754), .dinb(n9759), .dout(n17564));
  jor  g17309(.dina(n3749), .dinb(n10051), .dout(n17565));
  jand g17310(.dina(n17565), .dinb(n17564), .dout(n17566));
  jand g17311(.dina(n17566), .dinb(n17563), .dout(n17567));
  jand g17312(.dina(n17567), .dinb(n17562), .dout(n17568));
  jxor g17313(.dina(n17568), .dinb(n3410), .dout(n17569));
  jxor g17314(.dina(n17569), .dinb(n17561), .dout(n17570));
  jxor g17315(.dina(n17570), .dinb(n17439), .dout(n17571));
  jxor g17316(.dina(n17571), .dinb(n17430), .dout(n17572));
  jnot g17317(.din(n17572), .dout(n17573));
  jxor g17318(.dina(n17573), .dinb(n17425), .dout(f95 ));
  jand g17319(.dina(n17571), .dinb(n17430), .dout(n17575));
  jnot g17320(.din(n17575), .dout(n17576));
  jor  g17321(.dina(n17573), .dinb(n17425), .dout(n17577));
  jand g17322(.dina(n17577), .dinb(n17576), .dout(n17578));
  jor  g17323(.dina(n17438), .dinb(n17434), .dout(n17579));
  jand g17324(.dina(n17570), .dinb(n17439), .dout(n17580));
  jnot g17325(.din(n17580), .dout(n17581));
  jand g17326(.dina(n17581), .dinb(n17579), .dout(n17582));
  jnot g17327(.din(n17582), .dout(n17583));
  jand g17328(.dina(n17550), .dinb(n17445), .dout(n17584));
  jand g17329(.dina(n17559), .dinb(n17551), .dout(n17585));
  jor  g17330(.dina(n17585), .dinb(n17584), .dout(n17586));
  jand g17331(.dina(n17540), .dinb(n17448), .dout(n17587));
  jand g17332(.dina(n17549), .dinb(n17541), .dout(n17588));
  jor  g17333(.dina(n17588), .dinb(n17587), .dout(n17589));
  jand g17334(.dina(n17530), .dinb(n17451), .dout(n17590));
  jand g17335(.dina(n17539), .dinb(n17531), .dout(n17591));
  jor  g17336(.dina(n17591), .dinb(n17590), .dout(n17592));
  jor  g17337(.dina(n7844), .dinb(n5537), .dout(n17593));
  jor  g17338(.dina(n5315), .dinb(n7338), .dout(n17594));
  jor  g17339(.dina(n5534), .dinb(n7590), .dout(n17595));
  jor  g17340(.dina(n5539), .dinb(n7846), .dout(n17596));
  jand g17341(.dina(n17596), .dinb(n17595), .dout(n17597));
  jand g17342(.dina(n17597), .dinb(n17594), .dout(n17598));
  jand g17343(.dina(n17598), .dinb(n17593), .dout(n17599));
  jxor g17344(.dina(n17599), .dinb(n5111), .dout(n17600));
  jnot g17345(.din(n17600), .dout(n17601));
  jand g17346(.dina(n17520), .dinb(n17454), .dout(n17602));
  jand g17347(.dina(n17529), .dinb(n17521), .dout(n17603));
  jor  g17348(.dina(n17603), .dinb(n17602), .dout(n17604));
  jand g17349(.dina(n17510), .dinb(n17457), .dout(n17605));
  jand g17350(.dina(n17519), .dinb(n17511), .dout(n17606));
  jor  g17351(.dina(n17606), .dinb(n17605), .dout(n17607));
  jand g17352(.dina(n17500), .dinb(n17460), .dout(n17608));
  jand g17353(.dina(n17509), .dinb(n17501), .dout(n17609));
  jor  g17354(.dina(n17609), .dinb(n17608), .dout(n17610));
  jand g17355(.dina(n17490), .dinb(n17463), .dout(n17611));
  jand g17356(.dina(n17499), .dinb(n17491), .dout(n17612));
  jor  g17357(.dina(n17612), .dinb(n17611), .dout(n17613));
  jand g17358(.dina(n17480), .dinb(n17472), .dout(n17614));
  jand g17359(.dina(n17489), .dinb(n17481), .dout(n17615));
  jor  g17360(.dina(n17615), .dinb(n17614), .dout(n17616));
  jand g17361(.dina(n17470), .dinb(n17307), .dout(n17617));
  jand g17362(.dina(n17471), .dinb(n17466), .dout(n17618));
  jor  g17363(.dina(n17618), .dinb(n17617), .dout(n17619));
  jand g17364(.dina(n10594), .dinb(b32 ), .dout(n17620));
  jand g17365(.dina(n10129), .dinb(b33 ), .dout(n17621));
  jor  g17366(.dina(n17621), .dinb(n17620), .dout(n17622));
  jxor g17367(.dina(n17622), .dinb(n2918), .dout(n17623));
  jxor g17368(.dina(n17623), .dinb(n17469), .dout(n17624));
  jxor g17369(.dina(n17624), .dinb(n17619), .dout(n17625));
  jor  g17370(.dina(n10134), .dinb(n3871), .dout(n17626));
  jor  g17371(.dina(n9849), .dinb(n3522), .dout(n17627));
  jor  g17372(.dina(n10137), .dinb(n3698), .dout(n17628));
  jor  g17373(.dina(n10132), .dinb(n3873), .dout(n17629));
  jand g17374(.dina(n17629), .dinb(n17628), .dout(n17630));
  jand g17375(.dina(n17630), .dinb(n17627), .dout(n17631));
  jand g17376(.dina(n17631), .dinb(n17626), .dout(n17632));
  jxor g17377(.dina(n17632), .dinb(n9559), .dout(n17633));
  jxor g17378(.dina(n17633), .dinb(n17625), .dout(n17634));
  jor  g17379(.dina(n9271), .dinb(n4435), .dout(n17635));
  jor  g17380(.dina(n9003), .dinb(n4060), .dout(n17636));
  jor  g17381(.dina(n9273), .dinb(n4249), .dout(n17637));
  jor  g17382(.dina(n9268), .dinb(n4437), .dout(n17638));
  jand g17383(.dina(n17638), .dinb(n17637), .dout(n17639));
  jand g17384(.dina(n17639), .dinb(n17636), .dout(n17640));
  jand g17385(.dina(n17640), .dinb(n17635), .dout(n17641));
  jxor g17386(.dina(n17641), .dinb(n8729), .dout(n17642));
  jxor g17387(.dina(n17642), .dinb(n17634), .dout(n17643));
  jxor g17388(.dina(n17643), .dinb(n17616), .dout(n17644));
  jor  g17389(.dina(n8457), .dinb(n5038), .dout(n17645));
  jor  g17390(.dina(n8185), .dinb(n4637), .dout(n17646));
  jor  g17391(.dina(n8459), .dinb(n4839), .dout(n17647));
  jor  g17392(.dina(n8454), .dinb(n5040), .dout(n17648));
  jand g17393(.dina(n17648), .dinb(n17647), .dout(n17649));
  jand g17394(.dina(n17649), .dinb(n17646), .dout(n17650));
  jand g17395(.dina(n17650), .dinb(n17645), .dout(n17651));
  jxor g17396(.dina(n17651), .dinb(n7929), .dout(n17652));
  jxor g17397(.dina(n17652), .dinb(n17644), .dout(n17653));
  jxor g17398(.dina(n17653), .dinb(n17613), .dout(n17654));
  jor  g17399(.dina(n7660), .dinb(n5683), .dout(n17655));
  jor  g17400(.dina(n7415), .dinb(n5253), .dout(n17656));
  jor  g17401(.dina(n7657), .dinb(n5469), .dout(n17657));
  jor  g17402(.dina(n7662), .dinb(n5685), .dout(n17658));
  jand g17403(.dina(n17658), .dinb(n17657), .dout(n17659));
  jand g17404(.dina(n17659), .dinb(n17656), .dout(n17660));
  jand g17405(.dina(n17660), .dinb(n17655), .dout(n17661));
  jxor g17406(.dina(n17661), .dinb(n7166), .dout(n17662));
  jxor g17407(.dina(n17662), .dinb(n17654), .dout(n17663));
  jxor g17408(.dina(n17663), .dinb(n17610), .dout(n17664));
  jor  g17409(.dina(n6914), .dinb(n6364), .dout(n17665));
  jor  g17410(.dina(n6673), .dinb(n5911), .dout(n17666));
  jor  g17411(.dina(n6916), .dinb(n6366), .dout(n17667));
  jor  g17412(.dina(n6911), .dinb(n6139), .dout(n17668));
  jand g17413(.dina(n17668), .dinb(n17667), .dout(n17669));
  jand g17414(.dina(n17669), .dinb(n17666), .dout(n17670));
  jand g17415(.dina(n17670), .dinb(n17665), .dout(n17671));
  jxor g17416(.dina(n17671), .dinb(n6443), .dout(n17672));
  jxor g17417(.dina(n17672), .dinb(n17664), .dout(n17673));
  jxor g17418(.dina(n17673), .dinb(n17607), .dout(n17674));
  jnot g17419(.din(n17674), .dout(n17675));
  jor  g17420(.dina(n7084), .dinb(n6207), .dout(n17676));
  jor  g17421(.dina(n5975), .dinb(n6605), .dout(n17677));
  jor  g17422(.dina(n6210), .dinb(n6846), .dout(n17678));
  jor  g17423(.dina(n6205), .dinb(n7086), .dout(n17679));
  jand g17424(.dina(n17679), .dinb(n17678), .dout(n17680));
  jand g17425(.dina(n17680), .dinb(n17677), .dout(n17681));
  jand g17426(.dina(n17681), .dinb(n17676), .dout(n17682));
  jxor g17427(.dina(n17682), .dinb(n5759), .dout(n17683));
  jxor g17428(.dina(n17683), .dinb(n17675), .dout(n17684));
  jxor g17429(.dina(n17684), .dinb(n17604), .dout(n17685));
  jxor g17430(.dina(n17685), .dinb(n17601), .dout(n17686));
  jxor g17431(.dina(n17686), .dinb(n17592), .dout(n17687));
  jor  g17432(.dina(n8642), .dinb(n4902), .dout(n17688));
  jor  g17433(.dina(n4696), .dinb(n8111), .dout(n17689));
  jor  g17434(.dina(n4904), .dinb(n8378), .dout(n17690));
  jor  g17435(.dina(n4899), .dinb(n8644), .dout(n17691));
  jand g17436(.dina(n17691), .dinb(n17690), .dout(n17692));
  jand g17437(.dina(n17692), .dinb(n17689), .dout(n17693));
  jand g17438(.dina(n17693), .dinb(n17688), .dout(n17694));
  jxor g17439(.dina(n17694), .dinb(n4505), .dout(n17695));
  jxor g17440(.dina(n17695), .dinb(n17687), .dout(n17696));
  jxor g17441(.dina(n17696), .dinb(n17589), .dout(n17697));
  jor  g17442(.dina(n9473), .dinb(n4305), .dout(n17698));
  jor  g17443(.dina(n4116), .dinb(n8920), .dout(n17699));
  jor  g17444(.dina(n4308), .dinb(n9195), .dout(n17700));
  jor  g17445(.dina(n4303), .dinb(n9475), .dout(n17701));
  jand g17446(.dina(n17701), .dinb(n17700), .dout(n17702));
  jand g17447(.dina(n17702), .dinb(n17699), .dout(n17703));
  jand g17448(.dina(n17703), .dinb(n17698), .dout(n17704));
  jxor g17449(.dina(n17704), .dinb(n3938), .dout(n17705));
  jxor g17450(.dina(n17705), .dinb(n17697), .dout(n17706));
  jxor g17451(.dina(n17706), .dinb(n17586), .dout(n17707));
  jand g17452(.dina(n17560), .dinb(n17442), .dout(n17708));
  jand g17453(.dina(n17569), .dinb(n17561), .dout(n17709));
  jor  g17454(.dina(n17709), .dinb(n17708), .dout(n17710));
  jor  g17455(.dina(n10521), .dinb(n3751), .dout(n17711));
  jor  g17456(.dina(n3574), .dinb(n9759), .dout(n17712));
  jor  g17457(.dina(n3749), .dinb(n10523), .dout(n17713));
  jor  g17458(.dina(n3754), .dinb(n10051), .dout(n17714));
  jand g17459(.dina(n17714), .dinb(n17713), .dout(n17715));
  jand g17460(.dina(n17715), .dinb(n17712), .dout(n17716));
  jand g17461(.dina(n17716), .dinb(n17711), .dout(n17717));
  jxor g17462(.dina(n17717), .dinb(n3410), .dout(n17718));
  jxor g17463(.dina(n17718), .dinb(n17710), .dout(n17719));
  jxor g17464(.dina(n17719), .dinb(n17707), .dout(n17720));
  jxor g17465(.dina(n17720), .dinb(n17583), .dout(n17721));
  jnot g17466(.din(n17721), .dout(n17722));
  jxor g17467(.dina(n17722), .dinb(n17578), .dout(f96 ));
  jand g17468(.dina(n17720), .dinb(n17583), .dout(n17724));
  jnot g17469(.din(n17724), .dout(n17725));
  jor  g17470(.dina(n17722), .dinb(n17578), .dout(n17726));
  jand g17471(.dina(n17726), .dinb(n17725), .dout(n17727));
  jand g17472(.dina(n17718), .dinb(n17710), .dout(n17728));
  jand g17473(.dina(n17719), .dinb(n17707), .dout(n17729));
  jor  g17474(.dina(n17729), .dinb(n17728), .dout(n17730));
  jand g17475(.dina(n17705), .dinb(n17697), .dout(n17731));
  jand g17476(.dina(n17706), .dinb(n17586), .dout(n17732));
  jor  g17477(.dina(n17732), .dinb(n17731), .dout(n17733));
  jnot g17478(.din(n17733), .dout(n17734));
  jor  g17479(.dina(n3754), .dinb(n10523), .dout(n17735));
  jor  g17480(.dina(n10813), .dinb(n3751), .dout(n17736));
  jor  g17481(.dina(n3574), .dinb(n10051), .dout(n17737));
  jand g17482(.dina(n17737), .dinb(n17736), .dout(n17738));
  jand g17483(.dina(n17738), .dinb(n17735), .dout(n17739));
  jxor g17484(.dina(n17739), .dinb(a35 ), .dout(n17740));
  jxor g17485(.dina(n17740), .dinb(n17734), .dout(n17741));
  jand g17486(.dina(n17695), .dinb(n17687), .dout(n17742));
  jand g17487(.dina(n17696), .dinb(n17589), .dout(n17743));
  jor  g17488(.dina(n17743), .dinb(n17742), .dout(n17744));
  jor  g17489(.dina(n17685), .dinb(n17601), .dout(n17745));
  jand g17490(.dina(n17686), .dinb(n17592), .dout(n17746));
  jnot g17491(.din(n17746), .dout(n17747));
  jand g17492(.dina(n17747), .dinb(n17745), .dout(n17748));
  jnot g17493(.din(n17748), .dout(n17749));
  jand g17494(.dina(n17672), .dinb(n17664), .dout(n17750));
  jand g17495(.dina(n17673), .dinb(n17607), .dout(n17751));
  jor  g17496(.dina(n17751), .dinb(n17750), .dout(n17752));
  jand g17497(.dina(n17662), .dinb(n17654), .dout(n17753));
  jand g17498(.dina(n17663), .dinb(n17610), .dout(n17754));
  jor  g17499(.dina(n17754), .dinb(n17753), .dout(n17755));
  jand g17500(.dina(n17652), .dinb(n17644), .dout(n17756));
  jand g17501(.dina(n17653), .dinb(n17613), .dout(n17757));
  jor  g17502(.dina(n17757), .dinb(n17756), .dout(n17758));
  jand g17503(.dina(n17642), .dinb(n17634), .dout(n17759));
  jand g17504(.dina(n17643), .dinb(n17616), .dout(n17760));
  jor  g17505(.dina(n17760), .dinb(n17759), .dout(n17761));
  jand g17506(.dina(n17624), .dinb(n17619), .dout(n17762));
  jand g17507(.dina(n17633), .dinb(n17625), .dout(n17763));
  jor  g17508(.dina(n17763), .dinb(n17762), .dout(n17764));
  jand g17509(.dina(n10594), .dinb(b33 ), .dout(n17765));
  jand g17510(.dina(n10129), .dinb(b34 ), .dout(n17766));
  jor  g17511(.dina(n17766), .dinb(n17765), .dout(n17767));
  jnot g17512(.din(n17767), .dout(n17768));
  jand g17513(.dina(n17622), .dinb(n2918), .dout(n17769));
  jand g17514(.dina(n17623), .dinb(n17469), .dout(n17770));
  jor  g17515(.dina(n17770), .dinb(n17769), .dout(n17771));
  jxor g17516(.dina(n17771), .dinb(n17768), .dout(n17772));
  jor  g17517(.dina(n10134), .dinb(n4058), .dout(n17773));
  jor  g17518(.dina(n9849), .dinb(n3698), .dout(n17774));
  jor  g17519(.dina(n10132), .dinb(n4060), .dout(n17775));
  jor  g17520(.dina(n10137), .dinb(n3873), .dout(n17776));
  jand g17521(.dina(n17776), .dinb(n17775), .dout(n17777));
  jand g17522(.dina(n17777), .dinb(n17774), .dout(n17778));
  jand g17523(.dina(n17778), .dinb(n17773), .dout(n17779));
  jxor g17524(.dina(n17779), .dinb(n9559), .dout(n17780));
  jxor g17525(.dina(n17780), .dinb(n17772), .dout(n17781));
  jxor g17526(.dina(n17781), .dinb(n17764), .dout(n17782));
  jor  g17527(.dina(n9271), .dinb(n4635), .dout(n17783));
  jor  g17528(.dina(n9003), .dinb(n4249), .dout(n17784));
  jor  g17529(.dina(n9273), .dinb(n4437), .dout(n17785));
  jor  g17530(.dina(n9268), .dinb(n4637), .dout(n17786));
  jand g17531(.dina(n17786), .dinb(n17785), .dout(n17787));
  jand g17532(.dina(n17787), .dinb(n17784), .dout(n17788));
  jand g17533(.dina(n17788), .dinb(n17783), .dout(n17789));
  jxor g17534(.dina(n17789), .dinb(n8729), .dout(n17790));
  jxor g17535(.dina(n17790), .dinb(n17782), .dout(n17791));
  jxor g17536(.dina(n17791), .dinb(n17761), .dout(n17792));
  jor  g17537(.dina(n8457), .dinb(n5251), .dout(n17793));
  jor  g17538(.dina(n8185), .dinb(n4839), .dout(n17794));
  jor  g17539(.dina(n8454), .dinb(n5253), .dout(n17795));
  jor  g17540(.dina(n8459), .dinb(n5040), .dout(n17796));
  jand g17541(.dina(n17796), .dinb(n17795), .dout(n17797));
  jand g17542(.dina(n17797), .dinb(n17794), .dout(n17798));
  jand g17543(.dina(n17798), .dinb(n17793), .dout(n17799));
  jxor g17544(.dina(n17799), .dinb(n7929), .dout(n17800));
  jxor g17545(.dina(n17800), .dinb(n17792), .dout(n17801));
  jxor g17546(.dina(n17801), .dinb(n17758), .dout(n17802));
  jor  g17547(.dina(n7660), .dinb(n5909), .dout(n17803));
  jor  g17548(.dina(n7415), .dinb(n5469), .dout(n17804));
  jor  g17549(.dina(n7662), .dinb(n5911), .dout(n17805));
  jor  g17550(.dina(n7657), .dinb(n5685), .dout(n17806));
  jand g17551(.dina(n17806), .dinb(n17805), .dout(n17807));
  jand g17552(.dina(n17807), .dinb(n17804), .dout(n17808));
  jand g17553(.dina(n17808), .dinb(n17803), .dout(n17809));
  jxor g17554(.dina(n17809), .dinb(n7166), .dout(n17810));
  jxor g17555(.dina(n17810), .dinb(n17802), .dout(n17811));
  jxor g17556(.dina(n17811), .dinb(n17755), .dout(n17812));
  jor  g17557(.dina(n6603), .dinb(n6914), .dout(n17813));
  jor  g17558(.dina(n6673), .dinb(n6139), .dout(n17814));
  jor  g17559(.dina(n6911), .dinb(n6366), .dout(n17815));
  jor  g17560(.dina(n6916), .dinb(n6605), .dout(n17816));
  jand g17561(.dina(n17816), .dinb(n17815), .dout(n17817));
  jand g17562(.dina(n17817), .dinb(n17814), .dout(n17818));
  jand g17563(.dina(n17818), .dinb(n17813), .dout(n17819));
  jxor g17564(.dina(n17819), .dinb(n6443), .dout(n17820));
  jxor g17565(.dina(n17820), .dinb(n17812), .dout(n17821));
  jxor g17566(.dina(n17821), .dinb(n17752), .dout(n17822));
  jor  g17567(.dina(n7336), .dinb(n6207), .dout(n17823));
  jor  g17568(.dina(n5975), .dinb(n6846), .dout(n17824));
  jor  g17569(.dina(n6210), .dinb(n7086), .dout(n17825));
  jor  g17570(.dina(n6205), .dinb(n7338), .dout(n17826));
  jand g17571(.dina(n17826), .dinb(n17825), .dout(n17827));
  jand g17572(.dina(n17827), .dinb(n17824), .dout(n17828));
  jand g17573(.dina(n17828), .dinb(n17823), .dout(n17829));
  jxor g17574(.dina(n17829), .dinb(n5759), .dout(n17830));
  jxor g17575(.dina(n17830), .dinb(n17822), .dout(n17831));
  jnot g17576(.din(n17683), .dout(n17832));
  jand g17577(.dina(n17832), .dinb(n17675), .dout(n17833));
  jnot g17578(.din(n17833), .dout(n17834));
  jand g17579(.dina(n17683), .dinb(n17674), .dout(n17835));
  jor  g17580(.dina(n17835), .dinb(n17604), .dout(n17836));
  jand g17581(.dina(n17836), .dinb(n17834), .dout(n17837));
  jxor g17582(.dina(n17837), .dinb(n17831), .dout(n17838));
  jor  g17583(.dina(n8109), .dinb(n5537), .dout(n17839));
  jor  g17584(.dina(n5315), .dinb(n7590), .dout(n17840));
  jor  g17585(.dina(n5539), .dinb(n8111), .dout(n17841));
  jor  g17586(.dina(n5534), .dinb(n7846), .dout(n17842));
  jand g17587(.dina(n17842), .dinb(n17841), .dout(n17843));
  jand g17588(.dina(n17843), .dinb(n17840), .dout(n17844));
  jand g17589(.dina(n17844), .dinb(n17839), .dout(n17845));
  jxor g17590(.dina(n17845), .dinb(n5111), .dout(n17846));
  jxor g17591(.dina(n17846), .dinb(n17838), .dout(n17847));
  jxor g17592(.dina(n17847), .dinb(n17749), .dout(n17848));
  jor  g17593(.dina(n8918), .dinb(n4902), .dout(n17849));
  jor  g17594(.dina(n4696), .dinb(n8378), .dout(n17850));
  jor  g17595(.dina(n4904), .dinb(n8644), .dout(n17851));
  jor  g17596(.dina(n4899), .dinb(n8920), .dout(n17852));
  jand g17597(.dina(n17852), .dinb(n17851), .dout(n17853));
  jand g17598(.dina(n17853), .dinb(n17850), .dout(n17854));
  jand g17599(.dina(n17854), .dinb(n17849), .dout(n17855));
  jxor g17600(.dina(n17855), .dinb(n4505), .dout(n17856));
  jxor g17601(.dina(n17856), .dinb(n17848), .dout(n17857));
  jxor g17602(.dina(n17857), .dinb(n17744), .dout(n17858));
  jor  g17603(.dina(n9757), .dinb(n4305), .dout(n17859));
  jor  g17604(.dina(n4116), .dinb(n9195), .dout(n17860));
  jor  g17605(.dina(n4308), .dinb(n9475), .dout(n17861));
  jor  g17606(.dina(n4303), .dinb(n9759), .dout(n17862));
  jand g17607(.dina(n17862), .dinb(n17861), .dout(n17863));
  jand g17608(.dina(n17863), .dinb(n17860), .dout(n17864));
  jand g17609(.dina(n17864), .dinb(n17859), .dout(n17865));
  jxor g17610(.dina(n17865), .dinb(n3938), .dout(n17866));
  jxor g17611(.dina(n17866), .dinb(n17858), .dout(n17867));
  jxor g17612(.dina(n17867), .dinb(n17741), .dout(n17868));
  jxor g17613(.dina(n17868), .dinb(n17730), .dout(n17869));
  jnot g17614(.din(n17869), .dout(n17870));
  jxor g17615(.dina(n17870), .dinb(n17727), .dout(f97 ));
  jand g17616(.dina(n17868), .dinb(n17730), .dout(n17872));
  jnot g17617(.din(n17872), .dout(n17873));
  jor  g17618(.dina(n17870), .dinb(n17727), .dout(n17874));
  jand g17619(.dina(n17874), .dinb(n17873), .dout(n17875));
  jor  g17620(.dina(n17740), .dinb(n17734), .dout(n17876));
  jand g17621(.dina(n17867), .dinb(n17741), .dout(n17877));
  jnot g17622(.din(n17877), .dout(n17878));
  jand g17623(.dina(n17878), .dinb(n17876), .dout(n17879));
  jnot g17624(.din(n17879), .dout(n17880));
  jand g17625(.dina(n17857), .dinb(n17744), .dout(n17881));
  jand g17626(.dina(n17866), .dinb(n17858), .dout(n17882));
  jor  g17627(.dina(n17882), .dinb(n17881), .dout(n17883));
  jnot g17628(.din(n17883), .dout(n17884));
  jand g17629(.dina(n3575), .dinb(b63 ), .dout(n17885));
  jand g17630(.dina(n10832), .dinb(n3399), .dout(n17886));
  jor  g17631(.dina(n17886), .dinb(n17885), .dout(n17887));
  jxor g17632(.dina(n17887), .dinb(n3410), .dout(n17888));
  jxor g17633(.dina(n17888), .dinb(n17884), .dout(n17889));
  jand g17634(.dina(n17847), .dinb(n17749), .dout(n17890));
  jand g17635(.dina(n17856), .dinb(n17848), .dout(n17891));
  jor  g17636(.dina(n17891), .dinb(n17890), .dout(n17892));
  jand g17637(.dina(n17837), .dinb(n17831), .dout(n17893));
  jand g17638(.dina(n17846), .dinb(n17838), .dout(n17894));
  jor  g17639(.dina(n17894), .dinb(n17893), .dout(n17895));
  jand g17640(.dina(n17821), .dinb(n17752), .dout(n17896));
  jand g17641(.dina(n17830), .dinb(n17822), .dout(n17897));
  jor  g17642(.dina(n17897), .dinb(n17896), .dout(n17898));
  jand g17643(.dina(n17811), .dinb(n17755), .dout(n17899));
  jand g17644(.dina(n17820), .dinb(n17812), .dout(n17900));
  jor  g17645(.dina(n17900), .dinb(n17899), .dout(n17901));
  jand g17646(.dina(n17801), .dinb(n17758), .dout(n17902));
  jand g17647(.dina(n17810), .dinb(n17802), .dout(n17903));
  jor  g17648(.dina(n17903), .dinb(n17902), .dout(n17904));
  jand g17649(.dina(n17791), .dinb(n17761), .dout(n17905));
  jand g17650(.dina(n17800), .dinb(n17792), .dout(n17906));
  jor  g17651(.dina(n17906), .dinb(n17905), .dout(n17907));
  jand g17652(.dina(n17781), .dinb(n17764), .dout(n17908));
  jand g17653(.dina(n17790), .dinb(n17782), .dout(n17909));
  jor  g17654(.dina(n17909), .dinb(n17908), .dout(n17910));
  jand g17655(.dina(n17771), .dinb(n17768), .dout(n17911));
  jand g17656(.dina(n17780), .dinb(n17772), .dout(n17912));
  jor  g17657(.dina(n17912), .dinb(n17911), .dout(n17913));
  jand g17658(.dina(n10594), .dinb(b34 ), .dout(n17914));
  jand g17659(.dina(n10129), .dinb(b35 ), .dout(n17915));
  jor  g17660(.dina(n17915), .dinb(n17914), .dout(n17916));
  jnot g17661(.din(n17916), .dout(n17917));
  jxor g17662(.dina(n17917), .dinb(n17767), .dout(n17918));
  jxor g17663(.dina(n17918), .dinb(n17913), .dout(n17919));
  jor  g17664(.dina(n10134), .dinb(n4247), .dout(n17920));
  jor  g17665(.dina(n9849), .dinb(n3873), .dout(n17921));
  jor  g17666(.dina(n10132), .dinb(n4249), .dout(n17922));
  jor  g17667(.dina(n10137), .dinb(n4060), .dout(n17923));
  jand g17668(.dina(n17923), .dinb(n17922), .dout(n17924));
  jand g17669(.dina(n17924), .dinb(n17921), .dout(n17925));
  jand g17670(.dina(n17925), .dinb(n17920), .dout(n17926));
  jxor g17671(.dina(n17926), .dinb(n9559), .dout(n17927));
  jxor g17672(.dina(n17927), .dinb(n17919), .dout(n17928));
  jor  g17673(.dina(n9271), .dinb(n4837), .dout(n17929));
  jor  g17674(.dina(n9003), .dinb(n4437), .dout(n17930));
  jor  g17675(.dina(n9268), .dinb(n4839), .dout(n17931));
  jor  g17676(.dina(n9273), .dinb(n4637), .dout(n17932));
  jand g17677(.dina(n17932), .dinb(n17931), .dout(n17933));
  jand g17678(.dina(n17933), .dinb(n17930), .dout(n17934));
  jand g17679(.dina(n17934), .dinb(n17929), .dout(n17935));
  jxor g17680(.dina(n17935), .dinb(n8729), .dout(n17936));
  jxor g17681(.dina(n17936), .dinb(n17928), .dout(n17937));
  jxor g17682(.dina(n17937), .dinb(n17910), .dout(n17938));
  jor  g17683(.dina(n8457), .dinb(n5467), .dout(n17939));
  jor  g17684(.dina(n8185), .dinb(n5040), .dout(n17940));
  jor  g17685(.dina(n8459), .dinb(n5253), .dout(n17941));
  jor  g17686(.dina(n8454), .dinb(n5469), .dout(n17942));
  jand g17687(.dina(n17942), .dinb(n17941), .dout(n17943));
  jand g17688(.dina(n17943), .dinb(n17940), .dout(n17944));
  jand g17689(.dina(n17944), .dinb(n17939), .dout(n17945));
  jxor g17690(.dina(n17945), .dinb(n7929), .dout(n17946));
  jxor g17691(.dina(n17946), .dinb(n17938), .dout(n17947));
  jxor g17692(.dina(n17947), .dinb(n17907), .dout(n17948));
  jor  g17693(.dina(n7660), .dinb(n6137), .dout(n17949));
  jor  g17694(.dina(n7415), .dinb(n5685), .dout(n17950));
  jor  g17695(.dina(n7657), .dinb(n5911), .dout(n17951));
  jor  g17696(.dina(n7662), .dinb(n6139), .dout(n17952));
  jand g17697(.dina(n17952), .dinb(n17951), .dout(n17953));
  jand g17698(.dina(n17953), .dinb(n17950), .dout(n17954));
  jand g17699(.dina(n17954), .dinb(n17949), .dout(n17955));
  jxor g17700(.dina(n17955), .dinb(n7166), .dout(n17956));
  jxor g17701(.dina(n17956), .dinb(n17948), .dout(n17957));
  jxor g17702(.dina(n17957), .dinb(n17904), .dout(n17958));
  jor  g17703(.dina(n6844), .dinb(n6914), .dout(n17959));
  jor  g17704(.dina(n6673), .dinb(n6366), .dout(n17960));
  jor  g17705(.dina(n6911), .dinb(n6605), .dout(n17961));
  jor  g17706(.dina(n6916), .dinb(n6846), .dout(n17962));
  jand g17707(.dina(n17962), .dinb(n17961), .dout(n17963));
  jand g17708(.dina(n17963), .dinb(n17960), .dout(n17964));
  jand g17709(.dina(n17964), .dinb(n17959), .dout(n17965));
  jxor g17710(.dina(n17965), .dinb(n6443), .dout(n17966));
  jxor g17711(.dina(n17966), .dinb(n17958), .dout(n17967));
  jxor g17712(.dina(n17967), .dinb(n17901), .dout(n17968));
  jor  g17713(.dina(n7588), .dinb(n6207), .dout(n17969));
  jor  g17714(.dina(n5975), .dinb(n7086), .dout(n17970));
  jor  g17715(.dina(n6205), .dinb(n7590), .dout(n17971));
  jor  g17716(.dina(n6210), .dinb(n7338), .dout(n17972));
  jand g17717(.dina(n17972), .dinb(n17971), .dout(n17973));
  jand g17718(.dina(n17973), .dinb(n17970), .dout(n17974));
  jand g17719(.dina(n17974), .dinb(n17969), .dout(n17975));
  jxor g17720(.dina(n17975), .dinb(n5759), .dout(n17976));
  jxor g17721(.dina(n17976), .dinb(n17968), .dout(n17977));
  jxor g17722(.dina(n17977), .dinb(n17898), .dout(n17978));
  jor  g17723(.dina(n8376), .dinb(n5537), .dout(n17979));
  jor  g17724(.dina(n5315), .dinb(n7846), .dout(n17980));
  jor  g17725(.dina(n5539), .dinb(n8378), .dout(n17981));
  jor  g17726(.dina(n5534), .dinb(n8111), .dout(n17982));
  jand g17727(.dina(n17982), .dinb(n17981), .dout(n17983));
  jand g17728(.dina(n17983), .dinb(n17980), .dout(n17984));
  jand g17729(.dina(n17984), .dinb(n17979), .dout(n17985));
  jxor g17730(.dina(n17985), .dinb(n5111), .dout(n17986));
  jxor g17731(.dina(n17986), .dinb(n17978), .dout(n17987));
  jxor g17732(.dina(n17987), .dinb(n17895), .dout(n17988));
  jor  g17733(.dina(n9193), .dinb(n4902), .dout(n17989));
  jor  g17734(.dina(n4696), .dinb(n8644), .dout(n17990));
  jor  g17735(.dina(n4899), .dinb(n9195), .dout(n17991));
  jor  g17736(.dina(n4904), .dinb(n8920), .dout(n17992));
  jand g17737(.dina(n17992), .dinb(n17991), .dout(n17993));
  jand g17738(.dina(n17993), .dinb(n17990), .dout(n17994));
  jand g17739(.dina(n17994), .dinb(n17989), .dout(n17995));
  jxor g17740(.dina(n17995), .dinb(n4505), .dout(n17996));
  jxor g17741(.dina(n17996), .dinb(n17988), .dout(n17997));
  jxor g17742(.dina(n17997), .dinb(n17892), .dout(n17998));
  jor  g17743(.dina(n10049), .dinb(n4305), .dout(n17999));
  jor  g17744(.dina(n4116), .dinb(n9475), .dout(n18000));
  jor  g17745(.dina(n4303), .dinb(n10051), .dout(n18001));
  jor  g17746(.dina(n4308), .dinb(n9759), .dout(n18002));
  jand g17747(.dina(n18002), .dinb(n18001), .dout(n18003));
  jand g17748(.dina(n18003), .dinb(n18000), .dout(n18004));
  jand g17749(.dina(n18004), .dinb(n17999), .dout(n18005));
  jxor g17750(.dina(n18005), .dinb(n3938), .dout(n18006));
  jxor g17751(.dina(n18006), .dinb(n17998), .dout(n18007));
  jxor g17752(.dina(n18007), .dinb(n17889), .dout(n18008));
  jxor g17753(.dina(n18008), .dinb(n17880), .dout(n18009));
  jnot g17754(.din(n18009), .dout(n18010));
  jxor g17755(.dina(n18010), .dinb(n17875), .dout(f98 ));
  jand g17756(.dina(n18008), .dinb(n17880), .dout(n18012));
  jnot g17757(.din(n18012), .dout(n18013));
  jor  g17758(.dina(n18010), .dinb(n17875), .dout(n18014));
  jand g17759(.dina(n18014), .dinb(n18013), .dout(n18015));
  jand g17760(.dina(n17997), .dinb(n17892), .dout(n18016));
  jand g17761(.dina(n18006), .dinb(n17998), .dout(n18017));
  jor  g17762(.dina(n18017), .dinb(n18016), .dout(n18018));
  jand g17763(.dina(n17987), .dinb(n17895), .dout(n18019));
  jand g17764(.dina(n17996), .dinb(n17988), .dout(n18020));
  jor  g17765(.dina(n18020), .dinb(n18019), .dout(n18021));
  jand g17766(.dina(n17977), .dinb(n17898), .dout(n18022));
  jand g17767(.dina(n17986), .dinb(n17978), .dout(n18023));
  jor  g17768(.dina(n18023), .dinb(n18022), .dout(n18024));
  jand g17769(.dina(n17967), .dinb(n17901), .dout(n18025));
  jand g17770(.dina(n17976), .dinb(n17968), .dout(n18026));
  jor  g17771(.dina(n18026), .dinb(n18025), .dout(n18027));
  jand g17772(.dina(n17957), .dinb(n17904), .dout(n18028));
  jand g17773(.dina(n17966), .dinb(n17958), .dout(n18029));
  jor  g17774(.dina(n18029), .dinb(n18028), .dout(n18030));
  jand g17775(.dina(n17947), .dinb(n17907), .dout(n18031));
  jand g17776(.dina(n17956), .dinb(n17948), .dout(n18032));
  jor  g17777(.dina(n18032), .dinb(n18031), .dout(n18033));
  jand g17778(.dina(n17937), .dinb(n17910), .dout(n18034));
  jand g17779(.dina(n17946), .dinb(n17938), .dout(n18035));
  jor  g17780(.dina(n18035), .dinb(n18034), .dout(n18036));
  jand g17781(.dina(n17927), .dinb(n17919), .dout(n18037));
  jand g17782(.dina(n17936), .dinb(n17928), .dout(n18038));
  jor  g17783(.dina(n18038), .dinb(n18037), .dout(n18039));
  jand g17784(.dina(n17917), .dinb(n17767), .dout(n18040));
  jand g17785(.dina(n17918), .dinb(n17913), .dout(n18041));
  jor  g17786(.dina(n18041), .dinb(n18040), .dout(n18042));
  jand g17787(.dina(n10594), .dinb(b35 ), .dout(n18043));
  jand g17788(.dina(n10129), .dinb(b36 ), .dout(n18044));
  jor  g17789(.dina(n18044), .dinb(n18043), .dout(n18045));
  jxor g17790(.dina(n17916), .dinb(n3410), .dout(n18046));
  jxor g17791(.dina(n18046), .dinb(n18045), .dout(n18047));
  jxor g17792(.dina(n18047), .dinb(n18042), .dout(n18048));
  jor  g17793(.dina(n10134), .dinb(n4435), .dout(n18049));
  jor  g17794(.dina(n9849), .dinb(n4060), .dout(n18050));
  jor  g17795(.dina(n10132), .dinb(n4437), .dout(n18051));
  jor  g17796(.dina(n10137), .dinb(n4249), .dout(n18052));
  jand g17797(.dina(n18052), .dinb(n18051), .dout(n18053));
  jand g17798(.dina(n18053), .dinb(n18050), .dout(n18054));
  jand g17799(.dina(n18054), .dinb(n18049), .dout(n18055));
  jxor g17800(.dina(n18055), .dinb(n9559), .dout(n18056));
  jxor g17801(.dina(n18056), .dinb(n18048), .dout(n18057));
  jor  g17802(.dina(n9271), .dinb(n5038), .dout(n18058));
  jor  g17803(.dina(n9003), .dinb(n4637), .dout(n18059));
  jor  g17804(.dina(n9268), .dinb(n5040), .dout(n18060));
  jor  g17805(.dina(n9273), .dinb(n4839), .dout(n18061));
  jand g17806(.dina(n18061), .dinb(n18060), .dout(n18062));
  jand g17807(.dina(n18062), .dinb(n18059), .dout(n18063));
  jand g17808(.dina(n18063), .dinb(n18058), .dout(n18064));
  jxor g17809(.dina(n18064), .dinb(n8729), .dout(n18065));
  jxor g17810(.dina(n18065), .dinb(n18057), .dout(n18066));
  jxor g17811(.dina(n18066), .dinb(n18039), .dout(n18067));
  jor  g17812(.dina(n8457), .dinb(n5683), .dout(n18068));
  jor  g17813(.dina(n8185), .dinb(n5253), .dout(n18069));
  jor  g17814(.dina(n8454), .dinb(n5685), .dout(n18070));
  jor  g17815(.dina(n8459), .dinb(n5469), .dout(n18071));
  jand g17816(.dina(n18071), .dinb(n18070), .dout(n18072));
  jand g17817(.dina(n18072), .dinb(n18069), .dout(n18073));
  jand g17818(.dina(n18073), .dinb(n18068), .dout(n18074));
  jxor g17819(.dina(n18074), .dinb(n7929), .dout(n18075));
  jxor g17820(.dina(n18075), .dinb(n18067), .dout(n18076));
  jxor g17821(.dina(n18076), .dinb(n18036), .dout(n18077));
  jor  g17822(.dina(n7660), .dinb(n6364), .dout(n18078));
  jor  g17823(.dina(n7415), .dinb(n5911), .dout(n18079));
  jor  g17824(.dina(n7657), .dinb(n6139), .dout(n18080));
  jor  g17825(.dina(n7662), .dinb(n6366), .dout(n18081));
  jand g17826(.dina(n18081), .dinb(n18080), .dout(n18082));
  jand g17827(.dina(n18082), .dinb(n18079), .dout(n18083));
  jand g17828(.dina(n18083), .dinb(n18078), .dout(n18084));
  jxor g17829(.dina(n18084), .dinb(n7166), .dout(n18085));
  jxor g17830(.dina(n18085), .dinb(n18077), .dout(n18086));
  jxor g17831(.dina(n18086), .dinb(n18033), .dout(n18087));
  jor  g17832(.dina(n7084), .dinb(n6914), .dout(n18088));
  jor  g17833(.dina(n6673), .dinb(n6605), .dout(n18089));
  jor  g17834(.dina(n6916), .dinb(n7086), .dout(n18090));
  jor  g17835(.dina(n6911), .dinb(n6846), .dout(n18091));
  jand g17836(.dina(n18091), .dinb(n18090), .dout(n18092));
  jand g17837(.dina(n18092), .dinb(n18089), .dout(n18093));
  jand g17838(.dina(n18093), .dinb(n18088), .dout(n18094));
  jxor g17839(.dina(n18094), .dinb(n6443), .dout(n18095));
  jxor g17840(.dina(n18095), .dinb(n18087), .dout(n18096));
  jxor g17841(.dina(n18096), .dinb(n18030), .dout(n18097));
  jor  g17842(.dina(n7844), .dinb(n6207), .dout(n18098));
  jor  g17843(.dina(n5975), .dinb(n7338), .dout(n18099));
  jor  g17844(.dina(n6210), .dinb(n7590), .dout(n18100));
  jor  g17845(.dina(n6205), .dinb(n7846), .dout(n18101));
  jand g17846(.dina(n18101), .dinb(n18100), .dout(n18102));
  jand g17847(.dina(n18102), .dinb(n18099), .dout(n18103));
  jand g17848(.dina(n18103), .dinb(n18098), .dout(n18104));
  jxor g17849(.dina(n18104), .dinb(n5759), .dout(n18105));
  jxor g17850(.dina(n18105), .dinb(n18097), .dout(n18106));
  jxor g17851(.dina(n18106), .dinb(n18027), .dout(n18107));
  jor  g17852(.dina(n8642), .dinb(n5537), .dout(n18108));
  jor  g17853(.dina(n5315), .dinb(n8111), .dout(n18109));
  jor  g17854(.dina(n5539), .dinb(n8644), .dout(n18110));
  jor  g17855(.dina(n5534), .dinb(n8378), .dout(n18111));
  jand g17856(.dina(n18111), .dinb(n18110), .dout(n18112));
  jand g17857(.dina(n18112), .dinb(n18109), .dout(n18113));
  jand g17858(.dina(n18113), .dinb(n18108), .dout(n18114));
  jxor g17859(.dina(n18114), .dinb(n5111), .dout(n18115));
  jxor g17860(.dina(n18115), .dinb(n18107), .dout(n18116));
  jxor g17861(.dina(n18116), .dinb(n18024), .dout(n18117));
  jor  g17862(.dina(n9473), .dinb(n4902), .dout(n18118));
  jor  g17863(.dina(n4696), .dinb(n8920), .dout(n18119));
  jor  g17864(.dina(n4904), .dinb(n9195), .dout(n18120));
  jor  g17865(.dina(n4899), .dinb(n9475), .dout(n18121));
  jand g17866(.dina(n18121), .dinb(n18120), .dout(n18122));
  jand g17867(.dina(n18122), .dinb(n18119), .dout(n18123));
  jand g17868(.dina(n18123), .dinb(n18118), .dout(n18124));
  jxor g17869(.dina(n18124), .dinb(n4505), .dout(n18125));
  jxor g17870(.dina(n18125), .dinb(n18117), .dout(n18126));
  jxor g17871(.dina(n18126), .dinb(n18021), .dout(n18127));
  jor  g17872(.dina(n10521), .dinb(n4305), .dout(n18128));
  jor  g17873(.dina(n4116), .dinb(n9759), .dout(n18129));
  jor  g17874(.dina(n4303), .dinb(n10523), .dout(n18130));
  jor  g17875(.dina(n4308), .dinb(n10051), .dout(n18131));
  jand g17876(.dina(n18131), .dinb(n18130), .dout(n18132));
  jand g17877(.dina(n18132), .dinb(n18129), .dout(n18133));
  jand g17878(.dina(n18133), .dinb(n18128), .dout(n18134));
  jxor g17879(.dina(n18134), .dinb(n3938), .dout(n18135));
  jxor g17880(.dina(n18135), .dinb(n18127), .dout(n18136));
  jxor g17881(.dina(n18136), .dinb(n18018), .dout(n18137));
  jnot g17882(.din(n18137), .dout(n18138));
  jor  g17883(.dina(n17888), .dinb(n17884), .dout(n18139));
  jand g17884(.dina(n18007), .dinb(n17889), .dout(n18140));
  jnot g17885(.din(n18140), .dout(n18141));
  jand g17886(.dina(n18141), .dinb(n18139), .dout(n18142));
  jxor g17887(.dina(n18142), .dinb(n18138), .dout(n18143));
  jnot g17888(.din(n18143), .dout(n18144));
  jxor g17889(.dina(n18144), .dinb(n18015), .dout(f99 ));
  jand g17890(.dina(n18135), .dinb(n18127), .dout(n18146));
  jand g17891(.dina(n18136), .dinb(n18018), .dout(n18147));
  jor  g17892(.dina(n18147), .dinb(n18146), .dout(n18148));
  jand g17893(.dina(n18125), .dinb(n18117), .dout(n18149));
  jand g17894(.dina(n18126), .dinb(n18021), .dout(n18150));
  jor  g17895(.dina(n18150), .dinb(n18149), .dout(n18151));
  jnot g17896(.din(n18151), .dout(n18152));
  jor  g17897(.dina(n10813), .dinb(n4305), .dout(n18153));
  jor  g17898(.dina(n4116), .dinb(n10051), .dout(n18154));
  jor  g17899(.dina(n4308), .dinb(n10523), .dout(n18155));
  jand g17900(.dina(n18155), .dinb(n18154), .dout(n18156));
  jand g17901(.dina(n18156), .dinb(n18153), .dout(n18157));
  jxor g17902(.dina(n18157), .dinb(a38 ), .dout(n18158));
  jxor g17903(.dina(n18158), .dinb(n18152), .dout(n18159));
  jand g17904(.dina(n18115), .dinb(n18107), .dout(n18160));
  jand g17905(.dina(n18116), .dinb(n18024), .dout(n18161));
  jor  g17906(.dina(n18161), .dinb(n18160), .dout(n18162));
  jand g17907(.dina(n18105), .dinb(n18097), .dout(n18163));
  jand g17908(.dina(n18106), .dinb(n18027), .dout(n18164));
  jor  g17909(.dina(n18164), .dinb(n18163), .dout(n18165));
  jand g17910(.dina(n18095), .dinb(n18087), .dout(n18166));
  jand g17911(.dina(n18096), .dinb(n18030), .dout(n18167));
  jor  g17912(.dina(n18167), .dinb(n18166), .dout(n18168));
  jand g17913(.dina(n18085), .dinb(n18077), .dout(n18169));
  jand g17914(.dina(n18086), .dinb(n18033), .dout(n18170));
  jor  g17915(.dina(n18170), .dinb(n18169), .dout(n18171));
  jand g17916(.dina(n18075), .dinb(n18067), .dout(n18172));
  jand g17917(.dina(n18076), .dinb(n18036), .dout(n18173));
  jor  g17918(.dina(n18173), .dinb(n18172), .dout(n18174));
  jand g17919(.dina(n18065), .dinb(n18057), .dout(n18175));
  jand g17920(.dina(n18066), .dinb(n18039), .dout(n18176));
  jor  g17921(.dina(n18176), .dinb(n18175), .dout(n18177));
  jand g17922(.dina(n18047), .dinb(n18042), .dout(n18178));
  jand g17923(.dina(n18056), .dinb(n18048), .dout(n18179));
  jor  g17924(.dina(n18179), .dinb(n18178), .dout(n18180));
  jand g17925(.dina(n10594), .dinb(b36 ), .dout(n18181));
  jand g17926(.dina(n10129), .dinb(b37 ), .dout(n18182));
  jor  g17927(.dina(n18182), .dinb(n18181), .dout(n18183));
  jnot g17928(.din(n18183), .dout(n18184));
  jand g17929(.dina(n17916), .dinb(n3410), .dout(n18185));
  jand g17930(.dina(n18046), .dinb(n18045), .dout(n18186));
  jor  g17931(.dina(n18186), .dinb(n18185), .dout(n18187));
  jxor g17932(.dina(n18187), .dinb(n18184), .dout(n18188));
  jor  g17933(.dina(n10134), .dinb(n4635), .dout(n18189));
  jor  g17934(.dina(n9849), .dinb(n4249), .dout(n18190));
  jor  g17935(.dina(n10132), .dinb(n4637), .dout(n18191));
  jor  g17936(.dina(n10137), .dinb(n4437), .dout(n18192));
  jand g17937(.dina(n18192), .dinb(n18191), .dout(n18193));
  jand g17938(.dina(n18193), .dinb(n18190), .dout(n18194));
  jand g17939(.dina(n18194), .dinb(n18189), .dout(n18195));
  jxor g17940(.dina(n18195), .dinb(n9559), .dout(n18196));
  jxor g17941(.dina(n18196), .dinb(n18188), .dout(n18197));
  jxor g17942(.dina(n18197), .dinb(n18180), .dout(n18198));
  jor  g17943(.dina(n9271), .dinb(n5251), .dout(n18199));
  jor  g17944(.dina(n9003), .dinb(n4839), .dout(n18200));
  jor  g17945(.dina(n9268), .dinb(n5253), .dout(n18201));
  jor  g17946(.dina(n9273), .dinb(n5040), .dout(n18202));
  jand g17947(.dina(n18202), .dinb(n18201), .dout(n18203));
  jand g17948(.dina(n18203), .dinb(n18200), .dout(n18204));
  jand g17949(.dina(n18204), .dinb(n18199), .dout(n18205));
  jxor g17950(.dina(n18205), .dinb(n8729), .dout(n18206));
  jxor g17951(.dina(n18206), .dinb(n18198), .dout(n18207));
  jxor g17952(.dina(n18207), .dinb(n18177), .dout(n18208));
  jor  g17953(.dina(n8457), .dinb(n5909), .dout(n18209));
  jor  g17954(.dina(n8185), .dinb(n5469), .dout(n18210));
  jor  g17955(.dina(n8459), .dinb(n5685), .dout(n18211));
  jor  g17956(.dina(n8454), .dinb(n5911), .dout(n18212));
  jand g17957(.dina(n18212), .dinb(n18211), .dout(n18213));
  jand g17958(.dina(n18213), .dinb(n18210), .dout(n18214));
  jand g17959(.dina(n18214), .dinb(n18209), .dout(n18215));
  jxor g17960(.dina(n18215), .dinb(n7929), .dout(n18216));
  jxor g17961(.dina(n18216), .dinb(n18208), .dout(n18217));
  jxor g17962(.dina(n18217), .dinb(n18174), .dout(n18218));
  jor  g17963(.dina(n7660), .dinb(n6603), .dout(n18219));
  jor  g17964(.dina(n7415), .dinb(n6139), .dout(n18220));
  jor  g17965(.dina(n7662), .dinb(n6605), .dout(n18221));
  jor  g17966(.dina(n7657), .dinb(n6366), .dout(n18222));
  jand g17967(.dina(n18222), .dinb(n18221), .dout(n18223));
  jand g17968(.dina(n18223), .dinb(n18220), .dout(n18224));
  jand g17969(.dina(n18224), .dinb(n18219), .dout(n18225));
  jxor g17970(.dina(n18225), .dinb(n7166), .dout(n18226));
  jxor g17971(.dina(n18226), .dinb(n18218), .dout(n18227));
  jxor g17972(.dina(n18227), .dinb(n18171), .dout(n18228));
  jor  g17973(.dina(n7336), .dinb(n6914), .dout(n18229));
  jor  g17974(.dina(n6673), .dinb(n6846), .dout(n18230));
  jor  g17975(.dina(n6916), .dinb(n7338), .dout(n18231));
  jor  g17976(.dina(n6911), .dinb(n7086), .dout(n18232));
  jand g17977(.dina(n18232), .dinb(n18231), .dout(n18233));
  jand g17978(.dina(n18233), .dinb(n18230), .dout(n18234));
  jand g17979(.dina(n18234), .dinb(n18229), .dout(n18235));
  jxor g17980(.dina(n18235), .dinb(n6443), .dout(n18236));
  jxor g17981(.dina(n18236), .dinb(n18228), .dout(n18237));
  jxor g17982(.dina(n18237), .dinb(n18168), .dout(n18238));
  jor  g17983(.dina(n8109), .dinb(n6207), .dout(n18239));
  jor  g17984(.dina(n5975), .dinb(n7590), .dout(n18240));
  jor  g17985(.dina(n6210), .dinb(n7846), .dout(n18241));
  jor  g17986(.dina(n6205), .dinb(n8111), .dout(n18242));
  jand g17987(.dina(n18242), .dinb(n18241), .dout(n18243));
  jand g17988(.dina(n18243), .dinb(n18240), .dout(n18244));
  jand g17989(.dina(n18244), .dinb(n18239), .dout(n18245));
  jxor g17990(.dina(n18245), .dinb(n5759), .dout(n18246));
  jxor g17991(.dina(n18246), .dinb(n18238), .dout(n18247));
  jxor g17992(.dina(n18247), .dinb(n18165), .dout(n18248));
  jor  g17993(.dina(n8918), .dinb(n5537), .dout(n18249));
  jor  g17994(.dina(n5315), .dinb(n8378), .dout(n18250));
  jor  g17995(.dina(n5539), .dinb(n8920), .dout(n18251));
  jor  g17996(.dina(n5534), .dinb(n8644), .dout(n18252));
  jand g17997(.dina(n18252), .dinb(n18251), .dout(n18253));
  jand g17998(.dina(n18253), .dinb(n18250), .dout(n18254));
  jand g17999(.dina(n18254), .dinb(n18249), .dout(n18255));
  jxor g18000(.dina(n18255), .dinb(n5111), .dout(n18256));
  jxor g18001(.dina(n18256), .dinb(n18248), .dout(n18257));
  jxor g18002(.dina(n18257), .dinb(n18162), .dout(n18258));
  jor  g18003(.dina(n9757), .dinb(n4902), .dout(n18259));
  jor  g18004(.dina(n4696), .dinb(n9195), .dout(n18260));
  jor  g18005(.dina(n4904), .dinb(n9475), .dout(n18261));
  jor  g18006(.dina(n4899), .dinb(n9759), .dout(n18262));
  jand g18007(.dina(n18262), .dinb(n18261), .dout(n18263));
  jand g18008(.dina(n18263), .dinb(n18260), .dout(n18264));
  jand g18009(.dina(n18264), .dinb(n18259), .dout(n18265));
  jxor g18010(.dina(n18265), .dinb(n4505), .dout(n18266));
  jxor g18011(.dina(n18266), .dinb(n18258), .dout(n18267));
  jxor g18012(.dina(n18267), .dinb(n18159), .dout(n18268));
  jxor g18013(.dina(n18268), .dinb(n18148), .dout(n18269));
  jnot g18014(.din(n18269), .dout(n18270));
  jor  g18015(.dina(n18142), .dinb(n18138), .dout(n18271));
  jor  g18016(.dina(n18144), .dinb(n18015), .dout(n18272));
  jand g18017(.dina(n18272), .dinb(n18271), .dout(n18273));
  jxor g18018(.dina(n18273), .dinb(n18270), .dout(f100 ));
  jand g18019(.dina(n18268), .dinb(n18148), .dout(n18275));
  jnot g18020(.din(n18275), .dout(n18276));
  jor  g18021(.dina(n18273), .dinb(n18270), .dout(n18277));
  jand g18022(.dina(n18277), .dinb(n18276), .dout(n18278));
  jor  g18023(.dina(n18158), .dinb(n18152), .dout(n18279));
  jand g18024(.dina(n18267), .dinb(n18159), .dout(n18280));
  jnot g18025(.din(n18280), .dout(n18281));
  jand g18026(.dina(n18281), .dinb(n18279), .dout(n18282));
  jnot g18027(.din(n18282), .dout(n18283));
  jand g18028(.dina(n18257), .dinb(n18162), .dout(n18284));
  jand g18029(.dina(n18266), .dinb(n18258), .dout(n18285));
  jor  g18030(.dina(n18285), .dinb(n18284), .dout(n18286));
  jnot g18031(.din(n18286), .dout(n18287));
  jand g18032(.dina(n4117), .dinb(b63 ), .dout(n18288));
  jand g18033(.dina(n10832), .dinb(n3930), .dout(n18289));
  jor  g18034(.dina(n18289), .dinb(n18288), .dout(n18290));
  jxor g18035(.dina(n18290), .dinb(n3938), .dout(n18291));
  jxor g18036(.dina(n18291), .dinb(n18287), .dout(n18292));
  jand g18037(.dina(n18247), .dinb(n18165), .dout(n18293));
  jand g18038(.dina(n18256), .dinb(n18248), .dout(n18294));
  jor  g18039(.dina(n18294), .dinb(n18293), .dout(n18295));
  jand g18040(.dina(n18237), .dinb(n18168), .dout(n18296));
  jand g18041(.dina(n18246), .dinb(n18238), .dout(n18297));
  jor  g18042(.dina(n18297), .dinb(n18296), .dout(n18298));
  jand g18043(.dina(n18227), .dinb(n18171), .dout(n18299));
  jand g18044(.dina(n18236), .dinb(n18228), .dout(n18300));
  jor  g18045(.dina(n18300), .dinb(n18299), .dout(n18301));
  jand g18046(.dina(n18217), .dinb(n18174), .dout(n18302));
  jand g18047(.dina(n18226), .dinb(n18218), .dout(n18303));
  jor  g18048(.dina(n18303), .dinb(n18302), .dout(n18304));
  jand g18049(.dina(n18207), .dinb(n18177), .dout(n18305));
  jand g18050(.dina(n18216), .dinb(n18208), .dout(n18306));
  jor  g18051(.dina(n18306), .dinb(n18305), .dout(n18307));
  jand g18052(.dina(n18197), .dinb(n18180), .dout(n18308));
  jand g18053(.dina(n18206), .dinb(n18198), .dout(n18309));
  jor  g18054(.dina(n18309), .dinb(n18308), .dout(n18310));
  jand g18055(.dina(n18187), .dinb(n18184), .dout(n18311));
  jand g18056(.dina(n18196), .dinb(n18188), .dout(n18312));
  jor  g18057(.dina(n18312), .dinb(n18311), .dout(n18313));
  jand g18058(.dina(n10594), .dinb(b37 ), .dout(n18314));
  jand g18059(.dina(n10129), .dinb(b38 ), .dout(n18315));
  jor  g18060(.dina(n18315), .dinb(n18314), .dout(n18316));
  jxor g18061(.dina(n18316), .dinb(n18184), .dout(n18317));
  jxor g18062(.dina(n18317), .dinb(n18313), .dout(n18318));
  jor  g18063(.dina(n10134), .dinb(n4837), .dout(n18319));
  jor  g18064(.dina(n9849), .dinb(n4437), .dout(n18320));
  jor  g18065(.dina(n10137), .dinb(n4637), .dout(n18321));
  jor  g18066(.dina(n10132), .dinb(n4839), .dout(n18322));
  jand g18067(.dina(n18322), .dinb(n18321), .dout(n18323));
  jand g18068(.dina(n18323), .dinb(n18320), .dout(n18324));
  jand g18069(.dina(n18324), .dinb(n18319), .dout(n18325));
  jxor g18070(.dina(n18325), .dinb(n9559), .dout(n18326));
  jxor g18071(.dina(n18326), .dinb(n18318), .dout(n18327));
  jor  g18072(.dina(n9271), .dinb(n5467), .dout(n18328));
  jor  g18073(.dina(n9003), .dinb(n5040), .dout(n18329));
  jor  g18074(.dina(n9268), .dinb(n5469), .dout(n18330));
  jor  g18075(.dina(n9273), .dinb(n5253), .dout(n18331));
  jand g18076(.dina(n18331), .dinb(n18330), .dout(n18332));
  jand g18077(.dina(n18332), .dinb(n18329), .dout(n18333));
  jand g18078(.dina(n18333), .dinb(n18328), .dout(n18334));
  jxor g18079(.dina(n18334), .dinb(n8729), .dout(n18335));
  jxor g18080(.dina(n18335), .dinb(n18327), .dout(n18336));
  jxor g18081(.dina(n18336), .dinb(n18310), .dout(n18337));
  jor  g18082(.dina(n8457), .dinb(n6137), .dout(n18338));
  jor  g18083(.dina(n8185), .dinb(n5685), .dout(n18339));
  jor  g18084(.dina(n8459), .dinb(n5911), .dout(n18340));
  jor  g18085(.dina(n8454), .dinb(n6139), .dout(n18341));
  jand g18086(.dina(n18341), .dinb(n18340), .dout(n18342));
  jand g18087(.dina(n18342), .dinb(n18339), .dout(n18343));
  jand g18088(.dina(n18343), .dinb(n18338), .dout(n18344));
  jxor g18089(.dina(n18344), .dinb(n7929), .dout(n18345));
  jxor g18090(.dina(n18345), .dinb(n18337), .dout(n18346));
  jxor g18091(.dina(n18346), .dinb(n18307), .dout(n18347));
  jor  g18092(.dina(n7660), .dinb(n6844), .dout(n18348));
  jor  g18093(.dina(n7415), .dinb(n6366), .dout(n18349));
  jor  g18094(.dina(n7657), .dinb(n6605), .dout(n18350));
  jor  g18095(.dina(n7662), .dinb(n6846), .dout(n18351));
  jand g18096(.dina(n18351), .dinb(n18350), .dout(n18352));
  jand g18097(.dina(n18352), .dinb(n18349), .dout(n18353));
  jand g18098(.dina(n18353), .dinb(n18348), .dout(n18354));
  jxor g18099(.dina(n18354), .dinb(n7166), .dout(n18355));
  jxor g18100(.dina(n18355), .dinb(n18347), .dout(n18356));
  jxor g18101(.dina(n18356), .dinb(n18304), .dout(n18357));
  jor  g18102(.dina(n7588), .dinb(n6914), .dout(n18358));
  jor  g18103(.dina(n6673), .dinb(n7086), .dout(n18359));
  jor  g18104(.dina(n6911), .dinb(n7338), .dout(n18360));
  jor  g18105(.dina(n6916), .dinb(n7590), .dout(n18361));
  jand g18106(.dina(n18361), .dinb(n18360), .dout(n18362));
  jand g18107(.dina(n18362), .dinb(n18359), .dout(n18363));
  jand g18108(.dina(n18363), .dinb(n18358), .dout(n18364));
  jxor g18109(.dina(n18364), .dinb(n6443), .dout(n18365));
  jxor g18110(.dina(n18365), .dinb(n18357), .dout(n18366));
  jxor g18111(.dina(n18366), .dinb(n18301), .dout(n18367));
  jor  g18112(.dina(n8376), .dinb(n6207), .dout(n18368));
  jor  g18113(.dina(n5975), .dinb(n7846), .dout(n18369));
  jor  g18114(.dina(n6205), .dinb(n8378), .dout(n18370));
  jor  g18115(.dina(n6210), .dinb(n8111), .dout(n18371));
  jand g18116(.dina(n18371), .dinb(n18370), .dout(n18372));
  jand g18117(.dina(n18372), .dinb(n18369), .dout(n18373));
  jand g18118(.dina(n18373), .dinb(n18368), .dout(n18374));
  jxor g18119(.dina(n18374), .dinb(n5759), .dout(n18375));
  jxor g18120(.dina(n18375), .dinb(n18367), .dout(n18376));
  jxor g18121(.dina(n18376), .dinb(n18298), .dout(n18377));
  jor  g18122(.dina(n9193), .dinb(n5537), .dout(n18378));
  jor  g18123(.dina(n5315), .dinb(n8644), .dout(n18379));
  jor  g18124(.dina(n5534), .dinb(n8920), .dout(n18380));
  jor  g18125(.dina(n5539), .dinb(n9195), .dout(n18381));
  jand g18126(.dina(n18381), .dinb(n18380), .dout(n18382));
  jand g18127(.dina(n18382), .dinb(n18379), .dout(n18383));
  jand g18128(.dina(n18383), .dinb(n18378), .dout(n18384));
  jxor g18129(.dina(n18384), .dinb(n5111), .dout(n18385));
  jxor g18130(.dina(n18385), .dinb(n18377), .dout(n18386));
  jxor g18131(.dina(n18386), .dinb(n18295), .dout(n18387));
  jor  g18132(.dina(n10049), .dinb(n4902), .dout(n18388));
  jor  g18133(.dina(n4696), .dinb(n9475), .dout(n18389));
  jor  g18134(.dina(n4904), .dinb(n9759), .dout(n18390));
  jor  g18135(.dina(n4899), .dinb(n10051), .dout(n18391));
  jand g18136(.dina(n18391), .dinb(n18390), .dout(n18392));
  jand g18137(.dina(n18392), .dinb(n18389), .dout(n18393));
  jand g18138(.dina(n18393), .dinb(n18388), .dout(n18394));
  jxor g18139(.dina(n18394), .dinb(n4505), .dout(n18395));
  jxor g18140(.dina(n18395), .dinb(n18387), .dout(n18396));
  jxor g18141(.dina(n18396), .dinb(n18292), .dout(n18397));
  jxor g18142(.dina(n18397), .dinb(n18283), .dout(n18398));
  jnot g18143(.din(n18398), .dout(n18399));
  jxor g18144(.dina(n18399), .dinb(n18278), .dout(f101 ));
  jand g18145(.dina(n18397), .dinb(n18283), .dout(n18401));
  jnot g18146(.din(n18401), .dout(n18402));
  jor  g18147(.dina(n18399), .dinb(n18278), .dout(n18403));
  jand g18148(.dina(n18403), .dinb(n18402), .dout(n18404));
  jand g18149(.dina(n18386), .dinb(n18295), .dout(n18405));
  jand g18150(.dina(n18395), .dinb(n18387), .dout(n18406));
  jor  g18151(.dina(n18406), .dinb(n18405), .dout(n18407));
  jand g18152(.dina(n18376), .dinb(n18298), .dout(n18408));
  jand g18153(.dina(n18385), .dinb(n18377), .dout(n18409));
  jor  g18154(.dina(n18409), .dinb(n18408), .dout(n18410));
  jand g18155(.dina(n18366), .dinb(n18301), .dout(n18411));
  jand g18156(.dina(n18375), .dinb(n18367), .dout(n18412));
  jor  g18157(.dina(n18412), .dinb(n18411), .dout(n18413));
  jand g18158(.dina(n18356), .dinb(n18304), .dout(n18414));
  jand g18159(.dina(n18365), .dinb(n18357), .dout(n18415));
  jor  g18160(.dina(n18415), .dinb(n18414), .dout(n18416));
  jand g18161(.dina(n18346), .dinb(n18307), .dout(n18417));
  jand g18162(.dina(n18355), .dinb(n18347), .dout(n18418));
  jor  g18163(.dina(n18418), .dinb(n18417), .dout(n18419));
  jand g18164(.dina(n18336), .dinb(n18310), .dout(n18420));
  jand g18165(.dina(n18345), .dinb(n18337), .dout(n18421));
  jor  g18166(.dina(n18421), .dinb(n18420), .dout(n18422));
  jand g18167(.dina(n18326), .dinb(n18318), .dout(n18423));
  jand g18168(.dina(n18335), .dinb(n18327), .dout(n18424));
  jor  g18169(.dina(n18424), .dinb(n18423), .dout(n18425));
  jand g18170(.dina(n18316), .dinb(n18184), .dout(n18426));
  jand g18171(.dina(n18317), .dinb(n18313), .dout(n18427));
  jor  g18172(.dina(n18427), .dinb(n18426), .dout(n18428));
  jand g18173(.dina(n10594), .dinb(b38 ), .dout(n18429));
  jand g18174(.dina(n10129), .dinb(b39 ), .dout(n18430));
  jor  g18175(.dina(n18430), .dinb(n18429), .dout(n18431));
  jxor g18176(.dina(n18183), .dinb(n3938), .dout(n18432));
  jxor g18177(.dina(n18432), .dinb(n18431), .dout(n18433));
  jxor g18178(.dina(n18433), .dinb(n18428), .dout(n18434));
  jor  g18179(.dina(n10134), .dinb(n5038), .dout(n18435));
  jor  g18180(.dina(n9849), .dinb(n4637), .dout(n18436));
  jor  g18181(.dina(n10137), .dinb(n4839), .dout(n18437));
  jor  g18182(.dina(n10132), .dinb(n5040), .dout(n18438));
  jand g18183(.dina(n18438), .dinb(n18437), .dout(n18439));
  jand g18184(.dina(n18439), .dinb(n18436), .dout(n18440));
  jand g18185(.dina(n18440), .dinb(n18435), .dout(n18441));
  jxor g18186(.dina(n18441), .dinb(n9559), .dout(n18442));
  jxor g18187(.dina(n18442), .dinb(n18434), .dout(n18443));
  jor  g18188(.dina(n9271), .dinb(n5683), .dout(n18444));
  jor  g18189(.dina(n9003), .dinb(n5253), .dout(n18445));
  jor  g18190(.dina(n9273), .dinb(n5469), .dout(n18446));
  jor  g18191(.dina(n9268), .dinb(n5685), .dout(n18447));
  jand g18192(.dina(n18447), .dinb(n18446), .dout(n18448));
  jand g18193(.dina(n18448), .dinb(n18445), .dout(n18449));
  jand g18194(.dina(n18449), .dinb(n18444), .dout(n18450));
  jxor g18195(.dina(n18450), .dinb(n8729), .dout(n18451));
  jxor g18196(.dina(n18451), .dinb(n18443), .dout(n18452));
  jxor g18197(.dina(n18452), .dinb(n18425), .dout(n18453));
  jor  g18198(.dina(n8457), .dinb(n6364), .dout(n18454));
  jor  g18199(.dina(n8185), .dinb(n5911), .dout(n18455));
  jor  g18200(.dina(n8454), .dinb(n6366), .dout(n18456));
  jor  g18201(.dina(n8459), .dinb(n6139), .dout(n18457));
  jand g18202(.dina(n18457), .dinb(n18456), .dout(n18458));
  jand g18203(.dina(n18458), .dinb(n18455), .dout(n18459));
  jand g18204(.dina(n18459), .dinb(n18454), .dout(n18460));
  jxor g18205(.dina(n18460), .dinb(n7929), .dout(n18461));
  jxor g18206(.dina(n18461), .dinb(n18453), .dout(n18462));
  jxor g18207(.dina(n18462), .dinb(n18422), .dout(n18463));
  jor  g18208(.dina(n7660), .dinb(n7084), .dout(n18464));
  jor  g18209(.dina(n7415), .dinb(n6605), .dout(n18465));
  jor  g18210(.dina(n7662), .dinb(n7086), .dout(n18466));
  jor  g18211(.dina(n7657), .dinb(n6846), .dout(n18467));
  jand g18212(.dina(n18467), .dinb(n18466), .dout(n18468));
  jand g18213(.dina(n18468), .dinb(n18465), .dout(n18469));
  jand g18214(.dina(n18469), .dinb(n18464), .dout(n18470));
  jxor g18215(.dina(n18470), .dinb(n7166), .dout(n18471));
  jxor g18216(.dina(n18471), .dinb(n18463), .dout(n18472));
  jxor g18217(.dina(n18472), .dinb(n18419), .dout(n18473));
  jor  g18218(.dina(n7844), .dinb(n6914), .dout(n18474));
  jor  g18219(.dina(n6673), .dinb(n7338), .dout(n18475));
  jor  g18220(.dina(n6911), .dinb(n7590), .dout(n18476));
  jor  g18221(.dina(n6916), .dinb(n7846), .dout(n18477));
  jand g18222(.dina(n18477), .dinb(n18476), .dout(n18478));
  jand g18223(.dina(n18478), .dinb(n18475), .dout(n18479));
  jand g18224(.dina(n18479), .dinb(n18474), .dout(n18480));
  jxor g18225(.dina(n18480), .dinb(n6443), .dout(n18481));
  jxor g18226(.dina(n18481), .dinb(n18473), .dout(n18482));
  jxor g18227(.dina(n18482), .dinb(n18416), .dout(n18483));
  jor  g18228(.dina(n8642), .dinb(n6207), .dout(n18484));
  jor  g18229(.dina(n5975), .dinb(n8111), .dout(n18485));
  jor  g18230(.dina(n6205), .dinb(n8644), .dout(n18486));
  jor  g18231(.dina(n6210), .dinb(n8378), .dout(n18487));
  jand g18232(.dina(n18487), .dinb(n18486), .dout(n18488));
  jand g18233(.dina(n18488), .dinb(n18485), .dout(n18489));
  jand g18234(.dina(n18489), .dinb(n18484), .dout(n18490));
  jxor g18235(.dina(n18490), .dinb(n5759), .dout(n18491));
  jxor g18236(.dina(n18491), .dinb(n18483), .dout(n18492));
  jxor g18237(.dina(n18492), .dinb(n18413), .dout(n18493));
  jor  g18238(.dina(n9473), .dinb(n5537), .dout(n18494));
  jor  g18239(.dina(n5315), .dinb(n8920), .dout(n18495));
  jor  g18240(.dina(n5539), .dinb(n9475), .dout(n18496));
  jor  g18241(.dina(n5534), .dinb(n9195), .dout(n18497));
  jand g18242(.dina(n18497), .dinb(n18496), .dout(n18498));
  jand g18243(.dina(n18498), .dinb(n18495), .dout(n18499));
  jand g18244(.dina(n18499), .dinb(n18494), .dout(n18500));
  jxor g18245(.dina(n18500), .dinb(n5111), .dout(n18501));
  jxor g18246(.dina(n18501), .dinb(n18493), .dout(n18502));
  jxor g18247(.dina(n18502), .dinb(n18410), .dout(n18503));
  jor  g18248(.dina(n10521), .dinb(n4902), .dout(n18504));
  jor  g18249(.dina(n4696), .dinb(n9759), .dout(n18505));
  jor  g18250(.dina(n4899), .dinb(n10523), .dout(n18506));
  jor  g18251(.dina(n4904), .dinb(n10051), .dout(n18507));
  jand g18252(.dina(n18507), .dinb(n18506), .dout(n18508));
  jand g18253(.dina(n18508), .dinb(n18505), .dout(n18509));
  jand g18254(.dina(n18509), .dinb(n18504), .dout(n18510));
  jxor g18255(.dina(n18510), .dinb(n4505), .dout(n18511));
  jxor g18256(.dina(n18511), .dinb(n18503), .dout(n18512));
  jxor g18257(.dina(n18512), .dinb(n18407), .dout(n18513));
  jnot g18258(.din(n18513), .dout(n18514));
  jor  g18259(.dina(n18291), .dinb(n18287), .dout(n18515));
  jand g18260(.dina(n18396), .dinb(n18292), .dout(n18516));
  jnot g18261(.din(n18516), .dout(n18517));
  jand g18262(.dina(n18517), .dinb(n18515), .dout(n18518));
  jxor g18263(.dina(n18518), .dinb(n18514), .dout(n18519));
  jnot g18264(.din(n18519), .dout(n18520));
  jxor g18265(.dina(n18520), .dinb(n18404), .dout(f102 ));
  jand g18266(.dina(n18511), .dinb(n18503), .dout(n18522));
  jand g18267(.dina(n18512), .dinb(n18407), .dout(n18523));
  jor  g18268(.dina(n18523), .dinb(n18522), .dout(n18524));
  jand g18269(.dina(n18501), .dinb(n18493), .dout(n18525));
  jand g18270(.dina(n18502), .dinb(n18410), .dout(n18526));
  jor  g18271(.dina(n18526), .dinb(n18525), .dout(n18527));
  jnot g18272(.din(n18527), .dout(n18528));
  jor  g18273(.dina(n10813), .dinb(n4902), .dout(n18529));
  jor  g18274(.dina(n4696), .dinb(n10051), .dout(n18530));
  jor  g18275(.dina(n4904), .dinb(n10523), .dout(n18531));
  jand g18276(.dina(n18531), .dinb(n18530), .dout(n18532));
  jand g18277(.dina(n18532), .dinb(n18529), .dout(n18533));
  jxor g18278(.dina(n18533), .dinb(a41 ), .dout(n18534));
  jxor g18279(.dina(n18534), .dinb(n18528), .dout(n18535));
  jand g18280(.dina(n18491), .dinb(n18483), .dout(n18536));
  jand g18281(.dina(n18492), .dinb(n18413), .dout(n18537));
  jor  g18282(.dina(n18537), .dinb(n18536), .dout(n18538));
  jand g18283(.dina(n18481), .dinb(n18473), .dout(n18539));
  jand g18284(.dina(n18482), .dinb(n18416), .dout(n18540));
  jor  g18285(.dina(n18540), .dinb(n18539), .dout(n18541));
  jand g18286(.dina(n18471), .dinb(n18463), .dout(n18542));
  jand g18287(.dina(n18472), .dinb(n18419), .dout(n18543));
  jor  g18288(.dina(n18543), .dinb(n18542), .dout(n18544));
  jand g18289(.dina(n18461), .dinb(n18453), .dout(n18545));
  jand g18290(.dina(n18462), .dinb(n18422), .dout(n18546));
  jor  g18291(.dina(n18546), .dinb(n18545), .dout(n18547));
  jand g18292(.dina(n18451), .dinb(n18443), .dout(n18548));
  jand g18293(.dina(n18452), .dinb(n18425), .dout(n18549));
  jor  g18294(.dina(n18549), .dinb(n18548), .dout(n18550));
  jand g18295(.dina(n18433), .dinb(n18428), .dout(n18551));
  jand g18296(.dina(n18442), .dinb(n18434), .dout(n18552));
  jor  g18297(.dina(n18552), .dinb(n18551), .dout(n18553));
  jand g18298(.dina(n10594), .dinb(b39 ), .dout(n18554));
  jand g18299(.dina(n10129), .dinb(b40 ), .dout(n18555));
  jor  g18300(.dina(n18555), .dinb(n18554), .dout(n18556));
  jnot g18301(.din(n18556), .dout(n18557));
  jand g18302(.dina(n18183), .dinb(n3938), .dout(n18558));
  jand g18303(.dina(n18432), .dinb(n18431), .dout(n18559));
  jor  g18304(.dina(n18559), .dinb(n18558), .dout(n18560));
  jxor g18305(.dina(n18560), .dinb(n18557), .dout(n18561));
  jor  g18306(.dina(n10134), .dinb(n5251), .dout(n18562));
  jor  g18307(.dina(n9849), .dinb(n4839), .dout(n18563));
  jor  g18308(.dina(n10132), .dinb(n5253), .dout(n18564));
  jor  g18309(.dina(n10137), .dinb(n5040), .dout(n18565));
  jand g18310(.dina(n18565), .dinb(n18564), .dout(n18566));
  jand g18311(.dina(n18566), .dinb(n18563), .dout(n18567));
  jand g18312(.dina(n18567), .dinb(n18562), .dout(n18568));
  jxor g18313(.dina(n18568), .dinb(n9559), .dout(n18569));
  jxor g18314(.dina(n18569), .dinb(n18561), .dout(n18570));
  jxor g18315(.dina(n18570), .dinb(n18553), .dout(n18571));
  jor  g18316(.dina(n9271), .dinb(n5909), .dout(n18572));
  jor  g18317(.dina(n9003), .dinb(n5469), .dout(n18573));
  jor  g18318(.dina(n9268), .dinb(n5911), .dout(n18574));
  jor  g18319(.dina(n9273), .dinb(n5685), .dout(n18575));
  jand g18320(.dina(n18575), .dinb(n18574), .dout(n18576));
  jand g18321(.dina(n18576), .dinb(n18573), .dout(n18577));
  jand g18322(.dina(n18577), .dinb(n18572), .dout(n18578));
  jxor g18323(.dina(n18578), .dinb(n8729), .dout(n18579));
  jxor g18324(.dina(n18579), .dinb(n18571), .dout(n18580));
  jxor g18325(.dina(n18580), .dinb(n18550), .dout(n18581));
  jor  g18326(.dina(n8457), .dinb(n6603), .dout(n18582));
  jor  g18327(.dina(n8185), .dinb(n6139), .dout(n18583));
  jor  g18328(.dina(n8459), .dinb(n6366), .dout(n18584));
  jor  g18329(.dina(n8454), .dinb(n6605), .dout(n18585));
  jand g18330(.dina(n18585), .dinb(n18584), .dout(n18586));
  jand g18331(.dina(n18586), .dinb(n18583), .dout(n18587));
  jand g18332(.dina(n18587), .dinb(n18582), .dout(n18588));
  jxor g18333(.dina(n18588), .dinb(n7929), .dout(n18589));
  jxor g18334(.dina(n18589), .dinb(n18581), .dout(n18590));
  jxor g18335(.dina(n18590), .dinb(n18547), .dout(n18591));
  jor  g18336(.dina(n7336), .dinb(n7660), .dout(n18592));
  jor  g18337(.dina(n7415), .dinb(n6846), .dout(n18593));
  jor  g18338(.dina(n7662), .dinb(n7338), .dout(n18594));
  jor  g18339(.dina(n7657), .dinb(n7086), .dout(n18595));
  jand g18340(.dina(n18595), .dinb(n18594), .dout(n18596));
  jand g18341(.dina(n18596), .dinb(n18593), .dout(n18597));
  jand g18342(.dina(n18597), .dinb(n18592), .dout(n18598));
  jxor g18343(.dina(n18598), .dinb(n7166), .dout(n18599));
  jxor g18344(.dina(n18599), .dinb(n18591), .dout(n18600));
  jxor g18345(.dina(n18600), .dinb(n18544), .dout(n18601));
  jor  g18346(.dina(n8109), .dinb(n6914), .dout(n18602));
  jor  g18347(.dina(n6673), .dinb(n7590), .dout(n18603));
  jor  g18348(.dina(n6916), .dinb(n8111), .dout(n18604));
  jor  g18349(.dina(n6911), .dinb(n7846), .dout(n18605));
  jand g18350(.dina(n18605), .dinb(n18604), .dout(n18606));
  jand g18351(.dina(n18606), .dinb(n18603), .dout(n18607));
  jand g18352(.dina(n18607), .dinb(n18602), .dout(n18608));
  jxor g18353(.dina(n18608), .dinb(n6443), .dout(n18609));
  jxor g18354(.dina(n18609), .dinb(n18601), .dout(n18610));
  jxor g18355(.dina(n18610), .dinb(n18541), .dout(n18611));
  jor  g18356(.dina(n8918), .dinb(n6207), .dout(n18612));
  jor  g18357(.dina(n5975), .dinb(n8378), .dout(n18613));
  jor  g18358(.dina(n6210), .dinb(n8644), .dout(n18614));
  jor  g18359(.dina(n6205), .dinb(n8920), .dout(n18615));
  jand g18360(.dina(n18615), .dinb(n18614), .dout(n18616));
  jand g18361(.dina(n18616), .dinb(n18613), .dout(n18617));
  jand g18362(.dina(n18617), .dinb(n18612), .dout(n18618));
  jxor g18363(.dina(n18618), .dinb(n5759), .dout(n18619));
  jxor g18364(.dina(n18619), .dinb(n18611), .dout(n18620));
  jxor g18365(.dina(n18620), .dinb(n18538), .dout(n18621));
  jor  g18366(.dina(n9757), .dinb(n5537), .dout(n18622));
  jor  g18367(.dina(n5315), .dinb(n9195), .dout(n18623));
  jor  g18368(.dina(n5539), .dinb(n9759), .dout(n18624));
  jor  g18369(.dina(n5534), .dinb(n9475), .dout(n18625));
  jand g18370(.dina(n18625), .dinb(n18624), .dout(n18626));
  jand g18371(.dina(n18626), .dinb(n18623), .dout(n18627));
  jand g18372(.dina(n18627), .dinb(n18622), .dout(n18628));
  jxor g18373(.dina(n18628), .dinb(n5111), .dout(n18629));
  jxor g18374(.dina(n18629), .dinb(n18621), .dout(n18630));
  jxor g18375(.dina(n18630), .dinb(n18535), .dout(n18631));
  jxor g18376(.dina(n18631), .dinb(n18524), .dout(n18632));
  jnot g18377(.din(n18632), .dout(n18633));
  jor  g18378(.dina(n18518), .dinb(n18514), .dout(n18634));
  jor  g18379(.dina(n18520), .dinb(n18404), .dout(n18635));
  jand g18380(.dina(n18635), .dinb(n18634), .dout(n18636));
  jxor g18381(.dina(n18636), .dinb(n18633), .dout(f103 ));
  jand g18382(.dina(n18631), .dinb(n18524), .dout(n18638));
  jnot g18383(.din(n18638), .dout(n18639));
  jor  g18384(.dina(n18636), .dinb(n18633), .dout(n18640));
  jand g18385(.dina(n18640), .dinb(n18639), .dout(n18641));
  jor  g18386(.dina(n18534), .dinb(n18528), .dout(n18642));
  jand g18387(.dina(n18630), .dinb(n18535), .dout(n18643));
  jnot g18388(.din(n18643), .dout(n18644));
  jand g18389(.dina(n18644), .dinb(n18642), .dout(n18645));
  jnot g18390(.din(n18645), .dout(n18646));
  jand g18391(.dina(n18620), .dinb(n18538), .dout(n18647));
  jand g18392(.dina(n18629), .dinb(n18621), .dout(n18648));
  jor  g18393(.dina(n18648), .dinb(n18647), .dout(n18649));
  jnot g18394(.din(n18649), .dout(n18650));
  jand g18395(.dina(n4697), .dinb(b63 ), .dout(n18651));
  jand g18396(.dina(n10832), .dinb(n4494), .dout(n18652));
  jor  g18397(.dina(n18652), .dinb(n18651), .dout(n18653));
  jxor g18398(.dina(n18653), .dinb(n4505), .dout(n18654));
  jxor g18399(.dina(n18654), .dinb(n18650), .dout(n18655));
  jand g18400(.dina(n18610), .dinb(n18541), .dout(n18656));
  jand g18401(.dina(n18619), .dinb(n18611), .dout(n18657));
  jor  g18402(.dina(n18657), .dinb(n18656), .dout(n18658));
  jand g18403(.dina(n18600), .dinb(n18544), .dout(n18659));
  jand g18404(.dina(n18609), .dinb(n18601), .dout(n18660));
  jor  g18405(.dina(n18660), .dinb(n18659), .dout(n18661));
  jand g18406(.dina(n18590), .dinb(n18547), .dout(n18662));
  jand g18407(.dina(n18599), .dinb(n18591), .dout(n18663));
  jor  g18408(.dina(n18663), .dinb(n18662), .dout(n18664));
  jand g18409(.dina(n18580), .dinb(n18550), .dout(n18665));
  jand g18410(.dina(n18589), .dinb(n18581), .dout(n18666));
  jor  g18411(.dina(n18666), .dinb(n18665), .dout(n18667));
  jand g18412(.dina(n18570), .dinb(n18553), .dout(n18668));
  jand g18413(.dina(n18579), .dinb(n18571), .dout(n18669));
  jor  g18414(.dina(n18669), .dinb(n18668), .dout(n18670));
  jand g18415(.dina(n18560), .dinb(n18557), .dout(n18671));
  jand g18416(.dina(n18569), .dinb(n18561), .dout(n18672));
  jor  g18417(.dina(n18672), .dinb(n18671), .dout(n18673));
  jand g18418(.dina(n10594), .dinb(b40 ), .dout(n18674));
  jand g18419(.dina(n10129), .dinb(b41 ), .dout(n18675));
  jor  g18420(.dina(n18675), .dinb(n18674), .dout(n18676));
  jxor g18421(.dina(n18676), .dinb(n18557), .dout(n18677));
  jxor g18422(.dina(n18677), .dinb(n18673), .dout(n18678));
  jor  g18423(.dina(n10134), .dinb(n5467), .dout(n18679));
  jor  g18424(.dina(n9849), .dinb(n5040), .dout(n18680));
  jor  g18425(.dina(n10137), .dinb(n5253), .dout(n18681));
  jor  g18426(.dina(n10132), .dinb(n5469), .dout(n18682));
  jand g18427(.dina(n18682), .dinb(n18681), .dout(n18683));
  jand g18428(.dina(n18683), .dinb(n18680), .dout(n18684));
  jand g18429(.dina(n18684), .dinb(n18679), .dout(n18685));
  jxor g18430(.dina(n18685), .dinb(n9559), .dout(n18686));
  jxor g18431(.dina(n18686), .dinb(n18678), .dout(n18687));
  jor  g18432(.dina(n9271), .dinb(n6137), .dout(n18688));
  jor  g18433(.dina(n9003), .dinb(n5685), .dout(n18689));
  jor  g18434(.dina(n9273), .dinb(n5911), .dout(n18690));
  jor  g18435(.dina(n9268), .dinb(n6139), .dout(n18691));
  jand g18436(.dina(n18691), .dinb(n18690), .dout(n18692));
  jand g18437(.dina(n18692), .dinb(n18689), .dout(n18693));
  jand g18438(.dina(n18693), .dinb(n18688), .dout(n18694));
  jxor g18439(.dina(n18694), .dinb(n8729), .dout(n18695));
  jxor g18440(.dina(n18695), .dinb(n18687), .dout(n18696));
  jxor g18441(.dina(n18696), .dinb(n18670), .dout(n18697));
  jor  g18442(.dina(n8457), .dinb(n6844), .dout(n18698));
  jor  g18443(.dina(n8185), .dinb(n6366), .dout(n18699));
  jor  g18444(.dina(n8459), .dinb(n6605), .dout(n18700));
  jor  g18445(.dina(n8454), .dinb(n6846), .dout(n18701));
  jand g18446(.dina(n18701), .dinb(n18700), .dout(n18702));
  jand g18447(.dina(n18702), .dinb(n18699), .dout(n18703));
  jand g18448(.dina(n18703), .dinb(n18698), .dout(n18704));
  jxor g18449(.dina(n18704), .dinb(n7929), .dout(n18705));
  jxor g18450(.dina(n18705), .dinb(n18697), .dout(n18706));
  jxor g18451(.dina(n18706), .dinb(n18667), .dout(n18707));
  jor  g18452(.dina(n7588), .dinb(n7660), .dout(n18708));
  jor  g18453(.dina(n7415), .dinb(n7086), .dout(n18709));
  jor  g18454(.dina(n7657), .dinb(n7338), .dout(n18710));
  jor  g18455(.dina(n7662), .dinb(n7590), .dout(n18711));
  jand g18456(.dina(n18711), .dinb(n18710), .dout(n18712));
  jand g18457(.dina(n18712), .dinb(n18709), .dout(n18713));
  jand g18458(.dina(n18713), .dinb(n18708), .dout(n18714));
  jxor g18459(.dina(n18714), .dinb(n7166), .dout(n18715));
  jxor g18460(.dina(n18715), .dinb(n18707), .dout(n18716));
  jxor g18461(.dina(n18716), .dinb(n18664), .dout(n18717));
  jor  g18462(.dina(n8376), .dinb(n6914), .dout(n18718));
  jor  g18463(.dina(n6673), .dinb(n7846), .dout(n18719));
  jor  g18464(.dina(n6911), .dinb(n8111), .dout(n18720));
  jor  g18465(.dina(n6916), .dinb(n8378), .dout(n18721));
  jand g18466(.dina(n18721), .dinb(n18720), .dout(n18722));
  jand g18467(.dina(n18722), .dinb(n18719), .dout(n18723));
  jand g18468(.dina(n18723), .dinb(n18718), .dout(n18724));
  jxor g18469(.dina(n18724), .dinb(n6443), .dout(n18725));
  jxor g18470(.dina(n18725), .dinb(n18717), .dout(n18726));
  jxor g18471(.dina(n18726), .dinb(n18661), .dout(n18727));
  jor  g18472(.dina(n9193), .dinb(n6207), .dout(n18728));
  jor  g18473(.dina(n5975), .dinb(n8644), .dout(n18729));
  jor  g18474(.dina(n6205), .dinb(n9195), .dout(n18730));
  jor  g18475(.dina(n6210), .dinb(n8920), .dout(n18731));
  jand g18476(.dina(n18731), .dinb(n18730), .dout(n18732));
  jand g18477(.dina(n18732), .dinb(n18729), .dout(n18733));
  jand g18478(.dina(n18733), .dinb(n18728), .dout(n18734));
  jxor g18479(.dina(n18734), .dinb(n5759), .dout(n18735));
  jxor g18480(.dina(n18735), .dinb(n18727), .dout(n18736));
  jxor g18481(.dina(n18736), .dinb(n18658), .dout(n18737));
  jor  g18482(.dina(n10049), .dinb(n5537), .dout(n18738));
  jor  g18483(.dina(n5315), .dinb(n9475), .dout(n18739));
  jor  g18484(.dina(n5539), .dinb(n10051), .dout(n18740));
  jor  g18485(.dina(n5534), .dinb(n9759), .dout(n18741));
  jand g18486(.dina(n18741), .dinb(n18740), .dout(n18742));
  jand g18487(.dina(n18742), .dinb(n18739), .dout(n18743));
  jand g18488(.dina(n18743), .dinb(n18738), .dout(n18744));
  jxor g18489(.dina(n18744), .dinb(n5111), .dout(n18745));
  jxor g18490(.dina(n18745), .dinb(n18737), .dout(n18746));
  jxor g18491(.dina(n18746), .dinb(n18655), .dout(n18747));
  jxor g18492(.dina(n18747), .dinb(n18646), .dout(n18748));
  jnot g18493(.din(n18748), .dout(n18749));
  jxor g18494(.dina(n18749), .dinb(n18641), .dout(f104 ));
  jand g18495(.dina(n18747), .dinb(n18646), .dout(n18751));
  jnot g18496(.din(n18751), .dout(n18752));
  jor  g18497(.dina(n18749), .dinb(n18641), .dout(n18753));
  jand g18498(.dina(n18753), .dinb(n18752), .dout(n18754));
  jand g18499(.dina(n18736), .dinb(n18658), .dout(n18755));
  jand g18500(.dina(n18745), .dinb(n18737), .dout(n18756));
  jor  g18501(.dina(n18756), .dinb(n18755), .dout(n18757));
  jand g18502(.dina(n18726), .dinb(n18661), .dout(n18758));
  jand g18503(.dina(n18735), .dinb(n18727), .dout(n18759));
  jor  g18504(.dina(n18759), .dinb(n18758), .dout(n18760));
  jand g18505(.dina(n18716), .dinb(n18664), .dout(n18761));
  jand g18506(.dina(n18725), .dinb(n18717), .dout(n18762));
  jor  g18507(.dina(n18762), .dinb(n18761), .dout(n18763));
  jand g18508(.dina(n18706), .dinb(n18667), .dout(n18764));
  jand g18509(.dina(n18715), .dinb(n18707), .dout(n18765));
  jor  g18510(.dina(n18765), .dinb(n18764), .dout(n18766));
  jand g18511(.dina(n18696), .dinb(n18670), .dout(n18767));
  jand g18512(.dina(n18705), .dinb(n18697), .dout(n18768));
  jor  g18513(.dina(n18768), .dinb(n18767), .dout(n18769));
  jand g18514(.dina(n18686), .dinb(n18678), .dout(n18770));
  jand g18515(.dina(n18695), .dinb(n18687), .dout(n18771));
  jor  g18516(.dina(n18771), .dinb(n18770), .dout(n18772));
  jand g18517(.dina(n18676), .dinb(n18557), .dout(n18773));
  jand g18518(.dina(n18677), .dinb(n18673), .dout(n18774));
  jor  g18519(.dina(n18774), .dinb(n18773), .dout(n18775));
  jand g18520(.dina(n10594), .dinb(b41 ), .dout(n18776));
  jand g18521(.dina(n10129), .dinb(b42 ), .dout(n18777));
  jor  g18522(.dina(n18777), .dinb(n18776), .dout(n18778));
  jxor g18523(.dina(n18556), .dinb(n4505), .dout(n18779));
  jxor g18524(.dina(n18779), .dinb(n18778), .dout(n18780));
  jor  g18525(.dina(n10134), .dinb(n5683), .dout(n18781));
  jor  g18526(.dina(n9849), .dinb(n5253), .dout(n18782));
  jor  g18527(.dina(n10137), .dinb(n5469), .dout(n18783));
  jor  g18528(.dina(n10132), .dinb(n5685), .dout(n18784));
  jand g18529(.dina(n18784), .dinb(n18783), .dout(n18785));
  jand g18530(.dina(n18785), .dinb(n18782), .dout(n18786));
  jand g18531(.dina(n18786), .dinb(n18781), .dout(n18787));
  jxor g18532(.dina(n18787), .dinb(n9559), .dout(n18788));
  jxor g18533(.dina(n18788), .dinb(n18780), .dout(n18789));
  jxor g18534(.dina(n18789), .dinb(n18775), .dout(n18790));
  jor  g18535(.dina(n9271), .dinb(n6364), .dout(n18791));
  jor  g18536(.dina(n9003), .dinb(n5911), .dout(n18792));
  jor  g18537(.dina(n9273), .dinb(n6139), .dout(n18793));
  jor  g18538(.dina(n9268), .dinb(n6366), .dout(n18794));
  jand g18539(.dina(n18794), .dinb(n18793), .dout(n18795));
  jand g18540(.dina(n18795), .dinb(n18792), .dout(n18796));
  jand g18541(.dina(n18796), .dinb(n18791), .dout(n18797));
  jxor g18542(.dina(n18797), .dinb(n8729), .dout(n18798));
  jxor g18543(.dina(n18798), .dinb(n18790), .dout(n18799));
  jxor g18544(.dina(n18799), .dinb(n18772), .dout(n18800));
  jor  g18545(.dina(n8457), .dinb(n7084), .dout(n18801));
  jor  g18546(.dina(n8185), .dinb(n6605), .dout(n18802));
  jor  g18547(.dina(n8454), .dinb(n7086), .dout(n18803));
  jor  g18548(.dina(n8459), .dinb(n6846), .dout(n18804));
  jand g18549(.dina(n18804), .dinb(n18803), .dout(n18805));
  jand g18550(.dina(n18805), .dinb(n18802), .dout(n18806));
  jand g18551(.dina(n18806), .dinb(n18801), .dout(n18807));
  jxor g18552(.dina(n18807), .dinb(n7929), .dout(n18808));
  jxor g18553(.dina(n18808), .dinb(n18800), .dout(n18809));
  jxor g18554(.dina(n18809), .dinb(n18769), .dout(n18810));
  jor  g18555(.dina(n7844), .dinb(n7660), .dout(n18811));
  jor  g18556(.dina(n7415), .dinb(n7338), .dout(n18812));
  jor  g18557(.dina(n7662), .dinb(n7846), .dout(n18813));
  jor  g18558(.dina(n7657), .dinb(n7590), .dout(n18814));
  jand g18559(.dina(n18814), .dinb(n18813), .dout(n18815));
  jand g18560(.dina(n18815), .dinb(n18812), .dout(n18816));
  jand g18561(.dina(n18816), .dinb(n18811), .dout(n18817));
  jxor g18562(.dina(n18817), .dinb(n7166), .dout(n18818));
  jxor g18563(.dina(n18818), .dinb(n18810), .dout(n18819));
  jxor g18564(.dina(n18819), .dinb(n18766), .dout(n18820));
  jor  g18565(.dina(n8642), .dinb(n6914), .dout(n18821));
  jor  g18566(.dina(n6673), .dinb(n8111), .dout(n18822));
  jor  g18567(.dina(n6911), .dinb(n8378), .dout(n18823));
  jor  g18568(.dina(n6916), .dinb(n8644), .dout(n18824));
  jand g18569(.dina(n18824), .dinb(n18823), .dout(n18825));
  jand g18570(.dina(n18825), .dinb(n18822), .dout(n18826));
  jand g18571(.dina(n18826), .dinb(n18821), .dout(n18827));
  jxor g18572(.dina(n18827), .dinb(n6443), .dout(n18828));
  jxor g18573(.dina(n18828), .dinb(n18820), .dout(n18829));
  jxor g18574(.dina(n18829), .dinb(n18763), .dout(n18830));
  jor  g18575(.dina(n9473), .dinb(n6207), .dout(n18831));
  jor  g18576(.dina(n5975), .dinb(n8920), .dout(n18832));
  jor  g18577(.dina(n6210), .dinb(n9195), .dout(n18833));
  jor  g18578(.dina(n6205), .dinb(n9475), .dout(n18834));
  jand g18579(.dina(n18834), .dinb(n18833), .dout(n18835));
  jand g18580(.dina(n18835), .dinb(n18832), .dout(n18836));
  jand g18581(.dina(n18836), .dinb(n18831), .dout(n18837));
  jxor g18582(.dina(n18837), .dinb(n5759), .dout(n18838));
  jxor g18583(.dina(n18838), .dinb(n18830), .dout(n18839));
  jxor g18584(.dina(n18839), .dinb(n18760), .dout(n18840));
  jor  g18585(.dina(n10521), .dinb(n5537), .dout(n18841));
  jor  g18586(.dina(n5315), .dinb(n9759), .dout(n18842));
  jor  g18587(.dina(n5539), .dinb(n10523), .dout(n18843));
  jor  g18588(.dina(n5534), .dinb(n10051), .dout(n18844));
  jand g18589(.dina(n18844), .dinb(n18843), .dout(n18845));
  jand g18590(.dina(n18845), .dinb(n18842), .dout(n18846));
  jand g18591(.dina(n18846), .dinb(n18841), .dout(n18847));
  jxor g18592(.dina(n18847), .dinb(n5111), .dout(n18848));
  jxor g18593(.dina(n18848), .dinb(n18840), .dout(n18849));
  jxor g18594(.dina(n18849), .dinb(n18757), .dout(n18850));
  jnot g18595(.din(n18850), .dout(n18851));
  jor  g18596(.dina(n18654), .dinb(n18650), .dout(n18852));
  jand g18597(.dina(n18746), .dinb(n18655), .dout(n18853));
  jnot g18598(.din(n18853), .dout(n18854));
  jand g18599(.dina(n18854), .dinb(n18852), .dout(n18855));
  jxor g18600(.dina(n18855), .dinb(n18851), .dout(n18856));
  jnot g18601(.din(n18856), .dout(n18857));
  jxor g18602(.dina(n18857), .dinb(n18754), .dout(f105 ));
  jand g18603(.dina(n18848), .dinb(n18840), .dout(n18859));
  jand g18604(.dina(n18849), .dinb(n18757), .dout(n18860));
  jor  g18605(.dina(n18860), .dinb(n18859), .dout(n18861));
  jand g18606(.dina(n18838), .dinb(n18830), .dout(n18862));
  jand g18607(.dina(n18839), .dinb(n18760), .dout(n18863));
  jor  g18608(.dina(n18863), .dinb(n18862), .dout(n18864));
  jnot g18609(.din(n18864), .dout(n18865));
  jor  g18610(.dina(n10813), .dinb(n5537), .dout(n18866));
  jor  g18611(.dina(n5315), .dinb(n10051), .dout(n18867));
  jor  g18612(.dina(n5534), .dinb(n10523), .dout(n18868));
  jand g18613(.dina(n18868), .dinb(n18867), .dout(n18869));
  jand g18614(.dina(n18869), .dinb(n18866), .dout(n18870));
  jxor g18615(.dina(n18870), .dinb(a44 ), .dout(n18871));
  jxor g18616(.dina(n18871), .dinb(n18865), .dout(n18872));
  jand g18617(.dina(n18828), .dinb(n18820), .dout(n18873));
  jand g18618(.dina(n18829), .dinb(n18763), .dout(n18874));
  jor  g18619(.dina(n18874), .dinb(n18873), .dout(n18875));
  jand g18620(.dina(n18818), .dinb(n18810), .dout(n18876));
  jand g18621(.dina(n18819), .dinb(n18766), .dout(n18877));
  jor  g18622(.dina(n18877), .dinb(n18876), .dout(n18878));
  jand g18623(.dina(n18808), .dinb(n18800), .dout(n18879));
  jand g18624(.dina(n18809), .dinb(n18769), .dout(n18880));
  jor  g18625(.dina(n18880), .dinb(n18879), .dout(n18881));
  jand g18626(.dina(n18798), .dinb(n18790), .dout(n18882));
  jand g18627(.dina(n18799), .dinb(n18772), .dout(n18883));
  jor  g18628(.dina(n18883), .dinb(n18882), .dout(n18884));
  jand g18629(.dina(n18788), .dinb(n18780), .dout(n18885));
  jand g18630(.dina(n18789), .dinb(n18775), .dout(n18886));
  jor  g18631(.dina(n18886), .dinb(n18885), .dout(n18887));
  jand g18632(.dina(n10594), .dinb(b42 ), .dout(n18888));
  jand g18633(.dina(n10129), .dinb(b43 ), .dout(n18889));
  jor  g18634(.dina(n18889), .dinb(n18888), .dout(n18890));
  jnot g18635(.din(n18890), .dout(n18891));
  jand g18636(.dina(n18556), .dinb(n4505), .dout(n18892));
  jand g18637(.dina(n18779), .dinb(n18778), .dout(n18893));
  jor  g18638(.dina(n18893), .dinb(n18892), .dout(n18894));
  jxor g18639(.dina(n18894), .dinb(n18891), .dout(n18895));
  jor  g18640(.dina(n10134), .dinb(n5909), .dout(n18896));
  jor  g18641(.dina(n9849), .dinb(n5469), .dout(n18897));
  jor  g18642(.dina(n10137), .dinb(n5685), .dout(n18898));
  jor  g18643(.dina(n10132), .dinb(n5911), .dout(n18899));
  jand g18644(.dina(n18899), .dinb(n18898), .dout(n18900));
  jand g18645(.dina(n18900), .dinb(n18897), .dout(n18901));
  jand g18646(.dina(n18901), .dinb(n18896), .dout(n18902));
  jxor g18647(.dina(n18902), .dinb(n9559), .dout(n18903));
  jxor g18648(.dina(n18903), .dinb(n18895), .dout(n18904));
  jxor g18649(.dina(n18904), .dinb(n18887), .dout(n18905));
  jor  g18650(.dina(n9271), .dinb(n6603), .dout(n18906));
  jor  g18651(.dina(n9003), .dinb(n6139), .dout(n18907));
  jor  g18652(.dina(n9268), .dinb(n6605), .dout(n18908));
  jor  g18653(.dina(n9273), .dinb(n6366), .dout(n18909));
  jand g18654(.dina(n18909), .dinb(n18908), .dout(n18910));
  jand g18655(.dina(n18910), .dinb(n18907), .dout(n18911));
  jand g18656(.dina(n18911), .dinb(n18906), .dout(n18912));
  jxor g18657(.dina(n18912), .dinb(n8729), .dout(n18913));
  jxor g18658(.dina(n18913), .dinb(n18905), .dout(n18914));
  jxor g18659(.dina(n18914), .dinb(n18884), .dout(n18915));
  jor  g18660(.dina(n8457), .dinb(n7336), .dout(n18916));
  jor  g18661(.dina(n8185), .dinb(n6846), .dout(n18917));
  jor  g18662(.dina(n8454), .dinb(n7338), .dout(n18918));
  jor  g18663(.dina(n8459), .dinb(n7086), .dout(n18919));
  jand g18664(.dina(n18919), .dinb(n18918), .dout(n18920));
  jand g18665(.dina(n18920), .dinb(n18917), .dout(n18921));
  jand g18666(.dina(n18921), .dinb(n18916), .dout(n18922));
  jxor g18667(.dina(n18922), .dinb(n7929), .dout(n18923));
  jxor g18668(.dina(n18923), .dinb(n18915), .dout(n18924));
  jxor g18669(.dina(n18924), .dinb(n18881), .dout(n18925));
  jor  g18670(.dina(n8109), .dinb(n7660), .dout(n18926));
  jor  g18671(.dina(n7415), .dinb(n7590), .dout(n18927));
  jor  g18672(.dina(n7662), .dinb(n8111), .dout(n18928));
  jor  g18673(.dina(n7657), .dinb(n7846), .dout(n18929));
  jand g18674(.dina(n18929), .dinb(n18928), .dout(n18930));
  jand g18675(.dina(n18930), .dinb(n18927), .dout(n18931));
  jand g18676(.dina(n18931), .dinb(n18926), .dout(n18932));
  jxor g18677(.dina(n18932), .dinb(n7166), .dout(n18933));
  jxor g18678(.dina(n18933), .dinb(n18925), .dout(n18934));
  jxor g18679(.dina(n18934), .dinb(n18878), .dout(n18935));
  jor  g18680(.dina(n8918), .dinb(n6914), .dout(n18936));
  jor  g18681(.dina(n6673), .dinb(n8378), .dout(n18937));
  jor  g18682(.dina(n6911), .dinb(n8644), .dout(n18938));
  jor  g18683(.dina(n6916), .dinb(n8920), .dout(n18939));
  jand g18684(.dina(n18939), .dinb(n18938), .dout(n18940));
  jand g18685(.dina(n18940), .dinb(n18937), .dout(n18941));
  jand g18686(.dina(n18941), .dinb(n18936), .dout(n18942));
  jxor g18687(.dina(n18942), .dinb(n6443), .dout(n18943));
  jxor g18688(.dina(n18943), .dinb(n18935), .dout(n18944));
  jxor g18689(.dina(n18944), .dinb(n18875), .dout(n18945));
  jor  g18690(.dina(n9757), .dinb(n6207), .dout(n18946));
  jor  g18691(.dina(n5975), .dinb(n9195), .dout(n18947));
  jor  g18692(.dina(n6210), .dinb(n9475), .dout(n18948));
  jor  g18693(.dina(n6205), .dinb(n9759), .dout(n18949));
  jand g18694(.dina(n18949), .dinb(n18948), .dout(n18950));
  jand g18695(.dina(n18950), .dinb(n18947), .dout(n18951));
  jand g18696(.dina(n18951), .dinb(n18946), .dout(n18952));
  jxor g18697(.dina(n18952), .dinb(n5759), .dout(n18953));
  jxor g18698(.dina(n18953), .dinb(n18945), .dout(n18954));
  jxor g18699(.dina(n18954), .dinb(n18872), .dout(n18955));
  jxor g18700(.dina(n18955), .dinb(n18861), .dout(n18956));
  jnot g18701(.din(n18956), .dout(n18957));
  jor  g18702(.dina(n18855), .dinb(n18851), .dout(n18958));
  jor  g18703(.dina(n18857), .dinb(n18754), .dout(n18959));
  jand g18704(.dina(n18959), .dinb(n18958), .dout(n18960));
  jxor g18705(.dina(n18960), .dinb(n18957), .dout(f106 ));
  jand g18706(.dina(n18955), .dinb(n18861), .dout(n18962));
  jnot g18707(.din(n18962), .dout(n18963));
  jor  g18708(.dina(n18960), .dinb(n18957), .dout(n18964));
  jand g18709(.dina(n18964), .dinb(n18963), .dout(n18965));
  jor  g18710(.dina(n18871), .dinb(n18865), .dout(n18966));
  jand g18711(.dina(n18954), .dinb(n18872), .dout(n18967));
  jnot g18712(.din(n18967), .dout(n18968));
  jand g18713(.dina(n18968), .dinb(n18966), .dout(n18969));
  jnot g18714(.din(n18969), .dout(n18970));
  jand g18715(.dina(n18944), .dinb(n18875), .dout(n18971));
  jand g18716(.dina(n18953), .dinb(n18945), .dout(n18972));
  jor  g18717(.dina(n18972), .dinb(n18971), .dout(n18973));
  jnot g18718(.din(n18973), .dout(n18974));
  jand g18719(.dina(n5316), .dinb(b63 ), .dout(n18975));
  jand g18720(.dina(n10832), .dinb(n5100), .dout(n18976));
  jor  g18721(.dina(n18976), .dinb(n18975), .dout(n18977));
  jxor g18722(.dina(n18977), .dinb(n5111), .dout(n18978));
  jxor g18723(.dina(n18978), .dinb(n18974), .dout(n18979));
  jand g18724(.dina(n18934), .dinb(n18878), .dout(n18980));
  jand g18725(.dina(n18943), .dinb(n18935), .dout(n18981));
  jor  g18726(.dina(n18981), .dinb(n18980), .dout(n18982));
  jand g18727(.dina(n18924), .dinb(n18881), .dout(n18983));
  jand g18728(.dina(n18933), .dinb(n18925), .dout(n18984));
  jor  g18729(.dina(n18984), .dinb(n18983), .dout(n18985));
  jand g18730(.dina(n18914), .dinb(n18884), .dout(n18986));
  jand g18731(.dina(n18923), .dinb(n18915), .dout(n18987));
  jor  g18732(.dina(n18987), .dinb(n18986), .dout(n18988));
  jand g18733(.dina(n18904), .dinb(n18887), .dout(n18989));
  jand g18734(.dina(n18913), .dinb(n18905), .dout(n18990));
  jor  g18735(.dina(n18990), .dinb(n18989), .dout(n18991));
  jand g18736(.dina(n18894), .dinb(n18891), .dout(n18992));
  jand g18737(.dina(n18903), .dinb(n18895), .dout(n18993));
  jor  g18738(.dina(n18993), .dinb(n18992), .dout(n18994));
  jand g18739(.dina(n10594), .dinb(b43 ), .dout(n18995));
  jand g18740(.dina(n10129), .dinb(b44 ), .dout(n18996));
  jor  g18741(.dina(n18996), .dinb(n18995), .dout(n18997));
  jxor g18742(.dina(n18997), .dinb(n18891), .dout(n18998));
  jor  g18743(.dina(n10134), .dinb(n6137), .dout(n18999));
  jor  g18744(.dina(n9849), .dinb(n5685), .dout(n19000));
  jor  g18745(.dina(n10137), .dinb(n5911), .dout(n19001));
  jor  g18746(.dina(n10132), .dinb(n6139), .dout(n19002));
  jand g18747(.dina(n19002), .dinb(n19001), .dout(n19003));
  jand g18748(.dina(n19003), .dinb(n19000), .dout(n19004));
  jand g18749(.dina(n19004), .dinb(n18999), .dout(n19005));
  jxor g18750(.dina(n19005), .dinb(n9559), .dout(n19006));
  jxor g18751(.dina(n19006), .dinb(n18998), .dout(n19007));
  jxor g18752(.dina(n19007), .dinb(n18994), .dout(n19008));
  jor  g18753(.dina(n9271), .dinb(n6844), .dout(n19009));
  jor  g18754(.dina(n9003), .dinb(n6366), .dout(n19010));
  jor  g18755(.dina(n9268), .dinb(n6846), .dout(n19011));
  jor  g18756(.dina(n9273), .dinb(n6605), .dout(n19012));
  jand g18757(.dina(n19012), .dinb(n19011), .dout(n19013));
  jand g18758(.dina(n19013), .dinb(n19010), .dout(n19014));
  jand g18759(.dina(n19014), .dinb(n19009), .dout(n19015));
  jxor g18760(.dina(n19015), .dinb(n8729), .dout(n19016));
  jxor g18761(.dina(n19016), .dinb(n19008), .dout(n19017));
  jxor g18762(.dina(n19017), .dinb(n18991), .dout(n19018));
  jor  g18763(.dina(n8457), .dinb(n7588), .dout(n19019));
  jor  g18764(.dina(n8185), .dinb(n7086), .dout(n19020));
  jor  g18765(.dina(n8459), .dinb(n7338), .dout(n19021));
  jor  g18766(.dina(n8454), .dinb(n7590), .dout(n19022));
  jand g18767(.dina(n19022), .dinb(n19021), .dout(n19023));
  jand g18768(.dina(n19023), .dinb(n19020), .dout(n19024));
  jand g18769(.dina(n19024), .dinb(n19019), .dout(n19025));
  jxor g18770(.dina(n19025), .dinb(n7929), .dout(n19026));
  jxor g18771(.dina(n19026), .dinb(n19018), .dout(n19027));
  jxor g18772(.dina(n19027), .dinb(n18988), .dout(n19028));
  jor  g18773(.dina(n8376), .dinb(n7660), .dout(n19029));
  jor  g18774(.dina(n7415), .dinb(n7846), .dout(n19030));
  jor  g18775(.dina(n7657), .dinb(n8111), .dout(n19031));
  jor  g18776(.dina(n7662), .dinb(n8378), .dout(n19032));
  jand g18777(.dina(n19032), .dinb(n19031), .dout(n19033));
  jand g18778(.dina(n19033), .dinb(n19030), .dout(n19034));
  jand g18779(.dina(n19034), .dinb(n19029), .dout(n19035));
  jxor g18780(.dina(n19035), .dinb(n7166), .dout(n19036));
  jxor g18781(.dina(n19036), .dinb(n19028), .dout(n19037));
  jxor g18782(.dina(n19037), .dinb(n18985), .dout(n19038));
  jor  g18783(.dina(n9193), .dinb(n6914), .dout(n19039));
  jor  g18784(.dina(n6673), .dinb(n8644), .dout(n19040));
  jor  g18785(.dina(n6911), .dinb(n8920), .dout(n19041));
  jor  g18786(.dina(n6916), .dinb(n9195), .dout(n19042));
  jand g18787(.dina(n19042), .dinb(n19041), .dout(n19043));
  jand g18788(.dina(n19043), .dinb(n19040), .dout(n19044));
  jand g18789(.dina(n19044), .dinb(n19039), .dout(n19045));
  jxor g18790(.dina(n19045), .dinb(n6443), .dout(n19046));
  jxor g18791(.dina(n19046), .dinb(n19038), .dout(n19047));
  jxor g18792(.dina(n19047), .dinb(n18982), .dout(n19048));
  jor  g18793(.dina(n10049), .dinb(n6207), .dout(n19049));
  jor  g18794(.dina(n5975), .dinb(n9475), .dout(n19050));
  jor  g18795(.dina(n6210), .dinb(n9759), .dout(n19051));
  jor  g18796(.dina(n6205), .dinb(n10051), .dout(n19052));
  jand g18797(.dina(n19052), .dinb(n19051), .dout(n19053));
  jand g18798(.dina(n19053), .dinb(n19050), .dout(n19054));
  jand g18799(.dina(n19054), .dinb(n19049), .dout(n19055));
  jxor g18800(.dina(n19055), .dinb(n5759), .dout(n19056));
  jxor g18801(.dina(n19056), .dinb(n19048), .dout(n19057));
  jxor g18802(.dina(n19057), .dinb(n18979), .dout(n19058));
  jxor g18803(.dina(n19058), .dinb(n18970), .dout(n19059));
  jnot g18804(.din(n19059), .dout(n19060));
  jxor g18805(.dina(n19060), .dinb(n18965), .dout(f107 ));
  jand g18806(.dina(n19058), .dinb(n18970), .dout(n19062));
  jnot g18807(.din(n19062), .dout(n19063));
  jor  g18808(.dina(n19060), .dinb(n18965), .dout(n19064));
  jand g18809(.dina(n19064), .dinb(n19063), .dout(n19065));
  jand g18810(.dina(n19047), .dinb(n18982), .dout(n19066));
  jand g18811(.dina(n19056), .dinb(n19048), .dout(n19067));
  jor  g18812(.dina(n19067), .dinb(n19066), .dout(n19068));
  jand g18813(.dina(n19037), .dinb(n18985), .dout(n19069));
  jand g18814(.dina(n19046), .dinb(n19038), .dout(n19070));
  jor  g18815(.dina(n19070), .dinb(n19069), .dout(n19071));
  jand g18816(.dina(n19027), .dinb(n18988), .dout(n19072));
  jand g18817(.dina(n19036), .dinb(n19028), .dout(n19073));
  jor  g18818(.dina(n19073), .dinb(n19072), .dout(n19074));
  jand g18819(.dina(n19017), .dinb(n18991), .dout(n19075));
  jand g18820(.dina(n19026), .dinb(n19018), .dout(n19076));
  jor  g18821(.dina(n19076), .dinb(n19075), .dout(n19077));
  jand g18822(.dina(n19007), .dinb(n18994), .dout(n19078));
  jand g18823(.dina(n19016), .dinb(n19008), .dout(n19079));
  jor  g18824(.dina(n19079), .dinb(n19078), .dout(n19080));
  jand g18825(.dina(n18997), .dinb(n18891), .dout(n19081));
  jand g18826(.dina(n19006), .dinb(n18998), .dout(n19082));
  jor  g18827(.dina(n19082), .dinb(n19081), .dout(n19083));
  jand g18828(.dina(n10594), .dinb(b44 ), .dout(n19084));
  jand g18829(.dina(n10129), .dinb(b45 ), .dout(n19085));
  jor  g18830(.dina(n19085), .dinb(n19084), .dout(n19086));
  jxor g18831(.dina(n19086), .dinb(n5111), .dout(n19087));
  jxor g18832(.dina(n19087), .dinb(n18890), .dout(n19088));
  jxor g18833(.dina(n19088), .dinb(n19083), .dout(n19089));
  jor  g18834(.dina(n10134), .dinb(n6364), .dout(n19090));
  jor  g18835(.dina(n9849), .dinb(n5911), .dout(n19091));
  jor  g18836(.dina(n10137), .dinb(n6139), .dout(n19092));
  jor  g18837(.dina(n10132), .dinb(n6366), .dout(n19093));
  jand g18838(.dina(n19093), .dinb(n19092), .dout(n19094));
  jand g18839(.dina(n19094), .dinb(n19091), .dout(n19095));
  jand g18840(.dina(n19095), .dinb(n19090), .dout(n19096));
  jxor g18841(.dina(n19096), .dinb(n9559), .dout(n19097));
  jxor g18842(.dina(n19097), .dinb(n19089), .dout(n19098));
  jor  g18843(.dina(n9271), .dinb(n7084), .dout(n19099));
  jor  g18844(.dina(n9003), .dinb(n6605), .dout(n19100));
  jor  g18845(.dina(n9273), .dinb(n6846), .dout(n19101));
  jor  g18846(.dina(n9268), .dinb(n7086), .dout(n19102));
  jand g18847(.dina(n19102), .dinb(n19101), .dout(n19103));
  jand g18848(.dina(n19103), .dinb(n19100), .dout(n19104));
  jand g18849(.dina(n19104), .dinb(n19099), .dout(n19105));
  jxor g18850(.dina(n19105), .dinb(n8729), .dout(n19106));
  jxor g18851(.dina(n19106), .dinb(n19098), .dout(n19107));
  jxor g18852(.dina(n19107), .dinb(n19080), .dout(n19108));
  jor  g18853(.dina(n8457), .dinb(n7844), .dout(n19109));
  jor  g18854(.dina(n8185), .dinb(n7338), .dout(n19110));
  jor  g18855(.dina(n8454), .dinb(n7846), .dout(n19111));
  jor  g18856(.dina(n8459), .dinb(n7590), .dout(n19112));
  jand g18857(.dina(n19112), .dinb(n19111), .dout(n19113));
  jand g18858(.dina(n19113), .dinb(n19110), .dout(n19114));
  jand g18859(.dina(n19114), .dinb(n19109), .dout(n19115));
  jxor g18860(.dina(n19115), .dinb(n7929), .dout(n19116));
  jxor g18861(.dina(n19116), .dinb(n19108), .dout(n19117));
  jxor g18862(.dina(n19117), .dinb(n19077), .dout(n19118));
  jor  g18863(.dina(n8642), .dinb(n7660), .dout(n19119));
  jor  g18864(.dina(n7415), .dinb(n8111), .dout(n19120));
  jor  g18865(.dina(n7662), .dinb(n8644), .dout(n19121));
  jor  g18866(.dina(n7657), .dinb(n8378), .dout(n19122));
  jand g18867(.dina(n19122), .dinb(n19121), .dout(n19123));
  jand g18868(.dina(n19123), .dinb(n19120), .dout(n19124));
  jand g18869(.dina(n19124), .dinb(n19119), .dout(n19125));
  jxor g18870(.dina(n19125), .dinb(n7166), .dout(n19126));
  jxor g18871(.dina(n19126), .dinb(n19118), .dout(n19127));
  jxor g18872(.dina(n19127), .dinb(n19074), .dout(n19128));
  jor  g18873(.dina(n9473), .dinb(n6914), .dout(n19129));
  jor  g18874(.dina(n6673), .dinb(n8920), .dout(n19130));
  jor  g18875(.dina(n6911), .dinb(n9195), .dout(n19131));
  jor  g18876(.dina(n6916), .dinb(n9475), .dout(n19132));
  jand g18877(.dina(n19132), .dinb(n19131), .dout(n19133));
  jand g18878(.dina(n19133), .dinb(n19130), .dout(n19134));
  jand g18879(.dina(n19134), .dinb(n19129), .dout(n19135));
  jxor g18880(.dina(n19135), .dinb(n6443), .dout(n19136));
  jxor g18881(.dina(n19136), .dinb(n19128), .dout(n19137));
  jxor g18882(.dina(n19137), .dinb(n19071), .dout(n19138));
  jor  g18883(.dina(n10521), .dinb(n6207), .dout(n19139));
  jor  g18884(.dina(n5975), .dinb(n9759), .dout(n19140));
  jor  g18885(.dina(n6210), .dinb(n10051), .dout(n19141));
  jor  g18886(.dina(n6205), .dinb(n10523), .dout(n19142));
  jand g18887(.dina(n19142), .dinb(n19141), .dout(n19143));
  jand g18888(.dina(n19143), .dinb(n19140), .dout(n19144));
  jand g18889(.dina(n19144), .dinb(n19139), .dout(n19145));
  jxor g18890(.dina(n19145), .dinb(n5759), .dout(n19146));
  jxor g18891(.dina(n19146), .dinb(n19138), .dout(n19147));
  jxor g18892(.dina(n19147), .dinb(n19068), .dout(n19148));
  jnot g18893(.din(n19148), .dout(n19149));
  jor  g18894(.dina(n18978), .dinb(n18974), .dout(n19150));
  jand g18895(.dina(n19057), .dinb(n18979), .dout(n19151));
  jnot g18896(.din(n19151), .dout(n19152));
  jand g18897(.dina(n19152), .dinb(n19150), .dout(n19153));
  jxor g18898(.dina(n19153), .dinb(n19149), .dout(n19154));
  jnot g18899(.din(n19154), .dout(n19155));
  jxor g18900(.dina(n19155), .dinb(n19065), .dout(f108 ));
  jand g18901(.dina(n19146), .dinb(n19138), .dout(n19157));
  jand g18902(.dina(n19147), .dinb(n19068), .dout(n19158));
  jor  g18903(.dina(n19158), .dinb(n19157), .dout(n19159));
  jand g18904(.dina(n19136), .dinb(n19128), .dout(n19160));
  jand g18905(.dina(n19137), .dinb(n19071), .dout(n19161));
  jor  g18906(.dina(n19161), .dinb(n19160), .dout(n19162));
  jnot g18907(.din(n19162), .dout(n19163));
  jor  g18908(.dina(n6210), .dinb(n10523), .dout(n19164));
  jor  g18909(.dina(n10813), .dinb(n6207), .dout(n19165));
  jor  g18910(.dina(n5975), .dinb(n10051), .dout(n19166));
  jand g18911(.dina(n19166), .dinb(n19165), .dout(n19167));
  jand g18912(.dina(n19167), .dinb(n19164), .dout(n19168));
  jxor g18913(.dina(n19168), .dinb(a47 ), .dout(n19169));
  jxor g18914(.dina(n19169), .dinb(n19163), .dout(n19170));
  jand g18915(.dina(n19126), .dinb(n19118), .dout(n19171));
  jand g18916(.dina(n19127), .dinb(n19074), .dout(n19172));
  jor  g18917(.dina(n19172), .dinb(n19171), .dout(n19173));
  jand g18918(.dina(n19116), .dinb(n19108), .dout(n19174));
  jand g18919(.dina(n19117), .dinb(n19077), .dout(n19175));
  jor  g18920(.dina(n19175), .dinb(n19174), .dout(n19176));
  jand g18921(.dina(n19106), .dinb(n19098), .dout(n19177));
  jand g18922(.dina(n19107), .dinb(n19080), .dout(n19178));
  jor  g18923(.dina(n19178), .dinb(n19177), .dout(n19179));
  jand g18924(.dina(n19088), .dinb(n19083), .dout(n19180));
  jand g18925(.dina(n19097), .dinb(n19089), .dout(n19181));
  jor  g18926(.dina(n19181), .dinb(n19180), .dout(n19182));
  jand g18927(.dina(n10594), .dinb(b45 ), .dout(n19183));
  jand g18928(.dina(n10129), .dinb(b46 ), .dout(n19184));
  jor  g18929(.dina(n19184), .dinb(n19183), .dout(n19185));
  jnot g18930(.din(n19185), .dout(n19186));
  jand g18931(.dina(n19086), .dinb(n5111), .dout(n19187));
  jand g18932(.dina(n19087), .dinb(n18890), .dout(n19188));
  jor  g18933(.dina(n19188), .dinb(n19187), .dout(n19189));
  jxor g18934(.dina(n19189), .dinb(n19186), .dout(n19190));
  jor  g18935(.dina(n10134), .dinb(n6603), .dout(n19191));
  jor  g18936(.dina(n9849), .dinb(n6139), .dout(n19192));
  jor  g18937(.dina(n10137), .dinb(n6366), .dout(n19193));
  jor  g18938(.dina(n10132), .dinb(n6605), .dout(n19194));
  jand g18939(.dina(n19194), .dinb(n19193), .dout(n19195));
  jand g18940(.dina(n19195), .dinb(n19192), .dout(n19196));
  jand g18941(.dina(n19196), .dinb(n19191), .dout(n19197));
  jxor g18942(.dina(n19197), .dinb(n9559), .dout(n19198));
  jxor g18943(.dina(n19198), .dinb(n19190), .dout(n19199));
  jxor g18944(.dina(n19199), .dinb(n19182), .dout(n19200));
  jor  g18945(.dina(n9271), .dinb(n7336), .dout(n19201));
  jor  g18946(.dina(n9003), .dinb(n6846), .dout(n19202));
  jor  g18947(.dina(n9273), .dinb(n7086), .dout(n19203));
  jor  g18948(.dina(n9268), .dinb(n7338), .dout(n19204));
  jand g18949(.dina(n19204), .dinb(n19203), .dout(n19205));
  jand g18950(.dina(n19205), .dinb(n19202), .dout(n19206));
  jand g18951(.dina(n19206), .dinb(n19201), .dout(n19207));
  jxor g18952(.dina(n19207), .dinb(n8729), .dout(n19208));
  jxor g18953(.dina(n19208), .dinb(n19200), .dout(n19209));
  jxor g18954(.dina(n19209), .dinb(n19179), .dout(n19210));
  jor  g18955(.dina(n8109), .dinb(n8457), .dout(n19211));
  jor  g18956(.dina(n8185), .dinb(n7590), .dout(n19212));
  jor  g18957(.dina(n8459), .dinb(n7846), .dout(n19213));
  jor  g18958(.dina(n8454), .dinb(n8111), .dout(n19214));
  jand g18959(.dina(n19214), .dinb(n19213), .dout(n19215));
  jand g18960(.dina(n19215), .dinb(n19212), .dout(n19216));
  jand g18961(.dina(n19216), .dinb(n19211), .dout(n19217));
  jxor g18962(.dina(n19217), .dinb(n7929), .dout(n19218));
  jxor g18963(.dina(n19218), .dinb(n19210), .dout(n19219));
  jxor g18964(.dina(n19219), .dinb(n19176), .dout(n19220));
  jor  g18965(.dina(n8918), .dinb(n7660), .dout(n19221));
  jor  g18966(.dina(n7415), .dinb(n8378), .dout(n19222));
  jor  g18967(.dina(n7662), .dinb(n8920), .dout(n19223));
  jor  g18968(.dina(n7657), .dinb(n8644), .dout(n19224));
  jand g18969(.dina(n19224), .dinb(n19223), .dout(n19225));
  jand g18970(.dina(n19225), .dinb(n19222), .dout(n19226));
  jand g18971(.dina(n19226), .dinb(n19221), .dout(n19227));
  jxor g18972(.dina(n19227), .dinb(n7166), .dout(n19228));
  jxor g18973(.dina(n19228), .dinb(n19220), .dout(n19229));
  jxor g18974(.dina(n19229), .dinb(n19173), .dout(n19230));
  jor  g18975(.dina(n9757), .dinb(n6914), .dout(n19231));
  jor  g18976(.dina(n6673), .dinb(n9195), .dout(n19232));
  jor  g18977(.dina(n6911), .dinb(n9475), .dout(n19233));
  jor  g18978(.dina(n6916), .dinb(n9759), .dout(n19234));
  jand g18979(.dina(n19234), .dinb(n19233), .dout(n19235));
  jand g18980(.dina(n19235), .dinb(n19232), .dout(n19236));
  jand g18981(.dina(n19236), .dinb(n19231), .dout(n19237));
  jxor g18982(.dina(n19237), .dinb(n6443), .dout(n19238));
  jxor g18983(.dina(n19238), .dinb(n19230), .dout(n19239));
  jxor g18984(.dina(n19239), .dinb(n19170), .dout(n19240));
  jxor g18985(.dina(n19240), .dinb(n19159), .dout(n19241));
  jnot g18986(.din(n19241), .dout(n19242));
  jor  g18987(.dina(n19153), .dinb(n19149), .dout(n19243));
  jor  g18988(.dina(n19155), .dinb(n19065), .dout(n19244));
  jand g18989(.dina(n19244), .dinb(n19243), .dout(n19245));
  jxor g18990(.dina(n19245), .dinb(n19242), .dout(f109 ));
  jor  g18991(.dina(n19169), .dinb(n19163), .dout(n19247));
  jand g18992(.dina(n19239), .dinb(n19170), .dout(n19248));
  jnot g18993(.din(n19248), .dout(n19249));
  jand g18994(.dina(n19249), .dinb(n19247), .dout(n19250));
  jnot g18995(.din(n19250), .dout(n19251));
  jand g18996(.dina(n19229), .dinb(n19173), .dout(n19252));
  jand g18997(.dina(n19238), .dinb(n19230), .dout(n19253));
  jor  g18998(.dina(n19253), .dinb(n19252), .dout(n19254));
  jnot g18999(.din(n19254), .dout(n19255));
  jand g19000(.dina(n5976), .dinb(b63 ), .dout(n19256));
  jand g19001(.dina(n10832), .dinb(n5748), .dout(n19257));
  jor  g19002(.dina(n19257), .dinb(n19256), .dout(n19258));
  jxor g19003(.dina(n19258), .dinb(n5759), .dout(n19259));
  jxor g19004(.dina(n19259), .dinb(n19255), .dout(n19260));
  jand g19005(.dina(n19219), .dinb(n19176), .dout(n19261));
  jand g19006(.dina(n19228), .dinb(n19220), .dout(n19262));
  jor  g19007(.dina(n19262), .dinb(n19261), .dout(n19263));
  jand g19008(.dina(n19209), .dinb(n19179), .dout(n19264));
  jand g19009(.dina(n19218), .dinb(n19210), .dout(n19265));
  jor  g19010(.dina(n19265), .dinb(n19264), .dout(n19266));
  jand g19011(.dina(n19199), .dinb(n19182), .dout(n19267));
  jand g19012(.dina(n19208), .dinb(n19200), .dout(n19268));
  jor  g19013(.dina(n19268), .dinb(n19267), .dout(n19269));
  jand g19014(.dina(n19189), .dinb(n19186), .dout(n19270));
  jand g19015(.dina(n19198), .dinb(n19190), .dout(n19271));
  jor  g19016(.dina(n19271), .dinb(n19270), .dout(n19272));
  jand g19017(.dina(n10594), .dinb(b46 ), .dout(n19273));
  jand g19018(.dina(n10129), .dinb(b47 ), .dout(n19274));
  jor  g19019(.dina(n19274), .dinb(n19273), .dout(n19275));
  jnot g19020(.din(n19275), .dout(n19276));
  jxor g19021(.dina(n19276), .dinb(n19185), .dout(n19277));
  jxor g19022(.dina(n19277), .dinb(n19272), .dout(n19278));
  jor  g19023(.dina(n10134), .dinb(n6844), .dout(n19279));
  jor  g19024(.dina(n9849), .dinb(n6366), .dout(n19280));
  jor  g19025(.dina(n10132), .dinb(n6846), .dout(n19281));
  jor  g19026(.dina(n10137), .dinb(n6605), .dout(n19282));
  jand g19027(.dina(n19282), .dinb(n19281), .dout(n19283));
  jand g19028(.dina(n19283), .dinb(n19280), .dout(n19284));
  jand g19029(.dina(n19284), .dinb(n19279), .dout(n19285));
  jxor g19030(.dina(n19285), .dinb(n9559), .dout(n19286));
  jxor g19031(.dina(n19286), .dinb(n19278), .dout(n19287));
  jor  g19032(.dina(n9271), .dinb(n7588), .dout(n19288));
  jor  g19033(.dina(n9003), .dinb(n7086), .dout(n19289));
  jor  g19034(.dina(n9268), .dinb(n7590), .dout(n19290));
  jor  g19035(.dina(n9273), .dinb(n7338), .dout(n19291));
  jand g19036(.dina(n19291), .dinb(n19290), .dout(n19292));
  jand g19037(.dina(n19292), .dinb(n19289), .dout(n19293));
  jand g19038(.dina(n19293), .dinb(n19288), .dout(n19294));
  jxor g19039(.dina(n19294), .dinb(n8729), .dout(n19295));
  jxor g19040(.dina(n19295), .dinb(n19287), .dout(n19296));
  jxor g19041(.dina(n19296), .dinb(n19269), .dout(n19297));
  jor  g19042(.dina(n8376), .dinb(n8457), .dout(n19298));
  jor  g19043(.dina(n8185), .dinb(n7846), .dout(n19299));
  jor  g19044(.dina(n8459), .dinb(n8111), .dout(n19300));
  jor  g19045(.dina(n8454), .dinb(n8378), .dout(n19301));
  jand g19046(.dina(n19301), .dinb(n19300), .dout(n19302));
  jand g19047(.dina(n19302), .dinb(n19299), .dout(n19303));
  jand g19048(.dina(n19303), .dinb(n19298), .dout(n19304));
  jxor g19049(.dina(n19304), .dinb(n7929), .dout(n19305));
  jxor g19050(.dina(n19305), .dinb(n19297), .dout(n19306));
  jxor g19051(.dina(n19306), .dinb(n19266), .dout(n19307));
  jor  g19052(.dina(n9193), .dinb(n7660), .dout(n19308));
  jor  g19053(.dina(n7415), .dinb(n8644), .dout(n19309));
  jor  g19054(.dina(n7662), .dinb(n9195), .dout(n19310));
  jor  g19055(.dina(n7657), .dinb(n8920), .dout(n19311));
  jand g19056(.dina(n19311), .dinb(n19310), .dout(n19312));
  jand g19057(.dina(n19312), .dinb(n19309), .dout(n19313));
  jand g19058(.dina(n19313), .dinb(n19308), .dout(n19314));
  jxor g19059(.dina(n19314), .dinb(n7166), .dout(n19315));
  jxor g19060(.dina(n19315), .dinb(n19307), .dout(n19316));
  jxor g19061(.dina(n19316), .dinb(n19263), .dout(n19317));
  jor  g19062(.dina(n10049), .dinb(n6914), .dout(n19318));
  jor  g19063(.dina(n6673), .dinb(n9475), .dout(n19319));
  jor  g19064(.dina(n6916), .dinb(n10051), .dout(n19320));
  jor  g19065(.dina(n6911), .dinb(n9759), .dout(n19321));
  jand g19066(.dina(n19321), .dinb(n19320), .dout(n19322));
  jand g19067(.dina(n19322), .dinb(n19319), .dout(n19323));
  jand g19068(.dina(n19323), .dinb(n19318), .dout(n19324));
  jxor g19069(.dina(n19324), .dinb(n6443), .dout(n19325));
  jxor g19070(.dina(n19325), .dinb(n19317), .dout(n19326));
  jxor g19071(.dina(n19326), .dinb(n19260), .dout(n19327));
  jxor g19072(.dina(n19327), .dinb(n19251), .dout(n19328));
  jnot g19073(.din(n19328), .dout(n19329));
  jand g19074(.dina(n19240), .dinb(n19159), .dout(n19330));
  jnot g19075(.din(n19330), .dout(n19331));
  jor  g19076(.dina(n19245), .dinb(n19242), .dout(n19332));
  jand g19077(.dina(n19332), .dinb(n19331), .dout(n19333));
  jxor g19078(.dina(n19333), .dinb(n19329), .dout(f110 ));
  jand g19079(.dina(n19316), .dinb(n19263), .dout(n19335));
  jand g19080(.dina(n19325), .dinb(n19317), .dout(n19336));
  jor  g19081(.dina(n19336), .dinb(n19335), .dout(n19337));
  jand g19082(.dina(n19306), .dinb(n19266), .dout(n19338));
  jand g19083(.dina(n19315), .dinb(n19307), .dout(n19339));
  jor  g19084(.dina(n19339), .dinb(n19338), .dout(n19340));
  jand g19085(.dina(n19296), .dinb(n19269), .dout(n19341));
  jand g19086(.dina(n19305), .dinb(n19297), .dout(n19342));
  jor  g19087(.dina(n19342), .dinb(n19341), .dout(n19343));
  jand g19088(.dina(n19286), .dinb(n19278), .dout(n19344));
  jand g19089(.dina(n19295), .dinb(n19287), .dout(n19345));
  jor  g19090(.dina(n19345), .dinb(n19344), .dout(n19346));
  jand g19091(.dina(n19276), .dinb(n19185), .dout(n19347));
  jand g19092(.dina(n19277), .dinb(n19272), .dout(n19348));
  jor  g19093(.dina(n19348), .dinb(n19347), .dout(n19349));
  jand g19094(.dina(n10594), .dinb(b47 ), .dout(n19350));
  jand g19095(.dina(n10129), .dinb(b48 ), .dout(n19351));
  jor  g19096(.dina(n19351), .dinb(n19350), .dout(n19352));
  jxor g19097(.dina(n19275), .dinb(n5759), .dout(n19353));
  jxor g19098(.dina(n19353), .dinb(n19352), .dout(n19354));
  jor  g19099(.dina(n10134), .dinb(n7084), .dout(n19355));
  jor  g19100(.dina(n9849), .dinb(n6605), .dout(n19356));
  jor  g19101(.dina(n10137), .dinb(n6846), .dout(n19357));
  jor  g19102(.dina(n10132), .dinb(n7086), .dout(n19358));
  jand g19103(.dina(n19358), .dinb(n19357), .dout(n19359));
  jand g19104(.dina(n19359), .dinb(n19356), .dout(n19360));
  jand g19105(.dina(n19360), .dinb(n19355), .dout(n19361));
  jxor g19106(.dina(n19361), .dinb(n9559), .dout(n19362));
  jxor g19107(.dina(n19362), .dinb(n19354), .dout(n19363));
  jxor g19108(.dina(n19363), .dinb(n19349), .dout(n19364));
  jor  g19109(.dina(n9271), .dinb(n7844), .dout(n19365));
  jor  g19110(.dina(n9003), .dinb(n7338), .dout(n19366));
  jor  g19111(.dina(n9273), .dinb(n7590), .dout(n19367));
  jor  g19112(.dina(n9268), .dinb(n7846), .dout(n19368));
  jand g19113(.dina(n19368), .dinb(n19367), .dout(n19369));
  jand g19114(.dina(n19369), .dinb(n19366), .dout(n19370));
  jand g19115(.dina(n19370), .dinb(n19365), .dout(n19371));
  jxor g19116(.dina(n19371), .dinb(n8729), .dout(n19372));
  jxor g19117(.dina(n19372), .dinb(n19364), .dout(n19373));
  jxor g19118(.dina(n19373), .dinb(n19346), .dout(n19374));
  jor  g19119(.dina(n8642), .dinb(n8457), .dout(n19375));
  jor  g19120(.dina(n8185), .dinb(n8111), .dout(n19376));
  jor  g19121(.dina(n8454), .dinb(n8644), .dout(n19377));
  jor  g19122(.dina(n8459), .dinb(n8378), .dout(n19378));
  jand g19123(.dina(n19378), .dinb(n19377), .dout(n19379));
  jand g19124(.dina(n19379), .dinb(n19376), .dout(n19380));
  jand g19125(.dina(n19380), .dinb(n19375), .dout(n19381));
  jxor g19126(.dina(n19381), .dinb(n7929), .dout(n19382));
  jxor g19127(.dina(n19382), .dinb(n19374), .dout(n19383));
  jxor g19128(.dina(n19383), .dinb(n19343), .dout(n19384));
  jor  g19129(.dina(n9473), .dinb(n7660), .dout(n19385));
  jor  g19130(.dina(n7415), .dinb(n8920), .dout(n19386));
  jor  g19131(.dina(n7657), .dinb(n9195), .dout(n19387));
  jor  g19132(.dina(n7662), .dinb(n9475), .dout(n19388));
  jand g19133(.dina(n19388), .dinb(n19387), .dout(n19389));
  jand g19134(.dina(n19389), .dinb(n19386), .dout(n19390));
  jand g19135(.dina(n19390), .dinb(n19385), .dout(n19391));
  jxor g19136(.dina(n19391), .dinb(n7166), .dout(n19392));
  jxor g19137(.dina(n19392), .dinb(n19384), .dout(n19393));
  jxor g19138(.dina(n19393), .dinb(n19340), .dout(n19394));
  jor  g19139(.dina(n10521), .dinb(n6914), .dout(n19395));
  jor  g19140(.dina(n6673), .dinb(n9759), .dout(n19396));
  jor  g19141(.dina(n6916), .dinb(n10523), .dout(n19397));
  jor  g19142(.dina(n6911), .dinb(n10051), .dout(n19398));
  jand g19143(.dina(n19398), .dinb(n19397), .dout(n19399));
  jand g19144(.dina(n19399), .dinb(n19396), .dout(n19400));
  jand g19145(.dina(n19400), .dinb(n19395), .dout(n19401));
  jxor g19146(.dina(n19401), .dinb(n6443), .dout(n19402));
  jxor g19147(.dina(n19402), .dinb(n19394), .dout(n19403));
  jxor g19148(.dina(n19403), .dinb(n19337), .dout(n19404));
  jnot g19149(.din(n19404), .dout(n19405));
  jor  g19150(.dina(n19259), .dinb(n19255), .dout(n19406));
  jand g19151(.dina(n19326), .dinb(n19260), .dout(n19407));
  jnot g19152(.din(n19407), .dout(n19408));
  jand g19153(.dina(n19408), .dinb(n19406), .dout(n19409));
  jxor g19154(.dina(n19409), .dinb(n19405), .dout(n19410));
  jnot g19155(.din(n19410), .dout(n19411));
  jand g19156(.dina(n19327), .dinb(n19251), .dout(n19412));
  jnot g19157(.din(n19412), .dout(n19413));
  jor  g19158(.dina(n19333), .dinb(n19329), .dout(n19414));
  jand g19159(.dina(n19414), .dinb(n19413), .dout(n19415));
  jxor g19160(.dina(n19415), .dinb(n19411), .dout(f111 ));
  jand g19161(.dina(n19402), .dinb(n19394), .dout(n19417));
  jand g19162(.dina(n19403), .dinb(n19337), .dout(n19418));
  jor  g19163(.dina(n19418), .dinb(n19417), .dout(n19419));
  jand g19164(.dina(n19392), .dinb(n19384), .dout(n19420));
  jand g19165(.dina(n19393), .dinb(n19340), .dout(n19421));
  jor  g19166(.dina(n19421), .dinb(n19420), .dout(n19422));
  jand g19167(.dina(n19382), .dinb(n19374), .dout(n19423));
  jand g19168(.dina(n19383), .dinb(n19343), .dout(n19424));
  jor  g19169(.dina(n19424), .dinb(n19423), .dout(n19425));
  jand g19170(.dina(n19372), .dinb(n19364), .dout(n19426));
  jand g19171(.dina(n19373), .dinb(n19346), .dout(n19427));
  jor  g19172(.dina(n19427), .dinb(n19426), .dout(n19428));
  jand g19173(.dina(n19362), .dinb(n19354), .dout(n19429));
  jand g19174(.dina(n19363), .dinb(n19349), .dout(n19430));
  jor  g19175(.dina(n19430), .dinb(n19429), .dout(n19431));
  jand g19176(.dina(n10594), .dinb(b48 ), .dout(n19432));
  jand g19177(.dina(n10129), .dinb(b49 ), .dout(n19433));
  jor  g19178(.dina(n19433), .dinb(n19432), .dout(n19434));
  jnot g19179(.din(n19434), .dout(n19435));
  jand g19180(.dina(n19275), .dinb(n5759), .dout(n19436));
  jand g19181(.dina(n19353), .dinb(n19352), .dout(n19437));
  jor  g19182(.dina(n19437), .dinb(n19436), .dout(n19438));
  jxor g19183(.dina(n19438), .dinb(n19435), .dout(n19439));
  jor  g19184(.dina(n10134), .dinb(n7336), .dout(n19440));
  jor  g19185(.dina(n9849), .dinb(n6846), .dout(n19441));
  jor  g19186(.dina(n10137), .dinb(n7086), .dout(n19442));
  jor  g19187(.dina(n10132), .dinb(n7338), .dout(n19443));
  jand g19188(.dina(n19443), .dinb(n19442), .dout(n19444));
  jand g19189(.dina(n19444), .dinb(n19441), .dout(n19445));
  jand g19190(.dina(n19445), .dinb(n19440), .dout(n19446));
  jxor g19191(.dina(n19446), .dinb(n9559), .dout(n19447));
  jxor g19192(.dina(n19447), .dinb(n19439), .dout(n19448));
  jxor g19193(.dina(n19448), .dinb(n19431), .dout(n19449));
  jor  g19194(.dina(n9271), .dinb(n8109), .dout(n19450));
  jor  g19195(.dina(n9003), .dinb(n7590), .dout(n19451));
  jor  g19196(.dina(n9273), .dinb(n7846), .dout(n19452));
  jor  g19197(.dina(n9268), .dinb(n8111), .dout(n19453));
  jand g19198(.dina(n19453), .dinb(n19452), .dout(n19454));
  jand g19199(.dina(n19454), .dinb(n19451), .dout(n19455));
  jand g19200(.dina(n19455), .dinb(n19450), .dout(n19456));
  jxor g19201(.dina(n19456), .dinb(n8729), .dout(n19457));
  jxor g19202(.dina(n19457), .dinb(n19449), .dout(n19458));
  jxor g19203(.dina(n19458), .dinb(n19428), .dout(n19459));
  jor  g19204(.dina(n8918), .dinb(n8457), .dout(n19460));
  jor  g19205(.dina(n8185), .dinb(n8378), .dout(n19461));
  jor  g19206(.dina(n8454), .dinb(n8920), .dout(n19462));
  jor  g19207(.dina(n8459), .dinb(n8644), .dout(n19463));
  jand g19208(.dina(n19463), .dinb(n19462), .dout(n19464));
  jand g19209(.dina(n19464), .dinb(n19461), .dout(n19465));
  jand g19210(.dina(n19465), .dinb(n19460), .dout(n19466));
  jxor g19211(.dina(n19466), .dinb(n7929), .dout(n19467));
  jxor g19212(.dina(n19467), .dinb(n19459), .dout(n19468));
  jxor g19213(.dina(n19468), .dinb(n19425), .dout(n19469));
  jor  g19214(.dina(n9757), .dinb(n7660), .dout(n19470));
  jor  g19215(.dina(n7415), .dinb(n9195), .dout(n19471));
  jor  g19216(.dina(n7657), .dinb(n9475), .dout(n19472));
  jor  g19217(.dina(n7662), .dinb(n9759), .dout(n19473));
  jand g19218(.dina(n19473), .dinb(n19472), .dout(n19474));
  jand g19219(.dina(n19474), .dinb(n19471), .dout(n19475));
  jand g19220(.dina(n19475), .dinb(n19470), .dout(n19476));
  jxor g19221(.dina(n19476), .dinb(n7166), .dout(n19477));
  jxor g19222(.dina(n19477), .dinb(n19469), .dout(n19478));
  jxor g19223(.dina(n19478), .dinb(n19422), .dout(n19479));
  jnot g19224(.din(n19479), .dout(n19480));
  jor  g19225(.dina(n10813), .dinb(n6914), .dout(n19481));
  jor  g19226(.dina(n6673), .dinb(n10051), .dout(n19482));
  jor  g19227(.dina(n6911), .dinb(n10523), .dout(n19483));
  jand g19228(.dina(n19483), .dinb(n19482), .dout(n19484));
  jand g19229(.dina(n19484), .dinb(n19481), .dout(n19485));
  jxor g19230(.dina(n19485), .dinb(a50 ), .dout(n19486));
  jxor g19231(.dina(n19486), .dinb(n19480), .dout(n19487));
  jxor g19232(.dina(n19487), .dinb(n19419), .dout(n19488));
  jnot g19233(.din(n19488), .dout(n19489));
  jor  g19234(.dina(n19409), .dinb(n19405), .dout(n19490));
  jor  g19235(.dina(n19415), .dinb(n19411), .dout(n19491));
  jand g19236(.dina(n19491), .dinb(n19490), .dout(n19492));
  jxor g19237(.dina(n19492), .dinb(n19489), .dout(f112 ));
  jand g19238(.dina(n19478), .dinb(n19422), .dout(n19494));
  jnot g19239(.din(n19494), .dout(n19495));
  jor  g19240(.dina(n19486), .dinb(n19480), .dout(n19496));
  jand g19241(.dina(n19496), .dinb(n19495), .dout(n19497));
  jnot g19242(.din(n19497), .dout(n19498));
  jand g19243(.dina(n19468), .dinb(n19425), .dout(n19499));
  jand g19244(.dina(n19477), .dinb(n19469), .dout(n19500));
  jor  g19245(.dina(n19500), .dinb(n19499), .dout(n19501));
  jnot g19246(.din(n19501), .dout(n19502));
  jand g19247(.dina(n6674), .dinb(b63 ), .dout(n19503));
  jand g19248(.dina(n10832), .dinb(n6435), .dout(n19504));
  jor  g19249(.dina(n19504), .dinb(n19503), .dout(n19505));
  jxor g19250(.dina(n19505), .dinb(n6443), .dout(n19506));
  jxor g19251(.dina(n19506), .dinb(n19502), .dout(n19507));
  jand g19252(.dina(n19458), .dinb(n19428), .dout(n19508));
  jand g19253(.dina(n19467), .dinb(n19459), .dout(n19509));
  jor  g19254(.dina(n19509), .dinb(n19508), .dout(n19510));
  jand g19255(.dina(n19448), .dinb(n19431), .dout(n19511));
  jand g19256(.dina(n19457), .dinb(n19449), .dout(n19512));
  jor  g19257(.dina(n19512), .dinb(n19511), .dout(n19513));
  jand g19258(.dina(n19438), .dinb(n19435), .dout(n19514));
  jand g19259(.dina(n19447), .dinb(n19439), .dout(n19515));
  jor  g19260(.dina(n19515), .dinb(n19514), .dout(n19516));
  jand g19261(.dina(n10594), .dinb(b49 ), .dout(n19517));
  jand g19262(.dina(n10129), .dinb(b50 ), .dout(n19518));
  jor  g19263(.dina(n19518), .dinb(n19517), .dout(n19519));
  jxor g19264(.dina(n19519), .dinb(n19435), .dout(n19520));
  jor  g19265(.dina(n10134), .dinb(n7588), .dout(n19521));
  jor  g19266(.dina(n9849), .dinb(n7086), .dout(n19522));
  jor  g19267(.dina(n10132), .dinb(n7590), .dout(n19523));
  jor  g19268(.dina(n10137), .dinb(n7338), .dout(n19524));
  jand g19269(.dina(n19524), .dinb(n19523), .dout(n19525));
  jand g19270(.dina(n19525), .dinb(n19522), .dout(n19526));
  jand g19271(.dina(n19526), .dinb(n19521), .dout(n19527));
  jxor g19272(.dina(n19527), .dinb(n9559), .dout(n19528));
  jxor g19273(.dina(n19528), .dinb(n19520), .dout(n19529));
  jxor g19274(.dina(n19529), .dinb(n19516), .dout(n19530));
  jor  g19275(.dina(n9271), .dinb(n8376), .dout(n19531));
  jor  g19276(.dina(n9003), .dinb(n7846), .dout(n19532));
  jor  g19277(.dina(n9268), .dinb(n8378), .dout(n19533));
  jor  g19278(.dina(n9273), .dinb(n8111), .dout(n19534));
  jand g19279(.dina(n19534), .dinb(n19533), .dout(n19535));
  jand g19280(.dina(n19535), .dinb(n19532), .dout(n19536));
  jand g19281(.dina(n19536), .dinb(n19531), .dout(n19537));
  jxor g19282(.dina(n19537), .dinb(n8729), .dout(n19538));
  jxor g19283(.dina(n19538), .dinb(n19530), .dout(n19539));
  jxor g19284(.dina(n19539), .dinb(n19513), .dout(n19540));
  jor  g19285(.dina(n9193), .dinb(n8457), .dout(n19541));
  jor  g19286(.dina(n8185), .dinb(n8644), .dout(n19542));
  jor  g19287(.dina(n8454), .dinb(n9195), .dout(n19543));
  jor  g19288(.dina(n8459), .dinb(n8920), .dout(n19544));
  jand g19289(.dina(n19544), .dinb(n19543), .dout(n19545));
  jand g19290(.dina(n19545), .dinb(n19542), .dout(n19546));
  jand g19291(.dina(n19546), .dinb(n19541), .dout(n19547));
  jxor g19292(.dina(n19547), .dinb(n7929), .dout(n19548));
  jxor g19293(.dina(n19548), .dinb(n19540), .dout(n19549));
  jxor g19294(.dina(n19549), .dinb(n19510), .dout(n19550));
  jor  g19295(.dina(n10049), .dinb(n7660), .dout(n19551));
  jor  g19296(.dina(n7415), .dinb(n9475), .dout(n19552));
  jor  g19297(.dina(n7657), .dinb(n9759), .dout(n19553));
  jor  g19298(.dina(n7662), .dinb(n10051), .dout(n19554));
  jand g19299(.dina(n19554), .dinb(n19553), .dout(n19555));
  jand g19300(.dina(n19555), .dinb(n19552), .dout(n19556));
  jand g19301(.dina(n19556), .dinb(n19551), .dout(n19557));
  jxor g19302(.dina(n19557), .dinb(n7166), .dout(n19558));
  jxor g19303(.dina(n19558), .dinb(n19550), .dout(n19559));
  jxor g19304(.dina(n19559), .dinb(n19507), .dout(n19560));
  jxor g19305(.dina(n19560), .dinb(n19498), .dout(n19561));
  jnot g19306(.din(n19561), .dout(n19562));
  jand g19307(.dina(n19487), .dinb(n19419), .dout(n19563));
  jnot g19308(.din(n19563), .dout(n19564));
  jor  g19309(.dina(n19492), .dinb(n19489), .dout(n19565));
  jand g19310(.dina(n19565), .dinb(n19564), .dout(n19566));
  jxor g19311(.dina(n19566), .dinb(n19562), .dout(f113 ));
  jand g19312(.dina(n19549), .dinb(n19510), .dout(n19568));
  jand g19313(.dina(n19558), .dinb(n19550), .dout(n19569));
  jor  g19314(.dina(n19569), .dinb(n19568), .dout(n19570));
  jand g19315(.dina(n19539), .dinb(n19513), .dout(n19571));
  jand g19316(.dina(n19548), .dinb(n19540), .dout(n19572));
  jor  g19317(.dina(n19572), .dinb(n19571), .dout(n19573));
  jand g19318(.dina(n19529), .dinb(n19516), .dout(n19574));
  jand g19319(.dina(n19538), .dinb(n19530), .dout(n19575));
  jor  g19320(.dina(n19575), .dinb(n19574), .dout(n19576));
  jand g19321(.dina(n19519), .dinb(n19435), .dout(n19577));
  jand g19322(.dina(n19528), .dinb(n19520), .dout(n19578));
  jor  g19323(.dina(n19578), .dinb(n19577), .dout(n19579));
  jand g19324(.dina(n10594), .dinb(b50 ), .dout(n19580));
  jand g19325(.dina(n10129), .dinb(b51 ), .dout(n19581));
  jor  g19326(.dina(n19581), .dinb(n19580), .dout(n19582));
  jxor g19327(.dina(n19582), .dinb(n6443), .dout(n19583));
  jxor g19328(.dina(n19583), .dinb(n19434), .dout(n19584));
  jxor g19329(.dina(n19584), .dinb(n19579), .dout(n19585));
  jor  g19330(.dina(n10134), .dinb(n7844), .dout(n19586));
  jor  g19331(.dina(n9849), .dinb(n7338), .dout(n19587));
  jor  g19332(.dina(n10137), .dinb(n7590), .dout(n19588));
  jor  g19333(.dina(n10132), .dinb(n7846), .dout(n19589));
  jand g19334(.dina(n19589), .dinb(n19588), .dout(n19590));
  jand g19335(.dina(n19590), .dinb(n19587), .dout(n19591));
  jand g19336(.dina(n19591), .dinb(n19586), .dout(n19592));
  jxor g19337(.dina(n19592), .dinb(n9559), .dout(n19593));
  jxor g19338(.dina(n19593), .dinb(n19585), .dout(n19594));
  jor  g19339(.dina(n9271), .dinb(n8642), .dout(n19595));
  jor  g19340(.dina(n9003), .dinb(n8111), .dout(n19596));
  jor  g19341(.dina(n9273), .dinb(n8378), .dout(n19597));
  jor  g19342(.dina(n9268), .dinb(n8644), .dout(n19598));
  jand g19343(.dina(n19598), .dinb(n19597), .dout(n19599));
  jand g19344(.dina(n19599), .dinb(n19596), .dout(n19600));
  jand g19345(.dina(n19600), .dinb(n19595), .dout(n19601));
  jxor g19346(.dina(n19601), .dinb(n8729), .dout(n19602));
  jxor g19347(.dina(n19602), .dinb(n19594), .dout(n19603));
  jxor g19348(.dina(n19603), .dinb(n19576), .dout(n19604));
  jor  g19349(.dina(n9473), .dinb(n8457), .dout(n19605));
  jor  g19350(.dina(n8185), .dinb(n8920), .dout(n19606));
  jor  g19351(.dina(n8454), .dinb(n9475), .dout(n19607));
  jor  g19352(.dina(n8459), .dinb(n9195), .dout(n19608));
  jand g19353(.dina(n19608), .dinb(n19607), .dout(n19609));
  jand g19354(.dina(n19609), .dinb(n19606), .dout(n19610));
  jand g19355(.dina(n19610), .dinb(n19605), .dout(n19611));
  jxor g19356(.dina(n19611), .dinb(n7929), .dout(n19612));
  jxor g19357(.dina(n19612), .dinb(n19604), .dout(n19613));
  jxor g19358(.dina(n19613), .dinb(n19573), .dout(n19614));
  jor  g19359(.dina(n10521), .dinb(n7660), .dout(n19615));
  jor  g19360(.dina(n7415), .dinb(n9759), .dout(n19616));
  jor  g19361(.dina(n7662), .dinb(n10523), .dout(n19617));
  jor  g19362(.dina(n7657), .dinb(n10051), .dout(n19618));
  jand g19363(.dina(n19618), .dinb(n19617), .dout(n19619));
  jand g19364(.dina(n19619), .dinb(n19616), .dout(n19620));
  jand g19365(.dina(n19620), .dinb(n19615), .dout(n19621));
  jxor g19366(.dina(n19621), .dinb(n7166), .dout(n19622));
  jxor g19367(.dina(n19622), .dinb(n19614), .dout(n19623));
  jxor g19368(.dina(n19623), .dinb(n19570), .dout(n19624));
  jnot g19369(.din(n19624), .dout(n19625));
  jor  g19370(.dina(n19506), .dinb(n19502), .dout(n19626));
  jand g19371(.dina(n19559), .dinb(n19507), .dout(n19627));
  jnot g19372(.din(n19627), .dout(n19628));
  jand g19373(.dina(n19628), .dinb(n19626), .dout(n19629));
  jxor g19374(.dina(n19629), .dinb(n19625), .dout(n19630));
  jnot g19375(.din(n19630), .dout(n19631));
  jand g19376(.dina(n19560), .dinb(n19498), .dout(n19632));
  jnot g19377(.din(n19632), .dout(n19633));
  jor  g19378(.dina(n19566), .dinb(n19562), .dout(n19634));
  jand g19379(.dina(n19634), .dinb(n19633), .dout(n19635));
  jxor g19380(.dina(n19635), .dinb(n19631), .dout(f114 ));
  jand g19381(.dina(n19622), .dinb(n19614), .dout(n19637));
  jand g19382(.dina(n19623), .dinb(n19570), .dout(n19638));
  jor  g19383(.dina(n19638), .dinb(n19637), .dout(n19639));
  jand g19384(.dina(n19612), .dinb(n19604), .dout(n19640));
  jand g19385(.dina(n19613), .dinb(n19573), .dout(n19641));
  jor  g19386(.dina(n19641), .dinb(n19640), .dout(n19642));
  jand g19387(.dina(n19602), .dinb(n19594), .dout(n19643));
  jand g19388(.dina(n19603), .dinb(n19576), .dout(n19644));
  jor  g19389(.dina(n19644), .dinb(n19643), .dout(n19645));
  jand g19390(.dina(n19584), .dinb(n19579), .dout(n19646));
  jand g19391(.dina(n19593), .dinb(n19585), .dout(n19647));
  jor  g19392(.dina(n19647), .dinb(n19646), .dout(n19648));
  jand g19393(.dina(n10594), .dinb(b51 ), .dout(n19649));
  jand g19394(.dina(n10129), .dinb(b52 ), .dout(n19650));
  jor  g19395(.dina(n19650), .dinb(n19649), .dout(n19651));
  jnot g19396(.din(n19651), .dout(n19652));
  jand g19397(.dina(n19582), .dinb(n6443), .dout(n19653));
  jand g19398(.dina(n19583), .dinb(n19434), .dout(n19654));
  jor  g19399(.dina(n19654), .dinb(n19653), .dout(n19655));
  jxor g19400(.dina(n19655), .dinb(n19652), .dout(n19656));
  jor  g19401(.dina(n10134), .dinb(n8109), .dout(n19657));
  jor  g19402(.dina(n9849), .dinb(n7590), .dout(n19658));
  jor  g19403(.dina(n10132), .dinb(n8111), .dout(n19659));
  jor  g19404(.dina(n10137), .dinb(n7846), .dout(n19660));
  jand g19405(.dina(n19660), .dinb(n19659), .dout(n19661));
  jand g19406(.dina(n19661), .dinb(n19658), .dout(n19662));
  jand g19407(.dina(n19662), .dinb(n19657), .dout(n19663));
  jxor g19408(.dina(n19663), .dinb(n9559), .dout(n19664));
  jxor g19409(.dina(n19664), .dinb(n19656), .dout(n19665));
  jxor g19410(.dina(n19665), .dinb(n19648), .dout(n19666));
  jor  g19411(.dina(n8918), .dinb(n9271), .dout(n19667));
  jor  g19412(.dina(n9003), .dinb(n8378), .dout(n19668));
  jor  g19413(.dina(n9273), .dinb(n8644), .dout(n19669));
  jor  g19414(.dina(n9268), .dinb(n8920), .dout(n19670));
  jand g19415(.dina(n19670), .dinb(n19669), .dout(n19671));
  jand g19416(.dina(n19671), .dinb(n19668), .dout(n19672));
  jand g19417(.dina(n19672), .dinb(n19667), .dout(n19673));
  jxor g19418(.dina(n19673), .dinb(n8729), .dout(n19674));
  jxor g19419(.dina(n19674), .dinb(n19666), .dout(n19675));
  jxor g19420(.dina(n19675), .dinb(n19645), .dout(n19676));
  jor  g19421(.dina(n9757), .dinb(n8457), .dout(n19677));
  jor  g19422(.dina(n8185), .dinb(n9195), .dout(n19678));
  jor  g19423(.dina(n8459), .dinb(n9475), .dout(n19679));
  jor  g19424(.dina(n8454), .dinb(n9759), .dout(n19680));
  jand g19425(.dina(n19680), .dinb(n19679), .dout(n19681));
  jand g19426(.dina(n19681), .dinb(n19678), .dout(n19682));
  jand g19427(.dina(n19682), .dinb(n19677), .dout(n19683));
  jxor g19428(.dina(n19683), .dinb(n7929), .dout(n19684));
  jxor g19429(.dina(n19684), .dinb(n19676), .dout(n19685));
  jxor g19430(.dina(n19685), .dinb(n19642), .dout(n19686));
  jnot g19431(.din(n19686), .dout(n19687));
  jor  g19432(.dina(n10813), .dinb(n7660), .dout(n19688));
  jor  g19433(.dina(n7415), .dinb(n10051), .dout(n19689));
  jor  g19434(.dina(n7657), .dinb(n10523), .dout(n19690));
  jand g19435(.dina(n19690), .dinb(n19689), .dout(n19691));
  jand g19436(.dina(n19691), .dinb(n19688), .dout(n19692));
  jxor g19437(.dina(n19692), .dinb(a53 ), .dout(n19693));
  jxor g19438(.dina(n19693), .dinb(n19687), .dout(n19694));
  jxor g19439(.dina(n19694), .dinb(n19639), .dout(n19695));
  jnot g19440(.din(n19695), .dout(n19696));
  jor  g19441(.dina(n19629), .dinb(n19625), .dout(n19697));
  jor  g19442(.dina(n19635), .dinb(n19631), .dout(n19698));
  jand g19443(.dina(n19698), .dinb(n19697), .dout(n19699));
  jxor g19444(.dina(n19699), .dinb(n19696), .dout(f115 ));
  jand g19445(.dina(n19685), .dinb(n19642), .dout(n19701));
  jnot g19446(.din(n19701), .dout(n19702));
  jor  g19447(.dina(n19693), .dinb(n19687), .dout(n19703));
  jand g19448(.dina(n19703), .dinb(n19702), .dout(n19704));
  jnot g19449(.din(n19704), .dout(n19705));
  jand g19450(.dina(n19675), .dinb(n19645), .dout(n19706));
  jand g19451(.dina(n19684), .dinb(n19676), .dout(n19707));
  jor  g19452(.dina(n19707), .dinb(n19706), .dout(n19708));
  jnot g19453(.din(n19708), .dout(n19709));
  jand g19454(.dina(n7416), .dinb(b63 ), .dout(n19710));
  jand g19455(.dina(n10832), .dinb(n7155), .dout(n19711));
  jor  g19456(.dina(n19711), .dinb(n19710), .dout(n19712));
  jxor g19457(.dina(n19712), .dinb(n7166), .dout(n19713));
  jxor g19458(.dina(n19713), .dinb(n19709), .dout(n19714));
  jand g19459(.dina(n19665), .dinb(n19648), .dout(n19715));
  jand g19460(.dina(n19674), .dinb(n19666), .dout(n19716));
  jor  g19461(.dina(n19716), .dinb(n19715), .dout(n19717));
  jand g19462(.dina(n19655), .dinb(n19652), .dout(n19718));
  jand g19463(.dina(n19664), .dinb(n19656), .dout(n19719));
  jor  g19464(.dina(n19719), .dinb(n19718), .dout(n19720));
  jand g19465(.dina(n10594), .dinb(b52 ), .dout(n19721));
  jand g19466(.dina(n10129), .dinb(b53 ), .dout(n19722));
  jor  g19467(.dina(n19722), .dinb(n19721), .dout(n19723));
  jnot g19468(.din(n19723), .dout(n19724));
  jxor g19469(.dina(n19724), .dinb(n19651), .dout(n19725));
  jxor g19470(.dina(n19725), .dinb(n19720), .dout(n19726));
  jor  g19471(.dina(n10134), .dinb(n8376), .dout(n19727));
  jor  g19472(.dina(n9849), .dinb(n7846), .dout(n19728));
  jor  g19473(.dina(n10137), .dinb(n8111), .dout(n19729));
  jor  g19474(.dina(n10132), .dinb(n8378), .dout(n19730));
  jand g19475(.dina(n19730), .dinb(n19729), .dout(n19731));
  jand g19476(.dina(n19731), .dinb(n19728), .dout(n19732));
  jand g19477(.dina(n19732), .dinb(n19727), .dout(n19733));
  jxor g19478(.dina(n19733), .dinb(n9559), .dout(n19734));
  jxor g19479(.dina(n19734), .dinb(n19726), .dout(n19735));
  jor  g19480(.dina(n9193), .dinb(n9271), .dout(n19736));
  jor  g19481(.dina(n9003), .dinb(n8644), .dout(n19737));
  jor  g19482(.dina(n9273), .dinb(n8920), .dout(n19738));
  jor  g19483(.dina(n9268), .dinb(n9195), .dout(n19739));
  jand g19484(.dina(n19739), .dinb(n19738), .dout(n19740));
  jand g19485(.dina(n19740), .dinb(n19737), .dout(n19741));
  jand g19486(.dina(n19741), .dinb(n19736), .dout(n19742));
  jxor g19487(.dina(n19742), .dinb(n8729), .dout(n19743));
  jxor g19488(.dina(n19743), .dinb(n19735), .dout(n19744));
  jxor g19489(.dina(n19744), .dinb(n19717), .dout(n19745));
  jor  g19490(.dina(n10049), .dinb(n8457), .dout(n19746));
  jor  g19491(.dina(n8185), .dinb(n9475), .dout(n19747));
  jor  g19492(.dina(n8454), .dinb(n10051), .dout(n19748));
  jor  g19493(.dina(n8459), .dinb(n9759), .dout(n19749));
  jand g19494(.dina(n19749), .dinb(n19748), .dout(n19750));
  jand g19495(.dina(n19750), .dinb(n19747), .dout(n19751));
  jand g19496(.dina(n19751), .dinb(n19746), .dout(n19752));
  jxor g19497(.dina(n19752), .dinb(n7929), .dout(n19753));
  jxor g19498(.dina(n19753), .dinb(n19745), .dout(n19754));
  jxor g19499(.dina(n19754), .dinb(n19714), .dout(n19755));
  jxor g19500(.dina(n19755), .dinb(n19705), .dout(n19756));
  jnot g19501(.din(n19756), .dout(n19757));
  jand g19502(.dina(n19694), .dinb(n19639), .dout(n19758));
  jnot g19503(.din(n19758), .dout(n19759));
  jor  g19504(.dina(n19699), .dinb(n19696), .dout(n19760));
  jand g19505(.dina(n19760), .dinb(n19759), .dout(n19761));
  jxor g19506(.dina(n19761), .dinb(n19757), .dout(f116 ));
  jand g19507(.dina(n19755), .dinb(n19705), .dout(n19763));
  jnot g19508(.din(n19763), .dout(n19764));
  jor  g19509(.dina(n19761), .dinb(n19757), .dout(n19765));
  jand g19510(.dina(n19765), .dinb(n19764), .dout(n19766));
  jor  g19511(.dina(n19713), .dinb(n19709), .dout(n19767));
  jand g19512(.dina(n19754), .dinb(n19714), .dout(n19768));
  jnot g19513(.din(n19768), .dout(n19769));
  jand g19514(.dina(n19769), .dinb(n19767), .dout(n19770));
  jnot g19515(.din(n19770), .dout(n19771));
  jand g19516(.dina(n19744), .dinb(n19717), .dout(n19772));
  jand g19517(.dina(n19753), .dinb(n19745), .dout(n19773));
  jor  g19518(.dina(n19773), .dinb(n19772), .dout(n19774));
  jor  g19519(.dina(n10521), .dinb(n8457), .dout(n19775));
  jor  g19520(.dina(n8185), .dinb(n9759), .dout(n19776));
  jor  g19521(.dina(n8459), .dinb(n10051), .dout(n19777));
  jor  g19522(.dina(n8454), .dinb(n10523), .dout(n19778));
  jand g19523(.dina(n19778), .dinb(n19777), .dout(n19779));
  jand g19524(.dina(n19779), .dinb(n19776), .dout(n19780));
  jand g19525(.dina(n19780), .dinb(n19775), .dout(n19781));
  jxor g19526(.dina(n19781), .dinb(n7929), .dout(n19782));
  jxor g19527(.dina(n19782), .dinb(n19774), .dout(n19783));
  jand g19528(.dina(n19734), .dinb(n19726), .dout(n19784));
  jand g19529(.dina(n19743), .dinb(n19735), .dout(n19785));
  jor  g19530(.dina(n19785), .dinb(n19784), .dout(n19786));
  jand g19531(.dina(n19724), .dinb(n19651), .dout(n19787));
  jand g19532(.dina(n19725), .dinb(n19720), .dout(n19788));
  jor  g19533(.dina(n19788), .dinb(n19787), .dout(n19789));
  jand g19534(.dina(n10594), .dinb(b53 ), .dout(n19790));
  jand g19535(.dina(n10129), .dinb(b54 ), .dout(n19791));
  jor  g19536(.dina(n19791), .dinb(n19790), .dout(n19792));
  jxor g19537(.dina(n19723), .dinb(n7166), .dout(n19793));
  jxor g19538(.dina(n19793), .dinb(n19792), .dout(n19794));
  jor  g19539(.dina(n10134), .dinb(n8642), .dout(n19795));
  jor  g19540(.dina(n9849), .dinb(n8111), .dout(n19796));
  jor  g19541(.dina(n10137), .dinb(n8378), .dout(n19797));
  jor  g19542(.dina(n10132), .dinb(n8644), .dout(n19798));
  jand g19543(.dina(n19798), .dinb(n19797), .dout(n19799));
  jand g19544(.dina(n19799), .dinb(n19796), .dout(n19800));
  jand g19545(.dina(n19800), .dinb(n19795), .dout(n19801));
  jxor g19546(.dina(n19801), .dinb(n9559), .dout(n19802));
  jxor g19547(.dina(n19802), .dinb(n19794), .dout(n19803));
  jxor g19548(.dina(n19803), .dinb(n19789), .dout(n19804));
  jor  g19549(.dina(n9473), .dinb(n9271), .dout(n19805));
  jor  g19550(.dina(n9003), .dinb(n8920), .dout(n19806));
  jor  g19551(.dina(n9268), .dinb(n9475), .dout(n19807));
  jor  g19552(.dina(n9273), .dinb(n9195), .dout(n19808));
  jand g19553(.dina(n19808), .dinb(n19807), .dout(n19809));
  jand g19554(.dina(n19809), .dinb(n19806), .dout(n19810));
  jand g19555(.dina(n19810), .dinb(n19805), .dout(n19811));
  jxor g19556(.dina(n19811), .dinb(n8729), .dout(n19812));
  jxor g19557(.dina(n19812), .dinb(n19804), .dout(n19813));
  jxor g19558(.dina(n19813), .dinb(n19786), .dout(n19814));
  jxor g19559(.dina(n19814), .dinb(n19783), .dout(n19815));
  jxor g19560(.dina(n19815), .dinb(n19771), .dout(n19816));
  jnot g19561(.din(n19816), .dout(n19817));
  jxor g19562(.dina(n19817), .dinb(n19766), .dout(f117 ));
  jand g19563(.dina(n19815), .dinb(n19771), .dout(n19819));
  jnot g19564(.din(n19819), .dout(n19820));
  jor  g19565(.dina(n19817), .dinb(n19766), .dout(n19821));
  jand g19566(.dina(n19821), .dinb(n19820), .dout(n19822));
  jand g19567(.dina(n19782), .dinb(n19774), .dout(n19823));
  jand g19568(.dina(n19814), .dinb(n19783), .dout(n19824));
  jor  g19569(.dina(n19824), .dinb(n19823), .dout(n19825));
  jand g19570(.dina(n19812), .dinb(n19804), .dout(n19826));
  jand g19571(.dina(n19813), .dinb(n19786), .dout(n19827));
  jor  g19572(.dina(n19827), .dinb(n19826), .dout(n19828));
  jand g19573(.dina(n19802), .dinb(n19794), .dout(n19829));
  jand g19574(.dina(n19803), .dinb(n19789), .dout(n19830));
  jor  g19575(.dina(n19830), .dinb(n19829), .dout(n19831));
  jand g19576(.dina(n10594), .dinb(b54 ), .dout(n19832));
  jand g19577(.dina(n10129), .dinb(b55 ), .dout(n19833));
  jor  g19578(.dina(n19833), .dinb(n19832), .dout(n19834));
  jnot g19579(.din(n19834), .dout(n19835));
  jand g19580(.dina(n19723), .dinb(n7166), .dout(n19836));
  jand g19581(.dina(n19793), .dinb(n19792), .dout(n19837));
  jor  g19582(.dina(n19837), .dinb(n19836), .dout(n19838));
  jxor g19583(.dina(n19838), .dinb(n19835), .dout(n19839));
  jor  g19584(.dina(n10134), .dinb(n8918), .dout(n19840));
  jor  g19585(.dina(n9849), .dinb(n8378), .dout(n19841));
  jor  g19586(.dina(n10137), .dinb(n8644), .dout(n19842));
  jor  g19587(.dina(n10132), .dinb(n8920), .dout(n19843));
  jand g19588(.dina(n19843), .dinb(n19842), .dout(n19844));
  jand g19589(.dina(n19844), .dinb(n19841), .dout(n19845));
  jand g19590(.dina(n19845), .dinb(n19840), .dout(n19846));
  jxor g19591(.dina(n19846), .dinb(n9559), .dout(n19847));
  jxor g19592(.dina(n19847), .dinb(n19839), .dout(n19848));
  jxor g19593(.dina(n19848), .dinb(n19831), .dout(n19849));
  jor  g19594(.dina(n9757), .dinb(n9271), .dout(n19850));
  jor  g19595(.dina(n9003), .dinb(n9195), .dout(n19851));
  jor  g19596(.dina(n9268), .dinb(n9759), .dout(n19852));
  jor  g19597(.dina(n9273), .dinb(n9475), .dout(n19853));
  jand g19598(.dina(n19853), .dinb(n19852), .dout(n19854));
  jand g19599(.dina(n19854), .dinb(n19851), .dout(n19855));
  jand g19600(.dina(n19855), .dinb(n19850), .dout(n19856));
  jxor g19601(.dina(n19856), .dinb(n8729), .dout(n19857));
  jxor g19602(.dina(n19857), .dinb(n19849), .dout(n19858));
  jxor g19603(.dina(n19858), .dinb(n19828), .dout(n19859));
  jor  g19604(.dina(n10813), .dinb(n8457), .dout(n19860));
  jor  g19605(.dina(n8185), .dinb(n10051), .dout(n19861));
  jor  g19606(.dina(n8459), .dinb(n10523), .dout(n19862));
  jand g19607(.dina(n19862), .dinb(n19861), .dout(n19863));
  jand g19608(.dina(n19863), .dinb(n19860), .dout(n19864));
  jxor g19609(.dina(n19864), .dinb(n7929), .dout(n19865));
  jxor g19610(.dina(n19865), .dinb(n19859), .dout(n19866));
  jxor g19611(.dina(n19866), .dinb(n19825), .dout(n19867));
  jnot g19612(.din(n19867), .dout(n19868));
  jxor g19613(.dina(n19868), .dinb(n19822), .dout(f118 ));
  jand g19614(.dina(n19858), .dinb(n19828), .dout(n19870));
  jand g19615(.dina(n19865), .dinb(n19859), .dout(n19871));
  jor  g19616(.dina(n19871), .dinb(n19870), .dout(n19872));
  jand g19617(.dina(n19848), .dinb(n19831), .dout(n19873));
  jand g19618(.dina(n19857), .dinb(n19849), .dout(n19874));
  jor  g19619(.dina(n19874), .dinb(n19873), .dout(n19875));
  jnot g19620(.din(n19875), .dout(n19876));
  jand g19621(.dina(n8186), .dinb(b63 ), .dout(n19877));
  jand g19622(.dina(n10832), .dinb(n7918), .dout(n19878));
  jor  g19623(.dina(n19878), .dinb(n19877), .dout(n19879));
  jxor g19624(.dina(n19879), .dinb(n7929), .dout(n19880));
  jxor g19625(.dina(n19880), .dinb(n19876), .dout(n19881));
  jand g19626(.dina(n19838), .dinb(n19835), .dout(n19882));
  jand g19627(.dina(n19847), .dinb(n19839), .dout(n19883));
  jor  g19628(.dina(n19883), .dinb(n19882), .dout(n19884));
  jand g19629(.dina(n10594), .dinb(b55 ), .dout(n19885));
  jand g19630(.dina(n10129), .dinb(b56 ), .dout(n19886));
  jor  g19631(.dina(n19886), .dinb(n19885), .dout(n19887));
  jxor g19632(.dina(n19887), .dinb(n19835), .dout(n19888));
  jor  g19633(.dina(n10134), .dinb(n9193), .dout(n19889));
  jor  g19634(.dina(n9849), .dinb(n8644), .dout(n19890));
  jor  g19635(.dina(n10132), .dinb(n9195), .dout(n19891));
  jor  g19636(.dina(n10137), .dinb(n8920), .dout(n19892));
  jand g19637(.dina(n19892), .dinb(n19891), .dout(n19893));
  jand g19638(.dina(n19893), .dinb(n19890), .dout(n19894));
  jand g19639(.dina(n19894), .dinb(n19889), .dout(n19895));
  jxor g19640(.dina(n19895), .dinb(n9559), .dout(n19896));
  jxor g19641(.dina(n19896), .dinb(n19888), .dout(n19897));
  jxor g19642(.dina(n19897), .dinb(n19884), .dout(n19898));
  jor  g19643(.dina(n10049), .dinb(n9271), .dout(n19899));
  jor  g19644(.dina(n9003), .dinb(n9475), .dout(n19900));
  jor  g19645(.dina(n9273), .dinb(n9759), .dout(n19901));
  jor  g19646(.dina(n9268), .dinb(n10051), .dout(n19902));
  jand g19647(.dina(n19902), .dinb(n19901), .dout(n19903));
  jand g19648(.dina(n19903), .dinb(n19900), .dout(n19904));
  jand g19649(.dina(n19904), .dinb(n19899), .dout(n19905));
  jxor g19650(.dina(n19905), .dinb(n8729), .dout(n19906));
  jxor g19651(.dina(n19906), .dinb(n19898), .dout(n19907));
  jxor g19652(.dina(n19907), .dinb(n19881), .dout(n19908));
  jxor g19653(.dina(n19908), .dinb(n19872), .dout(n19909));
  jnot g19654(.din(n19909), .dout(n19910));
  jand g19655(.dina(n19866), .dinb(n19825), .dout(n19911));
  jnot g19656(.din(n19911), .dout(n19912));
  jor  g19657(.dina(n19868), .dinb(n19822), .dout(n19913));
  jand g19658(.dina(n19913), .dinb(n19912), .dout(n19914));
  jxor g19659(.dina(n19914), .dinb(n19910), .dout(f119 ));
  jor  g19660(.dina(n19880), .dinb(n19876), .dout(n19916));
  jand g19661(.dina(n19907), .dinb(n19881), .dout(n19917));
  jnot g19662(.din(n19917), .dout(n19918));
  jand g19663(.dina(n19918), .dinb(n19916), .dout(n19919));
  jnot g19664(.din(n19919), .dout(n19920));
  jand g19665(.dina(n19897), .dinb(n19884), .dout(n19921));
  jand g19666(.dina(n19906), .dinb(n19898), .dout(n19922));
  jor  g19667(.dina(n19922), .dinb(n19921), .dout(n19923));
  jor  g19668(.dina(n10521), .dinb(n9271), .dout(n19924));
  jor  g19669(.dina(n9003), .dinb(n9759), .dout(n19925));
  jor  g19670(.dina(n9273), .dinb(n10051), .dout(n19926));
  jor  g19671(.dina(n9268), .dinb(n10523), .dout(n19927));
  jand g19672(.dina(n19927), .dinb(n19926), .dout(n19928));
  jand g19673(.dina(n19928), .dinb(n19925), .dout(n19929));
  jand g19674(.dina(n19929), .dinb(n19924), .dout(n19930));
  jxor g19675(.dina(n19930), .dinb(n8729), .dout(n19931));
  jxor g19676(.dina(n19931), .dinb(n19923), .dout(n19932));
  jand g19677(.dina(n19887), .dinb(n19835), .dout(n19933));
  jand g19678(.dina(n19896), .dinb(n19888), .dout(n19934));
  jor  g19679(.dina(n19934), .dinb(n19933), .dout(n19935));
  jand g19680(.dina(n10594), .dinb(b56 ), .dout(n19936));
  jand g19681(.dina(n10129), .dinb(b57 ), .dout(n19937));
  jor  g19682(.dina(n19937), .dinb(n19936), .dout(n19938));
  jxor g19683(.dina(n19938), .dinb(n7929), .dout(n19939));
  jxor g19684(.dina(n19939), .dinb(n19834), .dout(n19940));
  jxor g19685(.dina(n19940), .dinb(n19935), .dout(n19941));
  jor  g19686(.dina(n10134), .dinb(n9473), .dout(n19942));
  jor  g19687(.dina(n9849), .dinb(n8920), .dout(n19943));
  jor  g19688(.dina(n10137), .dinb(n9195), .dout(n19944));
  jor  g19689(.dina(n10132), .dinb(n9475), .dout(n19945));
  jand g19690(.dina(n19945), .dinb(n19944), .dout(n19946));
  jand g19691(.dina(n19946), .dinb(n19943), .dout(n19947));
  jand g19692(.dina(n19947), .dinb(n19942), .dout(n19948));
  jxor g19693(.dina(n19948), .dinb(n9559), .dout(n19949));
  jxor g19694(.dina(n19949), .dinb(n19941), .dout(n19950));
  jxor g19695(.dina(n19950), .dinb(n19932), .dout(n19951));
  jxor g19696(.dina(n19951), .dinb(n19920), .dout(n19952));
  jnot g19697(.din(n19952), .dout(n19953));
  jand g19698(.dina(n19908), .dinb(n19872), .dout(n19954));
  jnot g19699(.din(n19954), .dout(n19955));
  jor  g19700(.dina(n19914), .dinb(n19910), .dout(n19956));
  jand g19701(.dina(n19956), .dinb(n19955), .dout(n19957));
  jxor g19702(.dina(n19957), .dinb(n19953), .dout(f120 ));
  jand g19703(.dina(n19931), .dinb(n19923), .dout(n19959));
  jand g19704(.dina(n19950), .dinb(n19932), .dout(n19960));
  jor  g19705(.dina(n19960), .dinb(n19959), .dout(n19961));
  jand g19706(.dina(n19940), .dinb(n19935), .dout(n19962));
  jand g19707(.dina(n19949), .dinb(n19941), .dout(n19963));
  jor  g19708(.dina(n19963), .dinb(n19962), .dout(n19964));
  jand g19709(.dina(n10594), .dinb(b57 ), .dout(n19965));
  jand g19710(.dina(n10129), .dinb(b58 ), .dout(n19966));
  jor  g19711(.dina(n19966), .dinb(n19965), .dout(n19967));
  jnot g19712(.din(n19967), .dout(n19968));
  jand g19713(.dina(n19938), .dinb(n7929), .dout(n19969));
  jand g19714(.dina(n19939), .dinb(n19834), .dout(n19970));
  jor  g19715(.dina(n19970), .dinb(n19969), .dout(n19971));
  jxor g19716(.dina(n19971), .dinb(n19968), .dout(n19972));
  jor  g19717(.dina(n9757), .dinb(n10134), .dout(n19973));
  jor  g19718(.dina(n9849), .dinb(n9195), .dout(n19974));
  jor  g19719(.dina(n10137), .dinb(n9475), .dout(n19975));
  jor  g19720(.dina(n10132), .dinb(n9759), .dout(n19976));
  jand g19721(.dina(n19976), .dinb(n19975), .dout(n19977));
  jand g19722(.dina(n19977), .dinb(n19974), .dout(n19978));
  jand g19723(.dina(n19978), .dinb(n19973), .dout(n19979));
  jxor g19724(.dina(n19979), .dinb(n9559), .dout(n19980));
  jxor g19725(.dina(n19980), .dinb(n19972), .dout(n19981));
  jxor g19726(.dina(n19981), .dinb(n19964), .dout(n19982));
  jnot g19727(.din(n19982), .dout(n19983));
  jor  g19728(.dina(n9273), .dinb(n10523), .dout(n19984));
  jor  g19729(.dina(n10813), .dinb(n9271), .dout(n19985));
  jor  g19730(.dina(n9003), .dinb(n10051), .dout(n19986));
  jand g19731(.dina(n19986), .dinb(n19985), .dout(n19987));
  jand g19732(.dina(n19987), .dinb(n19984), .dout(n19988));
  jxor g19733(.dina(n19988), .dinb(a59 ), .dout(n19989));
  jxor g19734(.dina(n19989), .dinb(n19983), .dout(n19990));
  jxor g19735(.dina(n19990), .dinb(n19961), .dout(n19991));
  jnot g19736(.din(n19991), .dout(n19992));
  jand g19737(.dina(n19951), .dinb(n19920), .dout(n19993));
  jnot g19738(.din(n19993), .dout(n19994));
  jor  g19739(.dina(n19957), .dinb(n19953), .dout(n19995));
  jand g19740(.dina(n19995), .dinb(n19994), .dout(n19996));
  jxor g19741(.dina(n19996), .dinb(n19992), .dout(f121 ));
  jand g19742(.dina(n19990), .dinb(n19961), .dout(n19998));
  jnot g19743(.din(n19998), .dout(n19999));
  jor  g19744(.dina(n19996), .dinb(n19992), .dout(n20000));
  jand g19745(.dina(n20000), .dinb(n19999), .dout(n20001));
  jand g19746(.dina(n19981), .dinb(n19964), .dout(n20002));
  jnot g19747(.din(n20002), .dout(n20003));
  jor  g19748(.dina(n19989), .dinb(n19983), .dout(n20004));
  jand g19749(.dina(n20004), .dinb(n20003), .dout(n20005));
  jnot g19750(.din(n20005), .dout(n20006));
  jor  g19751(.dina(n10049), .dinb(n10134), .dout(n20007));
  jor  g19752(.dina(n9849), .dinb(n9475), .dout(n20008));
  jor  g19753(.dina(n10132), .dinb(n10051), .dout(n20009));
  jor  g19754(.dina(n10137), .dinb(n9759), .dout(n20010));
  jand g19755(.dina(n20010), .dinb(n20009), .dout(n20011));
  jand g19756(.dina(n20011), .dinb(n20008), .dout(n20012));
  jand g19757(.dina(n20012), .dinb(n20007), .dout(n20013));
  jxor g19758(.dina(n20013), .dinb(n9559), .dout(n20014));
  jnot g19759(.din(n20014), .dout(n20015));
  jand g19760(.dina(n9004), .dinb(b63 ), .dout(n20016));
  jand g19761(.dina(n10832), .dinb(n8718), .dout(n20017));
  jor  g19762(.dina(n20017), .dinb(n20016), .dout(n20018));
  jxor g19763(.dina(n20018), .dinb(n8729), .dout(n20019));
  jxor g19764(.dina(n20019), .dinb(n20015), .dout(n20020));
  jand g19765(.dina(n19971), .dinb(n19968), .dout(n20021));
  jand g19766(.dina(n19980), .dinb(n19972), .dout(n20022));
  jor  g19767(.dina(n20022), .dinb(n20021), .dout(n20023));
  jand g19768(.dina(n10594), .dinb(b58 ), .dout(n20024));
  jand g19769(.dina(n10129), .dinb(b59 ), .dout(n20025));
  jor  g19770(.dina(n20025), .dinb(n20024), .dout(n20026));
  jnot g19771(.din(n20026), .dout(n20027));
  jxor g19772(.dina(n20027), .dinb(n19967), .dout(n20028));
  jxor g19773(.dina(n20028), .dinb(n20023), .dout(n20029));
  jxor g19774(.dina(n20029), .dinb(n20020), .dout(n20030));
  jxor g19775(.dina(n20030), .dinb(n20006), .dout(n20031));
  jnot g19776(.din(n20031), .dout(n20032));
  jxor g19777(.dina(n20032), .dinb(n20001), .dout(f122 ));
  jand g19778(.dina(n20030), .dinb(n20006), .dout(n20034));
  jnot g19779(.din(n20034), .dout(n20035));
  jor  g19780(.dina(n20032), .dinb(n20001), .dout(n20036));
  jand g19781(.dina(n20036), .dinb(n20035), .dout(n20037));
  jor  g19782(.dina(n20019), .dinb(n20015), .dout(n20038));
  jand g19783(.dina(n20029), .dinb(n20020), .dout(n20039));
  jnot g19784(.din(n20039), .dout(n20040));
  jand g19785(.dina(n20040), .dinb(n20038), .dout(n20041));
  jnot g19786(.din(n20041), .dout(n20042));
  jand g19787(.dina(n20027), .dinb(n19967), .dout(n20043));
  jand g19788(.dina(n20028), .dinb(n20023), .dout(n20044));
  jor  g19789(.dina(n20044), .dinb(n20043), .dout(n20045));
  jand g19790(.dina(n10594), .dinb(b59 ), .dout(n20046));
  jand g19791(.dina(n10129), .dinb(b60 ), .dout(n20047));
  jor  g19792(.dina(n20047), .dinb(n20046), .dout(n20048));
  jxor g19793(.dina(n20026), .dinb(n8729), .dout(n20049));
  jxor g19794(.dina(n20049), .dinb(n20048), .dout(n20050));
  jor  g19795(.dina(n10521), .dinb(n10134), .dout(n20051));
  jor  g19796(.dina(n9849), .dinb(n9759), .dout(n20052));
  jor  g19797(.dina(n10132), .dinb(n10523), .dout(n20053));
  jor  g19798(.dina(n10137), .dinb(n10051), .dout(n20054));
  jand g19799(.dina(n20054), .dinb(n20053), .dout(n20055));
  jand g19800(.dina(n20055), .dinb(n20052), .dout(n20056));
  jand g19801(.dina(n20056), .dinb(n20051), .dout(n20057));
  jxor g19802(.dina(n20057), .dinb(n9559), .dout(n20058));
  jxor g19803(.dina(n20058), .dinb(n20050), .dout(n20059));
  jxor g19804(.dina(n20059), .dinb(n20045), .dout(n20060));
  jxor g19805(.dina(n20060), .dinb(n20042), .dout(n20061));
  jnot g19806(.din(n20061), .dout(n20062));
  jxor g19807(.dina(n20062), .dinb(n20037), .dout(f123 ));
  jand g19808(.dina(n20060), .dinb(n20042), .dout(n20064));
  jnot g19809(.din(n20064), .dout(n20065));
  jor  g19810(.dina(n20062), .dinb(n20037), .dout(n20066));
  jand g19811(.dina(n20066), .dinb(n20065), .dout(n20067));
  jand g19812(.dina(n20058), .dinb(n20050), .dout(n20068));
  jand g19813(.dina(n20059), .dinb(n20045), .dout(n20069));
  jor  g19814(.dina(n20069), .dinb(n20068), .dout(n20070));
  jand g19815(.dina(n10594), .dinb(b60 ), .dout(n20071));
  jand g19816(.dina(n10129), .dinb(b61 ), .dout(n20072));
  jor  g19817(.dina(n20072), .dinb(n20071), .dout(n20073));
  jnot g19818(.din(n20073), .dout(n20074));
  jand g19819(.dina(n20026), .dinb(n8729), .dout(n20075));
  jand g19820(.dina(n20049), .dinb(n20048), .dout(n20076));
  jor  g19821(.dina(n20076), .dinb(n20075), .dout(n20077));
  jxor g19822(.dina(n20077), .dinb(n20074), .dout(n20078));
  jnot g19823(.din(n20078), .dout(n20079));
  jor  g19824(.dina(n10813), .dinb(n10134), .dout(n20080));
  jor  g19825(.dina(n9849), .dinb(n10051), .dout(n20081));
  jor  g19826(.dina(n10137), .dinb(n10523), .dout(n20082));
  jand g19827(.dina(n20082), .dinb(n20081), .dout(n20083));
  jand g19828(.dina(n20083), .dinb(n20080), .dout(n20084));
  jxor g19829(.dina(n20084), .dinb(a62 ), .dout(n20085));
  jxor g19830(.dina(n20085), .dinb(n20079), .dout(n20086));
  jxor g19831(.dina(n20086), .dinb(n20070), .dout(n20087));
  jnot g19832(.din(n20087), .dout(n20088));
  jxor g19833(.dina(n20088), .dinb(n20067), .dout(f124 ));
  jand g19834(.dina(n20086), .dinb(n20070), .dout(n20090));
  jnot g19835(.din(n20090), .dout(n20091));
  jor  g19836(.dina(n20088), .dinb(n20067), .dout(n20092));
  jand g19837(.dina(n20092), .dinb(n20091), .dout(n20093));
  jand g19838(.dina(n20077), .dinb(n20074), .dout(n20094));
  jnot g19839(.din(n20094), .dout(n20095));
  jor  g19840(.dina(n20085), .dinb(n20079), .dout(n20096));
  jand g19841(.dina(n20096), .dinb(n20095), .dout(n20097));
  jnot g19842(.din(n20097), .dout(n20098));
  jand g19843(.dina(n10594), .dinb(b61 ), .dout(n20099));
  jand g19844(.dina(n10129), .dinb(b62 ), .dout(n20100));
  jor  g19845(.dina(n20100), .dinb(n20099), .dout(n20101));
  jxor g19846(.dina(n20101), .dinb(n20074), .dout(n20102));
  jnot g19847(.din(n20102), .dout(n20103));
  jand g19848(.dina(n9850), .dinb(b63 ), .dout(n20104));
  jand g19849(.dina(n10832), .dinb(n9548), .dout(n20105));
  jor  g19850(.dina(n20105), .dinb(n20104), .dout(n20106));
  jxor g19851(.dina(n20106), .dinb(n9559), .dout(n20107));
  jxor g19852(.dina(n20107), .dinb(n20103), .dout(n20108));
  jxor g19853(.dina(n20108), .dinb(n20098), .dout(n20109));
  jnot g19854(.din(n20109), .dout(n20110));
  jxor g19855(.dina(n20110), .dinb(n20093), .dout(f125 ));
  jand g19856(.dina(n20108), .dinb(n20098), .dout(n20112));
  jnot g19857(.din(n20112), .dout(n20113));
  jor  g19858(.dina(n20110), .dinb(n20093), .dout(n20114));
  jand g19859(.dina(n20114), .dinb(n20113), .dout(n20115));
  jand g19860(.dina(n20101), .dinb(n20074), .dout(n20116));
  jnot g19861(.din(n20116), .dout(n20117));
  jor  g19862(.dina(n20107), .dinb(n20103), .dout(n20118));
  jand g19863(.dina(n20118), .dinb(n20117), .dout(n20119));
  jnot g19864(.din(a63 ), .dout(n20120));
  jor  g19865(.dina(b62 ), .dinb(n20120), .dout(n20121));
  jor  g19866(.dina(n20121), .dinb(n9559), .dout(n20122));
  jand g19867(.dina(a63 ), .dinb(n9559), .dout(n20123));
  jand g19868(.dina(n20123), .dinb(b63 ), .dout(n20124));
  jnot g19869(.din(n20124), .dout(n20125));
  jor  g19870(.dina(a63 ), .dinb(n9559), .dout(n20126));
  jor  g19871(.dina(n20126), .dinb(b63 ), .dout(n20127));
  jand g19872(.dina(n20127), .dinb(n20125), .dout(n20128));
  jand g19873(.dina(n20128), .dinb(n20122), .dout(n20129));
  jxor g19874(.dina(n20129), .dinb(n20073), .dout(n20130));
  jnot g19875(.din(n20130), .dout(n20131));
  jxor g19876(.dina(n20131), .dinb(n20119), .dout(n20132));
  jnot g19877(.din(n20132), .dout(n20133));
  jxor g19878(.dina(n20133), .dinb(n20115), .dout(f126 ));
  jor  g19879(.dina(n20131), .dinb(n20119), .dout(n20135));
  jor  g19880(.dina(n20133), .dinb(n20115), .dout(n20136));
  jand g19881(.dina(n20136), .dinb(n20135), .dout(n20137));
  jand g19882(.dina(n20129), .dinb(n20073), .dout(n20138));
  jor  g19883(.dina(n20138), .dinb(n20124), .dout(n20139));
  jand g19884(.dina(n10594), .dinb(b63 ), .dout(n20140));
  jxor g19885(.dina(n20140), .dinb(n20139), .dout(n20141));
  jxor g19886(.dina(n20141), .dinb(n20137), .dout(f127 ));
endmodule


