/*

c5315:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jdff: 6080
	jand: 606
	jor: 486

Summary:
	jxor: 112
	jspl: 279
	jspl3: 435
	jnot: 222
	jdff: 6080
	jand: 606
	jor: 486
*/

module c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [1:0] w_G1_2;
	wire [2:0] w_G4_0;
	wire [1:0] w_G11_0;
	wire [1:0] w_G14_0;
	wire [1:0] w_G17_0;
	wire [1:0] w_G20_0;
	wire [1:0] w_G37_0;
	wire [1:0] w_G40_0;
	wire [1:0] w_G43_0;
	wire [1:0] w_G46_0;
	wire [1:0] w_G49_0;
	wire [2:0] w_G54_0;
	wire [1:0] w_G61_0;
	wire [1:0] w_G64_0;
	wire [1:0] w_G67_0;
	wire [1:0] w_G70_0;
	wire [1:0] w_G73_0;
	wire [1:0] w_G76_0;
	wire [1:0] w_G91_0;
	wire [1:0] w_G100_0;
	wire [1:0] w_G103_0;
	wire [1:0] w_G106_0;
	wire [1:0] w_G109_0;
	wire [1:0] w_G123_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G137_2;
	wire [2:0] w_G137_3;
	wire [2:0] w_G137_4;
	wire [2:0] w_G137_5;
	wire [2:0] w_G137_6;
	wire [2:0] w_G137_7;
	wire [2:0] w_G137_8;
	wire [1:0] w_G137_9;
	wire [2:0] w_G141_0;
	wire [2:0] w_G141_1;
	wire [2:0] w_G141_2;
	wire [1:0] w_G146_0;
	wire [1:0] w_G149_0;
	wire [1:0] w_G152_0;
	wire [1:0] w_G155_0;
	wire [1:0] w_G158_0;
	wire [1:0] w_G161_0;
	wire [1:0] w_G164_0;
	wire [1:0] w_G167_0;
	wire [1:0] w_G170_0;
	wire [1:0] w_G173_0;
	wire [1:0] w_G182_0;
	wire [1:0] w_G185_0;
	wire [1:0] w_G188_0;
	wire [1:0] w_G191_0;
	wire [1:0] w_G194_0;
	wire [1:0] w_G197_0;
	wire [1:0] w_G200_0;
	wire [1:0] w_G203_0;
	wire [2:0] w_G206_0;
	wire [2:0] w_G206_1;
	wire [2:0] w_G210_0;
	wire [2:0] w_G210_1;
	wire [1:0] w_G210_2;
	wire [2:0] w_G218_0;
	wire [2:0] w_G218_1;
	wire [1:0] w_G218_2;
	wire [2:0] w_G226_0;
	wire [2:0] w_G226_1;
	wire [1:0] w_G226_2;
	wire [2:0] w_G234_0;
	wire [2:0] w_G234_1;
	wire [1:0] w_G234_2;
	wire [2:0] w_G242_0;
	wire [1:0] w_G242_1;
	wire [1:0] w_G245_0;
	wire [2:0] w_G248_0;
	wire [2:0] w_G248_1;
	wire [2:0] w_G248_2;
	wire [2:0] w_G248_3;
	wire [2:0] w_G248_4;
	wire [2:0] w_G248_5;
	wire [2:0] w_G251_0;
	wire [2:0] w_G251_1;
	wire [2:0] w_G251_2;
	wire [2:0] w_G251_3;
	wire [2:0] w_G251_4;
	wire [1:0] w_G251_5;
	wire [2:0] w_G254_0;
	wire [1:0] w_G254_1;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [1:0] w_G257_2;
	wire [2:0] w_G265_0;
	wire [2:0] w_G265_1;
	wire [2:0] w_G273_0;
	wire [2:0] w_G273_1;
	wire [1:0] w_G273_2;
	wire [2:0] w_G281_0;
	wire [2:0] w_G281_1;
	wire [1:0] w_G281_2;
	wire [1:0] w_G289_0;
	wire [2:0] w_G293_0;
	wire [2:0] w_G299_0;
	wire [2:0] w_G302_0;
	wire [2:0] w_G308_0;
	wire [2:0] w_G308_1;
	wire [2:0] w_G316_0;
	wire [1:0] w_G316_1;
	wire [2:0] w_G324_0;
	wire [2:0] w_G324_1;
	wire [1:0] w_G331_0;
	wire [2:0] w_G332_0;
	wire [2:0] w_G332_1;
	wire [2:0] w_G332_2;
	wire [2:0] w_G332_3;
	wire [2:0] w_G335_0;
	wire [1:0] w_G338_0;
	wire [2:0] w_G341_0;
	wire [2:0] w_G341_1;
	wire [2:0] w_G341_2;
	wire [1:0] w_G348_0;
	wire [2:0] w_G351_0;
	wire [2:0] w_G351_1;
	wire [2:0] w_G351_2;
	wire [1:0] w_G358_0;
	wire [2:0] w_G361_0;
	wire [1:0] w_G361_1;
	wire [1:0] w_G366_0;
	wire [1:0] w_G369_0;
	wire [2:0] w_G374_0;
	wire [2:0] w_G374_1;
	wire [2:0] w_G389_0;
	wire [2:0] w_G389_1;
	wire [2:0] w_G400_0;
	wire [2:0] w_G400_1;
	wire [2:0] w_G411_0;
	wire [2:0] w_G411_1;
	wire [1:0] w_G411_2;
	wire [2:0] w_G422_0;
	wire [1:0] w_G422_1;
	wire [2:0] w_G435_0;
	wire [2:0] w_G435_1;
	wire [2:0] w_G446_0;
	wire [2:0] w_G446_1;
	wire [2:0] w_G457_0;
	wire [2:0] w_G457_1;
	wire [2:0] w_G468_0;
	wire [2:0] w_G468_1;
	wire [2:0] w_G479_0;
	wire [2:0] w_G490_0;
	wire [1:0] w_G490_1;
	wire [2:0] w_G503_0;
	wire [2:0] w_G503_1;
	wire [1:0] w_G503_2;
	wire [2:0] w_G514_0;
	wire [2:0] w_G514_1;
	wire [1:0] w_G514_2;
	wire [2:0] w_G523_0;
	wire [2:0] w_G523_1;
	wire [2:0] w_G534_0;
	wire [2:0] w_G534_1;
	wire [1:0] w_G534_2;
	wire [2:0] w_G545_0;
	wire [2:0] w_G549_0;
	wire [1:0] w_G552_0;
	wire [1:0] w_G559_0;
	wire [1:0] w_G562_0;
	wire [2:0] w_G1497_0;
	wire [2:0] w_G1689_0;
	wire [2:0] w_G1689_1;
	wire [2:0] w_G1689_2;
	wire [2:0] w_G1689_3;
	wire [2:0] w_G1689_4;
	wire [1:0] w_G1689_5;
	wire [2:0] w_G1690_0;
	wire [1:0] w_G1690_1;
	wire [2:0] w_G1691_0;
	wire [2:0] w_G1691_1;
	wire [2:0] w_G1691_2;
	wire [2:0] w_G1691_3;
	wire [2:0] w_G1691_4;
	wire [1:0] w_G1691_5;
	wire [2:0] w_G1694_0;
	wire [1:0] w_G1694_1;
	wire [2:0] w_G2174_0;
	wire [2:0] w_G2358_0;
	wire [2:0] w_G2358_1;
	wire [2:0] w_G2358_2;
	wire [1:0] w_G3173_0;
	wire [2:0] w_G3546_0;
	wire [2:0] w_G3546_1;
	wire [2:0] w_G3546_2;
	wire [2:0] w_G3546_3;
	wire [2:0] w_G3546_4;
	wire [1:0] w_G3546_5;
	wire [2:0] w_G3548_0;
	wire [2:0] w_G3548_1;
	wire [2:0] w_G3548_2;
	wire [2:0] w_G3548_3;
	wire [2:0] w_G3548_4;
	wire [1:0] w_G3552_0;
	wire [1:0] w_G3717_0;
	wire [2:0] w_G3724_0;
	wire [2:0] w_G4087_0;
	wire [2:0] w_G4087_1;
	wire [2:0] w_G4087_2;
	wire [2:0] w_G4087_3;
	wire [2:0] w_G4087_4;
	wire [2:0] w_G4088_0;
	wire [2:0] w_G4088_1;
	wire [2:0] w_G4088_2;
	wire [2:0] w_G4088_3;
	wire [2:0] w_G4088_4;
	wire [2:0] w_G4088_5;
	wire [2:0] w_G4088_6;
	wire [2:0] w_G4088_7;
	wire [2:0] w_G4088_8;
	wire [2:0] w_G4088_9;
	wire [2:0] w_G4089_0;
	wire [2:0] w_G4089_1;
	wire [2:0] w_G4089_2;
	wire [2:0] w_G4089_3;
	wire [2:0] w_G4089_4;
	wire [2:0] w_G4089_5;
	wire [2:0] w_G4089_6;
	wire [2:0] w_G4089_7;
	wire [2:0] w_G4089_8;
	wire [2:0] w_G4089_9;
	wire [2:0] w_G4090_0;
	wire [2:0] w_G4090_1;
	wire [2:0] w_G4090_2;
	wire [2:0] w_G4090_3;
	wire [2:0] w_G4090_4;
	wire [2:0] w_G4091_0;
	wire [2:0] w_G4091_1;
	wire [2:0] w_G4091_2;
	wire [2:0] w_G4091_3;
	wire [2:0] w_G4091_4;
	wire [2:0] w_G4091_5;
	wire [1:0] w_G4091_6;
	wire [2:0] w_G4092_0;
	wire [2:0] w_G4092_1;
	wire [2:0] w_G4092_2;
	wire [2:0] w_G4092_3;
	wire [2:0] w_G4092_4;
	wire [2:0] w_G4092_5;
	wire [2:0] w_G4092_6;
	wire [2:0] w_G4092_7;
	wire [2:0] w_G4092_8;
	wire [2:0] w_G4092_9;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire [2:0] w_G809_0;
	wire [2:0] w_G809_1;
	wire [2:0] w_G809_2;
	wire [1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G623_0;
	wire G623_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G998_0;
	wire G998_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G865_0;
	wire G865_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire [1:0] w_n316_0;
	wire [1:0] w_n318_0;
	wire [2:0] w_n326_0;
	wire [2:0] w_n326_1;
	wire [1:0] w_n326_2;
	wire [1:0] w_n333_0;
	wire [1:0] w_n336_0;
	wire [1:0] w_n361_0;
	wire [1:0] w_n365_0;
	wire [2:0] w_n366_0;
	wire [2:0] w_n366_1;
	wire [2:0] w_n369_0;
	wire [2:0] w_n369_1;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [2:0] w_n374_0;
	wire [1:0] w_n374_1;
	wire [2:0] w_n375_0;
	wire [2:0] w_n375_1;
	wire [2:0] w_n375_2;
	wire [2:0] w_n375_3;
	wire [2:0] w_n375_4;
	wire [2:0] w_n377_0;
	wire [1:0] w_n377_1;
	wire [2:0] w_n378_0;
	wire [2:0] w_n378_1;
	wire [2:0] w_n378_2;
	wire [2:0] w_n378_3;
	wire [2:0] w_n378_4;
	wire [1:0] w_n386_0;
	wire [2:0] w_n387_0;
	wire [1:0] w_n387_1;
	wire [2:0] w_n389_0;
	wire [1:0] w_n389_1;
	wire [1:0] w_n397_0;
	wire [1:0] w_n401_0;
	wire [2:0] w_n402_0;
	wire [2:0] w_n406_0;
	wire [2:0] w_n406_1;
	wire [2:0] w_n406_2;
	wire [2:0] w_n406_3;
	wire [2:0] w_n406_4;
	wire [1:0] w_n406_5;
	wire [2:0] w_n408_0;
	wire [2:0] w_n408_1;
	wire [2:0] w_n408_2;
	wire [2:0] w_n408_3;
	wire [2:0] w_n408_4;
	wire [2:0] w_n408_5;
	wire [2:0] w_n412_0;
	wire [1:0] w_n414_0;
	wire [1:0] w_n415_0;
	wire [2:0] w_n423_0;
	wire [2:0] w_n425_0;
	wire [2:0] w_n428_0;
	wire [1:0] w_n428_1;
	wire [1:0] w_n429_0;
	wire [2:0] w_n433_0;
	wire [2:0] w_n435_0;
	wire [2:0] w_n435_1;
	wire [1:0] w_n435_2;
	wire [1:0] w_n437_0;
	wire [1:0] w_n445_0;
	wire [2:0] w_n449_0;
	wire [2:0] w_n449_1;
	wire [2:0] w_n451_0;
	wire [1:0] w_n459_0;
	wire [2:0] w_n460_0;
	wire [2:0] w_n460_1;
	wire [2:0] w_n462_0;
	wire [1:0] w_n470_0;
	wire [2:0] w_n471_0;
	wire [2:0] w_n471_1;
	wire [2:0] w_n473_0;
	wire [1:0] w_n473_1;
	wire [1:0] w_n481_0;
	wire [2:0] w_n483_0;
	wire [2:0] w_n483_1;
	wire [1:0] w_n483_2;
	wire [2:0] w_n485_0;
	wire [1:0] w_n485_1;
	wire [1:0] w_n493_0;
	wire [2:0] w_n494_0;
	wire [2:0] w_n494_1;
	wire [2:0] w_n496_0;
	wire [1:0] w_n496_1;
	wire [1:0] w_n504_0;
	wire [2:0] w_n507_0;
	wire [2:0] w_n507_1;
	wire [2:0] w_n509_0;
	wire [1:0] w_n517_0;
	wire [2:0] w_n518_0;
	wire [2:0] w_n518_1;
	wire [2:0] w_n520_0;
	wire [1:0] w_n528_0;
	wire [2:0] w_n530_0;
	wire [2:0] w_n530_1;
	wire [2:0] w_n532_0;
	wire [1:0] w_n532_1;
	wire [1:0] w_n540_0;
	wire [1:0] w_n543_0;
	wire [2:0] w_n551_0;
	wire [2:0] w_n556_0;
	wire [2:0] w_n556_1;
	wire [2:0] w_n556_2;
	wire [2:0] w_n556_3;
	wire [2:0] w_n556_4;
	wire [2:0] w_n556_5;
	wire [2:0] w_n556_6;
	wire [2:0] w_n556_7;
	wire [1:0] w_n556_8;
	wire [1:0] w_n557_0;
	wire [1:0] w_n559_0;
	wire [2:0] w_n560_0;
	wire [2:0] w_n561_0;
	wire [1:0] w_n561_1;
	wire [1:0] w_n562_0;
	wire [1:0] w_n564_0;
	wire [2:0] w_n565_0;
	wire [2:0] w_n566_0;
	wire [2:0] w_n567_0;
	wire [1:0] w_n569_0;
	wire [1:0] w_n571_0;
	wire [2:0] w_n572_0;
	wire [2:0] w_n573_0;
	wire [2:0] w_n574_0;
	wire [2:0] w_n578_0;
	wire [1:0] w_n578_1;
	wire [2:0] w_n579_0;
	wire [1:0] w_n579_1;
	wire [1:0] w_n581_0;
	wire [2:0] w_n586_0;
	wire [1:0] w_n586_1;
	wire [1:0] w_n587_0;
	wire [2:0] w_n588_0;
	wire [1:0] w_n588_1;
	wire [2:0] w_n591_0;
	wire [1:0] w_n591_1;
	wire [2:0] w_n592_0;
	wire [2:0] w_n596_0;
	wire [1:0] w_n596_1;
	wire [2:0] w_n597_0;
	wire [2:0] w_n601_0;
	wire [1:0] w_n601_1;
	wire [2:0] w_n602_0;
	wire [1:0] w_n603_0;
	wire [2:0] w_n607_0;
	wire [1:0] w_n607_1;
	wire [2:0] w_n608_0;
	wire [2:0] w_n609_0;
	wire [2:0] w_n611_0;
	wire [2:0] w_n613_0;
	wire [2:0] w_n613_1;
	wire [2:0] w_n613_2;
	wire [2:0] w_n613_3;
	wire [2:0] w_n613_4;
	wire [2:0] w_n613_5;
	wire [2:0] w_n617_0;
	wire [1:0] w_n617_1;
	wire [2:0] w_n618_0;
	wire [2:0] w_n619_0;
	wire [2:0] w_n619_1;
	wire [2:0] w_n620_0;
	wire [1:0] w_n620_1;
	wire [1:0] w_n621_0;
	wire [1:0] w_n623_0;
	wire [2:0] w_n624_0;
	wire [1:0] w_n625_0;
	wire [2:0] w_n627_0;
	wire [1:0] w_n627_1;
	wire [2:0] w_n628_0;
	wire [1:0] w_n631_0;
	wire [1:0] w_n632_0;
	wire [2:0] w_n635_0;
	wire [1:0] w_n635_1;
	wire [2:0] w_n636_0;
	wire [2:0] w_n637_0;
	wire [1:0] w_n638_0;
	wire [2:0] w_n639_0;
	wire [1:0] w_n640_0;
	wire [2:0] w_n641_0;
	wire [2:0] w_n641_1;
	wire [2:0] w_n644_0;
	wire [2:0] w_n648_0;
	wire [1:0] w_n648_1;
	wire [1:0] w_n649_0;
	wire [1:0] w_n650_0;
	wire [2:0] w_n653_0;
	wire [2:0] w_n654_0;
	wire [2:0] w_n654_1;
	wire [2:0] w_n654_2;
	wire [2:0] w_n658_0;
	wire [1:0] w_n658_1;
	wire [1:0] w_n659_0;
	wire [2:0] w_n660_0;
	wire [1:0] w_n660_1;
	wire [1:0] w_n661_0;
	wire [1:0] w_n670_0;
	wire [1:0] w_n680_0;
	wire [2:0] w_n682_0;
	wire [1:0] w_n684_0;
	wire [1:0] w_n685_0;
	wire [1:0] w_n686_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n689_0;
	wire [1:0] w_n690_0;
	wire [1:0] w_n692_0;
	wire [2:0] w_n694_0;
	wire [2:0] w_n695_0;
	wire [2:0] w_n699_0;
	wire [1:0] w_n701_0;
	wire [2:0] w_n703_0;
	wire [1:0] w_n704_0;
	wire [1:0] w_n709_0;
	wire [1:0] w_n710_0;
	wire [1:0] w_n711_0;
	wire [2:0] w_n713_0;
	wire [2:0] w_n715_0;
	wire [1:0] w_n717_0;
	wire [1:0] w_n719_0;
	wire [1:0] w_n720_0;
	wire [1:0] w_n721_0;
	wire [1:0] w_n722_0;
	wire [2:0] w_n725_0;
	wire [1:0] w_n726_0;
	wire [1:0] w_n728_0;
	wire [2:0] w_n733_0;
	wire [2:0] w_n735_0;
	wire [2:0] w_n737_0;
	wire [1:0] w_n737_1;
	wire [1:0] w_n738_0;
	wire [2:0] w_n742_0;
	wire [1:0] w_n745_0;
	wire [2:0] w_n746_0;
	wire [1:0] w_n747_0;
	wire [2:0] w_n749_0;
	wire [2:0] w_n749_1;
	wire [2:0] w_n749_2;
	wire [2:0] w_n749_3;
	wire [2:0] w_n749_4;
	wire [2:0] w_n749_5;
	wire [2:0] w_n749_6;
	wire [2:0] w_n749_7;
	wire [2:0] w_n749_8;
	wire [2:0] w_n749_9;
	wire [2:0] w_n749_10;
	wire [2:0] w_n749_11;
	wire [2:0] w_n749_12;
	wire [1:0] w_n749_13;
	wire [2:0] w_n750_0;
	wire [2:0] w_n750_1;
	wire [2:0] w_n750_2;
	wire [2:0] w_n750_3;
	wire [2:0] w_n750_4;
	wire [2:0] w_n750_5;
	wire [2:0] w_n750_6;
	wire [2:0] w_n750_7;
	wire [2:0] w_n750_8;
	wire [2:0] w_n753_0;
	wire [1:0] w_n753_1;
	wire [1:0] w_n755_0;
	wire [2:0] w_n763_0;
	wire [1:0] w_n767_0;
	wire [1:0] w_n779_0;
	wire [2:0] w_n786_0;
	wire [2:0] w_n788_0;
	wire [2:0] w_n790_0;
	wire [2:0] w_n792_0;
	wire [2:0] w_n795_0;
	wire [1:0] w_n795_1;
	wire [2:0] w_n797_0;
	wire [2:0] w_n797_1;
	wire [2:0] w_n797_2;
	wire [2:0] w_n797_3;
	wire [2:0] w_n797_4;
	wire [2:0] w_n797_5;
	wire [2:0] w_n797_6;
	wire [2:0] w_n797_7;
	wire [2:0] w_n797_8;
	wire [1:0] w_n797_9;
	wire [2:0] w_n798_0;
	wire [1:0] w_n798_1;
	wire [2:0] w_n800_0;
	wire [2:0] w_n800_1;
	wire [2:0] w_n800_2;
	wire [2:0] w_n800_3;
	wire [1:0] w_n800_4;
	wire [2:0] w_n801_0;
	wire [1:0] w_n801_1;
	wire [2:0] w_n814_0;
	wire [2:0] w_n819_0;
	wire [1:0] w_n821_0;
	wire [1:0] w_n824_0;
	wire [1:0] w_n827_0;
	wire [1:0] w_n836_0;
	wire [1:0] w_n847_0;
	wire [2:0] w_n852_0;
	wire [2:0] w_n852_1;
	wire [2:0] w_n852_2;
	wire [2:0] w_n852_3;
	wire [2:0] w_n852_4;
	wire [2:0] w_n852_5;
	wire [2:0] w_n852_6;
	wire [2:0] w_n852_7;
	wire [2:0] w_n852_8;
	wire [1:0] w_n852_9;
	wire [2:0] w_n854_0;
	wire [2:0] w_n854_1;
	wire [2:0] w_n854_2;
	wire [2:0] w_n854_3;
	wire [1:0] w_n854_4;
	wire [2:0] w_n865_0;
	wire [1:0] w_n867_0;
	wire [1:0] w_n868_0;
	wire [1:0] w_n870_0;
	wire [1:0] w_n871_0;
	wire [1:0] w_n880_0;
	wire [1:0] w_n890_0;
	wire [1:0] w_n901_0;
	wire [2:0] w_n923_0;
	wire [1:0] w_n935_0;
	wire [2:0] w_n938_0;
	wire [2:0] w_n940_0;
	wire [1:0] w_n940_1;
	wire [1:0] w_n944_0;
	wire [1:0] w_n949_0;
	wire [1:0] w_n953_0;
	wire [2:0] w_n954_0;
	wire [1:0] w_n957_0;
	wire [1:0] w_n962_0;
	wire [1:0] w_n964_0;
	wire [1:0] w_n969_0;
	wire [2:0] w_n977_0;
	wire [1:0] w_n981_0;
	wire [1:0] w_n986_0;
	wire [1:0] w_n989_0;
	wire [2:0] w_n993_0;
	wire [2:0] w_n993_1;
	wire [2:0] w_n993_2;
	wire [2:0] w_n993_3;
	wire [2:0] w_n993_4;
	wire [2:0] w_n994_0;
	wire [2:0] w_n994_1;
	wire [2:0] w_n994_2;
	wire [2:0] w_n994_3;
	wire [1:0] w_n994_4;
	wire [2:0] w_n996_0;
	wire [2:0] w_n996_1;
	wire [2:0] w_n996_2;
	wire [2:0] w_n996_3;
	wire [1:0] w_n996_4;
	wire [2:0] w_n999_0;
	wire [2:0] w_n999_1;
	wire [2:0] w_n999_2;
	wire [2:0] w_n999_3;
	wire [2:0] w_n1007_0;
	wire [2:0] w_n1007_1;
	wire [2:0] w_n1007_2;
	wire [2:0] w_n1007_3;
	wire [2:0] w_n1008_0;
	wire [2:0] w_n1008_1;
	wire [2:0] w_n1008_2;
	wire [2:0] w_n1008_3;
	wire [2:0] w_n1008_4;
	wire [2:0] w_n1012_0;
	wire [2:0] w_n1012_1;
	wire [2:0] w_n1012_2;
	wire [2:0] w_n1012_3;
	wire [1:0] w_n1012_4;
	wire [2:0] w_n1014_0;
	wire [2:0] w_n1014_1;
	wire [2:0] w_n1014_2;
	wire [2:0] w_n1014_3;
	wire [1:0] w_n1014_4;
	wire [2:0] w_n1019_0;
	wire [1:0] w_n1019_1;
	wire [2:0] w_n1021_0;
	wire [1:0] w_n1021_1;
	wire [2:0] w_n1030_0;
	wire [1:0] w_n1030_1;
	wire [2:0] w_n1032_0;
	wire [1:0] w_n1032_1;
	wire [2:0] w_n1041_0;
	wire [1:0] w_n1041_1;
	wire [2:0] w_n1043_0;
	wire [1:0] w_n1043_1;
	wire [2:0] w_n1052_0;
	wire [1:0] w_n1052_1;
	wire [2:0] w_n1054_0;
	wire [1:0] w_n1054_1;
	wire [1:0] w_n1177_0;
	wire [1:0] w_n1179_0;
	wire [2:0] w_n1196_0;
	wire [2:0] w_n1196_1;
	wire [2:0] w_n1201_0;
	wire [2:0] w_n1205_0;
	wire [2:0] w_n1205_1;
	wire [2:0] w_n1213_0;
	wire [2:0] w_n1213_1;
	wire [2:0] w_n1236_0;
	wire [2:0] w_n1236_1;
	wire [2:0] w_n1251_0;
	wire [2:0] w_n1251_1;
	wire [2:0] w_n1279_0;
	wire [1:0] w_n1279_1;
	wire [2:0] w_n1297_0;
	wire [1:0] w_n1297_1;
	wire [2:0] w_n1299_0;
	wire [1:0] w_n1299_1;
	wire [2:0] w_n1410_0;
	wire [2:0] w_n1412_0;
	wire [1:0] w_n1416_0;
	wire [1:0] w_n1422_0;
	wire [1:0] w_n1425_0;
	wire [1:0] w_n1428_0;
	wire [1:0] w_n1429_0;
	wire [1:0] w_n1451_0;
	wire [1:0] w_n1503_0;
	wire [1:0] w_n1504_0;
	wire [1:0] w_n1592_0;
	wire [1:0] w_n1593_0;
	wire [1:0] w_n1596_0;
	wire [1:0] w_n1599_0;
	wire [1:0] w_n1603_0;
	wire [1:0] w_n1605_0;
	wire [1:0] w_n1609_0;
	wire [2:0] w_n1611_0;
	wire [1:0] w_n1613_0;
	wire [1:0] w_n1615_0;
	wire [1:0] w_n1618_0;
	wire [1:0] w_n1633_0;
	wire [1:0] w_n1637_0;
	wire [1:0] w_n1643_0;
	wire [1:0] w_n1652_0;
	wire [1:0] w_n1665_0;
	wire [2:0] w_n1674_0;
	wire [1:0] w_n1675_0;
	wire [2:0] w_n1679_0;
	wire [1:0] w_n1680_0;
	wire [1:0] w_n1694_0;
	wire [1:0] w_n1695_0;
	wire [1:0] w_n1698_0;
	wire w_dff_B_zheJpM8a6_1;
	wire w_dff_B_AHgrt4gg1_0;
	wire w_dff_B_qYdKW0mJ1_1;
	wire w_dff_B_fb4w6OY08_1;
	wire w_dff_B_C8HPys6d9_2;
	wire w_dff_B_bn2KitwD0_1;
	wire w_dff_B_y0l8qKDv5_1;
	wire w_dff_B_rt3JmqTJ3_0;
	wire w_dff_B_yhLpS0385_1;
	wire w_dff_B_6QeaS1DH6_1;
	wire w_dff_B_mF2s9CBA5_0;
	wire w_dff_B_B3mKvrRi2_1;
	wire w_dff_A_r314CZIx0_0;
	wire w_dff_A_aWAYliXz7_0;
	wire w_dff_A_nO7XEJJZ0_0;
	wire w_dff_A_qdReZtOb3_0;
	wire w_dff_A_EQDWtB3Z5_1;
	wire w_dff_A_7SteU1572_1;
	wire w_dff_A_kGSLAakd1_1;
	wire w_dff_A_ISYTkH6Z2_1;
	wire w_dff_B_p6DqrFtN8_1;
	wire w_dff_B_F9C7J14E4_0;
	wire w_dff_B_R8DwcryY0_1;
	wire w_dff_B_NunCSItv5_1;
	wire w_dff_B_uJshMeGM7_1;
	wire w_dff_B_ujKs66H17_1;
	wire w_dff_A_Zx3hLzlE1_0;
	wire w_dff_A_5ZzhKa771_1;
	wire w_dff_A_418twjYf5_1;
	wire w_dff_A_gfj8NwyJ8_1;
	wire w_dff_A_EOYooCHi1_1;
	wire w_dff_A_97f50Gyd7_1;
	wire w_dff_A_YBfL4dKa4_2;
	wire w_dff_A_xkvQGNFG3_2;
	wire w_dff_A_vPHTtLPc4_2;
	wire w_dff_A_2t5NEtJb8_2;
	wire w_dff_B_oCKraORR2_1;
	wire w_dff_B_Aw4rgnp34_2;
	wire w_dff_B_WK3ML1VB5_2;
	wire w_dff_B_8622ALns4_2;
	wire w_dff_B_TlLd4l4R7_2;
	wire w_dff_B_mZyTBMf28_1;
	wire w_dff_B_Kt9ZlpMB8_1;
	wire w_dff_B_OFXwU7gD7_1;
	wire w_dff_B_RWLZ8jjJ7_1;
	wire w_dff_B_yrzte8g70_1;
	wire w_dff_B_zkPt8ae05_1;
	wire w_dff_B_GxGmzWvC4_1;
	wire w_dff_B_rxiWQAuY8_1;
	wire w_dff_B_QjFUmAcP5_1;
	wire w_dff_B_Vbora1Dg2_1;
	wire w_dff_B_8ZvMHrhM6_1;
	wire w_dff_A_MQXPV9BM5_1;
	wire w_dff_A_0MJbWzah7_1;
	wire w_dff_B_Vj7upYsK3_3;
	wire w_dff_B_BnjGn0yx4_2;
	wire w_dff_B_aNbiEs9k0_2;
	wire w_dff_B_1AgEg32t4_1;
	wire w_dff_B_UHgRrhal6_1;
	wire w_dff_A_BXfDRO4x4_0;
	wire w_dff_A_EHvls1S40_0;
	wire w_dff_A_lsaOxW2a0_0;
	wire w_dff_A_tWrpcTYi4_0;
	wire w_dff_A_BGwoNCKI6_0;
	wire w_dff_B_BKFKSKfn1_0;
	wire w_dff_B_cEkFTT688_0;
	wire w_dff_B_3TRYXpeV8_0;
	wire w_dff_B_kemvdtiQ3_0;
	wire w_dff_B_747LGKLP3_0;
	wire w_dff_B_OJj8kJAy1_0;
	wire w_dff_B_SjbGrnKe5_0;
	wire w_dff_B_Rgr8YSoU1_0;
	wire w_dff_B_olpJCSgP0_0;
	wire w_dff_B_RxKT6oOM6_0;
	wire w_dff_B_mrdx43LZ1_0;
	wire w_dff_A_hSru95eO1_1;
	wire w_dff_A_1Qrvskhk6_1;
	wire w_dff_A_lvNXFgN21_1;
	wire w_dff_A_BoKIMQyz7_1;
	wire w_dff_A_CF9HRJSa3_1;
	wire w_dff_A_rFDWPpvm6_1;
	wire w_dff_A_4fRtJ2Ld0_1;
	wire w_dff_A_VHKzP71n5_1;
	wire w_dff_A_hpnhSO6P5_1;
	wire w_dff_A_mEwAEQZs7_1;
	wire w_dff_B_zCBNTJbm1_0;
	wire w_dff_B_q0lgKwgL4_0;
	wire w_dff_B_tOxloe6R5_0;
	wire w_dff_B_KePzRO2j6_0;
	wire w_dff_B_6ejKKBRn3_0;
	wire w_dff_B_Ub1LOGCF4_0;
	wire w_dff_B_87aM68wY3_0;
	wire w_dff_B_oXpZxqun1_0;
	wire w_dff_B_k1ScRTkN0_0;
	wire w_dff_B_qqeTdjm71_0;
	wire w_dff_B_SC9aAKpH0_2;
	wire w_dff_B_fDqSVZGS8_0;
	wire w_dff_A_PSHJIkKu0_1;
	wire w_dff_A_xwnBkUym2_1;
	wire w_dff_A_llIZNsjG6_1;
	wire w_dff_A_N6HFh5Os7_1;
	wire w_dff_A_6qTt9jls3_1;
	wire w_dff_A_vTdWxZHE0_1;
	wire w_dff_A_ANUWJxK22_1;
	wire w_dff_A_NOjQBMsE7_1;
	wire w_dff_A_L6tmT5B07_1;
	wire w_dff_A_CnFrIYZc7_1;
	wire w_dff_B_mvtfbOKG2_0;
	wire w_dff_B_t6uc02AZ3_1;
	wire w_dff_B_E6nqMAx73_1;
	wire w_dff_B_F93TvI0b1_1;
	wire w_dff_B_ma5VyXQF8_0;
	wire w_dff_B_mseprEIa2_1;
	wire w_dff_B_aCYRy2Ew9_1;
	wire w_dff_B_tGoH7vJM5_1;
	wire w_dff_B_iCfsAdeF9_1;
	wire w_dff_B_vBhC3C0o8_1;
	wire w_dff_B_a9G33OtV7_1;
	wire w_dff_B_WvPKT57L9_1;
	wire w_dff_B_vy8eF0Ht1_1;
	wire w_dff_B_T9BagvzE4_1;
	wire w_dff_B_LWJuJS1r0_1;
	wire w_dff_B_OdbN9Vw01_1;
	wire w_dff_B_WEmpJA6T0_1;
	wire w_dff_B_ryhRjljt1_1;
	wire w_dff_B_gDqMrgC01_1;
	wire w_dff_B_8bHPYGMg2_1;
	wire w_dff_B_o6Ii1tFw3_1;
	wire w_dff_B_uZMLw7vn2_1;
	wire w_dff_B_F3veK4cD5_1;
	wire w_dff_B_PfKdQwpT6_1;
	wire w_dff_B_GP8W2Ox08_1;
	wire w_dff_B_uTGJv7LH8_1;
	wire w_dff_B_aNc5nfHR2_1;
	wire w_dff_B_a84F3n2V2_1;
	wire w_dff_B_CpMuQuO23_1;
	wire w_dff_B_a4g8dfkr9_1;
	wire w_dff_B_gD1qHAC90_1;
	wire w_dff_B_ScYqek9Z6_1;
	wire w_dff_B_gTsL1HLz8_1;
	wire w_dff_B_k6SjvXSa7_1;
	wire w_dff_B_pD7lTEdd0_0;
	wire w_dff_B_62L0GS0U4_0;
	wire w_dff_B_WldPV59z8_0;
	wire w_dff_B_pPDT1AQ16_0;
	wire w_dff_B_23bCwgkB6_0;
	wire w_dff_B_kfFsUcZl7_0;
	wire w_dff_B_5dojtcMA0_0;
	wire w_dff_B_ZaDQDCL62_0;
	wire w_dff_B_qIMYH9Qa7_0;
	wire w_dff_B_BSGKBOSb8_0;
	wire w_dff_B_2MIFHDv32_0;
	wire w_dff_B_f2GERJv18_1;
	wire w_dff_B_hqcGs7799_2;
	wire w_dff_B_1nqnb48u7_2;
	wire w_dff_B_FgmiDBhq7_2;
	wire w_dff_B_f4CK2JYY4_1;
	wire w_dff_B_XW9QjEk24_1;
	wire w_dff_B_VRgdXbNk2_1;
	wire w_dff_B_fBgsIMRS9_1;
	wire w_dff_B_CmOPjsED1_1;
	wire w_dff_B_8oO7MKjx3_1;
	wire w_dff_B_FJmefle53_1;
	wire w_dff_B_wWBhILXJ6_1;
	wire w_dff_B_0z2OHNJy6_0;
	wire w_dff_B_G5AviPzR2_1;
	wire w_dff_B_W6Ge03QS3_1;
	wire w_dff_A_pOxdtWsD6_0;
	wire w_dff_A_2mTScvy55_0;
	wire w_dff_B_Rm3ZK2Nx8_1;
	wire w_dff_B_4atA8eYM2_1;
	wire w_dff_B_PdZaLB6I9_1;
	wire w_dff_B_z6H0G1qN4_1;
	wire w_dff_B_MpnMFYaW1_1;
	wire w_dff_A_HyeU5No36_0;
	wire w_dff_A_OK5Px8QS4_0;
	wire w_dff_A_udCIlLJj0_0;
	wire w_dff_A_Nz7dAw6z6_0;
	wire w_dff_A_5MXuvVuT3_0;
	wire w_dff_A_k0Wk6R5K6_0;
	wire w_dff_A_uij7RR0U6_0;
	wire w_dff_A_zcM0sTcP0_0;
	wire w_dff_A_b00oFZC20_0;
	wire w_dff_A_wOYSOi314_0;
	wire w_dff_A_3vp1aYyX1_0;
	wire w_dff_B_v8h3GWND4_1;
	wire w_dff_B_fRNMjkG23_1;
	wire w_dff_B_7hi2OYhc7_0;
	wire w_dff_B_8CL04iFQ3_0;
	wire w_dff_B_s4wS4LRY2_0;
	wire w_dff_B_dn3hLhNJ1_0;
	wire w_dff_B_q7blMNJ18_0;
	wire w_dff_B_SblSu6v96_0;
	wire w_dff_B_OOjWpZ8N2_0;
	wire w_dff_B_e4us51jA8_0;
	wire w_dff_B_bF6LpzLO7_0;
	wire w_dff_B_0AVJ2yW95_0;
	wire w_dff_B_xzv5ohvN7_0;
	wire w_dff_B_WMSvK1lZ5_0;
	wire w_dff_B_c0siQ1Xo7_0;
	wire w_dff_B_zpsoaStt8_0;
	wire w_dff_B_wT1TZ09k6_0;
	wire w_dff_B_5gqfWVpb8_0;
	wire w_dff_B_neTZGdA48_1;
	wire w_dff_A_GnEUwN5J3_0;
	wire w_dff_A_WrQhqWRE5_0;
	wire w_dff_A_b8VkJsUx7_0;
	wire w_dff_A_5Zmgp9vf8_0;
	wire w_dff_A_dc2Ayljc6_0;
	wire w_dff_A_PlB2W2G97_0;
	wire w_dff_A_HaikhZZP3_0;
	wire w_dff_B_AB2s4cjT6_0;
	wire w_dff_B_4V624dSC0_0;
	wire w_dff_B_vSHwxjNt3_0;
	wire w_dff_B_FrnA06350_0;
	wire w_dff_B_gWo9ypdf2_0;
	wire w_dff_B_J5YxlibS3_0;
	wire w_dff_B_0U00ivlP3_0;
	wire w_dff_B_ytJmcFom0_0;
	wire w_dff_B_kNflGQzO7_0;
	wire w_dff_B_i46h3C6x0_0;
	wire w_dff_B_yCbYYlZM4_0;
	wire w_dff_B_YYFfSKoS8_0;
	wire w_dff_B_cJNGMVyF6_0;
	wire w_dff_B_aRCPDiZZ3_0;
	wire w_dff_B_lUb34adj1_0;
	wire w_dff_B_AiJxHKK30_1;
	wire w_dff_B_Cgqz8Wrk5_1;
	wire w_dff_A_7bUtwmem0_0;
	wire w_dff_A_jRn4hofL0_0;
	wire w_dff_A_VHpr4vki4_0;
	wire w_dff_A_lnf7rF5H4_0;
	wire w_dff_A_y6y09Jhf9_0;
	wire w_dff_A_alptRk5K0_0;
	wire w_dff_A_GXnVcBu23_0;
	wire w_dff_A_JaYRlBjm4_0;
	wire w_dff_A_ZbGSDWDX6_0;
	wire w_dff_A_ePEtkknh1_0;
	wire w_dff_A_MrNfuHpO4_0;
	wire w_dff_A_ni5jUwik3_0;
	wire w_dff_A_jc1ziRt50_0;
	wire w_dff_A_RHImzFgB8_0;
	wire w_dff_A_vhDY77Uo2_0;
	wire w_dff_A_uC3BmT1G3_2;
	wire w_dff_A_FRG6RNVF9_2;
	wire w_dff_A_CJZTRi2D7_2;
	wire w_dff_A_CN6zjNi78_2;
	wire w_dff_A_V9B0xiSf7_2;
	wire w_dff_A_ANwwNvdi7_2;
	wire w_dff_A_ymGeKsyE7_2;
	wire w_dff_A_HAG0qOwE3_2;
	wire w_dff_A_zXr0jjtr2_2;
	wire w_dff_A_Q3qG3HaV8_2;
	wire w_dff_A_xoeEYkuv6_2;
	wire w_dff_A_vUVoVSqV0_2;
	wire w_dff_A_zYbC1g8u3_2;
	wire w_dff_A_aeomzd4N3_2;
	wire w_dff_A_v3sdImXK4_2;
	wire w_dff_A_DjpfCeFM4_2;
	wire w_dff_A_5jc5QGIQ2_0;
	wire w_dff_A_sc1dwBSy1_0;
	wire w_dff_A_zk37MMkW3_0;
	wire w_dff_A_LaLxD0iW4_0;
	wire w_dff_A_EVGMUc7m3_0;
	wire w_dff_A_9n5u9eqE3_0;
	wire w_dff_A_kyf6Pxnx1_0;
	wire w_dff_A_4f8H9TnG9_0;
	wire w_dff_A_ip7iEMmh2_0;
	wire w_dff_A_eV7pVUD00_0;
	wire w_dff_A_3o7htMax4_0;
	wire w_dff_A_XVBPQJOj8_0;
	wire w_dff_A_2nbBza6c2_0;
	wire w_dff_A_If5rry6V3_2;
	wire w_dff_A_Fg0SGsut4_2;
	wire w_dff_A_uCwmK0434_2;
	wire w_dff_A_gJwoiWJP8_2;
	wire w_dff_A_iEW0y4j53_2;
	wire w_dff_A_eXTSK3Q03_2;
	wire w_dff_A_7LDOQc7k1_2;
	wire w_dff_A_S8yWeT8N2_2;
	wire w_dff_A_1CcmG2343_2;
	wire w_dff_A_oncGayq52_2;
	wire w_dff_A_ZYEJExNN1_2;
	wire w_dff_A_7JOIGxhs2_2;
	wire w_dff_A_JYf4Vl1q7_2;
	wire w_dff_A_JzxeJp815_2;
	wire w_dff_A_IzK3vsdV9_2;
	wire w_dff_B_6Bdj4B4U4_0;
	wire w_dff_B_O4dZeWzu8_0;
	wire w_dff_B_XdLfVSZa3_0;
	wire w_dff_B_AGuYI6W31_0;
	wire w_dff_B_JRyez78m4_0;
	wire w_dff_B_YWsugIs99_0;
	wire w_dff_B_LeXiBPKp7_0;
	wire w_dff_B_sWUguajH4_0;
	wire w_dff_B_1WYIyQsI4_0;
	wire w_dff_B_jfIJiS205_0;
	wire w_dff_B_54iNMhB09_0;
	wire w_dff_B_KABlnsFX8_0;
	wire w_dff_B_vv8Jq0650_0;
	wire w_dff_B_1CWlwn4L5_1;
	wire w_dff_A_61z1j6fq9_1;
	wire w_dff_A_j6YpSyXi4_1;
	wire w_dff_A_cRjUyetP3_1;
	wire w_dff_A_1W3Ck1436_1;
	wire w_dff_A_qx2BPPnp8_1;
	wire w_dff_A_cjUmcXkp1_1;
	wire w_dff_A_UhE6Z2CL7_1;
	wire w_dff_A_BX5AsIJI4_1;
	wire w_dff_A_viNjIyen4_1;
	wire w_dff_A_7DejEo559_1;
	wire w_dff_A_jxrR6EKm0_1;
	wire w_dff_A_EdaKIGxL6_1;
	wire w_dff_A_tjxL3j0M0_1;
	wire w_dff_A_2dQI5PSU5_1;
	wire w_dff_A_pn99vB4U9_1;
	wire w_dff_A_fPSn3NTK8_1;
	wire w_dff_A_hDK65s6C0_1;
	wire w_dff_A_w5738VEI4_1;
	wire w_dff_A_iucM0O0N7_1;
	wire w_dff_A_yTmAVrjS3_1;
	wire w_dff_A_Ct4zHAir9_1;
	wire w_dff_A_Pjsmd1b37_1;
	wire w_dff_A_2Q8jkmHO1_1;
	wire w_dff_A_wSVjyqq36_1;
	wire w_dff_A_NO74DbYq5_1;
	wire w_dff_B_3RD362Ma7_0;
	wire w_dff_B_ABqfpzg69_0;
	wire w_dff_B_UXtPxzaz2_0;
	wire w_dff_B_mcjsLtE48_0;
	wire w_dff_B_LeYyvyyl1_0;
	wire w_dff_B_yHPxfBZP8_0;
	wire w_dff_B_v9F355C89_0;
	wire w_dff_B_cA8qxjrA3_0;
	wire w_dff_B_1EiByaox8_0;
	wire w_dff_B_UpPZtJjT7_0;
	wire w_dff_B_vMRXBdSu0_0;
	wire w_dff_B_6y5qsEFA3_0;
	wire w_dff_B_Yz3a1iCD0_0;
	wire w_dff_B_lGrJQWgO6_0;
	wire w_dff_B_gGOmb6Bm4_1;
	wire w_dff_B_9mRNvP8I7_1;
	wire w_dff_B_CFdtmdKf5_1;
	wire w_dff_A_dHQr3Ovf9_0;
	wire w_dff_A_1zfdfJ0M9_2;
	wire w_dff_A_1ZfHs2xD5_2;
	wire w_dff_B_eH5w5cXP7_1;
	wire w_dff_B_kXMGvePy1_1;
	wire w_dff_B_fo2TNkQC5_1;
	wire w_dff_B_gKidYRAM0_1;
	wire w_dff_B_MJJtl3TZ6_1;
	wire w_dff_B_PGQTR6aG6_1;
	wire w_dff_B_8hMl1rn83_1;
	wire w_dff_B_oCnKrViL6_1;
	wire w_dff_B_U0pF2d0Q4_1;
	wire w_dff_B_sAkCvf2i1_1;
	wire w_dff_B_Xuc4zKOq6_1;
	wire w_dff_B_RgypynPF0_1;
	wire w_dff_B_kRcWTs473_1;
	wire w_dff_B_mbZ9vNCi8_1;
	wire w_dff_B_R05Mb3Zj5_1;
	wire w_dff_A_iDEZo0bi8_0;
	wire w_dff_A_GUJ3mcq12_0;
	wire w_dff_A_oDOfYQRV4_0;
	wire w_dff_A_2PV4RARu0_0;
	wire w_dff_A_AWzuBgCD8_0;
	wire w_dff_A_Uv1SmpKj6_0;
	wire w_dff_A_AerqLyH93_0;
	wire w_dff_A_F5luKNX98_0;
	wire w_dff_B_GERK1vqb5_1;
	wire w_dff_B_B0CHzlMz8_1;
	wire w_dff_B_dDPN7lR71_2;
	wire w_dff_B_v2rBuvSz1_1;
	wire w_dff_B_lKxiErD48_1;
	wire w_dff_B_gtujfV0o4_1;
	wire w_dff_B_0EuHrGhe6_1;
	wire w_dff_B_FLtnVVxT3_1;
	wire w_dff_B_BMfdatlS3_1;
	wire w_dff_B_SYDRlI0o9_1;
	wire w_dff_B_CAlsrD1v5_1;
	wire w_dff_B_YiHDiKMQ2_1;
	wire w_dff_B_cWIjwMMG6_1;
	wire w_dff_B_CEHtdWAg3_1;
	wire w_dff_B_bukuZ7MZ2_1;
	wire w_dff_B_O435alBe3_1;
	wire w_dff_B_LimWu8Tx3_1;
	wire w_dff_B_Lb1UTJyr6_0;
	wire w_dff_B_h7vnw1GH2_1;
	wire w_dff_B_0rjRKGPo7_1;
	wire w_dff_A_N9HelVsD7_1;
	wire w_dff_A_pxtHcMGG8_1;
	wire w_dff_A_XG7yHMMk8_1;
	wire w_dff_A_OV93YCTK4_1;
	wire w_dff_A_iLu1TPBr6_1;
	wire w_dff_A_Uv5qASFg5_1;
	wire w_dff_A_Wz3AUKzj7_1;
	wire w_dff_A_1q8jEL7r5_1;
	wire w_dff_A_Ia0vxgIO5_1;
	wire w_dff_A_bykttAQo3_1;
	wire w_dff_A_n88C7xSF6_1;
	wire w_dff_A_KrLRbemN7_1;
	wire w_dff_A_uhEqaxQP3_1;
	wire w_dff_A_n7XmxIk65_1;
	wire w_dff_A_hSbRJQCb8_1;
	wire w_dff_B_c1qR84vA7_2;
	wire w_dff_A_xjhFeVW48_1;
	wire w_dff_A_9xX7rbI98_1;
	wire w_dff_A_Grx4iNpn6_1;
	wire w_dff_A_eDRVwpQg3_1;
	wire w_dff_A_AaLsFLOJ9_1;
	wire w_dff_A_L2JRw27O9_1;
	wire w_dff_A_6if27TvK9_1;
	wire w_dff_A_GTRcu69w7_1;
	wire w_dff_A_DSNQ5J132_1;
	wire w_dff_A_6QIJxjfZ3_1;
	wire w_dff_A_xkF9HX0C0_1;
	wire w_dff_A_4NcFoFno2_1;
	wire w_dff_A_JOSlMOXr1_1;
	wire w_dff_A_HznXxpI56_1;
	wire w_dff_A_80tlyiIj1_1;
	wire w_dff_A_2ssKatZa8_1;
	wire w_dff_B_VQnQKQRU0_1;
	wire w_dff_B_aigW7DO80_1;
	wire w_dff_B_rONFTPY69_1;
	wire w_dff_B_evSSdnCp8_1;
	wire w_dff_B_N9oHBLAw4_1;
	wire w_dff_B_8S2wpDdz9_1;
	wire w_dff_B_CzwBVkD16_1;
	wire w_dff_B_o6snahXM1_1;
	wire w_dff_B_w5Qd7Bf83_1;
	wire w_dff_B_gpGkC0je6_1;
	wire w_dff_B_9aJWE6Au3_1;
	wire w_dff_B_4iclhfl35_1;
	wire w_dff_B_VStuxuLR3_1;
	wire w_dff_B_KOtNylFL9_1;
	wire w_dff_A_0b42GaHs4_0;
	wire w_dff_A_HasVrbxU8_0;
	wire w_dff_A_coAWXkyc8_0;
	wire w_dff_A_fBLIayiT8_0;
	wire w_dff_A_qvAmdHs83_0;
	wire w_dff_A_gqhERKaS8_0;
	wire w_dff_A_Qicp42AP9_0;
	wire w_dff_A_ginIMhxv5_0;
	wire w_dff_A_eexujbIh5_0;
	wire w_dff_A_KGVFU3zd0_0;
	wire w_dff_A_p4xrh6Df5_0;
	wire w_dff_A_8iaWdJjL1_0;
	wire w_dff_A_Ok4ajb1u1_2;
	wire w_dff_A_yRYfx1bf7_2;
	wire w_dff_A_lc7V1lKu0_2;
	wire w_dff_A_cbFSyLib9_2;
	wire w_dff_A_JmqDn6vc0_2;
	wire w_dff_A_Iy704UMF1_2;
	wire w_dff_A_yp9BvMpr8_2;
	wire w_dff_A_j6B03wjY9_2;
	wire w_dff_A_5QnVrgew1_2;
	wire w_dff_A_CcIk7B5N7_2;
	wire w_dff_A_ZIM4o9Ut8_2;
	wire w_dff_A_jbxI6xua1_2;
	wire w_dff_A_wEMJAAj20_2;
	wire w_dff_B_54uO2SaK2_2;
	wire w_dff_A_UZk809mu4_0;
	wire w_dff_A_VW7VbnnE2_0;
	wire w_dff_A_HYaYbMfj2_0;
	wire w_dff_A_89gHHQnH9_0;
	wire w_dff_A_NIac5FuB1_0;
	wire w_dff_A_g2GujtPk1_0;
	wire w_dff_A_PDkhJbq54_0;
	wire w_dff_A_hXanfFp21_0;
	wire w_dff_A_B4F0XnhH6_0;
	wire w_dff_A_C9wvEsN02_0;
	wire w_dff_A_1V4NTzXZ9_0;
	wire w_dff_A_c14cnpsO7_0;
	wire w_dff_A_oas7hLWv3_0;
	wire w_dff_A_nFqbBqfq5_2;
	wire w_dff_A_kdyrguMd8_2;
	wire w_dff_A_pgRJUIvr9_2;
	wire w_dff_A_WveXqnPt2_2;
	wire w_dff_A_d3hGncqQ2_2;
	wire w_dff_A_spm6nWV19_2;
	wire w_dff_A_BuoTJ5PJ1_2;
	wire w_dff_A_3SSokXxc4_2;
	wire w_dff_A_u8fD9G8y0_2;
	wire w_dff_A_mHf5WpV89_2;
	wire w_dff_A_OyoOkfum3_2;
	wire w_dff_A_vMo8Fad50_2;
	wire w_dff_A_rwJY1WPL1_2;
	wire w_dff_A_9KJNIPPm5_2;
	wire w_dff_A_caZmU7uz2_2;
	wire w_dff_B_gudhFVs46_0;
	wire w_dff_B_DqGdbygq5_0;
	wire w_dff_B_IvNO6U535_0;
	wire w_dff_B_b0fUwg5J6_0;
	wire w_dff_B_R84XIJoo9_0;
	wire w_dff_B_cUYTpxcm3_0;
	wire w_dff_B_oYPcxJV91_0;
	wire w_dff_B_txNPpcLf6_0;
	wire w_dff_B_Tgv9zwm00_0;
	wire w_dff_B_fn5qG8Ad1_0;
	wire w_dff_B_GFwzuDQT0_0;
	wire w_dff_B_MEU79m7I0_0;
	wire w_dff_B_7shZPb5S7_0;
	wire w_dff_B_vohdLkQS8_0;
	wire w_dff_A_3CliLQJe9_1;
	wire w_dff_A_sJEdiHEr5_2;
	wire w_dff_B_c7zUEjUl7_2;
	wire w_dff_B_Ydtt0Oin9_1;
	wire w_dff_B_X2YHWpL72_1;
	wire w_dff_B_w7zKmeRY0_1;
	wire w_dff_A_1o31NhMe6_2;
	wire w_dff_A_TfsvbHxf8_2;
	wire w_dff_B_vzT0zQNM9_0;
	wire w_dff_B_97mNUZED7_0;
	wire w_dff_B_NJ7VpaXy6_0;
	wire w_dff_B_X0LG8B3j2_0;
	wire w_dff_B_OY2u0qCL7_0;
	wire w_dff_B_XD2yctU06_0;
	wire w_dff_B_iY4Mz0ZL5_0;
	wire w_dff_B_0DFwfqhO9_0;
	wire w_dff_B_ZycPv5oO8_0;
	wire w_dff_B_rvyPFMQt5_0;
	wire w_dff_B_C8aP4go06_0;
	wire w_dff_B_VclQYvSf9_0;
	wire w_dff_B_UN6jiYz77_0;
	wire w_dff_B_kAtZXHiP9_0;
	wire w_dff_B_whG8IqYl2_0;
	wire w_dff_B_uHtD4vlp5_0;
	wire w_dff_B_YTrvBkwS9_1;
	wire w_dff_B_kIMNewnG9_0;
	wire w_dff_B_8hYkhCJR0_0;
	wire w_dff_B_nu4abJga0_0;
	wire w_dff_B_PJtGooSC0_0;
	wire w_dff_B_SgEkj2yl8_0;
	wire w_dff_B_Cs7V7OsT2_0;
	wire w_dff_B_c6oeIReX9_0;
	wire w_dff_B_BHwnXhEW7_0;
	wire w_dff_B_p2bxcDom7_0;
	wire w_dff_B_7Hydlfbz9_0;
	wire w_dff_B_MO8fuRYc6_0;
	wire w_dff_B_EiX5KooM5_0;
	wire w_dff_B_01lO3jCx5_0;
	wire w_dff_B_jKbWAgBq6_0;
	wire w_dff_A_8rINv8s73_0;
	wire w_dff_A_WMGHNPP52_0;
	wire w_dff_A_eJjTXKVm4_0;
	wire w_dff_A_38Agb6mp8_1;
	wire w_dff_A_xs2o5xqt0_1;
	wire w_dff_A_Pxi0wDm27_1;
	wire w_dff_A_8fIelWnw4_1;
	wire w_dff_A_62QZ4HDJ8_1;
	wire w_dff_A_JwLeYHrO6_1;
	wire w_dff_A_se7hXFni1_1;
	wire w_dff_A_tBVgznO13_0;
	wire w_dff_A_mkuxMxtW7_0;
	wire w_dff_A_3309tWKO4_0;
	wire w_dff_A_BAG2IICU2_0;
	wire w_dff_A_RaJD5xjh5_0;
	wire w_dff_A_PiOZqbeA7_1;
	wire w_dff_A_3FxU5nc13_1;
	wire w_dff_A_jMOXm3su3_1;
	wire w_dff_A_3pCUS7so0_1;
	wire w_dff_A_NOqqj6Mk0_1;
	wire w_dff_A_KmrKza565_1;
	wire w_dff_A_6BM9BGGk0_1;
	wire w_dff_B_hEqM9Hw33_0;
	wire w_dff_B_82pZnk8y6_0;
	wire w_dff_B_SzKpfUr24_0;
	wire w_dff_B_wsVCZe921_0;
	wire w_dff_B_l7FQPIQ24_0;
	wire w_dff_B_LRl3Xlgv4_0;
	wire w_dff_B_fonvdCnR0_0;
	wire w_dff_B_tXsp4Gnj1_0;
	wire w_dff_B_pn6eVVIs8_0;
	wire w_dff_B_TddAKzks3_0;
	wire w_dff_B_f2zBYRdW6_0;
	wire w_dff_B_yzIneDGH8_0;
	wire w_dff_B_zLZyw14N6_0;
	wire w_dff_B_HPK9lmlb8_1;
	wire w_dff_A_WB0fIQGN5_2;
	wire w_dff_A_KIUPQkRY8_2;
	wire w_dff_A_tbNmrbzc5_2;
	wire w_dff_B_IrZilIV99_0;
	wire w_dff_B_BHVBc84c2_0;
	wire w_dff_B_jXuyVCod4_0;
	wire w_dff_B_V7LK8I483_0;
	wire w_dff_B_YJWGexCA6_0;
	wire w_dff_B_uWr62opr2_0;
	wire w_dff_B_kuzGrrfn5_0;
	wire w_dff_B_hBm8z6RF3_0;
	wire w_dff_B_GHnnGyVa1_0;
	wire w_dff_B_P6iuIBXH4_0;
	wire w_dff_B_wzegfj990_0;
	wire w_dff_B_YUOZX00c4_0;
	wire w_dff_B_ytrX5FtM3_0;
	wire w_dff_B_1gDrkq6x2_0;
	wire w_dff_A_8lDlWQtO6_0;
	wire w_dff_A_VwRZDwaz7_0;
	wire w_dff_A_CC2qWIf52_1;
	wire w_dff_B_EqsrlkAY9_1;
	wire w_dff_B_jHZRUrdB5_1;
	wire w_dff_B_aBQHPIZc5_1;
	wire w_dff_B_GGtYoyhv6_1;
	wire w_dff_B_TQGPFfCw7_1;
	wire w_dff_B_v8xPUZ0R9_1;
	wire w_dff_B_TAsVhcUW7_1;
	wire w_dff_B_ZZS7ScBr7_1;
	wire w_dff_B_MBEZ6rRW8_1;
	wire w_dff_B_N0in5UnQ0_1;
	wire w_dff_B_fYRue3RB7_1;
	wire w_dff_B_ucU94RGc6_1;
	wire w_dff_B_VzIQXCFb0_1;
	wire w_dff_B_1KsPs9Jb0_1;
	wire w_dff_B_BlvpqnAG2_1;
	wire w_dff_B_7oZaUpvj9_1;
	wire w_dff_B_l8beA7pM1_1;
	wire w_dff_B_07b8zMqv5_1;
	wire w_dff_B_UtSEGdzN4_1;
	wire w_dff_B_0WME3dXU5_1;
	wire w_dff_B_Chuzd4SF0_1;
	wire w_dff_B_x9F0mnhp2_1;
	wire w_dff_B_5DvTuiwh8_1;
	wire w_dff_B_q6572KBE3_1;
	wire w_dff_B_jvNVoFVk8_1;
	wire w_dff_B_rT3rqSo23_1;
	wire w_dff_B_FPhCeDhE9_1;
	wire w_dff_B_D5DDbU3o9_1;
	wire w_dff_B_ROLApdNa1_1;
	wire w_dff_B_WKTjbkHm1_1;
	wire w_dff_B_nrtzlCTv5_1;
	wire w_dff_B_GmlogMg49_1;
	wire w_dff_B_06DKGFZm7_1;
	wire w_dff_B_Zah5riXS9_1;
	wire w_dff_B_A8p3AAgU4_1;
	wire w_dff_B_2UMaT1uP5_1;
	wire w_dff_B_2E2F5T8i2_1;
	wire w_dff_B_CC2gThHC7_1;
	wire w_dff_B_zk9vWeIP4_1;
	wire w_dff_B_fEbiifXh7_1;
	wire w_dff_B_PLgQJAgZ1_1;
	wire w_dff_B_AlFxG4ep9_1;
	wire w_dff_B_PVCJ2hWw0_1;
	wire w_dff_B_4eTKlpJq8_1;
	wire w_dff_B_W7L2ew7r4_0;
	wire w_dff_B_zBDlRoN46_0;
	wire w_dff_B_089RRlJP9_0;
	wire w_dff_B_JCYl6Vhl2_0;
	wire w_dff_B_BSCnZAbv7_0;
	wire w_dff_B_UIS0n0cy6_0;
	wire w_dff_B_w0Q4eRMQ9_1;
	wire w_dff_B_f9YYUJeb7_1;
	wire w_dff_B_Gez3os9P9_1;
	wire w_dff_B_O6iMNlxl3_1;
	wire w_dff_B_i9fWGNyT8_1;
	wire w_dff_B_X2fQecv99_1;
	wire w_dff_B_xAtnCFNh5_1;
	wire w_dff_B_CQYza13j0_1;
	wire w_dff_B_E1lXjz2A0_1;
	wire w_dff_B_YFG3Hif90_1;
	wire w_dff_B_0QZLWL4B4_1;
	wire w_dff_B_SOpIKrXM3_1;
	wire w_dff_B_qJMxlCiJ1_1;
	wire w_dff_B_unc3xdOr2_1;
	wire w_dff_B_WYWrfO6q3_1;
	wire w_dff_B_dLBtxQ8b9_1;
	wire w_dff_B_Mg9x6ze98_1;
	wire w_dff_B_5VSO5p555_1;
	wire w_dff_B_bhV7aBCh0_1;
	wire w_dff_B_xHA3HxgH1_0;
	wire w_dff_B_rfXfVhsf2_0;
	wire w_dff_B_YAiDbcMe4_0;
	wire w_dff_B_IQzoHech8_0;
	wire w_dff_B_OzL3IZBd2_0;
	wire w_dff_B_WLwaQdrP9_0;
	wire w_dff_B_7ogaCzHa8_1;
	wire w_dff_B_E4vL1V1K6_1;
	wire w_dff_B_wrJwdZHd9_1;
	wire w_dff_B_G7WvKJ7j7_1;
	wire w_dff_B_fV1F7oBh6_2;
	wire w_dff_B_3Dl9XxUb6_2;
	wire w_dff_B_Zm4pvZX48_2;
	wire w_dff_B_nbNfm5IV3_0;
	wire w_dff_B_0leJRDAP4_0;
	wire w_dff_B_VeiRMqA10_0;
	wire w_dff_B_GAdN59NS5_0;
	wire w_dff_B_D40llUlT4_0;
	wire w_dff_B_QejdSoeG8_0;
	wire w_dff_B_5Dl9fguZ6_0;
	wire w_dff_B_0CnjIi0W3_0;
	wire w_dff_B_WV9Yg7W70_0;
	wire w_dff_B_lv6Mg72Q9_0;
	wire w_dff_B_7fhbX3HY4_0;
	wire w_dff_B_J0McyiMk6_0;
	wire w_dff_B_y1UOWzRD6_0;
	wire w_dff_B_UGVHS3ko5_2;
	wire w_dff_B_lu2Jmb9Z9_2;
	wire w_dff_B_HOpJCSUc9_2;
	wire w_dff_B_pivs3WiK7_0;
	wire w_dff_B_u74rHInI8_1;
	wire w_dff_B_axjqmemQ7_1;
	wire w_dff_B_15dOJZD46_1;
	wire w_dff_B_d1IJW1IA7_1;
	wire w_dff_B_QFF1pcNc9_1;
	wire w_dff_B_Nwaz4MU14_1;
	wire w_dff_B_gsZrcHqF9_0;
	wire w_dff_B_i3OubGyD6_0;
	wire w_dff_B_24dM6nyX0_1;
	wire w_dff_B_GSMPQl2M4_1;
	wire w_dff_A_L34K2jlO5_0;
	wire w_dff_A_a2QCXQJn3_0;
	wire w_dff_B_0JWCdQHO9_1;
	wire w_dff_B_23LC9GOZ8_1;
	wire w_dff_B_IX2dHluj9_1;
	wire w_dff_A_L20R3OvP1_0;
	wire w_dff_A_kKypQXJj3_1;
	wire w_dff_A_eaZBJOnx8_1;
	wire w_dff_A_mbsEs87r4_1;
	wire w_dff_A_KOawNj8j2_1;
	wire w_dff_A_MiXGg6Hi7_1;
	wire w_dff_A_3SCYQOmj0_1;
	wire w_dff_B_pcbEym5T3_1;
	wire w_dff_B_LmUy60EZ2_1;
	wire w_dff_B_Tqqg0m4r6_1;
	wire w_dff_B_iOoWjQo79_1;
	wire w_dff_B_jhURF59J7_1;
	wire w_dff_B_OxIp23Sa1_1;
	wire w_dff_B_5iz5ATwb1_1;
	wire w_dff_B_4w5sM2TQ6_1;
	wire w_dff_B_J0DbFJi31_0;
	wire w_dff_B_vxSfaeuF8_0;
	wire w_dff_B_pv4rlYUd0_0;
	wire w_dff_B_QreqmqU37_0;
	wire w_dff_B_QIFB1MSw6_1;
	wire w_dff_B_SyeDNte46_1;
	wire w_dff_B_26RCtZf59_0;
	wire w_dff_B_V8ceVBG67_0;
	wire w_dff_B_Zajdvmtw0_0;
	wire w_dff_B_fqdV4id69_0;
	wire w_dff_A_cdVVsjCe9_0;
	wire w_dff_A_tIMtKK4g7_0;
	wire w_dff_A_k97jq2Wn5_0;
	wire w_dff_A_wja9FsvO5_0;
	wire w_dff_A_l8pysX0x7_0;
	wire w_dff_A_FuIfPWWe8_0;
	wire w_dff_A_WU9mHmMW4_0;
	wire w_dff_A_fxBZz2dK4_0;
	wire w_dff_A_qfAREajh4_0;
	wire w_dff_A_wJpX3Al28_0;
	wire w_dff_A_h5HoD7D52_2;
	wire w_dff_A_Lg6FT8AN9_2;
	wire w_dff_A_2NvsHdUV5_2;
	wire w_dff_B_Bo2dviGY1_1;
	wire w_dff_B_BIz860tW5_1;
	wire w_dff_A_sDoJ2deg5_1;
	wire w_dff_A_UctEwY1H7_1;
	wire w_dff_A_Kc8Z5IzR5_1;
	wire w_dff_A_XY0BUQfE6_1;
	wire w_dff_A_jG2qodlf0_2;
	wire w_dff_A_BPIqf5rI7_0;
	wire w_dff_A_QWfpafDM6_0;
	wire w_dff_A_bR76bPca5_1;
	wire w_dff_A_ue7qSbSQ9_1;
	wire w_dff_B_VCTn3SK60_0;
	wire w_dff_B_dm1VS66N0_0;
	wire w_dff_B_JCpG3cxf4_0;
	wire w_dff_B_Xir8SzCa5_0;
	wire w_dff_B_gENNqRjE4_0;
	wire w_dff_B_jM36jj2Z9_0;
	wire w_dff_B_nADyp6BT6_0;
	wire w_dff_B_3io3D0Hr7_0;
	wire w_dff_B_7rEfuANi1_0;
	wire w_dff_B_O1rvdU333_0;
	wire w_dff_B_hMrZ0uPE2_0;
	wire w_dff_B_uQSx3YNL7_0;
	wire w_dff_B_MkJiLRTw9_0;
	wire w_dff_B_FBUy87R54_2;
	wire w_dff_B_8QufpCzT9_2;
	wire w_dff_B_4ob1Ejiw3_2;
	wire w_dff_B_7TNR61dt0_1;
	wire w_dff_B_ynkkfbZU5_1;
	wire w_dff_B_Wi5oBCgA5_1;
	wire w_dff_B_WHUSTBAt3_1;
	wire w_dff_B_alWXNTHX7_1;
	wire w_dff_B_a6ZFEYDl6_1;
	wire w_dff_B_W9MvtiD98_1;
	wire w_dff_B_0ObkkvA53_1;
	wire w_dff_B_xf4nFuBp8_0;
	wire w_dff_B_D28aOgyg8_0;
	wire w_dff_B_Uja55WdY4_0;
	wire w_dff_B_WhjvR4bw5_1;
	wire w_dff_B_RgaHLtTI8_1;
	wire w_dff_B_N46Q13tX9_1;
	wire w_dff_B_TVfQ4Pp23_1;
	wire w_dff_B_d0O73iLt7_1;
	wire w_dff_B_PRLkGbq50_1;
	wire w_dff_B_d1hn19lt3_1;
	wire w_dff_B_tTJAqodU4_1;
	wire w_dff_B_euE0zI9h3_1;
	wire w_dff_B_HJcQ4XXB1_1;
	wire w_dff_B_tkO5Zrls7_1;
	wire w_dff_B_0m77Vsxo6_1;
	wire w_dff_B_j0sHRqff0_1;
	wire w_dff_B_bdLFoM7E2_1;
	wire w_dff_B_g0gNCxJa4_1;
	wire w_dff_A_KIDJxiBf7_0;
	wire w_dff_A_3cKzkmaC5_0;
	wire w_dff_A_Sdx6V3Sz3_0;
	wire w_dff_A_D0Gyjluq5_0;
	wire w_dff_A_SJ5wKky19_0;
	wire w_dff_B_a2IDp3261_1;
	wire w_dff_B_U9XiRrDq4_1;
	wire w_dff_B_s5MMWwXL4_1;
	wire w_dff_B_YHnInmKb8_1;
	wire w_dff_B_iO59QYdP1_0;
	wire w_dff_B_UI3T1w9Q6_0;
	wire w_dff_B_IyXndkve0_0;
	wire w_dff_B_lbZteEbc9_0;
	wire w_dff_B_LKoMlFcM0_0;
	wire w_dff_B_MALlDwj99_0;
	wire w_dff_B_wjbyFsUv4_0;
	wire w_dff_B_H1JCgz9B3_0;
	wire w_dff_B_rJO1WmZA8_0;
	wire w_dff_B_qeF7S8Vs7_0;
	wire w_dff_B_ILLp9iLJ9_0;
	wire w_dff_B_Hr3vt8wg1_0;
	wire w_dff_B_OTqproJZ7_0;
	wire w_dff_B_sFIvMDpm4_0;
	wire w_dff_B_C5Gn2Iqp1_2;
	wire w_dff_B_8LJWb9wq6_2;
	wire w_dff_B_4NUXgw828_2;
	wire w_dff_B_lpCaWUUQ1_1;
	wire w_dff_B_GOhy5pRA2_1;
	wire w_dff_B_rsoI9LAR9_1;
	wire w_dff_B_pnfwq5m68_1;
	wire w_dff_B_tvhdN1lp1_1;
	wire w_dff_B_DjSPTOBr9_1;
	wire w_dff_B_0h2uZ0XB6_1;
	wire w_dff_B_nuJyNRVB7_1;
	wire w_dff_B_uUyw6SBA8_0;
	wire w_dff_B_0i0gv2C88_0;
	wire w_dff_B_3Fv80fzf9_0;
	wire w_dff_B_V3cGInGs1_0;
	wire w_dff_B_zOGq44EE9_1;
	wire w_dff_B_XsWxfEym6_1;
	wire w_dff_A_eP7Rd7X16_2;
	wire w_dff_A_VfKayZhp7_2;
	wire w_dff_A_HTohEeBT0_2;
	wire w_dff_A_F0JhapCz1_0;
	wire w_dff_A_uKOnJYMr6_0;
	wire w_dff_A_hJYd0ebg5_0;
	wire w_dff_A_ALOmsiws4_0;
	wire w_dff_A_cxXdvzs87_0;
	wire w_dff_A_IkAbCPM81_1;
	wire w_dff_A_iToMPgUv9_2;
	wire w_dff_A_wM42BPhe6_2;
	wire w_dff_B_wNUOId764_1;
	wire w_dff_B_ztXtA0sx5_1;
	wire w_dff_A_MwqBT1ch8_0;
	wire w_dff_A_TFA1s4mL4_0;
	wire w_dff_A_2hbXSAaW4_1;
	wire w_dff_B_ef1jqy0p4_1;
	wire w_dff_B_eUK8pFhK0_1;
	wire w_dff_B_cpJWD3be5_1;
	wire w_dff_B_nHlm3X4o6_1;
	wire w_dff_B_o6Hv4IOT0_1;
	wire w_dff_B_upyi4HYX0_1;
	wire w_dff_B_2GZjt7VG3_1;
	wire w_dff_B_gaJd1ReL8_1;
	wire w_dff_B_Kz64QH1X3_1;
	wire w_dff_B_91QUffPM9_0;
	wire w_dff_B_yTyBLB759_0;
	wire w_dff_B_cbCql3jt1_0;
	wire w_dff_B_b3x1WAc13_0;
	wire w_dff_B_vl6j40Uh3_0;
	wire w_dff_B_ztQca1h34_0;
	wire w_dff_B_ub1rWXPF9_1;
	wire w_dff_A_09RYPLEY5_0;
	wire w_dff_A_NVDs0d1O7_1;
	wire w_dff_A_UPMtDmzk0_0;
	wire w_dff_A_NexaASTY3_2;
	wire w_dff_A_AnjC0Ijo8_1;
	wire w_dff_A_SwxSWY5E6_2;
	wire w_dff_A_XuWp6dEZ8_0;
	wire w_dff_A_K6H9YeB14_0;
	wire w_dff_A_I3fQUKHa0_0;
	wire w_dff_A_IqMxCBZb8_0;
	wire w_dff_A_PNbiSLXZ2_0;
	wire w_dff_A_GQD2edxX0_0;
	wire w_dff_A_XA3HZLVg6_0;
	wire w_dff_A_SuK89Nxe8_1;
	wire w_dff_A_DaXJgAHl0_1;
	wire w_dff_A_LTAqX0I66_2;
	wire w_dff_A_HiMulCm28_2;
	wire w_dff_A_QgVLGpdo9_2;
	wire w_dff_A_oF8Rkg9O6_2;
	wire w_dff_A_v65CWJYg0_2;
	wire w_dff_B_p4Mf3qHF5_3;
	wire w_dff_B_eHIEZXIz1_3;
	wire w_dff_A_64uspizJ6_0;
	wire w_dff_A_e4xWmsaF2_0;
	wire w_dff_A_HcMG7EVG3_0;
	wire w_dff_A_NGs4s4Vo9_0;
	wire w_dff_A_8F6JTJkA8_2;
	wire w_dff_A_VFM07rhN7_2;
	wire w_dff_A_jFYyJij92_2;
	wire w_dff_B_FQ5DCCzZ8_1;
	wire w_dff_B_JVMS83W53_1;
	wire w_dff_B_878hfwhA2_1;
	wire w_dff_B_dlQcxcXw5_1;
	wire w_dff_B_ggkqwLvQ9_1;
	wire w_dff_B_BuYMsqKl6_1;
	wire w_dff_B_xX9dfFky5_1;
	wire w_dff_B_a8L4tgbd2_1;
	wire w_dff_B_Q2chBNhn7_1;
	wire w_dff_B_HcL4UfEc1_1;
	wire w_dff_B_90w1LJGs7_1;
	wire w_dff_B_rtwK8WQK2_1;
	wire w_dff_B_Cp5HUqhv1_1;
	wire w_dff_B_awR0QHK92_1;
	wire w_dff_B_NukNxX8y4_1;
	wire w_dff_B_O7Wf56j41_1;
	wire w_dff_B_yFj93FxD3_1;
	wire w_dff_B_X4t6qNE25_1;
	wire w_dff_B_MBTv1AYc8_1;
	wire w_dff_B_QSIfbudR1_1;
	wire w_dff_B_IvTs3Xyw0_1;
	wire w_dff_B_aUrDXous6_1;
	wire w_dff_B_h2Z1q8qw5_1;
	wire w_dff_B_l2bDNCRO1_1;
	wire w_dff_B_74DlTyWW2_1;
	wire w_dff_B_GwvYsTUa7_1;
	wire w_dff_B_PmqqNJOO4_1;
	wire w_dff_B_pJUAKFgW4_1;
	wire w_dff_B_iXjaPqPW3_1;
	wire w_dff_B_JEENBjMl8_1;
	wire w_dff_B_okZtuIBU5_0;
	wire w_dff_B_34JMfYHQ5_0;
	wire w_dff_B_r0ShhH3K0_0;
	wire w_dff_B_00tyfqLR7_0;
	wire w_dff_B_1QfqCUSw9_0;
	wire w_dff_B_0ULmIPpw8_0;
	wire w_dff_B_6A3aoKRn7_0;
	wire w_dff_B_nxRAlrok4_0;
	wire w_dff_B_plC7k5TJ0_0;
	wire w_dff_B_eLQDXY4u6_0;
	wire w_dff_B_dTppWHvb1_0;
	wire w_dff_B_5qe7dsnQ1_0;
	wire w_dff_B_zflnnlws8_0;
	wire w_dff_B_I71IC8ty2_0;
	wire w_dff_B_2D6IMdj80_0;
	wire w_dff_B_VYAmWsj55_0;
	wire w_dff_B_JnpBMWfr7_1;
	wire w_dff_B_Kh4VdNXQ4_1;
	wire w_dff_B_GPiIhynG4_1;
	wire w_dff_B_TllRHp4q3_1;
	wire w_dff_B_sUH7TDOi9_1;
	wire w_dff_B_uaRH0Okv8_1;
	wire w_dff_B_mFXIpEUa0_1;
	wire w_dff_B_mx8dEiB92_1;
	wire w_dff_B_NEaFt02s3_1;
	wire w_dff_A_5zUNvNBm9_0;
	wire w_dff_A_mRIEnLgl0_0;
	wire w_dff_A_U72sNUkJ6_0;
	wire w_dff_A_8BHfggQZ0_0;
	wire w_dff_A_Fo2Mv4J16_0;
	wire w_dff_A_fcTc6bFA7_0;
	wire w_dff_A_2egfg4Gc8_0;
	wire w_dff_A_Twjnsnti9_0;
	wire w_dff_A_swfVtjcd7_0;
	wire w_dff_A_oT4WLw3O6_0;
	wire w_dff_A_ICC9pbgr6_0;
	wire w_dff_B_Q6fkFxpj8_2;
	wire w_dff_B_8LUOjPoT0_2;
	wire w_dff_B_aEjRTtTd9_2;
	wire w_dff_B_ZpVN6DKC2_2;
	wire w_dff_B_cYBHEi6R0_2;
	wire w_dff_A_5ks2fcuz9_0;
	wire w_dff_A_5EHyocmY4_1;
	wire w_dff_A_kfchUDvm4_2;
	wire w_dff_A_2Q8Xhje30_2;
	wire w_dff_A_ZCsVAV2w1_2;
	wire w_dff_A_dOM0HN591_2;
	wire w_dff_A_n00IHA5k6_0;
	wire w_dff_A_49KHGlqX7_0;
	wire w_dff_A_7TSw0oRm8_0;
	wire w_dff_A_nFLcoEgD4_0;
	wire w_dff_A_kMujjOwz8_0;
	wire w_dff_A_XV3EmB432_0;
	wire w_dff_A_xpomOwAB9_0;
	wire w_dff_A_Ac50fvil1_0;
	wire w_dff_A_1Lp7pGEt9_0;
	wire w_dff_A_zOiOBzm24_0;
	wire w_dff_A_vXobmQJ75_0;
	wire w_dff_B_cD0jNOOq0_1;
	wire w_dff_B_bwUTDkPc2_1;
	wire w_dff_B_uu0kXH8T2_1;
	wire w_dff_B_sGovDXq85_1;
	wire w_dff_B_MvEi3CGB6_1;
	wire w_dff_B_103t0hcc7_0;
	wire w_dff_B_Kz98kc4B3_0;
	wire w_dff_B_YG7YJKWX4_0;
	wire w_dff_B_7QKpzjzx6_0;
	wire w_dff_B_Mbqsu6jf8_0;
	wire w_dff_A_Ujmf1NMl0_0;
	wire w_dff_A_3Ccg3jVJ7_0;
	wire w_dff_B_hpGPWnPQ3_0;
	wire w_dff_B_cWFmm0rY8_1;
	wire w_dff_B_NKzmPQCu8_1;
	wire w_dff_B_ZGC8ArjM6_1;
	wire w_dff_B_jYQ8yJpf9_0;
	wire w_dff_B_6nFQBuEi0_1;
	wire w_dff_B_WrvP5RP93_0;
	wire w_dff_B_wEjuJzkp5_1;
	wire w_dff_B_YWgJBZQO1_1;
	wire w_dff_B_l0ah2yuI1_1;
	wire w_dff_B_j2Xx3lIg6_0;
	wire w_dff_B_8wHB2uIa9_0;
	wire w_dff_B_MvMuVnvU9_0;
	wire w_dff_B_i4RxXwLI4_0;
	wire w_dff_B_xUTfXL7O8_1;
	wire w_dff_A_ffeh8EW72_0;
	wire w_dff_A_HThBUF9J9_0;
	wire w_dff_A_xQepA7lE2_0;
	wire w_dff_A_TUtlYu8p7_0;
	wire w_dff_B_SIK51O1X2_1;
	wire w_dff_B_QMRvX1Xm5_1;
	wire w_dff_B_5BGTfmIR1_1;
	wire w_dff_B_SkgBOMHA8_1;
	wire w_dff_B_0pyGS53w1_1;
	wire w_dff_B_9KHWRPD95_1;
	wire w_dff_B_Er7mmR2p2_1;
	wire w_dff_B_Oyi3Kmkh2_1;
	wire w_dff_B_ZRijcHmZ5_1;
	wire w_dff_B_DuHaqnlu7_1;
	wire w_dff_B_6ycKs8Ul5_1;
	wire w_dff_B_JojlzJUQ4_1;
	wire w_dff_B_wjYXxjZn8_1;
	wire w_dff_B_xLZueeqH5_1;
	wire w_dff_B_9jmNcFPK6_1;
	wire w_dff_B_huTNExbU1_1;
	wire w_dff_B_dS1H8NTI7_1;
	wire w_dff_B_I12m6zPC5_1;
	wire w_dff_B_3ITbLQEB2_1;
	wire w_dff_B_4bd8CVAd1_1;
	wire w_dff_B_oNO33e4M9_1;
	wire w_dff_B_t6kyo3V09_1;
	wire w_dff_B_cUGmE2xi7_1;
	wire w_dff_B_t8Pisbq56_1;
	wire w_dff_B_aMRC4USe0_1;
	wire w_dff_B_E2Jbsujk9_1;
	wire w_dff_A_bZjkivdt3_2;
	wire w_dff_A_RUiGa3gj2_2;
	wire w_dff_A_1ZccmPtp3_2;
	wire w_dff_A_37x9uh2w9_2;
	wire w_dff_A_Fafs4uuO4_2;
	wire w_dff_A_uO8DG4fo7_2;
	wire w_dff_A_7m5Q2BUn5_2;
	wire w_dff_A_T30i9HG34_2;
	wire w_dff_A_f0wWj8nj2_2;
	wire w_dff_A_Um4hWMoT3_2;
	wire w_dff_A_lWXD2SPz5_2;
	wire w_dff_A_AeIzrj2Q0_2;
	wire w_dff_A_ItY1Ltvz6_2;
	wire w_dff_A_jpDXspEJ9_2;
	wire w_dff_A_5tUe9rvx5_2;
	wire w_dff_A_Yj10R95A7_2;
	wire w_dff_A_ZWJnLsyK3_2;
	wire w_dff_A_9TNq5Mf22_2;
	wire w_dff_A_6Be3uynq4_2;
	wire w_dff_A_36d3tN5Z3_2;
	wire w_dff_A_OQhmWYMb7_2;
	wire w_dff_A_aJTmaqrM1_2;
	wire w_dff_A_gat0Rh1U3_2;
	wire w_dff_A_FWefk98T1_2;
	wire w_dff_A_aqR0O6v62_2;
	wire w_dff_B_B45DUgTt2_0;
	wire w_dff_B_dejdAlZU0_0;
	wire w_dff_B_8PrbAwoS9_0;
	wire w_dff_B_ttBS6XoF1_0;
	wire w_dff_B_tJP0xN0h9_0;
	wire w_dff_B_i0LsO6C66_0;
	wire w_dff_B_IFnR1WK97_0;
	wire w_dff_B_SkSZD2h31_0;
	wire w_dff_B_izG3v0Ph6_0;
	wire w_dff_B_bFVLsN1s0_0;
	wire w_dff_B_7a3WPSu90_0;
	wire w_dff_B_x7a7Svar9_0;
	wire w_dff_B_URYZe7Nn6_0;
	wire w_dff_B_HLv28OkZ4_0;
	wire w_dff_B_Fc1eTT6o0_0;
	wire w_dff_B_VhsXr6N50_0;
	wire w_dff_B_aUw039ji2_0;
	wire w_dff_B_oY37qiuU8_0;
	wire w_dff_B_qhe0Dfjz0_0;
	wire w_dff_B_o5O3sxkA8_0;
	wire w_dff_B_nKOjYhof4_0;
	wire w_dff_B_GunH8rOf0_2;
	wire w_dff_B_TPgcoPC78_1;
	wire w_dff_B_FAOPZv5V7_1;
	wire w_dff_A_YatUVlqb4_0;
	wire w_dff_A_oaMnA73A3_0;
	wire w_dff_A_22uuCQQi7_0;
	wire w_dff_A_F8cigkBA4_0;
	wire w_dff_A_nnxMCx6P2_0;
	wire w_dff_A_G9Qpm1E87_0;
	wire w_dff_A_XucZTZjo5_0;
	wire w_dff_A_NELJFviY2_0;
	wire w_dff_A_w1TryHFu4_0;
	wire w_dff_A_WwSIhvIp1_0;
	wire w_dff_A_rOLPFYlk8_0;
	wire w_dff_A_fJyIdfnP4_0;
	wire w_dff_A_Tzb2EKum7_0;
	wire w_dff_A_ZZ8wciG30_0;
	wire w_dff_A_Nd1rsUZb0_0;
	wire w_dff_A_wcDu4QUg9_0;
	wire w_dff_A_8mFeL7In5_0;
	wire w_dff_A_MYGqcyeX0_0;
	wire w_dff_A_Cc5w5p4o8_0;
	wire w_dff_A_M62Dgl556_0;
	wire w_dff_A_uArWe7To1_2;
	wire w_dff_A_zj7dSgxe2_2;
	wire w_dff_A_6ZLfgkNP9_2;
	wire w_dff_A_EfRGGn2S9_2;
	wire w_dff_A_YHeqpXse7_2;
	wire w_dff_A_RYD1MbQy8_2;
	wire w_dff_A_r0Kp22jR4_2;
	wire w_dff_A_2fPKJ0f32_2;
	wire w_dff_A_DruDHhDh5_2;
	wire w_dff_A_k19TyxIt3_2;
	wire w_dff_A_I7AK9l4r1_2;
	wire w_dff_A_B5Y6mFqO3_0;
	wire w_dff_A_IyvYoxQS1_0;
	wire w_dff_A_IIJH541H5_0;
	wire w_dff_A_QnOub4wR5_0;
	wire w_dff_A_YUXrQRt75_0;
	wire w_dff_A_sw69g0bl1_0;
	wire w_dff_A_cVbZI1bH3_0;
	wire w_dff_A_oxJMVX9b7_0;
	wire w_dff_A_Fyv3BL9r0_0;
	wire w_dff_A_T5GIKLVB9_0;
	wire w_dff_A_65h5CQtB6_0;
	wire w_dff_A_wHmhoBTX2_0;
	wire w_dff_A_4vpslvjp9_0;
	wire w_dff_A_5Fv0ohq61_0;
	wire w_dff_A_ghGyuOvf7_0;
	wire w_dff_A_tAqmXO6k5_0;
	wire w_dff_A_qQ3ncG7g3_0;
	wire w_dff_A_TheF06gb3_0;
	wire w_dff_A_jNwxG6DG5_0;
	wire w_dff_A_ckOVcIE78_0;
	wire w_dff_A_ITruMqol5_2;
	wire w_dff_A_yTwjobei1_2;
	wire w_dff_A_74UCQE2E4_2;
	wire w_dff_A_7Vml2f5s0_2;
	wire w_dff_A_vTixQkao9_2;
	wire w_dff_A_e1eKY6Mv4_2;
	wire w_dff_A_4mvA1vTd7_2;
	wire w_dff_A_rywWiyIt8_2;
	wire w_dff_A_1SHa7NTa3_2;
	wire w_dff_A_vZqizPIh5_2;
	wire w_dff_A_MQ8GbLfP9_2;
	wire w_dff_A_H2fhytxY0_2;
	wire w_dff_A_yL7b2mlw7_2;
	wire w_dff_A_FCfSnQoz9_2;
	wire w_dff_B_sNyM61C42_0;
	wire w_dff_B_VUudYJUS1_0;
	wire w_dff_B_fQhLgF0i8_0;
	wire w_dff_B_fK7jVfCM7_0;
	wire w_dff_B_OzaYxBVF8_0;
	wire w_dff_B_Y7EpLbKs6_0;
	wire w_dff_B_88UUoN8p2_0;
	wire w_dff_B_kAZbV6ZR8_0;
	wire w_dff_B_eSvvKxEW5_0;
	wire w_dff_B_1vlxJ8pG3_0;
	wire w_dff_B_ijCYObGV6_0;
	wire w_dff_B_gzlnwjpf2_0;
	wire w_dff_B_06BbwClh5_0;
	wire w_dff_B_SxUfn8GP6_0;
	wire w_dff_B_9RDZ9AWw3_0;
	wire w_dff_B_Q1EKOq2A8_0;
	wire w_dff_B_L3aqFusI8_0;
	wire w_dff_B_L9TcNWmv1_0;
	wire w_dff_B_hCPLBj4e8_0;
	wire w_dff_B_ZrjqD6Vp2_0;
	wire w_dff_B_JUonUOeP4_1;
	wire w_dff_B_BqxIVWIf3_1;
	wire w_dff_A_XALJo0765_1;
	wire w_dff_A_xvhY1EeL9_1;
	wire w_dff_A_YScRzVKP1_1;
	wire w_dff_A_J7W4h7QO1_1;
	wire w_dff_A_CkVgemj40_1;
	wire w_dff_A_qQuHfedU1_1;
	wire w_dff_A_V9I5XJWd4_1;
	wire w_dff_A_jE6RT3ZK7_1;
	wire w_dff_A_PX3PcX5T5_1;
	wire w_dff_A_FipmS6DT5_1;
	wire w_dff_A_kCZkX5k74_1;
	wire w_dff_A_Z5RO2LRP8_1;
	wire w_dff_A_Wqyy6HN66_1;
	wire w_dff_A_6tdccHF38_1;
	wire w_dff_A_XIRbDcxe1_1;
	wire w_dff_A_Rs0yfhAM9_1;
	wire w_dff_A_ol22gvFD0_1;
	wire w_dff_A_bymHYt0J5_1;
	wire w_dff_A_ziN8tUle8_1;
	wire w_dff_A_ZRzb2x1z0_1;
	wire w_dff_A_wGhzLVgY6_1;
	wire w_dff_A_IWDv9ApJ2_1;
	wire w_dff_A_Glco3OWK0_1;
	wire w_dff_A_YSijWLRB0_1;
	wire w_dff_A_4V5FKOVv6_1;
	wire w_dff_A_UGlWfOtb2_1;
	wire w_dff_A_9lK2CwjN3_1;
	wire w_dff_A_ywXdEx3Y3_1;
	wire w_dff_A_8x00DkiB5_1;
	wire w_dff_A_ZAQPBO0B0_1;
	wire w_dff_A_C332n4v39_1;
	wire w_dff_A_eONCbjqm9_1;
	wire w_dff_A_QWegGdz06_1;
	wire w_dff_A_VNb1TNTD1_1;
	wire w_dff_A_YkE488Kg8_1;
	wire w_dff_A_64PowIwJ9_1;
	wire w_dff_A_Imr3ajC34_1;
	wire w_dff_A_FHmdRqKn5_1;
	wire w_dff_B_eYIAq1GA1_0;
	wire w_dff_B_QYBbsJPU9_0;
	wire w_dff_B_zGh82wrr9_0;
	wire w_dff_B_YsDCrJDR7_0;
	wire w_dff_B_O4Ev20zU0_0;
	wire w_dff_B_n2YgP0Z66_0;
	wire w_dff_B_fK8BoHQY7_0;
	wire w_dff_B_7mOewhfc0_0;
	wire w_dff_B_9irBfDwT6_0;
	wire w_dff_B_OKkB7sDT7_0;
	wire w_dff_B_aa85SRPe9_0;
	wire w_dff_B_fBLLpL2Z6_0;
	wire w_dff_B_sJfJuU600_0;
	wire w_dff_B_EfyyJG1Z1_0;
	wire w_dff_B_WZPliaLL8_0;
	wire w_dff_B_QuuTKFYE9_0;
	wire w_dff_B_qj1QhnIB5_0;
	wire w_dff_B_SbWZlCbF9_0;
	wire w_dff_B_vpNC1Scf1_0;
	wire w_dff_B_cWwYlpGe4_0;
	wire w_dff_B_XV8wNjjV6_1;
	wire w_dff_A_AEZVYED01_2;
	wire w_dff_B_Y9s8MDIv2_0;
	wire w_dff_B_kI4rUX5V0_0;
	wire w_dff_B_zaBMlB7G8_0;
	wire w_dff_B_q3PibDuZ6_0;
	wire w_dff_B_jy8nMNMh8_0;
	wire w_dff_B_t5fQrkdv1_0;
	wire w_dff_B_pIqRasak7_0;
	wire w_dff_B_kj977yMF8_0;
	wire w_dff_B_KXXa3ahS5_0;
	wire w_dff_B_rfPcbXZ02_0;
	wire w_dff_B_nC3fHxGw1_0;
	wire w_dff_B_nPD4e4Xh1_0;
	wire w_dff_B_7fMbkebf2_0;
	wire w_dff_B_TUi0c0967_0;
	wire w_dff_B_h4pD3d1Q3_0;
	wire w_dff_B_0LdIGTMp2_0;
	wire w_dff_B_YaPJtFmK6_0;
	wire w_dff_B_50Nw6W212_0;
	wire w_dff_B_wUvw5KZf0_0;
	wire w_dff_B_wqjCsreb5_1;
	wire w_dff_B_9UvqU0Mw7_1;
	wire w_dff_B_83ZWJmPx7_1;
	wire w_dff_A_4gCQgSGR6_0;
	wire w_dff_A_rlMoYNHS7_0;
	wire w_dff_A_0d8ehUXM9_0;
	wire w_dff_A_sgwSvJ3g2_0;
	wire w_dff_A_9XYPqs8J9_0;
	wire w_dff_A_MtXIsMij8_0;
	wire w_dff_A_vMmRTEqL0_0;
	wire w_dff_A_sKCqViBB7_0;
	wire w_dff_A_REnppv8d2_0;
	wire w_dff_A_9jtUpEyV1_0;
	wire w_dff_A_HdQVBbvz6_0;
	wire w_dff_A_O0Alu5EO1_0;
	wire w_dff_A_Ggo7q89V8_0;
	wire w_dff_A_YuMrfQl95_0;
	wire w_dff_A_xJSz6cr02_0;
	wire w_dff_A_J6eTM2V55_0;
	wire w_dff_A_K0qLzoO09_0;
	wire w_dff_A_Kyd6tigJ2_0;
	wire w_dff_A_VoakkPsj4_2;
	wire w_dff_A_za8zazYM5_2;
	wire w_dff_A_768eAWpu2_2;
	wire w_dff_A_JrluYIVV3_2;
	wire w_dff_A_wOmc1uPo2_2;
	wire w_dff_A_PpzZuoTb4_2;
	wire w_dff_A_aRnrflxL7_2;
	wire w_dff_A_MhQ7Nci84_2;
	wire w_dff_A_OKMVwSmv4_2;
	wire w_dff_A_TPybtCcY5_2;
	wire w_dff_A_mrGswC7c6_2;
	wire w_dff_A_Ls1thhwE1_2;
	wire w_dff_A_GFVJTBvp6_2;
	wire w_dff_A_CeD87hr09_2;
	wire w_dff_A_iyvt8MIR3_2;
	wire w_dff_A_nE0KVern0_2;
	wire w_dff_A_vfNadHEl0_2;
	wire w_dff_A_TmokUw5w2_2;
	wire w_dff_A_MKO4dv4O9_2;
	wire w_dff_A_PPOCxUvs9_0;
	wire w_dff_A_6XJVNJyQ8_0;
	wire w_dff_A_oLboJLN71_0;
	wire w_dff_A_JbqWqdSV6_0;
	wire w_dff_A_mPWSUyxJ4_0;
	wire w_dff_A_yrImN39F7_0;
	wire w_dff_A_2aiEzahd3_0;
	wire w_dff_A_95yoRKHZ7_0;
	wire w_dff_A_TZRiJMdD0_0;
	wire w_dff_A_fX256Ym36_0;
	wire w_dff_A_8ofDLLrF9_0;
	wire w_dff_A_jBVkFGap8_0;
	wire w_dff_A_HICobnjJ7_0;
	wire w_dff_A_ETtM8T6Z3_0;
	wire w_dff_A_JY1n396d6_0;
	wire w_dff_A_7AQRFNeS9_0;
	wire w_dff_A_7Swbm09q8_0;
	wire w_dff_A_g1Tf0iTQ7_2;
	wire w_dff_A_m70sggur0_2;
	wire w_dff_A_FDtVVnMn4_2;
	wire w_dff_A_KIXZiPsY5_2;
	wire w_dff_A_4kChQZ8h5_2;
	wire w_dff_A_nmwvYoTM2_2;
	wire w_dff_A_d5Ryocg67_2;
	wire w_dff_A_HMukPqrW3_2;
	wire w_dff_A_yVNf7jod6_2;
	wire w_dff_A_20b70NDv3_2;
	wire w_dff_A_7E1tYVwx3_2;
	wire w_dff_A_ZkvBa6zQ2_2;
	wire w_dff_A_sKkZe3G20_2;
	wire w_dff_A_jfcvFFFJ0_2;
	wire w_dff_A_ItTHYXAt0_2;
	wire w_dff_A_SIDaAc2k1_2;
	wire w_dff_A_CWC3y3JR5_2;
	wire w_dff_A_ZYuvNFx13_2;
	wire w_dff_A_TLCH7n487_2;
	wire w_dff_A_pjKoofEh2_2;
	wire w_dff_B_J60eXKgG2_0;
	wire w_dff_B_WSRhJrnt2_0;
	wire w_dff_B_j4bXQBwu5_0;
	wire w_dff_B_6bYcj14p9_0;
	wire w_dff_B_YRZTNHsg3_0;
	wire w_dff_B_VL9aqalw4_0;
	wire w_dff_B_3Wqpspjr2_0;
	wire w_dff_B_A3oFkFji7_0;
	wire w_dff_B_t2bE6uZk2_0;
	wire w_dff_B_etWH6cnO7_0;
	wire w_dff_B_HkX3qNgM9_0;
	wire w_dff_B_pkh93CVQ2_0;
	wire w_dff_B_xAMOHBZi3_0;
	wire w_dff_B_UsQFK8bR6_0;
	wire w_dff_B_XcDDGPAj4_0;
	wire w_dff_B_KFPTwAig1_0;
	wire w_dff_B_rmRVjMwl8_0;
	wire w_dff_B_ZH7tg8vm3_0;
	wire w_dff_B_qn1WiwTn9_0;
	wire w_dff_B_bsKDHyqd4_0;
	wire w_dff_B_1iiDpNCJ1_2;
	wire w_dff_B_ByI9NIUN9_1;
	wire w_dff_B_GERUinjS1_1;
	wire w_dff_A_DmdTJJ9j7_1;
	wire w_dff_A_qWlmct5i8_1;
	wire w_dff_A_RAE24eSo6_1;
	wire w_dff_A_I54Bc3Bz4_1;
	wire w_dff_A_apWsffSX3_1;
	wire w_dff_A_mrRvZvLn9_1;
	wire w_dff_A_D6ZeCKFF3_1;
	wire w_dff_A_jO3u9WTG8_1;
	wire w_dff_A_gbFroE9F2_1;
	wire w_dff_A_3hMaGZQG2_1;
	wire w_dff_A_BD36ye7G7_1;
	wire w_dff_A_Ei9yp1054_1;
	wire w_dff_A_U2v2jdlk9_1;
	wire w_dff_A_2kc4YKij9_1;
	wire w_dff_A_xd4xm3Fg1_1;
	wire w_dff_A_y4tLAUPo7_1;
	wire w_dff_A_MoUaTE9L8_1;
	wire w_dff_A_6oNJnF3U1_1;
	wire w_dff_A_4xcqPKm27_1;
	wire w_dff_A_UMninGSU0_2;
	wire w_dff_A_GC8pYjNn8_2;
	wire w_dff_A_axcAwmoL8_2;
	wire w_dff_A_hUEnJQpu2_2;
	wire w_dff_A_sNIPA7qp5_2;
	wire w_dff_A_PLhEKwZP8_2;
	wire w_dff_A_I4IF0Pxw3_2;
	wire w_dff_A_MKgQu3iE6_2;
	wire w_dff_A_YiZcyg1D0_2;
	wire w_dff_A_rCdV2gmw9_2;
	wire w_dff_A_i1gwYgew8_2;
	wire w_dff_A_PyK2QKkD6_2;
	wire w_dff_A_VXVyJfZ18_2;
	wire w_dff_A_05ATyDD63_2;
	wire w_dff_A_Gvdq3EKN6_2;
	wire w_dff_A_WHRqcrMG6_2;
	wire w_dff_A_qwruWkYt4_2;
	wire w_dff_A_VZe651fN8_2;
	wire w_dff_A_Il1SW8DM7_2;
	wire w_dff_A_tRYBKt5n9_2;
	wire w_dff_A_VkXPZzYQ4_1;
	wire w_dff_A_9g54clkG4_1;
	wire w_dff_A_zUaKOAz37_1;
	wire w_dff_A_uZQOUO5N9_1;
	wire w_dff_A_z4AncOV57_1;
	wire w_dff_A_lo1Qsoca6_1;
	wire w_dff_A_FIJSdwWl5_1;
	wire w_dff_A_ZT2pKGJ54_1;
	wire w_dff_A_xvTq5f9H3_1;
	wire w_dff_A_ohbwn4DH0_1;
	wire w_dff_A_Ap9v18aT1_1;
	wire w_dff_A_83ihjgF47_1;
	wire w_dff_A_LZeWXIrJ9_1;
	wire w_dff_A_tukI4Hbu1_1;
	wire w_dff_A_AwnaBnnP8_1;
	wire w_dff_A_p8ZPVSMX4_1;
	wire w_dff_A_aDy7lTlm0_1;
	wire w_dff_A_I1luDF322_1;
	wire w_dff_A_2M1RsakX4_1;
	wire w_dff_A_CT1pJcIv8_2;
	wire w_dff_A_QaHUIWPk4_2;
	wire w_dff_A_dY9oIj3R5_2;
	wire w_dff_A_SPvbf5KQ7_2;
	wire w_dff_A_r02y06yv6_2;
	wire w_dff_A_3qOMgvzZ8_2;
	wire w_dff_A_2fLrrPOJ2_2;
	wire w_dff_A_3H3bu0dK9_2;
	wire w_dff_A_EP9lU7jf9_2;
	wire w_dff_A_iH4ZRY9f4_2;
	wire w_dff_A_UaCf8izn3_2;
	wire w_dff_A_PKpybt2R3_2;
	wire w_dff_A_LeQzXgpj2_2;
	wire w_dff_A_qITQm8Z94_2;
	wire w_dff_A_4mAmj4Yt2_2;
	wire w_dff_A_ynEeKY1O4_2;
	wire w_dff_A_hLZQ4Cn07_2;
	wire w_dff_A_9QRPuVhF6_2;
	wire w_dff_A_hNiW7AmZ6_2;
	wire w_dff_A_hd8QYJlY8_2;
	wire w_dff_B_VgcngmYy7_0;
	wire w_dff_B_u3FmbG4H7_0;
	wire w_dff_B_PNQGyG9Z1_0;
	wire w_dff_B_ziHiVmR14_0;
	wire w_dff_B_c3tASEs72_0;
	wire w_dff_B_hrHc12Ln7_0;
	wire w_dff_B_SXtFyYYv4_0;
	wire w_dff_B_eWu49nh12_0;
	wire w_dff_B_nQcQNIhA2_0;
	wire w_dff_B_ur18KuvB7_0;
	wire w_dff_B_hcoQKYzl9_0;
	wire w_dff_B_Opo8cy6A0_0;
	wire w_dff_B_ers6BkD50_0;
	wire w_dff_B_SPvuNKpO4_0;
	wire w_dff_B_LPSobsfJ6_0;
	wire w_dff_B_6BADGxjz4_0;
	wire w_dff_B_U719I3d97_0;
	wire w_dff_B_9lWbF8ew9_0;
	wire w_dff_B_OKrlPkE78_0;
	wire w_dff_B_YZF84n0Q0_0;
	wire w_dff_A_oG5NCBMF8_2;
	wire w_dff_B_TggzarqU3_2;
	wire w_dff_B_P8Q07vcW5_1;
	wire w_dff_B_oWTo4IZ70_0;
	wire w_dff_B_MWkd3yfS8_0;
	wire w_dff_B_EiKIeVIS5_0;
	wire w_dff_B_PTXofejd0_0;
	wire w_dff_B_18fZtD3f9_0;
	wire w_dff_B_T60S0ktL9_0;
	wire w_dff_B_XeY8b9oO3_0;
	wire w_dff_B_CK4N7eof6_0;
	wire w_dff_B_GFi2iK3k4_0;
	wire w_dff_B_Cc6c2iMY4_0;
	wire w_dff_B_9IWprNb41_0;
	wire w_dff_B_FYCKJ5LT1_0;
	wire w_dff_B_W6vLBPDZ3_0;
	wire w_dff_B_X759oBYN0_0;
	wire w_dff_B_E7AYLJE73_0;
	wire w_dff_B_ODECBc4B5_0;
	wire w_dff_B_KHm83jYH8_0;
	wire w_dff_B_tLvTM9XN0_0;
	wire w_dff_B_wucxeoWg8_0;
	wire w_dff_B_g02a7w813_2;
	wire w_dff_B_wH6ZXEK84_1;
	wire w_dff_B_LV9tmisc5_1;
	wire w_dff_B_gCFCo7wU8_1;
	wire w_dff_A_5f3rJesb7_0;
	wire w_dff_A_GFGDxHB55_0;
	wire w_dff_A_UPwfE7ja2_0;
	wire w_dff_A_KaGLihMo7_0;
	wire w_dff_A_XPY1G27t6_0;
	wire w_dff_A_otABIdyQ9_0;
	wire w_dff_A_Z9P19O0e1_0;
	wire w_dff_A_Iop6I1MH0_0;
	wire w_dff_A_tg2Qaj433_0;
	wire w_dff_A_MkmjU6aP7_0;
	wire w_dff_A_uPChqG4i2_0;
	wire w_dff_A_pApaFv0r8_0;
	wire w_dff_A_0kcoK7jF6_0;
	wire w_dff_A_HUdzpgs96_0;
	wire w_dff_A_qBX1WSOm7_0;
	wire w_dff_A_pLczTBe23_0;
	wire w_dff_A_GNABojvH5_0;
	wire w_dff_A_ProXiB0p1_0;
	wire w_dff_A_ZArgnJNj4_2;
	wire w_dff_A_uFtIcpUa3_2;
	wire w_dff_A_ZViEz3Tc8_2;
	wire w_dff_A_cbDFD91B8_2;
	wire w_dff_A_1Rk7d5hL9_2;
	wire w_dff_A_vDMqAGR29_2;
	wire w_dff_A_Gz14ckvu9_2;
	wire w_dff_A_qMhmKxNO2_2;
	wire w_dff_A_9FNSNHVl3_2;
	wire w_dff_A_f7AAWilR6_2;
	wire w_dff_A_xAdEoUSC8_2;
	wire w_dff_A_DhdHWnMz4_2;
	wire w_dff_A_oK6VCFfR3_2;
	wire w_dff_A_tvwMDykL8_2;
	wire w_dff_A_89qTCW2n0_2;
	wire w_dff_A_uK5rKovo2_2;
	wire w_dff_A_Zq8Ea4cw1_2;
	wire w_dff_A_aKN8QaHX4_2;
	wire w_dff_A_w2NP7IaK8_2;
	wire w_dff_A_ZEpNc4jf7_0;
	wire w_dff_A_zcIJje8M8_0;
	wire w_dff_A_X20Sckfq9_0;
	wire w_dff_A_UUUjfqCD6_0;
	wire w_dff_A_VAI9XjON3_0;
	wire w_dff_A_N2x3levN2_0;
	wire w_dff_A_afVVJGMx7_0;
	wire w_dff_A_Qn49o1RX4_0;
	wire w_dff_A_NQColUxj0_0;
	wire w_dff_A_smWzWTeG8_0;
	wire w_dff_A_xdOE0AV27_0;
	wire w_dff_A_TCW1t95Q5_0;
	wire w_dff_A_YwgRfHf62_0;
	wire w_dff_A_G5kEngBQ4_0;
	wire w_dff_A_a4TUhWox8_0;
	wire w_dff_A_qzZ10NaD8_0;
	wire w_dff_A_bkjNZIKN0_0;
	wire w_dff_A_O9lhhJ3D8_2;
	wire w_dff_A_ZvCc4pju1_2;
	wire w_dff_A_k4Wijpaf9_2;
	wire w_dff_A_A80fwNxP5_2;
	wire w_dff_A_FOaS4qm72_2;
	wire w_dff_A_NEaqVqWG9_2;
	wire w_dff_A_4KKowJc26_2;
	wire w_dff_A_zFg4PUDz9_2;
	wire w_dff_A_GJLMnXCg4_2;
	wire w_dff_A_y6jj5itR9_2;
	wire w_dff_A_utr5CoJO4_2;
	wire w_dff_A_GWBbCcyn4_2;
	wire w_dff_A_Q9hckj7v5_2;
	wire w_dff_A_5gYJdO0q7_2;
	wire w_dff_A_JO0x2C7B1_2;
	wire w_dff_A_uVsnAcgH3_2;
	wire w_dff_A_833IOcGk4_2;
	wire w_dff_A_L1tVDxQ90_2;
	wire w_dff_A_nc6MxPa65_2;
	wire w_dff_A_fggixee15_2;
	wire w_dff_B_mZk8DadO8_0;
	wire w_dff_B_cVT2ypDr2_0;
	wire w_dff_B_v2xyDfLa6_0;
	wire w_dff_B_X6ceblqR4_0;
	wire w_dff_B_natTV8HQ5_0;
	wire w_dff_B_kRU1cT6X6_0;
	wire w_dff_B_kp5I4s5E8_0;
	wire w_dff_B_QOZYkWO01_0;
	wire w_dff_B_7OO2PNT44_0;
	wire w_dff_B_2u48I0ZQ2_0;
	wire w_dff_B_W3SHrZaa6_0;
	wire w_dff_B_yE3crgXW6_0;
	wire w_dff_B_yjJUCC3x5_0;
	wire w_dff_B_AuFJkS3l9_0;
	wire w_dff_B_fztX6vIt0_0;
	wire w_dff_B_RhWaCaTT4_0;
	wire w_dff_B_Jz9qHEXU8_0;
	wire w_dff_B_nFMKQL577_0;
	wire w_dff_B_ubgztRBW1_0;
	wire w_dff_B_zlsu6uTC2_1;
	wire w_dff_B_tXKxrf9s1_1;
	wire w_dff_B_ABsc0nYs4_1;
	wire w_dff_A_RDLo1Q703_0;
	wire w_dff_A_8gT6Xo5p5_0;
	wire w_dff_A_0pzcnxNl7_0;
	wire w_dff_A_smbNrJg58_0;
	wire w_dff_A_B9JONuk91_0;
	wire w_dff_A_gNqVIcRp2_0;
	wire w_dff_A_p5R2bQi48_1;
	wire w_dff_A_V4oXL9y83_0;
	wire w_dff_A_cnXsDLqu5_0;
	wire w_dff_A_o0ci5aYa7_0;
	wire w_dff_A_9L5JHhJU6_0;
	wire w_dff_A_qGxOKaZp3_1;
	wire w_dff_A_JUUW9lsD8_1;
	wire w_dff_A_BNNter448_0;
	wire w_dff_A_qZO2Lkdt2_0;
	wire w_dff_A_e6wOR5rI7_0;
	wire w_dff_A_oo6diNym5_0;
	wire w_dff_A_0adyCNG52_0;
	wire w_dff_A_iKHdrdEq0_0;
	wire w_dff_A_0CrxWVcA1_1;
	wire w_dff_B_2zwCAScy4_0;
	wire w_dff_B_Mx9K13cZ6_0;
	wire w_dff_B_nBvGElPF9_0;
	wire w_dff_B_VV1WvhOR8_0;
	wire w_dff_B_tcUsRVJQ0_0;
	wire w_dff_B_mkWUecon1_0;
	wire w_dff_B_GoHOyCPM4_0;
	wire w_dff_B_XvcaOzwA5_0;
	wire w_dff_B_VHn29TaX9_0;
	wire w_dff_B_BSC9Ld8P6_0;
	wire w_dff_B_Vb3IcSzo1_0;
	wire w_dff_B_Y9BEo8R88_0;
	wire w_dff_B_XydEaswq6_0;
	wire w_dff_B_oHanbBGp4_0;
	wire w_dff_B_W045XdAy6_0;
	wire w_dff_B_wmj0R0Sx4_0;
	wire w_dff_B_ihZKWXYs2_0;
	wire w_dff_B_AiOmB4mL5_0;
	wire w_dff_B_qz6367Se3_0;
	wire w_dff_B_GW0o3jnx6_0;
	wire w_dff_B_dPM72rwn1_1;
	wire w_dff_B_WqFWozgh4_1;
	wire w_dff_B_mZ5mP0hv6_1;
	wire w_dff_B_aYioYtRr2_1;
	wire w_dff_B_QxQXc6BT8_1;
	wire w_dff_B_jtKmuv6R5_1;
	wire w_dff_B_DkGma15y7_1;
	wire w_dff_B_5ayhU0Rg2_1;
	wire w_dff_B_JC05rPA08_1;
	wire w_dff_B_ATsFikNj9_1;
	wire w_dff_B_tZNoVLZI3_1;
	wire w_dff_B_cmuIQCN52_1;
	wire w_dff_B_HHTOpmCQ3_1;
	wire w_dff_B_HE99HN4o1_1;
	wire w_dff_B_uK9Hl7HN7_1;
	wire w_dff_B_MQ9FhYmA6_1;
	wire w_dff_B_QPBFYZcg9_1;
	wire w_dff_B_fYORsTpe3_1;
	wire w_dff_B_EcxWEDzd4_1;
	wire w_dff_B_2N7sWeEP9_1;
	wire w_dff_B_aM7Hh88Z6_1;
	wire w_dff_A_6ARgsfXK6_0;
	wire w_dff_A_2dPucS1o4_1;
	wire w_dff_B_n0fNFoP04_0;
	wire w_dff_B_HZpmXYVr6_1;
	wire w_dff_B_mZiglbwN2_1;
	wire w_dff_B_9SU1YpQd1_1;
	wire w_dff_B_QHJWhX3r1_1;
	wire w_dff_B_uaVPONxv7_1;
	wire w_dff_B_fHKgcpxq5_1;
	wire w_dff_B_jfhtiu9j5_1;
	wire w_dff_B_mtfiZGou8_1;
	wire w_dff_B_45DQP7MI3_1;
	wire w_dff_B_QZrZVwZg6_1;
	wire w_dff_B_yE8vwQXY9_1;
	wire w_dff_B_PiPz5vEE5_1;
	wire w_dff_B_9k9lo8dS9_1;
	wire w_dff_B_NOAdkUrY0_1;
	wire w_dff_B_Ri2MbYJE4_1;
	wire w_dff_B_EmsGaU8w7_1;
	wire w_dff_B_rmMndIEr1_1;
	wire w_dff_B_9XnAlZqg0_1;
	wire w_dff_B_qHZDVASq7_1;
	wire w_dff_B_9O0W9hO07_1;
	wire w_dff_B_ud4zDNMc5_1;
	wire w_dff_A_HJZRrLEG4_0;
	wire w_dff_A_zKLX45dN3_2;
	wire w_dff_A_UUwchZia9_0;
	wire w_dff_A_RlKZcSQj8_0;
	wire w_dff_A_Tli91gTS6_1;
	wire w_dff_A_8M2KqIGQ8_0;
	wire w_dff_A_8P8FX6qV1_0;
	wire w_dff_A_CckW1MhG9_0;
	wire w_dff_A_oe4XpMmv9_0;
	wire w_dff_A_7EZ4YDgG6_0;
	wire w_dff_A_VoSiUYyz2_0;
	wire w_dff_A_zN00DOpl0_0;
	wire w_dff_A_hFwu1MYn0_0;
	wire w_dff_A_Uh1Kfn9T3_0;
	wire w_dff_A_YtWZNf8k5_0;
	wire w_dff_A_qYXjQuKy8_0;
	wire w_dff_A_vDJTTgAp5_1;
	wire w_dff_A_DlPldBzq0_1;
	wire w_dff_A_8oSnNPd36_1;
	wire w_dff_A_3J7YtBlR4_1;
	wire w_dff_B_kltcvlBT9_3;
	wire w_dff_B_uQ3hNHun0_3;
	wire w_dff_B_DiW1C9fY2_3;
	wire w_dff_B_I17bN32S5_3;
	wire w_dff_B_hWSMz0cz6_3;
	wire w_dff_B_VEBeYxTG1_3;
	wire w_dff_B_HDZl0wU33_3;
	wire w_dff_B_nKJuCJj05_3;
	wire w_dff_B_gH9XOfcv5_3;
	wire w_dff_B_WuxwULkX2_0;
	wire w_dff_A_kcz5qDe10_0;
	wire w_dff_B_oNhKQnch1_0;
	wire w_dff_B_t98oNZmA4_0;
	wire w_dff_B_fXhRwIXX8_0;
	wire w_dff_B_eT2XgNwZ4_0;
	wire w_dff_B_x1vGDLVW9_0;
	wire w_dff_B_exUFEdiW6_0;
	wire w_dff_B_tP5Wgawe9_0;
	wire w_dff_B_o97lgQwU2_0;
	wire w_dff_B_ykrhYx5y7_0;
	wire w_dff_B_SPfTink03_0;
	wire w_dff_B_mG55dgay0_0;
	wire w_dff_B_j0r0l8Nh8_0;
	wire w_dff_B_OB95ABOx9_0;
	wire w_dff_B_jVDwKCqR3_0;
	wire w_dff_B_F7sHR3l28_0;
	wire w_dff_B_rEe3ADAP1_0;
	wire w_dff_B_BSFEM9Il6_0;
	wire w_dff_B_IFjCnL9p5_0;
	wire w_dff_B_LMyJSMy41_0;
	wire w_dff_B_3YGGGiVE7_2;
	wire w_dff_B_vpfIBe4U6_2;
	wire w_dff_B_sdn6Tn8o5_2;
	wire w_dff_B_3DPhSuQZ6_1;
	wire w_dff_B_Vx59He5A6_1;
	wire w_dff_B_kLo2r7RI9_1;
	wire w_dff_B_uAapR5Qn6_1;
	wire w_dff_B_dPcBdxqo8_1;
	wire w_dff_B_QuQvfOdS3_1;
	wire w_dff_B_RixEefj14_1;
	wire w_dff_B_sbpHS0em0_1;
	wire w_dff_B_b20BfPNH2_1;
	wire w_dff_B_sJ9orpA58_1;
	wire w_dff_B_AImiS8TP9_1;
	wire w_dff_B_oBDNuw0b4_1;
	wire w_dff_B_ZwxUGoIJ7_1;
	wire w_dff_B_5XWr8qUk4_1;
	wire w_dff_B_Ac9kbomT8_1;
	wire w_dff_B_z39GyPid4_1;
	wire w_dff_B_Q9Q1JZKq3_0;
	wire w_dff_B_vfijBjnP6_0;
	wire w_dff_B_IdzVWRJ20_0;
	wire w_dff_B_FuLaBeJw9_0;
	wire w_dff_B_j3URnBDD9_0;
	wire w_dff_B_5ta3wDFs3_0;
	wire w_dff_B_DMhh5lqb8_0;
	wire w_dff_B_oJEqyHun7_0;
	wire w_dff_B_LvgzSzjn0_0;
	wire w_dff_B_UlI2Nhbz5_1;
	wire w_dff_B_5spP29TG4_1;
	wire w_dff_B_rmvr7Zh08_1;
	wire w_dff_B_ZdKFumnR9_1;
	wire w_dff_A_U6838mNR2_0;
	wire w_dff_A_s7AfrquI6_0;
	wire w_dff_A_i5S6ZHBl3_0;
	wire w_dff_A_hhmWvY035_0;
	wire w_dff_A_pMfUvf6u9_0;
	wire w_dff_A_MkXZOu1o5_0;
	wire w_dff_A_FInBIvAe5_1;
	wire w_dff_B_QsVLWo5M4_1;
	wire w_dff_B_MLzapeKq4_1;
	wire w_dff_B_egi2egYW9_1;
	wire w_dff_B_2KP0CUQ02_1;
	wire w_dff_B_uV2F0mFV7_1;
	wire w_dff_B_K3fJ4o1u7_1;
	wire w_dff_B_O08tIw8b7_1;
	wire w_dff_B_g2qFy7mZ6_1;
	wire w_dff_B_zN12jrPW8_1;
	wire w_dff_B_xumPm5G10_1;
	wire w_dff_B_FP9SyRB59_1;
	wire w_dff_B_ApvnlSWa4_0;
	wire w_dff_B_AbYxge710_0;
	wire w_dff_B_NdOS22z31_0;
	wire w_dff_B_D2sojhaL3_0;
	wire w_dff_B_390DoZ1d2_0;
	wire w_dff_B_iqFcjq4L1_0;
	wire w_dff_B_GbydITx23_0;
	wire w_dff_A_gxZKuS240_1;
	wire w_dff_A_bVg8zjmE1_1;
	wire w_dff_A_VDh4o9zL3_1;
	wire w_dff_A_ZLXJuPVY7_1;
	wire w_dff_A_cgmkJVQL6_1;
	wire w_dff_B_MEDCZDtm7_1;
	wire w_dff_B_3ssWQ6XL7_1;
	wire w_dff_B_hrULTG3r5_1;
	wire w_dff_B_DXRqprTM4_1;
	wire w_dff_B_ARb2QoPd3_1;
	wire w_dff_B_9D7e0xVP8_1;
	wire w_dff_B_vtl9k3e31_1;
	wire w_dff_B_ppcvgk152_1;
	wire w_dff_A_LLViKpil3_0;
	wire w_dff_A_VYvhuAvX4_0;
	wire w_dff_A_xMrswLls9_0;
	wire w_dff_A_TIcULKQy2_0;
	wire w_dff_A_tSoCaoAp5_1;
	wire w_dff_A_AyyJTQSO9_1;
	wire w_dff_B_p2WWs4dO1_1;
	wire w_dff_B_hFkVxJ4x7_1;
	wire w_dff_B_z9pPafwW7_1;
	wire w_dff_B_7UeFKED25_1;
	wire w_dff_B_VKaHcStD9_1;
	wire w_dff_B_DKncdiQB2_1;
	wire w_dff_B_vnDkYqHq3_1;
	wire w_dff_B_WL1pQyqE5_1;
	wire w_dff_B_cwKcXo590_1;
	wire w_dff_B_ATwA34fK2_1;
	wire w_dff_B_ofV6NNc53_1;
	wire w_dff_B_2HI67dHS5_1;
	wire w_dff_B_ecLNolU72_1;
	wire w_dff_B_xtLdzSf50_1;
	wire w_dff_B_IgSpwvgU3_1;
	wire w_dff_B_iGh2f43X3_1;
	wire w_dff_B_cHymfyTx3_1;
	wire w_dff_B_V6AwSBvI4_1;
	wire w_dff_B_dEHTAsTF1_1;
	wire w_dff_B_6DI3sagl7_1;
	wire w_dff_B_BsGvu4lc8_1;
	wire w_dff_B_GhOkG0605_1;
	wire w_dff_B_HXUnzWRY4_1;
	wire w_dff_B_gEZPRPo12_1;
	wire w_dff_B_02CnrUPQ5_1;
	wire w_dff_B_hA8dwoGV0_1;
	wire w_dff_B_WuSlpCqL1_1;
	wire w_dff_B_2IAefZUF1_1;
	wire w_dff_B_XsGKdWxJ2_1;
	wire w_dff_B_jPyZcYFn7_1;
	wire w_dff_B_2dmljysv7_1;
	wire w_dff_B_aVrKJl0A3_1;
	wire w_dff_B_TerfcU185_1;
	wire w_dff_B_HkaWFrb58_1;
	wire w_dff_B_uuDGuNni8_1;
	wire w_dff_B_8VGlEAWL1_1;
	wire w_dff_B_C8xH7zdg3_1;
	wire w_dff_B_swYH9Qb04_1;
	wire w_dff_B_ISr2g28k4_1;
	wire w_dff_B_7CRJ4Ji20_1;
	wire w_dff_B_eRr7kqYR1_1;
	wire w_dff_B_0Zk4YnWz7_1;
	wire w_dff_B_KuMbj2xW9_1;
	wire w_dff_B_n7YbBHeH6_1;
	wire w_dff_B_qYFE3t1B0_1;
	wire w_dff_B_xh3eOoMT7_1;
	wire w_dff_B_sQBYefKu6_1;
	wire w_dff_B_UUPINPiN2_1;
	wire w_dff_B_G35Dpjh71_1;
	wire w_dff_B_JUdnOlon2_1;
	wire w_dff_B_wLOgCkTt1_1;
	wire w_dff_B_x6mYwETw3_1;
	wire w_dff_B_iLjUAyAc7_1;
	wire w_dff_B_4hANBpo36_1;
	wire w_dff_B_U77XHhe59_1;
	wire w_dff_B_R5eitxjB8_1;
	wire w_dff_B_U8buMZBn5_1;
	wire w_dff_B_DgmosfyD2_1;
	wire w_dff_B_wPc01Xff2_1;
	wire w_dff_B_o4O4XsoW3_1;
	wire w_dff_B_fh4ifOrf6_1;
	wire w_dff_B_Rjh3rheS3_1;
	wire w_dff_B_uMpaWiJB7_1;
	wire w_dff_B_YCPthgoq9_1;
	wire w_dff_B_bPsVyb8j1_1;
	wire w_dff_B_Fr8ZR9ph3_1;
	wire w_dff_B_in9njksg0_1;
	wire w_dff_B_L1bK1fbl9_1;
	wire w_dff_B_O0kiAZ539_1;
	wire w_dff_B_odToLabO9_1;
	wire w_dff_B_GWMxj4ZE5_1;
	wire w_dff_B_riJkI51u7_1;
	wire w_dff_B_UmXLvvYf4_1;
	wire w_dff_B_re8ILEbE4_1;
	wire w_dff_B_0ls9iHpe0_1;
	wire w_dff_B_N5C4SXT00_0;
	wire w_dff_B_PKVlJO5q2_0;
	wire w_dff_B_dBsGJJeR7_0;
	wire w_dff_B_YIbd9Jui4_0;
	wire w_dff_B_pivutCvQ4_0;
	wire w_dff_B_KOJPPlSy6_0;
	wire w_dff_B_oO6QsDMN6_0;
	wire w_dff_B_LNTsN6IM3_0;
	wire w_dff_B_8HibIQqz7_0;
	wire w_dff_B_K5sujEbX8_0;
	wire w_dff_B_toa6koN10_1;
	wire w_dff_B_6soc72gs1_1;
	wire w_dff_B_G8Mktwtq9_1;
	wire w_dff_B_n1mkz8xW1_1;
	wire w_dff_B_IqFng8PM3_1;
	wire w_dff_B_6GmatHib3_1;
	wire w_dff_B_SC9cXjYy2_1;
	wire w_dff_B_A7MjYjF48_1;
	wire w_dff_B_evwuM9UD2_1;
	wire w_dff_B_0ALb2b7X8_1;
	wire w_dff_B_2RwCbKtr9_1;
	wire w_dff_B_HwRS2yqS1_1;
	wire w_dff_B_vnzkMDfK1_1;
	wire w_dff_B_10NKltzk4_1;
	wire w_dff_B_N4OMMBhQ3_1;
	wire w_dff_B_Zit3e8cd9_1;
	wire w_dff_B_HLhD5N0M9_1;
	wire w_dff_B_ijBLdRBO8_0;
	wire w_dff_B_9aXorsj56_2;
	wire w_dff_B_H48A0kQm2_2;
	wire w_dff_B_VgeiRaJZ6_2;
	wire w_dff_B_AZvcbzd63_0;
	wire w_dff_B_TkkLXyD15_0;
	wire w_dff_B_qqqY8pEI5_0;
	wire w_dff_B_gDRjJvBD3_0;
	wire w_dff_B_ZVYnWGNU6_0;
	wire w_dff_B_cjBEo7AV0_0;
	wire w_dff_B_w6xcHZAP3_0;
	wire w_dff_B_pWYAyKHA0_0;
	wire w_dff_B_TEqgDbHD6_0;
	wire w_dff_B_3NlkGlqq2_0;
	wire w_dff_B_RQas0pJ69_0;
	wire w_dff_B_vU9Gs3iL9_0;
	wire w_dff_B_uGnDQR4r1_0;
	wire w_dff_B_vrEkEr026_0;
	wire w_dff_B_iQctaIDJ8_0;
	wire w_dff_B_nlPrNay41_0;
	wire w_dff_B_EoMrwKBg1_0;
	wire w_dff_B_SpQvWwNX4_0;
	wire w_dff_B_JnaAnNOS8_0;
	wire w_dff_B_exdElFVE8_0;
	wire w_dff_B_TbFIqqaD0_2;
	wire w_dff_B_m7hFPIXg9_2;
	wire w_dff_B_Rz0P6yzV7_2;
	wire w_dff_B_ssWr4pTK1_1;
	wire w_dff_B_yu53a9v41_1;
	wire w_dff_B_TGO8iULe2_1;
	wire w_dff_B_A37AbIAp2_1;
	wire w_dff_B_wvrreFmq1_1;
	wire w_dff_B_KTL9enEE4_1;
	wire w_dff_B_v4tyJpsv9_1;
	wire w_dff_B_0IwtZsoK9_1;
	wire w_dff_B_IfuORuYE1_1;
	wire w_dff_B_bLJBhXpd3_1;
	wire w_dff_B_pbdaXscH8_1;
	wire w_dff_B_34y1FdMT2_1;
	wire w_dff_B_RcYZ3R6z5_1;
	wire w_dff_B_FP5SvLkv9_1;
	wire w_dff_B_mHTpKiRG6_1;
	wire w_dff_B_ko9Gnr9s4_1;
	wire w_dff_B_uu31VkD16_0;
	wire w_dff_B_vatYfM3q5_0;
	wire w_dff_B_HTpWDVxP1_0;
	wire w_dff_B_4tC1GQv50_0;
	wire w_dff_B_uwRaskC55_0;
	wire w_dff_B_FdbOHdph3_0;
	wire w_dff_B_eC63qPAp6_0;
	wire w_dff_B_rvPwzAcj6_0;
	wire w_dff_B_TgL3nZaF8_0;
	wire w_dff_B_bhsRT5yD6_0;
	wire w_dff_A_P84LKBiu6_1;
	wire w_dff_A_o8CzVpOe9_1;
	wire w_dff_A_JxHJl6d94_1;
	wire w_dff_B_L640B3lG0_1;
	wire w_dff_B_qq3Zf2UL4_3;
	wire w_dff_B_35rSU6h96_1;
	wire w_dff_A_n93D60cc3_0;
	wire w_dff_A_ie8bqfPa0_0;
	wire w_dff_A_IBnOEhUf2_0;
	wire w_dff_A_a2aQVqUY5_0;
	wire w_dff_A_yxULFsEi1_0;
	wire w_dff_A_0D4zN2s97_0;
	wire w_dff_A_Ds3lcUdV8_0;
	wire w_dff_A_T2vrZu4X7_0;
	wire w_dff_A_Y41NaXej2_0;
	wire w_dff_A_1k0tT0x53_0;
	wire w_dff_A_tyqGwJg34_0;
	wire w_dff_A_xRxgL4oh5_1;
	wire w_dff_A_bR7YuVXX4_1;
	wire w_dff_B_7bcgBnsP3_1;
	wire w_dff_B_8323vT4Z2_1;
	wire w_dff_B_Svcea6JQ3_1;
	wire w_dff_B_G0ca0ANb6_1;
	wire w_dff_B_sZsrwk6p7_1;
	wire w_dff_B_pvf6Qcwc9_1;
	wire w_dff_A_GsAj6t7L0_0;
	wire w_dff_A_hcjprUEn9_0;
	wire w_dff_A_2coFkNWB2_1;
	wire w_dff_A_tJaTjfpf6_1;
	wire w_dff_A_cF2zdSL49_1;
	wire w_dff_B_nm3ztWNx6_1;
	wire w_dff_B_ceVZ87HC7_1;
	wire w_dff_A_rrVAIVQh7_0;
	wire w_dff_A_YblE7OkE0_1;
	wire w_dff_B_R2RYqGny3_1;
	wire w_dff_B_MR7DW47J8_1;
	wire w_dff_B_e5rhHoLf7_1;
	wire w_dff_B_HBkPwT7n1_1;
	wire w_dff_B_IPQI8ROY3_1;
	wire w_dff_B_Zpb95vKL1_1;
	wire w_dff_B_8pBTZIfu7_1;
	wire w_dff_B_IiSgUiam6_1;
	wire w_dff_B_4pWTaMZ64_1;
	wire w_dff_B_SfhaCR7j1_1;
	wire w_dff_B_QzW38vyZ3_1;
	wire w_dff_B_2MEIc2nO8_1;
	wire w_dff_B_bCxMWUCL1_1;
	wire w_dff_B_wYoQnzWD0_1;
	wire w_dff_B_UUBNS6RN1_1;
	wire w_dff_B_yO9CgMGc9_1;
	wire w_dff_B_sRx4mkvJ4_1;
	wire w_dff_B_D9MUkGsy8_1;
	wire w_dff_B_ZoKDbdFU1_1;
	wire w_dff_B_m6Kw7pPu6_1;
	wire w_dff_B_8tMERvoy0_1;
	wire w_dff_B_qeSXmeGi5_1;
	wire w_dff_B_RuRPskcX9_1;
	wire w_dff_B_56tmRObt7_1;
	wire w_dff_B_3RbHRXTT8_1;
	wire w_dff_B_dOvBVwnH4_1;
	wire w_dff_A_MQ68W1B17_0;
	wire w_dff_A_xrfi6bE16_0;
	wire w_dff_A_2dkfefY57_0;
	wire w_dff_A_DGoOqOG40_0;
	wire w_dff_A_spCwRyVo0_0;
	wire w_dff_A_gPwATUp97_0;
	wire w_dff_A_nmgjS8Xb6_0;
	wire w_dff_A_9iMpH7lA9_0;
	wire w_dff_A_Jw1AnA3z8_0;
	wire w_dff_A_YBqRgmnk3_1;
	wire w_dff_A_uzrKeSt25_1;
	wire w_dff_A_8DU6gyBa5_1;
	wire w_dff_A_Kx58S53e5_1;
	wire w_dff_A_jayGZ5ID5_1;
	wire w_dff_A_l4lB1dYV0_1;
	wire w_dff_A_UqJoYVA22_1;
	wire w_dff_A_Cj6H1oYe1_1;
	wire w_dff_A_ahJjgRGn7_1;
	wire w_dff_A_ymixlnCm8_1;
	wire w_dff_A_LYRoVFOK4_1;
	wire w_dff_A_mE7r4Qpk6_1;
	wire w_dff_A_8PseJUOO5_2;
	wire w_dff_A_SObhG7m44_2;
	wire w_dff_A_q08o9JDc0_2;
	wire w_dff_A_gO0CZgDl3_2;
	wire w_dff_A_syD6FuEI1_2;
	wire w_dff_A_isFRQLDD7_2;
	wire w_dff_A_Q8g3bbiG9_2;
	wire w_dff_A_SITtjx9A9_2;
	wire w_dff_A_SEsZpSUG7_2;
	wire w_dff_A_uj6YHgjT6_2;
	wire w_dff_B_GqNr4VAu7_1;
	wire w_dff_B_QiPIzaLg1_1;
	wire w_dff_A_8GZwz2KJ3_0;
	wire w_dff_A_hhdMewAI5_1;
	wire w_dff_A_VIwWP3qT5_0;
	wire w_dff_A_sutCKZEx3_0;
	wire w_dff_A_hCg5HeLP7_0;
	wire w_dff_A_ksZD6eyg6_0;
	wire w_dff_A_6UTAXgVo7_0;
	wire w_dff_A_rhf35aYN2_0;
	wire w_dff_A_SngXMl4h8_1;
	wire w_dff_A_TzB2tQIO0_1;
	wire w_dff_A_zH3xNstB7_1;
	wire w_dff_A_HbGjGKGn8_1;
	wire w_dff_A_HcCFGtfx4_1;
	wire w_dff_A_1sdCHrTZ4_1;
	wire w_dff_A_Wp9ZOKuG8_1;
	wire w_dff_B_wXvHJvZE3_0;
	wire w_dff_B_AqoFKCle4_0;
	wire w_dff_B_TdCBwaQ41_0;
	wire w_dff_B_cNU4RuQC6_0;
	wire w_dff_B_tYY4Xa7D4_0;
	wire w_dff_B_YS5Rfacl9_0;
	wire w_dff_B_g8mgNMtr4_0;
	wire w_dff_B_6oMTsNTo3_0;
	wire w_dff_B_VaYnM2Jn2_0;
	wire w_dff_B_w9OQaKfF7_0;
	wire w_dff_B_Y1szM2d48_0;
	wire w_dff_B_EVacmhTY0_0;
	wire w_dff_B_FhzvEcCL1_0;
	wire w_dff_B_xE0Vmuox9_0;
	wire w_dff_B_2r4vXc0i3_0;
	wire w_dff_B_Bn9goyHr5_0;
	wire w_dff_B_hWRH1XRT5_0;
	wire w_dff_B_A70fKCp26_0;
	wire w_dff_B_riE1MaDo8_0;
	wire w_dff_B_RcXC3ijD4_0;
	wire w_dff_B_6HB1p32S0_2;
	wire w_dff_B_hdwEuQoB3_2;
	wire w_dff_B_9a14oI2n7_2;
	wire w_dff_B_YE3uA6j95_1;
	wire w_dff_B_3Yhumh1w7_1;
	wire w_dff_B_X693vMg99_1;
	wire w_dff_B_ooVjqmHx5_1;
	wire w_dff_B_T2m38Ivc1_1;
	wire w_dff_B_FHpWsZqr2_1;
	wire w_dff_B_OCoJLNfz7_1;
	wire w_dff_B_pfMAzIb94_1;
	wire w_dff_B_tduQ2zyU3_1;
	wire w_dff_B_QocHKizL4_1;
	wire w_dff_B_gP2r9NcX1_1;
	wire w_dff_B_IbWYYQrg5_1;
	wire w_dff_B_1vD3Cpe86_1;
	wire w_dff_B_gJCNnDqk5_1;
	wire w_dff_B_wYESkZk22_1;
	wire w_dff_B_MwEejZKs4_1;
	wire w_dff_B_DLl6XSoQ4_0;
	wire w_dff_B_goRQgdUe3_0;
	wire w_dff_B_PRlc2US79_0;
	wire w_dff_B_QBrcBN801_0;
	wire w_dff_B_G0YE7U8x1_0;
	wire w_dff_B_JAlnbApl7_0;
	wire w_dff_B_rBBPpyKu4_0;
	wire w_dff_B_XKiMiVu94_0;
	wire w_dff_B_OET0gN4x9_0;
	wire w_dff_B_Qe4Fzh8e1_0;
	wire w_dff_B_JtQRx7758_0;
	wire w_dff_B_uUfT9kX12_0;
	wire w_dff_A_iTx9WcG79_1;
	wire w_dff_A_mBnuKcvg5_1;
	wire w_dff_A_94ZwdcIq1_2;
	wire w_dff_A_naL09aep2_2;
	wire w_dff_B_uoWfeqFs0_0;
	wire w_dff_B_vcCWrcpf7_0;
	wire w_dff_A_CGCniSRM1_0;
	wire w_dff_A_3XKYABDM8_0;
	wire w_dff_A_CzTllBbM8_0;
	wire w_dff_A_BHwiBTuq5_0;
	wire w_dff_A_Mu4bqUEB1_0;
	wire w_dff_A_x1a6zmGF5_0;
	wire w_dff_A_Q3rVDNb76_0;
	wire w_dff_A_xx0NPEfj7_0;
	wire w_dff_A_DMJLjAWC3_0;
	wire w_dff_A_cJWklolw2_1;
	wire w_dff_A_F7ldFdBy6_1;
	wire w_dff_A_rKJw0v9g3_1;
	wire w_dff_A_pnV8RWif9_1;
	wire w_dff_A_6uXU1W2I7_0;
	wire w_dff_A_tLZXFnJW9_2;
	wire w_dff_A_xNE3xJgf3_2;
	wire w_dff_A_9nmSpktc8_2;
	wire w_dff_A_CKzamNTm1_2;
	wire w_dff_A_LcIwscl35_2;
	wire w_dff_A_QYuWKXTJ8_2;
	wire w_dff_A_A3LVXdBy9_2;
	wire w_dff_A_paLvKvVC2_2;
	wire w_dff_A_5dsmW2Lf1_2;
	wire w_dff_A_RGEdYACW1_2;
	wire w_dff_A_soXo7ihW1_2;
	wire w_dff_A_JIgpSfBy7_2;
	wire w_dff_A_wJQXwZ5L1_2;
	wire w_dff_A_9Sq3Quiw6_2;
	wire w_dff_A_aufjJL5v8_0;
	wire w_dff_A_nINmy0MP3_0;
	wire w_dff_A_tKb3P4l32_0;
	wire w_dff_A_XGBsZiXQ1_2;
	wire w_dff_A_ympCL9KT2_2;
	wire w_dff_A_0EfxXLcI0_0;
	wire w_dff_A_gz7mNcrP8_0;
	wire w_dff_A_EXz1UC2q5_0;
	wire w_dff_A_Wr3c9Y7C9_0;
	wire w_dff_A_Qlxb89eu8_0;
	wire w_dff_A_uuMJeVJz7_0;
	wire w_dff_A_DPtnB4aD3_0;
	wire w_dff_A_oOqJZCNw0_0;
	wire w_dff_A_1grDYaM51_0;
	wire w_dff_A_jAzl1Tul2_1;
	wire w_dff_A_DLqRDtDr1_1;
	wire w_dff_B_I8dQ9LZl8_3;
	wire w_dff_B_LPjgQV3R1_3;
	wire w_dff_B_qJKGc85C8_3;
	wire w_dff_B_TsyjQJph9_3;
	wire w_dff_B_XtQIU3YD6_3;
	wire w_dff_B_sejIwKca4_3;
	wire w_dff_B_sFIaZoQx5_3;
	wire w_dff_B_bIbi6GKC1_3;
	wire w_dff_B_TCpHyeD96_3;
	wire w_dff_B_cROi7K2p8_3;
	wire w_dff_B_hRGElnj35_3;
	wire w_dff_B_amyy1rbg2_1;
	wire w_dff_B_uImP2r9Y7_1;
	wire w_dff_B_QA83R6Zu0_1;
	wire w_dff_B_eNf6nigZ6_1;
	wire w_dff_B_gL4Z7yot5_1;
	wire w_dff_B_bI5pD3sw3_1;
	wire w_dff_B_CyLly1rx7_1;
	wire w_dff_B_CH6wZtSF9_1;
	wire w_dff_B_lH0bQREE9_1;
	wire w_dff_B_27bVFTkF2_1;
	wire w_dff_B_2YTQ9NR07_1;
	wire w_dff_B_lZULK1WQ3_1;
	wire w_dff_B_8KE7QGNS8_1;
	wire w_dff_B_ePxNtX9s6_1;
	wire w_dff_B_ztTiXgTH8_1;
	wire w_dff_B_B4WLClEx0_1;
	wire w_dff_B_bNSu0CbU2_1;
	wire w_dff_B_jwehbJPO4_1;
	wire w_dff_B_0Vs4H8rV0_1;
	wire w_dff_B_wqEGCKr88_1;
	wire w_dff_B_DicT3vzA4_1;
	wire w_dff_B_9saAF3tT4_1;
	wire w_dff_B_gxf9qsTh2_1;
	wire w_dff_B_p0a6wSf96_1;
	wire w_dff_B_LzIyNZfT0_1;
	wire w_dff_B_AtBHc7Nr5_1;
	wire w_dff_B_7wsLq0fn9_1;
	wire w_dff_B_CrdZCWz15_1;
	wire w_dff_B_zNX5cKln3_1;
	wire w_dff_B_RHDk62kT6_1;
	wire w_dff_B_FlKAU1g28_1;
	wire w_dff_B_c6eV3Lj95_1;
	wire w_dff_B_YZM3O3dE1_1;
	wire w_dff_B_fyb1ZnLl0_1;
	wire w_dff_B_rqQWsDeM4_1;
	wire w_dff_B_TsL2Ppb41_1;
	wire w_dff_B_5E2anqwI9_1;
	wire w_dff_B_cJ47nVtA4_1;
	wire w_dff_B_A4cRV65P7_1;
	wire w_dff_B_Q5gAEA4b4_1;
	wire w_dff_B_2GHUucvT0_0;
	wire w_dff_B_JWZuuTxj3_1;
	wire w_dff_B_SZmFmjq37_1;
	wire w_dff_A_xUQ57v087_1;
	wire w_dff_B_hH0ckDwQ5_3;
	wire w_dff_B_YNp8mRoG2_3;
	wire w_dff_B_WEAVzPa68_3;
	wire w_dff_B_Iqy5LW3W3_3;
	wire w_dff_B_w06pBtwL9_3;
	wire w_dff_A_4TUwTOi88_0;
	wire w_dff_A_TLEHEiKi1_1;
	wire w_dff_A_k4Mc6obz5_1;
	wire w_dff_B_cCmWeS6q0_3;
	wire w_dff_B_c3hkSaUW6_3;
	wire w_dff_B_uxCjVNF17_3;
	wire w_dff_B_r2cDyF8a9_3;
	wire w_dff_B_cCrJqu9M4_3;
	wire w_dff_B_3w3pEc0O3_3;
	wire w_dff_B_Fp8ErwLW8_3;
	wire w_dff_B_RNvt37Yl6_3;
	wire w_dff_B_214luyp62_3;
	wire w_dff_B_BrGB2khJ2_3;
	wire w_dff_B_VYdMdNZN7_3;
	wire w_dff_B_nd5VjrdD3_3;
	wire w_dff_B_1f30x1bG4_3;
	wire w_dff_B_jTDJ0t9Z3_3;
	wire w_dff_B_cfmT20Li7_3;
	wire w_dff_A_CUy5sQBD5_0;
	wire w_dff_A_nexf5sNW3_0;
	wire w_dff_A_eJepZW6A4_0;
	wire w_dff_A_uSho9M3r2_0;
	wire w_dff_A_G9DbjvMO8_0;
	wire w_dff_A_1EefmUZz0_0;
	wire w_dff_A_zMTya1Hp5_1;
	wire w_dff_A_MtmE4Kbw7_1;
	wire w_dff_A_BUWK75vh2_1;
	wire w_dff_A_zvXr6Mlm4_1;
	wire w_dff_A_elzg1mGC6_1;
	wire w_dff_A_ggjRFm5I5_1;
	wire w_dff_A_TrhiBh0t8_0;
	wire w_dff_A_YV7CwGLn4_0;
	wire w_dff_A_MpHDPtHA6_0;
	wire w_dff_A_nGAJWrGH3_0;
	wire w_dff_A_SgjoVAQz5_0;
	wire w_dff_A_reBStM3D9_0;
	wire w_dff_A_UuKmZWsm8_0;
	wire w_dff_A_Xln8IGVO3_0;
	wire w_dff_A_WCnGhDnX8_0;
	wire w_dff_A_4jhB6L743_0;
	wire w_dff_A_idRuKuo31_0;
	wire w_dff_A_HZuQsZKv6_0;
	wire w_dff_A_2BnHsd3a5_0;
	wire w_dff_A_ILvPx3Bw2_0;
	wire w_dff_A_r9II7cxP0_1;
	wire w_dff_A_ylr9DSxj3_1;
	wire w_dff_B_R6hTYZ170_1;
	wire w_dff_B_x0JyqcE81_1;
	wire w_dff_B_8AWjwpun6_0;
	wire w_dff_B_SyI5cbYT6_0;
	wire w_dff_B_HtJ1tkWA4_0;
	wire w_dff_B_mkrlpxlu3_0;
	wire w_dff_B_Rsl7u3pY8_0;
	wire w_dff_B_OsXF8n4H2_0;
	wire w_dff_B_WX07blrw5_0;
	wire w_dff_B_AGJ2n9JF5_0;
	wire w_dff_B_oIZfdQ3t3_0;
	wire w_dff_B_0owryR163_0;
	wire w_dff_B_IEV8kL8x3_0;
	wire w_dff_B_IBCxfeT16_0;
	wire w_dff_B_HWXJRv2U3_0;
	wire w_dff_B_91Hm7drc8_0;
	wire w_dff_B_dTxkmirP4_0;
	wire w_dff_B_9DTG6AAB9_0;
	wire w_dff_B_2nAI3GlU6_0;
	wire w_dff_B_Vik9IfoL0_1;
	wire w_dff_B_VuECQi0n9_1;
	wire w_dff_B_dichDG2I4_1;
	wire w_dff_B_1p4irCzB1_0;
	wire w_dff_B_81zL4H8Z9_0;
	wire w_dff_B_kPiXskZA6_0;
	wire w_dff_B_QmSMmMpn5_0;
	wire w_dff_B_iw81HcQw0_0;
	wire w_dff_B_04dMJrY67_0;
	wire w_dff_B_ft4cY8BK5_0;
	wire w_dff_B_Ul80cRAF5_0;
	wire w_dff_B_HVbh6isF9_0;
	wire w_dff_B_VrASsSzX3_0;
	wire w_dff_B_tFw8L8ZE6_0;
	wire w_dff_B_OwOVWKcW5_0;
	wire w_dff_B_LNrbF8xU3_0;
	wire w_dff_B_n8iNjRAv9_0;
	wire w_dff_B_af7GzYc13_0;
	wire w_dff_B_eAEItApn7_0;
	wire w_dff_B_VLqBh0GW4_0;
	wire w_dff_B_YmPSEMOH6_1;
	wire w_dff_B_I52hihRt6_1;
	wire w_dff_B_2TsCaoR02_1;
	wire w_dff_A_8ObYxFQD0_0;
	wire w_dff_A_hoerIxgT4_0;
	wire w_dff_A_szTvRgYt2_0;
	wire w_dff_A_VendsrEd8_0;
	wire w_dff_A_ifR6nME50_0;
	wire w_dff_A_3CygBpVO8_1;
	wire w_dff_A_4NLguyDh3_1;
	wire w_dff_A_6lPGGltN3_1;
	wire w_dff_A_RhMIT62F1_1;
	wire w_dff_A_1J9UpE711_0;
	wire w_dff_A_QQJsqeN94_0;
	wire w_dff_A_MEQeOdlP0_0;
	wire w_dff_A_S4xEADRG4_0;
	wire w_dff_A_wMAhAGCw2_0;
	wire w_dff_A_xHRW5i751_1;
	wire w_dff_A_67FO2KtR2_1;
	wire w_dff_A_ueoFOx6y3_1;
	wire w_dff_A_ggGHQquF5_1;
	wire w_dff_A_cqBgmFZs1_0;
	wire w_dff_A_IMPRyMYe5_0;
	wire w_dff_A_UPfevPH08_0;
	wire w_dff_B_5e5zuS1a7_1;
	wire w_dff_B_cScKjOlA1_1;
	wire w_dff_B_Soo3aZbp8_1;
	wire w_dff_B_4kkelaZl7_1;
	wire w_dff_B_0CCn8k5K2_1;
	wire w_dff_B_6iKiU5vD1_1;
	wire w_dff_B_WyjygRrj8_1;
	wire w_dff_B_tmKQDly99_1;
	wire w_dff_B_B3u4WQN31_1;
	wire w_dff_B_0LXL32Ip2_1;
	wire w_dff_B_vi5kGt7H4_1;
	wire w_dff_B_srHVl0kn2_1;
	wire w_dff_B_fXDtazfX6_1;
	wire w_dff_B_cZm5gRNQ2_1;
	wire w_dff_B_CLiXq3ns6_1;
	wire w_dff_B_YfWEKviO1_1;
	wire w_dff_B_96Eip8xL8_1;
	wire w_dff_B_CxmjMu431_1;
	wire w_dff_B_P19xN8GO2_1;
	wire w_dff_B_RXiEFzrS9_1;
	wire w_dff_B_d7NXM7kH9_1;
	wire w_dff_B_l62URcUl6_1;
	wire w_dff_B_UuyVYPP90_1;
	wire w_dff_A_mKMkx3402_1;
	wire w_dff_A_shThLQD70_1;
	wire w_dff_A_w0BWLKlM7_1;
	wire w_dff_A_JK4DdP7w1_1;
	wire w_dff_A_3sjU6kPM0_1;
	wire w_dff_A_W06crO5J0_1;
	wire w_dff_A_aLNzTqI70_1;
	wire w_dff_A_T4z7Q8dh8_1;
	wire w_dff_A_WhiZjXB04_1;
	wire w_dff_A_S3qR5mKt8_1;
	wire w_dff_A_epKmczTI7_1;
	wire w_dff_A_BiVyAeaj8_1;
	wire w_dff_A_7AQuVPSb0_1;
	wire w_dff_A_uDMLZepB0_1;
	wire w_dff_A_2CAjTrrz1_2;
	wire w_dff_A_0jKcvtdD7_2;
	wire w_dff_A_6DLwqrha8_2;
	wire w_dff_A_cOUpg74E0_2;
	wire w_dff_A_hOCVYeko9_2;
	wire w_dff_A_FH4lGZ0e5_2;
	wire w_dff_A_q5y470NY4_2;
	wire w_dff_A_LSux8jAS9_2;
	wire w_dff_A_jk8k9AAV0_2;
	wire w_dff_A_BpvSD57Q4_2;
	wire w_dff_A_QaUtT28p8_1;
	wire w_dff_A_Cy1pQyLf6_1;
	wire w_dff_A_TQXjjSzL8_1;
	wire w_dff_A_WvDWmAAi1_1;
	wire w_dff_A_rKWZdJN14_1;
	wire w_dff_A_Nj8pWmv18_1;
	wire w_dff_A_el3opAui4_1;
	wire w_dff_A_PpPYDotE0_1;
	wire w_dff_A_KzQ1iZc55_1;
	wire w_dff_A_HbuwozZH6_1;
	wire w_dff_A_ZWMvM8Jk9_1;
	wire w_dff_A_72A47Qsx6_2;
	wire w_dff_A_cgRPNDmG7_2;
	wire w_dff_A_nqtTNS5b0_2;
	wire w_dff_A_S6rN69Ok5_2;
	wire w_dff_B_RepmlAMK5_3;
	wire w_dff_B_LWef8ZPO9_3;
	wire w_dff_B_rHb0Nf8Z9_3;
	wire w_dff_B_4rLMCRM48_3;
	wire w_dff_B_VnJsDzlZ0_3;
	wire w_dff_B_aeUcAszg5_3;
	wire w_dff_B_hjkqYJ0R5_3;
	wire w_dff_B_3fKYXCof6_3;
	wire w_dff_B_MwUyoqxu1_3;
	wire w_dff_A_s4mXJW8X6_0;
	wire w_dff_A_sg5nOhNJ8_1;
	wire w_dff_B_0OfVjyn06_1;
	wire w_dff_B_CZWc9HjP5_1;
	wire w_dff_A_C4fwjque9_0;
	wire w_dff_A_VtD9dtYE9_0;
	wire w_dff_A_Eo7AXJou5_0;
	wire w_dff_A_20lzqXXE1_0;
	wire w_dff_A_Rq61JYAI3_0;
	wire w_dff_A_Dpy9uMNc4_0;
	wire w_dff_A_V3Ovmbnu8_0;
	wire w_dff_A_t9JhJckN9_0;
	wire w_dff_A_9E4B0bnc0_0;
	wire w_dff_A_rQSOU49D5_0;
	wire w_dff_A_iCDC3FKU1_0;
	wire w_dff_A_hLzxzN376_0;
	wire w_dff_A_yDxUt3ZB4_0;
	wire w_dff_A_Ts7n3fiN4_0;
	wire w_dff_A_HRzarivN0_0;
	wire w_dff_A_I3ctsL385_0;
	wire w_dff_A_l32uxYpM6_0;
	wire w_dff_A_tbePrfwj9_0;
	wire w_dff_A_thC3xxEd2_0;
	wire w_dff_A_sX5Gxn2m6_0;
	wire w_dff_A_93XKIR4Z5_0;
	wire w_dff_A_qnlRfEJH3_0;
	wire w_dff_A_mExzMo0u8_1;
	wire w_dff_A_R1hUE9gF9_1;
	wire w_dff_A_ahiXVkYi4_1;
	wire w_dff_A_zH1Fmsaq0_1;
	wire w_dff_A_BP8l9MQe5_1;
	wire w_dff_A_geeYu1rM2_1;
	wire w_dff_A_1Kyrp0C55_1;
	wire w_dff_A_UUM8XIWb2_1;
	wire w_dff_A_rup8d4tL5_1;
	wire w_dff_A_cOZVQ2Qy5_1;
	wire w_dff_A_jiFySq680_1;
	wire w_dff_A_5ViwmFPS6_2;
	wire w_dff_A_z4gXNJDl6_1;
	wire w_dff_A_RCIjzLbv0_2;
	wire w_dff_A_pVl6RSdy0_0;
	wire w_dff_A_lG0fvDEl3_0;
	wire w_dff_A_pPnwH4os3_0;
	wire w_dff_A_UeNZaFw28_0;
	wire w_dff_A_yXrFLySN0_0;
	wire w_dff_A_m7aGkCFq7_0;
	wire w_dff_A_ektHuPxZ0_0;
	wire w_dff_A_ePg6tEvb3_0;
	wire w_dff_A_bYiS5xFi0_0;
	wire w_dff_A_OKbZz6mn5_0;
	wire w_dff_A_yMRX3B4B8_0;
	wire w_dff_A_xs7os9hb7_0;
	wire w_dff_A_dxsp55vT7_0;
	wire w_dff_A_zVzCJJkn9_0;
	wire w_dff_A_rPnQuvwW4_0;
	wire w_dff_A_AoVGNFxa4_0;
	wire w_dff_A_l5P2P98g9_0;
	wire w_dff_A_AzbpNtx49_0;
	wire w_dff_A_RYEMwVuI5_0;
	wire w_dff_A_cQSBFBQn1_0;
	wire w_dff_A_kKjm6x1T3_0;
	wire w_dff_A_rvtdpdSA9_0;
	wire w_dff_A_a1YkzlzF7_0;
	wire w_dff_B_HgJ8UPjT6_1;
	wire w_dff_B_YWLnt9UX1_1;
	wire w_dff_B_MPOY0pX70_1;
	wire w_dff_B_a62O9a6C9_1;
	wire w_dff_B_ZWfbfxKp9_1;
	wire w_dff_B_x72qEU6c5_1;
	wire w_dff_B_4TdQoK0d6_1;
	wire w_dff_B_VckQEQ0L1_1;
	wire w_dff_B_Wm1Zug195_1;
	wire w_dff_B_XN2ZOdsd8_1;
	wire w_dff_B_MiBFHln91_1;
	wire w_dff_B_SeNIhFYC4_1;
	wire w_dff_B_wbKTMj9v2_1;
	wire w_dff_B_mtPs3ggg7_1;
	wire w_dff_B_r5Hnzn2T6_1;
	wire w_dff_B_OBjHK4ED8_1;
	wire w_dff_B_7e4hA8VI6_1;
	wire w_dff_B_ABBur8aH1_1;
	wire w_dff_B_1aanQgeF5_1;
	wire w_dff_B_1zhas1ym0_1;
	wire w_dff_B_3yr8icmq5_1;
	wire w_dff_B_nzzW5EV01_1;
	wire w_dff_B_kT1rIe232_1;
	wire w_dff_A_4jVOEVBg2_1;
	wire w_dff_A_3Espyj9e2_1;
	wire w_dff_A_PjoTc44T1_1;
	wire w_dff_A_Pg61oTH26_1;
	wire w_dff_A_Cjwjtw2x4_1;
	wire w_dff_A_YGWF4hHO2_1;
	wire w_dff_A_bs99USbQ0_1;
	wire w_dff_A_staoFMI34_1;
	wire w_dff_A_dQmaPLvb6_1;
	wire w_dff_A_RCCUsXbQ6_1;
	wire w_dff_A_gWCrgGVr6_1;
	wire w_dff_A_4eNIcdzN6_1;
	wire w_dff_A_UdhofHLe6_1;
	wire w_dff_A_tYiNUfGA0_1;
	wire w_dff_A_vsaFAMqD6_2;
	wire w_dff_A_cPi1KRNX2_2;
	wire w_dff_A_Q2kYCTVY1_2;
	wire w_dff_A_NVDIreXF1_2;
	wire w_dff_A_e1ygDbgS2_2;
	wire w_dff_A_1wbVN6Ao6_2;
	wire w_dff_A_Qr4wcDax7_2;
	wire w_dff_A_otfdHdpE7_2;
	wire w_dff_A_WSJtnANh8_2;
	wire w_dff_A_jY9b8IVo4_2;
	wire w_dff_A_EpsawGem2_1;
	wire w_dff_A_yUKHhQlm8_1;
	wire w_dff_A_4qoWoKgS0_1;
	wire w_dff_A_1BgLTNUL3_1;
	wire w_dff_A_gQJlXu2F1_1;
	wire w_dff_A_hHTfZ0Hv9_1;
	wire w_dff_A_Kuwqft7N9_1;
	wire w_dff_A_0KwAEId78_1;
	wire w_dff_A_CWkbWoNy0_1;
	wire w_dff_A_DQyYBON80_1;
	wire w_dff_A_Jnct4fnW9_1;
	wire w_dff_A_xMfdpUh61_2;
	wire w_dff_A_eTq7qqbM5_2;
	wire w_dff_A_5whRubta6_2;
	wire w_dff_A_xl7ytOp19_2;
	wire w_dff_A_yKkjTM6S1_2;
	wire w_dff_B_EDGMNkaZ3_3;
	wire w_dff_B_XYvyIm6Z7_3;
	wire w_dff_B_5H2dPdpX3_3;
	wire w_dff_B_NagbFXfR8_3;
	wire w_dff_B_EiMOcFUM2_3;
	wire w_dff_B_SszUKQ7U8_3;
	wire w_dff_B_OOGxSDZl3_3;
	wire w_dff_B_ewRcziBi2_3;
	wire w_dff_B_d5G7vJYJ1_3;
	wire w_dff_A_ZKP47iAl5_0;
	wire w_dff_A_yU2mtP1v8_0;
	wire w_dff_A_wsrgcQzq2_1;
	wire w_dff_B_8HhfATdu6_1;
	wire w_dff_B_X3poD1NW2_1;
	wire w_dff_A_nnritehd3_0;
	wire w_dff_A_bFJAuPFw7_0;
	wire w_dff_A_cSVcj86P3_0;
	wire w_dff_A_ES1gNpws5_0;
	wire w_dff_A_uZ2MuqYv7_0;
	wire w_dff_A_SsgtXLWW5_0;
	wire w_dff_A_nRZzmmkZ5_0;
	wire w_dff_A_zPJl7H4M7_0;
	wire w_dff_A_mFBio6Xq5_0;
	wire w_dff_A_CMvuMxIf6_0;
	wire w_dff_A_r6ROu1PE9_0;
	wire w_dff_A_cKfaf0gZ1_0;
	wire w_dff_A_JwPA8TKO3_0;
	wire w_dff_A_xbm5mn4H7_0;
	wire w_dff_A_QvaSjINX6_0;
	wire w_dff_A_iWzEyBod0_0;
	wire w_dff_A_WMgA96Mm9_0;
	wire w_dff_A_OMsHxYZy4_0;
	wire w_dff_A_nOhZi9TO3_0;
	wire w_dff_A_Fodnh04C3_0;
	wire w_dff_A_ho5eJw8Q2_0;
	wire w_dff_A_ViaIf9gQ0_0;
	wire w_dff_A_49fwpllY0_1;
	wire w_dff_A_RyKlHmmw9_1;
	wire w_dff_A_fPv4t5mR7_1;
	wire w_dff_A_2udNlhav7_1;
	wire w_dff_A_xRSxyns32_1;
	wire w_dff_A_AXj1pz1W1_1;
	wire w_dff_A_5UMxVzrt3_1;
	wire w_dff_A_U6VoDHgm8_1;
	wire w_dff_A_U89a4rlK1_1;
	wire w_dff_B_usrkDEF45_2;
	wire w_dff_A_78NHFyP55_1;
	wire w_dff_A_UJNqLQE41_1;
	wire w_dff_A_8bKgs9nA1_2;
	wire w_dff_A_REUvvtvf3_1;
	wire w_dff_A_W5GRnw7Q9_2;
	wire w_dff_A_kYAyl4Es8_0;
	wire w_dff_A_xbX0qH2H3_0;
	wire w_dff_A_cFnGhN872_0;
	wire w_dff_A_iuIvA3rV3_0;
	wire w_dff_A_pqW3gnFS2_0;
	wire w_dff_A_TkTNPPh29_0;
	wire w_dff_A_XiUTjsH41_0;
	wire w_dff_A_gtbTygPp0_0;
	wire w_dff_A_gooogi1N5_0;
	wire w_dff_A_HBRPOocA4_0;
	wire w_dff_A_aCFXkw709_0;
	wire w_dff_A_ANDoUeuS0_0;
	wire w_dff_A_wekDcAyI7_0;
	wire w_dff_A_CTImzvee0_0;
	wire w_dff_A_Y9dxx01h4_0;
	wire w_dff_A_k1YFpIgV5_0;
	wire w_dff_A_OZ1jnFH57_0;
	wire w_dff_A_TGrAQ5lS2_0;
	wire w_dff_A_KiiWh2s00_0;
	wire w_dff_A_ENa69U1Q8_0;
	wire w_dff_A_63eRILzb9_0;
	wire w_dff_A_unOqZuzV5_0;
	wire w_dff_A_RKaJPw4R7_0;
	wire w_dff_B_V5IEzLUR7_1;
	wire w_dff_B_mPCpRXV06_1;
	wire w_dff_B_e5LCxlWi4_1;
	wire w_dff_B_zFn0wqg06_1;
	wire w_dff_B_qkSi2MYM9_1;
	wire w_dff_B_RFCJQDYN4_1;
	wire w_dff_B_aGSDuVwD1_1;
	wire w_dff_B_44izKsrk1_1;
	wire w_dff_B_E547pxtW2_1;
	wire w_dff_B_uiHgqJJs2_1;
	wire w_dff_B_tR5xXrwi6_1;
	wire w_dff_B_YeaBm7T12_1;
	wire w_dff_B_U7y8yZsP7_1;
	wire w_dff_B_tgNOku393_1;
	wire w_dff_B_QF3v6Wca2_1;
	wire w_dff_B_DdqiYxiA1_1;
	wire w_dff_B_HyoYCgQw7_1;
	wire w_dff_B_gshcjvz24_1;
	wire w_dff_B_xZjGJMqp0_1;
	wire w_dff_B_KDpoq9PG1_1;
	wire w_dff_B_KhEpIVJg3_1;
	wire w_dff_B_OfLo8Dwn5_1;
	wire w_dff_B_avnGWs4K3_1;
	wire w_dff_B_fI9Ko6vw1_1;
	wire w_dff_B_cGurmsCa7_1;
	wire w_dff_B_RNWimfls4_1;
	wire w_dff_B_0v12PZQq4_1;
	wire w_dff_B_ahKwhzbV6_1;
	wire w_dff_B_1CJMlBrW8_1;
	wire w_dff_B_MUvRWufT2_1;
	wire w_dff_B_mB18wU551_1;
	wire w_dff_B_BzJcBxKf6_1;
	wire w_dff_B_Rgw8ftP25_1;
	wire w_dff_B_6C5fKtuJ2_1;
	wire w_dff_B_TunFiVrq0_1;
	wire w_dff_B_dx4Mnm3x1_1;
	wire w_dff_B_n6thTjlm9_1;
	wire w_dff_B_7HXIOS9H0_1;
	wire w_dff_B_CFtJtP666_1;
	wire w_dff_B_MzpXaZU74_1;
	wire w_dff_B_2kJT5lgh8_1;
	wire w_dff_B_pxF6YiMo0_1;
	wire w_dff_B_j3YVEVL78_1;
	wire w_dff_B_CohgHBSY3_1;
	wire w_dff_B_wFekHFN83_1;
	wire w_dff_A_rVNUCMms5_0;
	wire w_dff_A_xttwV3ie8_0;
	wire w_dff_A_qSmVgy6h2_0;
	wire w_dff_A_f7GXBkXS7_0;
	wire w_dff_A_WmN2Cb3x5_0;
	wire w_dff_A_L4LmGRfS0_0;
	wire w_dff_A_hCZfusYl8_0;
	wire w_dff_A_UKfEVYh58_0;
	wire w_dff_A_iL6KFSsh0_0;
	wire w_dff_A_y2aSF4gJ6_0;
	wire w_dff_A_oK217UZV7_0;
	wire w_dff_A_mdEpUr4E1_0;
	wire w_dff_A_9Drrbq1Y8_0;
	wire w_dff_A_erbST0ow0_0;
	wire w_dff_A_qSpU3F0Z5_0;
	wire w_dff_A_5dPsLluu0_1;
	wire w_dff_A_bFvlcNX67_1;
	wire w_dff_A_T4R624mE2_1;
	wire w_dff_A_qFgXLMG63_1;
	wire w_dff_A_nm154Df46_1;
	wire w_dff_A_t7pXmoyr7_1;
	wire w_dff_A_n0TdrATN1_1;
	wire w_dff_A_mSYTnBfQ8_1;
	wire w_dff_A_7crUjiHr3_1;
	wire w_dff_A_NkslOwSe4_1;
	wire w_dff_A_u3Z345Or9_1;
	wire w_dff_A_TtrAxRY82_1;
	wire w_dff_A_txC9NkcK5_1;
	wire w_dff_A_XIzIFGDj1_1;
	wire w_dff_A_LSaItoaT7_1;
	wire w_dff_A_LkqS6dEE0_1;
	wire w_dff_A_ki2Ah21m4_1;
	wire w_dff_A_PAzOq7zy7_1;
	wire w_dff_A_zgxJgVYg7_1;
	wire w_dff_A_JWPUOYga0_1;
	wire w_dff_A_erRBw8ZA6_1;
	wire w_dff_A_H3IAuWaq0_1;
	wire w_dff_A_ujSvXf4I7_1;
	wire w_dff_A_QLQYgiUC5_1;
	wire w_dff_A_XdriLG8E9_1;
	wire w_dff_A_zLwyubXZ7_1;
	wire w_dff_A_RmDAx6AT3_1;
	wire w_dff_A_ly60JqnN4_1;
	wire w_dff_A_p5lmxcXw0_1;
	wire w_dff_A_82lobM707_1;
	wire w_dff_A_xn1HbwAj0_1;
	wire w_dff_A_bnPiJUJk7_2;
	wire w_dff_A_kDyCWJqk4_2;
	wire w_dff_A_vd3u4Ewu0_2;
	wire w_dff_A_MZ8MXjhX5_2;
	wire w_dff_A_1FKVDn6M2_2;
	wire w_dff_A_zyDbunfF3_2;
	wire w_dff_A_NGDH3qGO0_2;
	wire w_dff_A_ByRyP1HW5_2;
	wire w_dff_A_fzrE1owu5_2;
	wire w_dff_A_29yt73si3_2;
	wire w_dff_A_D2E6zgTh5_2;
	wire w_dff_A_oynphTOB3_2;
	wire w_dff_A_Rc4Jnk2v7_2;
	wire w_dff_A_PAIISbnq6_2;
	wire w_dff_A_YlBmGZHh2_2;
	wire w_dff_A_kXSJXCrt9_2;
	wire w_dff_A_22DRyuHC2_2;
	wire w_dff_A_yffEAbKz6_2;
	wire w_dff_A_8OLMbiwS5_2;
	wire w_dff_A_iBDS9ARQ2_2;
	wire w_dff_A_vCyZFVoO5_1;
	wire w_dff_A_nETcOfKL1_1;
	wire w_dff_A_ENashX1U6_1;
	wire w_dff_A_8ls4io8I3_1;
	wire w_dff_A_mq01duzk5_1;
	wire w_dff_A_0XkUD5EV1_1;
	wire w_dff_A_lwhZMMEm0_1;
	wire w_dff_A_WnNnlVG17_1;
	wire w_dff_A_KhjNfNI49_1;
	wire w_dff_A_H3VbJS9q1_1;
	wire w_dff_A_Awc6SkHf0_1;
	wire w_dff_A_nOo7LMw46_1;
	wire w_dff_A_nJijrz1b1_1;
	wire w_dff_A_PfiBgvRn6_1;
	wire w_dff_A_N2jZG2ad6_1;
	wire w_dff_A_crpsK3c79_1;
	wire w_dff_A_lw8G4GUT8_1;
	wire w_dff_A_NMehygOp9_1;
	wire w_dff_A_LgrVplrC2_2;
	wire w_dff_A_3gMgaEEW0_2;
	wire w_dff_A_y80IbRP17_2;
	wire w_dff_A_diOxwtbg9_2;
	wire w_dff_A_qqOvGl9I9_2;
	wire w_dff_A_T73MkNtP6_2;
	wire w_dff_A_aHvX8tWT8_2;
	wire w_dff_A_IZ0J4Get0_2;
	wire w_dff_A_9rRmXcKe0_2;
	wire w_dff_A_ADELT7Vs8_2;
	wire w_dff_A_olEYvere9_2;
	wire w_dff_A_c6VJc8HF5_1;
	wire w_dff_A_s0Hg9CDf6_1;
	wire w_dff_A_b7N5FImU1_1;
	wire w_dff_A_RpfOhTvr0_1;
	wire w_dff_A_UzgRR4S39_1;
	wire w_dff_A_v8lotj2U9_1;
	wire w_dff_A_n4rH0UBr1_1;
	wire w_dff_A_CrecUhpv0_1;
	wire w_dff_A_jmVhB9PT8_1;
	wire w_dff_A_LeyYPWqk5_1;
	wire w_dff_A_nqwXVtt81_1;
	wire w_dff_A_T4CLY8gb3_1;
	wire w_dff_A_CF1l3lga2_1;
	wire w_dff_A_pOBdfCEK3_1;
	wire w_dff_A_VCaThd1q3_1;
	wire w_dff_A_j2p6vO1V5_1;
	wire w_dff_A_H1aFAhHN5_1;
	wire w_dff_A_OkzwuYIS6_1;
	wire w_dff_A_Sgz9I38z2_1;
	wire w_dff_A_ngBRyqUN4_1;
	wire w_dff_A_4kfIcUqA6_1;
	wire w_dff_A_XLlFqoxv0_1;
	wire w_dff_A_jEYaMwoB4_1;
	wire w_dff_A_XlP6CFhZ0_1;
	wire w_dff_A_rNuAEmgB4_0;
	wire w_dff_A_bb7qMjrM9_0;
	wire w_dff_A_ygWYn2bj3_0;
	wire w_dff_A_d99eG6Th8_0;
	wire w_dff_A_aHLTcKNW6_0;
	wire w_dff_A_FvzwZuTH2_0;
	wire w_dff_A_WSVK0JUb1_0;
	wire w_dff_A_mbmiZXFa9_0;
	wire w_dff_A_b7Fpg7u54_0;
	wire w_dff_A_xKwHvcxb9_2;
	wire w_dff_A_Ls7O1bV69_2;
	wire w_dff_A_Z57ELrXu0_2;
	wire w_dff_A_l69HWdEl6_2;
	wire w_dff_A_shQhlWKM6_2;
	wire w_dff_A_5WLz3xtU3_2;
	wire w_dff_A_DBsOnch54_2;
	wire w_dff_A_mhquwqu78_2;
	wire w_dff_A_Y7xX38H71_2;
	wire w_dff_A_Xpbvfbj07_2;
	wire w_dff_A_LGSoJkVR4_2;
	wire w_dff_A_lFyJjsoJ0_2;
	wire w_dff_A_4W665TrL5_2;
	wire w_dff_A_vj2p8AEF5_2;
	wire w_dff_A_yvttYkk23_2;
	wire w_dff_A_6FdwXwMG7_2;
	wire w_dff_A_VkLc473u6_2;
	wire w_dff_A_4DUptWGz8_2;
	wire w_dff_A_xWT9hROC2_2;
	wire w_dff_A_UXWckWh10_2;
	wire w_dff_A_EV9tojrg9_2;
	wire w_dff_A_Kyriajg40_2;
	wire w_dff_A_yBqaRBxN0_1;
	wire w_dff_A_neSukdh07_1;
	wire w_dff_A_cJPdEet27_1;
	wire w_dff_A_ZQiGzv119_1;
	wire w_dff_A_crFJutxU7_1;
	wire w_dff_A_KKTRLcsr4_1;
	wire w_dff_A_wQQQCS093_1;
	wire w_dff_A_VmCq3Nf10_1;
	wire w_dff_A_g2h8skqp7_1;
	wire w_dff_A_IKmsPhYd5_1;
	wire w_dff_A_ubDseIHZ2_1;
	wire w_dff_A_YMi0R8rh5_1;
	wire w_dff_A_3nbfTjjo9_1;
	wire w_dff_A_wZuxnlWM7_1;
	wire w_dff_A_ZP6roR749_1;
	wire w_dff_A_HAouYHwE8_1;
	wire w_dff_A_ukfZl4yL8_1;
	wire w_dff_A_UarNc1l53_1;
	wire w_dff_A_v8UhOTPX0_1;
	wire w_dff_A_Nfc79ZMy5_2;
	wire w_dff_A_rvxLGAmG0_2;
	wire w_dff_A_vxQ2Vjw62_2;
	wire w_dff_A_aUrD6viN8_2;
	wire w_dff_A_9mzZP8q07_2;
	wire w_dff_A_5ozHnspx2_2;
	wire w_dff_A_pKXmSvw00_2;
	wire w_dff_A_S8Er80wL7_2;
	wire w_dff_A_DfSkNTJ80_2;
	wire w_dff_A_i6ApMTD60_2;
	wire w_dff_A_ot76YAmh8_2;
	wire w_dff_A_OyAR79sj4_2;
	wire w_dff_A_Xl6d13p94_2;
	wire w_dff_B_1kjSiEjw6_1;
	wire w_dff_B_0dlhkWcu6_1;
	wire w_dff_B_sunLTnWp9_1;
	wire w_dff_B_HHLt3znN7_1;
	wire w_dff_B_m77swa604_1;
	wire w_dff_B_9Y2rnsm06_1;
	wire w_dff_B_1RUThDct8_1;
	wire w_dff_B_jQatCG0n3_1;
	wire w_dff_B_7yHdn2Wc5_1;
	wire w_dff_B_NAohWdCa3_1;
	wire w_dff_B_HFvGyynk1_1;
	wire w_dff_B_81XKjS4J8_1;
	wire w_dff_B_uX0eNeH98_1;
	wire w_dff_B_ISoAeJD93_1;
	wire w_dff_B_sq8zqZoM7_1;
	wire w_dff_B_EblJsutN7_1;
	wire w_dff_B_GNHqy0OS0_1;
	wire w_dff_B_cHINSXlL4_1;
	wire w_dff_B_zEouXW107_1;
	wire w_dff_B_MC1CqQ0i9_1;
	wire w_dff_B_B2lM3Cwn0_1;
	wire w_dff_B_MWG9IqOL0_1;
	wire w_dff_B_C1gAIC6b5_1;
	wire w_dff_B_lK20VBSx8_1;
	wire w_dff_B_FLJHjwzx7_1;
	wire w_dff_B_rAdYT9FP7_1;
	wire w_dff_B_XRL9M5rQ4_1;
	wire w_dff_B_W2o8yhyI6_1;
	wire w_dff_B_TKjQU7uI1_1;
	wire w_dff_B_lE0OROBT1_1;
	wire w_dff_B_rVryp8kL2_1;
	wire w_dff_B_qXwJEIyb8_1;
	wire w_dff_B_obY4200g6_1;
	wire w_dff_B_u3VZ3E730_1;
	wire w_dff_B_UtmfcqAP0_1;
	wire w_dff_B_sJ4WLeyM0_1;
	wire w_dff_B_vPzjLQUq4_1;
	wire w_dff_B_ah0BjhyB9_1;
	wire w_dff_B_2TT76pLZ6_1;
	wire w_dff_B_YGxHVztd0_1;
	wire w_dff_B_7ZZJBXGH0_1;
	wire w_dff_B_ACDNcCPF8_1;
	wire w_dff_B_UFxbdRmG4_1;
	wire w_dff_B_GxSbALLt5_1;
	wire w_dff_B_b5XNq4Yj5_1;
	wire w_dff_B_wyGLOH1w5_0;
	wire w_dff_B_8xfjtWrt5_0;
	wire w_dff_B_18zmQWva2_0;
	wire w_dff_B_WMl50vtD4_0;
	wire w_dff_B_GePLgr399_0;
	wire w_dff_B_kC4npNCu9_0;
	wire w_dff_B_fX8Rrdkf8_0;
	wire w_dff_B_qWhNQUeJ7_0;
	wire w_dff_B_lRtGoqTU6_0;
	wire w_dff_B_79PgY89o7_0;
	wire w_dff_B_JXT4TP7N7_0;
	wire w_dff_B_1PXEBAQ64_0;
	wire w_dff_B_fiyiR4TN4_0;
	wire w_dff_B_Q69xA2qk9_0;
	wire w_dff_B_vcIYmIXm5_0;
	wire w_dff_B_NffOVg0X4_0;
	wire w_dff_B_WzZjOkoB0_0;
	wire w_dff_B_qJ6ZC2TC2_0;
	wire w_dff_B_RNrhA1g56_0;
	wire w_dff_B_YC3cl44O4_0;
	wire w_dff_B_6OMTBjEN4_0;
	wire w_dff_B_J3xMFMzu4_0;
	wire w_dff_B_9OHPeFdG6_0;
	wire w_dff_B_lw0hFDoO1_0;
	wire w_dff_B_5nvaracM7_0;
	wire w_dff_B_eHmpSaiz7_0;
	wire w_dff_B_ASVe7ABE1_0;
	wire w_dff_B_uBoKKbTs1_0;
	wire w_dff_B_qR3rCMT00_1;
	wire w_dff_B_pBSK8JsB7_1;
	wire w_dff_B_6UrklJ322_1;
	wire w_dff_A_NuoaZjgQ1_0;
	wire w_dff_B_txQzqDiA3_1;
	wire w_dff_B_8q75BwXS0_1;
	wire w_dff_A_0YSAPy1G7_1;
	wire w_dff_B_YFQvHGfJ1_0;
	wire w_dff_A_p0Cf2Y2O2_0;
	wire w_dff_B_0IfXNE3G0_1;
	wire w_dff_A_DA9kbywb7_0;
	wire w_dff_B_y3kByK1p7_2;
	wire w_dff_A_f0ymMM9S3_0;
	wire w_dff_A_OmWq2bZc5_0;
	wire w_dff_A_TVETGGw30_0;
	wire w_dff_B_1sRfBGLA1_1;
	wire w_dff_B_9RVLNSpN3_1;
	wire w_dff_B_SbN4iOHA4_1;
	wire w_dff_A_m2qxj6TM4_1;
	wire w_dff_B_WoUeSEXS3_1;
	wire w_dff_B_qaJGMqE42_1;
	wire w_dff_A_eRUhx5PH6_1;
	wire w_dff_B_Z90rQbll4_1;
	wire w_dff_A_MS4Ctbw94_0;
	wire w_dff_A_wgdFmCoQ5_0;
	wire w_dff_A_QST1B0gp0_0;
	wire w_dff_A_ADhn6bIm6_1;
	wire w_dff_A_SEGSm8Ks1_1;
	wire w_dff_A_nvpZD04T0_1;
	wire w_dff_A_qGz84Lul3_1;
	wire w_dff_A_lB6CdXag1_1;
	wire w_dff_A_yiuihqQH1_1;
	wire w_dff_A_1nueY5bw9_1;
	wire w_dff_A_ElibNCo56_1;
	wire w_dff_A_cqpGSbFZ2_1;
	wire w_dff_A_vsuBuerG9_1;
	wire w_dff_A_bzz8OX603_1;
	wire w_dff_A_KAFfH4199_1;
	wire w_dff_B_070zhp4a5_0;
	wire w_dff_A_g6zkyckM7_0;
	wire w_dff_A_JILC84RG8_0;
	wire w_dff_B_BRhfia9R7_0;
	wire w_dff_B_HxMFxo4U0_0;
	wire w_dff_B_fxt2xFq75_0;
	wire w_dff_B_tDfNTOYk1_1;
	wire w_dff_B_D9qgm0eL3_1;
	wire w_dff_B_M3EazxG68_1;
	wire w_dff_A_wjNFHBWa5_0;
	wire w_dff_A_wYgEsu1j2_0;
	wire w_dff_A_fqt9ow0n4_0;
	wire w_dff_A_XM2CG33k7_0;
	wire w_dff_A_8b9rerLI4_0;
	wire w_dff_A_Jl8lj5A05_0;
	wire w_dff_A_HJuIYKJ17_0;
	wire w_dff_A_7vTZhl8j5_0;
	wire w_dff_B_hdAH0NYh6_1;
	wire w_dff_B_jTV28bEn7_1;
	wire w_dff_B_4gd9p14e0_0;
	wire w_dff_B_rwnme35b7_0;
	wire w_dff_A_IjCUvMks7_0;
	wire w_dff_B_sbTVpKbU0_1;
	wire w_dff_A_4tqWAQzS3_2;
	wire w_dff_A_9PX4pKkY6_2;
	wire w_dff_A_9EDswMRN3_0;
	wire w_dff_A_GGPnnmZ95_0;
	wire w_dff_A_MvABrmes5_0;
	wire w_dff_A_GvO4Rd130_0;
	wire w_dff_A_SNNFvQ9E1_1;
	wire w_dff_B_BzB1UFcY7_3;
	wire w_dff_B_NvEx2L4N1_3;
	wire w_dff_A_OsoWLGTJ2_1;
	wire w_dff_A_WiJ4haWB9_1;
	wire w_dff_A_S2ZyZwVv3_1;
	wire w_dff_A_QwkIgFgX5_1;
	wire w_dff_A_DIC2YVHE3_1;
	wire w_dff_A_nyTJjvBJ0_1;
	wire w_dff_A_mg2hnIcf4_2;
	wire w_dff_A_8N7A6szk1_2;
	wire w_dff_A_JMEe3V9P9_2;
	wire w_dff_A_19B2iTki8_2;
	wire w_dff_A_BnrnhBTY2_2;
	wire w_dff_A_IoQihe982_2;
	wire w_dff_A_XgKPFoq79_2;
	wire w_dff_A_L66qirOK6_1;
	wire w_dff_A_rDB1eUaj8_1;
	wire w_dff_A_HDCz66Ce9_1;
	wire w_dff_A_rGUqccYP3_1;
	wire w_dff_A_TgplJfUF8_1;
	wire w_dff_A_hqzwr1cJ4_1;
	wire w_dff_A_67VDDRXs8_2;
	wire w_dff_A_pq0OAUj88_2;
	wire w_dff_A_xWm5OZUZ6_2;
	wire w_dff_A_Sed29K6s0_0;
	wire w_dff_B_V7dT85qn1_1;
	wire w_dff_A_qLkJq7Yp4_0;
	wire w_dff_B_83fBB4Zg2_1;
	wire w_dff_B_IwYH0tVS1_1;
	wire w_dff_B_74lelJ1H2_1;
	wire w_dff_B_aViG2jUQ5_1;
	wire w_dff_B_LvAdtN1b5_1;
	wire w_dff_A_i8yyIplH2_2;
	wire w_dff_A_l5PaLoW59_2;
	wire w_dff_A_AJqdgG8U3_2;
	wire w_dff_A_IuChjonL2_2;
	wire w_dff_A_uAsOX6ck7_2;
	wire w_dff_A_TEyNCykl0_2;
	wire w_dff_A_QATLQh7l7_2;
	wire w_dff_A_duxUuruZ6_2;
	wire w_dff_A_QjmHfwz06_2;
	wire w_dff_A_p6tyzjNY2_2;
	wire w_dff_A_ykCrhBdZ7_2;
	wire w_dff_A_zPf5536V2_2;
	wire w_dff_A_5ZcRhB5p2_2;
	wire w_dff_A_5SDxX0FA8_2;
	wire w_dff_A_eBOdeqzC9_2;
	wire w_dff_A_rLHjHBM64_1;
	wire w_dff_A_DT2oUB298_1;
	wire w_dff_A_Uym4fpnO9_1;
	wire w_dff_A_vTp8Jlp28_1;
	wire w_dff_A_lux5fZqY1_1;
	wire w_dff_A_WKhuoL1k8_1;
	wire w_dff_A_pAbX9eVw6_1;
	wire w_dff_A_NKvMMmvi2_1;
	wire w_dff_A_WPiyapb80_1;
	wire w_dff_A_5Cx11GKH9_1;
	wire w_dff_B_kj2qjmgO0_1;
	wire w_dff_B_B8tKFCJD3_1;
	wire w_dff_B_K3LAVPUE1_1;
	wire w_dff_B_6fn1E8pr1_1;
	wire w_dff_B_iqouE5Dq1_1;
	wire w_dff_B_mtGOdMAp0_1;
	wire w_dff_B_R8tE4bJQ6_1;
	wire w_dff_A_GKaXrJW94_1;
	wire w_dff_B_iPyaFyLN4_1;
	wire w_dff_B_QKPsNrL36_1;
	wire w_dff_B_4MwrLTNz6_1;
	wire w_dff_B_CS9FX0KI7_1;
	wire w_dff_B_HosoUUz22_1;
	wire w_dff_B_sAmJnBz90_1;
	wire w_dff_B_pKbLoEhn9_1;
	wire w_dff_A_K5I8OpjW7_1;
	wire w_dff_A_ECOYXRRD5_1;
	wire w_dff_A_wTccKRfM2_0;
	wire w_dff_A_jpK1YSoA7_0;
	wire w_dff_A_Of2A13lG7_0;
	wire w_dff_A_Ox40Ompz4_0;
	wire w_dff_A_MpFtsz1i4_1;
	wire w_dff_A_eJs5oGEJ3_1;
	wire w_dff_A_tfjwpnlU9_2;
	wire w_dff_B_wOVfCONj9_3;
	wire w_dff_A_aMYZnVF50_0;
	wire w_dff_A_riodS2C01_0;
	wire w_dff_A_KpExEhaJ8_0;
	wire w_dff_A_r33rlOjW2_1;
	wire w_dff_A_gNshOweR9_1;
	wire w_dff_A_Tc8l7UPY8_2;
	wire w_dff_B_4WThtRxK6_3;
	wire w_dff_B_juz86tgt3_3;
	wire w_dff_B_FKRt0SOf7_3;
	wire w_dff_B_PeEuHqG89_3;
	wire w_dff_B_N1UjULZ72_3;
	wire w_dff_B_X3lsKBLN1_3;
	wire w_dff_B_cAwO6GxZ7_3;
	wire w_dff_B_gba4Efgt3_3;
	wire w_dff_B_4AEnmj8c3_3;
	wire w_dff_B_t59Osa8H5_3;
	wire w_dff_A_v18HLLcD7_0;
	wire w_dff_A_tn4be7sx9_0;
	wire w_dff_A_WOCXykHj5_0;
	wire w_dff_A_Vfot0y3l7_0;
	wire w_dff_A_Qt41nr4G6_0;
	wire w_dff_A_ASigP1092_0;
	wire w_dff_A_8tMn8B7I1_0;
	wire w_dff_A_Gs9GXNQm0_0;
	wire w_dff_A_mzUlbWye1_0;
	wire w_dff_A_huMMXZVe7_0;
	wire w_dff_A_cNHhFBwc5_0;
	wire w_dff_A_gkfOwU5h4_0;
	wire w_dff_A_m2APYiOi5_0;
	wire w_dff_A_NGijUakd5_1;
	wire w_dff_A_MsgonRno8_1;
	wire w_dff_A_7gjxmdrv2_1;
	wire w_dff_A_iY2PWA2A5_1;
	wire w_dff_A_AUIfTuPs6_1;
	wire w_dff_A_jpX9c8Ra3_1;
	wire w_dff_A_dJaWcyFF0_1;
	wire w_dff_A_hUETWxeJ4_1;
	wire w_dff_A_129ujZau1_1;
	wire w_dff_A_aQ2sne377_1;
	wire w_dff_A_ezJhyCPW8_0;
	wire w_dff_B_tSgEasV35_0;
	wire w_dff_B_unjhe5ER1_0;
	wire w_dff_A_bkw6TpWq6_0;
	wire w_dff_A_PY9Lnkmo7_0;
	wire w_dff_A_s8jJaLwc5_0;
	wire w_dff_B_XuwBpfWG4_2;
	wire w_dff_A_ZC2btJ5m2_0;
	wire w_dff_A_H2HNYnEs5_0;
	wire w_dff_A_FUOC17pp8_0;
	wire w_dff_A_cYMiPkUq1_1;
	wire w_dff_A_vUuGiq4C9_1;
	wire w_dff_A_4eyTO76A5_1;
	wire w_dff_A_U3aJIZ4Z3_1;
	wire w_dff_A_MMWmBxtS2_1;
	wire w_dff_A_W2piALF04_1;
	wire w_dff_A_jYrslpcA9_1;
	wire w_dff_A_5GJOdGyi0_1;
	wire w_dff_A_pX4P1kdQ5_0;
	wire w_dff_A_feSviSIp1_0;
	wire w_dff_A_NlApwIhT5_0;
	wire w_dff_A_Sc2SMKNB7_0;
	wire w_dff_A_LBdEB4Xo8_2;
	wire w_dff_A_BFxkYivm6_2;
	wire w_dff_A_kZSg5MXX5_1;
	wire w_dff_A_S5Gh99jH1_1;
	wire w_dff_A_5uPZEH5K0_1;
	wire w_dff_A_kWMIyWPc4_1;
	wire w_dff_A_h8rFwdzc6_1;
	wire w_dff_B_XvG3bD4C6_1;
	wire w_dff_B_SfwD23T13_1;
	wire w_dff_A_hUotwwMm3_1;
	wire w_dff_A_cAGlh6xh6_1;
	wire w_dff_A_klRu9zIB9_1;
	wire w_dff_A_iGxtas971_1;
	wire w_dff_A_lqvx0U101_1;
	wire w_dff_A_aurhMe533_1;
	wire w_dff_A_hbkPjEYw5_1;
	wire w_dff_B_xm9n2cNj2_0;
	wire w_dff_B_ZekPhHNU8_1;
	wire w_dff_A_Sb7QOQec3_2;
	wire w_dff_A_Vl47BYZt6_1;
	wire w_dff_A_Uvjf0yqw3_1;
	wire w_dff_A_HEZv31Xe4_1;
	wire w_dff_A_JWxZI3X23_1;
	wire w_dff_A_CRcdYjRi2_2;
	wire w_dff_A_aBRlDjTD7_2;
	wire w_dff_A_JI7m7Q3p0_2;
	wire w_dff_A_iD7IMbK61_2;
	wire w_dff_A_IxvVKXhq0_0;
	wire w_dff_A_jDb5vWbQ6_0;
	wire w_dff_B_5zQTNqNL4_3;
	wire w_dff_A_xK9GoD8d5_0;
	wire w_dff_B_Q7E4iDB55_1;
	wire w_dff_B_CVVTHKpS5_1;
	wire w_dff_A_4q1hYdfh3_0;
	wire w_dff_A_PNkC3uu93_0;
	wire w_dff_B_jI44hNRp8_2;
	wire w_dff_A_buhOiGsc8_0;
	wire w_dff_A_Upu1yvLo5_0;
	wire w_dff_A_zu46DcNC2_0;
	wire w_dff_A_3kBbDxDQ4_1;
	wire w_dff_A_qv2urgCy8_1;
	wire w_dff_A_nmvMlbAs9_1;
	wire w_dff_A_PaFgiKnh5_1;
	wire w_dff_A_KT1GeWuA7_1;
	wire w_dff_A_0i8wc61A6_1;
	wire w_dff_A_2q2vU2484_1;
	wire w_dff_A_GroD6Vqu4_2;
	wire w_dff_A_Bf3qpHA62_2;
	wire w_dff_A_NW2y806O4_2;
	wire w_dff_A_jokAWxaH0_2;
	wire w_dff_A_q27zPIaQ0_2;
	wire w_dff_B_eEc63flA4_0;
	wire w_dff_B_iK4y7oQM2_1;
	wire w_dff_A_eWQJRtlK4_0;
	wire w_dff_A_6kitU1zB8_1;
	wire w_dff_B_dUa0MRE69_1;
	wire w_dff_A_1j4RLxNY6_0;
	wire w_dff_A_OfTuXaEp5_1;
	wire w_dff_A_8ywYSxFS9_1;
	wire w_dff_B_SfR3MZBx3_1;
	wire w_dff_A_Foq3VPLQ3_0;
	wire w_dff_A_JKLtRAxP4_0;
	wire w_dff_A_Fq3Yi8Dz9_2;
	wire w_dff_A_eb1XlFli1_0;
	wire w_dff_A_nvhxGLEV3_0;
	wire w_dff_A_L5VotdaR3_0;
	wire w_dff_A_NneLSLTL0_2;
	wire w_dff_A_5xH6wiIu1_0;
	wire w_dff_A_Hpe11eud5_1;
	wire w_dff_A_Tw4If2hQ9_2;
	wire w_dff_A_iyld7ep81_0;
	wire w_dff_A_p9XJx9lM5_0;
	wire w_dff_A_IDL7g5my3_0;
	wire w_dff_A_4v46mBNE5_2;
	wire w_dff_A_pNXeXqfn6_2;
	wire w_dff_A_MOvQLspi1_2;
	wire w_dff_A_tStlNfMY4_0;
	wire w_dff_A_Lpp4XiX75_0;
	wire w_dff_A_hcovNpaa2_0;
	wire w_dff_A_WSnSbauz7_1;
	wire w_dff_A_mbdOxSkR8_1;
	wire w_dff_A_Sl0epb350_2;
	wire w_dff_A_glcBLkLD3_0;
	wire w_dff_A_gkmhSzvi0_2;
	wire w_dff_B_84Cmest04_3;
	wire w_dff_A_V5DDT1wr1_0;
	wire w_dff_A_7TYcbolV4_0;
	wire w_dff_A_9mALEgny1_0;
	wire w_dff_A_1mS2KaGS0_1;
	wire w_dff_A_9OE3YKL51_1;
	wire w_dff_A_5pSo3KrS6_1;
	wire w_dff_A_USeJePYc5_1;
	wire w_dff_A_ihptJDIZ3_1;
	wire w_dff_A_Aw05G7vG7_1;
	wire w_dff_A_IChldhM89_2;
	wire w_dff_A_LSCJ1cll4_2;
	wire w_dff_A_3nvPKuqC5_2;
	wire w_dff_A_pwVsbGq33_1;
	wire w_dff_A_VU6hs2k22_1;
	wire w_dff_A_hQzJJwvS2_1;
	wire w_dff_A_ldf0b7vZ9_1;
	wire w_dff_A_5hhZrTyZ5_1;
	wire w_dff_A_IXDS5e1t1_1;
	wire w_dff_A_QJscMUJO4_1;
	wire w_dff_A_7ckStsVJ9_1;
	wire w_dff_A_tDgj3zKQ2_1;
	wire w_dff_A_Rw1rXM5c4_1;
	wire w_dff_A_xsATXNB53_1;
	wire w_dff_A_6D4cYah37_0;
	wire w_dff_A_zLCi2JRf0_0;
	wire w_dff_A_gqGYYdE64_0;
	wire w_dff_A_qQCaPRpQ6_2;
	wire w_dff_A_WkeJW0YD8_1;
	wire w_dff_A_ST5xq0FZ2_1;
	wire w_dff_A_lPWQYr1d8_1;
	wire w_dff_A_t6E3SN1s2_1;
	wire w_dff_A_IkVwVZtL1_1;
	wire w_dff_A_PRGlszqX1_1;
	wire w_dff_A_4IR1WgpV2_1;
	wire w_dff_A_oen9cJMi5_1;
	wire w_dff_A_lGvYCjGC7_1;
	wire w_dff_B_2P7cnQJX2_0;
	wire w_dff_A_TLSq3PvQ6_1;
	wire w_dff_A_S9P1YKLL9_1;
	wire w_dff_A_m0hJMGqo6_2;
	wire w_dff_A_HNdEweL63_0;
	wire w_dff_A_WCbEeCWh0_0;
	wire w_dff_A_hUPZcTEs3_0;
	wire w_dff_A_TkQf8VUZ5_0;
	wire w_dff_A_vLlAh7BJ3_2;
	wire w_dff_A_z10QLZuZ2_2;
	wire w_dff_A_InqCPwIB5_0;
	wire w_dff_A_oaUI5gpT5_0;
	wire w_dff_A_wNcPZAgX3_0;
	wire w_dff_A_QvcNGvMq9_0;
	wire w_dff_A_4xah8S4p1_0;
	wire w_dff_A_yRq5rjgp0_0;
	wire w_dff_A_uD75D0407_0;
	wire w_dff_A_gfuM77xF0_0;
	wire w_dff_A_CmPNRQtJ1_0;
	wire w_dff_A_svdtNH7T0_0;
	wire w_dff_A_wNWBEMgF1_0;
	wire w_dff_A_LeCjiudG4_0;
	wire w_dff_A_xmAUHCQt2_0;
	wire w_dff_A_4eBVXyyi9_0;
	wire w_dff_A_sGlV1iAw4_0;
	wire w_dff_A_FNNpIzeO2_0;
	wire w_dff_A_GSVGRiUH8_0;
	wire w_dff_A_HV17DwMK2_0;
	wire w_dff_A_g0ILb4HI3_0;
	wire w_dff_A_96sSh9NM1_0;
	wire w_dff_A_xqfXnHMP0_2;
	wire w_dff_A_eq1D3zvb3_2;
	wire w_dff_A_q2I5Dvgu0_2;
	wire w_dff_A_VHMWrw1t4_2;
	wire w_dff_B_gUbshfRD5_0;
	wire w_dff_B_jhkjn9Zl4_0;
	wire w_dff_B_Uoi2yFh10_0;
	wire w_dff_B_MVjIrnIv0_0;
	wire w_dff_B_Jm6O73Tk5_0;
	wire w_dff_B_x3Qlmyke3_0;
	wire w_dff_B_HrePYNtF4_0;
	wire w_dff_B_esu3p3g65_0;
	wire w_dff_B_ey1uRs3A9_0;
	wire w_dff_B_KILiCMsR7_0;
	wire w_dff_B_d5Jx423d6_0;
	wire w_dff_B_5Y5w8VxY9_0;
	wire w_dff_B_OsgGniXa9_0;
	wire w_dff_B_0347uEnU6_0;
	wire w_dff_B_v7oDXAX19_0;
	wire w_dff_B_lZt7TFpo7_0;
	wire w_dff_B_yjk0X1Kn2_0;
	wire w_dff_B_qYAwu6Vt6_0;
	wire w_dff_B_nPiJfuQE9_0;
	wire w_dff_B_0B4BLuop5_1;
	wire w_dff_B_OBGnQCwn1_1;
	wire w_dff_B_i9avABce2_1;
	wire w_dff_B_9tcoZrT43_1;
	wire w_dff_B_JS3lg73m1_1;
	wire w_dff_B_OtNKk3rR4_1;
	wire w_dff_B_m5hu5P1z5_1;
	wire w_dff_B_uWVyz5F21_1;
	wire w_dff_B_wuYXi2Et7_1;
	wire w_dff_B_7mRl6pvf8_1;
	wire w_dff_A_c3JiXYI61_2;
	wire w_dff_A_YA6qdyAm1_2;
	wire w_dff_A_ljs2Hp0w4_1;
	wire w_dff_B_U39WYkVf8_0;
	wire w_dff_B_SkQjwMPL6_1;
	wire w_dff_B_bhIyt8lL5_1;
	wire w_dff_B_G0JmWut19_1;
	wire w_dff_B_6F5f6ggu3_1;
	wire w_dff_B_gwOPQG2O0_1;
	wire w_dff_B_JKPtkImr4_1;
	wire w_dff_B_5EK2mvuK0_1;
	wire w_dff_B_UN3D2OQa0_0;
	wire w_dff_B_E9c8Q9st3_0;
	wire w_dff_A_lMfFZB3f7_1;
	wire w_dff_A_qN1R3Qou6_1;
	wire w_dff_A_uWkQqW285_1;
	wire w_dff_A_7StndMra4_1;
	wire w_dff_A_kjlwGibM2_1;
	wire w_dff_A_6jSZxBw04_1;
	wire w_dff_A_GfGyIHtP2_1;
	wire w_dff_A_ciDKAQsw9_1;
	wire w_dff_A_LBtMs73U2_1;
	wire w_dff_A_rg1LxCCa7_1;
	wire w_dff_A_U290aPjM7_1;
	wire w_dff_A_EQXPIS1N9_1;
	wire w_dff_A_w7y9CaQb5_1;
	wire w_dff_B_ePa9ZGLr2_2;
	wire w_dff_A_BTbKi5Jb9_2;
	wire w_dff_A_CH84g8MI4_2;
	wire w_dff_A_wVumRsB25_2;
	wire w_dff_A_y94MvvgY3_2;
	wire w_dff_A_Y4IRGbEd4_2;
	wire w_dff_B_HZ22xhO44_1;
	wire w_dff_B_c8tJW17L9_1;
	wire w_dff_B_bM6Z8sTg3_1;
	wire w_dff_B_C3TFEuEu2_1;
	wire w_dff_B_JjKRjUFL6_1;
	wire w_dff_A_stEpA5I53_1;
	wire w_dff_A_ltrH5PPd3_1;
	wire w_dff_A_DuemyRDn3_1;
	wire w_dff_A_qtKn5Lti2_1;
	wire w_dff_A_80AmkYVV1_1;
	wire w_dff_A_TpXMtvpr4_1;
	wire w_dff_A_OkWM4bmB6_1;
	wire w_dff_A_gA8xVCXm4_0;
	wire w_dff_A_uWVn8Rrn5_0;
	wire w_dff_A_nOmrw2Ua8_0;
	wire w_dff_A_NXxAqgyB4_0;
	wire w_dff_A_NdelxAfF1_0;
	wire w_dff_A_SZQgHzmo0_0;
	wire w_dff_A_KOwUvZYr6_0;
	wire w_dff_A_x46xDeyz9_0;
	wire w_dff_A_1IuIiZHH3_0;
	wire w_dff_A_5DSV6Ion8_0;
	wire w_dff_A_5Z60IyI02_0;
	wire w_dff_A_RoCQJvsK0_0;
	wire w_dff_A_EUXMbap50_0;
	wire w_dff_A_c6yKdYy39_0;
	wire w_dff_A_eYoFTxR21_0;
	wire w_dff_A_0btEpyaX9_0;
	wire w_dff_A_kwSz5bpb4_0;
	wire w_dff_B_7gkPcXSF8_2;
	wire w_dff_B_VeZvpyRk9_2;
	wire w_dff_A_y9p7nX1o0_1;
	wire w_dff_A_oL2g4Aja4_1;
	wire w_dff_A_4fdym84U1_1;
	wire w_dff_A_on1XCH9Z5_1;
	wire w_dff_A_AuzC6GbR3_1;
	wire w_dff_A_yOnSseSd2_1;
	wire w_dff_A_3c13K7Dr4_1;
	wire w_dff_A_A412UALn6_1;
	wire w_dff_A_KP6Onlmi6_1;
	wire w_dff_A_TDWXxzhw2_1;
	wire w_dff_A_Tmt5fEaE8_2;
	wire w_dff_B_kxUpVWOD1_0;
	wire w_dff_B_FNT2I8yG7_1;
	wire w_dff_A_JafzU21e9_0;
	wire w_dff_A_TJJFYm634_2;
	wire w_dff_A_gUId8wQW0_2;
	wire w_dff_A_OakfWlda1_2;
	wire w_dff_A_YJMKUC0n2_2;
	wire w_dff_B_jofkP0gt7_1;
	wire w_dff_B_tzD22bHC5_1;
	wire w_dff_A_hh2mcvLz5_0;
	wire w_dff_A_PLKQmBID7_0;
	wire w_dff_A_rsjm53rT8_0;
	wire w_dff_A_IhhqZhb00_2;
	wire w_dff_A_CVQrhsZZ8_2;
	wire w_dff_A_M19FBHYK2_2;
	wire w_dff_A_358nN0ZP7_2;
	wire w_dff_A_KDDCxiPb5_2;
	wire w_dff_A_KcfKXmrH4_2;
	wire w_dff_A_ZuWMt4rq6_2;
	wire w_dff_B_PBRYjV6g2_2;
	wire w_dff_A_4qAEFu3Q1_1;
	wire w_dff_B_sEJck0bU6_0;
	wire w_dff_B_jZXeDG7D1_1;
	wire w_dff_B_ZzFzfLkP7_0;
	wire w_dff_B_Ky2Cc9Hx3_1;
	wire w_dff_A_YX2jxMvL1_1;
	wire w_dff_A_OSrep8xP9_0;
	wire w_dff_A_iM2l6I6p5_0;
	wire w_dff_B_n2ov5BJX8_2;
	wire w_dff_B_jv55Wmyx7_2;
	wire w_dff_B_AW8r6ZLe9_2;
	wire w_dff_A_wNyQiAG10_0;
	wire w_dff_A_TacHl0VK9_0;
	wire w_dff_A_ZNAEuJrn7_0;
	wire w_dff_A_ugD9qJRX6_0;
	wire w_dff_A_LYdkwNnD8_1;
	wire w_dff_A_NJrYn3Gh1_1;
	wire w_dff_A_CvIrWNMh2_1;
	wire w_dff_A_FqhyJarJ1_1;
	wire w_dff_A_ocVvc1Do8_1;
	wire w_dff_A_UqjqprCo5_1;
	wire w_dff_A_rXYTpAJ86_2;
	wire w_dff_A_mo4gCKNG7_2;
	wire w_dff_A_i0jTaJLg0_2;
	wire w_dff_A_3NsMfUTc1_2;
	wire w_dff_A_IN7IVVj00_2;
	wire w_dff_A_SF6wwOlN4_2;
	wire w_dff_B_YFbsgk1z0_0;
	wire w_dff_B_kDISMzON5_0;
	wire w_dff_B_ADIfAWjU4_0;
	wire w_dff_B_x7MrCcHz2_0;
	wire w_dff_B_wfxsMGK99_0;
	wire w_dff_B_J5FNLLdD9_0;
	wire w_dff_B_oZBYRYpI6_0;
	wire w_dff_B_oBpoNX670_0;
	wire w_dff_B_IEWSCVWl1_0;
	wire w_dff_B_JSg1zwAr4_0;
	wire w_dff_B_G6Afcqu25_0;
	wire w_dff_B_FDhpUtO37_1;
	wire w_dff_B_zDJNFwb65_1;
	wire w_dff_B_DPIhoEAz3_1;
	wire w_dff_A_WVPlABGB7_0;
	wire w_dff_A_h9RHD1Wf3_0;
	wire w_dff_B_OSIpj3g87_2;
	wire w_dff_B_YdLpiqEO5_2;
	wire w_dff_B_yzs8FEqX4_2;
	wire w_dff_B_AlB55ZbM5_2;
	wire w_dff_B_Iaidy7DC6_2;
	wire w_dff_B_SsKWya6U1_2;
	wire w_dff_B_alvihZuQ4_2;
	wire w_dff_B_FA3jSb7Y0_2;
	wire w_dff_B_Q5W7Uo8m9_2;
	wire w_dff_B_YJZ1q6Pt9_2;
	wire w_dff_B_fQAwXlFt3_2;
	wire w_dff_B_D23ryYxv9_2;
	wire w_dff_A_DUQCjTfN9_0;
	wire w_dff_A_VYqd4jNF5_0;
	wire w_dff_A_MIM2syFJ0_0;
	wire w_dff_A_d8qdPqnj3_0;
	wire w_dff_A_wR4gVw5a5_0;
	wire w_dff_A_DaEx89iW2_0;
	wire w_dff_A_pW7PwdB17_0;
	wire w_dff_A_EZENiS5G4_0;
	wire w_dff_A_9HPwoaT46_0;
	wire w_dff_A_QunGUQS16_0;
	wire w_dff_A_Csaffvy12_0;
	wire w_dff_A_WSKbKUGS6_0;
	wire w_dff_A_6TlGoEjs4_0;
	wire w_dff_A_JnceUb9N1_0;
	wire w_dff_A_DIXrA4Ol2_0;
	wire w_dff_A_v8jUiXyq4_1;
	wire w_dff_A_JkE1apyh3_1;
	wire w_dff_A_Pl5Lvpbu9_1;
	wire w_dff_A_87EKpOGc5_1;
	wire w_dff_A_pCebwpN17_1;
	wire w_dff_A_eaMzEqWO4_1;
	wire w_dff_A_baz8KZBT4_1;
	wire w_dff_A_19Z73k5e8_1;
	wire w_dff_A_MXuOOcBD5_1;
	wire w_dff_A_QEqPepFN4_1;
	wire w_dff_A_sMBrycq73_1;
	wire w_dff_A_kMGXyWAW2_1;
	wire w_dff_B_tz7vm4622_1;
	wire w_dff_B_Is9FsIDa4_1;
	wire w_dff_B_AHzQ1bo01_0;
	wire w_dff_B_xjVLJxhP0_0;
	wire w_dff_B_TbBjUpTs8_0;
	wire w_dff_B_Q7Fir2LH9_0;
	wire w_dff_A_lOC6SxJh8_0;
	wire w_dff_A_sWAv6bEr5_0;
	wire w_dff_A_9dufPMrV9_0;
	wire w_dff_A_cwqlShOa0_0;
	wire w_dff_A_uS9qzP8y1_0;
	wire w_dff_A_rKYk0v846_0;
	wire w_dff_A_RQoPWnei5_2;
	wire w_dff_A_dGHbC1GY5_2;
	wire w_dff_A_IbaEiGjv0_2;
	wire w_dff_A_KIv1QUks9_2;
	wire w_dff_A_K2zayzws2_2;
	wire w_dff_A_ag8tbrgU9_1;
	wire w_dff_A_ucRjPzjK9_1;
	wire w_dff_A_6Du1Sg0U4_1;
	wire w_dff_A_cJouWD972_1;
	wire w_dff_B_0KfscTS83_0;
	wire w_dff_B_Cur9DqbV8_1;
	wire w_dff_B_NQuomSmT9_1;
	wire w_dff_B_dihszsxc3_1;
	wire w_dff_B_ZBZ2h3Xx8_1;
	wire w_dff_B_gJKpywDe3_1;
	wire w_dff_B_EEf1xN4e2_1;
	wire w_dff_A_45ISubVn8_1;
	wire w_dff_A_D0J2IDl14_1;
	wire w_dff_A_JglAYIaa8_1;
	wire w_dff_A_RI7rXPLc3_1;
	wire w_dff_A_B7oKu7HL8_1;
	wire w_dff_A_jkr9Psjl4_1;
	wire w_dff_A_afZGM9lt3_1;
	wire w_dff_A_t4w4FOuA7_0;
	wire w_dff_A_L6sGAcEm1_0;
	wire w_dff_A_bYjMFFCb7_1;
	wire w_dff_A_7jgF267z0_1;
	wire w_dff_A_0Db6W2Cs6_2;
	wire w_dff_A_Fg9V4URE0_2;
	wire w_dff_A_ImOe7M6h4_2;
	wire w_dff_A_C7zORkRV9_2;
	wire w_dff_B_Fapaexz99_0;
	wire w_dff_B_NKyFj8YE6_1;
	wire w_dff_A_rXySgHot6_1;
	wire w_dff_A_7iIMNZtS0_1;
	wire w_dff_A_CarUYmxb5_0;
	wire w_dff_A_eMdoammx6_0;
	wire w_dff_B_Vaz3kXuR5_0;
	wire w_dff_B_8Zp4ATZI9_0;
	wire w_dff_B_Ucp90mZP1_0;
	wire w_dff_A_UYNv0ANo9_0;
	wire w_dff_A_SdSKvjXD5_1;
	wire w_dff_A_VwBB50Uj6_1;
	wire w_dff_B_5KEEzPuo0_1;
	wire w_dff_A_Mo0cBftB0_0;
	wire w_dff_A_GzWpiUJQ3_1;
	wire w_dff_A_mYwDRUot2_1;
	wire w_dff_B_3wc4Nap28_1;
	wire w_dff_A_uhsIQN6V4_0;
	wire w_dff_A_A2GZ60vW9_0;
	wire w_dff_A_cSQndLGD4_1;
	wire w_dff_B_StTsmORO0_1;
	wire w_dff_A_0k8lOAaf5_0;
	wire w_dff_A_BgJsq9Jr0_0;
	wire w_dff_A_H1PaAqjw8_0;
	wire w_dff_A_BEGkXa3p6_1;
	wire w_dff_B_bwLRLfw68_1;
	wire w_dff_A_6ICbiHw30_0;
	wire w_dff_A_2d6Dcsjh5_0;
	wire w_dff_A_S32Xyl0Y1_0;
	wire w_dff_B_QkIf4nKc5_0;
	wire w_dff_B_RNCmrvdz4_1;
	wire w_dff_B_bsFFLQAk9_1;
	wire w_dff_A_omW0t1800_0;
	wire w_dff_A_bo21x2F13_1;
	wire w_dff_A_sxn8HzZ62_1;
	wire w_dff_B_258BLKiQ6_3;
	wire w_dff_A_x8EnYzKe3_0;
	wire w_dff_A_lIpRGklZ4_0;
	wire w_dff_A_JSUas53y4_0;
	wire w_dff_A_zRCf7qQ64_0;
	wire w_dff_A_H425gTGF7_1;
	wire w_dff_A_K7zQGfJv1_1;
	wire w_dff_A_rP4Wqp0u9_1;
	wire w_dff_A_ffHonvao3_1;
	wire w_dff_A_VWxaRlu41_1;
	wire w_dff_A_JYLhTTJa8_1;
	wire w_dff_A_OG0liO9r0_2;
	wire w_dff_A_UiraPyUx6_2;
	wire w_dff_A_7uH9SFkI4_2;
	wire w_dff_A_YnWKwscH0_2;
	wire w_dff_A_VsQiZBHr3_2;
	wire w_dff_B_UJdiGdRT3_1;
	wire w_dff_A_NUipEbn84_0;
	wire w_dff_A_yqjocQrS5_1;
	wire w_dff_A_oZTYeJI77_1;
	wire w_dff_B_Ue2RQK7M0_3;
	wire w_dff_A_2giIdlF59_0;
	wire w_dff_A_jOcXBYqR5_0;
	wire w_dff_A_a0tbMto75_0;
	wire w_dff_A_NyAn2Iwl2_0;
	wire w_dff_A_C9EHR4nj9_1;
	wire w_dff_A_gMChsRxG9_1;
	wire w_dff_A_zp28VQpV5_1;
	wire w_dff_B_gJhV3tqA0_1;
	wire w_dff_A_2dgVSwNM7_0;
	wire w_dff_A_200NXoVi2_1;
	wire w_dff_A_gqiZzrv91_1;
	wire w_dff_A_BoSwSDQu9_2;
	wire w_dff_A_HK9ADDy74_2;
	wire w_dff_A_9tsMg1EG3_2;
	wire w_dff_A_oN5HW0EJ7_2;
	wire w_dff_A_snz3ufaQ5_0;
	wire w_dff_B_zh9yCmRY4_1;
	wire w_dff_B_2COnfUBI7_1;
	wire w_dff_A_vLQ3zUm74_0;
	wire w_dff_A_7UYuPrNg3_2;
	wire w_dff_A_7ItgWThO1_2;
	wire w_dff_A_du6Mz9Sf0_2;
	wire w_dff_B_6xukRhGQ8_3;
	wire w_dff_A_YVqMVdyg0_0;
	wire w_dff_A_vTodZrR70_0;
	wire w_dff_A_4FNS6t941_0;
	wire w_dff_A_8ScpLo9y0_1;
	wire w_dff_A_bqMEHnsB8_1;
	wire w_dff_A_ihL37Hwh1_1;
	wire w_dff_A_G2By6A9Y4_2;
	wire w_dff_A_4vwKSeA09_2;
	wire w_dff_A_0X6XxiFk2_2;
	wire w_dff_A_RGIhfKH47_2;
	wire w_dff_A_YFIgcURp7_2;
	wire w_dff_B_sXS2qhCh4_1;
	wire w_dff_B_0MDGyf1J3_1;
	wire w_dff_B_mxxOHVf20_1;
	wire w_dff_A_tSgzqsuZ7_0;
	wire w_dff_A_c6yY6VmJ3_0;
	wire w_dff_A_cdMgZoFv3_0;
	wire w_dff_A_oZKcgZqF6_1;
	wire w_dff_A_H47IajYI2_1;
	wire w_dff_A_vPJtS8657_1;
	wire w_dff_A_RXlqpMv45_1;
	wire w_dff_A_CriMmbkp3_1;
	wire w_dff_A_DwvbHT6D0_1;
	wire w_dff_A_8yUT8lxV7_2;
	wire w_dff_A_REAC3s3q9_2;
	wire w_dff_A_f2gP5ZVl5_2;
	wire w_dff_A_1F6tAt515_0;
	wire w_dff_B_BsXdgS7b2_1;
	wire w_dff_B_Se3SyzF83_1;
	wire w_dff_B_6CGQjU6n3_1;
	wire w_dff_B_ak0qsddl7_1;
	wire w_dff_A_fMp54LYZ8_0;
	wire w_dff_A_4qNnXdDp7_1;
	wire w_dff_A_ZakBxiGE0_1;
	wire w_dff_A_QQ58oc3Q7_1;
	wire w_dff_B_4IsApSZi4_3;
	wire w_dff_A_vF4BLX0l8_0;
	wire w_dff_A_hDLByAA12_0;
	wire w_dff_A_DTh41GJm9_0;
	wire w_dff_A_wpZAXwbu1_0;
	wire w_dff_A_WMPP5CPu1_1;
	wire w_dff_A_fcXknSva2_1;
	wire w_dff_A_LDaXALsP2_1;
	wire w_dff_A_QrOT8bW25_1;
	wire w_dff_A_3hQrz8kn9_1;
	wire w_dff_A_BvM1Ub6G2_1;
	wire w_dff_A_vc9gITJm9_2;
	wire w_dff_A_rLV5VGiu1_2;
	wire w_dff_A_5PKAwhTq9_2;
	wire w_dff_A_VR5MfvCi8_2;
	wire w_dff_A_Vdnrw3Gg7_2;
	wire w_dff_B_K9GTT0wg4_1;
	wire w_dff_B_qUqFTHDw7_1;
	wire w_dff_A_9iZVWSZd3_0;
	wire w_dff_A_4nlF569f1_1;
	wire w_dff_A_nw1q9Y2Y4_1;
	wire w_dff_B_kmWkYj5y6_3;
	wire w_dff_A_IOBuc7UP6_0;
	wire w_dff_A_UXUCxW953_0;
	wire w_dff_A_0ZgOqPy23_0;
	wire w_dff_A_JzflguxI3_0;
	wire w_dff_A_ahzRbivf3_1;
	wire w_dff_A_sbbtQKiI3_1;
	wire w_dff_A_tMFfg7EN9_1;
	wire w_dff_A_YubtN7nb5_1;
	wire w_dff_A_WPD1xqto1_1;
	wire w_dff_A_4Ezae2bB4_1;
	wire w_dff_A_lj0sqnUK5_2;
	wire w_dff_A_p882NBI01_2;
	wire w_dff_A_BO0txMcK0_2;
	wire w_dff_A_spaQFyFL5_2;
	wire w_dff_A_UCUdfuzf8_2;
	wire w_dff_B_E6Ivhjnj0_1;
	wire w_dff_A_6GrVvIMI8_1;
	wire w_dff_A_WxCttBwT4_1;
	wire w_dff_A_MkVZMfz07_2;
	wire w_dff_B_Vi4jOAZY0_3;
	wire w_dff_A_fCpTHnQo3_0;
	wire w_dff_A_QdSxXu2G1_0;
	wire w_dff_A_O4E25Dpd2_0;
	wire w_dff_A_kQSqkvHw5_0;
	wire w_dff_A_CjFOTSwv9_1;
	wire w_dff_A_gPeqJYEJ5_1;
	wire w_dff_A_lS1IRETb5_1;
	wire w_dff_B_61LdT2ER1_1;
	wire w_dff_A_AN3A2DOu0_0;
	wire w_dff_A_AB26oXG68_0;
	wire w_dff_A_Xcenn3811_2;
	wire w_dff_A_ybWsuH9i4_1;
	wire w_dff_A_RyuxyeXw5_1;
	wire w_dff_A_plKmlqta5_2;
	wire w_dff_A_JfEtQdhX2_2;
	wire w_dff_A_LUYOThiy8_2;
	wire w_dff_A_UIuZFd6I2_2;
	wire w_dff_A_xejFgTk11_1;
	wire w_dff_A_oVA4nxdI7_2;
	wire w_dff_B_6LN4FPEo8_1;
	wire w_dff_B_84LvMF523_1;
	wire w_dff_A_SsgkcA2G8_0;
	wire w_dff_A_9TwE1wRF8_1;
	wire w_dff_A_IK6a6du75_1;
	wire w_dff_A_RObb8iE97_2;
	wire w_dff_A_dGVpQ0Fx4_2;
	wire w_dff_B_bVA2yGk26_3;
	wire w_dff_A_SHIZ7K8x2_0;
	wire w_dff_A_hbNxLAaW1_0;
	wire w_dff_A_DeB1ZDg64_0;
	wire w_dff_A_NCvTwNFW0_0;
	wire w_dff_A_XIfLBDJu3_1;
	wire w_dff_A_cggXNrML1_1;
	wire w_dff_A_ZHtEhEHW0_1;
	wire w_dff_A_ooErNWfW8_1;
	wire w_dff_A_g1La7HFk9_1;
	wire w_dff_A_4pKE69fy7_1;
	wire w_dff_A_fmwFvSQN3_2;
	wire w_dff_A_SDrAvg241_2;
	wire w_dff_A_N8zD4JvR7_2;
	wire w_dff_A_CHL3mOnJ1_2;
	wire w_dff_A_n0anY7p45_2;
	wire w_dff_A_SykPmhEG9_0;
	wire w_dff_A_dC6B2DkC2_1;
	wire w_dff_A_ep1c18em2_2;
	wire w_dff_B_Vrst2SN82_1;
	wire w_dff_B_Iy7RRtdp3_1;
	wire w_dff_A_HxChay362_0;
	wire w_dff_A_ag2tn0BI5_1;
	wire w_dff_A_wZ2op9mq3_2;
	wire w_dff_A_7MBIRTJ58_1;
	wire w_dff_A_eeLzT7dy9_1;
	wire w_dff_A_8KgFoi4m0_2;
	wire w_dff_A_kK2bVqdC6_2;
	wire w_dff_B_t2bDAX2O6_3;
	wire w_dff_A_lXLSYaYB8_0;
	wire w_dff_A_yK6I2eTU0_0;
	wire w_dff_A_vZS4jv8O6_0;
	wire w_dff_A_yiBZlk3W0_0;
	wire w_dff_A_VtORDEFH0_0;
	wire w_dff_A_IkiIFhRa1_0;
	wire w_dff_A_BVx3UiRc1_0;
	wire w_dff_A_buwzuigq6_2;
	wire w_dff_A_7JRegl3A8_2;
	wire w_dff_A_lV1aM1ki1_2;
	wire w_dff_A_XDgcLo2e7_1;
	wire w_dff_A_Xnc6CWE06_2;
	wire w_dff_A_A874vAr96_2;
	wire w_dff_A_QmFPONVY2_1;
	wire w_dff_A_rVnLMMcE5_1;
	wire w_dff_A_wIENmvx61_1;
	wire w_dff_A_mJkvDEot9_1;
	wire w_dff_A_LvXNHbYf9_1;
	wire w_dff_A_8x1s1C3x8_1;
	wire w_dff_A_xusRBEtk2_1;
	wire w_dff_A_1kC47ywc8_1;
	wire w_dff_A_SKrsXSo69_1;
	wire w_dff_A_aUNEpBAB7_1;
	wire w_dff_A_TZBFGHtN2_1;
	wire w_dff_A_tyeBYNT06_1;
	wire w_dff_A_GQEUk9Tg1_1;
	wire w_dff_A_SXDXHoG39_1;
	wire w_dff_A_K3YYi3n91_1;
	wire w_dff_A_8mp6hujI9_1;
	wire w_dff_A_18S8GhZa8_1;
	wire w_dff_A_FWMkj3kg1_2;
	wire w_dff_A_8tnFSRF75_2;
	wire w_dff_A_xA34DnvM7_2;
	wire w_dff_A_Jq8YDfEw5_2;
	wire w_dff_A_ldeQwlnR2_2;
	wire w_dff_A_bM15YuWf9_2;
	wire w_dff_A_Sfju9m4q5_2;
	wire w_dff_A_JmgRWSyj3_2;
	wire w_dff_A_qL7zN0U73_1;
	wire w_dff_A_4SBju4m50_1;
	wire w_dff_A_joNNIwb78_1;
	wire w_dff_A_gBzpWDv81_1;
	wire w_dff_A_wG3p4WJa2_2;
	wire w_dff_A_m8tm4q3K5_2;
	wire w_dff_A_nO0Ix8Q14_2;
	wire w_dff_A_hfKCLmh88_2;
	wire w_dff_A_2jP08G0W9_1;
	wire w_dff_A_P7w9oMCp7_1;
	wire w_dff_A_m1PNJ7gt1_2;
	wire w_dff_A_ulNocj2a9_2;
	wire w_dff_A_rpIbK18c5_2;
	wire w_dff_A_1PNMuPvk5_0;
	wire w_dff_A_L42a4hZQ2_0;
	wire w_dff_A_cgHyoynU1_0;
	wire w_dff_A_hg5jQ5yC8_0;
	wire w_dff_A_abu6zKXv4_0;
	wire w_dff_A_lOz16oa14_0;
	wire w_dff_A_jKkpTKZP7_0;
	wire w_dff_A_fQgA9Y8k2_0;
	wire w_dff_A_4bpCAS7U3_0;
	wire w_dff_A_Ya2MDvDg5_0;
	wire w_dff_A_ufVxp2va3_0;
	wire w_dff_A_acv2Moz75_0;
	wire w_dff_A_wCjJ2qrj9_0;
	wire w_dff_A_u33ZBVVq4_1;
	wire w_dff_A_7ygdSbNz5_1;
	wire w_dff_A_JjFCf3SU3_1;
	wire w_dff_A_4fSVkS468_1;
	wire w_dff_A_7ahHDM2d4_1;
	wire w_dff_A_f2bK6iJ99_1;
	wire w_dff_A_9pW0ku0l4_1;
	wire w_dff_A_SqUpkORK8_1;
	wire w_dff_A_e0IOgCa68_1;
	wire w_dff_A_MHTbhHOa0_1;
	wire w_dff_A_AoTVhK5r5_1;
	wire w_dff_A_QSj695yh7_1;
	wire w_dff_A_WF7BzBBr0_1;
	wire w_dff_A_15WhUGMC7_1;
	wire w_dff_A_xBOjaOlL7_1;
	wire w_dff_A_TkQwiBzn1_1;
	wire w_dff_A_L52SjsYQ4_1;
	wire w_dff_A_N2Pesr8z2_1;
	wire w_dff_A_XTCRzv6s1_1;
	wire w_dff_A_IS6nQ2ra3_1;
	wire w_dff_A_JDbvVLrP1_2;
	wire w_dff_A_vnLBKfjy6_2;
	wire w_dff_A_T7N0C8DA8_2;
	wire w_dff_A_G1CLjoIg1_2;
	wire w_dff_A_86ZiklER1_2;
	wire w_dff_A_bX3uCpoF3_2;
	wire w_dff_A_w8qgU3tT1_2;
	wire w_dff_A_Bwnsjr1H9_2;
	wire w_dff_A_La7wa7Bc6_2;
	wire w_dff_A_kHmuemLx6_2;
	wire w_dff_A_ZJlPIZyA0_2;
	wire w_dff_A_Hk6Fst9G4_2;
	wire w_dff_A_sl1auLmP0_2;
	wire w_dff_A_diD9t98R6_2;
	wire w_dff_A_Uyioptp97_2;
	wire w_dff_A_NYg3koBS9_2;
	wire w_dff_A_bT4QangZ4_2;
	wire w_dff_A_m6hxobLJ9_2;
	wire w_dff_A_mD33a3fK9_2;
	wire w_dff_A_LibtmzMl2_2;
	wire w_dff_A_xyW0CzY38_2;
	wire w_dff_A_LdmW8x0z3_2;
	wire w_dff_A_4TQbtAe49_2;
	wire w_dff_A_4kapq13Z7_2;
	wire w_dff_A_038Cfig42_2;
	wire w_dff_A_dCrUWxxP8_2;
	wire w_dff_A_GPjazOGn9_2;
	wire w_dff_A_QiMycBOG7_2;
	wire w_dff_A_zpumRBPU4_1;
	wire w_dff_A_tUyoymqM6_0;
	wire w_dff_A_leokNJoC3_0;
	wire w_dff_A_tMtAbBE44_0;
	wire w_dff_A_2zTBnVFY3_0;
	wire w_dff_A_RhfmZnRx8_0;
	wire w_dff_A_QsOMXu7T3_0;
	wire w_dff_A_cK0G9SQn9_0;
	wire w_dff_A_eKFeOMgR6_0;
	wire w_dff_A_CUrqyxfF2_0;
	wire w_dff_A_9gNR32xh3_0;
	wire w_dff_A_um0V0JMZ4_0;
	wire w_dff_A_u8FwNoFQ0_0;
	wire w_dff_A_hsJNcbhz1_0;
	wire w_dff_A_3qgpskuU3_0;
	wire w_dff_A_AOPqFoq74_0;
	wire w_dff_A_S6zvsmWW5_2;
	wire w_dff_A_qhKHZmkp2_2;
	wire w_dff_A_R5E4t7Wd7_2;
	wire w_dff_A_MGRmqino7_2;
	wire w_dff_A_GcTVFFyF2_2;
	wire w_dff_A_Tq99ZMKc7_2;
	wire w_dff_A_LJGOPbFW8_2;
	wire w_dff_A_Lbz5AVLt8_2;
	wire w_dff_A_4IbI5qIg8_2;
	wire w_dff_A_kzzigXOh3_2;
	wire w_dff_A_KvMsw2Wz1_1;
	wire w_dff_A_ABsvNh0q2_1;
	wire w_dff_A_9Ndf4BQT7_1;
	wire w_dff_A_6yGIbgJk9_1;
	wire w_dff_A_Bcdyjoly5_1;
	wire w_dff_A_jmAtlOM26_1;
	wire w_dff_A_sZMLoobE0_1;
	wire w_dff_A_OniJDID48_1;
	wire w_dff_A_cKvAUkTb6_1;
	wire w_dff_A_aX9q493N5_1;
	wire w_dff_A_hHg7xQvB7_1;
	wire w_dff_A_5H6tSYr47_1;
	wire w_dff_A_xWr7UH5Q3_1;
	wire w_dff_A_59QCt9ds9_1;
	wire w_dff_A_BO0euw167_1;
	wire w_dff_A_vBtuAjRG5_1;
	wire w_dff_A_fzWzgkzq4_1;
	wire w_dff_A_G1bb6GGQ8_1;
	wire w_dff_A_hqnH5O3V7_1;
	wire w_dff_A_XG3thPpc7_1;
	wire w_dff_A_6m7zhnEg7_1;
	wire w_dff_A_Q7TomOj72_2;
	wire w_dff_A_CKW59UZj8_2;
	wire w_dff_A_rQ78NIQ30_2;
	wire w_dff_A_ENqtAIKJ8_2;
	wire w_dff_A_l6YA0Qq68_2;
	wire w_dff_A_CgAlXiqs5_2;
	wire w_dff_A_CbNIir6s3_2;
	wire w_dff_A_6cSLp0Vr2_2;
	wire w_dff_A_Gi49wAiq8_2;
	wire w_dff_A_17q7hs9C8_2;
	wire w_dff_A_P09OghY97_2;
	wire w_dff_A_CXDKtMOS7_2;
	wire w_dff_A_HxlWNWNN4_2;
	wire w_dff_A_Gi4ay76v6_2;
	wire w_dff_A_73ILQWAl8_2;
	wire w_dff_A_RaJ5jN9j2_2;
	wire w_dff_A_GdkOIG3a5_2;
	wire w_dff_A_RVIUz57V5_2;
	wire w_dff_A_jtmbmHih5_2;
	wire w_dff_A_qDgDVAEX0_2;
	wire w_dff_A_n83Fldmf3_1;
	wire w_dff_A_7SnZt01m0_1;
	wire w_dff_A_1r6QYUXj7_1;
	wire w_dff_A_duODh0l13_1;
	wire w_dff_A_Qx5Aw0pp3_1;
	wire w_dff_A_S2krUQee6_1;
	wire w_dff_A_QHiPL11p7_1;
	wire w_dff_A_AQobxrTk8_1;
	wire w_dff_A_mBpcS1Uq1_1;
	wire w_dff_A_wfoOlIGA8_1;
	wire w_dff_A_N9vEfZbe5_1;
	wire w_dff_A_aRKS6wrS8_1;
	wire w_dff_A_iEHF2neW8_1;
	wire w_dff_A_CZMZSsPr3_1;
	wire w_dff_A_iJzWIcv50_1;
	wire w_dff_A_GCavndNK0_1;
	wire w_dff_A_cegOVNab9_1;
	wire w_dff_A_CjiMQbZv0_1;
	wire w_dff_A_EckuY08T7_2;
	wire w_dff_A_ZCFc1NNs1_2;
	wire w_dff_A_QrxlWYS79_2;
	wire w_dff_A_paxpOmvk8_2;
	wire w_dff_A_8Xwink375_2;
	wire w_dff_A_wDNAb4JQ6_2;
	wire w_dff_A_X9qoxXSa8_2;
	wire w_dff_A_MstGL8182_2;
	wire w_dff_A_yFbPnCGk3_2;
	wire w_dff_A_wo2T2kOp4_2;
	wire w_dff_A_R5JhrLx67_2;
	wire w_dff_A_Kd1woLoV1_1;
	wire w_dff_A_TL5yoWNt6_1;
	wire w_dff_A_p71EIynG9_1;
	wire w_dff_A_9FGJ1ogt3_1;
	wire w_dff_A_zyxbVRY35_1;
	wire w_dff_A_KNUNeVH45_1;
	wire w_dff_A_R4FSVQbU2_1;
	wire w_dff_A_IbRR8L6h1_1;
	wire w_dff_A_3RYyMW4v3_1;
	wire w_dff_B_vTTmgdXH3_2;
	wire w_dff_B_zUduTCUO7_2;
	wire w_dff_A_WvYQrlL30_1;
	wire w_dff_A_oxglm8aL4_1;
	wire w_dff_A_Uyau8rOH4_1;
	wire w_dff_A_iUWZmf4S8_1;
	wire w_dff_A_IQOPX7Yd0_1;
	wire w_dff_A_DSwvziJG4_1;
	wire w_dff_A_h0MFtjq21_1;
	wire w_dff_A_9yALk5ej3_1;
	wire w_dff_A_GwwbeOyA5_1;
	wire w_dff_A_5rOVFMcB6_1;
	wire w_dff_A_p6lVwuwY1_1;
	wire w_dff_A_DaDP6A9e5_1;
	wire w_dff_A_hCyIYmwG4_1;
	wire w_dff_A_cEKVsM0h0_1;
	wire w_dff_A_dTd3rY9p2_1;
	wire w_dff_A_XQXoc7ej7_1;
	wire w_dff_A_FtERhn0I3_1;
	wire w_dff_A_r7FVvO7W8_1;
	wire w_dff_A_Prm6Og5L4_1;
	wire w_dff_A_hG80psQJ5_1;
	wire w_dff_A_1jbPEVyJ8_1;
	wire w_dff_A_GUPV9wHc6_1;
	wire w_dff_A_maasZoqd6_1;
	wire w_dff_A_iSQ5fhzh9_2;
	wire w_dff_A_1zn0FW9l3_0;
	wire w_dff_A_sI0t8hvi3_0;
	wire w_dff_A_n8PzcbeJ9_0;
	wire w_dff_A_faxlmhbC2_0;
	wire w_dff_A_D5259ui21_0;
	wire w_dff_A_kDYYvRzI8_0;
	wire w_dff_A_4MzQigLh6_0;
	wire w_dff_A_BF833sLg1_0;
	wire w_dff_A_I2Ahqqac3_0;
	wire w_dff_A_wd0sOB1O0_0;
	wire w_dff_A_pnOQiB9S6_0;
	wire w_dff_A_ZjvMkhaB3_0;
	wire w_dff_A_0ZUkinzQ9_0;
	wire w_dff_A_B8nvlZ5P7_0;
	wire w_dff_A_pValhosE3_1;
	wire w_dff_A_qBUBGJnf6_1;
	wire w_dff_A_WwMkvTmg2_1;
	wire w_dff_A_0tZkGy2R5_1;
	wire w_dff_A_Q457IU110_1;
	wire w_dff_A_P1ZoAfh73_1;
	wire w_dff_A_8Bs1N5t89_1;
	wire w_dff_A_D82Fgav34_1;
	wire w_dff_A_gaZOFjBe1_1;
	wire w_dff_A_EKrQaWfW0_1;
	wire w_dff_A_kX03BD1P6_1;
	wire w_dff_A_UA9Pf4KL5_1;
	wire w_dff_A_zXcWcBZX6_1;
	wire w_dff_A_tb6fQmuU0_1;
	wire w_dff_A_q0m21wPi2_1;
	wire w_dff_A_QDiPIroo4_1;
	wire w_dff_A_PoiMz5Ac9_2;
	wire w_dff_A_JNKQLG351_2;
	wire w_dff_A_wXvvl4220_2;
	wire w_dff_A_eyUILGWx5_2;
	wire w_dff_A_ciRmbqC69_2;
	wire w_dff_A_toGPZZx61_2;
	wire w_dff_A_8BAYJSgG8_2;
	wire w_dff_A_0zVSTN7V4_2;
	wire w_dff_A_ZjiWu6AX5_2;
	wire w_dff_A_BCMNKDZn4_2;
	wire w_dff_A_y9X4lfj04_2;
	wire w_dff_A_oF5qS0QM0_2;
	wire w_dff_A_MJ2fc6d40_2;
	wire w_dff_A_QZHUGb6u4_2;
	wire w_dff_A_V1Ok5GXE1_2;
	wire w_dff_A_upmf6GZf8_2;
	wire w_dff_A_cG5jVoDi3_2;
	wire w_dff_A_JjpVs2l14_2;
	wire w_dff_A_0Zydq1sV2_2;
	wire w_dff_A_3bmgABKA0_2;
	wire w_dff_A_7LvYdvXl2_2;
	wire w_dff_A_eJwSTwYZ2_2;
	wire w_dff_A_UKG6o2On8_1;
	wire w_dff_A_FLatmz6y4_1;
	wire w_dff_A_Ofo6YQ9j5_1;
	wire w_dff_A_S7zuDv7J9_1;
	wire w_dff_A_2MDohQwi1_1;
	wire w_dff_A_OhKwQuUF8_1;
	wire w_dff_A_RXfymimW9_1;
	wire w_dff_A_6P6OGPYf9_1;
	wire w_dff_A_kcbGcgpW1_1;
	wire w_dff_A_eP5SoSc09_1;
	wire w_dff_A_9mEPYqNs0_1;
	wire w_dff_A_Oqh6KgFz0_1;
	wire w_dff_A_x0n7M0CU1_1;
	wire w_dff_A_VI9suVM74_1;
	wire w_dff_A_qhvw2oD49_1;
	wire w_dff_A_uRKIXgyP0_1;
	wire w_dff_A_1CLzg2rg9_1;
	wire w_dff_A_DdnqrwI38_1;
	wire w_dff_A_cCDNMOeN8_1;
	wire w_dff_A_ctaA7Ga85_2;
	wire w_dff_A_pvCPnmrF3_2;
	wire w_dff_A_FJqnepso1_2;
	wire w_dff_A_ZXqA7kjK0_2;
	wire w_dff_A_Sjj8KgGM0_2;
	wire w_dff_A_HVV6sDmd5_2;
	wire w_dff_A_nGmCrTM09_2;
	wire w_dff_A_iypFZ4u34_2;
	wire w_dff_A_AF0T8pOP5_2;
	wire w_dff_A_tZzpomHH7_2;
	wire w_dff_A_9twEvPVT9_2;
	wire w_dff_A_RuPJy40b7_2;
	wire w_dff_A_23j1qrul6_2;
	wire w_dff_B_2yHgIPs07_2;
	wire w_dff_B_9sooeByT0_2;
	wire w_dff_B_2NtVvx7U7_2;
	wire w_dff_B_ZxvMcgsl9_2;
	wire w_dff_B_66RmEDxR7_2;
	wire w_dff_B_2z3YppNc4_2;
	wire w_dff_B_7hBvI9OX1_2;
	wire w_dff_B_snZ0o9Go0_2;
	wire w_dff_B_Utc8l5Ed5_2;
	wire w_dff_B_NF5C1Nn97_2;
	wire w_dff_B_T2HUfdDr4_2;
	wire w_dff_B_nikbwyKM3_2;
	wire w_dff_B_Rep7RpYD2_2;
	wire w_dff_B_mPJEABN45_2;
	wire w_dff_B_28kfokIz3_2;
	wire w_dff_B_HT9O9xGS3_2;
	wire w_dff_B_Bl5IV9hL1_2;
	wire w_dff_B_exsyAiCG6_2;
	wire w_dff_B_sgULzQrm4_2;
	wire w_dff_B_wkl94Ujk6_2;
	wire w_dff_B_uJwmzMDo1_2;
	wire w_dff_B_u6C3mbq99_2;
	wire w_dff_B_X2NDuRZT2_2;
	wire w_dff_B_Tz5UtP4x1_2;
	wire w_dff_B_gBJalVQ91_2;
	wire w_dff_B_WbwCPc6t8_2;
	wire w_dff_B_ComM23HU8_2;
	wire w_dff_A_rx02fJcA4_2;
	wire w_dff_A_IjALdprk9_2;
	wire w_dff_A_Qh7WqTdm3_2;
	wire w_dff_A_sAIzt9Om2_2;
	wire w_dff_A_zjPgcxCe5_2;
	wire w_dff_A_EK5u4MGd4_2;
	wire w_dff_A_Qy0P7KGC3_2;
	wire w_dff_A_NpUXdRDf9_2;
	wire w_dff_A_U9QQQQ9q7_2;
	wire w_dff_A_o09nx3OJ9_2;
	wire w_dff_A_y4lPRZbD2_2;
	wire w_dff_A_hSUd2tAn6_2;
	wire w_dff_A_VwQ7Q4MO3_2;
	wire w_dff_A_dhOvOXiJ7_2;
	wire w_dff_A_k9OrDIyn6_2;
	wire w_dff_A_lz2J2iFq4_2;
	wire w_dff_A_X8bcnnpD2_2;
	wire w_dff_A_tgqHDiAc2_2;
	wire w_dff_A_wWrsynmd1_2;
	wire w_dff_A_isLajwhg1_2;
	wire w_dff_A_FyHF9BLE4_2;
	wire w_dff_A_xK66aRus4_2;
	wire w_dff_A_x6nZdfzX3_2;
	wire w_dff_A_sNwTwktN2_2;
	wire w_dff_A_A8BELJ2X6_0;
	wire w_dff_A_zKiWamOe3_0;
	wire w_dff_A_O5YFOKGR7_0;
	wire w_dff_A_mtujyeSZ6_0;
	wire w_dff_A_zW829UXt3_0;
	wire w_dff_A_GDujKmWD5_0;
	wire w_dff_A_wY8J6Gb31_0;
	wire w_dff_A_7KZUvj8u0_0;
	wire w_dff_A_BeQqMVqK0_0;
	wire w_dff_A_AfrDHYLP4_0;
	wire w_dff_A_JEuwzS7x6_0;
	wire w_dff_A_qjSc4dUF4_0;
	wire w_dff_A_151P5m3h8_0;
	wire w_dff_A_7k2fERvA4_0;
	wire w_dff_A_Z1q1Mqem2_0;
	wire w_dff_A_DRfSNG8T2_0;
	wire w_dff_A_kBbJ84pR7_0;
	wire w_dff_A_xRuhdLMe1_1;
	wire w_dff_A_aLpvP9LV1_1;
	wire w_dff_A_F0se0r0E0_1;
	wire w_dff_A_Csk56dO18_1;
	wire w_dff_A_troJ6RLa5_1;
	wire w_dff_A_9fKkWfc92_1;
	wire w_dff_A_26Jm6bKv9_1;
	wire w_dff_A_EsurVI7l9_1;
	wire w_dff_A_zkC8SsFR6_1;
	wire w_dff_A_1BWYzmuQ1_1;
	wire w_dff_A_UN5DTPSc9_1;
	wire w_dff_A_NW14Cpb48_1;
	wire w_dff_A_XdinJ2ua1_1;
	wire w_dff_A_596UulZT0_1;
	wire w_dff_A_4BTpAQXa4_1;
	wire w_dff_A_rVLNTSTJ6_1;
	wire w_dff_A_5W8qnzvR0_0;
	wire w_dff_A_DhSCiVOk5_0;
	wire w_dff_A_ZqmDPFpX7_0;
	wire w_dff_A_OlwTOGBO1_0;
	wire w_dff_A_3xkKmlGw6_0;
	wire w_dff_A_4Z7Y37RQ6_0;
	wire w_dff_A_2vtPyoSX7_0;
	wire w_dff_A_PIzinJ1w3_0;
	wire w_dff_A_fBhv2TTk2_0;
	wire w_dff_A_pw1HQgXf1_0;
	wire w_dff_A_bp4RaVkA5_0;
	wire w_dff_A_tkiJsETO3_0;
	wire w_dff_A_2jZ0Yaw72_0;
	wire w_dff_A_wKnrJxZZ7_0;
	wire w_dff_A_KHCyhPaf7_0;
	wire w_dff_A_g8dTMHiq0_0;
	wire w_dff_A_Cmuj7iFG0_0;
	wire w_dff_A_s01I0WgX4_0;
	wire w_dff_A_cmdd8QJ67_0;
	wire w_dff_A_7wJiYFI65_0;
	wire w_dff_A_qHkBqdhz5_0;
	wire w_dff_A_t4wnJ0ts3_0;
	wire w_dff_A_IxgCif1n3_0;
	wire w_dff_A_HWhrWMmM0_0;
	wire w_dff_A_rLl4xzb80_0;
	wire w_dff_A_36qrJKoI2_0;
	wire w_dff_A_T1lLeCux0_0;
	wire w_dff_A_66TVFEek2_1;
	wire w_dff_A_e6Tt3Oxu1_0;
	wire w_dff_A_vbjLKxae7_0;
	wire w_dff_A_3PHrQZBh9_0;
	wire w_dff_A_UD7NvugM4_0;
	wire w_dff_A_8wRcVrZn2_0;
	wire w_dff_A_GqtQunKv8_0;
	wire w_dff_A_4SX7KZ3w3_0;
	wire w_dff_A_88Cq0ZWY9_0;
	wire w_dff_A_8AS9GNjx5_0;
	wire w_dff_A_QHDwokZ27_0;
	wire w_dff_A_0vs2Z1sl0_0;
	wire w_dff_A_ZBBrLpEV9_0;
	wire w_dff_A_zbhioTiY5_0;
	wire w_dff_A_F3ynzS6p1_0;
	wire w_dff_A_i7kv418J8_0;
	wire w_dff_A_wjeJJvUX7_0;
	wire w_dff_A_991H8U6N3_0;
	wire w_dff_A_jIgKbxMV3_0;
	wire w_dff_A_DsI9Q1i31_0;
	wire w_dff_A_YgsK38Qp9_0;
	wire w_dff_A_ZNmpkZwe4_0;
	wire w_dff_A_zR3TTkFu2_0;
	wire w_dff_A_lPROXJ9D8_0;
	wire w_dff_A_Q1c3rkbg4_0;
	wire w_dff_A_UxRSzE180_0;
	wire w_dff_A_xVDouYFF1_0;
	wire w_dff_A_Kq4rLhGI3_0;
	wire w_dff_A_cOzPVBtM3_1;
	wire w_dff_A_72ZR4UTZ7_0;
	wire w_dff_A_Bf504nHY0_0;
	wire w_dff_A_f9QXljEo8_0;
	wire w_dff_A_eC9nqIBI8_0;
	wire w_dff_A_QRCuucQo4_0;
	wire w_dff_A_dsQe4pSS1_0;
	wire w_dff_A_Bb4uoTXu1_0;
	wire w_dff_A_HROEk1dt9_0;
	wire w_dff_A_XWlpIgNq2_0;
	wire w_dff_A_HE5m0u697_0;
	wire w_dff_A_PU03U1h99_0;
	wire w_dff_A_y5XCgYBi9_0;
	wire w_dff_A_X9rOq4NT7_0;
	wire w_dff_A_QjSIHy7p6_0;
	wire w_dff_A_vGBqmh7w4_0;
	wire w_dff_A_1IoinElv1_0;
	wire w_dff_A_YxVaFZGm1_0;
	wire w_dff_A_TTaP4J3h7_0;
	wire w_dff_A_0JrGIvkU7_0;
	wire w_dff_A_Povm8g0T8_0;
	wire w_dff_A_98x0DwU05_0;
	wire w_dff_A_J6FQE78K4_0;
	wire w_dff_A_c7QpQhh33_0;
	wire w_dff_A_r7UGk4pr6_0;
	wire w_dff_A_j0fGoIma0_0;
	wire w_dff_A_6ru6Hf1c0_0;
	wire w_dff_A_B6D4QjdY1_0;
	wire w_dff_A_ZBrec1Vu5_1;
	wire w_dff_A_9HjHzhb74_0;
	wire w_dff_A_0gQLt4rn2_0;
	wire w_dff_A_ZhY6jJLm8_0;
	wire w_dff_A_ZTcwPJYb6_0;
	wire w_dff_A_OmtjDjBq0_0;
	wire w_dff_A_LLOIkHnB4_0;
	wire w_dff_A_AsGV2thy5_0;
	wire w_dff_A_nNHQaBxV0_0;
	wire w_dff_A_PZ6END2h6_0;
	wire w_dff_A_NFJO4cCu4_0;
	wire w_dff_A_d7wBAC4s8_0;
	wire w_dff_A_Dcbnwu9o5_0;
	wire w_dff_A_iBrDHkMn3_0;
	wire w_dff_A_FOW0lCgf3_0;
	wire w_dff_A_geZbrlJo1_0;
	wire w_dff_A_rRuZsvsK4_0;
	wire w_dff_A_dsPzCTFW9_0;
	wire w_dff_A_9plZiwZc3_0;
	wire w_dff_A_XO8tngcP9_0;
	wire w_dff_A_LQamYGXh8_0;
	wire w_dff_A_i3kEDeyu6_0;
	wire w_dff_A_oaO3PXFu2_0;
	wire w_dff_A_HA5vElS69_0;
	wire w_dff_A_z1KxBbj12_0;
	wire w_dff_A_NEWGDjVD2_0;
	wire w_dff_A_LMxUAXnI3_0;
	wire w_dff_A_LWbmaDOx7_1;
	wire w_dff_A_G77qIhlB1_0;
	wire w_dff_A_ZH3LWzlQ5_0;
	wire w_dff_A_lFnt3W3e4_0;
	wire w_dff_A_ZA2xwnUC4_0;
	wire w_dff_A_CavUfkSL4_0;
	wire w_dff_A_ftBqPUNs2_0;
	wire w_dff_A_vMfyVpXQ3_0;
	wire w_dff_A_6bzKCMHS7_0;
	wire w_dff_A_81IYzGyB2_0;
	wire w_dff_A_iWBIU4cS1_0;
	wire w_dff_A_KpoOcQ1n0_0;
	wire w_dff_A_qGUqL9le2_0;
	wire w_dff_A_FY8epnLO2_0;
	wire w_dff_A_58mLI5xt3_0;
	wire w_dff_A_LOIpxovQ5_0;
	wire w_dff_A_U7TwF1Fc3_0;
	wire w_dff_A_anaQSJ0f6_0;
	wire w_dff_A_oc0T40gt3_0;
	wire w_dff_A_rG0LNEBt9_0;
	wire w_dff_A_vSmwMge69_0;
	wire w_dff_A_PtCPtguF5_0;
	wire w_dff_A_5qDUjCvt6_0;
	wire w_dff_A_hEjpu3F45_0;
	wire w_dff_A_Y4JP3PhZ8_0;
	wire w_dff_A_pczSir390_0;
	wire w_dff_A_0yq65Dyx6_0;
	wire w_dff_A_9M7VFoQ81_1;
	wire w_dff_A_Z1yuy3GJ8_0;
	wire w_dff_A_OJom6nUJ8_0;
	wire w_dff_A_6iUYxKgP2_0;
	wire w_dff_A_51N8aG8j0_0;
	wire w_dff_A_U51uCfT92_0;
	wire w_dff_A_wlNgaXLk5_0;
	wire w_dff_A_HJXjAIbc2_0;
	wire w_dff_A_0N9jKlA57_0;
	wire w_dff_A_Y0ccbfKC2_0;
	wire w_dff_A_OAc49W245_0;
	wire w_dff_A_GAlBH3L10_0;
	wire w_dff_A_PsPZevd36_0;
	wire w_dff_A_1WbWD7117_0;
	wire w_dff_A_pvVFRsvR6_0;
	wire w_dff_A_nqLPrIOh3_0;
	wire w_dff_A_fNSJmsjO5_0;
	wire w_dff_A_h2JhboCa1_0;
	wire w_dff_A_xI4VORAL7_0;
	wire w_dff_A_EDFjdaGP7_0;
	wire w_dff_A_cjoo9Vqa8_0;
	wire w_dff_A_sAlipV9a1_0;
	wire w_dff_A_PoJJFXU00_0;
	wire w_dff_A_cqVpYbPl9_0;
	wire w_dff_A_PzacCgIN6_0;
	wire w_dff_A_HG9QmtQO8_0;
	wire w_dff_A_wyoToT9J2_0;
	wire w_dff_A_ErVd9dvY1_1;
	wire w_dff_A_mQlTFZrd0_0;
	wire w_dff_A_6AC4U78P0_0;
	wire w_dff_A_z6lRIJMC3_0;
	wire w_dff_A_iwMok4iD9_0;
	wire w_dff_A_Mi1JnWHR1_0;
	wire w_dff_A_IMMCMqfQ5_0;
	wire w_dff_A_zvT66J7n0_0;
	wire w_dff_A_WDBcrvJJ8_0;
	wire w_dff_A_qXcma8tL2_0;
	wire w_dff_A_2fwqvAeD6_0;
	wire w_dff_A_YbE3af0v7_0;
	wire w_dff_A_doDlAHgH6_0;
	wire w_dff_A_HzYboDvG1_0;
	wire w_dff_A_iVrSmTkO0_0;
	wire w_dff_A_7E6Dxsf10_0;
	wire w_dff_A_QhCoLZ5E6_0;
	wire w_dff_A_Du10hnrC4_0;
	wire w_dff_A_VauC8AWi1_0;
	wire w_dff_A_zEDOjqZP2_0;
	wire w_dff_A_rsbtDTkc7_0;
	wire w_dff_A_OyM4Ma0l9_0;
	wire w_dff_A_WARWnHPy8_0;
	wire w_dff_A_zDAKdEI92_0;
	wire w_dff_A_tyEl8rog7_0;
	wire w_dff_A_1JraaIEI2_0;
	wire w_dff_A_k7cQgACV4_0;
	wire w_dff_A_KwFthaXT7_1;
	wire w_dff_A_oaR4YbRs8_0;
	wire w_dff_A_XZOVlZ2x5_0;
	wire w_dff_A_vnFPic539_0;
	wire w_dff_A_pkUTM2qt5_0;
	wire w_dff_A_DGSN06W86_0;
	wire w_dff_A_9iVrpYmB5_0;
	wire w_dff_A_07LJcw2a4_0;
	wire w_dff_A_APelAM7q8_0;
	wire w_dff_A_3raM8th58_0;
	wire w_dff_A_nR95UGcK1_0;
	wire w_dff_A_BYpW1t7u9_0;
	wire w_dff_A_W5GwHe6f1_0;
	wire w_dff_A_uWEDh6283_0;
	wire w_dff_A_jc1aaP861_0;
	wire w_dff_A_YAC5Br0L1_0;
	wire w_dff_A_8wLp2KdT5_0;
	wire w_dff_A_fNAlytst3_0;
	wire w_dff_A_gUrXzxCQ2_0;
	wire w_dff_A_EahSMhEL4_0;
	wire w_dff_A_zDoResQT0_0;
	wire w_dff_A_VxDRyiV39_0;
	wire w_dff_A_4zCX84kg7_0;
	wire w_dff_A_rT6o1Hc34_0;
	wire w_dff_A_GvWe8BoL4_0;
	wire w_dff_A_8cwhzSJf0_0;
	wire w_dff_A_GPIgC0h77_0;
	wire w_dff_A_IfMxj8Bd5_1;
	wire w_dff_A_KebsTOnD7_0;
	wire w_dff_A_wuINnOS62_0;
	wire w_dff_A_Ddm5GtEf5_0;
	wire w_dff_A_drb3WDHp9_0;
	wire w_dff_A_i1ZIJ60J7_0;
	wire w_dff_A_Ag1qUUy20_0;
	wire w_dff_A_BQ6YV57r3_0;
	wire w_dff_A_3LYRkJKU4_0;
	wire w_dff_A_Po1kKwBA1_0;
	wire w_dff_A_Rvwbnp683_0;
	wire w_dff_A_tlEXmYvm3_0;
	wire w_dff_A_Db40u4xW9_0;
	wire w_dff_A_udAuWS4M4_0;
	wire w_dff_A_DyuwXitL1_0;
	wire w_dff_A_eOu8vCrx4_0;
	wire w_dff_A_W6TKeSxX6_0;
	wire w_dff_A_giOXoufo4_0;
	wire w_dff_A_Q4P7yEMe0_0;
	wire w_dff_A_fR8qyBTb9_0;
	wire w_dff_A_idmUBCqj7_0;
	wire w_dff_A_AGAV1MQv2_0;
	wire w_dff_A_oT4cZ4Rn8_0;
	wire w_dff_A_wtVe6uhD5_0;
	wire w_dff_A_LGFMivYR5_0;
	wire w_dff_A_GmVoLtqC1_0;
	wire w_dff_A_PeTVeBSe3_0;
	wire w_dff_A_O2Tzkydk6_1;
	wire w_dff_A_O45zSPP70_0;
	wire w_dff_A_5EwzfoE47_0;
	wire w_dff_A_RHTKb1qR8_0;
	wire w_dff_A_oki8ZLtg1_0;
	wire w_dff_A_kJXcSCHo4_0;
	wire w_dff_A_UpkQRyx18_0;
	wire w_dff_A_woYCIYZu2_0;
	wire w_dff_A_gwBPAcOl9_0;
	wire w_dff_A_sfWtZCMB3_0;
	wire w_dff_A_cDUBZR605_0;
	wire w_dff_A_In1RWngt4_0;
	wire w_dff_A_VgIREoql1_0;
	wire w_dff_A_GbkU81ud2_0;
	wire w_dff_A_D4D9Vdl01_0;
	wire w_dff_A_me2yGOhm7_0;
	wire w_dff_A_fYmPdThD6_0;
	wire w_dff_A_TxJv3yc40_0;
	wire w_dff_A_a2sgY9XB8_0;
	wire w_dff_A_WzWtHhzQ2_0;
	wire w_dff_A_QRUzJfO15_0;
	wire w_dff_A_N1g9twN48_0;
	wire w_dff_A_GdTvfgpX7_0;
	wire w_dff_A_51vZNVEY9_0;
	wire w_dff_A_Dc3Yfork6_0;
	wire w_dff_A_zuz5rhrO4_0;
	wire w_dff_A_5RxE9owP5_0;
	wire w_dff_A_UzBVPGlV5_1;
	wire w_dff_A_ON8NVNbY4_0;
	wire w_dff_A_7qYTwD7H3_0;
	wire w_dff_A_8ZM378CX9_0;
	wire w_dff_A_kLEJLwSF4_0;
	wire w_dff_A_ZoBkBnAn7_0;
	wire w_dff_A_kAmwv8Rx0_0;
	wire w_dff_A_YnusH0PG2_0;
	wire w_dff_A_AJ24Mydj1_0;
	wire w_dff_A_Gcr3rltz5_0;
	wire w_dff_A_tRN5YyAv9_0;
	wire w_dff_A_Pp5CziCW6_0;
	wire w_dff_A_GzGihGTs2_0;
	wire w_dff_A_RWC9CCZz8_0;
	wire w_dff_A_qnxKGygg9_0;
	wire w_dff_A_IooDKUNC8_0;
	wire w_dff_A_TTKMYcMD7_0;
	wire w_dff_A_fkCUzq2r3_0;
	wire w_dff_A_fIkyIvQl3_0;
	wire w_dff_A_FxY7VJgL9_0;
	wire w_dff_A_MvJeQUfX4_0;
	wire w_dff_A_wqrGHSH05_0;
	wire w_dff_A_EJrXNefK2_0;
	wire w_dff_A_5VVAb7Yb0_0;
	wire w_dff_A_SW2Rxth20_0;
	wire w_dff_A_67BtqV7a7_0;
	wire w_dff_A_qIYPYWs10_0;
	wire w_dff_A_H84LiIAI2_1;
	wire w_dff_A_klJf9GTN0_0;
	wire w_dff_A_dLa3TJ7i4_0;
	wire w_dff_A_us5feTLe5_0;
	wire w_dff_A_PcnvCYzO8_0;
	wire w_dff_A_FmxEbqEg9_0;
	wire w_dff_A_kNP6ynXm5_0;
	wire w_dff_A_jC3WmOaw2_0;
	wire w_dff_A_BewFZWr49_0;
	wire w_dff_A_fVUUv8TZ4_0;
	wire w_dff_A_xqlq3lMV8_0;
	wire w_dff_A_d2VvDoEr3_0;
	wire w_dff_A_mKk4ipCh2_0;
	wire w_dff_A_xvkl5pjR3_0;
	wire w_dff_A_A885zRif6_0;
	wire w_dff_A_xoW5Fo8I8_0;
	wire w_dff_A_8xd8EdF42_0;
	wire w_dff_A_LzVFpbsl9_0;
	wire w_dff_A_slUyfZHg6_0;
	wire w_dff_A_DqBZnaXz4_0;
	wire w_dff_A_YoCQdpSa6_0;
	wire w_dff_A_KkuORzXV5_0;
	wire w_dff_A_azCJmzeU4_0;
	wire w_dff_A_6rjkUue98_0;
	wire w_dff_A_UGrUCVG39_0;
	wire w_dff_A_Di0Y2KWU5_0;
	wire w_dff_A_zJhJj7xq5_0;
	wire w_dff_A_PGzCSuv27_2;
	wire w_dff_A_nbzROnjq4_0;
	wire w_dff_A_31hQn1uG8_0;
	wire w_dff_A_emxNW8uW2_0;
	wire w_dff_A_xJvEIRen0_0;
	wire w_dff_A_7tKrWlig1_0;
	wire w_dff_A_iHYwScAp3_0;
	wire w_dff_A_FVq1fI5g5_0;
	wire w_dff_A_nhzoLx5Y0_0;
	wire w_dff_A_V4GACXBn5_0;
	wire w_dff_A_lSlGTfPR1_0;
	wire w_dff_A_ZjRbpGAA7_0;
	wire w_dff_A_I9jIwkzI9_0;
	wire w_dff_A_RKvvTUuK4_0;
	wire w_dff_A_q9XvF3KC9_0;
	wire w_dff_A_9LmIJdwi9_0;
	wire w_dff_A_v4j9H0yR1_0;
	wire w_dff_A_yUNbqcnn7_0;
	wire w_dff_A_saO0hVg49_0;
	wire w_dff_A_eX9IBP8q6_0;
	wire w_dff_A_G10u59Ef6_0;
	wire w_dff_A_7H2BZrwj8_0;
	wire w_dff_A_7x0Peckt6_0;
	wire w_dff_A_RzZRL4ze5_0;
	wire w_dff_A_rEvuMfh77_0;
	wire w_dff_A_NbQtXbDt9_0;
	wire w_dff_A_rjdsfxNx9_0;
	wire w_dff_A_hnSczvAh8_1;
	wire w_dff_A_Nbs4hPpN7_0;
	wire w_dff_A_dO1vHYcD4_0;
	wire w_dff_A_7fmWQpVy2_0;
	wire w_dff_A_SRUYm03Y0_0;
	wire w_dff_A_6fz4yv274_0;
	wire w_dff_A_Vo3Rhqdv9_0;
	wire w_dff_A_AsIlTvda8_0;
	wire w_dff_A_QkjBoflG7_0;
	wire w_dff_A_FNHLVngw2_0;
	wire w_dff_A_wysyuxlY7_0;
	wire w_dff_A_Bda6igyv2_0;
	wire w_dff_A_e0DYm3nv3_0;
	wire w_dff_A_dKlb3NNO0_0;
	wire w_dff_A_GuIx3jf61_0;
	wire w_dff_A_e25GyWQi9_0;
	wire w_dff_A_EeSk23ug7_0;
	wire w_dff_A_p5YU2Hlm6_0;
	wire w_dff_A_ZsExShIw2_0;
	wire w_dff_A_crsdc2Su0_0;
	wire w_dff_A_D10H6jgb4_0;
	wire w_dff_A_4gOFM9PK3_0;
	wire w_dff_A_iVGrjTjY9_0;
	wire w_dff_A_4fJQIBYF9_0;
	wire w_dff_A_cPBR0n1u7_0;
	wire w_dff_A_v65CSxwt7_0;
	wire w_dff_A_jlREcNb64_0;
	wire w_dff_A_E78jADKM5_1;
	wire w_dff_A_Os1MnMJ39_0;
	wire w_dff_A_TGsgyyYC2_0;
	wire w_dff_A_PjcRjUHK5_0;
	wire w_dff_A_Cxr7ye9u0_0;
	wire w_dff_A_oNqNQdg82_0;
	wire w_dff_A_9dSNBXjp7_0;
	wire w_dff_A_Ow9KclPc6_0;
	wire w_dff_A_vwhwAJIg3_0;
	wire w_dff_A_L0eOgLgU8_0;
	wire w_dff_A_l5MQNVHG6_0;
	wire w_dff_A_4Y9iyfRX8_0;
	wire w_dff_A_LRLQrrPQ7_0;
	wire w_dff_A_IyvFLNBx6_0;
	wire w_dff_A_HHMKFOdI6_0;
	wire w_dff_A_3KZgfooQ1_0;
	wire w_dff_A_v3IqwvLO4_0;
	wire w_dff_A_Sopqd15x4_0;
	wire w_dff_A_SjvWJzT00_0;
	wire w_dff_A_DNR58lFv5_0;
	wire w_dff_A_rOMVEJYf4_0;
	wire w_dff_A_CjUiSqz76_0;
	wire w_dff_A_U74x9EmH6_0;
	wire w_dff_A_yYU3lUVb7_0;
	wire w_dff_A_kucTH1T92_0;
	wire w_dff_A_5ygJ0C591_0;
	wire w_dff_A_nqMgHf3K7_0;
	wire w_dff_A_AVwe8LZD9_1;
	wire w_dff_A_PO7tgq5D9_0;
	wire w_dff_A_8MCDdNcp8_0;
	wire w_dff_A_cmQHrnNI5_0;
	wire w_dff_A_5PdJUxCH0_0;
	wire w_dff_A_9WfNcnOA4_0;
	wire w_dff_A_6UlGFyej0_0;
	wire w_dff_A_IzSs48DS6_0;
	wire w_dff_A_nyvPgYcF2_0;
	wire w_dff_A_teiwgbjW7_0;
	wire w_dff_A_KGjswTrX2_0;
	wire w_dff_A_i2u3Glm31_0;
	wire w_dff_A_XLqpSjFl1_0;
	wire w_dff_A_UcAqKqU75_0;
	wire w_dff_A_cp0D2UbL9_0;
	wire w_dff_A_1BBBmYvz5_0;
	wire w_dff_A_jCbprpTt4_0;
	wire w_dff_A_jvOE0Bcl4_0;
	wire w_dff_A_3Hmrvuz22_0;
	wire w_dff_A_mrvFK7Rw6_0;
	wire w_dff_A_gFFJRjsn5_0;
	wire w_dff_A_gCupuTys4_0;
	wire w_dff_A_hWfQPs7a0_0;
	wire w_dff_A_TxPodgNl0_0;
	wire w_dff_A_QFyiUs6Q1_0;
	wire w_dff_A_EAuEEzF05_0;
	wire w_dff_A_xp1vCgnp3_0;
	wire w_dff_A_8yW8rYSC0_1;
	wire w_dff_A_jWaUtTT72_0;
	wire w_dff_A_d8CCqeeI9_0;
	wire w_dff_A_7ZjhNA046_0;
	wire w_dff_A_cYXe9Txc3_0;
	wire w_dff_A_5zEpCGD84_0;
	wire w_dff_A_SrS0fT2L4_0;
	wire w_dff_A_CXkKXAno0_0;
	wire w_dff_A_OFEwH6rW2_0;
	wire w_dff_A_MmHuy6gC5_0;
	wire w_dff_A_YaAtkiWq9_0;
	wire w_dff_A_Ww66n3773_0;
	wire w_dff_A_SUUo5uWi6_0;
	wire w_dff_A_M7kAZ2C54_0;
	wire w_dff_A_9D3l8rqA9_0;
	wire w_dff_A_ZAOREYlY3_0;
	wire w_dff_A_dQvkqOqn5_0;
	wire w_dff_A_AjiYy8BX4_0;
	wire w_dff_A_KLBflqsX4_0;
	wire w_dff_A_SsSlhH227_0;
	wire w_dff_A_7uxBLpPp4_0;
	wire w_dff_A_CObSADYm1_0;
	wire w_dff_A_WIv7iNS84_0;
	wire w_dff_A_iSoCOx0I5_0;
	wire w_dff_A_lRdT4CJ46_0;
	wire w_dff_A_ekRwoShX9_0;
	wire w_dff_A_5JxwWsO02_0;
	wire w_dff_A_il5gzRQ12_2;
	wire w_dff_A_riEweXVy7_0;
	wire w_dff_A_JkSreVU53_0;
	wire w_dff_A_5hPsmtub3_0;
	wire w_dff_A_lc3etMdM7_0;
	wire w_dff_A_eIeDO3ks3_0;
	wire w_dff_A_jIV2dcNj9_0;
	wire w_dff_A_rTs8NITW9_0;
	wire w_dff_A_n4bOUqh09_0;
	wire w_dff_A_ytIRBICk7_0;
	wire w_dff_A_7Ptvir2R4_0;
	wire w_dff_A_h0wYJW9n1_0;
	wire w_dff_A_Mxj305Ms9_0;
	wire w_dff_A_wlrlNyfu2_0;
	wire w_dff_A_jxiveFpg2_0;
	wire w_dff_A_W1S3G9PT5_0;
	wire w_dff_A_e1JTv2eI4_0;
	wire w_dff_A_zJMi3bZE7_0;
	wire w_dff_A_ZLbLw1AG4_0;
	wire w_dff_A_tRbkvvAZ2_0;
	wire w_dff_A_HGapMj9y7_0;
	wire w_dff_A_ih1Xr53m3_0;
	wire w_dff_A_IuEaUu7G4_0;
	wire w_dff_A_OUk7o9UW8_0;
	wire w_dff_A_OUkKcXKL4_0;
	wire w_dff_A_2XUhHR2f1_0;
	wire w_dff_A_QWhXvLgw5_0;
	wire w_dff_A_5yZAzLY28_2;
	wire w_dff_A_tUbXQn0z4_0;
	wire w_dff_A_fz4Jpv666_0;
	wire w_dff_A_8nazHNcJ1_0;
	wire w_dff_A_uhe5p8Mq8_0;
	wire w_dff_A_Tkv499YQ4_0;
	wire w_dff_A_5olupmWL9_0;
	wire w_dff_A_M2ax1Wdn6_0;
	wire w_dff_A_TzNUu3ZK6_0;
	wire w_dff_A_wav0QNfw5_0;
	wire w_dff_A_ulKNR54U8_0;
	wire w_dff_A_7cjmnhhj8_0;
	wire w_dff_A_wzXXIedh6_0;
	wire w_dff_A_2ojMxaAV4_0;
	wire w_dff_A_mwMcFTOK1_0;
	wire w_dff_A_PoDZDGgX1_0;
	wire w_dff_A_stgsCdxf9_0;
	wire w_dff_A_5dYTDES71_0;
	wire w_dff_A_XDuiwhjT6_0;
	wire w_dff_A_xV9CNt115_0;
	wire w_dff_A_0LnJw27W4_0;
	wire w_dff_A_G1G1MDan4_0;
	wire w_dff_A_7TpO1Pdn4_0;
	wire w_dff_A_g0FEQjEd5_0;
	wire w_dff_A_xZlzbVAn2_0;
	wire w_dff_A_HI1Rh4ot5_0;
	wire w_dff_A_Dfh0sref6_2;
	wire w_dff_A_xwcyPH0a3_0;
	wire w_dff_A_pSo1dmi77_0;
	wire w_dff_A_DE5Y2rea6_0;
	wire w_dff_A_IkKvnjdu1_0;
	wire w_dff_A_zaEoPNvZ5_0;
	wire w_dff_A_U0d9brpo2_0;
	wire w_dff_A_pPlzUs7g2_0;
	wire w_dff_A_9jHMRoOV9_0;
	wire w_dff_A_YVRK1qKE8_0;
	wire w_dff_A_Oyf7yWf86_0;
	wire w_dff_A_7QbbRmnw9_0;
	wire w_dff_A_HPGJIieo8_0;
	wire w_dff_A_5BKg6cgW9_0;
	wire w_dff_A_x8z88Exm7_0;
	wire w_dff_A_gsCFFxp63_0;
	wire w_dff_A_tHM9M5NA1_0;
	wire w_dff_A_1SOcq7Q70_0;
	wire w_dff_A_S2q6Y5NH2_0;
	wire w_dff_A_IdBpOYNS3_0;
	wire w_dff_A_ROCzrkRF2_0;
	wire w_dff_A_QPo5Ne8z2_0;
	wire w_dff_A_7u2g0qVo5_0;
	wire w_dff_A_ocCrRWin3_0;
	wire w_dff_A_FrZTDCMc0_0;
	wire w_dff_A_WsxsxKl22_0;
	wire w_dff_A_9IakLXyU2_1;
	wire w_dff_A_rufGJAmd1_0;
	wire w_dff_A_QmbBvWQC0_0;
	wire w_dff_A_keuBOLpZ7_0;
	wire w_dff_A_z2hslrWB4_0;
	wire w_dff_A_RSMFuCRy1_0;
	wire w_dff_A_63x1gn8F8_0;
	wire w_dff_A_MuA5trTl3_0;
	wire w_dff_A_RHLYyt9m0_0;
	wire w_dff_A_hVrvFaWl3_0;
	wire w_dff_A_zJA8MhWX4_0;
	wire w_dff_A_pmT97wB52_0;
	wire w_dff_A_reTcRdcR2_0;
	wire w_dff_A_0fu0XvWa2_0;
	wire w_dff_A_sXXYdx8N5_0;
	wire w_dff_A_y8muQaPw3_0;
	wire w_dff_A_bel5rW7I8_0;
	wire w_dff_A_vL1ZCH203_0;
	wire w_dff_A_o40Ra72I2_0;
	wire w_dff_A_VL8Ea4yE8_0;
	wire w_dff_A_S5lDYPbk5_0;
	wire w_dff_A_NiYBZsHm1_0;
	wire w_dff_A_HC3Dwmbt3_0;
	wire w_dff_A_d6EH0yu26_0;
	wire w_dff_A_MORjDeJV8_0;
	wire w_dff_A_w8v0m3Q02_0;
	wire w_dff_A_7IidBGnj0_1;
	wire w_dff_A_4LFar5BP2_0;
	wire w_dff_A_4MZBsiiP3_0;
	wire w_dff_A_6GtuHvx63_0;
	wire w_dff_A_NozBF5TA0_0;
	wire w_dff_A_6bIEeuAb8_0;
	wire w_dff_A_MRTMuoUf8_0;
	wire w_dff_A_kJ6pB0zZ7_0;
	wire w_dff_A_zdH2Qkq25_0;
	wire w_dff_A_W2HfM4Lo4_0;
	wire w_dff_A_y4xyVCHZ3_0;
	wire w_dff_A_F34MBWH74_0;
	wire w_dff_A_71TPG1et7_0;
	wire w_dff_A_oLgXCcvY8_0;
	wire w_dff_A_zoFyNcDR9_0;
	wire w_dff_A_VkvV2lve3_0;
	wire w_dff_A_pb3KQtoy4_0;
	wire w_dff_A_HxOIOknW6_0;
	wire w_dff_A_nPf0dmm79_0;
	wire w_dff_A_Ae5euWha8_0;
	wire w_dff_A_kjlEW1Um4_0;
	wire w_dff_A_aEHGnoD38_0;
	wire w_dff_A_x2BWPgim7_0;
	wire w_dff_A_54R3MjDQ5_0;
	wire w_dff_A_2c6SKHDE7_0;
	wire w_dff_A_b28cF2pe2_0;
	wire w_dff_A_jchro18i2_0;
	wire w_dff_A_zHRMXs3k8_0;
	wire w_dff_A_hGDXCrDc6_1;
	wire w_dff_A_7iFwTMbE4_0;
	wire w_dff_A_pweeR05v0_0;
	wire w_dff_A_jsl0Mbs59_0;
	wire w_dff_A_MlmfdpkD6_0;
	wire w_dff_A_VzBw1px09_0;
	wire w_dff_A_6UL5Hx0P9_0;
	wire w_dff_A_wIHqwPWr9_0;
	wire w_dff_A_k9YT6nXx2_0;
	wire w_dff_A_5xY0XIJW0_0;
	wire w_dff_A_XnNjdOzZ6_0;
	wire w_dff_A_Se769BEq1_0;
	wire w_dff_A_ddGZYwbp8_0;
	wire w_dff_A_MSemvxeP2_0;
	wire w_dff_A_Kd6IDemI2_0;
	wire w_dff_A_PJCISWQ25_0;
	wire w_dff_A_Yr6uya6r5_0;
	wire w_dff_A_tmzvb0Nv3_0;
	wire w_dff_A_09sHDbOn8_0;
	wire w_dff_A_u5TMods47_0;
	wire w_dff_A_EKsT2u6v4_0;
	wire w_dff_A_6XqmmfcU9_0;
	wire w_dff_A_8l1yDHw52_0;
	wire w_dff_A_laH7v5ii6_0;
	wire w_dff_A_xgiFmAmt4_0;
	wire w_dff_A_SFt0XsSv2_0;
	wire w_dff_A_pmSOYl6a7_0;
	wire w_dff_A_vTi1v3ik7_0;
	wire w_dff_A_7dsw62mq4_1;
	wire w_dff_A_MuunuXcW0_0;
	wire w_dff_A_5vCTJySf5_0;
	wire w_dff_A_RYOJbis28_0;
	wire w_dff_A_MtY4ga2x0_0;
	wire w_dff_A_CJz1oVBS4_0;
	wire w_dff_A_bwPvtujk4_0;
	wire w_dff_A_lpXRc5bz2_0;
	wire w_dff_A_zfnB1HR61_0;
	wire w_dff_A_y3R5ZmfI6_0;
	wire w_dff_A_7qg4YaXB4_0;
	wire w_dff_A_HkNL83gj2_0;
	wire w_dff_A_Pkhy5hB22_0;
	wire w_dff_A_FC257lGZ0_0;
	wire w_dff_A_lsJRvMu18_0;
	wire w_dff_A_QvDMxXil1_0;
	wire w_dff_A_HNrVC0ug4_0;
	wire w_dff_A_gFdG6EaB9_0;
	wire w_dff_A_oKaXlgHz7_0;
	wire w_dff_A_NHR5rBU29_0;
	wire w_dff_A_2Bodj7jw8_0;
	wire w_dff_A_UW1p0P4r1_0;
	wire w_dff_A_8WY8intS6_0;
	wire w_dff_A_ZFGF9ZDk7_0;
	wire w_dff_A_3LOIkVtV0_0;
	wire w_dff_A_POEFWCQU0_0;
	wire w_dff_A_4DCfUm7D8_0;
	wire w_dff_A_8xI66C5M5_0;
	wire w_dff_A_c0W5v6CF5_1;
	wire w_dff_A_r5lRUBnq9_0;
	wire w_dff_A_kRSyerpV8_0;
	wire w_dff_A_mX1pyvFx8_0;
	wire w_dff_A_sTQLXnPG7_0;
	wire w_dff_A_RkEw0W1K6_0;
	wire w_dff_A_MD48YDDH5_0;
	wire w_dff_A_YmgMDCs35_0;
	wire w_dff_A_xPJJ0fCl7_0;
	wire w_dff_A_sz8RdjQS9_0;
	wire w_dff_A_qlyVixaW7_0;
	wire w_dff_A_iuztysXN0_0;
	wire w_dff_A_1ZpdAtcZ0_0;
	wire w_dff_A_cwRqYzhP6_0;
	wire w_dff_A_sEOzjlcf1_0;
	wire w_dff_A_mdxj7SA12_0;
	wire w_dff_A_St3EwTge7_0;
	wire w_dff_A_nox2nXZF0_0;
	wire w_dff_A_rsseIDFd5_0;
	wire w_dff_A_1dzeVR4x5_0;
	wire w_dff_A_4Rx18E6h1_0;
	wire w_dff_A_MYdC1wls7_0;
	wire w_dff_A_ABVQdonB3_0;
	wire w_dff_A_vGTmAkVD5_0;
	wire w_dff_A_P0VDaHoj4_0;
	wire w_dff_A_P1BRk2kJ4_0;
	wire w_dff_A_IffsPDLL1_0;
	wire w_dff_A_RqoeCGpI4_0;
	wire w_dff_A_acyZRsoC4_1;
	wire w_dff_A_HnbLRBsH4_0;
	wire w_dff_A_fR0Abpyz4_0;
	wire w_dff_A_eZWlfAxR4_0;
	wire w_dff_A_xjFOEtOy0_0;
	wire w_dff_A_zcA8IKaL5_0;
	wire w_dff_A_guublbGq9_0;
	wire w_dff_A_DHNFzFUI5_0;
	wire w_dff_A_WeLGNQIq5_0;
	wire w_dff_A_9W0MtKpL7_0;
	wire w_dff_A_jdrfZO7y6_0;
	wire w_dff_A_VRDWPNtr4_0;
	wire w_dff_A_LINeIFbt8_0;
	wire w_dff_A_AU7ahig87_0;
	wire w_dff_A_dJl9E4s11_0;
	wire w_dff_A_HBuQM9BI7_0;
	wire w_dff_A_C7tQtGoP0_0;
	wire w_dff_A_3PSg393z5_0;
	wire w_dff_A_QdgffaEX3_0;
	wire w_dff_A_CK0mp0d94_0;
	wire w_dff_A_Qw0w5TUn9_0;
	wire w_dff_A_4K2NvvMu6_0;
	wire w_dff_A_iomx5FVG3_0;
	wire w_dff_A_BYYqPllx1_0;
	wire w_dff_A_jO9zTWys7_0;
	wire w_dff_A_8sxygSq53_0;
	wire w_dff_A_BekpnsSZ5_0;
	wire w_dff_A_yTo56sWa6_0;
	wire w_dff_A_b5bppP9C3_1;
	wire w_dff_A_hnE3BRfa8_0;
	wire w_dff_A_czA4SQ235_0;
	wire w_dff_A_r37FywQz6_0;
	wire w_dff_A_ZyjzyN5B5_0;
	wire w_dff_A_DK3WwJLG1_0;
	wire w_dff_A_mg0rV9i28_0;
	wire w_dff_A_H1y6fXa81_0;
	wire w_dff_A_baiwRXhO1_0;
	wire w_dff_A_v9BqxDiH3_0;
	wire w_dff_A_JkIV7ZTq8_0;
	wire w_dff_A_zqlpA7yf2_0;
	wire w_dff_A_q2lKCze97_0;
	wire w_dff_A_MsLvlfxG9_0;
	wire w_dff_A_XmmkHZng5_0;
	wire w_dff_A_TFyeyPa05_0;
	wire w_dff_A_AcrGSD6c7_0;
	wire w_dff_A_Io1XcflI7_0;
	wire w_dff_A_2rpTxKuA7_0;
	wire w_dff_A_ZU6jxPRt4_0;
	wire w_dff_A_C80ll9O55_0;
	wire w_dff_A_WtOeLjFY5_0;
	wire w_dff_A_EBSmERs53_0;
	wire w_dff_A_R89C3gym6_0;
	wire w_dff_A_Up7ZdmrK2_0;
	wire w_dff_A_DWSKUaut1_0;
	wire w_dff_A_bClPVLyy4_0;
	wire w_dff_A_Cg0ajXrl8_2;
	wire w_dff_A_geKvccbu1_0;
	wire w_dff_A_N6XWPsdF4_0;
	wire w_dff_A_0rwvwVbQ9_0;
	wire w_dff_A_beL712qd1_0;
	wire w_dff_A_i8O7E6XR2_0;
	wire w_dff_A_JqarZ9RO6_0;
	wire w_dff_A_NOqzOnpU8_0;
	wire w_dff_A_KSvOr7C56_0;
	wire w_dff_A_HB9qGMTO4_0;
	wire w_dff_A_Nwewo1uX4_0;
	wire w_dff_A_epYu035e1_0;
	wire w_dff_A_0MoJMuhU0_0;
	wire w_dff_A_FUjHRh7t6_0;
	wire w_dff_A_6tA5NXI79_0;
	wire w_dff_A_j8AT1bTg5_0;
	wire w_dff_A_JUN2CzMo0_0;
	wire w_dff_A_KyawlIOu0_0;
	wire w_dff_A_zTdIvZ7q8_0;
	wire w_dff_A_vYhjTbvR1_0;
	wire w_dff_A_522ZjSav3_0;
	wire w_dff_A_yvvkBSnw3_0;
	wire w_dff_A_App9HfCg7_0;
	wire w_dff_A_5cR1rmsk3_0;
	wire w_dff_A_UkXn478t6_0;
	wire w_dff_A_a0LYu7n60_2;
	wire w_dff_A_ZeXevlTk5_0;
	wire w_dff_A_WDmciOda7_0;
	wire w_dff_A_WrQ06h0i6_0;
	wire w_dff_A_zsZpcWy06_0;
	wire w_dff_A_JXiXryOx2_0;
	wire w_dff_A_e3mYZuAI1_0;
	wire w_dff_A_MPf1c4C05_0;
	wire w_dff_A_XhAf601Y5_0;
	wire w_dff_A_3qWMNiSy2_0;
	wire w_dff_A_cczxyAGQ8_0;
	wire w_dff_A_cxV0sJJm4_0;
	wire w_dff_A_svYmSWiN7_0;
	wire w_dff_A_WbyHGIz05_0;
	wire w_dff_A_SIkVC4Oc5_0;
	wire w_dff_A_HiKZrVz16_0;
	wire w_dff_A_ZtkjIz6t9_0;
	wire w_dff_A_D1ehCP2g4_0;
	wire w_dff_A_19mRsXm90_0;
	wire w_dff_A_zcgssLyH6_0;
	wire w_dff_A_Y6WorKqY9_0;
	wire w_dff_A_WZUdXUac6_0;
	wire w_dff_A_BVHaAflh5_0;
	wire w_dff_A_9OeQf4eb6_0;
	wire w_dff_A_8tyub3pi3_0;
	wire w_dff_A_LqIS8KAc4_0;
	wire w_dff_A_4QLAB4kJ6_1;
	wire w_dff_A_CZMGzdzz1_0;
	wire w_dff_A_Ygeuxq6F1_0;
	wire w_dff_A_z1ji51ux9_0;
	wire w_dff_A_PyjhS6S69_0;
	wire w_dff_A_teiiGtEp3_0;
	wire w_dff_A_HYOg3Bkv0_0;
	wire w_dff_A_bSe9Pnpw0_0;
	wire w_dff_A_uVOTm3Ko8_0;
	wire w_dff_A_qFqMhNkT7_0;
	wire w_dff_A_IBqmQwFT7_0;
	wire w_dff_A_0TW2eqjN3_0;
	wire w_dff_A_JyQeqs1D0_0;
	wire w_dff_A_sZKe8kQL4_0;
	wire w_dff_A_ODDK0O692_0;
	wire w_dff_A_GD1Y1epJ9_0;
	wire w_dff_A_3d8b4sE41_0;
	wire w_dff_A_ul2CZcZb9_0;
	wire w_dff_A_Z6eb98ke2_0;
	wire w_dff_A_sxTzbnvi1_0;
	wire w_dff_A_ldl9McF27_0;
	wire w_dff_A_OmZtZWER0_0;
	wire w_dff_A_xunTitrv4_0;
	wire w_dff_A_qnVCCIDy9_0;
	wire w_dff_A_wsa53kUS7_0;
	wire w_dff_A_t9wlPRPO2_0;
	wire w_dff_A_77SON5gz3_0;
	wire w_dff_A_bPKViaZU8_0;
	wire w_dff_A_5y0biOwJ6_1;
	wire w_dff_A_CuP3HU3H8_0;
	wire w_dff_A_6wgO6idh6_0;
	wire w_dff_A_77yPZ8fE1_0;
	wire w_dff_A_33yENelA7_0;
	wire w_dff_A_8hleZckD4_0;
	wire w_dff_A_f6suGJYz6_0;
	wire w_dff_A_kY1TDHTo0_0;
	wire w_dff_A_Wja7P7eQ7_0;
	wire w_dff_A_p9zFzQ8H6_0;
	wire w_dff_A_YoR81gSB6_0;
	wire w_dff_A_wp3MD9zv8_0;
	wire w_dff_A_udm87nCJ5_0;
	wire w_dff_A_2c66gJNO3_0;
	wire w_dff_A_0pbHLEuH4_0;
	wire w_dff_A_u9PwAwCX0_0;
	wire w_dff_A_5syXSLwY7_0;
	wire w_dff_A_Tx9q6x1D7_0;
	wire w_dff_A_orBuZSoy1_0;
	wire w_dff_A_NvLUnGYQ0_0;
	wire w_dff_A_N7DRbtX59_0;
	wire w_dff_A_qc7W0tKd1_0;
	wire w_dff_A_dXj9QJZS2_0;
	wire w_dff_A_1MMrnxhe8_0;
	wire w_dff_A_30e7C8yc1_0;
	wire w_dff_A_BdDXYNqW2_0;
	wire w_dff_A_JCS8MAGB3_0;
	wire w_dff_A_8dGDKZ2C3_0;
	wire w_dff_A_S9WcFqMu6_1;
	wire w_dff_A_9C07X2mv9_0;
	wire w_dff_A_Wu1mNrHt8_0;
	wire w_dff_A_qdln7FBI9_0;
	wire w_dff_A_Hr9sj9h72_0;
	wire w_dff_A_FScjYHSM4_0;
	wire w_dff_A_TIFR0Jk78_0;
	wire w_dff_A_LCTuYaip1_0;
	wire w_dff_A_ZlS9lcro7_0;
	wire w_dff_A_6kbjqBFj3_0;
	wire w_dff_A_rPwsrr137_0;
	wire w_dff_A_qft6sav31_0;
	wire w_dff_A_izZgnMVf1_0;
	wire w_dff_A_OIyUcUvC0_0;
	wire w_dff_A_KIQgKCiW7_0;
	wire w_dff_A_vSzyXNyz4_0;
	wire w_dff_A_6idpLyrK4_0;
	wire w_dff_A_aQbxkq9u8_0;
	wire w_dff_A_FMX48Gvb7_0;
	wire w_dff_A_fAaUdg9x1_0;
	wire w_dff_A_hN3egfdk4_0;
	wire w_dff_A_5Elq8oQI6_0;
	wire w_dff_A_HKzzsOWF6_0;
	wire w_dff_A_dKdYD9LK0_0;
	wire w_dff_A_dQHTlihh4_0;
	wire w_dff_A_fiWm97NV6_0;
	wire w_dff_A_SAlkhw2R0_0;
	wire w_dff_A_S1wMbJWo4_0;
	wire w_dff_A_HDNNfVWU5_1;
	wire w_dff_A_6sfFDXGC5_0;
	wire w_dff_A_DJP4JRbb1_0;
	wire w_dff_A_LzIu2Qtx1_0;
	wire w_dff_A_nFTDqOIK6_0;
	wire w_dff_A_B4I7hajb7_0;
	wire w_dff_A_byCKrMao9_0;
	wire w_dff_A_vlrU0L6F8_0;
	wire w_dff_A_JaNHCmAC6_0;
	wire w_dff_A_qAoeGtu41_0;
	wire w_dff_A_KEXImDku0_0;
	wire w_dff_A_lYSxZKYt3_0;
	wire w_dff_A_xa7DKjyO9_0;
	wire w_dff_A_SJKwhtJY1_0;
	wire w_dff_A_rK2EIooO4_0;
	wire w_dff_A_zOOgChGn2_0;
	wire w_dff_A_XMT8fIlf2_0;
	wire w_dff_A_MiGnPugq5_0;
	wire w_dff_A_ih7JIhlA5_0;
	wire w_dff_A_aTYq7vq69_0;
	wire w_dff_A_mrxKdql00_0;
	wire w_dff_A_JbZu5Vcb3_0;
	wire w_dff_A_etlZr0Fc4_0;
	wire w_dff_A_y9Fhn2iO1_0;
	wire w_dff_A_aV9d9Ahv4_0;
	wire w_dff_A_HYY14ous9_0;
	wire w_dff_A_EtG2oFGJ4_0;
	wire w_dff_A_y1pevXfH0_0;
	wire w_dff_A_GoPIL2KR7_1;
	wire w_dff_A_DWu12fX50_0;
	wire w_dff_A_7LjJ3fMc4_0;
	wire w_dff_A_1tTXvfZ42_0;
	wire w_dff_A_fBX5UKo41_0;
	wire w_dff_A_pdI9saIx5_0;
	wire w_dff_A_ESBb8mrc3_0;
	wire w_dff_A_m7rtBfeA4_0;
	wire w_dff_A_xwILDn1Y5_0;
	wire w_dff_A_PSfK27IH3_0;
	wire w_dff_A_G2Uyhqqk9_0;
	wire w_dff_A_M75uakEJ4_0;
	wire w_dff_A_6ZQRETnL8_0;
	wire w_dff_A_un8jIdgZ8_0;
	wire w_dff_A_hd0DKlqA9_0;
	wire w_dff_A_auLaSAjA0_0;
	wire w_dff_A_1HORKG3D9_0;
	wire w_dff_A_KSJrzDiw1_0;
	wire w_dff_A_n25SCTnO0_0;
	wire w_dff_A_xX4znLr91_0;
	wire w_dff_A_H1vV2Uvp7_0;
	wire w_dff_A_mgzkWDKP1_0;
	wire w_dff_A_IdCbp0QU7_0;
	wire w_dff_A_NpQUEavQ7_0;
	wire w_dff_A_YT50ht6T6_0;
	wire w_dff_A_0bNf2yhJ3_0;
	wire w_dff_A_aMpuROvk1_0;
	wire w_dff_A_mn5ywUFE7_0;
	wire w_dff_A_ww1qOiDN8_1;
	wire w_dff_A_oZDkyHW71_0;
	wire w_dff_A_4TUklTGv5_0;
	wire w_dff_A_IPfPMvhA0_0;
	wire w_dff_A_CFG0Bizp2_0;
	wire w_dff_A_kQTupb4f6_0;
	wire w_dff_A_lKHZIYm71_0;
	wire w_dff_A_JSKTxqCl3_0;
	wire w_dff_A_sX3p9kSR5_0;
	wire w_dff_A_EJSc661k5_0;
	wire w_dff_A_5GxWJpKR5_0;
	wire w_dff_A_CFECPB2j4_0;
	wire w_dff_A_TI8ynnxC9_0;
	wire w_dff_A_2OFm0dyj1_0;
	wire w_dff_A_Ux3NbOna3_0;
	wire w_dff_A_xJiXxdQC3_0;
	wire w_dff_A_9pqRgPhB8_0;
	wire w_dff_A_8aRsQHeo5_0;
	wire w_dff_A_ZD7TQ8mt0_0;
	wire w_dff_A_zUb32NUd2_0;
	wire w_dff_A_wQqfaZfJ7_0;
	wire w_dff_A_o8ZTUgPI6_0;
	wire w_dff_A_pqDMTDRy9_0;
	wire w_dff_A_URQMZIQf7_0;
	wire w_dff_A_vxa3wBMC8_0;
	wire w_dff_A_0EEZoBeP8_0;
	wire w_dff_A_uNuYueNQ2_0;
	wire w_dff_A_W2A4HmRM0_2;
	wire w_dff_A_QaVnro5g8_0;
	wire w_dff_A_KxJUxQ7X3_0;
	wire w_dff_A_j47V9ViA0_0;
	wire w_dff_A_BQ7zS59F3_0;
	wire w_dff_A_CQFxXwSC1_0;
	wire w_dff_A_NcKCm2RQ7_0;
	wire w_dff_A_RXIdbIa09_0;
	wire w_dff_A_EHAXu3fA2_0;
	wire w_dff_A_yrCYcxV38_0;
	wire w_dff_A_cFaUsFTi2_0;
	wire w_dff_A_ejI6Ifvq5_0;
	wire w_dff_A_yZs6tPzz9_0;
	wire w_dff_A_gmhwfYOt8_0;
	wire w_dff_A_4QCUsUyT2_0;
	wire w_dff_A_JUk62hAx7_0;
	wire w_dff_A_s3nCDSrv4_0;
	wire w_dff_A_dJo9N0FU0_0;
	wire w_dff_A_u0ZNj4eS4_0;
	wire w_dff_A_Q69Txdew0_0;
	wire w_dff_A_hbpHU5w69_0;
	wire w_dff_A_7JiNTrmT1_0;
	wire w_dff_A_Tg0cR9NZ0_0;
	wire w_dff_A_7DowLR0a1_0;
	wire w_dff_A_pG90Hqzz7_2;
	wire w_dff_A_gGbUSuHi7_0;
	wire w_dff_A_387eAaDq7_0;
	wire w_dff_A_KfemJT5K1_0;
	wire w_dff_A_z0fXgH0Q6_0;
	wire w_dff_A_GlzAHUXK5_0;
	wire w_dff_A_EMUK8KtP2_0;
	wire w_dff_A_PQ5XnzNv5_0;
	wire w_dff_A_UELVUXQ85_0;
	wire w_dff_A_HOTDzVDX0_0;
	wire w_dff_A_C7LMqfjb6_0;
	wire w_dff_A_CppgYJzX3_0;
	wire w_dff_A_Au4xGyMt6_0;
	wire w_dff_A_vctVRZiB7_0;
	wire w_dff_A_eqlW5oT55_0;
	wire w_dff_A_uOzBKZdl6_0;
	wire w_dff_A_N2nUkNAX1_0;
	wire w_dff_A_l1Kldsk78_0;
	wire w_dff_A_cG5agdGi3_0;
	wire w_dff_A_lU5vq53o9_0;
	wire w_dff_A_s6joX8Qw8_0;
	wire w_dff_A_kxQeVdnn7_0;
	wire w_dff_A_A3I2hk9F6_0;
	wire w_dff_A_Zh1ey7W62_0;
	wire w_dff_A_m2Bez7pJ5_2;
	wire w_dff_A_IEGiFROW0_0;
	wire w_dff_A_xsR1Qmcl2_0;
	wire w_dff_A_yr3sTo9v8_0;
	wire w_dff_A_qCBLn4np1_0;
	wire w_dff_A_o7HPenKF7_0;
	wire w_dff_A_Mzx3jACP9_0;
	wire w_dff_A_w0Fn9rIC1_0;
	wire w_dff_A_PauUkWI95_0;
	wire w_dff_A_zI7cGY9U8_0;
	wire w_dff_A_HzI259gW3_0;
	wire w_dff_A_vX8f9ZFb7_0;
	wire w_dff_A_tvdyMFT33_0;
	wire w_dff_A_TbiC2r9n2_0;
	wire w_dff_A_tl90zuMQ3_0;
	wire w_dff_A_6ylJ5u3G3_0;
	wire w_dff_A_SuUos7Yg1_0;
	wire w_dff_A_xir742Vt1_0;
	wire w_dff_A_khCv8FGo2_0;
	wire w_dff_A_Xxsm5BjO1_0;
	wire w_dff_A_DBxV72Lx2_0;
	wire w_dff_A_cLLWsM2b5_0;
	wire w_dff_A_h8tZxkCY8_0;
	wire w_dff_A_0nS9Lz9c0_0;
	wire w_dff_A_nCW2wrlb6_2;
	wire w_dff_A_rm3mQbX44_0;
	wire w_dff_A_F0Di5moN0_0;
	wire w_dff_A_JQSx4VDl1_0;
	wire w_dff_A_abWIZwPH1_0;
	wire w_dff_A_NvYfZVb51_0;
	wire w_dff_A_589BAh5Y4_0;
	wire w_dff_A_lwOFuML74_0;
	wire w_dff_A_9948HUf75_0;
	wire w_dff_A_E8gbo8A65_0;
	wire w_dff_A_PB0uCKQX2_0;
	wire w_dff_A_E4NRKFz30_0;
	wire w_dff_A_rMFaMdjO9_0;
	wire w_dff_A_X69S294N0_0;
	wire w_dff_A_rVok3RTO5_0;
	wire w_dff_A_LS5SYU4S1_0;
	wire w_dff_A_z4NDDdqS8_0;
	wire w_dff_A_XKY1MtsD2_0;
	wire w_dff_A_z0QBkL9o7_0;
	wire w_dff_A_ZMnXw3W15_0;
	wire w_dff_A_mZT2myF72_0;
	wire w_dff_A_EB3YUvbq3_0;
	wire w_dff_A_FSklPrXv3_0;
	wire w_dff_A_ODiWA8Hz1_0;
	wire w_dff_A_E2aTN8uK4_0;
	wire w_dff_A_K0bgM94k1_2;
	wire w_dff_A_5rCS99ky1_0;
	wire w_dff_A_BSH08UoT0_0;
	wire w_dff_A_QrvB2chA9_0;
	wire w_dff_A_p5b4U0yj4_0;
	wire w_dff_A_mMmAh9ny7_0;
	wire w_dff_A_27XZIQsn8_0;
	wire w_dff_A_iZztC4bV1_0;
	wire w_dff_A_JFmtOsFX6_0;
	wire w_dff_A_UhOa6Xta4_0;
	wire w_dff_A_p6WqhNZ20_0;
	wire w_dff_A_3T0JLAE56_0;
	wire w_dff_A_fBcBcyuV8_0;
	wire w_dff_A_lzgitMHS2_0;
	wire w_dff_A_Dgr0O5x92_0;
	wire w_dff_A_BjZtKUNQ8_0;
	wire w_dff_A_gD4uF0fg7_0;
	wire w_dff_A_xngBk8al9_0;
	wire w_dff_A_k5uMO6GB6_0;
	wire w_dff_A_Ww1C57Rf7_0;
	wire w_dff_A_RtWKg3an9_0;
	wire w_dff_A_eDcIUdbT6_0;
	wire w_dff_A_LXKUm15T4_0;
	wire w_dff_A_ns2r2A0V2_2;
	wire w_dff_A_VtBd6G8p1_0;
	wire w_dff_A_73VoxK7z4_0;
	wire w_dff_A_idnZIVib4_0;
	wire w_dff_A_V1URt6g21_0;
	wire w_dff_A_ah69EgPr3_0;
	wire w_dff_A_Zr4hPuVN7_0;
	wire w_dff_A_DT8vc6qh1_0;
	wire w_dff_A_lgeWYzjY9_0;
	wire w_dff_A_tX91kvAs7_0;
	wire w_dff_A_AHmpaAUK4_0;
	wire w_dff_A_i54UaYFx6_0;
	wire w_dff_A_kRQ57SEZ2_0;
	wire w_dff_A_cMSEExtz6_0;
	wire w_dff_A_CjLEOFgY2_0;
	wire w_dff_A_Bzqt97gV6_0;
	wire w_dff_A_xJnbnE3e0_0;
	wire w_dff_A_trAH1DME2_0;
	wire w_dff_A_RWTfoV1Q4_0;
	wire w_dff_A_RPFYHpfd9_0;
	wire w_dff_A_99AewqOf5_0;
	wire w_dff_A_PREqOKbW0_0;
	wire w_dff_A_Yiu8GeYD4_0;
	wire w_dff_A_EboTNr2L1_2;
	wire w_dff_A_agnvmFPa9_0;
	wire w_dff_A_oLUkG5Md2_0;
	wire w_dff_A_XurTHM0r8_0;
	wire w_dff_A_5iFLZdds0_0;
	wire w_dff_A_zCqjhmeL4_0;
	wire w_dff_A_7cbJ3MdY6_0;
	wire w_dff_A_aHCI1Iem1_0;
	wire w_dff_A_Y3CTJq573_0;
	wire w_dff_A_LDLh5m0v8_0;
	wire w_dff_A_QFaYvZKE0_0;
	wire w_dff_A_JQOqABNp9_0;
	wire w_dff_A_ztmzWzrH5_0;
	wire w_dff_A_u1ToTu1r3_0;
	wire w_dff_A_93jyY1ri6_0;
	wire w_dff_A_R56LuyJI4_0;
	wire w_dff_A_FmbYh5YL4_0;
	wire w_dff_A_Y62OhfTG7_0;
	wire w_dff_A_xekOnK9u1_0;
	wire w_dff_A_CUwA76FH3_0;
	wire w_dff_A_5t41Rj8X3_0;
	wire w_dff_A_iImP5izh9_0;
	wire w_dff_A_vurdxdhW5_0;
	wire w_dff_A_irTx5kiE2_2;
	wire w_dff_A_qxO0PH441_0;
	wire w_dff_A_6Af8R8TV2_0;
	wire w_dff_A_PDemwxST6_0;
	wire w_dff_A_2tZQv2C57_0;
	wire w_dff_A_DgNsWwQf2_0;
	wire w_dff_A_YxBL8Wh46_0;
	wire w_dff_A_vKrnwEKv9_0;
	wire w_dff_A_U6qTqqy10_0;
	wire w_dff_A_2eqGKT7x7_0;
	wire w_dff_A_RsUMXBdf1_0;
	wire w_dff_A_I0NM0qeH8_0;
	wire w_dff_A_faklq2lQ6_0;
	wire w_dff_A_rJkfP4yh6_0;
	wire w_dff_A_Lp1MU6EB5_0;
	wire w_dff_A_3OkrusRu1_0;
	wire w_dff_A_zUACS2GE0_0;
	wire w_dff_A_JDIWKMuP2_0;
	wire w_dff_A_SJRFcrx57_0;
	wire w_dff_A_KrNVv2cv0_0;
	wire w_dff_A_knLz9pCg4_0;
	wire w_dff_A_YXskZwlQ4_0;
	wire w_dff_A_7sbpixWh0_0;
	wire w_dff_A_n5rTAWwz1_2;
	wire w_dff_A_OitPnp5b6_0;
	wire w_dff_A_Ulv1AIIe5_0;
	wire w_dff_A_cSCjgSiO6_0;
	wire w_dff_A_Rg3GDdbw3_0;
	wire w_dff_A_TFxvzmYG6_0;
	wire w_dff_A_6TOXXDxv9_0;
	wire w_dff_A_TYKCbDKs9_0;
	wire w_dff_A_WQlnJwOw5_0;
	wire w_dff_A_DktPXKxr7_0;
	wire w_dff_A_oCnjY3oC6_0;
	wire w_dff_A_krxf78v44_0;
	wire w_dff_A_QpOltkc82_0;
	wire w_dff_A_9XmaKbEu5_0;
	wire w_dff_A_Bg0I2PMk3_0;
	wire w_dff_A_DOtYBabN3_0;
	wire w_dff_A_S0xPbrrl1_0;
	wire w_dff_A_gr5JutjT0_0;
	wire w_dff_A_FXVMSB5l1_0;
	wire w_dff_A_WWiGWFJq0_0;
	wire w_dff_A_nrahmVjl6_2;
	wire w_dff_A_gJNmfqdw2_0;
	wire w_dff_A_r4LJK7Qq3_0;
	wire w_dff_A_xBT7N27k6_0;
	wire w_dff_A_77Cebwvq4_0;
	wire w_dff_A_DUBoqliQ4_0;
	wire w_dff_A_QpCZgQQK4_0;
	wire w_dff_A_kexmRSBR3_0;
	wire w_dff_A_FnWcXVaO8_0;
	wire w_dff_A_lTAyseaB6_0;
	wire w_dff_A_nTHi0pZl9_0;
	wire w_dff_A_i0wTYvHg5_0;
	wire w_dff_A_1MU40sgG8_0;
	wire w_dff_A_RLp9M79N2_0;
	wire w_dff_A_i7Iqz03p8_0;
	wire w_dff_A_HJXsng5R6_0;
	wire w_dff_A_nfrFDF2U4_0;
	wire w_dff_A_9oS0Va600_0;
	wire w_dff_A_RxNMsRf29_0;
	wire w_dff_A_RHR5feu64_2;
	wire w_dff_A_fF6Xt8aN2_0;
	wire w_dff_A_JqVYQZuN9_0;
	wire w_dff_A_H420Pagp6_0;
	wire w_dff_A_aXamRz1Q6_0;
	wire w_dff_A_lIoPnAyI0_0;
	wire w_dff_A_kvSIjSbT2_0;
	wire w_dff_A_up1A3Lm06_0;
	wire w_dff_A_DZlFkdvP0_0;
	wire w_dff_A_C85mTphH5_0;
	wire w_dff_A_6ePqGiPn9_0;
	wire w_dff_A_4aMRgxII0_0;
	wire w_dff_A_jPfzc2ib4_0;
	wire w_dff_A_ST4ndAa71_0;
	wire w_dff_A_cE1E5OSF7_0;
	wire w_dff_A_E2xsAdWp7_0;
	wire w_dff_A_zJENpbXn5_0;
	wire w_dff_A_QCJjv6qE4_2;
	wire w_dff_A_0noHcg101_0;
	wire w_dff_A_6wgbPrYP3_0;
	wire w_dff_A_2Ghlu4Eg8_0;
	wire w_dff_A_cKMaclMw9_0;
	wire w_dff_A_7gzxcZtL7_0;
	wire w_dff_A_05TkpdN03_0;
	wire w_dff_A_vBGTO0xF7_0;
	wire w_dff_A_gFNU69yT3_0;
	wire w_dff_A_lmAvD1OV4_0;
	wire w_dff_A_mDzFsg8Z9_0;
	wire w_dff_A_hF25cm8s4_0;
	wire w_dff_A_uC5iMHRi3_0;
	wire w_dff_A_GI4CL9851_0;
	wire w_dff_A_xZFobIqm7_0;
	wire w_dff_A_09bONyQn2_0;
	wire w_dff_A_vZUqpITH7_0;
	wire w_dff_A_Khh3TTeo2_0;
	wire w_dff_A_Dg5KC4an0_2;
	wire w_dff_A_eHVHO0sT1_0;
	wire w_dff_A_UCT4t5Rf2_0;
	wire w_dff_A_jZTUOCdY8_0;
	wire w_dff_A_66NDokpo9_0;
	wire w_dff_A_u2qcZ0eh1_0;
	wire w_dff_A_miumCsT48_0;
	wire w_dff_A_z3shtDXP9_0;
	wire w_dff_A_GgbdXAIj5_0;
	wire w_dff_A_2cWTen6x2_0;
	wire w_dff_A_S48hZHOi3_0;
	wire w_dff_A_uIOD6Wp56_0;
	wire w_dff_A_5S5U2Q2c1_0;
	wire w_dff_A_A0V4sbjp7_0;
	wire w_dff_A_Gb4QojF33_0;
	wire w_dff_A_OOOwFFxb5_0;
	wire w_dff_A_1qyQ6q1M1_0;
	wire w_dff_A_e0MEue5I5_0;
	wire w_dff_A_zX1uAcE31_2;
	wire w_dff_A_fw9UzGh89_0;
	wire w_dff_A_ZGTPVf9W2_0;
	wire w_dff_A_DGHH1tyM2_0;
	wire w_dff_A_pxCO5q8I4_0;
	wire w_dff_A_d4sdXjMy7_0;
	wire w_dff_A_tq84brqH5_0;
	wire w_dff_A_QzRkFl9R9_0;
	wire w_dff_A_qTlI0DBE0_0;
	wire w_dff_A_MhIHG7kR8_0;
	wire w_dff_A_SKHzLK3b9_0;
	wire w_dff_A_68nPV9O08_0;
	wire w_dff_A_c7OrDsHw1_0;
	wire w_dff_A_CL1eNI2R0_0;
	wire w_dff_A_2IPaDmAB2_0;
	wire w_dff_A_ZPU5Q32r8_0;
	wire w_dff_A_J06MSiW32_0;
	wire w_dff_A_hM9YJ7h17_1;
	wire w_dff_A_1zHWn9Mh3_0;
	wire w_dff_A_bncCssNd8_0;
	wire w_dff_A_HJk9iyZJ4_0;
	wire w_dff_A_nBradd275_0;
	wire w_dff_A_v4H21F0A9_0;
	wire w_dff_A_RAFoCmNz3_0;
	wire w_dff_A_ObdjxysS5_0;
	wire w_dff_A_mtTWLdfV8_0;
	wire w_dff_A_PFS7FIlM2_0;
	wire w_dff_A_iFjQS5Dp9_0;
	wire w_dff_A_KoroU8UW1_0;
	wire w_dff_A_X4pDVrFQ6_0;
	wire w_dff_A_cgDj8fhF2_0;
	wire w_dff_A_FVSw9pZ65_0;
	wire w_dff_A_covnFvY72_0;
	wire w_dff_A_LNodNHtu9_0;
	wire w_dff_A_wIdL56Et2_0;
	wire w_dff_A_qJbiZyYs6_0;
	wire w_dff_A_vp4rglR89_0;
	wire w_dff_A_v8mPjnKV5_0;
	wire w_dff_A_sBTcLB2d4_0;
	wire w_dff_A_E28C4AF21_0;
	wire w_dff_A_2qWiafb32_1;
	wire w_dff_A_SEkelveQ6_0;
	wire w_dff_A_syackUCF5_0;
	wire w_dff_A_mZEO4lcH5_0;
	wire w_dff_A_Qed4fNtD6_0;
	wire w_dff_A_dnkFVgsd9_0;
	wire w_dff_A_GzdROERb7_0;
	wire w_dff_A_H6pVIzM71_0;
	wire w_dff_A_fWCT3Tbj0_0;
	wire w_dff_A_LJittrPQ2_0;
	wire w_dff_A_O1Ysbbvb8_0;
	wire w_dff_A_wIAaI4lj1_0;
	wire w_dff_A_3AA3RUl77_0;
	wire w_dff_A_epUiVVul2_0;
	wire w_dff_A_SgiBcpn85_0;
	wire w_dff_A_lFX3JfSB8_0;
	wire w_dff_A_jsyb64pj3_0;
	wire w_dff_A_jstxn0x46_0;
	wire w_dff_A_g63k50sU5_0;
	wire w_dff_A_ugv7Mo1N1_0;
	wire w_dff_A_1rfbSUbt9_0;
	wire w_dff_A_Kyr4O1qO0_0;
	wire w_dff_A_yUdAOVuT6_0;
	wire w_dff_A_wVLt2fwl5_2;
	wire w_dff_A_PZCHGf947_0;
	wire w_dff_A_NJ11g6qr5_0;
	wire w_dff_A_mWohJyYd5_0;
	wire w_dff_A_EEbexcJG9_0;
	wire w_dff_A_7Wvr3adD9_0;
	wire w_dff_A_AnjeX9W55_0;
	wire w_dff_A_JeVX2hpH3_0;
	wire w_dff_A_mQ3pGYN86_0;
	wire w_dff_A_XYf36Z6f4_0;
	wire w_dff_A_DzdQewHO0_0;
	wire w_dff_A_RujkW4kl1_0;
	wire w_dff_A_6PA3kwT35_0;
	wire w_dff_A_zdVWXy3r7_0;
	wire w_dff_A_MzAOxEXW9_2;
	wire w_dff_A_9X3Pn8eE2_0;
	wire w_dff_A_qawLeH7P7_0;
	wire w_dff_A_9Rfmas5U0_0;
	wire w_dff_A_jEfDCNv94_0;
	wire w_dff_A_zk8pjiVS4_0;
	wire w_dff_A_OXsUkfJn6_0;
	wire w_dff_A_k4j8aSAO1_0;
	wire w_dff_A_ALiYrbV64_0;
	wire w_dff_A_hAvwYYuR6_0;
	wire w_dff_A_Ma8vgY6H1_0;
	wire w_dff_A_hY6M1ezZ6_0;
	wire w_dff_A_B1Joi4kL7_0;
	wire w_dff_A_tN8T7bLt9_0;
	wire w_dff_A_N8vkVn4P5_0;
	wire w_dff_A_J8PJIiZa7_2;
	wire w_dff_A_UMXLmLoQ3_0;
	wire w_dff_A_IwFPbbez8_0;
	wire w_dff_A_1NNzDRzd3_0;
	wire w_dff_A_LeKReWjO6_0;
	wire w_dff_A_l9rsI4ey3_0;
	wire w_dff_A_cndWKWAL7_0;
	wire w_dff_A_Vmg6RrNA6_0;
	wire w_dff_A_eLXdqB9e3_0;
	wire w_dff_A_3mfnXiYl9_0;
	wire w_dff_A_LGKsPkIc3_0;
	wire w_dff_A_DdYiOf791_0;
	wire w_dff_A_ZRvPIl9d4_0;
	wire w_dff_A_ApMhF7as7_0;
	wire w_dff_A_hRVgxDpe1_2;
	wire w_dff_A_3BKxgBZc2_0;
	wire w_dff_A_W9FL22ak9_0;
	wire w_dff_A_5VJjdRjV6_0;
	wire w_dff_A_UwkYKMji2_0;
	wire w_dff_A_ovQ3zXr26_0;
	wire w_dff_A_1T0kapjh0_0;
	wire w_dff_A_ajMJw7G86_0;
	wire w_dff_A_NGFkhBio2_0;
	wire w_dff_A_ONl7d8SL5_0;
	wire w_dff_A_11F9Sisx4_0;
	wire w_dff_A_dTEu4vA70_0;
	wire w_dff_A_54hU4fjU8_0;
	wire w_dff_A_1kwP5e1J8_0;
	wire w_dff_A_CGf1GCyk1_0;
	wire w_dff_A_SdU8Ychv1_1;
	wire w_dff_A_b59BOzON2_0;
	wire w_dff_A_5evS7cM61_0;
	wire w_dff_A_VQsZAgLQ5_0;
	wire w_dff_A_fvgTNHTg3_0;
	wire w_dff_A_LmxUshWR6_0;
	wire w_dff_A_YLOO6T3Q7_0;
	wire w_dff_A_FiQgZcED1_0;
	wire w_dff_A_TPFL85ES4_0;
	wire w_dff_A_VOrjK6ku2_0;
	wire w_dff_A_8MPjGdTR8_0;
	wire w_dff_A_sit0Az727_0;
	wire w_dff_A_adQgxcG27_0;
	wire w_dff_A_LCRA9Brj1_0;
	wire w_dff_A_T8BgQUx47_0;
	wire w_dff_A_UBPzdATJ5_0;
	wire w_dff_A_Z0mK3ixY2_0;
	wire w_dff_A_5IVW2f2u0_0;
	wire w_dff_A_j99qilMN7_0;
	wire w_dff_A_DUizNmRJ3_0;
	wire w_dff_A_a58wHPnb2_1;
	wire w_dff_A_wYn9j1Et6_0;
	wire w_dff_A_yI9ZSApH4_0;
	wire w_dff_A_lPSCcV8t7_0;
	wire w_dff_A_hDKu8tTO6_0;
	wire w_dff_A_TbUr0Iry2_0;
	wire w_dff_A_HCRNcGUn5_0;
	wire w_dff_A_S4LhQc787_0;
	wire w_dff_A_NTat5lOP9_0;
	wire w_dff_A_EaIYQwfe6_0;
	wire w_dff_A_tYebnlEB2_0;
	wire w_dff_A_WGg9h5RS3_0;
	wire w_dff_A_3wl6G3dr5_0;
	wire w_dff_A_EckDMSF67_0;
	wire w_dff_A_MQf5LBrF0_0;
	wire w_dff_A_32PGN2ft4_1;
	wire w_dff_A_0NT0t0jJ8_0;
	wire w_dff_A_WlYMB3uz7_0;
	wire w_dff_A_lAlYggaD6_0;
	wire w_dff_A_WclX20pc4_0;
	wire w_dff_A_6AHVoOgq9_0;
	wire w_dff_A_gD65qEXj8_0;
	wire w_dff_A_Te0haAZQ7_0;
	wire w_dff_A_x76ZPAeB7_0;
	wire w_dff_A_gLnDJxeA3_0;
	wire w_dff_A_469XsOUb1_0;
	wire w_dff_A_XgfTY49g7_0;
	wire w_dff_A_BWypaNZQ2_0;
	wire w_dff_A_pSruikRH1_0;
	wire w_dff_A_nYalfgC52_0;
	wire w_dff_A_hVbPYwVF4_0;
	wire w_dff_A_ePx9x8A67_0;
	wire w_dff_A_kyW7fDwR3_0;
	wire w_dff_A_3zZlppPo2_1;
	wire w_dff_A_8weYVMmf7_0;
	wire w_dff_A_46xYHbYS7_0;
	wire w_dff_A_O8QUlp923_0;
	wire w_dff_A_qHVTEQ9X1_0;
	wire w_dff_A_LIMCHDzK6_0;
	wire w_dff_A_5Tc8NSCd0_0;
	wire w_dff_A_fZyzX2971_0;
	wire w_dff_A_BjgDiEph7_0;
	wire w_dff_A_8ZxZ9coM0_0;
	wire w_dff_A_GoqX3tdp4_2;
	wire w_dff_A_I9xItxkS9_0;
	wire w_dff_A_uq9sOmXv4_0;
	wire w_dff_A_tNUsV5H25_0;
	wire w_dff_A_Z3uo7zSo0_0;
	wire w_dff_A_nrJ2TCgw8_0;
	wire w_dff_A_ct8DkuX10_0;
	wire w_dff_A_uiLP1dwA9_0;
	wire w_dff_A_ntBSl8Xl6_0;
	wire w_dff_A_HabsYJWC9_0;
	wire w_dff_A_4kUgOLuD8_0;
	wire w_dff_A_QtoxRyzn3_0;
	wire w_dff_A_2RuDNGB85_0;
	wire w_dff_A_cSpm6UOC1_0;
	wire w_dff_A_J4Jmmsg98_1;
	wire w_dff_A_fu8N7Iyj5_0;
	wire w_dff_A_q07gtgke8_0;
	wire w_dff_A_VMTIhTb74_0;
	wire w_dff_A_yxirF8vl7_0;
	wire w_dff_A_7IkhlJY36_0;
	wire w_dff_A_i5pzBwBT1_0;
	wire w_dff_A_K4J5kSOj3_0;
	wire w_dff_A_MEOPsBff9_0;
	wire w_dff_A_eYIqAtBs3_0;
	wire w_dff_A_SpvSlMBR6_0;
	wire w_dff_A_YM9XQKYJ3_0;
	wire w_dff_A_85IV5hjF4_0;
	wire w_dff_A_BZPX3kBd6_1;
	wire w_dff_A_MItrpGh65_0;
	wire w_dff_A_IUypSK960_0;
	wire w_dff_A_XzVI3ZSR3_0;
	wire w_dff_A_f9L7DiAN9_0;
	wire w_dff_A_a2K44Dff4_0;
	wire w_dff_A_Y41Fkdox8_0;
	wire w_dff_A_SPgIzt2E7_0;
	wire w_dff_A_9ssSqLAV8_0;
	wire w_dff_A_CXWCqIcV7_0;
	wire w_dff_A_srJsI7k85_0;
	wire w_dff_A_ADpst9c51_0;
	wire w_dff_A_rrDLn1se8_0;
	wire w_dff_A_hLae4ReT4_0;
	wire w_dff_A_YrJpRzMx9_1;
	wire w_dff_A_vPTUWUZ44_0;
	wire w_dff_A_4mbCgx3w6_0;
	wire w_dff_A_k7kLNezn5_0;
	wire w_dff_A_sSAHpwEj7_0;
	wire w_dff_A_JQ7IdnRW4_0;
	wire w_dff_A_k9QeNSBi3_0;
	wire w_dff_A_V72f7WbK2_0;
	wire w_dff_A_8SZzEg7y1_0;
	wire w_dff_A_ro2KrKeu3_0;
	wire w_dff_A_oIZkV3059_0;
	wire w_dff_A_Rr0bFvnv3_0;
	wire w_dff_A_JwJNc1rY2_0;
	wire w_dff_A_oEGW1y4M4_0;
	wire w_dff_A_jrRy5ZX90_0;
	wire w_dff_A_KAN7zrM39_0;
	wire w_dff_A_P2qeWm9N7_2;
	wire w_dff_A_cqLYJVgY1_0;
	wire w_dff_A_aNPxrL0N8_0;
	wire w_dff_A_JheEaVT01_0;
	wire w_dff_A_zC9WtCeW4_0;
	wire w_dff_A_zr3zYmsV5_0;
	wire w_dff_A_csHtLnaH5_0;
	wire w_dff_A_GLz5aASv1_0;
	wire w_dff_A_wxejWMT14_0;
	wire w_dff_A_lnS1CrEj9_0;
	wire w_dff_A_slRbJA7W9_0;
	wire w_dff_A_71s5LhIN8_0;
	wire w_dff_A_HatCxxBI5_0;
	wire w_dff_A_AKunThgh7_0;
	wire w_dff_A_mblDQHA37_1;
	wire w_dff_A_HJr4ozNT9_0;
	wire w_dff_A_t4aSr7M02_0;
	wire w_dff_A_Lzm1nq0E4_0;
	wire w_dff_A_qo1EGmtQ5_0;
	wire w_dff_A_dBBSXc9N2_0;
	wire w_dff_A_Npxmb5Lo1_0;
	wire w_dff_A_8xbCYDrK9_0;
	wire w_dff_A_V0v7UeVO0_0;
	wire w_dff_A_sl4C8Jhf8_0;
	wire w_dff_A_NMcB3cU60_0;
	wire w_dff_A_BrjD1oyV2_0;
	wire w_dff_A_woudQSwI3_0;
	wire w_dff_A_xLUN1R8u8_1;
	wire w_dff_A_1pgpu9CU4_0;
	wire w_dff_A_pHvWiNJH2_0;
	wire w_dff_A_TxSgeTzU5_0;
	wire w_dff_A_9IYKVSVY5_0;
	wire w_dff_A_2ko0mDBe5_0;
	wire w_dff_A_XQVLFwgm0_0;
	wire w_dff_A_byuaIsk05_0;
	wire w_dff_A_JfdV9wNw2_0;
	wire w_dff_A_UqtS7VJR7_0;
	wire w_dff_A_HLHm30nX3_0;
	wire w_dff_A_VkDpNVKu4_0;
	wire w_dff_A_4qsKLjYg6_0;
	wire w_dff_A_nXrFq2gP6_0;
	wire w_dff_A_GLd1uF4g4_0;
	wire w_dff_A_ze09dhrl2_1;
	wire w_dff_A_GY1YKhKI1_0;
	wire w_dff_A_0bLJJj1N7_0;
	wire w_dff_A_dpm6sj3J4_0;
	wire w_dff_A_q7zv4KAr1_0;
	wire w_dff_A_zNcILBaT1_0;
	wire w_dff_A_um3UCFwv5_0;
	wire w_dff_A_Rn2xYR6i9_0;
	wire w_dff_A_AEgbe3eT1_0;
	wire w_dff_A_uyPdBQa33_0;
	wire w_dff_A_HDBvyhYh9_0;
	wire w_dff_A_KnwHuFUu5_0;
	wire w_dff_A_paBzv8uy5_0;
	wire w_dff_A_NTj0Pi5f6_0;
	wire w_dff_A_WlVZTu3x2_0;
	wire w_dff_A_KkpLYZB45_0;
	wire w_dff_A_5ypKyrfN3_1;
	wire w_dff_A_bY06FGMf2_0;
	wire w_dff_A_58dvA11K9_0;
	wire w_dff_A_gAw9QXNE6_0;
	wire w_dff_A_ZYl6oI143_0;
	wire w_dff_A_wYcYkfCu7_0;
	wire w_dff_A_rhYpeoBP0_0;
	wire w_dff_A_DCkj2Yyc0_0;
	wire w_dff_A_aYqoDzMp9_0;
	wire w_dff_A_nD7vw8y92_0;
	wire w_dff_A_NVLplX6H2_0;
	wire w_dff_A_jwAkuYzq7_0;
	wire w_dff_A_dMmPU1zY1_0;
	wire w_dff_A_8mjvj9zO9_0;
	wire w_dff_A_0TjaEGZH2_0;
	wire w_dff_A_tib2Cl281_0;
	wire w_dff_A_nrb8HoE08_0;
	wire w_dff_A_neliHUfR6_1;
	wire w_dff_A_7ttjikvw7_0;
	wire w_dff_A_0eA05yF12_0;
	wire w_dff_A_f316JV8P5_0;
	wire w_dff_A_llQ1HV8w3_0;
	wire w_dff_A_qzEdIMsg0_0;
	wire w_dff_A_ooEUXoGn2_0;
	wire w_dff_A_x543VmWe4_0;
	wire w_dff_A_lAbSOpQ00_0;
	wire w_dff_A_28wg7lft1_0;
	wire w_dff_A_0Hr276hO9_0;
	wire w_dff_A_mnDWZTTI2_0;
	wire w_dff_A_CeiUXsYt1_0;
	wire w_dff_A_NlECMc2a2_0;
	wire w_dff_A_mLxXGnTj0_0;
	wire w_dff_A_X1wFQt2W8_0;
	wire w_dff_A_usXJEJZa3_0;
	wire w_dff_A_wdxWV2EP4_0;
	wire w_dff_A_WudY5Sp28_0;
	wire w_dff_A_pALQTfio4_0;
	wire w_dff_A_KTZtqfg71_1;
	wire w_dff_A_JQ0oYLoT5_0;
	wire w_dff_A_9Aue2sDH9_0;
	wire w_dff_A_xXSErffV0_0;
	wire w_dff_A_ElVZFpBl4_0;
	wire w_dff_A_efKfqH7a0_0;
	wire w_dff_A_v6ULwx0z3_0;
	wire w_dff_A_ZUq3jIUF3_0;
	wire w_dff_A_1ujXqndR2_0;
	wire w_dff_A_UtlVHKJ78_0;
	wire w_dff_A_fde4e3wZ3_0;
	wire w_dff_A_rt8TLl1A4_0;
	wire w_dff_A_zwAXs2pp4_0;
	wire w_dff_A_JqUsGe384_0;
	wire w_dff_A_PQrMPFrc2_0;
	wire w_dff_A_QsE1JNbt4_0;
	wire w_dff_A_tKPhJvgs8_0;
	wire w_dff_A_rPaLxlP80_0;
	wire w_dff_A_qJgPZP9y1_0;
	wire w_dff_A_oFxVWF266_2;
	wire w_dff_A_9wPjBMDI0_0;
	wire w_dff_A_Mjw2P9eH3_0;
	wire w_dff_A_ahniAdbA5_0;
	wire w_dff_A_cJf3CJ8Y8_0;
	wire w_dff_A_tw4viNqM8_0;
	wire w_dff_A_u2371pY15_0;
	wire w_dff_A_M2Ic8DYe9_0;
	wire w_dff_A_eSkGMLfB8_2;
	wire w_dff_A_Bjhe3bq82_0;
	wire w_dff_A_OMVhnJ9u7_0;
	wire w_dff_A_NftuWoC69_0;
	wire w_dff_A_1GsB7OMm0_0;
	wire w_dff_A_kw1x1V6S9_0;
	wire w_dff_A_9UfzsOYJ1_0;
	wire w_dff_A_IUyZibeU2_2;
	wire w_dff_A_cRRCAO2L6_0;
	wire w_dff_A_svkJMgjO6_0;
	wire w_dff_A_5ugU9kF67_0;
	wire w_dff_A_qqoXLBA01_0;
	wire w_dff_A_jqb47BX42_0;
	wire w_dff_A_lA1THRZE0_0;
	wire w_dff_A_mOyMGvcL5_0;
	wire w_dff_A_51ahXK5G8_0;
	wire w_dff_A_0HRDwkhQ6_0;
	wire w_dff_A_dIWxw3nm3_0;
	wire w_dff_A_PSgSGnz36_0;
	wire w_dff_A_cL0EQVCg1_2;
	wire w_dff_A_Dp0FxNQF2_0;
	wire w_dff_A_w9Ynxlfk2_0;
	wire w_dff_A_i95OBmFU3_0;
	wire w_dff_A_AX8U6Buc9_0;
	wire w_dff_A_2EiIwpA04_0;
	wire w_dff_A_W5mBCs2L4_0;
	wire w_dff_A_bLo8VeWw5_0;
	wire w_dff_A_kS2MxYg51_0;
	wire w_dff_A_6g9mpdPq0_0;
	wire w_dff_A_wlRpliVa4_0;
	wire w_dff_A_k7Y6xbUH1_0;
	wire w_dff_A_IGyoSSEu8_2;
	wire w_dff_A_fnYfrLi49_0;
	wire w_dff_A_07csGbv03_0;
	wire w_dff_A_V8THRWGJ7_0;
	wire w_dff_A_u1LgeGkp8_0;
	wire w_dff_A_O0C8QJB56_0;
	wire w_dff_A_6Seknxoa1_0;
	wire w_dff_A_gXRfmuoD9_0;
	wire w_dff_A_56RrwCqu2_2;
	wire w_dff_A_XSBLuAK12_0;
	wire w_dff_A_TkCiHhqg2_0;
	wire w_dff_A_iBUqbdgB6_0;
	wire w_dff_A_rqyikVq48_0;
	wire w_dff_A_rCYhtEKy0_0;
	wire w_dff_A_LoCEBRb97_0;
	wire w_dff_A_tQ2JJ1wQ9_0;
	wire w_dff_A_3qtcbthX2_0;
	wire w_dff_A_wwQGevd50_2;
	wire w_dff_A_LuCCvnEv7_0;
	wire w_dff_A_iOewLQyw8_0;
	wire w_dff_A_J6hqywOG7_0;
	wire w_dff_A_i38oytxA1_0;
	wire w_dff_A_EiYP8uzZ8_0;
	wire w_dff_A_JMo9xqPC4_0;
	wire w_dff_A_NHRKJE9o0_0;
	wire w_dff_A_vck6t0Ls7_0;
	wire w_dff_A_BCkQIoXj5_0;
	wire w_dff_A_zCFXhFnS0_0;
	wire w_dff_A_keQaPtPi2_2;
	wire w_dff_A_GuMAt2f15_0;
	wire w_dff_A_awe276pv0_0;
	wire w_dff_A_6vyJ4y485_0;
	wire w_dff_A_L2bcmLza9_0;
	wire w_dff_A_fUGivxGM4_0;
	wire w_dff_A_o0JrcGDO4_0;
	wire w_dff_A_cYm2RJ1k5_0;
	wire w_dff_A_uzM1zUeL4_0;
	wire w_dff_A_tIXEG92T5_0;
	wire w_dff_A_7oyN7Kg98_2;
	wire w_dff_A_yrqbt1aF4_0;
	wire w_dff_A_15HlcQp52_0;
	wire w_dff_A_1LRZ8Qgk5_0;
	wire w_dff_A_eh7ZjtDn5_0;
	wire w_dff_A_jjTVRLTX2_0;
	wire w_dff_A_Q9ukMb3J0_0;
	wire w_dff_A_GTOmaDn06_0;
	wire w_dff_A_HwrRny5T3_2;
	wire w_dff_A_IZXO5wd74_0;
	wire w_dff_A_R1pQn5dn0_0;
	wire w_dff_A_kWHmk5Ik3_0;
	wire w_dff_A_E7lF4cOj9_0;
	wire w_dff_A_LaEpSJrB2_0;
	wire w_dff_A_mT5BA4oI3_0;
	wire w_dff_A_erYO3d858_0;
	wire w_dff_A_KWCJk61z9_0;
	wire w_dff_A_hBJRCEio6_2;
	wire w_dff_A_4lWHOGkr7_0;
	wire w_dff_A_R7L5ePMw5_0;
	wire w_dff_A_EonOOZV55_0;
	wire w_dff_A_z2Y2UXP12_0;
	wire w_dff_A_6M29mEZe3_0;
	wire w_dff_A_35N0HQvi8_0;
	wire w_dff_A_nxmcxN7M2_0;
	wire w_dff_A_pkA0WnTx7_0;
	wire w_dff_A_UyNzVoq93_0;
	wire w_dff_A_YPP1kP491_0;
	wire w_dff_A_kRGQhKKq4_2;
	wire w_dff_A_WIc5xmtn9_0;
	wire w_dff_A_BZfoMNOJ8_0;
	wire w_dff_A_OKVU27gA8_0;
	wire w_dff_A_6M90IALQ6_0;
	wire w_dff_A_22v3171a1_0;
	wire w_dff_A_pnzLAGUv5_0;
	wire w_dff_A_MrILsDGm1_0;
	wire w_dff_A_QaFzE0QM7_0;
	wire w_dff_A_OZueif6j5_0;
	wire w_dff_A_wjAAGGZN0_2;
	wire w_dff_A_g6WAay8Z1_0;
	wire w_dff_A_JHpN8vBq4_0;
	wire w_dff_A_kPOWcMVs8_0;
	wire w_dff_A_reObvyOt0_0;
	wire w_dff_A_mX0XWHp30_0;
	wire w_dff_A_kFMhfeua5_0;
	wire w_dff_A_kbovglEb0_2;
	wire w_dff_A_kYSdAvvG4_0;
	wire w_dff_A_aF8eCFso6_0;
	wire w_dff_A_GjRz2egv7_0;
	wire w_dff_A_AwlHth9f5_0;
	wire w_dff_A_LviuiotL2_0;
	wire w_dff_A_AINrNPxn4_0;
	wire w_dff_A_rE8qxiW14_0;
	wire w_dff_A_u3zsD5KS2_0;
	wire w_dff_A_fxDlBdr66_0;
	wire w_dff_A_ss9SJ2Xo4_2;
	wire w_dff_A_P0Dx8lPm9_0;
	wire w_dff_A_0Etvfc4Q2_0;
	wire w_dff_A_qFpBRhTS2_0;
	wire w_dff_A_zdbF1X6j9_0;
	wire w_dff_A_4yIGQfuL3_0;
	wire w_dff_A_pXW0sItH6_0;
	wire w_dff_A_Ox42J1yh8_0;
	wire w_dff_A_pU10xJRe7_0;
	wire w_dff_A_sK2mi3pL2_0;
	wire w_dff_A_tBBw127J7_2;
	wire w_dff_A_oYjsusMY9_0;
	wire w_dff_A_CytBECid0_0;
	wire w_dff_A_IhNYKsG56_0;
	wire w_dff_A_1ual1f6d6_0;
	wire w_dff_A_cdKTJHI05_0;
	wire w_dff_A_FkZIukp17_0;
	wire w_dff_A_qzhJV5k79_0;
	wire w_dff_A_ogcvh6NP5_0;
	wire w_dff_A_FJ4eLE8y0_2;
	wire w_dff_A_PYdsn7pj3_0;
	wire w_dff_A_DHmYaf239_0;
	wire w_dff_A_7mmAos5b6_0;
	wire w_dff_A_9KSwdT595_0;
	wire w_dff_A_FoxYZBO38_0;
	wire w_dff_A_aPMm9gZk7_2;
	wire w_dff_A_3d66GSyw0_0;
	wire w_dff_A_6f2ZC6wu8_0;
	wire w_dff_A_G0NcBXiA6_0;
	wire w_dff_A_ray4PLmV4_0;
	wire w_dff_A_e1CuurEu2_0;
	wire w_dff_A_aZGTDgYD1_0;
	wire w_dff_A_fOOG70532_0;
	wire w_dff_A_HSBN9R1w9_0;
	wire w_dff_A_7QjQD5T44_0;
	wire w_dff_A_E416vl2P8_2;
	wire w_dff_A_P2jh8dN06_0;
	wire w_dff_A_crW3mDMJ7_0;
	wire w_dff_A_D00Sfr7D3_0;
	wire w_dff_A_sVFNQS8M3_0;
	wire w_dff_A_Q4v9FAB68_0;
	wire w_dff_A_ZWBjnRSv6_0;
	wire w_dff_A_Zk63SCOk5_0;
	wire w_dff_A_J6AimyZZ1_0;
	wire w_dff_A_gIpfvbWy7_0;
	wire w_dff_A_88KRnGpV7_2;
	wire w_dff_A_cYNTIumU9_0;
	wire w_dff_A_qeJVB7y90_0;
	wire w_dff_A_iwUG8mUG7_0;
	wire w_dff_A_Jeo8Nlfx1_0;
	wire w_dff_A_LXsOzG986_0;
	wire w_dff_A_UnA1ZE3e4_0;
	wire w_dff_A_Ur1W488X2_0;
	wire w_dff_A_DjupPxtm5_0;
	wire w_dff_A_oxuB7DjA9_2;
	wire w_dff_A_NxfNV3OH9_0;
	wire w_dff_A_OGGUHDmq4_0;
	wire w_dff_A_F598HQwd0_0;
	wire w_dff_A_rsCdqn5b3_0;
	wire w_dff_A_qIdEvIDR4_0;
	wire w_dff_A_RuC4hOr78_0;
	wire w_dff_A_jvwhkrDN8_2;
	wire w_dff_A_Y8d1aVOm5_0;
	wire w_dff_A_WaqFKYA54_0;
	wire w_dff_A_0kpxCFv33_0;
	wire w_dff_A_2ii10nXG5_0;
	wire w_dff_A_vgKVjSJ16_0;
	wire w_dff_A_2g2eiFvr1_0;
	wire w_dff_A_0BRhGLFc0_0;
	wire w_dff_A_j2omylgn7_0;
	wire w_dff_A_NIxKrJk80_0;
	wire w_dff_A_UrnIQvBs9_1;
	wire w_dff_A_z4hFqVTR2_0;
	wire w_dff_A_6GBVhRSQ7_0;
	wire w_dff_A_790Qc8Pg4_0;
	wire w_dff_A_SmfxvG303_0;
	wire w_dff_A_jqG8pdYj3_0;
	wire w_dff_A_piCXS0Pd0_0;
	wire w_dff_A_Fi5KrCYh7_1;
	wire w_dff_A_XU6G4Rnz6_0;
	wire w_dff_A_FOj9cwjG6_0;
	wire w_dff_A_7UcrxjYU9_0;
	wire w_dff_A_W1WjV6JE5_0;
	wire w_dff_A_4GH99eSJ4_0;
	wire w_dff_A_Acvk601o3_0;
	wire w_dff_A_w03832J53_0;
	wire w_dff_A_5bYRvP0i0_1;
	wire w_dff_A_sfPU4EOk3_0;
	wire w_dff_A_BlEsbe956_0;
	wire w_dff_A_h3Ni1l6T0_0;
	wire w_dff_A_EydOHUhY4_0;
	wire w_dff_A_7h98kp6x0_0;
	wire w_dff_A_whgDnFsH7_0;
	wire w_dff_A_RKhsEVmw6_1;
	wire w_dff_A_Ps8KofOz1_0;
	wire w_dff_A_uOYJOAMV8_0;
	wire w_dff_A_KzkGDMLA5_0;
	wire w_dff_A_N3n9LPEy2_0;
	wire w_dff_A_mA14aquq8_0;
	wire w_dff_A_GHyijkEL1_0;
	wire w_dff_A_V6fy43pr2_0;
	wire w_dff_A_R4gtxDkT9_0;
	wire w_dff_A_zcwqaNIL1_0;
	wire w_dff_A_P3klW2aS8_0;
	wire w_dff_A_grsRAp8K6_0;
	wire w_dff_A_vafD6ff48_2;
	wire w_dff_A_NHbc80Du1_0;
	wire w_dff_A_GjT1u7DS1_0;
	wire w_dff_A_egeNTtbU8_0;
	wire w_dff_A_lZi2bb4Y7_0;
	wire w_dff_A_WSu8YH2N6_0;
	wire w_dff_A_YgU5vIS79_0;
	wire w_dff_A_yLvlILzf0_0;
	wire w_dff_A_6H7heQwo1_0;
	wire w_dff_A_WDpuXTtO2_0;
	wire w_dff_A_iYgPbrkt8_0;
	wire w_dff_A_cJaLg3Re5_0;
	wire w_dff_A_wJrX1xWD4_0;
	wire w_dff_A_aeYc1dxD1_0;
	wire w_dff_A_GlxHJIEL1_0;
	wire w_dff_A_d4XYNGRD4_0;
	wire w_dff_A_sEelVtlB0_0;
	wire w_dff_A_MInp1sVP2_1;
	wire w_dff_A_spmEkXTn4_0;
	wire w_dff_A_jWlY2xyu9_0;
	wire w_dff_A_NOkych6E0_0;
	wire w_dff_A_4ojF5srM0_0;
	wire w_dff_A_Zf2BjFUE2_0;
	wire w_dff_A_cJBm3tzC8_1;
	wire w_dff_A_TTTwWwf34_0;
	wire w_dff_A_LhvBKKL64_0;
	wire w_dff_A_28qXxs1M3_0;
	wire w_dff_A_eFsPG5Va8_0;
	wire w_dff_A_Il93Y7Ju3_0;
	wire w_dff_A_so1IeFct6_0;
	wire w_dff_A_JRyMNrnF2_0;
	wire w_dff_A_G5tlOvfn8_0;
	wire w_dff_A_CZVTd2RE5_1;
	wire w_dff_A_wlNhtr8z1_0;
	wire w_dff_A_4ixODqpk9_0;
	wire w_dff_A_j3eFymXy2_0;
	wire w_dff_A_Z2ZM1x5n9_0;
	wire w_dff_A_okzo6YL03_0;
	wire w_dff_A_bM3xybTO2_0;
	wire w_dff_A_j23ZqMUB9_1;
	wire w_dff_A_BripIcQc4_0;
	wire w_dff_A_nkxwIEI26_0;
	wire w_dff_A_7thvBMRw5_0;
	wire w_dff_A_W4DvVmCP1_0;
	wire w_dff_A_Eda2cVrQ1_0;
	wire w_dff_A_raUYjNWG4_0;
	wire w_dff_A_NscxkqwB6_0;
	wire w_dff_A_Qz1Vf87J9_0;
	wire w_dff_A_0lvFX9Rn9_0;
	wire w_dff_A_2XGOUCxJ2_2;
	wire w_dff_A_L4YhNQt45_0;
	wire w_dff_A_LZr3Dsus0_0;
	wire w_dff_A_23BSm3Fp3_0;
	wire w_dff_A_fDdSOlMD0_2;
	wire w_dff_A_SN76x4gC2_0;
	wire w_dff_A_iJYymryz2_0;
	wire w_dff_A_5eIRg5hX3_2;
	wire w_dff_A_aaW5Ixtd9_0;
	wire w_dff_A_jYli0LbD5_0;
	wire w_dff_A_82A8IQ7J9_0;
	wire w_dff_A_sYyisCNw9_2;
	wire w_dff_A_uwf4jsWY1_0;
	wire w_dff_A_fvUwqR9F9_0;
	wire w_dff_A_igVS6zOD9_0;
	wire w_dff_A_jLaVIWAZ5_2;
	wire w_dff_A_zobrglLG5_0;
	wire w_dff_A_8BKcmYGu9_0;
	wire w_dff_A_CRzGPY5k9_0;
	wire w_dff_A_fMd2qyrI0_0;
	wire w_dff_A_jHQxUsEJ2_2;
	wire w_dff_A_VJVUz5976_0;
	wire w_dff_A_QSIPoHGe8_0;
	wire w_dff_A_W8Hw7NkO9_0;
	wire w_dff_A_nrcvRrKO0_2;
	wire w_dff_A_T2CRHUaN5_0;
	wire w_dff_A_CRb5XH6s3_0;
	wire w_dff_A_BeeoD6W52_0;
	wire w_dff_A_7DtcfDVl6_2;
	wire w_dff_A_SpizzXDb1_0;
	wire w_dff_A_9Ei9FrSA4_0;
	wire w_dff_A_uoq4p2iG1_0;
	wire w_dff_A_G8XakyhD1_0;
	wire w_dff_A_P32bXcZR1_2;
	wire w_dff_A_zJ9g5eMu7_0;
	wire w_dff_A_49XX6y1L1_0;
	wire w_dff_A_nB1rVZ1i2_0;
	wire w_dff_A_7lXH9BOj8_2;
	wire w_dff_A_O2WopYZH8_0;
	wire w_dff_A_BTztYjhw3_0;
	wire w_dff_A_6ondWxNN6_2;
	wire w_dff_A_RJ2UJ6Ua3_0;
	wire w_dff_A_SmIMZAQG8_0;
	wire w_dff_A_EW50mF6G8_2;
	wire w_dff_A_ToC18BX84_0;
	wire w_dff_A_qtIVFaz20_2;
	wire w_dff_A_sohk3fe49_0;
	wire w_dff_A_DL8HlS531_0;
	wire w_dff_A_Y83qaQXm3_0;
	wire w_dff_A_SZppPzwU8_2;
	wire w_dff_A_KWQ3KdOQ2_0;
	wire w_dff_A_DduDY9mV2_0;
	wire w_dff_A_EjeCPIAX3_2;
	wire w_dff_A_lSRPRseG4_0;
	wire w_dff_A_wmPkw9R00_0;
	wire w_dff_A_NyJ1LQKr6_2;
	wire w_dff_A_J5tMnEw31_0;
	wire w_dff_A_s8pDORCC1_0;
	wire w_dff_A_VYoWKH9V5_2;
	wire w_dff_A_iQeJaTKS7_0;
	wire w_dff_A_pjJjMj0F8_0;
	wire w_dff_A_Sd2CgZtn5_0;
	wire w_dff_A_PUbC0Vfa6_0;
	wire w_dff_A_uX9slJXe3_0;
	wire w_dff_A_6B9aVpnN0_2;
	wire w_dff_A_ZMGT75uD3_0;
	wire w_dff_A_C32bfpmL1_0;
	wire w_dff_A_jHkqsqtz0_0;
	wire w_dff_A_gPiOw7G95_0;
	wire w_dff_A_cscWtQnO0_0;
	wire w_dff_A_xjst1swX1_2;
	wire w_dff_A_73jqJqeU4_2;
	jnot g0000(.din(w_G545_0[2]),.dout(w_dff_A_ZBrec1Vu5_1),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(w_G366_0[1]),.dout(w_dff_A_9M7VFoQ81_1),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(w_dff_A_KwFthaXT7_1),.clk(gclk));
	jnot g0005(.din(w_G338_0[1]),.dout(w_dff_A_UzBVPGlV5_1),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(w_dff_A_PGzCSuv27_2),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(w_dff_A_hnSczvAh8_1),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(w_dff_A_E78jADKM5_1),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(w_dff_A_AVwe8LZD9_1),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(w_dff_A_8yW8rYSC0_1),.clk(gclk));
	jand g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(w_dff_A_il5gzRQ12_2),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_zheJpM8a6_1),.dout(w_dff_A_5yZAzLY28_2),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jor g0016(.dina(w_dff_B_AHgrt4gg1_0),.dinb(w_n316_0[1]),.dout(w_dff_A_Dfh0sref6_2),.clk(gclk));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(w_dff_A_9IakLXyU2_1),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jor g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_),.clk(gclk));
	jor g0022(.dina(w_G809_3[1]),.dinb(w_dff_B_qYdKW0mJ1_1),.dout(w_dff_A_Cg0ajXrl8_2),.clk(gclk));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jor g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330),.clk(gclk));
	jor g0030(.dina(n330),.dinb(w_dff_B_fb4w6OY08_1),.dout(w_dff_A_W2A4HmRM0_2),.clk(gclk));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jor g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336),.clk(gclk));
	jor g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(w_dff_A_pG90Hqzz7_2),.clk(gclk));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jor g0038(.dina(w_G809_2[1]),.dinb(w_dff_B_bn2KitwD0_1),.dout(w_dff_A_nCW2wrlb6_2),.clk(gclk));
	jand g0039(.dina(w_n326_1[2]),.dinb(w_dff_B_yhLpS0385_1),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jor g0041(.dina(w_dff_B_rt3JmqTJ3_0),.dinb(w_G809_2[0]),.dout(n342),.clk(gclk));
	jor g0042(.dina(n342),.dinb(w_dff_B_y0l8qKDv5_1),.dout(n343),.clk(gclk));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(w_dff_A_K0bgM94k1_2),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(w_dff_B_B3mKvrRi2_1),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jor g0046(.dina(w_dff_B_mF2s9CBA5_0),.dinb(w_G809_1[2]),.dout(n347),.clk(gclk));
	jor g0047(.dina(n347),.dinb(w_dff_B_6QeaS1DH6_1),.dout(n348),.clk(gclk));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(w_dff_A_ns2r2A0V2_2),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(w_dff_B_R8DwcryY0_1),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jor g0051(.dina(w_dff_B_F9C7J14E4_0),.dinb(w_G809_1[1]),.dout(n352),.clk(gclk));
	jor g0052(.dina(n352),.dinb(w_dff_B_p6DqrFtN8_1),.dout(n353),.clk(gclk));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(w_dff_A_EboTNr2L1_2),.clk(gclk));
	jand g0054(.dina(w_G2358_0[2]),.dinb(G80),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_n326_0[2]),.dinb(w_dff_B_ujKs66H17_1),.dout(n356),.clk(gclk));
	jor g0056(.dina(n356),.dinb(w_G809_1[0]),.dout(n357),.clk(gclk));
	jor g0057(.dina(n357),.dinb(w_dff_B_uJshMeGM7_1),.dout(n358),.clk(gclk));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(w_dff_A_irTx5kiE2_2),.clk(gclk));
	jand g0059(.dina(w_G3552_0[1]),.dinb(w_G514_2[1]),.dout(n360),.clk(gclk));
	jnot g0060(.din(w_G514_2[0]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G3546_5[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(n362),.dinb(w_n361_0[1]),.dout(n363),.clk(gclk));
	jor g0063(.dina(n363),.dinb(w_dff_B_ub1rWXPF9_1),.dout(n364),.clk(gclk));
	jnot g0064(.din(n364),.dout(n365),.clk(gclk));
	jnot g0065(.din(w_G251_5[1]),.dout(n366),.clk(gclk));
	jnot g0066(.din(w_G361_1[1]),.dout(n367),.clk(gclk));
	jand g0067(.dina(n367),.dinb(w_n366_1[2]),.dout(n368),.clk(gclk));
	jnot g0068(.din(w_G248_5[2]),.dout(n369),.clk(gclk));
	jand g0069(.dina(w_G361_1[0]),.dinb(w_n369_1[2]),.dout(n370),.clk(gclk));
	jor g0070(.dina(n370),.dinb(n368),.dout(n371),.clk(gclk));
	jnot g0071(.din(w_n371_0[1]),.dout(n372),.clk(gclk));
	jand g0072(.dina(w_n372_0[1]),.dinb(w_n365_0[1]),.dout(n373),.clk(gclk));
	jnot g0073(.din(w_G351_2[2]),.dout(n374),.clk(gclk));
	jnot g0074(.din(G3550),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_n375_4[2]),.dinb(w_n374_1[1]),.dout(n376),.clk(gclk));
	jnot g0076(.din(w_G534_2[1]),.dout(n377),.clk(gclk));
	jnot g0077(.din(w_G3552_0[0]),.dout(n378),.clk(gclk));
	jand g0078(.dina(w_n378_4[2]),.dinb(w_G351_2[1]),.dout(n379),.clk(gclk));
	jor g0079(.dina(n379),.dinb(w_n377_1[1]),.dout(n380),.clk(gclk));
	jor g0080(.dina(n380),.dinb(w_dff_B_SyeDNte46_1),.dout(n381),.clk(gclk));
	jand g0081(.dina(w_G3546_5[0]),.dinb(w_G351_2[0]),.dout(n382),.clk(gclk));
	jand g0082(.dina(w_G3548_4[2]),.dinb(w_n374_1[0]),.dout(n383),.clk(gclk));
	jor g0083(.dina(n383),.dinb(w_dff_B_QIFB1MSw6_1),.dout(n384),.clk(gclk));
	jor g0084(.dina(n384),.dinb(w_G534_2[0]),.dout(n385),.clk(gclk));
	jand g0085(.dina(n385),.dinb(n381),.dout(n386),.clk(gclk));
	jnot g0086(.din(w_G341_2[2]),.dout(n387),.clk(gclk));
	jand g0087(.dina(w_n375_4[1]),.dinb(w_n387_1[1]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G523_1[2]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n378_4[1]),.dinb(w_G341_2[1]),.dout(n390),.clk(gclk));
	jor g0090(.dina(n390),.dinb(w_n389_1[1]),.dout(n391),.clk(gclk));
	jor g0091(.dina(n391),.dinb(w_dff_B_U9XiRrDq4_1),.dout(n392),.clk(gclk));
	jand g0092(.dina(w_G3546_4[2]),.dinb(w_G341_2[0]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3548_4[1]),.dinb(w_n387_1[0]),.dout(n394),.clk(gclk));
	jor g0094(.dina(n394),.dinb(w_dff_B_a2IDp3261_1),.dout(n395),.clk(gclk));
	jor g0095(.dina(n395),.dinb(w_G523_1[1]),.dout(n396),.clk(gclk));
	jand g0096(.dina(n396),.dinb(n392),.dout(n397),.clk(gclk));
	jand g0097(.dina(w_n397_0[1]),.dinb(w_n386_0[1]),.dout(n398),.clk(gclk));
	jand g0098(.dina(n398),.dinb(w_dff_B_oCKraORR2_1),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G316_1[1]),.dinb(w_G248_5[1]),.dout(n400),.clk(gclk));
	jnot g0100(.din(w_G490_1[1]),.dout(n401),.clk(gclk));
	jnot g0101(.din(w_G316_1[0]),.dout(n402),.clk(gclk));
	jand g0102(.dina(w_n402_0[2]),.dinb(w_G251_5[0]),.dout(n403),.clk(gclk));
	jor g0103(.dina(n403),.dinb(w_n401_0[1]),.dout(n404),.clk(gclk));
	jor g0104(.dina(n404),.dinb(w_dff_B_8q75BwXS0_1),.dout(n405),.clk(gclk));
	jnot g0105(.din(w_G254_1[1]),.dout(n406),.clk(gclk));
	jand g0106(.dina(w_n402_0[1]),.dinb(w_n406_5[1]),.dout(n407),.clk(gclk));
	jnot g0107(.din(w_G242_1[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_G316_0[2]),.dinb(w_n408_5[2]),.dout(n409),.clk(gclk));
	jor g0109(.dina(n409),.dinb(n407),.dout(n410),.clk(gclk));
	jor g0110(.dina(n410),.dinb(w_G490_1[0]),.dout(n411),.clk(gclk));
	jand g0111(.dina(n411),.dinb(n405),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G308_1[2]),.dinb(w_G248_5[0]),.dout(n413),.clk(gclk));
	jnot g0113(.din(w_G479_0[2]),.dout(n414),.clk(gclk));
	jnot g0114(.din(w_G308_1[1]),.dout(n415),.clk(gclk));
	jand g0115(.dina(w_n415_0[1]),.dinb(w_G251_4[2]),.dout(n416),.clk(gclk));
	jor g0116(.dina(n416),.dinb(w_n414_0[1]),.dout(n417),.clk(gclk));
	jor g0117(.dina(n417),.dinb(w_dff_B_6UrklJ322_1),.dout(n418),.clk(gclk));
	jand g0118(.dina(w_n415_0[0]),.dinb(w_n406_5[0]),.dout(n419),.clk(gclk));
	jand g0119(.dina(w_G308_1[0]),.dinb(w_n408_5[1]),.dout(n420),.clk(gclk));
	jor g0120(.dina(n420),.dinb(n419),.dout(n421),.clk(gclk));
	jor g0121(.dina(n421),.dinb(w_G479_0[1]),.dout(n422),.clk(gclk));
	jand g0122(.dina(n422),.dinb(n418),.dout(n423),.clk(gclk));
	jand g0123(.dina(w_n423_0[2]),.dinb(w_n412_0[2]),.dout(n424),.clk(gclk));
	jnot g0124(.din(w_G293_0[2]),.dout(n425),.clk(gclk));
	jand g0125(.dina(w_n425_0[2]),.dinb(w_n406_4[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_G293_0[1]),.dinb(w_n408_5[0]),.dout(n427),.clk(gclk));
	jor g0127(.dina(n427),.dinb(n426),.dout(n428),.clk(gclk));
	jnot g0128(.din(w_G302_0[2]),.dout(n429),.clk(gclk));
	jand g0129(.dina(w_n429_0[1]),.dinb(w_n366_1[1]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G302_0[1]),.dinb(w_n369_1[1]),.dout(n431),.clk(gclk));
	jor g0131(.dina(n431),.dinb(n430),.dout(n432),.clk(gclk));
	jnot g0132(.din(n432),.dout(n433),.clk(gclk));
	jand g0133(.dina(w_n433_0[2]),.dinb(w_n428_1[1]),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G324_1[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n375_4[0]),.dinb(w_n435_2[1]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G503_2[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n378_4[0]),.dinb(w_G324_1[1]),.dout(n438),.clk(gclk));
	jor g0138(.dina(n438),.dinb(w_n437_0[1]),.dout(n439),.clk(gclk));
	jor g0139(.dina(n439),.dinb(w_dff_B_f9YYUJeb7_1),.dout(n440),.clk(gclk));
	jand g0140(.dina(w_G3546_4[1]),.dinb(w_G324_1[0]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3548_4[0]),.dinb(w_n435_2[0]),.dout(n442),.clk(gclk));
	jor g0142(.dina(n442),.dinb(w_dff_B_w0Q4eRMQ9_1),.dout(n443),.clk(gclk));
	jor g0143(.dina(n443),.dinb(w_G503_2[0]),.dout(n444),.clk(gclk));
	jand g0144(.dina(n444),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(n434),.dout(n446),.clk(gclk));
	jand g0146(.dina(n446),.dinb(n424),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(n399),.dout(w_dff_A_n5rTAWwz1_2),.clk(gclk));
	jnot g0148(.din(w_G210_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n375_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G457_1[2]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n378_3[2]),.dinb(w_G210_2[0]),.dout(n452),.clk(gclk));
	jor g0152(.dina(n452),.dinb(w_n451_0[2]),.dout(n453),.clk(gclk));
	jor g0153(.dina(n453),.dinb(w_dff_B_35rSU6h96_1),.dout(n454),.clk(gclk));
	jand g0154(.dina(w_G3546_4[0]),.dinb(w_G210_1[2]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n456),.clk(gclk));
	jor g0156(.dina(n456),.dinb(w_dff_B_L640B3lG0_1),.dout(n457),.clk(gclk));
	jor g0157(.dina(n457),.dinb(w_G457_1[1]),.dout(n458),.clk(gclk));
	jand g0158(.dina(n458),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n375_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n378_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jor g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464),.clk(gclk));
	jor g0164(.dina(n464),.dinb(w_dff_B_E4vL1V1K6_1),.dout(n465),.clk(gclk));
	jand g0165(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n467),.clk(gclk));
	jor g0167(.dina(n467),.dinb(w_dff_B_7ogaCzHa8_1),.dout(n468),.clk(gclk));
	jor g0168(.dina(n468),.dinb(w_G435_1[1]),.dout(n469),.clk(gclk));
	jand g0169(.dina(n469),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G273_2[1]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n375_3[0]),.dinb(w_n471_1[2]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G411_2[1]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n378_3[0]),.dinb(w_G273_2[0]),.dout(n474),.clk(gclk));
	jor g0174(.dina(n474),.dinb(w_n473_1[1]),.dout(n475),.clk(gclk));
	jor g0175(.dina(n475),.dinb(w_dff_B_GSMPQl2M4_1),.dout(n476),.clk(gclk));
	jand g0176(.dina(w_G3546_3[1]),.dinb(w_G273_1[2]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3548_3[0]),.dinb(w_n471_1[1]),.dout(n478),.clk(gclk));
	jor g0178(.dina(n478),.dinb(w_dff_B_24dM6nyX0_1),.dout(n479),.clk(gclk));
	jor g0179(.dina(n479),.dinb(w_G411_2[0]),.dout(n480),.clk(gclk));
	jand g0180(.dina(n480),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jnot g0182(.din(w_G265_1[2]),.dout(n483),.clk(gclk));
	jand g0183(.dina(w_n375_2[2]),.dinb(w_n483_2[1]),.dout(n484),.clk(gclk));
	jnot g0184(.din(w_G400_1[2]),.dout(n485),.clk(gclk));
	jand g0185(.dina(w_n378_2[2]),.dinb(w_G265_1[1]),.dout(n486),.clk(gclk));
	jor g0186(.dina(n486),.dinb(w_n485_1[1]),.dout(n487),.clk(gclk));
	jor g0187(.dina(n487),.dinb(w_dff_B_RgaHLtTI8_1),.dout(n488),.clk(gclk));
	jand g0188(.dina(w_G3546_3[0]),.dinb(w_G265_1[0]),.dout(n489),.clk(gclk));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n483_2[0]),.dout(n490),.clk(gclk));
	jor g0190(.dina(n490),.dinb(w_dff_B_WhjvR4bw5_1),.dout(n491),.clk(gclk));
	jor g0191(.dina(n491),.dinb(w_G400_1[1]),.dout(n492),.clk(gclk));
	jand g0192(.dina(n492),.dinb(n488),.dout(n493),.clk(gclk));
	jnot g0193(.din(w_G226_2[1]),.dout(n494),.clk(gclk));
	jand g0194(.dina(w_n375_2[1]),.dinb(w_n494_1[2]),.dout(n495),.clk(gclk));
	jnot g0195(.din(w_G422_1[1]),.dout(n496),.clk(gclk));
	jand g0196(.dina(w_n378_2[1]),.dinb(w_G226_2[0]),.dout(n497),.clk(gclk));
	jor g0197(.dina(n497),.dinb(w_n496_1[1]),.dout(n498),.clk(gclk));
	jor g0198(.dina(n498),.dinb(w_dff_B_5spP29TG4_1),.dout(n499),.clk(gclk));
	jand g0199(.dina(w_G3546_2[2]),.dinb(w_G226_1[2]),.dout(n500),.clk(gclk));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n494_1[1]),.dout(n501),.clk(gclk));
	jor g0201(.dina(n501),.dinb(w_dff_B_UlI2Nhbz5_1),.dout(n502),.clk(gclk));
	jor g0202(.dina(n502),.dinb(w_G422_1[0]),.dout(n503),.clk(gclk));
	jand g0203(.dina(n503),.dinb(n499),.dout(n504),.clk(gclk));
	jand g0204(.dina(w_n504_0[1]),.dinb(w_n493_0[1]),.dout(n505),.clk(gclk));
	jand g0205(.dina(n505),.dinb(n482),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[1]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n375_2[0]),.dinb(w_n507_1[2]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n378_2[0]),.dinb(w_G218_2[0]),.dout(n510),.clk(gclk));
	jor g0210(.dina(n510),.dinb(w_n509_0[2]),.dout(n511),.clk(gclk));
	jor g0211(.dina(n511),.dinb(w_dff_B_U8buMZBn5_1),.dout(n512),.clk(gclk));
	jand g0212(.dina(w_G3546_2[1]),.dinb(w_G218_1[2]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3548_2[0]),.dinb(w_n507_1[1]),.dout(n514),.clk(gclk));
	jor g0214(.dina(n514),.dinb(w_dff_B_R5eitxjB8_1),.dout(n515),.clk(gclk));
	jor g0215(.dina(n515),.dinb(w_G468_1[1]),.dout(n516),.clk(gclk));
	jand g0216(.dina(n516),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G257_2[1]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_n375_1[2]),.dinb(w_n518_1[2]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G389_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_n378_1[2]),.dinb(w_G257_2[0]),.dout(n521),.clk(gclk));
	jor g0221(.dina(n521),.dinb(w_n520_0[2]),.dout(n522),.clk(gclk));
	jor g0222(.dina(n522),.dinb(w_dff_B_XsWxfEym6_1),.dout(n523),.clk(gclk));
	jand g0223(.dina(w_G3546_2[0]),.dinb(w_G257_1[2]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_G3548_1[2]),.dinb(w_n518_1[1]),.dout(n525),.clk(gclk));
	jor g0225(.dina(n525),.dinb(w_dff_B_zOGq44EE9_1),.dout(n526),.clk(gclk));
	jor g0226(.dina(n526),.dinb(w_G389_1[1]),.dout(n527),.clk(gclk));
	jand g0227(.dina(n527),.dinb(n523),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[1]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G281_2[1]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n375_1[1]),.dinb(w_n530_1[2]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G374_1[2]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n378_1[1]),.dinb(w_G281_2[0]),.dout(n533),.clk(gclk));
	jor g0233(.dina(n533),.dinb(w_n532_1[1]),.dout(n534),.clk(gclk));
	jor g0234(.dina(n534),.dinb(w_dff_B_W6Ge03QS3_1),.dout(n535),.clk(gclk));
	jand g0235(.dina(w_G3546_1[2]),.dinb(w_G281_1[2]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3548_1[1]),.dinb(w_n530_1[1]),.dout(n537),.clk(gclk));
	jor g0237(.dina(n537),.dinb(w_dff_B_G5AviPzR2_1),.dout(n538),.clk(gclk));
	jor g0238(.dina(n538),.dinb(w_G374_1[1]),.dout(n539),.clk(gclk));
	jand g0239(.dina(n539),.dinb(n535),.dout(n540),.clk(gclk));
	jand g0240(.dina(w_G248_4[2]),.dinb(w_G206_1[2]),.dout(n541),.clk(gclk));
	jnot g0241(.din(w_G446_1[2]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G206_1[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_G251_4[1]),.dinb(w_n543_0[1]),.dout(n544),.clk(gclk));
	jor g0244(.dina(n544),.dinb(w_dff_B_mxxOHVf20_1),.dout(n545),.clk(gclk));
	jor g0245(.dina(n545),.dinb(w_dff_B_0MDGyf1J3_1),.dout(n546),.clk(gclk));
	jand g0246(.dina(w_n406_4[1]),.dinb(w_n543_0[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_n408_4[2]),.dinb(w_G206_1[0]),.dout(n548),.clk(gclk));
	jor g0248(.dina(n548),.dinb(n547),.dout(n549),.clk(gclk));
	jor g0249(.dina(n549),.dinb(w_G446_1[1]),.dout(n550),.clk(gclk));
	jand g0250(.dina(n550),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[2]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(n506),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_n459_0[1]),.dout(w_dff_A_nrahmVjl6_2),.clk(gclk));
	jnot g0255(.din(w_G335_0[2]),.dout(n556),.clk(gclk));
	jand g0256(.dina(w_n556_8[1]),.dinb(w_n530_1[0]),.dout(n557),.clk(gclk));
	jnot g0257(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jor g0258(.dina(w_n556_8[0]),.dinb(w_dff_B_StTsmORO0_1),.dout(n559),.clk(gclk));
	jand g0259(.dina(w_n559_0[1]),.dinb(n558),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_0[2]),.dinb(w_G374_1[0]),.dout(n561),.clk(gclk));
	jand g0261(.dina(w_n556_7[2]),.dinb(w_n471_1[0]),.dout(n562),.clk(gclk));
	jnot g0262(.din(w_n562_0[1]),.dout(n563),.clk(gclk));
	jor g0263(.dina(w_n556_7[1]),.dinb(w_dff_B_3wc4Nap28_1),.dout(n564),.clk(gclk));
	jand g0264(.dina(w_n564_0[1]),.dinb(n563),.dout(n565),.clk(gclk));
	jxor g0265(.dina(w_n565_0[2]),.dinb(w_G411_1[2]),.dout(n566),.clk(gclk));
	jand g0266(.dina(w_n566_0[2]),.dinb(w_n561_1[1]),.dout(n567),.clk(gclk));
	jnot g0267(.din(w_n567_0[2]),.dout(n568),.clk(gclk));
	jand g0268(.dina(w_n556_7[0]),.dinb(w_n483_1[2]),.dout(n569),.clk(gclk));
	jnot g0269(.din(w_n569_0[1]),.dout(n570),.clk(gclk));
	jor g0270(.dina(w_n556_6[2]),.dinb(w_dff_B_bwLRLfw68_1),.dout(n571),.clk(gclk));
	jand g0271(.dina(w_n571_0[1]),.dinb(n570),.dout(n572),.clk(gclk));
	jxor g0272(.dina(w_n572_0[2]),.dinb(w_G400_1[0]),.dout(n573),.clk(gclk));
	jnot g0273(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jand g0274(.dina(w_n556_6[1]),.dinb(w_n518_1[0]),.dout(n575),.clk(gclk));
	jnot g0275(.din(n575),.dout(n576),.clk(gclk));
	jor g0276(.dina(w_n556_6[0]),.dinb(w_dff_B_NKyFj8YE6_1),.dout(n577),.clk(gclk));
	jand g0277(.dina(w_dff_B_Fapaexz99_0),.dinb(n576),.dout(n578),.clk(gclk));
	jxor g0278(.dina(w_n578_1[1]),.dinb(w_n520_0[1]),.dout(n579),.clk(gclk));
	jor g0279(.dina(w_n579_1[1]),.dinb(w_n574_0[2]),.dout(n580),.clk(gclk));
	jor g0280(.dina(n580),.dinb(n568),.dout(n581),.clk(gclk));
	jnot g0281(.din(w_n581_0[1]),.dout(n582),.clk(gclk));
	jand g0282(.dina(w_n556_5[2]),.dinb(w_n460_1[0]),.dout(n583),.clk(gclk));
	jnot g0283(.din(n583),.dout(n584),.clk(gclk));
	jor g0284(.dina(w_n556_5[1]),.dinb(w_dff_B_Cur9DqbV8_1),.dout(n585),.clk(gclk));
	jand g0285(.dina(w_dff_B_0KfscTS83_0),.dinb(n584),.dout(n586),.clk(gclk));
	jxor g0286(.dina(w_n586_1[1]),.dinb(w_G435_1[0]),.dout(n587),.clk(gclk));
	jand g0287(.dina(w_n587_0[1]),.dinb(n582),.dout(n588),.clk(gclk));
	jor g0288(.dina(w_G335_0[1]),.dinb(w_G206_0[2]),.dout(n589),.clk(gclk));
	jor g0289(.dina(w_n556_5[0]),.dinb(w_dff_B_tzD22bHC5_1),.dout(n590),.clk(gclk));
	jand g0290(.dina(n590),.dinb(w_dff_B_jofkP0gt7_1),.dout(n591),.clk(gclk));
	jxor g0291(.dina(w_n591_1[1]),.dinb(w_G446_1[0]),.dout(n592),.clk(gclk));
	jand g0292(.dina(w_n556_4[2]),.dinb(w_n494_1[0]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jor g0294(.dina(w_n556_4[1]),.dinb(w_dff_B_Ky2Cc9Hx3_1),.dout(n595),.clk(gclk));
	jand g0295(.dina(w_dff_B_ZzFzfLkP7_0),.dinb(n594),.dout(n596),.clk(gclk));
	jxor g0296(.dina(w_n596_1[1]),.dinb(w_n496_1[0]),.dout(n597),.clk(gclk));
	jand g0297(.dina(w_n556_4[0]),.dinb(w_n507_1[0]),.dout(n598),.clk(gclk));
	jnot g0298(.din(n598),.dout(n599),.clk(gclk));
	jor g0299(.dina(w_n556_3[2]),.dinb(w_dff_B_jZXeDG7D1_1),.dout(n600),.clk(gclk));
	jand g0300(.dina(w_dff_B_sEJck0bU6_0),.dinb(n599),.dout(n601),.clk(gclk));
	jxor g0301(.dina(w_n601_1[1]),.dinb(w_n509_0[1]),.dout(n602),.clk(gclk));
	jor g0302(.dina(w_n602_0[2]),.dinb(w_n597_0[2]),.dout(n603),.clk(gclk));
	jand g0303(.dina(w_n556_3[1]),.dinb(w_n449_1[0]),.dout(n604),.clk(gclk));
	jnot g0304(.din(n604),.dout(n605),.clk(gclk));
	jor g0305(.dina(w_n556_3[0]),.dinb(w_dff_B_FNT2I8yG7_1),.dout(n606),.clk(gclk));
	jand g0306(.dina(w_dff_B_kxUpVWOD1_0),.dinb(n605),.dout(n607),.clk(gclk));
	jxor g0307(.dina(w_n607_1[1]),.dinb(w_n451_0[1]),.dout(n608),.clk(gclk));
	jor g0308(.dina(w_n608_0[2]),.dinb(w_n603_0[1]),.dout(n609),.clk(gclk));
	jnot g0309(.din(w_n609_0[2]),.dout(n610),.clk(gclk));
	jand g0310(.dina(n610),.dinb(w_n592_0[2]),.dout(n611),.clk(gclk));
	jand g0311(.dina(w_n611_0[2]),.dinb(w_n588_1[1]),.dout(w_dff_A_RHR5feu64_2),.clk(gclk));
	jnot g0312(.din(w_G332_3[2]),.dout(n613),.clk(gclk));
	jand g0313(.dina(w_n613_5[2]),.dinb(w_n435_1[2]),.dout(n614),.clk(gclk));
	jnot g0314(.din(n614),.dout(n615),.clk(gclk));
	jor g0315(.dina(w_n613_5[1]),.dinb(w_G331_0[1]),.dout(n616),.clk(gclk));
	jand g0316(.dina(w_dff_B_2P7cnQJX2_0),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_G503_1[2]),.dout(n618),.clk(gclk));
	jor g0318(.dina(w_G338_0[0]),.dinb(w_n613_5[0]),.dout(n619),.clk(gclk));
	jxor g0319(.dina(w_n619_1[2]),.dinb(w_G514_1[2]),.dout(n620),.clk(gclk));
	jor g0320(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n621),.clk(gclk));
	jor g0321(.dina(w_G348_0[0]),.dinb(w_n613_4[2]),.dout(n622),.clk(gclk));
	jand g0322(.dina(n622),.dinb(w_n621_0[1]),.dout(n623),.clk(gclk));
	jxor g0323(.dina(w_n623_0[1]),.dinb(w_G523_1[0]),.dout(n624),.clk(gclk));
	jor g0324(.dina(w_G351_1[2]),.dinb(w_G332_3[0]),.dout(n625),.clk(gclk));
	jor g0325(.dina(w_G358_0[0]),.dinb(w_n613_4[1]),.dout(n626),.clk(gclk));
	jand g0326(.dina(n626),.dinb(w_n625_0[1]),.dout(n627),.clk(gclk));
	jor g0327(.dina(w_n627_1[1]),.dinb(w_G534_1[2]),.dout(n628),.clk(gclk));
	jnot g0328(.din(w_n625_0[0]),.dout(n629),.clk(gclk));
	jand g0329(.dina(w_G612_0),.dinb(w_G332_2[2]),.dout(n630),.clk(gclk));
	jor g0330(.dina(n630),.dinb(n629),.dout(n631),.clk(gclk));
	jor g0331(.dina(w_n631_0[1]),.dinb(w_n377_1[0]),.dout(n632),.clk(gclk));
	jor g0332(.dina(w_G361_0[2]),.dinb(w_G332_2[1]),.dout(n633),.clk(gclk));
	jor g0333(.dina(w_G366_0[0]),.dinb(w_n613_4[0]),.dout(n634),.clk(gclk));
	jand g0334(.dina(n634),.dinb(w_dff_B_SfR3MZBx3_1),.dout(n635),.clk(gclk));
	jnot g0335(.din(w_n635_1[1]),.dout(n636),.clk(gclk));
	jand g0336(.dina(w_n636_0[2]),.dinb(w_n632_0[1]),.dout(n637),.clk(gclk));
	jand g0337(.dina(w_n637_0[2]),.dinb(w_n628_0[2]),.dout(n638),.clk(gclk));
	jand g0338(.dina(w_n638_0[1]),.dinb(w_n624_0[2]),.dout(n639),.clk(gclk));
	jand g0339(.dina(w_n639_0[2]),.dinb(w_n620_1[1]),.dout(n640),.clk(gclk));
	jand g0340(.dina(w_n640_0[1]),.dinb(w_n618_0[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n613_3[2]),.dinb(w_n425_0[1]),.dout(n642),.clk(gclk));
	jand g0342(.dina(w_G332_2[0]),.dinb(w_G593_0),.dout(n643),.clk(gclk));
	jor g0343(.dina(n643),.dinb(n642),.dout(n644),.clk(gclk));
	jand g0344(.dina(w_n613_3[1]),.dinb(w_n429_0[0]),.dout(n645),.clk(gclk));
	jnot g0345(.din(n645),.dout(n646),.clk(gclk));
	jor g0346(.dina(w_n613_3[0]),.dinb(w_dff_B_iK4y7oQM2_1),.dout(n647),.clk(gclk));
	jand g0347(.dina(w_dff_B_eEc63flA4_0),.dinb(n646),.dout(n648),.clk(gclk));
	jnot g0348(.din(w_n648_1[1]),.dout(n649),.clk(gclk));
	jand g0349(.dina(w_n649_0[1]),.dinb(w_n644_0[2]),.dout(n650),.clk(gclk));
	jor g0350(.dina(w_G332_1[2]),.dinb(w_G308_0[2]),.dout(n651),.clk(gclk));
	jor g0351(.dina(w_n613_2[2]),.dinb(w_dff_B_CVVTHKpS5_1),.dout(n652),.clk(gclk));
	jand g0352(.dina(n652),.dinb(w_dff_B_Q7E4iDB55_1),.dout(n653),.clk(gclk));
	jxor g0353(.dina(w_n653_0[2]),.dinb(w_G479_0[0]),.dout(n654),.clk(gclk));
	jand g0354(.dina(w_n613_2[1]),.dinb(w_n402_0[0]),.dout(n655),.clk(gclk));
	jnot g0355(.din(n655),.dout(n656),.clk(gclk));
	jor g0356(.dina(w_n613_2[0]),.dinb(w_dff_B_ZekPhHNU8_1),.dout(n657),.clk(gclk));
	jand g0357(.dina(w_dff_B_xm9n2cNj2_0),.dinb(n656),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_n658_1[1]),.dinb(w_G490_0[2]),.dout(n659),.clk(gclk));
	jand g0359(.dina(w_n659_0[1]),.dinb(w_n654_2[2]),.dout(n660),.clk(gclk));
	jand g0360(.dina(w_n660_1[1]),.dinb(w_n650_0[1]),.dout(n661),.clk(gclk));
	jand g0361(.dina(w_n661_0[1]),.dinb(w_n641_1[2]),.dout(w_dff_A_QCJjv6qE4_2),.clk(gclk));
	jxor g0362(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G302_0[0]),.dinb(w_n425_0[0]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(w_dff_B_cWFmm0rY8_1),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G369_0[1]),.dinb(w_G361_0[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(n666),.dinb(w_n435_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n668),.clk(gclk));
	jxor g0368(.dina(w_dff_B_hpGPWnPQ3_0),.dinb(n667),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n665),.dout(n670),.clk(gclk));
	jnot g0370(.din(w_n670_0[1]),.dout(w_dff_A_hM9YJ7h17_1),.clk(gclk));
	jxor g0371(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n672),.clk(gclk));
	jxor g0372(.dina(w_G273_1[1]),.dinb(w_n483_1[1]),.dout(n673),.clk(gclk));
	jxor g0373(.dina(n673),.dinb(w_dff_B_xUTfXL7O8_1),.dout(n674),.clk(gclk));
	jxor g0374(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n675),.clk(gclk));
	jxor g0375(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n676),.clk(gclk));
	jxor g0376(.dina(n676),.dinb(n675),.dout(n677),.clk(gclk));
	jxor g0377(.dina(w_G210_1[1]),.dinb(w_G206_0[1]),.dout(n678),.clk(gclk));
	jxor g0378(.dina(w_dff_B_i4RxXwLI4_0),.dinb(n677),.dout(n679),.clk(gclk));
	jxor g0379(.dina(n679),.dinb(n674),.dout(n680),.clk(gclk));
	jnot g0380(.din(w_n680_0[1]),.dout(w_dff_A_2qWiafb32_1),.clk(gclk));
	jand g0381(.dina(w_n586_1[0]),.dinb(w_G435_0[2]),.dout(n682),.clk(gclk));
	jnot g0382(.din(w_n586_0[2]),.dout(n683),.clk(gclk));
	jand g0383(.dina(n683),.dinb(w_n462_0[1]),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n684_0[1]),.dout(n685),.clk(gclk));
	jand g0385(.dina(w_n578_1[0]),.dinb(w_G389_1[0]),.dout(n686),.clk(gclk));
	jor g0386(.dina(w_n578_0[2]),.dinb(w_G389_0[2]),.dout(n687),.clk(gclk));
	jnot g0387(.din(w_n571_0[0]),.dout(n688),.clk(gclk));
	jor g0388(.dina(n688),.dinb(w_n569_0[0]),.dout(n689),.clk(gclk));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n485_1[0]),.dout(n690),.clk(gclk));
	jnot g0390(.din(w_n690_0[1]),.dout(n691),.clk(gclk));
	jand g0391(.dina(w_n560_0[1]),.dinb(w_G374_0[2]),.dout(n692),.clk(gclk));
	jor g0392(.dina(w_n565_0[1]),.dinb(w_G411_1[1]),.dout(n693),.clk(gclk));
	jand g0393(.dina(n693),.dinb(w_n692_0[1]),.dout(n694),.clk(gclk));
	jand g0394(.dina(w_n565_0[0]),.dinb(w_G411_1[0]),.dout(n695),.clk(gclk));
	jand g0395(.dina(w_n572_0[1]),.dinb(w_G400_0[2]),.dout(n696),.clk(gclk));
	jor g0396(.dina(n696),.dinb(w_n695_0[2]),.dout(n697),.clk(gclk));
	jor g0397(.dina(n697),.dinb(w_n694_0[2]),.dout(n698),.clk(gclk));
	jand g0398(.dina(n698),.dinb(w_dff_B_5KEEzPuo0_1),.dout(n699),.clk(gclk));
	jand g0399(.dina(w_n699_0[2]),.dinb(w_n687_0[1]),.dout(n700),.clk(gclk));
	jor g0400(.dina(n700),.dinb(w_n686_0[1]),.dout(n701),.clk(gclk));
	jand g0401(.dina(w_n701_0[1]),.dinb(w_n685_0[1]),.dout(n702),.clk(gclk));
	jor g0402(.dina(n702),.dinb(w_n682_0[2]),.dout(n703),.clk(gclk));
	jand g0403(.dina(w_n703_0[2]),.dinb(w_n611_0[1]),.dout(n704),.clk(gclk));
	jand g0404(.dina(w_n591_1[0]),.dinb(w_G446_0[2]),.dout(n705),.clk(gclk));
	jor g0405(.dina(w_n591_0[2]),.dinb(w_G446_0[1]),.dout(n706),.clk(gclk));
	jand g0406(.dina(w_n607_1[0]),.dinb(w_G457_1[0]),.dout(n707),.clk(gclk));
	jor g0407(.dina(w_n607_0[2]),.dinb(w_G457_0[2]),.dout(n708),.clk(gclk));
	jand g0408(.dina(w_n601_1[0]),.dinb(w_G468_1[0]),.dout(n709),.clk(gclk));
	jand g0409(.dina(w_n596_1[0]),.dinb(w_G422_0[2]),.dout(n710),.clk(gclk));
	jor g0410(.dina(w_n601_0[2]),.dinb(w_G468_0[2]),.dout(n711),.clk(gclk));
	jand g0411(.dina(w_n711_0[1]),.dinb(w_n710_0[1]),.dout(n712),.clk(gclk));
	jor g0412(.dina(n712),.dinb(w_n709_0[1]),.dout(n713),.clk(gclk));
	jand g0413(.dina(w_n713_0[2]),.dinb(w_dff_B_JjKRjUFL6_1),.dout(n714),.clk(gclk));
	jor g0414(.dina(n714),.dinb(w_dff_B_bM6Z8sTg3_1),.dout(n715),.clk(gclk));
	jand g0415(.dina(w_n715_0[2]),.dinb(w_dff_B_8ZvMHrhM6_1),.dout(n716),.clk(gclk));
	jor g0416(.dina(n716),.dinb(w_dff_B_zkPt8ae05_1),.dout(n717),.clk(gclk));
	jor g0417(.dina(w_n717_0[1]),.dinb(w_n704_0[1]),.dout(w_dff_A_wVLt2fwl5_2),.clk(gclk));
	jand g0418(.dina(w_n617_1[0]),.dinb(w_G503_1[1]),.dout(n719),.clk(gclk));
	jor g0419(.dina(w_n617_0[2]),.dinb(w_G503_1[0]),.dout(n720),.clk(gclk));
	jor g0420(.dina(w_n619_1[1]),.dinb(w_G514_1[1]),.dout(n721),.clk(gclk));
	jand g0421(.dina(w_n619_1[0]),.dinb(w_G514_1[0]),.dout(n722),.clk(gclk));
	jnot g0422(.din(w_n621_0[0]),.dout(n723),.clk(gclk));
	jand g0423(.dina(w_G599_0),.dinb(w_G332_1[1]),.dout(n724),.clk(gclk));
	jor g0424(.dina(n724),.dinb(n723),.dout(n725),.clk(gclk));
	jand g0425(.dina(w_n725_0[2]),.dinb(w_n389_1[0]),.dout(n726),.clk(gclk));
	jnot g0426(.din(w_n726_0[1]),.dout(n727),.clk(gclk));
	jand g0427(.dina(w_n635_1[0]),.dinb(w_n628_0[1]),.dout(n728),.clk(gclk));
	jand g0428(.dina(w_n623_0[0]),.dinb(w_G523_0[2]),.dout(n729),.clk(gclk));
	jand g0429(.dina(w_n627_1[0]),.dinb(w_G534_1[1]),.dout(n730),.clk(gclk));
	jor g0430(.dina(n730),.dinb(n729),.dout(n731),.clk(gclk));
	jor g0431(.dina(n731),.dinb(w_n728_0[1]),.dout(n732),.clk(gclk));
	jand g0432(.dina(n732),.dinb(w_dff_B_dUa0MRE69_1),.dout(n733),.clk(gclk));
	jor g0433(.dina(w_n733_0[2]),.dinb(w_n722_0[1]),.dout(n734),.clk(gclk));
	jand g0434(.dina(n734),.dinb(w_n721_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[2]),.dinb(w_n720_0[1]),.dout(n736),.clk(gclk));
	jor g0436(.dina(n736),.dinb(w_n719_0[1]),.dout(n737),.clk(gclk));
	jand g0437(.dina(w_n737_1[1]),.dinb(w_n660_1[0]),.dout(n738),.clk(gclk));
	jnot g0438(.din(w_n650_0[0]),.dout(n739),.clk(gclk));
	jnot g0439(.din(w_n653_0[1]),.dout(n740),.clk(gclk));
	jor g0440(.dina(n740),.dinb(w_n414_0[0]),.dout(n741),.clk(gclk));
	jand g0441(.dina(w_n658_1[0]),.dinb(w_G490_0[1]),.dout(n742),.clk(gclk));
	jand g0442(.dina(w_n742_0[2]),.dinb(w_n654_2[1]),.dout(n743),.clk(gclk));
	jnot g0443(.din(n743),.dout(n744),.clk(gclk));
	jand g0444(.dina(n744),.dinb(w_dff_B_SfwD23T13_1),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_n745_0[1]),.dout(n746),.clk(gclk));
	jor g0446(.dina(w_n746_0[2]),.dinb(w_dff_B_UHgRrhal6_1),.dout(n747),.clk(gclk));
	jor g0447(.dina(w_n747_0[1]),.dinb(w_n738_0[1]),.dout(w_dff_A_MzAOxEXW9_2),.clk(gclk));
	jnot g0448(.din(w_G4091_6[1]),.dout(n749),.clk(gclk));
	jand g0449(.dina(w_G4092_9[2]),.dinb(w_n749_13[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n750_8[2]),.dinb(w_dff_B_fRNMjkG23_1),.dout(n751),.clk(gclk));
	jnot g0451(.din(n751),.dout(n752),.clk(gclk));
	jnot g0452(.din(w_G54_0[2]),.dout(n753),.clk(gclk));
	jxor g0453(.dina(w_n635_0[2]),.dinb(w_n753_1[1]),.dout(n754),.clk(gclk));
	jnot g0454(.din(n754),.dout(n755),.clk(gclk));
	jand g0455(.dina(w_n755_0[1]),.dinb(w_G4091_6[0]),.dout(n756),.clk(gclk));
	jand g0456(.dina(w_n372_0[0]),.dinb(w_n749_13[0]),.dout(n757),.clk(gclk));
	jor g0457(.dina(n757),.dinb(w_G4092_9[1]),.dout(n758),.clk(gclk));
	jor g0458(.dina(n758),.dinb(n756),.dout(n759),.clk(gclk));
	jand g0459(.dina(n759),.dinb(w_dff_B_MpnMFYaW1_1),.dout(G822_fa_),.clk(gclk));
	jand g0460(.dina(w_n750_8[1]),.dinb(w_dff_B_BIz860tW5_1),.dout(n761),.clk(gclk));
	jnot g0461(.din(n761),.dout(n762),.clk(gclk));
	jxor g0462(.dina(w_n627_0[2]),.dinb(w_G534_1[0]),.dout(n763),.clk(gclk));
	jnot g0463(.din(w_n763_0[2]),.dout(n764),.clk(gclk));
	jand g0464(.dina(n764),.dinb(w_n635_0[1]),.dout(n765),.clk(gclk));
	jor g0465(.dina(n765),.dinb(w_n638_0[0]),.dout(n766),.clk(gclk));
	jnot g0466(.din(n766),.dout(n767),.clk(gclk));
	jand g0467(.dina(w_n767_0[1]),.dinb(w_n753_1[0]),.dout(n768),.clk(gclk));
	jand g0468(.dina(w_n763_0[1]),.dinb(w_G54_0[1]),.dout(n769),.clk(gclk));
	jor g0469(.dina(w_dff_B_fqdV4id69_0),.dinb(n768),.dout(n770),.clk(gclk));
	jand g0470(.dina(n770),.dinb(w_G4091_5[2]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n386_0[0]),.dinb(w_n749_12[2]),.dout(n772),.clk(gclk));
	jor g0472(.dina(n772),.dinb(w_G4092_9[0]),.dout(n773),.clk(gclk));
	jor g0473(.dina(w_dff_B_QreqmqU37_0),.dinb(n771),.dout(n774),.clk(gclk));
	jand g0474(.dina(n774),.dinb(w_dff_B_4w5sM2TQ6_1),.dout(G838_fa_),.clk(gclk));
	jand g0475(.dina(w_n750_8[0]),.dinb(w_dff_B_4atA8eYM2_1),.dout(n776),.clk(gclk));
	jnot g0476(.din(n776),.dout(n777),.clk(gclk));
	jxor g0477(.dina(w_n561_1[0]),.dinb(w_G4_0[2]),.dout(n778),.clk(gclk));
	jnot g0478(.din(n778),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n779_0[1]),.dinb(w_G4091_5[1]),.dout(n780),.clk(gclk));
	jand g0480(.dina(w_n540_0[0]),.dinb(w_n749_12[1]),.dout(n781),.clk(gclk));
	jor g0481(.dina(n781),.dinb(w_G4092_8[2]),.dout(n782),.clk(gclk));
	jor g0482(.dina(w_dff_B_0z2OHNJy6_0),.dinb(n780),.dout(n783),.clk(gclk));
	jand g0483(.dina(n783),.dinb(w_dff_B_wWBhILXJ6_1),.dout(G861_fa_),.clk(gclk));
	jand g0484(.dina(w_n641_1[1]),.dinb(w_G54_0[0]),.dout(n785),.clk(gclk));
	jor g0485(.dina(w_dff_B_vcCWrcpf7_0),.dinb(w_n737_1[0]),.dout(n786),.clk(gclk));
	jand g0486(.dina(w_n786_0[2]),.dinb(w_n660_0[2]),.dout(n787),.clk(gclk));
	jor g0487(.dina(n787),.dinb(w_n746_0[1]),.dout(n788),.clk(gclk));
	jnot g0488(.din(w_n788_0[2]),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n644_0[1]),.dout(n790),.clk(gclk));
	jxor g0490(.dina(w_n648_1[0]),.dinb(w_n790_0[2]),.dout(n791),.clk(gclk));
	jnot g0491(.din(n791),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_n792_0[2]),.dinb(n789),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n788_0[1]),.dinb(w_n790_0[1]),.dout(n794),.clk(gclk));
	jor g0494(.dina(w_dff_B_uoWfeqFs0_0),.dinb(n793),.dout(n795),.clk(gclk));
	jnot g0495(.din(w_n795_1[1]),.dout(G623_fa_),.clk(gclk));
	jnot g0496(.din(w_G4088_9[2]),.dout(n797),.clk(gclk));
	jnot g0497(.din(w_G861_0),.dout(n798),.clk(gclk));
	jor g0498(.dina(w_n798_1[1]),.dinb(w_n797_9[1]),.dout(n799),.clk(gclk));
	jnot g0499(.din(w_G4087_4[2]),.dout(n800),.clk(gclk));
	jnot g0500(.din(w_G822_0),.dout(n801),.clk(gclk));
	jor g0501(.dina(w_n801_1[1]),.dinb(w_G4088_9[1]),.dout(n802),.clk(gclk));
	jand g0502(.dina(n802),.dinb(w_n800_4[1]),.dout(n803),.clk(gclk));
	jand g0503(.dina(w_dff_B_mrdx43LZ1_0),.dinb(n799),.dout(n804),.clk(gclk));
	jor g0504(.dina(w_n797_9[0]),.dinb(w_G61_0[1]),.dout(n805),.clk(gclk));
	jor g0505(.dina(w_G4088_9[0]),.dinb(w_G11_0[1]),.dout(n806),.clk(gclk));
	jand g0506(.dina(n806),.dinb(w_G4087_4[1]),.dout(n807),.clk(gclk));
	jand g0507(.dina(n807),.dinb(n805),.dout(n808),.clk(gclk));
	jor g0508(.dina(w_dff_B_RxKT6oOM6_0),.dinb(n804),.dout(w_dff_A_GoqX3tdp4_2),.clk(gclk));
	jand g0509(.dina(w_n750_7[2]),.dinb(w_dff_B_E1lXjz2A0_1),.dout(n810),.clk(gclk));
	jnot g0510(.din(n810),.dout(n811),.clk(gclk));
	jnot g0511(.din(w_n721_0[0]),.dout(n812),.clk(gclk));
	jnot g0512(.din(w_n722_0[0]),.dout(n813),.clk(gclk));
	jand g0513(.dina(w_n631_0[0]),.dinb(w_n377_0[2]),.dout(n814),.clk(gclk));
	jor g0514(.dina(w_n636_0[1]),.dinb(w_n814_0[2]),.dout(n815),.clk(gclk));
	jor g0515(.dina(w_n725_0[1]),.dinb(w_n389_0[2]),.dout(n816),.clk(gclk));
	jand g0516(.dina(w_n632_0[0]),.dinb(n816),.dout(n817),.clk(gclk));
	jand g0517(.dina(n817),.dinb(n815),.dout(n818),.clk(gclk));
	jor g0518(.dina(n818),.dinb(w_n726_0[0]),.dout(n819),.clk(gclk));
	jand g0519(.dina(w_n819_0[2]),.dinb(w_dff_B_pKbLoEhn9_1),.dout(n820),.clk(gclk));
	jor g0520(.dina(n820),.dinb(w_dff_B_CS9FX0KI7_1),.dout(n821),.clk(gclk));
	jnot g0521(.din(w_n620_1[0]),.dout(n822),.clk(gclk));
	jnot g0522(.din(w_n639_0[1]),.dout(n823),.clk(gclk));
	jor g0523(.dina(n823),.dinb(w_n753_0[2]),.dout(n824),.clk(gclk));
	jor g0524(.dina(w_n824_0[1]),.dinb(w_dff_B_xAtnCFNh5_1),.dout(n825),.clk(gclk));
	jand g0525(.dina(n825),.dinb(w_n821_0[1]),.dout(n826),.clk(gclk));
	jxor g0526(.dina(n826),.dinb(w_n618_0[1]),.dout(n827),.clk(gclk));
	jand g0527(.dina(w_n827_0[1]),.dinb(w_G4091_5[0]),.dout(n828),.clk(gclk));
	jand g0528(.dina(w_n445_0[0]),.dinb(w_n749_12[0]),.dout(n829),.clk(gclk));
	jor g0529(.dina(n829),.dinb(w_G4092_8[1]),.dout(n830),.clk(gclk));
	jor g0530(.dina(w_dff_B_UIS0n0cy6_0),.dinb(n828),.dout(n831),.clk(gclk));
	jand g0531(.dina(n831),.dinb(w_dff_B_4eTKlpJq8_1),.dout(G832_fa_),.clk(gclk));
	jand g0532(.dina(w_n750_7[1]),.dinb(w_dff_B_JVMS83W53_1),.dout(n833),.clk(gclk));
	jnot g0533(.din(n833),.dout(n834),.clk(gclk));
	jand g0534(.dina(w_n824_0[0]),.dinb(w_n819_0[1]),.dout(n835),.clk(gclk));
	jxor g0535(.dina(n835),.dinb(w_n620_0[2]),.dout(n836),.clk(gclk));
	jand g0536(.dina(w_n836_0[1]),.dinb(w_G4091_4[2]),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_n365_0[0]),.dinb(w_n749_11[2]),.dout(n838),.clk(gclk));
	jor g0538(.dina(n838),.dinb(w_G4092_8[0]),.dout(n839),.clk(gclk));
	jor g0539(.dina(w_dff_B_ztQca1h34_0),.dinb(n837),.dout(n840),.clk(gclk));
	jand g0540(.dina(n840),.dinb(w_dff_B_Kz64QH1X3_1),.dout(G834_fa_),.clk(gclk));
	jand g0541(.dina(w_n750_7[0]),.dinb(w_dff_B_YHnInmKb8_1),.dout(n842),.clk(gclk));
	jnot g0542(.din(n842),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n397_0[0]),.dinb(w_n749_11[1]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_n637_0[1]),.dinb(w_n753_0[1]),.dout(n845),.clk(gclk));
	jor g0545(.dina(n845),.dinb(w_n814_0[1]),.dout(n846),.clk(gclk));
	jxor g0546(.dina(n846),.dinb(w_n624_0[1]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_0[1]),.dinb(w_G4091_4[1]),.dout(n848),.clk(gclk));
	jor g0548(.dina(n848),.dinb(w_G4092_7[2]),.dout(n849),.clk(gclk));
	jor g0549(.dina(n849),.dinb(w_dff_B_g0gNCxJa4_1),.dout(n850),.clk(gclk));
	jand g0550(.dina(n850),.dinb(w_dff_B_tkO5Zrls7_1),.dout(G836_fa_),.clk(gclk));
	jnot g0551(.din(w_G4089_9[2]),.dout(n852),.clk(gclk));
	jor g0552(.dina(w_n798_1[0]),.dinb(w_n852_9[1]),.dout(n853),.clk(gclk));
	jnot g0553(.din(w_G4090_4[2]),.dout(n854),.clk(gclk));
	jor g0554(.dina(w_n801_1[0]),.dinb(w_G4089_9[1]),.dout(n855),.clk(gclk));
	jand g0555(.dina(n855),.dinb(w_n854_4[1]),.dout(n856),.clk(gclk));
	jand g0556(.dina(w_dff_B_fDqSVZGS8_0),.dinb(n853),.dout(n857),.clk(gclk));
	jor g0557(.dina(w_n852_9[0]),.dinb(w_G61_0[0]),.dout(n858),.clk(gclk));
	jor g0558(.dina(w_G4089_9[0]),.dinb(w_G11_0[0]),.dout(n859),.clk(gclk));
	jand g0559(.dina(n859),.dinb(w_G4090_4[1]),.dout(n860),.clk(gclk));
	jand g0560(.dina(n860),.dinb(n858),.dout(n861),.clk(gclk));
	jor g0561(.dina(w_dff_B_qqeTdjm71_0),.dinb(n857),.dout(w_dff_A_P2qeWm9N7_2),.clk(gclk));
	jand g0562(.dina(w_n750_6[2]),.dinb(w_dff_B_G7WvKJ7j7_1),.dout(n863),.clk(gclk));
	jnot g0563(.din(n863),.dout(n864),.clk(gclk));
	jnot g0564(.din(w_n587_0[0]),.dout(n865),.clk(gclk));
	jnot g0565(.din(w_n579_1[0]),.dout(n866),.clk(gclk));
	jand g0566(.dina(w_n567_0[1]),.dinb(w_G4_0[1]),.dout(n867),.clk(gclk));
	jand g0567(.dina(w_n867_0[1]),.dinb(w_n573_0[1]),.dout(n868),.clk(gclk));
	jand g0568(.dina(w_n868_0[1]),.dinb(w_dff_B_SZmFmjq37_1),.dout(n869),.clk(gclk));
	jor g0569(.dina(w_dff_B_2GHUucvT0_0),.dinb(w_n701_0[0]),.dout(n870),.clk(gclk));
	jxor g0570(.dina(w_n870_0[1]),.dinb(w_n865_0[2]),.dout(n871),.clk(gclk));
	jand g0571(.dina(w_n871_0[1]),.dinb(w_G4091_4[0]),.dout(n872),.clk(gclk));
	jand g0572(.dina(w_n470_0[0]),.dinb(w_n749_11[0]),.dout(n873),.clk(gclk));
	jor g0573(.dina(n873),.dinb(w_G4092_7[1]),.dout(n874),.clk(gclk));
	jor g0574(.dina(w_dff_B_WLwaQdrP9_0),.dinb(n872),.dout(n875),.clk(gclk));
	jand g0575(.dina(n875),.dinb(w_dff_B_bhV7aBCh0_1),.dout(G871_fa_),.clk(gclk));
	jand g0576(.dina(w_n750_6[1]),.dinb(w_dff_B_ztXtA0sx5_1),.dout(n877),.clk(gclk));
	jnot g0577(.din(n877),.dout(n878),.clk(gclk));
	jor g0578(.dina(w_n868_0[0]),.dinb(w_n699_0[1]),.dout(n879),.clk(gclk));
	jxor g0579(.dina(n879),.dinb(w_n579_0[2]),.dout(n880),.clk(gclk));
	jand g0580(.dina(w_n880_0[1]),.dinb(w_G4091_3[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n528_0[0]),.dinb(w_n749_10[2]),.dout(n882),.clk(gclk));
	jor g0582(.dina(n882),.dinb(w_G4092_7[0]),.dout(n883),.clk(gclk));
	jor g0583(.dina(w_dff_B_V3cGInGs1_0),.dinb(n881),.dout(n884),.clk(gclk));
	jand g0584(.dina(n884),.dinb(w_dff_B_nuJyNRVB7_1),.dout(G873_fa_),.clk(gclk));
	jand g0585(.dina(w_n750_6[0]),.dinb(w_dff_B_TVfQ4Pp23_1),.dout(n886),.clk(gclk));
	jnot g0586(.din(n886),.dout(n887),.clk(gclk));
	jor g0587(.dina(w_n694_0[1]),.dinb(w_n695_0[1]),.dout(n888),.clk(gclk));
	jor g0588(.dina(n888),.dinb(w_n867_0[0]),.dout(n889),.clk(gclk));
	jxor g0589(.dina(n889),.dinb(w_n574_0[1]),.dout(n890),.clk(gclk));
	jand g0590(.dina(w_n890_0[1]),.dinb(w_G4091_3[1]),.dout(n891),.clk(gclk));
	jand g0591(.dina(w_n493_0[0]),.dinb(w_n749_10[1]),.dout(n892),.clk(gclk));
	jor g0592(.dina(n892),.dinb(w_G4092_6[2]),.dout(n893),.clk(gclk));
	jor g0593(.dina(w_dff_B_Uja55WdY4_0),.dinb(n891),.dout(n894),.clk(gclk));
	jand g0594(.dina(n894),.dinb(w_dff_B_0ObkkvA53_1),.dout(G875_fa_),.clk(gclk));
	jand g0595(.dina(w_n750_5[2]),.dinb(w_dff_B_IX2dHluj9_1),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jnot g0597(.din(w_n566_0[1]),.dout(n898),.clk(gclk));
	jand g0598(.dina(w_n561_0[2]),.dinb(w_G4_0[0]),.dout(n899),.clk(gclk));
	jor g0599(.dina(n899),.dinb(w_n692_0[0]),.dout(n900),.clk(gclk));
	jxor g0600(.dina(n900),.dinb(w_dff_B_0JWCdQHO9_1),.dout(n901),.clk(gclk));
	jand g0601(.dina(w_n901_0[1]),.dinb(w_G4091_3[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_n481_0[0]),.dinb(w_n749_10[0]),.dout(n903),.clk(gclk));
	jor g0603(.dina(n903),.dinb(w_G4092_6[1]),.dout(n904),.clk(gclk));
	jor g0604(.dina(w_dff_B_i3OubGyD6_0),.dinb(n902),.dout(n905),.clk(gclk));
	jand g0605(.dina(n905),.dinb(w_dff_B_Nwaz4MU14_1),.dout(G877_fa_),.clk(gclk));
	jnot g0606(.din(w_G331_0[0]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_n619_0[2]),.dout(n908),.clk(gclk));
	jand g0608(.dina(n908),.dinb(w_dff_B_l0ah2yuI1_1),.dout(n909),.clk(gclk));
	jand g0609(.dina(w_n619_0[1]),.dinb(w_n617_0[1]),.dout(n910),.clk(gclk));
	jor g0610(.dina(n910),.dinb(w_dff_B_wEjuJzkp5_1),.dout(n911),.clk(gclk));
	jxor g0611(.dina(n911),.dinb(w_n792_0[1]),.dout(n912),.clk(gclk));
	jor g0612(.dina(w_G369_0[0]),.dinb(w_G332_1[0]),.dout(n913),.clk(gclk));
	jor g0613(.dina(w_dff_B_WrvP5RP93_0),.dinb(w_n613_1[2]),.dout(n914),.clk(gclk));
	jand g0614(.dina(n914),.dinb(w_dff_B_6nFQBuEi0_1),.dout(n915),.clk(gclk));
	jxor g0615(.dina(w_dff_B_jYQ8yJpf9_0),.dinb(w_n636_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n627_0[1]),.dinb(w_n725_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(w_n658_0[2]),.dinb(w_n653_0[0]),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_dff_B_ZGC8ArjM6_1),.dout(n919),.clk(gclk));
	jxor g0619(.dina(n919),.dinb(w_dff_B_NKzmPQCu8_1),.dout(n920),.clk(gclk));
	jxor g0620(.dina(n920),.dinb(n912),.dout(G998_fa_),.clk(gclk));
	jnot g0621(.din(w_n564_0[0]),.dout(n922),.clk(gclk));
	jor g0622(.dina(n922),.dinb(w_n562_0[0]),.dout(n923),.clk(gclk));
	jxor g0623(.dina(w_n578_0[1]),.dinb(w_n923_0[2]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n572_0[0]),.dinb(w_n560_0[0]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jor g0626(.dina(w_G335_0[0]),.dinb(w_G289_0[0]),.dout(n927),.clk(gclk));
	jor g0627(.dina(w_n556_2[2]),.dinb(w_dff_B_0pyGS53w1_1),.dout(n928),.clk(gclk));
	jand g0628(.dina(n928),.dinb(w_dff_B_SkgBOMHA8_1),.dout(n929),.clk(gclk));
	jxor g0629(.dina(n929),.dinb(w_n591_0[1]),.dout(n930),.clk(gclk));
	jxor g0630(.dina(w_n596_0[2]),.dinb(w_n586_0[1]),.dout(n931),.clk(gclk));
	jxor g0631(.dina(w_n607_0[1]),.dinb(w_n601_0[1]),.dout(n932),.clk(gclk));
	jxor g0632(.dina(n932),.dinb(n931),.dout(n933),.clk(gclk));
	jxor g0633(.dina(n933),.dinb(w_dff_B_5BGTfmIR1_1),.dout(n934),.clk(gclk));
	jxor g0634(.dina(n934),.dinb(w_dff_B_SIK51O1X2_1),.dout(n935),.clk(gclk));
	jnot g0635(.din(w_n935_0[1]),.dout(w_dff_A_KTZtqfg71_1),.clk(gclk));
	jnot g0636(.din(w_n592_0[1]),.dout(n937),.clk(gclk));
	jnot g0637(.din(w_n715_0[1]),.dout(n938),.clk(gclk));
	jor g0638(.dina(w_n870_0[0]),.dinb(w_n682_0[1]),.dout(n939),.clk(gclk));
	jand g0639(.dina(n939),.dinb(w_n685_0[0]),.dout(n940),.clk(gclk));
	jnot g0640(.din(w_n940_1[1]),.dout(n941),.clk(gclk));
	jor g0641(.dina(n941),.dinb(w_n609_0[1]),.dout(n942),.clk(gclk));
	jand g0642(.dina(n942),.dinb(w_n938_0[2]),.dout(n943),.clk(gclk));
	jxor g0643(.dina(n943),.dinb(w_dff_B_Q5gAEA4b4_1),.dout(n944),.clk(gclk));
	jnot g0644(.din(w_n944_0[1]),.dout(n945),.clk(gclk));
	jnot g0645(.din(w_n603_0[0]),.dout(n946),.clk(gclk));
	jand g0646(.dina(w_n940_1[0]),.dinb(w_dff_B_pvf6Qcwc9_1),.dout(n947),.clk(gclk));
	jor g0647(.dina(n947),.dinb(w_n713_0[1]),.dout(n948),.clk(gclk));
	jxor g0648(.dina(n948),.dinb(w_n608_0[1]),.dout(n949),.clk(gclk));
	jand g0649(.dina(w_n949_0[1]),.dinb(n945),.dout(n950),.clk(gclk));
	jnot g0650(.din(w_n602_0[1]),.dout(n951),.clk(gclk));
	jnot g0651(.din(w_n596_0[1]),.dout(n952),.clk(gclk));
	jand g0652(.dina(n952),.dinb(w_n496_0[2]),.dout(n953),.clk(gclk));
	jnot g0653(.din(w_n953_0[1]),.dout(n954),.clk(gclk));
	jor g0654(.dina(w_n940_0[2]),.dinb(w_n710_0[0]),.dout(n955),.clk(gclk));
	jand g0655(.dina(n955),.dinb(w_n954_0[2]),.dout(n956),.clk(gclk));
	jxor g0656(.dina(n956),.dinb(w_dff_B_U77XHhe59_1),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n957_0[1]),.dout(n958),.clk(gclk));
	jand g0658(.dina(w_n890_0[0]),.dinb(w_n779_0[0]),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(w_n901_0[0]),.dout(n960),.clk(gclk));
	jand g0660(.dina(w_dff_B_ma5VyXQF8_0),.dinb(w_n871_0[0]),.dout(n961),.clk(gclk));
	jnot g0661(.din(w_n597_0[1]),.dout(n962),.clk(gclk));
	jxor g0662(.dina(w_n940_0[1]),.dinb(w_n962_0[1]),.dout(n963),.clk(gclk));
	jnot g0663(.din(n963),.dout(n964),.clk(gclk));
	jand g0664(.dina(w_n964_0[1]),.dinb(w_n880_0[0]),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(w_dff_B_F93TvI0b1_1),.dout(n966),.clk(gclk));
	jand g0666(.dina(n966),.dinb(n958),.dout(n967),.clk(gclk));
	jand g0667(.dina(w_dff_B_mvtfbOKG2_0),.dinb(n950),.dout(w_dff_A_oFxVWF266_2),.clk(gclk));
	jxor g0668(.dina(w_n788_0[0]),.dinb(w_n649_0[0]),.dout(n969),.clk(gclk));
	jnot g0669(.din(w_n969_0[1]),.dout(n970),.clk(gclk));
	jand g0670(.dina(n970),.dinb(w_n755_0[0]),.dout(n971),.clk(gclk));
	jand g0671(.dina(w_n836_0[0]),.dinb(w_G623_0),.dout(n972),.clk(gclk));
	jand g0672(.dina(n972),.dinb(w_dff_B_WvPKT57L9_1),.dout(n973),.clk(gclk));
	jand g0673(.dina(w_n827_0[0]),.dinb(w_n763_0[0]),.dout(n974),.clk(gclk));
	jand g0674(.dina(n974),.dinb(w_n847_0[0]),.dout(n975),.clk(gclk));
	jnot g0675(.din(w_n658_0[1]),.dout(n976),.clk(gclk));
	jand g0676(.dina(n976),.dinb(w_n401_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(w_n977_0[2]),.dinb(w_n654_2[0]),.dout(n978),.clk(gclk));
	jor g0678(.dina(w_n977_0[1]),.dinb(w_n654_1[2]),.dout(n979),.clk(gclk));
	jnot g0679(.din(n979),.dout(n980),.clk(gclk));
	jor g0680(.dina(w_n786_0[1]),.dinb(w_n742_0[1]),.dout(n981),.clk(gclk));
	jand g0681(.dina(w_n981_0[1]),.dinb(w_dff_B_N4OMMBhQ3_1),.dout(n982),.clk(gclk));
	jnot g0682(.din(w_n981_0[0]),.dout(n983),.clk(gclk));
	jand g0683(.dina(n983),.dinb(w_n654_1[1]),.dout(n984),.clk(gclk));
	jor g0684(.dina(n984),.dinb(w_dff_B_0ALb2b7X8_1),.dout(n985),.clk(gclk));
	jor g0685(.dina(n985),.dinb(w_dff_B_evwuM9UD2_1),.dout(n986),.clk(gclk));
	jnot g0686(.din(w_n986_0[1]),.dout(n987),.clk(gclk));
	jnot g0687(.din(w_n659_0[0]),.dout(n988),.clk(gclk));
	jxor g0688(.dina(w_n786_0[0]),.dinb(w_dff_B_9D7e0xVP8_1),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_n989_0[1]),.dinb(n987),.dout(n990),.clk(gclk));
	jand g0690(.dina(n990),.dinb(w_dff_B_vBhC3C0o8_1),.dout(n991),.clk(gclk));
	jand g0691(.dina(n991),.dinb(n973),.dout(w_dff_A_eSkGMLfB8_2),.clk(gclk));
	jnot g0692(.din(w_G1689_5[1]),.dout(n993),.clk(gclk));
	jand g0693(.dina(w_G1690_1[1]),.dinb(w_n993_4[2]),.dout(n994),.clk(gclk));
	jand g0694(.dina(w_n994_4[1]),.dinb(w_G182_0[1]),.dout(n995),.clk(gclk));
	jand g0695(.dina(w_G1690_1[0]),.dinb(w_G1689_5[0]),.dout(n996),.clk(gclk));
	jand g0696(.dina(w_n996_4[1]),.dinb(w_G185_0[1]),.dout(n997),.clk(gclk));
	jor g0697(.dina(w_n798_0[2]),.dinb(w_n993_4[1]),.dout(n998),.clk(gclk));
	jnot g0698(.din(w_G1690_0[2]),.dout(n999),.clk(gclk));
	jor g0699(.dina(w_n801_0[2]),.dinb(w_G1689_4[2]),.dout(n1000),.clk(gclk));
	jand g0700(.dina(n1000),.dinb(w_n999_3[2]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_dff_B_pD7lTEdd0_0),.dinb(n998),.dout(n1002),.clk(gclk));
	jor g0702(.dina(n1002),.dinb(w_dff_B_k6SjvXSa7_1),.dout(n1003),.clk(gclk));
	jor g0703(.dina(n1003),.dinb(w_dff_B_F3veK4cD5_1),.dout(n1004),.clk(gclk));
	jand g0704(.dina(n1004),.dinb(w_G137_9[1]),.dout(w_dff_A_IUyZibeU2_2),.clk(gclk));
	jor g0705(.dina(w_n801_0[1]),.dinb(w_G1691_5[1]),.dout(n1006),.clk(gclk));
	jnot g0706(.din(w_G1694_1[1]),.dout(n1007),.clk(gclk));
	jnot g0707(.din(w_G1691_5[0]),.dout(n1008),.clk(gclk));
	jor g0708(.dina(w_n798_0[1]),.dinb(w_n1008_4[2]),.dout(n1009),.clk(gclk));
	jand g0709(.dina(n1009),.dinb(w_n1007_3[2]),.dout(n1010),.clk(gclk));
	jand g0710(.dina(n1010),.dinb(w_dff_B_VRgdXbNk2_1),.dout(n1011),.clk(gclk));
	jand g0711(.dina(w_G1694_1[0]),.dinb(w_G1691_4[2]),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_4[1]),.dinb(w_G185_0[0]),.dout(n1013),.clk(gclk));
	jand g0713(.dina(w_G1694_0[2]),.dinb(w_n1008_4[1]),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_4[1]),.dinb(w_G182_0[0]),.dout(n1015),.clk(gclk));
	jor g0715(.dina(n1015),.dinb(w_dff_B_f2GERJv18_1),.dout(n1016),.clk(gclk));
	jor g0716(.dina(w_dff_B_2MIFHDv32_0),.dinb(n1011),.dout(n1017),.clk(gclk));
	jand g0717(.dina(n1017),.dinb(w_G137_9[0]),.dout(w_dff_A_cL0EQVCg1_2),.clk(gclk));
	jnot g0718(.din(w_G871_0),.dout(n1019),.clk(gclk));
	jor g0719(.dina(w_n1019_1[1]),.dinb(w_n797_8[2]),.dout(n1020),.clk(gclk));
	jnot g0720(.din(w_G832_0),.dout(n1021),.clk(gclk));
	jor g0721(.dina(w_n1021_1[1]),.dinb(w_G4088_8[2]),.dout(n1022),.clk(gclk));
	jand g0722(.dina(n1022),.dinb(w_n800_4[0]),.dout(n1023),.clk(gclk));
	jand g0723(.dina(n1023),.dinb(w_dff_B_neTZGdA48_1),.dout(n1024),.clk(gclk));
	jor g0724(.dina(w_n797_8[1]),.dinb(w_G37_0[1]),.dout(n1025),.clk(gclk));
	jor g0725(.dina(w_G4088_8[1]),.dinb(w_G43_0[1]),.dout(n1026),.clk(gclk));
	jand g0726(.dina(n1026),.dinb(w_G4087_4[0]),.dout(n1027),.clk(gclk));
	jand g0727(.dina(n1027),.dinb(n1025),.dout(n1028),.clk(gclk));
	jor g0728(.dina(w_dff_B_5gqfWVpb8_0),.dinb(n1024),.dout(w_dff_A_IGyoSSEu8_2),.clk(gclk));
	jnot g0729(.din(w_G873_0),.dout(n1030),.clk(gclk));
	jor g0730(.dina(w_n1030_1[1]),.dinb(w_n797_8[0]),.dout(n1031),.clk(gclk));
	jnot g0731(.din(w_G834_0),.dout(n1032),.clk(gclk));
	jor g0732(.dina(w_n1032_1[1]),.dinb(w_G4088_8[0]),.dout(n1033),.clk(gclk));
	jand g0733(.dina(n1033),.dinb(w_n800_3[2]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(n1034),.dinb(w_dff_B_Cgqz8Wrk5_1),.dout(n1035),.clk(gclk));
	jor g0735(.dina(w_n797_7[2]),.dinb(w_G20_0[1]),.dout(n1036),.clk(gclk));
	jor g0736(.dina(w_G4088_7[2]),.dinb(w_G76_0[1]),.dout(n1037),.clk(gclk));
	jand g0737(.dina(n1037),.dinb(w_G4087_3[2]),.dout(n1038),.clk(gclk));
	jand g0738(.dina(n1038),.dinb(n1036),.dout(n1039),.clk(gclk));
	jor g0739(.dina(w_dff_B_lUb34adj1_0),.dinb(n1035),.dout(w_dff_A_56RrwCqu2_2),.clk(gclk));
	jnot g0740(.din(w_G836_0),.dout(n1041),.clk(gclk));
	jor g0741(.dina(w_n1041_1[1]),.dinb(w_G4088_7[1]),.dout(n1042),.clk(gclk));
	jnot g0742(.din(w_G875_0),.dout(n1043),.clk(gclk));
	jor g0743(.dina(w_n1043_1[1]),.dinb(w_n797_7[1]),.dout(n1044),.clk(gclk));
	jand g0744(.dina(n1044),.dinb(w_n800_3[1]),.dout(n1045),.clk(gclk));
	jand g0745(.dina(n1045),.dinb(w_dff_B_1CWlwn4L5_1),.dout(n1046),.clk(gclk));
	jor g0746(.dina(w_n797_7[0]),.dinb(w_G17_0[1]),.dout(n1047),.clk(gclk));
	jor g0747(.dina(w_G4088_7[0]),.dinb(w_G73_0[1]),.dout(n1048),.clk(gclk));
	jand g0748(.dina(n1048),.dinb(w_G4087_3[1]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(n1049),.dinb(n1047),.dout(n1050),.clk(gclk));
	jor g0750(.dina(w_dff_B_vv8Jq0650_0),.dinb(n1046),.dout(w_dff_A_wwQGevd50_2),.clk(gclk));
	jnot g0751(.din(w_G877_0),.dout(n1052),.clk(gclk));
	jor g0752(.dina(w_n1052_1[1]),.dinb(w_n797_6[2]),.dout(n1053),.clk(gclk));
	jnot g0753(.din(w_G838_0),.dout(n1054),.clk(gclk));
	jor g0754(.dina(w_n1054_1[1]),.dinb(w_G4088_6[2]),.dout(n1055),.clk(gclk));
	jand g0755(.dina(n1055),.dinb(w_n800_3[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(n1056),.dinb(w_dff_B_CFdtmdKf5_1),.dout(n1057),.clk(gclk));
	jor g0757(.dina(w_n797_6[1]),.dinb(w_G70_0[1]),.dout(n1058),.clk(gclk));
	jor g0758(.dina(w_G4088_6[1]),.dinb(w_G67_0[1]),.dout(n1059),.clk(gclk));
	jand g0759(.dina(n1059),.dinb(w_G4087_3[0]),.dout(n1060),.clk(gclk));
	jand g0760(.dina(n1060),.dinb(n1058),.dout(n1061),.clk(gclk));
	jor g0761(.dina(w_dff_B_lGrJQWgO6_0),.dinb(n1057),.dout(w_dff_A_keQaPtPi2_2),.clk(gclk));
	jor g0762(.dina(w_G4089_8[2]),.dinb(w_G43_0[0]),.dout(n1063),.clk(gclk));
	jor g0763(.dina(w_n852_8[2]),.dinb(w_G37_0[0]),.dout(n1064),.clk(gclk));
	jand g0764(.dina(n1064),.dinb(w_G4090_4[0]),.dout(n1065),.clk(gclk));
	jand g0765(.dina(n1065),.dinb(w_dff_B_B0CHzlMz8_1),.dout(n1066),.clk(gclk));
	jor g0766(.dina(w_n1021_1[0]),.dinb(w_G4089_8[1]),.dout(n1067),.clk(gclk));
	jor g0767(.dina(w_n1019_1[0]),.dinb(w_n852_8[1]),.dout(n1068),.clk(gclk));
	jand g0768(.dina(n1068),.dinb(n1067),.dout(n1069),.clk(gclk));
	jand g0769(.dina(n1069),.dinb(w_n854_4[0]),.dout(n1070),.clk(gclk));
	jor g0770(.dina(n1070),.dinb(w_dff_B_R05Mb3Zj5_1),.dout(w_dff_A_7oyN7Kg98_2),.clk(gclk));
	jor g0771(.dina(w_G4089_8[0]),.dinb(w_G76_0[0]),.dout(n1072),.clk(gclk));
	jor g0772(.dina(w_n852_8[0]),.dinb(w_G20_0[0]),.dout(n1073),.clk(gclk));
	jand g0773(.dina(n1073),.dinb(w_G4090_3[2]),.dout(n1074),.clk(gclk));
	jand g0774(.dina(n1074),.dinb(w_dff_B_0rjRKGPo7_1),.dout(n1075),.clk(gclk));
	jor g0775(.dina(w_n1032_1[0]),.dinb(w_G4089_7[2]),.dout(n1076),.clk(gclk));
	jor g0776(.dina(w_n1030_1[0]),.dinb(w_n852_7[2]),.dout(n1077),.clk(gclk));
	jand g0777(.dina(w_dff_B_Lb1UTJyr6_0),.dinb(n1076),.dout(n1078),.clk(gclk));
	jand g0778(.dina(n1078),.dinb(w_n854_3[2]),.dout(n1079),.clk(gclk));
	jor g0779(.dina(n1079),.dinb(w_dff_B_LimWu8Tx3_1),.dout(w_dff_A_HwrRny5T3_2),.clk(gclk));
	jor g0780(.dina(w_G4089_7[1]),.dinb(w_G73_0[0]),.dout(n1081),.clk(gclk));
	jor g0781(.dina(w_n852_7[1]),.dinb(w_G17_0[0]),.dout(n1082),.clk(gclk));
	jand g0782(.dina(n1082),.dinb(w_G4090_3[1]),.dout(n1083),.clk(gclk));
	jand g0783(.dina(n1083),.dinb(w_dff_B_KOtNylFL9_1),.dout(n1084),.clk(gclk));
	jor g0784(.dina(w_n1043_1[0]),.dinb(w_n852_7[0]),.dout(n1085),.clk(gclk));
	jor g0785(.dina(w_n1041_1[0]),.dinb(w_G4089_7[0]),.dout(n1086),.clk(gclk));
	jand g0786(.dina(n1086),.dinb(n1085),.dout(n1087),.clk(gclk));
	jand g0787(.dina(n1087),.dinb(w_n854_3[1]),.dout(n1088),.clk(gclk));
	jor g0788(.dina(n1088),.dinb(w_dff_B_4iclhfl35_1),.dout(w_dff_A_hBJRCEio6_2),.clk(gclk));
	jor g0789(.dina(w_n1052_1[0]),.dinb(w_n852_6[2]),.dout(n1090),.clk(gclk));
	jor g0790(.dina(w_n1054_1[0]),.dinb(w_G4089_6[2]),.dout(n1091),.clk(gclk));
	jand g0791(.dina(n1091),.dinb(w_n854_3[0]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(n1092),.dinb(w_dff_B_w7zKmeRY0_1),.dout(n1093),.clk(gclk));
	jor g0793(.dina(w_n852_6[1]),.dinb(w_G70_0[0]),.dout(n1094),.clk(gclk));
	jor g0794(.dina(w_G4089_6[1]),.dinb(w_G67_0[0]),.dout(n1095),.clk(gclk));
	jand g0795(.dina(n1095),.dinb(w_G4090_3[0]),.dout(n1096),.clk(gclk));
	jand g0796(.dina(n1096),.dinb(n1094),.dout(n1097),.clk(gclk));
	jor g0797(.dina(w_dff_B_vohdLkQS8_0),.dinb(n1093),.dout(w_dff_A_kRGQhKKq4_2),.clk(gclk));
	jor g0798(.dina(w_n1021_0[2]),.dinb(w_G1689_4[1]),.dout(n1099),.clk(gclk));
	jor g0799(.dina(w_n1019_0[2]),.dinb(w_n993_4[0]),.dout(n1100),.clk(gclk));
	jand g0800(.dina(n1100),.dinb(w_n999_3[1]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(n1101),.dinb(w_dff_B_YTrvBkwS9_1),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n994_4[0]),.dinb(w_G200_0[1]),.dout(n1103),.clk(gclk));
	jand g0803(.dina(w_n996_4[0]),.dinb(w_G170_0[1]),.dout(n1104),.clk(gclk));
	jor g0804(.dina(w_dff_B_uHtD4vlp5_0),.dinb(n1103),.dout(n1105),.clk(gclk));
	jor g0805(.dina(w_dff_B_whG8IqYl2_0),.dinb(n1102),.dout(n1106),.clk(gclk));
	jand g0806(.dina(n1106),.dinb(w_G137_8[2]),.dout(w_dff_A_wjAAGGZN0_2),.clk(gclk));
	jor g0807(.dina(w_n1054_0[2]),.dinb(w_G1689_4[0]),.dout(n1108),.clk(gclk));
	jor g0808(.dina(w_n1052_0[2]),.dinb(w_n993_3[2]),.dout(n1109),.clk(gclk));
	jand g0809(.dina(n1109),.dinb(w_n999_3[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(w_dff_B_jKbWAgBq6_0),.dinb(n1108),.dout(n1111),.clk(gclk));
	jand g0811(.dina(w_n994_3[2]),.dinb(w_G188_0[1]),.dout(n1112),.clk(gclk));
	jand g0812(.dina(w_n996_3[2]),.dinb(w_G158_0[1]),.dout(n1113),.clk(gclk));
	jor g0813(.dina(w_dff_B_01lO3jCx5_0),.dinb(n1112),.dout(n1114),.clk(gclk));
	jor g0814(.dina(w_dff_B_EiX5KooM5_0),.dinb(n1111),.dout(n1115),.clk(gclk));
	jand g0815(.dina(n1115),.dinb(w_G137_8[1]),.dout(w_dff_A_kbovglEb0_2),.clk(gclk));
	jor g0816(.dina(w_n1041_0[2]),.dinb(w_G1689_3[2]),.dout(n1117),.clk(gclk));
	jor g0817(.dina(w_n1043_0[2]),.dinb(w_n993_3[1]),.dout(n1118),.clk(gclk));
	jand g0818(.dina(n1118),.dinb(w_n999_2[2]),.dout(n1119),.clk(gclk));
	jand g0819(.dina(n1119),.dinb(w_dff_B_HPK9lmlb8_1),.dout(n1120),.clk(gclk));
	jand g0820(.dina(w_n994_3[1]),.dinb(w_G155_0[1]),.dout(n1121),.clk(gclk));
	jand g0821(.dina(w_n996_3[1]),.dinb(w_G152_0[1]),.dout(n1122),.clk(gclk));
	jor g0822(.dina(w_dff_B_zLZyw14N6_0),.dinb(n1121),.dout(n1123),.clk(gclk));
	jor g0823(.dina(w_dff_B_yzIneDGH8_0),.dinb(n1120),.dout(n1124),.clk(gclk));
	jand g0824(.dina(n1124),.dinb(w_G137_8[0]),.dout(w_dff_A_ss9SJ2Xo4_2),.clk(gclk));
	jor g0825(.dina(w_n1032_0[2]),.dinb(w_G1689_3[1]),.dout(n1126),.clk(gclk));
	jor g0826(.dina(w_n1030_0[2]),.dinb(w_n993_3[0]),.dout(n1127),.clk(gclk));
	jand g0827(.dina(n1127),.dinb(w_n999_2[1]),.dout(n1128),.clk(gclk));
	jand g0828(.dina(n1128),.dinb(n1126),.dout(n1129),.clk(gclk));
	jand g0829(.dina(w_n994_3[0]),.dinb(w_G149_0[1]),.dout(n1130),.clk(gclk));
	jand g0830(.dina(w_n996_3[0]),.dinb(w_G146_0[1]),.dout(n1131),.clk(gclk));
	jor g0831(.dina(w_dff_B_1gDrkq6x2_0),.dinb(n1130),.dout(n1132),.clk(gclk));
	jor g0832(.dina(w_dff_B_ytrX5FtM3_0),.dinb(n1129),.dout(n1133),.clk(gclk));
	jand g0833(.dina(n1133),.dinb(w_G137_7[2]),.dout(w_dff_A_tBBw127J7_2),.clk(gclk));
	jand g0834(.dina(w_n1014_4[0]),.dinb(w_G200_0[0]),.dout(n1135),.clk(gclk));
	jand g0835(.dina(w_n1012_4[0]),.dinb(w_G170_0[0]),.dout(n1136),.clk(gclk));
	jor g0836(.dina(w_n1019_0[1]),.dinb(w_n1008_4[0]),.dout(n1137),.clk(gclk));
	jor g0837(.dina(w_n1021_0[1]),.dinb(w_G1691_4[1]),.dout(n1138),.clk(gclk));
	jand g0838(.dina(n1138),.dinb(n1137),.dout(n1139),.clk(gclk));
	jand g0839(.dina(n1139),.dinb(w_n1007_3[1]),.dout(n1140),.clk(gclk));
	jor g0840(.dina(n1140),.dinb(w_dff_B_Zah5riXS9_1),.dout(n1141),.clk(gclk));
	jor g0841(.dina(n1141),.dinb(w_dff_B_l8beA7pM1_1),.dout(n1142),.clk(gclk));
	jand g0842(.dina(n1142),.dinb(w_G137_7[1]),.dout(w_dff_A_FJ4eLE8y0_2),.clk(gclk));
	jor g0843(.dina(w_n1054_0[1]),.dinb(w_G1691_4[0]),.dout(n1144),.clk(gclk));
	jor g0844(.dina(w_n1052_0[1]),.dinb(w_n1008_3[2]),.dout(n1145),.clk(gclk));
	jand g0845(.dina(n1145),.dinb(w_n1007_3[0]),.dout(n1146),.clk(gclk));
	jand g0846(.dina(w_dff_B_pivs3WiK7_0),.dinb(n1144),.dout(n1147),.clk(gclk));
	jand g0847(.dina(w_n1014_3[2]),.dinb(w_G188_0[0]),.dout(n1148),.clk(gclk));
	jand g0848(.dina(w_n1012_3[2]),.dinb(w_G158_0[0]),.dout(n1149),.clk(gclk));
	jor g0849(.dina(w_dff_B_y1UOWzRD6_0),.dinb(n1148),.dout(n1150),.clk(gclk));
	jor g0850(.dina(w_dff_B_J0McyiMk6_0),.dinb(n1147),.dout(n1151),.clk(gclk));
	jand g0851(.dina(n1151),.dinb(w_G137_7[0]),.dout(w_dff_A_aPMm9gZk7_2),.clk(gclk));
	jor g0852(.dina(w_n1041_0[1]),.dinb(w_G1691_3[2]),.dout(n1153),.clk(gclk));
	jor g0853(.dina(w_n1043_0[1]),.dinb(w_n1008_3[1]),.dout(n1154),.clk(gclk));
	jand g0854(.dina(n1154),.dinb(w_n1007_2[2]),.dout(n1155),.clk(gclk));
	jand g0855(.dina(n1155),.dinb(w_dff_B_7TNR61dt0_1),.dout(n1156),.clk(gclk));
	jand g0856(.dina(w_n1014_3[1]),.dinb(w_G155_0[0]),.dout(n1157),.clk(gclk));
	jand g0857(.dina(w_n1012_3[1]),.dinb(w_G152_0[0]),.dout(n1158),.clk(gclk));
	jor g0858(.dina(w_dff_B_MkJiLRTw9_0),.dinb(n1157),.dout(n1159),.clk(gclk));
	jor g0859(.dina(w_dff_B_uQSx3YNL7_0),.dinb(n1156),.dout(n1160),.clk(gclk));
	jand g0860(.dina(n1160),.dinb(w_G137_6[2]),.dout(w_dff_A_E416vl2P8_2),.clk(gclk));
	jor g0861(.dina(w_n1032_0[1]),.dinb(w_G1691_3[1]),.dout(n1162),.clk(gclk));
	jor g0862(.dina(w_n1030_0[1]),.dinb(w_n1008_3[0]),.dout(n1163),.clk(gclk));
	jand g0863(.dina(n1163),.dinb(w_n1007_2[1]),.dout(n1164),.clk(gclk));
	jand g0864(.dina(n1164),.dinb(n1162),.dout(n1165),.clk(gclk));
	jand g0865(.dina(w_n1014_3[0]),.dinb(w_G149_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n1012_3[0]),.dinb(w_G146_0[0]),.dout(n1167),.clk(gclk));
	jor g0867(.dina(w_dff_B_sFIvMDpm4_0),.dinb(n1166),.dout(n1168),.clk(gclk));
	jor g0868(.dina(w_dff_B_OTqproJZ7_0),.dinb(n1165),.dout(n1169),.clk(gclk));
	jand g0869(.dina(n1169),.dinb(w_G137_6[1]),.dout(w_dff_A_88KRnGpV7_2),.clk(gclk));
	jnot g0870(.din(G135),.dout(n1171),.clk(gclk));
	jnot g0871(.din(G4115),.dout(n1172),.clk(gclk));
	jor g0872(.dina(n1172),.dinb(n1171),.dout(n1173),.clk(gclk));
	jnot g0873(.din(w_n428_1[0]),.dout(n1174),.clk(gclk));
	jor g0874(.dina(n1174),.dinb(w_G3724_0[2]),.dout(n1175),.clk(gclk));
	jnot g0875(.din(w_G3717_0[1]),.dout(n1176),.clk(gclk));
	jnot g0876(.din(w_G3724_0[1]),.dout(n1177),.clk(gclk));
	jxor g0877(.dina(w_n790_0[0]),.dinb(w_dff_B_sGovDXq85_1),.dout(n1178),.clk(gclk));
	jnot g0878(.din(n1178),.dout(n1179),.clk(gclk));
	jor g0879(.dina(w_n1179_0[1]),.dinb(w_n1177_0[1]),.dout(n1180),.clk(gclk));
	jand g0880(.dina(n1180),.dinb(w_dff_B_NEaFt02s3_1),.dout(n1181),.clk(gclk));
	jand g0881(.dina(n1181),.dinb(w_dff_B_GPiIhynG4_1),.dout(n1182),.clk(gclk));
	jor g0882(.dina(w_n795_1[0]),.dinb(w_n1177_0[0]),.dout(n1183),.clk(gclk));
	jor g0883(.dina(w_G3724_0[0]),.dinb(w_G123_0[1]),.dout(n1184),.clk(gclk));
	jand g0884(.dina(n1184),.dinb(w_G3717_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(w_dff_B_VYAmWsj55_0),.dinb(n1183),.dout(n1186),.clk(gclk));
	jor g0886(.dina(n1186),.dinb(w_dff_B_JEENBjMl8_1),.dout(n1187),.clk(gclk));
	jand g0887(.dina(n1187),.dinb(w_dff_B_QSIfbudR1_1),.dout(w_dff_A_oxuB7DjA9_2),.clk(gclk));
	jxor g0888(.dina(w_n1179_0[0]),.dinb(w_n795_0[2]),.dout(w_dff_A_jvwhkrDN8_2),.clk(gclk));
	jand g0889(.dina(w_n750_5[1]),.dinb(w_G123_0[0]),.dout(n1190),.clk(gclk));
	jor g0890(.dina(w_n795_0[1]),.dinb(w_n749_9[2]),.dout(n1191),.clk(gclk));
	jand g0891(.dina(w_n428_0[2]),.dinb(w_n749_9[1]),.dout(n1192),.clk(gclk));
	jor g0892(.dina(n1192),.dinb(w_G4092_6[0]),.dout(n1193),.clk(gclk));
	jnot g0893(.din(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_dff_B_uUfT9kX12_0),.dinb(n1191),.dout(n1195),.clk(gclk));
	jor g0895(.dina(n1195),.dinb(w_dff_B_MwEejZKs4_1),.dout(n1196),.clk(gclk));
	jnot g0896(.din(w_n1196_1[2]),.dout(w_dff_A_UrnIQvBs9_1),.clk(gclk));
	jand g0897(.dina(w_n750_5[0]),.dinb(w_dff_B_QiPIzaLg1_1),.dout(n1198),.clk(gclk));
	jand g0898(.dina(w_n433_0[1]),.dinb(w_n749_9[0]),.dout(n1199),.clk(gclk));
	jnot g0899(.din(n1199),.dout(n1200),.clk(gclk));
	jnot g0900(.din(w_G4092_5[2]),.dout(n1201),.clk(gclk));
	jor g0901(.dina(w_n969_0[0]),.dinb(w_n749_8[2]),.dout(n1202),.clk(gclk));
	jand g0902(.dina(n1202),.dinb(w_n1201_0[2]),.dout(n1203),.clk(gclk));
	jand g0903(.dina(n1203),.dinb(w_dff_B_dOvBVwnH4_1),.dout(n1204),.clk(gclk));
	jor g0904(.dina(n1204),.dinb(w_dff_B_UUBNS6RN1_1),.dout(n1205),.clk(gclk));
	jnot g0905(.din(w_n1205_1[2]),.dout(w_dff_A_Fi5KrCYh7_1),.clk(gclk));
	jand g0906(.dina(w_n750_4[2]),.dinb(w_dff_B_HLhD5N0M9_1),.dout(n1207),.clk(gclk));
	jor g0907(.dina(w_n986_0[0]),.dinb(w_n749_8[1]),.dout(n1208),.clk(gclk));
	jand g0908(.dina(w_n423_0[1]),.dinb(w_n749_8[0]),.dout(n1209),.clk(gclk));
	jor g0909(.dina(n1209),.dinb(w_G4092_5[1]),.dout(n1210),.clk(gclk));
	jnot g0910(.din(n1210),.dout(n1211),.clk(gclk));
	jand g0911(.dina(w_dff_B_K5sujEbX8_0),.dinb(n1208),.dout(n1212),.clk(gclk));
	jor g0912(.dina(n1212),.dinb(w_dff_B_0ls9iHpe0_1),.dout(n1213),.clk(gclk));
	jnot g0913(.din(w_n1213_1[2]),.dout(w_dff_A_5bYRvP0i0_1),.clk(gclk));
	jand g0914(.dina(w_n750_4[1]),.dinb(w_dff_B_ppcvgk152_1),.dout(n1215),.clk(gclk));
	jnot g0915(.din(n1215),.dout(n1216),.clk(gclk));
	jand g0916(.dina(w_n989_0[0]),.dinb(w_G4091_2[2]),.dout(n1217),.clk(gclk));
	jand g0917(.dina(w_n412_0[1]),.dinb(w_n749_7[2]),.dout(n1218),.clk(gclk));
	jor g0918(.dina(n1218),.dinb(w_G4092_5[0]),.dout(n1219),.clk(gclk));
	jor g0919(.dina(w_dff_B_GbydITx23_0),.dinb(n1217),.dout(n1220),.clk(gclk));
	jand g0920(.dina(n1220),.dinb(w_dff_B_FP9SyRB59_1),.dout(G830_fa_),.clk(gclk));
	jand g0921(.dina(w_n680_0[0]),.dinb(w_G245_0[0]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(w_dff_B_MvMuVnvU9_0),.dinb(w_n935_0[0]),.dout(n1223),.clk(gclk));
	jnot g0923(.din(w_G998_0),.dout(n1224),.clk(gclk));
	jand g0924(.dina(w_n318_0[0]),.dinb(w_G601_0),.dout(n1225),.clk(gclk));
	jand g0925(.dina(n1225),.dinb(w_G559_0[0]),.dout(n1226),.clk(gclk));
	jand g0926(.dina(w_dff_B_Mbqsu6jf8_0),.dinb(w_n670_0[0]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_dff_B_7QKpzjzx6_0),.dinb(n1224),.dout(n1228),.clk(gclk));
	jand g0928(.dina(n1228),.dinb(w_dff_B_MvEi3CGB6_1),.dout(w_dff_A_vafD6ff48_2),.clk(gclk));
	jand g0929(.dina(w_n750_4[0]),.dinb(w_dff_B_x0JyqcE81_1),.dout(n1230),.clk(gclk));
	jand g0930(.dina(w_n551_0[1]),.dinb(w_n749_7[1]),.dout(n1231),.clk(gclk));
	jnot g0931(.din(n1231),.dout(n1232),.clk(gclk));
	jor g0932(.dina(w_n944_0[0]),.dinb(w_n749_7[0]),.dout(n1233),.clk(gclk));
	jand g0933(.dina(n1233),.dinb(w_n1201_0[1]),.dout(n1234),.clk(gclk));
	jand g0934(.dina(n1234),.dinb(w_dff_B_zNX5cKln3_1),.dout(n1235),.clk(gclk));
	jor g0935(.dina(n1235),.dinb(w_dff_B_bNSu0CbU2_1),.dout(n1236),.clk(gclk));
	jnot g0936(.din(w_n1236_1[2]),.dout(w_dff_A_MInp1sVP2_1),.clk(gclk));
	jand g0937(.dina(w_n750_3[2]),.dinb(w_dff_B_ceVZ87HC7_1),.dout(n1238),.clk(gclk));
	jnot g0938(.din(n1238),.dout(n1239),.clk(gclk));
	jand g0939(.dina(w_n949_0[0]),.dinb(w_G4091_2[1]),.dout(n1240),.clk(gclk));
	jand g0940(.dina(w_n459_0[0]),.dinb(w_n749_6[2]),.dout(n1241),.clk(gclk));
	jor g0941(.dina(n1241),.dinb(w_G4092_4[2]),.dout(n1242),.clk(gclk));
	jor g0942(.dina(w_dff_B_bhsRT5yD6_0),.dinb(n1240),.dout(n1243),.clk(gclk));
	jand g0943(.dina(n1243),.dinb(w_dff_B_ko9Gnr9s4_1),.dout(G865_fa_),.clk(gclk));
	jand g0944(.dina(w_n750_3[1]),.dinb(w_dff_B_wPc01Xff2_1),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n517_0[0]),.dinb(w_n749_6[1]),.dout(n1246),.clk(gclk));
	jnot g0946(.din(n1246),.dout(n1247),.clk(gclk));
	jor g0947(.dina(w_n957_0[0]),.dinb(w_n749_6[0]),.dout(n1248),.clk(gclk));
	jand g0948(.dina(n1248),.dinb(w_n1201_0[0]),.dout(n1249),.clk(gclk));
	jand g0949(.dina(n1249),.dinb(w_dff_B_xh3eOoMT7_1),.dout(n1250),.clk(gclk));
	jor g0950(.dina(n1250),.dinb(w_dff_B_uuDGuNni8_1),.dout(n1251),.clk(gclk));
	jnot g0951(.din(w_n1251_1[2]),.dout(w_dff_A_CZVTd2RE5_1),.clk(gclk));
	jand g0952(.dina(w_n750_3[0]),.dinb(w_dff_B_ZdKFumnR9_1),.dout(n1253),.clk(gclk));
	jnot g0953(.din(n1253),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n964_0[0]),.dinb(w_G4091_2[0]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n504_0[0]),.dinb(w_n749_5[2]),.dout(n1256),.clk(gclk));
	jor g0956(.dina(n1256),.dinb(w_G4092_4[1]),.dout(n1257),.clk(gclk));
	jor g0957(.dina(w_dff_B_LvgzSzjn0_0),.dinb(n1255),.dout(n1258),.clk(gclk));
	jand g0958(.dina(n1258),.dinb(w_dff_B_z39GyPid4_1),.dout(G869_fa_),.clk(gclk));
	jor g0959(.dina(w_G4089_6[0]),.dinb(w_G109_0[1]),.dout(n1260),.clk(gclk));
	jor g0960(.dina(w_n852_6[0]),.dinb(w_G106_0[1]),.dout(n1261),.clk(gclk));
	jand g0961(.dina(n1261),.dinb(w_G4090_2[2]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(n1262),.dinb(w_dff_B_E2Jbsujk9_1),.dout(n1263),.clk(gclk));
	jor g0963(.dina(w_n1236_1[1]),.dinb(w_n852_5[2]),.dout(n1264),.clk(gclk));
	jor g0964(.dina(w_n1196_1[1]),.dinb(w_G4089_5[2]),.dout(n1265),.clk(gclk));
	jand g0965(.dina(n1265),.dinb(w_n854_2[2]),.dout(n1266),.clk(gclk));
	jand g0966(.dina(n1266),.dinb(n1264),.dout(n1267),.clk(gclk));
	jor g0967(.dina(n1267),.dinb(w_dff_B_t8Pisbq56_1),.dout(w_dff_A_2XGOUCxJ2_2),.clk(gclk));
	jor g0968(.dina(w_n1196_1[0]),.dinb(w_G4088_6[0]),.dout(n1269),.clk(gclk));
	jor g0969(.dina(w_n1236_1[0]),.dinb(w_n797_6[0]),.dout(n1270),.clk(gclk));
	jand g0970(.dina(n1270),.dinb(w_n800_2[2]),.dout(n1271),.clk(gclk));
	jand g0971(.dina(n1271),.dinb(w_dff_B_FAOPZv5V7_1),.dout(n1272),.clk(gclk));
	jor g0972(.dina(w_n797_5[2]),.dinb(w_G106_0[0]),.dout(n1273),.clk(gclk));
	jor g0973(.dina(w_G4088_5[2]),.dinb(w_G109_0[0]),.dout(n1274),.clk(gclk));
	jand g0974(.dina(n1274),.dinb(w_G4087_2[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(n1275),.dinb(n1273),.dout(n1276),.clk(gclk));
	jor g0976(.dina(w_dff_B_nKOjYhof4_0),.dinb(n1272),.dout(w_dff_A_fDdSOlMD0_2),.clk(gclk));
	jor g0977(.dina(w_n1205_1[1]),.dinb(w_G4088_5[1]),.dout(n1278),.clk(gclk));
	jnot g0978(.din(w_G865_0),.dout(n1279),.clk(gclk));
	jor g0979(.dina(w_n1279_1[1]),.dinb(w_n797_5[1]),.dout(n1280),.clk(gclk));
	jand g0980(.dina(n1280),.dinb(w_n800_2[1]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(n1281),.dinb(w_dff_B_BqxIVWIf3_1),.dout(n1282),.clk(gclk));
	jor g0982(.dina(w_n797_5[0]),.dinb(w_G49_0[1]),.dout(n1283),.clk(gclk));
	jor g0983(.dina(w_G4088_5[0]),.dinb(w_G46_0[1]),.dout(n1284),.clk(gclk));
	jand g0984(.dina(n1284),.dinb(w_G4087_2[1]),.dout(n1285),.clk(gclk));
	jand g0985(.dina(n1285),.dinb(n1283),.dout(n1286),.clk(gclk));
	jor g0986(.dina(w_dff_B_ZrjqD6Vp2_0),.dinb(n1282),.dout(w_dff_A_5eIRg5hX3_2),.clk(gclk));
	jor g0987(.dina(w_n1213_1[1]),.dinb(w_G4088_4[2]),.dout(n1288),.clk(gclk));
	jor g0988(.dina(w_n1251_1[1]),.dinb(w_n797_4[2]),.dout(n1289),.clk(gclk));
	jand g0989(.dina(n1289),.dinb(w_n800_2[0]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(n1290),.dinb(w_dff_B_XV8wNjjV6_1),.dout(n1291),.clk(gclk));
	jor g0991(.dina(w_n797_4[1]),.dinb(w_G103_0[1]),.dout(n1292),.clk(gclk));
	jor g0992(.dina(w_G4088_4[1]),.dinb(w_G100_0[1]),.dout(n1293),.clk(gclk));
	jand g0993(.dina(n1293),.dinb(w_G4087_2[0]),.dout(n1294),.clk(gclk));
	jand g0994(.dina(n1294),.dinb(n1292),.dout(n1295),.clk(gclk));
	jor g0995(.dina(w_dff_B_cWwYlpGe4_0),.dinb(n1291),.dout(w_dff_A_sYyisCNw9_2),.clk(gclk));
	jnot g0996(.din(w_G830_0),.dout(n1297),.clk(gclk));
	jor g0997(.dina(w_n1297_1[1]),.dinb(w_G4088_4[0]),.dout(n1298),.clk(gclk));
	jnot g0998(.din(w_G869_0),.dout(n1299),.clk(gclk));
	jor g0999(.dina(w_n1299_1[1]),.dinb(w_n797_4[0]),.dout(n1300),.clk(gclk));
	jand g1000(.dina(n1300),.dinb(w_n800_1[2]),.dout(n1301),.clk(gclk));
	jand g1001(.dina(n1301),.dinb(w_dff_B_83ZWJmPx7_1),.dout(n1302),.clk(gclk));
	jor g1002(.dina(w_n797_3[2]),.dinb(w_G40_0[1]),.dout(n1303),.clk(gclk));
	jor g1003(.dina(w_G4088_3[2]),.dinb(w_G91_0[1]),.dout(n1304),.clk(gclk));
	jand g1004(.dina(n1304),.dinb(w_G4087_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(n1305),.dinb(n1303),.dout(n1306),.clk(gclk));
	jor g1006(.dina(w_dff_B_wUvw5KZf0_0),.dinb(n1302),.dout(w_dff_A_jLaVIWAZ5_2),.clk(gclk));
	jor g1007(.dina(w_n1205_1[0]),.dinb(w_G4089_5[1]),.dout(n1308),.clk(gclk));
	jor g1008(.dina(w_n1279_1[0]),.dinb(w_n852_5[1]),.dout(n1309),.clk(gclk));
	jand g1009(.dina(n1309),.dinb(w_n854_2[1]),.dout(n1310),.clk(gclk));
	jand g1010(.dina(n1310),.dinb(w_dff_B_GERUinjS1_1),.dout(n1311),.clk(gclk));
	jor g1011(.dina(w_n852_5[0]),.dinb(w_G49_0[0]),.dout(n1312),.clk(gclk));
	jor g1012(.dina(w_G4089_5[0]),.dinb(w_G46_0[0]),.dout(n1313),.clk(gclk));
	jand g1013(.dina(n1313),.dinb(w_G4090_2[1]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(n1314),.dinb(n1312),.dout(n1315),.clk(gclk));
	jor g1015(.dina(w_dff_B_bsKDHyqd4_0),.dinb(n1311),.dout(w_dff_A_jHQxUsEJ2_2),.clk(gclk));
	jor g1016(.dina(w_n1213_1[0]),.dinb(w_G4089_4[2]),.dout(n1317),.clk(gclk));
	jor g1017(.dina(w_n1251_1[0]),.dinb(w_n852_4[2]),.dout(n1318),.clk(gclk));
	jand g1018(.dina(n1318),.dinb(w_n854_2[0]),.dout(n1319),.clk(gclk));
	jand g1019(.dina(n1319),.dinb(w_dff_B_P8Q07vcW5_1),.dout(n1320),.clk(gclk));
	jor g1020(.dina(w_n852_4[1]),.dinb(w_G103_0[0]),.dout(n1321),.clk(gclk));
	jor g1021(.dina(w_G4089_4[1]),.dinb(w_G100_0[0]),.dout(n1322),.clk(gclk));
	jand g1022(.dina(n1322),.dinb(w_G4090_2[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(n1323),.dinb(n1321),.dout(n1324),.clk(gclk));
	jor g1024(.dina(w_dff_B_YZF84n0Q0_0),.dinb(n1320),.dout(w_dff_A_nrcvRrKO0_2),.clk(gclk));
	jor g1025(.dina(w_n1297_1[0]),.dinb(w_G4089_4[0]),.dout(n1326),.clk(gclk));
	jor g1026(.dina(w_n1299_1[0]),.dinb(w_n852_4[0]),.dout(n1327),.clk(gclk));
	jand g1027(.dina(n1327),.dinb(w_n854_1[2]),.dout(n1328),.clk(gclk));
	jand g1028(.dina(n1328),.dinb(w_dff_B_gCFCo7wU8_1),.dout(n1329),.clk(gclk));
	jor g1029(.dina(w_n852_3[2]),.dinb(w_G40_0[0]),.dout(n1330),.clk(gclk));
	jor g1030(.dina(w_G4089_3[2]),.dinb(w_G91_0[0]),.dout(n1331),.clk(gclk));
	jand g1031(.dina(n1331),.dinb(w_G4090_1[2]),.dout(n1332),.clk(gclk));
	jand g1032(.dina(n1332),.dinb(n1330),.dout(n1333),.clk(gclk));
	jor g1033(.dina(w_dff_B_wucxeoWg8_0),.dinb(n1329),.dout(w_dff_A_7DtcfDVl6_2),.clk(gclk));
	jor g1034(.dina(w_n1297_0[2]),.dinb(w_G1689_3[0]),.dout(n1335),.clk(gclk));
	jor g1035(.dina(w_n1299_0[2]),.dinb(w_n993_2[2]),.dout(n1336),.clk(gclk));
	jand g1036(.dina(n1336),.dinb(w_n999_2[0]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(n1337),.dinb(w_dff_B_ABsc0nYs4_1),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n994_2[2]),.dinb(w_G203_0[1]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n996_2[2]),.dinb(w_G173_0[1]),.dout(n1340),.clk(gclk));
	jor g1040(.dina(w_dff_B_ubgztRBW1_0),.dinb(n1339),.dout(n1341),.clk(gclk));
	jor g1041(.dina(w_dff_B_nFMKQL577_0),.dinb(n1338),.dout(n1342),.clk(gclk));
	jand g1042(.dina(n1342),.dinb(w_G137_6[0]),.dout(w_dff_A_P32bXcZR1_2),.clk(gclk));
	jor g1043(.dina(w_n1251_0[2]),.dinb(w_n993_2[1]),.dout(n1344),.clk(gclk));
	jor g1044(.dina(w_n1213_0[2]),.dinb(w_G1689_2[2]),.dout(n1345),.clk(gclk));
	jand g1045(.dina(n1345),.dinb(w_n999_1[2]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(n1346),.dinb(w_dff_B_dPM72rwn1_1),.dout(n1347),.clk(gclk));
	jand g1047(.dina(w_n994_2[1]),.dinb(w_G197_0[1]),.dout(n1348),.clk(gclk));
	jand g1048(.dina(w_n996_2[1]),.dinb(w_G167_0[1]),.dout(n1349),.clk(gclk));
	jor g1049(.dina(w_dff_B_GW0o3jnx6_0),.dinb(n1348),.dout(n1350),.clk(gclk));
	jor g1050(.dina(w_dff_B_qz6367Se3_0),.dinb(n1347),.dout(n1351),.clk(gclk));
	jand g1051(.dina(n1351),.dinb(w_G137_5[2]),.dout(w_dff_A_7lXH9BOj8_2),.clk(gclk));
	jand g1052(.dina(w_n994_2[0]),.dinb(w_G194_0[1]),.dout(n1353),.clk(gclk));
	jand g1053(.dina(w_n996_2[0]),.dinb(w_G164_0[1]),.dout(n1354),.clk(gclk));
	jor g1054(.dina(w_dff_B_n0fNFoP04_0),.dinb(n1353),.dout(n1355),.clk(gclk));
	jor g1055(.dina(w_n1205_0[2]),.dinb(w_G1689_2[1]),.dout(n1356),.clk(gclk));
	jor g1056(.dina(w_n1279_0[2]),.dinb(w_n993_2[0]),.dout(n1357),.clk(gclk));
	jand g1057(.dina(n1357),.dinb(w_dff_B_aM7Hh88Z6_1),.dout(n1358),.clk(gclk));
	jand g1058(.dina(n1358),.dinb(w_n999_1[1]),.dout(n1359),.clk(gclk));
	jor g1059(.dina(n1359),.dinb(w_dff_B_2N7sWeEP9_1),.dout(n1360),.clk(gclk));
	jand g1060(.dina(n1360),.dinb(w_G137_5[1]),.dout(w_dff_A_6ondWxNN6_2),.clk(gclk));
	jand g1061(.dina(w_n994_1[2]),.dinb(w_G191_0[1]),.dout(n1362),.clk(gclk));
	jand g1062(.dina(w_n996_1[2]),.dinb(w_G161_0[1]),.dout(n1363),.clk(gclk));
	jor g1063(.dina(w_dff_B_WuxwULkX2_0),.dinb(n1362),.dout(n1364),.clk(gclk));
	jor g1064(.dina(w_n1196_0[2]),.dinb(w_G1689_2[0]),.dout(n1365),.clk(gclk));
	jor g1065(.dina(w_n1236_0[2]),.dinb(w_n993_1[2]),.dout(n1366),.clk(gclk));
	jand g1066(.dina(n1366),.dinb(w_dff_B_ud4zDNMc5_1),.dout(n1367),.clk(gclk));
	jand g1067(.dina(n1367),.dinb(w_n999_1[0]),.dout(n1368),.clk(gclk));
	jor g1068(.dina(n1368),.dinb(w_dff_B_9O0W9hO07_1),.dout(n1369),.clk(gclk));
	jand g1069(.dina(n1369),.dinb(w_G137_5[0]),.dout(w_dff_A_EW50mF6G8_2),.clk(gclk));
	jor g1070(.dina(w_n1297_0[1]),.dinb(w_G1691_3[0]),.dout(n1371),.clk(gclk));
	jor g1071(.dina(w_n1299_0[1]),.dinb(w_n1008_2[2]),.dout(n1372),.clk(gclk));
	jand g1072(.dina(n1372),.dinb(w_n1007_2[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(n1373),.dinb(w_dff_B_kLo2r7RI9_1),.dout(n1374),.clk(gclk));
	jand g1074(.dina(w_n1014_2[2]),.dinb(w_G203_0[0]),.dout(n1375),.clk(gclk));
	jand g1075(.dina(w_n1012_2[2]),.dinb(w_G173_0[0]),.dout(n1376),.clk(gclk));
	jor g1076(.dina(w_dff_B_LMyJSMy41_0),.dinb(n1375),.dout(n1377),.clk(gclk));
	jor g1077(.dina(w_dff_B_IFjCnL9p5_0),.dinb(n1374),.dout(n1378),.clk(gclk));
	jand g1078(.dina(n1378),.dinb(w_G137_4[2]),.dout(w_dff_A_qtIVFaz20_2),.clk(gclk));
	jand g1079(.dina(w_n1014_2[1]),.dinb(w_G197_0[0]),.dout(n1380),.clk(gclk));
	jand g1080(.dina(w_n1012_2[1]),.dinb(w_G167_0[0]),.dout(n1381),.clk(gclk));
	jor g1081(.dina(w_dff_B_ijBLdRBO8_0),.dinb(n1380),.dout(n1382),.clk(gclk));
	jor g1082(.dina(w_n1213_0[1]),.dinb(w_G1691_2[2]),.dout(n1383),.clk(gclk));
	jor g1083(.dina(w_n1251_0[1]),.dinb(w_n1008_2[1]),.dout(n1384),.clk(gclk));
	jand g1084(.dina(n1384),.dinb(n1383),.dout(n1385),.clk(gclk));
	jand g1085(.dina(n1385),.dinb(w_n1007_1[2]),.dout(n1386),.clk(gclk));
	jor g1086(.dina(n1386),.dinb(w_dff_B_dEHTAsTF1_1),.dout(n1387),.clk(gclk));
	jand g1087(.dina(n1387),.dinb(w_G137_4[1]),.dout(w_dff_A_SZppPzwU8_2),.clk(gclk));
	jor g1088(.dina(w_n1205_0[1]),.dinb(w_G1691_2[1]),.dout(n1389),.clk(gclk));
	jor g1089(.dina(w_n1279_0[1]),.dinb(w_n1008_2[0]),.dout(n1390),.clk(gclk));
	jand g1090(.dina(n1390),.dinb(w_n1007_1[1]),.dout(n1391),.clk(gclk));
	jand g1091(.dina(n1391),.dinb(w_dff_B_yu53a9v41_1),.dout(n1392),.clk(gclk));
	jand g1092(.dina(w_n1014_2[0]),.dinb(w_G194_0[0]),.dout(n1393),.clk(gclk));
	jand g1093(.dina(w_n1012_2[0]),.dinb(w_G164_0[0]),.dout(n1394),.clk(gclk));
	jor g1094(.dina(w_dff_B_exdElFVE8_0),.dinb(n1393),.dout(n1395),.clk(gclk));
	jor g1095(.dina(w_dff_B_JnaAnNOS8_0),.dinb(n1392),.dout(n1396),.clk(gclk));
	jand g1096(.dina(n1396),.dinb(w_G137_4[0]),.dout(w_dff_A_EjeCPIAX3_2),.clk(gclk));
	jor g1097(.dina(w_n1236_0[1]),.dinb(w_n1008_1[2]),.dout(n1398),.clk(gclk));
	jor g1098(.dina(w_n1196_0[1]),.dinb(w_G1691_2[0]),.dout(n1399),.clk(gclk));
	jand g1099(.dina(n1399),.dinb(w_n1007_1[0]),.dout(n1400),.clk(gclk));
	jand g1100(.dina(n1400),.dinb(n1398),.dout(n1401),.clk(gclk));
	jand g1101(.dina(w_n1014_1[2]),.dinb(w_G191_0[0]),.dout(n1402),.clk(gclk));
	jand g1102(.dina(w_n1012_1[2]),.dinb(w_G161_0[0]),.dout(n1403),.clk(gclk));
	jor g1103(.dina(w_dff_B_RcXC3ijD4_0),.dinb(n1402),.dout(n1404),.clk(gclk));
	jor g1104(.dina(w_dff_B_riE1MaDo8_0),.dinb(n1401),.dout(n1405),.clk(gclk));
	jand g1105(.dina(n1405),.dinb(w_G137_3[2]),.dout(w_dff_A_NyJ1LQKr6_2),.clk(gclk));
	jand g1106(.dina(w_n746_0[0]),.dinb(w_n648_0[2]),.dout(n1407),.clk(gclk));
	jxor g1107(.dina(w_n977_0[0]),.dinb(w_n654_1[0]),.dout(n1408),.clk(gclk));
	jxor g1108(.dina(n1408),.dinb(w_n644_0[0]),.dout(n1409),.clk(gclk));
	jxor g1109(.dina(w_dff_B_unjhe5ER1_0),.dinb(n1407),.dout(n1410),.clk(gclk));
	jor g1110(.dina(w_n1410_0[2]),.dinb(w_n737_0[2]),.dout(n1411),.clk(gclk));
	jnot g1111(.din(w_G2174_0[2]),.dout(n1412),.clk(gclk));
	jnot g1112(.din(w_n719_0[0]),.dout(n1413),.clk(gclk));
	jnot g1113(.din(w_n720_0[0]),.dout(n1414),.clk(gclk));
	jor g1114(.dina(w_n821_0[0]),.dinb(w_dff_B_R8tE4bJQ6_1),.dout(n1415),.clk(gclk));
	jand g1115(.dina(n1415),.dinb(w_dff_B_6fn1E8pr1_1),.dout(n1416),.clk(gclk));
	jxor g1116(.dina(w_n742_0[0]),.dinb(w_n654_0[2]),.dout(n1417),.clk(gclk));
	jxor g1117(.dina(n1417),.dinb(w_n792_0[0]),.dout(n1418),.clk(gclk));
	jnot g1118(.din(w_n660_0[1]),.dout(n1419),.clk(gclk));
	jand g1119(.dina(w_n745_0[0]),.dinb(w_n648_0[1]),.dout(n1420),.clk(gclk));
	jand g1120(.dina(n1420),.dinb(w_dff_B_LvAdtN1b5_1),.dout(n1421),.clk(gclk));
	jxor g1121(.dina(n1421),.dinb(w_dff_B_74lelJ1H2_1),.dout(n1422),.clk(gclk));
	jor g1122(.dina(w_n1422_0[1]),.dinb(w_n1416_0[1]),.dout(n1423),.clk(gclk));
	jand g1123(.dina(n1423),.dinb(w_n1412_0[2]),.dout(n1424),.clk(gclk));
	jand g1124(.dina(n1424),.dinb(w_dff_B_V7dT85qn1_1),.dout(n1425),.clk(gclk));
	jnot g1125(.din(w_n1425_0[1]),.dout(n1426),.clk(gclk));
	jnot g1126(.din(w_n641_1[0]),.dout(n1427),.clk(gclk));
	jand g1127(.dina(w_n1416_0[0]),.dinb(w_dff_B_sbTVpKbU0_1),.dout(n1428),.clk(gclk));
	jor g1128(.dina(w_n1428_0[1]),.dinb(w_n1422_0[0]),.dout(n1429),.clk(gclk));
	jnot g1129(.din(w_n1429_0[1]),.dout(n1430),.clk(gclk));
	jnot g1130(.din(w_n1410_0[1]),.dout(n1431),.clk(gclk));
	jand g1131(.dina(w_n1428_0[0]),.dinb(n1431),.dout(n1432),.clk(gclk));
	jor g1132(.dina(n1432),.dinb(w_n1412_0[1]),.dout(n1433),.clk(gclk));
	jor g1133(.dina(n1433),.dinb(n1430),.dout(n1434),.clk(gclk));
	jand g1134(.dina(n1434),.dinb(n1426),.dout(n1435),.clk(gclk));
	jor g1135(.dina(w_n728_0[0]),.dinb(w_n637_0[0]),.dout(n1436),.clk(gclk));
	jxor g1136(.dina(w_dff_B_rwnme35b7_0),.dinb(w_n733_0[1]),.dout(n1437),.clk(gclk));
	jxor g1137(.dina(w_dff_B_4gd9p14e0_0),.dinb(w_n735_0[1]),.dout(n1438),.clk(gclk));
	jor g1138(.dina(n1438),.dinb(w_G2174_0[1]),.dout(n1439),.clk(gclk));
	jor g1139(.dina(w_n735_0[0]),.dinb(w_n640_0[0]),.dout(n1440),.clk(gclk));
	jor g1140(.dina(w_n819_0[0]),.dinb(w_n628_0[0]),.dout(n1441),.clk(gclk));
	jor g1141(.dina(w_n733_0[0]),.dinb(w_n814_0[0]),.dout(n1442),.clk(gclk));
	jor g1142(.dina(n1442),.dinb(w_n639_0[0]),.dout(n1443),.clk(gclk));
	jand g1143(.dina(n1443),.dinb(w_dff_B_jTV28bEn7_1),.dout(n1444),.clk(gclk));
	jxor g1144(.dina(n1444),.dinb(n1440),.dout(n1445),.clk(gclk));
	jor g1145(.dina(n1445),.dinb(w_n1412_0[0]),.dout(n1446),.clk(gclk));
	jand g1146(.dina(n1446),.dinb(w_dff_B_hdAH0NYh6_1),.dout(n1447),.clk(gclk));
	jxor g1147(.dina(w_n620_0[1]),.dinb(w_n618_0[0]),.dout(n1448),.clk(gclk));
	jxor g1148(.dina(w_n767_0[0]),.dinb(w_n624_0[0]),.dout(n1449),.clk(gclk));
	jxor g1149(.dina(n1449),.dinb(w_dff_B_M3EazxG68_1),.dout(n1450),.clk(gclk));
	jxor g1150(.dina(w_dff_B_fxt2xFq75_0),.dinb(n1447),.dout(n1451),.clk(gclk));
	jnot g1151(.din(w_n1451_0[1]),.dout(n1452),.clk(gclk));
	jand g1152(.dina(w_dff_B_070zhp4a5_0),.dinb(n1435),.dout(n1453),.clk(gclk));
	jor g1153(.dina(w_n737_0[1]),.dinb(w_n641_0[2]),.dout(n1454),.clk(gclk));
	jor g1154(.dina(n1454),.dinb(w_n1410_0[0]),.dout(n1455),.clk(gclk));
	jand g1155(.dina(n1455),.dinb(w_G2174_0[0]),.dout(n1456),.clk(gclk));
	jand g1156(.dina(n1456),.dinb(w_n1429_0[0]),.dout(n1457),.clk(gclk));
	jor g1157(.dina(n1457),.dinb(w_n1425_0[0]),.dout(n1458),.clk(gclk));
	jand g1158(.dina(w_n1451_0[0]),.dinb(n1458),.dout(n1459),.clk(gclk));
	jor g1159(.dina(n1459),.dinb(w_n749_5[1]),.dout(n1460),.clk(gclk));
	jor g1160(.dina(n1460),.dinb(w_dff_B_Z90rQbll4_1),.dout(n1461),.clk(gclk));
	jand g1161(.dina(w_G351_1[0]),.dinb(w_G248_4[1]),.dout(n1462),.clk(gclk));
	jand g1162(.dina(w_n374_0[2]),.dinb(w_G251_4[0]),.dout(n1463),.clk(gclk));
	jor g1163(.dina(n1463),.dinb(w_n377_0[1]),.dout(n1464),.clk(gclk));
	jor g1164(.dina(n1464),.dinb(w_dff_B_qaJGMqE42_1),.dout(n1465),.clk(gclk));
	jand g1165(.dina(w_n374_0[1]),.dinb(w_n406_4[0]),.dout(n1466),.clk(gclk));
	jand g1166(.dina(w_G351_0[2]),.dinb(w_n408_4[1]),.dout(n1467),.clk(gclk));
	jor g1167(.dina(n1467),.dinb(n1466),.dout(n1468),.clk(gclk));
	jor g1168(.dina(n1468),.dinb(w_G534_0[2]),.dout(n1469),.clk(gclk));
	jand g1169(.dina(n1469),.dinb(n1465),.dout(n1470),.clk(gclk));
	jand g1170(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1471),.clk(gclk));
	jand g1171(.dina(w_n387_0[2]),.dinb(w_G251_3[2]),.dout(n1472),.clk(gclk));
	jor g1172(.dina(n1472),.dinb(w_n389_0[1]),.dout(n1473),.clk(gclk));
	jor g1173(.dina(n1473),.dinb(w_dff_B_SbN4iOHA4_1),.dout(n1474),.clk(gclk));
	jand g1174(.dina(w_n387_0[1]),.dinb(w_n406_3[2]),.dout(n1475),.clk(gclk));
	jand g1175(.dina(w_G341_0[2]),.dinb(w_n408_4[0]),.dout(n1476),.clk(gclk));
	jor g1176(.dina(n1476),.dinb(n1475),.dout(n1477),.clk(gclk));
	jor g1177(.dina(n1477),.dinb(w_G523_0[1]),.dout(n1478),.clk(gclk));
	jand g1178(.dina(n1478),.dinb(n1474),.dout(n1479),.clk(gclk));
	jxor g1179(.dina(n1479),.dinb(n1470),.dout(n1480),.clk(gclk));
	jor g1180(.dina(w_n435_1[0]),.dinb(w_n369_1[0]),.dout(n1481),.clk(gclk));
	jor g1181(.dina(w_G324_0[2]),.dinb(w_n366_1[0]),.dout(n1482),.clk(gclk));
	jand g1182(.dina(n1482),.dinb(w_G503_0[2]),.dout(n1483),.clk(gclk));
	jand g1183(.dina(n1483),.dinb(w_dff_B_1sRfBGLA1_1),.dout(n1484),.clk(gclk));
	jor g1184(.dina(w_G324_0[1]),.dinb(w_G254_1[0]),.dout(n1485),.clk(gclk));
	jor g1185(.dina(w_n435_0[2]),.dinb(w_G242_1[0]),.dout(n1486),.clk(gclk));
	jand g1186(.dina(n1486),.dinb(w_dff_B_0IfXNE3G0_1),.dout(n1487),.clk(gclk));
	jand g1187(.dina(n1487),.dinb(w_n437_0[0]),.dout(n1488),.clk(gclk));
	jor g1188(.dina(n1488),.dinb(n1484),.dout(n1489),.clk(gclk));
	jor g1189(.dina(w_G514_0[2]),.dinb(w_n408_3[2]),.dout(n1490),.clk(gclk));
	jor g1190(.dina(w_n361_0[0]),.dinb(w_G248_3[2]),.dout(n1491),.clk(gclk));
	jand g1191(.dina(n1491),.dinb(n1490),.dout(n1492),.clk(gclk));
	jxor g1192(.dina(n1492),.dinb(w_n371_0[0]),.dout(n1493),.clk(gclk));
	jxor g1193(.dina(w_dff_B_YFQvHGfJ1_0),.dinb(n1489),.dout(n1494),.clk(gclk));
	jxor g1194(.dina(n1494),.dinb(n1480),.dout(n1495),.clk(gclk));
	jxor g1195(.dina(w_n433_0[0]),.dinb(w_n428_0[1]),.dout(n1496),.clk(gclk));
	jxor g1196(.dina(w_n423_0[0]),.dinb(w_n412_0[0]),.dout(n1497),.clk(gclk));
	jxor g1197(.dina(n1497),.dinb(w_dff_B_qR3rCMT00_1),.dout(n1498),.clk(gclk));
	jxor g1198(.dina(n1498),.dinb(n1495),.dout(n1499),.clk(gclk));
	jand g1199(.dina(n1499),.dinb(w_n749_5[0]),.dout(n1500),.clk(gclk));
	jnot g1200(.din(n1500),.dout(n1501),.clk(gclk));
	jand g1201(.dina(w_dff_B_uBoKKbTs1_0),.dinb(n1461),.dout(n1502),.clk(gclk));
	jor g1202(.dina(n1502),.dinb(w_G4092_4[0]),.dout(n1503),.clk(gclk));
	jnot g1203(.din(w_n750_2[2]),.dout(n1504),.clk(gclk));
	jor g1204(.dina(w_n1504_0[1]),.dinb(w_dff_B_dichDG2I4_1),.dout(n1505),.clk(gclk));
	jand g1205(.dina(w_dff_B_2nAI3GlU6_0),.dinb(w_n1503_0[1]),.dout(w_dff_A_VYoWKH9V5_2),.clk(gclk));
	jand g1206(.dina(w_G273_1[0]),.dinb(w_G248_3[1]),.dout(n1507),.clk(gclk));
	jand g1207(.dina(w_n471_0[2]),.dinb(w_G251_3[1]),.dout(n1508),.clk(gclk));
	jor g1208(.dina(n1508),.dinb(w_n473_1[0]),.dout(n1509),.clk(gclk));
	jor g1209(.dina(n1509),.dinb(w_dff_B_Iy7RRtdp3_1),.dout(n1510),.clk(gclk));
	jand g1210(.dina(w_n471_0[1]),.dinb(w_n406_3[1]),.dout(n1511),.clk(gclk));
	jand g1211(.dina(w_G273_0[2]),.dinb(w_n408_3[1]),.dout(n1512),.clk(gclk));
	jor g1212(.dina(n1512),.dinb(n1511),.dout(n1513),.clk(gclk));
	jor g1213(.dina(n1513),.dinb(w_G411_0[2]),.dout(n1514),.clk(gclk));
	jand g1214(.dina(n1514),.dinb(n1510),.dout(n1515),.clk(gclk));
	jand g1215(.dina(w_G281_1[0]),.dinb(w_G248_3[0]),.dout(n1516),.clk(gclk));
	jand g1216(.dina(w_n530_0[2]),.dinb(w_G251_3[0]),.dout(n1517),.clk(gclk));
	jor g1217(.dina(n1517),.dinb(w_n532_1[0]),.dout(n1518),.clk(gclk));
	jor g1218(.dina(n1518),.dinb(w_dff_B_84LvMF523_1),.dout(n1519),.clk(gclk));
	jand g1219(.dina(w_n530_0[1]),.dinb(w_n406_3[0]),.dout(n1520),.clk(gclk));
	jand g1220(.dina(w_G281_0[2]),.dinb(w_n408_3[0]),.dout(n1521),.clk(gclk));
	jor g1221(.dina(n1521),.dinb(n1520),.dout(n1522),.clk(gclk));
	jor g1222(.dina(n1522),.dinb(w_G374_0[1]),.dout(n1523),.clk(gclk));
	jand g1223(.dina(n1523),.dinb(n1519),.dout(n1524),.clk(gclk));
	jxor g1224(.dina(n1524),.dinb(n1515),.dout(n1525),.clk(gclk));
	jor g1225(.dina(w_n483_1[0]),.dinb(w_n369_0[2]),.dout(n1526),.clk(gclk));
	jor g1226(.dina(w_G265_0[2]),.dinb(w_n366_0[2]),.dout(n1527),.clk(gclk));
	jand g1227(.dina(n1527),.dinb(w_G400_0[1]),.dout(n1528),.clk(gclk));
	jand g1228(.dina(n1528),.dinb(w_dff_B_61LdT2ER1_1),.dout(n1529),.clk(gclk));
	jor g1229(.dina(w_G265_0[1]),.dinb(w_G254_0[2]),.dout(n1530),.clk(gclk));
	jor g1230(.dina(w_n483_0[2]),.dinb(w_G242_0[2]),.dout(n1531),.clk(gclk));
	jand g1231(.dina(n1531),.dinb(w_dff_B_E6Ivhjnj0_1),.dout(n1532),.clk(gclk));
	jand g1232(.dina(n1532),.dinb(w_n485_0[2]),.dout(n1533),.clk(gclk));
	jor g1233(.dina(n1533),.dinb(n1529),.dout(n1534),.clk(gclk));
	jand g1234(.dina(w_G257_1[0]),.dinb(w_G248_2[2]),.dout(n1535),.clk(gclk));
	jand g1235(.dina(w_n518_0[2]),.dinb(w_G251_2[2]),.dout(n1536),.clk(gclk));
	jor g1236(.dina(n1536),.dinb(w_n520_0[0]),.dout(n1537),.clk(gclk));
	jor g1237(.dina(n1537),.dinb(w_dff_B_qUqFTHDw7_1),.dout(n1538),.clk(gclk));
	jand g1238(.dina(w_n518_0[1]),.dinb(w_n406_2[2]),.dout(n1539),.clk(gclk));
	jand g1239(.dina(w_G257_0[2]),.dinb(w_n408_2[2]),.dout(n1540),.clk(gclk));
	jor g1240(.dina(n1540),.dinb(n1539),.dout(n1541),.clk(gclk));
	jor g1241(.dina(n1541),.dinb(w_G389_0[1]),.dout(n1542),.clk(gclk));
	jand g1242(.dina(n1542),.dinb(n1538),.dout(n1543),.clk(gclk));
	jand g1243(.dina(w_G248_2[1]),.dinb(w_G234_1[0]),.dout(n1544),.clk(gclk));
	jand g1244(.dina(w_G251_2[1]),.dinb(w_n460_0[2]),.dout(n1545),.clk(gclk));
	jor g1245(.dina(n1545),.dinb(w_n462_0[0]),.dout(n1546),.clk(gclk));
	jor g1246(.dina(n1546),.dinb(w_dff_B_ak0qsddl7_1),.dout(n1547),.clk(gclk));
	jand g1247(.dina(w_n406_2[1]),.dinb(w_n460_0[1]),.dout(n1548),.clk(gclk));
	jand g1248(.dina(w_n408_2[1]),.dinb(w_G234_0[2]),.dout(n1549),.clk(gclk));
	jor g1249(.dina(n1549),.dinb(n1548),.dout(n1550),.clk(gclk));
	jor g1250(.dina(n1550),.dinb(w_G435_0[1]),.dout(n1551),.clk(gclk));
	jand g1251(.dina(n1551),.dinb(n1547),.dout(n1552),.clk(gclk));
	jxor g1252(.dina(n1552),.dinb(n1543),.dout(n1553),.clk(gclk));
	jxor g1253(.dina(n1553),.dinb(w_dff_B_Se3SyzF83_1),.dout(n1554),.clk(gclk));
	jxor g1254(.dina(n1554),.dinb(w_dff_B_BsXdgS7b2_1),.dout(n1555),.clk(gclk));
	jand g1255(.dina(w_G248_2[0]),.dinb(w_G226_1[0]),.dout(n1556),.clk(gclk));
	jand g1256(.dina(w_G251_2[0]),.dinb(w_n494_0[2]),.dout(n1557),.clk(gclk));
	jor g1257(.dina(n1557),.dinb(w_n496_0[1]),.dout(n1558),.clk(gclk));
	jor g1258(.dina(n1558),.dinb(w_dff_B_2COnfUBI7_1),.dout(n1559),.clk(gclk));
	jand g1259(.dina(w_n406_2[0]),.dinb(w_n494_0[1]),.dout(n1560),.clk(gclk));
	jand g1260(.dina(w_n408_2[0]),.dinb(w_G226_0[2]),.dout(n1561),.clk(gclk));
	jor g1261(.dina(n1561),.dinb(n1560),.dout(n1562),.clk(gclk));
	jor g1262(.dina(n1562),.dinb(w_G422_0[1]),.dout(n1563),.clk(gclk));
	jand g1263(.dina(n1563),.dinb(n1559),.dout(n1564),.clk(gclk));
	jxor g1264(.dina(n1564),.dinb(w_n551_0[0]),.dout(n1565),.clk(gclk));
	jor g1265(.dina(w_n369_0[1]),.dinb(w_n507_0[2]),.dout(n1566),.clk(gclk));
	jor g1266(.dina(w_n366_0[1]),.dinb(w_G218_1[0]),.dout(n1567),.clk(gclk));
	jand g1267(.dina(n1567),.dinb(w_G468_0[1]),.dout(n1568),.clk(gclk));
	jand g1268(.dina(n1568),.dinb(w_dff_B_gJhV3tqA0_1),.dout(n1569),.clk(gclk));
	jor g1269(.dina(w_G254_0[1]),.dinb(w_G218_0[2]),.dout(n1570),.clk(gclk));
	jor g1270(.dina(w_G242_0[1]),.dinb(w_n507_0[1]),.dout(n1571),.clk(gclk));
	jand g1271(.dina(n1571),.dinb(w_dff_B_UJdiGdRT3_1),.dout(n1572),.clk(gclk));
	jand g1272(.dina(n1572),.dinb(w_n509_0[0]),.dout(n1573),.clk(gclk));
	jor g1273(.dina(n1573),.dinb(n1569),.dout(n1574),.clk(gclk));
	jand g1274(.dina(w_G248_1[2]),.dinb(w_G210_1[0]),.dout(n1575),.clk(gclk));
	jand g1275(.dina(w_G251_1[2]),.dinb(w_n449_0[2]),.dout(n1576),.clk(gclk));
	jor g1276(.dina(n1576),.dinb(w_n451_0[0]),.dout(n1577),.clk(gclk));
	jor g1277(.dina(n1577),.dinb(w_dff_B_bsFFLQAk9_1),.dout(n1578),.clk(gclk));
	jand g1278(.dina(w_n406_1[2]),.dinb(w_n449_0[1]),.dout(n1579),.clk(gclk));
	jand g1279(.dina(w_n408_1[2]),.dinb(w_G210_0[2]),.dout(n1580),.clk(gclk));
	jor g1280(.dina(n1580),.dinb(n1579),.dout(n1581),.clk(gclk));
	jor g1281(.dina(n1581),.dinb(w_G457_0[1]),.dout(n1582),.clk(gclk));
	jand g1282(.dina(n1582),.dinb(n1578),.dout(n1583),.clk(gclk));
	jxor g1283(.dina(n1583),.dinb(n1574),.dout(n1584),.clk(gclk));
	jxor g1284(.dina(n1584),.dinb(n1565),.dout(n1585),.clk(gclk));
	jxor g1285(.dina(w_dff_B_QkIf4nKc5_0),.dinb(n1555),.dout(n1586),.clk(gclk));
	jand g1286(.dina(n1586),.dinb(w_n749_4[2]),.dout(n1587),.clk(gclk));
	jnot g1287(.din(n1587),.dout(n1588),.clk(gclk));
	jand g1288(.dina(w_n573_0[0]),.dinb(w_n567_0[0]),.dout(n1589),.clk(gclk));
	jor g1289(.dina(w_dff_B_Ucp90mZP1_0),.dinb(w_n699_0[0]),.dout(n1590),.clk(gclk));
	jnot g1290(.din(w_n559_0[0]),.dout(n1591),.clk(gclk));
	jor g1291(.dina(n1591),.dinb(w_n557_0[0]),.dout(n1592),.clk(gclk));
	jand g1292(.dina(w_n1592_0[1]),.dinb(w_n532_0[2]),.dout(n1593),.clk(gclk));
	jnot g1293(.din(w_n1593_0[1]),.dout(n1594),.clk(gclk));
	jor g1294(.dina(w_n695_0[0]),.dinb(n1594),.dout(n1595),.clk(gclk));
	jand g1295(.dina(w_n923_0[1]),.dinb(w_n473_0[2]),.dout(n1596),.clk(gclk));
	jor g1296(.dina(w_n1596_0[1]),.dinb(w_n1593_0[0]),.dout(n1597),.clk(gclk));
	jand g1297(.dina(w_dff_B_8Zp4ATZI9_0),.dinb(n1595),.dout(n1598),.clk(gclk));
	jxor g1298(.dina(w_dff_B_Vaz3kXuR5_0),.dinb(n1590),.dout(n1599),.clk(gclk));
	jnot g1299(.din(w_n1599_0[1]),.dout(n1600),.clk(gclk));
	jnot g1300(.din(w_n686_0[0]),.dout(n1601),.clk(gclk));
	jnot g1301(.din(w_n687_0[0]),.dout(n1602),.clk(gclk));
	jor g1302(.dina(w_n1592_0[0]),.dinb(w_n532_0[1]),.dout(n1603),.clk(gclk));
	jor g1303(.dina(w_n1596_0[0]),.dinb(w_n1603_0[1]),.dout(n1604),.clk(gclk));
	jor g1304(.dina(w_n923_0[0]),.dinb(w_n473_0[1]),.dout(n1605),.clk(gclk));
	jor g1305(.dina(w_n689_0[0]),.dinb(w_n485_0[1]),.dout(n1606),.clk(gclk));
	jand g1306(.dina(n1606),.dinb(w_n1605_0[1]),.dout(n1607),.clk(gclk));
	jand g1307(.dina(n1607),.dinb(n1604),.dout(n1608),.clk(gclk));
	jor g1308(.dina(n1608),.dinb(w_n690_0[0]),.dout(n1609),.clk(gclk));
	jor g1309(.dina(w_n1609_0[1]),.dinb(w_dff_B_EEf1xN4e2_1),.dout(n1610),.clk(gclk));
	jand g1310(.dina(n1610),.dinb(w_dff_B_ZBZ2h3Xx8_1),.dout(n1611),.clk(gclk));
	jand g1311(.dina(w_n1611_0[2]),.dinb(w_n581_0[0]),.dout(n1612),.clk(gclk));
	jxor g1312(.dina(w_n566_0[0]),.dinb(w_n561_0[1]),.dout(n1613),.clk(gclk));
	jxor g1313(.dina(w_n1613_0[1]),.dinb(w_n865_0[1]),.dout(n1614),.clk(gclk));
	jxor g1314(.dina(w_dff_B_Q7Fir2LH9_0),.dinb(n1612),.dout(n1615),.clk(gclk));
	jnot g1315(.din(w_n1615_0[1]),.dout(n1616),.clk(gclk));
	jand g1316(.dina(n1616),.dinb(w_dff_B_Is9FsIDa4_1),.dout(n1617),.clk(gclk));
	jnot g1317(.din(w_G1497_0[2]),.dout(n1618),.clk(gclk));
	jand g1318(.dina(w_n1615_0[0]),.dinb(w_n1599_0[0]),.dout(n1619),.clk(gclk));
	jor g1319(.dina(n1619),.dinb(w_n1618_0[1]),.dout(n1620),.clk(gclk));
	jor g1320(.dina(n1620),.dinb(n1617),.dout(n1621),.clk(gclk));
	jand g1321(.dina(w_n1605_0[0]),.dinb(w_n1603_0[0]),.dout(n1622),.clk(gclk));
	jor g1322(.dina(n1622),.dinb(w_n694_0[0]),.dout(n1623),.clk(gclk));
	jxor g1323(.dina(w_n1613_0[0]),.dinb(w_n1609_0[0]),.dout(n1624),.clk(gclk));
	jxor g1324(.dina(n1624),.dinb(w_dff_B_DPIhoEAz3_1),.dout(n1625),.clk(gclk));
	jxor g1325(.dina(w_n1611_0[1]),.dinb(w_n865_0[0]),.dout(n1626),.clk(gclk));
	jxor g1326(.dina(n1626),.dinb(w_dff_B_FDhpUtO37_1),.dout(n1627),.clk(gclk));
	jor g1327(.dina(n1627),.dinb(w_G1497_0[1]),.dout(n1628),.clk(gclk));
	jand g1328(.dina(w_dff_B_G6Afcqu25_0),.dinb(n1621),.dout(n1629),.clk(gclk));
	jxor g1329(.dina(w_n579_0[1]),.dinb(w_n574_0[0]),.dout(n1630),.clk(gclk));
	jxor g1330(.dina(w_dff_B_IEWSCVWl1_0),.dinb(n1629),.dout(n1631),.clk(gclk));
	jnot g1331(.din(w_n709_0[0]),.dout(n1632),.clk(gclk));
	jand g1332(.dina(n1632),.dinb(w_n953_0[0]),.dout(n1633),.clk(gclk));
	jand g1333(.dina(w_n711_0[0]),.dinb(w_n954_0[1]),.dout(n1634),.clk(gclk));
	jor g1334(.dina(n1634),.dinb(w_n1633_0[1]),.dout(n1635),.clk(gclk));
	jxor g1335(.dina(w_n608_0[0]),.dinb(w_n592_0[0]),.dout(n1636),.clk(gclk));
	jxor g1336(.dina(n1636),.dinb(w_n602_0[0]),.dout(n1637),.clk(gclk));
	jxor g1337(.dina(w_n1637_0[1]),.dinb(n1635),.dout(n1638),.clk(gclk));
	jor g1338(.dina(w_n938_0[1]),.dinb(w_n597_0[0]),.dout(n1639),.clk(gclk));
	jand g1339(.dina(w_n609_0[0]),.dinb(w_n962_0[0]),.dout(n1640),.clk(gclk));
	jor g1340(.dina(w_dff_B_E9c8Q9st3_0),.dinb(w_n715_0[0]),.dout(n1641),.clk(gclk));
	jand g1341(.dina(w_dff_B_UN3D2OQa0_0),.dinb(n1639),.dout(n1642),.clk(gclk));
	jxor g1342(.dina(n1642),.dinb(w_dff_B_5EK2mvuK0_1),.dout(n1643),.clk(gclk));
	jand g1343(.dina(w_n1643_0[1]),.dinb(w_n703_0[1]),.dout(n1644),.clk(gclk));
	jnot g1344(.din(w_n682_0[0]),.dout(n1645),.clk(gclk));
	jor g1345(.dina(w_n1611_0[0]),.dinb(w_n684_0[0]),.dout(n1646),.clk(gclk));
	jand g1346(.dina(n1646),.dinb(w_dff_B_gwOPQG2O0_1),.dout(n1647),.clk(gclk));
	jand g1347(.dina(w_n713_0[0]),.dinb(w_n954_0[0]),.dout(n1648),.clk(gclk));
	jor g1348(.dina(n1648),.dinb(w_n1633_0[0]),.dout(n1649),.clk(gclk));
	jxor g1349(.dina(w_dff_B_U39WYkVf8_0),.dinb(w_n938_0[0]),.dout(n1650),.clk(gclk));
	jxor g1350(.dina(n1650),.dinb(w_n1637_0[0]),.dout(n1651),.clk(gclk));
	jand g1351(.dina(n1651),.dinb(n1647),.dout(n1652),.clk(gclk));
	jor g1352(.dina(w_n1652_0[1]),.dinb(n1644),.dout(n1653),.clk(gclk));
	jor g1353(.dina(n1653),.dinb(w_G1497_0[0]),.dout(n1654),.clk(gclk));
	jnot g1354(.din(w_n588_1[0]),.dout(n1655),.clk(gclk));
	jand g1355(.dina(w_n1652_0[0]),.dinb(w_dff_B_7mRl6pvf8_1),.dout(n1656),.clk(gclk));
	jor g1356(.dina(w_n703_0[0]),.dinb(w_n588_0[2]),.dout(n1657),.clk(gclk));
	jand g1357(.dina(n1657),.dinb(w_n1643_0[0]),.dout(n1658),.clk(gclk));
	jor g1358(.dina(n1658),.dinb(n1656),.dout(n1659),.clk(gclk));
	jor g1359(.dina(n1659),.dinb(w_n1618_0[0]),.dout(n1660),.clk(gclk));
	jand g1360(.dina(n1660),.dinb(n1654),.dout(n1661),.clk(gclk));
	jxor g1361(.dina(n1661),.dinb(n1631),.dout(n1662),.clk(gclk));
	jor g1362(.dina(n1662),.dinb(w_n749_4[1]),.dout(n1663),.clk(gclk));
	jand g1363(.dina(n1663),.dinb(w_dff_B_uWVyz5F21_1),.dout(n1664),.clk(gclk));
	jor g1364(.dina(n1664),.dinb(w_G4092_3[2]),.dout(n1665),.clk(gclk));
	jor g1365(.dina(w_n1504_0[0]),.dinb(w_dff_B_2TsCaoR02_1),.dout(n1666),.clk(gclk));
	jand g1366(.dina(w_dff_B_VLqBh0GW4_0),.dinb(w_n1665_0[1]),.dout(w_dff_A_6B9aVpnN0_2),.clk(gclk));
	jor g1367(.dina(w_G4088_3[1]),.dinb(w_G14_0[1]),.dout(n1668),.clk(gclk));
	jor g1368(.dina(w_n797_3[1]),.dinb(w_G64_0[1]),.dout(n1669),.clk(gclk));
	jand g1369(.dina(n1669),.dinb(w_G4087_1[1]),.dout(n1670),.clk(gclk));
	jand g1370(.dina(n1670),.dinb(w_dff_B_CZWc9HjP5_1),.dout(n1671),.clk(gclk));
	jand g1371(.dina(w_G4092_3[1]),.dinb(G97),.dout(n1672),.clk(gclk));
	jnot g1372(.din(n1672),.dout(n1673),.clk(gclk));
	jand g1373(.dina(w_dff_B_nPiJfuQE9_0),.dinb(w_n1665_0[0]),.dout(n1674),.clk(gclk));
	jnot g1374(.din(w_n1674_0[2]),.dout(n1675),.clk(gclk));
	jor g1375(.dina(w_n1675_0[1]),.dinb(w_n797_3[0]),.dout(n1676),.clk(gclk));
	jand g1376(.dina(w_G4092_3[0]),.dinb(G94),.dout(n1677),.clk(gclk));
	jnot g1377(.din(n1677),.dout(n1678),.clk(gclk));
	jand g1378(.dina(w_dff_B_RNrhA1g56_0),.dinb(w_n1503_0[0]),.dout(n1679),.clk(gclk));
	jnot g1379(.din(w_n1679_0[2]),.dout(n1680),.clk(gclk));
	jor g1380(.dina(w_n1680_0[1]),.dinb(w_G4088_3[0]),.dout(n1681),.clk(gclk));
	jand g1381(.dina(n1681),.dinb(w_n800_1[1]),.dout(n1682),.clk(gclk));
	jand g1382(.dina(n1682),.dinb(w_dff_B_UuyVYPP90_1),.dout(n1683),.clk(gclk));
	jor g1383(.dina(n1683),.dinb(w_dff_B_l62URcUl6_1),.dout(w_dff_A_xjst1swX1_2),.clk(gclk));
	jor g1384(.dina(w_G4089_3[1]),.dinb(w_G14_0[0]),.dout(n1685),.clk(gclk));
	jor g1385(.dina(w_n852_3[1]),.dinb(w_G64_0[0]),.dout(n1686),.clk(gclk));
	jand g1386(.dina(n1686),.dinb(w_G4090_1[1]),.dout(n1687),.clk(gclk));
	jand g1387(.dina(n1687),.dinb(w_dff_B_X3poD1NW2_1),.dout(n1688),.clk(gclk));
	jor g1388(.dina(w_n1675_0[0]),.dinb(w_n852_3[0]),.dout(n1689),.clk(gclk));
	jor g1389(.dina(w_n1680_0[0]),.dinb(w_G4089_3[0]),.dout(n1690),.clk(gclk));
	jand g1390(.dina(n1690),.dinb(w_n854_1[1]),.dout(n1691),.clk(gclk));
	jand g1391(.dina(n1691),.dinb(w_dff_B_kT1rIe232_1),.dout(n1692),.clk(gclk));
	jor g1392(.dina(n1692),.dinb(w_dff_B_nzzW5EV01_1),.dout(w_dff_A_73jqJqeU4_2),.clk(gclk));
	jnot g1393(.din(w_G137_3[1]),.dout(n1694),.clk(gclk));
	jnot g1394(.din(G179),.dout(n1695),.clk(gclk));
	jnot g1395(.din(w_n996_1[1]),.dout(n1696),.clk(gclk));
	jor g1396(.dina(n1696),.dinb(w_n1695_0[1]),.dout(n1697),.clk(gclk));
	jnot g1397(.din(G176),.dout(n1698),.clk(gclk));
	jnot g1398(.din(w_n994_1[1]),.dout(n1699),.clk(gclk));
	jor g1399(.dina(n1699),.dinb(w_n1698_0[1]),.dout(n1700),.clk(gclk));
	jand g1400(.dina(w_n1674_0[1]),.dinb(w_G1689_1[2]),.dout(n1701),.clk(gclk));
	jand g1401(.dina(w_n1679_0[1]),.dinb(w_n993_1[1]),.dout(n1702),.clk(gclk));
	jor g1402(.dina(n1702),.dinb(w_G1690_0[1]),.dout(n1703),.clk(gclk));
	jor g1403(.dina(n1703),.dinb(w_dff_B_wFekHFN83_1),.dout(n1704),.clk(gclk));
	jand g1404(.dina(n1704),.dinb(w_dff_B_CohgHBSY3_1),.dout(n1705),.clk(gclk));
	jand g1405(.dina(n1705),.dinb(w_dff_B_avnGWs4K3_1),.dout(n1706),.clk(gclk));
	jor g1406(.dina(n1706),.dinb(w_n1694_0[1]),.dout(G658),.clk(gclk));
	jnot g1407(.din(w_n1012_1[1]),.dout(n1708),.clk(gclk));
	jor g1408(.dina(n1708),.dinb(w_n1695_0[0]),.dout(n1709),.clk(gclk));
	jnot g1409(.din(w_n1014_1[1]),.dout(n1710),.clk(gclk));
	jor g1410(.dina(n1710),.dinb(w_n1698_0[0]),.dout(n1711),.clk(gclk));
	jand g1411(.dina(w_n1674_0[0]),.dinb(w_G1691_1[2]),.dout(n1712),.clk(gclk));
	jand g1412(.dina(w_n1679_0[0]),.dinb(w_n1008_1[1]),.dout(n1713),.clk(gclk));
	jor g1413(.dina(n1713),.dinb(w_G1694_0[1]),.dout(n1714),.clk(gclk));
	jor g1414(.dina(n1714),.dinb(w_dff_B_b5XNq4Yj5_1),.dout(n1715),.clk(gclk));
	jand g1415(.dina(n1715),.dinb(w_dff_B_GxSbALLt5_1),.dout(n1716),.clk(gclk));
	jand g1416(.dina(n1716),.dinb(w_dff_B_C1gAIC6b5_1),.dout(n1717),.clk(gclk));
	jor g1417(.dina(n1717),.dinb(w_n1694_0[0]),.dout(G690),.clk(gclk));
	buf g1418(.din(w_G141_1[0]),.dout(w_dff_A_rVLNTSTJ6_1));
	buf g1419(.din(w_G293_0[0]),.dout(w_dff_A_66TVFEek2_1));
	buf g1420(.din(w_G3173_0[0]),.dout(w_dff_A_cOzPVBtM3_1));
	jnot g1421(.din(w_G545_0[1]),.dout(w_dff_A_IfMxj8Bd5_1),.clk(gclk));
	jnot g1422(.din(w_G545_0[0]),.dout(w_dff_A_O2Tzkydk6_1),.clk(gclk));
	buf g1423(.din(w_G137_3[0]),.dout(w_dff_A_7IidBGnj0_1));
	buf g1424(.din(w_G141_0[2]),.dout(w_dff_A_hGDXCrDc6_1));
	buf g1425(.din(w_G1_2[0]),.dout(w_dff_A_7dsw62mq4_1));
	buf g1426(.din(w_G549_0[1]),.dout(w_dff_A_c0W5v6CF5_1));
	buf g1427(.din(w_G299_0[1]),.dout(w_dff_A_acyZRsoC4_1));
	jnot g1428(.din(w_G549_0[0]),.dout(w_dff_A_b5bppP9C3_1),.clk(gclk));
	buf g1429(.din(w_G1_1[2]),.dout(w_dff_A_4QLAB4kJ6_1));
	buf g1430(.din(w_G1_1[1]),.dout(w_dff_A_5y0biOwJ6_1));
	buf g1431(.din(w_G1_1[0]),.dout(w_dff_A_S9WcFqMu6_1));
	buf g1432(.din(w_G1_0[2]),.dout(w_dff_A_HDNNfVWU5_1));
	buf g1433(.din(w_G299_0[0]),.dout(w_dff_A_GoPIL2KR7_1));
	jor g1434(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(w_dff_A_m2Bez7pJ5_2),.clk(gclk));
	jand g1435(.dina(w_n661_0[0]),.dinb(w_n641_0[1]),.dout(w_dff_A_Dg5KC4an0_2),.clk(gclk));
	jand g1436(.dina(w_n611_0[0]),.dinb(w_n588_0[1]),.dout(w_dff_A_zX1uAcE31_2),.clk(gclk));
	jor g1437(.dina(w_n717_0[0]),.dinb(w_n704_0[0]),.dout(w_dff_A_J8PJIiZa7_2),.clk(gclk));
	jor g1438(.dina(w_n747_0[0]),.dinb(w_n738_0[0]),.dout(w_dff_A_hRVgxDpe1_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_dff_A_xUQ57v087_1),.doutc(w_G4_0[2]),.din(w_dff_B_w06pBtwL9_3));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(G11));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(G14));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(w_dff_B_54uO2SaK2_2));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(w_dff_B_c1qR84vA7_2));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(w_dff_B_dDPN7lR71_2));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(w_dff_B_g02a7w813_2));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(G43));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(G46));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(w_dff_B_1iiDpNCJ1_2));
	jspl3 jspl3_w_G54_0(.douta(w_dff_A_DMJLjAWC3_0),.doutb(w_dff_A_pnV8RWif9_1),.doutc(w_G54_0[2]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(w_dff_B_SC9aAKpH0_2));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(w_dff_B_usrkDEF45_2));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(G67));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(w_dff_B_c7zUEjUl7_2));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(G73));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(G76));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(G91));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(G100));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(w_dff_B_TggzarqU3_2));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(w_dff_B_GunH8rOf0_2));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(G109));
	jspl jspl_w_G123_0(.douta(w_dff_A_nINmy0MP3_0),.doutb(w_G123_0[1]),.din(G123));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_kBbJ84pR7_0),.doutb(w_dff_A_4BTpAQXa4_1),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_rhf35aYN2_0),.doutb(w_dff_A_Wp9ZOKuG8_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_QWfpafDM6_0),.doutb(w_dff_A_ue7qSbSQ9_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_dff_A_sNwTwktN2_2),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_dff_A_8GZwz2KJ3_0),.doutb(w_dff_A_hhdMewAI5_1),.doutc(w_G137_4[2]),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_dff_A_kcz5qDe10_0),.doutb(w_G137_5[1]),.doutc(w_G137_5[2]),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_iKHdrdEq0_0),.doutb(w_dff_A_0CrxWVcA1_1),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_XY0BUQfE6_1),.doutc(w_dff_A_jG2qodlf0_2),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_G137_8[0]),.doutb(w_G137_8[1]),.doutc(w_dff_A_tbNmrbzc5_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_G137_9[0]),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_97f50Gyd7_1),.doutc(w_dff_A_2t5NEtJb8_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_qdReZtOb3_0),.doutb(w_dff_A_ISYTkH6Z2_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(w_dff_B_C5Gn2Iqp1_2));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(w_dff_B_4NUXgw828_2));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(w_dff_B_FBUy87R54_2));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(w_dff_B_4ob1Ejiw3_2));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(w_dff_B_UGVHS3ko5_2));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(w_dff_B_6HB1p32S0_2));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(w_dff_B_TbFIqqaD0_2));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(w_dff_B_9aXorsj56_2));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(w_dff_B_fV1F7oBh6_2));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(w_dff_B_3YGGGiVE7_2));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(w_dff_B_1nqnb48u7_2));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(w_dff_B_FgmiDBhq7_2));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(w_dff_B_HOpJCSUc9_2));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(w_dff_B_9a14oI2n7_2));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(w_dff_B_Rz0P6yzV7_2));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(w_dff_B_VgeiRaJZ6_2));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(w_dff_B_Zm4pvZX48_2));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(w_dff_B_sdn6Tn8o5_2));
	jspl3 jspl3_w_G206_0(.douta(w_G206_0[0]),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G206_1(.douta(w_dff_A_1F6tAt515_0),.doutb(w_G206_1[1]),.doutc(w_G206_1[2]),.din(w_G206_0[0]));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_dff_A_VsQiZBHr3_2),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_G210_1[1]),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl jspl_w_G210_2(.douta(w_dff_A_omW0t1800_0),.doutb(w_G210_2[1]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_dff_A_2dgVSwNM7_0),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl jspl_w_G218_2(.douta(w_dff_A_snz3ufaQ5_0),.doutb(w_G218_2[1]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_dff_A_YFIgcURp7_2),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_G226_1[0]),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl jspl_w_G226_2(.douta(w_dff_A_vLQ3zUm74_0),.doutb(w_G226_2[1]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_dff_A_Vdnrw3Gg7_2),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_dff_A_fMp54LYZ8_0),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_dff_A_dC6B2DkC2_1),.doutc(w_dff_A_ep1c18em2_2),.din(G242));
	jspl jspl_w_G242_1(.douta(w_dff_A_SykPmhEG9_0),.doutb(w_G242_1[1]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_dff_A_TUtlYu8p7_0),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_dff_A_A874vAr96_2),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl3 jspl3_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.doutc(w_G248_5[2]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_dff_A_ag2tn0BI5_1),.doutc(w_dff_A_wZ2op9mq3_2),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_dff_A_AB26oXG68_0),.doutb(w_G251_1[1]),.doutc(w_dff_A_Xcenn3811_2),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_G251_4[1]),.doutc(w_G251_4[2]),.din(w_G251_1[0]));
	jspl jspl_w_G251_5(.douta(w_dff_A_AN3A2DOu0_0),.doutb(w_G251_5[1]),.din(w_G251_1[1]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl jspl_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_dff_A_UCUdfuzf8_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_G257_1[0]),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl jspl_w_G257_2(.douta(w_dff_A_9iZVWSZd3_0),.doutb(w_G257_2[1]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_dff_A_oVA4nxdI7_2),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_dff_A_xejFgTk11_1),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_dff_A_Xnc6CWE06_2),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_dff_A_XDgcLo2e7_1),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl jspl_w_G273_2(.douta(w_dff_A_HxChay362_0),.doutb(w_G273_2[1]),.din(w_G273_0[1]));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_dff_A_n0anY7p45_2),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_dff_A_SsgkcA2G8_0),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_G289_0[0]),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_dff_A_kZSg5MXX5_1),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_dff_A_eWQJRtlK4_0),.doutb(w_dff_A_6kitU1zB8_1),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_dff_A_NuoaZjgQ1_0),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_dff_A_Sb7QOQec3_2),.din(G316));
	jspl jspl_w_G316_1(.douta(w_G316_1[0]),.doutb(w_G316_1[1]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_G324_0[1]),.doutc(w_dff_A_m0hJMGqo6_2),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_dff_A_S9P1YKLL9_1),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_dff_A_TLSq3PvQ6_1),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_dff_A_WSnSbauz7_1),.doutc(w_G332_1[2]),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_dff_A_JKLtRAxP4_0),.doutb(w_G332_2[1]),.doutc(w_dff_A_Fq3Yi8Dz9_2),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_G332_3[0]),.doutb(w_G332_3[1]),.doutc(w_G332_3[2]),.din(w_G332_0[2]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl jspl_w_G338_0(.douta(w_dff_A_6D4cYah37_0),.doutb(w_G338_0[1]),.din(G338));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_dff_A_Sl0epb350_2),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_dff_A_m2qxj6TM4_1),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_dff_A_hcovNpaa2_0),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_dff_A_Tw4If2hQ9_2),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_G351_1[0]),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_dff_A_eRUhx5PH6_1),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_dff_A_5xH6wiIu1_0),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_G361_0[1]),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G361_1(.douta(w_dff_A_p0Cf2Y2O2_0),.doutb(w_G361_1[1]),.din(w_G361_0[0]));
	jspl jspl_w_G366_0(.douta(w_dff_A_Foq3VPLQ3_0),.doutb(w_G366_0[1]),.din(G366));
	jspl jspl_w_G369_0(.douta(w_G369_0[0]),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_G374_0[0]),.doutb(w_dff_A_4pKE69fy7_1),.doutc(w_dff_A_CHL3mOnJ1_2),.din(G374));
	jspl3 jspl3_w_G374_1(.douta(w_dff_A_NCvTwNFW0_0),.doutb(w_dff_A_ZHtEhEHW0_1),.doutc(w_G374_1[2]),.din(w_G374_0[0]));
	jspl3 jspl3_w_G389_0(.douta(w_G389_0[0]),.doutb(w_dff_A_4Ezae2bB4_1),.doutc(w_dff_A_spaQFyFL5_2),.din(G389));
	jspl3 jspl3_w_G389_1(.douta(w_dff_A_JzflguxI3_0),.doutb(w_dff_A_tMFfg7EN9_1),.doutc(w_G389_1[2]),.din(w_G389_0[0]));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_dff_A_RyuxyeXw5_1),.doutc(w_dff_A_UIuZFd6I2_2),.din(G400));
	jspl3 jspl3_w_G400_1(.douta(w_dff_A_kQSqkvHw5_0),.doutb(w_dff_A_lS1IRETb5_1),.doutc(w_G400_1[2]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_dff_A_BVx3UiRc1_0),.doutb(w_G411_0[1]),.doutc(w_dff_A_lV1aM1ki1_2),.din(G411));
	jspl3 jspl3_w_G411_1(.douta(w_G411_1[0]),.doutb(w_G411_1[1]),.doutc(w_G411_1[2]),.din(w_G411_0[0]));
	jspl jspl_w_G411_2(.douta(w_dff_A_vZS4jv8O6_0),.doutb(w_G411_2[1]),.din(w_G411_0[1]));
	jspl3 jspl3_w_G422_0(.douta(w_G422_0[0]),.doutb(w_dff_A_ihL37Hwh1_1),.doutc(w_dff_A_RGIhfKH47_2),.din(G422));
	jspl jspl_w_G422_1(.douta(w_dff_A_4FNS6t941_0),.doutb(w_G422_1[1]),.din(w_G422_0[0]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_dff_A_BvM1Ub6G2_1),.doutc(w_dff_A_VR5MfvCi8_2),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_dff_A_wpZAXwbu1_0),.doutb(w_dff_A_LDaXALsP2_1),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_dff_A_DwvbHT6D0_1),.doutc(w_dff_A_f2gP5ZVl5_2),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_dff_A_cdMgZoFv3_0),.doutb(w_dff_A_vPJtS8657_1),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_G457_0[0]),.doutb(w_dff_A_JYLhTTJa8_1),.doutc(w_dff_A_YnWKwscH0_2),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_dff_A_zRCf7qQ64_0),.doutb(w_dff_A_rP4Wqp0u9_1),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_dff_A_gqiZzrv91_1),.doutc(w_dff_A_oN5HW0EJ7_2),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_dff_A_NyAn2Iwl2_0),.doutb(w_dff_A_zp28VQpV5_1),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_dff_A_zu46DcNC2_0),.doutb(w_dff_A_nmvMlbAs9_1),.doutc(w_G479_0[2]),.din(G479));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_dff_A_JWxZI3X23_1),.doutc(w_dff_A_iD7IMbK61_2),.din(G490));
	jspl jspl_w_G490_1(.douta(w_dff_A_FUOC17pp8_0),.doutb(w_G490_1[1]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_dff_A_TkQf8VUZ5_0),.doutb(w_G503_0[1]),.doutc(w_dff_A_z10QLZuZ2_2),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_G503_1[0]),.doutb(w_G503_1[1]),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl jspl_w_G503_2(.douta(w_dff_A_TVETGGw30_0),.doutb(w_G503_2[1]),.din(w_G503_0[1]));
	jspl3 jspl3_w_G514_0(.douta(w_dff_A_gqGYYdE64_0),.doutb(w_G514_0[1]),.doutc(w_dff_A_qQCaPRpQ6_2),.din(G514));
	jspl3 jspl3_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.doutc(w_G514_1[2]),.din(w_G514_0[0]));
	jspl jspl_w_G514_2(.douta(w_G514_2[0]),.doutb(w_G514_2[1]),.din(w_G514_0[1]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_dff_A_Aw05G7vG7_1),.doutc(w_dff_A_3nvPKuqC5_2),.din(G523));
	jspl3 jspl3_w_G523_1(.douta(w_dff_A_9mALEgny1_0),.doutb(w_dff_A_5pSo3KrS6_1),.doutc(w_G523_1[2]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_dff_A_IDL7g5my3_0),.doutb(w_G534_0[1]),.doutc(w_dff_A_MOvQLspi1_2),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_G534_1[0]),.doutb(w_G534_1[1]),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl jspl_w_G534_2(.douta(w_dff_A_KpExEhaJ8_0),.doutb(w_G534_2[1]),.din(w_G534_0[1]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_dff_A_3Ccg3jVJ7_0),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_dff_A_DIXrA4Ol2_0),.doutb(w_dff_A_kMGXyWAW2_1),.doutc(w_G1497_0[2]),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_dff_A_v8UhOTPX0_1),.doutc(w_dff_A_Xl6d13p94_2),.din(G1689));
	jspl3 jspl3_w_G1689_1(.douta(w_dff_A_b7Fpg7u54_0),.doutb(w_G1689_1[1]),.doutc(w_dff_A_Kyriajg40_2),.din(w_G1689_0[0]));
	jspl3 jspl3_w_G1689_2(.douta(w_dff_A_HJZRrLEG4_0),.doutb(w_G1689_2[1]),.doutc(w_dff_A_zKLX45dN3_2),.din(w_G1689_0[1]));
	jspl3 jspl3_w_G1689_3(.douta(w_dff_A_9L5JHhJU6_0),.doutb(w_dff_A_JUUW9lsD8_1),.doutc(w_G1689_3[2]),.din(w_G1689_0[2]));
	jspl3 jspl3_w_G1689_4(.douta(w_dff_A_RaJD5xjh5_0),.doutb(w_dff_A_6BM9BGGk0_1),.doutc(w_G1689_4[2]),.din(w_G1689_1[0]));
	jspl jspl_w_G1689_5(.douta(w_G1689_5[0]),.doutb(w_G1689_5[1]),.din(w_G1689_1[1]));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_dff_A_XlP6CFhZ0_1),.doutc(w_G1690_0[2]),.din(G1690));
	jspl jspl_w_G1690_1(.douta(w_G1690_1[0]),.doutb(w_dff_A_c6VJc8HF5_1),.din(w_G1690_0[0]));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_dff_A_cCDNMOeN8_1),.doutc(w_dff_A_23j1qrul6_2),.din(G1691));
	jspl3 jspl3_w_G1691_1(.douta(w_G1691_1[0]),.doutb(w_G1691_1[1]),.doutc(w_dff_A_eJwSTwYZ2_2),.din(w_G1691_0[0]));
	jspl3 jspl3_w_G1691_2(.douta(w_dff_A_tKb3P4l32_0),.doutb(w_G1691_2[1]),.doutc(w_dff_A_XGBsZiXQ1_2),.din(w_G1691_0[1]));
	jspl3 jspl3_w_G1691_3(.douta(w_dff_A_TIcULKQy2_0),.doutb(w_dff_A_AyyJTQSO9_1),.doutc(w_G1691_3[2]),.din(w_G1691_0[2]));
	jspl3 jspl3_w_G1691_4(.douta(w_dff_A_B8nvlZ5P7_0),.doutb(w_dff_A_QDiPIroo4_1),.doutc(w_G1691_4[2]),.din(w_G1691_1[0]));
	jspl jspl_w_G1691_5(.douta(w_G1691_5[0]),.doutb(w_dff_A_3RYyMW4v3_1),.din(w_G1691_1[1]));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_dff_A_maasZoqd6_1),.doutc(w_dff_A_iSQ5fhzh9_2),.din(G1694));
	jspl jspl_w_G1694_1(.douta(w_G1694_1[0]),.doutb(w_G1694_1[1]),.din(w_G1694_0[0]));
	jspl3 jspl3_w_G2174_0(.douta(w_dff_A_m2APYiOi5_0),.doutb(w_dff_A_aQ2sne377_1),.doutc(w_G2174_0[2]),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_dff_A_Zx3hLzlE1_0),.doutb(w_dff_A_5ZzhKa771_1),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(w_dff_B_qq3Zf2UL4_3));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_dff_A_5ks2fcuz9_0),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_G3724_0[0]),.doutb(w_G3724_0[1]),.doutc(w_dff_A_dOM0HN591_2),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_dff_A_z4gXNJDl6_1),.doutc(w_dff_A_RCIjzLbv0_2),.din(G4087));
	jspl3 jspl3_w_G4087_1(.douta(w_G4087_1[0]),.doutb(w_dff_A_jiFySq680_1),.doutc(w_dff_A_5ViwmFPS6_2),.din(w_G4087_0[0]));
	jspl3 jspl3_w_G4087_2(.douta(w_G4087_2[0]),.doutb(w_G4087_2[1]),.doutc(w_G4087_2[2]),.din(w_G4087_0[1]));
	jspl3 jspl3_w_G4087_3(.douta(w_G4087_3[0]),.doutb(w_G4087_3[1]),.doutc(w_G4087_3[2]),.din(w_G4087_0[2]));
	jspl3 jspl3_w_G4087_4(.douta(w_dff_A_s4mXJW8X6_0),.doutb(w_dff_A_sg5nOhNJ8_1),.doutc(w_G4087_4[2]),.din(w_G4087_1[0]));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_G4088_0[2]),.din(G4088));
	jspl3 jspl3_w_G4088_1(.douta(w_G4088_1[0]),.doutb(w_G4088_1[1]),.doutc(w_G4088_1[2]),.din(w_G4088_0[0]));
	jspl3 jspl3_w_G4088_2(.douta(w_G4088_2[0]),.doutb(w_G4088_2[1]),.doutc(w_G4088_2[2]),.din(w_G4088_0[1]));
	jspl3 jspl3_w_G4088_3(.douta(w_dff_A_a1YkzlzF7_0),.doutb(w_G4088_3[1]),.doutc(w_G4088_3[2]),.din(w_G4088_0[2]));
	jspl3 jspl3_w_G4088_4(.douta(w_dff_A_7Swbm09q8_0),.doutb(w_G4088_4[1]),.doutc(w_dff_A_pjKoofEh2_2),.din(w_G4088_1[0]));
	jspl3 jspl3_w_G4088_5(.douta(w_G4088_5[0]),.doutb(w_dff_A_FHmdRqKn5_1),.doutc(w_G4088_5[2]),.din(w_G4088_1[1]));
	jspl3 jspl3_w_G4088_6(.douta(w_dff_A_ckOVcIE78_0),.doutb(w_G4088_6[1]),.doutc(w_dff_A_FCfSnQoz9_2),.din(w_G4088_1[2]));
	jspl3 jspl3_w_G4088_7(.douta(w_G4088_7[0]),.doutb(w_dff_A_NO74DbYq5_1),.doutc(w_G4088_7[2]),.din(w_G4088_2[0]));
	jspl3 jspl3_w_G4088_8(.douta(w_dff_A_vhDY77Uo2_0),.doutb(w_G4088_8[1]),.doutc(w_dff_A_DjpfCeFM4_2),.din(w_G4088_2[1]));
	jspl3 jspl3_w_G4088_9(.douta(w_G4088_9[0]),.doutb(w_dff_A_rup8d4tL5_1),.doutc(w_G4088_9[2]),.din(w_G4088_2[2]));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_G4089_0[2]),.din(G4089));
	jspl3 jspl3_w_G4089_1(.douta(w_G4089_1[0]),.doutb(w_G4089_1[1]),.doutc(w_G4089_1[2]),.din(w_G4089_0[0]));
	jspl3 jspl3_w_G4089_2(.douta(w_G4089_2[0]),.doutb(w_G4089_2[1]),.doutc(w_G4089_2[2]),.din(w_G4089_0[1]));
	jspl3 jspl3_w_G4089_3(.douta(w_dff_A_RKaJPw4R7_0),.doutb(w_G4089_3[1]),.doutc(w_G4089_3[2]),.din(w_G4089_0[2]));
	jspl3 jspl3_w_G4089_4(.douta(w_dff_A_bkjNZIKN0_0),.doutb(w_G4089_4[1]),.doutc(w_dff_A_fggixee15_2),.din(w_G4089_1[0]));
	jspl3 jspl3_w_G4089_5(.douta(w_G4089_5[0]),.doutb(w_dff_A_2M1RsakX4_1),.doutc(w_dff_A_hd8QYJlY8_2),.din(w_G4089_1[1]));
	jspl3 jspl3_w_G4089_6(.douta(w_G4089_6[0]),.doutb(w_G4089_6[1]),.doutc(w_dff_A_aqR0O6v62_2),.din(w_G4089_1[2]));
	jspl3 jspl3_w_G4089_7(.douta(w_dff_A_oas7hLWv3_0),.doutb(w_G4089_7[1]),.doutc(w_dff_A_caZmU7uz2_2),.din(w_G4089_2[0]));
	jspl3 jspl3_w_G4089_8(.douta(w_G4089_8[0]),.doutb(w_dff_A_2ssKatZa8_1),.doutc(w_G4089_8[2]),.din(w_G4089_2[1]));
	jspl3 jspl3_w_G4089_9(.douta(w_G4089_9[0]),.doutb(w_dff_A_U89a4rlK1_1),.doutc(w_G4089_9[2]),.din(w_G4089_2[2]));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_dff_A_REUvvtvf3_1),.doutc(w_dff_A_W5GRnw7Q9_2),.din(G4090));
	jspl3 jspl3_w_G4090_1(.douta(w_G4090_1[0]),.doutb(w_dff_A_UJNqLQE41_1),.doutc(w_dff_A_8bKgs9nA1_2),.din(w_G4090_0[0]));
	jspl3 jspl3_w_G4090_2(.douta(w_G4090_2[0]),.doutb(w_G4090_2[1]),.doutc(w_dff_A_oG5NCBMF8_2),.din(w_G4090_0[1]));
	jspl3 jspl3_w_G4090_3(.douta(w_G4090_3[0]),.doutb(w_dff_A_3CliLQJe9_1),.doutc(w_dff_A_sJEdiHEr5_2),.din(w_G4090_0[2]));
	jspl3 jspl3_w_G4090_4(.douta(w_dff_A_yU2mtP1v8_0),.doutb(w_dff_A_wsrgcQzq2_1),.doutc(w_G4090_4[2]),.din(w_G4090_1[0]));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_dff_A_IS6nQ2ra3_1),.doutc(w_dff_A_Bwnsjr1H9_2),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_dff_A_wCjJ2qrj9_0),.doutb(w_dff_A_9pW0ku0l4_1),.doutc(w_G4091_1[2]),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_dff_A_hcjprUEn9_0),.doutb(w_dff_A_cF2zdSL49_1),.doutc(w_G4091_2[2]),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4091_3(.douta(w_G4091_3[0]),.doutb(w_dff_A_IkAbCPM81_1),.doutc(w_dff_A_wM42BPhe6_2),.din(w_G4091_0[2]));
	jspl3 jspl3_w_G4091_4(.douta(w_dff_A_NGs4s4Vo9_0),.doutb(w_G4091_4[1]),.doutc(w_dff_A_jFYyJij92_2),.din(w_G4091_1[0]));
	jspl3 jspl3_w_G4091_5(.douta(w_dff_A_wJpX3Al28_0),.doutb(w_G4091_5[1]),.doutc(w_dff_A_2NvsHdUV5_2),.din(w_G4091_1[1]));
	jspl jspl_w_G4091_6(.douta(w_dff_A_abu6zKXv4_0),.doutb(w_G4091_6[1]),.din(w_G4091_1[2]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_dff_A_zpumRBPU4_1),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_dff_A_96sSh9NM1_0),.doutb(w_G4092_1[1]),.doutc(w_dff_A_VHMWrw1t4_2),.din(w_G4092_0[0]));
	jspl3 jspl3_w_G4092_2(.douta(w_dff_A_wMAhAGCw2_0),.doutb(w_dff_A_ggGHQquF5_1),.doutc(w_G4092_2[2]),.din(w_G4092_0[1]));
	jspl3 jspl3_w_G4092_3(.douta(w_G4092_3[0]),.doutb(w_G4092_3[1]),.doutc(w_dff_A_QiMycBOG7_2),.din(w_G4092_0[2]));
	jspl3 jspl3_w_G4092_4(.douta(w_dff_A_4eBVXyyi9_0),.doutb(w_G4092_4[1]),.doutc(w_G4092_4[2]),.din(w_G4092_1[0]));
	jspl3 jspl3_w_G4092_5(.douta(w_dff_A_1EefmUZz0_0),.doutb(w_dff_A_ggjRFm5I5_1),.doutc(w_G4092_5[2]),.din(w_G4092_1[1]));
	jspl3 jspl3_w_G4092_6(.douta(w_G4092_6[0]),.doutb(w_dff_A_mBnuKcvg5_1),.doutc(w_dff_A_naL09aep2_2),.din(w_G4092_1[2]));
	jspl3 jspl3_w_G4092_7(.douta(w_G4092_7[0]),.doutb(w_G4092_7[1]),.doutc(w_dff_A_HTohEeBT0_2),.din(w_G4092_2[0]));
	jspl3 jspl3_w_G4092_8(.douta(w_G4092_8[0]),.doutb(w_dff_A_AnjC0Ijo8_1),.doutc(w_dff_A_SwxSWY5E6_2),.din(w_G4092_2[1]));
	jspl3 jspl3_w_G4092_9(.douta(w_dff_A_ifR6nME50_0),.doutb(w_dff_A_RhMIT62F1_1),.doutc(w_G4092_9[2]),.din(w_G4092_2[2]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(w_dff_A_LWbmaDOx7_1),.din(G599_fa_));
	jspl jspl_w_G601_0(.douta(w_G601_0),.doutb(w_dff_A_ErVd9dvY1_1),.din(G601_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(w_dff_A_H84LiIAI2_1),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_G809_1[0]),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_G809_2[2]),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_G809_3[0]),.doutb(w_G809_3[1]),.doutc(w_dff_A_a0LYu7n60_2),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(w_dff_A_ww1qOiDN8_1),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(w_dff_A_SdU8Ychv1_1),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(w_dff_A_a58wHPnb2_1),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(w_dff_A_32PGN2ft4_1),.din(G861_fa_));
	jspl jspl_w_G623_0(.douta(w_G623_0),.doutb(w_dff_A_3zZlppPo2_1),.din(G623_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(w_dff_A_J4Jmmsg98_1),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(w_dff_A_BZPX3kBd6_1),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(w_dff_A_YrJpRzMx9_1),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(w_dff_A_mblDQHA37_1),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(w_dff_A_xLUN1R8u8_1),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(w_dff_A_ze09dhrl2_1),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(w_dff_A_5ypKyrfN3_1),.din(G877_fa_));
	jspl jspl_w_G998_0(.douta(w_G998_0),.doutb(w_dff_A_neliHUfR6_1),.din(G998_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(w_dff_A_RKhsEVmw6_1),.din(G830_fa_));
	jspl jspl_w_G865_0(.douta(w_G865_0),.doutb(w_dff_A_cJBm3tzC8_1),.din(G865_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(w_dff_A_j23ZqMUB9_1),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(w_dff_B_C8HPys6d9_2));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.doutc(w_n369_0[2]),.din(n369));
	jspl3 jspl3_w_n369_1(.douta(w_n369_1[0]),.doutb(w_n369_1[1]),.doutc(w_n369_1[2]),.din(w_n369_0[0]));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl3 jspl3_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.doutc(w_n374_0[2]),.din(n374));
	jspl jspl_w_n374_1(.douta(w_n374_1[0]),.doutb(w_n374_1[1]),.din(w_n374_0[0]));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl3 jspl3_w_n375_1(.douta(w_n375_1[0]),.doutb(w_n375_1[1]),.doutc(w_n375_1[2]),.din(w_n375_0[0]));
	jspl3 jspl3_w_n375_2(.douta(w_n375_2[0]),.doutb(w_n375_2[1]),.doutc(w_n375_2[2]),.din(w_n375_0[1]));
	jspl3 jspl3_w_n375_3(.douta(w_n375_3[0]),.doutb(w_n375_3[1]),.doutc(w_n375_3[2]),.din(w_n375_0[2]));
	jspl3 jspl3_w_n375_4(.douta(w_n375_4[0]),.doutb(w_n375_4[1]),.doutc(w_n375_4[2]),.din(w_n375_1[0]));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_dff_A_tfjwpnlU9_2),.din(w_dff_B_wOVfCONj9_3));
	jspl jspl_w_n377_1(.douta(w_dff_A_wTccKRfM2_0),.doutb(w_n377_1[1]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.doutc(w_n378_0[2]),.din(n378));
	jspl3 jspl3_w_n378_1(.douta(w_n378_1[0]),.doutb(w_n378_1[1]),.doutc(w_n378_1[2]),.din(w_n378_0[0]));
	jspl3 jspl3_w_n378_2(.douta(w_n378_2[0]),.doutb(w_n378_2[1]),.doutc(w_n378_2[2]),.din(w_n378_0[1]));
	jspl3 jspl3_w_n378_3(.douta(w_n378_3[0]),.doutb(w_n378_3[1]),.doutc(w_n378_3[2]),.din(w_n378_0[2]));
	jspl3 jspl3_w_n378_4(.douta(w_n378_4[0]),.doutb(w_n378_4[1]),.doutc(w_n378_4[2]),.din(w_n378_1[0]));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_dff_A_gkmhSzvi0_2),.din(w_dff_B_84Cmest04_3));
	jspl jspl_w_n389_1(.douta(w_dff_A_glcBLkLD3_0),.doutb(w_n389_1[1]),.din(w_n389_0[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n401_0(.douta(w_dff_A_s8jJaLwc5_0),.doutb(w_n401_0[1]),.din(w_dff_B_XuwBpfWG4_2));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.doutc(w_n406_0[2]),.din(n406));
	jspl3 jspl3_w_n406_1(.douta(w_n406_1[0]),.doutb(w_n406_1[1]),.doutc(w_n406_1[2]),.din(w_n406_0[0]));
	jspl3 jspl3_w_n406_2(.douta(w_n406_2[0]),.doutb(w_n406_2[1]),.doutc(w_n406_2[2]),.din(w_n406_0[1]));
	jspl3 jspl3_w_n406_3(.douta(w_n406_3[0]),.doutb(w_n406_3[1]),.doutc(w_n406_3[2]),.din(w_n406_0[2]));
	jspl3 jspl3_w_n406_4(.douta(w_n406_4[0]),.doutb(w_n406_4[1]),.doutc(w_n406_4[2]),.din(w_n406_1[0]));
	jspl jspl_w_n406_5(.douta(w_n406_5[0]),.doutb(w_n406_5[1]),.din(w_n406_1[1]));
	jspl3 jspl3_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.doutc(w_n408_0[2]),.din(n408));
	jspl3 jspl3_w_n408_1(.douta(w_n408_1[0]),.doutb(w_n408_1[1]),.doutc(w_n408_1[2]),.din(w_n408_0[0]));
	jspl3 jspl3_w_n408_2(.douta(w_n408_2[0]),.doutb(w_n408_2[1]),.doutc(w_n408_2[2]),.din(w_n408_0[1]));
	jspl3 jspl3_w_n408_3(.douta(w_n408_3[0]),.doutb(w_n408_3[1]),.doutc(w_n408_3[2]),.din(w_n408_0[2]));
	jspl3 jspl3_w_n408_4(.douta(w_n408_4[0]),.doutb(w_n408_4[1]),.doutc(w_n408_4[2]),.din(w_n408_1[0]));
	jspl3 jspl3_w_n408_5(.douta(w_n408_5[0]),.doutb(w_n408_5[1]),.doutc(w_n408_5[2]),.din(w_n408_1[1]));
	jspl3 jspl3_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.doutc(w_n412_0[2]),.din(n412));
	jspl jspl_w_n414_0(.douta(w_dff_A_PNkC3uu93_0),.doutb(w_n414_0[1]),.din(w_dff_B_jI44hNRp8_2));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl3 jspl3_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.doutc(w_n423_0[2]),.din(n423));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_n425_0[2]),.din(n425));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_dff_A_0YSAPy1G7_1),.doutc(w_n428_0[2]),.din(n428));
	jspl jspl_w_n428_1(.douta(w_n428_1[0]),.doutb(w_dff_A_5EHyocmY4_1),.din(w_n428_0[0]));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl3 jspl3_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.doutc(w_n433_0[2]),.din(n433));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl jspl_w_n435_2(.douta(w_n435_2[0]),.doutb(w_n435_2[1]),.din(w_n435_0[1]));
	jspl jspl_w_n437_0(.douta(w_dff_A_DA9kbywb7_0),.doutb(w_n437_0[1]),.din(w_dff_B_y3kByK1p7_2));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_dff_A_sxn8HzZ62_1),.doutc(w_n451_0[2]),.din(w_dff_B_258BLKiQ6_3));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_dff_A_JxHJl6d94_1),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_QQ58oc3Q7_1),.doutc(w_n462_0[2]),.din(w_dff_B_4IsApSZi4_3));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl3 jspl3_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.doutc(w_n471_1[2]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_dff_A_eeLzT7dy9_1),.doutc(w_dff_A_kK2bVqdC6_2),.din(w_dff_B_t2bDAX2O6_3));
	jspl jspl_w_n473_1(.douta(w_n473_1[0]),.doutb(w_n473_1[1]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.doutc(w_n483_0[2]),.din(n483));
	jspl3 jspl3_w_n483_1(.douta(w_n483_1[0]),.doutb(w_n483_1[1]),.doutc(w_n483_1[2]),.din(w_n483_0[0]));
	jspl jspl_w_n483_2(.douta(w_n483_2[0]),.doutb(w_n483_2[1]),.din(w_n483_0[1]));
	jspl3 jspl3_w_n485_0(.douta(w_n485_0[0]),.doutb(w_dff_A_WxCttBwT4_1),.doutc(w_dff_A_MkVZMfz07_2),.din(w_dff_B_Vi4jOAZY0_3));
	jspl jspl_w_n485_1(.douta(w_dff_A_S32Xyl0Y1_0),.doutb(w_n485_1[1]),.din(w_n485_0[0]));
	jspl jspl_w_n493_0(.douta(w_n493_0[0]),.doutb(w_n493_0[1]),.din(n493));
	jspl3 jspl3_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.doutc(w_n494_0[2]),.din(n494));
	jspl3 jspl3_w_n494_1(.douta(w_n494_1[0]),.doutb(w_n494_1[1]),.doutc(w_n494_1[2]),.din(w_n494_0[0]));
	jspl3 jspl3_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.doutc(w_dff_A_du6Mz9Sf0_2),.din(w_dff_B_6xukRhGQ8_3));
	jspl jspl_w_n496_1(.douta(w_dff_A_eYoFTxR21_0),.doutb(w_n496_1[1]),.din(w_n496_0[0]));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl3 jspl3_w_n509_0(.douta(w_dff_A_NUipEbn84_0),.doutb(w_dff_A_oZTYeJI77_1),.doutc(w_n509_0[2]),.din(w_dff_B_Ue2RQK7M0_3));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl3 jspl3_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.doutc(w_n518_1[2]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n520_0(.douta(w_n520_0[0]),.doutb(w_dff_A_nw1q9Y2Y4_1),.doutc(w_n520_0[2]),.din(w_dff_B_kmWkYj5y6_3));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl3 jspl3_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.doutc(w_n530_1[2]),.din(w_n530_0[0]));
	jspl3 jspl3_w_n532_0(.douta(w_n532_0[0]),.doutb(w_dff_A_IK6a6du75_1),.doutc(w_dff_A_dGVpQ0Fx4_2),.din(w_dff_B_bVA2yGk26_3));
	jspl jspl_w_n532_1(.douta(w_n532_1[0]),.doutb(w_n532_1[1]),.din(w_n532_0[0]));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.doutc(w_n551_0[2]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl3 jspl3_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.doutc(w_n556_5[2]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n556_6(.douta(w_n556_6[0]),.doutb(w_n556_6[1]),.doutc(w_n556_6[2]),.din(w_n556_1[2]));
	jspl3 jspl3_w_n556_7(.douta(w_n556_7[0]),.doutb(w_n556_7[1]),.doutc(w_n556_7[2]),.din(w_n556_2[0]));
	jspl jspl_w_n556_8(.douta(w_n556_8[0]),.doutb(w_n556_8[1]),.din(w_n556_2[1]));
	jspl jspl_w_n557_0(.douta(w_dff_A_0k8lOAaf5_0),.doutb(w_n557_0[1]),.din(n557));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_dff_A_cSQndLGD4_1),.din(n559));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n561_1(.douta(w_n561_1[0]),.doutb(w_n561_1[1]),.din(w_n561_0[0]));
	jspl jspl_w_n562_0(.douta(w_dff_A_uhsIQN6V4_0),.doutb(w_n562_0[1]),.din(n562));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_dff_A_mYwDRUot2_1),.din(n564));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n569_0(.douta(w_dff_A_6ICbiHw30_0),.doutb(w_n569_0[1]),.din(n569));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_dff_A_BEGkXa3p6_1),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_dff_A_UYNv0ANo9_0),.doutb(w_dff_A_VwBB50Uj6_1),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_dff_A_7iIMNZtS0_1),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.doutc(w_n578_0[2]),.din(n578));
	jspl jspl_w_n578_1(.douta(w_n578_1[0]),.doutb(w_n578_1[1]),.din(w_n578_0[0]));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_dff_A_7jgF267z0_1),.doutc(w_dff_A_C7zORkRV9_2),.din(n579));
	jspl jspl_w_n579_1(.douta(w_n579_1[0]),.doutb(w_dff_A_bYjMFFCb7_1),.din(w_n579_0[0]));
	jspl jspl_w_n581_0(.douta(w_dff_A_L6sGAcEm1_0),.doutb(w_n581_0[1]),.din(n581));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n586_1(.douta(w_n586_1[0]),.doutb(w_n586_1[1]),.din(w_n586_0[0]));
	jspl jspl_w_n587_0(.douta(w_n587_0[0]),.doutb(w_dff_A_cJouWD972_1),.din(n587));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_dff_A_YA6qdyAm1_2),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.doutc(w_n591_0[2]),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_dff_A_JafzU21e9_0),.doutb(w_n592_0[1]),.doutc(w_dff_A_YJMKUC0n2_2),.din(n592));
	jspl3 jspl3_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl jspl_w_n596_1(.douta(w_n596_1[0]),.doutb(w_n596_1[1]),.din(w_n596_0[0]));
	jspl3 jspl3_w_n597_0(.douta(w_dff_A_EUXMbap50_0),.doutb(w_n597_0[1]),.doutc(w_n597_0[2]),.din(n597));
	jspl3 jspl3_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.doutc(w_n601_0[2]),.din(n601));
	jspl jspl_w_n601_1(.douta(w_n601_1[0]),.doutb(w_n601_1[1]),.din(w_n601_0[0]));
	jspl3 jspl3_w_n602_0(.douta(w_dff_A_hh2mcvLz5_0),.doutb(w_n602_0[1]),.doutc(w_n602_0[2]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n607_1(.douta(w_n607_1[0]),.doutb(w_n607_1[1]),.din(w_n607_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_dff_A_TDWXxzhw2_1),.doutc(w_dff_A_Tmt5fEaE8_2),.din(n608));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_dff_A_GfGyIHtP2_1),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n611_0(.douta(w_n611_0[0]),.doutb(w_dff_A_0MJbWzah7_1),.doutc(w_n611_0[2]),.din(w_dff_B_Vj7upYsK3_3));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.doutc(w_n613_1[2]),.din(w_n613_0[0]));
	jspl3 jspl3_w_n613_2(.douta(w_n613_2[0]),.doutb(w_n613_2[1]),.doutc(w_n613_2[2]),.din(w_n613_0[1]));
	jspl3 jspl3_w_n613_3(.douta(w_n613_3[0]),.doutb(w_n613_3[1]),.doutc(w_n613_3[2]),.din(w_n613_0[2]));
	jspl3 jspl3_w_n613_4(.douta(w_n613_4[0]),.doutb(w_n613_4[1]),.doutc(w_n613_4[2]),.din(w_n613_1[0]));
	jspl3 jspl3_w_n613_5(.douta(w_n613_5[0]),.doutb(w_n613_5[1]),.doutc(w_n613_5[2]),.din(w_n613_1[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_dff_A_hqzwr1cJ4_1),.doutc(w_dff_A_xWm5OZUZ6_2),.din(n618));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_dff_A_xsATXNB53_1),.doutc(w_n619_0[2]),.din(n619));
	jspl3 jspl3_w_n619_1(.douta(w_n619_1[0]),.doutb(w_n619_1[1]),.doutc(w_n619_1[2]),.din(w_n619_0[0]));
	jspl3 jspl3_w_n620_0(.douta(w_n620_0[0]),.doutb(w_dff_A_nyTJjvBJ0_1),.doutc(w_dff_A_XgKPFoq79_2),.din(n620));
	jspl jspl_w_n620_1(.douta(w_n620_1[0]),.doutb(w_dff_A_QwkIgFgX5_1),.din(w_n620_0[0]));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_dff_A_mbdOxSkR8_1),.din(n621));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_dff_A_GvO4Rd130_0),.doutb(w_dff_A_SNNFvQ9E1_1),.doutc(w_n624_0[2]),.din(w_dff_B_NvEx2L4N1_3));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_dff_A_Hpe11eud5_1),.din(n625));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl jspl_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n628_0(.douta(w_dff_A_L5VotdaR3_0),.doutb(w_n628_0[1]),.doutc(w_dff_A_NneLSLTL0_2),.din(n628));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_dff_A_8ywYSxFS9_1),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n635_1(.douta(w_dff_A_1j4RLxNY6_0),.doutb(w_n635_1[1]),.din(w_n635_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.doutc(w_n637_0[2]),.din(n637));
	jspl jspl_w_n638_0(.douta(w_n638_0[0]),.doutb(w_n638_0[1]),.din(n638));
	jspl3 jspl3_w_n639_0(.douta(w_dff_A_GGPnnmZ95_0),.doutb(w_n639_0[1]),.doutc(w_n639_0[2]),.din(n639));
	jspl jspl_w_n640_0(.douta(w_dff_A_9EDswMRN3_0),.doutb(w_n640_0[1]),.din(n640));
	jspl3 jspl3_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.doutc(w_dff_A_9PX4pKkY6_2),.din(n641));
	jspl3 jspl3_w_n641_1(.douta(w_n641_1[0]),.doutb(w_n641_1[1]),.doutc(w_n641_1[2]),.din(w_n641_0[0]));
	jspl3 jspl3_w_n644_0(.douta(w_dff_A_Sc2SMKNB7_0),.doutb(w_n644_0[1]),.doutc(w_dff_A_BFxkYivm6_2),.din(n644));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_dff_A_2q2vU2484_1),.doutc(w_dff_A_q27zPIaQ0_2),.din(n648));
	jspl jspl_w_n648_1(.douta(w_n648_1[0]),.doutb(w_n648_1[1]),.din(w_n648_0[0]));
	jspl jspl_w_n649_0(.douta(w_dff_A_Jw1AnA3z8_0),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n653_0(.douta(w_dff_A_xK9GoD8d5_0),.doutb(w_n653_0[1]),.doutc(w_n653_0[2]),.din(n653));
	jspl3 jspl3_w_n654_0(.douta(w_dff_A_jDb5vWbQ6_0),.doutb(w_n654_0[1]),.doutc(w_n654_0[2]),.din(w_dff_B_5zQTNqNL4_3));
	jspl3 jspl3_w_n654_1(.douta(w_n654_1[0]),.doutb(w_dff_A_5GJOdGyi0_1),.doutc(w_n654_1[2]),.din(w_n654_0[0]));
	jspl3 jspl3_w_n654_2(.douta(w_dff_A_IxvVKXhq0_0),.doutb(w_n654_2[1]),.doutc(w_n654_2[2]),.din(w_n654_0[1]));
	jspl3 jspl3_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.doutc(w_n658_0[2]),.din(n658));
	jspl jspl_w_n658_1(.douta(w_n658_1[0]),.doutb(w_n658_1[1]),.din(w_n658_0[0]));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_dff_A_TEyNCykl0_2),.din(n660));
	jspl jspl_w_n660_1(.douta(w_dff_A_BGwoNCKI6_0),.doutb(w_n660_1[1]),.din(w_n660_0[0]));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(w_dff_B_WK3ML1VB5_2));
	jspl jspl_w_n670_0(.douta(w_n670_0[0]),.doutb(w_n670_0[1]),.din(n670));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl3 jspl3_w_n682_0(.douta(w_n682_0[0]),.doutb(w_dff_A_UqjqprCo5_1),.doutc(w_dff_A_SF6wwOlN4_2),.din(n682));
	jspl jspl_w_n684_0(.douta(w_dff_A_ugD9qJRX6_0),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_dff_A_iM2l6I6p5_0),.doutb(w_n685_0[1]),.din(w_dff_B_AW8r6ZLe9_2));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_dff_A_afZGM9lt3_1),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_dff_A_JglAYIaa8_1),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_dff_A_H1PaAqjw8_0),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n692_0(.douta(w_dff_A_A2GZ60vW9_0),.doutb(w_n692_0[1]),.din(n692));
	jspl3 jspl3_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.doutc(w_n694_0[2]),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_dff_A_Mo0cBftB0_0),.doutb(w_dff_A_GzWpiUJQ3_1),.doutc(w_n695_0[2]),.din(n695));
	jspl3 jspl3_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.doutc(w_n699_0[2]),.din(n699));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_dff_A_YX2jxMvL1_1),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_dff_A_4qAEFu3Q1_1),.din(n709));
	jspl jspl_w_n710_0(.douta(w_dff_A_x46xDeyz9_0),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_dff_A_rsjm53rT8_0),.doutb(w_n711_0[1]),.din(n711));
	jspl3 jspl3_w_n713_0(.douta(w_n713_0[0]),.doutb(w_dff_A_OkWM4bmB6_1),.doutc(w_n713_0[2]),.din(n713));
	jspl3 jspl3_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.doutc(w_n715_0[2]),.din(n715));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(w_dff_B_TlLd4l4R7_2));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_dff_A_lGvYCjGC7_1),.din(n719));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_dff_A_t6E3SN1s2_1),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_dff_A_tDgj3zKQ2_1),.din(n721));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_dff_A_ldf0b7vZ9_1),.din(n722));
	jspl3 jspl3_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.doutc(w_n725_0[2]),.din(n725));
	jspl jspl_w_n726_0(.douta(w_dff_A_Lpp4XiX75_0),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.doutc(w_n733_0[2]),.din(n733));
	jspl3 jspl3_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.doutc(w_n735_0[2]),.din(n735));
	jspl3 jspl3_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl jspl_w_n737_1(.douta(w_n737_1[0]),.doutb(w_n737_1[1]),.din(w_n737_0[0]));
	jspl jspl_w_n738_0(.douta(w_n738_0[0]),.doutb(w_n738_0[1]),.din(n738));
	jspl3 jspl3_w_n742_0(.douta(w_n742_0[0]),.doutb(w_dff_A_hbkPjEYw5_1),.doutc(w_n742_0[2]),.din(n742));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_dff_A_h8rFwdzc6_1),.doutc(w_n746_0[2]),.din(n746));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(w_dff_B_aNbiEs9k0_2));
	jspl3 jspl3_w_n749_0(.douta(w_n749_0[0]),.doutb(w_dff_A_P7w9oMCp7_1),.doutc(w_dff_A_rpIbK18c5_2),.din(n749));
	jspl3 jspl3_w_n749_1(.douta(w_n749_1[0]),.doutb(w_dff_A_gBzpWDv81_1),.doutc(w_dff_A_hfKCLmh88_2),.din(w_n749_0[0]));
	jspl3 jspl3_w_n749_2(.douta(w_dff_A_ILvPx3Bw2_0),.doutb(w_dff_A_ylr9DSxj3_1),.doutc(w_n749_2[2]),.din(w_n749_0[1]));
	jspl3 jspl3_w_n749_3(.douta(w_dff_A_UPMtDmzk0_0),.doutb(w_n749_3[1]),.doutc(w_dff_A_NexaASTY3_2),.din(w_n749_0[2]));
	jspl3 jspl3_w_n749_4(.douta(w_n749_4[0]),.doutb(w_dff_A_18S8GhZa8_1),.doutc(w_dff_A_JmgRWSyj3_2),.din(w_n749_1[0]));
	jspl3 jspl3_w_n749_5(.douta(w_dff_A_QST1B0gp0_0),.doutb(w_dff_A_KAFfH4199_1),.doutc(w_n749_5[2]),.din(w_n749_1[1]));
	jspl3 jspl3_w_n749_6(.douta(w_dff_A_tyqGwJg34_0),.doutb(w_n749_6[1]),.doutc(w_n749_6[2]),.din(w_n749_1[2]));
	jspl3 jspl3_w_n749_7(.douta(w_dff_A_HZuQsZKv6_0),.doutb(w_n749_7[1]),.doutc(w_n749_7[2]),.din(w_n749_2[0]));
	jspl3 jspl3_w_n749_8(.douta(w_n749_8[0]),.doutb(w_dff_A_mE7r4Qpk6_1),.doutc(w_dff_A_uj6YHgjT6_2),.din(w_n749_2[1]));
	jspl3 jspl3_w_n749_9(.douta(w_dff_A_6uXU1W2I7_0),.doutb(w_n749_9[1]),.doutc(w_dff_A_9Sq3Quiw6_2),.din(w_n749_2[2]));
	jspl3 jspl3_w_n749_10(.douta(w_n749_10[0]),.doutb(w_n749_10[1]),.doutc(w_n749_10[2]),.din(w_n749_3[0]));
	jspl3 jspl3_w_n749_11(.douta(w_dff_A_09RYPLEY5_0),.doutb(w_dff_A_NVDs0d1O7_1),.doutc(w_n749_11[2]),.din(w_n749_3[1]));
	jspl3 jspl3_w_n749_12(.douta(w_n749_12[0]),.doutb(w_n749_12[1]),.doutc(w_n749_12[2]),.din(w_n749_3[2]));
	jspl jspl_w_n749_13(.douta(w_dff_A_UPfevPH08_0),.doutb(w_n749_13[1]),.din(w_n749_4[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.doutc(w_n750_0[2]),.din(n750));
	jspl3 jspl3_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.doutc(w_n750_1[2]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n750_2(.douta(w_n750_2[0]),.doutb(w_n750_2[1]),.doutc(w_n750_2[2]),.din(w_n750_0[1]));
	jspl3 jspl3_w_n750_3(.douta(w_n750_3[0]),.doutb(w_n750_3[1]),.doutc(w_n750_3[2]),.din(w_n750_0[2]));
	jspl3 jspl3_w_n750_4(.douta(w_n750_4[0]),.doutb(w_n750_4[1]),.doutc(w_n750_4[2]),.din(w_n750_1[0]));
	jspl3 jspl3_w_n750_5(.douta(w_n750_5[0]),.doutb(w_n750_5[1]),.doutc(w_n750_5[2]),.din(w_n750_1[1]));
	jspl3 jspl3_w_n750_6(.douta(w_n750_6[0]),.doutb(w_n750_6[1]),.doutc(w_n750_6[2]),.din(w_n750_1[2]));
	jspl3 jspl3_w_n750_7(.douta(w_n750_7[0]),.doutb(w_n750_7[1]),.doutc(w_n750_7[2]),.din(w_n750_2[0]));
	jspl3 jspl3_w_n750_8(.douta(w_n750_8[0]),.doutb(w_n750_8[1]),.doutc(w_n750_8[2]),.din(w_n750_2[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_dff_A_DaXJgAHl0_1),.doutc(w_dff_A_v65CWJYg0_2),.din(w_dff_B_eHIEZXIz1_3));
	jspl jspl_w_n753_1(.douta(w_dff_A_l8pysX0x7_0),.doutb(w_n753_1[1]),.din(w_n753_0[0]));
	jspl jspl_w_n755_0(.douta(w_dff_A_3vp1aYyX1_0),.doutb(w_n755_0[1]),.din(n755));
	jspl3 jspl3_w_n763_0(.douta(w_dff_A_7vTZhl8j5_0),.doutb(w_n763_0[1]),.doutc(w_n763_0[2]),.din(n763));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(n767));
	jspl jspl_w_n779_0(.douta(w_dff_A_2mTScvy55_0),.doutb(w_n779_0[1]),.din(n779));
	jspl3 jspl3_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.doutc(w_n786_0[2]),.din(n786));
	jspl3 jspl3_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.doutc(w_n788_0[2]),.din(n788));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_dff_A_5Cx11GKH9_1),.doutc(w_n790_0[2]),.din(n790));
	jspl3 jspl3_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.doutc(w_dff_A_eBOdeqzC9_2),.din(n792));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_n797_1[1]),.doutc(w_n797_1[2]),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_n797_2[2]),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_dff_A_qnlRfEJH3_0),.doutb(w_n797_3[1]),.doutc(w_n797_3[2]),.din(w_n797_0[2]));
	jspl3 jspl3_w_n797_4(.douta(w_dff_A_Kyd6tigJ2_0),.doutb(w_n797_4[1]),.doutc(w_dff_A_MKO4dv4O9_2),.din(w_n797_1[0]));
	jspl3 jspl3_w_n797_5(.douta(w_n797_5[0]),.doutb(w_dff_A_ziN8tUle8_1),.doutc(w_n797_5[2]),.din(w_n797_1[1]));
	jspl3 jspl3_w_n797_6(.douta(w_dff_A_M62Dgl556_0),.doutb(w_n797_6[1]),.doutc(w_dff_A_I7AK9l4r1_2),.din(w_n797_1[2]));
	jspl3 jspl3_w_n797_7(.douta(w_n797_7[0]),.doutb(w_dff_A_EdaKIGxL6_1),.doutc(w_n797_7[2]),.din(w_n797_2[0]));
	jspl3 jspl3_w_n797_8(.douta(w_dff_A_2nbBza6c2_0),.doutb(w_n797_8[1]),.doutc(w_dff_A_IzK3vsdV9_2),.din(w_n797_2[1]));
	jspl jspl_w_n797_9(.douta(w_n797_9[0]),.doutb(w_dff_A_mEwAEQZs7_1),.din(w_n797_2[2]));
	jspl3 jspl3_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.doutc(w_n798_0[2]),.din(n798));
	jspl jspl_w_n798_1(.douta(w_n798_1[0]),.doutb(w_n798_1[1]),.din(w_n798_0[0]));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_dff_A_ZWMvM8Jk9_1),.doutc(w_dff_A_S6rN69Ok5_2),.din(w_dff_B_MwUyoqxu1_3));
	jspl3 jspl3_w_n800_1(.douta(w_n800_1[0]),.doutb(w_dff_A_uDMLZepB0_1),.doutc(w_dff_A_BpvSD57Q4_2),.din(w_n800_0[0]));
	jspl3 jspl3_w_n800_2(.douta(w_n800_2[0]),.doutb(w_n800_2[1]),.doutc(w_dff_A_AEZVYED01_2),.din(w_n800_0[1]));
	jspl3 jspl3_w_n800_3(.douta(w_dff_A_dHQr3Ovf9_0),.doutb(w_n800_3[1]),.doutc(w_dff_A_1ZfHs2xD5_2),.din(w_n800_0[2]));
	jspl jspl_w_n800_4(.douta(w_dff_A_HaikhZZP3_0),.doutb(w_n800_4[1]),.din(w_n800_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl jspl_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n814_0(.douta(w_dff_A_Ox40Ompz4_0),.doutb(w_dff_A_eJs5oGEJ3_1),.doutc(w_n814_0[2]),.din(n814));
	jspl3 jspl3_w_n819_0(.douta(w_n819_0[0]),.doutb(w_dff_A_ECOYXRRD5_1),.doutc(w_n819_0[2]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_dff_A_GKaXrJW94_1),.din(n821));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n836_0(.douta(w_dff_A_XA3HZLVg6_0),.doutb(w_n836_0[1]),.din(n836));
	jspl jspl_w_n847_0(.douta(w_dff_A_SJ5wKky19_0),.doutb(w_n847_0[1]),.din(n847));
	jspl3 jspl3_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.doutc(w_n852_0[2]),.din(n852));
	jspl3 jspl3_w_n852_1(.douta(w_n852_1[0]),.doutb(w_n852_1[1]),.doutc(w_n852_1[2]),.din(w_n852_0[0]));
	jspl3 jspl3_w_n852_2(.douta(w_n852_2[0]),.doutb(w_n852_2[1]),.doutc(w_n852_2[2]),.din(w_n852_0[1]));
	jspl3 jspl3_w_n852_3(.douta(w_dff_A_ViaIf9gQ0_0),.doutb(w_n852_3[1]),.doutc(w_n852_3[2]),.din(w_n852_0[2]));
	jspl3 jspl3_w_n852_4(.douta(w_dff_A_ProXiB0p1_0),.doutb(w_n852_4[1]),.doutc(w_dff_A_w2NP7IaK8_2),.din(w_n852_1[0]));
	jspl3 jspl3_w_n852_5(.douta(w_n852_5[0]),.doutb(w_dff_A_4xcqPKm27_1),.doutc(w_dff_A_tRYBKt5n9_2),.din(w_n852_1[1]));
	jspl3 jspl3_w_n852_6(.douta(w_n852_6[0]),.doutb(w_n852_6[1]),.doutc(w_dff_A_lWXD2SPz5_2),.din(w_n852_1[2]));
	jspl3 jspl3_w_n852_7(.douta(w_dff_A_8iaWdJjL1_0),.doutb(w_n852_7[1]),.doutc(w_dff_A_wEMJAAj20_2),.din(w_n852_2[0]));
	jspl3 jspl3_w_n852_8(.douta(w_n852_8[0]),.doutb(w_dff_A_hSbRJQCb8_1),.doutc(w_n852_8[2]),.din(w_n852_2[1]));
	jspl jspl_w_n852_9(.douta(w_n852_9[0]),.doutb(w_dff_A_CnFrIYZc7_1),.din(w_n852_2[2]));
	jspl3 jspl3_w_n854_0(.douta(w_n854_0[0]),.doutb(w_dff_A_Jnct4fnW9_1),.doutc(w_dff_A_yKkjTM6S1_2),.din(w_dff_B_d5G7vJYJ1_3));
	jspl3 jspl3_w_n854_1(.douta(w_n854_1[0]),.doutb(w_dff_A_tYiNUfGA0_1),.doutc(w_dff_A_jY9b8IVo4_2),.din(w_n854_0[0]));
	jspl3 jspl3_w_n854_2(.douta(w_n854_2[0]),.doutb(w_n854_2[1]),.doutc(w_n854_2[2]),.din(w_n854_0[1]));
	jspl3 jspl3_w_n854_3(.douta(w_n854_3[0]),.doutb(w_n854_3[1]),.doutc(w_dff_A_TfsvbHxf8_2),.din(w_n854_0[2]));
	jspl jspl_w_n854_4(.douta(w_dff_A_F5luKNX98_0),.doutb(w_n854_4[1]),.din(w_n854_1[0]));
	jspl3 jspl3_w_n865_0(.douta(w_dff_A_rKYk0v846_0),.doutb(w_n865_0[1]),.doutc(w_dff_A_K2zayzws2_2),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n868_0(.douta(w_n868_0[0]),.doutb(w_n868_0[1]),.din(n868));
	jspl jspl_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.din(n870));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl jspl_w_n880_0(.douta(w_dff_A_cxXdvzs87_0),.doutb(w_n880_0[1]),.din(n880));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(n890));
	jspl jspl_w_n901_0(.douta(w_dff_A_a2QCXQJn3_0),.doutb(w_n901_0[1]),.din(n901));
	jspl3 jspl3_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.doutc(w_n923_0[2]),.din(n923));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl3 jspl3_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.doutc(w_dff_A_Y4IRGbEd4_2),.din(n938));
	jspl3 jspl3_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.doutc(w_n940_0[2]),.din(n940));
	jspl jspl_w_n940_1(.douta(w_n940_1[0]),.doutb(w_n940_1[1]),.din(w_n940_0[0]));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(n944));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_dff_A_bR7YuVXX4_1),.din(n949));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl3 jspl3_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.doutc(w_dff_A_ZuWMt4rq6_2),.din(n954));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_dff_A_w7y9CaQb5_1),.din(w_dff_B_ePa9ZGLr2_2));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl3 jspl3_w_n977_0(.douta(w_n977_0[0]),.doutb(w_n977_0[1]),.doutc(w_n977_0[2]),.din(n977));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_dff_A_cgmkJVQL6_1),.din(n989));
	jspl3 jspl3_w_n993_0(.douta(w_n993_0[0]),.doutb(w_dff_A_NMehygOp9_1),.doutc(w_dff_A_olEYvere9_2),.din(n993));
	jspl3 jspl3_w_n993_1(.douta(w_n993_1[0]),.doutb(w_dff_A_xn1HbwAj0_1),.doutc(w_dff_A_iBDS9ARQ2_2),.din(w_n993_0[0]));
	jspl3 jspl3_w_n993_2(.douta(w_dff_A_6ARgsfXK6_0),.doutb(w_dff_A_2dPucS1o4_1),.doutc(w_n993_2[2]),.din(w_n993_0[1]));
	jspl3 jspl3_w_n993_3(.douta(w_dff_A_VwRZDwaz7_0),.doutb(w_dff_A_CC2qWIf52_1),.doutc(w_n993_3[2]),.din(w_n993_0[2]));
	jspl3 jspl3_w_n993_4(.douta(w_dff_A_qSpU3F0Z5_0),.doutb(w_dff_A_NkslOwSe4_1),.doutc(w_n993_4[2]),.din(w_n993_1[0]));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n994_1(.douta(w_n994_1[0]),.doutb(w_n994_1[1]),.doutc(w_n994_1[2]),.din(w_n994_0[0]));
	jspl3 jspl3_w_n994_2(.douta(w_n994_2[0]),.doutb(w_n994_2[1]),.doutc(w_n994_2[2]),.din(w_n994_0[1]));
	jspl3 jspl3_w_n994_3(.douta(w_n994_3[0]),.doutb(w_n994_3[1]),.doutc(w_n994_3[2]),.din(w_n994_0[2]));
	jspl jspl_w_n994_4(.douta(w_n994_4[0]),.doutb(w_n994_4[1]),.din(w_n994_1[0]));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl3 jspl3_w_n996_1(.douta(w_n996_1[0]),.doutb(w_n996_1[1]),.doutc(w_n996_1[2]),.din(w_n996_0[0]));
	jspl3 jspl3_w_n996_2(.douta(w_n996_2[0]),.doutb(w_n996_2[1]),.doutc(w_n996_2[2]),.din(w_n996_0[1]));
	jspl3 jspl3_w_n996_3(.douta(w_n996_3[0]),.doutb(w_n996_3[1]),.doutc(w_n996_3[2]),.din(w_n996_0[2]));
	jspl jspl_w_n996_4(.douta(w_n996_4[0]),.doutb(w_n996_4[1]),.din(w_n996_1[0]));
	jspl3 jspl3_w_n999_0(.douta(w_dff_A_qYXjQuKy8_0),.doutb(w_dff_A_3J7YtBlR4_1),.doutc(w_n999_0[2]),.din(w_dff_B_gH9XOfcv5_3));
	jspl3 jspl3_w_n999_1(.douta(w_dff_A_RlKZcSQj8_0),.doutb(w_dff_A_Tli91gTS6_1),.doutc(w_n999_1[2]),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_dff_A_gNqVIcRp2_0),.doutb(w_dff_A_p5R2bQi48_1),.doutc(w_n999_2[2]),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_dff_A_eJjTXKVm4_0),.doutb(w_dff_A_se7hXFni1_1),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl3 jspl3_w_n1007_0(.douta(w_dff_A_1grDYaM51_0),.doutb(w_dff_A_DLqRDtDr1_1),.doutc(w_n1007_0[2]),.din(w_dff_B_hRGElnj35_3));
	jspl3 jspl3_w_n1007_1(.douta(w_n1007_1[0]),.doutb(w_n1007_1[1]),.doutc(w_dff_A_ympCL9KT2_2),.din(w_n1007_0[0]));
	jspl3 jspl3_w_n1007_2(.douta(w_dff_A_MkXZOu1o5_0),.doutb(w_dff_A_FInBIvAe5_1),.doutc(w_n1007_2[2]),.din(w_n1007_0[1]));
	jspl3 jspl3_w_n1007_3(.douta(w_dff_A_L20R3OvP1_0),.doutb(w_dff_A_3SCYQOmj0_1),.doutc(w_n1007_3[2]),.din(w_n1007_0[2]));
	jspl3 jspl3_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_dff_A_CjiMQbZv0_1),.doutc(w_dff_A_R5JhrLx67_2),.din(n1008));
	jspl3 jspl3_w_n1008_1(.douta(w_n1008_1[0]),.doutb(w_dff_A_6m7zhnEg7_1),.doutc(w_dff_A_qDgDVAEX0_2),.din(w_n1008_0[0]));
	jspl3 jspl3_w_n1008_2(.douta(w_dff_A_rrVAIVQh7_0),.doutb(w_dff_A_YblE7OkE0_1),.doutc(w_n1008_2[2]),.din(w_n1008_0[1]));
	jspl3 jspl3_w_n1008_3(.douta(w_dff_A_TFA1s4mL4_0),.doutb(w_dff_A_2hbXSAaW4_1),.doutc(w_n1008_3[2]),.din(w_n1008_0[2]));
	jspl3 jspl3_w_n1008_4(.douta(w_dff_A_AOPqFoq74_0),.doutb(w_n1008_4[1]),.doutc(w_dff_A_kzzigXOh3_2),.din(w_n1008_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl3 jspl3_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.doutc(w_n1012_1[2]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1012_2(.douta(w_n1012_2[0]),.doutb(w_n1012_2[1]),.doutc(w_n1012_2[2]),.din(w_n1012_0[1]));
	jspl3 jspl3_w_n1012_3(.douta(w_n1012_3[0]),.doutb(w_n1012_3[1]),.doutc(w_n1012_3[2]),.din(w_n1012_0[2]));
	jspl jspl_w_n1012_4(.douta(w_n1012_4[0]),.doutb(w_n1012_4[1]),.din(w_n1012_1[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl3 jspl3_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.doutc(w_n1014_1[2]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1014_2(.douta(w_n1014_2[0]),.doutb(w_n1014_2[1]),.doutc(w_n1014_2[2]),.din(w_n1014_0[1]));
	jspl3 jspl3_w_n1014_3(.douta(w_n1014_3[0]),.doutb(w_n1014_3[1]),.doutc(w_n1014_3[2]),.din(w_n1014_0[2]));
	jspl jspl_w_n1014_4(.douta(w_n1014_4[0]),.doutb(w_n1014_4[1]),.din(w_n1014_1[0]));
	jspl3 jspl3_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.doutc(w_n1019_0[2]),.din(n1019));
	jspl jspl_w_n1019_1(.douta(w_n1019_1[0]),.doutb(w_n1019_1[1]),.din(w_n1019_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl3 jspl3_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.doutc(w_n1043_0[2]),.din(n1043));
	jspl jspl_w_n1043_1(.douta(w_n1043_1[0]),.doutb(w_n1043_1[1]),.din(w_n1043_0[0]));
	jspl3 jspl3_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.doutc(w_n1052_0[2]),.din(n1052));
	jspl jspl_w_n1052_1(.douta(w_n1052_1[0]),.doutb(w_n1052_1[1]),.din(w_n1052_0[0]));
	jspl3 jspl3_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.doutc(w_n1054_0[2]),.din(n1054));
	jspl jspl_w_n1054_1(.douta(w_n1054_1[0]),.doutb(w_n1054_1[1]),.din(w_n1054_0[0]));
	jspl jspl_w_n1177_0(.douta(w_dff_A_ICC9pbgr6_0),.doutb(w_n1177_0[1]),.din(w_dff_B_cYBHEi6R0_2));
	jspl jspl_w_n1179_0(.douta(w_dff_A_vXobmQJ75_0),.doutb(w_n1179_0[1]),.din(n1179));
	jspl3 jspl3_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.doutc(w_n1196_0[2]),.din(n1196));
	jspl3 jspl3_w_n1196_1(.douta(w_n1196_1[0]),.doutb(w_n1196_1[1]),.doutc(w_n1196_1[2]),.din(w_n1196_0[0]));
	jspl3 jspl3_w_n1201_0(.douta(w_dff_A_4TUwTOi88_0),.doutb(w_dff_A_k4Mc6obz5_1),.doutc(w_n1201_0[2]),.din(w_dff_B_cfmT20Li7_3));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.doutc(w_n1213_0[2]),.din(n1213));
	jspl3 jspl3_w_n1213_1(.douta(w_n1213_1[0]),.doutb(w_n1213_1[1]),.doutc(w_n1213_1[2]),.din(w_n1213_0[0]));
	jspl3 jspl3_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.doutc(w_n1236_0[2]),.din(n1236));
	jspl3 jspl3_w_n1236_1(.douta(w_n1236_1[0]),.doutb(w_n1236_1[1]),.doutc(w_n1236_1[2]),.din(w_n1236_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl3 jspl3_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.doutc(w_n1251_1[2]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.doutc(w_n1279_0[2]),.din(n1279));
	jspl jspl_w_n1279_1(.douta(w_n1279_1[0]),.doutb(w_n1279_1[1]),.din(w_n1279_0[0]));
	jspl3 jspl3_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.doutc(w_n1297_0[2]),.din(n1297));
	jspl jspl_w_n1297_1(.douta(w_n1297_1[0]),.doutb(w_n1297_1[1]),.din(w_n1297_0[0]));
	jspl3 jspl3_w_n1299_0(.douta(w_n1299_0[0]),.doutb(w_n1299_0[1]),.doutc(w_n1299_0[2]),.din(n1299));
	jspl jspl_w_n1299_1(.douta(w_n1299_1[0]),.doutb(w_n1299_1[1]),.din(w_n1299_0[0]));
	jspl3 jspl3_w_n1410_0(.douta(w_dff_A_ezJhyCPW8_0),.doutb(w_n1410_0[1]),.doutc(w_n1410_0[2]),.din(n1410));
	jspl3 jspl3_w_n1412_0(.douta(w_n1412_0[0]),.doutb(w_dff_A_gNshOweR9_1),.doutc(w_dff_A_Tc8l7UPY8_2),.din(w_dff_B_t59Osa8H5_3));
	jspl jspl_w_n1416_0(.douta(w_n1416_0[0]),.doutb(w_n1416_0[1]),.din(n1416));
	jspl jspl_w_n1422_0(.douta(w_dff_A_qLkJq7Yp4_0),.doutb(w_n1422_0[1]),.din(n1422));
	jspl jspl_w_n1425_0(.douta(w_dff_A_Sed29K6s0_0),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(n1428));
	jspl jspl_w_n1429_0(.douta(w_dff_A_IjCUvMks7_0),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1451_0(.douta(w_dff_A_JILC84RG8_0),.doutb(w_n1451_0[1]),.din(n1451));
	jspl jspl_w_n1503_0(.douta(w_n1503_0[0]),.doutb(w_n1503_0[1]),.din(n1503));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1592_0(.douta(w_n1592_0[0]),.doutb(w_n1592_0[1]),.din(n1592));
	jspl jspl_w_n1593_0(.douta(w_n1593_0[0]),.doutb(w_n1593_0[1]),.din(n1593));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1599_0(.douta(w_dff_A_eMdoammx6_0),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_n1603_0[1]),.din(n1603));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl3 jspl3_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.doutc(w_n1611_0[2]),.din(n1611));
	jspl jspl_w_n1613_0(.douta(w_dff_A_sWAv6bEr5_0),.doutb(w_n1613_0[1]),.din(n1613));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(n1615));
	jspl jspl_w_n1618_0(.douta(w_dff_A_h9RHD1Wf3_0),.doutb(w_n1618_0[1]),.din(w_dff_B_D23ryYxv9_2));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(w_dff_B_PBRYjV6g2_2));
	jspl jspl_w_n1637_0(.douta(w_dff_A_kwSz5bpb4_0),.doutb(w_n1637_0[1]),.din(w_dff_B_VeZvpyRk9_2));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(n1643));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_dff_A_ljs2Hp0w4_1),.din(n1652));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl3 jspl3_w_n1674_0(.douta(w_n1674_0[0]),.doutb(w_n1674_0[1]),.doutc(w_n1674_0[2]),.din(n1674));
	jspl jspl_w_n1675_0(.douta(w_n1675_0[0]),.doutb(w_n1675_0[1]),.din(n1675));
	jspl3 jspl3_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.doutc(w_n1679_0[2]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(w_dff_B_ComM23HU8_2));
	jspl jspl_w_n1695_0(.douta(w_n1695_0[0]),.doutb(w_n1695_0[1]),.din(w_dff_B_2yHgIPs07_2));
	jspl jspl_w_n1698_0(.douta(w_n1698_0[0]),.doutb(w_n1698_0[1]),.din(w_dff_B_zUduTCUO7_2));
	jdff dff_B_zheJpM8a6_1(.din(G136),.dout(w_dff_B_zheJpM8a6_1),.clk(gclk));
	jdff dff_B_AHgrt4gg1_0(.din(G2824),.dout(w_dff_B_AHgrt4gg1_0),.clk(gclk));
	jdff dff_B_qYdKW0mJ1_1(.din(n320),.dout(w_dff_B_qYdKW0mJ1_1),.clk(gclk));
	jdff dff_B_fb4w6OY08_1(.din(n327),.dout(w_dff_B_fb4w6OY08_1),.clk(gclk));
	jdff dff_B_C8HPys6d9_2(.din(n333),.dout(w_dff_B_C8HPys6d9_2),.clk(gclk));
	jdff dff_B_bn2KitwD0_1(.din(n338),.dout(w_dff_B_bn2KitwD0_1),.clk(gclk));
	jdff dff_B_y0l8qKDv5_1(.din(n340),.dout(w_dff_B_y0l8qKDv5_1),.clk(gclk));
	jdff dff_B_rt3JmqTJ3_0(.din(n341),.dout(w_dff_B_rt3JmqTJ3_0),.clk(gclk));
	jdff dff_B_yhLpS0385_1(.din(G24),.dout(w_dff_B_yhLpS0385_1),.clk(gclk));
	jdff dff_B_6QeaS1DH6_1(.din(n345),.dout(w_dff_B_6QeaS1DH6_1),.clk(gclk));
	jdff dff_B_mF2s9CBA5_0(.din(n346),.dout(w_dff_B_mF2s9CBA5_0),.clk(gclk));
	jdff dff_B_B3mKvrRi2_1(.din(G26),.dout(w_dff_B_B3mKvrRi2_1),.clk(gclk));
	jdff dff_A_r314CZIx0_0(.dout(w_G141_2[0]),.din(w_dff_A_r314CZIx0_0),.clk(gclk));
	jdff dff_A_aWAYliXz7_0(.dout(w_dff_A_r314CZIx0_0),.din(w_dff_A_aWAYliXz7_0),.clk(gclk));
	jdff dff_A_nO7XEJJZ0_0(.dout(w_dff_A_aWAYliXz7_0),.din(w_dff_A_nO7XEJJZ0_0),.clk(gclk));
	jdff dff_A_qdReZtOb3_0(.dout(w_dff_A_nO7XEJJZ0_0),.din(w_dff_A_qdReZtOb3_0),.clk(gclk));
	jdff dff_A_EQDWtB3Z5_1(.dout(w_G141_2[1]),.din(w_dff_A_EQDWtB3Z5_1),.clk(gclk));
	jdff dff_A_7SteU1572_1(.dout(w_dff_A_EQDWtB3Z5_1),.din(w_dff_A_7SteU1572_1),.clk(gclk));
	jdff dff_A_kGSLAakd1_1(.dout(w_dff_A_7SteU1572_1),.din(w_dff_A_kGSLAakd1_1),.clk(gclk));
	jdff dff_A_ISYTkH6Z2_1(.dout(w_dff_A_kGSLAakd1_1),.din(w_dff_A_ISYTkH6Z2_1),.clk(gclk));
	jdff dff_B_p6DqrFtN8_1(.din(n350),.dout(w_dff_B_p6DqrFtN8_1),.clk(gclk));
	jdff dff_B_F9C7J14E4_0(.din(n351),.dout(w_dff_B_F9C7J14E4_0),.clk(gclk));
	jdff dff_B_R8DwcryY0_1(.din(G79),.dout(w_dff_B_R8DwcryY0_1),.clk(gclk));
	jdff dff_B_NunCSItv5_1(.din(n355),.dout(w_dff_B_NunCSItv5_1),.clk(gclk));
	jdff dff_B_uJshMeGM7_1(.din(w_dff_B_NunCSItv5_1),.dout(w_dff_B_uJshMeGM7_1),.clk(gclk));
	jdff dff_B_ujKs66H17_1(.din(G82),.dout(w_dff_B_ujKs66H17_1),.clk(gclk));
	jdff dff_A_Zx3hLzlE1_0(.dout(w_G2358_2[0]),.din(w_dff_A_Zx3hLzlE1_0),.clk(gclk));
	jdff dff_A_5ZzhKa771_1(.dout(w_G2358_2[1]),.din(w_dff_A_5ZzhKa771_1),.clk(gclk));
	jdff dff_A_418twjYf5_1(.dout(w_G141_1[1]),.din(w_dff_A_418twjYf5_1),.clk(gclk));
	jdff dff_A_gfj8NwyJ8_1(.dout(w_dff_A_418twjYf5_1),.din(w_dff_A_gfj8NwyJ8_1),.clk(gclk));
	jdff dff_A_EOYooCHi1_1(.dout(w_dff_A_gfj8NwyJ8_1),.din(w_dff_A_EOYooCHi1_1),.clk(gclk));
	jdff dff_A_97f50Gyd7_1(.dout(w_dff_A_EOYooCHi1_1),.din(w_dff_A_97f50Gyd7_1),.clk(gclk));
	jdff dff_A_YBfL4dKa4_2(.dout(w_G141_1[2]),.din(w_dff_A_YBfL4dKa4_2),.clk(gclk));
	jdff dff_A_xkvQGNFG3_2(.dout(w_dff_A_YBfL4dKa4_2),.din(w_dff_A_xkvQGNFG3_2),.clk(gclk));
	jdff dff_A_vPHTtLPc4_2(.dout(w_dff_A_xkvQGNFG3_2),.din(w_dff_A_vPHTtLPc4_2),.clk(gclk));
	jdff dff_A_2t5NEtJb8_2(.dout(w_dff_A_vPHTtLPc4_2),.din(w_dff_A_2t5NEtJb8_2),.clk(gclk));
	jdff dff_B_oCKraORR2_1(.din(n373),.dout(w_dff_B_oCKraORR2_1),.clk(gclk));
	jdff dff_B_Aw4rgnp34_2(.din(n661),.dout(w_dff_B_Aw4rgnp34_2),.clk(gclk));
	jdff dff_B_WK3ML1VB5_2(.din(w_dff_B_Aw4rgnp34_2),.dout(w_dff_B_WK3ML1VB5_2),.clk(gclk));
	jdff dff_B_8622ALns4_2(.din(n717),.dout(w_dff_B_8622ALns4_2),.clk(gclk));
	jdff dff_B_TlLd4l4R7_2(.din(w_dff_B_8622ALns4_2),.dout(w_dff_B_TlLd4l4R7_2),.clk(gclk));
	jdff dff_B_mZyTBMf28_1(.din(n705),.dout(w_dff_B_mZyTBMf28_1),.clk(gclk));
	jdff dff_B_Kt9ZlpMB8_1(.din(w_dff_B_mZyTBMf28_1),.dout(w_dff_B_Kt9ZlpMB8_1),.clk(gclk));
	jdff dff_B_OFXwU7gD7_1(.din(w_dff_B_Kt9ZlpMB8_1),.dout(w_dff_B_OFXwU7gD7_1),.clk(gclk));
	jdff dff_B_RWLZ8jjJ7_1(.din(w_dff_B_OFXwU7gD7_1),.dout(w_dff_B_RWLZ8jjJ7_1),.clk(gclk));
	jdff dff_B_yrzte8g70_1(.din(w_dff_B_RWLZ8jjJ7_1),.dout(w_dff_B_yrzte8g70_1),.clk(gclk));
	jdff dff_B_zkPt8ae05_1(.din(w_dff_B_yrzte8g70_1),.dout(w_dff_B_zkPt8ae05_1),.clk(gclk));
	jdff dff_B_GxGmzWvC4_1(.din(n706),.dout(w_dff_B_GxGmzWvC4_1),.clk(gclk));
	jdff dff_B_rxiWQAuY8_1(.din(w_dff_B_GxGmzWvC4_1),.dout(w_dff_B_rxiWQAuY8_1),.clk(gclk));
	jdff dff_B_QjFUmAcP5_1(.din(w_dff_B_rxiWQAuY8_1),.dout(w_dff_B_QjFUmAcP5_1),.clk(gclk));
	jdff dff_B_Vbora1Dg2_1(.din(w_dff_B_QjFUmAcP5_1),.dout(w_dff_B_Vbora1Dg2_1),.clk(gclk));
	jdff dff_B_8ZvMHrhM6_1(.din(w_dff_B_Vbora1Dg2_1),.dout(w_dff_B_8ZvMHrhM6_1),.clk(gclk));
	jdff dff_A_MQXPV9BM5_1(.dout(w_n611_0[1]),.din(w_dff_A_MQXPV9BM5_1),.clk(gclk));
	jdff dff_A_0MJbWzah7_1(.dout(w_dff_A_MQXPV9BM5_1),.din(w_dff_A_0MJbWzah7_1),.clk(gclk));
	jdff dff_B_Vj7upYsK3_3(.din(n611),.dout(w_dff_B_Vj7upYsK3_3),.clk(gclk));
	jdff dff_B_BnjGn0yx4_2(.din(n747),.dout(w_dff_B_BnjGn0yx4_2),.clk(gclk));
	jdff dff_B_aNbiEs9k0_2(.din(w_dff_B_BnjGn0yx4_2),.dout(w_dff_B_aNbiEs9k0_2),.clk(gclk));
	jdff dff_B_1AgEg32t4_1(.din(n739),.dout(w_dff_B_1AgEg32t4_1),.clk(gclk));
	jdff dff_B_UHgRrhal6_1(.din(w_dff_B_1AgEg32t4_1),.dout(w_dff_B_UHgRrhal6_1),.clk(gclk));
	jdff dff_A_BXfDRO4x4_0(.dout(w_n660_1[0]),.din(w_dff_A_BXfDRO4x4_0),.clk(gclk));
	jdff dff_A_EHvls1S40_0(.dout(w_dff_A_BXfDRO4x4_0),.din(w_dff_A_EHvls1S40_0),.clk(gclk));
	jdff dff_A_lsaOxW2a0_0(.dout(w_dff_A_EHvls1S40_0),.din(w_dff_A_lsaOxW2a0_0),.clk(gclk));
	jdff dff_A_tWrpcTYi4_0(.dout(w_dff_A_lsaOxW2a0_0),.din(w_dff_A_tWrpcTYi4_0),.clk(gclk));
	jdff dff_A_BGwoNCKI6_0(.dout(w_dff_A_tWrpcTYi4_0),.din(w_dff_A_BGwoNCKI6_0),.clk(gclk));
	jdff dff_B_BKFKSKfn1_0(.din(n808),.dout(w_dff_B_BKFKSKfn1_0),.clk(gclk));
	jdff dff_B_cEkFTT688_0(.din(w_dff_B_BKFKSKfn1_0),.dout(w_dff_B_cEkFTT688_0),.clk(gclk));
	jdff dff_B_3TRYXpeV8_0(.din(w_dff_B_cEkFTT688_0),.dout(w_dff_B_3TRYXpeV8_0),.clk(gclk));
	jdff dff_B_kemvdtiQ3_0(.din(w_dff_B_3TRYXpeV8_0),.dout(w_dff_B_kemvdtiQ3_0),.clk(gclk));
	jdff dff_B_747LGKLP3_0(.din(w_dff_B_kemvdtiQ3_0),.dout(w_dff_B_747LGKLP3_0),.clk(gclk));
	jdff dff_B_OJj8kJAy1_0(.din(w_dff_B_747LGKLP3_0),.dout(w_dff_B_OJj8kJAy1_0),.clk(gclk));
	jdff dff_B_SjbGrnKe5_0(.din(w_dff_B_OJj8kJAy1_0),.dout(w_dff_B_SjbGrnKe5_0),.clk(gclk));
	jdff dff_B_Rgr8YSoU1_0(.din(w_dff_B_SjbGrnKe5_0),.dout(w_dff_B_Rgr8YSoU1_0),.clk(gclk));
	jdff dff_B_olpJCSgP0_0(.din(w_dff_B_Rgr8YSoU1_0),.dout(w_dff_B_olpJCSgP0_0),.clk(gclk));
	jdff dff_B_RxKT6oOM6_0(.din(w_dff_B_olpJCSgP0_0),.dout(w_dff_B_RxKT6oOM6_0),.clk(gclk));
	jdff dff_B_mrdx43LZ1_0(.din(n803),.dout(w_dff_B_mrdx43LZ1_0),.clk(gclk));
	jdff dff_A_hSru95eO1_1(.dout(w_n797_9[1]),.din(w_dff_A_hSru95eO1_1),.clk(gclk));
	jdff dff_A_1Qrvskhk6_1(.dout(w_dff_A_hSru95eO1_1),.din(w_dff_A_1Qrvskhk6_1),.clk(gclk));
	jdff dff_A_lvNXFgN21_1(.dout(w_dff_A_1Qrvskhk6_1),.din(w_dff_A_lvNXFgN21_1),.clk(gclk));
	jdff dff_A_BoKIMQyz7_1(.dout(w_dff_A_lvNXFgN21_1),.din(w_dff_A_BoKIMQyz7_1),.clk(gclk));
	jdff dff_A_CF9HRJSa3_1(.dout(w_dff_A_BoKIMQyz7_1),.din(w_dff_A_CF9HRJSa3_1),.clk(gclk));
	jdff dff_A_rFDWPpvm6_1(.dout(w_dff_A_CF9HRJSa3_1),.din(w_dff_A_rFDWPpvm6_1),.clk(gclk));
	jdff dff_A_4fRtJ2Ld0_1(.dout(w_dff_A_rFDWPpvm6_1),.din(w_dff_A_4fRtJ2Ld0_1),.clk(gclk));
	jdff dff_A_VHKzP71n5_1(.dout(w_dff_A_4fRtJ2Ld0_1),.din(w_dff_A_VHKzP71n5_1),.clk(gclk));
	jdff dff_A_hpnhSO6P5_1(.dout(w_dff_A_VHKzP71n5_1),.din(w_dff_A_hpnhSO6P5_1),.clk(gclk));
	jdff dff_A_mEwAEQZs7_1(.dout(w_dff_A_hpnhSO6P5_1),.din(w_dff_A_mEwAEQZs7_1),.clk(gclk));
	jdff dff_B_zCBNTJbm1_0(.din(n861),.dout(w_dff_B_zCBNTJbm1_0),.clk(gclk));
	jdff dff_B_q0lgKwgL4_0(.din(w_dff_B_zCBNTJbm1_0),.dout(w_dff_B_q0lgKwgL4_0),.clk(gclk));
	jdff dff_B_tOxloe6R5_0(.din(w_dff_B_q0lgKwgL4_0),.dout(w_dff_B_tOxloe6R5_0),.clk(gclk));
	jdff dff_B_KePzRO2j6_0(.din(w_dff_B_tOxloe6R5_0),.dout(w_dff_B_KePzRO2j6_0),.clk(gclk));
	jdff dff_B_6ejKKBRn3_0(.din(w_dff_B_KePzRO2j6_0),.dout(w_dff_B_6ejKKBRn3_0),.clk(gclk));
	jdff dff_B_Ub1LOGCF4_0(.din(w_dff_B_6ejKKBRn3_0),.dout(w_dff_B_Ub1LOGCF4_0),.clk(gclk));
	jdff dff_B_87aM68wY3_0(.din(w_dff_B_Ub1LOGCF4_0),.dout(w_dff_B_87aM68wY3_0),.clk(gclk));
	jdff dff_B_oXpZxqun1_0(.din(w_dff_B_87aM68wY3_0),.dout(w_dff_B_oXpZxqun1_0),.clk(gclk));
	jdff dff_B_k1ScRTkN0_0(.din(w_dff_B_oXpZxqun1_0),.dout(w_dff_B_k1ScRTkN0_0),.clk(gclk));
	jdff dff_B_qqeTdjm71_0(.din(w_dff_B_k1ScRTkN0_0),.dout(w_dff_B_qqeTdjm71_0),.clk(gclk));
	jdff dff_B_SC9aAKpH0_2(.din(G61),.dout(w_dff_B_SC9aAKpH0_2),.clk(gclk));
	jdff dff_B_fDqSVZGS8_0(.din(n856),.dout(w_dff_B_fDqSVZGS8_0),.clk(gclk));
	jdff dff_A_PSHJIkKu0_1(.dout(w_n852_9[1]),.din(w_dff_A_PSHJIkKu0_1),.clk(gclk));
	jdff dff_A_xwnBkUym2_1(.dout(w_dff_A_PSHJIkKu0_1),.din(w_dff_A_xwnBkUym2_1),.clk(gclk));
	jdff dff_A_llIZNsjG6_1(.dout(w_dff_A_xwnBkUym2_1),.din(w_dff_A_llIZNsjG6_1),.clk(gclk));
	jdff dff_A_N6HFh5Os7_1(.dout(w_dff_A_llIZNsjG6_1),.din(w_dff_A_N6HFh5Os7_1),.clk(gclk));
	jdff dff_A_6qTt9jls3_1(.dout(w_dff_A_N6HFh5Os7_1),.din(w_dff_A_6qTt9jls3_1),.clk(gclk));
	jdff dff_A_vTdWxZHE0_1(.dout(w_dff_A_6qTt9jls3_1),.din(w_dff_A_vTdWxZHE0_1),.clk(gclk));
	jdff dff_A_ANUWJxK22_1(.dout(w_dff_A_vTdWxZHE0_1),.din(w_dff_A_ANUWJxK22_1),.clk(gclk));
	jdff dff_A_NOjQBMsE7_1(.dout(w_dff_A_ANUWJxK22_1),.din(w_dff_A_NOjQBMsE7_1),.clk(gclk));
	jdff dff_A_L6tmT5B07_1(.dout(w_dff_A_NOjQBMsE7_1),.din(w_dff_A_L6tmT5B07_1),.clk(gclk));
	jdff dff_A_CnFrIYZc7_1(.dout(w_dff_A_L6tmT5B07_1),.din(w_dff_A_CnFrIYZc7_1),.clk(gclk));
	jdff dff_B_mvtfbOKG2_0(.din(n967),.dout(w_dff_B_mvtfbOKG2_0),.clk(gclk));
	jdff dff_B_t6uc02AZ3_1(.din(n961),.dout(w_dff_B_t6uc02AZ3_1),.clk(gclk));
	jdff dff_B_E6nqMAx73_1(.din(w_dff_B_t6uc02AZ3_1),.dout(w_dff_B_E6nqMAx73_1),.clk(gclk));
	jdff dff_B_F93TvI0b1_1(.din(w_dff_B_E6nqMAx73_1),.dout(w_dff_B_F93TvI0b1_1),.clk(gclk));
	jdff dff_B_ma5VyXQF8_0(.din(n960),.dout(w_dff_B_ma5VyXQF8_0),.clk(gclk));
	jdff dff_B_mseprEIa2_1(.din(n975),.dout(w_dff_B_mseprEIa2_1),.clk(gclk));
	jdff dff_B_aCYRy2Ew9_1(.din(w_dff_B_mseprEIa2_1),.dout(w_dff_B_aCYRy2Ew9_1),.clk(gclk));
	jdff dff_B_tGoH7vJM5_1(.din(w_dff_B_aCYRy2Ew9_1),.dout(w_dff_B_tGoH7vJM5_1),.clk(gclk));
	jdff dff_B_iCfsAdeF9_1(.din(w_dff_B_tGoH7vJM5_1),.dout(w_dff_B_iCfsAdeF9_1),.clk(gclk));
	jdff dff_B_vBhC3C0o8_1(.din(w_dff_B_iCfsAdeF9_1),.dout(w_dff_B_vBhC3C0o8_1),.clk(gclk));
	jdff dff_B_a9G33OtV7_1(.din(n971),.dout(w_dff_B_a9G33OtV7_1),.clk(gclk));
	jdff dff_B_WvPKT57L9_1(.din(w_dff_B_a9G33OtV7_1),.dout(w_dff_B_WvPKT57L9_1),.clk(gclk));
	jdff dff_B_vy8eF0Ht1_1(.din(n995),.dout(w_dff_B_vy8eF0Ht1_1),.clk(gclk));
	jdff dff_B_T9BagvzE4_1(.din(w_dff_B_vy8eF0Ht1_1),.dout(w_dff_B_T9BagvzE4_1),.clk(gclk));
	jdff dff_B_LWJuJS1r0_1(.din(w_dff_B_T9BagvzE4_1),.dout(w_dff_B_LWJuJS1r0_1),.clk(gclk));
	jdff dff_B_OdbN9Vw01_1(.din(w_dff_B_LWJuJS1r0_1),.dout(w_dff_B_OdbN9Vw01_1),.clk(gclk));
	jdff dff_B_WEmpJA6T0_1(.din(w_dff_B_OdbN9Vw01_1),.dout(w_dff_B_WEmpJA6T0_1),.clk(gclk));
	jdff dff_B_ryhRjljt1_1(.din(w_dff_B_WEmpJA6T0_1),.dout(w_dff_B_ryhRjljt1_1),.clk(gclk));
	jdff dff_B_gDqMrgC01_1(.din(w_dff_B_ryhRjljt1_1),.dout(w_dff_B_gDqMrgC01_1),.clk(gclk));
	jdff dff_B_8bHPYGMg2_1(.din(w_dff_B_gDqMrgC01_1),.dout(w_dff_B_8bHPYGMg2_1),.clk(gclk));
	jdff dff_B_o6Ii1tFw3_1(.din(w_dff_B_8bHPYGMg2_1),.dout(w_dff_B_o6Ii1tFw3_1),.clk(gclk));
	jdff dff_B_uZMLw7vn2_1(.din(w_dff_B_o6Ii1tFw3_1),.dout(w_dff_B_uZMLw7vn2_1),.clk(gclk));
	jdff dff_B_F3veK4cD5_1(.din(w_dff_B_uZMLw7vn2_1),.dout(w_dff_B_F3veK4cD5_1),.clk(gclk));
	jdff dff_B_PfKdQwpT6_1(.din(n997),.dout(w_dff_B_PfKdQwpT6_1),.clk(gclk));
	jdff dff_B_GP8W2Ox08_1(.din(w_dff_B_PfKdQwpT6_1),.dout(w_dff_B_GP8W2Ox08_1),.clk(gclk));
	jdff dff_B_uTGJv7LH8_1(.din(w_dff_B_GP8W2Ox08_1),.dout(w_dff_B_uTGJv7LH8_1),.clk(gclk));
	jdff dff_B_aNc5nfHR2_1(.din(w_dff_B_uTGJv7LH8_1),.dout(w_dff_B_aNc5nfHR2_1),.clk(gclk));
	jdff dff_B_a84F3n2V2_1(.din(w_dff_B_aNc5nfHR2_1),.dout(w_dff_B_a84F3n2V2_1),.clk(gclk));
	jdff dff_B_CpMuQuO23_1(.din(w_dff_B_a84F3n2V2_1),.dout(w_dff_B_CpMuQuO23_1),.clk(gclk));
	jdff dff_B_a4g8dfkr9_1(.din(w_dff_B_CpMuQuO23_1),.dout(w_dff_B_a4g8dfkr9_1),.clk(gclk));
	jdff dff_B_gD1qHAC90_1(.din(w_dff_B_a4g8dfkr9_1),.dout(w_dff_B_gD1qHAC90_1),.clk(gclk));
	jdff dff_B_ScYqek9Z6_1(.din(w_dff_B_gD1qHAC90_1),.dout(w_dff_B_ScYqek9Z6_1),.clk(gclk));
	jdff dff_B_gTsL1HLz8_1(.din(w_dff_B_ScYqek9Z6_1),.dout(w_dff_B_gTsL1HLz8_1),.clk(gclk));
	jdff dff_B_k6SjvXSa7_1(.din(w_dff_B_gTsL1HLz8_1),.dout(w_dff_B_k6SjvXSa7_1),.clk(gclk));
	jdff dff_B_pD7lTEdd0_0(.din(n1001),.dout(w_dff_B_pD7lTEdd0_0),.clk(gclk));
	jdff dff_B_62L0GS0U4_0(.din(n1016),.dout(w_dff_B_62L0GS0U4_0),.clk(gclk));
	jdff dff_B_WldPV59z8_0(.din(w_dff_B_62L0GS0U4_0),.dout(w_dff_B_WldPV59z8_0),.clk(gclk));
	jdff dff_B_pPDT1AQ16_0(.din(w_dff_B_WldPV59z8_0),.dout(w_dff_B_pPDT1AQ16_0),.clk(gclk));
	jdff dff_B_23bCwgkB6_0(.din(w_dff_B_pPDT1AQ16_0),.dout(w_dff_B_23bCwgkB6_0),.clk(gclk));
	jdff dff_B_kfFsUcZl7_0(.din(w_dff_B_23bCwgkB6_0),.dout(w_dff_B_kfFsUcZl7_0),.clk(gclk));
	jdff dff_B_5dojtcMA0_0(.din(w_dff_B_kfFsUcZl7_0),.dout(w_dff_B_5dojtcMA0_0),.clk(gclk));
	jdff dff_B_ZaDQDCL62_0(.din(w_dff_B_5dojtcMA0_0),.dout(w_dff_B_ZaDQDCL62_0),.clk(gclk));
	jdff dff_B_qIMYH9Qa7_0(.din(w_dff_B_ZaDQDCL62_0),.dout(w_dff_B_qIMYH9Qa7_0),.clk(gclk));
	jdff dff_B_BSGKBOSb8_0(.din(w_dff_B_qIMYH9Qa7_0),.dout(w_dff_B_BSGKBOSb8_0),.clk(gclk));
	jdff dff_B_2MIFHDv32_0(.din(w_dff_B_BSGKBOSb8_0),.dout(w_dff_B_2MIFHDv32_0),.clk(gclk));
	jdff dff_B_f2GERJv18_1(.din(n1013),.dout(w_dff_B_f2GERJv18_1),.clk(gclk));
	jdff dff_B_hqcGs7799_2(.din(G182),.dout(w_dff_B_hqcGs7799_2),.clk(gclk));
	jdff dff_B_1nqnb48u7_2(.din(w_dff_B_hqcGs7799_2),.dout(w_dff_B_1nqnb48u7_2),.clk(gclk));
	jdff dff_B_FgmiDBhq7_2(.din(G185),.dout(w_dff_B_FgmiDBhq7_2),.clk(gclk));
	jdff dff_B_f4CK2JYY4_1(.din(n1006),.dout(w_dff_B_f4CK2JYY4_1),.clk(gclk));
	jdff dff_B_XW9QjEk24_1(.din(w_dff_B_f4CK2JYY4_1),.dout(w_dff_B_XW9QjEk24_1),.clk(gclk));
	jdff dff_B_VRgdXbNk2_1(.din(w_dff_B_XW9QjEk24_1),.dout(w_dff_B_VRgdXbNk2_1),.clk(gclk));
	jdff dff_B_fBgsIMRS9_1(.din(n777),.dout(w_dff_B_fBgsIMRS9_1),.clk(gclk));
	jdff dff_B_CmOPjsED1_1(.din(w_dff_B_fBgsIMRS9_1),.dout(w_dff_B_CmOPjsED1_1),.clk(gclk));
	jdff dff_B_8oO7MKjx3_1(.din(w_dff_B_CmOPjsED1_1),.dout(w_dff_B_8oO7MKjx3_1),.clk(gclk));
	jdff dff_B_FJmefle53_1(.din(w_dff_B_8oO7MKjx3_1),.dout(w_dff_B_FJmefle53_1),.clk(gclk));
	jdff dff_B_wWBhILXJ6_1(.din(w_dff_B_FJmefle53_1),.dout(w_dff_B_wWBhILXJ6_1),.clk(gclk));
	jdff dff_B_0z2OHNJy6_0(.din(n782),.dout(w_dff_B_0z2OHNJy6_0),.clk(gclk));
	jdff dff_B_G5AviPzR2_1(.din(n536),.dout(w_dff_B_G5AviPzR2_1),.clk(gclk));
	jdff dff_B_W6Ge03QS3_1(.din(n531),.dout(w_dff_B_W6Ge03QS3_1),.clk(gclk));
	jdff dff_A_pOxdtWsD6_0(.dout(w_n779_0[0]),.din(w_dff_A_pOxdtWsD6_0),.clk(gclk));
	jdff dff_A_2mTScvy55_0(.dout(w_dff_A_pOxdtWsD6_0),.din(w_dff_A_2mTScvy55_0),.clk(gclk));
	jdff dff_B_Rm3ZK2Nx8_1(.din(G117),.dout(w_dff_B_Rm3ZK2Nx8_1),.clk(gclk));
	jdff dff_B_4atA8eYM2_1(.din(w_dff_B_Rm3ZK2Nx8_1),.dout(w_dff_B_4atA8eYM2_1),.clk(gclk));
	jdff dff_B_PdZaLB6I9_1(.din(n752),.dout(w_dff_B_PdZaLB6I9_1),.clk(gclk));
	jdff dff_B_z6H0G1qN4_1(.din(w_dff_B_PdZaLB6I9_1),.dout(w_dff_B_z6H0G1qN4_1),.clk(gclk));
	jdff dff_B_MpnMFYaW1_1(.din(w_dff_B_z6H0G1qN4_1),.dout(w_dff_B_MpnMFYaW1_1),.clk(gclk));
	jdff dff_A_HyeU5No36_0(.dout(w_n755_0[0]),.din(w_dff_A_HyeU5No36_0),.clk(gclk));
	jdff dff_A_OK5Px8QS4_0(.dout(w_dff_A_HyeU5No36_0),.din(w_dff_A_OK5Px8QS4_0),.clk(gclk));
	jdff dff_A_udCIlLJj0_0(.dout(w_dff_A_OK5Px8QS4_0),.din(w_dff_A_udCIlLJj0_0),.clk(gclk));
	jdff dff_A_Nz7dAw6z6_0(.dout(w_dff_A_udCIlLJj0_0),.din(w_dff_A_Nz7dAw6z6_0),.clk(gclk));
	jdff dff_A_5MXuvVuT3_0(.dout(w_dff_A_Nz7dAw6z6_0),.din(w_dff_A_5MXuvVuT3_0),.clk(gclk));
	jdff dff_A_k0Wk6R5K6_0(.dout(w_dff_A_5MXuvVuT3_0),.din(w_dff_A_k0Wk6R5K6_0),.clk(gclk));
	jdff dff_A_uij7RR0U6_0(.dout(w_dff_A_k0Wk6R5K6_0),.din(w_dff_A_uij7RR0U6_0),.clk(gclk));
	jdff dff_A_zcM0sTcP0_0(.dout(w_dff_A_uij7RR0U6_0),.din(w_dff_A_zcM0sTcP0_0),.clk(gclk));
	jdff dff_A_b00oFZC20_0(.dout(w_dff_A_zcM0sTcP0_0),.din(w_dff_A_b00oFZC20_0),.clk(gclk));
	jdff dff_A_wOYSOi314_0(.dout(w_dff_A_b00oFZC20_0),.din(w_dff_A_wOYSOi314_0),.clk(gclk));
	jdff dff_A_3vp1aYyX1_0(.dout(w_dff_A_wOYSOi314_0),.din(w_dff_A_3vp1aYyX1_0),.clk(gclk));
	jdff dff_B_v8h3GWND4_1(.din(G131),.dout(w_dff_B_v8h3GWND4_1),.clk(gclk));
	jdff dff_B_fRNMjkG23_1(.din(w_dff_B_v8h3GWND4_1),.dout(w_dff_B_fRNMjkG23_1),.clk(gclk));
	jdff dff_B_7hi2OYhc7_0(.din(n1028),.dout(w_dff_B_7hi2OYhc7_0),.clk(gclk));
	jdff dff_B_8CL04iFQ3_0(.din(w_dff_B_7hi2OYhc7_0),.dout(w_dff_B_8CL04iFQ3_0),.clk(gclk));
	jdff dff_B_s4wS4LRY2_0(.din(w_dff_B_8CL04iFQ3_0),.dout(w_dff_B_s4wS4LRY2_0),.clk(gclk));
	jdff dff_B_dn3hLhNJ1_0(.din(w_dff_B_s4wS4LRY2_0),.dout(w_dff_B_dn3hLhNJ1_0),.clk(gclk));
	jdff dff_B_q7blMNJ18_0(.din(w_dff_B_dn3hLhNJ1_0),.dout(w_dff_B_q7blMNJ18_0),.clk(gclk));
	jdff dff_B_SblSu6v96_0(.din(w_dff_B_q7blMNJ18_0),.dout(w_dff_B_SblSu6v96_0),.clk(gclk));
	jdff dff_B_OOjWpZ8N2_0(.din(w_dff_B_SblSu6v96_0),.dout(w_dff_B_OOjWpZ8N2_0),.clk(gclk));
	jdff dff_B_e4us51jA8_0(.din(w_dff_B_OOjWpZ8N2_0),.dout(w_dff_B_e4us51jA8_0),.clk(gclk));
	jdff dff_B_bF6LpzLO7_0(.din(w_dff_B_e4us51jA8_0),.dout(w_dff_B_bF6LpzLO7_0),.clk(gclk));
	jdff dff_B_0AVJ2yW95_0(.din(w_dff_B_bF6LpzLO7_0),.dout(w_dff_B_0AVJ2yW95_0),.clk(gclk));
	jdff dff_B_xzv5ohvN7_0(.din(w_dff_B_0AVJ2yW95_0),.dout(w_dff_B_xzv5ohvN7_0),.clk(gclk));
	jdff dff_B_WMSvK1lZ5_0(.din(w_dff_B_xzv5ohvN7_0),.dout(w_dff_B_WMSvK1lZ5_0),.clk(gclk));
	jdff dff_B_c0siQ1Xo7_0(.din(w_dff_B_WMSvK1lZ5_0),.dout(w_dff_B_c0siQ1Xo7_0),.clk(gclk));
	jdff dff_B_zpsoaStt8_0(.din(w_dff_B_c0siQ1Xo7_0),.dout(w_dff_B_zpsoaStt8_0),.clk(gclk));
	jdff dff_B_wT1TZ09k6_0(.din(w_dff_B_zpsoaStt8_0),.dout(w_dff_B_wT1TZ09k6_0),.clk(gclk));
	jdff dff_B_5gqfWVpb8_0(.din(w_dff_B_wT1TZ09k6_0),.dout(w_dff_B_5gqfWVpb8_0),.clk(gclk));
	jdff dff_B_neTZGdA48_1(.din(n1020),.dout(w_dff_B_neTZGdA48_1),.clk(gclk));
	jdff dff_A_GnEUwN5J3_0(.dout(w_n800_4[0]),.din(w_dff_A_GnEUwN5J3_0),.clk(gclk));
	jdff dff_A_WrQhqWRE5_0(.dout(w_dff_A_GnEUwN5J3_0),.din(w_dff_A_WrQhqWRE5_0),.clk(gclk));
	jdff dff_A_b8VkJsUx7_0(.dout(w_dff_A_WrQhqWRE5_0),.din(w_dff_A_b8VkJsUx7_0),.clk(gclk));
	jdff dff_A_5Zmgp9vf8_0(.dout(w_dff_A_b8VkJsUx7_0),.din(w_dff_A_5Zmgp9vf8_0),.clk(gclk));
	jdff dff_A_dc2Ayljc6_0(.dout(w_dff_A_5Zmgp9vf8_0),.din(w_dff_A_dc2Ayljc6_0),.clk(gclk));
	jdff dff_A_PlB2W2G97_0(.dout(w_dff_A_dc2Ayljc6_0),.din(w_dff_A_PlB2W2G97_0),.clk(gclk));
	jdff dff_A_HaikhZZP3_0(.dout(w_dff_A_PlB2W2G97_0),.din(w_dff_A_HaikhZZP3_0),.clk(gclk));
	jdff dff_B_AB2s4cjT6_0(.din(n1039),.dout(w_dff_B_AB2s4cjT6_0),.clk(gclk));
	jdff dff_B_4V624dSC0_0(.din(w_dff_B_AB2s4cjT6_0),.dout(w_dff_B_4V624dSC0_0),.clk(gclk));
	jdff dff_B_vSHwxjNt3_0(.din(w_dff_B_4V624dSC0_0),.dout(w_dff_B_vSHwxjNt3_0),.clk(gclk));
	jdff dff_B_FrnA06350_0(.din(w_dff_B_vSHwxjNt3_0),.dout(w_dff_B_FrnA06350_0),.clk(gclk));
	jdff dff_B_gWo9ypdf2_0(.din(w_dff_B_FrnA06350_0),.dout(w_dff_B_gWo9ypdf2_0),.clk(gclk));
	jdff dff_B_J5YxlibS3_0(.din(w_dff_B_gWo9ypdf2_0),.dout(w_dff_B_J5YxlibS3_0),.clk(gclk));
	jdff dff_B_0U00ivlP3_0(.din(w_dff_B_J5YxlibS3_0),.dout(w_dff_B_0U00ivlP3_0),.clk(gclk));
	jdff dff_B_ytJmcFom0_0(.din(w_dff_B_0U00ivlP3_0),.dout(w_dff_B_ytJmcFom0_0),.clk(gclk));
	jdff dff_B_kNflGQzO7_0(.din(w_dff_B_ytJmcFom0_0),.dout(w_dff_B_kNflGQzO7_0),.clk(gclk));
	jdff dff_B_i46h3C6x0_0(.din(w_dff_B_kNflGQzO7_0),.dout(w_dff_B_i46h3C6x0_0),.clk(gclk));
	jdff dff_B_yCbYYlZM4_0(.din(w_dff_B_i46h3C6x0_0),.dout(w_dff_B_yCbYYlZM4_0),.clk(gclk));
	jdff dff_B_YYFfSKoS8_0(.din(w_dff_B_yCbYYlZM4_0),.dout(w_dff_B_YYFfSKoS8_0),.clk(gclk));
	jdff dff_B_cJNGMVyF6_0(.din(w_dff_B_YYFfSKoS8_0),.dout(w_dff_B_cJNGMVyF6_0),.clk(gclk));
	jdff dff_B_aRCPDiZZ3_0(.din(w_dff_B_cJNGMVyF6_0),.dout(w_dff_B_aRCPDiZZ3_0),.clk(gclk));
	jdff dff_B_lUb34adj1_0(.din(w_dff_B_aRCPDiZZ3_0),.dout(w_dff_B_lUb34adj1_0),.clk(gclk));
	jdff dff_B_AiJxHKK30_1(.din(n1031),.dout(w_dff_B_AiJxHKK30_1),.clk(gclk));
	jdff dff_B_Cgqz8Wrk5_1(.din(w_dff_B_AiJxHKK30_1),.dout(w_dff_B_Cgqz8Wrk5_1),.clk(gclk));
	jdff dff_A_7bUtwmem0_0(.dout(w_G4088_8[0]),.din(w_dff_A_7bUtwmem0_0),.clk(gclk));
	jdff dff_A_jRn4hofL0_0(.dout(w_dff_A_7bUtwmem0_0),.din(w_dff_A_jRn4hofL0_0),.clk(gclk));
	jdff dff_A_VHpr4vki4_0(.dout(w_dff_A_jRn4hofL0_0),.din(w_dff_A_VHpr4vki4_0),.clk(gclk));
	jdff dff_A_lnf7rF5H4_0(.dout(w_dff_A_VHpr4vki4_0),.din(w_dff_A_lnf7rF5H4_0),.clk(gclk));
	jdff dff_A_y6y09Jhf9_0(.dout(w_dff_A_lnf7rF5H4_0),.din(w_dff_A_y6y09Jhf9_0),.clk(gclk));
	jdff dff_A_alptRk5K0_0(.dout(w_dff_A_y6y09Jhf9_0),.din(w_dff_A_alptRk5K0_0),.clk(gclk));
	jdff dff_A_GXnVcBu23_0(.dout(w_dff_A_alptRk5K0_0),.din(w_dff_A_GXnVcBu23_0),.clk(gclk));
	jdff dff_A_JaYRlBjm4_0(.dout(w_dff_A_GXnVcBu23_0),.din(w_dff_A_JaYRlBjm4_0),.clk(gclk));
	jdff dff_A_ZbGSDWDX6_0(.dout(w_dff_A_JaYRlBjm4_0),.din(w_dff_A_ZbGSDWDX6_0),.clk(gclk));
	jdff dff_A_ePEtkknh1_0(.dout(w_dff_A_ZbGSDWDX6_0),.din(w_dff_A_ePEtkknh1_0),.clk(gclk));
	jdff dff_A_MrNfuHpO4_0(.dout(w_dff_A_ePEtkknh1_0),.din(w_dff_A_MrNfuHpO4_0),.clk(gclk));
	jdff dff_A_ni5jUwik3_0(.dout(w_dff_A_MrNfuHpO4_0),.din(w_dff_A_ni5jUwik3_0),.clk(gclk));
	jdff dff_A_jc1ziRt50_0(.dout(w_dff_A_ni5jUwik3_0),.din(w_dff_A_jc1ziRt50_0),.clk(gclk));
	jdff dff_A_RHImzFgB8_0(.dout(w_dff_A_jc1ziRt50_0),.din(w_dff_A_RHImzFgB8_0),.clk(gclk));
	jdff dff_A_vhDY77Uo2_0(.dout(w_dff_A_RHImzFgB8_0),.din(w_dff_A_vhDY77Uo2_0),.clk(gclk));
	jdff dff_A_uC3BmT1G3_2(.dout(w_G4088_8[2]),.din(w_dff_A_uC3BmT1G3_2),.clk(gclk));
	jdff dff_A_FRG6RNVF9_2(.dout(w_dff_A_uC3BmT1G3_2),.din(w_dff_A_FRG6RNVF9_2),.clk(gclk));
	jdff dff_A_CJZTRi2D7_2(.dout(w_dff_A_FRG6RNVF9_2),.din(w_dff_A_CJZTRi2D7_2),.clk(gclk));
	jdff dff_A_CN6zjNi78_2(.dout(w_dff_A_CJZTRi2D7_2),.din(w_dff_A_CN6zjNi78_2),.clk(gclk));
	jdff dff_A_V9B0xiSf7_2(.dout(w_dff_A_CN6zjNi78_2),.din(w_dff_A_V9B0xiSf7_2),.clk(gclk));
	jdff dff_A_ANwwNvdi7_2(.dout(w_dff_A_V9B0xiSf7_2),.din(w_dff_A_ANwwNvdi7_2),.clk(gclk));
	jdff dff_A_ymGeKsyE7_2(.dout(w_dff_A_ANwwNvdi7_2),.din(w_dff_A_ymGeKsyE7_2),.clk(gclk));
	jdff dff_A_HAG0qOwE3_2(.dout(w_dff_A_ymGeKsyE7_2),.din(w_dff_A_HAG0qOwE3_2),.clk(gclk));
	jdff dff_A_zXr0jjtr2_2(.dout(w_dff_A_HAG0qOwE3_2),.din(w_dff_A_zXr0jjtr2_2),.clk(gclk));
	jdff dff_A_Q3qG3HaV8_2(.dout(w_dff_A_zXr0jjtr2_2),.din(w_dff_A_Q3qG3HaV8_2),.clk(gclk));
	jdff dff_A_xoeEYkuv6_2(.dout(w_dff_A_Q3qG3HaV8_2),.din(w_dff_A_xoeEYkuv6_2),.clk(gclk));
	jdff dff_A_vUVoVSqV0_2(.dout(w_dff_A_xoeEYkuv6_2),.din(w_dff_A_vUVoVSqV0_2),.clk(gclk));
	jdff dff_A_zYbC1g8u3_2(.dout(w_dff_A_vUVoVSqV0_2),.din(w_dff_A_zYbC1g8u3_2),.clk(gclk));
	jdff dff_A_aeomzd4N3_2(.dout(w_dff_A_zYbC1g8u3_2),.din(w_dff_A_aeomzd4N3_2),.clk(gclk));
	jdff dff_A_v3sdImXK4_2(.dout(w_dff_A_aeomzd4N3_2),.din(w_dff_A_v3sdImXK4_2),.clk(gclk));
	jdff dff_A_DjpfCeFM4_2(.dout(w_dff_A_v3sdImXK4_2),.din(w_dff_A_DjpfCeFM4_2),.clk(gclk));
	jdff dff_A_5jc5QGIQ2_0(.dout(w_n797_8[0]),.din(w_dff_A_5jc5QGIQ2_0),.clk(gclk));
	jdff dff_A_sc1dwBSy1_0(.dout(w_dff_A_5jc5QGIQ2_0),.din(w_dff_A_sc1dwBSy1_0),.clk(gclk));
	jdff dff_A_zk37MMkW3_0(.dout(w_dff_A_sc1dwBSy1_0),.din(w_dff_A_zk37MMkW3_0),.clk(gclk));
	jdff dff_A_LaLxD0iW4_0(.dout(w_dff_A_zk37MMkW3_0),.din(w_dff_A_LaLxD0iW4_0),.clk(gclk));
	jdff dff_A_EVGMUc7m3_0(.dout(w_dff_A_LaLxD0iW4_0),.din(w_dff_A_EVGMUc7m3_0),.clk(gclk));
	jdff dff_A_9n5u9eqE3_0(.dout(w_dff_A_EVGMUc7m3_0),.din(w_dff_A_9n5u9eqE3_0),.clk(gclk));
	jdff dff_A_kyf6Pxnx1_0(.dout(w_dff_A_9n5u9eqE3_0),.din(w_dff_A_kyf6Pxnx1_0),.clk(gclk));
	jdff dff_A_4f8H9TnG9_0(.dout(w_dff_A_kyf6Pxnx1_0),.din(w_dff_A_4f8H9TnG9_0),.clk(gclk));
	jdff dff_A_ip7iEMmh2_0(.dout(w_dff_A_4f8H9TnG9_0),.din(w_dff_A_ip7iEMmh2_0),.clk(gclk));
	jdff dff_A_eV7pVUD00_0(.dout(w_dff_A_ip7iEMmh2_0),.din(w_dff_A_eV7pVUD00_0),.clk(gclk));
	jdff dff_A_3o7htMax4_0(.dout(w_dff_A_eV7pVUD00_0),.din(w_dff_A_3o7htMax4_0),.clk(gclk));
	jdff dff_A_XVBPQJOj8_0(.dout(w_dff_A_3o7htMax4_0),.din(w_dff_A_XVBPQJOj8_0),.clk(gclk));
	jdff dff_A_2nbBza6c2_0(.dout(w_dff_A_XVBPQJOj8_0),.din(w_dff_A_2nbBza6c2_0),.clk(gclk));
	jdff dff_A_If5rry6V3_2(.dout(w_n797_8[2]),.din(w_dff_A_If5rry6V3_2),.clk(gclk));
	jdff dff_A_Fg0SGsut4_2(.dout(w_dff_A_If5rry6V3_2),.din(w_dff_A_Fg0SGsut4_2),.clk(gclk));
	jdff dff_A_uCwmK0434_2(.dout(w_dff_A_Fg0SGsut4_2),.din(w_dff_A_uCwmK0434_2),.clk(gclk));
	jdff dff_A_gJwoiWJP8_2(.dout(w_dff_A_uCwmK0434_2),.din(w_dff_A_gJwoiWJP8_2),.clk(gclk));
	jdff dff_A_iEW0y4j53_2(.dout(w_dff_A_gJwoiWJP8_2),.din(w_dff_A_iEW0y4j53_2),.clk(gclk));
	jdff dff_A_eXTSK3Q03_2(.dout(w_dff_A_iEW0y4j53_2),.din(w_dff_A_eXTSK3Q03_2),.clk(gclk));
	jdff dff_A_7LDOQc7k1_2(.dout(w_dff_A_eXTSK3Q03_2),.din(w_dff_A_7LDOQc7k1_2),.clk(gclk));
	jdff dff_A_S8yWeT8N2_2(.dout(w_dff_A_7LDOQc7k1_2),.din(w_dff_A_S8yWeT8N2_2),.clk(gclk));
	jdff dff_A_1CcmG2343_2(.dout(w_dff_A_S8yWeT8N2_2),.din(w_dff_A_1CcmG2343_2),.clk(gclk));
	jdff dff_A_oncGayq52_2(.dout(w_dff_A_1CcmG2343_2),.din(w_dff_A_oncGayq52_2),.clk(gclk));
	jdff dff_A_ZYEJExNN1_2(.dout(w_dff_A_oncGayq52_2),.din(w_dff_A_ZYEJExNN1_2),.clk(gclk));
	jdff dff_A_7JOIGxhs2_2(.dout(w_dff_A_ZYEJExNN1_2),.din(w_dff_A_7JOIGxhs2_2),.clk(gclk));
	jdff dff_A_JYf4Vl1q7_2(.dout(w_dff_A_7JOIGxhs2_2),.din(w_dff_A_JYf4Vl1q7_2),.clk(gclk));
	jdff dff_A_JzxeJp815_2(.dout(w_dff_A_JYf4Vl1q7_2),.din(w_dff_A_JzxeJp815_2),.clk(gclk));
	jdff dff_A_IzK3vsdV9_2(.dout(w_dff_A_JzxeJp815_2),.din(w_dff_A_IzK3vsdV9_2),.clk(gclk));
	jdff dff_B_6Bdj4B4U4_0(.din(n1050),.dout(w_dff_B_6Bdj4B4U4_0),.clk(gclk));
	jdff dff_B_O4dZeWzu8_0(.din(w_dff_B_6Bdj4B4U4_0),.dout(w_dff_B_O4dZeWzu8_0),.clk(gclk));
	jdff dff_B_XdLfVSZa3_0(.din(w_dff_B_O4dZeWzu8_0),.dout(w_dff_B_XdLfVSZa3_0),.clk(gclk));
	jdff dff_B_AGuYI6W31_0(.din(w_dff_B_XdLfVSZa3_0),.dout(w_dff_B_AGuYI6W31_0),.clk(gclk));
	jdff dff_B_JRyez78m4_0(.din(w_dff_B_AGuYI6W31_0),.dout(w_dff_B_JRyez78m4_0),.clk(gclk));
	jdff dff_B_YWsugIs99_0(.din(w_dff_B_JRyez78m4_0),.dout(w_dff_B_YWsugIs99_0),.clk(gclk));
	jdff dff_B_LeXiBPKp7_0(.din(w_dff_B_YWsugIs99_0),.dout(w_dff_B_LeXiBPKp7_0),.clk(gclk));
	jdff dff_B_sWUguajH4_0(.din(w_dff_B_LeXiBPKp7_0),.dout(w_dff_B_sWUguajH4_0),.clk(gclk));
	jdff dff_B_1WYIyQsI4_0(.din(w_dff_B_sWUguajH4_0),.dout(w_dff_B_1WYIyQsI4_0),.clk(gclk));
	jdff dff_B_jfIJiS205_0(.din(w_dff_B_1WYIyQsI4_0),.dout(w_dff_B_jfIJiS205_0),.clk(gclk));
	jdff dff_B_54iNMhB09_0(.din(w_dff_B_jfIJiS205_0),.dout(w_dff_B_54iNMhB09_0),.clk(gclk));
	jdff dff_B_KABlnsFX8_0(.din(w_dff_B_54iNMhB09_0),.dout(w_dff_B_KABlnsFX8_0),.clk(gclk));
	jdff dff_B_vv8Jq0650_0(.din(w_dff_B_KABlnsFX8_0),.dout(w_dff_B_vv8Jq0650_0),.clk(gclk));
	jdff dff_B_1CWlwn4L5_1(.din(n1042),.dout(w_dff_B_1CWlwn4L5_1),.clk(gclk));
	jdff dff_A_61z1j6fq9_1(.dout(w_n797_7[1]),.din(w_dff_A_61z1j6fq9_1),.clk(gclk));
	jdff dff_A_j6YpSyXi4_1(.dout(w_dff_A_61z1j6fq9_1),.din(w_dff_A_j6YpSyXi4_1),.clk(gclk));
	jdff dff_A_cRjUyetP3_1(.dout(w_dff_A_j6YpSyXi4_1),.din(w_dff_A_cRjUyetP3_1),.clk(gclk));
	jdff dff_A_1W3Ck1436_1(.dout(w_dff_A_cRjUyetP3_1),.din(w_dff_A_1W3Ck1436_1),.clk(gclk));
	jdff dff_A_qx2BPPnp8_1(.dout(w_dff_A_1W3Ck1436_1),.din(w_dff_A_qx2BPPnp8_1),.clk(gclk));
	jdff dff_A_cjUmcXkp1_1(.dout(w_dff_A_qx2BPPnp8_1),.din(w_dff_A_cjUmcXkp1_1),.clk(gclk));
	jdff dff_A_UhE6Z2CL7_1(.dout(w_dff_A_cjUmcXkp1_1),.din(w_dff_A_UhE6Z2CL7_1),.clk(gclk));
	jdff dff_A_BX5AsIJI4_1(.dout(w_dff_A_UhE6Z2CL7_1),.din(w_dff_A_BX5AsIJI4_1),.clk(gclk));
	jdff dff_A_viNjIyen4_1(.dout(w_dff_A_BX5AsIJI4_1),.din(w_dff_A_viNjIyen4_1),.clk(gclk));
	jdff dff_A_7DejEo559_1(.dout(w_dff_A_viNjIyen4_1),.din(w_dff_A_7DejEo559_1),.clk(gclk));
	jdff dff_A_jxrR6EKm0_1(.dout(w_dff_A_7DejEo559_1),.din(w_dff_A_jxrR6EKm0_1),.clk(gclk));
	jdff dff_A_EdaKIGxL6_1(.dout(w_dff_A_jxrR6EKm0_1),.din(w_dff_A_EdaKIGxL6_1),.clk(gclk));
	jdff dff_A_tjxL3j0M0_1(.dout(w_G4088_7[1]),.din(w_dff_A_tjxL3j0M0_1),.clk(gclk));
	jdff dff_A_2dQI5PSU5_1(.dout(w_dff_A_tjxL3j0M0_1),.din(w_dff_A_2dQI5PSU5_1),.clk(gclk));
	jdff dff_A_pn99vB4U9_1(.dout(w_dff_A_2dQI5PSU5_1),.din(w_dff_A_pn99vB4U9_1),.clk(gclk));
	jdff dff_A_fPSn3NTK8_1(.dout(w_dff_A_pn99vB4U9_1),.din(w_dff_A_fPSn3NTK8_1),.clk(gclk));
	jdff dff_A_hDK65s6C0_1(.dout(w_dff_A_fPSn3NTK8_1),.din(w_dff_A_hDK65s6C0_1),.clk(gclk));
	jdff dff_A_w5738VEI4_1(.dout(w_dff_A_hDK65s6C0_1),.din(w_dff_A_w5738VEI4_1),.clk(gclk));
	jdff dff_A_iucM0O0N7_1(.dout(w_dff_A_w5738VEI4_1),.din(w_dff_A_iucM0O0N7_1),.clk(gclk));
	jdff dff_A_yTmAVrjS3_1(.dout(w_dff_A_iucM0O0N7_1),.din(w_dff_A_yTmAVrjS3_1),.clk(gclk));
	jdff dff_A_Ct4zHAir9_1(.dout(w_dff_A_yTmAVrjS3_1),.din(w_dff_A_Ct4zHAir9_1),.clk(gclk));
	jdff dff_A_Pjsmd1b37_1(.dout(w_dff_A_Ct4zHAir9_1),.din(w_dff_A_Pjsmd1b37_1),.clk(gclk));
	jdff dff_A_2Q8jkmHO1_1(.dout(w_dff_A_Pjsmd1b37_1),.din(w_dff_A_2Q8jkmHO1_1),.clk(gclk));
	jdff dff_A_wSVjyqq36_1(.dout(w_dff_A_2Q8jkmHO1_1),.din(w_dff_A_wSVjyqq36_1),.clk(gclk));
	jdff dff_A_NO74DbYq5_1(.dout(w_dff_A_wSVjyqq36_1),.din(w_dff_A_NO74DbYq5_1),.clk(gclk));
	jdff dff_B_3RD362Ma7_0(.din(n1061),.dout(w_dff_B_3RD362Ma7_0),.clk(gclk));
	jdff dff_B_ABqfpzg69_0(.din(w_dff_B_3RD362Ma7_0),.dout(w_dff_B_ABqfpzg69_0),.clk(gclk));
	jdff dff_B_UXtPxzaz2_0(.din(w_dff_B_ABqfpzg69_0),.dout(w_dff_B_UXtPxzaz2_0),.clk(gclk));
	jdff dff_B_mcjsLtE48_0(.din(w_dff_B_UXtPxzaz2_0),.dout(w_dff_B_mcjsLtE48_0),.clk(gclk));
	jdff dff_B_LeYyvyyl1_0(.din(w_dff_B_mcjsLtE48_0),.dout(w_dff_B_LeYyvyyl1_0),.clk(gclk));
	jdff dff_B_yHPxfBZP8_0(.din(w_dff_B_LeYyvyyl1_0),.dout(w_dff_B_yHPxfBZP8_0),.clk(gclk));
	jdff dff_B_v9F355C89_0(.din(w_dff_B_yHPxfBZP8_0),.dout(w_dff_B_v9F355C89_0),.clk(gclk));
	jdff dff_B_cA8qxjrA3_0(.din(w_dff_B_v9F355C89_0),.dout(w_dff_B_cA8qxjrA3_0),.clk(gclk));
	jdff dff_B_1EiByaox8_0(.din(w_dff_B_cA8qxjrA3_0),.dout(w_dff_B_1EiByaox8_0),.clk(gclk));
	jdff dff_B_UpPZtJjT7_0(.din(w_dff_B_1EiByaox8_0),.dout(w_dff_B_UpPZtJjT7_0),.clk(gclk));
	jdff dff_B_vMRXBdSu0_0(.din(w_dff_B_UpPZtJjT7_0),.dout(w_dff_B_vMRXBdSu0_0),.clk(gclk));
	jdff dff_B_6y5qsEFA3_0(.din(w_dff_B_vMRXBdSu0_0),.dout(w_dff_B_6y5qsEFA3_0),.clk(gclk));
	jdff dff_B_Yz3a1iCD0_0(.din(w_dff_B_6y5qsEFA3_0),.dout(w_dff_B_Yz3a1iCD0_0),.clk(gclk));
	jdff dff_B_lGrJQWgO6_0(.din(w_dff_B_Yz3a1iCD0_0),.dout(w_dff_B_lGrJQWgO6_0),.clk(gclk));
	jdff dff_B_gGOmb6Bm4_1(.din(n1053),.dout(w_dff_B_gGOmb6Bm4_1),.clk(gclk));
	jdff dff_B_9mRNvP8I7_1(.din(w_dff_B_gGOmb6Bm4_1),.dout(w_dff_B_9mRNvP8I7_1),.clk(gclk));
	jdff dff_B_CFdtmdKf5_1(.din(w_dff_B_9mRNvP8I7_1),.dout(w_dff_B_CFdtmdKf5_1),.clk(gclk));
	jdff dff_A_dHQr3Ovf9_0(.dout(w_n800_3[0]),.din(w_dff_A_dHQr3Ovf9_0),.clk(gclk));
	jdff dff_A_1zfdfJ0M9_2(.dout(w_n800_3[2]),.din(w_dff_A_1zfdfJ0M9_2),.clk(gclk));
	jdff dff_A_1ZfHs2xD5_2(.dout(w_dff_A_1zfdfJ0M9_2),.din(w_dff_A_1ZfHs2xD5_2),.clk(gclk));
	jdff dff_B_eH5w5cXP7_1(.din(n1066),.dout(w_dff_B_eH5w5cXP7_1),.clk(gclk));
	jdff dff_B_kXMGvePy1_1(.din(w_dff_B_eH5w5cXP7_1),.dout(w_dff_B_kXMGvePy1_1),.clk(gclk));
	jdff dff_B_fo2TNkQC5_1(.din(w_dff_B_kXMGvePy1_1),.dout(w_dff_B_fo2TNkQC5_1),.clk(gclk));
	jdff dff_B_gKidYRAM0_1(.din(w_dff_B_fo2TNkQC5_1),.dout(w_dff_B_gKidYRAM0_1),.clk(gclk));
	jdff dff_B_MJJtl3TZ6_1(.din(w_dff_B_gKidYRAM0_1),.dout(w_dff_B_MJJtl3TZ6_1),.clk(gclk));
	jdff dff_B_PGQTR6aG6_1(.din(w_dff_B_MJJtl3TZ6_1),.dout(w_dff_B_PGQTR6aG6_1),.clk(gclk));
	jdff dff_B_8hMl1rn83_1(.din(w_dff_B_PGQTR6aG6_1),.dout(w_dff_B_8hMl1rn83_1),.clk(gclk));
	jdff dff_B_oCnKrViL6_1(.din(w_dff_B_8hMl1rn83_1),.dout(w_dff_B_oCnKrViL6_1),.clk(gclk));
	jdff dff_B_U0pF2d0Q4_1(.din(w_dff_B_oCnKrViL6_1),.dout(w_dff_B_U0pF2d0Q4_1),.clk(gclk));
	jdff dff_B_sAkCvf2i1_1(.din(w_dff_B_U0pF2d0Q4_1),.dout(w_dff_B_sAkCvf2i1_1),.clk(gclk));
	jdff dff_B_Xuc4zKOq6_1(.din(w_dff_B_sAkCvf2i1_1),.dout(w_dff_B_Xuc4zKOq6_1),.clk(gclk));
	jdff dff_B_RgypynPF0_1(.din(w_dff_B_Xuc4zKOq6_1),.dout(w_dff_B_RgypynPF0_1),.clk(gclk));
	jdff dff_B_kRcWTs473_1(.din(w_dff_B_RgypynPF0_1),.dout(w_dff_B_kRcWTs473_1),.clk(gclk));
	jdff dff_B_mbZ9vNCi8_1(.din(w_dff_B_kRcWTs473_1),.dout(w_dff_B_mbZ9vNCi8_1),.clk(gclk));
	jdff dff_B_R05Mb3Zj5_1(.din(w_dff_B_mbZ9vNCi8_1),.dout(w_dff_B_R05Mb3Zj5_1),.clk(gclk));
	jdff dff_A_iDEZo0bi8_0(.dout(w_n854_4[0]),.din(w_dff_A_iDEZo0bi8_0),.clk(gclk));
	jdff dff_A_GUJ3mcq12_0(.dout(w_dff_A_iDEZo0bi8_0),.din(w_dff_A_GUJ3mcq12_0),.clk(gclk));
	jdff dff_A_oDOfYQRV4_0(.dout(w_dff_A_GUJ3mcq12_0),.din(w_dff_A_oDOfYQRV4_0),.clk(gclk));
	jdff dff_A_2PV4RARu0_0(.dout(w_dff_A_oDOfYQRV4_0),.din(w_dff_A_2PV4RARu0_0),.clk(gclk));
	jdff dff_A_AWzuBgCD8_0(.dout(w_dff_A_2PV4RARu0_0),.din(w_dff_A_AWzuBgCD8_0),.clk(gclk));
	jdff dff_A_Uv1SmpKj6_0(.dout(w_dff_A_AWzuBgCD8_0),.din(w_dff_A_Uv1SmpKj6_0),.clk(gclk));
	jdff dff_A_AerqLyH93_0(.dout(w_dff_A_Uv1SmpKj6_0),.din(w_dff_A_AerqLyH93_0),.clk(gclk));
	jdff dff_A_F5luKNX98_0(.dout(w_dff_A_AerqLyH93_0),.din(w_dff_A_F5luKNX98_0),.clk(gclk));
	jdff dff_B_GERK1vqb5_1(.din(n1063),.dout(w_dff_B_GERK1vqb5_1),.clk(gclk));
	jdff dff_B_B0CHzlMz8_1(.din(w_dff_B_GERK1vqb5_1),.dout(w_dff_B_B0CHzlMz8_1),.clk(gclk));
	jdff dff_B_dDPN7lR71_2(.din(G37),.dout(w_dff_B_dDPN7lR71_2),.clk(gclk));
	jdff dff_B_v2rBuvSz1_1(.din(n1075),.dout(w_dff_B_v2rBuvSz1_1),.clk(gclk));
	jdff dff_B_lKxiErD48_1(.din(w_dff_B_v2rBuvSz1_1),.dout(w_dff_B_lKxiErD48_1),.clk(gclk));
	jdff dff_B_gtujfV0o4_1(.din(w_dff_B_lKxiErD48_1),.dout(w_dff_B_gtujfV0o4_1),.clk(gclk));
	jdff dff_B_0EuHrGhe6_1(.din(w_dff_B_gtujfV0o4_1),.dout(w_dff_B_0EuHrGhe6_1),.clk(gclk));
	jdff dff_B_FLtnVVxT3_1(.din(w_dff_B_0EuHrGhe6_1),.dout(w_dff_B_FLtnVVxT3_1),.clk(gclk));
	jdff dff_B_BMfdatlS3_1(.din(w_dff_B_FLtnVVxT3_1),.dout(w_dff_B_BMfdatlS3_1),.clk(gclk));
	jdff dff_B_SYDRlI0o9_1(.din(w_dff_B_BMfdatlS3_1),.dout(w_dff_B_SYDRlI0o9_1),.clk(gclk));
	jdff dff_B_CAlsrD1v5_1(.din(w_dff_B_SYDRlI0o9_1),.dout(w_dff_B_CAlsrD1v5_1),.clk(gclk));
	jdff dff_B_YiHDiKMQ2_1(.din(w_dff_B_CAlsrD1v5_1),.dout(w_dff_B_YiHDiKMQ2_1),.clk(gclk));
	jdff dff_B_cWIjwMMG6_1(.din(w_dff_B_YiHDiKMQ2_1),.dout(w_dff_B_cWIjwMMG6_1),.clk(gclk));
	jdff dff_B_CEHtdWAg3_1(.din(w_dff_B_cWIjwMMG6_1),.dout(w_dff_B_CEHtdWAg3_1),.clk(gclk));
	jdff dff_B_bukuZ7MZ2_1(.din(w_dff_B_CEHtdWAg3_1),.dout(w_dff_B_bukuZ7MZ2_1),.clk(gclk));
	jdff dff_B_O435alBe3_1(.din(w_dff_B_bukuZ7MZ2_1),.dout(w_dff_B_O435alBe3_1),.clk(gclk));
	jdff dff_B_LimWu8Tx3_1(.din(w_dff_B_O435alBe3_1),.dout(w_dff_B_LimWu8Tx3_1),.clk(gclk));
	jdff dff_B_Lb1UTJyr6_0(.din(n1077),.dout(w_dff_B_Lb1UTJyr6_0),.clk(gclk));
	jdff dff_B_h7vnw1GH2_1(.din(n1072),.dout(w_dff_B_h7vnw1GH2_1),.clk(gclk));
	jdff dff_B_0rjRKGPo7_1(.din(w_dff_B_h7vnw1GH2_1),.dout(w_dff_B_0rjRKGPo7_1),.clk(gclk));
	jdff dff_A_N9HelVsD7_1(.dout(w_n852_8[1]),.din(w_dff_A_N9HelVsD7_1),.clk(gclk));
	jdff dff_A_pxtHcMGG8_1(.dout(w_dff_A_N9HelVsD7_1),.din(w_dff_A_pxtHcMGG8_1),.clk(gclk));
	jdff dff_A_XG7yHMMk8_1(.dout(w_dff_A_pxtHcMGG8_1),.din(w_dff_A_XG7yHMMk8_1),.clk(gclk));
	jdff dff_A_OV93YCTK4_1(.dout(w_dff_A_XG7yHMMk8_1),.din(w_dff_A_OV93YCTK4_1),.clk(gclk));
	jdff dff_A_iLu1TPBr6_1(.dout(w_dff_A_OV93YCTK4_1),.din(w_dff_A_iLu1TPBr6_1),.clk(gclk));
	jdff dff_A_Uv5qASFg5_1(.dout(w_dff_A_iLu1TPBr6_1),.din(w_dff_A_Uv5qASFg5_1),.clk(gclk));
	jdff dff_A_Wz3AUKzj7_1(.dout(w_dff_A_Uv5qASFg5_1),.din(w_dff_A_Wz3AUKzj7_1),.clk(gclk));
	jdff dff_A_1q8jEL7r5_1(.dout(w_dff_A_Wz3AUKzj7_1),.din(w_dff_A_1q8jEL7r5_1),.clk(gclk));
	jdff dff_A_Ia0vxgIO5_1(.dout(w_dff_A_1q8jEL7r5_1),.din(w_dff_A_Ia0vxgIO5_1),.clk(gclk));
	jdff dff_A_bykttAQo3_1(.dout(w_dff_A_Ia0vxgIO5_1),.din(w_dff_A_bykttAQo3_1),.clk(gclk));
	jdff dff_A_n88C7xSF6_1(.dout(w_dff_A_bykttAQo3_1),.din(w_dff_A_n88C7xSF6_1),.clk(gclk));
	jdff dff_A_KrLRbemN7_1(.dout(w_dff_A_n88C7xSF6_1),.din(w_dff_A_KrLRbemN7_1),.clk(gclk));
	jdff dff_A_uhEqaxQP3_1(.dout(w_dff_A_KrLRbemN7_1),.din(w_dff_A_uhEqaxQP3_1),.clk(gclk));
	jdff dff_A_n7XmxIk65_1(.dout(w_dff_A_uhEqaxQP3_1),.din(w_dff_A_n7XmxIk65_1),.clk(gclk));
	jdff dff_A_hSbRJQCb8_1(.dout(w_dff_A_n7XmxIk65_1),.din(w_dff_A_hSbRJQCb8_1),.clk(gclk));
	jdff dff_B_c1qR84vA7_2(.din(G20),.dout(w_dff_B_c1qR84vA7_2),.clk(gclk));
	jdff dff_A_xjhFeVW48_1(.dout(w_G4089_8[1]),.din(w_dff_A_xjhFeVW48_1),.clk(gclk));
	jdff dff_A_9xX7rbI98_1(.dout(w_dff_A_xjhFeVW48_1),.din(w_dff_A_9xX7rbI98_1),.clk(gclk));
	jdff dff_A_Grx4iNpn6_1(.dout(w_dff_A_9xX7rbI98_1),.din(w_dff_A_Grx4iNpn6_1),.clk(gclk));
	jdff dff_A_eDRVwpQg3_1(.dout(w_dff_A_Grx4iNpn6_1),.din(w_dff_A_eDRVwpQg3_1),.clk(gclk));
	jdff dff_A_AaLsFLOJ9_1(.dout(w_dff_A_eDRVwpQg3_1),.din(w_dff_A_AaLsFLOJ9_1),.clk(gclk));
	jdff dff_A_L2JRw27O9_1(.dout(w_dff_A_AaLsFLOJ9_1),.din(w_dff_A_L2JRw27O9_1),.clk(gclk));
	jdff dff_A_6if27TvK9_1(.dout(w_dff_A_L2JRw27O9_1),.din(w_dff_A_6if27TvK9_1),.clk(gclk));
	jdff dff_A_GTRcu69w7_1(.dout(w_dff_A_6if27TvK9_1),.din(w_dff_A_GTRcu69w7_1),.clk(gclk));
	jdff dff_A_DSNQ5J132_1(.dout(w_dff_A_GTRcu69w7_1),.din(w_dff_A_DSNQ5J132_1),.clk(gclk));
	jdff dff_A_6QIJxjfZ3_1(.dout(w_dff_A_DSNQ5J132_1),.din(w_dff_A_6QIJxjfZ3_1),.clk(gclk));
	jdff dff_A_xkF9HX0C0_1(.dout(w_dff_A_6QIJxjfZ3_1),.din(w_dff_A_xkF9HX0C0_1),.clk(gclk));
	jdff dff_A_4NcFoFno2_1(.dout(w_dff_A_xkF9HX0C0_1),.din(w_dff_A_4NcFoFno2_1),.clk(gclk));
	jdff dff_A_JOSlMOXr1_1(.dout(w_dff_A_4NcFoFno2_1),.din(w_dff_A_JOSlMOXr1_1),.clk(gclk));
	jdff dff_A_HznXxpI56_1(.dout(w_dff_A_JOSlMOXr1_1),.din(w_dff_A_HznXxpI56_1),.clk(gclk));
	jdff dff_A_80tlyiIj1_1(.dout(w_dff_A_HznXxpI56_1),.din(w_dff_A_80tlyiIj1_1),.clk(gclk));
	jdff dff_A_2ssKatZa8_1(.dout(w_dff_A_80tlyiIj1_1),.din(w_dff_A_2ssKatZa8_1),.clk(gclk));
	jdff dff_B_VQnQKQRU0_1(.din(n1084),.dout(w_dff_B_VQnQKQRU0_1),.clk(gclk));
	jdff dff_B_aigW7DO80_1(.din(w_dff_B_VQnQKQRU0_1),.dout(w_dff_B_aigW7DO80_1),.clk(gclk));
	jdff dff_B_rONFTPY69_1(.din(w_dff_B_aigW7DO80_1),.dout(w_dff_B_rONFTPY69_1),.clk(gclk));
	jdff dff_B_evSSdnCp8_1(.din(w_dff_B_rONFTPY69_1),.dout(w_dff_B_evSSdnCp8_1),.clk(gclk));
	jdff dff_B_N9oHBLAw4_1(.din(w_dff_B_evSSdnCp8_1),.dout(w_dff_B_N9oHBLAw4_1),.clk(gclk));
	jdff dff_B_8S2wpDdz9_1(.din(w_dff_B_N9oHBLAw4_1),.dout(w_dff_B_8S2wpDdz9_1),.clk(gclk));
	jdff dff_B_CzwBVkD16_1(.din(w_dff_B_8S2wpDdz9_1),.dout(w_dff_B_CzwBVkD16_1),.clk(gclk));
	jdff dff_B_o6snahXM1_1(.din(w_dff_B_CzwBVkD16_1),.dout(w_dff_B_o6snahXM1_1),.clk(gclk));
	jdff dff_B_w5Qd7Bf83_1(.din(w_dff_B_o6snahXM1_1),.dout(w_dff_B_w5Qd7Bf83_1),.clk(gclk));
	jdff dff_B_gpGkC0je6_1(.din(w_dff_B_w5Qd7Bf83_1),.dout(w_dff_B_gpGkC0je6_1),.clk(gclk));
	jdff dff_B_9aJWE6Au3_1(.din(w_dff_B_gpGkC0je6_1),.dout(w_dff_B_9aJWE6Au3_1),.clk(gclk));
	jdff dff_B_4iclhfl35_1(.din(w_dff_B_9aJWE6Au3_1),.dout(w_dff_B_4iclhfl35_1),.clk(gclk));
	jdff dff_B_VStuxuLR3_1(.din(n1081),.dout(w_dff_B_VStuxuLR3_1),.clk(gclk));
	jdff dff_B_KOtNylFL9_1(.din(w_dff_B_VStuxuLR3_1),.dout(w_dff_B_KOtNylFL9_1),.clk(gclk));
	jdff dff_A_0b42GaHs4_0(.dout(w_n852_7[0]),.din(w_dff_A_0b42GaHs4_0),.clk(gclk));
	jdff dff_A_HasVrbxU8_0(.dout(w_dff_A_0b42GaHs4_0),.din(w_dff_A_HasVrbxU8_0),.clk(gclk));
	jdff dff_A_coAWXkyc8_0(.dout(w_dff_A_HasVrbxU8_0),.din(w_dff_A_coAWXkyc8_0),.clk(gclk));
	jdff dff_A_fBLIayiT8_0(.dout(w_dff_A_coAWXkyc8_0),.din(w_dff_A_fBLIayiT8_0),.clk(gclk));
	jdff dff_A_qvAmdHs83_0(.dout(w_dff_A_fBLIayiT8_0),.din(w_dff_A_qvAmdHs83_0),.clk(gclk));
	jdff dff_A_gqhERKaS8_0(.dout(w_dff_A_qvAmdHs83_0),.din(w_dff_A_gqhERKaS8_0),.clk(gclk));
	jdff dff_A_Qicp42AP9_0(.dout(w_dff_A_gqhERKaS8_0),.din(w_dff_A_Qicp42AP9_0),.clk(gclk));
	jdff dff_A_ginIMhxv5_0(.dout(w_dff_A_Qicp42AP9_0),.din(w_dff_A_ginIMhxv5_0),.clk(gclk));
	jdff dff_A_eexujbIh5_0(.dout(w_dff_A_ginIMhxv5_0),.din(w_dff_A_eexujbIh5_0),.clk(gclk));
	jdff dff_A_KGVFU3zd0_0(.dout(w_dff_A_eexujbIh5_0),.din(w_dff_A_KGVFU3zd0_0),.clk(gclk));
	jdff dff_A_p4xrh6Df5_0(.dout(w_dff_A_KGVFU3zd0_0),.din(w_dff_A_p4xrh6Df5_0),.clk(gclk));
	jdff dff_A_8iaWdJjL1_0(.dout(w_dff_A_p4xrh6Df5_0),.din(w_dff_A_8iaWdJjL1_0),.clk(gclk));
	jdff dff_A_Ok4ajb1u1_2(.dout(w_n852_7[2]),.din(w_dff_A_Ok4ajb1u1_2),.clk(gclk));
	jdff dff_A_yRYfx1bf7_2(.dout(w_dff_A_Ok4ajb1u1_2),.din(w_dff_A_yRYfx1bf7_2),.clk(gclk));
	jdff dff_A_lc7V1lKu0_2(.dout(w_dff_A_yRYfx1bf7_2),.din(w_dff_A_lc7V1lKu0_2),.clk(gclk));
	jdff dff_A_cbFSyLib9_2(.dout(w_dff_A_lc7V1lKu0_2),.din(w_dff_A_cbFSyLib9_2),.clk(gclk));
	jdff dff_A_JmqDn6vc0_2(.dout(w_dff_A_cbFSyLib9_2),.din(w_dff_A_JmqDn6vc0_2),.clk(gclk));
	jdff dff_A_Iy704UMF1_2(.dout(w_dff_A_JmqDn6vc0_2),.din(w_dff_A_Iy704UMF1_2),.clk(gclk));
	jdff dff_A_yp9BvMpr8_2(.dout(w_dff_A_Iy704UMF1_2),.din(w_dff_A_yp9BvMpr8_2),.clk(gclk));
	jdff dff_A_j6B03wjY9_2(.dout(w_dff_A_yp9BvMpr8_2),.din(w_dff_A_j6B03wjY9_2),.clk(gclk));
	jdff dff_A_5QnVrgew1_2(.dout(w_dff_A_j6B03wjY9_2),.din(w_dff_A_5QnVrgew1_2),.clk(gclk));
	jdff dff_A_CcIk7B5N7_2(.dout(w_dff_A_5QnVrgew1_2),.din(w_dff_A_CcIk7B5N7_2),.clk(gclk));
	jdff dff_A_ZIM4o9Ut8_2(.dout(w_dff_A_CcIk7B5N7_2),.din(w_dff_A_ZIM4o9Ut8_2),.clk(gclk));
	jdff dff_A_jbxI6xua1_2(.dout(w_dff_A_ZIM4o9Ut8_2),.din(w_dff_A_jbxI6xua1_2),.clk(gclk));
	jdff dff_A_wEMJAAj20_2(.dout(w_dff_A_jbxI6xua1_2),.din(w_dff_A_wEMJAAj20_2),.clk(gclk));
	jdff dff_B_54uO2SaK2_2(.din(G17),.dout(w_dff_B_54uO2SaK2_2),.clk(gclk));
	jdff dff_A_UZk809mu4_0(.dout(w_G4089_7[0]),.din(w_dff_A_UZk809mu4_0),.clk(gclk));
	jdff dff_A_VW7VbnnE2_0(.dout(w_dff_A_UZk809mu4_0),.din(w_dff_A_VW7VbnnE2_0),.clk(gclk));
	jdff dff_A_HYaYbMfj2_0(.dout(w_dff_A_VW7VbnnE2_0),.din(w_dff_A_HYaYbMfj2_0),.clk(gclk));
	jdff dff_A_89gHHQnH9_0(.dout(w_dff_A_HYaYbMfj2_0),.din(w_dff_A_89gHHQnH9_0),.clk(gclk));
	jdff dff_A_NIac5FuB1_0(.dout(w_dff_A_89gHHQnH9_0),.din(w_dff_A_NIac5FuB1_0),.clk(gclk));
	jdff dff_A_g2GujtPk1_0(.dout(w_dff_A_NIac5FuB1_0),.din(w_dff_A_g2GujtPk1_0),.clk(gclk));
	jdff dff_A_PDkhJbq54_0(.dout(w_dff_A_g2GujtPk1_0),.din(w_dff_A_PDkhJbq54_0),.clk(gclk));
	jdff dff_A_hXanfFp21_0(.dout(w_dff_A_PDkhJbq54_0),.din(w_dff_A_hXanfFp21_0),.clk(gclk));
	jdff dff_A_B4F0XnhH6_0(.dout(w_dff_A_hXanfFp21_0),.din(w_dff_A_B4F0XnhH6_0),.clk(gclk));
	jdff dff_A_C9wvEsN02_0(.dout(w_dff_A_B4F0XnhH6_0),.din(w_dff_A_C9wvEsN02_0),.clk(gclk));
	jdff dff_A_1V4NTzXZ9_0(.dout(w_dff_A_C9wvEsN02_0),.din(w_dff_A_1V4NTzXZ9_0),.clk(gclk));
	jdff dff_A_c14cnpsO7_0(.dout(w_dff_A_1V4NTzXZ9_0),.din(w_dff_A_c14cnpsO7_0),.clk(gclk));
	jdff dff_A_oas7hLWv3_0(.dout(w_dff_A_c14cnpsO7_0),.din(w_dff_A_oas7hLWv3_0),.clk(gclk));
	jdff dff_A_nFqbBqfq5_2(.dout(w_G4089_7[2]),.din(w_dff_A_nFqbBqfq5_2),.clk(gclk));
	jdff dff_A_kdyrguMd8_2(.dout(w_dff_A_nFqbBqfq5_2),.din(w_dff_A_kdyrguMd8_2),.clk(gclk));
	jdff dff_A_pgRJUIvr9_2(.dout(w_dff_A_kdyrguMd8_2),.din(w_dff_A_pgRJUIvr9_2),.clk(gclk));
	jdff dff_A_WveXqnPt2_2(.dout(w_dff_A_pgRJUIvr9_2),.din(w_dff_A_WveXqnPt2_2),.clk(gclk));
	jdff dff_A_d3hGncqQ2_2(.dout(w_dff_A_WveXqnPt2_2),.din(w_dff_A_d3hGncqQ2_2),.clk(gclk));
	jdff dff_A_spm6nWV19_2(.dout(w_dff_A_d3hGncqQ2_2),.din(w_dff_A_spm6nWV19_2),.clk(gclk));
	jdff dff_A_BuoTJ5PJ1_2(.dout(w_dff_A_spm6nWV19_2),.din(w_dff_A_BuoTJ5PJ1_2),.clk(gclk));
	jdff dff_A_3SSokXxc4_2(.dout(w_dff_A_BuoTJ5PJ1_2),.din(w_dff_A_3SSokXxc4_2),.clk(gclk));
	jdff dff_A_u8fD9G8y0_2(.dout(w_dff_A_3SSokXxc4_2),.din(w_dff_A_u8fD9G8y0_2),.clk(gclk));
	jdff dff_A_mHf5WpV89_2(.dout(w_dff_A_u8fD9G8y0_2),.din(w_dff_A_mHf5WpV89_2),.clk(gclk));
	jdff dff_A_OyoOkfum3_2(.dout(w_dff_A_mHf5WpV89_2),.din(w_dff_A_OyoOkfum3_2),.clk(gclk));
	jdff dff_A_vMo8Fad50_2(.dout(w_dff_A_OyoOkfum3_2),.din(w_dff_A_vMo8Fad50_2),.clk(gclk));
	jdff dff_A_rwJY1WPL1_2(.dout(w_dff_A_vMo8Fad50_2),.din(w_dff_A_rwJY1WPL1_2),.clk(gclk));
	jdff dff_A_9KJNIPPm5_2(.dout(w_dff_A_rwJY1WPL1_2),.din(w_dff_A_9KJNIPPm5_2),.clk(gclk));
	jdff dff_A_caZmU7uz2_2(.dout(w_dff_A_9KJNIPPm5_2),.din(w_dff_A_caZmU7uz2_2),.clk(gclk));
	jdff dff_B_gudhFVs46_0(.din(n1097),.dout(w_dff_B_gudhFVs46_0),.clk(gclk));
	jdff dff_B_DqGdbygq5_0(.din(w_dff_B_gudhFVs46_0),.dout(w_dff_B_DqGdbygq5_0),.clk(gclk));
	jdff dff_B_IvNO6U535_0(.din(w_dff_B_DqGdbygq5_0),.dout(w_dff_B_IvNO6U535_0),.clk(gclk));
	jdff dff_B_b0fUwg5J6_0(.din(w_dff_B_IvNO6U535_0),.dout(w_dff_B_b0fUwg5J6_0),.clk(gclk));
	jdff dff_B_R84XIJoo9_0(.din(w_dff_B_b0fUwg5J6_0),.dout(w_dff_B_R84XIJoo9_0),.clk(gclk));
	jdff dff_B_cUYTpxcm3_0(.din(w_dff_B_R84XIJoo9_0),.dout(w_dff_B_cUYTpxcm3_0),.clk(gclk));
	jdff dff_B_oYPcxJV91_0(.din(w_dff_B_cUYTpxcm3_0),.dout(w_dff_B_oYPcxJV91_0),.clk(gclk));
	jdff dff_B_txNPpcLf6_0(.din(w_dff_B_oYPcxJV91_0),.dout(w_dff_B_txNPpcLf6_0),.clk(gclk));
	jdff dff_B_Tgv9zwm00_0(.din(w_dff_B_txNPpcLf6_0),.dout(w_dff_B_Tgv9zwm00_0),.clk(gclk));
	jdff dff_B_fn5qG8Ad1_0(.din(w_dff_B_Tgv9zwm00_0),.dout(w_dff_B_fn5qG8Ad1_0),.clk(gclk));
	jdff dff_B_GFwzuDQT0_0(.din(w_dff_B_fn5qG8Ad1_0),.dout(w_dff_B_GFwzuDQT0_0),.clk(gclk));
	jdff dff_B_MEU79m7I0_0(.din(w_dff_B_GFwzuDQT0_0),.dout(w_dff_B_MEU79m7I0_0),.clk(gclk));
	jdff dff_B_7shZPb5S7_0(.din(w_dff_B_MEU79m7I0_0),.dout(w_dff_B_7shZPb5S7_0),.clk(gclk));
	jdff dff_B_vohdLkQS8_0(.din(w_dff_B_7shZPb5S7_0),.dout(w_dff_B_vohdLkQS8_0),.clk(gclk));
	jdff dff_A_3CliLQJe9_1(.dout(w_G4090_3[1]),.din(w_dff_A_3CliLQJe9_1),.clk(gclk));
	jdff dff_A_sJEdiHEr5_2(.dout(w_G4090_3[2]),.din(w_dff_A_sJEdiHEr5_2),.clk(gclk));
	jdff dff_B_c7zUEjUl7_2(.din(G70),.dout(w_dff_B_c7zUEjUl7_2),.clk(gclk));
	jdff dff_B_Ydtt0Oin9_1(.din(n1090),.dout(w_dff_B_Ydtt0Oin9_1),.clk(gclk));
	jdff dff_B_X2YHWpL72_1(.din(w_dff_B_Ydtt0Oin9_1),.dout(w_dff_B_X2YHWpL72_1),.clk(gclk));
	jdff dff_B_w7zKmeRY0_1(.din(w_dff_B_X2YHWpL72_1),.dout(w_dff_B_w7zKmeRY0_1),.clk(gclk));
	jdff dff_A_1o31NhMe6_2(.dout(w_n854_3[2]),.din(w_dff_A_1o31NhMe6_2),.clk(gclk));
	jdff dff_A_TfsvbHxf8_2(.dout(w_dff_A_1o31NhMe6_2),.din(w_dff_A_TfsvbHxf8_2),.clk(gclk));
	jdff dff_B_vzT0zQNM9_0(.din(n1105),.dout(w_dff_B_vzT0zQNM9_0),.clk(gclk));
	jdff dff_B_97mNUZED7_0(.din(w_dff_B_vzT0zQNM9_0),.dout(w_dff_B_97mNUZED7_0),.clk(gclk));
	jdff dff_B_NJ7VpaXy6_0(.din(w_dff_B_97mNUZED7_0),.dout(w_dff_B_NJ7VpaXy6_0),.clk(gclk));
	jdff dff_B_X0LG8B3j2_0(.din(w_dff_B_NJ7VpaXy6_0),.dout(w_dff_B_X0LG8B3j2_0),.clk(gclk));
	jdff dff_B_OY2u0qCL7_0(.din(w_dff_B_X0LG8B3j2_0),.dout(w_dff_B_OY2u0qCL7_0),.clk(gclk));
	jdff dff_B_XD2yctU06_0(.din(w_dff_B_OY2u0qCL7_0),.dout(w_dff_B_XD2yctU06_0),.clk(gclk));
	jdff dff_B_iY4Mz0ZL5_0(.din(w_dff_B_XD2yctU06_0),.dout(w_dff_B_iY4Mz0ZL5_0),.clk(gclk));
	jdff dff_B_0DFwfqhO9_0(.din(w_dff_B_iY4Mz0ZL5_0),.dout(w_dff_B_0DFwfqhO9_0),.clk(gclk));
	jdff dff_B_ZycPv5oO8_0(.din(w_dff_B_0DFwfqhO9_0),.dout(w_dff_B_ZycPv5oO8_0),.clk(gclk));
	jdff dff_B_rvyPFMQt5_0(.din(w_dff_B_ZycPv5oO8_0),.dout(w_dff_B_rvyPFMQt5_0),.clk(gclk));
	jdff dff_B_C8aP4go06_0(.din(w_dff_B_rvyPFMQt5_0),.dout(w_dff_B_C8aP4go06_0),.clk(gclk));
	jdff dff_B_VclQYvSf9_0(.din(w_dff_B_C8aP4go06_0),.dout(w_dff_B_VclQYvSf9_0),.clk(gclk));
	jdff dff_B_UN6jiYz77_0(.din(w_dff_B_VclQYvSf9_0),.dout(w_dff_B_UN6jiYz77_0),.clk(gclk));
	jdff dff_B_kAtZXHiP9_0(.din(w_dff_B_UN6jiYz77_0),.dout(w_dff_B_kAtZXHiP9_0),.clk(gclk));
	jdff dff_B_whG8IqYl2_0(.din(w_dff_B_kAtZXHiP9_0),.dout(w_dff_B_whG8IqYl2_0),.clk(gclk));
	jdff dff_B_uHtD4vlp5_0(.din(n1104),.dout(w_dff_B_uHtD4vlp5_0),.clk(gclk));
	jdff dff_B_YTrvBkwS9_1(.din(n1099),.dout(w_dff_B_YTrvBkwS9_1),.clk(gclk));
	jdff dff_B_kIMNewnG9_0(.din(n1114),.dout(w_dff_B_kIMNewnG9_0),.clk(gclk));
	jdff dff_B_8hYkhCJR0_0(.din(w_dff_B_kIMNewnG9_0),.dout(w_dff_B_8hYkhCJR0_0),.clk(gclk));
	jdff dff_B_nu4abJga0_0(.din(w_dff_B_8hYkhCJR0_0),.dout(w_dff_B_nu4abJga0_0),.clk(gclk));
	jdff dff_B_PJtGooSC0_0(.din(w_dff_B_nu4abJga0_0),.dout(w_dff_B_PJtGooSC0_0),.clk(gclk));
	jdff dff_B_SgEkj2yl8_0(.din(w_dff_B_PJtGooSC0_0),.dout(w_dff_B_SgEkj2yl8_0),.clk(gclk));
	jdff dff_B_Cs7V7OsT2_0(.din(w_dff_B_SgEkj2yl8_0),.dout(w_dff_B_Cs7V7OsT2_0),.clk(gclk));
	jdff dff_B_c6oeIReX9_0(.din(w_dff_B_Cs7V7OsT2_0),.dout(w_dff_B_c6oeIReX9_0),.clk(gclk));
	jdff dff_B_BHwnXhEW7_0(.din(w_dff_B_c6oeIReX9_0),.dout(w_dff_B_BHwnXhEW7_0),.clk(gclk));
	jdff dff_B_p2bxcDom7_0(.din(w_dff_B_BHwnXhEW7_0),.dout(w_dff_B_p2bxcDom7_0),.clk(gclk));
	jdff dff_B_7Hydlfbz9_0(.din(w_dff_B_p2bxcDom7_0),.dout(w_dff_B_7Hydlfbz9_0),.clk(gclk));
	jdff dff_B_MO8fuRYc6_0(.din(w_dff_B_7Hydlfbz9_0),.dout(w_dff_B_MO8fuRYc6_0),.clk(gclk));
	jdff dff_B_EiX5KooM5_0(.din(w_dff_B_MO8fuRYc6_0),.dout(w_dff_B_EiX5KooM5_0),.clk(gclk));
	jdff dff_B_01lO3jCx5_0(.din(n1113),.dout(w_dff_B_01lO3jCx5_0),.clk(gclk));
	jdff dff_B_jKbWAgBq6_0(.din(n1110),.dout(w_dff_B_jKbWAgBq6_0),.clk(gclk));
	jdff dff_A_8rINv8s73_0(.dout(w_n999_3[0]),.din(w_dff_A_8rINv8s73_0),.clk(gclk));
	jdff dff_A_WMGHNPP52_0(.dout(w_dff_A_8rINv8s73_0),.din(w_dff_A_WMGHNPP52_0),.clk(gclk));
	jdff dff_A_eJjTXKVm4_0(.dout(w_dff_A_WMGHNPP52_0),.din(w_dff_A_eJjTXKVm4_0),.clk(gclk));
	jdff dff_A_38Agb6mp8_1(.dout(w_n999_3[1]),.din(w_dff_A_38Agb6mp8_1),.clk(gclk));
	jdff dff_A_xs2o5xqt0_1(.dout(w_dff_A_38Agb6mp8_1),.din(w_dff_A_xs2o5xqt0_1),.clk(gclk));
	jdff dff_A_Pxi0wDm27_1(.dout(w_dff_A_xs2o5xqt0_1),.din(w_dff_A_Pxi0wDm27_1),.clk(gclk));
	jdff dff_A_8fIelWnw4_1(.dout(w_dff_A_Pxi0wDm27_1),.din(w_dff_A_8fIelWnw4_1),.clk(gclk));
	jdff dff_A_62QZ4HDJ8_1(.dout(w_dff_A_8fIelWnw4_1),.din(w_dff_A_62QZ4HDJ8_1),.clk(gclk));
	jdff dff_A_JwLeYHrO6_1(.dout(w_dff_A_62QZ4HDJ8_1),.din(w_dff_A_JwLeYHrO6_1),.clk(gclk));
	jdff dff_A_se7hXFni1_1(.dout(w_dff_A_JwLeYHrO6_1),.din(w_dff_A_se7hXFni1_1),.clk(gclk));
	jdff dff_A_tBVgznO13_0(.dout(w_G1689_4[0]),.din(w_dff_A_tBVgznO13_0),.clk(gclk));
	jdff dff_A_mkuxMxtW7_0(.dout(w_dff_A_tBVgznO13_0),.din(w_dff_A_mkuxMxtW7_0),.clk(gclk));
	jdff dff_A_3309tWKO4_0(.dout(w_dff_A_mkuxMxtW7_0),.din(w_dff_A_3309tWKO4_0),.clk(gclk));
	jdff dff_A_BAG2IICU2_0(.dout(w_dff_A_3309tWKO4_0),.din(w_dff_A_BAG2IICU2_0),.clk(gclk));
	jdff dff_A_RaJD5xjh5_0(.dout(w_dff_A_BAG2IICU2_0),.din(w_dff_A_RaJD5xjh5_0),.clk(gclk));
	jdff dff_A_PiOZqbeA7_1(.dout(w_G1689_4[1]),.din(w_dff_A_PiOZqbeA7_1),.clk(gclk));
	jdff dff_A_3FxU5nc13_1(.dout(w_dff_A_PiOZqbeA7_1),.din(w_dff_A_3FxU5nc13_1),.clk(gclk));
	jdff dff_A_jMOXm3su3_1(.dout(w_dff_A_3FxU5nc13_1),.din(w_dff_A_jMOXm3su3_1),.clk(gclk));
	jdff dff_A_3pCUS7so0_1(.dout(w_dff_A_jMOXm3su3_1),.din(w_dff_A_3pCUS7so0_1),.clk(gclk));
	jdff dff_A_NOqqj6Mk0_1(.dout(w_dff_A_3pCUS7so0_1),.din(w_dff_A_NOqqj6Mk0_1),.clk(gclk));
	jdff dff_A_KmrKza565_1(.dout(w_dff_A_NOqqj6Mk0_1),.din(w_dff_A_KmrKza565_1),.clk(gclk));
	jdff dff_A_6BM9BGGk0_1(.dout(w_dff_A_KmrKza565_1),.din(w_dff_A_6BM9BGGk0_1),.clk(gclk));
	jdff dff_B_hEqM9Hw33_0(.din(n1123),.dout(w_dff_B_hEqM9Hw33_0),.clk(gclk));
	jdff dff_B_82pZnk8y6_0(.din(w_dff_B_hEqM9Hw33_0),.dout(w_dff_B_82pZnk8y6_0),.clk(gclk));
	jdff dff_B_SzKpfUr24_0(.din(w_dff_B_82pZnk8y6_0),.dout(w_dff_B_SzKpfUr24_0),.clk(gclk));
	jdff dff_B_wsVCZe921_0(.din(w_dff_B_SzKpfUr24_0),.dout(w_dff_B_wsVCZe921_0),.clk(gclk));
	jdff dff_B_l7FQPIQ24_0(.din(w_dff_B_wsVCZe921_0),.dout(w_dff_B_l7FQPIQ24_0),.clk(gclk));
	jdff dff_B_LRl3Xlgv4_0(.din(w_dff_B_l7FQPIQ24_0),.dout(w_dff_B_LRl3Xlgv4_0),.clk(gclk));
	jdff dff_B_fonvdCnR0_0(.din(w_dff_B_LRl3Xlgv4_0),.dout(w_dff_B_fonvdCnR0_0),.clk(gclk));
	jdff dff_B_tXsp4Gnj1_0(.din(w_dff_B_fonvdCnR0_0),.dout(w_dff_B_tXsp4Gnj1_0),.clk(gclk));
	jdff dff_B_pn6eVVIs8_0(.din(w_dff_B_tXsp4Gnj1_0),.dout(w_dff_B_pn6eVVIs8_0),.clk(gclk));
	jdff dff_B_TddAKzks3_0(.din(w_dff_B_pn6eVVIs8_0),.dout(w_dff_B_TddAKzks3_0),.clk(gclk));
	jdff dff_B_f2zBYRdW6_0(.din(w_dff_B_TddAKzks3_0),.dout(w_dff_B_f2zBYRdW6_0),.clk(gclk));
	jdff dff_B_yzIneDGH8_0(.din(w_dff_B_f2zBYRdW6_0),.dout(w_dff_B_yzIneDGH8_0),.clk(gclk));
	jdff dff_B_zLZyw14N6_0(.din(n1122),.dout(w_dff_B_zLZyw14N6_0),.clk(gclk));
	jdff dff_B_HPK9lmlb8_1(.din(n1117),.dout(w_dff_B_HPK9lmlb8_1),.clk(gclk));
	jdff dff_A_WB0fIQGN5_2(.dout(w_G137_8[2]),.din(w_dff_A_WB0fIQGN5_2),.clk(gclk));
	jdff dff_A_KIUPQkRY8_2(.dout(w_dff_A_WB0fIQGN5_2),.din(w_dff_A_KIUPQkRY8_2),.clk(gclk));
	jdff dff_A_tbNmrbzc5_2(.dout(w_dff_A_KIUPQkRY8_2),.din(w_dff_A_tbNmrbzc5_2),.clk(gclk));
	jdff dff_B_IrZilIV99_0(.din(n1132),.dout(w_dff_B_IrZilIV99_0),.clk(gclk));
	jdff dff_B_BHVBc84c2_0(.din(w_dff_B_IrZilIV99_0),.dout(w_dff_B_BHVBc84c2_0),.clk(gclk));
	jdff dff_B_jXuyVCod4_0(.din(w_dff_B_BHVBc84c2_0),.dout(w_dff_B_jXuyVCod4_0),.clk(gclk));
	jdff dff_B_V7LK8I483_0(.din(w_dff_B_jXuyVCod4_0),.dout(w_dff_B_V7LK8I483_0),.clk(gclk));
	jdff dff_B_YJWGexCA6_0(.din(w_dff_B_V7LK8I483_0),.dout(w_dff_B_YJWGexCA6_0),.clk(gclk));
	jdff dff_B_uWr62opr2_0(.din(w_dff_B_YJWGexCA6_0),.dout(w_dff_B_uWr62opr2_0),.clk(gclk));
	jdff dff_B_kuzGrrfn5_0(.din(w_dff_B_uWr62opr2_0),.dout(w_dff_B_kuzGrrfn5_0),.clk(gclk));
	jdff dff_B_hBm8z6RF3_0(.din(w_dff_B_kuzGrrfn5_0),.dout(w_dff_B_hBm8z6RF3_0),.clk(gclk));
	jdff dff_B_GHnnGyVa1_0(.din(w_dff_B_hBm8z6RF3_0),.dout(w_dff_B_GHnnGyVa1_0),.clk(gclk));
	jdff dff_B_P6iuIBXH4_0(.din(w_dff_B_GHnnGyVa1_0),.dout(w_dff_B_P6iuIBXH4_0),.clk(gclk));
	jdff dff_B_wzegfj990_0(.din(w_dff_B_P6iuIBXH4_0),.dout(w_dff_B_wzegfj990_0),.clk(gclk));
	jdff dff_B_YUOZX00c4_0(.din(w_dff_B_wzegfj990_0),.dout(w_dff_B_YUOZX00c4_0),.clk(gclk));
	jdff dff_B_ytrX5FtM3_0(.din(w_dff_B_YUOZX00c4_0),.dout(w_dff_B_ytrX5FtM3_0),.clk(gclk));
	jdff dff_B_1gDrkq6x2_0(.din(n1131),.dout(w_dff_B_1gDrkq6x2_0),.clk(gclk));
	jdff dff_A_8lDlWQtO6_0(.dout(w_n993_3[0]),.din(w_dff_A_8lDlWQtO6_0),.clk(gclk));
	jdff dff_A_VwRZDwaz7_0(.dout(w_dff_A_8lDlWQtO6_0),.din(w_dff_A_VwRZDwaz7_0),.clk(gclk));
	jdff dff_A_CC2qWIf52_1(.dout(w_n993_3[1]),.din(w_dff_A_CC2qWIf52_1),.clk(gclk));
	jdff dff_B_EqsrlkAY9_1(.din(n1135),.dout(w_dff_B_EqsrlkAY9_1),.clk(gclk));
	jdff dff_B_jHZRUrdB5_1(.din(w_dff_B_EqsrlkAY9_1),.dout(w_dff_B_jHZRUrdB5_1),.clk(gclk));
	jdff dff_B_aBQHPIZc5_1(.din(w_dff_B_jHZRUrdB5_1),.dout(w_dff_B_aBQHPIZc5_1),.clk(gclk));
	jdff dff_B_GGtYoyhv6_1(.din(w_dff_B_aBQHPIZc5_1),.dout(w_dff_B_GGtYoyhv6_1),.clk(gclk));
	jdff dff_B_TQGPFfCw7_1(.din(w_dff_B_GGtYoyhv6_1),.dout(w_dff_B_TQGPFfCw7_1),.clk(gclk));
	jdff dff_B_v8xPUZ0R9_1(.din(w_dff_B_TQGPFfCw7_1),.dout(w_dff_B_v8xPUZ0R9_1),.clk(gclk));
	jdff dff_B_TAsVhcUW7_1(.din(w_dff_B_v8xPUZ0R9_1),.dout(w_dff_B_TAsVhcUW7_1),.clk(gclk));
	jdff dff_B_ZZS7ScBr7_1(.din(w_dff_B_TAsVhcUW7_1),.dout(w_dff_B_ZZS7ScBr7_1),.clk(gclk));
	jdff dff_B_MBEZ6rRW8_1(.din(w_dff_B_ZZS7ScBr7_1),.dout(w_dff_B_MBEZ6rRW8_1),.clk(gclk));
	jdff dff_B_N0in5UnQ0_1(.din(w_dff_B_MBEZ6rRW8_1),.dout(w_dff_B_N0in5UnQ0_1),.clk(gclk));
	jdff dff_B_fYRue3RB7_1(.din(w_dff_B_N0in5UnQ0_1),.dout(w_dff_B_fYRue3RB7_1),.clk(gclk));
	jdff dff_B_ucU94RGc6_1(.din(w_dff_B_fYRue3RB7_1),.dout(w_dff_B_ucU94RGc6_1),.clk(gclk));
	jdff dff_B_VzIQXCFb0_1(.din(w_dff_B_ucU94RGc6_1),.dout(w_dff_B_VzIQXCFb0_1),.clk(gclk));
	jdff dff_B_1KsPs9Jb0_1(.din(w_dff_B_VzIQXCFb0_1),.dout(w_dff_B_1KsPs9Jb0_1),.clk(gclk));
	jdff dff_B_BlvpqnAG2_1(.din(w_dff_B_1KsPs9Jb0_1),.dout(w_dff_B_BlvpqnAG2_1),.clk(gclk));
	jdff dff_B_7oZaUpvj9_1(.din(w_dff_B_BlvpqnAG2_1),.dout(w_dff_B_7oZaUpvj9_1),.clk(gclk));
	jdff dff_B_l8beA7pM1_1(.din(w_dff_B_7oZaUpvj9_1),.dout(w_dff_B_l8beA7pM1_1),.clk(gclk));
	jdff dff_B_07b8zMqv5_1(.din(n1136),.dout(w_dff_B_07b8zMqv5_1),.clk(gclk));
	jdff dff_B_UtSEGdzN4_1(.din(w_dff_B_07b8zMqv5_1),.dout(w_dff_B_UtSEGdzN4_1),.clk(gclk));
	jdff dff_B_0WME3dXU5_1(.din(w_dff_B_UtSEGdzN4_1),.dout(w_dff_B_0WME3dXU5_1),.clk(gclk));
	jdff dff_B_Chuzd4SF0_1(.din(w_dff_B_0WME3dXU5_1),.dout(w_dff_B_Chuzd4SF0_1),.clk(gclk));
	jdff dff_B_x9F0mnhp2_1(.din(w_dff_B_Chuzd4SF0_1),.dout(w_dff_B_x9F0mnhp2_1),.clk(gclk));
	jdff dff_B_5DvTuiwh8_1(.din(w_dff_B_x9F0mnhp2_1),.dout(w_dff_B_5DvTuiwh8_1),.clk(gclk));
	jdff dff_B_q6572KBE3_1(.din(w_dff_B_5DvTuiwh8_1),.dout(w_dff_B_q6572KBE3_1),.clk(gclk));
	jdff dff_B_jvNVoFVk8_1(.din(w_dff_B_q6572KBE3_1),.dout(w_dff_B_jvNVoFVk8_1),.clk(gclk));
	jdff dff_B_rT3rqSo23_1(.din(w_dff_B_jvNVoFVk8_1),.dout(w_dff_B_rT3rqSo23_1),.clk(gclk));
	jdff dff_B_FPhCeDhE9_1(.din(w_dff_B_rT3rqSo23_1),.dout(w_dff_B_FPhCeDhE9_1),.clk(gclk));
	jdff dff_B_D5DDbU3o9_1(.din(w_dff_B_FPhCeDhE9_1),.dout(w_dff_B_D5DDbU3o9_1),.clk(gclk));
	jdff dff_B_ROLApdNa1_1(.din(w_dff_B_D5DDbU3o9_1),.dout(w_dff_B_ROLApdNa1_1),.clk(gclk));
	jdff dff_B_WKTjbkHm1_1(.din(w_dff_B_ROLApdNa1_1),.dout(w_dff_B_WKTjbkHm1_1),.clk(gclk));
	jdff dff_B_nrtzlCTv5_1(.din(w_dff_B_WKTjbkHm1_1),.dout(w_dff_B_nrtzlCTv5_1),.clk(gclk));
	jdff dff_B_GmlogMg49_1(.din(w_dff_B_nrtzlCTv5_1),.dout(w_dff_B_GmlogMg49_1),.clk(gclk));
	jdff dff_B_06DKGFZm7_1(.din(w_dff_B_GmlogMg49_1),.dout(w_dff_B_06DKGFZm7_1),.clk(gclk));
	jdff dff_B_Zah5riXS9_1(.din(w_dff_B_06DKGFZm7_1),.dout(w_dff_B_Zah5riXS9_1),.clk(gclk));
	jdff dff_B_A8p3AAgU4_1(.din(n811),.dout(w_dff_B_A8p3AAgU4_1),.clk(gclk));
	jdff dff_B_2UMaT1uP5_1(.din(w_dff_B_A8p3AAgU4_1),.dout(w_dff_B_2UMaT1uP5_1),.clk(gclk));
	jdff dff_B_2E2F5T8i2_1(.din(w_dff_B_2UMaT1uP5_1),.dout(w_dff_B_2E2F5T8i2_1),.clk(gclk));
	jdff dff_B_CC2gThHC7_1(.din(w_dff_B_2E2F5T8i2_1),.dout(w_dff_B_CC2gThHC7_1),.clk(gclk));
	jdff dff_B_zk9vWeIP4_1(.din(w_dff_B_CC2gThHC7_1),.dout(w_dff_B_zk9vWeIP4_1),.clk(gclk));
	jdff dff_B_fEbiifXh7_1(.din(w_dff_B_zk9vWeIP4_1),.dout(w_dff_B_fEbiifXh7_1),.clk(gclk));
	jdff dff_B_PLgQJAgZ1_1(.din(w_dff_B_fEbiifXh7_1),.dout(w_dff_B_PLgQJAgZ1_1),.clk(gclk));
	jdff dff_B_AlFxG4ep9_1(.din(w_dff_B_PLgQJAgZ1_1),.dout(w_dff_B_AlFxG4ep9_1),.clk(gclk));
	jdff dff_B_PVCJ2hWw0_1(.din(w_dff_B_AlFxG4ep9_1),.dout(w_dff_B_PVCJ2hWw0_1),.clk(gclk));
	jdff dff_B_4eTKlpJq8_1(.din(w_dff_B_PVCJ2hWw0_1),.dout(w_dff_B_4eTKlpJq8_1),.clk(gclk));
	jdff dff_B_W7L2ew7r4_0(.din(n830),.dout(w_dff_B_W7L2ew7r4_0),.clk(gclk));
	jdff dff_B_zBDlRoN46_0(.din(w_dff_B_W7L2ew7r4_0),.dout(w_dff_B_zBDlRoN46_0),.clk(gclk));
	jdff dff_B_089RRlJP9_0(.din(w_dff_B_zBDlRoN46_0),.dout(w_dff_B_089RRlJP9_0),.clk(gclk));
	jdff dff_B_JCYl6Vhl2_0(.din(w_dff_B_089RRlJP9_0),.dout(w_dff_B_JCYl6Vhl2_0),.clk(gclk));
	jdff dff_B_BSCnZAbv7_0(.din(w_dff_B_JCYl6Vhl2_0),.dout(w_dff_B_BSCnZAbv7_0),.clk(gclk));
	jdff dff_B_UIS0n0cy6_0(.din(w_dff_B_BSCnZAbv7_0),.dout(w_dff_B_UIS0n0cy6_0),.clk(gclk));
	jdff dff_B_w0Q4eRMQ9_1(.din(n441),.dout(w_dff_B_w0Q4eRMQ9_1),.clk(gclk));
	jdff dff_B_f9YYUJeb7_1(.din(n436),.dout(w_dff_B_f9YYUJeb7_1),.clk(gclk));
	jdff dff_B_Gez3os9P9_1(.din(n822),.dout(w_dff_B_Gez3os9P9_1),.clk(gclk));
	jdff dff_B_O6iMNlxl3_1(.din(w_dff_B_Gez3os9P9_1),.dout(w_dff_B_O6iMNlxl3_1),.clk(gclk));
	jdff dff_B_i9fWGNyT8_1(.din(w_dff_B_O6iMNlxl3_1),.dout(w_dff_B_i9fWGNyT8_1),.clk(gclk));
	jdff dff_B_X2fQecv99_1(.din(w_dff_B_i9fWGNyT8_1),.dout(w_dff_B_X2fQecv99_1),.clk(gclk));
	jdff dff_B_xAtnCFNh5_1(.din(w_dff_B_X2fQecv99_1),.dout(w_dff_B_xAtnCFNh5_1),.clk(gclk));
	jdff dff_B_CQYza13j0_1(.din(G52),.dout(w_dff_B_CQYza13j0_1),.clk(gclk));
	jdff dff_B_E1lXjz2A0_1(.din(w_dff_B_CQYza13j0_1),.dout(w_dff_B_E1lXjz2A0_1),.clk(gclk));
	jdff dff_B_YFG3Hif90_1(.din(n864),.dout(w_dff_B_YFG3Hif90_1),.clk(gclk));
	jdff dff_B_0QZLWL4B4_1(.din(w_dff_B_YFG3Hif90_1),.dout(w_dff_B_0QZLWL4B4_1),.clk(gclk));
	jdff dff_B_SOpIKrXM3_1(.din(w_dff_B_0QZLWL4B4_1),.dout(w_dff_B_SOpIKrXM3_1),.clk(gclk));
	jdff dff_B_qJMxlCiJ1_1(.din(w_dff_B_SOpIKrXM3_1),.dout(w_dff_B_qJMxlCiJ1_1),.clk(gclk));
	jdff dff_B_unc3xdOr2_1(.din(w_dff_B_qJMxlCiJ1_1),.dout(w_dff_B_unc3xdOr2_1),.clk(gclk));
	jdff dff_B_WYWrfO6q3_1(.din(w_dff_B_unc3xdOr2_1),.dout(w_dff_B_WYWrfO6q3_1),.clk(gclk));
	jdff dff_B_dLBtxQ8b9_1(.din(w_dff_B_WYWrfO6q3_1),.dout(w_dff_B_dLBtxQ8b9_1),.clk(gclk));
	jdff dff_B_Mg9x6ze98_1(.din(w_dff_B_dLBtxQ8b9_1),.dout(w_dff_B_Mg9x6ze98_1),.clk(gclk));
	jdff dff_B_5VSO5p555_1(.din(w_dff_B_Mg9x6ze98_1),.dout(w_dff_B_5VSO5p555_1),.clk(gclk));
	jdff dff_B_bhV7aBCh0_1(.din(w_dff_B_5VSO5p555_1),.dout(w_dff_B_bhV7aBCh0_1),.clk(gclk));
	jdff dff_B_xHA3HxgH1_0(.din(n874),.dout(w_dff_B_xHA3HxgH1_0),.clk(gclk));
	jdff dff_B_rfXfVhsf2_0(.din(w_dff_B_xHA3HxgH1_0),.dout(w_dff_B_rfXfVhsf2_0),.clk(gclk));
	jdff dff_B_YAiDbcMe4_0(.din(w_dff_B_rfXfVhsf2_0),.dout(w_dff_B_YAiDbcMe4_0),.clk(gclk));
	jdff dff_B_IQzoHech8_0(.din(w_dff_B_YAiDbcMe4_0),.dout(w_dff_B_IQzoHech8_0),.clk(gclk));
	jdff dff_B_OzL3IZBd2_0(.din(w_dff_B_IQzoHech8_0),.dout(w_dff_B_OzL3IZBd2_0),.clk(gclk));
	jdff dff_B_WLwaQdrP9_0(.din(w_dff_B_OzL3IZBd2_0),.dout(w_dff_B_WLwaQdrP9_0),.clk(gclk));
	jdff dff_B_7ogaCzHa8_1(.din(n466),.dout(w_dff_B_7ogaCzHa8_1),.clk(gclk));
	jdff dff_B_E4vL1V1K6_1(.din(n461),.dout(w_dff_B_E4vL1V1K6_1),.clk(gclk));
	jdff dff_B_wrJwdZHd9_1(.din(G122),.dout(w_dff_B_wrJwdZHd9_1),.clk(gclk));
	jdff dff_B_G7WvKJ7j7_1(.din(w_dff_B_wrJwdZHd9_1),.dout(w_dff_B_G7WvKJ7j7_1),.clk(gclk));
	jdff dff_B_fV1F7oBh6_2(.din(G170),.dout(w_dff_B_fV1F7oBh6_2),.clk(gclk));
	jdff dff_B_3Dl9XxUb6_2(.din(G200),.dout(w_dff_B_3Dl9XxUb6_2),.clk(gclk));
	jdff dff_B_Zm4pvZX48_2(.din(w_dff_B_3Dl9XxUb6_2),.dout(w_dff_B_Zm4pvZX48_2),.clk(gclk));
	jdff dff_B_nbNfm5IV3_0(.din(n1150),.dout(w_dff_B_nbNfm5IV3_0),.clk(gclk));
	jdff dff_B_0leJRDAP4_0(.din(w_dff_B_nbNfm5IV3_0),.dout(w_dff_B_0leJRDAP4_0),.clk(gclk));
	jdff dff_B_VeiRMqA10_0(.din(w_dff_B_0leJRDAP4_0),.dout(w_dff_B_VeiRMqA10_0),.clk(gclk));
	jdff dff_B_GAdN59NS5_0(.din(w_dff_B_VeiRMqA10_0),.dout(w_dff_B_GAdN59NS5_0),.clk(gclk));
	jdff dff_B_D40llUlT4_0(.din(w_dff_B_GAdN59NS5_0),.dout(w_dff_B_D40llUlT4_0),.clk(gclk));
	jdff dff_B_QejdSoeG8_0(.din(w_dff_B_D40llUlT4_0),.dout(w_dff_B_QejdSoeG8_0),.clk(gclk));
	jdff dff_B_5Dl9fguZ6_0(.din(w_dff_B_QejdSoeG8_0),.dout(w_dff_B_5Dl9fguZ6_0),.clk(gclk));
	jdff dff_B_0CnjIi0W3_0(.din(w_dff_B_5Dl9fguZ6_0),.dout(w_dff_B_0CnjIi0W3_0),.clk(gclk));
	jdff dff_B_WV9Yg7W70_0(.din(w_dff_B_0CnjIi0W3_0),.dout(w_dff_B_WV9Yg7W70_0),.clk(gclk));
	jdff dff_B_lv6Mg72Q9_0(.din(w_dff_B_WV9Yg7W70_0),.dout(w_dff_B_lv6Mg72Q9_0),.clk(gclk));
	jdff dff_B_7fhbX3HY4_0(.din(w_dff_B_lv6Mg72Q9_0),.dout(w_dff_B_7fhbX3HY4_0),.clk(gclk));
	jdff dff_B_J0McyiMk6_0(.din(w_dff_B_7fhbX3HY4_0),.dout(w_dff_B_J0McyiMk6_0),.clk(gclk));
	jdff dff_B_y1UOWzRD6_0(.din(n1149),.dout(w_dff_B_y1UOWzRD6_0),.clk(gclk));
	jdff dff_B_UGVHS3ko5_2(.din(G158),.dout(w_dff_B_UGVHS3ko5_2),.clk(gclk));
	jdff dff_B_lu2Jmb9Z9_2(.din(G188),.dout(w_dff_B_lu2Jmb9Z9_2),.clk(gclk));
	jdff dff_B_HOpJCSUc9_2(.din(w_dff_B_lu2Jmb9Z9_2),.dout(w_dff_B_HOpJCSUc9_2),.clk(gclk));
	jdff dff_B_pivs3WiK7_0(.din(n1146),.dout(w_dff_B_pivs3WiK7_0),.clk(gclk));
	jdff dff_B_u74rHInI8_1(.din(n897),.dout(w_dff_B_u74rHInI8_1),.clk(gclk));
	jdff dff_B_axjqmemQ7_1(.din(w_dff_B_u74rHInI8_1),.dout(w_dff_B_axjqmemQ7_1),.clk(gclk));
	jdff dff_B_15dOJZD46_1(.din(w_dff_B_axjqmemQ7_1),.dout(w_dff_B_15dOJZD46_1),.clk(gclk));
	jdff dff_B_d1IJW1IA7_1(.din(w_dff_B_15dOJZD46_1),.dout(w_dff_B_d1IJW1IA7_1),.clk(gclk));
	jdff dff_B_QFF1pcNc9_1(.din(w_dff_B_d1IJW1IA7_1),.dout(w_dff_B_QFF1pcNc9_1),.clk(gclk));
	jdff dff_B_Nwaz4MU14_1(.din(w_dff_B_QFF1pcNc9_1),.dout(w_dff_B_Nwaz4MU14_1),.clk(gclk));
	jdff dff_B_gsZrcHqF9_0(.din(n904),.dout(w_dff_B_gsZrcHqF9_0),.clk(gclk));
	jdff dff_B_i3OubGyD6_0(.din(w_dff_B_gsZrcHqF9_0),.dout(w_dff_B_i3OubGyD6_0),.clk(gclk));
	jdff dff_B_24dM6nyX0_1(.din(n477),.dout(w_dff_B_24dM6nyX0_1),.clk(gclk));
	jdff dff_B_GSMPQl2M4_1(.din(n472),.dout(w_dff_B_GSMPQl2M4_1),.clk(gclk));
	jdff dff_A_L34K2jlO5_0(.dout(w_n901_0[0]),.din(w_dff_A_L34K2jlO5_0),.clk(gclk));
	jdff dff_A_a2QCXQJn3_0(.dout(w_dff_A_L34K2jlO5_0),.din(w_dff_A_a2QCXQJn3_0),.clk(gclk));
	jdff dff_B_0JWCdQHO9_1(.din(n898),.dout(w_dff_B_0JWCdQHO9_1),.clk(gclk));
	jdff dff_B_23LC9GOZ8_1(.din(G126),.dout(w_dff_B_23LC9GOZ8_1),.clk(gclk));
	jdff dff_B_IX2dHluj9_1(.din(w_dff_B_23LC9GOZ8_1),.dout(w_dff_B_IX2dHluj9_1),.clk(gclk));
	jdff dff_A_L20R3OvP1_0(.dout(w_n1007_3[0]),.din(w_dff_A_L20R3OvP1_0),.clk(gclk));
	jdff dff_A_kKypQXJj3_1(.dout(w_n1007_3[1]),.din(w_dff_A_kKypQXJj3_1),.clk(gclk));
	jdff dff_A_eaZBJOnx8_1(.dout(w_dff_A_kKypQXJj3_1),.din(w_dff_A_eaZBJOnx8_1),.clk(gclk));
	jdff dff_A_mbsEs87r4_1(.dout(w_dff_A_eaZBJOnx8_1),.din(w_dff_A_mbsEs87r4_1),.clk(gclk));
	jdff dff_A_KOawNj8j2_1(.dout(w_dff_A_mbsEs87r4_1),.din(w_dff_A_KOawNj8j2_1),.clk(gclk));
	jdff dff_A_MiXGg6Hi7_1(.dout(w_dff_A_KOawNj8j2_1),.din(w_dff_A_MiXGg6Hi7_1),.clk(gclk));
	jdff dff_A_3SCYQOmj0_1(.dout(w_dff_A_MiXGg6Hi7_1),.din(w_dff_A_3SCYQOmj0_1),.clk(gclk));
	jdff dff_B_pcbEym5T3_1(.din(n762),.dout(w_dff_B_pcbEym5T3_1),.clk(gclk));
	jdff dff_B_LmUy60EZ2_1(.din(w_dff_B_pcbEym5T3_1),.dout(w_dff_B_LmUy60EZ2_1),.clk(gclk));
	jdff dff_B_Tqqg0m4r6_1(.din(w_dff_B_LmUy60EZ2_1),.dout(w_dff_B_Tqqg0m4r6_1),.clk(gclk));
	jdff dff_B_iOoWjQo79_1(.din(w_dff_B_Tqqg0m4r6_1),.dout(w_dff_B_iOoWjQo79_1),.clk(gclk));
	jdff dff_B_jhURF59J7_1(.din(w_dff_B_iOoWjQo79_1),.dout(w_dff_B_jhURF59J7_1),.clk(gclk));
	jdff dff_B_OxIp23Sa1_1(.din(w_dff_B_jhURF59J7_1),.dout(w_dff_B_OxIp23Sa1_1),.clk(gclk));
	jdff dff_B_5iz5ATwb1_1(.din(w_dff_B_OxIp23Sa1_1),.dout(w_dff_B_5iz5ATwb1_1),.clk(gclk));
	jdff dff_B_4w5sM2TQ6_1(.din(w_dff_B_5iz5ATwb1_1),.dout(w_dff_B_4w5sM2TQ6_1),.clk(gclk));
	jdff dff_B_J0DbFJi31_0(.din(n773),.dout(w_dff_B_J0DbFJi31_0),.clk(gclk));
	jdff dff_B_vxSfaeuF8_0(.din(w_dff_B_J0DbFJi31_0),.dout(w_dff_B_vxSfaeuF8_0),.clk(gclk));
	jdff dff_B_pv4rlYUd0_0(.din(w_dff_B_vxSfaeuF8_0),.dout(w_dff_B_pv4rlYUd0_0),.clk(gclk));
	jdff dff_B_QreqmqU37_0(.din(w_dff_B_pv4rlYUd0_0),.dout(w_dff_B_QreqmqU37_0),.clk(gclk));
	jdff dff_B_QIFB1MSw6_1(.din(n382),.dout(w_dff_B_QIFB1MSw6_1),.clk(gclk));
	jdff dff_B_SyeDNte46_1(.din(n376),.dout(w_dff_B_SyeDNte46_1),.clk(gclk));
	jdff dff_B_26RCtZf59_0(.din(n769),.dout(w_dff_B_26RCtZf59_0),.clk(gclk));
	jdff dff_B_V8ceVBG67_0(.din(w_dff_B_26RCtZf59_0),.dout(w_dff_B_V8ceVBG67_0),.clk(gclk));
	jdff dff_B_Zajdvmtw0_0(.din(w_dff_B_V8ceVBG67_0),.dout(w_dff_B_Zajdvmtw0_0),.clk(gclk));
	jdff dff_B_fqdV4id69_0(.din(w_dff_B_Zajdvmtw0_0),.dout(w_dff_B_fqdV4id69_0),.clk(gclk));
	jdff dff_A_cdVVsjCe9_0(.dout(w_n753_1[0]),.din(w_dff_A_cdVVsjCe9_0),.clk(gclk));
	jdff dff_A_tIMtKK4g7_0(.dout(w_dff_A_cdVVsjCe9_0),.din(w_dff_A_tIMtKK4g7_0),.clk(gclk));
	jdff dff_A_k97jq2Wn5_0(.dout(w_dff_A_tIMtKK4g7_0),.din(w_dff_A_k97jq2Wn5_0),.clk(gclk));
	jdff dff_A_wja9FsvO5_0(.dout(w_dff_A_k97jq2Wn5_0),.din(w_dff_A_wja9FsvO5_0),.clk(gclk));
	jdff dff_A_l8pysX0x7_0(.dout(w_dff_A_wja9FsvO5_0),.din(w_dff_A_l8pysX0x7_0),.clk(gclk));
	jdff dff_A_FuIfPWWe8_0(.dout(w_G4091_5[0]),.din(w_dff_A_FuIfPWWe8_0),.clk(gclk));
	jdff dff_A_WU9mHmMW4_0(.dout(w_dff_A_FuIfPWWe8_0),.din(w_dff_A_WU9mHmMW4_0),.clk(gclk));
	jdff dff_A_fxBZz2dK4_0(.dout(w_dff_A_WU9mHmMW4_0),.din(w_dff_A_fxBZz2dK4_0),.clk(gclk));
	jdff dff_A_qfAREajh4_0(.dout(w_dff_A_fxBZz2dK4_0),.din(w_dff_A_qfAREajh4_0),.clk(gclk));
	jdff dff_A_wJpX3Al28_0(.dout(w_dff_A_qfAREajh4_0),.din(w_dff_A_wJpX3Al28_0),.clk(gclk));
	jdff dff_A_h5HoD7D52_2(.dout(w_G4091_5[2]),.din(w_dff_A_h5HoD7D52_2),.clk(gclk));
	jdff dff_A_Lg6FT8AN9_2(.dout(w_dff_A_h5HoD7D52_2),.din(w_dff_A_Lg6FT8AN9_2),.clk(gclk));
	jdff dff_A_2NvsHdUV5_2(.dout(w_dff_A_Lg6FT8AN9_2),.din(w_dff_A_2NvsHdUV5_2),.clk(gclk));
	jdff dff_B_Bo2dviGY1_1(.din(G129),.dout(w_dff_B_Bo2dviGY1_1),.clk(gclk));
	jdff dff_B_BIz860tW5_1(.din(w_dff_B_Bo2dviGY1_1),.dout(w_dff_B_BIz860tW5_1),.clk(gclk));
	jdff dff_A_sDoJ2deg5_1(.dout(w_G137_7[1]),.din(w_dff_A_sDoJ2deg5_1),.clk(gclk));
	jdff dff_A_UctEwY1H7_1(.dout(w_dff_A_sDoJ2deg5_1),.din(w_dff_A_UctEwY1H7_1),.clk(gclk));
	jdff dff_A_Kc8Z5IzR5_1(.dout(w_dff_A_UctEwY1H7_1),.din(w_dff_A_Kc8Z5IzR5_1),.clk(gclk));
	jdff dff_A_XY0BUQfE6_1(.dout(w_dff_A_Kc8Z5IzR5_1),.din(w_dff_A_XY0BUQfE6_1),.clk(gclk));
	jdff dff_A_jG2qodlf0_2(.dout(w_G137_7[2]),.din(w_dff_A_jG2qodlf0_2),.clk(gclk));
	jdff dff_A_BPIqf5rI7_0(.dout(w_G137_2[0]),.din(w_dff_A_BPIqf5rI7_0),.clk(gclk));
	jdff dff_A_QWfpafDM6_0(.dout(w_dff_A_BPIqf5rI7_0),.din(w_dff_A_QWfpafDM6_0),.clk(gclk));
	jdff dff_A_bR76bPca5_1(.dout(w_G137_2[1]),.din(w_dff_A_bR76bPca5_1),.clk(gclk));
	jdff dff_A_ue7qSbSQ9_1(.dout(w_dff_A_bR76bPca5_1),.din(w_dff_A_ue7qSbSQ9_1),.clk(gclk));
	jdff dff_B_VCTn3SK60_0(.din(n1159),.dout(w_dff_B_VCTn3SK60_0),.clk(gclk));
	jdff dff_B_dm1VS66N0_0(.din(w_dff_B_VCTn3SK60_0),.dout(w_dff_B_dm1VS66N0_0),.clk(gclk));
	jdff dff_B_JCpG3cxf4_0(.din(w_dff_B_dm1VS66N0_0),.dout(w_dff_B_JCpG3cxf4_0),.clk(gclk));
	jdff dff_B_Xir8SzCa5_0(.din(w_dff_B_JCpG3cxf4_0),.dout(w_dff_B_Xir8SzCa5_0),.clk(gclk));
	jdff dff_B_gENNqRjE4_0(.din(w_dff_B_Xir8SzCa5_0),.dout(w_dff_B_gENNqRjE4_0),.clk(gclk));
	jdff dff_B_jM36jj2Z9_0(.din(w_dff_B_gENNqRjE4_0),.dout(w_dff_B_jM36jj2Z9_0),.clk(gclk));
	jdff dff_B_nADyp6BT6_0(.din(w_dff_B_jM36jj2Z9_0),.dout(w_dff_B_nADyp6BT6_0),.clk(gclk));
	jdff dff_B_3io3D0Hr7_0(.din(w_dff_B_nADyp6BT6_0),.dout(w_dff_B_3io3D0Hr7_0),.clk(gclk));
	jdff dff_B_7rEfuANi1_0(.din(w_dff_B_3io3D0Hr7_0),.dout(w_dff_B_7rEfuANi1_0),.clk(gclk));
	jdff dff_B_O1rvdU333_0(.din(w_dff_B_7rEfuANi1_0),.dout(w_dff_B_O1rvdU333_0),.clk(gclk));
	jdff dff_B_hMrZ0uPE2_0(.din(w_dff_B_O1rvdU333_0),.dout(w_dff_B_hMrZ0uPE2_0),.clk(gclk));
	jdff dff_B_uQSx3YNL7_0(.din(w_dff_B_hMrZ0uPE2_0),.dout(w_dff_B_uQSx3YNL7_0),.clk(gclk));
	jdff dff_B_MkJiLRTw9_0(.din(n1158),.dout(w_dff_B_MkJiLRTw9_0),.clk(gclk));
	jdff dff_B_FBUy87R54_2(.din(G152),.dout(w_dff_B_FBUy87R54_2),.clk(gclk));
	jdff dff_B_8QufpCzT9_2(.din(G155),.dout(w_dff_B_8QufpCzT9_2),.clk(gclk));
	jdff dff_B_4ob1Ejiw3_2(.din(w_dff_B_8QufpCzT9_2),.dout(w_dff_B_4ob1Ejiw3_2),.clk(gclk));
	jdff dff_B_7TNR61dt0_1(.din(n1153),.dout(w_dff_B_7TNR61dt0_1),.clk(gclk));
	jdff dff_B_ynkkfbZU5_1(.din(n887),.dout(w_dff_B_ynkkfbZU5_1),.clk(gclk));
	jdff dff_B_Wi5oBCgA5_1(.din(w_dff_B_ynkkfbZU5_1),.dout(w_dff_B_Wi5oBCgA5_1),.clk(gclk));
	jdff dff_B_WHUSTBAt3_1(.din(w_dff_B_Wi5oBCgA5_1),.dout(w_dff_B_WHUSTBAt3_1),.clk(gclk));
	jdff dff_B_alWXNTHX7_1(.din(w_dff_B_WHUSTBAt3_1),.dout(w_dff_B_alWXNTHX7_1),.clk(gclk));
	jdff dff_B_a6ZFEYDl6_1(.din(w_dff_B_alWXNTHX7_1),.dout(w_dff_B_a6ZFEYDl6_1),.clk(gclk));
	jdff dff_B_W9MvtiD98_1(.din(w_dff_B_a6ZFEYDl6_1),.dout(w_dff_B_W9MvtiD98_1),.clk(gclk));
	jdff dff_B_0ObkkvA53_1(.din(w_dff_B_W9MvtiD98_1),.dout(w_dff_B_0ObkkvA53_1),.clk(gclk));
	jdff dff_B_xf4nFuBp8_0(.din(n893),.dout(w_dff_B_xf4nFuBp8_0),.clk(gclk));
	jdff dff_B_D28aOgyg8_0(.din(w_dff_B_xf4nFuBp8_0),.dout(w_dff_B_D28aOgyg8_0),.clk(gclk));
	jdff dff_B_Uja55WdY4_0(.din(w_dff_B_D28aOgyg8_0),.dout(w_dff_B_Uja55WdY4_0),.clk(gclk));
	jdff dff_B_WhjvR4bw5_1(.din(n489),.dout(w_dff_B_WhjvR4bw5_1),.clk(gclk));
	jdff dff_B_RgaHLtTI8_1(.din(n484),.dout(w_dff_B_RgaHLtTI8_1),.clk(gclk));
	jdff dff_B_N46Q13tX9_1(.din(G127),.dout(w_dff_B_N46Q13tX9_1),.clk(gclk));
	jdff dff_B_TVfQ4Pp23_1(.din(w_dff_B_N46Q13tX9_1),.dout(w_dff_B_TVfQ4Pp23_1),.clk(gclk));
	jdff dff_B_d0O73iLt7_1(.din(n843),.dout(w_dff_B_d0O73iLt7_1),.clk(gclk));
	jdff dff_B_PRLkGbq50_1(.din(w_dff_B_d0O73iLt7_1),.dout(w_dff_B_PRLkGbq50_1),.clk(gclk));
	jdff dff_B_d1hn19lt3_1(.din(w_dff_B_PRLkGbq50_1),.dout(w_dff_B_d1hn19lt3_1),.clk(gclk));
	jdff dff_B_tTJAqodU4_1(.din(w_dff_B_d1hn19lt3_1),.dout(w_dff_B_tTJAqodU4_1),.clk(gclk));
	jdff dff_B_euE0zI9h3_1(.din(w_dff_B_tTJAqodU4_1),.dout(w_dff_B_euE0zI9h3_1),.clk(gclk));
	jdff dff_B_HJcQ4XXB1_1(.din(w_dff_B_euE0zI9h3_1),.dout(w_dff_B_HJcQ4XXB1_1),.clk(gclk));
	jdff dff_B_tkO5Zrls7_1(.din(w_dff_B_HJcQ4XXB1_1),.dout(w_dff_B_tkO5Zrls7_1),.clk(gclk));
	jdff dff_B_0m77Vsxo6_1(.din(n844),.dout(w_dff_B_0m77Vsxo6_1),.clk(gclk));
	jdff dff_B_j0sHRqff0_1(.din(w_dff_B_0m77Vsxo6_1),.dout(w_dff_B_j0sHRqff0_1),.clk(gclk));
	jdff dff_B_bdLFoM7E2_1(.din(w_dff_B_j0sHRqff0_1),.dout(w_dff_B_bdLFoM7E2_1),.clk(gclk));
	jdff dff_B_g0gNCxJa4_1(.din(w_dff_B_bdLFoM7E2_1),.dout(w_dff_B_g0gNCxJa4_1),.clk(gclk));
	jdff dff_A_KIDJxiBf7_0(.dout(w_n847_0[0]),.din(w_dff_A_KIDJxiBf7_0),.clk(gclk));
	jdff dff_A_3cKzkmaC5_0(.dout(w_dff_A_KIDJxiBf7_0),.din(w_dff_A_3cKzkmaC5_0),.clk(gclk));
	jdff dff_A_Sdx6V3Sz3_0(.dout(w_dff_A_3cKzkmaC5_0),.din(w_dff_A_Sdx6V3Sz3_0),.clk(gclk));
	jdff dff_A_D0Gyjluq5_0(.dout(w_dff_A_Sdx6V3Sz3_0),.din(w_dff_A_D0Gyjluq5_0),.clk(gclk));
	jdff dff_A_SJ5wKky19_0(.dout(w_dff_A_D0Gyjluq5_0),.din(w_dff_A_SJ5wKky19_0),.clk(gclk));
	jdff dff_B_a2IDp3261_1(.din(n393),.dout(w_dff_B_a2IDp3261_1),.clk(gclk));
	jdff dff_B_U9XiRrDq4_1(.din(n388),.dout(w_dff_B_U9XiRrDq4_1),.clk(gclk));
	jdff dff_B_s5MMWwXL4_1(.din(G119),.dout(w_dff_B_s5MMWwXL4_1),.clk(gclk));
	jdff dff_B_YHnInmKb8_1(.din(w_dff_B_s5MMWwXL4_1),.dout(w_dff_B_YHnInmKb8_1),.clk(gclk));
	jdff dff_B_iO59QYdP1_0(.din(n1168),.dout(w_dff_B_iO59QYdP1_0),.clk(gclk));
	jdff dff_B_UI3T1w9Q6_0(.din(w_dff_B_iO59QYdP1_0),.dout(w_dff_B_UI3T1w9Q6_0),.clk(gclk));
	jdff dff_B_IyXndkve0_0(.din(w_dff_B_UI3T1w9Q6_0),.dout(w_dff_B_IyXndkve0_0),.clk(gclk));
	jdff dff_B_lbZteEbc9_0(.din(w_dff_B_IyXndkve0_0),.dout(w_dff_B_lbZteEbc9_0),.clk(gclk));
	jdff dff_B_LKoMlFcM0_0(.din(w_dff_B_lbZteEbc9_0),.dout(w_dff_B_LKoMlFcM0_0),.clk(gclk));
	jdff dff_B_MALlDwj99_0(.din(w_dff_B_LKoMlFcM0_0),.dout(w_dff_B_MALlDwj99_0),.clk(gclk));
	jdff dff_B_wjbyFsUv4_0(.din(w_dff_B_MALlDwj99_0),.dout(w_dff_B_wjbyFsUv4_0),.clk(gclk));
	jdff dff_B_H1JCgz9B3_0(.din(w_dff_B_wjbyFsUv4_0),.dout(w_dff_B_H1JCgz9B3_0),.clk(gclk));
	jdff dff_B_rJO1WmZA8_0(.din(w_dff_B_H1JCgz9B3_0),.dout(w_dff_B_rJO1WmZA8_0),.clk(gclk));
	jdff dff_B_qeF7S8Vs7_0(.din(w_dff_B_rJO1WmZA8_0),.dout(w_dff_B_qeF7S8Vs7_0),.clk(gclk));
	jdff dff_B_ILLp9iLJ9_0(.din(w_dff_B_qeF7S8Vs7_0),.dout(w_dff_B_ILLp9iLJ9_0),.clk(gclk));
	jdff dff_B_Hr3vt8wg1_0(.din(w_dff_B_ILLp9iLJ9_0),.dout(w_dff_B_Hr3vt8wg1_0),.clk(gclk));
	jdff dff_B_OTqproJZ7_0(.din(w_dff_B_Hr3vt8wg1_0),.dout(w_dff_B_OTqproJZ7_0),.clk(gclk));
	jdff dff_B_sFIvMDpm4_0(.din(n1167),.dout(w_dff_B_sFIvMDpm4_0),.clk(gclk));
	jdff dff_B_C5Gn2Iqp1_2(.din(G146),.dout(w_dff_B_C5Gn2Iqp1_2),.clk(gclk));
	jdff dff_B_8LJWb9wq6_2(.din(G149),.dout(w_dff_B_8LJWb9wq6_2),.clk(gclk));
	jdff dff_B_4NUXgw828_2(.din(w_dff_B_8LJWb9wq6_2),.dout(w_dff_B_4NUXgw828_2),.clk(gclk));
	jdff dff_B_lpCaWUUQ1_1(.din(n878),.dout(w_dff_B_lpCaWUUQ1_1),.clk(gclk));
	jdff dff_B_GOhy5pRA2_1(.din(w_dff_B_lpCaWUUQ1_1),.dout(w_dff_B_GOhy5pRA2_1),.clk(gclk));
	jdff dff_B_rsoI9LAR9_1(.din(w_dff_B_GOhy5pRA2_1),.dout(w_dff_B_rsoI9LAR9_1),.clk(gclk));
	jdff dff_B_pnfwq5m68_1(.din(w_dff_B_rsoI9LAR9_1),.dout(w_dff_B_pnfwq5m68_1),.clk(gclk));
	jdff dff_B_tvhdN1lp1_1(.din(w_dff_B_pnfwq5m68_1),.dout(w_dff_B_tvhdN1lp1_1),.clk(gclk));
	jdff dff_B_DjSPTOBr9_1(.din(w_dff_B_tvhdN1lp1_1),.dout(w_dff_B_DjSPTOBr9_1),.clk(gclk));
	jdff dff_B_0h2uZ0XB6_1(.din(w_dff_B_DjSPTOBr9_1),.dout(w_dff_B_0h2uZ0XB6_1),.clk(gclk));
	jdff dff_B_nuJyNRVB7_1(.din(w_dff_B_0h2uZ0XB6_1),.dout(w_dff_B_nuJyNRVB7_1),.clk(gclk));
	jdff dff_B_uUyw6SBA8_0(.din(n883),.dout(w_dff_B_uUyw6SBA8_0),.clk(gclk));
	jdff dff_B_0i0gv2C88_0(.din(w_dff_B_uUyw6SBA8_0),.dout(w_dff_B_0i0gv2C88_0),.clk(gclk));
	jdff dff_B_3Fv80fzf9_0(.din(w_dff_B_0i0gv2C88_0),.dout(w_dff_B_3Fv80fzf9_0),.clk(gclk));
	jdff dff_B_V3cGInGs1_0(.din(w_dff_B_3Fv80fzf9_0),.dout(w_dff_B_V3cGInGs1_0),.clk(gclk));
	jdff dff_B_zOGq44EE9_1(.din(n524),.dout(w_dff_B_zOGq44EE9_1),.clk(gclk));
	jdff dff_B_XsWxfEym6_1(.din(n519),.dout(w_dff_B_XsWxfEym6_1),.clk(gclk));
	jdff dff_A_eP7Rd7X16_2(.dout(w_G4092_7[2]),.din(w_dff_A_eP7Rd7X16_2),.clk(gclk));
	jdff dff_A_VfKayZhp7_2(.dout(w_dff_A_eP7Rd7X16_2),.din(w_dff_A_VfKayZhp7_2),.clk(gclk));
	jdff dff_A_HTohEeBT0_2(.dout(w_dff_A_VfKayZhp7_2),.din(w_dff_A_HTohEeBT0_2),.clk(gclk));
	jdff dff_A_F0JhapCz1_0(.dout(w_n880_0[0]),.din(w_dff_A_F0JhapCz1_0),.clk(gclk));
	jdff dff_A_uKOnJYMr6_0(.dout(w_dff_A_F0JhapCz1_0),.din(w_dff_A_uKOnJYMr6_0),.clk(gclk));
	jdff dff_A_hJYd0ebg5_0(.dout(w_dff_A_uKOnJYMr6_0),.din(w_dff_A_hJYd0ebg5_0),.clk(gclk));
	jdff dff_A_ALOmsiws4_0(.dout(w_dff_A_hJYd0ebg5_0),.din(w_dff_A_ALOmsiws4_0),.clk(gclk));
	jdff dff_A_cxXdvzs87_0(.dout(w_dff_A_ALOmsiws4_0),.din(w_dff_A_cxXdvzs87_0),.clk(gclk));
	jdff dff_A_IkAbCPM81_1(.dout(w_G4091_3[1]),.din(w_dff_A_IkAbCPM81_1),.clk(gclk));
	jdff dff_A_iToMPgUv9_2(.dout(w_G4091_3[2]),.din(w_dff_A_iToMPgUv9_2),.clk(gclk));
	jdff dff_A_wM42BPhe6_2(.dout(w_dff_A_iToMPgUv9_2),.din(w_dff_A_wM42BPhe6_2),.clk(gclk));
	jdff dff_B_wNUOId764_1(.din(G128),.dout(w_dff_B_wNUOId764_1),.clk(gclk));
	jdff dff_B_ztXtA0sx5_1(.din(w_dff_B_wNUOId764_1),.dout(w_dff_B_ztXtA0sx5_1),.clk(gclk));
	jdff dff_A_MwqBT1ch8_0(.dout(w_n1008_3[0]),.din(w_dff_A_MwqBT1ch8_0),.clk(gclk));
	jdff dff_A_TFA1s4mL4_0(.dout(w_dff_A_MwqBT1ch8_0),.din(w_dff_A_TFA1s4mL4_0),.clk(gclk));
	jdff dff_A_2hbXSAaW4_1(.dout(w_n1008_3[1]),.din(w_dff_A_2hbXSAaW4_1),.clk(gclk));
	jdff dff_B_ef1jqy0p4_1(.din(n834),.dout(w_dff_B_ef1jqy0p4_1),.clk(gclk));
	jdff dff_B_eUK8pFhK0_1(.din(w_dff_B_ef1jqy0p4_1),.dout(w_dff_B_eUK8pFhK0_1),.clk(gclk));
	jdff dff_B_cpJWD3be5_1(.din(w_dff_B_eUK8pFhK0_1),.dout(w_dff_B_cpJWD3be5_1),.clk(gclk));
	jdff dff_B_nHlm3X4o6_1(.din(w_dff_B_cpJWD3be5_1),.dout(w_dff_B_nHlm3X4o6_1),.clk(gclk));
	jdff dff_B_o6Hv4IOT0_1(.din(w_dff_B_nHlm3X4o6_1),.dout(w_dff_B_o6Hv4IOT0_1),.clk(gclk));
	jdff dff_B_upyi4HYX0_1(.din(w_dff_B_o6Hv4IOT0_1),.dout(w_dff_B_upyi4HYX0_1),.clk(gclk));
	jdff dff_B_2GZjt7VG3_1(.din(w_dff_B_upyi4HYX0_1),.dout(w_dff_B_2GZjt7VG3_1),.clk(gclk));
	jdff dff_B_gaJd1ReL8_1(.din(w_dff_B_2GZjt7VG3_1),.dout(w_dff_B_gaJd1ReL8_1),.clk(gclk));
	jdff dff_B_Kz64QH1X3_1(.din(w_dff_B_gaJd1ReL8_1),.dout(w_dff_B_Kz64QH1X3_1),.clk(gclk));
	jdff dff_B_91QUffPM9_0(.din(n839),.dout(w_dff_B_91QUffPM9_0),.clk(gclk));
	jdff dff_B_yTyBLB759_0(.din(w_dff_B_91QUffPM9_0),.dout(w_dff_B_yTyBLB759_0),.clk(gclk));
	jdff dff_B_cbCql3jt1_0(.din(w_dff_B_yTyBLB759_0),.dout(w_dff_B_cbCql3jt1_0),.clk(gclk));
	jdff dff_B_b3x1WAc13_0(.din(w_dff_B_cbCql3jt1_0),.dout(w_dff_B_b3x1WAc13_0),.clk(gclk));
	jdff dff_B_vl6j40Uh3_0(.din(w_dff_B_b3x1WAc13_0),.dout(w_dff_B_vl6j40Uh3_0),.clk(gclk));
	jdff dff_B_ztQca1h34_0(.din(w_dff_B_vl6j40Uh3_0),.dout(w_dff_B_ztQca1h34_0),.clk(gclk));
	jdff dff_B_ub1rWXPF9_1(.din(n360),.dout(w_dff_B_ub1rWXPF9_1),.clk(gclk));
	jdff dff_A_09RYPLEY5_0(.dout(w_n749_11[0]),.din(w_dff_A_09RYPLEY5_0),.clk(gclk));
	jdff dff_A_NVDs0d1O7_1(.dout(w_n749_11[1]),.din(w_dff_A_NVDs0d1O7_1),.clk(gclk));
	jdff dff_A_UPMtDmzk0_0(.dout(w_n749_3[0]),.din(w_dff_A_UPMtDmzk0_0),.clk(gclk));
	jdff dff_A_NexaASTY3_2(.dout(w_n749_3[2]),.din(w_dff_A_NexaASTY3_2),.clk(gclk));
	jdff dff_A_AnjC0Ijo8_1(.dout(w_G4092_8[1]),.din(w_dff_A_AnjC0Ijo8_1),.clk(gclk));
	jdff dff_A_SwxSWY5E6_2(.dout(w_G4092_8[2]),.din(w_dff_A_SwxSWY5E6_2),.clk(gclk));
	jdff dff_A_XuWp6dEZ8_0(.dout(w_n836_0[0]),.din(w_dff_A_XuWp6dEZ8_0),.clk(gclk));
	jdff dff_A_K6H9YeB14_0(.dout(w_dff_A_XuWp6dEZ8_0),.din(w_dff_A_K6H9YeB14_0),.clk(gclk));
	jdff dff_A_I3fQUKHa0_0(.dout(w_dff_A_K6H9YeB14_0),.din(w_dff_A_I3fQUKHa0_0),.clk(gclk));
	jdff dff_A_IqMxCBZb8_0(.dout(w_dff_A_I3fQUKHa0_0),.din(w_dff_A_IqMxCBZb8_0),.clk(gclk));
	jdff dff_A_PNbiSLXZ2_0(.dout(w_dff_A_IqMxCBZb8_0),.din(w_dff_A_PNbiSLXZ2_0),.clk(gclk));
	jdff dff_A_GQD2edxX0_0(.dout(w_dff_A_PNbiSLXZ2_0),.din(w_dff_A_GQD2edxX0_0),.clk(gclk));
	jdff dff_A_XA3HZLVg6_0(.dout(w_dff_A_GQD2edxX0_0),.din(w_dff_A_XA3HZLVg6_0),.clk(gclk));
	jdff dff_A_SuK89Nxe8_1(.dout(w_n753_0[1]),.din(w_dff_A_SuK89Nxe8_1),.clk(gclk));
	jdff dff_A_DaXJgAHl0_1(.dout(w_dff_A_SuK89Nxe8_1),.din(w_dff_A_DaXJgAHl0_1),.clk(gclk));
	jdff dff_A_LTAqX0I66_2(.dout(w_n753_0[2]),.din(w_dff_A_LTAqX0I66_2),.clk(gclk));
	jdff dff_A_HiMulCm28_2(.dout(w_dff_A_LTAqX0I66_2),.din(w_dff_A_HiMulCm28_2),.clk(gclk));
	jdff dff_A_QgVLGpdo9_2(.dout(w_dff_A_HiMulCm28_2),.din(w_dff_A_QgVLGpdo9_2),.clk(gclk));
	jdff dff_A_oF8Rkg9O6_2(.dout(w_dff_A_QgVLGpdo9_2),.din(w_dff_A_oF8Rkg9O6_2),.clk(gclk));
	jdff dff_A_v65CWJYg0_2(.dout(w_dff_A_oF8Rkg9O6_2),.din(w_dff_A_v65CWJYg0_2),.clk(gclk));
	jdff dff_B_p4Mf3qHF5_3(.din(n753),.dout(w_dff_B_p4Mf3qHF5_3),.clk(gclk));
	jdff dff_B_eHIEZXIz1_3(.din(w_dff_B_p4Mf3qHF5_3),.dout(w_dff_B_eHIEZXIz1_3),.clk(gclk));
	jdff dff_A_64uspizJ6_0(.dout(w_G4091_4[0]),.din(w_dff_A_64uspizJ6_0),.clk(gclk));
	jdff dff_A_e4xWmsaF2_0(.dout(w_dff_A_64uspizJ6_0),.din(w_dff_A_e4xWmsaF2_0),.clk(gclk));
	jdff dff_A_HcMG7EVG3_0(.dout(w_dff_A_e4xWmsaF2_0),.din(w_dff_A_HcMG7EVG3_0),.clk(gclk));
	jdff dff_A_NGs4s4Vo9_0(.dout(w_dff_A_HcMG7EVG3_0),.din(w_dff_A_NGs4s4Vo9_0),.clk(gclk));
	jdff dff_A_8F6JTJkA8_2(.dout(w_G4091_4[2]),.din(w_dff_A_8F6JTJkA8_2),.clk(gclk));
	jdff dff_A_VFM07rhN7_2(.dout(w_dff_A_8F6JTJkA8_2),.din(w_dff_A_VFM07rhN7_2),.clk(gclk));
	jdff dff_A_jFYyJij92_2(.dout(w_dff_A_VFM07rhN7_2),.din(w_dff_A_jFYyJij92_2),.clk(gclk));
	jdff dff_B_FQ5DCCzZ8_1(.din(G130),.dout(w_dff_B_FQ5DCCzZ8_1),.clk(gclk));
	jdff dff_B_JVMS83W53_1(.din(w_dff_B_FQ5DCCzZ8_1),.dout(w_dff_B_JVMS83W53_1),.clk(gclk));
	jdff dff_B_878hfwhA2_1(.din(n1173),.dout(w_dff_B_878hfwhA2_1),.clk(gclk));
	jdff dff_B_dlQcxcXw5_1(.din(w_dff_B_878hfwhA2_1),.dout(w_dff_B_dlQcxcXw5_1),.clk(gclk));
	jdff dff_B_ggkqwLvQ9_1(.din(w_dff_B_dlQcxcXw5_1),.dout(w_dff_B_ggkqwLvQ9_1),.clk(gclk));
	jdff dff_B_BuYMsqKl6_1(.din(w_dff_B_ggkqwLvQ9_1),.dout(w_dff_B_BuYMsqKl6_1),.clk(gclk));
	jdff dff_B_xX9dfFky5_1(.din(w_dff_B_BuYMsqKl6_1),.dout(w_dff_B_xX9dfFky5_1),.clk(gclk));
	jdff dff_B_a8L4tgbd2_1(.din(w_dff_B_xX9dfFky5_1),.dout(w_dff_B_a8L4tgbd2_1),.clk(gclk));
	jdff dff_B_Q2chBNhn7_1(.din(w_dff_B_a8L4tgbd2_1),.dout(w_dff_B_Q2chBNhn7_1),.clk(gclk));
	jdff dff_B_HcL4UfEc1_1(.din(w_dff_B_Q2chBNhn7_1),.dout(w_dff_B_HcL4UfEc1_1),.clk(gclk));
	jdff dff_B_90w1LJGs7_1(.din(w_dff_B_HcL4UfEc1_1),.dout(w_dff_B_90w1LJGs7_1),.clk(gclk));
	jdff dff_B_rtwK8WQK2_1(.din(w_dff_B_90w1LJGs7_1),.dout(w_dff_B_rtwK8WQK2_1),.clk(gclk));
	jdff dff_B_Cp5HUqhv1_1(.din(w_dff_B_rtwK8WQK2_1),.dout(w_dff_B_Cp5HUqhv1_1),.clk(gclk));
	jdff dff_B_awR0QHK92_1(.din(w_dff_B_Cp5HUqhv1_1),.dout(w_dff_B_awR0QHK92_1),.clk(gclk));
	jdff dff_B_NukNxX8y4_1(.din(w_dff_B_awR0QHK92_1),.dout(w_dff_B_NukNxX8y4_1),.clk(gclk));
	jdff dff_B_O7Wf56j41_1(.din(w_dff_B_NukNxX8y4_1),.dout(w_dff_B_O7Wf56j41_1),.clk(gclk));
	jdff dff_B_yFj93FxD3_1(.din(w_dff_B_O7Wf56j41_1),.dout(w_dff_B_yFj93FxD3_1),.clk(gclk));
	jdff dff_B_X4t6qNE25_1(.din(w_dff_B_yFj93FxD3_1),.dout(w_dff_B_X4t6qNE25_1),.clk(gclk));
	jdff dff_B_MBTv1AYc8_1(.din(w_dff_B_X4t6qNE25_1),.dout(w_dff_B_MBTv1AYc8_1),.clk(gclk));
	jdff dff_B_QSIfbudR1_1(.din(w_dff_B_MBTv1AYc8_1),.dout(w_dff_B_QSIfbudR1_1),.clk(gclk));
	jdff dff_B_IvTs3Xyw0_1(.din(n1182),.dout(w_dff_B_IvTs3Xyw0_1),.clk(gclk));
	jdff dff_B_aUrDXous6_1(.din(w_dff_B_IvTs3Xyw0_1),.dout(w_dff_B_aUrDXous6_1),.clk(gclk));
	jdff dff_B_h2Z1q8qw5_1(.din(w_dff_B_aUrDXous6_1),.dout(w_dff_B_h2Z1q8qw5_1),.clk(gclk));
	jdff dff_B_l2bDNCRO1_1(.din(w_dff_B_h2Z1q8qw5_1),.dout(w_dff_B_l2bDNCRO1_1),.clk(gclk));
	jdff dff_B_74DlTyWW2_1(.din(w_dff_B_l2bDNCRO1_1),.dout(w_dff_B_74DlTyWW2_1),.clk(gclk));
	jdff dff_B_GwvYsTUa7_1(.din(w_dff_B_74DlTyWW2_1),.dout(w_dff_B_GwvYsTUa7_1),.clk(gclk));
	jdff dff_B_PmqqNJOO4_1(.din(w_dff_B_GwvYsTUa7_1),.dout(w_dff_B_PmqqNJOO4_1),.clk(gclk));
	jdff dff_B_pJUAKFgW4_1(.din(w_dff_B_PmqqNJOO4_1),.dout(w_dff_B_pJUAKFgW4_1),.clk(gclk));
	jdff dff_B_iXjaPqPW3_1(.din(w_dff_B_pJUAKFgW4_1),.dout(w_dff_B_iXjaPqPW3_1),.clk(gclk));
	jdff dff_B_JEENBjMl8_1(.din(w_dff_B_iXjaPqPW3_1),.dout(w_dff_B_JEENBjMl8_1),.clk(gclk));
	jdff dff_B_okZtuIBU5_0(.din(n1185),.dout(w_dff_B_okZtuIBU5_0),.clk(gclk));
	jdff dff_B_34JMfYHQ5_0(.din(w_dff_B_okZtuIBU5_0),.dout(w_dff_B_34JMfYHQ5_0),.clk(gclk));
	jdff dff_B_r0ShhH3K0_0(.din(w_dff_B_34JMfYHQ5_0),.dout(w_dff_B_r0ShhH3K0_0),.clk(gclk));
	jdff dff_B_00tyfqLR7_0(.din(w_dff_B_r0ShhH3K0_0),.dout(w_dff_B_00tyfqLR7_0),.clk(gclk));
	jdff dff_B_1QfqCUSw9_0(.din(w_dff_B_00tyfqLR7_0),.dout(w_dff_B_1QfqCUSw9_0),.clk(gclk));
	jdff dff_B_0ULmIPpw8_0(.din(w_dff_B_1QfqCUSw9_0),.dout(w_dff_B_0ULmIPpw8_0),.clk(gclk));
	jdff dff_B_6A3aoKRn7_0(.din(w_dff_B_0ULmIPpw8_0),.dout(w_dff_B_6A3aoKRn7_0),.clk(gclk));
	jdff dff_B_nxRAlrok4_0(.din(w_dff_B_6A3aoKRn7_0),.dout(w_dff_B_nxRAlrok4_0),.clk(gclk));
	jdff dff_B_plC7k5TJ0_0(.din(w_dff_B_nxRAlrok4_0),.dout(w_dff_B_plC7k5TJ0_0),.clk(gclk));
	jdff dff_B_eLQDXY4u6_0(.din(w_dff_B_plC7k5TJ0_0),.dout(w_dff_B_eLQDXY4u6_0),.clk(gclk));
	jdff dff_B_dTppWHvb1_0(.din(w_dff_B_eLQDXY4u6_0),.dout(w_dff_B_dTppWHvb1_0),.clk(gclk));
	jdff dff_B_5qe7dsnQ1_0(.din(w_dff_B_dTppWHvb1_0),.dout(w_dff_B_5qe7dsnQ1_0),.clk(gclk));
	jdff dff_B_zflnnlws8_0(.din(w_dff_B_5qe7dsnQ1_0),.dout(w_dff_B_zflnnlws8_0),.clk(gclk));
	jdff dff_B_I71IC8ty2_0(.din(w_dff_B_zflnnlws8_0),.dout(w_dff_B_I71IC8ty2_0),.clk(gclk));
	jdff dff_B_2D6IMdj80_0(.din(w_dff_B_I71IC8ty2_0),.dout(w_dff_B_2D6IMdj80_0),.clk(gclk));
	jdff dff_B_VYAmWsj55_0(.din(w_dff_B_2D6IMdj80_0),.dout(w_dff_B_VYAmWsj55_0),.clk(gclk));
	jdff dff_B_JnpBMWfr7_1(.din(n1175),.dout(w_dff_B_JnpBMWfr7_1),.clk(gclk));
	jdff dff_B_Kh4VdNXQ4_1(.din(w_dff_B_JnpBMWfr7_1),.dout(w_dff_B_Kh4VdNXQ4_1),.clk(gclk));
	jdff dff_B_GPiIhynG4_1(.din(w_dff_B_Kh4VdNXQ4_1),.dout(w_dff_B_GPiIhynG4_1),.clk(gclk));
	jdff dff_B_TllRHp4q3_1(.din(n1176),.dout(w_dff_B_TllRHp4q3_1),.clk(gclk));
	jdff dff_B_sUH7TDOi9_1(.din(w_dff_B_TllRHp4q3_1),.dout(w_dff_B_sUH7TDOi9_1),.clk(gclk));
	jdff dff_B_uaRH0Okv8_1(.din(w_dff_B_sUH7TDOi9_1),.dout(w_dff_B_uaRH0Okv8_1),.clk(gclk));
	jdff dff_B_mFXIpEUa0_1(.din(w_dff_B_uaRH0Okv8_1),.dout(w_dff_B_mFXIpEUa0_1),.clk(gclk));
	jdff dff_B_mx8dEiB92_1(.din(w_dff_B_mFXIpEUa0_1),.dout(w_dff_B_mx8dEiB92_1),.clk(gclk));
	jdff dff_B_NEaFt02s3_1(.din(w_dff_B_mx8dEiB92_1),.dout(w_dff_B_NEaFt02s3_1),.clk(gclk));
	jdff dff_A_5zUNvNBm9_0(.dout(w_n1177_0[0]),.din(w_dff_A_5zUNvNBm9_0),.clk(gclk));
	jdff dff_A_mRIEnLgl0_0(.dout(w_dff_A_5zUNvNBm9_0),.din(w_dff_A_mRIEnLgl0_0),.clk(gclk));
	jdff dff_A_U72sNUkJ6_0(.dout(w_dff_A_mRIEnLgl0_0),.din(w_dff_A_U72sNUkJ6_0),.clk(gclk));
	jdff dff_A_8BHfggQZ0_0(.dout(w_dff_A_U72sNUkJ6_0),.din(w_dff_A_8BHfggQZ0_0),.clk(gclk));
	jdff dff_A_Fo2Mv4J16_0(.dout(w_dff_A_8BHfggQZ0_0),.din(w_dff_A_Fo2Mv4J16_0),.clk(gclk));
	jdff dff_A_fcTc6bFA7_0(.dout(w_dff_A_Fo2Mv4J16_0),.din(w_dff_A_fcTc6bFA7_0),.clk(gclk));
	jdff dff_A_2egfg4Gc8_0(.dout(w_dff_A_fcTc6bFA7_0),.din(w_dff_A_2egfg4Gc8_0),.clk(gclk));
	jdff dff_A_Twjnsnti9_0(.dout(w_dff_A_2egfg4Gc8_0),.din(w_dff_A_Twjnsnti9_0),.clk(gclk));
	jdff dff_A_swfVtjcd7_0(.dout(w_dff_A_Twjnsnti9_0),.din(w_dff_A_swfVtjcd7_0),.clk(gclk));
	jdff dff_A_oT4WLw3O6_0(.dout(w_dff_A_swfVtjcd7_0),.din(w_dff_A_oT4WLw3O6_0),.clk(gclk));
	jdff dff_A_ICC9pbgr6_0(.dout(w_dff_A_oT4WLw3O6_0),.din(w_dff_A_ICC9pbgr6_0),.clk(gclk));
	jdff dff_B_Q6fkFxpj8_2(.din(n1177),.dout(w_dff_B_Q6fkFxpj8_2),.clk(gclk));
	jdff dff_B_8LUOjPoT0_2(.din(w_dff_B_Q6fkFxpj8_2),.dout(w_dff_B_8LUOjPoT0_2),.clk(gclk));
	jdff dff_B_aEjRTtTd9_2(.din(w_dff_B_8LUOjPoT0_2),.dout(w_dff_B_aEjRTtTd9_2),.clk(gclk));
	jdff dff_B_ZpVN6DKC2_2(.din(w_dff_B_aEjRTtTd9_2),.dout(w_dff_B_ZpVN6DKC2_2),.clk(gclk));
	jdff dff_B_cYBHEi6R0_2(.din(w_dff_B_ZpVN6DKC2_2),.dout(w_dff_B_cYBHEi6R0_2),.clk(gclk));
	jdff dff_A_5ks2fcuz9_0(.dout(w_G3717_0[0]),.din(w_dff_A_5ks2fcuz9_0),.clk(gclk));
	jdff dff_A_5EHyocmY4_1(.dout(w_n428_1[1]),.din(w_dff_A_5EHyocmY4_1),.clk(gclk));
	jdff dff_A_kfchUDvm4_2(.dout(w_G3724_0[2]),.din(w_dff_A_kfchUDvm4_2),.clk(gclk));
	jdff dff_A_2Q8Xhje30_2(.dout(w_dff_A_kfchUDvm4_2),.din(w_dff_A_2Q8Xhje30_2),.clk(gclk));
	jdff dff_A_ZCsVAV2w1_2(.dout(w_dff_A_2Q8Xhje30_2),.din(w_dff_A_ZCsVAV2w1_2),.clk(gclk));
	jdff dff_A_dOM0HN591_2(.dout(w_dff_A_ZCsVAV2w1_2),.din(w_dff_A_dOM0HN591_2),.clk(gclk));
	jdff dff_A_n00IHA5k6_0(.dout(w_n1179_0[0]),.din(w_dff_A_n00IHA5k6_0),.clk(gclk));
	jdff dff_A_49KHGlqX7_0(.dout(w_dff_A_n00IHA5k6_0),.din(w_dff_A_49KHGlqX7_0),.clk(gclk));
	jdff dff_A_7TSw0oRm8_0(.dout(w_dff_A_49KHGlqX7_0),.din(w_dff_A_7TSw0oRm8_0),.clk(gclk));
	jdff dff_A_nFLcoEgD4_0(.dout(w_dff_A_7TSw0oRm8_0),.din(w_dff_A_nFLcoEgD4_0),.clk(gclk));
	jdff dff_A_kMujjOwz8_0(.dout(w_dff_A_nFLcoEgD4_0),.din(w_dff_A_kMujjOwz8_0),.clk(gclk));
	jdff dff_A_XV3EmB432_0(.dout(w_dff_A_kMujjOwz8_0),.din(w_dff_A_XV3EmB432_0),.clk(gclk));
	jdff dff_A_xpomOwAB9_0(.dout(w_dff_A_XV3EmB432_0),.din(w_dff_A_xpomOwAB9_0),.clk(gclk));
	jdff dff_A_Ac50fvil1_0(.dout(w_dff_A_xpomOwAB9_0),.din(w_dff_A_Ac50fvil1_0),.clk(gclk));
	jdff dff_A_1Lp7pGEt9_0(.dout(w_dff_A_Ac50fvil1_0),.din(w_dff_A_1Lp7pGEt9_0),.clk(gclk));
	jdff dff_A_zOiOBzm24_0(.dout(w_dff_A_1Lp7pGEt9_0),.din(w_dff_A_zOiOBzm24_0),.clk(gclk));
	jdff dff_A_vXobmQJ75_0(.dout(w_dff_A_zOiOBzm24_0),.din(w_dff_A_vXobmQJ75_0),.clk(gclk));
	jdff dff_B_cD0jNOOq0_1(.din(G132),.dout(w_dff_B_cD0jNOOq0_1),.clk(gclk));
	jdff dff_B_bwUTDkPc2_1(.din(w_dff_B_cD0jNOOq0_1),.dout(w_dff_B_bwUTDkPc2_1),.clk(gclk));
	jdff dff_B_uu0kXH8T2_1(.din(w_dff_B_bwUTDkPc2_1),.dout(w_dff_B_uu0kXH8T2_1),.clk(gclk));
	jdff dff_B_sGovDXq85_1(.din(w_dff_B_uu0kXH8T2_1),.dout(w_dff_B_sGovDXq85_1),.clk(gclk));
	jdff dff_B_MvEi3CGB6_1(.din(n1223),.dout(w_dff_B_MvEi3CGB6_1),.clk(gclk));
	jdff dff_B_103t0hcc7_0(.din(n1227),.dout(w_dff_B_103t0hcc7_0),.clk(gclk));
	jdff dff_B_Kz98kc4B3_0(.din(w_dff_B_103t0hcc7_0),.dout(w_dff_B_Kz98kc4B3_0),.clk(gclk));
	jdff dff_B_YG7YJKWX4_0(.din(w_dff_B_Kz98kc4B3_0),.dout(w_dff_B_YG7YJKWX4_0),.clk(gclk));
	jdff dff_B_7QKpzjzx6_0(.din(w_dff_B_YG7YJKWX4_0),.dout(w_dff_B_7QKpzjzx6_0),.clk(gclk));
	jdff dff_B_Mbqsu6jf8_0(.din(n1226),.dout(w_dff_B_Mbqsu6jf8_0),.clk(gclk));
	jdff dff_A_Ujmf1NMl0_0(.dout(w_G559_0[0]),.din(w_dff_A_Ujmf1NMl0_0),.clk(gclk));
	jdff dff_A_3Ccg3jVJ7_0(.dout(w_dff_A_Ujmf1NMl0_0),.din(w_dff_A_3Ccg3jVJ7_0),.clk(gclk));
	jdff dff_B_hpGPWnPQ3_0(.din(n668),.dout(w_dff_B_hpGPWnPQ3_0),.clk(gclk));
	jdff dff_B_cWFmm0rY8_1(.din(n663),.dout(w_dff_B_cWFmm0rY8_1),.clk(gclk));
	jdff dff_B_NKzmPQCu8_1(.din(n916),.dout(w_dff_B_NKzmPQCu8_1),.clk(gclk));
	jdff dff_B_ZGC8ArjM6_1(.din(n917),.dout(w_dff_B_ZGC8ArjM6_1),.clk(gclk));
	jdff dff_B_jYQ8yJpf9_0(.din(n915),.dout(w_dff_B_jYQ8yJpf9_0),.clk(gclk));
	jdff dff_B_6nFQBuEi0_1(.din(n913),.dout(w_dff_B_6nFQBuEi0_1),.clk(gclk));
	jdff dff_B_WrvP5RP93_0(.din(G372),.dout(w_dff_B_WrvP5RP93_0),.clk(gclk));
	jdff dff_B_wEjuJzkp5_1(.din(n909),.dout(w_dff_B_wEjuJzkp5_1),.clk(gclk));
	jdff dff_B_YWgJBZQO1_1(.din(n907),.dout(w_dff_B_YWgJBZQO1_1),.clk(gclk));
	jdff dff_B_l0ah2yuI1_1(.din(w_dff_B_YWgJBZQO1_1),.dout(w_dff_B_l0ah2yuI1_1),.clk(gclk));
	jdff dff_B_j2Xx3lIg6_0(.din(n1222),.dout(w_dff_B_j2Xx3lIg6_0),.clk(gclk));
	jdff dff_B_8wHB2uIa9_0(.din(w_dff_B_j2Xx3lIg6_0),.dout(w_dff_B_8wHB2uIa9_0),.clk(gclk));
	jdff dff_B_MvMuVnvU9_0(.din(w_dff_B_8wHB2uIa9_0),.dout(w_dff_B_MvMuVnvU9_0),.clk(gclk));
	jdff dff_B_i4RxXwLI4_0(.din(n678),.dout(w_dff_B_i4RxXwLI4_0),.clk(gclk));
	jdff dff_B_xUTfXL7O8_1(.din(n672),.dout(w_dff_B_xUTfXL7O8_1),.clk(gclk));
	jdff dff_A_ffeh8EW72_0(.dout(w_G245_0[0]),.din(w_dff_A_ffeh8EW72_0),.clk(gclk));
	jdff dff_A_HThBUF9J9_0(.dout(w_dff_A_ffeh8EW72_0),.din(w_dff_A_HThBUF9J9_0),.clk(gclk));
	jdff dff_A_xQepA7lE2_0(.dout(w_dff_A_HThBUF9J9_0),.din(w_dff_A_xQepA7lE2_0),.clk(gclk));
	jdff dff_A_TUtlYu8p7_0(.dout(w_dff_A_xQepA7lE2_0),.din(w_dff_A_TUtlYu8p7_0),.clk(gclk));
	jdff dff_B_SIK51O1X2_1(.din(n926),.dout(w_dff_B_SIK51O1X2_1),.clk(gclk));
	jdff dff_B_QMRvX1Xm5_1(.din(n930),.dout(w_dff_B_QMRvX1Xm5_1),.clk(gclk));
	jdff dff_B_5BGTfmIR1_1(.din(w_dff_B_QMRvX1Xm5_1),.dout(w_dff_B_5BGTfmIR1_1),.clk(gclk));
	jdff dff_B_SkgBOMHA8_1(.din(n927),.dout(w_dff_B_SkgBOMHA8_1),.clk(gclk));
	jdff dff_B_0pyGS53w1_1(.din(G292),.dout(w_dff_B_0pyGS53w1_1),.clk(gclk));
	jdff dff_B_9KHWRPD95_1(.din(n1263),.dout(w_dff_B_9KHWRPD95_1),.clk(gclk));
	jdff dff_B_Er7mmR2p2_1(.din(w_dff_B_9KHWRPD95_1),.dout(w_dff_B_Er7mmR2p2_1),.clk(gclk));
	jdff dff_B_Oyi3Kmkh2_1(.din(w_dff_B_Er7mmR2p2_1),.dout(w_dff_B_Oyi3Kmkh2_1),.clk(gclk));
	jdff dff_B_ZRijcHmZ5_1(.din(w_dff_B_Oyi3Kmkh2_1),.dout(w_dff_B_ZRijcHmZ5_1),.clk(gclk));
	jdff dff_B_DuHaqnlu7_1(.din(w_dff_B_ZRijcHmZ5_1),.dout(w_dff_B_DuHaqnlu7_1),.clk(gclk));
	jdff dff_B_6ycKs8Ul5_1(.din(w_dff_B_DuHaqnlu7_1),.dout(w_dff_B_6ycKs8Ul5_1),.clk(gclk));
	jdff dff_B_JojlzJUQ4_1(.din(w_dff_B_6ycKs8Ul5_1),.dout(w_dff_B_JojlzJUQ4_1),.clk(gclk));
	jdff dff_B_wjYXxjZn8_1(.din(w_dff_B_JojlzJUQ4_1),.dout(w_dff_B_wjYXxjZn8_1),.clk(gclk));
	jdff dff_B_xLZueeqH5_1(.din(w_dff_B_wjYXxjZn8_1),.dout(w_dff_B_xLZueeqH5_1),.clk(gclk));
	jdff dff_B_9jmNcFPK6_1(.din(w_dff_B_xLZueeqH5_1),.dout(w_dff_B_9jmNcFPK6_1),.clk(gclk));
	jdff dff_B_huTNExbU1_1(.din(w_dff_B_9jmNcFPK6_1),.dout(w_dff_B_huTNExbU1_1),.clk(gclk));
	jdff dff_B_dS1H8NTI7_1(.din(w_dff_B_huTNExbU1_1),.dout(w_dff_B_dS1H8NTI7_1),.clk(gclk));
	jdff dff_B_I12m6zPC5_1(.din(w_dff_B_dS1H8NTI7_1),.dout(w_dff_B_I12m6zPC5_1),.clk(gclk));
	jdff dff_B_3ITbLQEB2_1(.din(w_dff_B_I12m6zPC5_1),.dout(w_dff_B_3ITbLQEB2_1),.clk(gclk));
	jdff dff_B_4bd8CVAd1_1(.din(w_dff_B_3ITbLQEB2_1),.dout(w_dff_B_4bd8CVAd1_1),.clk(gclk));
	jdff dff_B_oNO33e4M9_1(.din(w_dff_B_4bd8CVAd1_1),.dout(w_dff_B_oNO33e4M9_1),.clk(gclk));
	jdff dff_B_t6kyo3V09_1(.din(w_dff_B_oNO33e4M9_1),.dout(w_dff_B_t6kyo3V09_1),.clk(gclk));
	jdff dff_B_cUGmE2xi7_1(.din(w_dff_B_t6kyo3V09_1),.dout(w_dff_B_cUGmE2xi7_1),.clk(gclk));
	jdff dff_B_t8Pisbq56_1(.din(w_dff_B_cUGmE2xi7_1),.dout(w_dff_B_t8Pisbq56_1),.clk(gclk));
	jdff dff_B_aMRC4USe0_1(.din(n1260),.dout(w_dff_B_aMRC4USe0_1),.clk(gclk));
	jdff dff_B_E2Jbsujk9_1(.din(w_dff_B_aMRC4USe0_1),.dout(w_dff_B_E2Jbsujk9_1),.clk(gclk));
	jdff dff_A_bZjkivdt3_2(.dout(w_n852_6[2]),.din(w_dff_A_bZjkivdt3_2),.clk(gclk));
	jdff dff_A_RUiGa3gj2_2(.dout(w_dff_A_bZjkivdt3_2),.din(w_dff_A_RUiGa3gj2_2),.clk(gclk));
	jdff dff_A_1ZccmPtp3_2(.dout(w_dff_A_RUiGa3gj2_2),.din(w_dff_A_1ZccmPtp3_2),.clk(gclk));
	jdff dff_A_37x9uh2w9_2(.dout(w_dff_A_1ZccmPtp3_2),.din(w_dff_A_37x9uh2w9_2),.clk(gclk));
	jdff dff_A_Fafs4uuO4_2(.dout(w_dff_A_37x9uh2w9_2),.din(w_dff_A_Fafs4uuO4_2),.clk(gclk));
	jdff dff_A_uO8DG4fo7_2(.dout(w_dff_A_Fafs4uuO4_2),.din(w_dff_A_uO8DG4fo7_2),.clk(gclk));
	jdff dff_A_7m5Q2BUn5_2(.dout(w_dff_A_uO8DG4fo7_2),.din(w_dff_A_7m5Q2BUn5_2),.clk(gclk));
	jdff dff_A_T30i9HG34_2(.dout(w_dff_A_7m5Q2BUn5_2),.din(w_dff_A_T30i9HG34_2),.clk(gclk));
	jdff dff_A_f0wWj8nj2_2(.dout(w_dff_A_T30i9HG34_2),.din(w_dff_A_f0wWj8nj2_2),.clk(gclk));
	jdff dff_A_Um4hWMoT3_2(.dout(w_dff_A_f0wWj8nj2_2),.din(w_dff_A_Um4hWMoT3_2),.clk(gclk));
	jdff dff_A_lWXD2SPz5_2(.dout(w_dff_A_Um4hWMoT3_2),.din(w_dff_A_lWXD2SPz5_2),.clk(gclk));
	jdff dff_A_AeIzrj2Q0_2(.dout(w_G4089_6[2]),.din(w_dff_A_AeIzrj2Q0_2),.clk(gclk));
	jdff dff_A_ItY1Ltvz6_2(.dout(w_dff_A_AeIzrj2Q0_2),.din(w_dff_A_ItY1Ltvz6_2),.clk(gclk));
	jdff dff_A_jpDXspEJ9_2(.dout(w_dff_A_ItY1Ltvz6_2),.din(w_dff_A_jpDXspEJ9_2),.clk(gclk));
	jdff dff_A_5tUe9rvx5_2(.dout(w_dff_A_jpDXspEJ9_2),.din(w_dff_A_5tUe9rvx5_2),.clk(gclk));
	jdff dff_A_Yj10R95A7_2(.dout(w_dff_A_5tUe9rvx5_2),.din(w_dff_A_Yj10R95A7_2),.clk(gclk));
	jdff dff_A_ZWJnLsyK3_2(.dout(w_dff_A_Yj10R95A7_2),.din(w_dff_A_ZWJnLsyK3_2),.clk(gclk));
	jdff dff_A_9TNq5Mf22_2(.dout(w_dff_A_ZWJnLsyK3_2),.din(w_dff_A_9TNq5Mf22_2),.clk(gclk));
	jdff dff_A_6Be3uynq4_2(.dout(w_dff_A_9TNq5Mf22_2),.din(w_dff_A_6Be3uynq4_2),.clk(gclk));
	jdff dff_A_36d3tN5Z3_2(.dout(w_dff_A_6Be3uynq4_2),.din(w_dff_A_36d3tN5Z3_2),.clk(gclk));
	jdff dff_A_OQhmWYMb7_2(.dout(w_dff_A_36d3tN5Z3_2),.din(w_dff_A_OQhmWYMb7_2),.clk(gclk));
	jdff dff_A_aJTmaqrM1_2(.dout(w_dff_A_OQhmWYMb7_2),.din(w_dff_A_aJTmaqrM1_2),.clk(gclk));
	jdff dff_A_gat0Rh1U3_2(.dout(w_dff_A_aJTmaqrM1_2),.din(w_dff_A_gat0Rh1U3_2),.clk(gclk));
	jdff dff_A_FWefk98T1_2(.dout(w_dff_A_gat0Rh1U3_2),.din(w_dff_A_FWefk98T1_2),.clk(gclk));
	jdff dff_A_aqR0O6v62_2(.dout(w_dff_A_FWefk98T1_2),.din(w_dff_A_aqR0O6v62_2),.clk(gclk));
	jdff dff_B_B45DUgTt2_0(.din(n1276),.dout(w_dff_B_B45DUgTt2_0),.clk(gclk));
	jdff dff_B_dejdAlZU0_0(.din(w_dff_B_B45DUgTt2_0),.dout(w_dff_B_dejdAlZU0_0),.clk(gclk));
	jdff dff_B_8PrbAwoS9_0(.din(w_dff_B_dejdAlZU0_0),.dout(w_dff_B_8PrbAwoS9_0),.clk(gclk));
	jdff dff_B_ttBS6XoF1_0(.din(w_dff_B_8PrbAwoS9_0),.dout(w_dff_B_ttBS6XoF1_0),.clk(gclk));
	jdff dff_B_tJP0xN0h9_0(.din(w_dff_B_ttBS6XoF1_0),.dout(w_dff_B_tJP0xN0h9_0),.clk(gclk));
	jdff dff_B_i0LsO6C66_0(.din(w_dff_B_tJP0xN0h9_0),.dout(w_dff_B_i0LsO6C66_0),.clk(gclk));
	jdff dff_B_IFnR1WK97_0(.din(w_dff_B_i0LsO6C66_0),.dout(w_dff_B_IFnR1WK97_0),.clk(gclk));
	jdff dff_B_SkSZD2h31_0(.din(w_dff_B_IFnR1WK97_0),.dout(w_dff_B_SkSZD2h31_0),.clk(gclk));
	jdff dff_B_izG3v0Ph6_0(.din(w_dff_B_SkSZD2h31_0),.dout(w_dff_B_izG3v0Ph6_0),.clk(gclk));
	jdff dff_B_bFVLsN1s0_0(.din(w_dff_B_izG3v0Ph6_0),.dout(w_dff_B_bFVLsN1s0_0),.clk(gclk));
	jdff dff_B_7a3WPSu90_0(.din(w_dff_B_bFVLsN1s0_0),.dout(w_dff_B_7a3WPSu90_0),.clk(gclk));
	jdff dff_B_x7a7Svar9_0(.din(w_dff_B_7a3WPSu90_0),.dout(w_dff_B_x7a7Svar9_0),.clk(gclk));
	jdff dff_B_URYZe7Nn6_0(.din(w_dff_B_x7a7Svar9_0),.dout(w_dff_B_URYZe7Nn6_0),.clk(gclk));
	jdff dff_B_HLv28OkZ4_0(.din(w_dff_B_URYZe7Nn6_0),.dout(w_dff_B_HLv28OkZ4_0),.clk(gclk));
	jdff dff_B_Fc1eTT6o0_0(.din(w_dff_B_HLv28OkZ4_0),.dout(w_dff_B_Fc1eTT6o0_0),.clk(gclk));
	jdff dff_B_VhsXr6N50_0(.din(w_dff_B_Fc1eTT6o0_0),.dout(w_dff_B_VhsXr6N50_0),.clk(gclk));
	jdff dff_B_aUw039ji2_0(.din(w_dff_B_VhsXr6N50_0),.dout(w_dff_B_aUw039ji2_0),.clk(gclk));
	jdff dff_B_oY37qiuU8_0(.din(w_dff_B_aUw039ji2_0),.dout(w_dff_B_oY37qiuU8_0),.clk(gclk));
	jdff dff_B_qhe0Dfjz0_0(.din(w_dff_B_oY37qiuU8_0),.dout(w_dff_B_qhe0Dfjz0_0),.clk(gclk));
	jdff dff_B_o5O3sxkA8_0(.din(w_dff_B_qhe0Dfjz0_0),.dout(w_dff_B_o5O3sxkA8_0),.clk(gclk));
	jdff dff_B_nKOjYhof4_0(.din(w_dff_B_o5O3sxkA8_0),.dout(w_dff_B_nKOjYhof4_0),.clk(gclk));
	jdff dff_B_GunH8rOf0_2(.din(G106),.dout(w_dff_B_GunH8rOf0_2),.clk(gclk));
	jdff dff_B_TPgcoPC78_1(.din(n1269),.dout(w_dff_B_TPgcoPC78_1),.clk(gclk));
	jdff dff_B_FAOPZv5V7_1(.din(w_dff_B_TPgcoPC78_1),.dout(w_dff_B_FAOPZv5V7_1),.clk(gclk));
	jdff dff_A_YatUVlqb4_0(.dout(w_n797_6[0]),.din(w_dff_A_YatUVlqb4_0),.clk(gclk));
	jdff dff_A_oaMnA73A3_0(.dout(w_dff_A_YatUVlqb4_0),.din(w_dff_A_oaMnA73A3_0),.clk(gclk));
	jdff dff_A_22uuCQQi7_0(.dout(w_dff_A_oaMnA73A3_0),.din(w_dff_A_22uuCQQi7_0),.clk(gclk));
	jdff dff_A_F8cigkBA4_0(.dout(w_dff_A_22uuCQQi7_0),.din(w_dff_A_F8cigkBA4_0),.clk(gclk));
	jdff dff_A_nnxMCx6P2_0(.dout(w_dff_A_F8cigkBA4_0),.din(w_dff_A_nnxMCx6P2_0),.clk(gclk));
	jdff dff_A_G9Qpm1E87_0(.dout(w_dff_A_nnxMCx6P2_0),.din(w_dff_A_G9Qpm1E87_0),.clk(gclk));
	jdff dff_A_XucZTZjo5_0(.dout(w_dff_A_G9Qpm1E87_0),.din(w_dff_A_XucZTZjo5_0),.clk(gclk));
	jdff dff_A_NELJFviY2_0(.dout(w_dff_A_XucZTZjo5_0),.din(w_dff_A_NELJFviY2_0),.clk(gclk));
	jdff dff_A_w1TryHFu4_0(.dout(w_dff_A_NELJFviY2_0),.din(w_dff_A_w1TryHFu4_0),.clk(gclk));
	jdff dff_A_WwSIhvIp1_0(.dout(w_dff_A_w1TryHFu4_0),.din(w_dff_A_WwSIhvIp1_0),.clk(gclk));
	jdff dff_A_rOLPFYlk8_0(.dout(w_dff_A_WwSIhvIp1_0),.din(w_dff_A_rOLPFYlk8_0),.clk(gclk));
	jdff dff_A_fJyIdfnP4_0(.dout(w_dff_A_rOLPFYlk8_0),.din(w_dff_A_fJyIdfnP4_0),.clk(gclk));
	jdff dff_A_Tzb2EKum7_0(.dout(w_dff_A_fJyIdfnP4_0),.din(w_dff_A_Tzb2EKum7_0),.clk(gclk));
	jdff dff_A_ZZ8wciG30_0(.dout(w_dff_A_Tzb2EKum7_0),.din(w_dff_A_ZZ8wciG30_0),.clk(gclk));
	jdff dff_A_Nd1rsUZb0_0(.dout(w_dff_A_ZZ8wciG30_0),.din(w_dff_A_Nd1rsUZb0_0),.clk(gclk));
	jdff dff_A_wcDu4QUg9_0(.dout(w_dff_A_Nd1rsUZb0_0),.din(w_dff_A_wcDu4QUg9_0),.clk(gclk));
	jdff dff_A_8mFeL7In5_0(.dout(w_dff_A_wcDu4QUg9_0),.din(w_dff_A_8mFeL7In5_0),.clk(gclk));
	jdff dff_A_MYGqcyeX0_0(.dout(w_dff_A_8mFeL7In5_0),.din(w_dff_A_MYGqcyeX0_0),.clk(gclk));
	jdff dff_A_Cc5w5p4o8_0(.dout(w_dff_A_MYGqcyeX0_0),.din(w_dff_A_Cc5w5p4o8_0),.clk(gclk));
	jdff dff_A_M62Dgl556_0(.dout(w_dff_A_Cc5w5p4o8_0),.din(w_dff_A_M62Dgl556_0),.clk(gclk));
	jdff dff_A_uArWe7To1_2(.dout(w_n797_6[2]),.din(w_dff_A_uArWe7To1_2),.clk(gclk));
	jdff dff_A_zj7dSgxe2_2(.dout(w_dff_A_uArWe7To1_2),.din(w_dff_A_zj7dSgxe2_2),.clk(gclk));
	jdff dff_A_6ZLfgkNP9_2(.dout(w_dff_A_zj7dSgxe2_2),.din(w_dff_A_6ZLfgkNP9_2),.clk(gclk));
	jdff dff_A_EfRGGn2S9_2(.dout(w_dff_A_6ZLfgkNP9_2),.din(w_dff_A_EfRGGn2S9_2),.clk(gclk));
	jdff dff_A_YHeqpXse7_2(.dout(w_dff_A_EfRGGn2S9_2),.din(w_dff_A_YHeqpXse7_2),.clk(gclk));
	jdff dff_A_RYD1MbQy8_2(.dout(w_dff_A_YHeqpXse7_2),.din(w_dff_A_RYD1MbQy8_2),.clk(gclk));
	jdff dff_A_r0Kp22jR4_2(.dout(w_dff_A_RYD1MbQy8_2),.din(w_dff_A_r0Kp22jR4_2),.clk(gclk));
	jdff dff_A_2fPKJ0f32_2(.dout(w_dff_A_r0Kp22jR4_2),.din(w_dff_A_2fPKJ0f32_2),.clk(gclk));
	jdff dff_A_DruDHhDh5_2(.dout(w_dff_A_2fPKJ0f32_2),.din(w_dff_A_DruDHhDh5_2),.clk(gclk));
	jdff dff_A_k19TyxIt3_2(.dout(w_dff_A_DruDHhDh5_2),.din(w_dff_A_k19TyxIt3_2),.clk(gclk));
	jdff dff_A_I7AK9l4r1_2(.dout(w_dff_A_k19TyxIt3_2),.din(w_dff_A_I7AK9l4r1_2),.clk(gclk));
	jdff dff_A_B5Y6mFqO3_0(.dout(w_G4088_6[0]),.din(w_dff_A_B5Y6mFqO3_0),.clk(gclk));
	jdff dff_A_IyvYoxQS1_0(.dout(w_dff_A_B5Y6mFqO3_0),.din(w_dff_A_IyvYoxQS1_0),.clk(gclk));
	jdff dff_A_IIJH541H5_0(.dout(w_dff_A_IyvYoxQS1_0),.din(w_dff_A_IIJH541H5_0),.clk(gclk));
	jdff dff_A_QnOub4wR5_0(.dout(w_dff_A_IIJH541H5_0),.din(w_dff_A_QnOub4wR5_0),.clk(gclk));
	jdff dff_A_YUXrQRt75_0(.dout(w_dff_A_QnOub4wR5_0),.din(w_dff_A_YUXrQRt75_0),.clk(gclk));
	jdff dff_A_sw69g0bl1_0(.dout(w_dff_A_YUXrQRt75_0),.din(w_dff_A_sw69g0bl1_0),.clk(gclk));
	jdff dff_A_cVbZI1bH3_0(.dout(w_dff_A_sw69g0bl1_0),.din(w_dff_A_cVbZI1bH3_0),.clk(gclk));
	jdff dff_A_oxJMVX9b7_0(.dout(w_dff_A_cVbZI1bH3_0),.din(w_dff_A_oxJMVX9b7_0),.clk(gclk));
	jdff dff_A_Fyv3BL9r0_0(.dout(w_dff_A_oxJMVX9b7_0),.din(w_dff_A_Fyv3BL9r0_0),.clk(gclk));
	jdff dff_A_T5GIKLVB9_0(.dout(w_dff_A_Fyv3BL9r0_0),.din(w_dff_A_T5GIKLVB9_0),.clk(gclk));
	jdff dff_A_65h5CQtB6_0(.dout(w_dff_A_T5GIKLVB9_0),.din(w_dff_A_65h5CQtB6_0),.clk(gclk));
	jdff dff_A_wHmhoBTX2_0(.dout(w_dff_A_65h5CQtB6_0),.din(w_dff_A_wHmhoBTX2_0),.clk(gclk));
	jdff dff_A_4vpslvjp9_0(.dout(w_dff_A_wHmhoBTX2_0),.din(w_dff_A_4vpslvjp9_0),.clk(gclk));
	jdff dff_A_5Fv0ohq61_0(.dout(w_dff_A_4vpslvjp9_0),.din(w_dff_A_5Fv0ohq61_0),.clk(gclk));
	jdff dff_A_ghGyuOvf7_0(.dout(w_dff_A_5Fv0ohq61_0),.din(w_dff_A_ghGyuOvf7_0),.clk(gclk));
	jdff dff_A_tAqmXO6k5_0(.dout(w_dff_A_ghGyuOvf7_0),.din(w_dff_A_tAqmXO6k5_0),.clk(gclk));
	jdff dff_A_qQ3ncG7g3_0(.dout(w_dff_A_tAqmXO6k5_0),.din(w_dff_A_qQ3ncG7g3_0),.clk(gclk));
	jdff dff_A_TheF06gb3_0(.dout(w_dff_A_qQ3ncG7g3_0),.din(w_dff_A_TheF06gb3_0),.clk(gclk));
	jdff dff_A_jNwxG6DG5_0(.dout(w_dff_A_TheF06gb3_0),.din(w_dff_A_jNwxG6DG5_0),.clk(gclk));
	jdff dff_A_ckOVcIE78_0(.dout(w_dff_A_jNwxG6DG5_0),.din(w_dff_A_ckOVcIE78_0),.clk(gclk));
	jdff dff_A_ITruMqol5_2(.dout(w_G4088_6[2]),.din(w_dff_A_ITruMqol5_2),.clk(gclk));
	jdff dff_A_yTwjobei1_2(.dout(w_dff_A_ITruMqol5_2),.din(w_dff_A_yTwjobei1_2),.clk(gclk));
	jdff dff_A_74UCQE2E4_2(.dout(w_dff_A_yTwjobei1_2),.din(w_dff_A_74UCQE2E4_2),.clk(gclk));
	jdff dff_A_7Vml2f5s0_2(.dout(w_dff_A_74UCQE2E4_2),.din(w_dff_A_7Vml2f5s0_2),.clk(gclk));
	jdff dff_A_vTixQkao9_2(.dout(w_dff_A_7Vml2f5s0_2),.din(w_dff_A_vTixQkao9_2),.clk(gclk));
	jdff dff_A_e1eKY6Mv4_2(.dout(w_dff_A_vTixQkao9_2),.din(w_dff_A_e1eKY6Mv4_2),.clk(gclk));
	jdff dff_A_4mvA1vTd7_2(.dout(w_dff_A_e1eKY6Mv4_2),.din(w_dff_A_4mvA1vTd7_2),.clk(gclk));
	jdff dff_A_rywWiyIt8_2(.dout(w_dff_A_4mvA1vTd7_2),.din(w_dff_A_rywWiyIt8_2),.clk(gclk));
	jdff dff_A_1SHa7NTa3_2(.dout(w_dff_A_rywWiyIt8_2),.din(w_dff_A_1SHa7NTa3_2),.clk(gclk));
	jdff dff_A_vZqizPIh5_2(.dout(w_dff_A_1SHa7NTa3_2),.din(w_dff_A_vZqizPIh5_2),.clk(gclk));
	jdff dff_A_MQ8GbLfP9_2(.dout(w_dff_A_vZqizPIh5_2),.din(w_dff_A_MQ8GbLfP9_2),.clk(gclk));
	jdff dff_A_H2fhytxY0_2(.dout(w_dff_A_MQ8GbLfP9_2),.din(w_dff_A_H2fhytxY0_2),.clk(gclk));
	jdff dff_A_yL7b2mlw7_2(.dout(w_dff_A_H2fhytxY0_2),.din(w_dff_A_yL7b2mlw7_2),.clk(gclk));
	jdff dff_A_FCfSnQoz9_2(.dout(w_dff_A_yL7b2mlw7_2),.din(w_dff_A_FCfSnQoz9_2),.clk(gclk));
	jdff dff_B_sNyM61C42_0(.din(n1286),.dout(w_dff_B_sNyM61C42_0),.clk(gclk));
	jdff dff_B_VUudYJUS1_0(.din(w_dff_B_sNyM61C42_0),.dout(w_dff_B_VUudYJUS1_0),.clk(gclk));
	jdff dff_B_fQhLgF0i8_0(.din(w_dff_B_VUudYJUS1_0),.dout(w_dff_B_fQhLgF0i8_0),.clk(gclk));
	jdff dff_B_fK7jVfCM7_0(.din(w_dff_B_fQhLgF0i8_0),.dout(w_dff_B_fK7jVfCM7_0),.clk(gclk));
	jdff dff_B_OzaYxBVF8_0(.din(w_dff_B_fK7jVfCM7_0),.dout(w_dff_B_OzaYxBVF8_0),.clk(gclk));
	jdff dff_B_Y7EpLbKs6_0(.din(w_dff_B_OzaYxBVF8_0),.dout(w_dff_B_Y7EpLbKs6_0),.clk(gclk));
	jdff dff_B_88UUoN8p2_0(.din(w_dff_B_Y7EpLbKs6_0),.dout(w_dff_B_88UUoN8p2_0),.clk(gclk));
	jdff dff_B_kAZbV6ZR8_0(.din(w_dff_B_88UUoN8p2_0),.dout(w_dff_B_kAZbV6ZR8_0),.clk(gclk));
	jdff dff_B_eSvvKxEW5_0(.din(w_dff_B_kAZbV6ZR8_0),.dout(w_dff_B_eSvvKxEW5_0),.clk(gclk));
	jdff dff_B_1vlxJ8pG3_0(.din(w_dff_B_eSvvKxEW5_0),.dout(w_dff_B_1vlxJ8pG3_0),.clk(gclk));
	jdff dff_B_ijCYObGV6_0(.din(w_dff_B_1vlxJ8pG3_0),.dout(w_dff_B_ijCYObGV6_0),.clk(gclk));
	jdff dff_B_gzlnwjpf2_0(.din(w_dff_B_ijCYObGV6_0),.dout(w_dff_B_gzlnwjpf2_0),.clk(gclk));
	jdff dff_B_06BbwClh5_0(.din(w_dff_B_gzlnwjpf2_0),.dout(w_dff_B_06BbwClh5_0),.clk(gclk));
	jdff dff_B_SxUfn8GP6_0(.din(w_dff_B_06BbwClh5_0),.dout(w_dff_B_SxUfn8GP6_0),.clk(gclk));
	jdff dff_B_9RDZ9AWw3_0(.din(w_dff_B_SxUfn8GP6_0),.dout(w_dff_B_9RDZ9AWw3_0),.clk(gclk));
	jdff dff_B_Q1EKOq2A8_0(.din(w_dff_B_9RDZ9AWw3_0),.dout(w_dff_B_Q1EKOq2A8_0),.clk(gclk));
	jdff dff_B_L3aqFusI8_0(.din(w_dff_B_Q1EKOq2A8_0),.dout(w_dff_B_L3aqFusI8_0),.clk(gclk));
	jdff dff_B_L9TcNWmv1_0(.din(w_dff_B_L3aqFusI8_0),.dout(w_dff_B_L9TcNWmv1_0),.clk(gclk));
	jdff dff_B_hCPLBj4e8_0(.din(w_dff_B_L9TcNWmv1_0),.dout(w_dff_B_hCPLBj4e8_0),.clk(gclk));
	jdff dff_B_ZrjqD6Vp2_0(.din(w_dff_B_hCPLBj4e8_0),.dout(w_dff_B_ZrjqD6Vp2_0),.clk(gclk));
	jdff dff_B_JUonUOeP4_1(.din(n1278),.dout(w_dff_B_JUonUOeP4_1),.clk(gclk));
	jdff dff_B_BqxIVWIf3_1(.din(w_dff_B_JUonUOeP4_1),.dout(w_dff_B_BqxIVWIf3_1),.clk(gclk));
	jdff dff_A_XALJo0765_1(.dout(w_n797_5[1]),.din(w_dff_A_XALJo0765_1),.clk(gclk));
	jdff dff_A_xvhY1EeL9_1(.dout(w_dff_A_XALJo0765_1),.din(w_dff_A_xvhY1EeL9_1),.clk(gclk));
	jdff dff_A_YScRzVKP1_1(.dout(w_dff_A_xvhY1EeL9_1),.din(w_dff_A_YScRzVKP1_1),.clk(gclk));
	jdff dff_A_J7W4h7QO1_1(.dout(w_dff_A_YScRzVKP1_1),.din(w_dff_A_J7W4h7QO1_1),.clk(gclk));
	jdff dff_A_CkVgemj40_1(.dout(w_dff_A_J7W4h7QO1_1),.din(w_dff_A_CkVgemj40_1),.clk(gclk));
	jdff dff_A_qQuHfedU1_1(.dout(w_dff_A_CkVgemj40_1),.din(w_dff_A_qQuHfedU1_1),.clk(gclk));
	jdff dff_A_V9I5XJWd4_1(.dout(w_dff_A_qQuHfedU1_1),.din(w_dff_A_V9I5XJWd4_1),.clk(gclk));
	jdff dff_A_jE6RT3ZK7_1(.dout(w_dff_A_V9I5XJWd4_1),.din(w_dff_A_jE6RT3ZK7_1),.clk(gclk));
	jdff dff_A_PX3PcX5T5_1(.dout(w_dff_A_jE6RT3ZK7_1),.din(w_dff_A_PX3PcX5T5_1),.clk(gclk));
	jdff dff_A_FipmS6DT5_1(.dout(w_dff_A_PX3PcX5T5_1),.din(w_dff_A_FipmS6DT5_1),.clk(gclk));
	jdff dff_A_kCZkX5k74_1(.dout(w_dff_A_FipmS6DT5_1),.din(w_dff_A_kCZkX5k74_1),.clk(gclk));
	jdff dff_A_Z5RO2LRP8_1(.dout(w_dff_A_kCZkX5k74_1),.din(w_dff_A_Z5RO2LRP8_1),.clk(gclk));
	jdff dff_A_Wqyy6HN66_1(.dout(w_dff_A_Z5RO2LRP8_1),.din(w_dff_A_Wqyy6HN66_1),.clk(gclk));
	jdff dff_A_6tdccHF38_1(.dout(w_dff_A_Wqyy6HN66_1),.din(w_dff_A_6tdccHF38_1),.clk(gclk));
	jdff dff_A_XIRbDcxe1_1(.dout(w_dff_A_6tdccHF38_1),.din(w_dff_A_XIRbDcxe1_1),.clk(gclk));
	jdff dff_A_Rs0yfhAM9_1(.dout(w_dff_A_XIRbDcxe1_1),.din(w_dff_A_Rs0yfhAM9_1),.clk(gclk));
	jdff dff_A_ol22gvFD0_1(.dout(w_dff_A_Rs0yfhAM9_1),.din(w_dff_A_ol22gvFD0_1),.clk(gclk));
	jdff dff_A_bymHYt0J5_1(.dout(w_dff_A_ol22gvFD0_1),.din(w_dff_A_bymHYt0J5_1),.clk(gclk));
	jdff dff_A_ziN8tUle8_1(.dout(w_dff_A_bymHYt0J5_1),.din(w_dff_A_ziN8tUle8_1),.clk(gclk));
	jdff dff_A_ZRzb2x1z0_1(.dout(w_G4088_5[1]),.din(w_dff_A_ZRzb2x1z0_1),.clk(gclk));
	jdff dff_A_wGhzLVgY6_1(.dout(w_dff_A_ZRzb2x1z0_1),.din(w_dff_A_wGhzLVgY6_1),.clk(gclk));
	jdff dff_A_IWDv9ApJ2_1(.dout(w_dff_A_wGhzLVgY6_1),.din(w_dff_A_IWDv9ApJ2_1),.clk(gclk));
	jdff dff_A_Glco3OWK0_1(.dout(w_dff_A_IWDv9ApJ2_1),.din(w_dff_A_Glco3OWK0_1),.clk(gclk));
	jdff dff_A_YSijWLRB0_1(.dout(w_dff_A_Glco3OWK0_1),.din(w_dff_A_YSijWLRB0_1),.clk(gclk));
	jdff dff_A_4V5FKOVv6_1(.dout(w_dff_A_YSijWLRB0_1),.din(w_dff_A_4V5FKOVv6_1),.clk(gclk));
	jdff dff_A_UGlWfOtb2_1(.dout(w_dff_A_4V5FKOVv6_1),.din(w_dff_A_UGlWfOtb2_1),.clk(gclk));
	jdff dff_A_9lK2CwjN3_1(.dout(w_dff_A_UGlWfOtb2_1),.din(w_dff_A_9lK2CwjN3_1),.clk(gclk));
	jdff dff_A_ywXdEx3Y3_1(.dout(w_dff_A_9lK2CwjN3_1),.din(w_dff_A_ywXdEx3Y3_1),.clk(gclk));
	jdff dff_A_8x00DkiB5_1(.dout(w_dff_A_ywXdEx3Y3_1),.din(w_dff_A_8x00DkiB5_1),.clk(gclk));
	jdff dff_A_ZAQPBO0B0_1(.dout(w_dff_A_8x00DkiB5_1),.din(w_dff_A_ZAQPBO0B0_1),.clk(gclk));
	jdff dff_A_C332n4v39_1(.dout(w_dff_A_ZAQPBO0B0_1),.din(w_dff_A_C332n4v39_1),.clk(gclk));
	jdff dff_A_eONCbjqm9_1(.dout(w_dff_A_C332n4v39_1),.din(w_dff_A_eONCbjqm9_1),.clk(gclk));
	jdff dff_A_QWegGdz06_1(.dout(w_dff_A_eONCbjqm9_1),.din(w_dff_A_QWegGdz06_1),.clk(gclk));
	jdff dff_A_VNb1TNTD1_1(.dout(w_dff_A_QWegGdz06_1),.din(w_dff_A_VNb1TNTD1_1),.clk(gclk));
	jdff dff_A_YkE488Kg8_1(.dout(w_dff_A_VNb1TNTD1_1),.din(w_dff_A_YkE488Kg8_1),.clk(gclk));
	jdff dff_A_64PowIwJ9_1(.dout(w_dff_A_YkE488Kg8_1),.din(w_dff_A_64PowIwJ9_1),.clk(gclk));
	jdff dff_A_Imr3ajC34_1(.dout(w_dff_A_64PowIwJ9_1),.din(w_dff_A_Imr3ajC34_1),.clk(gclk));
	jdff dff_A_FHmdRqKn5_1(.dout(w_dff_A_Imr3ajC34_1),.din(w_dff_A_FHmdRqKn5_1),.clk(gclk));
	jdff dff_B_eYIAq1GA1_0(.din(n1295),.dout(w_dff_B_eYIAq1GA1_0),.clk(gclk));
	jdff dff_B_QYBbsJPU9_0(.din(w_dff_B_eYIAq1GA1_0),.dout(w_dff_B_QYBbsJPU9_0),.clk(gclk));
	jdff dff_B_zGh82wrr9_0(.din(w_dff_B_QYBbsJPU9_0),.dout(w_dff_B_zGh82wrr9_0),.clk(gclk));
	jdff dff_B_YsDCrJDR7_0(.din(w_dff_B_zGh82wrr9_0),.dout(w_dff_B_YsDCrJDR7_0),.clk(gclk));
	jdff dff_B_O4Ev20zU0_0(.din(w_dff_B_YsDCrJDR7_0),.dout(w_dff_B_O4Ev20zU0_0),.clk(gclk));
	jdff dff_B_n2YgP0Z66_0(.din(w_dff_B_O4Ev20zU0_0),.dout(w_dff_B_n2YgP0Z66_0),.clk(gclk));
	jdff dff_B_fK8BoHQY7_0(.din(w_dff_B_n2YgP0Z66_0),.dout(w_dff_B_fK8BoHQY7_0),.clk(gclk));
	jdff dff_B_7mOewhfc0_0(.din(w_dff_B_fK8BoHQY7_0),.dout(w_dff_B_7mOewhfc0_0),.clk(gclk));
	jdff dff_B_9irBfDwT6_0(.din(w_dff_B_7mOewhfc0_0),.dout(w_dff_B_9irBfDwT6_0),.clk(gclk));
	jdff dff_B_OKkB7sDT7_0(.din(w_dff_B_9irBfDwT6_0),.dout(w_dff_B_OKkB7sDT7_0),.clk(gclk));
	jdff dff_B_aa85SRPe9_0(.din(w_dff_B_OKkB7sDT7_0),.dout(w_dff_B_aa85SRPe9_0),.clk(gclk));
	jdff dff_B_fBLLpL2Z6_0(.din(w_dff_B_aa85SRPe9_0),.dout(w_dff_B_fBLLpL2Z6_0),.clk(gclk));
	jdff dff_B_sJfJuU600_0(.din(w_dff_B_fBLLpL2Z6_0),.dout(w_dff_B_sJfJuU600_0),.clk(gclk));
	jdff dff_B_EfyyJG1Z1_0(.din(w_dff_B_sJfJuU600_0),.dout(w_dff_B_EfyyJG1Z1_0),.clk(gclk));
	jdff dff_B_WZPliaLL8_0(.din(w_dff_B_EfyyJG1Z1_0),.dout(w_dff_B_WZPliaLL8_0),.clk(gclk));
	jdff dff_B_QuuTKFYE9_0(.din(w_dff_B_WZPliaLL8_0),.dout(w_dff_B_QuuTKFYE9_0),.clk(gclk));
	jdff dff_B_qj1QhnIB5_0(.din(w_dff_B_QuuTKFYE9_0),.dout(w_dff_B_qj1QhnIB5_0),.clk(gclk));
	jdff dff_B_SbWZlCbF9_0(.din(w_dff_B_qj1QhnIB5_0),.dout(w_dff_B_SbWZlCbF9_0),.clk(gclk));
	jdff dff_B_vpNC1Scf1_0(.din(w_dff_B_SbWZlCbF9_0),.dout(w_dff_B_vpNC1Scf1_0),.clk(gclk));
	jdff dff_B_cWwYlpGe4_0(.din(w_dff_B_vpNC1Scf1_0),.dout(w_dff_B_cWwYlpGe4_0),.clk(gclk));
	jdff dff_B_XV8wNjjV6_1(.din(n1288),.dout(w_dff_B_XV8wNjjV6_1),.clk(gclk));
	jdff dff_A_AEZVYED01_2(.dout(w_n800_2[2]),.din(w_dff_A_AEZVYED01_2),.clk(gclk));
	jdff dff_B_Y9s8MDIv2_0(.din(n1306),.dout(w_dff_B_Y9s8MDIv2_0),.clk(gclk));
	jdff dff_B_kI4rUX5V0_0(.din(w_dff_B_Y9s8MDIv2_0),.dout(w_dff_B_kI4rUX5V0_0),.clk(gclk));
	jdff dff_B_zaBMlB7G8_0(.din(w_dff_B_kI4rUX5V0_0),.dout(w_dff_B_zaBMlB7G8_0),.clk(gclk));
	jdff dff_B_q3PibDuZ6_0(.din(w_dff_B_zaBMlB7G8_0),.dout(w_dff_B_q3PibDuZ6_0),.clk(gclk));
	jdff dff_B_jy8nMNMh8_0(.din(w_dff_B_q3PibDuZ6_0),.dout(w_dff_B_jy8nMNMh8_0),.clk(gclk));
	jdff dff_B_t5fQrkdv1_0(.din(w_dff_B_jy8nMNMh8_0),.dout(w_dff_B_t5fQrkdv1_0),.clk(gclk));
	jdff dff_B_pIqRasak7_0(.din(w_dff_B_t5fQrkdv1_0),.dout(w_dff_B_pIqRasak7_0),.clk(gclk));
	jdff dff_B_kj977yMF8_0(.din(w_dff_B_pIqRasak7_0),.dout(w_dff_B_kj977yMF8_0),.clk(gclk));
	jdff dff_B_KXXa3ahS5_0(.din(w_dff_B_kj977yMF8_0),.dout(w_dff_B_KXXa3ahS5_0),.clk(gclk));
	jdff dff_B_rfPcbXZ02_0(.din(w_dff_B_KXXa3ahS5_0),.dout(w_dff_B_rfPcbXZ02_0),.clk(gclk));
	jdff dff_B_nC3fHxGw1_0(.din(w_dff_B_rfPcbXZ02_0),.dout(w_dff_B_nC3fHxGw1_0),.clk(gclk));
	jdff dff_B_nPD4e4Xh1_0(.din(w_dff_B_nC3fHxGw1_0),.dout(w_dff_B_nPD4e4Xh1_0),.clk(gclk));
	jdff dff_B_7fMbkebf2_0(.din(w_dff_B_nPD4e4Xh1_0),.dout(w_dff_B_7fMbkebf2_0),.clk(gclk));
	jdff dff_B_TUi0c0967_0(.din(w_dff_B_7fMbkebf2_0),.dout(w_dff_B_TUi0c0967_0),.clk(gclk));
	jdff dff_B_h4pD3d1Q3_0(.din(w_dff_B_TUi0c0967_0),.dout(w_dff_B_h4pD3d1Q3_0),.clk(gclk));
	jdff dff_B_0LdIGTMp2_0(.din(w_dff_B_h4pD3d1Q3_0),.dout(w_dff_B_0LdIGTMp2_0),.clk(gclk));
	jdff dff_B_YaPJtFmK6_0(.din(w_dff_B_0LdIGTMp2_0),.dout(w_dff_B_YaPJtFmK6_0),.clk(gclk));
	jdff dff_B_50Nw6W212_0(.din(w_dff_B_YaPJtFmK6_0),.dout(w_dff_B_50Nw6W212_0),.clk(gclk));
	jdff dff_B_wUvw5KZf0_0(.din(w_dff_B_50Nw6W212_0),.dout(w_dff_B_wUvw5KZf0_0),.clk(gclk));
	jdff dff_B_wqjCsreb5_1(.din(n1298),.dout(w_dff_B_wqjCsreb5_1),.clk(gclk));
	jdff dff_B_9UvqU0Mw7_1(.din(w_dff_B_wqjCsreb5_1),.dout(w_dff_B_9UvqU0Mw7_1),.clk(gclk));
	jdff dff_B_83ZWJmPx7_1(.din(w_dff_B_9UvqU0Mw7_1),.dout(w_dff_B_83ZWJmPx7_1),.clk(gclk));
	jdff dff_A_4gCQgSGR6_0(.dout(w_n797_4[0]),.din(w_dff_A_4gCQgSGR6_0),.clk(gclk));
	jdff dff_A_rlMoYNHS7_0(.dout(w_dff_A_4gCQgSGR6_0),.din(w_dff_A_rlMoYNHS7_0),.clk(gclk));
	jdff dff_A_0d8ehUXM9_0(.dout(w_dff_A_rlMoYNHS7_0),.din(w_dff_A_0d8ehUXM9_0),.clk(gclk));
	jdff dff_A_sgwSvJ3g2_0(.dout(w_dff_A_0d8ehUXM9_0),.din(w_dff_A_sgwSvJ3g2_0),.clk(gclk));
	jdff dff_A_9XYPqs8J9_0(.dout(w_dff_A_sgwSvJ3g2_0),.din(w_dff_A_9XYPqs8J9_0),.clk(gclk));
	jdff dff_A_MtXIsMij8_0(.dout(w_dff_A_9XYPqs8J9_0),.din(w_dff_A_MtXIsMij8_0),.clk(gclk));
	jdff dff_A_vMmRTEqL0_0(.dout(w_dff_A_MtXIsMij8_0),.din(w_dff_A_vMmRTEqL0_0),.clk(gclk));
	jdff dff_A_sKCqViBB7_0(.dout(w_dff_A_vMmRTEqL0_0),.din(w_dff_A_sKCqViBB7_0),.clk(gclk));
	jdff dff_A_REnppv8d2_0(.dout(w_dff_A_sKCqViBB7_0),.din(w_dff_A_REnppv8d2_0),.clk(gclk));
	jdff dff_A_9jtUpEyV1_0(.dout(w_dff_A_REnppv8d2_0),.din(w_dff_A_9jtUpEyV1_0),.clk(gclk));
	jdff dff_A_HdQVBbvz6_0(.dout(w_dff_A_9jtUpEyV1_0),.din(w_dff_A_HdQVBbvz6_0),.clk(gclk));
	jdff dff_A_O0Alu5EO1_0(.dout(w_dff_A_HdQVBbvz6_0),.din(w_dff_A_O0Alu5EO1_0),.clk(gclk));
	jdff dff_A_Ggo7q89V8_0(.dout(w_dff_A_O0Alu5EO1_0),.din(w_dff_A_Ggo7q89V8_0),.clk(gclk));
	jdff dff_A_YuMrfQl95_0(.dout(w_dff_A_Ggo7q89V8_0),.din(w_dff_A_YuMrfQl95_0),.clk(gclk));
	jdff dff_A_xJSz6cr02_0(.dout(w_dff_A_YuMrfQl95_0),.din(w_dff_A_xJSz6cr02_0),.clk(gclk));
	jdff dff_A_J6eTM2V55_0(.dout(w_dff_A_xJSz6cr02_0),.din(w_dff_A_J6eTM2V55_0),.clk(gclk));
	jdff dff_A_K0qLzoO09_0(.dout(w_dff_A_J6eTM2V55_0),.din(w_dff_A_K0qLzoO09_0),.clk(gclk));
	jdff dff_A_Kyd6tigJ2_0(.dout(w_dff_A_K0qLzoO09_0),.din(w_dff_A_Kyd6tigJ2_0),.clk(gclk));
	jdff dff_A_VoakkPsj4_2(.dout(w_n797_4[2]),.din(w_dff_A_VoakkPsj4_2),.clk(gclk));
	jdff dff_A_za8zazYM5_2(.dout(w_dff_A_VoakkPsj4_2),.din(w_dff_A_za8zazYM5_2),.clk(gclk));
	jdff dff_A_768eAWpu2_2(.dout(w_dff_A_za8zazYM5_2),.din(w_dff_A_768eAWpu2_2),.clk(gclk));
	jdff dff_A_JrluYIVV3_2(.dout(w_dff_A_768eAWpu2_2),.din(w_dff_A_JrluYIVV3_2),.clk(gclk));
	jdff dff_A_wOmc1uPo2_2(.dout(w_dff_A_JrluYIVV3_2),.din(w_dff_A_wOmc1uPo2_2),.clk(gclk));
	jdff dff_A_PpzZuoTb4_2(.dout(w_dff_A_wOmc1uPo2_2),.din(w_dff_A_PpzZuoTb4_2),.clk(gclk));
	jdff dff_A_aRnrflxL7_2(.dout(w_dff_A_PpzZuoTb4_2),.din(w_dff_A_aRnrflxL7_2),.clk(gclk));
	jdff dff_A_MhQ7Nci84_2(.dout(w_dff_A_aRnrflxL7_2),.din(w_dff_A_MhQ7Nci84_2),.clk(gclk));
	jdff dff_A_OKMVwSmv4_2(.dout(w_dff_A_MhQ7Nci84_2),.din(w_dff_A_OKMVwSmv4_2),.clk(gclk));
	jdff dff_A_TPybtCcY5_2(.dout(w_dff_A_OKMVwSmv4_2),.din(w_dff_A_TPybtCcY5_2),.clk(gclk));
	jdff dff_A_mrGswC7c6_2(.dout(w_dff_A_TPybtCcY5_2),.din(w_dff_A_mrGswC7c6_2),.clk(gclk));
	jdff dff_A_Ls1thhwE1_2(.dout(w_dff_A_mrGswC7c6_2),.din(w_dff_A_Ls1thhwE1_2),.clk(gclk));
	jdff dff_A_GFVJTBvp6_2(.dout(w_dff_A_Ls1thhwE1_2),.din(w_dff_A_GFVJTBvp6_2),.clk(gclk));
	jdff dff_A_CeD87hr09_2(.dout(w_dff_A_GFVJTBvp6_2),.din(w_dff_A_CeD87hr09_2),.clk(gclk));
	jdff dff_A_iyvt8MIR3_2(.dout(w_dff_A_CeD87hr09_2),.din(w_dff_A_iyvt8MIR3_2),.clk(gclk));
	jdff dff_A_nE0KVern0_2(.dout(w_dff_A_iyvt8MIR3_2),.din(w_dff_A_nE0KVern0_2),.clk(gclk));
	jdff dff_A_vfNadHEl0_2(.dout(w_dff_A_nE0KVern0_2),.din(w_dff_A_vfNadHEl0_2),.clk(gclk));
	jdff dff_A_TmokUw5w2_2(.dout(w_dff_A_vfNadHEl0_2),.din(w_dff_A_TmokUw5w2_2),.clk(gclk));
	jdff dff_A_MKO4dv4O9_2(.dout(w_dff_A_TmokUw5w2_2),.din(w_dff_A_MKO4dv4O9_2),.clk(gclk));
	jdff dff_A_PPOCxUvs9_0(.dout(w_G4088_4[0]),.din(w_dff_A_PPOCxUvs9_0),.clk(gclk));
	jdff dff_A_6XJVNJyQ8_0(.dout(w_dff_A_PPOCxUvs9_0),.din(w_dff_A_6XJVNJyQ8_0),.clk(gclk));
	jdff dff_A_oLboJLN71_0(.dout(w_dff_A_6XJVNJyQ8_0),.din(w_dff_A_oLboJLN71_0),.clk(gclk));
	jdff dff_A_JbqWqdSV6_0(.dout(w_dff_A_oLboJLN71_0),.din(w_dff_A_JbqWqdSV6_0),.clk(gclk));
	jdff dff_A_mPWSUyxJ4_0(.dout(w_dff_A_JbqWqdSV6_0),.din(w_dff_A_mPWSUyxJ4_0),.clk(gclk));
	jdff dff_A_yrImN39F7_0(.dout(w_dff_A_mPWSUyxJ4_0),.din(w_dff_A_yrImN39F7_0),.clk(gclk));
	jdff dff_A_2aiEzahd3_0(.dout(w_dff_A_yrImN39F7_0),.din(w_dff_A_2aiEzahd3_0),.clk(gclk));
	jdff dff_A_95yoRKHZ7_0(.dout(w_dff_A_2aiEzahd3_0),.din(w_dff_A_95yoRKHZ7_0),.clk(gclk));
	jdff dff_A_TZRiJMdD0_0(.dout(w_dff_A_95yoRKHZ7_0),.din(w_dff_A_TZRiJMdD0_0),.clk(gclk));
	jdff dff_A_fX256Ym36_0(.dout(w_dff_A_TZRiJMdD0_0),.din(w_dff_A_fX256Ym36_0),.clk(gclk));
	jdff dff_A_8ofDLLrF9_0(.dout(w_dff_A_fX256Ym36_0),.din(w_dff_A_8ofDLLrF9_0),.clk(gclk));
	jdff dff_A_jBVkFGap8_0(.dout(w_dff_A_8ofDLLrF9_0),.din(w_dff_A_jBVkFGap8_0),.clk(gclk));
	jdff dff_A_HICobnjJ7_0(.dout(w_dff_A_jBVkFGap8_0),.din(w_dff_A_HICobnjJ7_0),.clk(gclk));
	jdff dff_A_ETtM8T6Z3_0(.dout(w_dff_A_HICobnjJ7_0),.din(w_dff_A_ETtM8T6Z3_0),.clk(gclk));
	jdff dff_A_JY1n396d6_0(.dout(w_dff_A_ETtM8T6Z3_0),.din(w_dff_A_JY1n396d6_0),.clk(gclk));
	jdff dff_A_7AQRFNeS9_0(.dout(w_dff_A_JY1n396d6_0),.din(w_dff_A_7AQRFNeS9_0),.clk(gclk));
	jdff dff_A_7Swbm09q8_0(.dout(w_dff_A_7AQRFNeS9_0),.din(w_dff_A_7Swbm09q8_0),.clk(gclk));
	jdff dff_A_g1Tf0iTQ7_2(.dout(w_G4088_4[2]),.din(w_dff_A_g1Tf0iTQ7_2),.clk(gclk));
	jdff dff_A_m70sggur0_2(.dout(w_dff_A_g1Tf0iTQ7_2),.din(w_dff_A_m70sggur0_2),.clk(gclk));
	jdff dff_A_FDtVVnMn4_2(.dout(w_dff_A_m70sggur0_2),.din(w_dff_A_FDtVVnMn4_2),.clk(gclk));
	jdff dff_A_KIXZiPsY5_2(.dout(w_dff_A_FDtVVnMn4_2),.din(w_dff_A_KIXZiPsY5_2),.clk(gclk));
	jdff dff_A_4kChQZ8h5_2(.dout(w_dff_A_KIXZiPsY5_2),.din(w_dff_A_4kChQZ8h5_2),.clk(gclk));
	jdff dff_A_nmwvYoTM2_2(.dout(w_dff_A_4kChQZ8h5_2),.din(w_dff_A_nmwvYoTM2_2),.clk(gclk));
	jdff dff_A_d5Ryocg67_2(.dout(w_dff_A_nmwvYoTM2_2),.din(w_dff_A_d5Ryocg67_2),.clk(gclk));
	jdff dff_A_HMukPqrW3_2(.dout(w_dff_A_d5Ryocg67_2),.din(w_dff_A_HMukPqrW3_2),.clk(gclk));
	jdff dff_A_yVNf7jod6_2(.dout(w_dff_A_HMukPqrW3_2),.din(w_dff_A_yVNf7jod6_2),.clk(gclk));
	jdff dff_A_20b70NDv3_2(.dout(w_dff_A_yVNf7jod6_2),.din(w_dff_A_20b70NDv3_2),.clk(gclk));
	jdff dff_A_7E1tYVwx3_2(.dout(w_dff_A_20b70NDv3_2),.din(w_dff_A_7E1tYVwx3_2),.clk(gclk));
	jdff dff_A_ZkvBa6zQ2_2(.dout(w_dff_A_7E1tYVwx3_2),.din(w_dff_A_ZkvBa6zQ2_2),.clk(gclk));
	jdff dff_A_sKkZe3G20_2(.dout(w_dff_A_ZkvBa6zQ2_2),.din(w_dff_A_sKkZe3G20_2),.clk(gclk));
	jdff dff_A_jfcvFFFJ0_2(.dout(w_dff_A_sKkZe3G20_2),.din(w_dff_A_jfcvFFFJ0_2),.clk(gclk));
	jdff dff_A_ItTHYXAt0_2(.dout(w_dff_A_jfcvFFFJ0_2),.din(w_dff_A_ItTHYXAt0_2),.clk(gclk));
	jdff dff_A_SIDaAc2k1_2(.dout(w_dff_A_ItTHYXAt0_2),.din(w_dff_A_SIDaAc2k1_2),.clk(gclk));
	jdff dff_A_CWC3y3JR5_2(.dout(w_dff_A_SIDaAc2k1_2),.din(w_dff_A_CWC3y3JR5_2),.clk(gclk));
	jdff dff_A_ZYuvNFx13_2(.dout(w_dff_A_CWC3y3JR5_2),.din(w_dff_A_ZYuvNFx13_2),.clk(gclk));
	jdff dff_A_TLCH7n487_2(.dout(w_dff_A_ZYuvNFx13_2),.din(w_dff_A_TLCH7n487_2),.clk(gclk));
	jdff dff_A_pjKoofEh2_2(.dout(w_dff_A_TLCH7n487_2),.din(w_dff_A_pjKoofEh2_2),.clk(gclk));
	jdff dff_B_J60eXKgG2_0(.din(n1315),.dout(w_dff_B_J60eXKgG2_0),.clk(gclk));
	jdff dff_B_WSRhJrnt2_0(.din(w_dff_B_J60eXKgG2_0),.dout(w_dff_B_WSRhJrnt2_0),.clk(gclk));
	jdff dff_B_j4bXQBwu5_0(.din(w_dff_B_WSRhJrnt2_0),.dout(w_dff_B_j4bXQBwu5_0),.clk(gclk));
	jdff dff_B_6bYcj14p9_0(.din(w_dff_B_j4bXQBwu5_0),.dout(w_dff_B_6bYcj14p9_0),.clk(gclk));
	jdff dff_B_YRZTNHsg3_0(.din(w_dff_B_6bYcj14p9_0),.dout(w_dff_B_YRZTNHsg3_0),.clk(gclk));
	jdff dff_B_VL9aqalw4_0(.din(w_dff_B_YRZTNHsg3_0),.dout(w_dff_B_VL9aqalw4_0),.clk(gclk));
	jdff dff_B_3Wqpspjr2_0(.din(w_dff_B_VL9aqalw4_0),.dout(w_dff_B_3Wqpspjr2_0),.clk(gclk));
	jdff dff_B_A3oFkFji7_0(.din(w_dff_B_3Wqpspjr2_0),.dout(w_dff_B_A3oFkFji7_0),.clk(gclk));
	jdff dff_B_t2bE6uZk2_0(.din(w_dff_B_A3oFkFji7_0),.dout(w_dff_B_t2bE6uZk2_0),.clk(gclk));
	jdff dff_B_etWH6cnO7_0(.din(w_dff_B_t2bE6uZk2_0),.dout(w_dff_B_etWH6cnO7_0),.clk(gclk));
	jdff dff_B_HkX3qNgM9_0(.din(w_dff_B_etWH6cnO7_0),.dout(w_dff_B_HkX3qNgM9_0),.clk(gclk));
	jdff dff_B_pkh93CVQ2_0(.din(w_dff_B_HkX3qNgM9_0),.dout(w_dff_B_pkh93CVQ2_0),.clk(gclk));
	jdff dff_B_xAMOHBZi3_0(.din(w_dff_B_pkh93CVQ2_0),.dout(w_dff_B_xAMOHBZi3_0),.clk(gclk));
	jdff dff_B_UsQFK8bR6_0(.din(w_dff_B_xAMOHBZi3_0),.dout(w_dff_B_UsQFK8bR6_0),.clk(gclk));
	jdff dff_B_XcDDGPAj4_0(.din(w_dff_B_UsQFK8bR6_0),.dout(w_dff_B_XcDDGPAj4_0),.clk(gclk));
	jdff dff_B_KFPTwAig1_0(.din(w_dff_B_XcDDGPAj4_0),.dout(w_dff_B_KFPTwAig1_0),.clk(gclk));
	jdff dff_B_rmRVjMwl8_0(.din(w_dff_B_KFPTwAig1_0),.dout(w_dff_B_rmRVjMwl8_0),.clk(gclk));
	jdff dff_B_ZH7tg8vm3_0(.din(w_dff_B_rmRVjMwl8_0),.dout(w_dff_B_ZH7tg8vm3_0),.clk(gclk));
	jdff dff_B_qn1WiwTn9_0(.din(w_dff_B_ZH7tg8vm3_0),.dout(w_dff_B_qn1WiwTn9_0),.clk(gclk));
	jdff dff_B_bsKDHyqd4_0(.din(w_dff_B_qn1WiwTn9_0),.dout(w_dff_B_bsKDHyqd4_0),.clk(gclk));
	jdff dff_B_1iiDpNCJ1_2(.din(G49),.dout(w_dff_B_1iiDpNCJ1_2),.clk(gclk));
	jdff dff_B_ByI9NIUN9_1(.din(n1308),.dout(w_dff_B_ByI9NIUN9_1),.clk(gclk));
	jdff dff_B_GERUinjS1_1(.din(w_dff_B_ByI9NIUN9_1),.dout(w_dff_B_GERUinjS1_1),.clk(gclk));
	jdff dff_A_DmdTJJ9j7_1(.dout(w_n852_5[1]),.din(w_dff_A_DmdTJJ9j7_1),.clk(gclk));
	jdff dff_A_qWlmct5i8_1(.dout(w_dff_A_DmdTJJ9j7_1),.din(w_dff_A_qWlmct5i8_1),.clk(gclk));
	jdff dff_A_RAE24eSo6_1(.dout(w_dff_A_qWlmct5i8_1),.din(w_dff_A_RAE24eSo6_1),.clk(gclk));
	jdff dff_A_I54Bc3Bz4_1(.dout(w_dff_A_RAE24eSo6_1),.din(w_dff_A_I54Bc3Bz4_1),.clk(gclk));
	jdff dff_A_apWsffSX3_1(.dout(w_dff_A_I54Bc3Bz4_1),.din(w_dff_A_apWsffSX3_1),.clk(gclk));
	jdff dff_A_mrRvZvLn9_1(.dout(w_dff_A_apWsffSX3_1),.din(w_dff_A_mrRvZvLn9_1),.clk(gclk));
	jdff dff_A_D6ZeCKFF3_1(.dout(w_dff_A_mrRvZvLn9_1),.din(w_dff_A_D6ZeCKFF3_1),.clk(gclk));
	jdff dff_A_jO3u9WTG8_1(.dout(w_dff_A_D6ZeCKFF3_1),.din(w_dff_A_jO3u9WTG8_1),.clk(gclk));
	jdff dff_A_gbFroE9F2_1(.dout(w_dff_A_jO3u9WTG8_1),.din(w_dff_A_gbFroE9F2_1),.clk(gclk));
	jdff dff_A_3hMaGZQG2_1(.dout(w_dff_A_gbFroE9F2_1),.din(w_dff_A_3hMaGZQG2_1),.clk(gclk));
	jdff dff_A_BD36ye7G7_1(.dout(w_dff_A_3hMaGZQG2_1),.din(w_dff_A_BD36ye7G7_1),.clk(gclk));
	jdff dff_A_Ei9yp1054_1(.dout(w_dff_A_BD36ye7G7_1),.din(w_dff_A_Ei9yp1054_1),.clk(gclk));
	jdff dff_A_U2v2jdlk9_1(.dout(w_dff_A_Ei9yp1054_1),.din(w_dff_A_U2v2jdlk9_1),.clk(gclk));
	jdff dff_A_2kc4YKij9_1(.dout(w_dff_A_U2v2jdlk9_1),.din(w_dff_A_2kc4YKij9_1),.clk(gclk));
	jdff dff_A_xd4xm3Fg1_1(.dout(w_dff_A_2kc4YKij9_1),.din(w_dff_A_xd4xm3Fg1_1),.clk(gclk));
	jdff dff_A_y4tLAUPo7_1(.dout(w_dff_A_xd4xm3Fg1_1),.din(w_dff_A_y4tLAUPo7_1),.clk(gclk));
	jdff dff_A_MoUaTE9L8_1(.dout(w_dff_A_y4tLAUPo7_1),.din(w_dff_A_MoUaTE9L8_1),.clk(gclk));
	jdff dff_A_6oNJnF3U1_1(.dout(w_dff_A_MoUaTE9L8_1),.din(w_dff_A_6oNJnF3U1_1),.clk(gclk));
	jdff dff_A_4xcqPKm27_1(.dout(w_dff_A_6oNJnF3U1_1),.din(w_dff_A_4xcqPKm27_1),.clk(gclk));
	jdff dff_A_UMninGSU0_2(.dout(w_n852_5[2]),.din(w_dff_A_UMninGSU0_2),.clk(gclk));
	jdff dff_A_GC8pYjNn8_2(.dout(w_dff_A_UMninGSU0_2),.din(w_dff_A_GC8pYjNn8_2),.clk(gclk));
	jdff dff_A_axcAwmoL8_2(.dout(w_dff_A_GC8pYjNn8_2),.din(w_dff_A_axcAwmoL8_2),.clk(gclk));
	jdff dff_A_hUEnJQpu2_2(.dout(w_dff_A_axcAwmoL8_2),.din(w_dff_A_hUEnJQpu2_2),.clk(gclk));
	jdff dff_A_sNIPA7qp5_2(.dout(w_dff_A_hUEnJQpu2_2),.din(w_dff_A_sNIPA7qp5_2),.clk(gclk));
	jdff dff_A_PLhEKwZP8_2(.dout(w_dff_A_sNIPA7qp5_2),.din(w_dff_A_PLhEKwZP8_2),.clk(gclk));
	jdff dff_A_I4IF0Pxw3_2(.dout(w_dff_A_PLhEKwZP8_2),.din(w_dff_A_I4IF0Pxw3_2),.clk(gclk));
	jdff dff_A_MKgQu3iE6_2(.dout(w_dff_A_I4IF0Pxw3_2),.din(w_dff_A_MKgQu3iE6_2),.clk(gclk));
	jdff dff_A_YiZcyg1D0_2(.dout(w_dff_A_MKgQu3iE6_2),.din(w_dff_A_YiZcyg1D0_2),.clk(gclk));
	jdff dff_A_rCdV2gmw9_2(.dout(w_dff_A_YiZcyg1D0_2),.din(w_dff_A_rCdV2gmw9_2),.clk(gclk));
	jdff dff_A_i1gwYgew8_2(.dout(w_dff_A_rCdV2gmw9_2),.din(w_dff_A_i1gwYgew8_2),.clk(gclk));
	jdff dff_A_PyK2QKkD6_2(.dout(w_dff_A_i1gwYgew8_2),.din(w_dff_A_PyK2QKkD6_2),.clk(gclk));
	jdff dff_A_VXVyJfZ18_2(.dout(w_dff_A_PyK2QKkD6_2),.din(w_dff_A_VXVyJfZ18_2),.clk(gclk));
	jdff dff_A_05ATyDD63_2(.dout(w_dff_A_VXVyJfZ18_2),.din(w_dff_A_05ATyDD63_2),.clk(gclk));
	jdff dff_A_Gvdq3EKN6_2(.dout(w_dff_A_05ATyDD63_2),.din(w_dff_A_Gvdq3EKN6_2),.clk(gclk));
	jdff dff_A_WHRqcrMG6_2(.dout(w_dff_A_Gvdq3EKN6_2),.din(w_dff_A_WHRqcrMG6_2),.clk(gclk));
	jdff dff_A_qwruWkYt4_2(.dout(w_dff_A_WHRqcrMG6_2),.din(w_dff_A_qwruWkYt4_2),.clk(gclk));
	jdff dff_A_VZe651fN8_2(.dout(w_dff_A_qwruWkYt4_2),.din(w_dff_A_VZe651fN8_2),.clk(gclk));
	jdff dff_A_Il1SW8DM7_2(.dout(w_dff_A_VZe651fN8_2),.din(w_dff_A_Il1SW8DM7_2),.clk(gclk));
	jdff dff_A_tRYBKt5n9_2(.dout(w_dff_A_Il1SW8DM7_2),.din(w_dff_A_tRYBKt5n9_2),.clk(gclk));
	jdff dff_A_VkXPZzYQ4_1(.dout(w_G4089_5[1]),.din(w_dff_A_VkXPZzYQ4_1),.clk(gclk));
	jdff dff_A_9g54clkG4_1(.dout(w_dff_A_VkXPZzYQ4_1),.din(w_dff_A_9g54clkG4_1),.clk(gclk));
	jdff dff_A_zUaKOAz37_1(.dout(w_dff_A_9g54clkG4_1),.din(w_dff_A_zUaKOAz37_1),.clk(gclk));
	jdff dff_A_uZQOUO5N9_1(.dout(w_dff_A_zUaKOAz37_1),.din(w_dff_A_uZQOUO5N9_1),.clk(gclk));
	jdff dff_A_z4AncOV57_1(.dout(w_dff_A_uZQOUO5N9_1),.din(w_dff_A_z4AncOV57_1),.clk(gclk));
	jdff dff_A_lo1Qsoca6_1(.dout(w_dff_A_z4AncOV57_1),.din(w_dff_A_lo1Qsoca6_1),.clk(gclk));
	jdff dff_A_FIJSdwWl5_1(.dout(w_dff_A_lo1Qsoca6_1),.din(w_dff_A_FIJSdwWl5_1),.clk(gclk));
	jdff dff_A_ZT2pKGJ54_1(.dout(w_dff_A_FIJSdwWl5_1),.din(w_dff_A_ZT2pKGJ54_1),.clk(gclk));
	jdff dff_A_xvTq5f9H3_1(.dout(w_dff_A_ZT2pKGJ54_1),.din(w_dff_A_xvTq5f9H3_1),.clk(gclk));
	jdff dff_A_ohbwn4DH0_1(.dout(w_dff_A_xvTq5f9H3_1),.din(w_dff_A_ohbwn4DH0_1),.clk(gclk));
	jdff dff_A_Ap9v18aT1_1(.dout(w_dff_A_ohbwn4DH0_1),.din(w_dff_A_Ap9v18aT1_1),.clk(gclk));
	jdff dff_A_83ihjgF47_1(.dout(w_dff_A_Ap9v18aT1_1),.din(w_dff_A_83ihjgF47_1),.clk(gclk));
	jdff dff_A_LZeWXIrJ9_1(.dout(w_dff_A_83ihjgF47_1),.din(w_dff_A_LZeWXIrJ9_1),.clk(gclk));
	jdff dff_A_tukI4Hbu1_1(.dout(w_dff_A_LZeWXIrJ9_1),.din(w_dff_A_tukI4Hbu1_1),.clk(gclk));
	jdff dff_A_AwnaBnnP8_1(.dout(w_dff_A_tukI4Hbu1_1),.din(w_dff_A_AwnaBnnP8_1),.clk(gclk));
	jdff dff_A_p8ZPVSMX4_1(.dout(w_dff_A_AwnaBnnP8_1),.din(w_dff_A_p8ZPVSMX4_1),.clk(gclk));
	jdff dff_A_aDy7lTlm0_1(.dout(w_dff_A_p8ZPVSMX4_1),.din(w_dff_A_aDy7lTlm0_1),.clk(gclk));
	jdff dff_A_I1luDF322_1(.dout(w_dff_A_aDy7lTlm0_1),.din(w_dff_A_I1luDF322_1),.clk(gclk));
	jdff dff_A_2M1RsakX4_1(.dout(w_dff_A_I1luDF322_1),.din(w_dff_A_2M1RsakX4_1),.clk(gclk));
	jdff dff_A_CT1pJcIv8_2(.dout(w_G4089_5[2]),.din(w_dff_A_CT1pJcIv8_2),.clk(gclk));
	jdff dff_A_QaHUIWPk4_2(.dout(w_dff_A_CT1pJcIv8_2),.din(w_dff_A_QaHUIWPk4_2),.clk(gclk));
	jdff dff_A_dY9oIj3R5_2(.dout(w_dff_A_QaHUIWPk4_2),.din(w_dff_A_dY9oIj3R5_2),.clk(gclk));
	jdff dff_A_SPvbf5KQ7_2(.dout(w_dff_A_dY9oIj3R5_2),.din(w_dff_A_SPvbf5KQ7_2),.clk(gclk));
	jdff dff_A_r02y06yv6_2(.dout(w_dff_A_SPvbf5KQ7_2),.din(w_dff_A_r02y06yv6_2),.clk(gclk));
	jdff dff_A_3qOMgvzZ8_2(.dout(w_dff_A_r02y06yv6_2),.din(w_dff_A_3qOMgvzZ8_2),.clk(gclk));
	jdff dff_A_2fLrrPOJ2_2(.dout(w_dff_A_3qOMgvzZ8_2),.din(w_dff_A_2fLrrPOJ2_2),.clk(gclk));
	jdff dff_A_3H3bu0dK9_2(.dout(w_dff_A_2fLrrPOJ2_2),.din(w_dff_A_3H3bu0dK9_2),.clk(gclk));
	jdff dff_A_EP9lU7jf9_2(.dout(w_dff_A_3H3bu0dK9_2),.din(w_dff_A_EP9lU7jf9_2),.clk(gclk));
	jdff dff_A_iH4ZRY9f4_2(.dout(w_dff_A_EP9lU7jf9_2),.din(w_dff_A_iH4ZRY9f4_2),.clk(gclk));
	jdff dff_A_UaCf8izn3_2(.dout(w_dff_A_iH4ZRY9f4_2),.din(w_dff_A_UaCf8izn3_2),.clk(gclk));
	jdff dff_A_PKpybt2R3_2(.dout(w_dff_A_UaCf8izn3_2),.din(w_dff_A_PKpybt2R3_2),.clk(gclk));
	jdff dff_A_LeQzXgpj2_2(.dout(w_dff_A_PKpybt2R3_2),.din(w_dff_A_LeQzXgpj2_2),.clk(gclk));
	jdff dff_A_qITQm8Z94_2(.dout(w_dff_A_LeQzXgpj2_2),.din(w_dff_A_qITQm8Z94_2),.clk(gclk));
	jdff dff_A_4mAmj4Yt2_2(.dout(w_dff_A_qITQm8Z94_2),.din(w_dff_A_4mAmj4Yt2_2),.clk(gclk));
	jdff dff_A_ynEeKY1O4_2(.dout(w_dff_A_4mAmj4Yt2_2),.din(w_dff_A_ynEeKY1O4_2),.clk(gclk));
	jdff dff_A_hLZQ4Cn07_2(.dout(w_dff_A_ynEeKY1O4_2),.din(w_dff_A_hLZQ4Cn07_2),.clk(gclk));
	jdff dff_A_9QRPuVhF6_2(.dout(w_dff_A_hLZQ4Cn07_2),.din(w_dff_A_9QRPuVhF6_2),.clk(gclk));
	jdff dff_A_hNiW7AmZ6_2(.dout(w_dff_A_9QRPuVhF6_2),.din(w_dff_A_hNiW7AmZ6_2),.clk(gclk));
	jdff dff_A_hd8QYJlY8_2(.dout(w_dff_A_hNiW7AmZ6_2),.din(w_dff_A_hd8QYJlY8_2),.clk(gclk));
	jdff dff_B_VgcngmYy7_0(.din(n1324),.dout(w_dff_B_VgcngmYy7_0),.clk(gclk));
	jdff dff_B_u3FmbG4H7_0(.din(w_dff_B_VgcngmYy7_0),.dout(w_dff_B_u3FmbG4H7_0),.clk(gclk));
	jdff dff_B_PNQGyG9Z1_0(.din(w_dff_B_u3FmbG4H7_0),.dout(w_dff_B_PNQGyG9Z1_0),.clk(gclk));
	jdff dff_B_ziHiVmR14_0(.din(w_dff_B_PNQGyG9Z1_0),.dout(w_dff_B_ziHiVmR14_0),.clk(gclk));
	jdff dff_B_c3tASEs72_0(.din(w_dff_B_ziHiVmR14_0),.dout(w_dff_B_c3tASEs72_0),.clk(gclk));
	jdff dff_B_hrHc12Ln7_0(.din(w_dff_B_c3tASEs72_0),.dout(w_dff_B_hrHc12Ln7_0),.clk(gclk));
	jdff dff_B_SXtFyYYv4_0(.din(w_dff_B_hrHc12Ln7_0),.dout(w_dff_B_SXtFyYYv4_0),.clk(gclk));
	jdff dff_B_eWu49nh12_0(.din(w_dff_B_SXtFyYYv4_0),.dout(w_dff_B_eWu49nh12_0),.clk(gclk));
	jdff dff_B_nQcQNIhA2_0(.din(w_dff_B_eWu49nh12_0),.dout(w_dff_B_nQcQNIhA2_0),.clk(gclk));
	jdff dff_B_ur18KuvB7_0(.din(w_dff_B_nQcQNIhA2_0),.dout(w_dff_B_ur18KuvB7_0),.clk(gclk));
	jdff dff_B_hcoQKYzl9_0(.din(w_dff_B_ur18KuvB7_0),.dout(w_dff_B_hcoQKYzl9_0),.clk(gclk));
	jdff dff_B_Opo8cy6A0_0(.din(w_dff_B_hcoQKYzl9_0),.dout(w_dff_B_Opo8cy6A0_0),.clk(gclk));
	jdff dff_B_ers6BkD50_0(.din(w_dff_B_Opo8cy6A0_0),.dout(w_dff_B_ers6BkD50_0),.clk(gclk));
	jdff dff_B_SPvuNKpO4_0(.din(w_dff_B_ers6BkD50_0),.dout(w_dff_B_SPvuNKpO4_0),.clk(gclk));
	jdff dff_B_LPSobsfJ6_0(.din(w_dff_B_SPvuNKpO4_0),.dout(w_dff_B_LPSobsfJ6_0),.clk(gclk));
	jdff dff_B_6BADGxjz4_0(.din(w_dff_B_LPSobsfJ6_0),.dout(w_dff_B_6BADGxjz4_0),.clk(gclk));
	jdff dff_B_U719I3d97_0(.din(w_dff_B_6BADGxjz4_0),.dout(w_dff_B_U719I3d97_0),.clk(gclk));
	jdff dff_B_9lWbF8ew9_0(.din(w_dff_B_U719I3d97_0),.dout(w_dff_B_9lWbF8ew9_0),.clk(gclk));
	jdff dff_B_OKrlPkE78_0(.din(w_dff_B_9lWbF8ew9_0),.dout(w_dff_B_OKrlPkE78_0),.clk(gclk));
	jdff dff_B_YZF84n0Q0_0(.din(w_dff_B_OKrlPkE78_0),.dout(w_dff_B_YZF84n0Q0_0),.clk(gclk));
	jdff dff_A_oG5NCBMF8_2(.dout(w_G4090_2[2]),.din(w_dff_A_oG5NCBMF8_2),.clk(gclk));
	jdff dff_B_TggzarqU3_2(.din(G103),.dout(w_dff_B_TggzarqU3_2),.clk(gclk));
	jdff dff_B_P8Q07vcW5_1(.din(n1317),.dout(w_dff_B_P8Q07vcW5_1),.clk(gclk));
	jdff dff_B_oWTo4IZ70_0(.din(n1333),.dout(w_dff_B_oWTo4IZ70_0),.clk(gclk));
	jdff dff_B_MWkd3yfS8_0(.din(w_dff_B_oWTo4IZ70_0),.dout(w_dff_B_MWkd3yfS8_0),.clk(gclk));
	jdff dff_B_EiKIeVIS5_0(.din(w_dff_B_MWkd3yfS8_0),.dout(w_dff_B_EiKIeVIS5_0),.clk(gclk));
	jdff dff_B_PTXofejd0_0(.din(w_dff_B_EiKIeVIS5_0),.dout(w_dff_B_PTXofejd0_0),.clk(gclk));
	jdff dff_B_18fZtD3f9_0(.din(w_dff_B_PTXofejd0_0),.dout(w_dff_B_18fZtD3f9_0),.clk(gclk));
	jdff dff_B_T60S0ktL9_0(.din(w_dff_B_18fZtD3f9_0),.dout(w_dff_B_T60S0ktL9_0),.clk(gclk));
	jdff dff_B_XeY8b9oO3_0(.din(w_dff_B_T60S0ktL9_0),.dout(w_dff_B_XeY8b9oO3_0),.clk(gclk));
	jdff dff_B_CK4N7eof6_0(.din(w_dff_B_XeY8b9oO3_0),.dout(w_dff_B_CK4N7eof6_0),.clk(gclk));
	jdff dff_B_GFi2iK3k4_0(.din(w_dff_B_CK4N7eof6_0),.dout(w_dff_B_GFi2iK3k4_0),.clk(gclk));
	jdff dff_B_Cc6c2iMY4_0(.din(w_dff_B_GFi2iK3k4_0),.dout(w_dff_B_Cc6c2iMY4_0),.clk(gclk));
	jdff dff_B_9IWprNb41_0(.din(w_dff_B_Cc6c2iMY4_0),.dout(w_dff_B_9IWprNb41_0),.clk(gclk));
	jdff dff_B_FYCKJ5LT1_0(.din(w_dff_B_9IWprNb41_0),.dout(w_dff_B_FYCKJ5LT1_0),.clk(gclk));
	jdff dff_B_W6vLBPDZ3_0(.din(w_dff_B_FYCKJ5LT1_0),.dout(w_dff_B_W6vLBPDZ3_0),.clk(gclk));
	jdff dff_B_X759oBYN0_0(.din(w_dff_B_W6vLBPDZ3_0),.dout(w_dff_B_X759oBYN0_0),.clk(gclk));
	jdff dff_B_E7AYLJE73_0(.din(w_dff_B_X759oBYN0_0),.dout(w_dff_B_E7AYLJE73_0),.clk(gclk));
	jdff dff_B_ODECBc4B5_0(.din(w_dff_B_E7AYLJE73_0),.dout(w_dff_B_ODECBc4B5_0),.clk(gclk));
	jdff dff_B_KHm83jYH8_0(.din(w_dff_B_ODECBc4B5_0),.dout(w_dff_B_KHm83jYH8_0),.clk(gclk));
	jdff dff_B_tLvTM9XN0_0(.din(w_dff_B_KHm83jYH8_0),.dout(w_dff_B_tLvTM9XN0_0),.clk(gclk));
	jdff dff_B_wucxeoWg8_0(.din(w_dff_B_tLvTM9XN0_0),.dout(w_dff_B_wucxeoWg8_0),.clk(gclk));
	jdff dff_B_g02a7w813_2(.din(G40),.dout(w_dff_B_g02a7w813_2),.clk(gclk));
	jdff dff_B_wH6ZXEK84_1(.din(n1326),.dout(w_dff_B_wH6ZXEK84_1),.clk(gclk));
	jdff dff_B_LV9tmisc5_1(.din(w_dff_B_wH6ZXEK84_1),.dout(w_dff_B_LV9tmisc5_1),.clk(gclk));
	jdff dff_B_gCFCo7wU8_1(.din(w_dff_B_LV9tmisc5_1),.dout(w_dff_B_gCFCo7wU8_1),.clk(gclk));
	jdff dff_A_5f3rJesb7_0(.dout(w_n852_4[0]),.din(w_dff_A_5f3rJesb7_0),.clk(gclk));
	jdff dff_A_GFGDxHB55_0(.dout(w_dff_A_5f3rJesb7_0),.din(w_dff_A_GFGDxHB55_0),.clk(gclk));
	jdff dff_A_UPwfE7ja2_0(.dout(w_dff_A_GFGDxHB55_0),.din(w_dff_A_UPwfE7ja2_0),.clk(gclk));
	jdff dff_A_KaGLihMo7_0(.dout(w_dff_A_UPwfE7ja2_0),.din(w_dff_A_KaGLihMo7_0),.clk(gclk));
	jdff dff_A_XPY1G27t6_0(.dout(w_dff_A_KaGLihMo7_0),.din(w_dff_A_XPY1G27t6_0),.clk(gclk));
	jdff dff_A_otABIdyQ9_0(.dout(w_dff_A_XPY1G27t6_0),.din(w_dff_A_otABIdyQ9_0),.clk(gclk));
	jdff dff_A_Z9P19O0e1_0(.dout(w_dff_A_otABIdyQ9_0),.din(w_dff_A_Z9P19O0e1_0),.clk(gclk));
	jdff dff_A_Iop6I1MH0_0(.dout(w_dff_A_Z9P19O0e1_0),.din(w_dff_A_Iop6I1MH0_0),.clk(gclk));
	jdff dff_A_tg2Qaj433_0(.dout(w_dff_A_Iop6I1MH0_0),.din(w_dff_A_tg2Qaj433_0),.clk(gclk));
	jdff dff_A_MkmjU6aP7_0(.dout(w_dff_A_tg2Qaj433_0),.din(w_dff_A_MkmjU6aP7_0),.clk(gclk));
	jdff dff_A_uPChqG4i2_0(.dout(w_dff_A_MkmjU6aP7_0),.din(w_dff_A_uPChqG4i2_0),.clk(gclk));
	jdff dff_A_pApaFv0r8_0(.dout(w_dff_A_uPChqG4i2_0),.din(w_dff_A_pApaFv0r8_0),.clk(gclk));
	jdff dff_A_0kcoK7jF6_0(.dout(w_dff_A_pApaFv0r8_0),.din(w_dff_A_0kcoK7jF6_0),.clk(gclk));
	jdff dff_A_HUdzpgs96_0(.dout(w_dff_A_0kcoK7jF6_0),.din(w_dff_A_HUdzpgs96_0),.clk(gclk));
	jdff dff_A_qBX1WSOm7_0(.dout(w_dff_A_HUdzpgs96_0),.din(w_dff_A_qBX1WSOm7_0),.clk(gclk));
	jdff dff_A_pLczTBe23_0(.dout(w_dff_A_qBX1WSOm7_0),.din(w_dff_A_pLczTBe23_0),.clk(gclk));
	jdff dff_A_GNABojvH5_0(.dout(w_dff_A_pLczTBe23_0),.din(w_dff_A_GNABojvH5_0),.clk(gclk));
	jdff dff_A_ProXiB0p1_0(.dout(w_dff_A_GNABojvH5_0),.din(w_dff_A_ProXiB0p1_0),.clk(gclk));
	jdff dff_A_ZArgnJNj4_2(.dout(w_n852_4[2]),.din(w_dff_A_ZArgnJNj4_2),.clk(gclk));
	jdff dff_A_uFtIcpUa3_2(.dout(w_dff_A_ZArgnJNj4_2),.din(w_dff_A_uFtIcpUa3_2),.clk(gclk));
	jdff dff_A_ZViEz3Tc8_2(.dout(w_dff_A_uFtIcpUa3_2),.din(w_dff_A_ZViEz3Tc8_2),.clk(gclk));
	jdff dff_A_cbDFD91B8_2(.dout(w_dff_A_ZViEz3Tc8_2),.din(w_dff_A_cbDFD91B8_2),.clk(gclk));
	jdff dff_A_1Rk7d5hL9_2(.dout(w_dff_A_cbDFD91B8_2),.din(w_dff_A_1Rk7d5hL9_2),.clk(gclk));
	jdff dff_A_vDMqAGR29_2(.dout(w_dff_A_1Rk7d5hL9_2),.din(w_dff_A_vDMqAGR29_2),.clk(gclk));
	jdff dff_A_Gz14ckvu9_2(.dout(w_dff_A_vDMqAGR29_2),.din(w_dff_A_Gz14ckvu9_2),.clk(gclk));
	jdff dff_A_qMhmKxNO2_2(.dout(w_dff_A_Gz14ckvu9_2),.din(w_dff_A_qMhmKxNO2_2),.clk(gclk));
	jdff dff_A_9FNSNHVl3_2(.dout(w_dff_A_qMhmKxNO2_2),.din(w_dff_A_9FNSNHVl3_2),.clk(gclk));
	jdff dff_A_f7AAWilR6_2(.dout(w_dff_A_9FNSNHVl3_2),.din(w_dff_A_f7AAWilR6_2),.clk(gclk));
	jdff dff_A_xAdEoUSC8_2(.dout(w_dff_A_f7AAWilR6_2),.din(w_dff_A_xAdEoUSC8_2),.clk(gclk));
	jdff dff_A_DhdHWnMz4_2(.dout(w_dff_A_xAdEoUSC8_2),.din(w_dff_A_DhdHWnMz4_2),.clk(gclk));
	jdff dff_A_oK6VCFfR3_2(.dout(w_dff_A_DhdHWnMz4_2),.din(w_dff_A_oK6VCFfR3_2),.clk(gclk));
	jdff dff_A_tvwMDykL8_2(.dout(w_dff_A_oK6VCFfR3_2),.din(w_dff_A_tvwMDykL8_2),.clk(gclk));
	jdff dff_A_89qTCW2n0_2(.dout(w_dff_A_tvwMDykL8_2),.din(w_dff_A_89qTCW2n0_2),.clk(gclk));
	jdff dff_A_uK5rKovo2_2(.dout(w_dff_A_89qTCW2n0_2),.din(w_dff_A_uK5rKovo2_2),.clk(gclk));
	jdff dff_A_Zq8Ea4cw1_2(.dout(w_dff_A_uK5rKovo2_2),.din(w_dff_A_Zq8Ea4cw1_2),.clk(gclk));
	jdff dff_A_aKN8QaHX4_2(.dout(w_dff_A_Zq8Ea4cw1_2),.din(w_dff_A_aKN8QaHX4_2),.clk(gclk));
	jdff dff_A_w2NP7IaK8_2(.dout(w_dff_A_aKN8QaHX4_2),.din(w_dff_A_w2NP7IaK8_2),.clk(gclk));
	jdff dff_A_ZEpNc4jf7_0(.dout(w_G4089_4[0]),.din(w_dff_A_ZEpNc4jf7_0),.clk(gclk));
	jdff dff_A_zcIJje8M8_0(.dout(w_dff_A_ZEpNc4jf7_0),.din(w_dff_A_zcIJje8M8_0),.clk(gclk));
	jdff dff_A_X20Sckfq9_0(.dout(w_dff_A_zcIJje8M8_0),.din(w_dff_A_X20Sckfq9_0),.clk(gclk));
	jdff dff_A_UUUjfqCD6_0(.dout(w_dff_A_X20Sckfq9_0),.din(w_dff_A_UUUjfqCD6_0),.clk(gclk));
	jdff dff_A_VAI9XjON3_0(.dout(w_dff_A_UUUjfqCD6_0),.din(w_dff_A_VAI9XjON3_0),.clk(gclk));
	jdff dff_A_N2x3levN2_0(.dout(w_dff_A_VAI9XjON3_0),.din(w_dff_A_N2x3levN2_0),.clk(gclk));
	jdff dff_A_afVVJGMx7_0(.dout(w_dff_A_N2x3levN2_0),.din(w_dff_A_afVVJGMx7_0),.clk(gclk));
	jdff dff_A_Qn49o1RX4_0(.dout(w_dff_A_afVVJGMx7_0),.din(w_dff_A_Qn49o1RX4_0),.clk(gclk));
	jdff dff_A_NQColUxj0_0(.dout(w_dff_A_Qn49o1RX4_0),.din(w_dff_A_NQColUxj0_0),.clk(gclk));
	jdff dff_A_smWzWTeG8_0(.dout(w_dff_A_NQColUxj0_0),.din(w_dff_A_smWzWTeG8_0),.clk(gclk));
	jdff dff_A_xdOE0AV27_0(.dout(w_dff_A_smWzWTeG8_0),.din(w_dff_A_xdOE0AV27_0),.clk(gclk));
	jdff dff_A_TCW1t95Q5_0(.dout(w_dff_A_xdOE0AV27_0),.din(w_dff_A_TCW1t95Q5_0),.clk(gclk));
	jdff dff_A_YwgRfHf62_0(.dout(w_dff_A_TCW1t95Q5_0),.din(w_dff_A_YwgRfHf62_0),.clk(gclk));
	jdff dff_A_G5kEngBQ4_0(.dout(w_dff_A_YwgRfHf62_0),.din(w_dff_A_G5kEngBQ4_0),.clk(gclk));
	jdff dff_A_a4TUhWox8_0(.dout(w_dff_A_G5kEngBQ4_0),.din(w_dff_A_a4TUhWox8_0),.clk(gclk));
	jdff dff_A_qzZ10NaD8_0(.dout(w_dff_A_a4TUhWox8_0),.din(w_dff_A_qzZ10NaD8_0),.clk(gclk));
	jdff dff_A_bkjNZIKN0_0(.dout(w_dff_A_qzZ10NaD8_0),.din(w_dff_A_bkjNZIKN0_0),.clk(gclk));
	jdff dff_A_O9lhhJ3D8_2(.dout(w_G4089_4[2]),.din(w_dff_A_O9lhhJ3D8_2),.clk(gclk));
	jdff dff_A_ZvCc4pju1_2(.dout(w_dff_A_O9lhhJ3D8_2),.din(w_dff_A_ZvCc4pju1_2),.clk(gclk));
	jdff dff_A_k4Wijpaf9_2(.dout(w_dff_A_ZvCc4pju1_2),.din(w_dff_A_k4Wijpaf9_2),.clk(gclk));
	jdff dff_A_A80fwNxP5_2(.dout(w_dff_A_k4Wijpaf9_2),.din(w_dff_A_A80fwNxP5_2),.clk(gclk));
	jdff dff_A_FOaS4qm72_2(.dout(w_dff_A_A80fwNxP5_2),.din(w_dff_A_FOaS4qm72_2),.clk(gclk));
	jdff dff_A_NEaqVqWG9_2(.dout(w_dff_A_FOaS4qm72_2),.din(w_dff_A_NEaqVqWG9_2),.clk(gclk));
	jdff dff_A_4KKowJc26_2(.dout(w_dff_A_NEaqVqWG9_2),.din(w_dff_A_4KKowJc26_2),.clk(gclk));
	jdff dff_A_zFg4PUDz9_2(.dout(w_dff_A_4KKowJc26_2),.din(w_dff_A_zFg4PUDz9_2),.clk(gclk));
	jdff dff_A_GJLMnXCg4_2(.dout(w_dff_A_zFg4PUDz9_2),.din(w_dff_A_GJLMnXCg4_2),.clk(gclk));
	jdff dff_A_y6jj5itR9_2(.dout(w_dff_A_GJLMnXCg4_2),.din(w_dff_A_y6jj5itR9_2),.clk(gclk));
	jdff dff_A_utr5CoJO4_2(.dout(w_dff_A_y6jj5itR9_2),.din(w_dff_A_utr5CoJO4_2),.clk(gclk));
	jdff dff_A_GWBbCcyn4_2(.dout(w_dff_A_utr5CoJO4_2),.din(w_dff_A_GWBbCcyn4_2),.clk(gclk));
	jdff dff_A_Q9hckj7v5_2(.dout(w_dff_A_GWBbCcyn4_2),.din(w_dff_A_Q9hckj7v5_2),.clk(gclk));
	jdff dff_A_5gYJdO0q7_2(.dout(w_dff_A_Q9hckj7v5_2),.din(w_dff_A_5gYJdO0q7_2),.clk(gclk));
	jdff dff_A_JO0x2C7B1_2(.dout(w_dff_A_5gYJdO0q7_2),.din(w_dff_A_JO0x2C7B1_2),.clk(gclk));
	jdff dff_A_uVsnAcgH3_2(.dout(w_dff_A_JO0x2C7B1_2),.din(w_dff_A_uVsnAcgH3_2),.clk(gclk));
	jdff dff_A_833IOcGk4_2(.dout(w_dff_A_uVsnAcgH3_2),.din(w_dff_A_833IOcGk4_2),.clk(gclk));
	jdff dff_A_L1tVDxQ90_2(.dout(w_dff_A_833IOcGk4_2),.din(w_dff_A_L1tVDxQ90_2),.clk(gclk));
	jdff dff_A_nc6MxPa65_2(.dout(w_dff_A_L1tVDxQ90_2),.din(w_dff_A_nc6MxPa65_2),.clk(gclk));
	jdff dff_A_fggixee15_2(.dout(w_dff_A_nc6MxPa65_2),.din(w_dff_A_fggixee15_2),.clk(gclk));
	jdff dff_B_mZk8DadO8_0(.din(n1341),.dout(w_dff_B_mZk8DadO8_0),.clk(gclk));
	jdff dff_B_cVT2ypDr2_0(.din(w_dff_B_mZk8DadO8_0),.dout(w_dff_B_cVT2ypDr2_0),.clk(gclk));
	jdff dff_B_v2xyDfLa6_0(.din(w_dff_B_cVT2ypDr2_0),.dout(w_dff_B_v2xyDfLa6_0),.clk(gclk));
	jdff dff_B_X6ceblqR4_0(.din(w_dff_B_v2xyDfLa6_0),.dout(w_dff_B_X6ceblqR4_0),.clk(gclk));
	jdff dff_B_natTV8HQ5_0(.din(w_dff_B_X6ceblqR4_0),.dout(w_dff_B_natTV8HQ5_0),.clk(gclk));
	jdff dff_B_kRU1cT6X6_0(.din(w_dff_B_natTV8HQ5_0),.dout(w_dff_B_kRU1cT6X6_0),.clk(gclk));
	jdff dff_B_kp5I4s5E8_0(.din(w_dff_B_kRU1cT6X6_0),.dout(w_dff_B_kp5I4s5E8_0),.clk(gclk));
	jdff dff_B_QOZYkWO01_0(.din(w_dff_B_kp5I4s5E8_0),.dout(w_dff_B_QOZYkWO01_0),.clk(gclk));
	jdff dff_B_7OO2PNT44_0(.din(w_dff_B_QOZYkWO01_0),.dout(w_dff_B_7OO2PNT44_0),.clk(gclk));
	jdff dff_B_2u48I0ZQ2_0(.din(w_dff_B_7OO2PNT44_0),.dout(w_dff_B_2u48I0ZQ2_0),.clk(gclk));
	jdff dff_B_W3SHrZaa6_0(.din(w_dff_B_2u48I0ZQ2_0),.dout(w_dff_B_W3SHrZaa6_0),.clk(gclk));
	jdff dff_B_yE3crgXW6_0(.din(w_dff_B_W3SHrZaa6_0),.dout(w_dff_B_yE3crgXW6_0),.clk(gclk));
	jdff dff_B_yjJUCC3x5_0(.din(w_dff_B_yE3crgXW6_0),.dout(w_dff_B_yjJUCC3x5_0),.clk(gclk));
	jdff dff_B_AuFJkS3l9_0(.din(w_dff_B_yjJUCC3x5_0),.dout(w_dff_B_AuFJkS3l9_0),.clk(gclk));
	jdff dff_B_fztX6vIt0_0(.din(w_dff_B_AuFJkS3l9_0),.dout(w_dff_B_fztX6vIt0_0),.clk(gclk));
	jdff dff_B_RhWaCaTT4_0(.din(w_dff_B_fztX6vIt0_0),.dout(w_dff_B_RhWaCaTT4_0),.clk(gclk));
	jdff dff_B_Jz9qHEXU8_0(.din(w_dff_B_RhWaCaTT4_0),.dout(w_dff_B_Jz9qHEXU8_0),.clk(gclk));
	jdff dff_B_nFMKQL577_0(.din(w_dff_B_Jz9qHEXU8_0),.dout(w_dff_B_nFMKQL577_0),.clk(gclk));
	jdff dff_B_ubgztRBW1_0(.din(n1340),.dout(w_dff_B_ubgztRBW1_0),.clk(gclk));
	jdff dff_B_zlsu6uTC2_1(.din(n1335),.dout(w_dff_B_zlsu6uTC2_1),.clk(gclk));
	jdff dff_B_tXKxrf9s1_1(.din(w_dff_B_zlsu6uTC2_1),.dout(w_dff_B_tXKxrf9s1_1),.clk(gclk));
	jdff dff_B_ABsc0nYs4_1(.din(w_dff_B_tXKxrf9s1_1),.dout(w_dff_B_ABsc0nYs4_1),.clk(gclk));
	jdff dff_A_RDLo1Q703_0(.dout(w_n999_2[0]),.din(w_dff_A_RDLo1Q703_0),.clk(gclk));
	jdff dff_A_8gT6Xo5p5_0(.dout(w_dff_A_RDLo1Q703_0),.din(w_dff_A_8gT6Xo5p5_0),.clk(gclk));
	jdff dff_A_0pzcnxNl7_0(.dout(w_dff_A_8gT6Xo5p5_0),.din(w_dff_A_0pzcnxNl7_0),.clk(gclk));
	jdff dff_A_smbNrJg58_0(.dout(w_dff_A_0pzcnxNl7_0),.din(w_dff_A_smbNrJg58_0),.clk(gclk));
	jdff dff_A_B9JONuk91_0(.dout(w_dff_A_smbNrJg58_0),.din(w_dff_A_B9JONuk91_0),.clk(gclk));
	jdff dff_A_gNqVIcRp2_0(.dout(w_dff_A_B9JONuk91_0),.din(w_dff_A_gNqVIcRp2_0),.clk(gclk));
	jdff dff_A_p5R2bQi48_1(.dout(w_n999_2[1]),.din(w_dff_A_p5R2bQi48_1),.clk(gclk));
	jdff dff_A_V4oXL9y83_0(.dout(w_G1689_3[0]),.din(w_dff_A_V4oXL9y83_0),.clk(gclk));
	jdff dff_A_cnXsDLqu5_0(.dout(w_dff_A_V4oXL9y83_0),.din(w_dff_A_cnXsDLqu5_0),.clk(gclk));
	jdff dff_A_o0ci5aYa7_0(.dout(w_dff_A_cnXsDLqu5_0),.din(w_dff_A_o0ci5aYa7_0),.clk(gclk));
	jdff dff_A_9L5JHhJU6_0(.dout(w_dff_A_o0ci5aYa7_0),.din(w_dff_A_9L5JHhJU6_0),.clk(gclk));
	jdff dff_A_qGxOKaZp3_1(.dout(w_G1689_3[1]),.din(w_dff_A_qGxOKaZp3_1),.clk(gclk));
	jdff dff_A_JUUW9lsD8_1(.dout(w_dff_A_qGxOKaZp3_1),.din(w_dff_A_JUUW9lsD8_1),.clk(gclk));
	jdff dff_A_BNNter448_0(.dout(w_G137_6[0]),.din(w_dff_A_BNNter448_0),.clk(gclk));
	jdff dff_A_qZO2Lkdt2_0(.dout(w_dff_A_BNNter448_0),.din(w_dff_A_qZO2Lkdt2_0),.clk(gclk));
	jdff dff_A_e6wOR5rI7_0(.dout(w_dff_A_qZO2Lkdt2_0),.din(w_dff_A_e6wOR5rI7_0),.clk(gclk));
	jdff dff_A_oo6diNym5_0(.dout(w_dff_A_e6wOR5rI7_0),.din(w_dff_A_oo6diNym5_0),.clk(gclk));
	jdff dff_A_0adyCNG52_0(.dout(w_dff_A_oo6diNym5_0),.din(w_dff_A_0adyCNG52_0),.clk(gclk));
	jdff dff_A_iKHdrdEq0_0(.dout(w_dff_A_0adyCNG52_0),.din(w_dff_A_iKHdrdEq0_0),.clk(gclk));
	jdff dff_A_0CrxWVcA1_1(.dout(w_G137_6[1]),.din(w_dff_A_0CrxWVcA1_1),.clk(gclk));
	jdff dff_B_2zwCAScy4_0(.din(n1350),.dout(w_dff_B_2zwCAScy4_0),.clk(gclk));
	jdff dff_B_Mx9K13cZ6_0(.din(w_dff_B_2zwCAScy4_0),.dout(w_dff_B_Mx9K13cZ6_0),.clk(gclk));
	jdff dff_B_nBvGElPF9_0(.din(w_dff_B_Mx9K13cZ6_0),.dout(w_dff_B_nBvGElPF9_0),.clk(gclk));
	jdff dff_B_VV1WvhOR8_0(.din(w_dff_B_nBvGElPF9_0),.dout(w_dff_B_VV1WvhOR8_0),.clk(gclk));
	jdff dff_B_tcUsRVJQ0_0(.din(w_dff_B_VV1WvhOR8_0),.dout(w_dff_B_tcUsRVJQ0_0),.clk(gclk));
	jdff dff_B_mkWUecon1_0(.din(w_dff_B_tcUsRVJQ0_0),.dout(w_dff_B_mkWUecon1_0),.clk(gclk));
	jdff dff_B_GoHOyCPM4_0(.din(w_dff_B_mkWUecon1_0),.dout(w_dff_B_GoHOyCPM4_0),.clk(gclk));
	jdff dff_B_XvcaOzwA5_0(.din(w_dff_B_GoHOyCPM4_0),.dout(w_dff_B_XvcaOzwA5_0),.clk(gclk));
	jdff dff_B_VHn29TaX9_0(.din(w_dff_B_XvcaOzwA5_0),.dout(w_dff_B_VHn29TaX9_0),.clk(gclk));
	jdff dff_B_BSC9Ld8P6_0(.din(w_dff_B_VHn29TaX9_0),.dout(w_dff_B_BSC9Ld8P6_0),.clk(gclk));
	jdff dff_B_Vb3IcSzo1_0(.din(w_dff_B_BSC9Ld8P6_0),.dout(w_dff_B_Vb3IcSzo1_0),.clk(gclk));
	jdff dff_B_Y9BEo8R88_0(.din(w_dff_B_Vb3IcSzo1_0),.dout(w_dff_B_Y9BEo8R88_0),.clk(gclk));
	jdff dff_B_XydEaswq6_0(.din(w_dff_B_Y9BEo8R88_0),.dout(w_dff_B_XydEaswq6_0),.clk(gclk));
	jdff dff_B_oHanbBGp4_0(.din(w_dff_B_XydEaswq6_0),.dout(w_dff_B_oHanbBGp4_0),.clk(gclk));
	jdff dff_B_W045XdAy6_0(.din(w_dff_B_oHanbBGp4_0),.dout(w_dff_B_W045XdAy6_0),.clk(gclk));
	jdff dff_B_wmj0R0Sx4_0(.din(w_dff_B_W045XdAy6_0),.dout(w_dff_B_wmj0R0Sx4_0),.clk(gclk));
	jdff dff_B_ihZKWXYs2_0(.din(w_dff_B_wmj0R0Sx4_0),.dout(w_dff_B_ihZKWXYs2_0),.clk(gclk));
	jdff dff_B_AiOmB4mL5_0(.din(w_dff_B_ihZKWXYs2_0),.dout(w_dff_B_AiOmB4mL5_0),.clk(gclk));
	jdff dff_B_qz6367Se3_0(.din(w_dff_B_AiOmB4mL5_0),.dout(w_dff_B_qz6367Se3_0),.clk(gclk));
	jdff dff_B_GW0o3jnx6_0(.din(n1349),.dout(w_dff_B_GW0o3jnx6_0),.clk(gclk));
	jdff dff_B_dPM72rwn1_1(.din(n1344),.dout(w_dff_B_dPM72rwn1_1),.clk(gclk));
	jdff dff_B_WqFWozgh4_1(.din(n1355),.dout(w_dff_B_WqFWozgh4_1),.clk(gclk));
	jdff dff_B_mZ5mP0hv6_1(.din(w_dff_B_WqFWozgh4_1),.dout(w_dff_B_mZ5mP0hv6_1),.clk(gclk));
	jdff dff_B_aYioYtRr2_1(.din(w_dff_B_mZ5mP0hv6_1),.dout(w_dff_B_aYioYtRr2_1),.clk(gclk));
	jdff dff_B_QxQXc6BT8_1(.din(w_dff_B_aYioYtRr2_1),.dout(w_dff_B_QxQXc6BT8_1),.clk(gclk));
	jdff dff_B_jtKmuv6R5_1(.din(w_dff_B_QxQXc6BT8_1),.dout(w_dff_B_jtKmuv6R5_1),.clk(gclk));
	jdff dff_B_DkGma15y7_1(.din(w_dff_B_jtKmuv6R5_1),.dout(w_dff_B_DkGma15y7_1),.clk(gclk));
	jdff dff_B_5ayhU0Rg2_1(.din(w_dff_B_DkGma15y7_1),.dout(w_dff_B_5ayhU0Rg2_1),.clk(gclk));
	jdff dff_B_JC05rPA08_1(.din(w_dff_B_5ayhU0Rg2_1),.dout(w_dff_B_JC05rPA08_1),.clk(gclk));
	jdff dff_B_ATsFikNj9_1(.din(w_dff_B_JC05rPA08_1),.dout(w_dff_B_ATsFikNj9_1),.clk(gclk));
	jdff dff_B_tZNoVLZI3_1(.din(w_dff_B_ATsFikNj9_1),.dout(w_dff_B_tZNoVLZI3_1),.clk(gclk));
	jdff dff_B_cmuIQCN52_1(.din(w_dff_B_tZNoVLZI3_1),.dout(w_dff_B_cmuIQCN52_1),.clk(gclk));
	jdff dff_B_HHTOpmCQ3_1(.din(w_dff_B_cmuIQCN52_1),.dout(w_dff_B_HHTOpmCQ3_1),.clk(gclk));
	jdff dff_B_HE99HN4o1_1(.din(w_dff_B_HHTOpmCQ3_1),.dout(w_dff_B_HE99HN4o1_1),.clk(gclk));
	jdff dff_B_uK9Hl7HN7_1(.din(w_dff_B_HE99HN4o1_1),.dout(w_dff_B_uK9Hl7HN7_1),.clk(gclk));
	jdff dff_B_MQ9FhYmA6_1(.din(w_dff_B_uK9Hl7HN7_1),.dout(w_dff_B_MQ9FhYmA6_1),.clk(gclk));
	jdff dff_B_QPBFYZcg9_1(.din(w_dff_B_MQ9FhYmA6_1),.dout(w_dff_B_QPBFYZcg9_1),.clk(gclk));
	jdff dff_B_fYORsTpe3_1(.din(w_dff_B_QPBFYZcg9_1),.dout(w_dff_B_fYORsTpe3_1),.clk(gclk));
	jdff dff_B_EcxWEDzd4_1(.din(w_dff_B_fYORsTpe3_1),.dout(w_dff_B_EcxWEDzd4_1),.clk(gclk));
	jdff dff_B_2N7sWeEP9_1(.din(w_dff_B_EcxWEDzd4_1),.dout(w_dff_B_2N7sWeEP9_1),.clk(gclk));
	jdff dff_B_aM7Hh88Z6_1(.din(n1356),.dout(w_dff_B_aM7Hh88Z6_1),.clk(gclk));
	jdff dff_A_6ARgsfXK6_0(.dout(w_n993_2[0]),.din(w_dff_A_6ARgsfXK6_0),.clk(gclk));
	jdff dff_A_2dPucS1o4_1(.dout(w_n993_2[1]),.din(w_dff_A_2dPucS1o4_1),.clk(gclk));
	jdff dff_B_n0fNFoP04_0(.din(n1354),.dout(w_dff_B_n0fNFoP04_0),.clk(gclk));
	jdff dff_B_HZpmXYVr6_1(.din(n1364),.dout(w_dff_B_HZpmXYVr6_1),.clk(gclk));
	jdff dff_B_mZiglbwN2_1(.din(w_dff_B_HZpmXYVr6_1),.dout(w_dff_B_mZiglbwN2_1),.clk(gclk));
	jdff dff_B_9SU1YpQd1_1(.din(w_dff_B_mZiglbwN2_1),.dout(w_dff_B_9SU1YpQd1_1),.clk(gclk));
	jdff dff_B_QHJWhX3r1_1(.din(w_dff_B_9SU1YpQd1_1),.dout(w_dff_B_QHJWhX3r1_1),.clk(gclk));
	jdff dff_B_uaVPONxv7_1(.din(w_dff_B_QHJWhX3r1_1),.dout(w_dff_B_uaVPONxv7_1),.clk(gclk));
	jdff dff_B_fHKgcpxq5_1(.din(w_dff_B_uaVPONxv7_1),.dout(w_dff_B_fHKgcpxq5_1),.clk(gclk));
	jdff dff_B_jfhtiu9j5_1(.din(w_dff_B_fHKgcpxq5_1),.dout(w_dff_B_jfhtiu9j5_1),.clk(gclk));
	jdff dff_B_mtfiZGou8_1(.din(w_dff_B_jfhtiu9j5_1),.dout(w_dff_B_mtfiZGou8_1),.clk(gclk));
	jdff dff_B_45DQP7MI3_1(.din(w_dff_B_mtfiZGou8_1),.dout(w_dff_B_45DQP7MI3_1),.clk(gclk));
	jdff dff_B_QZrZVwZg6_1(.din(w_dff_B_45DQP7MI3_1),.dout(w_dff_B_QZrZVwZg6_1),.clk(gclk));
	jdff dff_B_yE8vwQXY9_1(.din(w_dff_B_QZrZVwZg6_1),.dout(w_dff_B_yE8vwQXY9_1),.clk(gclk));
	jdff dff_B_PiPz5vEE5_1(.din(w_dff_B_yE8vwQXY9_1),.dout(w_dff_B_PiPz5vEE5_1),.clk(gclk));
	jdff dff_B_9k9lo8dS9_1(.din(w_dff_B_PiPz5vEE5_1),.dout(w_dff_B_9k9lo8dS9_1),.clk(gclk));
	jdff dff_B_NOAdkUrY0_1(.din(w_dff_B_9k9lo8dS9_1),.dout(w_dff_B_NOAdkUrY0_1),.clk(gclk));
	jdff dff_B_Ri2MbYJE4_1(.din(w_dff_B_NOAdkUrY0_1),.dout(w_dff_B_Ri2MbYJE4_1),.clk(gclk));
	jdff dff_B_EmsGaU8w7_1(.din(w_dff_B_Ri2MbYJE4_1),.dout(w_dff_B_EmsGaU8w7_1),.clk(gclk));
	jdff dff_B_rmMndIEr1_1(.din(w_dff_B_EmsGaU8w7_1),.dout(w_dff_B_rmMndIEr1_1),.clk(gclk));
	jdff dff_B_9XnAlZqg0_1(.din(w_dff_B_rmMndIEr1_1),.dout(w_dff_B_9XnAlZqg0_1),.clk(gclk));
	jdff dff_B_qHZDVASq7_1(.din(w_dff_B_9XnAlZqg0_1),.dout(w_dff_B_qHZDVASq7_1),.clk(gclk));
	jdff dff_B_9O0W9hO07_1(.din(w_dff_B_qHZDVASq7_1),.dout(w_dff_B_9O0W9hO07_1),.clk(gclk));
	jdff dff_B_ud4zDNMc5_1(.din(n1365),.dout(w_dff_B_ud4zDNMc5_1),.clk(gclk));
	jdff dff_A_HJZRrLEG4_0(.dout(w_G1689_2[0]),.din(w_dff_A_HJZRrLEG4_0),.clk(gclk));
	jdff dff_A_zKLX45dN3_2(.dout(w_G1689_2[2]),.din(w_dff_A_zKLX45dN3_2),.clk(gclk));
	jdff dff_A_UUwchZia9_0(.dout(w_n999_1[0]),.din(w_dff_A_UUwchZia9_0),.clk(gclk));
	jdff dff_A_RlKZcSQj8_0(.dout(w_dff_A_UUwchZia9_0),.din(w_dff_A_RlKZcSQj8_0),.clk(gclk));
	jdff dff_A_Tli91gTS6_1(.dout(w_n999_1[1]),.din(w_dff_A_Tli91gTS6_1),.clk(gclk));
	jdff dff_A_8M2KqIGQ8_0(.dout(w_n999_0[0]),.din(w_dff_A_8M2KqIGQ8_0),.clk(gclk));
	jdff dff_A_8P8FX6qV1_0(.dout(w_dff_A_8M2KqIGQ8_0),.din(w_dff_A_8P8FX6qV1_0),.clk(gclk));
	jdff dff_A_CckW1MhG9_0(.dout(w_dff_A_8P8FX6qV1_0),.din(w_dff_A_CckW1MhG9_0),.clk(gclk));
	jdff dff_A_oe4XpMmv9_0(.dout(w_dff_A_CckW1MhG9_0),.din(w_dff_A_oe4XpMmv9_0),.clk(gclk));
	jdff dff_A_7EZ4YDgG6_0(.dout(w_dff_A_oe4XpMmv9_0),.din(w_dff_A_7EZ4YDgG6_0),.clk(gclk));
	jdff dff_A_VoSiUYyz2_0(.dout(w_dff_A_7EZ4YDgG6_0),.din(w_dff_A_VoSiUYyz2_0),.clk(gclk));
	jdff dff_A_zN00DOpl0_0(.dout(w_dff_A_VoSiUYyz2_0),.din(w_dff_A_zN00DOpl0_0),.clk(gclk));
	jdff dff_A_hFwu1MYn0_0(.dout(w_dff_A_zN00DOpl0_0),.din(w_dff_A_hFwu1MYn0_0),.clk(gclk));
	jdff dff_A_Uh1Kfn9T3_0(.dout(w_dff_A_hFwu1MYn0_0),.din(w_dff_A_Uh1Kfn9T3_0),.clk(gclk));
	jdff dff_A_YtWZNf8k5_0(.dout(w_dff_A_Uh1Kfn9T3_0),.din(w_dff_A_YtWZNf8k5_0),.clk(gclk));
	jdff dff_A_qYXjQuKy8_0(.dout(w_dff_A_YtWZNf8k5_0),.din(w_dff_A_qYXjQuKy8_0),.clk(gclk));
	jdff dff_A_vDJTTgAp5_1(.dout(w_n999_0[1]),.din(w_dff_A_vDJTTgAp5_1),.clk(gclk));
	jdff dff_A_DlPldBzq0_1(.dout(w_dff_A_vDJTTgAp5_1),.din(w_dff_A_DlPldBzq0_1),.clk(gclk));
	jdff dff_A_8oSnNPd36_1(.dout(w_dff_A_DlPldBzq0_1),.din(w_dff_A_8oSnNPd36_1),.clk(gclk));
	jdff dff_A_3J7YtBlR4_1(.dout(w_dff_A_8oSnNPd36_1),.din(w_dff_A_3J7YtBlR4_1),.clk(gclk));
	jdff dff_B_kltcvlBT9_3(.din(n999),.dout(w_dff_B_kltcvlBT9_3),.clk(gclk));
	jdff dff_B_uQ3hNHun0_3(.din(w_dff_B_kltcvlBT9_3),.dout(w_dff_B_uQ3hNHun0_3),.clk(gclk));
	jdff dff_B_DiW1C9fY2_3(.din(w_dff_B_uQ3hNHun0_3),.dout(w_dff_B_DiW1C9fY2_3),.clk(gclk));
	jdff dff_B_I17bN32S5_3(.din(w_dff_B_DiW1C9fY2_3),.dout(w_dff_B_I17bN32S5_3),.clk(gclk));
	jdff dff_B_hWSMz0cz6_3(.din(w_dff_B_I17bN32S5_3),.dout(w_dff_B_hWSMz0cz6_3),.clk(gclk));
	jdff dff_B_VEBeYxTG1_3(.din(w_dff_B_hWSMz0cz6_3),.dout(w_dff_B_VEBeYxTG1_3),.clk(gclk));
	jdff dff_B_HDZl0wU33_3(.din(w_dff_B_VEBeYxTG1_3),.dout(w_dff_B_HDZl0wU33_3),.clk(gclk));
	jdff dff_B_nKJuCJj05_3(.din(w_dff_B_HDZl0wU33_3),.dout(w_dff_B_nKJuCJj05_3),.clk(gclk));
	jdff dff_B_gH9XOfcv5_3(.din(w_dff_B_nKJuCJj05_3),.dout(w_dff_B_gH9XOfcv5_3),.clk(gclk));
	jdff dff_B_WuxwULkX2_0(.din(n1363),.dout(w_dff_B_WuxwULkX2_0),.clk(gclk));
	jdff dff_A_kcz5qDe10_0(.dout(w_G137_5[0]),.din(w_dff_A_kcz5qDe10_0),.clk(gclk));
	jdff dff_B_oNhKQnch1_0(.din(n1377),.dout(w_dff_B_oNhKQnch1_0),.clk(gclk));
	jdff dff_B_t98oNZmA4_0(.din(w_dff_B_oNhKQnch1_0),.dout(w_dff_B_t98oNZmA4_0),.clk(gclk));
	jdff dff_B_fXhRwIXX8_0(.din(w_dff_B_t98oNZmA4_0),.dout(w_dff_B_fXhRwIXX8_0),.clk(gclk));
	jdff dff_B_eT2XgNwZ4_0(.din(w_dff_B_fXhRwIXX8_0),.dout(w_dff_B_eT2XgNwZ4_0),.clk(gclk));
	jdff dff_B_x1vGDLVW9_0(.din(w_dff_B_eT2XgNwZ4_0),.dout(w_dff_B_x1vGDLVW9_0),.clk(gclk));
	jdff dff_B_exUFEdiW6_0(.din(w_dff_B_x1vGDLVW9_0),.dout(w_dff_B_exUFEdiW6_0),.clk(gclk));
	jdff dff_B_tP5Wgawe9_0(.din(w_dff_B_exUFEdiW6_0),.dout(w_dff_B_tP5Wgawe9_0),.clk(gclk));
	jdff dff_B_o97lgQwU2_0(.din(w_dff_B_tP5Wgawe9_0),.dout(w_dff_B_o97lgQwU2_0),.clk(gclk));
	jdff dff_B_ykrhYx5y7_0(.din(w_dff_B_o97lgQwU2_0),.dout(w_dff_B_ykrhYx5y7_0),.clk(gclk));
	jdff dff_B_SPfTink03_0(.din(w_dff_B_ykrhYx5y7_0),.dout(w_dff_B_SPfTink03_0),.clk(gclk));
	jdff dff_B_mG55dgay0_0(.din(w_dff_B_SPfTink03_0),.dout(w_dff_B_mG55dgay0_0),.clk(gclk));
	jdff dff_B_j0r0l8Nh8_0(.din(w_dff_B_mG55dgay0_0),.dout(w_dff_B_j0r0l8Nh8_0),.clk(gclk));
	jdff dff_B_OB95ABOx9_0(.din(w_dff_B_j0r0l8Nh8_0),.dout(w_dff_B_OB95ABOx9_0),.clk(gclk));
	jdff dff_B_jVDwKCqR3_0(.din(w_dff_B_OB95ABOx9_0),.dout(w_dff_B_jVDwKCqR3_0),.clk(gclk));
	jdff dff_B_F7sHR3l28_0(.din(w_dff_B_jVDwKCqR3_0),.dout(w_dff_B_F7sHR3l28_0),.clk(gclk));
	jdff dff_B_rEe3ADAP1_0(.din(w_dff_B_F7sHR3l28_0),.dout(w_dff_B_rEe3ADAP1_0),.clk(gclk));
	jdff dff_B_BSFEM9Il6_0(.din(w_dff_B_rEe3ADAP1_0),.dout(w_dff_B_BSFEM9Il6_0),.clk(gclk));
	jdff dff_B_IFjCnL9p5_0(.din(w_dff_B_BSFEM9Il6_0),.dout(w_dff_B_IFjCnL9p5_0),.clk(gclk));
	jdff dff_B_LMyJSMy41_0(.din(n1376),.dout(w_dff_B_LMyJSMy41_0),.clk(gclk));
	jdff dff_B_3YGGGiVE7_2(.din(G173),.dout(w_dff_B_3YGGGiVE7_2),.clk(gclk));
	jdff dff_B_vpfIBe4U6_2(.din(G203),.dout(w_dff_B_vpfIBe4U6_2),.clk(gclk));
	jdff dff_B_sdn6Tn8o5_2(.din(w_dff_B_vpfIBe4U6_2),.dout(w_dff_B_sdn6Tn8o5_2),.clk(gclk));
	jdff dff_B_3DPhSuQZ6_1(.din(n1371),.dout(w_dff_B_3DPhSuQZ6_1),.clk(gclk));
	jdff dff_B_Vx59He5A6_1(.din(w_dff_B_3DPhSuQZ6_1),.dout(w_dff_B_Vx59He5A6_1),.clk(gclk));
	jdff dff_B_kLo2r7RI9_1(.din(w_dff_B_Vx59He5A6_1),.dout(w_dff_B_kLo2r7RI9_1),.clk(gclk));
	jdff dff_B_uAapR5Qn6_1(.din(n1254),.dout(w_dff_B_uAapR5Qn6_1),.clk(gclk));
	jdff dff_B_dPcBdxqo8_1(.din(w_dff_B_uAapR5Qn6_1),.dout(w_dff_B_dPcBdxqo8_1),.clk(gclk));
	jdff dff_B_QuQvfOdS3_1(.din(w_dff_B_dPcBdxqo8_1),.dout(w_dff_B_QuQvfOdS3_1),.clk(gclk));
	jdff dff_B_RixEefj14_1(.din(w_dff_B_QuQvfOdS3_1),.dout(w_dff_B_RixEefj14_1),.clk(gclk));
	jdff dff_B_sbpHS0em0_1(.din(w_dff_B_RixEefj14_1),.dout(w_dff_B_sbpHS0em0_1),.clk(gclk));
	jdff dff_B_b20BfPNH2_1(.din(w_dff_B_sbpHS0em0_1),.dout(w_dff_B_b20BfPNH2_1),.clk(gclk));
	jdff dff_B_sJ9orpA58_1(.din(w_dff_B_b20BfPNH2_1),.dout(w_dff_B_sJ9orpA58_1),.clk(gclk));
	jdff dff_B_AImiS8TP9_1(.din(w_dff_B_sJ9orpA58_1),.dout(w_dff_B_AImiS8TP9_1),.clk(gclk));
	jdff dff_B_oBDNuw0b4_1(.din(w_dff_B_AImiS8TP9_1),.dout(w_dff_B_oBDNuw0b4_1),.clk(gclk));
	jdff dff_B_ZwxUGoIJ7_1(.din(w_dff_B_oBDNuw0b4_1),.dout(w_dff_B_ZwxUGoIJ7_1),.clk(gclk));
	jdff dff_B_5XWr8qUk4_1(.din(w_dff_B_ZwxUGoIJ7_1),.dout(w_dff_B_5XWr8qUk4_1),.clk(gclk));
	jdff dff_B_Ac9kbomT8_1(.din(w_dff_B_5XWr8qUk4_1),.dout(w_dff_B_Ac9kbomT8_1),.clk(gclk));
	jdff dff_B_z39GyPid4_1(.din(w_dff_B_Ac9kbomT8_1),.dout(w_dff_B_z39GyPid4_1),.clk(gclk));
	jdff dff_B_Q9Q1JZKq3_0(.din(n1257),.dout(w_dff_B_Q9Q1JZKq3_0),.clk(gclk));
	jdff dff_B_vfijBjnP6_0(.din(w_dff_B_Q9Q1JZKq3_0),.dout(w_dff_B_vfijBjnP6_0),.clk(gclk));
	jdff dff_B_IdzVWRJ20_0(.din(w_dff_B_vfijBjnP6_0),.dout(w_dff_B_IdzVWRJ20_0),.clk(gclk));
	jdff dff_B_FuLaBeJw9_0(.din(w_dff_B_IdzVWRJ20_0),.dout(w_dff_B_FuLaBeJw9_0),.clk(gclk));
	jdff dff_B_j3URnBDD9_0(.din(w_dff_B_FuLaBeJw9_0),.dout(w_dff_B_j3URnBDD9_0),.clk(gclk));
	jdff dff_B_5ta3wDFs3_0(.din(w_dff_B_j3URnBDD9_0),.dout(w_dff_B_5ta3wDFs3_0),.clk(gclk));
	jdff dff_B_DMhh5lqb8_0(.din(w_dff_B_5ta3wDFs3_0),.dout(w_dff_B_DMhh5lqb8_0),.clk(gclk));
	jdff dff_B_oJEqyHun7_0(.din(w_dff_B_DMhh5lqb8_0),.dout(w_dff_B_oJEqyHun7_0),.clk(gclk));
	jdff dff_B_LvgzSzjn0_0(.din(w_dff_B_oJEqyHun7_0),.dout(w_dff_B_LvgzSzjn0_0),.clk(gclk));
	jdff dff_B_UlI2Nhbz5_1(.din(n500),.dout(w_dff_B_UlI2Nhbz5_1),.clk(gclk));
	jdff dff_B_5spP29TG4_1(.din(n495),.dout(w_dff_B_5spP29TG4_1),.clk(gclk));
	jdff dff_B_rmvr7Zh08_1(.din(G113),.dout(w_dff_B_rmvr7Zh08_1),.clk(gclk));
	jdff dff_B_ZdKFumnR9_1(.din(w_dff_B_rmvr7Zh08_1),.dout(w_dff_B_ZdKFumnR9_1),.clk(gclk));
	jdff dff_A_U6838mNR2_0(.dout(w_n1007_2[0]),.din(w_dff_A_U6838mNR2_0),.clk(gclk));
	jdff dff_A_s7AfrquI6_0(.dout(w_dff_A_U6838mNR2_0),.din(w_dff_A_s7AfrquI6_0),.clk(gclk));
	jdff dff_A_i5S6ZHBl3_0(.dout(w_dff_A_s7AfrquI6_0),.din(w_dff_A_i5S6ZHBl3_0),.clk(gclk));
	jdff dff_A_hhmWvY035_0(.dout(w_dff_A_i5S6ZHBl3_0),.din(w_dff_A_hhmWvY035_0),.clk(gclk));
	jdff dff_A_pMfUvf6u9_0(.dout(w_dff_A_hhmWvY035_0),.din(w_dff_A_pMfUvf6u9_0),.clk(gclk));
	jdff dff_A_MkXZOu1o5_0(.dout(w_dff_A_pMfUvf6u9_0),.din(w_dff_A_MkXZOu1o5_0),.clk(gclk));
	jdff dff_A_FInBIvAe5_1(.dout(w_n1007_2[1]),.din(w_dff_A_FInBIvAe5_1),.clk(gclk));
	jdff dff_B_QsVLWo5M4_1(.din(n1216),.dout(w_dff_B_QsVLWo5M4_1),.clk(gclk));
	jdff dff_B_MLzapeKq4_1(.din(w_dff_B_QsVLWo5M4_1),.dout(w_dff_B_MLzapeKq4_1),.clk(gclk));
	jdff dff_B_egi2egYW9_1(.din(w_dff_B_MLzapeKq4_1),.dout(w_dff_B_egi2egYW9_1),.clk(gclk));
	jdff dff_B_2KP0CUQ02_1(.din(w_dff_B_egi2egYW9_1),.dout(w_dff_B_2KP0CUQ02_1),.clk(gclk));
	jdff dff_B_uV2F0mFV7_1(.din(w_dff_B_2KP0CUQ02_1),.dout(w_dff_B_uV2F0mFV7_1),.clk(gclk));
	jdff dff_B_K3fJ4o1u7_1(.din(w_dff_B_uV2F0mFV7_1),.dout(w_dff_B_K3fJ4o1u7_1),.clk(gclk));
	jdff dff_B_O08tIw8b7_1(.din(w_dff_B_K3fJ4o1u7_1),.dout(w_dff_B_O08tIw8b7_1),.clk(gclk));
	jdff dff_B_g2qFy7mZ6_1(.din(w_dff_B_O08tIw8b7_1),.dout(w_dff_B_g2qFy7mZ6_1),.clk(gclk));
	jdff dff_B_zN12jrPW8_1(.din(w_dff_B_g2qFy7mZ6_1),.dout(w_dff_B_zN12jrPW8_1),.clk(gclk));
	jdff dff_B_xumPm5G10_1(.din(w_dff_B_zN12jrPW8_1),.dout(w_dff_B_xumPm5G10_1),.clk(gclk));
	jdff dff_B_FP9SyRB59_1(.din(w_dff_B_xumPm5G10_1),.dout(w_dff_B_FP9SyRB59_1),.clk(gclk));
	jdff dff_B_ApvnlSWa4_0(.din(n1219),.dout(w_dff_B_ApvnlSWa4_0),.clk(gclk));
	jdff dff_B_AbYxge710_0(.din(w_dff_B_ApvnlSWa4_0),.dout(w_dff_B_AbYxge710_0),.clk(gclk));
	jdff dff_B_NdOS22z31_0(.din(w_dff_B_AbYxge710_0),.dout(w_dff_B_NdOS22z31_0),.clk(gclk));
	jdff dff_B_D2sojhaL3_0(.din(w_dff_B_NdOS22z31_0),.dout(w_dff_B_D2sojhaL3_0),.clk(gclk));
	jdff dff_B_390DoZ1d2_0(.din(w_dff_B_D2sojhaL3_0),.dout(w_dff_B_390DoZ1d2_0),.clk(gclk));
	jdff dff_B_iqFcjq4L1_0(.din(w_dff_B_390DoZ1d2_0),.dout(w_dff_B_iqFcjq4L1_0),.clk(gclk));
	jdff dff_B_GbydITx23_0(.din(w_dff_B_iqFcjq4L1_0),.dout(w_dff_B_GbydITx23_0),.clk(gclk));
	jdff dff_A_gxZKuS240_1(.dout(w_n989_0[1]),.din(w_dff_A_gxZKuS240_1),.clk(gclk));
	jdff dff_A_bVg8zjmE1_1(.dout(w_dff_A_gxZKuS240_1),.din(w_dff_A_bVg8zjmE1_1),.clk(gclk));
	jdff dff_A_VDh4o9zL3_1(.dout(w_dff_A_bVg8zjmE1_1),.din(w_dff_A_VDh4o9zL3_1),.clk(gclk));
	jdff dff_A_ZLXJuPVY7_1(.dout(w_dff_A_VDh4o9zL3_1),.din(w_dff_A_ZLXJuPVY7_1),.clk(gclk));
	jdff dff_A_cgmkJVQL6_1(.dout(w_dff_A_ZLXJuPVY7_1),.din(w_dff_A_cgmkJVQL6_1),.clk(gclk));
	jdff dff_B_MEDCZDtm7_1(.din(n988),.dout(w_dff_B_MEDCZDtm7_1),.clk(gclk));
	jdff dff_B_3ssWQ6XL7_1(.din(w_dff_B_MEDCZDtm7_1),.dout(w_dff_B_3ssWQ6XL7_1),.clk(gclk));
	jdff dff_B_hrULTG3r5_1(.din(w_dff_B_3ssWQ6XL7_1),.dout(w_dff_B_hrULTG3r5_1),.clk(gclk));
	jdff dff_B_DXRqprTM4_1(.din(w_dff_B_hrULTG3r5_1),.dout(w_dff_B_DXRqprTM4_1),.clk(gclk));
	jdff dff_B_ARb2QoPd3_1(.din(w_dff_B_DXRqprTM4_1),.dout(w_dff_B_ARb2QoPd3_1),.clk(gclk));
	jdff dff_B_9D7e0xVP8_1(.din(w_dff_B_ARb2QoPd3_1),.dout(w_dff_B_9D7e0xVP8_1),.clk(gclk));
	jdff dff_B_vtl9k3e31_1(.din(G112),.dout(w_dff_B_vtl9k3e31_1),.clk(gclk));
	jdff dff_B_ppcvgk152_1(.din(w_dff_B_vtl9k3e31_1),.dout(w_dff_B_ppcvgk152_1),.clk(gclk));
	jdff dff_A_LLViKpil3_0(.dout(w_G1691_3[0]),.din(w_dff_A_LLViKpil3_0),.clk(gclk));
	jdff dff_A_VYvhuAvX4_0(.dout(w_dff_A_LLViKpil3_0),.din(w_dff_A_VYvhuAvX4_0),.clk(gclk));
	jdff dff_A_xMrswLls9_0(.dout(w_dff_A_VYvhuAvX4_0),.din(w_dff_A_xMrswLls9_0),.clk(gclk));
	jdff dff_A_TIcULKQy2_0(.dout(w_dff_A_xMrswLls9_0),.din(w_dff_A_TIcULKQy2_0),.clk(gclk));
	jdff dff_A_tSoCaoAp5_1(.dout(w_G1691_3[1]),.din(w_dff_A_tSoCaoAp5_1),.clk(gclk));
	jdff dff_A_AyyJTQSO9_1(.dout(w_dff_A_tSoCaoAp5_1),.din(w_dff_A_AyyJTQSO9_1),.clk(gclk));
	jdff dff_B_p2WWs4dO1_1(.din(n1382),.dout(w_dff_B_p2WWs4dO1_1),.clk(gclk));
	jdff dff_B_hFkVxJ4x7_1(.din(w_dff_B_p2WWs4dO1_1),.dout(w_dff_B_hFkVxJ4x7_1),.clk(gclk));
	jdff dff_B_z9pPafwW7_1(.din(w_dff_B_hFkVxJ4x7_1),.dout(w_dff_B_z9pPafwW7_1),.clk(gclk));
	jdff dff_B_7UeFKED25_1(.din(w_dff_B_z9pPafwW7_1),.dout(w_dff_B_7UeFKED25_1),.clk(gclk));
	jdff dff_B_VKaHcStD9_1(.din(w_dff_B_7UeFKED25_1),.dout(w_dff_B_VKaHcStD9_1),.clk(gclk));
	jdff dff_B_DKncdiQB2_1(.din(w_dff_B_VKaHcStD9_1),.dout(w_dff_B_DKncdiQB2_1),.clk(gclk));
	jdff dff_B_vnDkYqHq3_1(.din(w_dff_B_DKncdiQB2_1),.dout(w_dff_B_vnDkYqHq3_1),.clk(gclk));
	jdff dff_B_WL1pQyqE5_1(.din(w_dff_B_vnDkYqHq3_1),.dout(w_dff_B_WL1pQyqE5_1),.clk(gclk));
	jdff dff_B_cwKcXo590_1(.din(w_dff_B_WL1pQyqE5_1),.dout(w_dff_B_cwKcXo590_1),.clk(gclk));
	jdff dff_B_ATwA34fK2_1(.din(w_dff_B_cwKcXo590_1),.dout(w_dff_B_ATwA34fK2_1),.clk(gclk));
	jdff dff_B_ofV6NNc53_1(.din(w_dff_B_ATwA34fK2_1),.dout(w_dff_B_ofV6NNc53_1),.clk(gclk));
	jdff dff_B_2HI67dHS5_1(.din(w_dff_B_ofV6NNc53_1),.dout(w_dff_B_2HI67dHS5_1),.clk(gclk));
	jdff dff_B_ecLNolU72_1(.din(w_dff_B_2HI67dHS5_1),.dout(w_dff_B_ecLNolU72_1),.clk(gclk));
	jdff dff_B_xtLdzSf50_1(.din(w_dff_B_ecLNolU72_1),.dout(w_dff_B_xtLdzSf50_1),.clk(gclk));
	jdff dff_B_IgSpwvgU3_1(.din(w_dff_B_xtLdzSf50_1),.dout(w_dff_B_IgSpwvgU3_1),.clk(gclk));
	jdff dff_B_iGh2f43X3_1(.din(w_dff_B_IgSpwvgU3_1),.dout(w_dff_B_iGh2f43X3_1),.clk(gclk));
	jdff dff_B_cHymfyTx3_1(.din(w_dff_B_iGh2f43X3_1),.dout(w_dff_B_cHymfyTx3_1),.clk(gclk));
	jdff dff_B_V6AwSBvI4_1(.din(w_dff_B_cHymfyTx3_1),.dout(w_dff_B_V6AwSBvI4_1),.clk(gclk));
	jdff dff_B_dEHTAsTF1_1(.din(w_dff_B_V6AwSBvI4_1),.dout(w_dff_B_dEHTAsTF1_1),.clk(gclk));
	jdff dff_B_6DI3sagl7_1(.din(n1245),.dout(w_dff_B_6DI3sagl7_1),.clk(gclk));
	jdff dff_B_BsGvu4lc8_1(.din(w_dff_B_6DI3sagl7_1),.dout(w_dff_B_BsGvu4lc8_1),.clk(gclk));
	jdff dff_B_GhOkG0605_1(.din(w_dff_B_BsGvu4lc8_1),.dout(w_dff_B_GhOkG0605_1),.clk(gclk));
	jdff dff_B_HXUnzWRY4_1(.din(w_dff_B_GhOkG0605_1),.dout(w_dff_B_HXUnzWRY4_1),.clk(gclk));
	jdff dff_B_gEZPRPo12_1(.din(w_dff_B_HXUnzWRY4_1),.dout(w_dff_B_gEZPRPo12_1),.clk(gclk));
	jdff dff_B_02CnrUPQ5_1(.din(w_dff_B_gEZPRPo12_1),.dout(w_dff_B_02CnrUPQ5_1),.clk(gclk));
	jdff dff_B_hA8dwoGV0_1(.din(w_dff_B_02CnrUPQ5_1),.dout(w_dff_B_hA8dwoGV0_1),.clk(gclk));
	jdff dff_B_WuSlpCqL1_1(.din(w_dff_B_hA8dwoGV0_1),.dout(w_dff_B_WuSlpCqL1_1),.clk(gclk));
	jdff dff_B_2IAefZUF1_1(.din(w_dff_B_WuSlpCqL1_1),.dout(w_dff_B_2IAefZUF1_1),.clk(gclk));
	jdff dff_B_XsGKdWxJ2_1(.din(w_dff_B_2IAefZUF1_1),.dout(w_dff_B_XsGKdWxJ2_1),.clk(gclk));
	jdff dff_B_jPyZcYFn7_1(.din(w_dff_B_XsGKdWxJ2_1),.dout(w_dff_B_jPyZcYFn7_1),.clk(gclk));
	jdff dff_B_2dmljysv7_1(.din(w_dff_B_jPyZcYFn7_1),.dout(w_dff_B_2dmljysv7_1),.clk(gclk));
	jdff dff_B_aVrKJl0A3_1(.din(w_dff_B_2dmljysv7_1),.dout(w_dff_B_aVrKJl0A3_1),.clk(gclk));
	jdff dff_B_TerfcU185_1(.din(w_dff_B_aVrKJl0A3_1),.dout(w_dff_B_TerfcU185_1),.clk(gclk));
	jdff dff_B_HkaWFrb58_1(.din(w_dff_B_TerfcU185_1),.dout(w_dff_B_HkaWFrb58_1),.clk(gclk));
	jdff dff_B_uuDGuNni8_1(.din(w_dff_B_HkaWFrb58_1),.dout(w_dff_B_uuDGuNni8_1),.clk(gclk));
	jdff dff_B_8VGlEAWL1_1(.din(n1247),.dout(w_dff_B_8VGlEAWL1_1),.clk(gclk));
	jdff dff_B_C8xH7zdg3_1(.din(w_dff_B_8VGlEAWL1_1),.dout(w_dff_B_C8xH7zdg3_1),.clk(gclk));
	jdff dff_B_swYH9Qb04_1(.din(w_dff_B_C8xH7zdg3_1),.dout(w_dff_B_swYH9Qb04_1),.clk(gclk));
	jdff dff_B_ISr2g28k4_1(.din(w_dff_B_swYH9Qb04_1),.dout(w_dff_B_ISr2g28k4_1),.clk(gclk));
	jdff dff_B_7CRJ4Ji20_1(.din(w_dff_B_ISr2g28k4_1),.dout(w_dff_B_7CRJ4Ji20_1),.clk(gclk));
	jdff dff_B_eRr7kqYR1_1(.din(w_dff_B_7CRJ4Ji20_1),.dout(w_dff_B_eRr7kqYR1_1),.clk(gclk));
	jdff dff_B_0Zk4YnWz7_1(.din(w_dff_B_eRr7kqYR1_1),.dout(w_dff_B_0Zk4YnWz7_1),.clk(gclk));
	jdff dff_B_KuMbj2xW9_1(.din(w_dff_B_0Zk4YnWz7_1),.dout(w_dff_B_KuMbj2xW9_1),.clk(gclk));
	jdff dff_B_n7YbBHeH6_1(.din(w_dff_B_KuMbj2xW9_1),.dout(w_dff_B_n7YbBHeH6_1),.clk(gclk));
	jdff dff_B_qYFE3t1B0_1(.din(w_dff_B_n7YbBHeH6_1),.dout(w_dff_B_qYFE3t1B0_1),.clk(gclk));
	jdff dff_B_xh3eOoMT7_1(.din(w_dff_B_qYFE3t1B0_1),.dout(w_dff_B_xh3eOoMT7_1),.clk(gclk));
	jdff dff_B_sQBYefKu6_1(.din(n951),.dout(w_dff_B_sQBYefKu6_1),.clk(gclk));
	jdff dff_B_UUPINPiN2_1(.din(w_dff_B_sQBYefKu6_1),.dout(w_dff_B_UUPINPiN2_1),.clk(gclk));
	jdff dff_B_G35Dpjh71_1(.din(w_dff_B_UUPINPiN2_1),.dout(w_dff_B_G35Dpjh71_1),.clk(gclk));
	jdff dff_B_JUdnOlon2_1(.din(w_dff_B_G35Dpjh71_1),.dout(w_dff_B_JUdnOlon2_1),.clk(gclk));
	jdff dff_B_wLOgCkTt1_1(.din(w_dff_B_JUdnOlon2_1),.dout(w_dff_B_wLOgCkTt1_1),.clk(gclk));
	jdff dff_B_x6mYwETw3_1(.din(w_dff_B_wLOgCkTt1_1),.dout(w_dff_B_x6mYwETw3_1),.clk(gclk));
	jdff dff_B_iLjUAyAc7_1(.din(w_dff_B_x6mYwETw3_1),.dout(w_dff_B_iLjUAyAc7_1),.clk(gclk));
	jdff dff_B_4hANBpo36_1(.din(w_dff_B_iLjUAyAc7_1),.dout(w_dff_B_4hANBpo36_1),.clk(gclk));
	jdff dff_B_U77XHhe59_1(.din(w_dff_B_4hANBpo36_1),.dout(w_dff_B_U77XHhe59_1),.clk(gclk));
	jdff dff_B_R5eitxjB8_1(.din(n513),.dout(w_dff_B_R5eitxjB8_1),.clk(gclk));
	jdff dff_B_U8buMZBn5_1(.din(n508),.dout(w_dff_B_U8buMZBn5_1),.clk(gclk));
	jdff dff_B_DgmosfyD2_1(.din(G53),.dout(w_dff_B_DgmosfyD2_1),.clk(gclk));
	jdff dff_B_wPc01Xff2_1(.din(w_dff_B_DgmosfyD2_1),.dout(w_dff_B_wPc01Xff2_1),.clk(gclk));
	jdff dff_B_o4O4XsoW3_1(.din(n1207),.dout(w_dff_B_o4O4XsoW3_1),.clk(gclk));
	jdff dff_B_fh4ifOrf6_1(.din(w_dff_B_o4O4XsoW3_1),.dout(w_dff_B_fh4ifOrf6_1),.clk(gclk));
	jdff dff_B_Rjh3rheS3_1(.din(w_dff_B_fh4ifOrf6_1),.dout(w_dff_B_Rjh3rheS3_1),.clk(gclk));
	jdff dff_B_uMpaWiJB7_1(.din(w_dff_B_Rjh3rheS3_1),.dout(w_dff_B_uMpaWiJB7_1),.clk(gclk));
	jdff dff_B_YCPthgoq9_1(.din(w_dff_B_uMpaWiJB7_1),.dout(w_dff_B_YCPthgoq9_1),.clk(gclk));
	jdff dff_B_bPsVyb8j1_1(.din(w_dff_B_YCPthgoq9_1),.dout(w_dff_B_bPsVyb8j1_1),.clk(gclk));
	jdff dff_B_Fr8ZR9ph3_1(.din(w_dff_B_bPsVyb8j1_1),.dout(w_dff_B_Fr8ZR9ph3_1),.clk(gclk));
	jdff dff_B_in9njksg0_1(.din(w_dff_B_Fr8ZR9ph3_1),.dout(w_dff_B_in9njksg0_1),.clk(gclk));
	jdff dff_B_L1bK1fbl9_1(.din(w_dff_B_in9njksg0_1),.dout(w_dff_B_L1bK1fbl9_1),.clk(gclk));
	jdff dff_B_O0kiAZ539_1(.din(w_dff_B_L1bK1fbl9_1),.dout(w_dff_B_O0kiAZ539_1),.clk(gclk));
	jdff dff_B_odToLabO9_1(.din(w_dff_B_O0kiAZ539_1),.dout(w_dff_B_odToLabO9_1),.clk(gclk));
	jdff dff_B_GWMxj4ZE5_1(.din(w_dff_B_odToLabO9_1),.dout(w_dff_B_GWMxj4ZE5_1),.clk(gclk));
	jdff dff_B_riJkI51u7_1(.din(w_dff_B_GWMxj4ZE5_1),.dout(w_dff_B_riJkI51u7_1),.clk(gclk));
	jdff dff_B_UmXLvvYf4_1(.din(w_dff_B_riJkI51u7_1),.dout(w_dff_B_UmXLvvYf4_1),.clk(gclk));
	jdff dff_B_re8ILEbE4_1(.din(w_dff_B_UmXLvvYf4_1),.dout(w_dff_B_re8ILEbE4_1),.clk(gclk));
	jdff dff_B_0ls9iHpe0_1(.din(w_dff_B_re8ILEbE4_1),.dout(w_dff_B_0ls9iHpe0_1),.clk(gclk));
	jdff dff_B_N5C4SXT00_0(.din(n1211),.dout(w_dff_B_N5C4SXT00_0),.clk(gclk));
	jdff dff_B_PKVlJO5q2_0(.din(w_dff_B_N5C4SXT00_0),.dout(w_dff_B_PKVlJO5q2_0),.clk(gclk));
	jdff dff_B_dBsGJJeR7_0(.din(w_dff_B_PKVlJO5q2_0),.dout(w_dff_B_dBsGJJeR7_0),.clk(gclk));
	jdff dff_B_YIbd9Jui4_0(.din(w_dff_B_dBsGJJeR7_0),.dout(w_dff_B_YIbd9Jui4_0),.clk(gclk));
	jdff dff_B_pivutCvQ4_0(.din(w_dff_B_YIbd9Jui4_0),.dout(w_dff_B_pivutCvQ4_0),.clk(gclk));
	jdff dff_B_KOJPPlSy6_0(.din(w_dff_B_pivutCvQ4_0),.dout(w_dff_B_KOJPPlSy6_0),.clk(gclk));
	jdff dff_B_oO6QsDMN6_0(.din(w_dff_B_KOJPPlSy6_0),.dout(w_dff_B_oO6QsDMN6_0),.clk(gclk));
	jdff dff_B_LNTsN6IM3_0(.din(w_dff_B_oO6QsDMN6_0),.dout(w_dff_B_LNTsN6IM3_0),.clk(gclk));
	jdff dff_B_8HibIQqz7_0(.din(w_dff_B_LNTsN6IM3_0),.dout(w_dff_B_8HibIQqz7_0),.clk(gclk));
	jdff dff_B_K5sujEbX8_0(.din(w_dff_B_8HibIQqz7_0),.dout(w_dff_B_K5sujEbX8_0),.clk(gclk));
	jdff dff_B_toa6koN10_1(.din(n978),.dout(w_dff_B_toa6koN10_1),.clk(gclk));
	jdff dff_B_6soc72gs1_1(.din(w_dff_B_toa6koN10_1),.dout(w_dff_B_6soc72gs1_1),.clk(gclk));
	jdff dff_B_G8Mktwtq9_1(.din(w_dff_B_6soc72gs1_1),.dout(w_dff_B_G8Mktwtq9_1),.clk(gclk));
	jdff dff_B_n1mkz8xW1_1(.din(w_dff_B_G8Mktwtq9_1),.dout(w_dff_B_n1mkz8xW1_1),.clk(gclk));
	jdff dff_B_IqFng8PM3_1(.din(w_dff_B_n1mkz8xW1_1),.dout(w_dff_B_IqFng8PM3_1),.clk(gclk));
	jdff dff_B_6GmatHib3_1(.din(w_dff_B_IqFng8PM3_1),.dout(w_dff_B_6GmatHib3_1),.clk(gclk));
	jdff dff_B_SC9cXjYy2_1(.din(w_dff_B_6GmatHib3_1),.dout(w_dff_B_SC9cXjYy2_1),.clk(gclk));
	jdff dff_B_A7MjYjF48_1(.din(w_dff_B_SC9cXjYy2_1),.dout(w_dff_B_A7MjYjF48_1),.clk(gclk));
	jdff dff_B_evwuM9UD2_1(.din(w_dff_B_A7MjYjF48_1),.dout(w_dff_B_evwuM9UD2_1),.clk(gclk));
	jdff dff_B_0ALb2b7X8_1(.din(n982),.dout(w_dff_B_0ALb2b7X8_1),.clk(gclk));
	jdff dff_B_2RwCbKtr9_1(.din(n980),.dout(w_dff_B_2RwCbKtr9_1),.clk(gclk));
	jdff dff_B_HwRS2yqS1_1(.din(w_dff_B_2RwCbKtr9_1),.dout(w_dff_B_HwRS2yqS1_1),.clk(gclk));
	jdff dff_B_vnzkMDfK1_1(.din(w_dff_B_HwRS2yqS1_1),.dout(w_dff_B_vnzkMDfK1_1),.clk(gclk));
	jdff dff_B_10NKltzk4_1(.din(w_dff_B_vnzkMDfK1_1),.dout(w_dff_B_10NKltzk4_1),.clk(gclk));
	jdff dff_B_N4OMMBhQ3_1(.din(w_dff_B_10NKltzk4_1),.dout(w_dff_B_N4OMMBhQ3_1),.clk(gclk));
	jdff dff_B_Zit3e8cd9_1(.din(G116),.dout(w_dff_B_Zit3e8cd9_1),.clk(gclk));
	jdff dff_B_HLhD5N0M9_1(.din(w_dff_B_Zit3e8cd9_1),.dout(w_dff_B_HLhD5N0M9_1),.clk(gclk));
	jdff dff_B_ijBLdRBO8_0(.din(n1381),.dout(w_dff_B_ijBLdRBO8_0),.clk(gclk));
	jdff dff_B_9aXorsj56_2(.din(G167),.dout(w_dff_B_9aXorsj56_2),.clk(gclk));
	jdff dff_B_H48A0kQm2_2(.din(G197),.dout(w_dff_B_H48A0kQm2_2),.clk(gclk));
	jdff dff_B_VgeiRaJZ6_2(.din(w_dff_B_H48A0kQm2_2),.dout(w_dff_B_VgeiRaJZ6_2),.clk(gclk));
	jdff dff_B_AZvcbzd63_0(.din(n1395),.dout(w_dff_B_AZvcbzd63_0),.clk(gclk));
	jdff dff_B_TkkLXyD15_0(.din(w_dff_B_AZvcbzd63_0),.dout(w_dff_B_TkkLXyD15_0),.clk(gclk));
	jdff dff_B_qqqY8pEI5_0(.din(w_dff_B_TkkLXyD15_0),.dout(w_dff_B_qqqY8pEI5_0),.clk(gclk));
	jdff dff_B_gDRjJvBD3_0(.din(w_dff_B_qqqY8pEI5_0),.dout(w_dff_B_gDRjJvBD3_0),.clk(gclk));
	jdff dff_B_ZVYnWGNU6_0(.din(w_dff_B_gDRjJvBD3_0),.dout(w_dff_B_ZVYnWGNU6_0),.clk(gclk));
	jdff dff_B_cjBEo7AV0_0(.din(w_dff_B_ZVYnWGNU6_0),.dout(w_dff_B_cjBEo7AV0_0),.clk(gclk));
	jdff dff_B_w6xcHZAP3_0(.din(w_dff_B_cjBEo7AV0_0),.dout(w_dff_B_w6xcHZAP3_0),.clk(gclk));
	jdff dff_B_pWYAyKHA0_0(.din(w_dff_B_w6xcHZAP3_0),.dout(w_dff_B_pWYAyKHA0_0),.clk(gclk));
	jdff dff_B_TEqgDbHD6_0(.din(w_dff_B_pWYAyKHA0_0),.dout(w_dff_B_TEqgDbHD6_0),.clk(gclk));
	jdff dff_B_3NlkGlqq2_0(.din(w_dff_B_TEqgDbHD6_0),.dout(w_dff_B_3NlkGlqq2_0),.clk(gclk));
	jdff dff_B_RQas0pJ69_0(.din(w_dff_B_3NlkGlqq2_0),.dout(w_dff_B_RQas0pJ69_0),.clk(gclk));
	jdff dff_B_vU9Gs3iL9_0(.din(w_dff_B_RQas0pJ69_0),.dout(w_dff_B_vU9Gs3iL9_0),.clk(gclk));
	jdff dff_B_uGnDQR4r1_0(.din(w_dff_B_vU9Gs3iL9_0),.dout(w_dff_B_uGnDQR4r1_0),.clk(gclk));
	jdff dff_B_vrEkEr026_0(.din(w_dff_B_uGnDQR4r1_0),.dout(w_dff_B_vrEkEr026_0),.clk(gclk));
	jdff dff_B_iQctaIDJ8_0(.din(w_dff_B_vrEkEr026_0),.dout(w_dff_B_iQctaIDJ8_0),.clk(gclk));
	jdff dff_B_nlPrNay41_0(.din(w_dff_B_iQctaIDJ8_0),.dout(w_dff_B_nlPrNay41_0),.clk(gclk));
	jdff dff_B_EoMrwKBg1_0(.din(w_dff_B_nlPrNay41_0),.dout(w_dff_B_EoMrwKBg1_0),.clk(gclk));
	jdff dff_B_SpQvWwNX4_0(.din(w_dff_B_EoMrwKBg1_0),.dout(w_dff_B_SpQvWwNX4_0),.clk(gclk));
	jdff dff_B_JnaAnNOS8_0(.din(w_dff_B_SpQvWwNX4_0),.dout(w_dff_B_JnaAnNOS8_0),.clk(gclk));
	jdff dff_B_exdElFVE8_0(.din(n1394),.dout(w_dff_B_exdElFVE8_0),.clk(gclk));
	jdff dff_B_TbFIqqaD0_2(.din(G164),.dout(w_dff_B_TbFIqqaD0_2),.clk(gclk));
	jdff dff_B_m7hFPIXg9_2(.din(G194),.dout(w_dff_B_m7hFPIXg9_2),.clk(gclk));
	jdff dff_B_Rz0P6yzV7_2(.din(w_dff_B_m7hFPIXg9_2),.dout(w_dff_B_Rz0P6yzV7_2),.clk(gclk));
	jdff dff_B_ssWr4pTK1_1(.din(n1389),.dout(w_dff_B_ssWr4pTK1_1),.clk(gclk));
	jdff dff_B_yu53a9v41_1(.din(w_dff_B_ssWr4pTK1_1),.dout(w_dff_B_yu53a9v41_1),.clk(gclk));
	jdff dff_B_TGO8iULe2_1(.din(n1239),.dout(w_dff_B_TGO8iULe2_1),.clk(gclk));
	jdff dff_B_A37AbIAp2_1(.din(w_dff_B_TGO8iULe2_1),.dout(w_dff_B_A37AbIAp2_1),.clk(gclk));
	jdff dff_B_wvrreFmq1_1(.din(w_dff_B_A37AbIAp2_1),.dout(w_dff_B_wvrreFmq1_1),.clk(gclk));
	jdff dff_B_KTL9enEE4_1(.din(w_dff_B_wvrreFmq1_1),.dout(w_dff_B_KTL9enEE4_1),.clk(gclk));
	jdff dff_B_v4tyJpsv9_1(.din(w_dff_B_KTL9enEE4_1),.dout(w_dff_B_v4tyJpsv9_1),.clk(gclk));
	jdff dff_B_0IwtZsoK9_1(.din(w_dff_B_v4tyJpsv9_1),.dout(w_dff_B_0IwtZsoK9_1),.clk(gclk));
	jdff dff_B_IfuORuYE1_1(.din(w_dff_B_0IwtZsoK9_1),.dout(w_dff_B_IfuORuYE1_1),.clk(gclk));
	jdff dff_B_bLJBhXpd3_1(.din(w_dff_B_IfuORuYE1_1),.dout(w_dff_B_bLJBhXpd3_1),.clk(gclk));
	jdff dff_B_pbdaXscH8_1(.din(w_dff_B_bLJBhXpd3_1),.dout(w_dff_B_pbdaXscH8_1),.clk(gclk));
	jdff dff_B_34y1FdMT2_1(.din(w_dff_B_pbdaXscH8_1),.dout(w_dff_B_34y1FdMT2_1),.clk(gclk));
	jdff dff_B_RcYZ3R6z5_1(.din(w_dff_B_34y1FdMT2_1),.dout(w_dff_B_RcYZ3R6z5_1),.clk(gclk));
	jdff dff_B_FP5SvLkv9_1(.din(w_dff_B_RcYZ3R6z5_1),.dout(w_dff_B_FP5SvLkv9_1),.clk(gclk));
	jdff dff_B_mHTpKiRG6_1(.din(w_dff_B_FP5SvLkv9_1),.dout(w_dff_B_mHTpKiRG6_1),.clk(gclk));
	jdff dff_B_ko9Gnr9s4_1(.din(w_dff_B_mHTpKiRG6_1),.dout(w_dff_B_ko9Gnr9s4_1),.clk(gclk));
	jdff dff_B_uu31VkD16_0(.din(n1242),.dout(w_dff_B_uu31VkD16_0),.clk(gclk));
	jdff dff_B_vatYfM3q5_0(.din(w_dff_B_uu31VkD16_0),.dout(w_dff_B_vatYfM3q5_0),.clk(gclk));
	jdff dff_B_HTpWDVxP1_0(.din(w_dff_B_vatYfM3q5_0),.dout(w_dff_B_HTpWDVxP1_0),.clk(gclk));
	jdff dff_B_4tC1GQv50_0(.din(w_dff_B_HTpWDVxP1_0),.dout(w_dff_B_4tC1GQv50_0),.clk(gclk));
	jdff dff_B_uwRaskC55_0(.din(w_dff_B_4tC1GQv50_0),.dout(w_dff_B_uwRaskC55_0),.clk(gclk));
	jdff dff_B_FdbOHdph3_0(.din(w_dff_B_uwRaskC55_0),.dout(w_dff_B_FdbOHdph3_0),.clk(gclk));
	jdff dff_B_eC63qPAp6_0(.din(w_dff_B_FdbOHdph3_0),.dout(w_dff_B_eC63qPAp6_0),.clk(gclk));
	jdff dff_B_rvPwzAcj6_0(.din(w_dff_B_eC63qPAp6_0),.dout(w_dff_B_rvPwzAcj6_0),.clk(gclk));
	jdff dff_B_TgL3nZaF8_0(.din(w_dff_B_rvPwzAcj6_0),.dout(w_dff_B_TgL3nZaF8_0),.clk(gclk));
	jdff dff_B_bhsRT5yD6_0(.din(w_dff_B_TgL3nZaF8_0),.dout(w_dff_B_bhsRT5yD6_0),.clk(gclk));
	jdff dff_A_P84LKBiu6_1(.dout(w_n459_0[1]),.din(w_dff_A_P84LKBiu6_1),.clk(gclk));
	jdff dff_A_o8CzVpOe9_1(.dout(w_dff_A_P84LKBiu6_1),.din(w_dff_A_o8CzVpOe9_1),.clk(gclk));
	jdff dff_A_JxHJl6d94_1(.dout(w_dff_A_o8CzVpOe9_1),.din(w_dff_A_JxHJl6d94_1),.clk(gclk));
	jdff dff_B_L640B3lG0_1(.din(n455),.dout(w_dff_B_L640B3lG0_1),.clk(gclk));
	jdff dff_B_qq3Zf2UL4_3(.din(G3548),.dout(w_dff_B_qq3Zf2UL4_3),.clk(gclk));
	jdff dff_B_35rSU6h96_1(.din(n450),.dout(w_dff_B_35rSU6h96_1),.clk(gclk));
	jdff dff_A_n93D60cc3_0(.dout(w_n749_6[0]),.din(w_dff_A_n93D60cc3_0),.clk(gclk));
	jdff dff_A_ie8bqfPa0_0(.dout(w_dff_A_n93D60cc3_0),.din(w_dff_A_ie8bqfPa0_0),.clk(gclk));
	jdff dff_A_IBnOEhUf2_0(.dout(w_dff_A_ie8bqfPa0_0),.din(w_dff_A_IBnOEhUf2_0),.clk(gclk));
	jdff dff_A_a2aQVqUY5_0(.dout(w_dff_A_IBnOEhUf2_0),.din(w_dff_A_a2aQVqUY5_0),.clk(gclk));
	jdff dff_A_yxULFsEi1_0(.dout(w_dff_A_a2aQVqUY5_0),.din(w_dff_A_yxULFsEi1_0),.clk(gclk));
	jdff dff_A_0D4zN2s97_0(.dout(w_dff_A_yxULFsEi1_0),.din(w_dff_A_0D4zN2s97_0),.clk(gclk));
	jdff dff_A_Ds3lcUdV8_0(.dout(w_dff_A_0D4zN2s97_0),.din(w_dff_A_Ds3lcUdV8_0),.clk(gclk));
	jdff dff_A_T2vrZu4X7_0(.dout(w_dff_A_Ds3lcUdV8_0),.din(w_dff_A_T2vrZu4X7_0),.clk(gclk));
	jdff dff_A_Y41NaXej2_0(.dout(w_dff_A_T2vrZu4X7_0),.din(w_dff_A_Y41NaXej2_0),.clk(gclk));
	jdff dff_A_1k0tT0x53_0(.dout(w_dff_A_Y41NaXej2_0),.din(w_dff_A_1k0tT0x53_0),.clk(gclk));
	jdff dff_A_tyqGwJg34_0(.dout(w_dff_A_1k0tT0x53_0),.din(w_dff_A_tyqGwJg34_0),.clk(gclk));
	jdff dff_A_xRxgL4oh5_1(.dout(w_n949_0[1]),.din(w_dff_A_xRxgL4oh5_1),.clk(gclk));
	jdff dff_A_bR7YuVXX4_1(.dout(w_dff_A_xRxgL4oh5_1),.din(w_dff_A_bR7YuVXX4_1),.clk(gclk));
	jdff dff_B_7bcgBnsP3_1(.din(n946),.dout(w_dff_B_7bcgBnsP3_1),.clk(gclk));
	jdff dff_B_8323vT4Z2_1(.din(w_dff_B_7bcgBnsP3_1),.dout(w_dff_B_8323vT4Z2_1),.clk(gclk));
	jdff dff_B_Svcea6JQ3_1(.din(w_dff_B_8323vT4Z2_1),.dout(w_dff_B_Svcea6JQ3_1),.clk(gclk));
	jdff dff_B_G0ca0ANb6_1(.din(w_dff_B_Svcea6JQ3_1),.dout(w_dff_B_G0ca0ANb6_1),.clk(gclk));
	jdff dff_B_sZsrwk6p7_1(.din(w_dff_B_G0ca0ANb6_1),.dout(w_dff_B_sZsrwk6p7_1),.clk(gclk));
	jdff dff_B_pvf6Qcwc9_1(.din(w_dff_B_sZsrwk6p7_1),.dout(w_dff_B_pvf6Qcwc9_1),.clk(gclk));
	jdff dff_A_GsAj6t7L0_0(.dout(w_G4091_2[0]),.din(w_dff_A_GsAj6t7L0_0),.clk(gclk));
	jdff dff_A_hcjprUEn9_0(.dout(w_dff_A_GsAj6t7L0_0),.din(w_dff_A_hcjprUEn9_0),.clk(gclk));
	jdff dff_A_2coFkNWB2_1(.dout(w_G4091_2[1]),.din(w_dff_A_2coFkNWB2_1),.clk(gclk));
	jdff dff_A_tJaTjfpf6_1(.dout(w_dff_A_2coFkNWB2_1),.din(w_dff_A_tJaTjfpf6_1),.clk(gclk));
	jdff dff_A_cF2zdSL49_1(.dout(w_dff_A_tJaTjfpf6_1),.din(w_dff_A_cF2zdSL49_1),.clk(gclk));
	jdff dff_B_nm3ztWNx6_1(.din(G114),.dout(w_dff_B_nm3ztWNx6_1),.clk(gclk));
	jdff dff_B_ceVZ87HC7_1(.din(w_dff_B_nm3ztWNx6_1),.dout(w_dff_B_ceVZ87HC7_1),.clk(gclk));
	jdff dff_A_rrVAIVQh7_0(.dout(w_n1008_2[0]),.din(w_dff_A_rrVAIVQh7_0),.clk(gclk));
	jdff dff_A_YblE7OkE0_1(.dout(w_n1008_2[1]),.din(w_dff_A_YblE7OkE0_1),.clk(gclk));
	jdff dff_B_R2RYqGny3_1(.din(n1198),.dout(w_dff_B_R2RYqGny3_1),.clk(gclk));
	jdff dff_B_MR7DW47J8_1(.din(w_dff_B_R2RYqGny3_1),.dout(w_dff_B_MR7DW47J8_1),.clk(gclk));
	jdff dff_B_e5rhHoLf7_1(.din(w_dff_B_MR7DW47J8_1),.dout(w_dff_B_e5rhHoLf7_1),.clk(gclk));
	jdff dff_B_HBkPwT7n1_1(.din(w_dff_B_e5rhHoLf7_1),.dout(w_dff_B_HBkPwT7n1_1),.clk(gclk));
	jdff dff_B_IPQI8ROY3_1(.din(w_dff_B_HBkPwT7n1_1),.dout(w_dff_B_IPQI8ROY3_1),.clk(gclk));
	jdff dff_B_Zpb95vKL1_1(.din(w_dff_B_IPQI8ROY3_1),.dout(w_dff_B_Zpb95vKL1_1),.clk(gclk));
	jdff dff_B_8pBTZIfu7_1(.din(w_dff_B_Zpb95vKL1_1),.dout(w_dff_B_8pBTZIfu7_1),.clk(gclk));
	jdff dff_B_IiSgUiam6_1(.din(w_dff_B_8pBTZIfu7_1),.dout(w_dff_B_IiSgUiam6_1),.clk(gclk));
	jdff dff_B_4pWTaMZ64_1(.din(w_dff_B_IiSgUiam6_1),.dout(w_dff_B_4pWTaMZ64_1),.clk(gclk));
	jdff dff_B_SfhaCR7j1_1(.din(w_dff_B_4pWTaMZ64_1),.dout(w_dff_B_SfhaCR7j1_1),.clk(gclk));
	jdff dff_B_QzW38vyZ3_1(.din(w_dff_B_SfhaCR7j1_1),.dout(w_dff_B_QzW38vyZ3_1),.clk(gclk));
	jdff dff_B_2MEIc2nO8_1(.din(w_dff_B_QzW38vyZ3_1),.dout(w_dff_B_2MEIc2nO8_1),.clk(gclk));
	jdff dff_B_bCxMWUCL1_1(.din(w_dff_B_2MEIc2nO8_1),.dout(w_dff_B_bCxMWUCL1_1),.clk(gclk));
	jdff dff_B_wYoQnzWD0_1(.din(w_dff_B_bCxMWUCL1_1),.dout(w_dff_B_wYoQnzWD0_1),.clk(gclk));
	jdff dff_B_UUBNS6RN1_1(.din(w_dff_B_wYoQnzWD0_1),.dout(w_dff_B_UUBNS6RN1_1),.clk(gclk));
	jdff dff_B_yO9CgMGc9_1(.din(n1200),.dout(w_dff_B_yO9CgMGc9_1),.clk(gclk));
	jdff dff_B_sRx4mkvJ4_1(.din(w_dff_B_yO9CgMGc9_1),.dout(w_dff_B_sRx4mkvJ4_1),.clk(gclk));
	jdff dff_B_D9MUkGsy8_1(.din(w_dff_B_sRx4mkvJ4_1),.dout(w_dff_B_D9MUkGsy8_1),.clk(gclk));
	jdff dff_B_ZoKDbdFU1_1(.din(w_dff_B_D9MUkGsy8_1),.dout(w_dff_B_ZoKDbdFU1_1),.clk(gclk));
	jdff dff_B_m6Kw7pPu6_1(.din(w_dff_B_ZoKDbdFU1_1),.dout(w_dff_B_m6Kw7pPu6_1),.clk(gclk));
	jdff dff_B_8tMERvoy0_1(.din(w_dff_B_m6Kw7pPu6_1),.dout(w_dff_B_8tMERvoy0_1),.clk(gclk));
	jdff dff_B_qeSXmeGi5_1(.din(w_dff_B_8tMERvoy0_1),.dout(w_dff_B_qeSXmeGi5_1),.clk(gclk));
	jdff dff_B_RuRPskcX9_1(.din(w_dff_B_qeSXmeGi5_1),.dout(w_dff_B_RuRPskcX9_1),.clk(gclk));
	jdff dff_B_56tmRObt7_1(.din(w_dff_B_RuRPskcX9_1),.dout(w_dff_B_56tmRObt7_1),.clk(gclk));
	jdff dff_B_3RbHRXTT8_1(.din(w_dff_B_56tmRObt7_1),.dout(w_dff_B_3RbHRXTT8_1),.clk(gclk));
	jdff dff_B_dOvBVwnH4_1(.din(w_dff_B_3RbHRXTT8_1),.dout(w_dff_B_dOvBVwnH4_1),.clk(gclk));
	jdff dff_A_MQ68W1B17_0(.dout(w_n649_0[0]),.din(w_dff_A_MQ68W1B17_0),.clk(gclk));
	jdff dff_A_xrfi6bE16_0(.dout(w_dff_A_MQ68W1B17_0),.din(w_dff_A_xrfi6bE16_0),.clk(gclk));
	jdff dff_A_2dkfefY57_0(.dout(w_dff_A_xrfi6bE16_0),.din(w_dff_A_2dkfefY57_0),.clk(gclk));
	jdff dff_A_DGoOqOG40_0(.dout(w_dff_A_2dkfefY57_0),.din(w_dff_A_DGoOqOG40_0),.clk(gclk));
	jdff dff_A_spCwRyVo0_0(.dout(w_dff_A_DGoOqOG40_0),.din(w_dff_A_spCwRyVo0_0),.clk(gclk));
	jdff dff_A_gPwATUp97_0(.dout(w_dff_A_spCwRyVo0_0),.din(w_dff_A_gPwATUp97_0),.clk(gclk));
	jdff dff_A_nmgjS8Xb6_0(.dout(w_dff_A_gPwATUp97_0),.din(w_dff_A_nmgjS8Xb6_0),.clk(gclk));
	jdff dff_A_9iMpH7lA9_0(.dout(w_dff_A_nmgjS8Xb6_0),.din(w_dff_A_9iMpH7lA9_0),.clk(gclk));
	jdff dff_A_Jw1AnA3z8_0(.dout(w_dff_A_9iMpH7lA9_0),.din(w_dff_A_Jw1AnA3z8_0),.clk(gclk));
	jdff dff_A_YBqRgmnk3_1(.dout(w_n749_8[1]),.din(w_dff_A_YBqRgmnk3_1),.clk(gclk));
	jdff dff_A_uzrKeSt25_1(.dout(w_dff_A_YBqRgmnk3_1),.din(w_dff_A_uzrKeSt25_1),.clk(gclk));
	jdff dff_A_8DU6gyBa5_1(.dout(w_dff_A_uzrKeSt25_1),.din(w_dff_A_8DU6gyBa5_1),.clk(gclk));
	jdff dff_A_Kx58S53e5_1(.dout(w_dff_A_8DU6gyBa5_1),.din(w_dff_A_Kx58S53e5_1),.clk(gclk));
	jdff dff_A_jayGZ5ID5_1(.dout(w_dff_A_Kx58S53e5_1),.din(w_dff_A_jayGZ5ID5_1),.clk(gclk));
	jdff dff_A_l4lB1dYV0_1(.dout(w_dff_A_jayGZ5ID5_1),.din(w_dff_A_l4lB1dYV0_1),.clk(gclk));
	jdff dff_A_UqJoYVA22_1(.dout(w_dff_A_l4lB1dYV0_1),.din(w_dff_A_UqJoYVA22_1),.clk(gclk));
	jdff dff_A_Cj6H1oYe1_1(.dout(w_dff_A_UqJoYVA22_1),.din(w_dff_A_Cj6H1oYe1_1),.clk(gclk));
	jdff dff_A_ahJjgRGn7_1(.dout(w_dff_A_Cj6H1oYe1_1),.din(w_dff_A_ahJjgRGn7_1),.clk(gclk));
	jdff dff_A_ymixlnCm8_1(.dout(w_dff_A_ahJjgRGn7_1),.din(w_dff_A_ymixlnCm8_1),.clk(gclk));
	jdff dff_A_LYRoVFOK4_1(.dout(w_dff_A_ymixlnCm8_1),.din(w_dff_A_LYRoVFOK4_1),.clk(gclk));
	jdff dff_A_mE7r4Qpk6_1(.dout(w_dff_A_LYRoVFOK4_1),.din(w_dff_A_mE7r4Qpk6_1),.clk(gclk));
	jdff dff_A_8PseJUOO5_2(.dout(w_n749_8[2]),.din(w_dff_A_8PseJUOO5_2),.clk(gclk));
	jdff dff_A_SObhG7m44_2(.dout(w_dff_A_8PseJUOO5_2),.din(w_dff_A_SObhG7m44_2),.clk(gclk));
	jdff dff_A_q08o9JDc0_2(.dout(w_dff_A_SObhG7m44_2),.din(w_dff_A_q08o9JDc0_2),.clk(gclk));
	jdff dff_A_gO0CZgDl3_2(.dout(w_dff_A_q08o9JDc0_2),.din(w_dff_A_gO0CZgDl3_2),.clk(gclk));
	jdff dff_A_syD6FuEI1_2(.dout(w_dff_A_gO0CZgDl3_2),.din(w_dff_A_syD6FuEI1_2),.clk(gclk));
	jdff dff_A_isFRQLDD7_2(.dout(w_dff_A_syD6FuEI1_2),.din(w_dff_A_isFRQLDD7_2),.clk(gclk));
	jdff dff_A_Q8g3bbiG9_2(.dout(w_dff_A_isFRQLDD7_2),.din(w_dff_A_Q8g3bbiG9_2),.clk(gclk));
	jdff dff_A_SITtjx9A9_2(.dout(w_dff_A_Q8g3bbiG9_2),.din(w_dff_A_SITtjx9A9_2),.clk(gclk));
	jdff dff_A_SEsZpSUG7_2(.dout(w_dff_A_SITtjx9A9_2),.din(w_dff_A_SEsZpSUG7_2),.clk(gclk));
	jdff dff_A_uj6YHgjT6_2(.dout(w_dff_A_SEsZpSUG7_2),.din(w_dff_A_uj6YHgjT6_2),.clk(gclk));
	jdff dff_B_GqNr4VAu7_1(.din(G121),.dout(w_dff_B_GqNr4VAu7_1),.clk(gclk));
	jdff dff_B_QiPIzaLg1_1(.din(w_dff_B_GqNr4VAu7_1),.dout(w_dff_B_QiPIzaLg1_1),.clk(gclk));
	jdff dff_A_8GZwz2KJ3_0(.dout(w_G137_4[0]),.din(w_dff_A_8GZwz2KJ3_0),.clk(gclk));
	jdff dff_A_hhdMewAI5_1(.dout(w_G137_4[1]),.din(w_dff_A_hhdMewAI5_1),.clk(gclk));
	jdff dff_A_VIwWP3qT5_0(.dout(w_G137_1[0]),.din(w_dff_A_VIwWP3qT5_0),.clk(gclk));
	jdff dff_A_sutCKZEx3_0(.dout(w_dff_A_VIwWP3qT5_0),.din(w_dff_A_sutCKZEx3_0),.clk(gclk));
	jdff dff_A_hCg5HeLP7_0(.dout(w_dff_A_sutCKZEx3_0),.din(w_dff_A_hCg5HeLP7_0),.clk(gclk));
	jdff dff_A_ksZD6eyg6_0(.dout(w_dff_A_hCg5HeLP7_0),.din(w_dff_A_ksZD6eyg6_0),.clk(gclk));
	jdff dff_A_6UTAXgVo7_0(.dout(w_dff_A_ksZD6eyg6_0),.din(w_dff_A_6UTAXgVo7_0),.clk(gclk));
	jdff dff_A_rhf35aYN2_0(.dout(w_dff_A_6UTAXgVo7_0),.din(w_dff_A_rhf35aYN2_0),.clk(gclk));
	jdff dff_A_SngXMl4h8_1(.dout(w_G137_1[1]),.din(w_dff_A_SngXMl4h8_1),.clk(gclk));
	jdff dff_A_TzB2tQIO0_1(.dout(w_dff_A_SngXMl4h8_1),.din(w_dff_A_TzB2tQIO0_1),.clk(gclk));
	jdff dff_A_zH3xNstB7_1(.dout(w_dff_A_TzB2tQIO0_1),.din(w_dff_A_zH3xNstB7_1),.clk(gclk));
	jdff dff_A_HbGjGKGn8_1(.dout(w_dff_A_zH3xNstB7_1),.din(w_dff_A_HbGjGKGn8_1),.clk(gclk));
	jdff dff_A_HcCFGtfx4_1(.dout(w_dff_A_HbGjGKGn8_1),.din(w_dff_A_HcCFGtfx4_1),.clk(gclk));
	jdff dff_A_1sdCHrTZ4_1(.dout(w_dff_A_HcCFGtfx4_1),.din(w_dff_A_1sdCHrTZ4_1),.clk(gclk));
	jdff dff_A_Wp9ZOKuG8_1(.dout(w_dff_A_1sdCHrTZ4_1),.din(w_dff_A_Wp9ZOKuG8_1),.clk(gclk));
	jdff dff_B_wXvHJvZE3_0(.din(n1404),.dout(w_dff_B_wXvHJvZE3_0),.clk(gclk));
	jdff dff_B_AqoFKCle4_0(.din(w_dff_B_wXvHJvZE3_0),.dout(w_dff_B_AqoFKCle4_0),.clk(gclk));
	jdff dff_B_TdCBwaQ41_0(.din(w_dff_B_AqoFKCle4_0),.dout(w_dff_B_TdCBwaQ41_0),.clk(gclk));
	jdff dff_B_cNU4RuQC6_0(.din(w_dff_B_TdCBwaQ41_0),.dout(w_dff_B_cNU4RuQC6_0),.clk(gclk));
	jdff dff_B_tYY4Xa7D4_0(.din(w_dff_B_cNU4RuQC6_0),.dout(w_dff_B_tYY4Xa7D4_0),.clk(gclk));
	jdff dff_B_YS5Rfacl9_0(.din(w_dff_B_tYY4Xa7D4_0),.dout(w_dff_B_YS5Rfacl9_0),.clk(gclk));
	jdff dff_B_g8mgNMtr4_0(.din(w_dff_B_YS5Rfacl9_0),.dout(w_dff_B_g8mgNMtr4_0),.clk(gclk));
	jdff dff_B_6oMTsNTo3_0(.din(w_dff_B_g8mgNMtr4_0),.dout(w_dff_B_6oMTsNTo3_0),.clk(gclk));
	jdff dff_B_VaYnM2Jn2_0(.din(w_dff_B_6oMTsNTo3_0),.dout(w_dff_B_VaYnM2Jn2_0),.clk(gclk));
	jdff dff_B_w9OQaKfF7_0(.din(w_dff_B_VaYnM2Jn2_0),.dout(w_dff_B_w9OQaKfF7_0),.clk(gclk));
	jdff dff_B_Y1szM2d48_0(.din(w_dff_B_w9OQaKfF7_0),.dout(w_dff_B_Y1szM2d48_0),.clk(gclk));
	jdff dff_B_EVacmhTY0_0(.din(w_dff_B_Y1szM2d48_0),.dout(w_dff_B_EVacmhTY0_0),.clk(gclk));
	jdff dff_B_FhzvEcCL1_0(.din(w_dff_B_EVacmhTY0_0),.dout(w_dff_B_FhzvEcCL1_0),.clk(gclk));
	jdff dff_B_xE0Vmuox9_0(.din(w_dff_B_FhzvEcCL1_0),.dout(w_dff_B_xE0Vmuox9_0),.clk(gclk));
	jdff dff_B_2r4vXc0i3_0(.din(w_dff_B_xE0Vmuox9_0),.dout(w_dff_B_2r4vXc0i3_0),.clk(gclk));
	jdff dff_B_Bn9goyHr5_0(.din(w_dff_B_2r4vXc0i3_0),.dout(w_dff_B_Bn9goyHr5_0),.clk(gclk));
	jdff dff_B_hWRH1XRT5_0(.din(w_dff_B_Bn9goyHr5_0),.dout(w_dff_B_hWRH1XRT5_0),.clk(gclk));
	jdff dff_B_A70fKCp26_0(.din(w_dff_B_hWRH1XRT5_0),.dout(w_dff_B_A70fKCp26_0),.clk(gclk));
	jdff dff_B_riE1MaDo8_0(.din(w_dff_B_A70fKCp26_0),.dout(w_dff_B_riE1MaDo8_0),.clk(gclk));
	jdff dff_B_RcXC3ijD4_0(.din(n1403),.dout(w_dff_B_RcXC3ijD4_0),.clk(gclk));
	jdff dff_B_6HB1p32S0_2(.din(G161),.dout(w_dff_B_6HB1p32S0_2),.clk(gclk));
	jdff dff_B_hdwEuQoB3_2(.din(G191),.dout(w_dff_B_hdwEuQoB3_2),.clk(gclk));
	jdff dff_B_9a14oI2n7_2(.din(w_dff_B_hdwEuQoB3_2),.dout(w_dff_B_9a14oI2n7_2),.clk(gclk));
	jdff dff_B_YE3uA6j95_1(.din(n1190),.dout(w_dff_B_YE3uA6j95_1),.clk(gclk));
	jdff dff_B_3Yhumh1w7_1(.din(w_dff_B_YE3uA6j95_1),.dout(w_dff_B_3Yhumh1w7_1),.clk(gclk));
	jdff dff_B_X693vMg99_1(.din(w_dff_B_3Yhumh1w7_1),.dout(w_dff_B_X693vMg99_1),.clk(gclk));
	jdff dff_B_ooVjqmHx5_1(.din(w_dff_B_X693vMg99_1),.dout(w_dff_B_ooVjqmHx5_1),.clk(gclk));
	jdff dff_B_T2m38Ivc1_1(.din(w_dff_B_ooVjqmHx5_1),.dout(w_dff_B_T2m38Ivc1_1),.clk(gclk));
	jdff dff_B_FHpWsZqr2_1(.din(w_dff_B_T2m38Ivc1_1),.dout(w_dff_B_FHpWsZqr2_1),.clk(gclk));
	jdff dff_B_OCoJLNfz7_1(.din(w_dff_B_FHpWsZqr2_1),.dout(w_dff_B_OCoJLNfz7_1),.clk(gclk));
	jdff dff_B_pfMAzIb94_1(.din(w_dff_B_OCoJLNfz7_1),.dout(w_dff_B_pfMAzIb94_1),.clk(gclk));
	jdff dff_B_tduQ2zyU3_1(.din(w_dff_B_pfMAzIb94_1),.dout(w_dff_B_tduQ2zyU3_1),.clk(gclk));
	jdff dff_B_QocHKizL4_1(.din(w_dff_B_tduQ2zyU3_1),.dout(w_dff_B_QocHKizL4_1),.clk(gclk));
	jdff dff_B_gP2r9NcX1_1(.din(w_dff_B_QocHKizL4_1),.dout(w_dff_B_gP2r9NcX1_1),.clk(gclk));
	jdff dff_B_IbWYYQrg5_1(.din(w_dff_B_gP2r9NcX1_1),.dout(w_dff_B_IbWYYQrg5_1),.clk(gclk));
	jdff dff_B_1vD3Cpe86_1(.din(w_dff_B_IbWYYQrg5_1),.dout(w_dff_B_1vD3Cpe86_1),.clk(gclk));
	jdff dff_B_gJCNnDqk5_1(.din(w_dff_B_1vD3Cpe86_1),.dout(w_dff_B_gJCNnDqk5_1),.clk(gclk));
	jdff dff_B_wYESkZk22_1(.din(w_dff_B_gJCNnDqk5_1),.dout(w_dff_B_wYESkZk22_1),.clk(gclk));
	jdff dff_B_MwEejZKs4_1(.din(w_dff_B_wYESkZk22_1),.dout(w_dff_B_MwEejZKs4_1),.clk(gclk));
	jdff dff_B_DLl6XSoQ4_0(.din(n1194),.dout(w_dff_B_DLl6XSoQ4_0),.clk(gclk));
	jdff dff_B_goRQgdUe3_0(.din(w_dff_B_DLl6XSoQ4_0),.dout(w_dff_B_goRQgdUe3_0),.clk(gclk));
	jdff dff_B_PRlc2US79_0(.din(w_dff_B_goRQgdUe3_0),.dout(w_dff_B_PRlc2US79_0),.clk(gclk));
	jdff dff_B_QBrcBN801_0(.din(w_dff_B_PRlc2US79_0),.dout(w_dff_B_QBrcBN801_0),.clk(gclk));
	jdff dff_B_G0YE7U8x1_0(.din(w_dff_B_QBrcBN801_0),.dout(w_dff_B_G0YE7U8x1_0),.clk(gclk));
	jdff dff_B_JAlnbApl7_0(.din(w_dff_B_G0YE7U8x1_0),.dout(w_dff_B_JAlnbApl7_0),.clk(gclk));
	jdff dff_B_rBBPpyKu4_0(.din(w_dff_B_JAlnbApl7_0),.dout(w_dff_B_rBBPpyKu4_0),.clk(gclk));
	jdff dff_B_XKiMiVu94_0(.din(w_dff_B_rBBPpyKu4_0),.dout(w_dff_B_XKiMiVu94_0),.clk(gclk));
	jdff dff_B_OET0gN4x9_0(.din(w_dff_B_XKiMiVu94_0),.dout(w_dff_B_OET0gN4x9_0),.clk(gclk));
	jdff dff_B_Qe4Fzh8e1_0(.din(w_dff_B_OET0gN4x9_0),.dout(w_dff_B_Qe4Fzh8e1_0),.clk(gclk));
	jdff dff_B_JtQRx7758_0(.din(w_dff_B_Qe4Fzh8e1_0),.dout(w_dff_B_JtQRx7758_0),.clk(gclk));
	jdff dff_B_uUfT9kX12_0(.din(w_dff_B_JtQRx7758_0),.dout(w_dff_B_uUfT9kX12_0),.clk(gclk));
	jdff dff_A_iTx9WcG79_1(.dout(w_G4092_6[1]),.din(w_dff_A_iTx9WcG79_1),.clk(gclk));
	jdff dff_A_mBnuKcvg5_1(.dout(w_dff_A_iTx9WcG79_1),.din(w_dff_A_mBnuKcvg5_1),.clk(gclk));
	jdff dff_A_94ZwdcIq1_2(.dout(w_G4092_6[2]),.din(w_dff_A_94ZwdcIq1_2),.clk(gclk));
	jdff dff_A_naL09aep2_2(.dout(w_dff_A_94ZwdcIq1_2),.din(w_dff_A_naL09aep2_2),.clk(gclk));
	jdff dff_B_uoWfeqFs0_0(.din(n794),.dout(w_dff_B_uoWfeqFs0_0),.clk(gclk));
	jdff dff_B_vcCWrcpf7_0(.din(n785),.dout(w_dff_B_vcCWrcpf7_0),.clk(gclk));
	jdff dff_A_CGCniSRM1_0(.dout(w_G54_0[0]),.din(w_dff_A_CGCniSRM1_0),.clk(gclk));
	jdff dff_A_3XKYABDM8_0(.dout(w_dff_A_CGCniSRM1_0),.din(w_dff_A_3XKYABDM8_0),.clk(gclk));
	jdff dff_A_CzTllBbM8_0(.dout(w_dff_A_3XKYABDM8_0),.din(w_dff_A_CzTllBbM8_0),.clk(gclk));
	jdff dff_A_BHwiBTuq5_0(.dout(w_dff_A_CzTllBbM8_0),.din(w_dff_A_BHwiBTuq5_0),.clk(gclk));
	jdff dff_A_Mu4bqUEB1_0(.dout(w_dff_A_BHwiBTuq5_0),.din(w_dff_A_Mu4bqUEB1_0),.clk(gclk));
	jdff dff_A_x1a6zmGF5_0(.dout(w_dff_A_Mu4bqUEB1_0),.din(w_dff_A_x1a6zmGF5_0),.clk(gclk));
	jdff dff_A_Q3rVDNb76_0(.dout(w_dff_A_x1a6zmGF5_0),.din(w_dff_A_Q3rVDNb76_0),.clk(gclk));
	jdff dff_A_xx0NPEfj7_0(.dout(w_dff_A_Q3rVDNb76_0),.din(w_dff_A_xx0NPEfj7_0),.clk(gclk));
	jdff dff_A_DMJLjAWC3_0(.dout(w_dff_A_xx0NPEfj7_0),.din(w_dff_A_DMJLjAWC3_0),.clk(gclk));
	jdff dff_A_cJWklolw2_1(.dout(w_G54_0[1]),.din(w_dff_A_cJWklolw2_1),.clk(gclk));
	jdff dff_A_F7ldFdBy6_1(.dout(w_dff_A_cJWklolw2_1),.din(w_dff_A_F7ldFdBy6_1),.clk(gclk));
	jdff dff_A_rKJw0v9g3_1(.dout(w_dff_A_F7ldFdBy6_1),.din(w_dff_A_rKJw0v9g3_1),.clk(gclk));
	jdff dff_A_pnV8RWif9_1(.dout(w_dff_A_rKJw0v9g3_1),.din(w_dff_A_pnV8RWif9_1),.clk(gclk));
	jdff dff_A_6uXU1W2I7_0(.dout(w_n749_9[0]),.din(w_dff_A_6uXU1W2I7_0),.clk(gclk));
	jdff dff_A_tLZXFnJW9_2(.dout(w_n749_9[2]),.din(w_dff_A_tLZXFnJW9_2),.clk(gclk));
	jdff dff_A_xNE3xJgf3_2(.dout(w_dff_A_tLZXFnJW9_2),.din(w_dff_A_xNE3xJgf3_2),.clk(gclk));
	jdff dff_A_9nmSpktc8_2(.dout(w_dff_A_xNE3xJgf3_2),.din(w_dff_A_9nmSpktc8_2),.clk(gclk));
	jdff dff_A_CKzamNTm1_2(.dout(w_dff_A_9nmSpktc8_2),.din(w_dff_A_CKzamNTm1_2),.clk(gclk));
	jdff dff_A_LcIwscl35_2(.dout(w_dff_A_CKzamNTm1_2),.din(w_dff_A_LcIwscl35_2),.clk(gclk));
	jdff dff_A_QYuWKXTJ8_2(.dout(w_dff_A_LcIwscl35_2),.din(w_dff_A_QYuWKXTJ8_2),.clk(gclk));
	jdff dff_A_A3LVXdBy9_2(.dout(w_dff_A_QYuWKXTJ8_2),.din(w_dff_A_A3LVXdBy9_2),.clk(gclk));
	jdff dff_A_paLvKvVC2_2(.dout(w_dff_A_A3LVXdBy9_2),.din(w_dff_A_paLvKvVC2_2),.clk(gclk));
	jdff dff_A_5dsmW2Lf1_2(.dout(w_dff_A_paLvKvVC2_2),.din(w_dff_A_5dsmW2Lf1_2),.clk(gclk));
	jdff dff_A_RGEdYACW1_2(.dout(w_dff_A_5dsmW2Lf1_2),.din(w_dff_A_RGEdYACW1_2),.clk(gclk));
	jdff dff_A_soXo7ihW1_2(.dout(w_dff_A_RGEdYACW1_2),.din(w_dff_A_soXo7ihW1_2),.clk(gclk));
	jdff dff_A_JIgpSfBy7_2(.dout(w_dff_A_soXo7ihW1_2),.din(w_dff_A_JIgpSfBy7_2),.clk(gclk));
	jdff dff_A_wJQXwZ5L1_2(.dout(w_dff_A_JIgpSfBy7_2),.din(w_dff_A_wJQXwZ5L1_2),.clk(gclk));
	jdff dff_A_9Sq3Quiw6_2(.dout(w_dff_A_wJQXwZ5L1_2),.din(w_dff_A_9Sq3Quiw6_2),.clk(gclk));
	jdff dff_A_aufjJL5v8_0(.dout(w_G123_0[0]),.din(w_dff_A_aufjJL5v8_0),.clk(gclk));
	jdff dff_A_nINmy0MP3_0(.dout(w_dff_A_aufjJL5v8_0),.din(w_dff_A_nINmy0MP3_0),.clk(gclk));
	jdff dff_A_tKb3P4l32_0(.dout(w_G1691_2[0]),.din(w_dff_A_tKb3P4l32_0),.clk(gclk));
	jdff dff_A_XGBsZiXQ1_2(.dout(w_G1691_2[2]),.din(w_dff_A_XGBsZiXQ1_2),.clk(gclk));
	jdff dff_A_ympCL9KT2_2(.dout(w_n1007_1[2]),.din(w_dff_A_ympCL9KT2_2),.clk(gclk));
	jdff dff_A_0EfxXLcI0_0(.dout(w_n1007_0[0]),.din(w_dff_A_0EfxXLcI0_0),.clk(gclk));
	jdff dff_A_gz7mNcrP8_0(.dout(w_dff_A_0EfxXLcI0_0),.din(w_dff_A_gz7mNcrP8_0),.clk(gclk));
	jdff dff_A_EXz1UC2q5_0(.dout(w_dff_A_gz7mNcrP8_0),.din(w_dff_A_EXz1UC2q5_0),.clk(gclk));
	jdff dff_A_Wr3c9Y7C9_0(.dout(w_dff_A_EXz1UC2q5_0),.din(w_dff_A_Wr3c9Y7C9_0),.clk(gclk));
	jdff dff_A_Qlxb89eu8_0(.dout(w_dff_A_Wr3c9Y7C9_0),.din(w_dff_A_Qlxb89eu8_0),.clk(gclk));
	jdff dff_A_uuMJeVJz7_0(.dout(w_dff_A_Qlxb89eu8_0),.din(w_dff_A_uuMJeVJz7_0),.clk(gclk));
	jdff dff_A_DPtnB4aD3_0(.dout(w_dff_A_uuMJeVJz7_0),.din(w_dff_A_DPtnB4aD3_0),.clk(gclk));
	jdff dff_A_oOqJZCNw0_0(.dout(w_dff_A_DPtnB4aD3_0),.din(w_dff_A_oOqJZCNw0_0),.clk(gclk));
	jdff dff_A_1grDYaM51_0(.dout(w_dff_A_oOqJZCNw0_0),.din(w_dff_A_1grDYaM51_0),.clk(gclk));
	jdff dff_A_jAzl1Tul2_1(.dout(w_n1007_0[1]),.din(w_dff_A_jAzl1Tul2_1),.clk(gclk));
	jdff dff_A_DLqRDtDr1_1(.dout(w_dff_A_jAzl1Tul2_1),.din(w_dff_A_DLqRDtDr1_1),.clk(gclk));
	jdff dff_B_I8dQ9LZl8_3(.din(n1007),.dout(w_dff_B_I8dQ9LZl8_3),.clk(gclk));
	jdff dff_B_LPjgQV3R1_3(.din(w_dff_B_I8dQ9LZl8_3),.dout(w_dff_B_LPjgQV3R1_3),.clk(gclk));
	jdff dff_B_qJKGc85C8_3(.din(w_dff_B_LPjgQV3R1_3),.dout(w_dff_B_qJKGc85C8_3),.clk(gclk));
	jdff dff_B_TsyjQJph9_3(.din(w_dff_B_qJKGc85C8_3),.dout(w_dff_B_TsyjQJph9_3),.clk(gclk));
	jdff dff_B_XtQIU3YD6_3(.din(w_dff_B_TsyjQJph9_3),.dout(w_dff_B_XtQIU3YD6_3),.clk(gclk));
	jdff dff_B_sejIwKca4_3(.din(w_dff_B_XtQIU3YD6_3),.dout(w_dff_B_sejIwKca4_3),.clk(gclk));
	jdff dff_B_sFIaZoQx5_3(.din(w_dff_B_sejIwKca4_3),.dout(w_dff_B_sFIaZoQx5_3),.clk(gclk));
	jdff dff_B_bIbi6GKC1_3(.din(w_dff_B_sFIaZoQx5_3),.dout(w_dff_B_bIbi6GKC1_3),.clk(gclk));
	jdff dff_B_TCpHyeD96_3(.din(w_dff_B_bIbi6GKC1_3),.dout(w_dff_B_TCpHyeD96_3),.clk(gclk));
	jdff dff_B_cROi7K2p8_3(.din(w_dff_B_TCpHyeD96_3),.dout(w_dff_B_cROi7K2p8_3),.clk(gclk));
	jdff dff_B_hRGElnj35_3(.din(w_dff_B_cROi7K2p8_3),.dout(w_dff_B_hRGElnj35_3),.clk(gclk));
	jdff dff_B_amyy1rbg2_1(.din(n1230),.dout(w_dff_B_amyy1rbg2_1),.clk(gclk));
	jdff dff_B_uImP2r9Y7_1(.din(w_dff_B_amyy1rbg2_1),.dout(w_dff_B_uImP2r9Y7_1),.clk(gclk));
	jdff dff_B_QA83R6Zu0_1(.din(w_dff_B_uImP2r9Y7_1),.dout(w_dff_B_QA83R6Zu0_1),.clk(gclk));
	jdff dff_B_eNf6nigZ6_1(.din(w_dff_B_QA83R6Zu0_1),.dout(w_dff_B_eNf6nigZ6_1),.clk(gclk));
	jdff dff_B_gL4Z7yot5_1(.din(w_dff_B_eNf6nigZ6_1),.dout(w_dff_B_gL4Z7yot5_1),.clk(gclk));
	jdff dff_B_bI5pD3sw3_1(.din(w_dff_B_gL4Z7yot5_1),.dout(w_dff_B_bI5pD3sw3_1),.clk(gclk));
	jdff dff_B_CyLly1rx7_1(.din(w_dff_B_bI5pD3sw3_1),.dout(w_dff_B_CyLly1rx7_1),.clk(gclk));
	jdff dff_B_CH6wZtSF9_1(.din(w_dff_B_CyLly1rx7_1),.dout(w_dff_B_CH6wZtSF9_1),.clk(gclk));
	jdff dff_B_lH0bQREE9_1(.din(w_dff_B_CH6wZtSF9_1),.dout(w_dff_B_lH0bQREE9_1),.clk(gclk));
	jdff dff_B_27bVFTkF2_1(.din(w_dff_B_lH0bQREE9_1),.dout(w_dff_B_27bVFTkF2_1),.clk(gclk));
	jdff dff_B_2YTQ9NR07_1(.din(w_dff_B_27bVFTkF2_1),.dout(w_dff_B_2YTQ9NR07_1),.clk(gclk));
	jdff dff_B_lZULK1WQ3_1(.din(w_dff_B_2YTQ9NR07_1),.dout(w_dff_B_lZULK1WQ3_1),.clk(gclk));
	jdff dff_B_8KE7QGNS8_1(.din(w_dff_B_lZULK1WQ3_1),.dout(w_dff_B_8KE7QGNS8_1),.clk(gclk));
	jdff dff_B_ePxNtX9s6_1(.din(w_dff_B_8KE7QGNS8_1),.dout(w_dff_B_ePxNtX9s6_1),.clk(gclk));
	jdff dff_B_ztTiXgTH8_1(.din(w_dff_B_ePxNtX9s6_1),.dout(w_dff_B_ztTiXgTH8_1),.clk(gclk));
	jdff dff_B_B4WLClEx0_1(.din(w_dff_B_ztTiXgTH8_1),.dout(w_dff_B_B4WLClEx0_1),.clk(gclk));
	jdff dff_B_bNSu0CbU2_1(.din(w_dff_B_B4WLClEx0_1),.dout(w_dff_B_bNSu0CbU2_1),.clk(gclk));
	jdff dff_B_jwehbJPO4_1(.din(n1232),.dout(w_dff_B_jwehbJPO4_1),.clk(gclk));
	jdff dff_B_0Vs4H8rV0_1(.din(w_dff_B_jwehbJPO4_1),.dout(w_dff_B_0Vs4H8rV0_1),.clk(gclk));
	jdff dff_B_wqEGCKr88_1(.din(w_dff_B_0Vs4H8rV0_1),.dout(w_dff_B_wqEGCKr88_1),.clk(gclk));
	jdff dff_B_DicT3vzA4_1(.din(w_dff_B_wqEGCKr88_1),.dout(w_dff_B_DicT3vzA4_1),.clk(gclk));
	jdff dff_B_9saAF3tT4_1(.din(w_dff_B_DicT3vzA4_1),.dout(w_dff_B_9saAF3tT4_1),.clk(gclk));
	jdff dff_B_gxf9qsTh2_1(.din(w_dff_B_9saAF3tT4_1),.dout(w_dff_B_gxf9qsTh2_1),.clk(gclk));
	jdff dff_B_p0a6wSf96_1(.din(w_dff_B_gxf9qsTh2_1),.dout(w_dff_B_p0a6wSf96_1),.clk(gclk));
	jdff dff_B_LzIyNZfT0_1(.din(w_dff_B_p0a6wSf96_1),.dout(w_dff_B_LzIyNZfT0_1),.clk(gclk));
	jdff dff_B_AtBHc7Nr5_1(.din(w_dff_B_LzIyNZfT0_1),.dout(w_dff_B_AtBHc7Nr5_1),.clk(gclk));
	jdff dff_B_7wsLq0fn9_1(.din(w_dff_B_AtBHc7Nr5_1),.dout(w_dff_B_7wsLq0fn9_1),.clk(gclk));
	jdff dff_B_CrdZCWz15_1(.din(w_dff_B_7wsLq0fn9_1),.dout(w_dff_B_CrdZCWz15_1),.clk(gclk));
	jdff dff_B_zNX5cKln3_1(.din(w_dff_B_CrdZCWz15_1),.dout(w_dff_B_zNX5cKln3_1),.clk(gclk));
	jdff dff_B_RHDk62kT6_1(.din(n937),.dout(w_dff_B_RHDk62kT6_1),.clk(gclk));
	jdff dff_B_FlKAU1g28_1(.din(w_dff_B_RHDk62kT6_1),.dout(w_dff_B_FlKAU1g28_1),.clk(gclk));
	jdff dff_B_c6eV3Lj95_1(.din(w_dff_B_FlKAU1g28_1),.dout(w_dff_B_c6eV3Lj95_1),.clk(gclk));
	jdff dff_B_YZM3O3dE1_1(.din(w_dff_B_c6eV3Lj95_1),.dout(w_dff_B_YZM3O3dE1_1),.clk(gclk));
	jdff dff_B_fyb1ZnLl0_1(.din(w_dff_B_YZM3O3dE1_1),.dout(w_dff_B_fyb1ZnLl0_1),.clk(gclk));
	jdff dff_B_rqQWsDeM4_1(.din(w_dff_B_fyb1ZnLl0_1),.dout(w_dff_B_rqQWsDeM4_1),.clk(gclk));
	jdff dff_B_TsL2Ppb41_1(.din(w_dff_B_rqQWsDeM4_1),.dout(w_dff_B_TsL2Ppb41_1),.clk(gclk));
	jdff dff_B_5E2anqwI9_1(.din(w_dff_B_TsL2Ppb41_1),.dout(w_dff_B_5E2anqwI9_1),.clk(gclk));
	jdff dff_B_cJ47nVtA4_1(.din(w_dff_B_5E2anqwI9_1),.dout(w_dff_B_cJ47nVtA4_1),.clk(gclk));
	jdff dff_B_A4cRV65P7_1(.din(w_dff_B_cJ47nVtA4_1),.dout(w_dff_B_A4cRV65P7_1),.clk(gclk));
	jdff dff_B_Q5gAEA4b4_1(.din(w_dff_B_A4cRV65P7_1),.dout(w_dff_B_Q5gAEA4b4_1),.clk(gclk));
	jdff dff_B_2GHUucvT0_0(.din(n869),.dout(w_dff_B_2GHUucvT0_0),.clk(gclk));
	jdff dff_B_JWZuuTxj3_1(.din(n866),.dout(w_dff_B_JWZuuTxj3_1),.clk(gclk));
	jdff dff_B_SZmFmjq37_1(.din(w_dff_B_JWZuuTxj3_1),.dout(w_dff_B_SZmFmjq37_1),.clk(gclk));
	jdff dff_A_xUQ57v087_1(.dout(w_G4_0[1]),.din(w_dff_A_xUQ57v087_1),.clk(gclk));
	jdff dff_B_hH0ckDwQ5_3(.din(G4),.dout(w_dff_B_hH0ckDwQ5_3),.clk(gclk));
	jdff dff_B_YNp8mRoG2_3(.din(w_dff_B_hH0ckDwQ5_3),.dout(w_dff_B_YNp8mRoG2_3),.clk(gclk));
	jdff dff_B_WEAVzPa68_3(.din(w_dff_B_YNp8mRoG2_3),.dout(w_dff_B_WEAVzPa68_3),.clk(gclk));
	jdff dff_B_Iqy5LW3W3_3(.din(w_dff_B_WEAVzPa68_3),.dout(w_dff_B_Iqy5LW3W3_3),.clk(gclk));
	jdff dff_B_w06pBtwL9_3(.din(w_dff_B_Iqy5LW3W3_3),.dout(w_dff_B_w06pBtwL9_3),.clk(gclk));
	jdff dff_A_4TUwTOi88_0(.dout(w_n1201_0[0]),.din(w_dff_A_4TUwTOi88_0),.clk(gclk));
	jdff dff_A_TLEHEiKi1_1(.dout(w_n1201_0[1]),.din(w_dff_A_TLEHEiKi1_1),.clk(gclk));
	jdff dff_A_k4Mc6obz5_1(.dout(w_dff_A_TLEHEiKi1_1),.din(w_dff_A_k4Mc6obz5_1),.clk(gclk));
	jdff dff_B_cCmWeS6q0_3(.din(n1201),.dout(w_dff_B_cCmWeS6q0_3),.clk(gclk));
	jdff dff_B_c3hkSaUW6_3(.din(w_dff_B_cCmWeS6q0_3),.dout(w_dff_B_c3hkSaUW6_3),.clk(gclk));
	jdff dff_B_uxCjVNF17_3(.din(w_dff_B_c3hkSaUW6_3),.dout(w_dff_B_uxCjVNF17_3),.clk(gclk));
	jdff dff_B_r2cDyF8a9_3(.din(w_dff_B_uxCjVNF17_3),.dout(w_dff_B_r2cDyF8a9_3),.clk(gclk));
	jdff dff_B_cCrJqu9M4_3(.din(w_dff_B_r2cDyF8a9_3),.dout(w_dff_B_cCrJqu9M4_3),.clk(gclk));
	jdff dff_B_3w3pEc0O3_3(.din(w_dff_B_cCrJqu9M4_3),.dout(w_dff_B_3w3pEc0O3_3),.clk(gclk));
	jdff dff_B_Fp8ErwLW8_3(.din(w_dff_B_3w3pEc0O3_3),.dout(w_dff_B_Fp8ErwLW8_3),.clk(gclk));
	jdff dff_B_RNvt37Yl6_3(.din(w_dff_B_Fp8ErwLW8_3),.dout(w_dff_B_RNvt37Yl6_3),.clk(gclk));
	jdff dff_B_214luyp62_3(.din(w_dff_B_RNvt37Yl6_3),.dout(w_dff_B_214luyp62_3),.clk(gclk));
	jdff dff_B_BrGB2khJ2_3(.din(w_dff_B_214luyp62_3),.dout(w_dff_B_BrGB2khJ2_3),.clk(gclk));
	jdff dff_B_VYdMdNZN7_3(.din(w_dff_B_BrGB2khJ2_3),.dout(w_dff_B_VYdMdNZN7_3),.clk(gclk));
	jdff dff_B_nd5VjrdD3_3(.din(w_dff_B_VYdMdNZN7_3),.dout(w_dff_B_nd5VjrdD3_3),.clk(gclk));
	jdff dff_B_1f30x1bG4_3(.din(w_dff_B_nd5VjrdD3_3),.dout(w_dff_B_1f30x1bG4_3),.clk(gclk));
	jdff dff_B_jTDJ0t9Z3_3(.din(w_dff_B_1f30x1bG4_3),.dout(w_dff_B_jTDJ0t9Z3_3),.clk(gclk));
	jdff dff_B_cfmT20Li7_3(.din(w_dff_B_jTDJ0t9Z3_3),.dout(w_dff_B_cfmT20Li7_3),.clk(gclk));
	jdff dff_A_CUy5sQBD5_0(.dout(w_G4092_5[0]),.din(w_dff_A_CUy5sQBD5_0),.clk(gclk));
	jdff dff_A_nexf5sNW3_0(.dout(w_dff_A_CUy5sQBD5_0),.din(w_dff_A_nexf5sNW3_0),.clk(gclk));
	jdff dff_A_eJepZW6A4_0(.dout(w_dff_A_nexf5sNW3_0),.din(w_dff_A_eJepZW6A4_0),.clk(gclk));
	jdff dff_A_uSho9M3r2_0(.dout(w_dff_A_eJepZW6A4_0),.din(w_dff_A_uSho9M3r2_0),.clk(gclk));
	jdff dff_A_G9DbjvMO8_0(.dout(w_dff_A_uSho9M3r2_0),.din(w_dff_A_G9DbjvMO8_0),.clk(gclk));
	jdff dff_A_1EefmUZz0_0(.dout(w_dff_A_G9DbjvMO8_0),.din(w_dff_A_1EefmUZz0_0),.clk(gclk));
	jdff dff_A_zMTya1Hp5_1(.dout(w_G4092_5[1]),.din(w_dff_A_zMTya1Hp5_1),.clk(gclk));
	jdff dff_A_MtmE4Kbw7_1(.dout(w_dff_A_zMTya1Hp5_1),.din(w_dff_A_MtmE4Kbw7_1),.clk(gclk));
	jdff dff_A_BUWK75vh2_1(.dout(w_dff_A_MtmE4Kbw7_1),.din(w_dff_A_BUWK75vh2_1),.clk(gclk));
	jdff dff_A_zvXr6Mlm4_1(.dout(w_dff_A_BUWK75vh2_1),.din(w_dff_A_zvXr6Mlm4_1),.clk(gclk));
	jdff dff_A_elzg1mGC6_1(.dout(w_dff_A_zvXr6Mlm4_1),.din(w_dff_A_elzg1mGC6_1),.clk(gclk));
	jdff dff_A_ggjRFm5I5_1(.dout(w_dff_A_elzg1mGC6_1),.din(w_dff_A_ggjRFm5I5_1),.clk(gclk));
	jdff dff_A_TrhiBh0t8_0(.dout(w_n749_7[0]),.din(w_dff_A_TrhiBh0t8_0),.clk(gclk));
	jdff dff_A_YV7CwGLn4_0(.dout(w_dff_A_TrhiBh0t8_0),.din(w_dff_A_YV7CwGLn4_0),.clk(gclk));
	jdff dff_A_MpHDPtHA6_0(.dout(w_dff_A_YV7CwGLn4_0),.din(w_dff_A_MpHDPtHA6_0),.clk(gclk));
	jdff dff_A_nGAJWrGH3_0(.dout(w_dff_A_MpHDPtHA6_0),.din(w_dff_A_nGAJWrGH3_0),.clk(gclk));
	jdff dff_A_SgjoVAQz5_0(.dout(w_dff_A_nGAJWrGH3_0),.din(w_dff_A_SgjoVAQz5_0),.clk(gclk));
	jdff dff_A_reBStM3D9_0(.dout(w_dff_A_SgjoVAQz5_0),.din(w_dff_A_reBStM3D9_0),.clk(gclk));
	jdff dff_A_UuKmZWsm8_0(.dout(w_dff_A_reBStM3D9_0),.din(w_dff_A_UuKmZWsm8_0),.clk(gclk));
	jdff dff_A_Xln8IGVO3_0(.dout(w_dff_A_UuKmZWsm8_0),.din(w_dff_A_Xln8IGVO3_0),.clk(gclk));
	jdff dff_A_WCnGhDnX8_0(.dout(w_dff_A_Xln8IGVO3_0),.din(w_dff_A_WCnGhDnX8_0),.clk(gclk));
	jdff dff_A_4jhB6L743_0(.dout(w_dff_A_WCnGhDnX8_0),.din(w_dff_A_4jhB6L743_0),.clk(gclk));
	jdff dff_A_idRuKuo31_0(.dout(w_dff_A_4jhB6L743_0),.din(w_dff_A_idRuKuo31_0),.clk(gclk));
	jdff dff_A_HZuQsZKv6_0(.dout(w_dff_A_idRuKuo31_0),.din(w_dff_A_HZuQsZKv6_0),.clk(gclk));
	jdff dff_A_2BnHsd3a5_0(.dout(w_n749_2[0]),.din(w_dff_A_2BnHsd3a5_0),.clk(gclk));
	jdff dff_A_ILvPx3Bw2_0(.dout(w_dff_A_2BnHsd3a5_0),.din(w_dff_A_ILvPx3Bw2_0),.clk(gclk));
	jdff dff_A_r9II7cxP0_1(.dout(w_n749_2[1]),.din(w_dff_A_r9II7cxP0_1),.clk(gclk));
	jdff dff_A_ylr9DSxj3_1(.dout(w_dff_A_r9II7cxP0_1),.din(w_dff_A_ylr9DSxj3_1),.clk(gclk));
	jdff dff_B_R6hTYZ170_1(.din(G115),.dout(w_dff_B_R6hTYZ170_1),.clk(gclk));
	jdff dff_B_x0JyqcE81_1(.din(w_dff_B_R6hTYZ170_1),.dout(w_dff_B_x0JyqcE81_1),.clk(gclk));
	jdff dff_B_8AWjwpun6_0(.din(n1505),.dout(w_dff_B_8AWjwpun6_0),.clk(gclk));
	jdff dff_B_SyI5cbYT6_0(.din(w_dff_B_8AWjwpun6_0),.dout(w_dff_B_SyI5cbYT6_0),.clk(gclk));
	jdff dff_B_HtJ1tkWA4_0(.din(w_dff_B_SyI5cbYT6_0),.dout(w_dff_B_HtJ1tkWA4_0),.clk(gclk));
	jdff dff_B_mkrlpxlu3_0(.din(w_dff_B_HtJ1tkWA4_0),.dout(w_dff_B_mkrlpxlu3_0),.clk(gclk));
	jdff dff_B_Rsl7u3pY8_0(.din(w_dff_B_mkrlpxlu3_0),.dout(w_dff_B_Rsl7u3pY8_0),.clk(gclk));
	jdff dff_B_OsXF8n4H2_0(.din(w_dff_B_Rsl7u3pY8_0),.dout(w_dff_B_OsXF8n4H2_0),.clk(gclk));
	jdff dff_B_WX07blrw5_0(.din(w_dff_B_OsXF8n4H2_0),.dout(w_dff_B_WX07blrw5_0),.clk(gclk));
	jdff dff_B_AGJ2n9JF5_0(.din(w_dff_B_WX07blrw5_0),.dout(w_dff_B_AGJ2n9JF5_0),.clk(gclk));
	jdff dff_B_oIZfdQ3t3_0(.din(w_dff_B_AGJ2n9JF5_0),.dout(w_dff_B_oIZfdQ3t3_0),.clk(gclk));
	jdff dff_B_0owryR163_0(.din(w_dff_B_oIZfdQ3t3_0),.dout(w_dff_B_0owryR163_0),.clk(gclk));
	jdff dff_B_IEV8kL8x3_0(.din(w_dff_B_0owryR163_0),.dout(w_dff_B_IEV8kL8x3_0),.clk(gclk));
	jdff dff_B_IBCxfeT16_0(.din(w_dff_B_IEV8kL8x3_0),.dout(w_dff_B_IBCxfeT16_0),.clk(gclk));
	jdff dff_B_HWXJRv2U3_0(.din(w_dff_B_IBCxfeT16_0),.dout(w_dff_B_HWXJRv2U3_0),.clk(gclk));
	jdff dff_B_91Hm7drc8_0(.din(w_dff_B_HWXJRv2U3_0),.dout(w_dff_B_91Hm7drc8_0),.clk(gclk));
	jdff dff_B_dTxkmirP4_0(.din(w_dff_B_91Hm7drc8_0),.dout(w_dff_B_dTxkmirP4_0),.clk(gclk));
	jdff dff_B_9DTG6AAB9_0(.din(w_dff_B_dTxkmirP4_0),.dout(w_dff_B_9DTG6AAB9_0),.clk(gclk));
	jdff dff_B_2nAI3GlU6_0(.din(w_dff_B_9DTG6AAB9_0),.dout(w_dff_B_2nAI3GlU6_0),.clk(gclk));
	jdff dff_B_Vik9IfoL0_1(.din(G120),.dout(w_dff_B_Vik9IfoL0_1),.clk(gclk));
	jdff dff_B_VuECQi0n9_1(.din(w_dff_B_Vik9IfoL0_1),.dout(w_dff_B_VuECQi0n9_1),.clk(gclk));
	jdff dff_B_dichDG2I4_1(.din(w_dff_B_VuECQi0n9_1),.dout(w_dff_B_dichDG2I4_1),.clk(gclk));
	jdff dff_B_1p4irCzB1_0(.din(n1666),.dout(w_dff_B_1p4irCzB1_0),.clk(gclk));
	jdff dff_B_81zL4H8Z9_0(.din(w_dff_B_1p4irCzB1_0),.dout(w_dff_B_81zL4H8Z9_0),.clk(gclk));
	jdff dff_B_kPiXskZA6_0(.din(w_dff_B_81zL4H8Z9_0),.dout(w_dff_B_kPiXskZA6_0),.clk(gclk));
	jdff dff_B_QmSMmMpn5_0(.din(w_dff_B_kPiXskZA6_0),.dout(w_dff_B_QmSMmMpn5_0),.clk(gclk));
	jdff dff_B_iw81HcQw0_0(.din(w_dff_B_QmSMmMpn5_0),.dout(w_dff_B_iw81HcQw0_0),.clk(gclk));
	jdff dff_B_04dMJrY67_0(.din(w_dff_B_iw81HcQw0_0),.dout(w_dff_B_04dMJrY67_0),.clk(gclk));
	jdff dff_B_ft4cY8BK5_0(.din(w_dff_B_04dMJrY67_0),.dout(w_dff_B_ft4cY8BK5_0),.clk(gclk));
	jdff dff_B_Ul80cRAF5_0(.din(w_dff_B_ft4cY8BK5_0),.dout(w_dff_B_Ul80cRAF5_0),.clk(gclk));
	jdff dff_B_HVbh6isF9_0(.din(w_dff_B_Ul80cRAF5_0),.dout(w_dff_B_HVbh6isF9_0),.clk(gclk));
	jdff dff_B_VrASsSzX3_0(.din(w_dff_B_HVbh6isF9_0),.dout(w_dff_B_VrASsSzX3_0),.clk(gclk));
	jdff dff_B_tFw8L8ZE6_0(.din(w_dff_B_VrASsSzX3_0),.dout(w_dff_B_tFw8L8ZE6_0),.clk(gclk));
	jdff dff_B_OwOVWKcW5_0(.din(w_dff_B_tFw8L8ZE6_0),.dout(w_dff_B_OwOVWKcW5_0),.clk(gclk));
	jdff dff_B_LNrbF8xU3_0(.din(w_dff_B_OwOVWKcW5_0),.dout(w_dff_B_LNrbF8xU3_0),.clk(gclk));
	jdff dff_B_n8iNjRAv9_0(.din(w_dff_B_LNrbF8xU3_0),.dout(w_dff_B_n8iNjRAv9_0),.clk(gclk));
	jdff dff_B_af7GzYc13_0(.din(w_dff_B_n8iNjRAv9_0),.dout(w_dff_B_af7GzYc13_0),.clk(gclk));
	jdff dff_B_eAEItApn7_0(.din(w_dff_B_af7GzYc13_0),.dout(w_dff_B_eAEItApn7_0),.clk(gclk));
	jdff dff_B_VLqBh0GW4_0(.din(w_dff_B_eAEItApn7_0),.dout(w_dff_B_VLqBh0GW4_0),.clk(gclk));
	jdff dff_B_YmPSEMOH6_1(.din(G118),.dout(w_dff_B_YmPSEMOH6_1),.clk(gclk));
	jdff dff_B_I52hihRt6_1(.din(w_dff_B_YmPSEMOH6_1),.dout(w_dff_B_I52hihRt6_1),.clk(gclk));
	jdff dff_B_2TsCaoR02_1(.din(w_dff_B_I52hihRt6_1),.dout(w_dff_B_2TsCaoR02_1),.clk(gclk));
	jdff dff_A_8ObYxFQD0_0(.dout(w_G4092_9[0]),.din(w_dff_A_8ObYxFQD0_0),.clk(gclk));
	jdff dff_A_hoerIxgT4_0(.dout(w_dff_A_8ObYxFQD0_0),.din(w_dff_A_hoerIxgT4_0),.clk(gclk));
	jdff dff_A_szTvRgYt2_0(.dout(w_dff_A_hoerIxgT4_0),.din(w_dff_A_szTvRgYt2_0),.clk(gclk));
	jdff dff_A_VendsrEd8_0(.dout(w_dff_A_szTvRgYt2_0),.din(w_dff_A_VendsrEd8_0),.clk(gclk));
	jdff dff_A_ifR6nME50_0(.dout(w_dff_A_VendsrEd8_0),.din(w_dff_A_ifR6nME50_0),.clk(gclk));
	jdff dff_A_3CygBpVO8_1(.dout(w_G4092_9[1]),.din(w_dff_A_3CygBpVO8_1),.clk(gclk));
	jdff dff_A_4NLguyDh3_1(.dout(w_dff_A_3CygBpVO8_1),.din(w_dff_A_4NLguyDh3_1),.clk(gclk));
	jdff dff_A_6lPGGltN3_1(.dout(w_dff_A_4NLguyDh3_1),.din(w_dff_A_6lPGGltN3_1),.clk(gclk));
	jdff dff_A_RhMIT62F1_1(.dout(w_dff_A_6lPGGltN3_1),.din(w_dff_A_RhMIT62F1_1),.clk(gclk));
	jdff dff_A_1J9UpE711_0(.dout(w_G4092_2[0]),.din(w_dff_A_1J9UpE711_0),.clk(gclk));
	jdff dff_A_QQJsqeN94_0(.dout(w_dff_A_1J9UpE711_0),.din(w_dff_A_QQJsqeN94_0),.clk(gclk));
	jdff dff_A_MEQeOdlP0_0(.dout(w_dff_A_QQJsqeN94_0),.din(w_dff_A_MEQeOdlP0_0),.clk(gclk));
	jdff dff_A_S4xEADRG4_0(.dout(w_dff_A_MEQeOdlP0_0),.din(w_dff_A_S4xEADRG4_0),.clk(gclk));
	jdff dff_A_wMAhAGCw2_0(.dout(w_dff_A_S4xEADRG4_0),.din(w_dff_A_wMAhAGCw2_0),.clk(gclk));
	jdff dff_A_xHRW5i751_1(.dout(w_G4092_2[1]),.din(w_dff_A_xHRW5i751_1),.clk(gclk));
	jdff dff_A_67FO2KtR2_1(.dout(w_dff_A_xHRW5i751_1),.din(w_dff_A_67FO2KtR2_1),.clk(gclk));
	jdff dff_A_ueoFOx6y3_1(.dout(w_dff_A_67FO2KtR2_1),.din(w_dff_A_ueoFOx6y3_1),.clk(gclk));
	jdff dff_A_ggGHQquF5_1(.dout(w_dff_A_ueoFOx6y3_1),.din(w_dff_A_ggGHQquF5_1),.clk(gclk));
	jdff dff_A_cqBgmFZs1_0(.dout(w_n749_13[0]),.din(w_dff_A_cqBgmFZs1_0),.clk(gclk));
	jdff dff_A_IMPRyMYe5_0(.dout(w_dff_A_cqBgmFZs1_0),.din(w_dff_A_IMPRyMYe5_0),.clk(gclk));
	jdff dff_A_UPfevPH08_0(.dout(w_dff_A_IMPRyMYe5_0),.din(w_dff_A_UPfevPH08_0),.clk(gclk));
	jdff dff_B_5e5zuS1a7_1(.din(n1671),.dout(w_dff_B_5e5zuS1a7_1),.clk(gclk));
	jdff dff_B_cScKjOlA1_1(.din(w_dff_B_5e5zuS1a7_1),.dout(w_dff_B_cScKjOlA1_1),.clk(gclk));
	jdff dff_B_Soo3aZbp8_1(.din(w_dff_B_cScKjOlA1_1),.dout(w_dff_B_Soo3aZbp8_1),.clk(gclk));
	jdff dff_B_4kkelaZl7_1(.din(w_dff_B_Soo3aZbp8_1),.dout(w_dff_B_4kkelaZl7_1),.clk(gclk));
	jdff dff_B_0CCn8k5K2_1(.din(w_dff_B_4kkelaZl7_1),.dout(w_dff_B_0CCn8k5K2_1),.clk(gclk));
	jdff dff_B_6iKiU5vD1_1(.din(w_dff_B_0CCn8k5K2_1),.dout(w_dff_B_6iKiU5vD1_1),.clk(gclk));
	jdff dff_B_WyjygRrj8_1(.din(w_dff_B_6iKiU5vD1_1),.dout(w_dff_B_WyjygRrj8_1),.clk(gclk));
	jdff dff_B_tmKQDly99_1(.din(w_dff_B_WyjygRrj8_1),.dout(w_dff_B_tmKQDly99_1),.clk(gclk));
	jdff dff_B_B3u4WQN31_1(.din(w_dff_B_tmKQDly99_1),.dout(w_dff_B_B3u4WQN31_1),.clk(gclk));
	jdff dff_B_0LXL32Ip2_1(.din(w_dff_B_B3u4WQN31_1),.dout(w_dff_B_0LXL32Ip2_1),.clk(gclk));
	jdff dff_B_vi5kGt7H4_1(.din(w_dff_B_0LXL32Ip2_1),.dout(w_dff_B_vi5kGt7H4_1),.clk(gclk));
	jdff dff_B_srHVl0kn2_1(.din(w_dff_B_vi5kGt7H4_1),.dout(w_dff_B_srHVl0kn2_1),.clk(gclk));
	jdff dff_B_fXDtazfX6_1(.din(w_dff_B_srHVl0kn2_1),.dout(w_dff_B_fXDtazfX6_1),.clk(gclk));
	jdff dff_B_cZm5gRNQ2_1(.din(w_dff_B_fXDtazfX6_1),.dout(w_dff_B_cZm5gRNQ2_1),.clk(gclk));
	jdff dff_B_CLiXq3ns6_1(.din(w_dff_B_cZm5gRNQ2_1),.dout(w_dff_B_CLiXq3ns6_1),.clk(gclk));
	jdff dff_B_YfWEKviO1_1(.din(w_dff_B_CLiXq3ns6_1),.dout(w_dff_B_YfWEKviO1_1),.clk(gclk));
	jdff dff_B_96Eip8xL8_1(.din(w_dff_B_YfWEKviO1_1),.dout(w_dff_B_96Eip8xL8_1),.clk(gclk));
	jdff dff_B_CxmjMu431_1(.din(w_dff_B_96Eip8xL8_1),.dout(w_dff_B_CxmjMu431_1),.clk(gclk));
	jdff dff_B_P19xN8GO2_1(.din(w_dff_B_CxmjMu431_1),.dout(w_dff_B_P19xN8GO2_1),.clk(gclk));
	jdff dff_B_RXiEFzrS9_1(.din(w_dff_B_P19xN8GO2_1),.dout(w_dff_B_RXiEFzrS9_1),.clk(gclk));
	jdff dff_B_d7NXM7kH9_1(.din(w_dff_B_RXiEFzrS9_1),.dout(w_dff_B_d7NXM7kH9_1),.clk(gclk));
	jdff dff_B_l62URcUl6_1(.din(w_dff_B_d7NXM7kH9_1),.dout(w_dff_B_l62URcUl6_1),.clk(gclk));
	jdff dff_B_UuyVYPP90_1(.din(n1676),.dout(w_dff_B_UuyVYPP90_1),.clk(gclk));
	jdff dff_A_mKMkx3402_1(.dout(w_n800_1[1]),.din(w_dff_A_mKMkx3402_1),.clk(gclk));
	jdff dff_A_shThLQD70_1(.dout(w_dff_A_mKMkx3402_1),.din(w_dff_A_shThLQD70_1),.clk(gclk));
	jdff dff_A_w0BWLKlM7_1(.dout(w_dff_A_shThLQD70_1),.din(w_dff_A_w0BWLKlM7_1),.clk(gclk));
	jdff dff_A_JK4DdP7w1_1(.dout(w_dff_A_w0BWLKlM7_1),.din(w_dff_A_JK4DdP7w1_1),.clk(gclk));
	jdff dff_A_3sjU6kPM0_1(.dout(w_dff_A_JK4DdP7w1_1),.din(w_dff_A_3sjU6kPM0_1),.clk(gclk));
	jdff dff_A_W06crO5J0_1(.dout(w_dff_A_3sjU6kPM0_1),.din(w_dff_A_W06crO5J0_1),.clk(gclk));
	jdff dff_A_aLNzTqI70_1(.dout(w_dff_A_W06crO5J0_1),.din(w_dff_A_aLNzTqI70_1),.clk(gclk));
	jdff dff_A_T4z7Q8dh8_1(.dout(w_dff_A_aLNzTqI70_1),.din(w_dff_A_T4z7Q8dh8_1),.clk(gclk));
	jdff dff_A_WhiZjXB04_1(.dout(w_dff_A_T4z7Q8dh8_1),.din(w_dff_A_WhiZjXB04_1),.clk(gclk));
	jdff dff_A_S3qR5mKt8_1(.dout(w_dff_A_WhiZjXB04_1),.din(w_dff_A_S3qR5mKt8_1),.clk(gclk));
	jdff dff_A_epKmczTI7_1(.dout(w_dff_A_S3qR5mKt8_1),.din(w_dff_A_epKmczTI7_1),.clk(gclk));
	jdff dff_A_BiVyAeaj8_1(.dout(w_dff_A_epKmczTI7_1),.din(w_dff_A_BiVyAeaj8_1),.clk(gclk));
	jdff dff_A_7AQuVPSb0_1(.dout(w_dff_A_BiVyAeaj8_1),.din(w_dff_A_7AQuVPSb0_1),.clk(gclk));
	jdff dff_A_uDMLZepB0_1(.dout(w_dff_A_7AQuVPSb0_1),.din(w_dff_A_uDMLZepB0_1),.clk(gclk));
	jdff dff_A_2CAjTrrz1_2(.dout(w_n800_1[2]),.din(w_dff_A_2CAjTrrz1_2),.clk(gclk));
	jdff dff_A_0jKcvtdD7_2(.dout(w_dff_A_2CAjTrrz1_2),.din(w_dff_A_0jKcvtdD7_2),.clk(gclk));
	jdff dff_A_6DLwqrha8_2(.dout(w_dff_A_0jKcvtdD7_2),.din(w_dff_A_6DLwqrha8_2),.clk(gclk));
	jdff dff_A_cOUpg74E0_2(.dout(w_dff_A_6DLwqrha8_2),.din(w_dff_A_cOUpg74E0_2),.clk(gclk));
	jdff dff_A_hOCVYeko9_2(.dout(w_dff_A_cOUpg74E0_2),.din(w_dff_A_hOCVYeko9_2),.clk(gclk));
	jdff dff_A_FH4lGZ0e5_2(.dout(w_dff_A_hOCVYeko9_2),.din(w_dff_A_FH4lGZ0e5_2),.clk(gclk));
	jdff dff_A_q5y470NY4_2(.dout(w_dff_A_FH4lGZ0e5_2),.din(w_dff_A_q5y470NY4_2),.clk(gclk));
	jdff dff_A_LSux8jAS9_2(.dout(w_dff_A_q5y470NY4_2),.din(w_dff_A_LSux8jAS9_2),.clk(gclk));
	jdff dff_A_jk8k9AAV0_2(.dout(w_dff_A_LSux8jAS9_2),.din(w_dff_A_jk8k9AAV0_2),.clk(gclk));
	jdff dff_A_BpvSD57Q4_2(.dout(w_dff_A_jk8k9AAV0_2),.din(w_dff_A_BpvSD57Q4_2),.clk(gclk));
	jdff dff_A_QaUtT28p8_1(.dout(w_n800_0[1]),.din(w_dff_A_QaUtT28p8_1),.clk(gclk));
	jdff dff_A_Cy1pQyLf6_1(.dout(w_dff_A_QaUtT28p8_1),.din(w_dff_A_Cy1pQyLf6_1),.clk(gclk));
	jdff dff_A_TQXjjSzL8_1(.dout(w_dff_A_Cy1pQyLf6_1),.din(w_dff_A_TQXjjSzL8_1),.clk(gclk));
	jdff dff_A_WvDWmAAi1_1(.dout(w_dff_A_TQXjjSzL8_1),.din(w_dff_A_WvDWmAAi1_1),.clk(gclk));
	jdff dff_A_rKWZdJN14_1(.dout(w_dff_A_WvDWmAAi1_1),.din(w_dff_A_rKWZdJN14_1),.clk(gclk));
	jdff dff_A_Nj8pWmv18_1(.dout(w_dff_A_rKWZdJN14_1),.din(w_dff_A_Nj8pWmv18_1),.clk(gclk));
	jdff dff_A_el3opAui4_1(.dout(w_dff_A_Nj8pWmv18_1),.din(w_dff_A_el3opAui4_1),.clk(gclk));
	jdff dff_A_PpPYDotE0_1(.dout(w_dff_A_el3opAui4_1),.din(w_dff_A_PpPYDotE0_1),.clk(gclk));
	jdff dff_A_KzQ1iZc55_1(.dout(w_dff_A_PpPYDotE0_1),.din(w_dff_A_KzQ1iZc55_1),.clk(gclk));
	jdff dff_A_HbuwozZH6_1(.dout(w_dff_A_KzQ1iZc55_1),.din(w_dff_A_HbuwozZH6_1),.clk(gclk));
	jdff dff_A_ZWMvM8Jk9_1(.dout(w_dff_A_HbuwozZH6_1),.din(w_dff_A_ZWMvM8Jk9_1),.clk(gclk));
	jdff dff_A_72A47Qsx6_2(.dout(w_n800_0[2]),.din(w_dff_A_72A47Qsx6_2),.clk(gclk));
	jdff dff_A_cgRPNDmG7_2(.dout(w_dff_A_72A47Qsx6_2),.din(w_dff_A_cgRPNDmG7_2),.clk(gclk));
	jdff dff_A_nqtTNS5b0_2(.dout(w_dff_A_cgRPNDmG7_2),.din(w_dff_A_nqtTNS5b0_2),.clk(gclk));
	jdff dff_A_S6rN69Ok5_2(.dout(w_dff_A_nqtTNS5b0_2),.din(w_dff_A_S6rN69Ok5_2),.clk(gclk));
	jdff dff_B_RepmlAMK5_3(.din(n800),.dout(w_dff_B_RepmlAMK5_3),.clk(gclk));
	jdff dff_B_LWef8ZPO9_3(.din(w_dff_B_RepmlAMK5_3),.dout(w_dff_B_LWef8ZPO9_3),.clk(gclk));
	jdff dff_B_rHb0Nf8Z9_3(.din(w_dff_B_LWef8ZPO9_3),.dout(w_dff_B_rHb0Nf8Z9_3),.clk(gclk));
	jdff dff_B_4rLMCRM48_3(.din(w_dff_B_rHb0Nf8Z9_3),.dout(w_dff_B_4rLMCRM48_3),.clk(gclk));
	jdff dff_B_VnJsDzlZ0_3(.din(w_dff_B_4rLMCRM48_3),.dout(w_dff_B_VnJsDzlZ0_3),.clk(gclk));
	jdff dff_B_aeUcAszg5_3(.din(w_dff_B_VnJsDzlZ0_3),.dout(w_dff_B_aeUcAszg5_3),.clk(gclk));
	jdff dff_B_hjkqYJ0R5_3(.din(w_dff_B_aeUcAszg5_3),.dout(w_dff_B_hjkqYJ0R5_3),.clk(gclk));
	jdff dff_B_3fKYXCof6_3(.din(w_dff_B_hjkqYJ0R5_3),.dout(w_dff_B_3fKYXCof6_3),.clk(gclk));
	jdff dff_B_MwUyoqxu1_3(.din(w_dff_B_3fKYXCof6_3),.dout(w_dff_B_MwUyoqxu1_3),.clk(gclk));
	jdff dff_A_s4mXJW8X6_0(.dout(w_G4087_4[0]),.din(w_dff_A_s4mXJW8X6_0),.clk(gclk));
	jdff dff_A_sg5nOhNJ8_1(.dout(w_G4087_4[1]),.din(w_dff_A_sg5nOhNJ8_1),.clk(gclk));
	jdff dff_B_0OfVjyn06_1(.din(n1668),.dout(w_dff_B_0OfVjyn06_1),.clk(gclk));
	jdff dff_B_CZWc9HjP5_1(.din(w_dff_B_0OfVjyn06_1),.dout(w_dff_B_CZWc9HjP5_1),.clk(gclk));
	jdff dff_A_C4fwjque9_0(.dout(w_n797_3[0]),.din(w_dff_A_C4fwjque9_0),.clk(gclk));
	jdff dff_A_VtD9dtYE9_0(.dout(w_dff_A_C4fwjque9_0),.din(w_dff_A_VtD9dtYE9_0),.clk(gclk));
	jdff dff_A_Eo7AXJou5_0(.dout(w_dff_A_VtD9dtYE9_0),.din(w_dff_A_Eo7AXJou5_0),.clk(gclk));
	jdff dff_A_20lzqXXE1_0(.dout(w_dff_A_Eo7AXJou5_0),.din(w_dff_A_20lzqXXE1_0),.clk(gclk));
	jdff dff_A_Rq61JYAI3_0(.dout(w_dff_A_20lzqXXE1_0),.din(w_dff_A_Rq61JYAI3_0),.clk(gclk));
	jdff dff_A_Dpy9uMNc4_0(.dout(w_dff_A_Rq61JYAI3_0),.din(w_dff_A_Dpy9uMNc4_0),.clk(gclk));
	jdff dff_A_V3Ovmbnu8_0(.dout(w_dff_A_Dpy9uMNc4_0),.din(w_dff_A_V3Ovmbnu8_0),.clk(gclk));
	jdff dff_A_t9JhJckN9_0(.dout(w_dff_A_V3Ovmbnu8_0),.din(w_dff_A_t9JhJckN9_0),.clk(gclk));
	jdff dff_A_9E4B0bnc0_0(.dout(w_dff_A_t9JhJckN9_0),.din(w_dff_A_9E4B0bnc0_0),.clk(gclk));
	jdff dff_A_rQSOU49D5_0(.dout(w_dff_A_9E4B0bnc0_0),.din(w_dff_A_rQSOU49D5_0),.clk(gclk));
	jdff dff_A_iCDC3FKU1_0(.dout(w_dff_A_rQSOU49D5_0),.din(w_dff_A_iCDC3FKU1_0),.clk(gclk));
	jdff dff_A_hLzxzN376_0(.dout(w_dff_A_iCDC3FKU1_0),.din(w_dff_A_hLzxzN376_0),.clk(gclk));
	jdff dff_A_yDxUt3ZB4_0(.dout(w_dff_A_hLzxzN376_0),.din(w_dff_A_yDxUt3ZB4_0),.clk(gclk));
	jdff dff_A_Ts7n3fiN4_0(.dout(w_dff_A_yDxUt3ZB4_0),.din(w_dff_A_Ts7n3fiN4_0),.clk(gclk));
	jdff dff_A_HRzarivN0_0(.dout(w_dff_A_Ts7n3fiN4_0),.din(w_dff_A_HRzarivN0_0),.clk(gclk));
	jdff dff_A_I3ctsL385_0(.dout(w_dff_A_HRzarivN0_0),.din(w_dff_A_I3ctsL385_0),.clk(gclk));
	jdff dff_A_l32uxYpM6_0(.dout(w_dff_A_I3ctsL385_0),.din(w_dff_A_l32uxYpM6_0),.clk(gclk));
	jdff dff_A_tbePrfwj9_0(.dout(w_dff_A_l32uxYpM6_0),.din(w_dff_A_tbePrfwj9_0),.clk(gclk));
	jdff dff_A_thC3xxEd2_0(.dout(w_dff_A_tbePrfwj9_0),.din(w_dff_A_thC3xxEd2_0),.clk(gclk));
	jdff dff_A_sX5Gxn2m6_0(.dout(w_dff_A_thC3xxEd2_0),.din(w_dff_A_sX5Gxn2m6_0),.clk(gclk));
	jdff dff_A_93XKIR4Z5_0(.dout(w_dff_A_sX5Gxn2m6_0),.din(w_dff_A_93XKIR4Z5_0),.clk(gclk));
	jdff dff_A_qnlRfEJH3_0(.dout(w_dff_A_93XKIR4Z5_0),.din(w_dff_A_qnlRfEJH3_0),.clk(gclk));
	jdff dff_A_mExzMo0u8_1(.dout(w_G4088_9[1]),.din(w_dff_A_mExzMo0u8_1),.clk(gclk));
	jdff dff_A_R1hUE9gF9_1(.dout(w_dff_A_mExzMo0u8_1),.din(w_dff_A_R1hUE9gF9_1),.clk(gclk));
	jdff dff_A_ahiXVkYi4_1(.dout(w_dff_A_R1hUE9gF9_1),.din(w_dff_A_ahiXVkYi4_1),.clk(gclk));
	jdff dff_A_zH1Fmsaq0_1(.dout(w_dff_A_ahiXVkYi4_1),.din(w_dff_A_zH1Fmsaq0_1),.clk(gclk));
	jdff dff_A_BP8l9MQe5_1(.dout(w_dff_A_zH1Fmsaq0_1),.din(w_dff_A_BP8l9MQe5_1),.clk(gclk));
	jdff dff_A_geeYu1rM2_1(.dout(w_dff_A_BP8l9MQe5_1),.din(w_dff_A_geeYu1rM2_1),.clk(gclk));
	jdff dff_A_1Kyrp0C55_1(.dout(w_dff_A_geeYu1rM2_1),.din(w_dff_A_1Kyrp0C55_1),.clk(gclk));
	jdff dff_A_UUM8XIWb2_1(.dout(w_dff_A_1Kyrp0C55_1),.din(w_dff_A_UUM8XIWb2_1),.clk(gclk));
	jdff dff_A_rup8d4tL5_1(.dout(w_dff_A_UUM8XIWb2_1),.din(w_dff_A_rup8d4tL5_1),.clk(gclk));
	jdff dff_A_cOZVQ2Qy5_1(.dout(w_G4087_1[1]),.din(w_dff_A_cOZVQ2Qy5_1),.clk(gclk));
	jdff dff_A_jiFySq680_1(.dout(w_dff_A_cOZVQ2Qy5_1),.din(w_dff_A_jiFySq680_1),.clk(gclk));
	jdff dff_A_5ViwmFPS6_2(.dout(w_G4087_1[2]),.din(w_dff_A_5ViwmFPS6_2),.clk(gclk));
	jdff dff_A_z4gXNJDl6_1(.dout(w_G4087_0[1]),.din(w_dff_A_z4gXNJDl6_1),.clk(gclk));
	jdff dff_A_RCIjzLbv0_2(.dout(w_G4087_0[2]),.din(w_dff_A_RCIjzLbv0_2),.clk(gclk));
	jdff dff_A_pVl6RSdy0_0(.dout(w_G4088_3[0]),.din(w_dff_A_pVl6RSdy0_0),.clk(gclk));
	jdff dff_A_lG0fvDEl3_0(.dout(w_dff_A_pVl6RSdy0_0),.din(w_dff_A_lG0fvDEl3_0),.clk(gclk));
	jdff dff_A_pPnwH4os3_0(.dout(w_dff_A_lG0fvDEl3_0),.din(w_dff_A_pPnwH4os3_0),.clk(gclk));
	jdff dff_A_UeNZaFw28_0(.dout(w_dff_A_pPnwH4os3_0),.din(w_dff_A_UeNZaFw28_0),.clk(gclk));
	jdff dff_A_yXrFLySN0_0(.dout(w_dff_A_UeNZaFw28_0),.din(w_dff_A_yXrFLySN0_0),.clk(gclk));
	jdff dff_A_m7aGkCFq7_0(.dout(w_dff_A_yXrFLySN0_0),.din(w_dff_A_m7aGkCFq7_0),.clk(gclk));
	jdff dff_A_ektHuPxZ0_0(.dout(w_dff_A_m7aGkCFq7_0),.din(w_dff_A_ektHuPxZ0_0),.clk(gclk));
	jdff dff_A_ePg6tEvb3_0(.dout(w_dff_A_ektHuPxZ0_0),.din(w_dff_A_ePg6tEvb3_0),.clk(gclk));
	jdff dff_A_bYiS5xFi0_0(.dout(w_dff_A_ePg6tEvb3_0),.din(w_dff_A_bYiS5xFi0_0),.clk(gclk));
	jdff dff_A_OKbZz6mn5_0(.dout(w_dff_A_bYiS5xFi0_0),.din(w_dff_A_OKbZz6mn5_0),.clk(gclk));
	jdff dff_A_yMRX3B4B8_0(.dout(w_dff_A_OKbZz6mn5_0),.din(w_dff_A_yMRX3B4B8_0),.clk(gclk));
	jdff dff_A_xs7os9hb7_0(.dout(w_dff_A_yMRX3B4B8_0),.din(w_dff_A_xs7os9hb7_0),.clk(gclk));
	jdff dff_A_dxsp55vT7_0(.dout(w_dff_A_xs7os9hb7_0),.din(w_dff_A_dxsp55vT7_0),.clk(gclk));
	jdff dff_A_zVzCJJkn9_0(.dout(w_dff_A_dxsp55vT7_0),.din(w_dff_A_zVzCJJkn9_0),.clk(gclk));
	jdff dff_A_rPnQuvwW4_0(.dout(w_dff_A_zVzCJJkn9_0),.din(w_dff_A_rPnQuvwW4_0),.clk(gclk));
	jdff dff_A_AoVGNFxa4_0(.dout(w_dff_A_rPnQuvwW4_0),.din(w_dff_A_AoVGNFxa4_0),.clk(gclk));
	jdff dff_A_l5P2P98g9_0(.dout(w_dff_A_AoVGNFxa4_0),.din(w_dff_A_l5P2P98g9_0),.clk(gclk));
	jdff dff_A_AzbpNtx49_0(.dout(w_dff_A_l5P2P98g9_0),.din(w_dff_A_AzbpNtx49_0),.clk(gclk));
	jdff dff_A_RYEMwVuI5_0(.dout(w_dff_A_AzbpNtx49_0),.din(w_dff_A_RYEMwVuI5_0),.clk(gclk));
	jdff dff_A_cQSBFBQn1_0(.dout(w_dff_A_RYEMwVuI5_0),.din(w_dff_A_cQSBFBQn1_0),.clk(gclk));
	jdff dff_A_kKjm6x1T3_0(.dout(w_dff_A_cQSBFBQn1_0),.din(w_dff_A_kKjm6x1T3_0),.clk(gclk));
	jdff dff_A_rvtdpdSA9_0(.dout(w_dff_A_kKjm6x1T3_0),.din(w_dff_A_rvtdpdSA9_0),.clk(gclk));
	jdff dff_A_a1YkzlzF7_0(.dout(w_dff_A_rvtdpdSA9_0),.din(w_dff_A_a1YkzlzF7_0),.clk(gclk));
	jdff dff_B_HgJ8UPjT6_1(.din(n1688),.dout(w_dff_B_HgJ8UPjT6_1),.clk(gclk));
	jdff dff_B_YWLnt9UX1_1(.din(w_dff_B_HgJ8UPjT6_1),.dout(w_dff_B_YWLnt9UX1_1),.clk(gclk));
	jdff dff_B_MPOY0pX70_1(.din(w_dff_B_YWLnt9UX1_1),.dout(w_dff_B_MPOY0pX70_1),.clk(gclk));
	jdff dff_B_a62O9a6C9_1(.din(w_dff_B_MPOY0pX70_1),.dout(w_dff_B_a62O9a6C9_1),.clk(gclk));
	jdff dff_B_ZWfbfxKp9_1(.din(w_dff_B_a62O9a6C9_1),.dout(w_dff_B_ZWfbfxKp9_1),.clk(gclk));
	jdff dff_B_x72qEU6c5_1(.din(w_dff_B_ZWfbfxKp9_1),.dout(w_dff_B_x72qEU6c5_1),.clk(gclk));
	jdff dff_B_4TdQoK0d6_1(.din(w_dff_B_x72qEU6c5_1),.dout(w_dff_B_4TdQoK0d6_1),.clk(gclk));
	jdff dff_B_VckQEQ0L1_1(.din(w_dff_B_4TdQoK0d6_1),.dout(w_dff_B_VckQEQ0L1_1),.clk(gclk));
	jdff dff_B_Wm1Zug195_1(.din(w_dff_B_VckQEQ0L1_1),.dout(w_dff_B_Wm1Zug195_1),.clk(gclk));
	jdff dff_B_XN2ZOdsd8_1(.din(w_dff_B_Wm1Zug195_1),.dout(w_dff_B_XN2ZOdsd8_1),.clk(gclk));
	jdff dff_B_MiBFHln91_1(.din(w_dff_B_XN2ZOdsd8_1),.dout(w_dff_B_MiBFHln91_1),.clk(gclk));
	jdff dff_B_SeNIhFYC4_1(.din(w_dff_B_MiBFHln91_1),.dout(w_dff_B_SeNIhFYC4_1),.clk(gclk));
	jdff dff_B_wbKTMj9v2_1(.din(w_dff_B_SeNIhFYC4_1),.dout(w_dff_B_wbKTMj9v2_1),.clk(gclk));
	jdff dff_B_mtPs3ggg7_1(.din(w_dff_B_wbKTMj9v2_1),.dout(w_dff_B_mtPs3ggg7_1),.clk(gclk));
	jdff dff_B_r5Hnzn2T6_1(.din(w_dff_B_mtPs3ggg7_1),.dout(w_dff_B_r5Hnzn2T6_1),.clk(gclk));
	jdff dff_B_OBjHK4ED8_1(.din(w_dff_B_r5Hnzn2T6_1),.dout(w_dff_B_OBjHK4ED8_1),.clk(gclk));
	jdff dff_B_7e4hA8VI6_1(.din(w_dff_B_OBjHK4ED8_1),.dout(w_dff_B_7e4hA8VI6_1),.clk(gclk));
	jdff dff_B_ABBur8aH1_1(.din(w_dff_B_7e4hA8VI6_1),.dout(w_dff_B_ABBur8aH1_1),.clk(gclk));
	jdff dff_B_1aanQgeF5_1(.din(w_dff_B_ABBur8aH1_1),.dout(w_dff_B_1aanQgeF5_1),.clk(gclk));
	jdff dff_B_1zhas1ym0_1(.din(w_dff_B_1aanQgeF5_1),.dout(w_dff_B_1zhas1ym0_1),.clk(gclk));
	jdff dff_B_3yr8icmq5_1(.din(w_dff_B_1zhas1ym0_1),.dout(w_dff_B_3yr8icmq5_1),.clk(gclk));
	jdff dff_B_nzzW5EV01_1(.din(w_dff_B_3yr8icmq5_1),.dout(w_dff_B_nzzW5EV01_1),.clk(gclk));
	jdff dff_B_kT1rIe232_1(.din(n1689),.dout(w_dff_B_kT1rIe232_1),.clk(gclk));
	jdff dff_A_4jVOEVBg2_1(.dout(w_n854_1[1]),.din(w_dff_A_4jVOEVBg2_1),.clk(gclk));
	jdff dff_A_3Espyj9e2_1(.dout(w_dff_A_4jVOEVBg2_1),.din(w_dff_A_3Espyj9e2_1),.clk(gclk));
	jdff dff_A_PjoTc44T1_1(.dout(w_dff_A_3Espyj9e2_1),.din(w_dff_A_PjoTc44T1_1),.clk(gclk));
	jdff dff_A_Pg61oTH26_1(.dout(w_dff_A_PjoTc44T1_1),.din(w_dff_A_Pg61oTH26_1),.clk(gclk));
	jdff dff_A_Cjwjtw2x4_1(.dout(w_dff_A_Pg61oTH26_1),.din(w_dff_A_Cjwjtw2x4_1),.clk(gclk));
	jdff dff_A_YGWF4hHO2_1(.dout(w_dff_A_Cjwjtw2x4_1),.din(w_dff_A_YGWF4hHO2_1),.clk(gclk));
	jdff dff_A_bs99USbQ0_1(.dout(w_dff_A_YGWF4hHO2_1),.din(w_dff_A_bs99USbQ0_1),.clk(gclk));
	jdff dff_A_staoFMI34_1(.dout(w_dff_A_bs99USbQ0_1),.din(w_dff_A_staoFMI34_1),.clk(gclk));
	jdff dff_A_dQmaPLvb6_1(.dout(w_dff_A_staoFMI34_1),.din(w_dff_A_dQmaPLvb6_1),.clk(gclk));
	jdff dff_A_RCCUsXbQ6_1(.dout(w_dff_A_dQmaPLvb6_1),.din(w_dff_A_RCCUsXbQ6_1),.clk(gclk));
	jdff dff_A_gWCrgGVr6_1(.dout(w_dff_A_RCCUsXbQ6_1),.din(w_dff_A_gWCrgGVr6_1),.clk(gclk));
	jdff dff_A_4eNIcdzN6_1(.dout(w_dff_A_gWCrgGVr6_1),.din(w_dff_A_4eNIcdzN6_1),.clk(gclk));
	jdff dff_A_UdhofHLe6_1(.dout(w_dff_A_4eNIcdzN6_1),.din(w_dff_A_UdhofHLe6_1),.clk(gclk));
	jdff dff_A_tYiNUfGA0_1(.dout(w_dff_A_UdhofHLe6_1),.din(w_dff_A_tYiNUfGA0_1),.clk(gclk));
	jdff dff_A_vsaFAMqD6_2(.dout(w_n854_1[2]),.din(w_dff_A_vsaFAMqD6_2),.clk(gclk));
	jdff dff_A_cPi1KRNX2_2(.dout(w_dff_A_vsaFAMqD6_2),.din(w_dff_A_cPi1KRNX2_2),.clk(gclk));
	jdff dff_A_Q2kYCTVY1_2(.dout(w_dff_A_cPi1KRNX2_2),.din(w_dff_A_Q2kYCTVY1_2),.clk(gclk));
	jdff dff_A_NVDIreXF1_2(.dout(w_dff_A_Q2kYCTVY1_2),.din(w_dff_A_NVDIreXF1_2),.clk(gclk));
	jdff dff_A_e1ygDbgS2_2(.dout(w_dff_A_NVDIreXF1_2),.din(w_dff_A_e1ygDbgS2_2),.clk(gclk));
	jdff dff_A_1wbVN6Ao6_2(.dout(w_dff_A_e1ygDbgS2_2),.din(w_dff_A_1wbVN6Ao6_2),.clk(gclk));
	jdff dff_A_Qr4wcDax7_2(.dout(w_dff_A_1wbVN6Ao6_2),.din(w_dff_A_Qr4wcDax7_2),.clk(gclk));
	jdff dff_A_otfdHdpE7_2(.dout(w_dff_A_Qr4wcDax7_2),.din(w_dff_A_otfdHdpE7_2),.clk(gclk));
	jdff dff_A_WSJtnANh8_2(.dout(w_dff_A_otfdHdpE7_2),.din(w_dff_A_WSJtnANh8_2),.clk(gclk));
	jdff dff_A_jY9b8IVo4_2(.dout(w_dff_A_WSJtnANh8_2),.din(w_dff_A_jY9b8IVo4_2),.clk(gclk));
	jdff dff_A_EpsawGem2_1(.dout(w_n854_0[1]),.din(w_dff_A_EpsawGem2_1),.clk(gclk));
	jdff dff_A_yUKHhQlm8_1(.dout(w_dff_A_EpsawGem2_1),.din(w_dff_A_yUKHhQlm8_1),.clk(gclk));
	jdff dff_A_4qoWoKgS0_1(.dout(w_dff_A_yUKHhQlm8_1),.din(w_dff_A_4qoWoKgS0_1),.clk(gclk));
	jdff dff_A_1BgLTNUL3_1(.dout(w_dff_A_4qoWoKgS0_1),.din(w_dff_A_1BgLTNUL3_1),.clk(gclk));
	jdff dff_A_gQJlXu2F1_1(.dout(w_dff_A_1BgLTNUL3_1),.din(w_dff_A_gQJlXu2F1_1),.clk(gclk));
	jdff dff_A_hHTfZ0Hv9_1(.dout(w_dff_A_gQJlXu2F1_1),.din(w_dff_A_hHTfZ0Hv9_1),.clk(gclk));
	jdff dff_A_Kuwqft7N9_1(.dout(w_dff_A_hHTfZ0Hv9_1),.din(w_dff_A_Kuwqft7N9_1),.clk(gclk));
	jdff dff_A_0KwAEId78_1(.dout(w_dff_A_Kuwqft7N9_1),.din(w_dff_A_0KwAEId78_1),.clk(gclk));
	jdff dff_A_CWkbWoNy0_1(.dout(w_dff_A_0KwAEId78_1),.din(w_dff_A_CWkbWoNy0_1),.clk(gclk));
	jdff dff_A_DQyYBON80_1(.dout(w_dff_A_CWkbWoNy0_1),.din(w_dff_A_DQyYBON80_1),.clk(gclk));
	jdff dff_A_Jnct4fnW9_1(.dout(w_dff_A_DQyYBON80_1),.din(w_dff_A_Jnct4fnW9_1),.clk(gclk));
	jdff dff_A_xMfdpUh61_2(.dout(w_n854_0[2]),.din(w_dff_A_xMfdpUh61_2),.clk(gclk));
	jdff dff_A_eTq7qqbM5_2(.dout(w_dff_A_xMfdpUh61_2),.din(w_dff_A_eTq7qqbM5_2),.clk(gclk));
	jdff dff_A_5whRubta6_2(.dout(w_dff_A_eTq7qqbM5_2),.din(w_dff_A_5whRubta6_2),.clk(gclk));
	jdff dff_A_xl7ytOp19_2(.dout(w_dff_A_5whRubta6_2),.din(w_dff_A_xl7ytOp19_2),.clk(gclk));
	jdff dff_A_yKkjTM6S1_2(.dout(w_dff_A_xl7ytOp19_2),.din(w_dff_A_yKkjTM6S1_2),.clk(gclk));
	jdff dff_B_EDGMNkaZ3_3(.din(n854),.dout(w_dff_B_EDGMNkaZ3_3),.clk(gclk));
	jdff dff_B_XYvyIm6Z7_3(.din(w_dff_B_EDGMNkaZ3_3),.dout(w_dff_B_XYvyIm6Z7_3),.clk(gclk));
	jdff dff_B_5H2dPdpX3_3(.din(w_dff_B_XYvyIm6Z7_3),.dout(w_dff_B_5H2dPdpX3_3),.clk(gclk));
	jdff dff_B_NagbFXfR8_3(.din(w_dff_B_5H2dPdpX3_3),.dout(w_dff_B_NagbFXfR8_3),.clk(gclk));
	jdff dff_B_EiMOcFUM2_3(.din(w_dff_B_NagbFXfR8_3),.dout(w_dff_B_EiMOcFUM2_3),.clk(gclk));
	jdff dff_B_SszUKQ7U8_3(.din(w_dff_B_EiMOcFUM2_3),.dout(w_dff_B_SszUKQ7U8_3),.clk(gclk));
	jdff dff_B_OOGxSDZl3_3(.din(w_dff_B_SszUKQ7U8_3),.dout(w_dff_B_OOGxSDZl3_3),.clk(gclk));
	jdff dff_B_ewRcziBi2_3(.din(w_dff_B_OOGxSDZl3_3),.dout(w_dff_B_ewRcziBi2_3),.clk(gclk));
	jdff dff_B_d5G7vJYJ1_3(.din(w_dff_B_ewRcziBi2_3),.dout(w_dff_B_d5G7vJYJ1_3),.clk(gclk));
	jdff dff_A_ZKP47iAl5_0(.dout(w_G4090_4[0]),.din(w_dff_A_ZKP47iAl5_0),.clk(gclk));
	jdff dff_A_yU2mtP1v8_0(.dout(w_dff_A_ZKP47iAl5_0),.din(w_dff_A_yU2mtP1v8_0),.clk(gclk));
	jdff dff_A_wsrgcQzq2_1(.dout(w_G4090_4[1]),.din(w_dff_A_wsrgcQzq2_1),.clk(gclk));
	jdff dff_B_8HhfATdu6_1(.din(n1685),.dout(w_dff_B_8HhfATdu6_1),.clk(gclk));
	jdff dff_B_X3poD1NW2_1(.din(w_dff_B_8HhfATdu6_1),.dout(w_dff_B_X3poD1NW2_1),.clk(gclk));
	jdff dff_A_nnritehd3_0(.dout(w_n852_3[0]),.din(w_dff_A_nnritehd3_0),.clk(gclk));
	jdff dff_A_bFJAuPFw7_0(.dout(w_dff_A_nnritehd3_0),.din(w_dff_A_bFJAuPFw7_0),.clk(gclk));
	jdff dff_A_cSVcj86P3_0(.dout(w_dff_A_bFJAuPFw7_0),.din(w_dff_A_cSVcj86P3_0),.clk(gclk));
	jdff dff_A_ES1gNpws5_0(.dout(w_dff_A_cSVcj86P3_0),.din(w_dff_A_ES1gNpws5_0),.clk(gclk));
	jdff dff_A_uZ2MuqYv7_0(.dout(w_dff_A_ES1gNpws5_0),.din(w_dff_A_uZ2MuqYv7_0),.clk(gclk));
	jdff dff_A_SsgtXLWW5_0(.dout(w_dff_A_uZ2MuqYv7_0),.din(w_dff_A_SsgtXLWW5_0),.clk(gclk));
	jdff dff_A_nRZzmmkZ5_0(.dout(w_dff_A_SsgtXLWW5_0),.din(w_dff_A_nRZzmmkZ5_0),.clk(gclk));
	jdff dff_A_zPJl7H4M7_0(.dout(w_dff_A_nRZzmmkZ5_0),.din(w_dff_A_zPJl7H4M7_0),.clk(gclk));
	jdff dff_A_mFBio6Xq5_0(.dout(w_dff_A_zPJl7H4M7_0),.din(w_dff_A_mFBio6Xq5_0),.clk(gclk));
	jdff dff_A_CMvuMxIf6_0(.dout(w_dff_A_mFBio6Xq5_0),.din(w_dff_A_CMvuMxIf6_0),.clk(gclk));
	jdff dff_A_r6ROu1PE9_0(.dout(w_dff_A_CMvuMxIf6_0),.din(w_dff_A_r6ROu1PE9_0),.clk(gclk));
	jdff dff_A_cKfaf0gZ1_0(.dout(w_dff_A_r6ROu1PE9_0),.din(w_dff_A_cKfaf0gZ1_0),.clk(gclk));
	jdff dff_A_JwPA8TKO3_0(.dout(w_dff_A_cKfaf0gZ1_0),.din(w_dff_A_JwPA8TKO3_0),.clk(gclk));
	jdff dff_A_xbm5mn4H7_0(.dout(w_dff_A_JwPA8TKO3_0),.din(w_dff_A_xbm5mn4H7_0),.clk(gclk));
	jdff dff_A_QvaSjINX6_0(.dout(w_dff_A_xbm5mn4H7_0),.din(w_dff_A_QvaSjINX6_0),.clk(gclk));
	jdff dff_A_iWzEyBod0_0(.dout(w_dff_A_QvaSjINX6_0),.din(w_dff_A_iWzEyBod0_0),.clk(gclk));
	jdff dff_A_WMgA96Mm9_0(.dout(w_dff_A_iWzEyBod0_0),.din(w_dff_A_WMgA96Mm9_0),.clk(gclk));
	jdff dff_A_OMsHxYZy4_0(.dout(w_dff_A_WMgA96Mm9_0),.din(w_dff_A_OMsHxYZy4_0),.clk(gclk));
	jdff dff_A_nOhZi9TO3_0(.dout(w_dff_A_OMsHxYZy4_0),.din(w_dff_A_nOhZi9TO3_0),.clk(gclk));
	jdff dff_A_Fodnh04C3_0(.dout(w_dff_A_nOhZi9TO3_0),.din(w_dff_A_Fodnh04C3_0),.clk(gclk));
	jdff dff_A_ho5eJw8Q2_0(.dout(w_dff_A_Fodnh04C3_0),.din(w_dff_A_ho5eJw8Q2_0),.clk(gclk));
	jdff dff_A_ViaIf9gQ0_0(.dout(w_dff_A_ho5eJw8Q2_0),.din(w_dff_A_ViaIf9gQ0_0),.clk(gclk));
	jdff dff_A_49fwpllY0_1(.dout(w_G4089_9[1]),.din(w_dff_A_49fwpllY0_1),.clk(gclk));
	jdff dff_A_RyKlHmmw9_1(.dout(w_dff_A_49fwpllY0_1),.din(w_dff_A_RyKlHmmw9_1),.clk(gclk));
	jdff dff_A_fPv4t5mR7_1(.dout(w_dff_A_RyKlHmmw9_1),.din(w_dff_A_fPv4t5mR7_1),.clk(gclk));
	jdff dff_A_2udNlhav7_1(.dout(w_dff_A_fPv4t5mR7_1),.din(w_dff_A_2udNlhav7_1),.clk(gclk));
	jdff dff_A_xRSxyns32_1(.dout(w_dff_A_2udNlhav7_1),.din(w_dff_A_xRSxyns32_1),.clk(gclk));
	jdff dff_A_AXj1pz1W1_1(.dout(w_dff_A_xRSxyns32_1),.din(w_dff_A_AXj1pz1W1_1),.clk(gclk));
	jdff dff_A_5UMxVzrt3_1(.dout(w_dff_A_AXj1pz1W1_1),.din(w_dff_A_5UMxVzrt3_1),.clk(gclk));
	jdff dff_A_U6VoDHgm8_1(.dout(w_dff_A_5UMxVzrt3_1),.din(w_dff_A_U6VoDHgm8_1),.clk(gclk));
	jdff dff_A_U89a4rlK1_1(.dout(w_dff_A_U6VoDHgm8_1),.din(w_dff_A_U89a4rlK1_1),.clk(gclk));
	jdff dff_B_usrkDEF45_2(.din(G64),.dout(w_dff_B_usrkDEF45_2),.clk(gclk));
	jdff dff_A_78NHFyP55_1(.dout(w_G4090_1[1]),.din(w_dff_A_78NHFyP55_1),.clk(gclk));
	jdff dff_A_UJNqLQE41_1(.dout(w_dff_A_78NHFyP55_1),.din(w_dff_A_UJNqLQE41_1),.clk(gclk));
	jdff dff_A_8bKgs9nA1_2(.dout(w_G4090_1[2]),.din(w_dff_A_8bKgs9nA1_2),.clk(gclk));
	jdff dff_A_REUvvtvf3_1(.dout(w_G4090_0[1]),.din(w_dff_A_REUvvtvf3_1),.clk(gclk));
	jdff dff_A_W5GRnw7Q9_2(.dout(w_G4090_0[2]),.din(w_dff_A_W5GRnw7Q9_2),.clk(gclk));
	jdff dff_A_kYAyl4Es8_0(.dout(w_G4089_3[0]),.din(w_dff_A_kYAyl4Es8_0),.clk(gclk));
	jdff dff_A_xbX0qH2H3_0(.dout(w_dff_A_kYAyl4Es8_0),.din(w_dff_A_xbX0qH2H3_0),.clk(gclk));
	jdff dff_A_cFnGhN872_0(.dout(w_dff_A_xbX0qH2H3_0),.din(w_dff_A_cFnGhN872_0),.clk(gclk));
	jdff dff_A_iuIvA3rV3_0(.dout(w_dff_A_cFnGhN872_0),.din(w_dff_A_iuIvA3rV3_0),.clk(gclk));
	jdff dff_A_pqW3gnFS2_0(.dout(w_dff_A_iuIvA3rV3_0),.din(w_dff_A_pqW3gnFS2_0),.clk(gclk));
	jdff dff_A_TkTNPPh29_0(.dout(w_dff_A_pqW3gnFS2_0),.din(w_dff_A_TkTNPPh29_0),.clk(gclk));
	jdff dff_A_XiUTjsH41_0(.dout(w_dff_A_TkTNPPh29_0),.din(w_dff_A_XiUTjsH41_0),.clk(gclk));
	jdff dff_A_gtbTygPp0_0(.dout(w_dff_A_XiUTjsH41_0),.din(w_dff_A_gtbTygPp0_0),.clk(gclk));
	jdff dff_A_gooogi1N5_0(.dout(w_dff_A_gtbTygPp0_0),.din(w_dff_A_gooogi1N5_0),.clk(gclk));
	jdff dff_A_HBRPOocA4_0(.dout(w_dff_A_gooogi1N5_0),.din(w_dff_A_HBRPOocA4_0),.clk(gclk));
	jdff dff_A_aCFXkw709_0(.dout(w_dff_A_HBRPOocA4_0),.din(w_dff_A_aCFXkw709_0),.clk(gclk));
	jdff dff_A_ANDoUeuS0_0(.dout(w_dff_A_aCFXkw709_0),.din(w_dff_A_ANDoUeuS0_0),.clk(gclk));
	jdff dff_A_wekDcAyI7_0(.dout(w_dff_A_ANDoUeuS0_0),.din(w_dff_A_wekDcAyI7_0),.clk(gclk));
	jdff dff_A_CTImzvee0_0(.dout(w_dff_A_wekDcAyI7_0),.din(w_dff_A_CTImzvee0_0),.clk(gclk));
	jdff dff_A_Y9dxx01h4_0(.dout(w_dff_A_CTImzvee0_0),.din(w_dff_A_Y9dxx01h4_0),.clk(gclk));
	jdff dff_A_k1YFpIgV5_0(.dout(w_dff_A_Y9dxx01h4_0),.din(w_dff_A_k1YFpIgV5_0),.clk(gclk));
	jdff dff_A_OZ1jnFH57_0(.dout(w_dff_A_k1YFpIgV5_0),.din(w_dff_A_OZ1jnFH57_0),.clk(gclk));
	jdff dff_A_TGrAQ5lS2_0(.dout(w_dff_A_OZ1jnFH57_0),.din(w_dff_A_TGrAQ5lS2_0),.clk(gclk));
	jdff dff_A_KiiWh2s00_0(.dout(w_dff_A_TGrAQ5lS2_0),.din(w_dff_A_KiiWh2s00_0),.clk(gclk));
	jdff dff_A_ENa69U1Q8_0(.dout(w_dff_A_KiiWh2s00_0),.din(w_dff_A_ENa69U1Q8_0),.clk(gclk));
	jdff dff_A_63eRILzb9_0(.dout(w_dff_A_ENa69U1Q8_0),.din(w_dff_A_63eRILzb9_0),.clk(gclk));
	jdff dff_A_unOqZuzV5_0(.dout(w_dff_A_63eRILzb9_0),.din(w_dff_A_unOqZuzV5_0),.clk(gclk));
	jdff dff_A_RKaJPw4R7_0(.dout(w_dff_A_unOqZuzV5_0),.din(w_dff_A_RKaJPw4R7_0),.clk(gclk));
	jdff dff_B_V5IEzLUR7_1(.din(n1697),.dout(w_dff_B_V5IEzLUR7_1),.clk(gclk));
	jdff dff_B_mPCpRXV06_1(.din(w_dff_B_V5IEzLUR7_1),.dout(w_dff_B_mPCpRXV06_1),.clk(gclk));
	jdff dff_B_e5LCxlWi4_1(.din(w_dff_B_mPCpRXV06_1),.dout(w_dff_B_e5LCxlWi4_1),.clk(gclk));
	jdff dff_B_zFn0wqg06_1(.din(w_dff_B_e5LCxlWi4_1),.dout(w_dff_B_zFn0wqg06_1),.clk(gclk));
	jdff dff_B_qkSi2MYM9_1(.din(w_dff_B_zFn0wqg06_1),.dout(w_dff_B_qkSi2MYM9_1),.clk(gclk));
	jdff dff_B_RFCJQDYN4_1(.din(w_dff_B_qkSi2MYM9_1),.dout(w_dff_B_RFCJQDYN4_1),.clk(gclk));
	jdff dff_B_aGSDuVwD1_1(.din(w_dff_B_RFCJQDYN4_1),.dout(w_dff_B_aGSDuVwD1_1),.clk(gclk));
	jdff dff_B_44izKsrk1_1(.din(w_dff_B_aGSDuVwD1_1),.dout(w_dff_B_44izKsrk1_1),.clk(gclk));
	jdff dff_B_E547pxtW2_1(.din(w_dff_B_44izKsrk1_1),.dout(w_dff_B_E547pxtW2_1),.clk(gclk));
	jdff dff_B_uiHgqJJs2_1(.din(w_dff_B_E547pxtW2_1),.dout(w_dff_B_uiHgqJJs2_1),.clk(gclk));
	jdff dff_B_tR5xXrwi6_1(.din(w_dff_B_uiHgqJJs2_1),.dout(w_dff_B_tR5xXrwi6_1),.clk(gclk));
	jdff dff_B_YeaBm7T12_1(.din(w_dff_B_tR5xXrwi6_1),.dout(w_dff_B_YeaBm7T12_1),.clk(gclk));
	jdff dff_B_U7y8yZsP7_1(.din(w_dff_B_YeaBm7T12_1),.dout(w_dff_B_U7y8yZsP7_1),.clk(gclk));
	jdff dff_B_tgNOku393_1(.din(w_dff_B_U7y8yZsP7_1),.dout(w_dff_B_tgNOku393_1),.clk(gclk));
	jdff dff_B_QF3v6Wca2_1(.din(w_dff_B_tgNOku393_1),.dout(w_dff_B_QF3v6Wca2_1),.clk(gclk));
	jdff dff_B_DdqiYxiA1_1(.din(w_dff_B_QF3v6Wca2_1),.dout(w_dff_B_DdqiYxiA1_1),.clk(gclk));
	jdff dff_B_HyoYCgQw7_1(.din(w_dff_B_DdqiYxiA1_1),.dout(w_dff_B_HyoYCgQw7_1),.clk(gclk));
	jdff dff_B_gshcjvz24_1(.din(w_dff_B_HyoYCgQw7_1),.dout(w_dff_B_gshcjvz24_1),.clk(gclk));
	jdff dff_B_xZjGJMqp0_1(.din(w_dff_B_gshcjvz24_1),.dout(w_dff_B_xZjGJMqp0_1),.clk(gclk));
	jdff dff_B_KDpoq9PG1_1(.din(w_dff_B_xZjGJMqp0_1),.dout(w_dff_B_KDpoq9PG1_1),.clk(gclk));
	jdff dff_B_KhEpIVJg3_1(.din(w_dff_B_KDpoq9PG1_1),.dout(w_dff_B_KhEpIVJg3_1),.clk(gclk));
	jdff dff_B_OfLo8Dwn5_1(.din(w_dff_B_KhEpIVJg3_1),.dout(w_dff_B_OfLo8Dwn5_1),.clk(gclk));
	jdff dff_B_avnGWs4K3_1(.din(w_dff_B_OfLo8Dwn5_1),.dout(w_dff_B_avnGWs4K3_1),.clk(gclk));
	jdff dff_B_fI9Ko6vw1_1(.din(n1700),.dout(w_dff_B_fI9Ko6vw1_1),.clk(gclk));
	jdff dff_B_cGurmsCa7_1(.din(w_dff_B_fI9Ko6vw1_1),.dout(w_dff_B_cGurmsCa7_1),.clk(gclk));
	jdff dff_B_RNWimfls4_1(.din(w_dff_B_cGurmsCa7_1),.dout(w_dff_B_RNWimfls4_1),.clk(gclk));
	jdff dff_B_0v12PZQq4_1(.din(w_dff_B_RNWimfls4_1),.dout(w_dff_B_0v12PZQq4_1),.clk(gclk));
	jdff dff_B_ahKwhzbV6_1(.din(w_dff_B_0v12PZQq4_1),.dout(w_dff_B_ahKwhzbV6_1),.clk(gclk));
	jdff dff_B_1CJMlBrW8_1(.din(w_dff_B_ahKwhzbV6_1),.dout(w_dff_B_1CJMlBrW8_1),.clk(gclk));
	jdff dff_B_MUvRWufT2_1(.din(w_dff_B_1CJMlBrW8_1),.dout(w_dff_B_MUvRWufT2_1),.clk(gclk));
	jdff dff_B_mB18wU551_1(.din(w_dff_B_MUvRWufT2_1),.dout(w_dff_B_mB18wU551_1),.clk(gclk));
	jdff dff_B_BzJcBxKf6_1(.din(w_dff_B_mB18wU551_1),.dout(w_dff_B_BzJcBxKf6_1),.clk(gclk));
	jdff dff_B_Rgw8ftP25_1(.din(w_dff_B_BzJcBxKf6_1),.dout(w_dff_B_Rgw8ftP25_1),.clk(gclk));
	jdff dff_B_6C5fKtuJ2_1(.din(w_dff_B_Rgw8ftP25_1),.dout(w_dff_B_6C5fKtuJ2_1),.clk(gclk));
	jdff dff_B_TunFiVrq0_1(.din(w_dff_B_6C5fKtuJ2_1),.dout(w_dff_B_TunFiVrq0_1),.clk(gclk));
	jdff dff_B_dx4Mnm3x1_1(.din(w_dff_B_TunFiVrq0_1),.dout(w_dff_B_dx4Mnm3x1_1),.clk(gclk));
	jdff dff_B_n6thTjlm9_1(.din(w_dff_B_dx4Mnm3x1_1),.dout(w_dff_B_n6thTjlm9_1),.clk(gclk));
	jdff dff_B_7HXIOS9H0_1(.din(w_dff_B_n6thTjlm9_1),.dout(w_dff_B_7HXIOS9H0_1),.clk(gclk));
	jdff dff_B_CFtJtP666_1(.din(w_dff_B_7HXIOS9H0_1),.dout(w_dff_B_CFtJtP666_1),.clk(gclk));
	jdff dff_B_MzpXaZU74_1(.din(w_dff_B_CFtJtP666_1),.dout(w_dff_B_MzpXaZU74_1),.clk(gclk));
	jdff dff_B_2kJT5lgh8_1(.din(w_dff_B_MzpXaZU74_1),.dout(w_dff_B_2kJT5lgh8_1),.clk(gclk));
	jdff dff_B_pxF6YiMo0_1(.din(w_dff_B_2kJT5lgh8_1),.dout(w_dff_B_pxF6YiMo0_1),.clk(gclk));
	jdff dff_B_j3YVEVL78_1(.din(w_dff_B_pxF6YiMo0_1),.dout(w_dff_B_j3YVEVL78_1),.clk(gclk));
	jdff dff_B_CohgHBSY3_1(.din(w_dff_B_j3YVEVL78_1),.dout(w_dff_B_CohgHBSY3_1),.clk(gclk));
	jdff dff_B_wFekHFN83_1(.din(n1701),.dout(w_dff_B_wFekHFN83_1),.clk(gclk));
	jdff dff_A_rVNUCMms5_0(.dout(w_n993_4[0]),.din(w_dff_A_rVNUCMms5_0),.clk(gclk));
	jdff dff_A_xttwV3ie8_0(.dout(w_dff_A_rVNUCMms5_0),.din(w_dff_A_xttwV3ie8_0),.clk(gclk));
	jdff dff_A_qSmVgy6h2_0(.dout(w_dff_A_xttwV3ie8_0),.din(w_dff_A_qSmVgy6h2_0),.clk(gclk));
	jdff dff_A_f7GXBkXS7_0(.dout(w_dff_A_qSmVgy6h2_0),.din(w_dff_A_f7GXBkXS7_0),.clk(gclk));
	jdff dff_A_WmN2Cb3x5_0(.dout(w_dff_A_f7GXBkXS7_0),.din(w_dff_A_WmN2Cb3x5_0),.clk(gclk));
	jdff dff_A_L4LmGRfS0_0(.dout(w_dff_A_WmN2Cb3x5_0),.din(w_dff_A_L4LmGRfS0_0),.clk(gclk));
	jdff dff_A_hCZfusYl8_0(.dout(w_dff_A_L4LmGRfS0_0),.din(w_dff_A_hCZfusYl8_0),.clk(gclk));
	jdff dff_A_UKfEVYh58_0(.dout(w_dff_A_hCZfusYl8_0),.din(w_dff_A_UKfEVYh58_0),.clk(gclk));
	jdff dff_A_iL6KFSsh0_0(.dout(w_dff_A_UKfEVYh58_0),.din(w_dff_A_iL6KFSsh0_0),.clk(gclk));
	jdff dff_A_y2aSF4gJ6_0(.dout(w_dff_A_iL6KFSsh0_0),.din(w_dff_A_y2aSF4gJ6_0),.clk(gclk));
	jdff dff_A_oK217UZV7_0(.dout(w_dff_A_y2aSF4gJ6_0),.din(w_dff_A_oK217UZV7_0),.clk(gclk));
	jdff dff_A_mdEpUr4E1_0(.dout(w_dff_A_oK217UZV7_0),.din(w_dff_A_mdEpUr4E1_0),.clk(gclk));
	jdff dff_A_9Drrbq1Y8_0(.dout(w_dff_A_mdEpUr4E1_0),.din(w_dff_A_9Drrbq1Y8_0),.clk(gclk));
	jdff dff_A_erbST0ow0_0(.dout(w_dff_A_9Drrbq1Y8_0),.din(w_dff_A_erbST0ow0_0),.clk(gclk));
	jdff dff_A_qSpU3F0Z5_0(.dout(w_dff_A_erbST0ow0_0),.din(w_dff_A_qSpU3F0Z5_0),.clk(gclk));
	jdff dff_A_5dPsLluu0_1(.dout(w_n993_4[1]),.din(w_dff_A_5dPsLluu0_1),.clk(gclk));
	jdff dff_A_bFvlcNX67_1(.dout(w_dff_A_5dPsLluu0_1),.din(w_dff_A_bFvlcNX67_1),.clk(gclk));
	jdff dff_A_T4R624mE2_1(.dout(w_dff_A_bFvlcNX67_1),.din(w_dff_A_T4R624mE2_1),.clk(gclk));
	jdff dff_A_qFgXLMG63_1(.dout(w_dff_A_T4R624mE2_1),.din(w_dff_A_qFgXLMG63_1),.clk(gclk));
	jdff dff_A_nm154Df46_1(.dout(w_dff_A_qFgXLMG63_1),.din(w_dff_A_nm154Df46_1),.clk(gclk));
	jdff dff_A_t7pXmoyr7_1(.dout(w_dff_A_nm154Df46_1),.din(w_dff_A_t7pXmoyr7_1),.clk(gclk));
	jdff dff_A_n0TdrATN1_1(.dout(w_dff_A_t7pXmoyr7_1),.din(w_dff_A_n0TdrATN1_1),.clk(gclk));
	jdff dff_A_mSYTnBfQ8_1(.dout(w_dff_A_n0TdrATN1_1),.din(w_dff_A_mSYTnBfQ8_1),.clk(gclk));
	jdff dff_A_7crUjiHr3_1(.dout(w_dff_A_mSYTnBfQ8_1),.din(w_dff_A_7crUjiHr3_1),.clk(gclk));
	jdff dff_A_NkslOwSe4_1(.dout(w_dff_A_7crUjiHr3_1),.din(w_dff_A_NkslOwSe4_1),.clk(gclk));
	jdff dff_A_u3Z345Or9_1(.dout(w_n993_1[1]),.din(w_dff_A_u3Z345Or9_1),.clk(gclk));
	jdff dff_A_TtrAxRY82_1(.dout(w_dff_A_u3Z345Or9_1),.din(w_dff_A_TtrAxRY82_1),.clk(gclk));
	jdff dff_A_txC9NkcK5_1(.dout(w_dff_A_TtrAxRY82_1),.din(w_dff_A_txC9NkcK5_1),.clk(gclk));
	jdff dff_A_XIzIFGDj1_1(.dout(w_dff_A_txC9NkcK5_1),.din(w_dff_A_XIzIFGDj1_1),.clk(gclk));
	jdff dff_A_LSaItoaT7_1(.dout(w_dff_A_XIzIFGDj1_1),.din(w_dff_A_LSaItoaT7_1),.clk(gclk));
	jdff dff_A_LkqS6dEE0_1(.dout(w_dff_A_LSaItoaT7_1),.din(w_dff_A_LkqS6dEE0_1),.clk(gclk));
	jdff dff_A_ki2Ah21m4_1(.dout(w_dff_A_LkqS6dEE0_1),.din(w_dff_A_ki2Ah21m4_1),.clk(gclk));
	jdff dff_A_PAzOq7zy7_1(.dout(w_dff_A_ki2Ah21m4_1),.din(w_dff_A_PAzOq7zy7_1),.clk(gclk));
	jdff dff_A_zgxJgVYg7_1(.dout(w_dff_A_PAzOq7zy7_1),.din(w_dff_A_zgxJgVYg7_1),.clk(gclk));
	jdff dff_A_JWPUOYga0_1(.dout(w_dff_A_zgxJgVYg7_1),.din(w_dff_A_JWPUOYga0_1),.clk(gclk));
	jdff dff_A_erRBw8ZA6_1(.dout(w_dff_A_JWPUOYga0_1),.din(w_dff_A_erRBw8ZA6_1),.clk(gclk));
	jdff dff_A_H3IAuWaq0_1(.dout(w_dff_A_erRBw8ZA6_1),.din(w_dff_A_H3IAuWaq0_1),.clk(gclk));
	jdff dff_A_ujSvXf4I7_1(.dout(w_dff_A_H3IAuWaq0_1),.din(w_dff_A_ujSvXf4I7_1),.clk(gclk));
	jdff dff_A_QLQYgiUC5_1(.dout(w_dff_A_ujSvXf4I7_1),.din(w_dff_A_QLQYgiUC5_1),.clk(gclk));
	jdff dff_A_XdriLG8E9_1(.dout(w_dff_A_QLQYgiUC5_1),.din(w_dff_A_XdriLG8E9_1),.clk(gclk));
	jdff dff_A_zLwyubXZ7_1(.dout(w_dff_A_XdriLG8E9_1),.din(w_dff_A_zLwyubXZ7_1),.clk(gclk));
	jdff dff_A_RmDAx6AT3_1(.dout(w_dff_A_zLwyubXZ7_1),.din(w_dff_A_RmDAx6AT3_1),.clk(gclk));
	jdff dff_A_ly60JqnN4_1(.dout(w_dff_A_RmDAx6AT3_1),.din(w_dff_A_ly60JqnN4_1),.clk(gclk));
	jdff dff_A_p5lmxcXw0_1(.dout(w_dff_A_ly60JqnN4_1),.din(w_dff_A_p5lmxcXw0_1),.clk(gclk));
	jdff dff_A_82lobM707_1(.dout(w_dff_A_p5lmxcXw0_1),.din(w_dff_A_82lobM707_1),.clk(gclk));
	jdff dff_A_xn1HbwAj0_1(.dout(w_dff_A_82lobM707_1),.din(w_dff_A_xn1HbwAj0_1),.clk(gclk));
	jdff dff_A_bnPiJUJk7_2(.dout(w_n993_1[2]),.din(w_dff_A_bnPiJUJk7_2),.clk(gclk));
	jdff dff_A_kDyCWJqk4_2(.dout(w_dff_A_bnPiJUJk7_2),.din(w_dff_A_kDyCWJqk4_2),.clk(gclk));
	jdff dff_A_vd3u4Ewu0_2(.dout(w_dff_A_kDyCWJqk4_2),.din(w_dff_A_vd3u4Ewu0_2),.clk(gclk));
	jdff dff_A_MZ8MXjhX5_2(.dout(w_dff_A_vd3u4Ewu0_2),.din(w_dff_A_MZ8MXjhX5_2),.clk(gclk));
	jdff dff_A_1FKVDn6M2_2(.dout(w_dff_A_MZ8MXjhX5_2),.din(w_dff_A_1FKVDn6M2_2),.clk(gclk));
	jdff dff_A_zyDbunfF3_2(.dout(w_dff_A_1FKVDn6M2_2),.din(w_dff_A_zyDbunfF3_2),.clk(gclk));
	jdff dff_A_NGDH3qGO0_2(.dout(w_dff_A_zyDbunfF3_2),.din(w_dff_A_NGDH3qGO0_2),.clk(gclk));
	jdff dff_A_ByRyP1HW5_2(.dout(w_dff_A_NGDH3qGO0_2),.din(w_dff_A_ByRyP1HW5_2),.clk(gclk));
	jdff dff_A_fzrE1owu5_2(.dout(w_dff_A_ByRyP1HW5_2),.din(w_dff_A_fzrE1owu5_2),.clk(gclk));
	jdff dff_A_29yt73si3_2(.dout(w_dff_A_fzrE1owu5_2),.din(w_dff_A_29yt73si3_2),.clk(gclk));
	jdff dff_A_D2E6zgTh5_2(.dout(w_dff_A_29yt73si3_2),.din(w_dff_A_D2E6zgTh5_2),.clk(gclk));
	jdff dff_A_oynphTOB3_2(.dout(w_dff_A_D2E6zgTh5_2),.din(w_dff_A_oynphTOB3_2),.clk(gclk));
	jdff dff_A_Rc4Jnk2v7_2(.dout(w_dff_A_oynphTOB3_2),.din(w_dff_A_Rc4Jnk2v7_2),.clk(gclk));
	jdff dff_A_PAIISbnq6_2(.dout(w_dff_A_Rc4Jnk2v7_2),.din(w_dff_A_PAIISbnq6_2),.clk(gclk));
	jdff dff_A_YlBmGZHh2_2(.dout(w_dff_A_PAIISbnq6_2),.din(w_dff_A_YlBmGZHh2_2),.clk(gclk));
	jdff dff_A_kXSJXCrt9_2(.dout(w_dff_A_YlBmGZHh2_2),.din(w_dff_A_kXSJXCrt9_2),.clk(gclk));
	jdff dff_A_22DRyuHC2_2(.dout(w_dff_A_kXSJXCrt9_2),.din(w_dff_A_22DRyuHC2_2),.clk(gclk));
	jdff dff_A_yffEAbKz6_2(.dout(w_dff_A_22DRyuHC2_2),.din(w_dff_A_yffEAbKz6_2),.clk(gclk));
	jdff dff_A_8OLMbiwS5_2(.dout(w_dff_A_yffEAbKz6_2),.din(w_dff_A_8OLMbiwS5_2),.clk(gclk));
	jdff dff_A_iBDS9ARQ2_2(.dout(w_dff_A_8OLMbiwS5_2),.din(w_dff_A_iBDS9ARQ2_2),.clk(gclk));
	jdff dff_A_vCyZFVoO5_1(.dout(w_n993_0[1]),.din(w_dff_A_vCyZFVoO5_1),.clk(gclk));
	jdff dff_A_nETcOfKL1_1(.dout(w_dff_A_vCyZFVoO5_1),.din(w_dff_A_nETcOfKL1_1),.clk(gclk));
	jdff dff_A_ENashX1U6_1(.dout(w_dff_A_nETcOfKL1_1),.din(w_dff_A_ENashX1U6_1),.clk(gclk));
	jdff dff_A_8ls4io8I3_1(.dout(w_dff_A_ENashX1U6_1),.din(w_dff_A_8ls4io8I3_1),.clk(gclk));
	jdff dff_A_mq01duzk5_1(.dout(w_dff_A_8ls4io8I3_1),.din(w_dff_A_mq01duzk5_1),.clk(gclk));
	jdff dff_A_0XkUD5EV1_1(.dout(w_dff_A_mq01duzk5_1),.din(w_dff_A_0XkUD5EV1_1),.clk(gclk));
	jdff dff_A_lwhZMMEm0_1(.dout(w_dff_A_0XkUD5EV1_1),.din(w_dff_A_lwhZMMEm0_1),.clk(gclk));
	jdff dff_A_WnNnlVG17_1(.dout(w_dff_A_lwhZMMEm0_1),.din(w_dff_A_WnNnlVG17_1),.clk(gclk));
	jdff dff_A_KhjNfNI49_1(.dout(w_dff_A_WnNnlVG17_1),.din(w_dff_A_KhjNfNI49_1),.clk(gclk));
	jdff dff_A_H3VbJS9q1_1(.dout(w_dff_A_KhjNfNI49_1),.din(w_dff_A_H3VbJS9q1_1),.clk(gclk));
	jdff dff_A_Awc6SkHf0_1(.dout(w_dff_A_H3VbJS9q1_1),.din(w_dff_A_Awc6SkHf0_1),.clk(gclk));
	jdff dff_A_nOo7LMw46_1(.dout(w_dff_A_Awc6SkHf0_1),.din(w_dff_A_nOo7LMw46_1),.clk(gclk));
	jdff dff_A_nJijrz1b1_1(.dout(w_dff_A_nOo7LMw46_1),.din(w_dff_A_nJijrz1b1_1),.clk(gclk));
	jdff dff_A_PfiBgvRn6_1(.dout(w_dff_A_nJijrz1b1_1),.din(w_dff_A_PfiBgvRn6_1),.clk(gclk));
	jdff dff_A_N2jZG2ad6_1(.dout(w_dff_A_PfiBgvRn6_1),.din(w_dff_A_N2jZG2ad6_1),.clk(gclk));
	jdff dff_A_crpsK3c79_1(.dout(w_dff_A_N2jZG2ad6_1),.din(w_dff_A_crpsK3c79_1),.clk(gclk));
	jdff dff_A_lw8G4GUT8_1(.dout(w_dff_A_crpsK3c79_1),.din(w_dff_A_lw8G4GUT8_1),.clk(gclk));
	jdff dff_A_NMehygOp9_1(.dout(w_dff_A_lw8G4GUT8_1),.din(w_dff_A_NMehygOp9_1),.clk(gclk));
	jdff dff_A_LgrVplrC2_2(.dout(w_n993_0[2]),.din(w_dff_A_LgrVplrC2_2),.clk(gclk));
	jdff dff_A_3gMgaEEW0_2(.dout(w_dff_A_LgrVplrC2_2),.din(w_dff_A_3gMgaEEW0_2),.clk(gclk));
	jdff dff_A_y80IbRP17_2(.dout(w_dff_A_3gMgaEEW0_2),.din(w_dff_A_y80IbRP17_2),.clk(gclk));
	jdff dff_A_diOxwtbg9_2(.dout(w_dff_A_y80IbRP17_2),.din(w_dff_A_diOxwtbg9_2),.clk(gclk));
	jdff dff_A_qqOvGl9I9_2(.dout(w_dff_A_diOxwtbg9_2),.din(w_dff_A_qqOvGl9I9_2),.clk(gclk));
	jdff dff_A_T73MkNtP6_2(.dout(w_dff_A_qqOvGl9I9_2),.din(w_dff_A_T73MkNtP6_2),.clk(gclk));
	jdff dff_A_aHvX8tWT8_2(.dout(w_dff_A_T73MkNtP6_2),.din(w_dff_A_aHvX8tWT8_2),.clk(gclk));
	jdff dff_A_IZ0J4Get0_2(.dout(w_dff_A_aHvX8tWT8_2),.din(w_dff_A_IZ0J4Get0_2),.clk(gclk));
	jdff dff_A_9rRmXcKe0_2(.dout(w_dff_A_IZ0J4Get0_2),.din(w_dff_A_9rRmXcKe0_2),.clk(gclk));
	jdff dff_A_ADELT7Vs8_2(.dout(w_dff_A_9rRmXcKe0_2),.din(w_dff_A_ADELT7Vs8_2),.clk(gclk));
	jdff dff_A_olEYvere9_2(.dout(w_dff_A_ADELT7Vs8_2),.din(w_dff_A_olEYvere9_2),.clk(gclk));
	jdff dff_A_c6VJc8HF5_1(.dout(w_G1690_1[1]),.din(w_dff_A_c6VJc8HF5_1),.clk(gclk));
	jdff dff_A_s0Hg9CDf6_1(.dout(w_G1690_0[1]),.din(w_dff_A_s0Hg9CDf6_1),.clk(gclk));
	jdff dff_A_b7N5FImU1_1(.dout(w_dff_A_s0Hg9CDf6_1),.din(w_dff_A_b7N5FImU1_1),.clk(gclk));
	jdff dff_A_RpfOhTvr0_1(.dout(w_dff_A_b7N5FImU1_1),.din(w_dff_A_RpfOhTvr0_1),.clk(gclk));
	jdff dff_A_UzgRR4S39_1(.dout(w_dff_A_RpfOhTvr0_1),.din(w_dff_A_UzgRR4S39_1),.clk(gclk));
	jdff dff_A_v8lotj2U9_1(.dout(w_dff_A_UzgRR4S39_1),.din(w_dff_A_v8lotj2U9_1),.clk(gclk));
	jdff dff_A_n4rH0UBr1_1(.dout(w_dff_A_v8lotj2U9_1),.din(w_dff_A_n4rH0UBr1_1),.clk(gclk));
	jdff dff_A_CrecUhpv0_1(.dout(w_dff_A_n4rH0UBr1_1),.din(w_dff_A_CrecUhpv0_1),.clk(gclk));
	jdff dff_A_jmVhB9PT8_1(.dout(w_dff_A_CrecUhpv0_1),.din(w_dff_A_jmVhB9PT8_1),.clk(gclk));
	jdff dff_A_LeyYPWqk5_1(.dout(w_dff_A_jmVhB9PT8_1),.din(w_dff_A_LeyYPWqk5_1),.clk(gclk));
	jdff dff_A_nqwXVtt81_1(.dout(w_dff_A_LeyYPWqk5_1),.din(w_dff_A_nqwXVtt81_1),.clk(gclk));
	jdff dff_A_T4CLY8gb3_1(.dout(w_dff_A_nqwXVtt81_1),.din(w_dff_A_T4CLY8gb3_1),.clk(gclk));
	jdff dff_A_CF1l3lga2_1(.dout(w_dff_A_T4CLY8gb3_1),.din(w_dff_A_CF1l3lga2_1),.clk(gclk));
	jdff dff_A_pOBdfCEK3_1(.dout(w_dff_A_CF1l3lga2_1),.din(w_dff_A_pOBdfCEK3_1),.clk(gclk));
	jdff dff_A_VCaThd1q3_1(.dout(w_dff_A_pOBdfCEK3_1),.din(w_dff_A_VCaThd1q3_1),.clk(gclk));
	jdff dff_A_j2p6vO1V5_1(.dout(w_dff_A_VCaThd1q3_1),.din(w_dff_A_j2p6vO1V5_1),.clk(gclk));
	jdff dff_A_H1aFAhHN5_1(.dout(w_dff_A_j2p6vO1V5_1),.din(w_dff_A_H1aFAhHN5_1),.clk(gclk));
	jdff dff_A_OkzwuYIS6_1(.dout(w_dff_A_H1aFAhHN5_1),.din(w_dff_A_OkzwuYIS6_1),.clk(gclk));
	jdff dff_A_Sgz9I38z2_1(.dout(w_dff_A_OkzwuYIS6_1),.din(w_dff_A_Sgz9I38z2_1),.clk(gclk));
	jdff dff_A_ngBRyqUN4_1(.dout(w_dff_A_Sgz9I38z2_1),.din(w_dff_A_ngBRyqUN4_1),.clk(gclk));
	jdff dff_A_4kfIcUqA6_1(.dout(w_dff_A_ngBRyqUN4_1),.din(w_dff_A_4kfIcUqA6_1),.clk(gclk));
	jdff dff_A_XLlFqoxv0_1(.dout(w_dff_A_4kfIcUqA6_1),.din(w_dff_A_XLlFqoxv0_1),.clk(gclk));
	jdff dff_A_jEYaMwoB4_1(.dout(w_dff_A_XLlFqoxv0_1),.din(w_dff_A_jEYaMwoB4_1),.clk(gclk));
	jdff dff_A_XlP6CFhZ0_1(.dout(w_dff_A_jEYaMwoB4_1),.din(w_dff_A_XlP6CFhZ0_1),.clk(gclk));
	jdff dff_A_rNuAEmgB4_0(.dout(w_G1689_1[0]),.din(w_dff_A_rNuAEmgB4_0),.clk(gclk));
	jdff dff_A_bb7qMjrM9_0(.dout(w_dff_A_rNuAEmgB4_0),.din(w_dff_A_bb7qMjrM9_0),.clk(gclk));
	jdff dff_A_ygWYn2bj3_0(.dout(w_dff_A_bb7qMjrM9_0),.din(w_dff_A_ygWYn2bj3_0),.clk(gclk));
	jdff dff_A_d99eG6Th8_0(.dout(w_dff_A_ygWYn2bj3_0),.din(w_dff_A_d99eG6Th8_0),.clk(gclk));
	jdff dff_A_aHLTcKNW6_0(.dout(w_dff_A_d99eG6Th8_0),.din(w_dff_A_aHLTcKNW6_0),.clk(gclk));
	jdff dff_A_FvzwZuTH2_0(.dout(w_dff_A_aHLTcKNW6_0),.din(w_dff_A_FvzwZuTH2_0),.clk(gclk));
	jdff dff_A_WSVK0JUb1_0(.dout(w_dff_A_FvzwZuTH2_0),.din(w_dff_A_WSVK0JUb1_0),.clk(gclk));
	jdff dff_A_mbmiZXFa9_0(.dout(w_dff_A_WSVK0JUb1_0),.din(w_dff_A_mbmiZXFa9_0),.clk(gclk));
	jdff dff_A_b7Fpg7u54_0(.dout(w_dff_A_mbmiZXFa9_0),.din(w_dff_A_b7Fpg7u54_0),.clk(gclk));
	jdff dff_A_xKwHvcxb9_2(.dout(w_G1689_1[2]),.din(w_dff_A_xKwHvcxb9_2),.clk(gclk));
	jdff dff_A_Ls7O1bV69_2(.dout(w_dff_A_xKwHvcxb9_2),.din(w_dff_A_Ls7O1bV69_2),.clk(gclk));
	jdff dff_A_Z57ELrXu0_2(.dout(w_dff_A_Ls7O1bV69_2),.din(w_dff_A_Z57ELrXu0_2),.clk(gclk));
	jdff dff_A_l69HWdEl6_2(.dout(w_dff_A_Z57ELrXu0_2),.din(w_dff_A_l69HWdEl6_2),.clk(gclk));
	jdff dff_A_shQhlWKM6_2(.dout(w_dff_A_l69HWdEl6_2),.din(w_dff_A_shQhlWKM6_2),.clk(gclk));
	jdff dff_A_5WLz3xtU3_2(.dout(w_dff_A_shQhlWKM6_2),.din(w_dff_A_5WLz3xtU3_2),.clk(gclk));
	jdff dff_A_DBsOnch54_2(.dout(w_dff_A_5WLz3xtU3_2),.din(w_dff_A_DBsOnch54_2),.clk(gclk));
	jdff dff_A_mhquwqu78_2(.dout(w_dff_A_DBsOnch54_2),.din(w_dff_A_mhquwqu78_2),.clk(gclk));
	jdff dff_A_Y7xX38H71_2(.dout(w_dff_A_mhquwqu78_2),.din(w_dff_A_Y7xX38H71_2),.clk(gclk));
	jdff dff_A_Xpbvfbj07_2(.dout(w_dff_A_Y7xX38H71_2),.din(w_dff_A_Xpbvfbj07_2),.clk(gclk));
	jdff dff_A_LGSoJkVR4_2(.dout(w_dff_A_Xpbvfbj07_2),.din(w_dff_A_LGSoJkVR4_2),.clk(gclk));
	jdff dff_A_lFyJjsoJ0_2(.dout(w_dff_A_LGSoJkVR4_2),.din(w_dff_A_lFyJjsoJ0_2),.clk(gclk));
	jdff dff_A_4W665TrL5_2(.dout(w_dff_A_lFyJjsoJ0_2),.din(w_dff_A_4W665TrL5_2),.clk(gclk));
	jdff dff_A_vj2p8AEF5_2(.dout(w_dff_A_4W665TrL5_2),.din(w_dff_A_vj2p8AEF5_2),.clk(gclk));
	jdff dff_A_yvttYkk23_2(.dout(w_dff_A_vj2p8AEF5_2),.din(w_dff_A_yvttYkk23_2),.clk(gclk));
	jdff dff_A_6FdwXwMG7_2(.dout(w_dff_A_yvttYkk23_2),.din(w_dff_A_6FdwXwMG7_2),.clk(gclk));
	jdff dff_A_VkLc473u6_2(.dout(w_dff_A_6FdwXwMG7_2),.din(w_dff_A_VkLc473u6_2),.clk(gclk));
	jdff dff_A_4DUptWGz8_2(.dout(w_dff_A_VkLc473u6_2),.din(w_dff_A_4DUptWGz8_2),.clk(gclk));
	jdff dff_A_xWT9hROC2_2(.dout(w_dff_A_4DUptWGz8_2),.din(w_dff_A_xWT9hROC2_2),.clk(gclk));
	jdff dff_A_UXWckWh10_2(.dout(w_dff_A_xWT9hROC2_2),.din(w_dff_A_UXWckWh10_2),.clk(gclk));
	jdff dff_A_EV9tojrg9_2(.dout(w_dff_A_UXWckWh10_2),.din(w_dff_A_EV9tojrg9_2),.clk(gclk));
	jdff dff_A_Kyriajg40_2(.dout(w_dff_A_EV9tojrg9_2),.din(w_dff_A_Kyriajg40_2),.clk(gclk));
	jdff dff_A_yBqaRBxN0_1(.dout(w_G1689_0[1]),.din(w_dff_A_yBqaRBxN0_1),.clk(gclk));
	jdff dff_A_neSukdh07_1(.dout(w_dff_A_yBqaRBxN0_1),.din(w_dff_A_neSukdh07_1),.clk(gclk));
	jdff dff_A_cJPdEet27_1(.dout(w_dff_A_neSukdh07_1),.din(w_dff_A_cJPdEet27_1),.clk(gclk));
	jdff dff_A_ZQiGzv119_1(.dout(w_dff_A_cJPdEet27_1),.din(w_dff_A_ZQiGzv119_1),.clk(gclk));
	jdff dff_A_crFJutxU7_1(.dout(w_dff_A_ZQiGzv119_1),.din(w_dff_A_crFJutxU7_1),.clk(gclk));
	jdff dff_A_KKTRLcsr4_1(.dout(w_dff_A_crFJutxU7_1),.din(w_dff_A_KKTRLcsr4_1),.clk(gclk));
	jdff dff_A_wQQQCS093_1(.dout(w_dff_A_KKTRLcsr4_1),.din(w_dff_A_wQQQCS093_1),.clk(gclk));
	jdff dff_A_VmCq3Nf10_1(.dout(w_dff_A_wQQQCS093_1),.din(w_dff_A_VmCq3Nf10_1),.clk(gclk));
	jdff dff_A_g2h8skqp7_1(.dout(w_dff_A_VmCq3Nf10_1),.din(w_dff_A_g2h8skqp7_1),.clk(gclk));
	jdff dff_A_IKmsPhYd5_1(.dout(w_dff_A_g2h8skqp7_1),.din(w_dff_A_IKmsPhYd5_1),.clk(gclk));
	jdff dff_A_ubDseIHZ2_1(.dout(w_dff_A_IKmsPhYd5_1),.din(w_dff_A_ubDseIHZ2_1),.clk(gclk));
	jdff dff_A_YMi0R8rh5_1(.dout(w_dff_A_ubDseIHZ2_1),.din(w_dff_A_YMi0R8rh5_1),.clk(gclk));
	jdff dff_A_3nbfTjjo9_1(.dout(w_dff_A_YMi0R8rh5_1),.din(w_dff_A_3nbfTjjo9_1),.clk(gclk));
	jdff dff_A_wZuxnlWM7_1(.dout(w_dff_A_3nbfTjjo9_1),.din(w_dff_A_wZuxnlWM7_1),.clk(gclk));
	jdff dff_A_ZP6roR749_1(.dout(w_dff_A_wZuxnlWM7_1),.din(w_dff_A_ZP6roR749_1),.clk(gclk));
	jdff dff_A_HAouYHwE8_1(.dout(w_dff_A_ZP6roR749_1),.din(w_dff_A_HAouYHwE8_1),.clk(gclk));
	jdff dff_A_ukfZl4yL8_1(.dout(w_dff_A_HAouYHwE8_1),.din(w_dff_A_ukfZl4yL8_1),.clk(gclk));
	jdff dff_A_UarNc1l53_1(.dout(w_dff_A_ukfZl4yL8_1),.din(w_dff_A_UarNc1l53_1),.clk(gclk));
	jdff dff_A_v8UhOTPX0_1(.dout(w_dff_A_UarNc1l53_1),.din(w_dff_A_v8UhOTPX0_1),.clk(gclk));
	jdff dff_A_Nfc79ZMy5_2(.dout(w_G1689_0[2]),.din(w_dff_A_Nfc79ZMy5_2),.clk(gclk));
	jdff dff_A_rvxLGAmG0_2(.dout(w_dff_A_Nfc79ZMy5_2),.din(w_dff_A_rvxLGAmG0_2),.clk(gclk));
	jdff dff_A_vxQ2Vjw62_2(.dout(w_dff_A_rvxLGAmG0_2),.din(w_dff_A_vxQ2Vjw62_2),.clk(gclk));
	jdff dff_A_aUrD6viN8_2(.dout(w_dff_A_vxQ2Vjw62_2),.din(w_dff_A_aUrD6viN8_2),.clk(gclk));
	jdff dff_A_9mzZP8q07_2(.dout(w_dff_A_aUrD6viN8_2),.din(w_dff_A_9mzZP8q07_2),.clk(gclk));
	jdff dff_A_5ozHnspx2_2(.dout(w_dff_A_9mzZP8q07_2),.din(w_dff_A_5ozHnspx2_2),.clk(gclk));
	jdff dff_A_pKXmSvw00_2(.dout(w_dff_A_5ozHnspx2_2),.din(w_dff_A_pKXmSvw00_2),.clk(gclk));
	jdff dff_A_S8Er80wL7_2(.dout(w_dff_A_pKXmSvw00_2),.din(w_dff_A_S8Er80wL7_2),.clk(gclk));
	jdff dff_A_DfSkNTJ80_2(.dout(w_dff_A_S8Er80wL7_2),.din(w_dff_A_DfSkNTJ80_2),.clk(gclk));
	jdff dff_A_i6ApMTD60_2(.dout(w_dff_A_DfSkNTJ80_2),.din(w_dff_A_i6ApMTD60_2),.clk(gclk));
	jdff dff_A_ot76YAmh8_2(.dout(w_dff_A_i6ApMTD60_2),.din(w_dff_A_ot76YAmh8_2),.clk(gclk));
	jdff dff_A_OyAR79sj4_2(.dout(w_dff_A_ot76YAmh8_2),.din(w_dff_A_OyAR79sj4_2),.clk(gclk));
	jdff dff_A_Xl6d13p94_2(.dout(w_dff_A_OyAR79sj4_2),.din(w_dff_A_Xl6d13p94_2),.clk(gclk));
	jdff dff_B_1kjSiEjw6_1(.din(n1709),.dout(w_dff_B_1kjSiEjw6_1),.clk(gclk));
	jdff dff_B_0dlhkWcu6_1(.din(w_dff_B_1kjSiEjw6_1),.dout(w_dff_B_0dlhkWcu6_1),.clk(gclk));
	jdff dff_B_sunLTnWp9_1(.din(w_dff_B_0dlhkWcu6_1),.dout(w_dff_B_sunLTnWp9_1),.clk(gclk));
	jdff dff_B_HHLt3znN7_1(.din(w_dff_B_sunLTnWp9_1),.dout(w_dff_B_HHLt3znN7_1),.clk(gclk));
	jdff dff_B_m77swa604_1(.din(w_dff_B_HHLt3znN7_1),.dout(w_dff_B_m77swa604_1),.clk(gclk));
	jdff dff_B_9Y2rnsm06_1(.din(w_dff_B_m77swa604_1),.dout(w_dff_B_9Y2rnsm06_1),.clk(gclk));
	jdff dff_B_1RUThDct8_1(.din(w_dff_B_9Y2rnsm06_1),.dout(w_dff_B_1RUThDct8_1),.clk(gclk));
	jdff dff_B_jQatCG0n3_1(.din(w_dff_B_1RUThDct8_1),.dout(w_dff_B_jQatCG0n3_1),.clk(gclk));
	jdff dff_B_7yHdn2Wc5_1(.din(w_dff_B_jQatCG0n3_1),.dout(w_dff_B_7yHdn2Wc5_1),.clk(gclk));
	jdff dff_B_NAohWdCa3_1(.din(w_dff_B_7yHdn2Wc5_1),.dout(w_dff_B_NAohWdCa3_1),.clk(gclk));
	jdff dff_B_HFvGyynk1_1(.din(w_dff_B_NAohWdCa3_1),.dout(w_dff_B_HFvGyynk1_1),.clk(gclk));
	jdff dff_B_81XKjS4J8_1(.din(w_dff_B_HFvGyynk1_1),.dout(w_dff_B_81XKjS4J8_1),.clk(gclk));
	jdff dff_B_uX0eNeH98_1(.din(w_dff_B_81XKjS4J8_1),.dout(w_dff_B_uX0eNeH98_1),.clk(gclk));
	jdff dff_B_ISoAeJD93_1(.din(w_dff_B_uX0eNeH98_1),.dout(w_dff_B_ISoAeJD93_1),.clk(gclk));
	jdff dff_B_sq8zqZoM7_1(.din(w_dff_B_ISoAeJD93_1),.dout(w_dff_B_sq8zqZoM7_1),.clk(gclk));
	jdff dff_B_EblJsutN7_1(.din(w_dff_B_sq8zqZoM7_1),.dout(w_dff_B_EblJsutN7_1),.clk(gclk));
	jdff dff_B_GNHqy0OS0_1(.din(w_dff_B_EblJsutN7_1),.dout(w_dff_B_GNHqy0OS0_1),.clk(gclk));
	jdff dff_B_cHINSXlL4_1(.din(w_dff_B_GNHqy0OS0_1),.dout(w_dff_B_cHINSXlL4_1),.clk(gclk));
	jdff dff_B_zEouXW107_1(.din(w_dff_B_cHINSXlL4_1),.dout(w_dff_B_zEouXW107_1),.clk(gclk));
	jdff dff_B_MC1CqQ0i9_1(.din(w_dff_B_zEouXW107_1),.dout(w_dff_B_MC1CqQ0i9_1),.clk(gclk));
	jdff dff_B_B2lM3Cwn0_1(.din(w_dff_B_MC1CqQ0i9_1),.dout(w_dff_B_B2lM3Cwn0_1),.clk(gclk));
	jdff dff_B_MWG9IqOL0_1(.din(w_dff_B_B2lM3Cwn0_1),.dout(w_dff_B_MWG9IqOL0_1),.clk(gclk));
	jdff dff_B_C1gAIC6b5_1(.din(w_dff_B_MWG9IqOL0_1),.dout(w_dff_B_C1gAIC6b5_1),.clk(gclk));
	jdff dff_B_lK20VBSx8_1(.din(n1711),.dout(w_dff_B_lK20VBSx8_1),.clk(gclk));
	jdff dff_B_FLJHjwzx7_1(.din(w_dff_B_lK20VBSx8_1),.dout(w_dff_B_FLJHjwzx7_1),.clk(gclk));
	jdff dff_B_rAdYT9FP7_1(.din(w_dff_B_FLJHjwzx7_1),.dout(w_dff_B_rAdYT9FP7_1),.clk(gclk));
	jdff dff_B_XRL9M5rQ4_1(.din(w_dff_B_rAdYT9FP7_1),.dout(w_dff_B_XRL9M5rQ4_1),.clk(gclk));
	jdff dff_B_W2o8yhyI6_1(.din(w_dff_B_XRL9M5rQ4_1),.dout(w_dff_B_W2o8yhyI6_1),.clk(gclk));
	jdff dff_B_TKjQU7uI1_1(.din(w_dff_B_W2o8yhyI6_1),.dout(w_dff_B_TKjQU7uI1_1),.clk(gclk));
	jdff dff_B_lE0OROBT1_1(.din(w_dff_B_TKjQU7uI1_1),.dout(w_dff_B_lE0OROBT1_1),.clk(gclk));
	jdff dff_B_rVryp8kL2_1(.din(w_dff_B_lE0OROBT1_1),.dout(w_dff_B_rVryp8kL2_1),.clk(gclk));
	jdff dff_B_qXwJEIyb8_1(.din(w_dff_B_rVryp8kL2_1),.dout(w_dff_B_qXwJEIyb8_1),.clk(gclk));
	jdff dff_B_obY4200g6_1(.din(w_dff_B_qXwJEIyb8_1),.dout(w_dff_B_obY4200g6_1),.clk(gclk));
	jdff dff_B_u3VZ3E730_1(.din(w_dff_B_obY4200g6_1),.dout(w_dff_B_u3VZ3E730_1),.clk(gclk));
	jdff dff_B_UtmfcqAP0_1(.din(w_dff_B_u3VZ3E730_1),.dout(w_dff_B_UtmfcqAP0_1),.clk(gclk));
	jdff dff_B_sJ4WLeyM0_1(.din(w_dff_B_UtmfcqAP0_1),.dout(w_dff_B_sJ4WLeyM0_1),.clk(gclk));
	jdff dff_B_vPzjLQUq4_1(.din(w_dff_B_sJ4WLeyM0_1),.dout(w_dff_B_vPzjLQUq4_1),.clk(gclk));
	jdff dff_B_ah0BjhyB9_1(.din(w_dff_B_vPzjLQUq4_1),.dout(w_dff_B_ah0BjhyB9_1),.clk(gclk));
	jdff dff_B_2TT76pLZ6_1(.din(w_dff_B_ah0BjhyB9_1),.dout(w_dff_B_2TT76pLZ6_1),.clk(gclk));
	jdff dff_B_YGxHVztd0_1(.din(w_dff_B_2TT76pLZ6_1),.dout(w_dff_B_YGxHVztd0_1),.clk(gclk));
	jdff dff_B_7ZZJBXGH0_1(.din(w_dff_B_YGxHVztd0_1),.dout(w_dff_B_7ZZJBXGH0_1),.clk(gclk));
	jdff dff_B_ACDNcCPF8_1(.din(w_dff_B_7ZZJBXGH0_1),.dout(w_dff_B_ACDNcCPF8_1),.clk(gclk));
	jdff dff_B_UFxbdRmG4_1(.din(w_dff_B_ACDNcCPF8_1),.dout(w_dff_B_UFxbdRmG4_1),.clk(gclk));
	jdff dff_B_GxSbALLt5_1(.din(w_dff_B_UFxbdRmG4_1),.dout(w_dff_B_GxSbALLt5_1),.clk(gclk));
	jdff dff_B_b5XNq4Yj5_1(.din(n1712),.dout(w_dff_B_b5XNq4Yj5_1),.clk(gclk));
	jdff dff_B_wyGLOH1w5_0(.din(n1678),.dout(w_dff_B_wyGLOH1w5_0),.clk(gclk));
	jdff dff_B_8xfjtWrt5_0(.din(w_dff_B_wyGLOH1w5_0),.dout(w_dff_B_8xfjtWrt5_0),.clk(gclk));
	jdff dff_B_18zmQWva2_0(.din(w_dff_B_8xfjtWrt5_0),.dout(w_dff_B_18zmQWva2_0),.clk(gclk));
	jdff dff_B_WMl50vtD4_0(.din(w_dff_B_18zmQWva2_0),.dout(w_dff_B_WMl50vtD4_0),.clk(gclk));
	jdff dff_B_GePLgr399_0(.din(w_dff_B_WMl50vtD4_0),.dout(w_dff_B_GePLgr399_0),.clk(gclk));
	jdff dff_B_kC4npNCu9_0(.din(w_dff_B_GePLgr399_0),.dout(w_dff_B_kC4npNCu9_0),.clk(gclk));
	jdff dff_B_fX8Rrdkf8_0(.din(w_dff_B_kC4npNCu9_0),.dout(w_dff_B_fX8Rrdkf8_0),.clk(gclk));
	jdff dff_B_qWhNQUeJ7_0(.din(w_dff_B_fX8Rrdkf8_0),.dout(w_dff_B_qWhNQUeJ7_0),.clk(gclk));
	jdff dff_B_lRtGoqTU6_0(.din(w_dff_B_qWhNQUeJ7_0),.dout(w_dff_B_lRtGoqTU6_0),.clk(gclk));
	jdff dff_B_79PgY89o7_0(.din(w_dff_B_lRtGoqTU6_0),.dout(w_dff_B_79PgY89o7_0),.clk(gclk));
	jdff dff_B_JXT4TP7N7_0(.din(w_dff_B_79PgY89o7_0),.dout(w_dff_B_JXT4TP7N7_0),.clk(gclk));
	jdff dff_B_1PXEBAQ64_0(.din(w_dff_B_JXT4TP7N7_0),.dout(w_dff_B_1PXEBAQ64_0),.clk(gclk));
	jdff dff_B_fiyiR4TN4_0(.din(w_dff_B_1PXEBAQ64_0),.dout(w_dff_B_fiyiR4TN4_0),.clk(gclk));
	jdff dff_B_Q69xA2qk9_0(.din(w_dff_B_fiyiR4TN4_0),.dout(w_dff_B_Q69xA2qk9_0),.clk(gclk));
	jdff dff_B_vcIYmIXm5_0(.din(w_dff_B_Q69xA2qk9_0),.dout(w_dff_B_vcIYmIXm5_0),.clk(gclk));
	jdff dff_B_NffOVg0X4_0(.din(w_dff_B_vcIYmIXm5_0),.dout(w_dff_B_NffOVg0X4_0),.clk(gclk));
	jdff dff_B_WzZjOkoB0_0(.din(w_dff_B_NffOVg0X4_0),.dout(w_dff_B_WzZjOkoB0_0),.clk(gclk));
	jdff dff_B_qJ6ZC2TC2_0(.din(w_dff_B_WzZjOkoB0_0),.dout(w_dff_B_qJ6ZC2TC2_0),.clk(gclk));
	jdff dff_B_RNrhA1g56_0(.din(w_dff_B_qJ6ZC2TC2_0),.dout(w_dff_B_RNrhA1g56_0),.clk(gclk));
	jdff dff_B_YC3cl44O4_0(.din(n1501),.dout(w_dff_B_YC3cl44O4_0),.clk(gclk));
	jdff dff_B_6OMTBjEN4_0(.din(w_dff_B_YC3cl44O4_0),.dout(w_dff_B_6OMTBjEN4_0),.clk(gclk));
	jdff dff_B_J3xMFMzu4_0(.din(w_dff_B_6OMTBjEN4_0),.dout(w_dff_B_J3xMFMzu4_0),.clk(gclk));
	jdff dff_B_9OHPeFdG6_0(.din(w_dff_B_J3xMFMzu4_0),.dout(w_dff_B_9OHPeFdG6_0),.clk(gclk));
	jdff dff_B_lw0hFDoO1_0(.din(w_dff_B_9OHPeFdG6_0),.dout(w_dff_B_lw0hFDoO1_0),.clk(gclk));
	jdff dff_B_5nvaracM7_0(.din(w_dff_B_lw0hFDoO1_0),.dout(w_dff_B_5nvaracM7_0),.clk(gclk));
	jdff dff_B_eHmpSaiz7_0(.din(w_dff_B_5nvaracM7_0),.dout(w_dff_B_eHmpSaiz7_0),.clk(gclk));
	jdff dff_B_ASVe7ABE1_0(.din(w_dff_B_eHmpSaiz7_0),.dout(w_dff_B_ASVe7ABE1_0),.clk(gclk));
	jdff dff_B_uBoKKbTs1_0(.din(w_dff_B_ASVe7ABE1_0),.dout(w_dff_B_uBoKKbTs1_0),.clk(gclk));
	jdff dff_B_qR3rCMT00_1(.din(n1496),.dout(w_dff_B_qR3rCMT00_1),.clk(gclk));
	jdff dff_B_pBSK8JsB7_1(.din(n413),.dout(w_dff_B_pBSK8JsB7_1),.clk(gclk));
	jdff dff_B_6UrklJ322_1(.din(w_dff_B_pBSK8JsB7_1),.dout(w_dff_B_6UrklJ322_1),.clk(gclk));
	jdff dff_A_NuoaZjgQ1_0(.dout(w_G308_1[0]),.din(w_dff_A_NuoaZjgQ1_0),.clk(gclk));
	jdff dff_B_txQzqDiA3_1(.din(n400),.dout(w_dff_B_txQzqDiA3_1),.clk(gclk));
	jdff dff_B_8q75BwXS0_1(.din(w_dff_B_txQzqDiA3_1),.dout(w_dff_B_8q75BwXS0_1),.clk(gclk));
	jdff dff_A_0YSAPy1G7_1(.dout(w_n428_0[1]),.din(w_dff_A_0YSAPy1G7_1),.clk(gclk));
	jdff dff_B_YFQvHGfJ1_0(.din(n1493),.dout(w_dff_B_YFQvHGfJ1_0),.clk(gclk));
	jdff dff_A_p0Cf2Y2O2_0(.dout(w_G361_1[0]),.din(w_dff_A_p0Cf2Y2O2_0),.clk(gclk));
	jdff dff_B_0IfXNE3G0_1(.din(n1485),.dout(w_dff_B_0IfXNE3G0_1),.clk(gclk));
	jdff dff_A_DA9kbywb7_0(.dout(w_n437_0[0]),.din(w_dff_A_DA9kbywb7_0),.clk(gclk));
	jdff dff_B_y3kByK1p7_2(.din(n437),.dout(w_dff_B_y3kByK1p7_2),.clk(gclk));
	jdff dff_A_f0ymMM9S3_0(.dout(w_G503_2[0]),.din(w_dff_A_f0ymMM9S3_0),.clk(gclk));
	jdff dff_A_OmWq2bZc5_0(.dout(w_dff_A_f0ymMM9S3_0),.din(w_dff_A_OmWq2bZc5_0),.clk(gclk));
	jdff dff_A_TVETGGw30_0(.dout(w_dff_A_OmWq2bZc5_0),.din(w_dff_A_TVETGGw30_0),.clk(gclk));
	jdff dff_B_1sRfBGLA1_1(.din(n1481),.dout(w_dff_B_1sRfBGLA1_1),.clk(gclk));
	jdff dff_B_9RVLNSpN3_1(.din(n1471),.dout(w_dff_B_9RVLNSpN3_1),.clk(gclk));
	jdff dff_B_SbN4iOHA4_1(.din(w_dff_B_9RVLNSpN3_1),.dout(w_dff_B_SbN4iOHA4_1),.clk(gclk));
	jdff dff_A_m2qxj6TM4_1(.dout(w_G341_2[1]),.din(w_dff_A_m2qxj6TM4_1),.clk(gclk));
	jdff dff_B_WoUeSEXS3_1(.din(n1462),.dout(w_dff_B_WoUeSEXS3_1),.clk(gclk));
	jdff dff_B_qaJGMqE42_1(.din(w_dff_B_WoUeSEXS3_1),.dout(w_dff_B_qaJGMqE42_1),.clk(gclk));
	jdff dff_A_eRUhx5PH6_1(.dout(w_G351_2[1]),.din(w_dff_A_eRUhx5PH6_1),.clk(gclk));
	jdff dff_B_Z90rQbll4_1(.din(n1453),.dout(w_dff_B_Z90rQbll4_1),.clk(gclk));
	jdff dff_A_MS4Ctbw94_0(.dout(w_n749_5[0]),.din(w_dff_A_MS4Ctbw94_0),.clk(gclk));
	jdff dff_A_wgdFmCoQ5_0(.dout(w_dff_A_MS4Ctbw94_0),.din(w_dff_A_wgdFmCoQ5_0),.clk(gclk));
	jdff dff_A_QST1B0gp0_0(.dout(w_dff_A_wgdFmCoQ5_0),.din(w_dff_A_QST1B0gp0_0),.clk(gclk));
	jdff dff_A_ADhn6bIm6_1(.dout(w_n749_5[1]),.din(w_dff_A_ADhn6bIm6_1),.clk(gclk));
	jdff dff_A_SEGSm8Ks1_1(.dout(w_dff_A_ADhn6bIm6_1),.din(w_dff_A_SEGSm8Ks1_1),.clk(gclk));
	jdff dff_A_nvpZD04T0_1(.dout(w_dff_A_SEGSm8Ks1_1),.din(w_dff_A_nvpZD04T0_1),.clk(gclk));
	jdff dff_A_qGz84Lul3_1(.dout(w_dff_A_nvpZD04T0_1),.din(w_dff_A_qGz84Lul3_1),.clk(gclk));
	jdff dff_A_lB6CdXag1_1(.dout(w_dff_A_qGz84Lul3_1),.din(w_dff_A_lB6CdXag1_1),.clk(gclk));
	jdff dff_A_yiuihqQH1_1(.dout(w_dff_A_lB6CdXag1_1),.din(w_dff_A_yiuihqQH1_1),.clk(gclk));
	jdff dff_A_1nueY5bw9_1(.dout(w_dff_A_yiuihqQH1_1),.din(w_dff_A_1nueY5bw9_1),.clk(gclk));
	jdff dff_A_ElibNCo56_1(.dout(w_dff_A_1nueY5bw9_1),.din(w_dff_A_ElibNCo56_1),.clk(gclk));
	jdff dff_A_cqpGSbFZ2_1(.dout(w_dff_A_ElibNCo56_1),.din(w_dff_A_cqpGSbFZ2_1),.clk(gclk));
	jdff dff_A_vsuBuerG9_1(.dout(w_dff_A_cqpGSbFZ2_1),.din(w_dff_A_vsuBuerG9_1),.clk(gclk));
	jdff dff_A_bzz8OX603_1(.dout(w_dff_A_vsuBuerG9_1),.din(w_dff_A_bzz8OX603_1),.clk(gclk));
	jdff dff_A_KAFfH4199_1(.dout(w_dff_A_bzz8OX603_1),.din(w_dff_A_KAFfH4199_1),.clk(gclk));
	jdff dff_B_070zhp4a5_0(.din(n1452),.dout(w_dff_B_070zhp4a5_0),.clk(gclk));
	jdff dff_A_g6zkyckM7_0(.dout(w_n1451_0[0]),.din(w_dff_A_g6zkyckM7_0),.clk(gclk));
	jdff dff_A_JILC84RG8_0(.dout(w_dff_A_g6zkyckM7_0),.din(w_dff_A_JILC84RG8_0),.clk(gclk));
	jdff dff_B_BRhfia9R7_0(.din(n1450),.dout(w_dff_B_BRhfia9R7_0),.clk(gclk));
	jdff dff_B_HxMFxo4U0_0(.din(w_dff_B_BRhfia9R7_0),.dout(w_dff_B_HxMFxo4U0_0),.clk(gclk));
	jdff dff_B_fxt2xFq75_0(.din(w_dff_B_HxMFxo4U0_0),.dout(w_dff_B_fxt2xFq75_0),.clk(gclk));
	jdff dff_B_tDfNTOYk1_1(.din(n1448),.dout(w_dff_B_tDfNTOYk1_1),.clk(gclk));
	jdff dff_B_D9qgm0eL3_1(.din(w_dff_B_tDfNTOYk1_1),.dout(w_dff_B_D9qgm0eL3_1),.clk(gclk));
	jdff dff_B_M3EazxG68_1(.din(w_dff_B_D9qgm0eL3_1),.dout(w_dff_B_M3EazxG68_1),.clk(gclk));
	jdff dff_A_wjNFHBWa5_0(.dout(w_n763_0[0]),.din(w_dff_A_wjNFHBWa5_0),.clk(gclk));
	jdff dff_A_wYgEsu1j2_0(.dout(w_dff_A_wjNFHBWa5_0),.din(w_dff_A_wYgEsu1j2_0),.clk(gclk));
	jdff dff_A_fqt9ow0n4_0(.dout(w_dff_A_wYgEsu1j2_0),.din(w_dff_A_fqt9ow0n4_0),.clk(gclk));
	jdff dff_A_XM2CG33k7_0(.dout(w_dff_A_fqt9ow0n4_0),.din(w_dff_A_XM2CG33k7_0),.clk(gclk));
	jdff dff_A_8b9rerLI4_0(.dout(w_dff_A_XM2CG33k7_0),.din(w_dff_A_8b9rerLI4_0),.clk(gclk));
	jdff dff_A_Jl8lj5A05_0(.dout(w_dff_A_8b9rerLI4_0),.din(w_dff_A_Jl8lj5A05_0),.clk(gclk));
	jdff dff_A_HJuIYKJ17_0(.dout(w_dff_A_Jl8lj5A05_0),.din(w_dff_A_HJuIYKJ17_0),.clk(gclk));
	jdff dff_A_7vTZhl8j5_0(.dout(w_dff_A_HJuIYKJ17_0),.din(w_dff_A_7vTZhl8j5_0),.clk(gclk));
	jdff dff_B_hdAH0NYh6_1(.din(n1439),.dout(w_dff_B_hdAH0NYh6_1),.clk(gclk));
	jdff dff_B_jTV28bEn7_1(.din(n1441),.dout(w_dff_B_jTV28bEn7_1),.clk(gclk));
	jdff dff_B_4gd9p14e0_0(.din(n1437),.dout(w_dff_B_4gd9p14e0_0),.clk(gclk));
	jdff dff_B_rwnme35b7_0(.din(n1436),.dout(w_dff_B_rwnme35b7_0),.clk(gclk));
	jdff dff_A_IjCUvMks7_0(.dout(w_n1429_0[0]),.din(w_dff_A_IjCUvMks7_0),.clk(gclk));
	jdff dff_B_sbTVpKbU0_1(.din(n1427),.dout(w_dff_B_sbTVpKbU0_1),.clk(gclk));
	jdff dff_A_4tqWAQzS3_2(.dout(w_n641_0[2]),.din(w_dff_A_4tqWAQzS3_2),.clk(gclk));
	jdff dff_A_9PX4pKkY6_2(.dout(w_dff_A_4tqWAQzS3_2),.din(w_dff_A_9PX4pKkY6_2),.clk(gclk));
	jdff dff_A_9EDswMRN3_0(.dout(w_n640_0[0]),.din(w_dff_A_9EDswMRN3_0),.clk(gclk));
	jdff dff_A_GGPnnmZ95_0(.dout(w_n639_0[0]),.din(w_dff_A_GGPnnmZ95_0),.clk(gclk));
	jdff dff_A_MvABrmes5_0(.dout(w_n624_0[0]),.din(w_dff_A_MvABrmes5_0),.clk(gclk));
	jdff dff_A_GvO4Rd130_0(.dout(w_dff_A_MvABrmes5_0),.din(w_dff_A_GvO4Rd130_0),.clk(gclk));
	jdff dff_A_SNNFvQ9E1_1(.dout(w_n624_0[1]),.din(w_dff_A_SNNFvQ9E1_1),.clk(gclk));
	jdff dff_B_BzB1UFcY7_3(.din(n624),.dout(w_dff_B_BzB1UFcY7_3),.clk(gclk));
	jdff dff_B_NvEx2L4N1_3(.din(w_dff_B_BzB1UFcY7_3),.dout(w_dff_B_NvEx2L4N1_3),.clk(gclk));
	jdff dff_A_OsoWLGTJ2_1(.dout(w_n620_1[1]),.din(w_dff_A_OsoWLGTJ2_1),.clk(gclk));
	jdff dff_A_WiJ4haWB9_1(.dout(w_dff_A_OsoWLGTJ2_1),.din(w_dff_A_WiJ4haWB9_1),.clk(gclk));
	jdff dff_A_S2ZyZwVv3_1(.dout(w_dff_A_WiJ4haWB9_1),.din(w_dff_A_S2ZyZwVv3_1),.clk(gclk));
	jdff dff_A_QwkIgFgX5_1(.dout(w_dff_A_S2ZyZwVv3_1),.din(w_dff_A_QwkIgFgX5_1),.clk(gclk));
	jdff dff_A_DIC2YVHE3_1(.dout(w_n620_0[1]),.din(w_dff_A_DIC2YVHE3_1),.clk(gclk));
	jdff dff_A_nyTJjvBJ0_1(.dout(w_dff_A_DIC2YVHE3_1),.din(w_dff_A_nyTJjvBJ0_1),.clk(gclk));
	jdff dff_A_mg2hnIcf4_2(.dout(w_n620_0[2]),.din(w_dff_A_mg2hnIcf4_2),.clk(gclk));
	jdff dff_A_8N7A6szk1_2(.dout(w_dff_A_mg2hnIcf4_2),.din(w_dff_A_8N7A6szk1_2),.clk(gclk));
	jdff dff_A_JMEe3V9P9_2(.dout(w_dff_A_8N7A6szk1_2),.din(w_dff_A_JMEe3V9P9_2),.clk(gclk));
	jdff dff_A_19B2iTki8_2(.dout(w_dff_A_JMEe3V9P9_2),.din(w_dff_A_19B2iTki8_2),.clk(gclk));
	jdff dff_A_BnrnhBTY2_2(.dout(w_dff_A_19B2iTki8_2),.din(w_dff_A_BnrnhBTY2_2),.clk(gclk));
	jdff dff_A_IoQihe982_2(.dout(w_dff_A_BnrnhBTY2_2),.din(w_dff_A_IoQihe982_2),.clk(gclk));
	jdff dff_A_XgKPFoq79_2(.dout(w_dff_A_IoQihe982_2),.din(w_dff_A_XgKPFoq79_2),.clk(gclk));
	jdff dff_A_L66qirOK6_1(.dout(w_n618_0[1]),.din(w_dff_A_L66qirOK6_1),.clk(gclk));
	jdff dff_A_rDB1eUaj8_1(.dout(w_dff_A_L66qirOK6_1),.din(w_dff_A_rDB1eUaj8_1),.clk(gclk));
	jdff dff_A_HDCz66Ce9_1(.dout(w_dff_A_rDB1eUaj8_1),.din(w_dff_A_HDCz66Ce9_1),.clk(gclk));
	jdff dff_A_rGUqccYP3_1(.dout(w_dff_A_HDCz66Ce9_1),.din(w_dff_A_rGUqccYP3_1),.clk(gclk));
	jdff dff_A_TgplJfUF8_1(.dout(w_dff_A_rGUqccYP3_1),.din(w_dff_A_TgplJfUF8_1),.clk(gclk));
	jdff dff_A_hqzwr1cJ4_1(.dout(w_dff_A_TgplJfUF8_1),.din(w_dff_A_hqzwr1cJ4_1),.clk(gclk));
	jdff dff_A_67VDDRXs8_2(.dout(w_n618_0[2]),.din(w_dff_A_67VDDRXs8_2),.clk(gclk));
	jdff dff_A_pq0OAUj88_2(.dout(w_dff_A_67VDDRXs8_2),.din(w_dff_A_pq0OAUj88_2),.clk(gclk));
	jdff dff_A_xWm5OZUZ6_2(.dout(w_dff_A_pq0OAUj88_2),.din(w_dff_A_xWm5OZUZ6_2),.clk(gclk));
	jdff dff_A_Sed29K6s0_0(.dout(w_n1425_0[0]),.din(w_dff_A_Sed29K6s0_0),.clk(gclk));
	jdff dff_B_V7dT85qn1_1(.din(n1411),.dout(w_dff_B_V7dT85qn1_1),.clk(gclk));
	jdff dff_A_qLkJq7Yp4_0(.dout(w_n1422_0[0]),.din(w_dff_A_qLkJq7Yp4_0),.clk(gclk));
	jdff dff_B_83fBB4Zg2_1(.din(n1418),.dout(w_dff_B_83fBB4Zg2_1),.clk(gclk));
	jdff dff_B_IwYH0tVS1_1(.din(w_dff_B_83fBB4Zg2_1),.dout(w_dff_B_IwYH0tVS1_1),.clk(gclk));
	jdff dff_B_74lelJ1H2_1(.din(w_dff_B_IwYH0tVS1_1),.dout(w_dff_B_74lelJ1H2_1),.clk(gclk));
	jdff dff_B_aViG2jUQ5_1(.din(n1419),.dout(w_dff_B_aViG2jUQ5_1),.clk(gclk));
	jdff dff_B_LvAdtN1b5_1(.din(w_dff_B_aViG2jUQ5_1),.dout(w_dff_B_LvAdtN1b5_1),.clk(gclk));
	jdff dff_A_i8yyIplH2_2(.dout(w_n660_0[2]),.din(w_dff_A_i8yyIplH2_2),.clk(gclk));
	jdff dff_A_l5PaLoW59_2(.dout(w_dff_A_i8yyIplH2_2),.din(w_dff_A_l5PaLoW59_2),.clk(gclk));
	jdff dff_A_AJqdgG8U3_2(.dout(w_dff_A_l5PaLoW59_2),.din(w_dff_A_AJqdgG8U3_2),.clk(gclk));
	jdff dff_A_IuChjonL2_2(.dout(w_dff_A_AJqdgG8U3_2),.din(w_dff_A_IuChjonL2_2),.clk(gclk));
	jdff dff_A_uAsOX6ck7_2(.dout(w_dff_A_IuChjonL2_2),.din(w_dff_A_uAsOX6ck7_2),.clk(gclk));
	jdff dff_A_TEyNCykl0_2(.dout(w_dff_A_uAsOX6ck7_2),.din(w_dff_A_TEyNCykl0_2),.clk(gclk));
	jdff dff_A_QATLQh7l7_2(.dout(w_n792_0[2]),.din(w_dff_A_QATLQh7l7_2),.clk(gclk));
	jdff dff_A_duxUuruZ6_2(.dout(w_dff_A_QATLQh7l7_2),.din(w_dff_A_duxUuruZ6_2),.clk(gclk));
	jdff dff_A_QjmHfwz06_2(.dout(w_dff_A_duxUuruZ6_2),.din(w_dff_A_QjmHfwz06_2),.clk(gclk));
	jdff dff_A_p6tyzjNY2_2(.dout(w_dff_A_QjmHfwz06_2),.din(w_dff_A_p6tyzjNY2_2),.clk(gclk));
	jdff dff_A_ykCrhBdZ7_2(.dout(w_dff_A_p6tyzjNY2_2),.din(w_dff_A_ykCrhBdZ7_2),.clk(gclk));
	jdff dff_A_zPf5536V2_2(.dout(w_dff_A_ykCrhBdZ7_2),.din(w_dff_A_zPf5536V2_2),.clk(gclk));
	jdff dff_A_5ZcRhB5p2_2(.dout(w_dff_A_zPf5536V2_2),.din(w_dff_A_5ZcRhB5p2_2),.clk(gclk));
	jdff dff_A_5SDxX0FA8_2(.dout(w_dff_A_5ZcRhB5p2_2),.din(w_dff_A_5SDxX0FA8_2),.clk(gclk));
	jdff dff_A_eBOdeqzC9_2(.dout(w_dff_A_5SDxX0FA8_2),.din(w_dff_A_eBOdeqzC9_2),.clk(gclk));
	jdff dff_A_rLHjHBM64_1(.dout(w_n790_0[1]),.din(w_dff_A_rLHjHBM64_1),.clk(gclk));
	jdff dff_A_DT2oUB298_1(.dout(w_dff_A_rLHjHBM64_1),.din(w_dff_A_DT2oUB298_1),.clk(gclk));
	jdff dff_A_Uym4fpnO9_1(.dout(w_dff_A_DT2oUB298_1),.din(w_dff_A_Uym4fpnO9_1),.clk(gclk));
	jdff dff_A_vTp8Jlp28_1(.dout(w_dff_A_Uym4fpnO9_1),.din(w_dff_A_vTp8Jlp28_1),.clk(gclk));
	jdff dff_A_lux5fZqY1_1(.dout(w_dff_A_vTp8Jlp28_1),.din(w_dff_A_lux5fZqY1_1),.clk(gclk));
	jdff dff_A_WKhuoL1k8_1(.dout(w_dff_A_lux5fZqY1_1),.din(w_dff_A_WKhuoL1k8_1),.clk(gclk));
	jdff dff_A_pAbX9eVw6_1(.dout(w_dff_A_WKhuoL1k8_1),.din(w_dff_A_pAbX9eVw6_1),.clk(gclk));
	jdff dff_A_NKvMMmvi2_1(.dout(w_dff_A_pAbX9eVw6_1),.din(w_dff_A_NKvMMmvi2_1),.clk(gclk));
	jdff dff_A_WPiyapb80_1(.dout(w_dff_A_NKvMMmvi2_1),.din(w_dff_A_WPiyapb80_1),.clk(gclk));
	jdff dff_A_5Cx11GKH9_1(.dout(w_dff_A_WPiyapb80_1),.din(w_dff_A_5Cx11GKH9_1),.clk(gclk));
	jdff dff_B_kj2qjmgO0_1(.din(n1413),.dout(w_dff_B_kj2qjmgO0_1),.clk(gclk));
	jdff dff_B_B8tKFCJD3_1(.din(w_dff_B_kj2qjmgO0_1),.dout(w_dff_B_B8tKFCJD3_1),.clk(gclk));
	jdff dff_B_K3LAVPUE1_1(.din(w_dff_B_B8tKFCJD3_1),.dout(w_dff_B_K3LAVPUE1_1),.clk(gclk));
	jdff dff_B_6fn1E8pr1_1(.din(w_dff_B_K3LAVPUE1_1),.dout(w_dff_B_6fn1E8pr1_1),.clk(gclk));
	jdff dff_B_iqouE5Dq1_1(.din(n1414),.dout(w_dff_B_iqouE5Dq1_1),.clk(gclk));
	jdff dff_B_mtGOdMAp0_1(.din(w_dff_B_iqouE5Dq1_1),.dout(w_dff_B_mtGOdMAp0_1),.clk(gclk));
	jdff dff_B_R8tE4bJQ6_1(.din(w_dff_B_mtGOdMAp0_1),.dout(w_dff_B_R8tE4bJQ6_1),.clk(gclk));
	jdff dff_A_GKaXrJW94_1(.dout(w_n821_0[1]),.din(w_dff_A_GKaXrJW94_1),.clk(gclk));
	jdff dff_B_iPyaFyLN4_1(.din(n812),.dout(w_dff_B_iPyaFyLN4_1),.clk(gclk));
	jdff dff_B_QKPsNrL36_1(.din(w_dff_B_iPyaFyLN4_1),.dout(w_dff_B_QKPsNrL36_1),.clk(gclk));
	jdff dff_B_4MwrLTNz6_1(.din(w_dff_B_QKPsNrL36_1),.dout(w_dff_B_4MwrLTNz6_1),.clk(gclk));
	jdff dff_B_CS9FX0KI7_1(.din(w_dff_B_4MwrLTNz6_1),.dout(w_dff_B_CS9FX0KI7_1),.clk(gclk));
	jdff dff_B_HosoUUz22_1(.din(n813),.dout(w_dff_B_HosoUUz22_1),.clk(gclk));
	jdff dff_B_sAmJnBz90_1(.din(w_dff_B_HosoUUz22_1),.dout(w_dff_B_sAmJnBz90_1),.clk(gclk));
	jdff dff_B_pKbLoEhn9_1(.din(w_dff_B_sAmJnBz90_1),.dout(w_dff_B_pKbLoEhn9_1),.clk(gclk));
	jdff dff_A_K5I8OpjW7_1(.dout(w_n819_0[1]),.din(w_dff_A_K5I8OpjW7_1),.clk(gclk));
	jdff dff_A_ECOYXRRD5_1(.dout(w_dff_A_K5I8OpjW7_1),.din(w_dff_A_ECOYXRRD5_1),.clk(gclk));
	jdff dff_A_wTccKRfM2_0(.dout(w_n377_1[0]),.din(w_dff_A_wTccKRfM2_0),.clk(gclk));
	jdff dff_A_jpK1YSoA7_0(.dout(w_n814_0[0]),.din(w_dff_A_jpK1YSoA7_0),.clk(gclk));
	jdff dff_A_Of2A13lG7_0(.dout(w_dff_A_jpK1YSoA7_0),.din(w_dff_A_Of2A13lG7_0),.clk(gclk));
	jdff dff_A_Ox40Ompz4_0(.dout(w_dff_A_Of2A13lG7_0),.din(w_dff_A_Ox40Ompz4_0),.clk(gclk));
	jdff dff_A_MpFtsz1i4_1(.dout(w_n814_0[1]),.din(w_dff_A_MpFtsz1i4_1),.clk(gclk));
	jdff dff_A_eJs5oGEJ3_1(.dout(w_dff_A_MpFtsz1i4_1),.din(w_dff_A_eJs5oGEJ3_1),.clk(gclk));
	jdff dff_A_tfjwpnlU9_2(.dout(w_n377_0[2]),.din(w_dff_A_tfjwpnlU9_2),.clk(gclk));
	jdff dff_B_wOVfCONj9_3(.din(n377),.dout(w_dff_B_wOVfCONj9_3),.clk(gclk));
	jdff dff_A_aMYZnVF50_0(.dout(w_G534_2[0]),.din(w_dff_A_aMYZnVF50_0),.clk(gclk));
	jdff dff_A_riodS2C01_0(.dout(w_dff_A_aMYZnVF50_0),.din(w_dff_A_riodS2C01_0),.clk(gclk));
	jdff dff_A_KpExEhaJ8_0(.dout(w_dff_A_riodS2C01_0),.din(w_dff_A_KpExEhaJ8_0),.clk(gclk));
	jdff dff_A_r33rlOjW2_1(.dout(w_n1412_0[1]),.din(w_dff_A_r33rlOjW2_1),.clk(gclk));
	jdff dff_A_gNshOweR9_1(.dout(w_dff_A_r33rlOjW2_1),.din(w_dff_A_gNshOweR9_1),.clk(gclk));
	jdff dff_A_Tc8l7UPY8_2(.dout(w_n1412_0[2]),.din(w_dff_A_Tc8l7UPY8_2),.clk(gclk));
	jdff dff_B_4WThtRxK6_3(.din(n1412),.dout(w_dff_B_4WThtRxK6_3),.clk(gclk));
	jdff dff_B_juz86tgt3_3(.din(w_dff_B_4WThtRxK6_3),.dout(w_dff_B_juz86tgt3_3),.clk(gclk));
	jdff dff_B_FKRt0SOf7_3(.din(w_dff_B_juz86tgt3_3),.dout(w_dff_B_FKRt0SOf7_3),.clk(gclk));
	jdff dff_B_PeEuHqG89_3(.din(w_dff_B_FKRt0SOf7_3),.dout(w_dff_B_PeEuHqG89_3),.clk(gclk));
	jdff dff_B_N1UjULZ72_3(.din(w_dff_B_PeEuHqG89_3),.dout(w_dff_B_N1UjULZ72_3),.clk(gclk));
	jdff dff_B_X3lsKBLN1_3(.din(w_dff_B_N1UjULZ72_3),.dout(w_dff_B_X3lsKBLN1_3),.clk(gclk));
	jdff dff_B_cAwO6GxZ7_3(.din(w_dff_B_X3lsKBLN1_3),.dout(w_dff_B_cAwO6GxZ7_3),.clk(gclk));
	jdff dff_B_gba4Efgt3_3(.din(w_dff_B_cAwO6GxZ7_3),.dout(w_dff_B_gba4Efgt3_3),.clk(gclk));
	jdff dff_B_4AEnmj8c3_3(.din(w_dff_B_gba4Efgt3_3),.dout(w_dff_B_4AEnmj8c3_3),.clk(gclk));
	jdff dff_B_t59Osa8H5_3(.din(w_dff_B_4AEnmj8c3_3),.dout(w_dff_B_t59Osa8H5_3),.clk(gclk));
	jdff dff_A_v18HLLcD7_0(.dout(w_G2174_0[0]),.din(w_dff_A_v18HLLcD7_0),.clk(gclk));
	jdff dff_A_tn4be7sx9_0(.dout(w_dff_A_v18HLLcD7_0),.din(w_dff_A_tn4be7sx9_0),.clk(gclk));
	jdff dff_A_WOCXykHj5_0(.dout(w_dff_A_tn4be7sx9_0),.din(w_dff_A_WOCXykHj5_0),.clk(gclk));
	jdff dff_A_Vfot0y3l7_0(.dout(w_dff_A_WOCXykHj5_0),.din(w_dff_A_Vfot0y3l7_0),.clk(gclk));
	jdff dff_A_Qt41nr4G6_0(.dout(w_dff_A_Vfot0y3l7_0),.din(w_dff_A_Qt41nr4G6_0),.clk(gclk));
	jdff dff_A_ASigP1092_0(.dout(w_dff_A_Qt41nr4G6_0),.din(w_dff_A_ASigP1092_0),.clk(gclk));
	jdff dff_A_8tMn8B7I1_0(.dout(w_dff_A_ASigP1092_0),.din(w_dff_A_8tMn8B7I1_0),.clk(gclk));
	jdff dff_A_Gs9GXNQm0_0(.dout(w_dff_A_8tMn8B7I1_0),.din(w_dff_A_Gs9GXNQm0_0),.clk(gclk));
	jdff dff_A_mzUlbWye1_0(.dout(w_dff_A_Gs9GXNQm0_0),.din(w_dff_A_mzUlbWye1_0),.clk(gclk));
	jdff dff_A_huMMXZVe7_0(.dout(w_dff_A_mzUlbWye1_0),.din(w_dff_A_huMMXZVe7_0),.clk(gclk));
	jdff dff_A_cNHhFBwc5_0(.dout(w_dff_A_huMMXZVe7_0),.din(w_dff_A_cNHhFBwc5_0),.clk(gclk));
	jdff dff_A_gkfOwU5h4_0(.dout(w_dff_A_cNHhFBwc5_0),.din(w_dff_A_gkfOwU5h4_0),.clk(gclk));
	jdff dff_A_m2APYiOi5_0(.dout(w_dff_A_gkfOwU5h4_0),.din(w_dff_A_m2APYiOi5_0),.clk(gclk));
	jdff dff_A_NGijUakd5_1(.dout(w_G2174_0[1]),.din(w_dff_A_NGijUakd5_1),.clk(gclk));
	jdff dff_A_MsgonRno8_1(.dout(w_dff_A_NGijUakd5_1),.din(w_dff_A_MsgonRno8_1),.clk(gclk));
	jdff dff_A_7gjxmdrv2_1(.dout(w_dff_A_MsgonRno8_1),.din(w_dff_A_7gjxmdrv2_1),.clk(gclk));
	jdff dff_A_iY2PWA2A5_1(.dout(w_dff_A_7gjxmdrv2_1),.din(w_dff_A_iY2PWA2A5_1),.clk(gclk));
	jdff dff_A_AUIfTuPs6_1(.dout(w_dff_A_iY2PWA2A5_1),.din(w_dff_A_AUIfTuPs6_1),.clk(gclk));
	jdff dff_A_jpX9c8Ra3_1(.dout(w_dff_A_AUIfTuPs6_1),.din(w_dff_A_jpX9c8Ra3_1),.clk(gclk));
	jdff dff_A_dJaWcyFF0_1(.dout(w_dff_A_jpX9c8Ra3_1),.din(w_dff_A_dJaWcyFF0_1),.clk(gclk));
	jdff dff_A_hUETWxeJ4_1(.dout(w_dff_A_dJaWcyFF0_1),.din(w_dff_A_hUETWxeJ4_1),.clk(gclk));
	jdff dff_A_129ujZau1_1(.dout(w_dff_A_hUETWxeJ4_1),.din(w_dff_A_129ujZau1_1),.clk(gclk));
	jdff dff_A_aQ2sne377_1(.dout(w_dff_A_129ujZau1_1),.din(w_dff_A_aQ2sne377_1),.clk(gclk));
	jdff dff_A_ezJhyCPW8_0(.dout(w_n1410_0[0]),.din(w_dff_A_ezJhyCPW8_0),.clk(gclk));
	jdff dff_B_tSgEasV35_0(.din(n1409),.dout(w_dff_B_tSgEasV35_0),.clk(gclk));
	jdff dff_B_unjhe5ER1_0(.din(w_dff_B_tSgEasV35_0),.dout(w_dff_B_unjhe5ER1_0),.clk(gclk));
	jdff dff_A_bkw6TpWq6_0(.dout(w_n401_0[0]),.din(w_dff_A_bkw6TpWq6_0),.clk(gclk));
	jdff dff_A_PY9Lnkmo7_0(.dout(w_dff_A_bkw6TpWq6_0),.din(w_dff_A_PY9Lnkmo7_0),.clk(gclk));
	jdff dff_A_s8jJaLwc5_0(.dout(w_dff_A_PY9Lnkmo7_0),.din(w_dff_A_s8jJaLwc5_0),.clk(gclk));
	jdff dff_B_XuwBpfWG4_2(.din(n401),.dout(w_dff_B_XuwBpfWG4_2),.clk(gclk));
	jdff dff_A_ZC2btJ5m2_0(.dout(w_G490_1[0]),.din(w_dff_A_ZC2btJ5m2_0),.clk(gclk));
	jdff dff_A_H2HNYnEs5_0(.dout(w_dff_A_ZC2btJ5m2_0),.din(w_dff_A_H2HNYnEs5_0),.clk(gclk));
	jdff dff_A_FUOC17pp8_0(.dout(w_dff_A_H2HNYnEs5_0),.din(w_dff_A_FUOC17pp8_0),.clk(gclk));
	jdff dff_A_cYMiPkUq1_1(.dout(w_n654_1[1]),.din(w_dff_A_cYMiPkUq1_1),.clk(gclk));
	jdff dff_A_vUuGiq4C9_1(.dout(w_dff_A_cYMiPkUq1_1),.din(w_dff_A_vUuGiq4C9_1),.clk(gclk));
	jdff dff_A_4eyTO76A5_1(.dout(w_dff_A_vUuGiq4C9_1),.din(w_dff_A_4eyTO76A5_1),.clk(gclk));
	jdff dff_A_U3aJIZ4Z3_1(.dout(w_dff_A_4eyTO76A5_1),.din(w_dff_A_U3aJIZ4Z3_1),.clk(gclk));
	jdff dff_A_MMWmBxtS2_1(.dout(w_dff_A_U3aJIZ4Z3_1),.din(w_dff_A_MMWmBxtS2_1),.clk(gclk));
	jdff dff_A_W2piALF04_1(.dout(w_dff_A_MMWmBxtS2_1),.din(w_dff_A_W2piALF04_1),.clk(gclk));
	jdff dff_A_jYrslpcA9_1(.dout(w_dff_A_W2piALF04_1),.din(w_dff_A_jYrslpcA9_1),.clk(gclk));
	jdff dff_A_5GJOdGyi0_1(.dout(w_dff_A_jYrslpcA9_1),.din(w_dff_A_5GJOdGyi0_1),.clk(gclk));
	jdff dff_A_pX4P1kdQ5_0(.dout(w_n644_0[0]),.din(w_dff_A_pX4P1kdQ5_0),.clk(gclk));
	jdff dff_A_feSviSIp1_0(.dout(w_dff_A_pX4P1kdQ5_0),.din(w_dff_A_feSviSIp1_0),.clk(gclk));
	jdff dff_A_NlApwIhT5_0(.dout(w_dff_A_feSviSIp1_0),.din(w_dff_A_NlApwIhT5_0),.clk(gclk));
	jdff dff_A_Sc2SMKNB7_0(.dout(w_dff_A_NlApwIhT5_0),.din(w_dff_A_Sc2SMKNB7_0),.clk(gclk));
	jdff dff_A_LBdEB4Xo8_2(.dout(w_n644_0[2]),.din(w_dff_A_LBdEB4Xo8_2),.clk(gclk));
	jdff dff_A_BFxkYivm6_2(.dout(w_dff_A_LBdEB4Xo8_2),.din(w_dff_A_BFxkYivm6_2),.clk(gclk));
	jdff dff_A_kZSg5MXX5_1(.dout(w_G293_0[1]),.din(w_dff_A_kZSg5MXX5_1),.clk(gclk));
	jdff dff_A_S5Gh99jH1_1(.dout(w_n746_0[1]),.din(w_dff_A_S5Gh99jH1_1),.clk(gclk));
	jdff dff_A_5uPZEH5K0_1(.dout(w_dff_A_S5Gh99jH1_1),.din(w_dff_A_5uPZEH5K0_1),.clk(gclk));
	jdff dff_A_kWMIyWPc4_1(.dout(w_dff_A_5uPZEH5K0_1),.din(w_dff_A_kWMIyWPc4_1),.clk(gclk));
	jdff dff_A_h8rFwdzc6_1(.dout(w_dff_A_kWMIyWPc4_1),.din(w_dff_A_h8rFwdzc6_1),.clk(gclk));
	jdff dff_B_XvG3bD4C6_1(.din(n741),.dout(w_dff_B_XvG3bD4C6_1),.clk(gclk));
	jdff dff_B_SfwD23T13_1(.din(w_dff_B_XvG3bD4C6_1),.dout(w_dff_B_SfwD23T13_1),.clk(gclk));
	jdff dff_A_hUotwwMm3_1(.dout(w_n742_0[1]),.din(w_dff_A_hUotwwMm3_1),.clk(gclk));
	jdff dff_A_cAGlh6xh6_1(.dout(w_dff_A_hUotwwMm3_1),.din(w_dff_A_cAGlh6xh6_1),.clk(gclk));
	jdff dff_A_klRu9zIB9_1(.dout(w_dff_A_cAGlh6xh6_1),.din(w_dff_A_klRu9zIB9_1),.clk(gclk));
	jdff dff_A_iGxtas971_1(.dout(w_dff_A_klRu9zIB9_1),.din(w_dff_A_iGxtas971_1),.clk(gclk));
	jdff dff_A_lqvx0U101_1(.dout(w_dff_A_iGxtas971_1),.din(w_dff_A_lqvx0U101_1),.clk(gclk));
	jdff dff_A_aurhMe533_1(.dout(w_dff_A_lqvx0U101_1),.din(w_dff_A_aurhMe533_1),.clk(gclk));
	jdff dff_A_hbkPjEYw5_1(.dout(w_dff_A_aurhMe533_1),.din(w_dff_A_hbkPjEYw5_1),.clk(gclk));
	jdff dff_B_xm9n2cNj2_0(.din(n657),.dout(w_dff_B_xm9n2cNj2_0),.clk(gclk));
	jdff dff_B_ZekPhHNU8_1(.din(G323),.dout(w_dff_B_ZekPhHNU8_1),.clk(gclk));
	jdff dff_A_Sb7QOQec3_2(.dout(w_G316_0[2]),.din(w_dff_A_Sb7QOQec3_2),.clk(gclk));
	jdff dff_A_Vl47BYZt6_1(.dout(w_G490_0[1]),.din(w_dff_A_Vl47BYZt6_1),.clk(gclk));
	jdff dff_A_Uvjf0yqw3_1(.dout(w_dff_A_Vl47BYZt6_1),.din(w_dff_A_Uvjf0yqw3_1),.clk(gclk));
	jdff dff_A_HEZv31Xe4_1(.dout(w_dff_A_Uvjf0yqw3_1),.din(w_dff_A_HEZv31Xe4_1),.clk(gclk));
	jdff dff_A_JWxZI3X23_1(.dout(w_dff_A_HEZv31Xe4_1),.din(w_dff_A_JWxZI3X23_1),.clk(gclk));
	jdff dff_A_CRcdYjRi2_2(.dout(w_G490_0[2]),.din(w_dff_A_CRcdYjRi2_2),.clk(gclk));
	jdff dff_A_aBRlDjTD7_2(.dout(w_dff_A_CRcdYjRi2_2),.din(w_dff_A_aBRlDjTD7_2),.clk(gclk));
	jdff dff_A_JI7m7Q3p0_2(.dout(w_dff_A_aBRlDjTD7_2),.din(w_dff_A_JI7m7Q3p0_2),.clk(gclk));
	jdff dff_A_iD7IMbK61_2(.dout(w_dff_A_JI7m7Q3p0_2),.din(w_dff_A_iD7IMbK61_2),.clk(gclk));
	jdff dff_A_IxvVKXhq0_0(.dout(w_n654_2[0]),.din(w_dff_A_IxvVKXhq0_0),.clk(gclk));
	jdff dff_A_jDb5vWbQ6_0(.dout(w_n654_0[0]),.din(w_dff_A_jDb5vWbQ6_0),.clk(gclk));
	jdff dff_B_5zQTNqNL4_3(.din(n654),.dout(w_dff_B_5zQTNqNL4_3),.clk(gclk));
	jdff dff_A_xK9GoD8d5_0(.dout(w_n653_0[0]),.din(w_dff_A_xK9GoD8d5_0),.clk(gclk));
	jdff dff_B_Q7E4iDB55_1(.din(n651),.dout(w_dff_B_Q7E4iDB55_1),.clk(gclk));
	jdff dff_B_CVVTHKpS5_1(.din(G315),.dout(w_dff_B_CVVTHKpS5_1),.clk(gclk));
	jdff dff_A_4q1hYdfh3_0(.dout(w_n414_0[0]),.din(w_dff_A_4q1hYdfh3_0),.clk(gclk));
	jdff dff_A_PNkC3uu93_0(.dout(w_dff_A_4q1hYdfh3_0),.din(w_dff_A_PNkC3uu93_0),.clk(gclk));
	jdff dff_B_jI44hNRp8_2(.din(n414),.dout(w_dff_B_jI44hNRp8_2),.clk(gclk));
	jdff dff_A_buhOiGsc8_0(.dout(w_G479_0[0]),.din(w_dff_A_buhOiGsc8_0),.clk(gclk));
	jdff dff_A_Upu1yvLo5_0(.dout(w_dff_A_buhOiGsc8_0),.din(w_dff_A_Upu1yvLo5_0),.clk(gclk));
	jdff dff_A_zu46DcNC2_0(.dout(w_dff_A_Upu1yvLo5_0),.din(w_dff_A_zu46DcNC2_0),.clk(gclk));
	jdff dff_A_3kBbDxDQ4_1(.dout(w_G479_0[1]),.din(w_dff_A_3kBbDxDQ4_1),.clk(gclk));
	jdff dff_A_qv2urgCy8_1(.dout(w_dff_A_3kBbDxDQ4_1),.din(w_dff_A_qv2urgCy8_1),.clk(gclk));
	jdff dff_A_nmvMlbAs9_1(.dout(w_dff_A_qv2urgCy8_1),.din(w_dff_A_nmvMlbAs9_1),.clk(gclk));
	jdff dff_A_PaFgiKnh5_1(.dout(w_n648_0[1]),.din(w_dff_A_PaFgiKnh5_1),.clk(gclk));
	jdff dff_A_KT1GeWuA7_1(.dout(w_dff_A_PaFgiKnh5_1),.din(w_dff_A_KT1GeWuA7_1),.clk(gclk));
	jdff dff_A_0i8wc61A6_1(.dout(w_dff_A_KT1GeWuA7_1),.din(w_dff_A_0i8wc61A6_1),.clk(gclk));
	jdff dff_A_2q2vU2484_1(.dout(w_dff_A_0i8wc61A6_1),.din(w_dff_A_2q2vU2484_1),.clk(gclk));
	jdff dff_A_GroD6Vqu4_2(.dout(w_n648_0[2]),.din(w_dff_A_GroD6Vqu4_2),.clk(gclk));
	jdff dff_A_Bf3qpHA62_2(.dout(w_dff_A_GroD6Vqu4_2),.din(w_dff_A_Bf3qpHA62_2),.clk(gclk));
	jdff dff_A_NW2y806O4_2(.dout(w_dff_A_Bf3qpHA62_2),.din(w_dff_A_NW2y806O4_2),.clk(gclk));
	jdff dff_A_jokAWxaH0_2(.dout(w_dff_A_NW2y806O4_2),.din(w_dff_A_jokAWxaH0_2),.clk(gclk));
	jdff dff_A_q27zPIaQ0_2(.dout(w_dff_A_jokAWxaH0_2),.din(w_dff_A_q27zPIaQ0_2),.clk(gclk));
	jdff dff_B_eEc63flA4_0(.din(n647),.dout(w_dff_B_eEc63flA4_0),.clk(gclk));
	jdff dff_B_iK4y7oQM2_1(.din(G307),.dout(w_dff_B_iK4y7oQM2_1),.clk(gclk));
	jdff dff_A_eWQJRtlK4_0(.dout(w_G302_0[0]),.din(w_dff_A_eWQJRtlK4_0),.clk(gclk));
	jdff dff_A_6kitU1zB8_1(.dout(w_G302_0[1]),.din(w_dff_A_6kitU1zB8_1),.clk(gclk));
	jdff dff_B_dUa0MRE69_1(.din(n727),.dout(w_dff_B_dUa0MRE69_1),.clk(gclk));
	jdff dff_A_1j4RLxNY6_0(.dout(w_n635_1[0]),.din(w_dff_A_1j4RLxNY6_0),.clk(gclk));
	jdff dff_A_OfTuXaEp5_1(.dout(w_n635_0[1]),.din(w_dff_A_OfTuXaEp5_1),.clk(gclk));
	jdff dff_A_8ywYSxFS9_1(.dout(w_dff_A_OfTuXaEp5_1),.din(w_dff_A_8ywYSxFS9_1),.clk(gclk));
	jdff dff_B_SfR3MZBx3_1(.din(n633),.dout(w_dff_B_SfR3MZBx3_1),.clk(gclk));
	jdff dff_A_Foq3VPLQ3_0(.dout(w_G366_0[0]),.din(w_dff_A_Foq3VPLQ3_0),.clk(gclk));
	jdff dff_A_JKLtRAxP4_0(.dout(w_G332_2[0]),.din(w_dff_A_JKLtRAxP4_0),.clk(gclk));
	jdff dff_A_Fq3Yi8Dz9_2(.dout(w_G332_2[2]),.din(w_dff_A_Fq3Yi8Dz9_2),.clk(gclk));
	jdff dff_A_eb1XlFli1_0(.dout(w_n628_0[0]),.din(w_dff_A_eb1XlFli1_0),.clk(gclk));
	jdff dff_A_nvhxGLEV3_0(.dout(w_dff_A_eb1XlFli1_0),.din(w_dff_A_nvhxGLEV3_0),.clk(gclk));
	jdff dff_A_L5VotdaR3_0(.dout(w_dff_A_nvhxGLEV3_0),.din(w_dff_A_L5VotdaR3_0),.clk(gclk));
	jdff dff_A_NneLSLTL0_2(.dout(w_n628_0[2]),.din(w_dff_A_NneLSLTL0_2),.clk(gclk));
	jdff dff_A_5xH6wiIu1_0(.dout(w_G358_0[0]),.din(w_dff_A_5xH6wiIu1_0),.clk(gclk));
	jdff dff_A_Hpe11eud5_1(.dout(w_n625_0[1]),.din(w_dff_A_Hpe11eud5_1),.clk(gclk));
	jdff dff_A_Tw4If2hQ9_2(.dout(w_G351_0[2]),.din(w_dff_A_Tw4If2hQ9_2),.clk(gclk));
	jdff dff_A_iyld7ep81_0(.dout(w_G534_0[0]),.din(w_dff_A_iyld7ep81_0),.clk(gclk));
	jdff dff_A_p9XJx9lM5_0(.dout(w_dff_A_iyld7ep81_0),.din(w_dff_A_p9XJx9lM5_0),.clk(gclk));
	jdff dff_A_IDL7g5my3_0(.dout(w_dff_A_p9XJx9lM5_0),.din(w_dff_A_IDL7g5my3_0),.clk(gclk));
	jdff dff_A_4v46mBNE5_2(.dout(w_G534_0[2]),.din(w_dff_A_4v46mBNE5_2),.clk(gclk));
	jdff dff_A_pNXeXqfn6_2(.dout(w_dff_A_4v46mBNE5_2),.din(w_dff_A_pNXeXqfn6_2),.clk(gclk));
	jdff dff_A_MOvQLspi1_2(.dout(w_dff_A_pNXeXqfn6_2),.din(w_dff_A_MOvQLspi1_2),.clk(gclk));
	jdff dff_A_tStlNfMY4_0(.dout(w_n726_0[0]),.din(w_dff_A_tStlNfMY4_0),.clk(gclk));
	jdff dff_A_Lpp4XiX75_0(.dout(w_dff_A_tStlNfMY4_0),.din(w_dff_A_Lpp4XiX75_0),.clk(gclk));
	jdff dff_A_hcovNpaa2_0(.dout(w_G348_0[0]),.din(w_dff_A_hcovNpaa2_0),.clk(gclk));
	jdff dff_A_WSnSbauz7_1(.dout(w_G332_1[1]),.din(w_dff_A_WSnSbauz7_1),.clk(gclk));
	jdff dff_A_mbdOxSkR8_1(.dout(w_n621_0[1]),.din(w_dff_A_mbdOxSkR8_1),.clk(gclk));
	jdff dff_A_Sl0epb350_2(.dout(w_G341_0[2]),.din(w_dff_A_Sl0epb350_2),.clk(gclk));
	jdff dff_A_glcBLkLD3_0(.dout(w_n389_1[0]),.din(w_dff_A_glcBLkLD3_0),.clk(gclk));
	jdff dff_A_gkmhSzvi0_2(.dout(w_n389_0[2]),.din(w_dff_A_gkmhSzvi0_2),.clk(gclk));
	jdff dff_B_84Cmest04_3(.din(n389),.dout(w_dff_B_84Cmest04_3),.clk(gclk));
	jdff dff_A_V5DDT1wr1_0(.dout(w_G523_1[0]),.din(w_dff_A_V5DDT1wr1_0),.clk(gclk));
	jdff dff_A_7TYcbolV4_0(.dout(w_dff_A_V5DDT1wr1_0),.din(w_dff_A_7TYcbolV4_0),.clk(gclk));
	jdff dff_A_9mALEgny1_0(.dout(w_dff_A_7TYcbolV4_0),.din(w_dff_A_9mALEgny1_0),.clk(gclk));
	jdff dff_A_1mS2KaGS0_1(.dout(w_G523_1[1]),.din(w_dff_A_1mS2KaGS0_1),.clk(gclk));
	jdff dff_A_9OE3YKL51_1(.dout(w_dff_A_1mS2KaGS0_1),.din(w_dff_A_9OE3YKL51_1),.clk(gclk));
	jdff dff_A_5pSo3KrS6_1(.dout(w_dff_A_9OE3YKL51_1),.din(w_dff_A_5pSo3KrS6_1),.clk(gclk));
	jdff dff_A_USeJePYc5_1(.dout(w_G523_0[1]),.din(w_dff_A_USeJePYc5_1),.clk(gclk));
	jdff dff_A_ihptJDIZ3_1(.dout(w_dff_A_USeJePYc5_1),.din(w_dff_A_ihptJDIZ3_1),.clk(gclk));
	jdff dff_A_Aw05G7vG7_1(.dout(w_dff_A_ihptJDIZ3_1),.din(w_dff_A_Aw05G7vG7_1),.clk(gclk));
	jdff dff_A_IChldhM89_2(.dout(w_G523_0[2]),.din(w_dff_A_IChldhM89_2),.clk(gclk));
	jdff dff_A_LSCJ1cll4_2(.dout(w_dff_A_IChldhM89_2),.din(w_dff_A_LSCJ1cll4_2),.clk(gclk));
	jdff dff_A_3nvPKuqC5_2(.dout(w_dff_A_LSCJ1cll4_2),.din(w_dff_A_3nvPKuqC5_2),.clk(gclk));
	jdff dff_A_pwVsbGq33_1(.dout(w_n722_0[1]),.din(w_dff_A_pwVsbGq33_1),.clk(gclk));
	jdff dff_A_VU6hs2k22_1(.dout(w_dff_A_pwVsbGq33_1),.din(w_dff_A_VU6hs2k22_1),.clk(gclk));
	jdff dff_A_hQzJJwvS2_1(.dout(w_dff_A_VU6hs2k22_1),.din(w_dff_A_hQzJJwvS2_1),.clk(gclk));
	jdff dff_A_ldf0b7vZ9_1(.dout(w_dff_A_hQzJJwvS2_1),.din(w_dff_A_ldf0b7vZ9_1),.clk(gclk));
	jdff dff_A_5hhZrTyZ5_1(.dout(w_n721_0[1]),.din(w_dff_A_5hhZrTyZ5_1),.clk(gclk));
	jdff dff_A_IXDS5e1t1_1(.dout(w_dff_A_5hhZrTyZ5_1),.din(w_dff_A_IXDS5e1t1_1),.clk(gclk));
	jdff dff_A_QJscMUJO4_1(.dout(w_dff_A_IXDS5e1t1_1),.din(w_dff_A_QJscMUJO4_1),.clk(gclk));
	jdff dff_A_7ckStsVJ9_1(.dout(w_dff_A_QJscMUJO4_1),.din(w_dff_A_7ckStsVJ9_1),.clk(gclk));
	jdff dff_A_tDgj3zKQ2_1(.dout(w_dff_A_7ckStsVJ9_1),.din(w_dff_A_tDgj3zKQ2_1),.clk(gclk));
	jdff dff_A_Rw1rXM5c4_1(.dout(w_n619_0[1]),.din(w_dff_A_Rw1rXM5c4_1),.clk(gclk));
	jdff dff_A_xsATXNB53_1(.dout(w_dff_A_Rw1rXM5c4_1),.din(w_dff_A_xsATXNB53_1),.clk(gclk));
	jdff dff_A_6D4cYah37_0(.dout(w_G338_0[0]),.din(w_dff_A_6D4cYah37_0),.clk(gclk));
	jdff dff_A_zLCi2JRf0_0(.dout(w_G514_0[0]),.din(w_dff_A_zLCi2JRf0_0),.clk(gclk));
	jdff dff_A_gqGYYdE64_0(.dout(w_dff_A_zLCi2JRf0_0),.din(w_dff_A_gqGYYdE64_0),.clk(gclk));
	jdff dff_A_qQCaPRpQ6_2(.dout(w_G514_0[2]),.din(w_dff_A_qQCaPRpQ6_2),.clk(gclk));
	jdff dff_A_WkeJW0YD8_1(.dout(w_n720_0[1]),.din(w_dff_A_WkeJW0YD8_1),.clk(gclk));
	jdff dff_A_ST5xq0FZ2_1(.dout(w_dff_A_WkeJW0YD8_1),.din(w_dff_A_ST5xq0FZ2_1),.clk(gclk));
	jdff dff_A_lPWQYr1d8_1(.dout(w_dff_A_ST5xq0FZ2_1),.din(w_dff_A_lPWQYr1d8_1),.clk(gclk));
	jdff dff_A_t6E3SN1s2_1(.dout(w_dff_A_lPWQYr1d8_1),.din(w_dff_A_t6E3SN1s2_1),.clk(gclk));
	jdff dff_A_IkVwVZtL1_1(.dout(w_n719_0[1]),.din(w_dff_A_IkVwVZtL1_1),.clk(gclk));
	jdff dff_A_PRGlszqX1_1(.dout(w_dff_A_IkVwVZtL1_1),.din(w_dff_A_PRGlszqX1_1),.clk(gclk));
	jdff dff_A_4IR1WgpV2_1(.dout(w_dff_A_PRGlszqX1_1),.din(w_dff_A_4IR1WgpV2_1),.clk(gclk));
	jdff dff_A_oen9cJMi5_1(.dout(w_dff_A_4IR1WgpV2_1),.din(w_dff_A_oen9cJMi5_1),.clk(gclk));
	jdff dff_A_lGvYCjGC7_1(.dout(w_dff_A_oen9cJMi5_1),.din(w_dff_A_lGvYCjGC7_1),.clk(gclk));
	jdff dff_B_2P7cnQJX2_0(.din(n616),.dout(w_dff_B_2P7cnQJX2_0),.clk(gclk));
	jdff dff_A_TLSq3PvQ6_1(.dout(w_G331_0[1]),.din(w_dff_A_TLSq3PvQ6_1),.clk(gclk));
	jdff dff_A_S9P1YKLL9_1(.dout(w_G324_1[1]),.din(w_dff_A_S9P1YKLL9_1),.clk(gclk));
	jdff dff_A_m0hJMGqo6_2(.dout(w_G324_0[2]),.din(w_dff_A_m0hJMGqo6_2),.clk(gclk));
	jdff dff_A_HNdEweL63_0(.dout(w_G503_0[0]),.din(w_dff_A_HNdEweL63_0),.clk(gclk));
	jdff dff_A_WCbEeCWh0_0(.dout(w_dff_A_HNdEweL63_0),.din(w_dff_A_WCbEeCWh0_0),.clk(gclk));
	jdff dff_A_hUPZcTEs3_0(.dout(w_dff_A_WCbEeCWh0_0),.din(w_dff_A_hUPZcTEs3_0),.clk(gclk));
	jdff dff_A_TkQf8VUZ5_0(.dout(w_dff_A_hUPZcTEs3_0),.din(w_dff_A_TkQf8VUZ5_0),.clk(gclk));
	jdff dff_A_vLlAh7BJ3_2(.dout(w_G503_0[2]),.din(w_dff_A_vLlAh7BJ3_2),.clk(gclk));
	jdff dff_A_z10QLZuZ2_2(.dout(w_dff_A_vLlAh7BJ3_2),.din(w_dff_A_z10QLZuZ2_2),.clk(gclk));
	jdff dff_A_InqCPwIB5_0(.dout(w_G4092_4[0]),.din(w_dff_A_InqCPwIB5_0),.clk(gclk));
	jdff dff_A_oaUI5gpT5_0(.dout(w_dff_A_InqCPwIB5_0),.din(w_dff_A_oaUI5gpT5_0),.clk(gclk));
	jdff dff_A_wNcPZAgX3_0(.dout(w_dff_A_oaUI5gpT5_0),.din(w_dff_A_wNcPZAgX3_0),.clk(gclk));
	jdff dff_A_QvcNGvMq9_0(.dout(w_dff_A_wNcPZAgX3_0),.din(w_dff_A_QvcNGvMq9_0),.clk(gclk));
	jdff dff_A_4xah8S4p1_0(.dout(w_dff_A_QvcNGvMq9_0),.din(w_dff_A_4xah8S4p1_0),.clk(gclk));
	jdff dff_A_yRq5rjgp0_0(.dout(w_dff_A_4xah8S4p1_0),.din(w_dff_A_yRq5rjgp0_0),.clk(gclk));
	jdff dff_A_uD75D0407_0(.dout(w_dff_A_yRq5rjgp0_0),.din(w_dff_A_uD75D0407_0),.clk(gclk));
	jdff dff_A_gfuM77xF0_0(.dout(w_dff_A_uD75D0407_0),.din(w_dff_A_gfuM77xF0_0),.clk(gclk));
	jdff dff_A_CmPNRQtJ1_0(.dout(w_dff_A_gfuM77xF0_0),.din(w_dff_A_CmPNRQtJ1_0),.clk(gclk));
	jdff dff_A_svdtNH7T0_0(.dout(w_dff_A_CmPNRQtJ1_0),.din(w_dff_A_svdtNH7T0_0),.clk(gclk));
	jdff dff_A_wNWBEMgF1_0(.dout(w_dff_A_svdtNH7T0_0),.din(w_dff_A_wNWBEMgF1_0),.clk(gclk));
	jdff dff_A_LeCjiudG4_0(.dout(w_dff_A_wNWBEMgF1_0),.din(w_dff_A_LeCjiudG4_0),.clk(gclk));
	jdff dff_A_xmAUHCQt2_0(.dout(w_dff_A_LeCjiudG4_0),.din(w_dff_A_xmAUHCQt2_0),.clk(gclk));
	jdff dff_A_4eBVXyyi9_0(.dout(w_dff_A_xmAUHCQt2_0),.din(w_dff_A_4eBVXyyi9_0),.clk(gclk));
	jdff dff_A_sGlV1iAw4_0(.dout(w_G4092_1[0]),.din(w_dff_A_sGlV1iAw4_0),.clk(gclk));
	jdff dff_A_FNNpIzeO2_0(.dout(w_dff_A_sGlV1iAw4_0),.din(w_dff_A_FNNpIzeO2_0),.clk(gclk));
	jdff dff_A_GSVGRiUH8_0(.dout(w_dff_A_FNNpIzeO2_0),.din(w_dff_A_GSVGRiUH8_0),.clk(gclk));
	jdff dff_A_HV17DwMK2_0(.dout(w_dff_A_GSVGRiUH8_0),.din(w_dff_A_HV17DwMK2_0),.clk(gclk));
	jdff dff_A_g0ILb4HI3_0(.dout(w_dff_A_HV17DwMK2_0),.din(w_dff_A_g0ILb4HI3_0),.clk(gclk));
	jdff dff_A_96sSh9NM1_0(.dout(w_dff_A_g0ILb4HI3_0),.din(w_dff_A_96sSh9NM1_0),.clk(gclk));
	jdff dff_A_xqfXnHMP0_2(.dout(w_G4092_1[2]),.din(w_dff_A_xqfXnHMP0_2),.clk(gclk));
	jdff dff_A_eq1D3zvb3_2(.dout(w_dff_A_xqfXnHMP0_2),.din(w_dff_A_eq1D3zvb3_2),.clk(gclk));
	jdff dff_A_q2I5Dvgu0_2(.dout(w_dff_A_eq1D3zvb3_2),.din(w_dff_A_q2I5Dvgu0_2),.clk(gclk));
	jdff dff_A_VHMWrw1t4_2(.dout(w_dff_A_q2I5Dvgu0_2),.din(w_dff_A_VHMWrw1t4_2),.clk(gclk));
	jdff dff_B_gUbshfRD5_0(.din(n1673),.dout(w_dff_B_gUbshfRD5_0),.clk(gclk));
	jdff dff_B_jhkjn9Zl4_0(.din(w_dff_B_gUbshfRD5_0),.dout(w_dff_B_jhkjn9Zl4_0),.clk(gclk));
	jdff dff_B_Uoi2yFh10_0(.din(w_dff_B_jhkjn9Zl4_0),.dout(w_dff_B_Uoi2yFh10_0),.clk(gclk));
	jdff dff_B_MVjIrnIv0_0(.din(w_dff_B_Uoi2yFh10_0),.dout(w_dff_B_MVjIrnIv0_0),.clk(gclk));
	jdff dff_B_Jm6O73Tk5_0(.din(w_dff_B_MVjIrnIv0_0),.dout(w_dff_B_Jm6O73Tk5_0),.clk(gclk));
	jdff dff_B_x3Qlmyke3_0(.din(w_dff_B_Jm6O73Tk5_0),.dout(w_dff_B_x3Qlmyke3_0),.clk(gclk));
	jdff dff_B_HrePYNtF4_0(.din(w_dff_B_x3Qlmyke3_0),.dout(w_dff_B_HrePYNtF4_0),.clk(gclk));
	jdff dff_B_esu3p3g65_0(.din(w_dff_B_HrePYNtF4_0),.dout(w_dff_B_esu3p3g65_0),.clk(gclk));
	jdff dff_B_ey1uRs3A9_0(.din(w_dff_B_esu3p3g65_0),.dout(w_dff_B_ey1uRs3A9_0),.clk(gclk));
	jdff dff_B_KILiCMsR7_0(.din(w_dff_B_ey1uRs3A9_0),.dout(w_dff_B_KILiCMsR7_0),.clk(gclk));
	jdff dff_B_d5Jx423d6_0(.din(w_dff_B_KILiCMsR7_0),.dout(w_dff_B_d5Jx423d6_0),.clk(gclk));
	jdff dff_B_5Y5w8VxY9_0(.din(w_dff_B_d5Jx423d6_0),.dout(w_dff_B_5Y5w8VxY9_0),.clk(gclk));
	jdff dff_B_OsgGniXa9_0(.din(w_dff_B_5Y5w8VxY9_0),.dout(w_dff_B_OsgGniXa9_0),.clk(gclk));
	jdff dff_B_0347uEnU6_0(.din(w_dff_B_OsgGniXa9_0),.dout(w_dff_B_0347uEnU6_0),.clk(gclk));
	jdff dff_B_v7oDXAX19_0(.din(w_dff_B_0347uEnU6_0),.dout(w_dff_B_v7oDXAX19_0),.clk(gclk));
	jdff dff_B_lZt7TFpo7_0(.din(w_dff_B_v7oDXAX19_0),.dout(w_dff_B_lZt7TFpo7_0),.clk(gclk));
	jdff dff_B_yjk0X1Kn2_0(.din(w_dff_B_lZt7TFpo7_0),.dout(w_dff_B_yjk0X1Kn2_0),.clk(gclk));
	jdff dff_B_qYAwu6Vt6_0(.din(w_dff_B_yjk0X1Kn2_0),.dout(w_dff_B_qYAwu6Vt6_0),.clk(gclk));
	jdff dff_B_nPiJfuQE9_0(.din(w_dff_B_qYAwu6Vt6_0),.dout(w_dff_B_nPiJfuQE9_0),.clk(gclk));
	jdff dff_B_0B4BLuop5_1(.din(n1588),.dout(w_dff_B_0B4BLuop5_1),.clk(gclk));
	jdff dff_B_OBGnQCwn1_1(.din(w_dff_B_0B4BLuop5_1),.dout(w_dff_B_OBGnQCwn1_1),.clk(gclk));
	jdff dff_B_i9avABce2_1(.din(w_dff_B_OBGnQCwn1_1),.dout(w_dff_B_i9avABce2_1),.clk(gclk));
	jdff dff_B_9tcoZrT43_1(.din(w_dff_B_i9avABce2_1),.dout(w_dff_B_9tcoZrT43_1),.clk(gclk));
	jdff dff_B_JS3lg73m1_1(.din(w_dff_B_9tcoZrT43_1),.dout(w_dff_B_JS3lg73m1_1),.clk(gclk));
	jdff dff_B_OtNKk3rR4_1(.din(w_dff_B_JS3lg73m1_1),.dout(w_dff_B_OtNKk3rR4_1),.clk(gclk));
	jdff dff_B_m5hu5P1z5_1(.din(w_dff_B_OtNKk3rR4_1),.dout(w_dff_B_m5hu5P1z5_1),.clk(gclk));
	jdff dff_B_uWVyz5F21_1(.din(w_dff_B_m5hu5P1z5_1),.dout(w_dff_B_uWVyz5F21_1),.clk(gclk));
	jdff dff_B_wuYXi2Et7_1(.din(n1655),.dout(w_dff_B_wuYXi2Et7_1),.clk(gclk));
	jdff dff_B_7mRl6pvf8_1(.din(w_dff_B_wuYXi2Et7_1),.dout(w_dff_B_7mRl6pvf8_1),.clk(gclk));
	jdff dff_A_c3JiXYI61_2(.dout(w_n588_0[2]),.din(w_dff_A_c3JiXYI61_2),.clk(gclk));
	jdff dff_A_YA6qdyAm1_2(.dout(w_dff_A_c3JiXYI61_2),.din(w_dff_A_YA6qdyAm1_2),.clk(gclk));
	jdff dff_A_ljs2Hp0w4_1(.dout(w_n1652_0[1]),.din(w_dff_A_ljs2Hp0w4_1),.clk(gclk));
	jdff dff_B_U39WYkVf8_0(.din(n1649),.dout(w_dff_B_U39WYkVf8_0),.clk(gclk));
	jdff dff_B_SkQjwMPL6_1(.din(n1645),.dout(w_dff_B_SkQjwMPL6_1),.clk(gclk));
	jdff dff_B_bhIyt8lL5_1(.din(w_dff_B_SkQjwMPL6_1),.dout(w_dff_B_bhIyt8lL5_1),.clk(gclk));
	jdff dff_B_G0JmWut19_1(.din(w_dff_B_bhIyt8lL5_1),.dout(w_dff_B_G0JmWut19_1),.clk(gclk));
	jdff dff_B_6F5f6ggu3_1(.din(w_dff_B_G0JmWut19_1),.dout(w_dff_B_6F5f6ggu3_1),.clk(gclk));
	jdff dff_B_gwOPQG2O0_1(.din(w_dff_B_6F5f6ggu3_1),.dout(w_dff_B_gwOPQG2O0_1),.clk(gclk));
	jdff dff_B_JKPtkImr4_1(.din(n1638),.dout(w_dff_B_JKPtkImr4_1),.clk(gclk));
	jdff dff_B_5EK2mvuK0_1(.din(w_dff_B_JKPtkImr4_1),.dout(w_dff_B_5EK2mvuK0_1),.clk(gclk));
	jdff dff_B_UN3D2OQa0_0(.din(n1641),.dout(w_dff_B_UN3D2OQa0_0),.clk(gclk));
	jdff dff_B_E9c8Q9st3_0(.din(n1640),.dout(w_dff_B_E9c8Q9st3_0),.clk(gclk));
	jdff dff_A_lMfFZB3f7_1(.dout(w_n609_0[1]),.din(w_dff_A_lMfFZB3f7_1),.clk(gclk));
	jdff dff_A_qN1R3Qou6_1(.dout(w_dff_A_lMfFZB3f7_1),.din(w_dff_A_qN1R3Qou6_1),.clk(gclk));
	jdff dff_A_uWkQqW285_1(.dout(w_dff_A_qN1R3Qou6_1),.din(w_dff_A_uWkQqW285_1),.clk(gclk));
	jdff dff_A_7StndMra4_1(.dout(w_dff_A_uWkQqW285_1),.din(w_dff_A_7StndMra4_1),.clk(gclk));
	jdff dff_A_kjlwGibM2_1(.dout(w_dff_A_7StndMra4_1),.din(w_dff_A_kjlwGibM2_1),.clk(gclk));
	jdff dff_A_6jSZxBw04_1(.dout(w_dff_A_kjlwGibM2_1),.din(w_dff_A_6jSZxBw04_1),.clk(gclk));
	jdff dff_A_GfGyIHtP2_1(.dout(w_dff_A_6jSZxBw04_1),.din(w_dff_A_GfGyIHtP2_1),.clk(gclk));
	jdff dff_A_ciDKAQsw9_1(.dout(w_n962_0[1]),.din(w_dff_A_ciDKAQsw9_1),.clk(gclk));
	jdff dff_A_LBtMs73U2_1(.dout(w_dff_A_ciDKAQsw9_1),.din(w_dff_A_LBtMs73U2_1),.clk(gclk));
	jdff dff_A_rg1LxCCa7_1(.dout(w_dff_A_LBtMs73U2_1),.din(w_dff_A_rg1LxCCa7_1),.clk(gclk));
	jdff dff_A_U290aPjM7_1(.dout(w_dff_A_rg1LxCCa7_1),.din(w_dff_A_U290aPjM7_1),.clk(gclk));
	jdff dff_A_EQXPIS1N9_1(.dout(w_dff_A_U290aPjM7_1),.din(w_dff_A_EQXPIS1N9_1),.clk(gclk));
	jdff dff_A_w7y9CaQb5_1(.dout(w_dff_A_EQXPIS1N9_1),.din(w_dff_A_w7y9CaQb5_1),.clk(gclk));
	jdff dff_B_ePa9ZGLr2_2(.din(n962),.dout(w_dff_B_ePa9ZGLr2_2),.clk(gclk));
	jdff dff_A_BTbKi5Jb9_2(.dout(w_n938_0[2]),.din(w_dff_A_BTbKi5Jb9_2),.clk(gclk));
	jdff dff_A_CH84g8MI4_2(.dout(w_dff_A_BTbKi5Jb9_2),.din(w_dff_A_CH84g8MI4_2),.clk(gclk));
	jdff dff_A_wVumRsB25_2(.dout(w_dff_A_CH84g8MI4_2),.din(w_dff_A_wVumRsB25_2),.clk(gclk));
	jdff dff_A_y94MvvgY3_2(.dout(w_dff_A_wVumRsB25_2),.din(w_dff_A_y94MvvgY3_2),.clk(gclk));
	jdff dff_A_Y4IRGbEd4_2(.dout(w_dff_A_y94MvvgY3_2),.din(w_dff_A_Y4IRGbEd4_2),.clk(gclk));
	jdff dff_B_HZ22xhO44_1(.din(n707),.dout(w_dff_B_HZ22xhO44_1),.clk(gclk));
	jdff dff_B_c8tJW17L9_1(.din(w_dff_B_HZ22xhO44_1),.dout(w_dff_B_c8tJW17L9_1),.clk(gclk));
	jdff dff_B_bM6Z8sTg3_1(.din(w_dff_B_c8tJW17L9_1),.dout(w_dff_B_bM6Z8sTg3_1),.clk(gclk));
	jdff dff_B_C3TFEuEu2_1(.din(n708),.dout(w_dff_B_C3TFEuEu2_1),.clk(gclk));
	jdff dff_B_JjKRjUFL6_1(.din(w_dff_B_C3TFEuEu2_1),.dout(w_dff_B_JjKRjUFL6_1),.clk(gclk));
	jdff dff_A_stEpA5I53_1(.dout(w_n713_0[1]),.din(w_dff_A_stEpA5I53_1),.clk(gclk));
	jdff dff_A_ltrH5PPd3_1(.dout(w_dff_A_stEpA5I53_1),.din(w_dff_A_ltrH5PPd3_1),.clk(gclk));
	jdff dff_A_DuemyRDn3_1(.dout(w_dff_A_ltrH5PPd3_1),.din(w_dff_A_DuemyRDn3_1),.clk(gclk));
	jdff dff_A_qtKn5Lti2_1(.dout(w_dff_A_DuemyRDn3_1),.din(w_dff_A_qtKn5Lti2_1),.clk(gclk));
	jdff dff_A_80AmkYVV1_1(.dout(w_dff_A_qtKn5Lti2_1),.din(w_dff_A_80AmkYVV1_1),.clk(gclk));
	jdff dff_A_TpXMtvpr4_1(.dout(w_dff_A_80AmkYVV1_1),.din(w_dff_A_TpXMtvpr4_1),.clk(gclk));
	jdff dff_A_OkWM4bmB6_1(.dout(w_dff_A_TpXMtvpr4_1),.din(w_dff_A_OkWM4bmB6_1),.clk(gclk));
	jdff dff_A_gA8xVCXm4_0(.dout(w_n710_0[0]),.din(w_dff_A_gA8xVCXm4_0),.clk(gclk));
	jdff dff_A_uWVn8Rrn5_0(.dout(w_dff_A_gA8xVCXm4_0),.din(w_dff_A_uWVn8Rrn5_0),.clk(gclk));
	jdff dff_A_nOmrw2Ua8_0(.dout(w_dff_A_uWVn8Rrn5_0),.din(w_dff_A_nOmrw2Ua8_0),.clk(gclk));
	jdff dff_A_NXxAqgyB4_0(.dout(w_dff_A_nOmrw2Ua8_0),.din(w_dff_A_NXxAqgyB4_0),.clk(gclk));
	jdff dff_A_NdelxAfF1_0(.dout(w_dff_A_NXxAqgyB4_0),.din(w_dff_A_NdelxAfF1_0),.clk(gclk));
	jdff dff_A_SZQgHzmo0_0(.dout(w_dff_A_NdelxAfF1_0),.din(w_dff_A_SZQgHzmo0_0),.clk(gclk));
	jdff dff_A_KOwUvZYr6_0(.dout(w_dff_A_SZQgHzmo0_0),.din(w_dff_A_KOwUvZYr6_0),.clk(gclk));
	jdff dff_A_x46xDeyz9_0(.dout(w_dff_A_KOwUvZYr6_0),.din(w_dff_A_x46xDeyz9_0),.clk(gclk));
	jdff dff_A_1IuIiZHH3_0(.dout(w_n597_0[0]),.din(w_dff_A_1IuIiZHH3_0),.clk(gclk));
	jdff dff_A_5DSV6Ion8_0(.dout(w_dff_A_1IuIiZHH3_0),.din(w_dff_A_5DSV6Ion8_0),.clk(gclk));
	jdff dff_A_5Z60IyI02_0(.dout(w_dff_A_5DSV6Ion8_0),.din(w_dff_A_5Z60IyI02_0),.clk(gclk));
	jdff dff_A_RoCQJvsK0_0(.dout(w_dff_A_5Z60IyI02_0),.din(w_dff_A_RoCQJvsK0_0),.clk(gclk));
	jdff dff_A_EUXMbap50_0(.dout(w_dff_A_RoCQJvsK0_0),.din(w_dff_A_EUXMbap50_0),.clk(gclk));
	jdff dff_A_c6yKdYy39_0(.dout(w_n496_1[0]),.din(w_dff_A_c6yKdYy39_0),.clk(gclk));
	jdff dff_A_eYoFTxR21_0(.dout(w_dff_A_c6yKdYy39_0),.din(w_dff_A_eYoFTxR21_0),.clk(gclk));
	jdff dff_A_0btEpyaX9_0(.dout(w_n1637_0[0]),.din(w_dff_A_0btEpyaX9_0),.clk(gclk));
	jdff dff_A_kwSz5bpb4_0(.dout(w_dff_A_0btEpyaX9_0),.din(w_dff_A_kwSz5bpb4_0),.clk(gclk));
	jdff dff_B_7gkPcXSF8_2(.din(n1637),.dout(w_dff_B_7gkPcXSF8_2),.clk(gclk));
	jdff dff_B_VeZvpyRk9_2(.din(w_dff_B_7gkPcXSF8_2),.dout(w_dff_B_VeZvpyRk9_2),.clk(gclk));
	jdff dff_A_y9p7nX1o0_1(.dout(w_n608_0[1]),.din(w_dff_A_y9p7nX1o0_1),.clk(gclk));
	jdff dff_A_oL2g4Aja4_1(.dout(w_dff_A_y9p7nX1o0_1),.din(w_dff_A_oL2g4Aja4_1),.clk(gclk));
	jdff dff_A_4fdym84U1_1(.dout(w_dff_A_oL2g4Aja4_1),.din(w_dff_A_4fdym84U1_1),.clk(gclk));
	jdff dff_A_on1XCH9Z5_1(.dout(w_dff_A_4fdym84U1_1),.din(w_dff_A_on1XCH9Z5_1),.clk(gclk));
	jdff dff_A_AuzC6GbR3_1(.dout(w_dff_A_on1XCH9Z5_1),.din(w_dff_A_AuzC6GbR3_1),.clk(gclk));
	jdff dff_A_yOnSseSd2_1(.dout(w_dff_A_AuzC6GbR3_1),.din(w_dff_A_yOnSseSd2_1),.clk(gclk));
	jdff dff_A_3c13K7Dr4_1(.dout(w_dff_A_yOnSseSd2_1),.din(w_dff_A_3c13K7Dr4_1),.clk(gclk));
	jdff dff_A_A412UALn6_1(.dout(w_dff_A_3c13K7Dr4_1),.din(w_dff_A_A412UALn6_1),.clk(gclk));
	jdff dff_A_KP6Onlmi6_1(.dout(w_dff_A_A412UALn6_1),.din(w_dff_A_KP6Onlmi6_1),.clk(gclk));
	jdff dff_A_TDWXxzhw2_1(.dout(w_dff_A_KP6Onlmi6_1),.din(w_dff_A_TDWXxzhw2_1),.clk(gclk));
	jdff dff_A_Tmt5fEaE8_2(.dout(w_n608_0[2]),.din(w_dff_A_Tmt5fEaE8_2),.clk(gclk));
	jdff dff_B_kxUpVWOD1_0(.din(n606),.dout(w_dff_B_kxUpVWOD1_0),.clk(gclk));
	jdff dff_B_FNT2I8yG7_1(.din(G217),.dout(w_dff_B_FNT2I8yG7_1),.clk(gclk));
	jdff dff_A_JafzU21e9_0(.dout(w_n592_0[0]),.din(w_dff_A_JafzU21e9_0),.clk(gclk));
	jdff dff_A_TJJFYm634_2(.dout(w_n592_0[2]),.din(w_dff_A_TJJFYm634_2),.clk(gclk));
	jdff dff_A_gUId8wQW0_2(.dout(w_dff_A_TJJFYm634_2),.din(w_dff_A_gUId8wQW0_2),.clk(gclk));
	jdff dff_A_OakfWlda1_2(.dout(w_dff_A_gUId8wQW0_2),.din(w_dff_A_OakfWlda1_2),.clk(gclk));
	jdff dff_A_YJMKUC0n2_2(.dout(w_dff_A_OakfWlda1_2),.din(w_dff_A_YJMKUC0n2_2),.clk(gclk));
	jdff dff_B_jofkP0gt7_1(.din(n589),.dout(w_dff_B_jofkP0gt7_1),.clk(gclk));
	jdff dff_B_tzD22bHC5_1(.din(G209),.dout(w_dff_B_tzD22bHC5_1),.clk(gclk));
	jdff dff_A_hh2mcvLz5_0(.dout(w_n602_0[0]),.din(w_dff_A_hh2mcvLz5_0),.clk(gclk));
	jdff dff_A_PLKQmBID7_0(.dout(w_n711_0[0]),.din(w_dff_A_PLKQmBID7_0),.clk(gclk));
	jdff dff_A_rsjm53rT8_0(.dout(w_dff_A_PLKQmBID7_0),.din(w_dff_A_rsjm53rT8_0),.clk(gclk));
	jdff dff_A_IhhqZhb00_2(.dout(w_n954_0[2]),.din(w_dff_A_IhhqZhb00_2),.clk(gclk));
	jdff dff_A_CVQrhsZZ8_2(.dout(w_dff_A_IhhqZhb00_2),.din(w_dff_A_CVQrhsZZ8_2),.clk(gclk));
	jdff dff_A_M19FBHYK2_2(.dout(w_dff_A_CVQrhsZZ8_2),.din(w_dff_A_M19FBHYK2_2),.clk(gclk));
	jdff dff_A_358nN0ZP7_2(.dout(w_dff_A_M19FBHYK2_2),.din(w_dff_A_358nN0ZP7_2),.clk(gclk));
	jdff dff_A_KDDCxiPb5_2(.dout(w_dff_A_358nN0ZP7_2),.din(w_dff_A_KDDCxiPb5_2),.clk(gclk));
	jdff dff_A_KcfKXmrH4_2(.dout(w_dff_A_KDDCxiPb5_2),.din(w_dff_A_KcfKXmrH4_2),.clk(gclk));
	jdff dff_A_ZuWMt4rq6_2(.dout(w_dff_A_KcfKXmrH4_2),.din(w_dff_A_ZuWMt4rq6_2),.clk(gclk));
	jdff dff_B_PBRYjV6g2_2(.din(n1633),.dout(w_dff_B_PBRYjV6g2_2),.clk(gclk));
	jdff dff_A_4qAEFu3Q1_1(.dout(w_n709_0[1]),.din(w_dff_A_4qAEFu3Q1_1),.clk(gclk));
	jdff dff_B_sEJck0bU6_0(.din(n600),.dout(w_dff_B_sEJck0bU6_0),.clk(gclk));
	jdff dff_B_jZXeDG7D1_1(.din(G225),.dout(w_dff_B_jZXeDG7D1_1),.clk(gclk));
	jdff dff_B_ZzFzfLkP7_0(.din(n595),.dout(w_dff_B_ZzFzfLkP7_0),.clk(gclk));
	jdff dff_B_Ky2Cc9Hx3_1(.din(G233),.dout(w_dff_B_Ky2Cc9Hx3_1),.clk(gclk));
	jdff dff_A_YX2jxMvL1_1(.dout(w_n703_0[1]),.din(w_dff_A_YX2jxMvL1_1),.clk(gclk));
	jdff dff_A_OSrep8xP9_0(.dout(w_n685_0[0]),.din(w_dff_A_OSrep8xP9_0),.clk(gclk));
	jdff dff_A_iM2l6I6p5_0(.dout(w_dff_A_OSrep8xP9_0),.din(w_dff_A_iM2l6I6p5_0),.clk(gclk));
	jdff dff_B_n2ov5BJX8_2(.din(n685),.dout(w_dff_B_n2ov5BJX8_2),.clk(gclk));
	jdff dff_B_jv55Wmyx7_2(.din(w_dff_B_n2ov5BJX8_2),.dout(w_dff_B_jv55Wmyx7_2),.clk(gclk));
	jdff dff_B_AW8r6ZLe9_2(.din(w_dff_B_jv55Wmyx7_2),.dout(w_dff_B_AW8r6ZLe9_2),.clk(gclk));
	jdff dff_A_wNyQiAG10_0(.dout(w_n684_0[0]),.din(w_dff_A_wNyQiAG10_0),.clk(gclk));
	jdff dff_A_TacHl0VK9_0(.dout(w_dff_A_wNyQiAG10_0),.din(w_dff_A_TacHl0VK9_0),.clk(gclk));
	jdff dff_A_ZNAEuJrn7_0(.dout(w_dff_A_TacHl0VK9_0),.din(w_dff_A_ZNAEuJrn7_0),.clk(gclk));
	jdff dff_A_ugD9qJRX6_0(.dout(w_dff_A_ZNAEuJrn7_0),.din(w_dff_A_ugD9qJRX6_0),.clk(gclk));
	jdff dff_A_LYdkwNnD8_1(.dout(w_n682_0[1]),.din(w_dff_A_LYdkwNnD8_1),.clk(gclk));
	jdff dff_A_NJrYn3Gh1_1(.dout(w_dff_A_LYdkwNnD8_1),.din(w_dff_A_NJrYn3Gh1_1),.clk(gclk));
	jdff dff_A_CvIrWNMh2_1(.dout(w_dff_A_NJrYn3Gh1_1),.din(w_dff_A_CvIrWNMh2_1),.clk(gclk));
	jdff dff_A_FqhyJarJ1_1(.dout(w_dff_A_CvIrWNMh2_1),.din(w_dff_A_FqhyJarJ1_1),.clk(gclk));
	jdff dff_A_ocVvc1Do8_1(.dout(w_dff_A_FqhyJarJ1_1),.din(w_dff_A_ocVvc1Do8_1),.clk(gclk));
	jdff dff_A_UqjqprCo5_1(.dout(w_dff_A_ocVvc1Do8_1),.din(w_dff_A_UqjqprCo5_1),.clk(gclk));
	jdff dff_A_rXYTpAJ86_2(.dout(w_n682_0[2]),.din(w_dff_A_rXYTpAJ86_2),.clk(gclk));
	jdff dff_A_mo4gCKNG7_2(.dout(w_dff_A_rXYTpAJ86_2),.din(w_dff_A_mo4gCKNG7_2),.clk(gclk));
	jdff dff_A_i0jTaJLg0_2(.dout(w_dff_A_mo4gCKNG7_2),.din(w_dff_A_i0jTaJLg0_2),.clk(gclk));
	jdff dff_A_3NsMfUTc1_2(.dout(w_dff_A_i0jTaJLg0_2),.din(w_dff_A_3NsMfUTc1_2),.clk(gclk));
	jdff dff_A_IN7IVVj00_2(.dout(w_dff_A_3NsMfUTc1_2),.din(w_dff_A_IN7IVVj00_2),.clk(gclk));
	jdff dff_A_SF6wwOlN4_2(.dout(w_dff_A_IN7IVVj00_2),.din(w_dff_A_SF6wwOlN4_2),.clk(gclk));
	jdff dff_B_YFbsgk1z0_0(.din(n1630),.dout(w_dff_B_YFbsgk1z0_0),.clk(gclk));
	jdff dff_B_kDISMzON5_0(.din(w_dff_B_YFbsgk1z0_0),.dout(w_dff_B_kDISMzON5_0),.clk(gclk));
	jdff dff_B_ADIfAWjU4_0(.din(w_dff_B_kDISMzON5_0),.dout(w_dff_B_ADIfAWjU4_0),.clk(gclk));
	jdff dff_B_x7MrCcHz2_0(.din(w_dff_B_ADIfAWjU4_0),.dout(w_dff_B_x7MrCcHz2_0),.clk(gclk));
	jdff dff_B_wfxsMGK99_0(.din(w_dff_B_x7MrCcHz2_0),.dout(w_dff_B_wfxsMGK99_0),.clk(gclk));
	jdff dff_B_J5FNLLdD9_0(.din(w_dff_B_wfxsMGK99_0),.dout(w_dff_B_J5FNLLdD9_0),.clk(gclk));
	jdff dff_B_oZBYRYpI6_0(.din(w_dff_B_J5FNLLdD9_0),.dout(w_dff_B_oZBYRYpI6_0),.clk(gclk));
	jdff dff_B_oBpoNX670_0(.din(w_dff_B_oZBYRYpI6_0),.dout(w_dff_B_oBpoNX670_0),.clk(gclk));
	jdff dff_B_IEWSCVWl1_0(.din(w_dff_B_oBpoNX670_0),.dout(w_dff_B_IEWSCVWl1_0),.clk(gclk));
	jdff dff_B_JSg1zwAr4_0(.din(n1628),.dout(w_dff_B_JSg1zwAr4_0),.clk(gclk));
	jdff dff_B_G6Afcqu25_0(.din(w_dff_B_JSg1zwAr4_0),.dout(w_dff_B_G6Afcqu25_0),.clk(gclk));
	jdff dff_B_FDhpUtO37_1(.din(n1625),.dout(w_dff_B_FDhpUtO37_1),.clk(gclk));
	jdff dff_B_zDJNFwb65_1(.din(n1623),.dout(w_dff_B_zDJNFwb65_1),.clk(gclk));
	jdff dff_B_DPIhoEAz3_1(.din(w_dff_B_zDJNFwb65_1),.dout(w_dff_B_DPIhoEAz3_1),.clk(gclk));
	jdff dff_A_WVPlABGB7_0(.dout(w_n1618_0[0]),.din(w_dff_A_WVPlABGB7_0),.clk(gclk));
	jdff dff_A_h9RHD1Wf3_0(.dout(w_dff_A_WVPlABGB7_0),.din(w_dff_A_h9RHD1Wf3_0),.clk(gclk));
	jdff dff_B_OSIpj3g87_2(.din(n1618),.dout(w_dff_B_OSIpj3g87_2),.clk(gclk));
	jdff dff_B_YdLpiqEO5_2(.din(w_dff_B_OSIpj3g87_2),.dout(w_dff_B_YdLpiqEO5_2),.clk(gclk));
	jdff dff_B_yzs8FEqX4_2(.din(w_dff_B_YdLpiqEO5_2),.dout(w_dff_B_yzs8FEqX4_2),.clk(gclk));
	jdff dff_B_AlB55ZbM5_2(.din(w_dff_B_yzs8FEqX4_2),.dout(w_dff_B_AlB55ZbM5_2),.clk(gclk));
	jdff dff_B_Iaidy7DC6_2(.din(w_dff_B_AlB55ZbM5_2),.dout(w_dff_B_Iaidy7DC6_2),.clk(gclk));
	jdff dff_B_SsKWya6U1_2(.din(w_dff_B_Iaidy7DC6_2),.dout(w_dff_B_SsKWya6U1_2),.clk(gclk));
	jdff dff_B_alvihZuQ4_2(.din(w_dff_B_SsKWya6U1_2),.dout(w_dff_B_alvihZuQ4_2),.clk(gclk));
	jdff dff_B_FA3jSb7Y0_2(.din(w_dff_B_alvihZuQ4_2),.dout(w_dff_B_FA3jSb7Y0_2),.clk(gclk));
	jdff dff_B_Q5W7Uo8m9_2(.din(w_dff_B_FA3jSb7Y0_2),.dout(w_dff_B_Q5W7Uo8m9_2),.clk(gclk));
	jdff dff_B_YJZ1q6Pt9_2(.din(w_dff_B_Q5W7Uo8m9_2),.dout(w_dff_B_YJZ1q6Pt9_2),.clk(gclk));
	jdff dff_B_fQAwXlFt3_2(.din(w_dff_B_YJZ1q6Pt9_2),.dout(w_dff_B_fQAwXlFt3_2),.clk(gclk));
	jdff dff_B_D23ryYxv9_2(.din(w_dff_B_fQAwXlFt3_2),.dout(w_dff_B_D23ryYxv9_2),.clk(gclk));
	jdff dff_A_DUQCjTfN9_0(.dout(w_G1497_0[0]),.din(w_dff_A_DUQCjTfN9_0),.clk(gclk));
	jdff dff_A_VYqd4jNF5_0(.dout(w_dff_A_DUQCjTfN9_0),.din(w_dff_A_VYqd4jNF5_0),.clk(gclk));
	jdff dff_A_MIM2syFJ0_0(.dout(w_dff_A_VYqd4jNF5_0),.din(w_dff_A_MIM2syFJ0_0),.clk(gclk));
	jdff dff_A_d8qdPqnj3_0(.dout(w_dff_A_MIM2syFJ0_0),.din(w_dff_A_d8qdPqnj3_0),.clk(gclk));
	jdff dff_A_wR4gVw5a5_0(.dout(w_dff_A_d8qdPqnj3_0),.din(w_dff_A_wR4gVw5a5_0),.clk(gclk));
	jdff dff_A_DaEx89iW2_0(.dout(w_dff_A_wR4gVw5a5_0),.din(w_dff_A_DaEx89iW2_0),.clk(gclk));
	jdff dff_A_pW7PwdB17_0(.dout(w_dff_A_DaEx89iW2_0),.din(w_dff_A_pW7PwdB17_0),.clk(gclk));
	jdff dff_A_EZENiS5G4_0(.dout(w_dff_A_pW7PwdB17_0),.din(w_dff_A_EZENiS5G4_0),.clk(gclk));
	jdff dff_A_9HPwoaT46_0(.dout(w_dff_A_EZENiS5G4_0),.din(w_dff_A_9HPwoaT46_0),.clk(gclk));
	jdff dff_A_QunGUQS16_0(.dout(w_dff_A_9HPwoaT46_0),.din(w_dff_A_QunGUQS16_0),.clk(gclk));
	jdff dff_A_Csaffvy12_0(.dout(w_dff_A_QunGUQS16_0),.din(w_dff_A_Csaffvy12_0),.clk(gclk));
	jdff dff_A_WSKbKUGS6_0(.dout(w_dff_A_Csaffvy12_0),.din(w_dff_A_WSKbKUGS6_0),.clk(gclk));
	jdff dff_A_6TlGoEjs4_0(.dout(w_dff_A_WSKbKUGS6_0),.din(w_dff_A_6TlGoEjs4_0),.clk(gclk));
	jdff dff_A_JnceUb9N1_0(.dout(w_dff_A_6TlGoEjs4_0),.din(w_dff_A_JnceUb9N1_0),.clk(gclk));
	jdff dff_A_DIXrA4Ol2_0(.dout(w_dff_A_JnceUb9N1_0),.din(w_dff_A_DIXrA4Ol2_0),.clk(gclk));
	jdff dff_A_v8jUiXyq4_1(.dout(w_G1497_0[1]),.din(w_dff_A_v8jUiXyq4_1),.clk(gclk));
	jdff dff_A_JkE1apyh3_1(.dout(w_dff_A_v8jUiXyq4_1),.din(w_dff_A_JkE1apyh3_1),.clk(gclk));
	jdff dff_A_Pl5Lvpbu9_1(.dout(w_dff_A_JkE1apyh3_1),.din(w_dff_A_Pl5Lvpbu9_1),.clk(gclk));
	jdff dff_A_87EKpOGc5_1(.dout(w_dff_A_Pl5Lvpbu9_1),.din(w_dff_A_87EKpOGc5_1),.clk(gclk));
	jdff dff_A_pCebwpN17_1(.dout(w_dff_A_87EKpOGc5_1),.din(w_dff_A_pCebwpN17_1),.clk(gclk));
	jdff dff_A_eaMzEqWO4_1(.dout(w_dff_A_pCebwpN17_1),.din(w_dff_A_eaMzEqWO4_1),.clk(gclk));
	jdff dff_A_baz8KZBT4_1(.dout(w_dff_A_eaMzEqWO4_1),.din(w_dff_A_baz8KZBT4_1),.clk(gclk));
	jdff dff_A_19Z73k5e8_1(.dout(w_dff_A_baz8KZBT4_1),.din(w_dff_A_19Z73k5e8_1),.clk(gclk));
	jdff dff_A_MXuOOcBD5_1(.dout(w_dff_A_19Z73k5e8_1),.din(w_dff_A_MXuOOcBD5_1),.clk(gclk));
	jdff dff_A_QEqPepFN4_1(.dout(w_dff_A_MXuOOcBD5_1),.din(w_dff_A_QEqPepFN4_1),.clk(gclk));
	jdff dff_A_sMBrycq73_1(.dout(w_dff_A_QEqPepFN4_1),.din(w_dff_A_sMBrycq73_1),.clk(gclk));
	jdff dff_A_kMGXyWAW2_1(.dout(w_dff_A_sMBrycq73_1),.din(w_dff_A_kMGXyWAW2_1),.clk(gclk));
	jdff dff_B_tz7vm4622_1(.din(n1600),.dout(w_dff_B_tz7vm4622_1),.clk(gclk));
	jdff dff_B_Is9FsIDa4_1(.din(w_dff_B_tz7vm4622_1),.dout(w_dff_B_Is9FsIDa4_1),.clk(gclk));
	jdff dff_B_AHzQ1bo01_0(.din(n1614),.dout(w_dff_B_AHzQ1bo01_0),.clk(gclk));
	jdff dff_B_xjVLJxhP0_0(.din(w_dff_B_AHzQ1bo01_0),.dout(w_dff_B_xjVLJxhP0_0),.clk(gclk));
	jdff dff_B_TbBjUpTs8_0(.din(w_dff_B_xjVLJxhP0_0),.dout(w_dff_B_TbBjUpTs8_0),.clk(gclk));
	jdff dff_B_Q7Fir2LH9_0(.din(w_dff_B_TbBjUpTs8_0),.dout(w_dff_B_Q7Fir2LH9_0),.clk(gclk));
	jdff dff_A_lOC6SxJh8_0(.dout(w_n1613_0[0]),.din(w_dff_A_lOC6SxJh8_0),.clk(gclk));
	jdff dff_A_sWAv6bEr5_0(.dout(w_dff_A_lOC6SxJh8_0),.din(w_dff_A_sWAv6bEr5_0),.clk(gclk));
	jdff dff_A_9dufPMrV9_0(.dout(w_n865_0[0]),.din(w_dff_A_9dufPMrV9_0),.clk(gclk));
	jdff dff_A_cwqlShOa0_0(.dout(w_dff_A_9dufPMrV9_0),.din(w_dff_A_cwqlShOa0_0),.clk(gclk));
	jdff dff_A_uS9qzP8y1_0(.dout(w_dff_A_cwqlShOa0_0),.din(w_dff_A_uS9qzP8y1_0),.clk(gclk));
	jdff dff_A_rKYk0v846_0(.dout(w_dff_A_uS9qzP8y1_0),.din(w_dff_A_rKYk0v846_0),.clk(gclk));
	jdff dff_A_RQoPWnei5_2(.dout(w_n865_0[2]),.din(w_dff_A_RQoPWnei5_2),.clk(gclk));
	jdff dff_A_dGHbC1GY5_2(.dout(w_dff_A_RQoPWnei5_2),.din(w_dff_A_dGHbC1GY5_2),.clk(gclk));
	jdff dff_A_IbaEiGjv0_2(.dout(w_dff_A_dGHbC1GY5_2),.din(w_dff_A_IbaEiGjv0_2),.clk(gclk));
	jdff dff_A_KIv1QUks9_2(.dout(w_dff_A_IbaEiGjv0_2),.din(w_dff_A_KIv1QUks9_2),.clk(gclk));
	jdff dff_A_K2zayzws2_2(.dout(w_dff_A_KIv1QUks9_2),.din(w_dff_A_K2zayzws2_2),.clk(gclk));
	jdff dff_A_ag8tbrgU9_1(.dout(w_n587_0[1]),.din(w_dff_A_ag8tbrgU9_1),.clk(gclk));
	jdff dff_A_ucRjPzjK9_1(.dout(w_dff_A_ag8tbrgU9_1),.din(w_dff_A_ucRjPzjK9_1),.clk(gclk));
	jdff dff_A_6Du1Sg0U4_1(.dout(w_dff_A_ucRjPzjK9_1),.din(w_dff_A_6Du1Sg0U4_1),.clk(gclk));
	jdff dff_A_cJouWD972_1(.dout(w_dff_A_6Du1Sg0U4_1),.din(w_dff_A_cJouWD972_1),.clk(gclk));
	jdff dff_B_0KfscTS83_0(.din(n585),.dout(w_dff_B_0KfscTS83_0),.clk(gclk));
	jdff dff_B_Cur9DqbV8_1(.din(G241),.dout(w_dff_B_Cur9DqbV8_1),.clk(gclk));
	jdff dff_B_NQuomSmT9_1(.din(n1601),.dout(w_dff_B_NQuomSmT9_1),.clk(gclk));
	jdff dff_B_dihszsxc3_1(.din(w_dff_B_NQuomSmT9_1),.dout(w_dff_B_dihszsxc3_1),.clk(gclk));
	jdff dff_B_ZBZ2h3Xx8_1(.din(w_dff_B_dihszsxc3_1),.dout(w_dff_B_ZBZ2h3Xx8_1),.clk(gclk));
	jdff dff_B_gJKpywDe3_1(.din(n1602),.dout(w_dff_B_gJKpywDe3_1),.clk(gclk));
	jdff dff_B_EEf1xN4e2_1(.din(w_dff_B_gJKpywDe3_1),.dout(w_dff_B_EEf1xN4e2_1),.clk(gclk));
	jdff dff_A_45ISubVn8_1(.dout(w_n687_0[1]),.din(w_dff_A_45ISubVn8_1),.clk(gclk));
	jdff dff_A_D0J2IDl14_1(.dout(w_dff_A_45ISubVn8_1),.din(w_dff_A_D0J2IDl14_1),.clk(gclk));
	jdff dff_A_JglAYIaa8_1(.dout(w_dff_A_D0J2IDl14_1),.din(w_dff_A_JglAYIaa8_1),.clk(gclk));
	jdff dff_A_RI7rXPLc3_1(.dout(w_n686_0[1]),.din(w_dff_A_RI7rXPLc3_1),.clk(gclk));
	jdff dff_A_B7oKu7HL8_1(.dout(w_dff_A_RI7rXPLc3_1),.din(w_dff_A_B7oKu7HL8_1),.clk(gclk));
	jdff dff_A_jkr9Psjl4_1(.dout(w_dff_A_B7oKu7HL8_1),.din(w_dff_A_jkr9Psjl4_1),.clk(gclk));
	jdff dff_A_afZGM9lt3_1(.dout(w_dff_A_jkr9Psjl4_1),.din(w_dff_A_afZGM9lt3_1),.clk(gclk));
	jdff dff_A_t4w4FOuA7_0(.dout(w_n581_0[0]),.din(w_dff_A_t4w4FOuA7_0),.clk(gclk));
	jdff dff_A_L6sGAcEm1_0(.dout(w_dff_A_t4w4FOuA7_0),.din(w_dff_A_L6sGAcEm1_0),.clk(gclk));
	jdff dff_A_bYjMFFCb7_1(.dout(w_n579_1[1]),.din(w_dff_A_bYjMFFCb7_1),.clk(gclk));
	jdff dff_A_7jgF267z0_1(.dout(w_n579_0[1]),.din(w_dff_A_7jgF267z0_1),.clk(gclk));
	jdff dff_A_0Db6W2Cs6_2(.dout(w_n579_0[2]),.din(w_dff_A_0Db6W2Cs6_2),.clk(gclk));
	jdff dff_A_Fg9V4URE0_2(.dout(w_dff_A_0Db6W2Cs6_2),.din(w_dff_A_Fg9V4URE0_2),.clk(gclk));
	jdff dff_A_ImOe7M6h4_2(.dout(w_dff_A_Fg9V4URE0_2),.din(w_dff_A_ImOe7M6h4_2),.clk(gclk));
	jdff dff_A_C7zORkRV9_2(.dout(w_dff_A_ImOe7M6h4_2),.din(w_dff_A_C7zORkRV9_2),.clk(gclk));
	jdff dff_B_Fapaexz99_0(.din(n577),.dout(w_dff_B_Fapaexz99_0),.clk(gclk));
	jdff dff_B_NKyFj8YE6_1(.din(G264),.dout(w_dff_B_NKyFj8YE6_1),.clk(gclk));
	jdff dff_A_rXySgHot6_1(.dout(w_n574_0[1]),.din(w_dff_A_rXySgHot6_1),.clk(gclk));
	jdff dff_A_7iIMNZtS0_1(.dout(w_dff_A_rXySgHot6_1),.din(w_dff_A_7iIMNZtS0_1),.clk(gclk));
	jdff dff_A_CarUYmxb5_0(.dout(w_n1599_0[0]),.din(w_dff_A_CarUYmxb5_0),.clk(gclk));
	jdff dff_A_eMdoammx6_0(.dout(w_dff_A_CarUYmxb5_0),.din(w_dff_A_eMdoammx6_0),.clk(gclk));
	jdff dff_B_Vaz3kXuR5_0(.din(n1598),.dout(w_dff_B_Vaz3kXuR5_0),.clk(gclk));
	jdff dff_B_8Zp4ATZI9_0(.din(n1597),.dout(w_dff_B_8Zp4ATZI9_0),.clk(gclk));
	jdff dff_B_Ucp90mZP1_0(.din(n1589),.dout(w_dff_B_Ucp90mZP1_0),.clk(gclk));
	jdff dff_A_UYNv0ANo9_0(.dout(w_n573_0[0]),.din(w_dff_A_UYNv0ANo9_0),.clk(gclk));
	jdff dff_A_SdSKvjXD5_1(.dout(w_n573_0[1]),.din(w_dff_A_SdSKvjXD5_1),.clk(gclk));
	jdff dff_A_VwBB50Uj6_1(.dout(w_dff_A_SdSKvjXD5_1),.din(w_dff_A_VwBB50Uj6_1),.clk(gclk));
	jdff dff_B_5KEEzPuo0_1(.din(n691),.dout(w_dff_B_5KEEzPuo0_1),.clk(gclk));
	jdff dff_A_Mo0cBftB0_0(.dout(w_n695_0[0]),.din(w_dff_A_Mo0cBftB0_0),.clk(gclk));
	jdff dff_A_GzWpiUJQ3_1(.dout(w_n695_0[1]),.din(w_dff_A_GzWpiUJQ3_1),.clk(gclk));
	jdff dff_A_mYwDRUot2_1(.dout(w_n564_0[1]),.din(w_dff_A_mYwDRUot2_1),.clk(gclk));
	jdff dff_B_3wc4Nap28_1(.din(G280),.dout(w_dff_B_3wc4Nap28_1),.clk(gclk));
	jdff dff_A_uhsIQN6V4_0(.dout(w_n562_0[0]),.din(w_dff_A_uhsIQN6V4_0),.clk(gclk));
	jdff dff_A_A2GZ60vW9_0(.dout(w_n692_0[0]),.din(w_dff_A_A2GZ60vW9_0),.clk(gclk));
	jdff dff_A_cSQndLGD4_1(.dout(w_n559_0[1]),.din(w_dff_A_cSQndLGD4_1),.clk(gclk));
	jdff dff_B_StTsmORO0_1(.din(G288),.dout(w_dff_B_StTsmORO0_1),.clk(gclk));
	jdff dff_A_0k8lOAaf5_0(.dout(w_n557_0[0]),.din(w_dff_A_0k8lOAaf5_0),.clk(gclk));
	jdff dff_A_BgJsq9Jr0_0(.dout(w_n690_0[0]),.din(w_dff_A_BgJsq9Jr0_0),.clk(gclk));
	jdff dff_A_H1PaAqjw8_0(.dout(w_dff_A_BgJsq9Jr0_0),.din(w_dff_A_H1PaAqjw8_0),.clk(gclk));
	jdff dff_A_BEGkXa3p6_1(.dout(w_n571_0[1]),.din(w_dff_A_BEGkXa3p6_1),.clk(gclk));
	jdff dff_B_bwLRLfw68_1(.din(G272),.dout(w_dff_B_bwLRLfw68_1),.clk(gclk));
	jdff dff_A_6ICbiHw30_0(.dout(w_n569_0[0]),.din(w_dff_A_6ICbiHw30_0),.clk(gclk));
	jdff dff_A_2d6Dcsjh5_0(.dout(w_n485_1[0]),.din(w_dff_A_2d6Dcsjh5_0),.clk(gclk));
	jdff dff_A_S32Xyl0Y1_0(.dout(w_dff_A_2d6Dcsjh5_0),.din(w_dff_A_S32Xyl0Y1_0),.clk(gclk));
	jdff dff_B_QkIf4nKc5_0(.din(n1585),.dout(w_dff_B_QkIf4nKc5_0),.clk(gclk));
	jdff dff_B_RNCmrvdz4_1(.din(n1575),.dout(w_dff_B_RNCmrvdz4_1),.clk(gclk));
	jdff dff_B_bsFFLQAk9_1(.din(w_dff_B_RNCmrvdz4_1),.dout(w_dff_B_bsFFLQAk9_1),.clk(gclk));
	jdff dff_A_omW0t1800_0(.dout(w_G210_2[0]),.din(w_dff_A_omW0t1800_0),.clk(gclk));
	jdff dff_A_bo21x2F13_1(.dout(w_n451_0[1]),.din(w_dff_A_bo21x2F13_1),.clk(gclk));
	jdff dff_A_sxn8HzZ62_1(.dout(w_dff_A_bo21x2F13_1),.din(w_dff_A_sxn8HzZ62_1),.clk(gclk));
	jdff dff_B_258BLKiQ6_3(.din(n451),.dout(w_dff_B_258BLKiQ6_3),.clk(gclk));
	jdff dff_A_x8EnYzKe3_0(.dout(w_G457_1[0]),.din(w_dff_A_x8EnYzKe3_0),.clk(gclk));
	jdff dff_A_lIpRGklZ4_0(.dout(w_dff_A_x8EnYzKe3_0),.din(w_dff_A_lIpRGklZ4_0),.clk(gclk));
	jdff dff_A_JSUas53y4_0(.dout(w_dff_A_lIpRGklZ4_0),.din(w_dff_A_JSUas53y4_0),.clk(gclk));
	jdff dff_A_zRCf7qQ64_0(.dout(w_dff_A_JSUas53y4_0),.din(w_dff_A_zRCf7qQ64_0),.clk(gclk));
	jdff dff_A_H425gTGF7_1(.dout(w_G457_1[1]),.din(w_dff_A_H425gTGF7_1),.clk(gclk));
	jdff dff_A_K7zQGfJv1_1(.dout(w_dff_A_H425gTGF7_1),.din(w_dff_A_K7zQGfJv1_1),.clk(gclk));
	jdff dff_A_rP4Wqp0u9_1(.dout(w_dff_A_K7zQGfJv1_1),.din(w_dff_A_rP4Wqp0u9_1),.clk(gclk));
	jdff dff_A_ffHonvao3_1(.dout(w_G457_0[1]),.din(w_dff_A_ffHonvao3_1),.clk(gclk));
	jdff dff_A_VWxaRlu41_1(.dout(w_dff_A_ffHonvao3_1),.din(w_dff_A_VWxaRlu41_1),.clk(gclk));
	jdff dff_A_JYLhTTJa8_1(.dout(w_dff_A_VWxaRlu41_1),.din(w_dff_A_JYLhTTJa8_1),.clk(gclk));
	jdff dff_A_OG0liO9r0_2(.dout(w_G457_0[2]),.din(w_dff_A_OG0liO9r0_2),.clk(gclk));
	jdff dff_A_UiraPyUx6_2(.dout(w_dff_A_OG0liO9r0_2),.din(w_dff_A_UiraPyUx6_2),.clk(gclk));
	jdff dff_A_7uH9SFkI4_2(.dout(w_dff_A_UiraPyUx6_2),.din(w_dff_A_7uH9SFkI4_2),.clk(gclk));
	jdff dff_A_YnWKwscH0_2(.dout(w_dff_A_7uH9SFkI4_2),.din(w_dff_A_YnWKwscH0_2),.clk(gclk));
	jdff dff_A_VsQiZBHr3_2(.dout(w_G210_0[2]),.din(w_dff_A_VsQiZBHr3_2),.clk(gclk));
	jdff dff_B_UJdiGdRT3_1(.din(n1570),.dout(w_dff_B_UJdiGdRT3_1),.clk(gclk));
	jdff dff_A_NUipEbn84_0(.dout(w_n509_0[0]),.din(w_dff_A_NUipEbn84_0),.clk(gclk));
	jdff dff_A_yqjocQrS5_1(.dout(w_n509_0[1]),.din(w_dff_A_yqjocQrS5_1),.clk(gclk));
	jdff dff_A_oZTYeJI77_1(.dout(w_dff_A_yqjocQrS5_1),.din(w_dff_A_oZTYeJI77_1),.clk(gclk));
	jdff dff_B_Ue2RQK7M0_3(.din(n509),.dout(w_dff_B_Ue2RQK7M0_3),.clk(gclk));
	jdff dff_A_2giIdlF59_0(.dout(w_G468_1[0]),.din(w_dff_A_2giIdlF59_0),.clk(gclk));
	jdff dff_A_jOcXBYqR5_0(.dout(w_dff_A_2giIdlF59_0),.din(w_dff_A_jOcXBYqR5_0),.clk(gclk));
	jdff dff_A_a0tbMto75_0(.dout(w_dff_A_jOcXBYqR5_0),.din(w_dff_A_a0tbMto75_0),.clk(gclk));
	jdff dff_A_NyAn2Iwl2_0(.dout(w_dff_A_a0tbMto75_0),.din(w_dff_A_NyAn2Iwl2_0),.clk(gclk));
	jdff dff_A_C9EHR4nj9_1(.dout(w_G468_1[1]),.din(w_dff_A_C9EHR4nj9_1),.clk(gclk));
	jdff dff_A_gMChsRxG9_1(.dout(w_dff_A_C9EHR4nj9_1),.din(w_dff_A_gMChsRxG9_1),.clk(gclk));
	jdff dff_A_zp28VQpV5_1(.dout(w_dff_A_gMChsRxG9_1),.din(w_dff_A_zp28VQpV5_1),.clk(gclk));
	jdff dff_B_gJhV3tqA0_1(.din(n1566),.dout(w_dff_B_gJhV3tqA0_1),.clk(gclk));
	jdff dff_A_2dgVSwNM7_0(.dout(w_G218_1[0]),.din(w_dff_A_2dgVSwNM7_0),.clk(gclk));
	jdff dff_A_200NXoVi2_1(.dout(w_G468_0[1]),.din(w_dff_A_200NXoVi2_1),.clk(gclk));
	jdff dff_A_gqiZzrv91_1(.dout(w_dff_A_200NXoVi2_1),.din(w_dff_A_gqiZzrv91_1),.clk(gclk));
	jdff dff_A_BoSwSDQu9_2(.dout(w_G468_0[2]),.din(w_dff_A_BoSwSDQu9_2),.clk(gclk));
	jdff dff_A_HK9ADDy74_2(.dout(w_dff_A_BoSwSDQu9_2),.din(w_dff_A_HK9ADDy74_2),.clk(gclk));
	jdff dff_A_9tsMg1EG3_2(.dout(w_dff_A_HK9ADDy74_2),.din(w_dff_A_9tsMg1EG3_2),.clk(gclk));
	jdff dff_A_oN5HW0EJ7_2(.dout(w_dff_A_9tsMg1EG3_2),.din(w_dff_A_oN5HW0EJ7_2),.clk(gclk));
	jdff dff_A_snz3ufaQ5_0(.dout(w_G218_2[0]),.din(w_dff_A_snz3ufaQ5_0),.clk(gclk));
	jdff dff_B_zh9yCmRY4_1(.din(n1556),.dout(w_dff_B_zh9yCmRY4_1),.clk(gclk));
	jdff dff_B_2COnfUBI7_1(.din(w_dff_B_zh9yCmRY4_1),.dout(w_dff_B_2COnfUBI7_1),.clk(gclk));
	jdff dff_A_vLQ3zUm74_0(.dout(w_G226_2[0]),.din(w_dff_A_vLQ3zUm74_0),.clk(gclk));
	jdff dff_A_7UYuPrNg3_2(.dout(w_n496_0[2]),.din(w_dff_A_7UYuPrNg3_2),.clk(gclk));
	jdff dff_A_7ItgWThO1_2(.dout(w_dff_A_7UYuPrNg3_2),.din(w_dff_A_7ItgWThO1_2),.clk(gclk));
	jdff dff_A_du6Mz9Sf0_2(.dout(w_dff_A_7ItgWThO1_2),.din(w_dff_A_du6Mz9Sf0_2),.clk(gclk));
	jdff dff_B_6xukRhGQ8_3(.din(n496),.dout(w_dff_B_6xukRhGQ8_3),.clk(gclk));
	jdff dff_A_YVqMVdyg0_0(.dout(w_G422_1[0]),.din(w_dff_A_YVqMVdyg0_0),.clk(gclk));
	jdff dff_A_vTodZrR70_0(.dout(w_dff_A_YVqMVdyg0_0),.din(w_dff_A_vTodZrR70_0),.clk(gclk));
	jdff dff_A_4FNS6t941_0(.dout(w_dff_A_vTodZrR70_0),.din(w_dff_A_4FNS6t941_0),.clk(gclk));
	jdff dff_A_8ScpLo9y0_1(.dout(w_G422_0[1]),.din(w_dff_A_8ScpLo9y0_1),.clk(gclk));
	jdff dff_A_bqMEHnsB8_1(.dout(w_dff_A_8ScpLo9y0_1),.din(w_dff_A_bqMEHnsB8_1),.clk(gclk));
	jdff dff_A_ihL37Hwh1_1(.dout(w_dff_A_bqMEHnsB8_1),.din(w_dff_A_ihL37Hwh1_1),.clk(gclk));
	jdff dff_A_G2By6A9Y4_2(.dout(w_G422_0[2]),.din(w_dff_A_G2By6A9Y4_2),.clk(gclk));
	jdff dff_A_4vwKSeA09_2(.dout(w_dff_A_G2By6A9Y4_2),.din(w_dff_A_4vwKSeA09_2),.clk(gclk));
	jdff dff_A_0X6XxiFk2_2(.dout(w_dff_A_4vwKSeA09_2),.din(w_dff_A_0X6XxiFk2_2),.clk(gclk));
	jdff dff_A_RGIhfKH47_2(.dout(w_dff_A_0X6XxiFk2_2),.din(w_dff_A_RGIhfKH47_2),.clk(gclk));
	jdff dff_A_YFIgcURp7_2(.dout(w_G226_0[2]),.din(w_dff_A_YFIgcURp7_2),.clk(gclk));
	jdff dff_B_sXS2qhCh4_1(.din(n541),.dout(w_dff_B_sXS2qhCh4_1),.clk(gclk));
	jdff dff_B_0MDGyf1J3_1(.din(w_dff_B_sXS2qhCh4_1),.dout(w_dff_B_0MDGyf1J3_1),.clk(gclk));
	jdff dff_B_mxxOHVf20_1(.din(n542),.dout(w_dff_B_mxxOHVf20_1),.clk(gclk));
	jdff dff_A_tSgzqsuZ7_0(.dout(w_G446_1[0]),.din(w_dff_A_tSgzqsuZ7_0),.clk(gclk));
	jdff dff_A_c6yY6VmJ3_0(.dout(w_dff_A_tSgzqsuZ7_0),.din(w_dff_A_c6yY6VmJ3_0),.clk(gclk));
	jdff dff_A_cdMgZoFv3_0(.dout(w_dff_A_c6yY6VmJ3_0),.din(w_dff_A_cdMgZoFv3_0),.clk(gclk));
	jdff dff_A_oZKcgZqF6_1(.dout(w_G446_1[1]),.din(w_dff_A_oZKcgZqF6_1),.clk(gclk));
	jdff dff_A_H47IajYI2_1(.dout(w_dff_A_oZKcgZqF6_1),.din(w_dff_A_H47IajYI2_1),.clk(gclk));
	jdff dff_A_vPJtS8657_1(.dout(w_dff_A_H47IajYI2_1),.din(w_dff_A_vPJtS8657_1),.clk(gclk));
	jdff dff_A_RXlqpMv45_1(.dout(w_G446_0[1]),.din(w_dff_A_RXlqpMv45_1),.clk(gclk));
	jdff dff_A_CriMmbkp3_1(.dout(w_dff_A_RXlqpMv45_1),.din(w_dff_A_CriMmbkp3_1),.clk(gclk));
	jdff dff_A_DwvbHT6D0_1(.dout(w_dff_A_CriMmbkp3_1),.din(w_dff_A_DwvbHT6D0_1),.clk(gclk));
	jdff dff_A_8yUT8lxV7_2(.dout(w_G446_0[2]),.din(w_dff_A_8yUT8lxV7_2),.clk(gclk));
	jdff dff_A_REAC3s3q9_2(.dout(w_dff_A_8yUT8lxV7_2),.din(w_dff_A_REAC3s3q9_2),.clk(gclk));
	jdff dff_A_f2gP5ZVl5_2(.dout(w_dff_A_REAC3s3q9_2),.din(w_dff_A_f2gP5ZVl5_2),.clk(gclk));
	jdff dff_A_1F6tAt515_0(.dout(w_G206_1[0]),.din(w_dff_A_1F6tAt515_0),.clk(gclk));
	jdff dff_B_BsXdgS7b2_1(.din(n1525),.dout(w_dff_B_BsXdgS7b2_1),.clk(gclk));
	jdff dff_B_Se3SyzF83_1(.din(n1534),.dout(w_dff_B_Se3SyzF83_1),.clk(gclk));
	jdff dff_B_6CGQjU6n3_1(.din(n1544),.dout(w_dff_B_6CGQjU6n3_1),.clk(gclk));
	jdff dff_B_ak0qsddl7_1(.din(w_dff_B_6CGQjU6n3_1),.dout(w_dff_B_ak0qsddl7_1),.clk(gclk));
	jdff dff_A_fMp54LYZ8_0(.dout(w_G234_2[0]),.din(w_dff_A_fMp54LYZ8_0),.clk(gclk));
	jdff dff_A_4qNnXdDp7_1(.dout(w_n462_0[1]),.din(w_dff_A_4qNnXdDp7_1),.clk(gclk));
	jdff dff_A_ZakBxiGE0_1(.dout(w_dff_A_4qNnXdDp7_1),.din(w_dff_A_ZakBxiGE0_1),.clk(gclk));
	jdff dff_A_QQ58oc3Q7_1(.dout(w_dff_A_ZakBxiGE0_1),.din(w_dff_A_QQ58oc3Q7_1),.clk(gclk));
	jdff dff_B_4IsApSZi4_3(.din(n462),.dout(w_dff_B_4IsApSZi4_3),.clk(gclk));
	jdff dff_A_vF4BLX0l8_0(.dout(w_G435_1[0]),.din(w_dff_A_vF4BLX0l8_0),.clk(gclk));
	jdff dff_A_hDLByAA12_0(.dout(w_dff_A_vF4BLX0l8_0),.din(w_dff_A_hDLByAA12_0),.clk(gclk));
	jdff dff_A_DTh41GJm9_0(.dout(w_dff_A_hDLByAA12_0),.din(w_dff_A_DTh41GJm9_0),.clk(gclk));
	jdff dff_A_wpZAXwbu1_0(.dout(w_dff_A_DTh41GJm9_0),.din(w_dff_A_wpZAXwbu1_0),.clk(gclk));
	jdff dff_A_WMPP5CPu1_1(.dout(w_G435_1[1]),.din(w_dff_A_WMPP5CPu1_1),.clk(gclk));
	jdff dff_A_fcXknSva2_1(.dout(w_dff_A_WMPP5CPu1_1),.din(w_dff_A_fcXknSva2_1),.clk(gclk));
	jdff dff_A_LDaXALsP2_1(.dout(w_dff_A_fcXknSva2_1),.din(w_dff_A_LDaXALsP2_1),.clk(gclk));
	jdff dff_A_QrOT8bW25_1(.dout(w_G435_0[1]),.din(w_dff_A_QrOT8bW25_1),.clk(gclk));
	jdff dff_A_3hQrz8kn9_1(.dout(w_dff_A_QrOT8bW25_1),.din(w_dff_A_3hQrz8kn9_1),.clk(gclk));
	jdff dff_A_BvM1Ub6G2_1(.dout(w_dff_A_3hQrz8kn9_1),.din(w_dff_A_BvM1Ub6G2_1),.clk(gclk));
	jdff dff_A_vc9gITJm9_2(.dout(w_G435_0[2]),.din(w_dff_A_vc9gITJm9_2),.clk(gclk));
	jdff dff_A_rLV5VGiu1_2(.dout(w_dff_A_vc9gITJm9_2),.din(w_dff_A_rLV5VGiu1_2),.clk(gclk));
	jdff dff_A_5PKAwhTq9_2(.dout(w_dff_A_rLV5VGiu1_2),.din(w_dff_A_5PKAwhTq9_2),.clk(gclk));
	jdff dff_A_VR5MfvCi8_2(.dout(w_dff_A_5PKAwhTq9_2),.din(w_dff_A_VR5MfvCi8_2),.clk(gclk));
	jdff dff_A_Vdnrw3Gg7_2(.dout(w_G234_0[2]),.din(w_dff_A_Vdnrw3Gg7_2),.clk(gclk));
	jdff dff_B_K9GTT0wg4_1(.din(n1535),.dout(w_dff_B_K9GTT0wg4_1),.clk(gclk));
	jdff dff_B_qUqFTHDw7_1(.din(w_dff_B_K9GTT0wg4_1),.dout(w_dff_B_qUqFTHDw7_1),.clk(gclk));
	jdff dff_A_9iZVWSZd3_0(.dout(w_G257_2[0]),.din(w_dff_A_9iZVWSZd3_0),.clk(gclk));
	jdff dff_A_4nlF569f1_1(.dout(w_n520_0[1]),.din(w_dff_A_4nlF569f1_1),.clk(gclk));
	jdff dff_A_nw1q9Y2Y4_1(.dout(w_dff_A_4nlF569f1_1),.din(w_dff_A_nw1q9Y2Y4_1),.clk(gclk));
	jdff dff_B_kmWkYj5y6_3(.din(n520),.dout(w_dff_B_kmWkYj5y6_3),.clk(gclk));
	jdff dff_A_IOBuc7UP6_0(.dout(w_G389_1[0]),.din(w_dff_A_IOBuc7UP6_0),.clk(gclk));
	jdff dff_A_UXUCxW953_0(.dout(w_dff_A_IOBuc7UP6_0),.din(w_dff_A_UXUCxW953_0),.clk(gclk));
	jdff dff_A_0ZgOqPy23_0(.dout(w_dff_A_UXUCxW953_0),.din(w_dff_A_0ZgOqPy23_0),.clk(gclk));
	jdff dff_A_JzflguxI3_0(.dout(w_dff_A_0ZgOqPy23_0),.din(w_dff_A_JzflguxI3_0),.clk(gclk));
	jdff dff_A_ahzRbivf3_1(.dout(w_G389_1[1]),.din(w_dff_A_ahzRbivf3_1),.clk(gclk));
	jdff dff_A_sbbtQKiI3_1(.dout(w_dff_A_ahzRbivf3_1),.din(w_dff_A_sbbtQKiI3_1),.clk(gclk));
	jdff dff_A_tMFfg7EN9_1(.dout(w_dff_A_sbbtQKiI3_1),.din(w_dff_A_tMFfg7EN9_1),.clk(gclk));
	jdff dff_A_YubtN7nb5_1(.dout(w_G389_0[1]),.din(w_dff_A_YubtN7nb5_1),.clk(gclk));
	jdff dff_A_WPD1xqto1_1(.dout(w_dff_A_YubtN7nb5_1),.din(w_dff_A_WPD1xqto1_1),.clk(gclk));
	jdff dff_A_4Ezae2bB4_1(.dout(w_dff_A_WPD1xqto1_1),.din(w_dff_A_4Ezae2bB4_1),.clk(gclk));
	jdff dff_A_lj0sqnUK5_2(.dout(w_G389_0[2]),.din(w_dff_A_lj0sqnUK5_2),.clk(gclk));
	jdff dff_A_p882NBI01_2(.dout(w_dff_A_lj0sqnUK5_2),.din(w_dff_A_p882NBI01_2),.clk(gclk));
	jdff dff_A_BO0txMcK0_2(.dout(w_dff_A_p882NBI01_2),.din(w_dff_A_BO0txMcK0_2),.clk(gclk));
	jdff dff_A_spaQFyFL5_2(.dout(w_dff_A_BO0txMcK0_2),.din(w_dff_A_spaQFyFL5_2),.clk(gclk));
	jdff dff_A_UCUdfuzf8_2(.dout(w_G257_0[2]),.din(w_dff_A_UCUdfuzf8_2),.clk(gclk));
	jdff dff_B_E6Ivhjnj0_1(.din(n1530),.dout(w_dff_B_E6Ivhjnj0_1),.clk(gclk));
	jdff dff_A_6GrVvIMI8_1(.dout(w_n485_0[1]),.din(w_dff_A_6GrVvIMI8_1),.clk(gclk));
	jdff dff_A_WxCttBwT4_1(.dout(w_dff_A_6GrVvIMI8_1),.din(w_dff_A_WxCttBwT4_1),.clk(gclk));
	jdff dff_A_MkVZMfz07_2(.dout(w_n485_0[2]),.din(w_dff_A_MkVZMfz07_2),.clk(gclk));
	jdff dff_B_Vi4jOAZY0_3(.din(n485),.dout(w_dff_B_Vi4jOAZY0_3),.clk(gclk));
	jdff dff_A_fCpTHnQo3_0(.dout(w_G400_1[0]),.din(w_dff_A_fCpTHnQo3_0),.clk(gclk));
	jdff dff_A_QdSxXu2G1_0(.dout(w_dff_A_fCpTHnQo3_0),.din(w_dff_A_QdSxXu2G1_0),.clk(gclk));
	jdff dff_A_O4E25Dpd2_0(.dout(w_dff_A_QdSxXu2G1_0),.din(w_dff_A_O4E25Dpd2_0),.clk(gclk));
	jdff dff_A_kQSqkvHw5_0(.dout(w_dff_A_O4E25Dpd2_0),.din(w_dff_A_kQSqkvHw5_0),.clk(gclk));
	jdff dff_A_CjFOTSwv9_1(.dout(w_G400_1[1]),.din(w_dff_A_CjFOTSwv9_1),.clk(gclk));
	jdff dff_A_gPeqJYEJ5_1(.dout(w_dff_A_CjFOTSwv9_1),.din(w_dff_A_gPeqJYEJ5_1),.clk(gclk));
	jdff dff_A_lS1IRETb5_1(.dout(w_dff_A_gPeqJYEJ5_1),.din(w_dff_A_lS1IRETb5_1),.clk(gclk));
	jdff dff_B_61LdT2ER1_1(.din(n1526),.dout(w_dff_B_61LdT2ER1_1),.clk(gclk));
	jdff dff_A_AN3A2DOu0_0(.dout(w_G251_5[0]),.din(w_dff_A_AN3A2DOu0_0),.clk(gclk));
	jdff dff_A_AB26oXG68_0(.dout(w_G251_1[0]),.din(w_dff_A_AB26oXG68_0),.clk(gclk));
	jdff dff_A_Xcenn3811_2(.dout(w_G251_1[2]),.din(w_dff_A_Xcenn3811_2),.clk(gclk));
	jdff dff_A_ybWsuH9i4_1(.dout(w_G400_0[1]),.din(w_dff_A_ybWsuH9i4_1),.clk(gclk));
	jdff dff_A_RyuxyeXw5_1(.dout(w_dff_A_ybWsuH9i4_1),.din(w_dff_A_RyuxyeXw5_1),.clk(gclk));
	jdff dff_A_plKmlqta5_2(.dout(w_G400_0[2]),.din(w_dff_A_plKmlqta5_2),.clk(gclk));
	jdff dff_A_JfEtQdhX2_2(.dout(w_dff_A_plKmlqta5_2),.din(w_dff_A_JfEtQdhX2_2),.clk(gclk));
	jdff dff_A_LUYOThiy8_2(.dout(w_dff_A_JfEtQdhX2_2),.din(w_dff_A_LUYOThiy8_2),.clk(gclk));
	jdff dff_A_UIuZFd6I2_2(.dout(w_dff_A_LUYOThiy8_2),.din(w_dff_A_UIuZFd6I2_2),.clk(gclk));
	jdff dff_A_xejFgTk11_1(.dout(w_G265_1[1]),.din(w_dff_A_xejFgTk11_1),.clk(gclk));
	jdff dff_A_oVA4nxdI7_2(.dout(w_G265_0[2]),.din(w_dff_A_oVA4nxdI7_2),.clk(gclk));
	jdff dff_B_6LN4FPEo8_1(.din(n1516),.dout(w_dff_B_6LN4FPEo8_1),.clk(gclk));
	jdff dff_B_84LvMF523_1(.din(w_dff_B_6LN4FPEo8_1),.dout(w_dff_B_84LvMF523_1),.clk(gclk));
	jdff dff_A_SsgkcA2G8_0(.dout(w_G281_2[0]),.din(w_dff_A_SsgkcA2G8_0),.clk(gclk));
	jdff dff_A_9TwE1wRF8_1(.dout(w_n532_0[1]),.din(w_dff_A_9TwE1wRF8_1),.clk(gclk));
	jdff dff_A_IK6a6du75_1(.dout(w_dff_A_9TwE1wRF8_1),.din(w_dff_A_IK6a6du75_1),.clk(gclk));
	jdff dff_A_RObb8iE97_2(.dout(w_n532_0[2]),.din(w_dff_A_RObb8iE97_2),.clk(gclk));
	jdff dff_A_dGVpQ0Fx4_2(.dout(w_dff_A_RObb8iE97_2),.din(w_dff_A_dGVpQ0Fx4_2),.clk(gclk));
	jdff dff_B_bVA2yGk26_3(.din(n532),.dout(w_dff_B_bVA2yGk26_3),.clk(gclk));
	jdff dff_A_SHIZ7K8x2_0(.dout(w_G374_1[0]),.din(w_dff_A_SHIZ7K8x2_0),.clk(gclk));
	jdff dff_A_hbNxLAaW1_0(.dout(w_dff_A_SHIZ7K8x2_0),.din(w_dff_A_hbNxLAaW1_0),.clk(gclk));
	jdff dff_A_DeB1ZDg64_0(.dout(w_dff_A_hbNxLAaW1_0),.din(w_dff_A_DeB1ZDg64_0),.clk(gclk));
	jdff dff_A_NCvTwNFW0_0(.dout(w_dff_A_DeB1ZDg64_0),.din(w_dff_A_NCvTwNFW0_0),.clk(gclk));
	jdff dff_A_XIfLBDJu3_1(.dout(w_G374_1[1]),.din(w_dff_A_XIfLBDJu3_1),.clk(gclk));
	jdff dff_A_cggXNrML1_1(.dout(w_dff_A_XIfLBDJu3_1),.din(w_dff_A_cggXNrML1_1),.clk(gclk));
	jdff dff_A_ZHtEhEHW0_1(.dout(w_dff_A_cggXNrML1_1),.din(w_dff_A_ZHtEhEHW0_1),.clk(gclk));
	jdff dff_A_ooErNWfW8_1(.dout(w_G374_0[1]),.din(w_dff_A_ooErNWfW8_1),.clk(gclk));
	jdff dff_A_g1La7HFk9_1(.dout(w_dff_A_ooErNWfW8_1),.din(w_dff_A_g1La7HFk9_1),.clk(gclk));
	jdff dff_A_4pKE69fy7_1(.dout(w_dff_A_g1La7HFk9_1),.din(w_dff_A_4pKE69fy7_1),.clk(gclk));
	jdff dff_A_fmwFvSQN3_2(.dout(w_G374_0[2]),.din(w_dff_A_fmwFvSQN3_2),.clk(gclk));
	jdff dff_A_SDrAvg241_2(.dout(w_dff_A_fmwFvSQN3_2),.din(w_dff_A_SDrAvg241_2),.clk(gclk));
	jdff dff_A_N8zD4JvR7_2(.dout(w_dff_A_SDrAvg241_2),.din(w_dff_A_N8zD4JvR7_2),.clk(gclk));
	jdff dff_A_CHL3mOnJ1_2(.dout(w_dff_A_N8zD4JvR7_2),.din(w_dff_A_CHL3mOnJ1_2),.clk(gclk));
	jdff dff_A_n0anY7p45_2(.dout(w_G281_0[2]),.din(w_dff_A_n0anY7p45_2),.clk(gclk));
	jdff dff_A_SykPmhEG9_0(.dout(w_G242_1[0]),.din(w_dff_A_SykPmhEG9_0),.clk(gclk));
	jdff dff_A_dC6B2DkC2_1(.dout(w_G242_0[1]),.din(w_dff_A_dC6B2DkC2_1),.clk(gclk));
	jdff dff_A_ep1c18em2_2(.dout(w_G242_0[2]),.din(w_dff_A_ep1c18em2_2),.clk(gclk));
	jdff dff_B_Vrst2SN82_1(.din(n1507),.dout(w_dff_B_Vrst2SN82_1),.clk(gclk));
	jdff dff_B_Iy7RRtdp3_1(.din(w_dff_B_Vrst2SN82_1),.dout(w_dff_B_Iy7RRtdp3_1),.clk(gclk));
	jdff dff_A_HxChay362_0(.dout(w_G273_2[0]),.din(w_dff_A_HxChay362_0),.clk(gclk));
	jdff dff_A_ag2tn0BI5_1(.dout(w_G251_0[1]),.din(w_dff_A_ag2tn0BI5_1),.clk(gclk));
	jdff dff_A_wZ2op9mq3_2(.dout(w_G251_0[2]),.din(w_dff_A_wZ2op9mq3_2),.clk(gclk));
	jdff dff_A_7MBIRTJ58_1(.dout(w_n473_0[1]),.din(w_dff_A_7MBIRTJ58_1),.clk(gclk));
	jdff dff_A_eeLzT7dy9_1(.dout(w_dff_A_7MBIRTJ58_1),.din(w_dff_A_eeLzT7dy9_1),.clk(gclk));
	jdff dff_A_8KgFoi4m0_2(.dout(w_n473_0[2]),.din(w_dff_A_8KgFoi4m0_2),.clk(gclk));
	jdff dff_A_kK2bVqdC6_2(.dout(w_dff_A_8KgFoi4m0_2),.din(w_dff_A_kK2bVqdC6_2),.clk(gclk));
	jdff dff_B_t2bDAX2O6_3(.din(n473),.dout(w_dff_B_t2bDAX2O6_3),.clk(gclk));
	jdff dff_A_lXLSYaYB8_0(.dout(w_G411_2[0]),.din(w_dff_A_lXLSYaYB8_0),.clk(gclk));
	jdff dff_A_yK6I2eTU0_0(.dout(w_dff_A_lXLSYaYB8_0),.din(w_dff_A_yK6I2eTU0_0),.clk(gclk));
	jdff dff_A_vZS4jv8O6_0(.dout(w_dff_A_yK6I2eTU0_0),.din(w_dff_A_vZS4jv8O6_0),.clk(gclk));
	jdff dff_A_yiBZlk3W0_0(.dout(w_G411_0[0]),.din(w_dff_A_yiBZlk3W0_0),.clk(gclk));
	jdff dff_A_VtORDEFH0_0(.dout(w_dff_A_yiBZlk3W0_0),.din(w_dff_A_VtORDEFH0_0),.clk(gclk));
	jdff dff_A_IkiIFhRa1_0(.dout(w_dff_A_VtORDEFH0_0),.din(w_dff_A_IkiIFhRa1_0),.clk(gclk));
	jdff dff_A_BVx3UiRc1_0(.dout(w_dff_A_IkiIFhRa1_0),.din(w_dff_A_BVx3UiRc1_0),.clk(gclk));
	jdff dff_A_buwzuigq6_2(.dout(w_G411_0[2]),.din(w_dff_A_buwzuigq6_2),.clk(gclk));
	jdff dff_A_7JRegl3A8_2(.dout(w_dff_A_buwzuigq6_2),.din(w_dff_A_7JRegl3A8_2),.clk(gclk));
	jdff dff_A_lV1aM1ki1_2(.dout(w_dff_A_7JRegl3A8_2),.din(w_dff_A_lV1aM1ki1_2),.clk(gclk));
	jdff dff_A_XDgcLo2e7_1(.dout(w_G273_1[1]),.din(w_dff_A_XDgcLo2e7_1),.clk(gclk));
	jdff dff_A_Xnc6CWE06_2(.dout(w_G273_0[2]),.din(w_dff_A_Xnc6CWE06_2),.clk(gclk));
	jdff dff_A_A874vAr96_2(.dout(w_G248_3[2]),.din(w_dff_A_A874vAr96_2),.clk(gclk));
	jdff dff_A_QmFPONVY2_1(.dout(w_n749_4[1]),.din(w_dff_A_QmFPONVY2_1),.clk(gclk));
	jdff dff_A_rVnLMMcE5_1(.dout(w_dff_A_QmFPONVY2_1),.din(w_dff_A_rVnLMMcE5_1),.clk(gclk));
	jdff dff_A_wIENmvx61_1(.dout(w_dff_A_rVnLMMcE5_1),.din(w_dff_A_wIENmvx61_1),.clk(gclk));
	jdff dff_A_mJkvDEot9_1(.dout(w_dff_A_wIENmvx61_1),.din(w_dff_A_mJkvDEot9_1),.clk(gclk));
	jdff dff_A_LvXNHbYf9_1(.dout(w_dff_A_mJkvDEot9_1),.din(w_dff_A_LvXNHbYf9_1),.clk(gclk));
	jdff dff_A_8x1s1C3x8_1(.dout(w_dff_A_LvXNHbYf9_1),.din(w_dff_A_8x1s1C3x8_1),.clk(gclk));
	jdff dff_A_xusRBEtk2_1(.dout(w_dff_A_8x1s1C3x8_1),.din(w_dff_A_xusRBEtk2_1),.clk(gclk));
	jdff dff_A_1kC47ywc8_1(.dout(w_dff_A_xusRBEtk2_1),.din(w_dff_A_1kC47ywc8_1),.clk(gclk));
	jdff dff_A_SKrsXSo69_1(.dout(w_dff_A_1kC47ywc8_1),.din(w_dff_A_SKrsXSo69_1),.clk(gclk));
	jdff dff_A_aUNEpBAB7_1(.dout(w_dff_A_SKrsXSo69_1),.din(w_dff_A_aUNEpBAB7_1),.clk(gclk));
	jdff dff_A_TZBFGHtN2_1(.dout(w_dff_A_aUNEpBAB7_1),.din(w_dff_A_TZBFGHtN2_1),.clk(gclk));
	jdff dff_A_tyeBYNT06_1(.dout(w_dff_A_TZBFGHtN2_1),.din(w_dff_A_tyeBYNT06_1),.clk(gclk));
	jdff dff_A_GQEUk9Tg1_1(.dout(w_dff_A_tyeBYNT06_1),.din(w_dff_A_GQEUk9Tg1_1),.clk(gclk));
	jdff dff_A_SXDXHoG39_1(.dout(w_dff_A_GQEUk9Tg1_1),.din(w_dff_A_SXDXHoG39_1),.clk(gclk));
	jdff dff_A_K3YYi3n91_1(.dout(w_dff_A_SXDXHoG39_1),.din(w_dff_A_K3YYi3n91_1),.clk(gclk));
	jdff dff_A_8mp6hujI9_1(.dout(w_dff_A_K3YYi3n91_1),.din(w_dff_A_8mp6hujI9_1),.clk(gclk));
	jdff dff_A_18S8GhZa8_1(.dout(w_dff_A_8mp6hujI9_1),.din(w_dff_A_18S8GhZa8_1),.clk(gclk));
	jdff dff_A_FWMkj3kg1_2(.dout(w_n749_4[2]),.din(w_dff_A_FWMkj3kg1_2),.clk(gclk));
	jdff dff_A_8tnFSRF75_2(.dout(w_dff_A_FWMkj3kg1_2),.din(w_dff_A_8tnFSRF75_2),.clk(gclk));
	jdff dff_A_xA34DnvM7_2(.dout(w_dff_A_8tnFSRF75_2),.din(w_dff_A_xA34DnvM7_2),.clk(gclk));
	jdff dff_A_Jq8YDfEw5_2(.dout(w_dff_A_xA34DnvM7_2),.din(w_dff_A_Jq8YDfEw5_2),.clk(gclk));
	jdff dff_A_ldeQwlnR2_2(.dout(w_dff_A_Jq8YDfEw5_2),.din(w_dff_A_ldeQwlnR2_2),.clk(gclk));
	jdff dff_A_bM15YuWf9_2(.dout(w_dff_A_ldeQwlnR2_2),.din(w_dff_A_bM15YuWf9_2),.clk(gclk));
	jdff dff_A_Sfju9m4q5_2(.dout(w_dff_A_bM15YuWf9_2),.din(w_dff_A_Sfju9m4q5_2),.clk(gclk));
	jdff dff_A_JmgRWSyj3_2(.dout(w_dff_A_Sfju9m4q5_2),.din(w_dff_A_JmgRWSyj3_2),.clk(gclk));
	jdff dff_A_qL7zN0U73_1(.dout(w_n749_1[1]),.din(w_dff_A_qL7zN0U73_1),.clk(gclk));
	jdff dff_A_4SBju4m50_1(.dout(w_dff_A_qL7zN0U73_1),.din(w_dff_A_4SBju4m50_1),.clk(gclk));
	jdff dff_A_joNNIwb78_1(.dout(w_dff_A_4SBju4m50_1),.din(w_dff_A_joNNIwb78_1),.clk(gclk));
	jdff dff_A_gBzpWDv81_1(.dout(w_dff_A_joNNIwb78_1),.din(w_dff_A_gBzpWDv81_1),.clk(gclk));
	jdff dff_A_wG3p4WJa2_2(.dout(w_n749_1[2]),.din(w_dff_A_wG3p4WJa2_2),.clk(gclk));
	jdff dff_A_m8tm4q3K5_2(.dout(w_dff_A_wG3p4WJa2_2),.din(w_dff_A_m8tm4q3K5_2),.clk(gclk));
	jdff dff_A_nO0Ix8Q14_2(.dout(w_dff_A_m8tm4q3K5_2),.din(w_dff_A_nO0Ix8Q14_2),.clk(gclk));
	jdff dff_A_hfKCLmh88_2(.dout(w_dff_A_nO0Ix8Q14_2),.din(w_dff_A_hfKCLmh88_2),.clk(gclk));
	jdff dff_A_2jP08G0W9_1(.dout(w_n749_0[1]),.din(w_dff_A_2jP08G0W9_1),.clk(gclk));
	jdff dff_A_P7w9oMCp7_1(.dout(w_dff_A_2jP08G0W9_1),.din(w_dff_A_P7w9oMCp7_1),.clk(gclk));
	jdff dff_A_m1PNJ7gt1_2(.dout(w_n749_0[2]),.din(w_dff_A_m1PNJ7gt1_2),.clk(gclk));
	jdff dff_A_ulNocj2a9_2(.dout(w_dff_A_m1PNJ7gt1_2),.din(w_dff_A_ulNocj2a9_2),.clk(gclk));
	jdff dff_A_rpIbK18c5_2(.dout(w_dff_A_ulNocj2a9_2),.din(w_dff_A_rpIbK18c5_2),.clk(gclk));
	jdff dff_A_1PNMuPvk5_0(.dout(w_G4091_6[0]),.din(w_dff_A_1PNMuPvk5_0),.clk(gclk));
	jdff dff_A_L42a4hZQ2_0(.dout(w_dff_A_1PNMuPvk5_0),.din(w_dff_A_L42a4hZQ2_0),.clk(gclk));
	jdff dff_A_cgHyoynU1_0(.dout(w_dff_A_L42a4hZQ2_0),.din(w_dff_A_cgHyoynU1_0),.clk(gclk));
	jdff dff_A_hg5jQ5yC8_0(.dout(w_dff_A_cgHyoynU1_0),.din(w_dff_A_hg5jQ5yC8_0),.clk(gclk));
	jdff dff_A_abu6zKXv4_0(.dout(w_dff_A_hg5jQ5yC8_0),.din(w_dff_A_abu6zKXv4_0),.clk(gclk));
	jdff dff_A_lOz16oa14_0(.dout(w_G4091_1[0]),.din(w_dff_A_lOz16oa14_0),.clk(gclk));
	jdff dff_A_jKkpTKZP7_0(.dout(w_dff_A_lOz16oa14_0),.din(w_dff_A_jKkpTKZP7_0),.clk(gclk));
	jdff dff_A_fQgA9Y8k2_0(.dout(w_dff_A_jKkpTKZP7_0),.din(w_dff_A_fQgA9Y8k2_0),.clk(gclk));
	jdff dff_A_4bpCAS7U3_0(.dout(w_dff_A_fQgA9Y8k2_0),.din(w_dff_A_4bpCAS7U3_0),.clk(gclk));
	jdff dff_A_Ya2MDvDg5_0(.dout(w_dff_A_4bpCAS7U3_0),.din(w_dff_A_Ya2MDvDg5_0),.clk(gclk));
	jdff dff_A_ufVxp2va3_0(.dout(w_dff_A_Ya2MDvDg5_0),.din(w_dff_A_ufVxp2va3_0),.clk(gclk));
	jdff dff_A_acv2Moz75_0(.dout(w_dff_A_ufVxp2va3_0),.din(w_dff_A_acv2Moz75_0),.clk(gclk));
	jdff dff_A_wCjJ2qrj9_0(.dout(w_dff_A_acv2Moz75_0),.din(w_dff_A_wCjJ2qrj9_0),.clk(gclk));
	jdff dff_A_u33ZBVVq4_1(.dout(w_G4091_1[1]),.din(w_dff_A_u33ZBVVq4_1),.clk(gclk));
	jdff dff_A_7ygdSbNz5_1(.dout(w_dff_A_u33ZBVVq4_1),.din(w_dff_A_7ygdSbNz5_1),.clk(gclk));
	jdff dff_A_JjFCf3SU3_1(.dout(w_dff_A_7ygdSbNz5_1),.din(w_dff_A_JjFCf3SU3_1),.clk(gclk));
	jdff dff_A_4fSVkS468_1(.dout(w_dff_A_JjFCf3SU3_1),.din(w_dff_A_4fSVkS468_1),.clk(gclk));
	jdff dff_A_7ahHDM2d4_1(.dout(w_dff_A_4fSVkS468_1),.din(w_dff_A_7ahHDM2d4_1),.clk(gclk));
	jdff dff_A_f2bK6iJ99_1(.dout(w_dff_A_7ahHDM2d4_1),.din(w_dff_A_f2bK6iJ99_1),.clk(gclk));
	jdff dff_A_9pW0ku0l4_1(.dout(w_dff_A_f2bK6iJ99_1),.din(w_dff_A_9pW0ku0l4_1),.clk(gclk));
	jdff dff_A_SqUpkORK8_1(.dout(w_G4091_0[1]),.din(w_dff_A_SqUpkORK8_1),.clk(gclk));
	jdff dff_A_e0IOgCa68_1(.dout(w_dff_A_SqUpkORK8_1),.din(w_dff_A_e0IOgCa68_1),.clk(gclk));
	jdff dff_A_MHTbhHOa0_1(.dout(w_dff_A_e0IOgCa68_1),.din(w_dff_A_MHTbhHOa0_1),.clk(gclk));
	jdff dff_A_AoTVhK5r5_1(.dout(w_dff_A_MHTbhHOa0_1),.din(w_dff_A_AoTVhK5r5_1),.clk(gclk));
	jdff dff_A_QSj695yh7_1(.dout(w_dff_A_AoTVhK5r5_1),.din(w_dff_A_QSj695yh7_1),.clk(gclk));
	jdff dff_A_WF7BzBBr0_1(.dout(w_dff_A_QSj695yh7_1),.din(w_dff_A_WF7BzBBr0_1),.clk(gclk));
	jdff dff_A_15WhUGMC7_1(.dout(w_dff_A_WF7BzBBr0_1),.din(w_dff_A_15WhUGMC7_1),.clk(gclk));
	jdff dff_A_xBOjaOlL7_1(.dout(w_dff_A_15WhUGMC7_1),.din(w_dff_A_xBOjaOlL7_1),.clk(gclk));
	jdff dff_A_TkQwiBzn1_1(.dout(w_dff_A_xBOjaOlL7_1),.din(w_dff_A_TkQwiBzn1_1),.clk(gclk));
	jdff dff_A_L52SjsYQ4_1(.dout(w_dff_A_TkQwiBzn1_1),.din(w_dff_A_L52SjsYQ4_1),.clk(gclk));
	jdff dff_A_N2Pesr8z2_1(.dout(w_dff_A_L52SjsYQ4_1),.din(w_dff_A_N2Pesr8z2_1),.clk(gclk));
	jdff dff_A_XTCRzv6s1_1(.dout(w_dff_A_N2Pesr8z2_1),.din(w_dff_A_XTCRzv6s1_1),.clk(gclk));
	jdff dff_A_IS6nQ2ra3_1(.dout(w_dff_A_XTCRzv6s1_1),.din(w_dff_A_IS6nQ2ra3_1),.clk(gclk));
	jdff dff_A_JDbvVLrP1_2(.dout(w_G4091_0[2]),.din(w_dff_A_JDbvVLrP1_2),.clk(gclk));
	jdff dff_A_vnLBKfjy6_2(.dout(w_dff_A_JDbvVLrP1_2),.din(w_dff_A_vnLBKfjy6_2),.clk(gclk));
	jdff dff_A_T7N0C8DA8_2(.dout(w_dff_A_vnLBKfjy6_2),.din(w_dff_A_T7N0C8DA8_2),.clk(gclk));
	jdff dff_A_G1CLjoIg1_2(.dout(w_dff_A_T7N0C8DA8_2),.din(w_dff_A_G1CLjoIg1_2),.clk(gclk));
	jdff dff_A_86ZiklER1_2(.dout(w_dff_A_G1CLjoIg1_2),.din(w_dff_A_86ZiklER1_2),.clk(gclk));
	jdff dff_A_bX3uCpoF3_2(.dout(w_dff_A_86ZiklER1_2),.din(w_dff_A_bX3uCpoF3_2),.clk(gclk));
	jdff dff_A_w8qgU3tT1_2(.dout(w_dff_A_bX3uCpoF3_2),.din(w_dff_A_w8qgU3tT1_2),.clk(gclk));
	jdff dff_A_Bwnsjr1H9_2(.dout(w_dff_A_w8qgU3tT1_2),.din(w_dff_A_Bwnsjr1H9_2),.clk(gclk));
	jdff dff_A_La7wa7Bc6_2(.dout(w_G4092_3[2]),.din(w_dff_A_La7wa7Bc6_2),.clk(gclk));
	jdff dff_A_kHmuemLx6_2(.dout(w_dff_A_La7wa7Bc6_2),.din(w_dff_A_kHmuemLx6_2),.clk(gclk));
	jdff dff_A_ZJlPIZyA0_2(.dout(w_dff_A_kHmuemLx6_2),.din(w_dff_A_ZJlPIZyA0_2),.clk(gclk));
	jdff dff_A_Hk6Fst9G4_2(.dout(w_dff_A_ZJlPIZyA0_2),.din(w_dff_A_Hk6Fst9G4_2),.clk(gclk));
	jdff dff_A_sl1auLmP0_2(.dout(w_dff_A_Hk6Fst9G4_2),.din(w_dff_A_sl1auLmP0_2),.clk(gclk));
	jdff dff_A_diD9t98R6_2(.dout(w_dff_A_sl1auLmP0_2),.din(w_dff_A_diD9t98R6_2),.clk(gclk));
	jdff dff_A_Uyioptp97_2(.dout(w_dff_A_diD9t98R6_2),.din(w_dff_A_Uyioptp97_2),.clk(gclk));
	jdff dff_A_NYg3koBS9_2(.dout(w_dff_A_Uyioptp97_2),.din(w_dff_A_NYg3koBS9_2),.clk(gclk));
	jdff dff_A_bT4QangZ4_2(.dout(w_dff_A_NYg3koBS9_2),.din(w_dff_A_bT4QangZ4_2),.clk(gclk));
	jdff dff_A_m6hxobLJ9_2(.dout(w_dff_A_bT4QangZ4_2),.din(w_dff_A_m6hxobLJ9_2),.clk(gclk));
	jdff dff_A_mD33a3fK9_2(.dout(w_dff_A_m6hxobLJ9_2),.din(w_dff_A_mD33a3fK9_2),.clk(gclk));
	jdff dff_A_LibtmzMl2_2(.dout(w_dff_A_mD33a3fK9_2),.din(w_dff_A_LibtmzMl2_2),.clk(gclk));
	jdff dff_A_xyW0CzY38_2(.dout(w_dff_A_LibtmzMl2_2),.din(w_dff_A_xyW0CzY38_2),.clk(gclk));
	jdff dff_A_LdmW8x0z3_2(.dout(w_dff_A_xyW0CzY38_2),.din(w_dff_A_LdmW8x0z3_2),.clk(gclk));
	jdff dff_A_4TQbtAe49_2(.dout(w_dff_A_LdmW8x0z3_2),.din(w_dff_A_4TQbtAe49_2),.clk(gclk));
	jdff dff_A_4kapq13Z7_2(.dout(w_dff_A_4TQbtAe49_2),.din(w_dff_A_4kapq13Z7_2),.clk(gclk));
	jdff dff_A_038Cfig42_2(.dout(w_dff_A_4kapq13Z7_2),.din(w_dff_A_038Cfig42_2),.clk(gclk));
	jdff dff_A_dCrUWxxP8_2(.dout(w_dff_A_038Cfig42_2),.din(w_dff_A_dCrUWxxP8_2),.clk(gclk));
	jdff dff_A_GPjazOGn9_2(.dout(w_dff_A_dCrUWxxP8_2),.din(w_dff_A_GPjazOGn9_2),.clk(gclk));
	jdff dff_A_QiMycBOG7_2(.dout(w_dff_A_GPjazOGn9_2),.din(w_dff_A_QiMycBOG7_2),.clk(gclk));
	jdff dff_A_zpumRBPU4_1(.dout(w_G4092_0[1]),.din(w_dff_A_zpumRBPU4_1),.clk(gclk));
	jdff dff_A_tUyoymqM6_0(.dout(w_n1008_4[0]),.din(w_dff_A_tUyoymqM6_0),.clk(gclk));
	jdff dff_A_leokNJoC3_0(.dout(w_dff_A_tUyoymqM6_0),.din(w_dff_A_leokNJoC3_0),.clk(gclk));
	jdff dff_A_tMtAbBE44_0(.dout(w_dff_A_leokNJoC3_0),.din(w_dff_A_tMtAbBE44_0),.clk(gclk));
	jdff dff_A_2zTBnVFY3_0(.dout(w_dff_A_tMtAbBE44_0),.din(w_dff_A_2zTBnVFY3_0),.clk(gclk));
	jdff dff_A_RhfmZnRx8_0(.dout(w_dff_A_2zTBnVFY3_0),.din(w_dff_A_RhfmZnRx8_0),.clk(gclk));
	jdff dff_A_QsOMXu7T3_0(.dout(w_dff_A_RhfmZnRx8_0),.din(w_dff_A_QsOMXu7T3_0),.clk(gclk));
	jdff dff_A_cK0G9SQn9_0(.dout(w_dff_A_QsOMXu7T3_0),.din(w_dff_A_cK0G9SQn9_0),.clk(gclk));
	jdff dff_A_eKFeOMgR6_0(.dout(w_dff_A_cK0G9SQn9_0),.din(w_dff_A_eKFeOMgR6_0),.clk(gclk));
	jdff dff_A_CUrqyxfF2_0(.dout(w_dff_A_eKFeOMgR6_0),.din(w_dff_A_CUrqyxfF2_0),.clk(gclk));
	jdff dff_A_9gNR32xh3_0(.dout(w_dff_A_CUrqyxfF2_0),.din(w_dff_A_9gNR32xh3_0),.clk(gclk));
	jdff dff_A_um0V0JMZ4_0(.dout(w_dff_A_9gNR32xh3_0),.din(w_dff_A_um0V0JMZ4_0),.clk(gclk));
	jdff dff_A_u8FwNoFQ0_0(.dout(w_dff_A_um0V0JMZ4_0),.din(w_dff_A_u8FwNoFQ0_0),.clk(gclk));
	jdff dff_A_hsJNcbhz1_0(.dout(w_dff_A_u8FwNoFQ0_0),.din(w_dff_A_hsJNcbhz1_0),.clk(gclk));
	jdff dff_A_3qgpskuU3_0(.dout(w_dff_A_hsJNcbhz1_0),.din(w_dff_A_3qgpskuU3_0),.clk(gclk));
	jdff dff_A_AOPqFoq74_0(.dout(w_dff_A_3qgpskuU3_0),.din(w_dff_A_AOPqFoq74_0),.clk(gclk));
	jdff dff_A_S6zvsmWW5_2(.dout(w_n1008_4[2]),.din(w_dff_A_S6zvsmWW5_2),.clk(gclk));
	jdff dff_A_qhKHZmkp2_2(.dout(w_dff_A_S6zvsmWW5_2),.din(w_dff_A_qhKHZmkp2_2),.clk(gclk));
	jdff dff_A_R5E4t7Wd7_2(.dout(w_dff_A_qhKHZmkp2_2),.din(w_dff_A_R5E4t7Wd7_2),.clk(gclk));
	jdff dff_A_MGRmqino7_2(.dout(w_dff_A_R5E4t7Wd7_2),.din(w_dff_A_MGRmqino7_2),.clk(gclk));
	jdff dff_A_GcTVFFyF2_2(.dout(w_dff_A_MGRmqino7_2),.din(w_dff_A_GcTVFFyF2_2),.clk(gclk));
	jdff dff_A_Tq99ZMKc7_2(.dout(w_dff_A_GcTVFFyF2_2),.din(w_dff_A_Tq99ZMKc7_2),.clk(gclk));
	jdff dff_A_LJGOPbFW8_2(.dout(w_dff_A_Tq99ZMKc7_2),.din(w_dff_A_LJGOPbFW8_2),.clk(gclk));
	jdff dff_A_Lbz5AVLt8_2(.dout(w_dff_A_LJGOPbFW8_2),.din(w_dff_A_Lbz5AVLt8_2),.clk(gclk));
	jdff dff_A_4IbI5qIg8_2(.dout(w_dff_A_Lbz5AVLt8_2),.din(w_dff_A_4IbI5qIg8_2),.clk(gclk));
	jdff dff_A_kzzigXOh3_2(.dout(w_dff_A_4IbI5qIg8_2),.din(w_dff_A_kzzigXOh3_2),.clk(gclk));
	jdff dff_A_KvMsw2Wz1_1(.dout(w_n1008_1[1]),.din(w_dff_A_KvMsw2Wz1_1),.clk(gclk));
	jdff dff_A_ABsvNh0q2_1(.dout(w_dff_A_KvMsw2Wz1_1),.din(w_dff_A_ABsvNh0q2_1),.clk(gclk));
	jdff dff_A_9Ndf4BQT7_1(.dout(w_dff_A_ABsvNh0q2_1),.din(w_dff_A_9Ndf4BQT7_1),.clk(gclk));
	jdff dff_A_6yGIbgJk9_1(.dout(w_dff_A_9Ndf4BQT7_1),.din(w_dff_A_6yGIbgJk9_1),.clk(gclk));
	jdff dff_A_Bcdyjoly5_1(.dout(w_dff_A_6yGIbgJk9_1),.din(w_dff_A_Bcdyjoly5_1),.clk(gclk));
	jdff dff_A_jmAtlOM26_1(.dout(w_dff_A_Bcdyjoly5_1),.din(w_dff_A_jmAtlOM26_1),.clk(gclk));
	jdff dff_A_sZMLoobE0_1(.dout(w_dff_A_jmAtlOM26_1),.din(w_dff_A_sZMLoobE0_1),.clk(gclk));
	jdff dff_A_OniJDID48_1(.dout(w_dff_A_sZMLoobE0_1),.din(w_dff_A_OniJDID48_1),.clk(gclk));
	jdff dff_A_cKvAUkTb6_1(.dout(w_dff_A_OniJDID48_1),.din(w_dff_A_cKvAUkTb6_1),.clk(gclk));
	jdff dff_A_aX9q493N5_1(.dout(w_dff_A_cKvAUkTb6_1),.din(w_dff_A_aX9q493N5_1),.clk(gclk));
	jdff dff_A_hHg7xQvB7_1(.dout(w_dff_A_aX9q493N5_1),.din(w_dff_A_hHg7xQvB7_1),.clk(gclk));
	jdff dff_A_5H6tSYr47_1(.dout(w_dff_A_hHg7xQvB7_1),.din(w_dff_A_5H6tSYr47_1),.clk(gclk));
	jdff dff_A_xWr7UH5Q3_1(.dout(w_dff_A_5H6tSYr47_1),.din(w_dff_A_xWr7UH5Q3_1),.clk(gclk));
	jdff dff_A_59QCt9ds9_1(.dout(w_dff_A_xWr7UH5Q3_1),.din(w_dff_A_59QCt9ds9_1),.clk(gclk));
	jdff dff_A_BO0euw167_1(.dout(w_dff_A_59QCt9ds9_1),.din(w_dff_A_BO0euw167_1),.clk(gclk));
	jdff dff_A_vBtuAjRG5_1(.dout(w_dff_A_BO0euw167_1),.din(w_dff_A_vBtuAjRG5_1),.clk(gclk));
	jdff dff_A_fzWzgkzq4_1(.dout(w_dff_A_vBtuAjRG5_1),.din(w_dff_A_fzWzgkzq4_1),.clk(gclk));
	jdff dff_A_G1bb6GGQ8_1(.dout(w_dff_A_fzWzgkzq4_1),.din(w_dff_A_G1bb6GGQ8_1),.clk(gclk));
	jdff dff_A_hqnH5O3V7_1(.dout(w_dff_A_G1bb6GGQ8_1),.din(w_dff_A_hqnH5O3V7_1),.clk(gclk));
	jdff dff_A_XG3thPpc7_1(.dout(w_dff_A_hqnH5O3V7_1),.din(w_dff_A_XG3thPpc7_1),.clk(gclk));
	jdff dff_A_6m7zhnEg7_1(.dout(w_dff_A_XG3thPpc7_1),.din(w_dff_A_6m7zhnEg7_1),.clk(gclk));
	jdff dff_A_Q7TomOj72_2(.dout(w_n1008_1[2]),.din(w_dff_A_Q7TomOj72_2),.clk(gclk));
	jdff dff_A_CKW59UZj8_2(.dout(w_dff_A_Q7TomOj72_2),.din(w_dff_A_CKW59UZj8_2),.clk(gclk));
	jdff dff_A_rQ78NIQ30_2(.dout(w_dff_A_CKW59UZj8_2),.din(w_dff_A_rQ78NIQ30_2),.clk(gclk));
	jdff dff_A_ENqtAIKJ8_2(.dout(w_dff_A_rQ78NIQ30_2),.din(w_dff_A_ENqtAIKJ8_2),.clk(gclk));
	jdff dff_A_l6YA0Qq68_2(.dout(w_dff_A_ENqtAIKJ8_2),.din(w_dff_A_l6YA0Qq68_2),.clk(gclk));
	jdff dff_A_CgAlXiqs5_2(.dout(w_dff_A_l6YA0Qq68_2),.din(w_dff_A_CgAlXiqs5_2),.clk(gclk));
	jdff dff_A_CbNIir6s3_2(.dout(w_dff_A_CgAlXiqs5_2),.din(w_dff_A_CbNIir6s3_2),.clk(gclk));
	jdff dff_A_6cSLp0Vr2_2(.dout(w_dff_A_CbNIir6s3_2),.din(w_dff_A_6cSLp0Vr2_2),.clk(gclk));
	jdff dff_A_Gi49wAiq8_2(.dout(w_dff_A_6cSLp0Vr2_2),.din(w_dff_A_Gi49wAiq8_2),.clk(gclk));
	jdff dff_A_17q7hs9C8_2(.dout(w_dff_A_Gi49wAiq8_2),.din(w_dff_A_17q7hs9C8_2),.clk(gclk));
	jdff dff_A_P09OghY97_2(.dout(w_dff_A_17q7hs9C8_2),.din(w_dff_A_P09OghY97_2),.clk(gclk));
	jdff dff_A_CXDKtMOS7_2(.dout(w_dff_A_P09OghY97_2),.din(w_dff_A_CXDKtMOS7_2),.clk(gclk));
	jdff dff_A_HxlWNWNN4_2(.dout(w_dff_A_CXDKtMOS7_2),.din(w_dff_A_HxlWNWNN4_2),.clk(gclk));
	jdff dff_A_Gi4ay76v6_2(.dout(w_dff_A_HxlWNWNN4_2),.din(w_dff_A_Gi4ay76v6_2),.clk(gclk));
	jdff dff_A_73ILQWAl8_2(.dout(w_dff_A_Gi4ay76v6_2),.din(w_dff_A_73ILQWAl8_2),.clk(gclk));
	jdff dff_A_RaJ5jN9j2_2(.dout(w_dff_A_73ILQWAl8_2),.din(w_dff_A_RaJ5jN9j2_2),.clk(gclk));
	jdff dff_A_GdkOIG3a5_2(.dout(w_dff_A_RaJ5jN9j2_2),.din(w_dff_A_GdkOIG3a5_2),.clk(gclk));
	jdff dff_A_RVIUz57V5_2(.dout(w_dff_A_GdkOIG3a5_2),.din(w_dff_A_RVIUz57V5_2),.clk(gclk));
	jdff dff_A_jtmbmHih5_2(.dout(w_dff_A_RVIUz57V5_2),.din(w_dff_A_jtmbmHih5_2),.clk(gclk));
	jdff dff_A_qDgDVAEX0_2(.dout(w_dff_A_jtmbmHih5_2),.din(w_dff_A_qDgDVAEX0_2),.clk(gclk));
	jdff dff_A_n83Fldmf3_1(.dout(w_n1008_0[1]),.din(w_dff_A_n83Fldmf3_1),.clk(gclk));
	jdff dff_A_7SnZt01m0_1(.dout(w_dff_A_n83Fldmf3_1),.din(w_dff_A_7SnZt01m0_1),.clk(gclk));
	jdff dff_A_1r6QYUXj7_1(.dout(w_dff_A_7SnZt01m0_1),.din(w_dff_A_1r6QYUXj7_1),.clk(gclk));
	jdff dff_A_duODh0l13_1(.dout(w_dff_A_1r6QYUXj7_1),.din(w_dff_A_duODh0l13_1),.clk(gclk));
	jdff dff_A_Qx5Aw0pp3_1(.dout(w_dff_A_duODh0l13_1),.din(w_dff_A_Qx5Aw0pp3_1),.clk(gclk));
	jdff dff_A_S2krUQee6_1(.dout(w_dff_A_Qx5Aw0pp3_1),.din(w_dff_A_S2krUQee6_1),.clk(gclk));
	jdff dff_A_QHiPL11p7_1(.dout(w_dff_A_S2krUQee6_1),.din(w_dff_A_QHiPL11p7_1),.clk(gclk));
	jdff dff_A_AQobxrTk8_1(.dout(w_dff_A_QHiPL11p7_1),.din(w_dff_A_AQobxrTk8_1),.clk(gclk));
	jdff dff_A_mBpcS1Uq1_1(.dout(w_dff_A_AQobxrTk8_1),.din(w_dff_A_mBpcS1Uq1_1),.clk(gclk));
	jdff dff_A_wfoOlIGA8_1(.dout(w_dff_A_mBpcS1Uq1_1),.din(w_dff_A_wfoOlIGA8_1),.clk(gclk));
	jdff dff_A_N9vEfZbe5_1(.dout(w_dff_A_wfoOlIGA8_1),.din(w_dff_A_N9vEfZbe5_1),.clk(gclk));
	jdff dff_A_aRKS6wrS8_1(.dout(w_dff_A_N9vEfZbe5_1),.din(w_dff_A_aRKS6wrS8_1),.clk(gclk));
	jdff dff_A_iEHF2neW8_1(.dout(w_dff_A_aRKS6wrS8_1),.din(w_dff_A_iEHF2neW8_1),.clk(gclk));
	jdff dff_A_CZMZSsPr3_1(.dout(w_dff_A_iEHF2neW8_1),.din(w_dff_A_CZMZSsPr3_1),.clk(gclk));
	jdff dff_A_iJzWIcv50_1(.dout(w_dff_A_CZMZSsPr3_1),.din(w_dff_A_iJzWIcv50_1),.clk(gclk));
	jdff dff_A_GCavndNK0_1(.dout(w_dff_A_iJzWIcv50_1),.din(w_dff_A_GCavndNK0_1),.clk(gclk));
	jdff dff_A_cegOVNab9_1(.dout(w_dff_A_GCavndNK0_1),.din(w_dff_A_cegOVNab9_1),.clk(gclk));
	jdff dff_A_CjiMQbZv0_1(.dout(w_dff_A_cegOVNab9_1),.din(w_dff_A_CjiMQbZv0_1),.clk(gclk));
	jdff dff_A_EckuY08T7_2(.dout(w_n1008_0[2]),.din(w_dff_A_EckuY08T7_2),.clk(gclk));
	jdff dff_A_ZCFc1NNs1_2(.dout(w_dff_A_EckuY08T7_2),.din(w_dff_A_ZCFc1NNs1_2),.clk(gclk));
	jdff dff_A_QrxlWYS79_2(.dout(w_dff_A_ZCFc1NNs1_2),.din(w_dff_A_QrxlWYS79_2),.clk(gclk));
	jdff dff_A_paxpOmvk8_2(.dout(w_dff_A_QrxlWYS79_2),.din(w_dff_A_paxpOmvk8_2),.clk(gclk));
	jdff dff_A_8Xwink375_2(.dout(w_dff_A_paxpOmvk8_2),.din(w_dff_A_8Xwink375_2),.clk(gclk));
	jdff dff_A_wDNAb4JQ6_2(.dout(w_dff_A_8Xwink375_2),.din(w_dff_A_wDNAb4JQ6_2),.clk(gclk));
	jdff dff_A_X9qoxXSa8_2(.dout(w_dff_A_wDNAb4JQ6_2),.din(w_dff_A_X9qoxXSa8_2),.clk(gclk));
	jdff dff_A_MstGL8182_2(.dout(w_dff_A_X9qoxXSa8_2),.din(w_dff_A_MstGL8182_2),.clk(gclk));
	jdff dff_A_yFbPnCGk3_2(.dout(w_dff_A_MstGL8182_2),.din(w_dff_A_yFbPnCGk3_2),.clk(gclk));
	jdff dff_A_wo2T2kOp4_2(.dout(w_dff_A_yFbPnCGk3_2),.din(w_dff_A_wo2T2kOp4_2),.clk(gclk));
	jdff dff_A_R5JhrLx67_2(.dout(w_dff_A_wo2T2kOp4_2),.din(w_dff_A_R5JhrLx67_2),.clk(gclk));
	jdff dff_A_Kd1woLoV1_1(.dout(w_G1691_5[1]),.din(w_dff_A_Kd1woLoV1_1),.clk(gclk));
	jdff dff_A_TL5yoWNt6_1(.dout(w_dff_A_Kd1woLoV1_1),.din(w_dff_A_TL5yoWNt6_1),.clk(gclk));
	jdff dff_A_p71EIynG9_1(.dout(w_dff_A_TL5yoWNt6_1),.din(w_dff_A_p71EIynG9_1),.clk(gclk));
	jdff dff_A_9FGJ1ogt3_1(.dout(w_dff_A_p71EIynG9_1),.din(w_dff_A_9FGJ1ogt3_1),.clk(gclk));
	jdff dff_A_zyxbVRY35_1(.dout(w_dff_A_9FGJ1ogt3_1),.din(w_dff_A_zyxbVRY35_1),.clk(gclk));
	jdff dff_A_KNUNeVH45_1(.dout(w_dff_A_zyxbVRY35_1),.din(w_dff_A_KNUNeVH45_1),.clk(gclk));
	jdff dff_A_R4FSVQbU2_1(.dout(w_dff_A_KNUNeVH45_1),.din(w_dff_A_R4FSVQbU2_1),.clk(gclk));
	jdff dff_A_IbRR8L6h1_1(.dout(w_dff_A_R4FSVQbU2_1),.din(w_dff_A_IbRR8L6h1_1),.clk(gclk));
	jdff dff_A_3RYyMW4v3_1(.dout(w_dff_A_IbRR8L6h1_1),.din(w_dff_A_3RYyMW4v3_1),.clk(gclk));
	jdff dff_B_vTTmgdXH3_2(.din(n1698),.dout(w_dff_B_vTTmgdXH3_2),.clk(gclk));
	jdff dff_B_zUduTCUO7_2(.din(w_dff_B_vTTmgdXH3_2),.dout(w_dff_B_zUduTCUO7_2),.clk(gclk));
	jdff dff_A_WvYQrlL30_1(.dout(w_G1694_0[1]),.din(w_dff_A_WvYQrlL30_1),.clk(gclk));
	jdff dff_A_oxglm8aL4_1(.dout(w_dff_A_WvYQrlL30_1),.din(w_dff_A_oxglm8aL4_1),.clk(gclk));
	jdff dff_A_Uyau8rOH4_1(.dout(w_dff_A_oxglm8aL4_1),.din(w_dff_A_Uyau8rOH4_1),.clk(gclk));
	jdff dff_A_iUWZmf4S8_1(.dout(w_dff_A_Uyau8rOH4_1),.din(w_dff_A_iUWZmf4S8_1),.clk(gclk));
	jdff dff_A_IQOPX7Yd0_1(.dout(w_dff_A_iUWZmf4S8_1),.din(w_dff_A_IQOPX7Yd0_1),.clk(gclk));
	jdff dff_A_DSwvziJG4_1(.dout(w_dff_A_IQOPX7Yd0_1),.din(w_dff_A_DSwvziJG4_1),.clk(gclk));
	jdff dff_A_h0MFtjq21_1(.dout(w_dff_A_DSwvziJG4_1),.din(w_dff_A_h0MFtjq21_1),.clk(gclk));
	jdff dff_A_9yALk5ej3_1(.dout(w_dff_A_h0MFtjq21_1),.din(w_dff_A_9yALk5ej3_1),.clk(gclk));
	jdff dff_A_GwwbeOyA5_1(.dout(w_dff_A_9yALk5ej3_1),.din(w_dff_A_GwwbeOyA5_1),.clk(gclk));
	jdff dff_A_5rOVFMcB6_1(.dout(w_dff_A_GwwbeOyA5_1),.din(w_dff_A_5rOVFMcB6_1),.clk(gclk));
	jdff dff_A_p6lVwuwY1_1(.dout(w_dff_A_5rOVFMcB6_1),.din(w_dff_A_p6lVwuwY1_1),.clk(gclk));
	jdff dff_A_DaDP6A9e5_1(.dout(w_dff_A_p6lVwuwY1_1),.din(w_dff_A_DaDP6A9e5_1),.clk(gclk));
	jdff dff_A_hCyIYmwG4_1(.dout(w_dff_A_DaDP6A9e5_1),.din(w_dff_A_hCyIYmwG4_1),.clk(gclk));
	jdff dff_A_cEKVsM0h0_1(.dout(w_dff_A_hCyIYmwG4_1),.din(w_dff_A_cEKVsM0h0_1),.clk(gclk));
	jdff dff_A_dTd3rY9p2_1(.dout(w_dff_A_cEKVsM0h0_1),.din(w_dff_A_dTd3rY9p2_1),.clk(gclk));
	jdff dff_A_XQXoc7ej7_1(.dout(w_dff_A_dTd3rY9p2_1),.din(w_dff_A_XQXoc7ej7_1),.clk(gclk));
	jdff dff_A_FtERhn0I3_1(.dout(w_dff_A_XQXoc7ej7_1),.din(w_dff_A_FtERhn0I3_1),.clk(gclk));
	jdff dff_A_r7FVvO7W8_1(.dout(w_dff_A_FtERhn0I3_1),.din(w_dff_A_r7FVvO7W8_1),.clk(gclk));
	jdff dff_A_Prm6Og5L4_1(.dout(w_dff_A_r7FVvO7W8_1),.din(w_dff_A_Prm6Og5L4_1),.clk(gclk));
	jdff dff_A_hG80psQJ5_1(.dout(w_dff_A_Prm6Og5L4_1),.din(w_dff_A_hG80psQJ5_1),.clk(gclk));
	jdff dff_A_1jbPEVyJ8_1(.dout(w_dff_A_hG80psQJ5_1),.din(w_dff_A_1jbPEVyJ8_1),.clk(gclk));
	jdff dff_A_GUPV9wHc6_1(.dout(w_dff_A_1jbPEVyJ8_1),.din(w_dff_A_GUPV9wHc6_1),.clk(gclk));
	jdff dff_A_maasZoqd6_1(.dout(w_dff_A_GUPV9wHc6_1),.din(w_dff_A_maasZoqd6_1),.clk(gclk));
	jdff dff_A_iSQ5fhzh9_2(.dout(w_G1694_0[2]),.din(w_dff_A_iSQ5fhzh9_2),.clk(gclk));
	jdff dff_A_1zn0FW9l3_0(.dout(w_G1691_4[0]),.din(w_dff_A_1zn0FW9l3_0),.clk(gclk));
	jdff dff_A_sI0t8hvi3_0(.dout(w_dff_A_1zn0FW9l3_0),.din(w_dff_A_sI0t8hvi3_0),.clk(gclk));
	jdff dff_A_n8PzcbeJ9_0(.dout(w_dff_A_sI0t8hvi3_0),.din(w_dff_A_n8PzcbeJ9_0),.clk(gclk));
	jdff dff_A_faxlmhbC2_0(.dout(w_dff_A_n8PzcbeJ9_0),.din(w_dff_A_faxlmhbC2_0),.clk(gclk));
	jdff dff_A_D5259ui21_0(.dout(w_dff_A_faxlmhbC2_0),.din(w_dff_A_D5259ui21_0),.clk(gclk));
	jdff dff_A_kDYYvRzI8_0(.dout(w_dff_A_D5259ui21_0),.din(w_dff_A_kDYYvRzI8_0),.clk(gclk));
	jdff dff_A_4MzQigLh6_0(.dout(w_dff_A_kDYYvRzI8_0),.din(w_dff_A_4MzQigLh6_0),.clk(gclk));
	jdff dff_A_BF833sLg1_0(.dout(w_dff_A_4MzQigLh6_0),.din(w_dff_A_BF833sLg1_0),.clk(gclk));
	jdff dff_A_I2Ahqqac3_0(.dout(w_dff_A_BF833sLg1_0),.din(w_dff_A_I2Ahqqac3_0),.clk(gclk));
	jdff dff_A_wd0sOB1O0_0(.dout(w_dff_A_I2Ahqqac3_0),.din(w_dff_A_wd0sOB1O0_0),.clk(gclk));
	jdff dff_A_pnOQiB9S6_0(.dout(w_dff_A_wd0sOB1O0_0),.din(w_dff_A_pnOQiB9S6_0),.clk(gclk));
	jdff dff_A_ZjvMkhaB3_0(.dout(w_dff_A_pnOQiB9S6_0),.din(w_dff_A_ZjvMkhaB3_0),.clk(gclk));
	jdff dff_A_0ZUkinzQ9_0(.dout(w_dff_A_ZjvMkhaB3_0),.din(w_dff_A_0ZUkinzQ9_0),.clk(gclk));
	jdff dff_A_B8nvlZ5P7_0(.dout(w_dff_A_0ZUkinzQ9_0),.din(w_dff_A_B8nvlZ5P7_0),.clk(gclk));
	jdff dff_A_pValhosE3_1(.dout(w_G1691_4[1]),.din(w_dff_A_pValhosE3_1),.clk(gclk));
	jdff dff_A_qBUBGJnf6_1(.dout(w_dff_A_pValhosE3_1),.din(w_dff_A_qBUBGJnf6_1),.clk(gclk));
	jdff dff_A_WwMkvTmg2_1(.dout(w_dff_A_qBUBGJnf6_1),.din(w_dff_A_WwMkvTmg2_1),.clk(gclk));
	jdff dff_A_0tZkGy2R5_1(.dout(w_dff_A_WwMkvTmg2_1),.din(w_dff_A_0tZkGy2R5_1),.clk(gclk));
	jdff dff_A_Q457IU110_1(.dout(w_dff_A_0tZkGy2R5_1),.din(w_dff_A_Q457IU110_1),.clk(gclk));
	jdff dff_A_P1ZoAfh73_1(.dout(w_dff_A_Q457IU110_1),.din(w_dff_A_P1ZoAfh73_1),.clk(gclk));
	jdff dff_A_8Bs1N5t89_1(.dout(w_dff_A_P1ZoAfh73_1),.din(w_dff_A_8Bs1N5t89_1),.clk(gclk));
	jdff dff_A_D82Fgav34_1(.dout(w_dff_A_8Bs1N5t89_1),.din(w_dff_A_D82Fgav34_1),.clk(gclk));
	jdff dff_A_gaZOFjBe1_1(.dout(w_dff_A_D82Fgav34_1),.din(w_dff_A_gaZOFjBe1_1),.clk(gclk));
	jdff dff_A_EKrQaWfW0_1(.dout(w_dff_A_gaZOFjBe1_1),.din(w_dff_A_EKrQaWfW0_1),.clk(gclk));
	jdff dff_A_kX03BD1P6_1(.dout(w_dff_A_EKrQaWfW0_1),.din(w_dff_A_kX03BD1P6_1),.clk(gclk));
	jdff dff_A_UA9Pf4KL5_1(.dout(w_dff_A_kX03BD1P6_1),.din(w_dff_A_UA9Pf4KL5_1),.clk(gclk));
	jdff dff_A_zXcWcBZX6_1(.dout(w_dff_A_UA9Pf4KL5_1),.din(w_dff_A_zXcWcBZX6_1),.clk(gclk));
	jdff dff_A_tb6fQmuU0_1(.dout(w_dff_A_zXcWcBZX6_1),.din(w_dff_A_tb6fQmuU0_1),.clk(gclk));
	jdff dff_A_q0m21wPi2_1(.dout(w_dff_A_tb6fQmuU0_1),.din(w_dff_A_q0m21wPi2_1),.clk(gclk));
	jdff dff_A_QDiPIroo4_1(.dout(w_dff_A_q0m21wPi2_1),.din(w_dff_A_QDiPIroo4_1),.clk(gclk));
	jdff dff_A_PoiMz5Ac9_2(.dout(w_G1691_1[2]),.din(w_dff_A_PoiMz5Ac9_2),.clk(gclk));
	jdff dff_A_JNKQLG351_2(.dout(w_dff_A_PoiMz5Ac9_2),.din(w_dff_A_JNKQLG351_2),.clk(gclk));
	jdff dff_A_wXvvl4220_2(.dout(w_dff_A_JNKQLG351_2),.din(w_dff_A_wXvvl4220_2),.clk(gclk));
	jdff dff_A_eyUILGWx5_2(.dout(w_dff_A_wXvvl4220_2),.din(w_dff_A_eyUILGWx5_2),.clk(gclk));
	jdff dff_A_ciRmbqC69_2(.dout(w_dff_A_eyUILGWx5_2),.din(w_dff_A_ciRmbqC69_2),.clk(gclk));
	jdff dff_A_toGPZZx61_2(.dout(w_dff_A_ciRmbqC69_2),.din(w_dff_A_toGPZZx61_2),.clk(gclk));
	jdff dff_A_8BAYJSgG8_2(.dout(w_dff_A_toGPZZx61_2),.din(w_dff_A_8BAYJSgG8_2),.clk(gclk));
	jdff dff_A_0zVSTN7V4_2(.dout(w_dff_A_8BAYJSgG8_2),.din(w_dff_A_0zVSTN7V4_2),.clk(gclk));
	jdff dff_A_ZjiWu6AX5_2(.dout(w_dff_A_0zVSTN7V4_2),.din(w_dff_A_ZjiWu6AX5_2),.clk(gclk));
	jdff dff_A_BCMNKDZn4_2(.dout(w_dff_A_ZjiWu6AX5_2),.din(w_dff_A_BCMNKDZn4_2),.clk(gclk));
	jdff dff_A_y9X4lfj04_2(.dout(w_dff_A_BCMNKDZn4_2),.din(w_dff_A_y9X4lfj04_2),.clk(gclk));
	jdff dff_A_oF5qS0QM0_2(.dout(w_dff_A_y9X4lfj04_2),.din(w_dff_A_oF5qS0QM0_2),.clk(gclk));
	jdff dff_A_MJ2fc6d40_2(.dout(w_dff_A_oF5qS0QM0_2),.din(w_dff_A_MJ2fc6d40_2),.clk(gclk));
	jdff dff_A_QZHUGb6u4_2(.dout(w_dff_A_MJ2fc6d40_2),.din(w_dff_A_QZHUGb6u4_2),.clk(gclk));
	jdff dff_A_V1Ok5GXE1_2(.dout(w_dff_A_QZHUGb6u4_2),.din(w_dff_A_V1Ok5GXE1_2),.clk(gclk));
	jdff dff_A_upmf6GZf8_2(.dout(w_dff_A_V1Ok5GXE1_2),.din(w_dff_A_upmf6GZf8_2),.clk(gclk));
	jdff dff_A_cG5jVoDi3_2(.dout(w_dff_A_upmf6GZf8_2),.din(w_dff_A_cG5jVoDi3_2),.clk(gclk));
	jdff dff_A_JjpVs2l14_2(.dout(w_dff_A_cG5jVoDi3_2),.din(w_dff_A_JjpVs2l14_2),.clk(gclk));
	jdff dff_A_0Zydq1sV2_2(.dout(w_dff_A_JjpVs2l14_2),.din(w_dff_A_0Zydq1sV2_2),.clk(gclk));
	jdff dff_A_3bmgABKA0_2(.dout(w_dff_A_0Zydq1sV2_2),.din(w_dff_A_3bmgABKA0_2),.clk(gclk));
	jdff dff_A_7LvYdvXl2_2(.dout(w_dff_A_3bmgABKA0_2),.din(w_dff_A_7LvYdvXl2_2),.clk(gclk));
	jdff dff_A_eJwSTwYZ2_2(.dout(w_dff_A_7LvYdvXl2_2),.din(w_dff_A_eJwSTwYZ2_2),.clk(gclk));
	jdff dff_A_UKG6o2On8_1(.dout(w_G1691_0[1]),.din(w_dff_A_UKG6o2On8_1),.clk(gclk));
	jdff dff_A_FLatmz6y4_1(.dout(w_dff_A_UKG6o2On8_1),.din(w_dff_A_FLatmz6y4_1),.clk(gclk));
	jdff dff_A_Ofo6YQ9j5_1(.dout(w_dff_A_FLatmz6y4_1),.din(w_dff_A_Ofo6YQ9j5_1),.clk(gclk));
	jdff dff_A_S7zuDv7J9_1(.dout(w_dff_A_Ofo6YQ9j5_1),.din(w_dff_A_S7zuDv7J9_1),.clk(gclk));
	jdff dff_A_2MDohQwi1_1(.dout(w_dff_A_S7zuDv7J9_1),.din(w_dff_A_2MDohQwi1_1),.clk(gclk));
	jdff dff_A_OhKwQuUF8_1(.dout(w_dff_A_2MDohQwi1_1),.din(w_dff_A_OhKwQuUF8_1),.clk(gclk));
	jdff dff_A_RXfymimW9_1(.dout(w_dff_A_OhKwQuUF8_1),.din(w_dff_A_RXfymimW9_1),.clk(gclk));
	jdff dff_A_6P6OGPYf9_1(.dout(w_dff_A_RXfymimW9_1),.din(w_dff_A_6P6OGPYf9_1),.clk(gclk));
	jdff dff_A_kcbGcgpW1_1(.dout(w_dff_A_6P6OGPYf9_1),.din(w_dff_A_kcbGcgpW1_1),.clk(gclk));
	jdff dff_A_eP5SoSc09_1(.dout(w_dff_A_kcbGcgpW1_1),.din(w_dff_A_eP5SoSc09_1),.clk(gclk));
	jdff dff_A_9mEPYqNs0_1(.dout(w_dff_A_eP5SoSc09_1),.din(w_dff_A_9mEPYqNs0_1),.clk(gclk));
	jdff dff_A_Oqh6KgFz0_1(.dout(w_dff_A_9mEPYqNs0_1),.din(w_dff_A_Oqh6KgFz0_1),.clk(gclk));
	jdff dff_A_x0n7M0CU1_1(.dout(w_dff_A_Oqh6KgFz0_1),.din(w_dff_A_x0n7M0CU1_1),.clk(gclk));
	jdff dff_A_VI9suVM74_1(.dout(w_dff_A_x0n7M0CU1_1),.din(w_dff_A_VI9suVM74_1),.clk(gclk));
	jdff dff_A_qhvw2oD49_1(.dout(w_dff_A_VI9suVM74_1),.din(w_dff_A_qhvw2oD49_1),.clk(gclk));
	jdff dff_A_uRKIXgyP0_1(.dout(w_dff_A_qhvw2oD49_1),.din(w_dff_A_uRKIXgyP0_1),.clk(gclk));
	jdff dff_A_1CLzg2rg9_1(.dout(w_dff_A_uRKIXgyP0_1),.din(w_dff_A_1CLzg2rg9_1),.clk(gclk));
	jdff dff_A_DdnqrwI38_1(.dout(w_dff_A_1CLzg2rg9_1),.din(w_dff_A_DdnqrwI38_1),.clk(gclk));
	jdff dff_A_cCDNMOeN8_1(.dout(w_dff_A_DdnqrwI38_1),.din(w_dff_A_cCDNMOeN8_1),.clk(gclk));
	jdff dff_A_ctaA7Ga85_2(.dout(w_G1691_0[2]),.din(w_dff_A_ctaA7Ga85_2),.clk(gclk));
	jdff dff_A_pvCPnmrF3_2(.dout(w_dff_A_ctaA7Ga85_2),.din(w_dff_A_pvCPnmrF3_2),.clk(gclk));
	jdff dff_A_FJqnepso1_2(.dout(w_dff_A_pvCPnmrF3_2),.din(w_dff_A_FJqnepso1_2),.clk(gclk));
	jdff dff_A_ZXqA7kjK0_2(.dout(w_dff_A_FJqnepso1_2),.din(w_dff_A_ZXqA7kjK0_2),.clk(gclk));
	jdff dff_A_Sjj8KgGM0_2(.dout(w_dff_A_ZXqA7kjK0_2),.din(w_dff_A_Sjj8KgGM0_2),.clk(gclk));
	jdff dff_A_HVV6sDmd5_2(.dout(w_dff_A_Sjj8KgGM0_2),.din(w_dff_A_HVV6sDmd5_2),.clk(gclk));
	jdff dff_A_nGmCrTM09_2(.dout(w_dff_A_HVV6sDmd5_2),.din(w_dff_A_nGmCrTM09_2),.clk(gclk));
	jdff dff_A_iypFZ4u34_2(.dout(w_dff_A_nGmCrTM09_2),.din(w_dff_A_iypFZ4u34_2),.clk(gclk));
	jdff dff_A_AF0T8pOP5_2(.dout(w_dff_A_iypFZ4u34_2),.din(w_dff_A_AF0T8pOP5_2),.clk(gclk));
	jdff dff_A_tZzpomHH7_2(.dout(w_dff_A_AF0T8pOP5_2),.din(w_dff_A_tZzpomHH7_2),.clk(gclk));
	jdff dff_A_9twEvPVT9_2(.dout(w_dff_A_tZzpomHH7_2),.din(w_dff_A_9twEvPVT9_2),.clk(gclk));
	jdff dff_A_RuPJy40b7_2(.dout(w_dff_A_9twEvPVT9_2),.din(w_dff_A_RuPJy40b7_2),.clk(gclk));
	jdff dff_A_23j1qrul6_2(.dout(w_dff_A_RuPJy40b7_2),.din(w_dff_A_23j1qrul6_2),.clk(gclk));
	jdff dff_B_2yHgIPs07_2(.din(n1695),.dout(w_dff_B_2yHgIPs07_2),.clk(gclk));
	jdff dff_B_9sooeByT0_2(.din(n1694),.dout(w_dff_B_9sooeByT0_2),.clk(gclk));
	jdff dff_B_2NtVvx7U7_2(.din(w_dff_B_9sooeByT0_2),.dout(w_dff_B_2NtVvx7U7_2),.clk(gclk));
	jdff dff_B_ZxvMcgsl9_2(.din(w_dff_B_2NtVvx7U7_2),.dout(w_dff_B_ZxvMcgsl9_2),.clk(gclk));
	jdff dff_B_66RmEDxR7_2(.din(w_dff_B_ZxvMcgsl9_2),.dout(w_dff_B_66RmEDxR7_2),.clk(gclk));
	jdff dff_B_2z3YppNc4_2(.din(w_dff_B_66RmEDxR7_2),.dout(w_dff_B_2z3YppNc4_2),.clk(gclk));
	jdff dff_B_7hBvI9OX1_2(.din(w_dff_B_2z3YppNc4_2),.dout(w_dff_B_7hBvI9OX1_2),.clk(gclk));
	jdff dff_B_snZ0o9Go0_2(.din(w_dff_B_7hBvI9OX1_2),.dout(w_dff_B_snZ0o9Go0_2),.clk(gclk));
	jdff dff_B_Utc8l5Ed5_2(.din(w_dff_B_snZ0o9Go0_2),.dout(w_dff_B_Utc8l5Ed5_2),.clk(gclk));
	jdff dff_B_NF5C1Nn97_2(.din(w_dff_B_Utc8l5Ed5_2),.dout(w_dff_B_NF5C1Nn97_2),.clk(gclk));
	jdff dff_B_T2HUfdDr4_2(.din(w_dff_B_NF5C1Nn97_2),.dout(w_dff_B_T2HUfdDr4_2),.clk(gclk));
	jdff dff_B_nikbwyKM3_2(.din(w_dff_B_T2HUfdDr4_2),.dout(w_dff_B_nikbwyKM3_2),.clk(gclk));
	jdff dff_B_Rep7RpYD2_2(.din(w_dff_B_nikbwyKM3_2),.dout(w_dff_B_Rep7RpYD2_2),.clk(gclk));
	jdff dff_B_mPJEABN45_2(.din(w_dff_B_Rep7RpYD2_2),.dout(w_dff_B_mPJEABN45_2),.clk(gclk));
	jdff dff_B_28kfokIz3_2(.din(w_dff_B_mPJEABN45_2),.dout(w_dff_B_28kfokIz3_2),.clk(gclk));
	jdff dff_B_HT9O9xGS3_2(.din(w_dff_B_28kfokIz3_2),.dout(w_dff_B_HT9O9xGS3_2),.clk(gclk));
	jdff dff_B_Bl5IV9hL1_2(.din(w_dff_B_HT9O9xGS3_2),.dout(w_dff_B_Bl5IV9hL1_2),.clk(gclk));
	jdff dff_B_exsyAiCG6_2(.din(w_dff_B_Bl5IV9hL1_2),.dout(w_dff_B_exsyAiCG6_2),.clk(gclk));
	jdff dff_B_sgULzQrm4_2(.din(w_dff_B_exsyAiCG6_2),.dout(w_dff_B_sgULzQrm4_2),.clk(gclk));
	jdff dff_B_wkl94Ujk6_2(.din(w_dff_B_sgULzQrm4_2),.dout(w_dff_B_wkl94Ujk6_2),.clk(gclk));
	jdff dff_B_uJwmzMDo1_2(.din(w_dff_B_wkl94Ujk6_2),.dout(w_dff_B_uJwmzMDo1_2),.clk(gclk));
	jdff dff_B_u6C3mbq99_2(.din(w_dff_B_uJwmzMDo1_2),.dout(w_dff_B_u6C3mbq99_2),.clk(gclk));
	jdff dff_B_X2NDuRZT2_2(.din(w_dff_B_u6C3mbq99_2),.dout(w_dff_B_X2NDuRZT2_2),.clk(gclk));
	jdff dff_B_Tz5UtP4x1_2(.din(w_dff_B_X2NDuRZT2_2),.dout(w_dff_B_Tz5UtP4x1_2),.clk(gclk));
	jdff dff_B_gBJalVQ91_2(.din(w_dff_B_Tz5UtP4x1_2),.dout(w_dff_B_gBJalVQ91_2),.clk(gclk));
	jdff dff_B_WbwCPc6t8_2(.din(w_dff_B_gBJalVQ91_2),.dout(w_dff_B_WbwCPc6t8_2),.clk(gclk));
	jdff dff_B_ComM23HU8_2(.din(w_dff_B_WbwCPc6t8_2),.dout(w_dff_B_ComM23HU8_2),.clk(gclk));
	jdff dff_A_rx02fJcA4_2(.dout(w_G137_3[2]),.din(w_dff_A_rx02fJcA4_2),.clk(gclk));
	jdff dff_A_IjALdprk9_2(.dout(w_dff_A_rx02fJcA4_2),.din(w_dff_A_IjALdprk9_2),.clk(gclk));
	jdff dff_A_Qh7WqTdm3_2(.dout(w_dff_A_IjALdprk9_2),.din(w_dff_A_Qh7WqTdm3_2),.clk(gclk));
	jdff dff_A_sAIzt9Om2_2(.dout(w_dff_A_Qh7WqTdm3_2),.din(w_dff_A_sAIzt9Om2_2),.clk(gclk));
	jdff dff_A_zjPgcxCe5_2(.dout(w_dff_A_sAIzt9Om2_2),.din(w_dff_A_zjPgcxCe5_2),.clk(gclk));
	jdff dff_A_EK5u4MGd4_2(.dout(w_dff_A_zjPgcxCe5_2),.din(w_dff_A_EK5u4MGd4_2),.clk(gclk));
	jdff dff_A_Qy0P7KGC3_2(.dout(w_dff_A_EK5u4MGd4_2),.din(w_dff_A_Qy0P7KGC3_2),.clk(gclk));
	jdff dff_A_NpUXdRDf9_2(.dout(w_dff_A_Qy0P7KGC3_2),.din(w_dff_A_NpUXdRDf9_2),.clk(gclk));
	jdff dff_A_U9QQQQ9q7_2(.dout(w_dff_A_NpUXdRDf9_2),.din(w_dff_A_U9QQQQ9q7_2),.clk(gclk));
	jdff dff_A_o09nx3OJ9_2(.dout(w_dff_A_U9QQQQ9q7_2),.din(w_dff_A_o09nx3OJ9_2),.clk(gclk));
	jdff dff_A_y4lPRZbD2_2(.dout(w_dff_A_o09nx3OJ9_2),.din(w_dff_A_y4lPRZbD2_2),.clk(gclk));
	jdff dff_A_hSUd2tAn6_2(.dout(w_dff_A_y4lPRZbD2_2),.din(w_dff_A_hSUd2tAn6_2),.clk(gclk));
	jdff dff_A_VwQ7Q4MO3_2(.dout(w_dff_A_hSUd2tAn6_2),.din(w_dff_A_VwQ7Q4MO3_2),.clk(gclk));
	jdff dff_A_dhOvOXiJ7_2(.dout(w_dff_A_VwQ7Q4MO3_2),.din(w_dff_A_dhOvOXiJ7_2),.clk(gclk));
	jdff dff_A_k9OrDIyn6_2(.dout(w_dff_A_dhOvOXiJ7_2),.din(w_dff_A_k9OrDIyn6_2),.clk(gclk));
	jdff dff_A_lz2J2iFq4_2(.dout(w_dff_A_k9OrDIyn6_2),.din(w_dff_A_lz2J2iFq4_2),.clk(gclk));
	jdff dff_A_X8bcnnpD2_2(.dout(w_dff_A_lz2J2iFq4_2),.din(w_dff_A_X8bcnnpD2_2),.clk(gclk));
	jdff dff_A_tgqHDiAc2_2(.dout(w_dff_A_X8bcnnpD2_2),.din(w_dff_A_tgqHDiAc2_2),.clk(gclk));
	jdff dff_A_wWrsynmd1_2(.dout(w_dff_A_tgqHDiAc2_2),.din(w_dff_A_wWrsynmd1_2),.clk(gclk));
	jdff dff_A_isLajwhg1_2(.dout(w_dff_A_wWrsynmd1_2),.din(w_dff_A_isLajwhg1_2),.clk(gclk));
	jdff dff_A_FyHF9BLE4_2(.dout(w_dff_A_isLajwhg1_2),.din(w_dff_A_FyHF9BLE4_2),.clk(gclk));
	jdff dff_A_xK66aRus4_2(.dout(w_dff_A_FyHF9BLE4_2),.din(w_dff_A_xK66aRus4_2),.clk(gclk));
	jdff dff_A_x6nZdfzX3_2(.dout(w_dff_A_xK66aRus4_2),.din(w_dff_A_x6nZdfzX3_2),.clk(gclk));
	jdff dff_A_sNwTwktN2_2(.dout(w_dff_A_x6nZdfzX3_2),.din(w_dff_A_sNwTwktN2_2),.clk(gclk));
	jdff dff_A_A8BELJ2X6_0(.dout(w_G137_0[0]),.din(w_dff_A_A8BELJ2X6_0),.clk(gclk));
	jdff dff_A_zKiWamOe3_0(.dout(w_dff_A_A8BELJ2X6_0),.din(w_dff_A_zKiWamOe3_0),.clk(gclk));
	jdff dff_A_O5YFOKGR7_0(.dout(w_dff_A_zKiWamOe3_0),.din(w_dff_A_O5YFOKGR7_0),.clk(gclk));
	jdff dff_A_mtujyeSZ6_0(.dout(w_dff_A_O5YFOKGR7_0),.din(w_dff_A_mtujyeSZ6_0),.clk(gclk));
	jdff dff_A_zW829UXt3_0(.dout(w_dff_A_mtujyeSZ6_0),.din(w_dff_A_zW829UXt3_0),.clk(gclk));
	jdff dff_A_GDujKmWD5_0(.dout(w_dff_A_zW829UXt3_0),.din(w_dff_A_GDujKmWD5_0),.clk(gclk));
	jdff dff_A_wY8J6Gb31_0(.dout(w_dff_A_GDujKmWD5_0),.din(w_dff_A_wY8J6Gb31_0),.clk(gclk));
	jdff dff_A_7KZUvj8u0_0(.dout(w_dff_A_wY8J6Gb31_0),.din(w_dff_A_7KZUvj8u0_0),.clk(gclk));
	jdff dff_A_BeQqMVqK0_0(.dout(w_dff_A_7KZUvj8u0_0),.din(w_dff_A_BeQqMVqK0_0),.clk(gclk));
	jdff dff_A_AfrDHYLP4_0(.dout(w_dff_A_BeQqMVqK0_0),.din(w_dff_A_AfrDHYLP4_0),.clk(gclk));
	jdff dff_A_JEuwzS7x6_0(.dout(w_dff_A_AfrDHYLP4_0),.din(w_dff_A_JEuwzS7x6_0),.clk(gclk));
	jdff dff_A_qjSc4dUF4_0(.dout(w_dff_A_JEuwzS7x6_0),.din(w_dff_A_qjSc4dUF4_0),.clk(gclk));
	jdff dff_A_151P5m3h8_0(.dout(w_dff_A_qjSc4dUF4_0),.din(w_dff_A_151P5m3h8_0),.clk(gclk));
	jdff dff_A_7k2fERvA4_0(.dout(w_dff_A_151P5m3h8_0),.din(w_dff_A_7k2fERvA4_0),.clk(gclk));
	jdff dff_A_Z1q1Mqem2_0(.dout(w_dff_A_7k2fERvA4_0),.din(w_dff_A_Z1q1Mqem2_0),.clk(gclk));
	jdff dff_A_DRfSNG8T2_0(.dout(w_dff_A_Z1q1Mqem2_0),.din(w_dff_A_DRfSNG8T2_0),.clk(gclk));
	jdff dff_A_kBbJ84pR7_0(.dout(w_dff_A_DRfSNG8T2_0),.din(w_dff_A_kBbJ84pR7_0),.clk(gclk));
	jdff dff_A_xRuhdLMe1_1(.dout(w_G137_0[1]),.din(w_dff_A_xRuhdLMe1_1),.clk(gclk));
	jdff dff_A_aLpvP9LV1_1(.dout(w_dff_A_xRuhdLMe1_1),.din(w_dff_A_aLpvP9LV1_1),.clk(gclk));
	jdff dff_A_F0se0r0E0_1(.dout(w_dff_A_aLpvP9LV1_1),.din(w_dff_A_F0se0r0E0_1),.clk(gclk));
	jdff dff_A_Csk56dO18_1(.dout(w_dff_A_F0se0r0E0_1),.din(w_dff_A_Csk56dO18_1),.clk(gclk));
	jdff dff_A_troJ6RLa5_1(.dout(w_dff_A_Csk56dO18_1),.din(w_dff_A_troJ6RLa5_1),.clk(gclk));
	jdff dff_A_9fKkWfc92_1(.dout(w_dff_A_troJ6RLa5_1),.din(w_dff_A_9fKkWfc92_1),.clk(gclk));
	jdff dff_A_26Jm6bKv9_1(.dout(w_dff_A_9fKkWfc92_1),.din(w_dff_A_26Jm6bKv9_1),.clk(gclk));
	jdff dff_A_EsurVI7l9_1(.dout(w_dff_A_26Jm6bKv9_1),.din(w_dff_A_EsurVI7l9_1),.clk(gclk));
	jdff dff_A_zkC8SsFR6_1(.dout(w_dff_A_EsurVI7l9_1),.din(w_dff_A_zkC8SsFR6_1),.clk(gclk));
	jdff dff_A_1BWYzmuQ1_1(.dout(w_dff_A_zkC8SsFR6_1),.din(w_dff_A_1BWYzmuQ1_1),.clk(gclk));
	jdff dff_A_UN5DTPSc9_1(.dout(w_dff_A_1BWYzmuQ1_1),.din(w_dff_A_UN5DTPSc9_1),.clk(gclk));
	jdff dff_A_NW14Cpb48_1(.dout(w_dff_A_UN5DTPSc9_1),.din(w_dff_A_NW14Cpb48_1),.clk(gclk));
	jdff dff_A_XdinJ2ua1_1(.dout(w_dff_A_NW14Cpb48_1),.din(w_dff_A_XdinJ2ua1_1),.clk(gclk));
	jdff dff_A_596UulZT0_1(.dout(w_dff_A_XdinJ2ua1_1),.din(w_dff_A_596UulZT0_1),.clk(gclk));
	jdff dff_A_4BTpAQXa4_1(.dout(w_dff_A_596UulZT0_1),.din(w_dff_A_4BTpAQXa4_1),.clk(gclk));
	jdff dff_A_rVLNTSTJ6_1(.dout(w_dff_A_5W8qnzvR0_0),.din(w_dff_A_rVLNTSTJ6_1),.clk(gclk));
	jdff dff_A_5W8qnzvR0_0(.dout(w_dff_A_DhSCiVOk5_0),.din(w_dff_A_5W8qnzvR0_0),.clk(gclk));
	jdff dff_A_DhSCiVOk5_0(.dout(w_dff_A_ZqmDPFpX7_0),.din(w_dff_A_DhSCiVOk5_0),.clk(gclk));
	jdff dff_A_ZqmDPFpX7_0(.dout(w_dff_A_OlwTOGBO1_0),.din(w_dff_A_ZqmDPFpX7_0),.clk(gclk));
	jdff dff_A_OlwTOGBO1_0(.dout(w_dff_A_3xkKmlGw6_0),.din(w_dff_A_OlwTOGBO1_0),.clk(gclk));
	jdff dff_A_3xkKmlGw6_0(.dout(w_dff_A_4Z7Y37RQ6_0),.din(w_dff_A_3xkKmlGw6_0),.clk(gclk));
	jdff dff_A_4Z7Y37RQ6_0(.dout(w_dff_A_2vtPyoSX7_0),.din(w_dff_A_4Z7Y37RQ6_0),.clk(gclk));
	jdff dff_A_2vtPyoSX7_0(.dout(w_dff_A_PIzinJ1w3_0),.din(w_dff_A_2vtPyoSX7_0),.clk(gclk));
	jdff dff_A_PIzinJ1w3_0(.dout(w_dff_A_fBhv2TTk2_0),.din(w_dff_A_PIzinJ1w3_0),.clk(gclk));
	jdff dff_A_fBhv2TTk2_0(.dout(w_dff_A_pw1HQgXf1_0),.din(w_dff_A_fBhv2TTk2_0),.clk(gclk));
	jdff dff_A_pw1HQgXf1_0(.dout(w_dff_A_bp4RaVkA5_0),.din(w_dff_A_pw1HQgXf1_0),.clk(gclk));
	jdff dff_A_bp4RaVkA5_0(.dout(w_dff_A_tkiJsETO3_0),.din(w_dff_A_bp4RaVkA5_0),.clk(gclk));
	jdff dff_A_tkiJsETO3_0(.dout(w_dff_A_2jZ0Yaw72_0),.din(w_dff_A_tkiJsETO3_0),.clk(gclk));
	jdff dff_A_2jZ0Yaw72_0(.dout(w_dff_A_wKnrJxZZ7_0),.din(w_dff_A_2jZ0Yaw72_0),.clk(gclk));
	jdff dff_A_wKnrJxZZ7_0(.dout(w_dff_A_KHCyhPaf7_0),.din(w_dff_A_wKnrJxZZ7_0),.clk(gclk));
	jdff dff_A_KHCyhPaf7_0(.dout(w_dff_A_g8dTMHiq0_0),.din(w_dff_A_KHCyhPaf7_0),.clk(gclk));
	jdff dff_A_g8dTMHiq0_0(.dout(w_dff_A_Cmuj7iFG0_0),.din(w_dff_A_g8dTMHiq0_0),.clk(gclk));
	jdff dff_A_Cmuj7iFG0_0(.dout(w_dff_A_s01I0WgX4_0),.din(w_dff_A_Cmuj7iFG0_0),.clk(gclk));
	jdff dff_A_s01I0WgX4_0(.dout(w_dff_A_cmdd8QJ67_0),.din(w_dff_A_s01I0WgX4_0),.clk(gclk));
	jdff dff_A_cmdd8QJ67_0(.dout(w_dff_A_7wJiYFI65_0),.din(w_dff_A_cmdd8QJ67_0),.clk(gclk));
	jdff dff_A_7wJiYFI65_0(.dout(w_dff_A_qHkBqdhz5_0),.din(w_dff_A_7wJiYFI65_0),.clk(gclk));
	jdff dff_A_qHkBqdhz5_0(.dout(w_dff_A_t4wnJ0ts3_0),.din(w_dff_A_qHkBqdhz5_0),.clk(gclk));
	jdff dff_A_t4wnJ0ts3_0(.dout(w_dff_A_IxgCif1n3_0),.din(w_dff_A_t4wnJ0ts3_0),.clk(gclk));
	jdff dff_A_IxgCif1n3_0(.dout(w_dff_A_HWhrWMmM0_0),.din(w_dff_A_IxgCif1n3_0),.clk(gclk));
	jdff dff_A_HWhrWMmM0_0(.dout(w_dff_A_rLl4xzb80_0),.din(w_dff_A_HWhrWMmM0_0),.clk(gclk));
	jdff dff_A_rLl4xzb80_0(.dout(w_dff_A_36qrJKoI2_0),.din(w_dff_A_rLl4xzb80_0),.clk(gclk));
	jdff dff_A_36qrJKoI2_0(.dout(w_dff_A_T1lLeCux0_0),.din(w_dff_A_36qrJKoI2_0),.clk(gclk));
	jdff dff_A_T1lLeCux0_0(.dout(G144),.din(w_dff_A_T1lLeCux0_0),.clk(gclk));
	jdff dff_A_66TVFEek2_1(.dout(w_dff_A_e6Tt3Oxu1_0),.din(w_dff_A_66TVFEek2_1),.clk(gclk));
	jdff dff_A_e6Tt3Oxu1_0(.dout(w_dff_A_vbjLKxae7_0),.din(w_dff_A_e6Tt3Oxu1_0),.clk(gclk));
	jdff dff_A_vbjLKxae7_0(.dout(w_dff_A_3PHrQZBh9_0),.din(w_dff_A_vbjLKxae7_0),.clk(gclk));
	jdff dff_A_3PHrQZBh9_0(.dout(w_dff_A_UD7NvugM4_0),.din(w_dff_A_3PHrQZBh9_0),.clk(gclk));
	jdff dff_A_UD7NvugM4_0(.dout(w_dff_A_8wRcVrZn2_0),.din(w_dff_A_UD7NvugM4_0),.clk(gclk));
	jdff dff_A_8wRcVrZn2_0(.dout(w_dff_A_GqtQunKv8_0),.din(w_dff_A_8wRcVrZn2_0),.clk(gclk));
	jdff dff_A_GqtQunKv8_0(.dout(w_dff_A_4SX7KZ3w3_0),.din(w_dff_A_GqtQunKv8_0),.clk(gclk));
	jdff dff_A_4SX7KZ3w3_0(.dout(w_dff_A_88Cq0ZWY9_0),.din(w_dff_A_4SX7KZ3w3_0),.clk(gclk));
	jdff dff_A_88Cq0ZWY9_0(.dout(w_dff_A_8AS9GNjx5_0),.din(w_dff_A_88Cq0ZWY9_0),.clk(gclk));
	jdff dff_A_8AS9GNjx5_0(.dout(w_dff_A_QHDwokZ27_0),.din(w_dff_A_8AS9GNjx5_0),.clk(gclk));
	jdff dff_A_QHDwokZ27_0(.dout(w_dff_A_0vs2Z1sl0_0),.din(w_dff_A_QHDwokZ27_0),.clk(gclk));
	jdff dff_A_0vs2Z1sl0_0(.dout(w_dff_A_ZBBrLpEV9_0),.din(w_dff_A_0vs2Z1sl0_0),.clk(gclk));
	jdff dff_A_ZBBrLpEV9_0(.dout(w_dff_A_zbhioTiY5_0),.din(w_dff_A_ZBBrLpEV9_0),.clk(gclk));
	jdff dff_A_zbhioTiY5_0(.dout(w_dff_A_F3ynzS6p1_0),.din(w_dff_A_zbhioTiY5_0),.clk(gclk));
	jdff dff_A_F3ynzS6p1_0(.dout(w_dff_A_i7kv418J8_0),.din(w_dff_A_F3ynzS6p1_0),.clk(gclk));
	jdff dff_A_i7kv418J8_0(.dout(w_dff_A_wjeJJvUX7_0),.din(w_dff_A_i7kv418J8_0),.clk(gclk));
	jdff dff_A_wjeJJvUX7_0(.dout(w_dff_A_991H8U6N3_0),.din(w_dff_A_wjeJJvUX7_0),.clk(gclk));
	jdff dff_A_991H8U6N3_0(.dout(w_dff_A_jIgKbxMV3_0),.din(w_dff_A_991H8U6N3_0),.clk(gclk));
	jdff dff_A_jIgKbxMV3_0(.dout(w_dff_A_DsI9Q1i31_0),.din(w_dff_A_jIgKbxMV3_0),.clk(gclk));
	jdff dff_A_DsI9Q1i31_0(.dout(w_dff_A_YgsK38Qp9_0),.din(w_dff_A_DsI9Q1i31_0),.clk(gclk));
	jdff dff_A_YgsK38Qp9_0(.dout(w_dff_A_ZNmpkZwe4_0),.din(w_dff_A_YgsK38Qp9_0),.clk(gclk));
	jdff dff_A_ZNmpkZwe4_0(.dout(w_dff_A_zR3TTkFu2_0),.din(w_dff_A_ZNmpkZwe4_0),.clk(gclk));
	jdff dff_A_zR3TTkFu2_0(.dout(w_dff_A_lPROXJ9D8_0),.din(w_dff_A_zR3TTkFu2_0),.clk(gclk));
	jdff dff_A_lPROXJ9D8_0(.dout(w_dff_A_Q1c3rkbg4_0),.din(w_dff_A_lPROXJ9D8_0),.clk(gclk));
	jdff dff_A_Q1c3rkbg4_0(.dout(w_dff_A_UxRSzE180_0),.din(w_dff_A_Q1c3rkbg4_0),.clk(gclk));
	jdff dff_A_UxRSzE180_0(.dout(w_dff_A_xVDouYFF1_0),.din(w_dff_A_UxRSzE180_0),.clk(gclk));
	jdff dff_A_xVDouYFF1_0(.dout(w_dff_A_Kq4rLhGI3_0),.din(w_dff_A_xVDouYFF1_0),.clk(gclk));
	jdff dff_A_Kq4rLhGI3_0(.dout(G298),.din(w_dff_A_Kq4rLhGI3_0),.clk(gclk));
	jdff dff_A_cOzPVBtM3_1(.dout(w_dff_A_72ZR4UTZ7_0),.din(w_dff_A_cOzPVBtM3_1),.clk(gclk));
	jdff dff_A_72ZR4UTZ7_0(.dout(w_dff_A_Bf504nHY0_0),.din(w_dff_A_72ZR4UTZ7_0),.clk(gclk));
	jdff dff_A_Bf504nHY0_0(.dout(w_dff_A_f9QXljEo8_0),.din(w_dff_A_Bf504nHY0_0),.clk(gclk));
	jdff dff_A_f9QXljEo8_0(.dout(w_dff_A_eC9nqIBI8_0),.din(w_dff_A_f9QXljEo8_0),.clk(gclk));
	jdff dff_A_eC9nqIBI8_0(.dout(w_dff_A_QRCuucQo4_0),.din(w_dff_A_eC9nqIBI8_0),.clk(gclk));
	jdff dff_A_QRCuucQo4_0(.dout(w_dff_A_dsQe4pSS1_0),.din(w_dff_A_QRCuucQo4_0),.clk(gclk));
	jdff dff_A_dsQe4pSS1_0(.dout(w_dff_A_Bb4uoTXu1_0),.din(w_dff_A_dsQe4pSS1_0),.clk(gclk));
	jdff dff_A_Bb4uoTXu1_0(.dout(w_dff_A_HROEk1dt9_0),.din(w_dff_A_Bb4uoTXu1_0),.clk(gclk));
	jdff dff_A_HROEk1dt9_0(.dout(w_dff_A_XWlpIgNq2_0),.din(w_dff_A_HROEk1dt9_0),.clk(gclk));
	jdff dff_A_XWlpIgNq2_0(.dout(w_dff_A_HE5m0u697_0),.din(w_dff_A_XWlpIgNq2_0),.clk(gclk));
	jdff dff_A_HE5m0u697_0(.dout(w_dff_A_PU03U1h99_0),.din(w_dff_A_HE5m0u697_0),.clk(gclk));
	jdff dff_A_PU03U1h99_0(.dout(w_dff_A_y5XCgYBi9_0),.din(w_dff_A_PU03U1h99_0),.clk(gclk));
	jdff dff_A_y5XCgYBi9_0(.dout(w_dff_A_X9rOq4NT7_0),.din(w_dff_A_y5XCgYBi9_0),.clk(gclk));
	jdff dff_A_X9rOq4NT7_0(.dout(w_dff_A_QjSIHy7p6_0),.din(w_dff_A_X9rOq4NT7_0),.clk(gclk));
	jdff dff_A_QjSIHy7p6_0(.dout(w_dff_A_vGBqmh7w4_0),.din(w_dff_A_QjSIHy7p6_0),.clk(gclk));
	jdff dff_A_vGBqmh7w4_0(.dout(w_dff_A_1IoinElv1_0),.din(w_dff_A_vGBqmh7w4_0),.clk(gclk));
	jdff dff_A_1IoinElv1_0(.dout(w_dff_A_YxVaFZGm1_0),.din(w_dff_A_1IoinElv1_0),.clk(gclk));
	jdff dff_A_YxVaFZGm1_0(.dout(w_dff_A_TTaP4J3h7_0),.din(w_dff_A_YxVaFZGm1_0),.clk(gclk));
	jdff dff_A_TTaP4J3h7_0(.dout(w_dff_A_0JrGIvkU7_0),.din(w_dff_A_TTaP4J3h7_0),.clk(gclk));
	jdff dff_A_0JrGIvkU7_0(.dout(w_dff_A_Povm8g0T8_0),.din(w_dff_A_0JrGIvkU7_0),.clk(gclk));
	jdff dff_A_Povm8g0T8_0(.dout(w_dff_A_98x0DwU05_0),.din(w_dff_A_Povm8g0T8_0),.clk(gclk));
	jdff dff_A_98x0DwU05_0(.dout(w_dff_A_J6FQE78K4_0),.din(w_dff_A_98x0DwU05_0),.clk(gclk));
	jdff dff_A_J6FQE78K4_0(.dout(w_dff_A_c7QpQhh33_0),.din(w_dff_A_J6FQE78K4_0),.clk(gclk));
	jdff dff_A_c7QpQhh33_0(.dout(w_dff_A_r7UGk4pr6_0),.din(w_dff_A_c7QpQhh33_0),.clk(gclk));
	jdff dff_A_r7UGk4pr6_0(.dout(w_dff_A_j0fGoIma0_0),.din(w_dff_A_r7UGk4pr6_0),.clk(gclk));
	jdff dff_A_j0fGoIma0_0(.dout(w_dff_A_6ru6Hf1c0_0),.din(w_dff_A_j0fGoIma0_0),.clk(gclk));
	jdff dff_A_6ru6Hf1c0_0(.dout(w_dff_A_B6D4QjdY1_0),.din(w_dff_A_6ru6Hf1c0_0),.clk(gclk));
	jdff dff_A_B6D4QjdY1_0(.dout(G973),.din(w_dff_A_B6D4QjdY1_0),.clk(gclk));
	jdff dff_A_ZBrec1Vu5_1(.dout(w_dff_A_9HjHzhb74_0),.din(w_dff_A_ZBrec1Vu5_1),.clk(gclk));
	jdff dff_A_9HjHzhb74_0(.dout(w_dff_A_0gQLt4rn2_0),.din(w_dff_A_9HjHzhb74_0),.clk(gclk));
	jdff dff_A_0gQLt4rn2_0(.dout(w_dff_A_ZhY6jJLm8_0),.din(w_dff_A_0gQLt4rn2_0),.clk(gclk));
	jdff dff_A_ZhY6jJLm8_0(.dout(w_dff_A_ZTcwPJYb6_0),.din(w_dff_A_ZhY6jJLm8_0),.clk(gclk));
	jdff dff_A_ZTcwPJYb6_0(.dout(w_dff_A_OmtjDjBq0_0),.din(w_dff_A_ZTcwPJYb6_0),.clk(gclk));
	jdff dff_A_OmtjDjBq0_0(.dout(w_dff_A_LLOIkHnB4_0),.din(w_dff_A_OmtjDjBq0_0),.clk(gclk));
	jdff dff_A_LLOIkHnB4_0(.dout(w_dff_A_AsGV2thy5_0),.din(w_dff_A_LLOIkHnB4_0),.clk(gclk));
	jdff dff_A_AsGV2thy5_0(.dout(w_dff_A_nNHQaBxV0_0),.din(w_dff_A_AsGV2thy5_0),.clk(gclk));
	jdff dff_A_nNHQaBxV0_0(.dout(w_dff_A_PZ6END2h6_0),.din(w_dff_A_nNHQaBxV0_0),.clk(gclk));
	jdff dff_A_PZ6END2h6_0(.dout(w_dff_A_NFJO4cCu4_0),.din(w_dff_A_PZ6END2h6_0),.clk(gclk));
	jdff dff_A_NFJO4cCu4_0(.dout(w_dff_A_d7wBAC4s8_0),.din(w_dff_A_NFJO4cCu4_0),.clk(gclk));
	jdff dff_A_d7wBAC4s8_0(.dout(w_dff_A_Dcbnwu9o5_0),.din(w_dff_A_d7wBAC4s8_0),.clk(gclk));
	jdff dff_A_Dcbnwu9o5_0(.dout(w_dff_A_iBrDHkMn3_0),.din(w_dff_A_Dcbnwu9o5_0),.clk(gclk));
	jdff dff_A_iBrDHkMn3_0(.dout(w_dff_A_FOW0lCgf3_0),.din(w_dff_A_iBrDHkMn3_0),.clk(gclk));
	jdff dff_A_FOW0lCgf3_0(.dout(w_dff_A_geZbrlJo1_0),.din(w_dff_A_FOW0lCgf3_0),.clk(gclk));
	jdff dff_A_geZbrlJo1_0(.dout(w_dff_A_rRuZsvsK4_0),.din(w_dff_A_geZbrlJo1_0),.clk(gclk));
	jdff dff_A_rRuZsvsK4_0(.dout(w_dff_A_dsPzCTFW9_0),.din(w_dff_A_rRuZsvsK4_0),.clk(gclk));
	jdff dff_A_dsPzCTFW9_0(.dout(w_dff_A_9plZiwZc3_0),.din(w_dff_A_dsPzCTFW9_0),.clk(gclk));
	jdff dff_A_9plZiwZc3_0(.dout(w_dff_A_XO8tngcP9_0),.din(w_dff_A_9plZiwZc3_0),.clk(gclk));
	jdff dff_A_XO8tngcP9_0(.dout(w_dff_A_LQamYGXh8_0),.din(w_dff_A_XO8tngcP9_0),.clk(gclk));
	jdff dff_A_LQamYGXh8_0(.dout(w_dff_A_i3kEDeyu6_0),.din(w_dff_A_LQamYGXh8_0),.clk(gclk));
	jdff dff_A_i3kEDeyu6_0(.dout(w_dff_A_oaO3PXFu2_0),.din(w_dff_A_i3kEDeyu6_0),.clk(gclk));
	jdff dff_A_oaO3PXFu2_0(.dout(w_dff_A_HA5vElS69_0),.din(w_dff_A_oaO3PXFu2_0),.clk(gclk));
	jdff dff_A_HA5vElS69_0(.dout(w_dff_A_z1KxBbj12_0),.din(w_dff_A_HA5vElS69_0),.clk(gclk));
	jdff dff_A_z1KxBbj12_0(.dout(w_dff_A_NEWGDjVD2_0),.din(w_dff_A_z1KxBbj12_0),.clk(gclk));
	jdff dff_A_NEWGDjVD2_0(.dout(w_dff_A_LMxUAXnI3_0),.din(w_dff_A_NEWGDjVD2_0),.clk(gclk));
	jdff dff_A_LMxUAXnI3_0(.dout(G594),.din(w_dff_A_LMxUAXnI3_0),.clk(gclk));
	jdff dff_A_LWbmaDOx7_1(.dout(w_dff_A_G77qIhlB1_0),.din(w_dff_A_LWbmaDOx7_1),.clk(gclk));
	jdff dff_A_G77qIhlB1_0(.dout(w_dff_A_ZH3LWzlQ5_0),.din(w_dff_A_G77qIhlB1_0),.clk(gclk));
	jdff dff_A_ZH3LWzlQ5_0(.dout(w_dff_A_lFnt3W3e4_0),.din(w_dff_A_ZH3LWzlQ5_0),.clk(gclk));
	jdff dff_A_lFnt3W3e4_0(.dout(w_dff_A_ZA2xwnUC4_0),.din(w_dff_A_lFnt3W3e4_0),.clk(gclk));
	jdff dff_A_ZA2xwnUC4_0(.dout(w_dff_A_CavUfkSL4_0),.din(w_dff_A_ZA2xwnUC4_0),.clk(gclk));
	jdff dff_A_CavUfkSL4_0(.dout(w_dff_A_ftBqPUNs2_0),.din(w_dff_A_CavUfkSL4_0),.clk(gclk));
	jdff dff_A_ftBqPUNs2_0(.dout(w_dff_A_vMfyVpXQ3_0),.din(w_dff_A_ftBqPUNs2_0),.clk(gclk));
	jdff dff_A_vMfyVpXQ3_0(.dout(w_dff_A_6bzKCMHS7_0),.din(w_dff_A_vMfyVpXQ3_0),.clk(gclk));
	jdff dff_A_6bzKCMHS7_0(.dout(w_dff_A_81IYzGyB2_0),.din(w_dff_A_6bzKCMHS7_0),.clk(gclk));
	jdff dff_A_81IYzGyB2_0(.dout(w_dff_A_iWBIU4cS1_0),.din(w_dff_A_81IYzGyB2_0),.clk(gclk));
	jdff dff_A_iWBIU4cS1_0(.dout(w_dff_A_KpoOcQ1n0_0),.din(w_dff_A_iWBIU4cS1_0),.clk(gclk));
	jdff dff_A_KpoOcQ1n0_0(.dout(w_dff_A_qGUqL9le2_0),.din(w_dff_A_KpoOcQ1n0_0),.clk(gclk));
	jdff dff_A_qGUqL9le2_0(.dout(w_dff_A_FY8epnLO2_0),.din(w_dff_A_qGUqL9le2_0),.clk(gclk));
	jdff dff_A_FY8epnLO2_0(.dout(w_dff_A_58mLI5xt3_0),.din(w_dff_A_FY8epnLO2_0),.clk(gclk));
	jdff dff_A_58mLI5xt3_0(.dout(w_dff_A_LOIpxovQ5_0),.din(w_dff_A_58mLI5xt3_0),.clk(gclk));
	jdff dff_A_LOIpxovQ5_0(.dout(w_dff_A_U7TwF1Fc3_0),.din(w_dff_A_LOIpxovQ5_0),.clk(gclk));
	jdff dff_A_U7TwF1Fc3_0(.dout(w_dff_A_anaQSJ0f6_0),.din(w_dff_A_U7TwF1Fc3_0),.clk(gclk));
	jdff dff_A_anaQSJ0f6_0(.dout(w_dff_A_oc0T40gt3_0),.din(w_dff_A_anaQSJ0f6_0),.clk(gclk));
	jdff dff_A_oc0T40gt3_0(.dout(w_dff_A_rG0LNEBt9_0),.din(w_dff_A_oc0T40gt3_0),.clk(gclk));
	jdff dff_A_rG0LNEBt9_0(.dout(w_dff_A_vSmwMge69_0),.din(w_dff_A_rG0LNEBt9_0),.clk(gclk));
	jdff dff_A_vSmwMge69_0(.dout(w_dff_A_PtCPtguF5_0),.din(w_dff_A_vSmwMge69_0),.clk(gclk));
	jdff dff_A_PtCPtguF5_0(.dout(w_dff_A_5qDUjCvt6_0),.din(w_dff_A_PtCPtguF5_0),.clk(gclk));
	jdff dff_A_5qDUjCvt6_0(.dout(w_dff_A_hEjpu3F45_0),.din(w_dff_A_5qDUjCvt6_0),.clk(gclk));
	jdff dff_A_hEjpu3F45_0(.dout(w_dff_A_Y4JP3PhZ8_0),.din(w_dff_A_hEjpu3F45_0),.clk(gclk));
	jdff dff_A_Y4JP3PhZ8_0(.dout(w_dff_A_pczSir390_0),.din(w_dff_A_Y4JP3PhZ8_0),.clk(gclk));
	jdff dff_A_pczSir390_0(.dout(w_dff_A_0yq65Dyx6_0),.din(w_dff_A_pczSir390_0),.clk(gclk));
	jdff dff_A_0yq65Dyx6_0(.dout(G599),.din(w_dff_A_0yq65Dyx6_0),.clk(gclk));
	jdff dff_A_9M7VFoQ81_1(.dout(w_dff_A_Z1yuy3GJ8_0),.din(w_dff_A_9M7VFoQ81_1),.clk(gclk));
	jdff dff_A_Z1yuy3GJ8_0(.dout(w_dff_A_OJom6nUJ8_0),.din(w_dff_A_Z1yuy3GJ8_0),.clk(gclk));
	jdff dff_A_OJom6nUJ8_0(.dout(w_dff_A_6iUYxKgP2_0),.din(w_dff_A_OJom6nUJ8_0),.clk(gclk));
	jdff dff_A_6iUYxKgP2_0(.dout(w_dff_A_51N8aG8j0_0),.din(w_dff_A_6iUYxKgP2_0),.clk(gclk));
	jdff dff_A_51N8aG8j0_0(.dout(w_dff_A_U51uCfT92_0),.din(w_dff_A_51N8aG8j0_0),.clk(gclk));
	jdff dff_A_U51uCfT92_0(.dout(w_dff_A_wlNgaXLk5_0),.din(w_dff_A_U51uCfT92_0),.clk(gclk));
	jdff dff_A_wlNgaXLk5_0(.dout(w_dff_A_HJXjAIbc2_0),.din(w_dff_A_wlNgaXLk5_0),.clk(gclk));
	jdff dff_A_HJXjAIbc2_0(.dout(w_dff_A_0N9jKlA57_0),.din(w_dff_A_HJXjAIbc2_0),.clk(gclk));
	jdff dff_A_0N9jKlA57_0(.dout(w_dff_A_Y0ccbfKC2_0),.din(w_dff_A_0N9jKlA57_0),.clk(gclk));
	jdff dff_A_Y0ccbfKC2_0(.dout(w_dff_A_OAc49W245_0),.din(w_dff_A_Y0ccbfKC2_0),.clk(gclk));
	jdff dff_A_OAc49W245_0(.dout(w_dff_A_GAlBH3L10_0),.din(w_dff_A_OAc49W245_0),.clk(gclk));
	jdff dff_A_GAlBH3L10_0(.dout(w_dff_A_PsPZevd36_0),.din(w_dff_A_GAlBH3L10_0),.clk(gclk));
	jdff dff_A_PsPZevd36_0(.dout(w_dff_A_1WbWD7117_0),.din(w_dff_A_PsPZevd36_0),.clk(gclk));
	jdff dff_A_1WbWD7117_0(.dout(w_dff_A_pvVFRsvR6_0),.din(w_dff_A_1WbWD7117_0),.clk(gclk));
	jdff dff_A_pvVFRsvR6_0(.dout(w_dff_A_nqLPrIOh3_0),.din(w_dff_A_pvVFRsvR6_0),.clk(gclk));
	jdff dff_A_nqLPrIOh3_0(.dout(w_dff_A_fNSJmsjO5_0),.din(w_dff_A_nqLPrIOh3_0),.clk(gclk));
	jdff dff_A_fNSJmsjO5_0(.dout(w_dff_A_h2JhboCa1_0),.din(w_dff_A_fNSJmsjO5_0),.clk(gclk));
	jdff dff_A_h2JhboCa1_0(.dout(w_dff_A_xI4VORAL7_0),.din(w_dff_A_h2JhboCa1_0),.clk(gclk));
	jdff dff_A_xI4VORAL7_0(.dout(w_dff_A_EDFjdaGP7_0),.din(w_dff_A_xI4VORAL7_0),.clk(gclk));
	jdff dff_A_EDFjdaGP7_0(.dout(w_dff_A_cjoo9Vqa8_0),.din(w_dff_A_EDFjdaGP7_0),.clk(gclk));
	jdff dff_A_cjoo9Vqa8_0(.dout(w_dff_A_sAlipV9a1_0),.din(w_dff_A_cjoo9Vqa8_0),.clk(gclk));
	jdff dff_A_sAlipV9a1_0(.dout(w_dff_A_PoJJFXU00_0),.din(w_dff_A_sAlipV9a1_0),.clk(gclk));
	jdff dff_A_PoJJFXU00_0(.dout(w_dff_A_cqVpYbPl9_0),.din(w_dff_A_PoJJFXU00_0),.clk(gclk));
	jdff dff_A_cqVpYbPl9_0(.dout(w_dff_A_PzacCgIN6_0),.din(w_dff_A_cqVpYbPl9_0),.clk(gclk));
	jdff dff_A_PzacCgIN6_0(.dout(w_dff_A_HG9QmtQO8_0),.din(w_dff_A_PzacCgIN6_0),.clk(gclk));
	jdff dff_A_HG9QmtQO8_0(.dout(w_dff_A_wyoToT9J2_0),.din(w_dff_A_HG9QmtQO8_0),.clk(gclk));
	jdff dff_A_wyoToT9J2_0(.dout(G600),.din(w_dff_A_wyoToT9J2_0),.clk(gclk));
	jdff dff_A_ErVd9dvY1_1(.dout(w_dff_A_mQlTFZrd0_0),.din(w_dff_A_ErVd9dvY1_1),.clk(gclk));
	jdff dff_A_mQlTFZrd0_0(.dout(w_dff_A_6AC4U78P0_0),.din(w_dff_A_mQlTFZrd0_0),.clk(gclk));
	jdff dff_A_6AC4U78P0_0(.dout(w_dff_A_z6lRIJMC3_0),.din(w_dff_A_6AC4U78P0_0),.clk(gclk));
	jdff dff_A_z6lRIJMC3_0(.dout(w_dff_A_iwMok4iD9_0),.din(w_dff_A_z6lRIJMC3_0),.clk(gclk));
	jdff dff_A_iwMok4iD9_0(.dout(w_dff_A_Mi1JnWHR1_0),.din(w_dff_A_iwMok4iD9_0),.clk(gclk));
	jdff dff_A_Mi1JnWHR1_0(.dout(w_dff_A_IMMCMqfQ5_0),.din(w_dff_A_Mi1JnWHR1_0),.clk(gclk));
	jdff dff_A_IMMCMqfQ5_0(.dout(w_dff_A_zvT66J7n0_0),.din(w_dff_A_IMMCMqfQ5_0),.clk(gclk));
	jdff dff_A_zvT66J7n0_0(.dout(w_dff_A_WDBcrvJJ8_0),.din(w_dff_A_zvT66J7n0_0),.clk(gclk));
	jdff dff_A_WDBcrvJJ8_0(.dout(w_dff_A_qXcma8tL2_0),.din(w_dff_A_WDBcrvJJ8_0),.clk(gclk));
	jdff dff_A_qXcma8tL2_0(.dout(w_dff_A_2fwqvAeD6_0),.din(w_dff_A_qXcma8tL2_0),.clk(gclk));
	jdff dff_A_2fwqvAeD6_0(.dout(w_dff_A_YbE3af0v7_0),.din(w_dff_A_2fwqvAeD6_0),.clk(gclk));
	jdff dff_A_YbE3af0v7_0(.dout(w_dff_A_doDlAHgH6_0),.din(w_dff_A_YbE3af0v7_0),.clk(gclk));
	jdff dff_A_doDlAHgH6_0(.dout(w_dff_A_HzYboDvG1_0),.din(w_dff_A_doDlAHgH6_0),.clk(gclk));
	jdff dff_A_HzYboDvG1_0(.dout(w_dff_A_iVrSmTkO0_0),.din(w_dff_A_HzYboDvG1_0),.clk(gclk));
	jdff dff_A_iVrSmTkO0_0(.dout(w_dff_A_7E6Dxsf10_0),.din(w_dff_A_iVrSmTkO0_0),.clk(gclk));
	jdff dff_A_7E6Dxsf10_0(.dout(w_dff_A_QhCoLZ5E6_0),.din(w_dff_A_7E6Dxsf10_0),.clk(gclk));
	jdff dff_A_QhCoLZ5E6_0(.dout(w_dff_A_Du10hnrC4_0),.din(w_dff_A_QhCoLZ5E6_0),.clk(gclk));
	jdff dff_A_Du10hnrC4_0(.dout(w_dff_A_VauC8AWi1_0),.din(w_dff_A_Du10hnrC4_0),.clk(gclk));
	jdff dff_A_VauC8AWi1_0(.dout(w_dff_A_zEDOjqZP2_0),.din(w_dff_A_VauC8AWi1_0),.clk(gclk));
	jdff dff_A_zEDOjqZP2_0(.dout(w_dff_A_rsbtDTkc7_0),.din(w_dff_A_zEDOjqZP2_0),.clk(gclk));
	jdff dff_A_rsbtDTkc7_0(.dout(w_dff_A_OyM4Ma0l9_0),.din(w_dff_A_rsbtDTkc7_0),.clk(gclk));
	jdff dff_A_OyM4Ma0l9_0(.dout(w_dff_A_WARWnHPy8_0),.din(w_dff_A_OyM4Ma0l9_0),.clk(gclk));
	jdff dff_A_WARWnHPy8_0(.dout(w_dff_A_zDAKdEI92_0),.din(w_dff_A_WARWnHPy8_0),.clk(gclk));
	jdff dff_A_zDAKdEI92_0(.dout(w_dff_A_tyEl8rog7_0),.din(w_dff_A_zDAKdEI92_0),.clk(gclk));
	jdff dff_A_tyEl8rog7_0(.dout(w_dff_A_1JraaIEI2_0),.din(w_dff_A_tyEl8rog7_0),.clk(gclk));
	jdff dff_A_1JraaIEI2_0(.dout(w_dff_A_k7cQgACV4_0),.din(w_dff_A_1JraaIEI2_0),.clk(gclk));
	jdff dff_A_k7cQgACV4_0(.dout(G601),.din(w_dff_A_k7cQgACV4_0),.clk(gclk));
	jdff dff_A_KwFthaXT7_1(.dout(w_dff_A_oaR4YbRs8_0),.din(w_dff_A_KwFthaXT7_1),.clk(gclk));
	jdff dff_A_oaR4YbRs8_0(.dout(w_dff_A_XZOVlZ2x5_0),.din(w_dff_A_oaR4YbRs8_0),.clk(gclk));
	jdff dff_A_XZOVlZ2x5_0(.dout(w_dff_A_vnFPic539_0),.din(w_dff_A_XZOVlZ2x5_0),.clk(gclk));
	jdff dff_A_vnFPic539_0(.dout(w_dff_A_pkUTM2qt5_0),.din(w_dff_A_vnFPic539_0),.clk(gclk));
	jdff dff_A_pkUTM2qt5_0(.dout(w_dff_A_DGSN06W86_0),.din(w_dff_A_pkUTM2qt5_0),.clk(gclk));
	jdff dff_A_DGSN06W86_0(.dout(w_dff_A_9iVrpYmB5_0),.din(w_dff_A_DGSN06W86_0),.clk(gclk));
	jdff dff_A_9iVrpYmB5_0(.dout(w_dff_A_07LJcw2a4_0),.din(w_dff_A_9iVrpYmB5_0),.clk(gclk));
	jdff dff_A_07LJcw2a4_0(.dout(w_dff_A_APelAM7q8_0),.din(w_dff_A_07LJcw2a4_0),.clk(gclk));
	jdff dff_A_APelAM7q8_0(.dout(w_dff_A_3raM8th58_0),.din(w_dff_A_APelAM7q8_0),.clk(gclk));
	jdff dff_A_3raM8th58_0(.dout(w_dff_A_nR95UGcK1_0),.din(w_dff_A_3raM8th58_0),.clk(gclk));
	jdff dff_A_nR95UGcK1_0(.dout(w_dff_A_BYpW1t7u9_0),.din(w_dff_A_nR95UGcK1_0),.clk(gclk));
	jdff dff_A_BYpW1t7u9_0(.dout(w_dff_A_W5GwHe6f1_0),.din(w_dff_A_BYpW1t7u9_0),.clk(gclk));
	jdff dff_A_W5GwHe6f1_0(.dout(w_dff_A_uWEDh6283_0),.din(w_dff_A_W5GwHe6f1_0),.clk(gclk));
	jdff dff_A_uWEDh6283_0(.dout(w_dff_A_jc1aaP861_0),.din(w_dff_A_uWEDh6283_0),.clk(gclk));
	jdff dff_A_jc1aaP861_0(.dout(w_dff_A_YAC5Br0L1_0),.din(w_dff_A_jc1aaP861_0),.clk(gclk));
	jdff dff_A_YAC5Br0L1_0(.dout(w_dff_A_8wLp2KdT5_0),.din(w_dff_A_YAC5Br0L1_0),.clk(gclk));
	jdff dff_A_8wLp2KdT5_0(.dout(w_dff_A_fNAlytst3_0),.din(w_dff_A_8wLp2KdT5_0),.clk(gclk));
	jdff dff_A_fNAlytst3_0(.dout(w_dff_A_gUrXzxCQ2_0),.din(w_dff_A_fNAlytst3_0),.clk(gclk));
	jdff dff_A_gUrXzxCQ2_0(.dout(w_dff_A_EahSMhEL4_0),.din(w_dff_A_gUrXzxCQ2_0),.clk(gclk));
	jdff dff_A_EahSMhEL4_0(.dout(w_dff_A_zDoResQT0_0),.din(w_dff_A_EahSMhEL4_0),.clk(gclk));
	jdff dff_A_zDoResQT0_0(.dout(w_dff_A_VxDRyiV39_0),.din(w_dff_A_zDoResQT0_0),.clk(gclk));
	jdff dff_A_VxDRyiV39_0(.dout(w_dff_A_4zCX84kg7_0),.din(w_dff_A_VxDRyiV39_0),.clk(gclk));
	jdff dff_A_4zCX84kg7_0(.dout(w_dff_A_rT6o1Hc34_0),.din(w_dff_A_4zCX84kg7_0),.clk(gclk));
	jdff dff_A_rT6o1Hc34_0(.dout(w_dff_A_GvWe8BoL4_0),.din(w_dff_A_rT6o1Hc34_0),.clk(gclk));
	jdff dff_A_GvWe8BoL4_0(.dout(w_dff_A_8cwhzSJf0_0),.din(w_dff_A_GvWe8BoL4_0),.clk(gclk));
	jdff dff_A_8cwhzSJf0_0(.dout(w_dff_A_GPIgC0h77_0),.din(w_dff_A_8cwhzSJf0_0),.clk(gclk));
	jdff dff_A_GPIgC0h77_0(.dout(G602),.din(w_dff_A_GPIgC0h77_0),.clk(gclk));
	jdff dff_A_IfMxj8Bd5_1(.dout(w_dff_A_KebsTOnD7_0),.din(w_dff_A_IfMxj8Bd5_1),.clk(gclk));
	jdff dff_A_KebsTOnD7_0(.dout(w_dff_A_wuINnOS62_0),.din(w_dff_A_KebsTOnD7_0),.clk(gclk));
	jdff dff_A_wuINnOS62_0(.dout(w_dff_A_Ddm5GtEf5_0),.din(w_dff_A_wuINnOS62_0),.clk(gclk));
	jdff dff_A_Ddm5GtEf5_0(.dout(w_dff_A_drb3WDHp9_0),.din(w_dff_A_Ddm5GtEf5_0),.clk(gclk));
	jdff dff_A_drb3WDHp9_0(.dout(w_dff_A_i1ZIJ60J7_0),.din(w_dff_A_drb3WDHp9_0),.clk(gclk));
	jdff dff_A_i1ZIJ60J7_0(.dout(w_dff_A_Ag1qUUy20_0),.din(w_dff_A_i1ZIJ60J7_0),.clk(gclk));
	jdff dff_A_Ag1qUUy20_0(.dout(w_dff_A_BQ6YV57r3_0),.din(w_dff_A_Ag1qUUy20_0),.clk(gclk));
	jdff dff_A_BQ6YV57r3_0(.dout(w_dff_A_3LYRkJKU4_0),.din(w_dff_A_BQ6YV57r3_0),.clk(gclk));
	jdff dff_A_3LYRkJKU4_0(.dout(w_dff_A_Po1kKwBA1_0),.din(w_dff_A_3LYRkJKU4_0),.clk(gclk));
	jdff dff_A_Po1kKwBA1_0(.dout(w_dff_A_Rvwbnp683_0),.din(w_dff_A_Po1kKwBA1_0),.clk(gclk));
	jdff dff_A_Rvwbnp683_0(.dout(w_dff_A_tlEXmYvm3_0),.din(w_dff_A_Rvwbnp683_0),.clk(gclk));
	jdff dff_A_tlEXmYvm3_0(.dout(w_dff_A_Db40u4xW9_0),.din(w_dff_A_tlEXmYvm3_0),.clk(gclk));
	jdff dff_A_Db40u4xW9_0(.dout(w_dff_A_udAuWS4M4_0),.din(w_dff_A_Db40u4xW9_0),.clk(gclk));
	jdff dff_A_udAuWS4M4_0(.dout(w_dff_A_DyuwXitL1_0),.din(w_dff_A_udAuWS4M4_0),.clk(gclk));
	jdff dff_A_DyuwXitL1_0(.dout(w_dff_A_eOu8vCrx4_0),.din(w_dff_A_DyuwXitL1_0),.clk(gclk));
	jdff dff_A_eOu8vCrx4_0(.dout(w_dff_A_W6TKeSxX6_0),.din(w_dff_A_eOu8vCrx4_0),.clk(gclk));
	jdff dff_A_W6TKeSxX6_0(.dout(w_dff_A_giOXoufo4_0),.din(w_dff_A_W6TKeSxX6_0),.clk(gclk));
	jdff dff_A_giOXoufo4_0(.dout(w_dff_A_Q4P7yEMe0_0),.din(w_dff_A_giOXoufo4_0),.clk(gclk));
	jdff dff_A_Q4P7yEMe0_0(.dout(w_dff_A_fR8qyBTb9_0),.din(w_dff_A_Q4P7yEMe0_0),.clk(gclk));
	jdff dff_A_fR8qyBTb9_0(.dout(w_dff_A_idmUBCqj7_0),.din(w_dff_A_fR8qyBTb9_0),.clk(gclk));
	jdff dff_A_idmUBCqj7_0(.dout(w_dff_A_AGAV1MQv2_0),.din(w_dff_A_idmUBCqj7_0),.clk(gclk));
	jdff dff_A_AGAV1MQv2_0(.dout(w_dff_A_oT4cZ4Rn8_0),.din(w_dff_A_AGAV1MQv2_0),.clk(gclk));
	jdff dff_A_oT4cZ4Rn8_0(.dout(w_dff_A_wtVe6uhD5_0),.din(w_dff_A_oT4cZ4Rn8_0),.clk(gclk));
	jdff dff_A_wtVe6uhD5_0(.dout(w_dff_A_LGFMivYR5_0),.din(w_dff_A_wtVe6uhD5_0),.clk(gclk));
	jdff dff_A_LGFMivYR5_0(.dout(w_dff_A_GmVoLtqC1_0),.din(w_dff_A_LGFMivYR5_0),.clk(gclk));
	jdff dff_A_GmVoLtqC1_0(.dout(w_dff_A_PeTVeBSe3_0),.din(w_dff_A_GmVoLtqC1_0),.clk(gclk));
	jdff dff_A_PeTVeBSe3_0(.dout(G603),.din(w_dff_A_PeTVeBSe3_0),.clk(gclk));
	jdff dff_A_O2Tzkydk6_1(.dout(w_dff_A_O45zSPP70_0),.din(w_dff_A_O2Tzkydk6_1),.clk(gclk));
	jdff dff_A_O45zSPP70_0(.dout(w_dff_A_5EwzfoE47_0),.din(w_dff_A_O45zSPP70_0),.clk(gclk));
	jdff dff_A_5EwzfoE47_0(.dout(w_dff_A_RHTKb1qR8_0),.din(w_dff_A_5EwzfoE47_0),.clk(gclk));
	jdff dff_A_RHTKb1qR8_0(.dout(w_dff_A_oki8ZLtg1_0),.din(w_dff_A_RHTKb1qR8_0),.clk(gclk));
	jdff dff_A_oki8ZLtg1_0(.dout(w_dff_A_kJXcSCHo4_0),.din(w_dff_A_oki8ZLtg1_0),.clk(gclk));
	jdff dff_A_kJXcSCHo4_0(.dout(w_dff_A_UpkQRyx18_0),.din(w_dff_A_kJXcSCHo4_0),.clk(gclk));
	jdff dff_A_UpkQRyx18_0(.dout(w_dff_A_woYCIYZu2_0),.din(w_dff_A_UpkQRyx18_0),.clk(gclk));
	jdff dff_A_woYCIYZu2_0(.dout(w_dff_A_gwBPAcOl9_0),.din(w_dff_A_woYCIYZu2_0),.clk(gclk));
	jdff dff_A_gwBPAcOl9_0(.dout(w_dff_A_sfWtZCMB3_0),.din(w_dff_A_gwBPAcOl9_0),.clk(gclk));
	jdff dff_A_sfWtZCMB3_0(.dout(w_dff_A_cDUBZR605_0),.din(w_dff_A_sfWtZCMB3_0),.clk(gclk));
	jdff dff_A_cDUBZR605_0(.dout(w_dff_A_In1RWngt4_0),.din(w_dff_A_cDUBZR605_0),.clk(gclk));
	jdff dff_A_In1RWngt4_0(.dout(w_dff_A_VgIREoql1_0),.din(w_dff_A_In1RWngt4_0),.clk(gclk));
	jdff dff_A_VgIREoql1_0(.dout(w_dff_A_GbkU81ud2_0),.din(w_dff_A_VgIREoql1_0),.clk(gclk));
	jdff dff_A_GbkU81ud2_0(.dout(w_dff_A_D4D9Vdl01_0),.din(w_dff_A_GbkU81ud2_0),.clk(gclk));
	jdff dff_A_D4D9Vdl01_0(.dout(w_dff_A_me2yGOhm7_0),.din(w_dff_A_D4D9Vdl01_0),.clk(gclk));
	jdff dff_A_me2yGOhm7_0(.dout(w_dff_A_fYmPdThD6_0),.din(w_dff_A_me2yGOhm7_0),.clk(gclk));
	jdff dff_A_fYmPdThD6_0(.dout(w_dff_A_TxJv3yc40_0),.din(w_dff_A_fYmPdThD6_0),.clk(gclk));
	jdff dff_A_TxJv3yc40_0(.dout(w_dff_A_a2sgY9XB8_0),.din(w_dff_A_TxJv3yc40_0),.clk(gclk));
	jdff dff_A_a2sgY9XB8_0(.dout(w_dff_A_WzWtHhzQ2_0),.din(w_dff_A_a2sgY9XB8_0),.clk(gclk));
	jdff dff_A_WzWtHhzQ2_0(.dout(w_dff_A_QRUzJfO15_0),.din(w_dff_A_WzWtHhzQ2_0),.clk(gclk));
	jdff dff_A_QRUzJfO15_0(.dout(w_dff_A_N1g9twN48_0),.din(w_dff_A_QRUzJfO15_0),.clk(gclk));
	jdff dff_A_N1g9twN48_0(.dout(w_dff_A_GdTvfgpX7_0),.din(w_dff_A_N1g9twN48_0),.clk(gclk));
	jdff dff_A_GdTvfgpX7_0(.dout(w_dff_A_51vZNVEY9_0),.din(w_dff_A_GdTvfgpX7_0),.clk(gclk));
	jdff dff_A_51vZNVEY9_0(.dout(w_dff_A_Dc3Yfork6_0),.din(w_dff_A_51vZNVEY9_0),.clk(gclk));
	jdff dff_A_Dc3Yfork6_0(.dout(w_dff_A_zuz5rhrO4_0),.din(w_dff_A_Dc3Yfork6_0),.clk(gclk));
	jdff dff_A_zuz5rhrO4_0(.dout(w_dff_A_5RxE9owP5_0),.din(w_dff_A_zuz5rhrO4_0),.clk(gclk));
	jdff dff_A_5RxE9owP5_0(.dout(G604),.din(w_dff_A_5RxE9owP5_0),.clk(gclk));
	jdff dff_A_UzBVPGlV5_1(.dout(w_dff_A_ON8NVNbY4_0),.din(w_dff_A_UzBVPGlV5_1),.clk(gclk));
	jdff dff_A_ON8NVNbY4_0(.dout(w_dff_A_7qYTwD7H3_0),.din(w_dff_A_ON8NVNbY4_0),.clk(gclk));
	jdff dff_A_7qYTwD7H3_0(.dout(w_dff_A_8ZM378CX9_0),.din(w_dff_A_7qYTwD7H3_0),.clk(gclk));
	jdff dff_A_8ZM378CX9_0(.dout(w_dff_A_kLEJLwSF4_0),.din(w_dff_A_8ZM378CX9_0),.clk(gclk));
	jdff dff_A_kLEJLwSF4_0(.dout(w_dff_A_ZoBkBnAn7_0),.din(w_dff_A_kLEJLwSF4_0),.clk(gclk));
	jdff dff_A_ZoBkBnAn7_0(.dout(w_dff_A_kAmwv8Rx0_0),.din(w_dff_A_ZoBkBnAn7_0),.clk(gclk));
	jdff dff_A_kAmwv8Rx0_0(.dout(w_dff_A_YnusH0PG2_0),.din(w_dff_A_kAmwv8Rx0_0),.clk(gclk));
	jdff dff_A_YnusH0PG2_0(.dout(w_dff_A_AJ24Mydj1_0),.din(w_dff_A_YnusH0PG2_0),.clk(gclk));
	jdff dff_A_AJ24Mydj1_0(.dout(w_dff_A_Gcr3rltz5_0),.din(w_dff_A_AJ24Mydj1_0),.clk(gclk));
	jdff dff_A_Gcr3rltz5_0(.dout(w_dff_A_tRN5YyAv9_0),.din(w_dff_A_Gcr3rltz5_0),.clk(gclk));
	jdff dff_A_tRN5YyAv9_0(.dout(w_dff_A_Pp5CziCW6_0),.din(w_dff_A_tRN5YyAv9_0),.clk(gclk));
	jdff dff_A_Pp5CziCW6_0(.dout(w_dff_A_GzGihGTs2_0),.din(w_dff_A_Pp5CziCW6_0),.clk(gclk));
	jdff dff_A_GzGihGTs2_0(.dout(w_dff_A_RWC9CCZz8_0),.din(w_dff_A_GzGihGTs2_0),.clk(gclk));
	jdff dff_A_RWC9CCZz8_0(.dout(w_dff_A_qnxKGygg9_0),.din(w_dff_A_RWC9CCZz8_0),.clk(gclk));
	jdff dff_A_qnxKGygg9_0(.dout(w_dff_A_IooDKUNC8_0),.din(w_dff_A_qnxKGygg9_0),.clk(gclk));
	jdff dff_A_IooDKUNC8_0(.dout(w_dff_A_TTKMYcMD7_0),.din(w_dff_A_IooDKUNC8_0),.clk(gclk));
	jdff dff_A_TTKMYcMD7_0(.dout(w_dff_A_fkCUzq2r3_0),.din(w_dff_A_TTKMYcMD7_0),.clk(gclk));
	jdff dff_A_fkCUzq2r3_0(.dout(w_dff_A_fIkyIvQl3_0),.din(w_dff_A_fkCUzq2r3_0),.clk(gclk));
	jdff dff_A_fIkyIvQl3_0(.dout(w_dff_A_FxY7VJgL9_0),.din(w_dff_A_fIkyIvQl3_0),.clk(gclk));
	jdff dff_A_FxY7VJgL9_0(.dout(w_dff_A_MvJeQUfX4_0),.din(w_dff_A_FxY7VJgL9_0),.clk(gclk));
	jdff dff_A_MvJeQUfX4_0(.dout(w_dff_A_wqrGHSH05_0),.din(w_dff_A_MvJeQUfX4_0),.clk(gclk));
	jdff dff_A_wqrGHSH05_0(.dout(w_dff_A_EJrXNefK2_0),.din(w_dff_A_wqrGHSH05_0),.clk(gclk));
	jdff dff_A_EJrXNefK2_0(.dout(w_dff_A_5VVAb7Yb0_0),.din(w_dff_A_EJrXNefK2_0),.clk(gclk));
	jdff dff_A_5VVAb7Yb0_0(.dout(w_dff_A_SW2Rxth20_0),.din(w_dff_A_5VVAb7Yb0_0),.clk(gclk));
	jdff dff_A_SW2Rxth20_0(.dout(w_dff_A_67BtqV7a7_0),.din(w_dff_A_SW2Rxth20_0),.clk(gclk));
	jdff dff_A_67BtqV7a7_0(.dout(w_dff_A_qIYPYWs10_0),.din(w_dff_A_67BtqV7a7_0),.clk(gclk));
	jdff dff_A_qIYPYWs10_0(.dout(G611),.din(w_dff_A_qIYPYWs10_0),.clk(gclk));
	jdff dff_A_H84LiIAI2_1(.dout(w_dff_A_klJf9GTN0_0),.din(w_dff_A_H84LiIAI2_1),.clk(gclk));
	jdff dff_A_klJf9GTN0_0(.dout(w_dff_A_dLa3TJ7i4_0),.din(w_dff_A_klJf9GTN0_0),.clk(gclk));
	jdff dff_A_dLa3TJ7i4_0(.dout(w_dff_A_us5feTLe5_0),.din(w_dff_A_dLa3TJ7i4_0),.clk(gclk));
	jdff dff_A_us5feTLe5_0(.dout(w_dff_A_PcnvCYzO8_0),.din(w_dff_A_us5feTLe5_0),.clk(gclk));
	jdff dff_A_PcnvCYzO8_0(.dout(w_dff_A_FmxEbqEg9_0),.din(w_dff_A_PcnvCYzO8_0),.clk(gclk));
	jdff dff_A_FmxEbqEg9_0(.dout(w_dff_A_kNP6ynXm5_0),.din(w_dff_A_FmxEbqEg9_0),.clk(gclk));
	jdff dff_A_kNP6ynXm5_0(.dout(w_dff_A_jC3WmOaw2_0),.din(w_dff_A_kNP6ynXm5_0),.clk(gclk));
	jdff dff_A_jC3WmOaw2_0(.dout(w_dff_A_BewFZWr49_0),.din(w_dff_A_jC3WmOaw2_0),.clk(gclk));
	jdff dff_A_BewFZWr49_0(.dout(w_dff_A_fVUUv8TZ4_0),.din(w_dff_A_BewFZWr49_0),.clk(gclk));
	jdff dff_A_fVUUv8TZ4_0(.dout(w_dff_A_xqlq3lMV8_0),.din(w_dff_A_fVUUv8TZ4_0),.clk(gclk));
	jdff dff_A_xqlq3lMV8_0(.dout(w_dff_A_d2VvDoEr3_0),.din(w_dff_A_xqlq3lMV8_0),.clk(gclk));
	jdff dff_A_d2VvDoEr3_0(.dout(w_dff_A_mKk4ipCh2_0),.din(w_dff_A_d2VvDoEr3_0),.clk(gclk));
	jdff dff_A_mKk4ipCh2_0(.dout(w_dff_A_xvkl5pjR3_0),.din(w_dff_A_mKk4ipCh2_0),.clk(gclk));
	jdff dff_A_xvkl5pjR3_0(.dout(w_dff_A_A885zRif6_0),.din(w_dff_A_xvkl5pjR3_0),.clk(gclk));
	jdff dff_A_A885zRif6_0(.dout(w_dff_A_xoW5Fo8I8_0),.din(w_dff_A_A885zRif6_0),.clk(gclk));
	jdff dff_A_xoW5Fo8I8_0(.dout(w_dff_A_8xd8EdF42_0),.din(w_dff_A_xoW5Fo8I8_0),.clk(gclk));
	jdff dff_A_8xd8EdF42_0(.dout(w_dff_A_LzVFpbsl9_0),.din(w_dff_A_8xd8EdF42_0),.clk(gclk));
	jdff dff_A_LzVFpbsl9_0(.dout(w_dff_A_slUyfZHg6_0),.din(w_dff_A_LzVFpbsl9_0),.clk(gclk));
	jdff dff_A_slUyfZHg6_0(.dout(w_dff_A_DqBZnaXz4_0),.din(w_dff_A_slUyfZHg6_0),.clk(gclk));
	jdff dff_A_DqBZnaXz4_0(.dout(w_dff_A_YoCQdpSa6_0),.din(w_dff_A_DqBZnaXz4_0),.clk(gclk));
	jdff dff_A_YoCQdpSa6_0(.dout(w_dff_A_KkuORzXV5_0),.din(w_dff_A_YoCQdpSa6_0),.clk(gclk));
	jdff dff_A_KkuORzXV5_0(.dout(w_dff_A_azCJmzeU4_0),.din(w_dff_A_KkuORzXV5_0),.clk(gclk));
	jdff dff_A_azCJmzeU4_0(.dout(w_dff_A_6rjkUue98_0),.din(w_dff_A_azCJmzeU4_0),.clk(gclk));
	jdff dff_A_6rjkUue98_0(.dout(w_dff_A_UGrUCVG39_0),.din(w_dff_A_6rjkUue98_0),.clk(gclk));
	jdff dff_A_UGrUCVG39_0(.dout(w_dff_A_Di0Y2KWU5_0),.din(w_dff_A_UGrUCVG39_0),.clk(gclk));
	jdff dff_A_Di0Y2KWU5_0(.dout(w_dff_A_zJhJj7xq5_0),.din(w_dff_A_Di0Y2KWU5_0),.clk(gclk));
	jdff dff_A_zJhJj7xq5_0(.dout(G612),.din(w_dff_A_zJhJj7xq5_0),.clk(gclk));
	jdff dff_A_PGzCSuv27_2(.dout(w_dff_A_nbzROnjq4_0),.din(w_dff_A_PGzCSuv27_2),.clk(gclk));
	jdff dff_A_nbzROnjq4_0(.dout(w_dff_A_31hQn1uG8_0),.din(w_dff_A_nbzROnjq4_0),.clk(gclk));
	jdff dff_A_31hQn1uG8_0(.dout(w_dff_A_emxNW8uW2_0),.din(w_dff_A_31hQn1uG8_0),.clk(gclk));
	jdff dff_A_emxNW8uW2_0(.dout(w_dff_A_xJvEIRen0_0),.din(w_dff_A_emxNW8uW2_0),.clk(gclk));
	jdff dff_A_xJvEIRen0_0(.dout(w_dff_A_7tKrWlig1_0),.din(w_dff_A_xJvEIRen0_0),.clk(gclk));
	jdff dff_A_7tKrWlig1_0(.dout(w_dff_A_iHYwScAp3_0),.din(w_dff_A_7tKrWlig1_0),.clk(gclk));
	jdff dff_A_iHYwScAp3_0(.dout(w_dff_A_FVq1fI5g5_0),.din(w_dff_A_iHYwScAp3_0),.clk(gclk));
	jdff dff_A_FVq1fI5g5_0(.dout(w_dff_A_nhzoLx5Y0_0),.din(w_dff_A_FVq1fI5g5_0),.clk(gclk));
	jdff dff_A_nhzoLx5Y0_0(.dout(w_dff_A_V4GACXBn5_0),.din(w_dff_A_nhzoLx5Y0_0),.clk(gclk));
	jdff dff_A_V4GACXBn5_0(.dout(w_dff_A_lSlGTfPR1_0),.din(w_dff_A_V4GACXBn5_0),.clk(gclk));
	jdff dff_A_lSlGTfPR1_0(.dout(w_dff_A_ZjRbpGAA7_0),.din(w_dff_A_lSlGTfPR1_0),.clk(gclk));
	jdff dff_A_ZjRbpGAA7_0(.dout(w_dff_A_I9jIwkzI9_0),.din(w_dff_A_ZjRbpGAA7_0),.clk(gclk));
	jdff dff_A_I9jIwkzI9_0(.dout(w_dff_A_RKvvTUuK4_0),.din(w_dff_A_I9jIwkzI9_0),.clk(gclk));
	jdff dff_A_RKvvTUuK4_0(.dout(w_dff_A_q9XvF3KC9_0),.din(w_dff_A_RKvvTUuK4_0),.clk(gclk));
	jdff dff_A_q9XvF3KC9_0(.dout(w_dff_A_9LmIJdwi9_0),.din(w_dff_A_q9XvF3KC9_0),.clk(gclk));
	jdff dff_A_9LmIJdwi9_0(.dout(w_dff_A_v4j9H0yR1_0),.din(w_dff_A_9LmIJdwi9_0),.clk(gclk));
	jdff dff_A_v4j9H0yR1_0(.dout(w_dff_A_yUNbqcnn7_0),.din(w_dff_A_v4j9H0yR1_0),.clk(gclk));
	jdff dff_A_yUNbqcnn7_0(.dout(w_dff_A_saO0hVg49_0),.din(w_dff_A_yUNbqcnn7_0),.clk(gclk));
	jdff dff_A_saO0hVg49_0(.dout(w_dff_A_eX9IBP8q6_0),.din(w_dff_A_saO0hVg49_0),.clk(gclk));
	jdff dff_A_eX9IBP8q6_0(.dout(w_dff_A_G10u59Ef6_0),.din(w_dff_A_eX9IBP8q6_0),.clk(gclk));
	jdff dff_A_G10u59Ef6_0(.dout(w_dff_A_7H2BZrwj8_0),.din(w_dff_A_G10u59Ef6_0),.clk(gclk));
	jdff dff_A_7H2BZrwj8_0(.dout(w_dff_A_7x0Peckt6_0),.din(w_dff_A_7H2BZrwj8_0),.clk(gclk));
	jdff dff_A_7x0Peckt6_0(.dout(w_dff_A_RzZRL4ze5_0),.din(w_dff_A_7x0Peckt6_0),.clk(gclk));
	jdff dff_A_RzZRL4ze5_0(.dout(w_dff_A_rEvuMfh77_0),.din(w_dff_A_RzZRL4ze5_0),.clk(gclk));
	jdff dff_A_rEvuMfh77_0(.dout(w_dff_A_NbQtXbDt9_0),.din(w_dff_A_rEvuMfh77_0),.clk(gclk));
	jdff dff_A_NbQtXbDt9_0(.dout(w_dff_A_rjdsfxNx9_0),.din(w_dff_A_NbQtXbDt9_0),.clk(gclk));
	jdff dff_A_rjdsfxNx9_0(.dout(G810),.din(w_dff_A_rjdsfxNx9_0),.clk(gclk));
	jdff dff_A_hnSczvAh8_1(.dout(w_dff_A_Nbs4hPpN7_0),.din(w_dff_A_hnSczvAh8_1),.clk(gclk));
	jdff dff_A_Nbs4hPpN7_0(.dout(w_dff_A_dO1vHYcD4_0),.din(w_dff_A_Nbs4hPpN7_0),.clk(gclk));
	jdff dff_A_dO1vHYcD4_0(.dout(w_dff_A_7fmWQpVy2_0),.din(w_dff_A_dO1vHYcD4_0),.clk(gclk));
	jdff dff_A_7fmWQpVy2_0(.dout(w_dff_A_SRUYm03Y0_0),.din(w_dff_A_7fmWQpVy2_0),.clk(gclk));
	jdff dff_A_SRUYm03Y0_0(.dout(w_dff_A_6fz4yv274_0),.din(w_dff_A_SRUYm03Y0_0),.clk(gclk));
	jdff dff_A_6fz4yv274_0(.dout(w_dff_A_Vo3Rhqdv9_0),.din(w_dff_A_6fz4yv274_0),.clk(gclk));
	jdff dff_A_Vo3Rhqdv9_0(.dout(w_dff_A_AsIlTvda8_0),.din(w_dff_A_Vo3Rhqdv9_0),.clk(gclk));
	jdff dff_A_AsIlTvda8_0(.dout(w_dff_A_QkjBoflG7_0),.din(w_dff_A_AsIlTvda8_0),.clk(gclk));
	jdff dff_A_QkjBoflG7_0(.dout(w_dff_A_FNHLVngw2_0),.din(w_dff_A_QkjBoflG7_0),.clk(gclk));
	jdff dff_A_FNHLVngw2_0(.dout(w_dff_A_wysyuxlY7_0),.din(w_dff_A_FNHLVngw2_0),.clk(gclk));
	jdff dff_A_wysyuxlY7_0(.dout(w_dff_A_Bda6igyv2_0),.din(w_dff_A_wysyuxlY7_0),.clk(gclk));
	jdff dff_A_Bda6igyv2_0(.dout(w_dff_A_e0DYm3nv3_0),.din(w_dff_A_Bda6igyv2_0),.clk(gclk));
	jdff dff_A_e0DYm3nv3_0(.dout(w_dff_A_dKlb3NNO0_0),.din(w_dff_A_e0DYm3nv3_0),.clk(gclk));
	jdff dff_A_dKlb3NNO0_0(.dout(w_dff_A_GuIx3jf61_0),.din(w_dff_A_dKlb3NNO0_0),.clk(gclk));
	jdff dff_A_GuIx3jf61_0(.dout(w_dff_A_e25GyWQi9_0),.din(w_dff_A_GuIx3jf61_0),.clk(gclk));
	jdff dff_A_e25GyWQi9_0(.dout(w_dff_A_EeSk23ug7_0),.din(w_dff_A_e25GyWQi9_0),.clk(gclk));
	jdff dff_A_EeSk23ug7_0(.dout(w_dff_A_p5YU2Hlm6_0),.din(w_dff_A_EeSk23ug7_0),.clk(gclk));
	jdff dff_A_p5YU2Hlm6_0(.dout(w_dff_A_ZsExShIw2_0),.din(w_dff_A_p5YU2Hlm6_0),.clk(gclk));
	jdff dff_A_ZsExShIw2_0(.dout(w_dff_A_crsdc2Su0_0),.din(w_dff_A_ZsExShIw2_0),.clk(gclk));
	jdff dff_A_crsdc2Su0_0(.dout(w_dff_A_D10H6jgb4_0),.din(w_dff_A_crsdc2Su0_0),.clk(gclk));
	jdff dff_A_D10H6jgb4_0(.dout(w_dff_A_4gOFM9PK3_0),.din(w_dff_A_D10H6jgb4_0),.clk(gclk));
	jdff dff_A_4gOFM9PK3_0(.dout(w_dff_A_iVGrjTjY9_0),.din(w_dff_A_4gOFM9PK3_0),.clk(gclk));
	jdff dff_A_iVGrjTjY9_0(.dout(w_dff_A_4fJQIBYF9_0),.din(w_dff_A_iVGrjTjY9_0),.clk(gclk));
	jdff dff_A_4fJQIBYF9_0(.dout(w_dff_A_cPBR0n1u7_0),.din(w_dff_A_4fJQIBYF9_0),.clk(gclk));
	jdff dff_A_cPBR0n1u7_0(.dout(w_dff_A_v65CSxwt7_0),.din(w_dff_A_cPBR0n1u7_0),.clk(gclk));
	jdff dff_A_v65CSxwt7_0(.dout(w_dff_A_jlREcNb64_0),.din(w_dff_A_v65CSxwt7_0),.clk(gclk));
	jdff dff_A_jlREcNb64_0(.dout(G848),.din(w_dff_A_jlREcNb64_0),.clk(gclk));
	jdff dff_A_E78jADKM5_1(.dout(w_dff_A_Os1MnMJ39_0),.din(w_dff_A_E78jADKM5_1),.clk(gclk));
	jdff dff_A_Os1MnMJ39_0(.dout(w_dff_A_TGsgyyYC2_0),.din(w_dff_A_Os1MnMJ39_0),.clk(gclk));
	jdff dff_A_TGsgyyYC2_0(.dout(w_dff_A_PjcRjUHK5_0),.din(w_dff_A_TGsgyyYC2_0),.clk(gclk));
	jdff dff_A_PjcRjUHK5_0(.dout(w_dff_A_Cxr7ye9u0_0),.din(w_dff_A_PjcRjUHK5_0),.clk(gclk));
	jdff dff_A_Cxr7ye9u0_0(.dout(w_dff_A_oNqNQdg82_0),.din(w_dff_A_Cxr7ye9u0_0),.clk(gclk));
	jdff dff_A_oNqNQdg82_0(.dout(w_dff_A_9dSNBXjp7_0),.din(w_dff_A_oNqNQdg82_0),.clk(gclk));
	jdff dff_A_9dSNBXjp7_0(.dout(w_dff_A_Ow9KclPc6_0),.din(w_dff_A_9dSNBXjp7_0),.clk(gclk));
	jdff dff_A_Ow9KclPc6_0(.dout(w_dff_A_vwhwAJIg3_0),.din(w_dff_A_Ow9KclPc6_0),.clk(gclk));
	jdff dff_A_vwhwAJIg3_0(.dout(w_dff_A_L0eOgLgU8_0),.din(w_dff_A_vwhwAJIg3_0),.clk(gclk));
	jdff dff_A_L0eOgLgU8_0(.dout(w_dff_A_l5MQNVHG6_0),.din(w_dff_A_L0eOgLgU8_0),.clk(gclk));
	jdff dff_A_l5MQNVHG6_0(.dout(w_dff_A_4Y9iyfRX8_0),.din(w_dff_A_l5MQNVHG6_0),.clk(gclk));
	jdff dff_A_4Y9iyfRX8_0(.dout(w_dff_A_LRLQrrPQ7_0),.din(w_dff_A_4Y9iyfRX8_0),.clk(gclk));
	jdff dff_A_LRLQrrPQ7_0(.dout(w_dff_A_IyvFLNBx6_0),.din(w_dff_A_LRLQrrPQ7_0),.clk(gclk));
	jdff dff_A_IyvFLNBx6_0(.dout(w_dff_A_HHMKFOdI6_0),.din(w_dff_A_IyvFLNBx6_0),.clk(gclk));
	jdff dff_A_HHMKFOdI6_0(.dout(w_dff_A_3KZgfooQ1_0),.din(w_dff_A_HHMKFOdI6_0),.clk(gclk));
	jdff dff_A_3KZgfooQ1_0(.dout(w_dff_A_v3IqwvLO4_0),.din(w_dff_A_3KZgfooQ1_0),.clk(gclk));
	jdff dff_A_v3IqwvLO4_0(.dout(w_dff_A_Sopqd15x4_0),.din(w_dff_A_v3IqwvLO4_0),.clk(gclk));
	jdff dff_A_Sopqd15x4_0(.dout(w_dff_A_SjvWJzT00_0),.din(w_dff_A_Sopqd15x4_0),.clk(gclk));
	jdff dff_A_SjvWJzT00_0(.dout(w_dff_A_DNR58lFv5_0),.din(w_dff_A_SjvWJzT00_0),.clk(gclk));
	jdff dff_A_DNR58lFv5_0(.dout(w_dff_A_rOMVEJYf4_0),.din(w_dff_A_DNR58lFv5_0),.clk(gclk));
	jdff dff_A_rOMVEJYf4_0(.dout(w_dff_A_CjUiSqz76_0),.din(w_dff_A_rOMVEJYf4_0),.clk(gclk));
	jdff dff_A_CjUiSqz76_0(.dout(w_dff_A_U74x9EmH6_0),.din(w_dff_A_CjUiSqz76_0),.clk(gclk));
	jdff dff_A_U74x9EmH6_0(.dout(w_dff_A_yYU3lUVb7_0),.din(w_dff_A_U74x9EmH6_0),.clk(gclk));
	jdff dff_A_yYU3lUVb7_0(.dout(w_dff_A_kucTH1T92_0),.din(w_dff_A_yYU3lUVb7_0),.clk(gclk));
	jdff dff_A_kucTH1T92_0(.dout(w_dff_A_5ygJ0C591_0),.din(w_dff_A_kucTH1T92_0),.clk(gclk));
	jdff dff_A_5ygJ0C591_0(.dout(w_dff_A_nqMgHf3K7_0),.din(w_dff_A_5ygJ0C591_0),.clk(gclk));
	jdff dff_A_nqMgHf3K7_0(.dout(G849),.din(w_dff_A_nqMgHf3K7_0),.clk(gclk));
	jdff dff_A_AVwe8LZD9_1(.dout(w_dff_A_PO7tgq5D9_0),.din(w_dff_A_AVwe8LZD9_1),.clk(gclk));
	jdff dff_A_PO7tgq5D9_0(.dout(w_dff_A_8MCDdNcp8_0),.din(w_dff_A_PO7tgq5D9_0),.clk(gclk));
	jdff dff_A_8MCDdNcp8_0(.dout(w_dff_A_cmQHrnNI5_0),.din(w_dff_A_8MCDdNcp8_0),.clk(gclk));
	jdff dff_A_cmQHrnNI5_0(.dout(w_dff_A_5PdJUxCH0_0),.din(w_dff_A_cmQHrnNI5_0),.clk(gclk));
	jdff dff_A_5PdJUxCH0_0(.dout(w_dff_A_9WfNcnOA4_0),.din(w_dff_A_5PdJUxCH0_0),.clk(gclk));
	jdff dff_A_9WfNcnOA4_0(.dout(w_dff_A_6UlGFyej0_0),.din(w_dff_A_9WfNcnOA4_0),.clk(gclk));
	jdff dff_A_6UlGFyej0_0(.dout(w_dff_A_IzSs48DS6_0),.din(w_dff_A_6UlGFyej0_0),.clk(gclk));
	jdff dff_A_IzSs48DS6_0(.dout(w_dff_A_nyvPgYcF2_0),.din(w_dff_A_IzSs48DS6_0),.clk(gclk));
	jdff dff_A_nyvPgYcF2_0(.dout(w_dff_A_teiwgbjW7_0),.din(w_dff_A_nyvPgYcF2_0),.clk(gclk));
	jdff dff_A_teiwgbjW7_0(.dout(w_dff_A_KGjswTrX2_0),.din(w_dff_A_teiwgbjW7_0),.clk(gclk));
	jdff dff_A_KGjswTrX2_0(.dout(w_dff_A_i2u3Glm31_0),.din(w_dff_A_KGjswTrX2_0),.clk(gclk));
	jdff dff_A_i2u3Glm31_0(.dout(w_dff_A_XLqpSjFl1_0),.din(w_dff_A_i2u3Glm31_0),.clk(gclk));
	jdff dff_A_XLqpSjFl1_0(.dout(w_dff_A_UcAqKqU75_0),.din(w_dff_A_XLqpSjFl1_0),.clk(gclk));
	jdff dff_A_UcAqKqU75_0(.dout(w_dff_A_cp0D2UbL9_0),.din(w_dff_A_UcAqKqU75_0),.clk(gclk));
	jdff dff_A_cp0D2UbL9_0(.dout(w_dff_A_1BBBmYvz5_0),.din(w_dff_A_cp0D2UbL9_0),.clk(gclk));
	jdff dff_A_1BBBmYvz5_0(.dout(w_dff_A_jCbprpTt4_0),.din(w_dff_A_1BBBmYvz5_0),.clk(gclk));
	jdff dff_A_jCbprpTt4_0(.dout(w_dff_A_jvOE0Bcl4_0),.din(w_dff_A_jCbprpTt4_0),.clk(gclk));
	jdff dff_A_jvOE0Bcl4_0(.dout(w_dff_A_3Hmrvuz22_0),.din(w_dff_A_jvOE0Bcl4_0),.clk(gclk));
	jdff dff_A_3Hmrvuz22_0(.dout(w_dff_A_mrvFK7Rw6_0),.din(w_dff_A_3Hmrvuz22_0),.clk(gclk));
	jdff dff_A_mrvFK7Rw6_0(.dout(w_dff_A_gFFJRjsn5_0),.din(w_dff_A_mrvFK7Rw6_0),.clk(gclk));
	jdff dff_A_gFFJRjsn5_0(.dout(w_dff_A_gCupuTys4_0),.din(w_dff_A_gFFJRjsn5_0),.clk(gclk));
	jdff dff_A_gCupuTys4_0(.dout(w_dff_A_hWfQPs7a0_0),.din(w_dff_A_gCupuTys4_0),.clk(gclk));
	jdff dff_A_hWfQPs7a0_0(.dout(w_dff_A_TxPodgNl0_0),.din(w_dff_A_hWfQPs7a0_0),.clk(gclk));
	jdff dff_A_TxPodgNl0_0(.dout(w_dff_A_QFyiUs6Q1_0),.din(w_dff_A_TxPodgNl0_0),.clk(gclk));
	jdff dff_A_QFyiUs6Q1_0(.dout(w_dff_A_EAuEEzF05_0),.din(w_dff_A_QFyiUs6Q1_0),.clk(gclk));
	jdff dff_A_EAuEEzF05_0(.dout(w_dff_A_xp1vCgnp3_0),.din(w_dff_A_EAuEEzF05_0),.clk(gclk));
	jdff dff_A_xp1vCgnp3_0(.dout(G850),.din(w_dff_A_xp1vCgnp3_0),.clk(gclk));
	jdff dff_A_8yW8rYSC0_1(.dout(w_dff_A_jWaUtTT72_0),.din(w_dff_A_8yW8rYSC0_1),.clk(gclk));
	jdff dff_A_jWaUtTT72_0(.dout(w_dff_A_d8CCqeeI9_0),.din(w_dff_A_jWaUtTT72_0),.clk(gclk));
	jdff dff_A_d8CCqeeI9_0(.dout(w_dff_A_7ZjhNA046_0),.din(w_dff_A_d8CCqeeI9_0),.clk(gclk));
	jdff dff_A_7ZjhNA046_0(.dout(w_dff_A_cYXe9Txc3_0),.din(w_dff_A_7ZjhNA046_0),.clk(gclk));
	jdff dff_A_cYXe9Txc3_0(.dout(w_dff_A_5zEpCGD84_0),.din(w_dff_A_cYXe9Txc3_0),.clk(gclk));
	jdff dff_A_5zEpCGD84_0(.dout(w_dff_A_SrS0fT2L4_0),.din(w_dff_A_5zEpCGD84_0),.clk(gclk));
	jdff dff_A_SrS0fT2L4_0(.dout(w_dff_A_CXkKXAno0_0),.din(w_dff_A_SrS0fT2L4_0),.clk(gclk));
	jdff dff_A_CXkKXAno0_0(.dout(w_dff_A_OFEwH6rW2_0),.din(w_dff_A_CXkKXAno0_0),.clk(gclk));
	jdff dff_A_OFEwH6rW2_0(.dout(w_dff_A_MmHuy6gC5_0),.din(w_dff_A_OFEwH6rW2_0),.clk(gclk));
	jdff dff_A_MmHuy6gC5_0(.dout(w_dff_A_YaAtkiWq9_0),.din(w_dff_A_MmHuy6gC5_0),.clk(gclk));
	jdff dff_A_YaAtkiWq9_0(.dout(w_dff_A_Ww66n3773_0),.din(w_dff_A_YaAtkiWq9_0),.clk(gclk));
	jdff dff_A_Ww66n3773_0(.dout(w_dff_A_SUUo5uWi6_0),.din(w_dff_A_Ww66n3773_0),.clk(gclk));
	jdff dff_A_SUUo5uWi6_0(.dout(w_dff_A_M7kAZ2C54_0),.din(w_dff_A_SUUo5uWi6_0),.clk(gclk));
	jdff dff_A_M7kAZ2C54_0(.dout(w_dff_A_9D3l8rqA9_0),.din(w_dff_A_M7kAZ2C54_0),.clk(gclk));
	jdff dff_A_9D3l8rqA9_0(.dout(w_dff_A_ZAOREYlY3_0),.din(w_dff_A_9D3l8rqA9_0),.clk(gclk));
	jdff dff_A_ZAOREYlY3_0(.dout(w_dff_A_dQvkqOqn5_0),.din(w_dff_A_ZAOREYlY3_0),.clk(gclk));
	jdff dff_A_dQvkqOqn5_0(.dout(w_dff_A_AjiYy8BX4_0),.din(w_dff_A_dQvkqOqn5_0),.clk(gclk));
	jdff dff_A_AjiYy8BX4_0(.dout(w_dff_A_KLBflqsX4_0),.din(w_dff_A_AjiYy8BX4_0),.clk(gclk));
	jdff dff_A_KLBflqsX4_0(.dout(w_dff_A_SsSlhH227_0),.din(w_dff_A_KLBflqsX4_0),.clk(gclk));
	jdff dff_A_SsSlhH227_0(.dout(w_dff_A_7uxBLpPp4_0),.din(w_dff_A_SsSlhH227_0),.clk(gclk));
	jdff dff_A_7uxBLpPp4_0(.dout(w_dff_A_CObSADYm1_0),.din(w_dff_A_7uxBLpPp4_0),.clk(gclk));
	jdff dff_A_CObSADYm1_0(.dout(w_dff_A_WIv7iNS84_0),.din(w_dff_A_CObSADYm1_0),.clk(gclk));
	jdff dff_A_WIv7iNS84_0(.dout(w_dff_A_iSoCOx0I5_0),.din(w_dff_A_WIv7iNS84_0),.clk(gclk));
	jdff dff_A_iSoCOx0I5_0(.dout(w_dff_A_lRdT4CJ46_0),.din(w_dff_A_iSoCOx0I5_0),.clk(gclk));
	jdff dff_A_lRdT4CJ46_0(.dout(w_dff_A_ekRwoShX9_0),.din(w_dff_A_lRdT4CJ46_0),.clk(gclk));
	jdff dff_A_ekRwoShX9_0(.dout(w_dff_A_5JxwWsO02_0),.din(w_dff_A_ekRwoShX9_0),.clk(gclk));
	jdff dff_A_5JxwWsO02_0(.dout(G851),.din(w_dff_A_5JxwWsO02_0),.clk(gclk));
	jdff dff_A_il5gzRQ12_2(.dout(w_dff_A_riEweXVy7_0),.din(w_dff_A_il5gzRQ12_2),.clk(gclk));
	jdff dff_A_riEweXVy7_0(.dout(w_dff_A_JkSreVU53_0),.din(w_dff_A_riEweXVy7_0),.clk(gclk));
	jdff dff_A_JkSreVU53_0(.dout(w_dff_A_5hPsmtub3_0),.din(w_dff_A_JkSreVU53_0),.clk(gclk));
	jdff dff_A_5hPsmtub3_0(.dout(w_dff_A_lc3etMdM7_0),.din(w_dff_A_5hPsmtub3_0),.clk(gclk));
	jdff dff_A_lc3etMdM7_0(.dout(w_dff_A_eIeDO3ks3_0),.din(w_dff_A_lc3etMdM7_0),.clk(gclk));
	jdff dff_A_eIeDO3ks3_0(.dout(w_dff_A_jIV2dcNj9_0),.din(w_dff_A_eIeDO3ks3_0),.clk(gclk));
	jdff dff_A_jIV2dcNj9_0(.dout(w_dff_A_rTs8NITW9_0),.din(w_dff_A_jIV2dcNj9_0),.clk(gclk));
	jdff dff_A_rTs8NITW9_0(.dout(w_dff_A_n4bOUqh09_0),.din(w_dff_A_rTs8NITW9_0),.clk(gclk));
	jdff dff_A_n4bOUqh09_0(.dout(w_dff_A_ytIRBICk7_0),.din(w_dff_A_n4bOUqh09_0),.clk(gclk));
	jdff dff_A_ytIRBICk7_0(.dout(w_dff_A_7Ptvir2R4_0),.din(w_dff_A_ytIRBICk7_0),.clk(gclk));
	jdff dff_A_7Ptvir2R4_0(.dout(w_dff_A_h0wYJW9n1_0),.din(w_dff_A_7Ptvir2R4_0),.clk(gclk));
	jdff dff_A_h0wYJW9n1_0(.dout(w_dff_A_Mxj305Ms9_0),.din(w_dff_A_h0wYJW9n1_0),.clk(gclk));
	jdff dff_A_Mxj305Ms9_0(.dout(w_dff_A_wlrlNyfu2_0),.din(w_dff_A_Mxj305Ms9_0),.clk(gclk));
	jdff dff_A_wlrlNyfu2_0(.dout(w_dff_A_jxiveFpg2_0),.din(w_dff_A_wlrlNyfu2_0),.clk(gclk));
	jdff dff_A_jxiveFpg2_0(.dout(w_dff_A_W1S3G9PT5_0),.din(w_dff_A_jxiveFpg2_0),.clk(gclk));
	jdff dff_A_W1S3G9PT5_0(.dout(w_dff_A_e1JTv2eI4_0),.din(w_dff_A_W1S3G9PT5_0),.clk(gclk));
	jdff dff_A_e1JTv2eI4_0(.dout(w_dff_A_zJMi3bZE7_0),.din(w_dff_A_e1JTv2eI4_0),.clk(gclk));
	jdff dff_A_zJMi3bZE7_0(.dout(w_dff_A_ZLbLw1AG4_0),.din(w_dff_A_zJMi3bZE7_0),.clk(gclk));
	jdff dff_A_ZLbLw1AG4_0(.dout(w_dff_A_tRbkvvAZ2_0),.din(w_dff_A_ZLbLw1AG4_0),.clk(gclk));
	jdff dff_A_tRbkvvAZ2_0(.dout(w_dff_A_HGapMj9y7_0),.din(w_dff_A_tRbkvvAZ2_0),.clk(gclk));
	jdff dff_A_HGapMj9y7_0(.dout(w_dff_A_ih1Xr53m3_0),.din(w_dff_A_HGapMj9y7_0),.clk(gclk));
	jdff dff_A_ih1Xr53m3_0(.dout(w_dff_A_IuEaUu7G4_0),.din(w_dff_A_ih1Xr53m3_0),.clk(gclk));
	jdff dff_A_IuEaUu7G4_0(.dout(w_dff_A_OUk7o9UW8_0),.din(w_dff_A_IuEaUu7G4_0),.clk(gclk));
	jdff dff_A_OUk7o9UW8_0(.dout(w_dff_A_OUkKcXKL4_0),.din(w_dff_A_OUk7o9UW8_0),.clk(gclk));
	jdff dff_A_OUkKcXKL4_0(.dout(w_dff_A_2XUhHR2f1_0),.din(w_dff_A_OUkKcXKL4_0),.clk(gclk));
	jdff dff_A_2XUhHR2f1_0(.dout(w_dff_A_QWhXvLgw5_0),.din(w_dff_A_2XUhHR2f1_0),.clk(gclk));
	jdff dff_A_QWhXvLgw5_0(.dout(G634),.din(w_dff_A_QWhXvLgw5_0),.clk(gclk));
	jdff dff_A_5yZAzLY28_2(.dout(w_dff_A_tUbXQn0z4_0),.din(w_dff_A_5yZAzLY28_2),.clk(gclk));
	jdff dff_A_tUbXQn0z4_0(.dout(w_dff_A_fz4Jpv666_0),.din(w_dff_A_tUbXQn0z4_0),.clk(gclk));
	jdff dff_A_fz4Jpv666_0(.dout(w_dff_A_8nazHNcJ1_0),.din(w_dff_A_fz4Jpv666_0),.clk(gclk));
	jdff dff_A_8nazHNcJ1_0(.dout(w_dff_A_uhe5p8Mq8_0),.din(w_dff_A_8nazHNcJ1_0),.clk(gclk));
	jdff dff_A_uhe5p8Mq8_0(.dout(w_dff_A_Tkv499YQ4_0),.din(w_dff_A_uhe5p8Mq8_0),.clk(gclk));
	jdff dff_A_Tkv499YQ4_0(.dout(w_dff_A_5olupmWL9_0),.din(w_dff_A_Tkv499YQ4_0),.clk(gclk));
	jdff dff_A_5olupmWL9_0(.dout(w_dff_A_M2ax1Wdn6_0),.din(w_dff_A_5olupmWL9_0),.clk(gclk));
	jdff dff_A_M2ax1Wdn6_0(.dout(w_dff_A_TzNUu3ZK6_0),.din(w_dff_A_M2ax1Wdn6_0),.clk(gclk));
	jdff dff_A_TzNUu3ZK6_0(.dout(w_dff_A_wav0QNfw5_0),.din(w_dff_A_TzNUu3ZK6_0),.clk(gclk));
	jdff dff_A_wav0QNfw5_0(.dout(w_dff_A_ulKNR54U8_0),.din(w_dff_A_wav0QNfw5_0),.clk(gclk));
	jdff dff_A_ulKNR54U8_0(.dout(w_dff_A_7cjmnhhj8_0),.din(w_dff_A_ulKNR54U8_0),.clk(gclk));
	jdff dff_A_7cjmnhhj8_0(.dout(w_dff_A_wzXXIedh6_0),.din(w_dff_A_7cjmnhhj8_0),.clk(gclk));
	jdff dff_A_wzXXIedh6_0(.dout(w_dff_A_2ojMxaAV4_0),.din(w_dff_A_wzXXIedh6_0),.clk(gclk));
	jdff dff_A_2ojMxaAV4_0(.dout(w_dff_A_mwMcFTOK1_0),.din(w_dff_A_2ojMxaAV4_0),.clk(gclk));
	jdff dff_A_mwMcFTOK1_0(.dout(w_dff_A_PoDZDGgX1_0),.din(w_dff_A_mwMcFTOK1_0),.clk(gclk));
	jdff dff_A_PoDZDGgX1_0(.dout(w_dff_A_stgsCdxf9_0),.din(w_dff_A_PoDZDGgX1_0),.clk(gclk));
	jdff dff_A_stgsCdxf9_0(.dout(w_dff_A_5dYTDES71_0),.din(w_dff_A_stgsCdxf9_0),.clk(gclk));
	jdff dff_A_5dYTDES71_0(.dout(w_dff_A_XDuiwhjT6_0),.din(w_dff_A_5dYTDES71_0),.clk(gclk));
	jdff dff_A_XDuiwhjT6_0(.dout(w_dff_A_xV9CNt115_0),.din(w_dff_A_XDuiwhjT6_0),.clk(gclk));
	jdff dff_A_xV9CNt115_0(.dout(w_dff_A_0LnJw27W4_0),.din(w_dff_A_xV9CNt115_0),.clk(gclk));
	jdff dff_A_0LnJw27W4_0(.dout(w_dff_A_G1G1MDan4_0),.din(w_dff_A_0LnJw27W4_0),.clk(gclk));
	jdff dff_A_G1G1MDan4_0(.dout(w_dff_A_7TpO1Pdn4_0),.din(w_dff_A_G1G1MDan4_0),.clk(gclk));
	jdff dff_A_7TpO1Pdn4_0(.dout(w_dff_A_g0FEQjEd5_0),.din(w_dff_A_7TpO1Pdn4_0),.clk(gclk));
	jdff dff_A_g0FEQjEd5_0(.dout(w_dff_A_xZlzbVAn2_0),.din(w_dff_A_g0FEQjEd5_0),.clk(gclk));
	jdff dff_A_xZlzbVAn2_0(.dout(w_dff_A_HI1Rh4ot5_0),.din(w_dff_A_xZlzbVAn2_0),.clk(gclk));
	jdff dff_A_HI1Rh4ot5_0(.dout(G815),.din(w_dff_A_HI1Rh4ot5_0),.clk(gclk));
	jdff dff_A_Dfh0sref6_2(.dout(w_dff_A_xwcyPH0a3_0),.din(w_dff_A_Dfh0sref6_2),.clk(gclk));
	jdff dff_A_xwcyPH0a3_0(.dout(w_dff_A_pSo1dmi77_0),.din(w_dff_A_xwcyPH0a3_0),.clk(gclk));
	jdff dff_A_pSo1dmi77_0(.dout(w_dff_A_DE5Y2rea6_0),.din(w_dff_A_pSo1dmi77_0),.clk(gclk));
	jdff dff_A_DE5Y2rea6_0(.dout(w_dff_A_IkKvnjdu1_0),.din(w_dff_A_DE5Y2rea6_0),.clk(gclk));
	jdff dff_A_IkKvnjdu1_0(.dout(w_dff_A_zaEoPNvZ5_0),.din(w_dff_A_IkKvnjdu1_0),.clk(gclk));
	jdff dff_A_zaEoPNvZ5_0(.dout(w_dff_A_U0d9brpo2_0),.din(w_dff_A_zaEoPNvZ5_0),.clk(gclk));
	jdff dff_A_U0d9brpo2_0(.dout(w_dff_A_pPlzUs7g2_0),.din(w_dff_A_U0d9brpo2_0),.clk(gclk));
	jdff dff_A_pPlzUs7g2_0(.dout(w_dff_A_9jHMRoOV9_0),.din(w_dff_A_pPlzUs7g2_0),.clk(gclk));
	jdff dff_A_9jHMRoOV9_0(.dout(w_dff_A_YVRK1qKE8_0),.din(w_dff_A_9jHMRoOV9_0),.clk(gclk));
	jdff dff_A_YVRK1qKE8_0(.dout(w_dff_A_Oyf7yWf86_0),.din(w_dff_A_YVRK1qKE8_0),.clk(gclk));
	jdff dff_A_Oyf7yWf86_0(.dout(w_dff_A_7QbbRmnw9_0),.din(w_dff_A_Oyf7yWf86_0),.clk(gclk));
	jdff dff_A_7QbbRmnw9_0(.dout(w_dff_A_HPGJIieo8_0),.din(w_dff_A_7QbbRmnw9_0),.clk(gclk));
	jdff dff_A_HPGJIieo8_0(.dout(w_dff_A_5BKg6cgW9_0),.din(w_dff_A_HPGJIieo8_0),.clk(gclk));
	jdff dff_A_5BKg6cgW9_0(.dout(w_dff_A_x8z88Exm7_0),.din(w_dff_A_5BKg6cgW9_0),.clk(gclk));
	jdff dff_A_x8z88Exm7_0(.dout(w_dff_A_gsCFFxp63_0),.din(w_dff_A_x8z88Exm7_0),.clk(gclk));
	jdff dff_A_gsCFFxp63_0(.dout(w_dff_A_tHM9M5NA1_0),.din(w_dff_A_gsCFFxp63_0),.clk(gclk));
	jdff dff_A_tHM9M5NA1_0(.dout(w_dff_A_1SOcq7Q70_0),.din(w_dff_A_tHM9M5NA1_0),.clk(gclk));
	jdff dff_A_1SOcq7Q70_0(.dout(w_dff_A_S2q6Y5NH2_0),.din(w_dff_A_1SOcq7Q70_0),.clk(gclk));
	jdff dff_A_S2q6Y5NH2_0(.dout(w_dff_A_IdBpOYNS3_0),.din(w_dff_A_S2q6Y5NH2_0),.clk(gclk));
	jdff dff_A_IdBpOYNS3_0(.dout(w_dff_A_ROCzrkRF2_0),.din(w_dff_A_IdBpOYNS3_0),.clk(gclk));
	jdff dff_A_ROCzrkRF2_0(.dout(w_dff_A_QPo5Ne8z2_0),.din(w_dff_A_ROCzrkRF2_0),.clk(gclk));
	jdff dff_A_QPo5Ne8z2_0(.dout(w_dff_A_7u2g0qVo5_0),.din(w_dff_A_QPo5Ne8z2_0),.clk(gclk));
	jdff dff_A_7u2g0qVo5_0(.dout(w_dff_A_ocCrRWin3_0),.din(w_dff_A_7u2g0qVo5_0),.clk(gclk));
	jdff dff_A_ocCrRWin3_0(.dout(w_dff_A_FrZTDCMc0_0),.din(w_dff_A_ocCrRWin3_0),.clk(gclk));
	jdff dff_A_FrZTDCMc0_0(.dout(w_dff_A_WsxsxKl22_0),.din(w_dff_A_FrZTDCMc0_0),.clk(gclk));
	jdff dff_A_WsxsxKl22_0(.dout(G845),.din(w_dff_A_WsxsxKl22_0),.clk(gclk));
	jdff dff_A_9IakLXyU2_1(.dout(w_dff_A_rufGJAmd1_0),.din(w_dff_A_9IakLXyU2_1),.clk(gclk));
	jdff dff_A_rufGJAmd1_0(.dout(w_dff_A_QmbBvWQC0_0),.din(w_dff_A_rufGJAmd1_0),.clk(gclk));
	jdff dff_A_QmbBvWQC0_0(.dout(w_dff_A_keuBOLpZ7_0),.din(w_dff_A_QmbBvWQC0_0),.clk(gclk));
	jdff dff_A_keuBOLpZ7_0(.dout(w_dff_A_z2hslrWB4_0),.din(w_dff_A_keuBOLpZ7_0),.clk(gclk));
	jdff dff_A_z2hslrWB4_0(.dout(w_dff_A_RSMFuCRy1_0),.din(w_dff_A_z2hslrWB4_0),.clk(gclk));
	jdff dff_A_RSMFuCRy1_0(.dout(w_dff_A_63x1gn8F8_0),.din(w_dff_A_RSMFuCRy1_0),.clk(gclk));
	jdff dff_A_63x1gn8F8_0(.dout(w_dff_A_MuA5trTl3_0),.din(w_dff_A_63x1gn8F8_0),.clk(gclk));
	jdff dff_A_MuA5trTl3_0(.dout(w_dff_A_RHLYyt9m0_0),.din(w_dff_A_MuA5trTl3_0),.clk(gclk));
	jdff dff_A_RHLYyt9m0_0(.dout(w_dff_A_hVrvFaWl3_0),.din(w_dff_A_RHLYyt9m0_0),.clk(gclk));
	jdff dff_A_hVrvFaWl3_0(.dout(w_dff_A_zJA8MhWX4_0),.din(w_dff_A_hVrvFaWl3_0),.clk(gclk));
	jdff dff_A_zJA8MhWX4_0(.dout(w_dff_A_pmT97wB52_0),.din(w_dff_A_zJA8MhWX4_0),.clk(gclk));
	jdff dff_A_pmT97wB52_0(.dout(w_dff_A_reTcRdcR2_0),.din(w_dff_A_pmT97wB52_0),.clk(gclk));
	jdff dff_A_reTcRdcR2_0(.dout(w_dff_A_0fu0XvWa2_0),.din(w_dff_A_reTcRdcR2_0),.clk(gclk));
	jdff dff_A_0fu0XvWa2_0(.dout(w_dff_A_sXXYdx8N5_0),.din(w_dff_A_0fu0XvWa2_0),.clk(gclk));
	jdff dff_A_sXXYdx8N5_0(.dout(w_dff_A_y8muQaPw3_0),.din(w_dff_A_sXXYdx8N5_0),.clk(gclk));
	jdff dff_A_y8muQaPw3_0(.dout(w_dff_A_bel5rW7I8_0),.din(w_dff_A_y8muQaPw3_0),.clk(gclk));
	jdff dff_A_bel5rW7I8_0(.dout(w_dff_A_vL1ZCH203_0),.din(w_dff_A_bel5rW7I8_0),.clk(gclk));
	jdff dff_A_vL1ZCH203_0(.dout(w_dff_A_o40Ra72I2_0),.din(w_dff_A_vL1ZCH203_0),.clk(gclk));
	jdff dff_A_o40Ra72I2_0(.dout(w_dff_A_VL8Ea4yE8_0),.din(w_dff_A_o40Ra72I2_0),.clk(gclk));
	jdff dff_A_VL8Ea4yE8_0(.dout(w_dff_A_S5lDYPbk5_0),.din(w_dff_A_VL8Ea4yE8_0),.clk(gclk));
	jdff dff_A_S5lDYPbk5_0(.dout(w_dff_A_NiYBZsHm1_0),.din(w_dff_A_S5lDYPbk5_0),.clk(gclk));
	jdff dff_A_NiYBZsHm1_0(.dout(w_dff_A_HC3Dwmbt3_0),.din(w_dff_A_NiYBZsHm1_0),.clk(gclk));
	jdff dff_A_HC3Dwmbt3_0(.dout(w_dff_A_d6EH0yu26_0),.din(w_dff_A_HC3Dwmbt3_0),.clk(gclk));
	jdff dff_A_d6EH0yu26_0(.dout(w_dff_A_MORjDeJV8_0),.din(w_dff_A_d6EH0yu26_0),.clk(gclk));
	jdff dff_A_MORjDeJV8_0(.dout(w_dff_A_w8v0m3Q02_0),.din(w_dff_A_MORjDeJV8_0),.clk(gclk));
	jdff dff_A_w8v0m3Q02_0(.dout(G847),.din(w_dff_A_w8v0m3Q02_0),.clk(gclk));
	jdff dff_A_7IidBGnj0_1(.dout(w_dff_A_4LFar5BP2_0),.din(w_dff_A_7IidBGnj0_1),.clk(gclk));
	jdff dff_A_4LFar5BP2_0(.dout(w_dff_A_4MZBsiiP3_0),.din(w_dff_A_4LFar5BP2_0),.clk(gclk));
	jdff dff_A_4MZBsiiP3_0(.dout(w_dff_A_6GtuHvx63_0),.din(w_dff_A_4MZBsiiP3_0),.clk(gclk));
	jdff dff_A_6GtuHvx63_0(.dout(w_dff_A_NozBF5TA0_0),.din(w_dff_A_6GtuHvx63_0),.clk(gclk));
	jdff dff_A_NozBF5TA0_0(.dout(w_dff_A_6bIEeuAb8_0),.din(w_dff_A_NozBF5TA0_0),.clk(gclk));
	jdff dff_A_6bIEeuAb8_0(.dout(w_dff_A_MRTMuoUf8_0),.din(w_dff_A_6bIEeuAb8_0),.clk(gclk));
	jdff dff_A_MRTMuoUf8_0(.dout(w_dff_A_kJ6pB0zZ7_0),.din(w_dff_A_MRTMuoUf8_0),.clk(gclk));
	jdff dff_A_kJ6pB0zZ7_0(.dout(w_dff_A_zdH2Qkq25_0),.din(w_dff_A_kJ6pB0zZ7_0),.clk(gclk));
	jdff dff_A_zdH2Qkq25_0(.dout(w_dff_A_W2HfM4Lo4_0),.din(w_dff_A_zdH2Qkq25_0),.clk(gclk));
	jdff dff_A_W2HfM4Lo4_0(.dout(w_dff_A_y4xyVCHZ3_0),.din(w_dff_A_W2HfM4Lo4_0),.clk(gclk));
	jdff dff_A_y4xyVCHZ3_0(.dout(w_dff_A_F34MBWH74_0),.din(w_dff_A_y4xyVCHZ3_0),.clk(gclk));
	jdff dff_A_F34MBWH74_0(.dout(w_dff_A_71TPG1et7_0),.din(w_dff_A_F34MBWH74_0),.clk(gclk));
	jdff dff_A_71TPG1et7_0(.dout(w_dff_A_oLgXCcvY8_0),.din(w_dff_A_71TPG1et7_0),.clk(gclk));
	jdff dff_A_oLgXCcvY8_0(.dout(w_dff_A_zoFyNcDR9_0),.din(w_dff_A_oLgXCcvY8_0),.clk(gclk));
	jdff dff_A_zoFyNcDR9_0(.dout(w_dff_A_VkvV2lve3_0),.din(w_dff_A_zoFyNcDR9_0),.clk(gclk));
	jdff dff_A_VkvV2lve3_0(.dout(w_dff_A_pb3KQtoy4_0),.din(w_dff_A_VkvV2lve3_0),.clk(gclk));
	jdff dff_A_pb3KQtoy4_0(.dout(w_dff_A_HxOIOknW6_0),.din(w_dff_A_pb3KQtoy4_0),.clk(gclk));
	jdff dff_A_HxOIOknW6_0(.dout(w_dff_A_nPf0dmm79_0),.din(w_dff_A_HxOIOknW6_0),.clk(gclk));
	jdff dff_A_nPf0dmm79_0(.dout(w_dff_A_Ae5euWha8_0),.din(w_dff_A_nPf0dmm79_0),.clk(gclk));
	jdff dff_A_Ae5euWha8_0(.dout(w_dff_A_kjlEW1Um4_0),.din(w_dff_A_Ae5euWha8_0),.clk(gclk));
	jdff dff_A_kjlEW1Um4_0(.dout(w_dff_A_aEHGnoD38_0),.din(w_dff_A_kjlEW1Um4_0),.clk(gclk));
	jdff dff_A_aEHGnoD38_0(.dout(w_dff_A_x2BWPgim7_0),.din(w_dff_A_aEHGnoD38_0),.clk(gclk));
	jdff dff_A_x2BWPgim7_0(.dout(w_dff_A_54R3MjDQ5_0),.din(w_dff_A_x2BWPgim7_0),.clk(gclk));
	jdff dff_A_54R3MjDQ5_0(.dout(w_dff_A_2c6SKHDE7_0),.din(w_dff_A_54R3MjDQ5_0),.clk(gclk));
	jdff dff_A_2c6SKHDE7_0(.dout(w_dff_A_b28cF2pe2_0),.din(w_dff_A_2c6SKHDE7_0),.clk(gclk));
	jdff dff_A_b28cF2pe2_0(.dout(w_dff_A_jchro18i2_0),.din(w_dff_A_b28cF2pe2_0),.clk(gclk));
	jdff dff_A_jchro18i2_0(.dout(w_dff_A_zHRMXs3k8_0),.din(w_dff_A_jchro18i2_0),.clk(gclk));
	jdff dff_A_zHRMXs3k8_0(.dout(G926),.din(w_dff_A_zHRMXs3k8_0),.clk(gclk));
	jdff dff_A_hGDXCrDc6_1(.dout(w_dff_A_7iFwTMbE4_0),.din(w_dff_A_hGDXCrDc6_1),.clk(gclk));
	jdff dff_A_7iFwTMbE4_0(.dout(w_dff_A_pweeR05v0_0),.din(w_dff_A_7iFwTMbE4_0),.clk(gclk));
	jdff dff_A_pweeR05v0_0(.dout(w_dff_A_jsl0Mbs59_0),.din(w_dff_A_pweeR05v0_0),.clk(gclk));
	jdff dff_A_jsl0Mbs59_0(.dout(w_dff_A_MlmfdpkD6_0),.din(w_dff_A_jsl0Mbs59_0),.clk(gclk));
	jdff dff_A_MlmfdpkD6_0(.dout(w_dff_A_VzBw1px09_0),.din(w_dff_A_MlmfdpkD6_0),.clk(gclk));
	jdff dff_A_VzBw1px09_0(.dout(w_dff_A_6UL5Hx0P9_0),.din(w_dff_A_VzBw1px09_0),.clk(gclk));
	jdff dff_A_6UL5Hx0P9_0(.dout(w_dff_A_wIHqwPWr9_0),.din(w_dff_A_6UL5Hx0P9_0),.clk(gclk));
	jdff dff_A_wIHqwPWr9_0(.dout(w_dff_A_k9YT6nXx2_0),.din(w_dff_A_wIHqwPWr9_0),.clk(gclk));
	jdff dff_A_k9YT6nXx2_0(.dout(w_dff_A_5xY0XIJW0_0),.din(w_dff_A_k9YT6nXx2_0),.clk(gclk));
	jdff dff_A_5xY0XIJW0_0(.dout(w_dff_A_XnNjdOzZ6_0),.din(w_dff_A_5xY0XIJW0_0),.clk(gclk));
	jdff dff_A_XnNjdOzZ6_0(.dout(w_dff_A_Se769BEq1_0),.din(w_dff_A_XnNjdOzZ6_0),.clk(gclk));
	jdff dff_A_Se769BEq1_0(.dout(w_dff_A_ddGZYwbp8_0),.din(w_dff_A_Se769BEq1_0),.clk(gclk));
	jdff dff_A_ddGZYwbp8_0(.dout(w_dff_A_MSemvxeP2_0),.din(w_dff_A_ddGZYwbp8_0),.clk(gclk));
	jdff dff_A_MSemvxeP2_0(.dout(w_dff_A_Kd6IDemI2_0),.din(w_dff_A_MSemvxeP2_0),.clk(gclk));
	jdff dff_A_Kd6IDemI2_0(.dout(w_dff_A_PJCISWQ25_0),.din(w_dff_A_Kd6IDemI2_0),.clk(gclk));
	jdff dff_A_PJCISWQ25_0(.dout(w_dff_A_Yr6uya6r5_0),.din(w_dff_A_PJCISWQ25_0),.clk(gclk));
	jdff dff_A_Yr6uya6r5_0(.dout(w_dff_A_tmzvb0Nv3_0),.din(w_dff_A_Yr6uya6r5_0),.clk(gclk));
	jdff dff_A_tmzvb0Nv3_0(.dout(w_dff_A_09sHDbOn8_0),.din(w_dff_A_tmzvb0Nv3_0),.clk(gclk));
	jdff dff_A_09sHDbOn8_0(.dout(w_dff_A_u5TMods47_0),.din(w_dff_A_09sHDbOn8_0),.clk(gclk));
	jdff dff_A_u5TMods47_0(.dout(w_dff_A_EKsT2u6v4_0),.din(w_dff_A_u5TMods47_0),.clk(gclk));
	jdff dff_A_EKsT2u6v4_0(.dout(w_dff_A_6XqmmfcU9_0),.din(w_dff_A_EKsT2u6v4_0),.clk(gclk));
	jdff dff_A_6XqmmfcU9_0(.dout(w_dff_A_8l1yDHw52_0),.din(w_dff_A_6XqmmfcU9_0),.clk(gclk));
	jdff dff_A_8l1yDHw52_0(.dout(w_dff_A_laH7v5ii6_0),.din(w_dff_A_8l1yDHw52_0),.clk(gclk));
	jdff dff_A_laH7v5ii6_0(.dout(w_dff_A_xgiFmAmt4_0),.din(w_dff_A_laH7v5ii6_0),.clk(gclk));
	jdff dff_A_xgiFmAmt4_0(.dout(w_dff_A_SFt0XsSv2_0),.din(w_dff_A_xgiFmAmt4_0),.clk(gclk));
	jdff dff_A_SFt0XsSv2_0(.dout(w_dff_A_pmSOYl6a7_0),.din(w_dff_A_SFt0XsSv2_0),.clk(gclk));
	jdff dff_A_pmSOYl6a7_0(.dout(w_dff_A_vTi1v3ik7_0),.din(w_dff_A_pmSOYl6a7_0),.clk(gclk));
	jdff dff_A_vTi1v3ik7_0(.dout(G923),.din(w_dff_A_vTi1v3ik7_0),.clk(gclk));
	jdff dff_A_7dsw62mq4_1(.dout(w_dff_A_MuunuXcW0_0),.din(w_dff_A_7dsw62mq4_1),.clk(gclk));
	jdff dff_A_MuunuXcW0_0(.dout(w_dff_A_5vCTJySf5_0),.din(w_dff_A_MuunuXcW0_0),.clk(gclk));
	jdff dff_A_5vCTJySf5_0(.dout(w_dff_A_RYOJbis28_0),.din(w_dff_A_5vCTJySf5_0),.clk(gclk));
	jdff dff_A_RYOJbis28_0(.dout(w_dff_A_MtY4ga2x0_0),.din(w_dff_A_RYOJbis28_0),.clk(gclk));
	jdff dff_A_MtY4ga2x0_0(.dout(w_dff_A_CJz1oVBS4_0),.din(w_dff_A_MtY4ga2x0_0),.clk(gclk));
	jdff dff_A_CJz1oVBS4_0(.dout(w_dff_A_bwPvtujk4_0),.din(w_dff_A_CJz1oVBS4_0),.clk(gclk));
	jdff dff_A_bwPvtujk4_0(.dout(w_dff_A_lpXRc5bz2_0),.din(w_dff_A_bwPvtujk4_0),.clk(gclk));
	jdff dff_A_lpXRc5bz2_0(.dout(w_dff_A_zfnB1HR61_0),.din(w_dff_A_lpXRc5bz2_0),.clk(gclk));
	jdff dff_A_zfnB1HR61_0(.dout(w_dff_A_y3R5ZmfI6_0),.din(w_dff_A_zfnB1HR61_0),.clk(gclk));
	jdff dff_A_y3R5ZmfI6_0(.dout(w_dff_A_7qg4YaXB4_0),.din(w_dff_A_y3R5ZmfI6_0),.clk(gclk));
	jdff dff_A_7qg4YaXB4_0(.dout(w_dff_A_HkNL83gj2_0),.din(w_dff_A_7qg4YaXB4_0),.clk(gclk));
	jdff dff_A_HkNL83gj2_0(.dout(w_dff_A_Pkhy5hB22_0),.din(w_dff_A_HkNL83gj2_0),.clk(gclk));
	jdff dff_A_Pkhy5hB22_0(.dout(w_dff_A_FC257lGZ0_0),.din(w_dff_A_Pkhy5hB22_0),.clk(gclk));
	jdff dff_A_FC257lGZ0_0(.dout(w_dff_A_lsJRvMu18_0),.din(w_dff_A_FC257lGZ0_0),.clk(gclk));
	jdff dff_A_lsJRvMu18_0(.dout(w_dff_A_QvDMxXil1_0),.din(w_dff_A_lsJRvMu18_0),.clk(gclk));
	jdff dff_A_QvDMxXil1_0(.dout(w_dff_A_HNrVC0ug4_0),.din(w_dff_A_QvDMxXil1_0),.clk(gclk));
	jdff dff_A_HNrVC0ug4_0(.dout(w_dff_A_gFdG6EaB9_0),.din(w_dff_A_HNrVC0ug4_0),.clk(gclk));
	jdff dff_A_gFdG6EaB9_0(.dout(w_dff_A_oKaXlgHz7_0),.din(w_dff_A_gFdG6EaB9_0),.clk(gclk));
	jdff dff_A_oKaXlgHz7_0(.dout(w_dff_A_NHR5rBU29_0),.din(w_dff_A_oKaXlgHz7_0),.clk(gclk));
	jdff dff_A_NHR5rBU29_0(.dout(w_dff_A_2Bodj7jw8_0),.din(w_dff_A_NHR5rBU29_0),.clk(gclk));
	jdff dff_A_2Bodj7jw8_0(.dout(w_dff_A_UW1p0P4r1_0),.din(w_dff_A_2Bodj7jw8_0),.clk(gclk));
	jdff dff_A_UW1p0P4r1_0(.dout(w_dff_A_8WY8intS6_0),.din(w_dff_A_UW1p0P4r1_0),.clk(gclk));
	jdff dff_A_8WY8intS6_0(.dout(w_dff_A_ZFGF9ZDk7_0),.din(w_dff_A_8WY8intS6_0),.clk(gclk));
	jdff dff_A_ZFGF9ZDk7_0(.dout(w_dff_A_3LOIkVtV0_0),.din(w_dff_A_ZFGF9ZDk7_0),.clk(gclk));
	jdff dff_A_3LOIkVtV0_0(.dout(w_dff_A_POEFWCQU0_0),.din(w_dff_A_3LOIkVtV0_0),.clk(gclk));
	jdff dff_A_POEFWCQU0_0(.dout(w_dff_A_4DCfUm7D8_0),.din(w_dff_A_POEFWCQU0_0),.clk(gclk));
	jdff dff_A_4DCfUm7D8_0(.dout(w_dff_A_8xI66C5M5_0),.din(w_dff_A_4DCfUm7D8_0),.clk(gclk));
	jdff dff_A_8xI66C5M5_0(.dout(G921),.din(w_dff_A_8xI66C5M5_0),.clk(gclk));
	jdff dff_A_c0W5v6CF5_1(.dout(w_dff_A_r5lRUBnq9_0),.din(w_dff_A_c0W5v6CF5_1),.clk(gclk));
	jdff dff_A_r5lRUBnq9_0(.dout(w_dff_A_kRSyerpV8_0),.din(w_dff_A_r5lRUBnq9_0),.clk(gclk));
	jdff dff_A_kRSyerpV8_0(.dout(w_dff_A_mX1pyvFx8_0),.din(w_dff_A_kRSyerpV8_0),.clk(gclk));
	jdff dff_A_mX1pyvFx8_0(.dout(w_dff_A_sTQLXnPG7_0),.din(w_dff_A_mX1pyvFx8_0),.clk(gclk));
	jdff dff_A_sTQLXnPG7_0(.dout(w_dff_A_RkEw0W1K6_0),.din(w_dff_A_sTQLXnPG7_0),.clk(gclk));
	jdff dff_A_RkEw0W1K6_0(.dout(w_dff_A_MD48YDDH5_0),.din(w_dff_A_RkEw0W1K6_0),.clk(gclk));
	jdff dff_A_MD48YDDH5_0(.dout(w_dff_A_YmgMDCs35_0),.din(w_dff_A_MD48YDDH5_0),.clk(gclk));
	jdff dff_A_YmgMDCs35_0(.dout(w_dff_A_xPJJ0fCl7_0),.din(w_dff_A_YmgMDCs35_0),.clk(gclk));
	jdff dff_A_xPJJ0fCl7_0(.dout(w_dff_A_sz8RdjQS9_0),.din(w_dff_A_xPJJ0fCl7_0),.clk(gclk));
	jdff dff_A_sz8RdjQS9_0(.dout(w_dff_A_qlyVixaW7_0),.din(w_dff_A_sz8RdjQS9_0),.clk(gclk));
	jdff dff_A_qlyVixaW7_0(.dout(w_dff_A_iuztysXN0_0),.din(w_dff_A_qlyVixaW7_0),.clk(gclk));
	jdff dff_A_iuztysXN0_0(.dout(w_dff_A_1ZpdAtcZ0_0),.din(w_dff_A_iuztysXN0_0),.clk(gclk));
	jdff dff_A_1ZpdAtcZ0_0(.dout(w_dff_A_cwRqYzhP6_0),.din(w_dff_A_1ZpdAtcZ0_0),.clk(gclk));
	jdff dff_A_cwRqYzhP6_0(.dout(w_dff_A_sEOzjlcf1_0),.din(w_dff_A_cwRqYzhP6_0),.clk(gclk));
	jdff dff_A_sEOzjlcf1_0(.dout(w_dff_A_mdxj7SA12_0),.din(w_dff_A_sEOzjlcf1_0),.clk(gclk));
	jdff dff_A_mdxj7SA12_0(.dout(w_dff_A_St3EwTge7_0),.din(w_dff_A_mdxj7SA12_0),.clk(gclk));
	jdff dff_A_St3EwTge7_0(.dout(w_dff_A_nox2nXZF0_0),.din(w_dff_A_St3EwTge7_0),.clk(gclk));
	jdff dff_A_nox2nXZF0_0(.dout(w_dff_A_rsseIDFd5_0),.din(w_dff_A_nox2nXZF0_0),.clk(gclk));
	jdff dff_A_rsseIDFd5_0(.dout(w_dff_A_1dzeVR4x5_0),.din(w_dff_A_rsseIDFd5_0),.clk(gclk));
	jdff dff_A_1dzeVR4x5_0(.dout(w_dff_A_4Rx18E6h1_0),.din(w_dff_A_1dzeVR4x5_0),.clk(gclk));
	jdff dff_A_4Rx18E6h1_0(.dout(w_dff_A_MYdC1wls7_0),.din(w_dff_A_4Rx18E6h1_0),.clk(gclk));
	jdff dff_A_MYdC1wls7_0(.dout(w_dff_A_ABVQdonB3_0),.din(w_dff_A_MYdC1wls7_0),.clk(gclk));
	jdff dff_A_ABVQdonB3_0(.dout(w_dff_A_vGTmAkVD5_0),.din(w_dff_A_ABVQdonB3_0),.clk(gclk));
	jdff dff_A_vGTmAkVD5_0(.dout(w_dff_A_P0VDaHoj4_0),.din(w_dff_A_vGTmAkVD5_0),.clk(gclk));
	jdff dff_A_P0VDaHoj4_0(.dout(w_dff_A_P1BRk2kJ4_0),.din(w_dff_A_P0VDaHoj4_0),.clk(gclk));
	jdff dff_A_P1BRk2kJ4_0(.dout(w_dff_A_IffsPDLL1_0),.din(w_dff_A_P1BRk2kJ4_0),.clk(gclk));
	jdff dff_A_IffsPDLL1_0(.dout(w_dff_A_RqoeCGpI4_0),.din(w_dff_A_IffsPDLL1_0),.clk(gclk));
	jdff dff_A_RqoeCGpI4_0(.dout(G892),.din(w_dff_A_RqoeCGpI4_0),.clk(gclk));
	jdff dff_A_acyZRsoC4_1(.dout(w_dff_A_HnbLRBsH4_0),.din(w_dff_A_acyZRsoC4_1),.clk(gclk));
	jdff dff_A_HnbLRBsH4_0(.dout(w_dff_A_fR0Abpyz4_0),.din(w_dff_A_HnbLRBsH4_0),.clk(gclk));
	jdff dff_A_fR0Abpyz4_0(.dout(w_dff_A_eZWlfAxR4_0),.din(w_dff_A_fR0Abpyz4_0),.clk(gclk));
	jdff dff_A_eZWlfAxR4_0(.dout(w_dff_A_xjFOEtOy0_0),.din(w_dff_A_eZWlfAxR4_0),.clk(gclk));
	jdff dff_A_xjFOEtOy0_0(.dout(w_dff_A_zcA8IKaL5_0),.din(w_dff_A_xjFOEtOy0_0),.clk(gclk));
	jdff dff_A_zcA8IKaL5_0(.dout(w_dff_A_guublbGq9_0),.din(w_dff_A_zcA8IKaL5_0),.clk(gclk));
	jdff dff_A_guublbGq9_0(.dout(w_dff_A_DHNFzFUI5_0),.din(w_dff_A_guublbGq9_0),.clk(gclk));
	jdff dff_A_DHNFzFUI5_0(.dout(w_dff_A_WeLGNQIq5_0),.din(w_dff_A_DHNFzFUI5_0),.clk(gclk));
	jdff dff_A_WeLGNQIq5_0(.dout(w_dff_A_9W0MtKpL7_0),.din(w_dff_A_WeLGNQIq5_0),.clk(gclk));
	jdff dff_A_9W0MtKpL7_0(.dout(w_dff_A_jdrfZO7y6_0),.din(w_dff_A_9W0MtKpL7_0),.clk(gclk));
	jdff dff_A_jdrfZO7y6_0(.dout(w_dff_A_VRDWPNtr4_0),.din(w_dff_A_jdrfZO7y6_0),.clk(gclk));
	jdff dff_A_VRDWPNtr4_0(.dout(w_dff_A_LINeIFbt8_0),.din(w_dff_A_VRDWPNtr4_0),.clk(gclk));
	jdff dff_A_LINeIFbt8_0(.dout(w_dff_A_AU7ahig87_0),.din(w_dff_A_LINeIFbt8_0),.clk(gclk));
	jdff dff_A_AU7ahig87_0(.dout(w_dff_A_dJl9E4s11_0),.din(w_dff_A_AU7ahig87_0),.clk(gclk));
	jdff dff_A_dJl9E4s11_0(.dout(w_dff_A_HBuQM9BI7_0),.din(w_dff_A_dJl9E4s11_0),.clk(gclk));
	jdff dff_A_HBuQM9BI7_0(.dout(w_dff_A_C7tQtGoP0_0),.din(w_dff_A_HBuQM9BI7_0),.clk(gclk));
	jdff dff_A_C7tQtGoP0_0(.dout(w_dff_A_3PSg393z5_0),.din(w_dff_A_C7tQtGoP0_0),.clk(gclk));
	jdff dff_A_3PSg393z5_0(.dout(w_dff_A_QdgffaEX3_0),.din(w_dff_A_3PSg393z5_0),.clk(gclk));
	jdff dff_A_QdgffaEX3_0(.dout(w_dff_A_CK0mp0d94_0),.din(w_dff_A_QdgffaEX3_0),.clk(gclk));
	jdff dff_A_CK0mp0d94_0(.dout(w_dff_A_Qw0w5TUn9_0),.din(w_dff_A_CK0mp0d94_0),.clk(gclk));
	jdff dff_A_Qw0w5TUn9_0(.dout(w_dff_A_4K2NvvMu6_0),.din(w_dff_A_Qw0w5TUn9_0),.clk(gclk));
	jdff dff_A_4K2NvvMu6_0(.dout(w_dff_A_iomx5FVG3_0),.din(w_dff_A_4K2NvvMu6_0),.clk(gclk));
	jdff dff_A_iomx5FVG3_0(.dout(w_dff_A_BYYqPllx1_0),.din(w_dff_A_iomx5FVG3_0),.clk(gclk));
	jdff dff_A_BYYqPllx1_0(.dout(w_dff_A_jO9zTWys7_0),.din(w_dff_A_BYYqPllx1_0),.clk(gclk));
	jdff dff_A_jO9zTWys7_0(.dout(w_dff_A_8sxygSq53_0),.din(w_dff_A_jO9zTWys7_0),.clk(gclk));
	jdff dff_A_8sxygSq53_0(.dout(w_dff_A_BekpnsSZ5_0),.din(w_dff_A_8sxygSq53_0),.clk(gclk));
	jdff dff_A_BekpnsSZ5_0(.dout(w_dff_A_yTo56sWa6_0),.din(w_dff_A_BekpnsSZ5_0),.clk(gclk));
	jdff dff_A_yTo56sWa6_0(.dout(G887),.din(w_dff_A_yTo56sWa6_0),.clk(gclk));
	jdff dff_A_b5bppP9C3_1(.dout(w_dff_A_hnE3BRfa8_0),.din(w_dff_A_b5bppP9C3_1),.clk(gclk));
	jdff dff_A_hnE3BRfa8_0(.dout(w_dff_A_czA4SQ235_0),.din(w_dff_A_hnE3BRfa8_0),.clk(gclk));
	jdff dff_A_czA4SQ235_0(.dout(w_dff_A_r37FywQz6_0),.din(w_dff_A_czA4SQ235_0),.clk(gclk));
	jdff dff_A_r37FywQz6_0(.dout(w_dff_A_ZyjzyN5B5_0),.din(w_dff_A_r37FywQz6_0),.clk(gclk));
	jdff dff_A_ZyjzyN5B5_0(.dout(w_dff_A_DK3WwJLG1_0),.din(w_dff_A_ZyjzyN5B5_0),.clk(gclk));
	jdff dff_A_DK3WwJLG1_0(.dout(w_dff_A_mg0rV9i28_0),.din(w_dff_A_DK3WwJLG1_0),.clk(gclk));
	jdff dff_A_mg0rV9i28_0(.dout(w_dff_A_H1y6fXa81_0),.din(w_dff_A_mg0rV9i28_0),.clk(gclk));
	jdff dff_A_H1y6fXa81_0(.dout(w_dff_A_baiwRXhO1_0),.din(w_dff_A_H1y6fXa81_0),.clk(gclk));
	jdff dff_A_baiwRXhO1_0(.dout(w_dff_A_v9BqxDiH3_0),.din(w_dff_A_baiwRXhO1_0),.clk(gclk));
	jdff dff_A_v9BqxDiH3_0(.dout(w_dff_A_JkIV7ZTq8_0),.din(w_dff_A_v9BqxDiH3_0),.clk(gclk));
	jdff dff_A_JkIV7ZTq8_0(.dout(w_dff_A_zqlpA7yf2_0),.din(w_dff_A_JkIV7ZTq8_0),.clk(gclk));
	jdff dff_A_zqlpA7yf2_0(.dout(w_dff_A_q2lKCze97_0),.din(w_dff_A_zqlpA7yf2_0),.clk(gclk));
	jdff dff_A_q2lKCze97_0(.dout(w_dff_A_MsLvlfxG9_0),.din(w_dff_A_q2lKCze97_0),.clk(gclk));
	jdff dff_A_MsLvlfxG9_0(.dout(w_dff_A_XmmkHZng5_0),.din(w_dff_A_MsLvlfxG9_0),.clk(gclk));
	jdff dff_A_XmmkHZng5_0(.dout(w_dff_A_TFyeyPa05_0),.din(w_dff_A_XmmkHZng5_0),.clk(gclk));
	jdff dff_A_TFyeyPa05_0(.dout(w_dff_A_AcrGSD6c7_0),.din(w_dff_A_TFyeyPa05_0),.clk(gclk));
	jdff dff_A_AcrGSD6c7_0(.dout(w_dff_A_Io1XcflI7_0),.din(w_dff_A_AcrGSD6c7_0),.clk(gclk));
	jdff dff_A_Io1XcflI7_0(.dout(w_dff_A_2rpTxKuA7_0),.din(w_dff_A_Io1XcflI7_0),.clk(gclk));
	jdff dff_A_2rpTxKuA7_0(.dout(w_dff_A_ZU6jxPRt4_0),.din(w_dff_A_2rpTxKuA7_0),.clk(gclk));
	jdff dff_A_ZU6jxPRt4_0(.dout(w_dff_A_C80ll9O55_0),.din(w_dff_A_ZU6jxPRt4_0),.clk(gclk));
	jdff dff_A_C80ll9O55_0(.dout(w_dff_A_WtOeLjFY5_0),.din(w_dff_A_C80ll9O55_0),.clk(gclk));
	jdff dff_A_WtOeLjFY5_0(.dout(w_dff_A_EBSmERs53_0),.din(w_dff_A_WtOeLjFY5_0),.clk(gclk));
	jdff dff_A_EBSmERs53_0(.dout(w_dff_A_R89C3gym6_0),.din(w_dff_A_EBSmERs53_0),.clk(gclk));
	jdff dff_A_R89C3gym6_0(.dout(w_dff_A_Up7ZdmrK2_0),.din(w_dff_A_R89C3gym6_0),.clk(gclk));
	jdff dff_A_Up7ZdmrK2_0(.dout(w_dff_A_DWSKUaut1_0),.din(w_dff_A_Up7ZdmrK2_0),.clk(gclk));
	jdff dff_A_DWSKUaut1_0(.dout(w_dff_A_bClPVLyy4_0),.din(w_dff_A_DWSKUaut1_0),.clk(gclk));
	jdff dff_A_bClPVLyy4_0(.dout(G606),.din(w_dff_A_bClPVLyy4_0),.clk(gclk));
	jdff dff_A_Cg0ajXrl8_2(.dout(w_dff_A_geKvccbu1_0),.din(w_dff_A_Cg0ajXrl8_2),.clk(gclk));
	jdff dff_A_geKvccbu1_0(.dout(w_dff_A_N6XWPsdF4_0),.din(w_dff_A_geKvccbu1_0),.clk(gclk));
	jdff dff_A_N6XWPsdF4_0(.dout(w_dff_A_0rwvwVbQ9_0),.din(w_dff_A_N6XWPsdF4_0),.clk(gclk));
	jdff dff_A_0rwvwVbQ9_0(.dout(w_dff_A_beL712qd1_0),.din(w_dff_A_0rwvwVbQ9_0),.clk(gclk));
	jdff dff_A_beL712qd1_0(.dout(w_dff_A_i8O7E6XR2_0),.din(w_dff_A_beL712qd1_0),.clk(gclk));
	jdff dff_A_i8O7E6XR2_0(.dout(w_dff_A_JqarZ9RO6_0),.din(w_dff_A_i8O7E6XR2_0),.clk(gclk));
	jdff dff_A_JqarZ9RO6_0(.dout(w_dff_A_NOqzOnpU8_0),.din(w_dff_A_JqarZ9RO6_0),.clk(gclk));
	jdff dff_A_NOqzOnpU8_0(.dout(w_dff_A_KSvOr7C56_0),.din(w_dff_A_NOqzOnpU8_0),.clk(gclk));
	jdff dff_A_KSvOr7C56_0(.dout(w_dff_A_HB9qGMTO4_0),.din(w_dff_A_KSvOr7C56_0),.clk(gclk));
	jdff dff_A_HB9qGMTO4_0(.dout(w_dff_A_Nwewo1uX4_0),.din(w_dff_A_HB9qGMTO4_0),.clk(gclk));
	jdff dff_A_Nwewo1uX4_0(.dout(w_dff_A_epYu035e1_0),.din(w_dff_A_Nwewo1uX4_0),.clk(gclk));
	jdff dff_A_epYu035e1_0(.dout(w_dff_A_0MoJMuhU0_0),.din(w_dff_A_epYu035e1_0),.clk(gclk));
	jdff dff_A_0MoJMuhU0_0(.dout(w_dff_A_FUjHRh7t6_0),.din(w_dff_A_0MoJMuhU0_0),.clk(gclk));
	jdff dff_A_FUjHRh7t6_0(.dout(w_dff_A_6tA5NXI79_0),.din(w_dff_A_FUjHRh7t6_0),.clk(gclk));
	jdff dff_A_6tA5NXI79_0(.dout(w_dff_A_j8AT1bTg5_0),.din(w_dff_A_6tA5NXI79_0),.clk(gclk));
	jdff dff_A_j8AT1bTg5_0(.dout(w_dff_A_JUN2CzMo0_0),.din(w_dff_A_j8AT1bTg5_0),.clk(gclk));
	jdff dff_A_JUN2CzMo0_0(.dout(w_dff_A_KyawlIOu0_0),.din(w_dff_A_JUN2CzMo0_0),.clk(gclk));
	jdff dff_A_KyawlIOu0_0(.dout(w_dff_A_zTdIvZ7q8_0),.din(w_dff_A_KyawlIOu0_0),.clk(gclk));
	jdff dff_A_zTdIvZ7q8_0(.dout(w_dff_A_vYhjTbvR1_0),.din(w_dff_A_zTdIvZ7q8_0),.clk(gclk));
	jdff dff_A_vYhjTbvR1_0(.dout(w_dff_A_522ZjSav3_0),.din(w_dff_A_vYhjTbvR1_0),.clk(gclk));
	jdff dff_A_522ZjSav3_0(.dout(w_dff_A_yvvkBSnw3_0),.din(w_dff_A_522ZjSav3_0),.clk(gclk));
	jdff dff_A_yvvkBSnw3_0(.dout(w_dff_A_App9HfCg7_0),.din(w_dff_A_yvvkBSnw3_0),.clk(gclk));
	jdff dff_A_App9HfCg7_0(.dout(w_dff_A_5cR1rmsk3_0),.din(w_dff_A_App9HfCg7_0),.clk(gclk));
	jdff dff_A_5cR1rmsk3_0(.dout(w_dff_A_UkXn478t6_0),.din(w_dff_A_5cR1rmsk3_0),.clk(gclk));
	jdff dff_A_UkXn478t6_0(.dout(G656),.din(w_dff_A_UkXn478t6_0),.clk(gclk));
	jdff dff_A_a0LYu7n60_2(.dout(w_dff_A_ZeXevlTk5_0),.din(w_dff_A_a0LYu7n60_2),.clk(gclk));
	jdff dff_A_ZeXevlTk5_0(.dout(w_dff_A_WDmciOda7_0),.din(w_dff_A_ZeXevlTk5_0),.clk(gclk));
	jdff dff_A_WDmciOda7_0(.dout(w_dff_A_WrQ06h0i6_0),.din(w_dff_A_WDmciOda7_0),.clk(gclk));
	jdff dff_A_WrQ06h0i6_0(.dout(w_dff_A_zsZpcWy06_0),.din(w_dff_A_WrQ06h0i6_0),.clk(gclk));
	jdff dff_A_zsZpcWy06_0(.dout(w_dff_A_JXiXryOx2_0),.din(w_dff_A_zsZpcWy06_0),.clk(gclk));
	jdff dff_A_JXiXryOx2_0(.dout(w_dff_A_e3mYZuAI1_0),.din(w_dff_A_JXiXryOx2_0),.clk(gclk));
	jdff dff_A_e3mYZuAI1_0(.dout(w_dff_A_MPf1c4C05_0),.din(w_dff_A_e3mYZuAI1_0),.clk(gclk));
	jdff dff_A_MPf1c4C05_0(.dout(w_dff_A_XhAf601Y5_0),.din(w_dff_A_MPf1c4C05_0),.clk(gclk));
	jdff dff_A_XhAf601Y5_0(.dout(w_dff_A_3qWMNiSy2_0),.din(w_dff_A_XhAf601Y5_0),.clk(gclk));
	jdff dff_A_3qWMNiSy2_0(.dout(w_dff_A_cczxyAGQ8_0),.din(w_dff_A_3qWMNiSy2_0),.clk(gclk));
	jdff dff_A_cczxyAGQ8_0(.dout(w_dff_A_cxV0sJJm4_0),.din(w_dff_A_cczxyAGQ8_0),.clk(gclk));
	jdff dff_A_cxV0sJJm4_0(.dout(w_dff_A_svYmSWiN7_0),.din(w_dff_A_cxV0sJJm4_0),.clk(gclk));
	jdff dff_A_svYmSWiN7_0(.dout(w_dff_A_WbyHGIz05_0),.din(w_dff_A_svYmSWiN7_0),.clk(gclk));
	jdff dff_A_WbyHGIz05_0(.dout(w_dff_A_SIkVC4Oc5_0),.din(w_dff_A_WbyHGIz05_0),.clk(gclk));
	jdff dff_A_SIkVC4Oc5_0(.dout(w_dff_A_HiKZrVz16_0),.din(w_dff_A_SIkVC4Oc5_0),.clk(gclk));
	jdff dff_A_HiKZrVz16_0(.dout(w_dff_A_ZtkjIz6t9_0),.din(w_dff_A_HiKZrVz16_0),.clk(gclk));
	jdff dff_A_ZtkjIz6t9_0(.dout(w_dff_A_D1ehCP2g4_0),.din(w_dff_A_ZtkjIz6t9_0),.clk(gclk));
	jdff dff_A_D1ehCP2g4_0(.dout(w_dff_A_19mRsXm90_0),.din(w_dff_A_D1ehCP2g4_0),.clk(gclk));
	jdff dff_A_19mRsXm90_0(.dout(w_dff_A_zcgssLyH6_0),.din(w_dff_A_19mRsXm90_0),.clk(gclk));
	jdff dff_A_zcgssLyH6_0(.dout(w_dff_A_Y6WorKqY9_0),.din(w_dff_A_zcgssLyH6_0),.clk(gclk));
	jdff dff_A_Y6WorKqY9_0(.dout(w_dff_A_WZUdXUac6_0),.din(w_dff_A_Y6WorKqY9_0),.clk(gclk));
	jdff dff_A_WZUdXUac6_0(.dout(w_dff_A_BVHaAflh5_0),.din(w_dff_A_WZUdXUac6_0),.clk(gclk));
	jdff dff_A_BVHaAflh5_0(.dout(w_dff_A_9OeQf4eb6_0),.din(w_dff_A_BVHaAflh5_0),.clk(gclk));
	jdff dff_A_9OeQf4eb6_0(.dout(w_dff_A_8tyub3pi3_0),.din(w_dff_A_9OeQf4eb6_0),.clk(gclk));
	jdff dff_A_8tyub3pi3_0(.dout(w_dff_A_LqIS8KAc4_0),.din(w_dff_A_8tyub3pi3_0),.clk(gclk));
	jdff dff_A_LqIS8KAc4_0(.dout(G809),.din(w_dff_A_LqIS8KAc4_0),.clk(gclk));
	jdff dff_A_4QLAB4kJ6_1(.dout(w_dff_A_CZMGzdzz1_0),.din(w_dff_A_4QLAB4kJ6_1),.clk(gclk));
	jdff dff_A_CZMGzdzz1_0(.dout(w_dff_A_Ygeuxq6F1_0),.din(w_dff_A_CZMGzdzz1_0),.clk(gclk));
	jdff dff_A_Ygeuxq6F1_0(.dout(w_dff_A_z1ji51ux9_0),.din(w_dff_A_Ygeuxq6F1_0),.clk(gclk));
	jdff dff_A_z1ji51ux9_0(.dout(w_dff_A_PyjhS6S69_0),.din(w_dff_A_z1ji51ux9_0),.clk(gclk));
	jdff dff_A_PyjhS6S69_0(.dout(w_dff_A_teiiGtEp3_0),.din(w_dff_A_PyjhS6S69_0),.clk(gclk));
	jdff dff_A_teiiGtEp3_0(.dout(w_dff_A_HYOg3Bkv0_0),.din(w_dff_A_teiiGtEp3_0),.clk(gclk));
	jdff dff_A_HYOg3Bkv0_0(.dout(w_dff_A_bSe9Pnpw0_0),.din(w_dff_A_HYOg3Bkv0_0),.clk(gclk));
	jdff dff_A_bSe9Pnpw0_0(.dout(w_dff_A_uVOTm3Ko8_0),.din(w_dff_A_bSe9Pnpw0_0),.clk(gclk));
	jdff dff_A_uVOTm3Ko8_0(.dout(w_dff_A_qFqMhNkT7_0),.din(w_dff_A_uVOTm3Ko8_0),.clk(gclk));
	jdff dff_A_qFqMhNkT7_0(.dout(w_dff_A_IBqmQwFT7_0),.din(w_dff_A_qFqMhNkT7_0),.clk(gclk));
	jdff dff_A_IBqmQwFT7_0(.dout(w_dff_A_0TW2eqjN3_0),.din(w_dff_A_IBqmQwFT7_0),.clk(gclk));
	jdff dff_A_0TW2eqjN3_0(.dout(w_dff_A_JyQeqs1D0_0),.din(w_dff_A_0TW2eqjN3_0),.clk(gclk));
	jdff dff_A_JyQeqs1D0_0(.dout(w_dff_A_sZKe8kQL4_0),.din(w_dff_A_JyQeqs1D0_0),.clk(gclk));
	jdff dff_A_sZKe8kQL4_0(.dout(w_dff_A_ODDK0O692_0),.din(w_dff_A_sZKe8kQL4_0),.clk(gclk));
	jdff dff_A_ODDK0O692_0(.dout(w_dff_A_GD1Y1epJ9_0),.din(w_dff_A_ODDK0O692_0),.clk(gclk));
	jdff dff_A_GD1Y1epJ9_0(.dout(w_dff_A_3d8b4sE41_0),.din(w_dff_A_GD1Y1epJ9_0),.clk(gclk));
	jdff dff_A_3d8b4sE41_0(.dout(w_dff_A_ul2CZcZb9_0),.din(w_dff_A_3d8b4sE41_0),.clk(gclk));
	jdff dff_A_ul2CZcZb9_0(.dout(w_dff_A_Z6eb98ke2_0),.din(w_dff_A_ul2CZcZb9_0),.clk(gclk));
	jdff dff_A_Z6eb98ke2_0(.dout(w_dff_A_sxTzbnvi1_0),.din(w_dff_A_Z6eb98ke2_0),.clk(gclk));
	jdff dff_A_sxTzbnvi1_0(.dout(w_dff_A_ldl9McF27_0),.din(w_dff_A_sxTzbnvi1_0),.clk(gclk));
	jdff dff_A_ldl9McF27_0(.dout(w_dff_A_OmZtZWER0_0),.din(w_dff_A_ldl9McF27_0),.clk(gclk));
	jdff dff_A_OmZtZWER0_0(.dout(w_dff_A_xunTitrv4_0),.din(w_dff_A_OmZtZWER0_0),.clk(gclk));
	jdff dff_A_xunTitrv4_0(.dout(w_dff_A_qnVCCIDy9_0),.din(w_dff_A_xunTitrv4_0),.clk(gclk));
	jdff dff_A_qnVCCIDy9_0(.dout(w_dff_A_wsa53kUS7_0),.din(w_dff_A_qnVCCIDy9_0),.clk(gclk));
	jdff dff_A_wsa53kUS7_0(.dout(w_dff_A_t9wlPRPO2_0),.din(w_dff_A_wsa53kUS7_0),.clk(gclk));
	jdff dff_A_t9wlPRPO2_0(.dout(w_dff_A_77SON5gz3_0),.din(w_dff_A_t9wlPRPO2_0),.clk(gclk));
	jdff dff_A_77SON5gz3_0(.dout(w_dff_A_bPKViaZU8_0),.din(w_dff_A_77SON5gz3_0),.clk(gclk));
	jdff dff_A_bPKViaZU8_0(.dout(G993),.din(w_dff_A_bPKViaZU8_0),.clk(gclk));
	jdff dff_A_5y0biOwJ6_1(.dout(w_dff_A_CuP3HU3H8_0),.din(w_dff_A_5y0biOwJ6_1),.clk(gclk));
	jdff dff_A_CuP3HU3H8_0(.dout(w_dff_A_6wgO6idh6_0),.din(w_dff_A_CuP3HU3H8_0),.clk(gclk));
	jdff dff_A_6wgO6idh6_0(.dout(w_dff_A_77yPZ8fE1_0),.din(w_dff_A_6wgO6idh6_0),.clk(gclk));
	jdff dff_A_77yPZ8fE1_0(.dout(w_dff_A_33yENelA7_0),.din(w_dff_A_77yPZ8fE1_0),.clk(gclk));
	jdff dff_A_33yENelA7_0(.dout(w_dff_A_8hleZckD4_0),.din(w_dff_A_33yENelA7_0),.clk(gclk));
	jdff dff_A_8hleZckD4_0(.dout(w_dff_A_f6suGJYz6_0),.din(w_dff_A_8hleZckD4_0),.clk(gclk));
	jdff dff_A_f6suGJYz6_0(.dout(w_dff_A_kY1TDHTo0_0),.din(w_dff_A_f6suGJYz6_0),.clk(gclk));
	jdff dff_A_kY1TDHTo0_0(.dout(w_dff_A_Wja7P7eQ7_0),.din(w_dff_A_kY1TDHTo0_0),.clk(gclk));
	jdff dff_A_Wja7P7eQ7_0(.dout(w_dff_A_p9zFzQ8H6_0),.din(w_dff_A_Wja7P7eQ7_0),.clk(gclk));
	jdff dff_A_p9zFzQ8H6_0(.dout(w_dff_A_YoR81gSB6_0),.din(w_dff_A_p9zFzQ8H6_0),.clk(gclk));
	jdff dff_A_YoR81gSB6_0(.dout(w_dff_A_wp3MD9zv8_0),.din(w_dff_A_YoR81gSB6_0),.clk(gclk));
	jdff dff_A_wp3MD9zv8_0(.dout(w_dff_A_udm87nCJ5_0),.din(w_dff_A_wp3MD9zv8_0),.clk(gclk));
	jdff dff_A_udm87nCJ5_0(.dout(w_dff_A_2c66gJNO3_0),.din(w_dff_A_udm87nCJ5_0),.clk(gclk));
	jdff dff_A_2c66gJNO3_0(.dout(w_dff_A_0pbHLEuH4_0),.din(w_dff_A_2c66gJNO3_0),.clk(gclk));
	jdff dff_A_0pbHLEuH4_0(.dout(w_dff_A_u9PwAwCX0_0),.din(w_dff_A_0pbHLEuH4_0),.clk(gclk));
	jdff dff_A_u9PwAwCX0_0(.dout(w_dff_A_5syXSLwY7_0),.din(w_dff_A_u9PwAwCX0_0),.clk(gclk));
	jdff dff_A_5syXSLwY7_0(.dout(w_dff_A_Tx9q6x1D7_0),.din(w_dff_A_5syXSLwY7_0),.clk(gclk));
	jdff dff_A_Tx9q6x1D7_0(.dout(w_dff_A_orBuZSoy1_0),.din(w_dff_A_Tx9q6x1D7_0),.clk(gclk));
	jdff dff_A_orBuZSoy1_0(.dout(w_dff_A_NvLUnGYQ0_0),.din(w_dff_A_orBuZSoy1_0),.clk(gclk));
	jdff dff_A_NvLUnGYQ0_0(.dout(w_dff_A_N7DRbtX59_0),.din(w_dff_A_NvLUnGYQ0_0),.clk(gclk));
	jdff dff_A_N7DRbtX59_0(.dout(w_dff_A_qc7W0tKd1_0),.din(w_dff_A_N7DRbtX59_0),.clk(gclk));
	jdff dff_A_qc7W0tKd1_0(.dout(w_dff_A_dXj9QJZS2_0),.din(w_dff_A_qc7W0tKd1_0),.clk(gclk));
	jdff dff_A_dXj9QJZS2_0(.dout(w_dff_A_1MMrnxhe8_0),.din(w_dff_A_dXj9QJZS2_0),.clk(gclk));
	jdff dff_A_1MMrnxhe8_0(.dout(w_dff_A_30e7C8yc1_0),.din(w_dff_A_1MMrnxhe8_0),.clk(gclk));
	jdff dff_A_30e7C8yc1_0(.dout(w_dff_A_BdDXYNqW2_0),.din(w_dff_A_30e7C8yc1_0),.clk(gclk));
	jdff dff_A_BdDXYNqW2_0(.dout(w_dff_A_JCS8MAGB3_0),.din(w_dff_A_BdDXYNqW2_0),.clk(gclk));
	jdff dff_A_JCS8MAGB3_0(.dout(w_dff_A_8dGDKZ2C3_0),.din(w_dff_A_JCS8MAGB3_0),.clk(gclk));
	jdff dff_A_8dGDKZ2C3_0(.dout(G978),.din(w_dff_A_8dGDKZ2C3_0),.clk(gclk));
	jdff dff_A_S9WcFqMu6_1(.dout(w_dff_A_9C07X2mv9_0),.din(w_dff_A_S9WcFqMu6_1),.clk(gclk));
	jdff dff_A_9C07X2mv9_0(.dout(w_dff_A_Wu1mNrHt8_0),.din(w_dff_A_9C07X2mv9_0),.clk(gclk));
	jdff dff_A_Wu1mNrHt8_0(.dout(w_dff_A_qdln7FBI9_0),.din(w_dff_A_Wu1mNrHt8_0),.clk(gclk));
	jdff dff_A_qdln7FBI9_0(.dout(w_dff_A_Hr9sj9h72_0),.din(w_dff_A_qdln7FBI9_0),.clk(gclk));
	jdff dff_A_Hr9sj9h72_0(.dout(w_dff_A_FScjYHSM4_0),.din(w_dff_A_Hr9sj9h72_0),.clk(gclk));
	jdff dff_A_FScjYHSM4_0(.dout(w_dff_A_TIFR0Jk78_0),.din(w_dff_A_FScjYHSM4_0),.clk(gclk));
	jdff dff_A_TIFR0Jk78_0(.dout(w_dff_A_LCTuYaip1_0),.din(w_dff_A_TIFR0Jk78_0),.clk(gclk));
	jdff dff_A_LCTuYaip1_0(.dout(w_dff_A_ZlS9lcro7_0),.din(w_dff_A_LCTuYaip1_0),.clk(gclk));
	jdff dff_A_ZlS9lcro7_0(.dout(w_dff_A_6kbjqBFj3_0),.din(w_dff_A_ZlS9lcro7_0),.clk(gclk));
	jdff dff_A_6kbjqBFj3_0(.dout(w_dff_A_rPwsrr137_0),.din(w_dff_A_6kbjqBFj3_0),.clk(gclk));
	jdff dff_A_rPwsrr137_0(.dout(w_dff_A_qft6sav31_0),.din(w_dff_A_rPwsrr137_0),.clk(gclk));
	jdff dff_A_qft6sav31_0(.dout(w_dff_A_izZgnMVf1_0),.din(w_dff_A_qft6sav31_0),.clk(gclk));
	jdff dff_A_izZgnMVf1_0(.dout(w_dff_A_OIyUcUvC0_0),.din(w_dff_A_izZgnMVf1_0),.clk(gclk));
	jdff dff_A_OIyUcUvC0_0(.dout(w_dff_A_KIQgKCiW7_0),.din(w_dff_A_OIyUcUvC0_0),.clk(gclk));
	jdff dff_A_KIQgKCiW7_0(.dout(w_dff_A_vSzyXNyz4_0),.din(w_dff_A_KIQgKCiW7_0),.clk(gclk));
	jdff dff_A_vSzyXNyz4_0(.dout(w_dff_A_6idpLyrK4_0),.din(w_dff_A_vSzyXNyz4_0),.clk(gclk));
	jdff dff_A_6idpLyrK4_0(.dout(w_dff_A_aQbxkq9u8_0),.din(w_dff_A_6idpLyrK4_0),.clk(gclk));
	jdff dff_A_aQbxkq9u8_0(.dout(w_dff_A_FMX48Gvb7_0),.din(w_dff_A_aQbxkq9u8_0),.clk(gclk));
	jdff dff_A_FMX48Gvb7_0(.dout(w_dff_A_fAaUdg9x1_0),.din(w_dff_A_FMX48Gvb7_0),.clk(gclk));
	jdff dff_A_fAaUdg9x1_0(.dout(w_dff_A_hN3egfdk4_0),.din(w_dff_A_fAaUdg9x1_0),.clk(gclk));
	jdff dff_A_hN3egfdk4_0(.dout(w_dff_A_5Elq8oQI6_0),.din(w_dff_A_hN3egfdk4_0),.clk(gclk));
	jdff dff_A_5Elq8oQI6_0(.dout(w_dff_A_HKzzsOWF6_0),.din(w_dff_A_5Elq8oQI6_0),.clk(gclk));
	jdff dff_A_HKzzsOWF6_0(.dout(w_dff_A_dKdYD9LK0_0),.din(w_dff_A_HKzzsOWF6_0),.clk(gclk));
	jdff dff_A_dKdYD9LK0_0(.dout(w_dff_A_dQHTlihh4_0),.din(w_dff_A_dKdYD9LK0_0),.clk(gclk));
	jdff dff_A_dQHTlihh4_0(.dout(w_dff_A_fiWm97NV6_0),.din(w_dff_A_dQHTlihh4_0),.clk(gclk));
	jdff dff_A_fiWm97NV6_0(.dout(w_dff_A_SAlkhw2R0_0),.din(w_dff_A_fiWm97NV6_0),.clk(gclk));
	jdff dff_A_SAlkhw2R0_0(.dout(w_dff_A_S1wMbJWo4_0),.din(w_dff_A_SAlkhw2R0_0),.clk(gclk));
	jdff dff_A_S1wMbJWo4_0(.dout(G949),.din(w_dff_A_S1wMbJWo4_0),.clk(gclk));
	jdff dff_A_HDNNfVWU5_1(.dout(w_dff_A_6sfFDXGC5_0),.din(w_dff_A_HDNNfVWU5_1),.clk(gclk));
	jdff dff_A_6sfFDXGC5_0(.dout(w_dff_A_DJP4JRbb1_0),.din(w_dff_A_6sfFDXGC5_0),.clk(gclk));
	jdff dff_A_DJP4JRbb1_0(.dout(w_dff_A_LzIu2Qtx1_0),.din(w_dff_A_DJP4JRbb1_0),.clk(gclk));
	jdff dff_A_LzIu2Qtx1_0(.dout(w_dff_A_nFTDqOIK6_0),.din(w_dff_A_LzIu2Qtx1_0),.clk(gclk));
	jdff dff_A_nFTDqOIK6_0(.dout(w_dff_A_B4I7hajb7_0),.din(w_dff_A_nFTDqOIK6_0),.clk(gclk));
	jdff dff_A_B4I7hajb7_0(.dout(w_dff_A_byCKrMao9_0),.din(w_dff_A_B4I7hajb7_0),.clk(gclk));
	jdff dff_A_byCKrMao9_0(.dout(w_dff_A_vlrU0L6F8_0),.din(w_dff_A_byCKrMao9_0),.clk(gclk));
	jdff dff_A_vlrU0L6F8_0(.dout(w_dff_A_JaNHCmAC6_0),.din(w_dff_A_vlrU0L6F8_0),.clk(gclk));
	jdff dff_A_JaNHCmAC6_0(.dout(w_dff_A_qAoeGtu41_0),.din(w_dff_A_JaNHCmAC6_0),.clk(gclk));
	jdff dff_A_qAoeGtu41_0(.dout(w_dff_A_KEXImDku0_0),.din(w_dff_A_qAoeGtu41_0),.clk(gclk));
	jdff dff_A_KEXImDku0_0(.dout(w_dff_A_lYSxZKYt3_0),.din(w_dff_A_KEXImDku0_0),.clk(gclk));
	jdff dff_A_lYSxZKYt3_0(.dout(w_dff_A_xa7DKjyO9_0),.din(w_dff_A_lYSxZKYt3_0),.clk(gclk));
	jdff dff_A_xa7DKjyO9_0(.dout(w_dff_A_SJKwhtJY1_0),.din(w_dff_A_xa7DKjyO9_0),.clk(gclk));
	jdff dff_A_SJKwhtJY1_0(.dout(w_dff_A_rK2EIooO4_0),.din(w_dff_A_SJKwhtJY1_0),.clk(gclk));
	jdff dff_A_rK2EIooO4_0(.dout(w_dff_A_zOOgChGn2_0),.din(w_dff_A_rK2EIooO4_0),.clk(gclk));
	jdff dff_A_zOOgChGn2_0(.dout(w_dff_A_XMT8fIlf2_0),.din(w_dff_A_zOOgChGn2_0),.clk(gclk));
	jdff dff_A_XMT8fIlf2_0(.dout(w_dff_A_MiGnPugq5_0),.din(w_dff_A_XMT8fIlf2_0),.clk(gclk));
	jdff dff_A_MiGnPugq5_0(.dout(w_dff_A_ih7JIhlA5_0),.din(w_dff_A_MiGnPugq5_0),.clk(gclk));
	jdff dff_A_ih7JIhlA5_0(.dout(w_dff_A_aTYq7vq69_0),.din(w_dff_A_ih7JIhlA5_0),.clk(gclk));
	jdff dff_A_aTYq7vq69_0(.dout(w_dff_A_mrxKdql00_0),.din(w_dff_A_aTYq7vq69_0),.clk(gclk));
	jdff dff_A_mrxKdql00_0(.dout(w_dff_A_JbZu5Vcb3_0),.din(w_dff_A_mrxKdql00_0),.clk(gclk));
	jdff dff_A_JbZu5Vcb3_0(.dout(w_dff_A_etlZr0Fc4_0),.din(w_dff_A_JbZu5Vcb3_0),.clk(gclk));
	jdff dff_A_etlZr0Fc4_0(.dout(w_dff_A_y9Fhn2iO1_0),.din(w_dff_A_etlZr0Fc4_0),.clk(gclk));
	jdff dff_A_y9Fhn2iO1_0(.dout(w_dff_A_aV9d9Ahv4_0),.din(w_dff_A_y9Fhn2iO1_0),.clk(gclk));
	jdff dff_A_aV9d9Ahv4_0(.dout(w_dff_A_HYY14ous9_0),.din(w_dff_A_aV9d9Ahv4_0),.clk(gclk));
	jdff dff_A_HYY14ous9_0(.dout(w_dff_A_EtG2oFGJ4_0),.din(w_dff_A_HYY14ous9_0),.clk(gclk));
	jdff dff_A_EtG2oFGJ4_0(.dout(w_dff_A_y1pevXfH0_0),.din(w_dff_A_EtG2oFGJ4_0),.clk(gclk));
	jdff dff_A_y1pevXfH0_0(.dout(G939),.din(w_dff_A_y1pevXfH0_0),.clk(gclk));
	jdff dff_A_GoPIL2KR7_1(.dout(w_dff_A_DWu12fX50_0),.din(w_dff_A_GoPIL2KR7_1),.clk(gclk));
	jdff dff_A_DWu12fX50_0(.dout(w_dff_A_7LjJ3fMc4_0),.din(w_dff_A_DWu12fX50_0),.clk(gclk));
	jdff dff_A_7LjJ3fMc4_0(.dout(w_dff_A_1tTXvfZ42_0),.din(w_dff_A_7LjJ3fMc4_0),.clk(gclk));
	jdff dff_A_1tTXvfZ42_0(.dout(w_dff_A_fBX5UKo41_0),.din(w_dff_A_1tTXvfZ42_0),.clk(gclk));
	jdff dff_A_fBX5UKo41_0(.dout(w_dff_A_pdI9saIx5_0),.din(w_dff_A_fBX5UKo41_0),.clk(gclk));
	jdff dff_A_pdI9saIx5_0(.dout(w_dff_A_ESBb8mrc3_0),.din(w_dff_A_pdI9saIx5_0),.clk(gclk));
	jdff dff_A_ESBb8mrc3_0(.dout(w_dff_A_m7rtBfeA4_0),.din(w_dff_A_ESBb8mrc3_0),.clk(gclk));
	jdff dff_A_m7rtBfeA4_0(.dout(w_dff_A_xwILDn1Y5_0),.din(w_dff_A_m7rtBfeA4_0),.clk(gclk));
	jdff dff_A_xwILDn1Y5_0(.dout(w_dff_A_PSfK27IH3_0),.din(w_dff_A_xwILDn1Y5_0),.clk(gclk));
	jdff dff_A_PSfK27IH3_0(.dout(w_dff_A_G2Uyhqqk9_0),.din(w_dff_A_PSfK27IH3_0),.clk(gclk));
	jdff dff_A_G2Uyhqqk9_0(.dout(w_dff_A_M75uakEJ4_0),.din(w_dff_A_G2Uyhqqk9_0),.clk(gclk));
	jdff dff_A_M75uakEJ4_0(.dout(w_dff_A_6ZQRETnL8_0),.din(w_dff_A_M75uakEJ4_0),.clk(gclk));
	jdff dff_A_6ZQRETnL8_0(.dout(w_dff_A_un8jIdgZ8_0),.din(w_dff_A_6ZQRETnL8_0),.clk(gclk));
	jdff dff_A_un8jIdgZ8_0(.dout(w_dff_A_hd0DKlqA9_0),.din(w_dff_A_un8jIdgZ8_0),.clk(gclk));
	jdff dff_A_hd0DKlqA9_0(.dout(w_dff_A_auLaSAjA0_0),.din(w_dff_A_hd0DKlqA9_0),.clk(gclk));
	jdff dff_A_auLaSAjA0_0(.dout(w_dff_A_1HORKG3D9_0),.din(w_dff_A_auLaSAjA0_0),.clk(gclk));
	jdff dff_A_1HORKG3D9_0(.dout(w_dff_A_KSJrzDiw1_0),.din(w_dff_A_1HORKG3D9_0),.clk(gclk));
	jdff dff_A_KSJrzDiw1_0(.dout(w_dff_A_n25SCTnO0_0),.din(w_dff_A_KSJrzDiw1_0),.clk(gclk));
	jdff dff_A_n25SCTnO0_0(.dout(w_dff_A_xX4znLr91_0),.din(w_dff_A_n25SCTnO0_0),.clk(gclk));
	jdff dff_A_xX4znLr91_0(.dout(w_dff_A_H1vV2Uvp7_0),.din(w_dff_A_xX4znLr91_0),.clk(gclk));
	jdff dff_A_H1vV2Uvp7_0(.dout(w_dff_A_mgzkWDKP1_0),.din(w_dff_A_H1vV2Uvp7_0),.clk(gclk));
	jdff dff_A_mgzkWDKP1_0(.dout(w_dff_A_IdCbp0QU7_0),.din(w_dff_A_mgzkWDKP1_0),.clk(gclk));
	jdff dff_A_IdCbp0QU7_0(.dout(w_dff_A_NpQUEavQ7_0),.din(w_dff_A_IdCbp0QU7_0),.clk(gclk));
	jdff dff_A_NpQUEavQ7_0(.dout(w_dff_A_YT50ht6T6_0),.din(w_dff_A_NpQUEavQ7_0),.clk(gclk));
	jdff dff_A_YT50ht6T6_0(.dout(w_dff_A_0bNf2yhJ3_0),.din(w_dff_A_YT50ht6T6_0),.clk(gclk));
	jdff dff_A_0bNf2yhJ3_0(.dout(w_dff_A_aMpuROvk1_0),.din(w_dff_A_0bNf2yhJ3_0),.clk(gclk));
	jdff dff_A_aMpuROvk1_0(.dout(w_dff_A_mn5ywUFE7_0),.din(w_dff_A_aMpuROvk1_0),.clk(gclk));
	jdff dff_A_mn5ywUFE7_0(.dout(G889),.din(w_dff_A_mn5ywUFE7_0),.clk(gclk));
	jdff dff_A_ww1qOiDN8_1(.dout(w_dff_A_oZDkyHW71_0),.din(w_dff_A_ww1qOiDN8_1),.clk(gclk));
	jdff dff_A_oZDkyHW71_0(.dout(w_dff_A_4TUklTGv5_0),.din(w_dff_A_oZDkyHW71_0),.clk(gclk));
	jdff dff_A_4TUklTGv5_0(.dout(w_dff_A_IPfPMvhA0_0),.din(w_dff_A_4TUklTGv5_0),.clk(gclk));
	jdff dff_A_IPfPMvhA0_0(.dout(w_dff_A_CFG0Bizp2_0),.din(w_dff_A_IPfPMvhA0_0),.clk(gclk));
	jdff dff_A_CFG0Bizp2_0(.dout(w_dff_A_kQTupb4f6_0),.din(w_dff_A_CFG0Bizp2_0),.clk(gclk));
	jdff dff_A_kQTupb4f6_0(.dout(w_dff_A_lKHZIYm71_0),.din(w_dff_A_kQTupb4f6_0),.clk(gclk));
	jdff dff_A_lKHZIYm71_0(.dout(w_dff_A_JSKTxqCl3_0),.din(w_dff_A_lKHZIYm71_0),.clk(gclk));
	jdff dff_A_JSKTxqCl3_0(.dout(w_dff_A_sX3p9kSR5_0),.din(w_dff_A_JSKTxqCl3_0),.clk(gclk));
	jdff dff_A_sX3p9kSR5_0(.dout(w_dff_A_EJSc661k5_0),.din(w_dff_A_sX3p9kSR5_0),.clk(gclk));
	jdff dff_A_EJSc661k5_0(.dout(w_dff_A_5GxWJpKR5_0),.din(w_dff_A_EJSc661k5_0),.clk(gclk));
	jdff dff_A_5GxWJpKR5_0(.dout(w_dff_A_CFECPB2j4_0),.din(w_dff_A_5GxWJpKR5_0),.clk(gclk));
	jdff dff_A_CFECPB2j4_0(.dout(w_dff_A_TI8ynnxC9_0),.din(w_dff_A_CFECPB2j4_0),.clk(gclk));
	jdff dff_A_TI8ynnxC9_0(.dout(w_dff_A_2OFm0dyj1_0),.din(w_dff_A_TI8ynnxC9_0),.clk(gclk));
	jdff dff_A_2OFm0dyj1_0(.dout(w_dff_A_Ux3NbOna3_0),.din(w_dff_A_2OFm0dyj1_0),.clk(gclk));
	jdff dff_A_Ux3NbOna3_0(.dout(w_dff_A_xJiXxdQC3_0),.din(w_dff_A_Ux3NbOna3_0),.clk(gclk));
	jdff dff_A_xJiXxdQC3_0(.dout(w_dff_A_9pqRgPhB8_0),.din(w_dff_A_xJiXxdQC3_0),.clk(gclk));
	jdff dff_A_9pqRgPhB8_0(.dout(w_dff_A_8aRsQHeo5_0),.din(w_dff_A_9pqRgPhB8_0),.clk(gclk));
	jdff dff_A_8aRsQHeo5_0(.dout(w_dff_A_ZD7TQ8mt0_0),.din(w_dff_A_8aRsQHeo5_0),.clk(gclk));
	jdff dff_A_ZD7TQ8mt0_0(.dout(w_dff_A_zUb32NUd2_0),.din(w_dff_A_ZD7TQ8mt0_0),.clk(gclk));
	jdff dff_A_zUb32NUd2_0(.dout(w_dff_A_wQqfaZfJ7_0),.din(w_dff_A_zUb32NUd2_0),.clk(gclk));
	jdff dff_A_wQqfaZfJ7_0(.dout(w_dff_A_o8ZTUgPI6_0),.din(w_dff_A_wQqfaZfJ7_0),.clk(gclk));
	jdff dff_A_o8ZTUgPI6_0(.dout(w_dff_A_pqDMTDRy9_0),.din(w_dff_A_o8ZTUgPI6_0),.clk(gclk));
	jdff dff_A_pqDMTDRy9_0(.dout(w_dff_A_URQMZIQf7_0),.din(w_dff_A_pqDMTDRy9_0),.clk(gclk));
	jdff dff_A_URQMZIQf7_0(.dout(w_dff_A_vxa3wBMC8_0),.din(w_dff_A_URQMZIQf7_0),.clk(gclk));
	jdff dff_A_vxa3wBMC8_0(.dout(w_dff_A_0EEZoBeP8_0),.din(w_dff_A_vxa3wBMC8_0),.clk(gclk));
	jdff dff_A_0EEZoBeP8_0(.dout(w_dff_A_uNuYueNQ2_0),.din(w_dff_A_0EEZoBeP8_0),.clk(gclk));
	jdff dff_A_uNuYueNQ2_0(.dout(G593),.din(w_dff_A_uNuYueNQ2_0),.clk(gclk));
	jdff dff_A_W2A4HmRM0_2(.dout(w_dff_A_QaVnro5g8_0),.din(w_dff_A_W2A4HmRM0_2),.clk(gclk));
	jdff dff_A_QaVnro5g8_0(.dout(w_dff_A_KxJUxQ7X3_0),.din(w_dff_A_QaVnro5g8_0),.clk(gclk));
	jdff dff_A_KxJUxQ7X3_0(.dout(w_dff_A_j47V9ViA0_0),.din(w_dff_A_KxJUxQ7X3_0),.clk(gclk));
	jdff dff_A_j47V9ViA0_0(.dout(w_dff_A_BQ7zS59F3_0),.din(w_dff_A_j47V9ViA0_0),.clk(gclk));
	jdff dff_A_BQ7zS59F3_0(.dout(w_dff_A_CQFxXwSC1_0),.din(w_dff_A_BQ7zS59F3_0),.clk(gclk));
	jdff dff_A_CQFxXwSC1_0(.dout(w_dff_A_NcKCm2RQ7_0),.din(w_dff_A_CQFxXwSC1_0),.clk(gclk));
	jdff dff_A_NcKCm2RQ7_0(.dout(w_dff_A_RXIdbIa09_0),.din(w_dff_A_NcKCm2RQ7_0),.clk(gclk));
	jdff dff_A_RXIdbIa09_0(.dout(w_dff_A_EHAXu3fA2_0),.din(w_dff_A_RXIdbIa09_0),.clk(gclk));
	jdff dff_A_EHAXu3fA2_0(.dout(w_dff_A_yrCYcxV38_0),.din(w_dff_A_EHAXu3fA2_0),.clk(gclk));
	jdff dff_A_yrCYcxV38_0(.dout(w_dff_A_cFaUsFTi2_0),.din(w_dff_A_yrCYcxV38_0),.clk(gclk));
	jdff dff_A_cFaUsFTi2_0(.dout(w_dff_A_ejI6Ifvq5_0),.din(w_dff_A_cFaUsFTi2_0),.clk(gclk));
	jdff dff_A_ejI6Ifvq5_0(.dout(w_dff_A_yZs6tPzz9_0),.din(w_dff_A_ejI6Ifvq5_0),.clk(gclk));
	jdff dff_A_yZs6tPzz9_0(.dout(w_dff_A_gmhwfYOt8_0),.din(w_dff_A_yZs6tPzz9_0),.clk(gclk));
	jdff dff_A_gmhwfYOt8_0(.dout(w_dff_A_4QCUsUyT2_0),.din(w_dff_A_gmhwfYOt8_0),.clk(gclk));
	jdff dff_A_4QCUsUyT2_0(.dout(w_dff_A_JUk62hAx7_0),.din(w_dff_A_4QCUsUyT2_0),.clk(gclk));
	jdff dff_A_JUk62hAx7_0(.dout(w_dff_A_s3nCDSrv4_0),.din(w_dff_A_JUk62hAx7_0),.clk(gclk));
	jdff dff_A_s3nCDSrv4_0(.dout(w_dff_A_dJo9N0FU0_0),.din(w_dff_A_s3nCDSrv4_0),.clk(gclk));
	jdff dff_A_dJo9N0FU0_0(.dout(w_dff_A_u0ZNj4eS4_0),.din(w_dff_A_dJo9N0FU0_0),.clk(gclk));
	jdff dff_A_u0ZNj4eS4_0(.dout(w_dff_A_Q69Txdew0_0),.din(w_dff_A_u0ZNj4eS4_0),.clk(gclk));
	jdff dff_A_Q69Txdew0_0(.dout(w_dff_A_hbpHU5w69_0),.din(w_dff_A_Q69Txdew0_0),.clk(gclk));
	jdff dff_A_hbpHU5w69_0(.dout(w_dff_A_7JiNTrmT1_0),.din(w_dff_A_hbpHU5w69_0),.clk(gclk));
	jdff dff_A_7JiNTrmT1_0(.dout(w_dff_A_Tg0cR9NZ0_0),.din(w_dff_A_7JiNTrmT1_0),.clk(gclk));
	jdff dff_A_Tg0cR9NZ0_0(.dout(w_dff_A_7DowLR0a1_0),.din(w_dff_A_Tg0cR9NZ0_0),.clk(gclk));
	jdff dff_A_7DowLR0a1_0(.dout(G636),.din(w_dff_A_7DowLR0a1_0),.clk(gclk));
	jdff dff_A_pG90Hqzz7_2(.dout(w_dff_A_gGbUSuHi7_0),.din(w_dff_A_pG90Hqzz7_2),.clk(gclk));
	jdff dff_A_gGbUSuHi7_0(.dout(w_dff_A_387eAaDq7_0),.din(w_dff_A_gGbUSuHi7_0),.clk(gclk));
	jdff dff_A_387eAaDq7_0(.dout(w_dff_A_KfemJT5K1_0),.din(w_dff_A_387eAaDq7_0),.clk(gclk));
	jdff dff_A_KfemJT5K1_0(.dout(w_dff_A_z0fXgH0Q6_0),.din(w_dff_A_KfemJT5K1_0),.clk(gclk));
	jdff dff_A_z0fXgH0Q6_0(.dout(w_dff_A_GlzAHUXK5_0),.din(w_dff_A_z0fXgH0Q6_0),.clk(gclk));
	jdff dff_A_GlzAHUXK5_0(.dout(w_dff_A_EMUK8KtP2_0),.din(w_dff_A_GlzAHUXK5_0),.clk(gclk));
	jdff dff_A_EMUK8KtP2_0(.dout(w_dff_A_PQ5XnzNv5_0),.din(w_dff_A_EMUK8KtP2_0),.clk(gclk));
	jdff dff_A_PQ5XnzNv5_0(.dout(w_dff_A_UELVUXQ85_0),.din(w_dff_A_PQ5XnzNv5_0),.clk(gclk));
	jdff dff_A_UELVUXQ85_0(.dout(w_dff_A_HOTDzVDX0_0),.din(w_dff_A_UELVUXQ85_0),.clk(gclk));
	jdff dff_A_HOTDzVDX0_0(.dout(w_dff_A_C7LMqfjb6_0),.din(w_dff_A_HOTDzVDX0_0),.clk(gclk));
	jdff dff_A_C7LMqfjb6_0(.dout(w_dff_A_CppgYJzX3_0),.din(w_dff_A_C7LMqfjb6_0),.clk(gclk));
	jdff dff_A_CppgYJzX3_0(.dout(w_dff_A_Au4xGyMt6_0),.din(w_dff_A_CppgYJzX3_0),.clk(gclk));
	jdff dff_A_Au4xGyMt6_0(.dout(w_dff_A_vctVRZiB7_0),.din(w_dff_A_Au4xGyMt6_0),.clk(gclk));
	jdff dff_A_vctVRZiB7_0(.dout(w_dff_A_eqlW5oT55_0),.din(w_dff_A_vctVRZiB7_0),.clk(gclk));
	jdff dff_A_eqlW5oT55_0(.dout(w_dff_A_uOzBKZdl6_0),.din(w_dff_A_eqlW5oT55_0),.clk(gclk));
	jdff dff_A_uOzBKZdl6_0(.dout(w_dff_A_N2nUkNAX1_0),.din(w_dff_A_uOzBKZdl6_0),.clk(gclk));
	jdff dff_A_N2nUkNAX1_0(.dout(w_dff_A_l1Kldsk78_0),.din(w_dff_A_N2nUkNAX1_0),.clk(gclk));
	jdff dff_A_l1Kldsk78_0(.dout(w_dff_A_cG5agdGi3_0),.din(w_dff_A_l1Kldsk78_0),.clk(gclk));
	jdff dff_A_cG5agdGi3_0(.dout(w_dff_A_lU5vq53o9_0),.din(w_dff_A_cG5agdGi3_0),.clk(gclk));
	jdff dff_A_lU5vq53o9_0(.dout(w_dff_A_s6joX8Qw8_0),.din(w_dff_A_lU5vq53o9_0),.clk(gclk));
	jdff dff_A_s6joX8Qw8_0(.dout(w_dff_A_kxQeVdnn7_0),.din(w_dff_A_s6joX8Qw8_0),.clk(gclk));
	jdff dff_A_kxQeVdnn7_0(.dout(w_dff_A_A3I2hk9F6_0),.din(w_dff_A_kxQeVdnn7_0),.clk(gclk));
	jdff dff_A_A3I2hk9F6_0(.dout(w_dff_A_Zh1ey7W62_0),.din(w_dff_A_A3I2hk9F6_0),.clk(gclk));
	jdff dff_A_Zh1ey7W62_0(.dout(G704),.din(w_dff_A_Zh1ey7W62_0),.clk(gclk));
	jdff dff_A_m2Bez7pJ5_2(.dout(w_dff_A_IEGiFROW0_0),.din(w_dff_A_m2Bez7pJ5_2),.clk(gclk));
	jdff dff_A_IEGiFROW0_0(.dout(w_dff_A_xsR1Qmcl2_0),.din(w_dff_A_IEGiFROW0_0),.clk(gclk));
	jdff dff_A_xsR1Qmcl2_0(.dout(w_dff_A_yr3sTo9v8_0),.din(w_dff_A_xsR1Qmcl2_0),.clk(gclk));
	jdff dff_A_yr3sTo9v8_0(.dout(w_dff_A_qCBLn4np1_0),.din(w_dff_A_yr3sTo9v8_0),.clk(gclk));
	jdff dff_A_qCBLn4np1_0(.dout(w_dff_A_o7HPenKF7_0),.din(w_dff_A_qCBLn4np1_0),.clk(gclk));
	jdff dff_A_o7HPenKF7_0(.dout(w_dff_A_Mzx3jACP9_0),.din(w_dff_A_o7HPenKF7_0),.clk(gclk));
	jdff dff_A_Mzx3jACP9_0(.dout(w_dff_A_w0Fn9rIC1_0),.din(w_dff_A_Mzx3jACP9_0),.clk(gclk));
	jdff dff_A_w0Fn9rIC1_0(.dout(w_dff_A_PauUkWI95_0),.din(w_dff_A_w0Fn9rIC1_0),.clk(gclk));
	jdff dff_A_PauUkWI95_0(.dout(w_dff_A_zI7cGY9U8_0),.din(w_dff_A_PauUkWI95_0),.clk(gclk));
	jdff dff_A_zI7cGY9U8_0(.dout(w_dff_A_HzI259gW3_0),.din(w_dff_A_zI7cGY9U8_0),.clk(gclk));
	jdff dff_A_HzI259gW3_0(.dout(w_dff_A_vX8f9ZFb7_0),.din(w_dff_A_HzI259gW3_0),.clk(gclk));
	jdff dff_A_vX8f9ZFb7_0(.dout(w_dff_A_tvdyMFT33_0),.din(w_dff_A_vX8f9ZFb7_0),.clk(gclk));
	jdff dff_A_tvdyMFT33_0(.dout(w_dff_A_TbiC2r9n2_0),.din(w_dff_A_tvdyMFT33_0),.clk(gclk));
	jdff dff_A_TbiC2r9n2_0(.dout(w_dff_A_tl90zuMQ3_0),.din(w_dff_A_TbiC2r9n2_0),.clk(gclk));
	jdff dff_A_tl90zuMQ3_0(.dout(w_dff_A_6ylJ5u3G3_0),.din(w_dff_A_tl90zuMQ3_0),.clk(gclk));
	jdff dff_A_6ylJ5u3G3_0(.dout(w_dff_A_SuUos7Yg1_0),.din(w_dff_A_6ylJ5u3G3_0),.clk(gclk));
	jdff dff_A_SuUos7Yg1_0(.dout(w_dff_A_xir742Vt1_0),.din(w_dff_A_SuUos7Yg1_0),.clk(gclk));
	jdff dff_A_xir742Vt1_0(.dout(w_dff_A_khCv8FGo2_0),.din(w_dff_A_xir742Vt1_0),.clk(gclk));
	jdff dff_A_khCv8FGo2_0(.dout(w_dff_A_Xxsm5BjO1_0),.din(w_dff_A_khCv8FGo2_0),.clk(gclk));
	jdff dff_A_Xxsm5BjO1_0(.dout(w_dff_A_DBxV72Lx2_0),.din(w_dff_A_Xxsm5BjO1_0),.clk(gclk));
	jdff dff_A_DBxV72Lx2_0(.dout(w_dff_A_cLLWsM2b5_0),.din(w_dff_A_DBxV72Lx2_0),.clk(gclk));
	jdff dff_A_cLLWsM2b5_0(.dout(w_dff_A_h8tZxkCY8_0),.din(w_dff_A_cLLWsM2b5_0),.clk(gclk));
	jdff dff_A_h8tZxkCY8_0(.dout(w_dff_A_0nS9Lz9c0_0),.din(w_dff_A_h8tZxkCY8_0),.clk(gclk));
	jdff dff_A_0nS9Lz9c0_0(.dout(G717),.din(w_dff_A_0nS9Lz9c0_0),.clk(gclk));
	jdff dff_A_nCW2wrlb6_2(.dout(w_dff_A_rm3mQbX44_0),.din(w_dff_A_nCW2wrlb6_2),.clk(gclk));
	jdff dff_A_rm3mQbX44_0(.dout(w_dff_A_F0Di5moN0_0),.din(w_dff_A_rm3mQbX44_0),.clk(gclk));
	jdff dff_A_F0Di5moN0_0(.dout(w_dff_A_JQSx4VDl1_0),.din(w_dff_A_F0Di5moN0_0),.clk(gclk));
	jdff dff_A_JQSx4VDl1_0(.dout(w_dff_A_abWIZwPH1_0),.din(w_dff_A_JQSx4VDl1_0),.clk(gclk));
	jdff dff_A_abWIZwPH1_0(.dout(w_dff_A_NvYfZVb51_0),.din(w_dff_A_abWIZwPH1_0),.clk(gclk));
	jdff dff_A_NvYfZVb51_0(.dout(w_dff_A_589BAh5Y4_0),.din(w_dff_A_NvYfZVb51_0),.clk(gclk));
	jdff dff_A_589BAh5Y4_0(.dout(w_dff_A_lwOFuML74_0),.din(w_dff_A_589BAh5Y4_0),.clk(gclk));
	jdff dff_A_lwOFuML74_0(.dout(w_dff_A_9948HUf75_0),.din(w_dff_A_lwOFuML74_0),.clk(gclk));
	jdff dff_A_9948HUf75_0(.dout(w_dff_A_E8gbo8A65_0),.din(w_dff_A_9948HUf75_0),.clk(gclk));
	jdff dff_A_E8gbo8A65_0(.dout(w_dff_A_PB0uCKQX2_0),.din(w_dff_A_E8gbo8A65_0),.clk(gclk));
	jdff dff_A_PB0uCKQX2_0(.dout(w_dff_A_E4NRKFz30_0),.din(w_dff_A_PB0uCKQX2_0),.clk(gclk));
	jdff dff_A_E4NRKFz30_0(.dout(w_dff_A_rMFaMdjO9_0),.din(w_dff_A_E4NRKFz30_0),.clk(gclk));
	jdff dff_A_rMFaMdjO9_0(.dout(w_dff_A_X69S294N0_0),.din(w_dff_A_rMFaMdjO9_0),.clk(gclk));
	jdff dff_A_X69S294N0_0(.dout(w_dff_A_rVok3RTO5_0),.din(w_dff_A_X69S294N0_0),.clk(gclk));
	jdff dff_A_rVok3RTO5_0(.dout(w_dff_A_LS5SYU4S1_0),.din(w_dff_A_rVok3RTO5_0),.clk(gclk));
	jdff dff_A_LS5SYU4S1_0(.dout(w_dff_A_z4NDDdqS8_0),.din(w_dff_A_LS5SYU4S1_0),.clk(gclk));
	jdff dff_A_z4NDDdqS8_0(.dout(w_dff_A_XKY1MtsD2_0),.din(w_dff_A_z4NDDdqS8_0),.clk(gclk));
	jdff dff_A_XKY1MtsD2_0(.dout(w_dff_A_z0QBkL9o7_0),.din(w_dff_A_XKY1MtsD2_0),.clk(gclk));
	jdff dff_A_z0QBkL9o7_0(.dout(w_dff_A_ZMnXw3W15_0),.din(w_dff_A_z0QBkL9o7_0),.clk(gclk));
	jdff dff_A_ZMnXw3W15_0(.dout(w_dff_A_mZT2myF72_0),.din(w_dff_A_ZMnXw3W15_0),.clk(gclk));
	jdff dff_A_mZT2myF72_0(.dout(w_dff_A_EB3YUvbq3_0),.din(w_dff_A_mZT2myF72_0),.clk(gclk));
	jdff dff_A_EB3YUvbq3_0(.dout(w_dff_A_FSklPrXv3_0),.din(w_dff_A_EB3YUvbq3_0),.clk(gclk));
	jdff dff_A_FSklPrXv3_0(.dout(w_dff_A_ODiWA8Hz1_0),.din(w_dff_A_FSklPrXv3_0),.clk(gclk));
	jdff dff_A_ODiWA8Hz1_0(.dout(w_dff_A_E2aTN8uK4_0),.din(w_dff_A_ODiWA8Hz1_0),.clk(gclk));
	jdff dff_A_E2aTN8uK4_0(.dout(G820),.din(w_dff_A_E2aTN8uK4_0),.clk(gclk));
	jdff dff_A_K0bgM94k1_2(.dout(w_dff_A_5rCS99ky1_0),.din(w_dff_A_K0bgM94k1_2),.clk(gclk));
	jdff dff_A_5rCS99ky1_0(.dout(w_dff_A_BSH08UoT0_0),.din(w_dff_A_5rCS99ky1_0),.clk(gclk));
	jdff dff_A_BSH08UoT0_0(.dout(w_dff_A_QrvB2chA9_0),.din(w_dff_A_BSH08UoT0_0),.clk(gclk));
	jdff dff_A_QrvB2chA9_0(.dout(w_dff_A_p5b4U0yj4_0),.din(w_dff_A_QrvB2chA9_0),.clk(gclk));
	jdff dff_A_p5b4U0yj4_0(.dout(w_dff_A_mMmAh9ny7_0),.din(w_dff_A_p5b4U0yj4_0),.clk(gclk));
	jdff dff_A_mMmAh9ny7_0(.dout(w_dff_A_27XZIQsn8_0),.din(w_dff_A_mMmAh9ny7_0),.clk(gclk));
	jdff dff_A_27XZIQsn8_0(.dout(w_dff_A_iZztC4bV1_0),.din(w_dff_A_27XZIQsn8_0),.clk(gclk));
	jdff dff_A_iZztC4bV1_0(.dout(w_dff_A_JFmtOsFX6_0),.din(w_dff_A_iZztC4bV1_0),.clk(gclk));
	jdff dff_A_JFmtOsFX6_0(.dout(w_dff_A_UhOa6Xta4_0),.din(w_dff_A_JFmtOsFX6_0),.clk(gclk));
	jdff dff_A_UhOa6Xta4_0(.dout(w_dff_A_p6WqhNZ20_0),.din(w_dff_A_UhOa6Xta4_0),.clk(gclk));
	jdff dff_A_p6WqhNZ20_0(.dout(w_dff_A_3T0JLAE56_0),.din(w_dff_A_p6WqhNZ20_0),.clk(gclk));
	jdff dff_A_3T0JLAE56_0(.dout(w_dff_A_fBcBcyuV8_0),.din(w_dff_A_3T0JLAE56_0),.clk(gclk));
	jdff dff_A_fBcBcyuV8_0(.dout(w_dff_A_lzgitMHS2_0),.din(w_dff_A_fBcBcyuV8_0),.clk(gclk));
	jdff dff_A_lzgitMHS2_0(.dout(w_dff_A_Dgr0O5x92_0),.din(w_dff_A_lzgitMHS2_0),.clk(gclk));
	jdff dff_A_Dgr0O5x92_0(.dout(w_dff_A_BjZtKUNQ8_0),.din(w_dff_A_Dgr0O5x92_0),.clk(gclk));
	jdff dff_A_BjZtKUNQ8_0(.dout(w_dff_A_gD4uF0fg7_0),.din(w_dff_A_BjZtKUNQ8_0),.clk(gclk));
	jdff dff_A_gD4uF0fg7_0(.dout(w_dff_A_xngBk8al9_0),.din(w_dff_A_gD4uF0fg7_0),.clk(gclk));
	jdff dff_A_xngBk8al9_0(.dout(w_dff_A_k5uMO6GB6_0),.din(w_dff_A_xngBk8al9_0),.clk(gclk));
	jdff dff_A_k5uMO6GB6_0(.dout(w_dff_A_Ww1C57Rf7_0),.din(w_dff_A_k5uMO6GB6_0),.clk(gclk));
	jdff dff_A_Ww1C57Rf7_0(.dout(w_dff_A_RtWKg3an9_0),.din(w_dff_A_Ww1C57Rf7_0),.clk(gclk));
	jdff dff_A_RtWKg3an9_0(.dout(w_dff_A_eDcIUdbT6_0),.din(w_dff_A_RtWKg3an9_0),.clk(gclk));
	jdff dff_A_eDcIUdbT6_0(.dout(w_dff_A_LXKUm15T4_0),.din(w_dff_A_eDcIUdbT6_0),.clk(gclk));
	jdff dff_A_LXKUm15T4_0(.dout(G639),.din(w_dff_A_LXKUm15T4_0),.clk(gclk));
	jdff dff_A_ns2r2A0V2_2(.dout(w_dff_A_VtBd6G8p1_0),.din(w_dff_A_ns2r2A0V2_2),.clk(gclk));
	jdff dff_A_VtBd6G8p1_0(.dout(w_dff_A_73VoxK7z4_0),.din(w_dff_A_VtBd6G8p1_0),.clk(gclk));
	jdff dff_A_73VoxK7z4_0(.dout(w_dff_A_idnZIVib4_0),.din(w_dff_A_73VoxK7z4_0),.clk(gclk));
	jdff dff_A_idnZIVib4_0(.dout(w_dff_A_V1URt6g21_0),.din(w_dff_A_idnZIVib4_0),.clk(gclk));
	jdff dff_A_V1URt6g21_0(.dout(w_dff_A_ah69EgPr3_0),.din(w_dff_A_V1URt6g21_0),.clk(gclk));
	jdff dff_A_ah69EgPr3_0(.dout(w_dff_A_Zr4hPuVN7_0),.din(w_dff_A_ah69EgPr3_0),.clk(gclk));
	jdff dff_A_Zr4hPuVN7_0(.dout(w_dff_A_DT8vc6qh1_0),.din(w_dff_A_Zr4hPuVN7_0),.clk(gclk));
	jdff dff_A_DT8vc6qh1_0(.dout(w_dff_A_lgeWYzjY9_0),.din(w_dff_A_DT8vc6qh1_0),.clk(gclk));
	jdff dff_A_lgeWYzjY9_0(.dout(w_dff_A_tX91kvAs7_0),.din(w_dff_A_lgeWYzjY9_0),.clk(gclk));
	jdff dff_A_tX91kvAs7_0(.dout(w_dff_A_AHmpaAUK4_0),.din(w_dff_A_tX91kvAs7_0),.clk(gclk));
	jdff dff_A_AHmpaAUK4_0(.dout(w_dff_A_i54UaYFx6_0),.din(w_dff_A_AHmpaAUK4_0),.clk(gclk));
	jdff dff_A_i54UaYFx6_0(.dout(w_dff_A_kRQ57SEZ2_0),.din(w_dff_A_i54UaYFx6_0),.clk(gclk));
	jdff dff_A_kRQ57SEZ2_0(.dout(w_dff_A_cMSEExtz6_0),.din(w_dff_A_kRQ57SEZ2_0),.clk(gclk));
	jdff dff_A_cMSEExtz6_0(.dout(w_dff_A_CjLEOFgY2_0),.din(w_dff_A_cMSEExtz6_0),.clk(gclk));
	jdff dff_A_CjLEOFgY2_0(.dout(w_dff_A_Bzqt97gV6_0),.din(w_dff_A_CjLEOFgY2_0),.clk(gclk));
	jdff dff_A_Bzqt97gV6_0(.dout(w_dff_A_xJnbnE3e0_0),.din(w_dff_A_Bzqt97gV6_0),.clk(gclk));
	jdff dff_A_xJnbnE3e0_0(.dout(w_dff_A_trAH1DME2_0),.din(w_dff_A_xJnbnE3e0_0),.clk(gclk));
	jdff dff_A_trAH1DME2_0(.dout(w_dff_A_RWTfoV1Q4_0),.din(w_dff_A_trAH1DME2_0),.clk(gclk));
	jdff dff_A_RWTfoV1Q4_0(.dout(w_dff_A_RPFYHpfd9_0),.din(w_dff_A_RWTfoV1Q4_0),.clk(gclk));
	jdff dff_A_RPFYHpfd9_0(.dout(w_dff_A_99AewqOf5_0),.din(w_dff_A_RPFYHpfd9_0),.clk(gclk));
	jdff dff_A_99AewqOf5_0(.dout(w_dff_A_PREqOKbW0_0),.din(w_dff_A_99AewqOf5_0),.clk(gclk));
	jdff dff_A_PREqOKbW0_0(.dout(w_dff_A_Yiu8GeYD4_0),.din(w_dff_A_PREqOKbW0_0),.clk(gclk));
	jdff dff_A_Yiu8GeYD4_0(.dout(G673),.din(w_dff_A_Yiu8GeYD4_0),.clk(gclk));
	jdff dff_A_EboTNr2L1_2(.dout(w_dff_A_agnvmFPa9_0),.din(w_dff_A_EboTNr2L1_2),.clk(gclk));
	jdff dff_A_agnvmFPa9_0(.dout(w_dff_A_oLUkG5Md2_0),.din(w_dff_A_agnvmFPa9_0),.clk(gclk));
	jdff dff_A_oLUkG5Md2_0(.dout(w_dff_A_XurTHM0r8_0),.din(w_dff_A_oLUkG5Md2_0),.clk(gclk));
	jdff dff_A_XurTHM0r8_0(.dout(w_dff_A_5iFLZdds0_0),.din(w_dff_A_XurTHM0r8_0),.clk(gclk));
	jdff dff_A_5iFLZdds0_0(.dout(w_dff_A_zCqjhmeL4_0),.din(w_dff_A_5iFLZdds0_0),.clk(gclk));
	jdff dff_A_zCqjhmeL4_0(.dout(w_dff_A_7cbJ3MdY6_0),.din(w_dff_A_zCqjhmeL4_0),.clk(gclk));
	jdff dff_A_7cbJ3MdY6_0(.dout(w_dff_A_aHCI1Iem1_0),.din(w_dff_A_7cbJ3MdY6_0),.clk(gclk));
	jdff dff_A_aHCI1Iem1_0(.dout(w_dff_A_Y3CTJq573_0),.din(w_dff_A_aHCI1Iem1_0),.clk(gclk));
	jdff dff_A_Y3CTJq573_0(.dout(w_dff_A_LDLh5m0v8_0),.din(w_dff_A_Y3CTJq573_0),.clk(gclk));
	jdff dff_A_LDLh5m0v8_0(.dout(w_dff_A_QFaYvZKE0_0),.din(w_dff_A_LDLh5m0v8_0),.clk(gclk));
	jdff dff_A_QFaYvZKE0_0(.dout(w_dff_A_JQOqABNp9_0),.din(w_dff_A_QFaYvZKE0_0),.clk(gclk));
	jdff dff_A_JQOqABNp9_0(.dout(w_dff_A_ztmzWzrH5_0),.din(w_dff_A_JQOqABNp9_0),.clk(gclk));
	jdff dff_A_ztmzWzrH5_0(.dout(w_dff_A_u1ToTu1r3_0),.din(w_dff_A_ztmzWzrH5_0),.clk(gclk));
	jdff dff_A_u1ToTu1r3_0(.dout(w_dff_A_93jyY1ri6_0),.din(w_dff_A_u1ToTu1r3_0),.clk(gclk));
	jdff dff_A_93jyY1ri6_0(.dout(w_dff_A_R56LuyJI4_0),.din(w_dff_A_93jyY1ri6_0),.clk(gclk));
	jdff dff_A_R56LuyJI4_0(.dout(w_dff_A_FmbYh5YL4_0),.din(w_dff_A_R56LuyJI4_0),.clk(gclk));
	jdff dff_A_FmbYh5YL4_0(.dout(w_dff_A_Y62OhfTG7_0),.din(w_dff_A_FmbYh5YL4_0),.clk(gclk));
	jdff dff_A_Y62OhfTG7_0(.dout(w_dff_A_xekOnK9u1_0),.din(w_dff_A_Y62OhfTG7_0),.clk(gclk));
	jdff dff_A_xekOnK9u1_0(.dout(w_dff_A_CUwA76FH3_0),.din(w_dff_A_xekOnK9u1_0),.clk(gclk));
	jdff dff_A_CUwA76FH3_0(.dout(w_dff_A_5t41Rj8X3_0),.din(w_dff_A_CUwA76FH3_0),.clk(gclk));
	jdff dff_A_5t41Rj8X3_0(.dout(w_dff_A_iImP5izh9_0),.din(w_dff_A_5t41Rj8X3_0),.clk(gclk));
	jdff dff_A_iImP5izh9_0(.dout(w_dff_A_vurdxdhW5_0),.din(w_dff_A_iImP5izh9_0),.clk(gclk));
	jdff dff_A_vurdxdhW5_0(.dout(G707),.din(w_dff_A_vurdxdhW5_0),.clk(gclk));
	jdff dff_A_irTx5kiE2_2(.dout(w_dff_A_qxO0PH441_0),.din(w_dff_A_irTx5kiE2_2),.clk(gclk));
	jdff dff_A_qxO0PH441_0(.dout(w_dff_A_6Af8R8TV2_0),.din(w_dff_A_qxO0PH441_0),.clk(gclk));
	jdff dff_A_6Af8R8TV2_0(.dout(w_dff_A_PDemwxST6_0),.din(w_dff_A_6Af8R8TV2_0),.clk(gclk));
	jdff dff_A_PDemwxST6_0(.dout(w_dff_A_2tZQv2C57_0),.din(w_dff_A_PDemwxST6_0),.clk(gclk));
	jdff dff_A_2tZQv2C57_0(.dout(w_dff_A_DgNsWwQf2_0),.din(w_dff_A_2tZQv2C57_0),.clk(gclk));
	jdff dff_A_DgNsWwQf2_0(.dout(w_dff_A_YxBL8Wh46_0),.din(w_dff_A_DgNsWwQf2_0),.clk(gclk));
	jdff dff_A_YxBL8Wh46_0(.dout(w_dff_A_vKrnwEKv9_0),.din(w_dff_A_YxBL8Wh46_0),.clk(gclk));
	jdff dff_A_vKrnwEKv9_0(.dout(w_dff_A_U6qTqqy10_0),.din(w_dff_A_vKrnwEKv9_0),.clk(gclk));
	jdff dff_A_U6qTqqy10_0(.dout(w_dff_A_2eqGKT7x7_0),.din(w_dff_A_U6qTqqy10_0),.clk(gclk));
	jdff dff_A_2eqGKT7x7_0(.dout(w_dff_A_RsUMXBdf1_0),.din(w_dff_A_2eqGKT7x7_0),.clk(gclk));
	jdff dff_A_RsUMXBdf1_0(.dout(w_dff_A_I0NM0qeH8_0),.din(w_dff_A_RsUMXBdf1_0),.clk(gclk));
	jdff dff_A_I0NM0qeH8_0(.dout(w_dff_A_faklq2lQ6_0),.din(w_dff_A_I0NM0qeH8_0),.clk(gclk));
	jdff dff_A_faklq2lQ6_0(.dout(w_dff_A_rJkfP4yh6_0),.din(w_dff_A_faklq2lQ6_0),.clk(gclk));
	jdff dff_A_rJkfP4yh6_0(.dout(w_dff_A_Lp1MU6EB5_0),.din(w_dff_A_rJkfP4yh6_0),.clk(gclk));
	jdff dff_A_Lp1MU6EB5_0(.dout(w_dff_A_3OkrusRu1_0),.din(w_dff_A_Lp1MU6EB5_0),.clk(gclk));
	jdff dff_A_3OkrusRu1_0(.dout(w_dff_A_zUACS2GE0_0),.din(w_dff_A_3OkrusRu1_0),.clk(gclk));
	jdff dff_A_zUACS2GE0_0(.dout(w_dff_A_JDIWKMuP2_0),.din(w_dff_A_zUACS2GE0_0),.clk(gclk));
	jdff dff_A_JDIWKMuP2_0(.dout(w_dff_A_SJRFcrx57_0),.din(w_dff_A_JDIWKMuP2_0),.clk(gclk));
	jdff dff_A_SJRFcrx57_0(.dout(w_dff_A_KrNVv2cv0_0),.din(w_dff_A_SJRFcrx57_0),.clk(gclk));
	jdff dff_A_KrNVv2cv0_0(.dout(w_dff_A_knLz9pCg4_0),.din(w_dff_A_KrNVv2cv0_0),.clk(gclk));
	jdff dff_A_knLz9pCg4_0(.dout(w_dff_A_YXskZwlQ4_0),.din(w_dff_A_knLz9pCg4_0),.clk(gclk));
	jdff dff_A_YXskZwlQ4_0(.dout(w_dff_A_7sbpixWh0_0),.din(w_dff_A_YXskZwlQ4_0),.clk(gclk));
	jdff dff_A_7sbpixWh0_0(.dout(G715),.din(w_dff_A_7sbpixWh0_0),.clk(gclk));
	jdff dff_A_n5rTAWwz1_2(.dout(w_dff_A_OitPnp5b6_0),.din(w_dff_A_n5rTAWwz1_2),.clk(gclk));
	jdff dff_A_OitPnp5b6_0(.dout(w_dff_A_Ulv1AIIe5_0),.din(w_dff_A_OitPnp5b6_0),.clk(gclk));
	jdff dff_A_Ulv1AIIe5_0(.dout(w_dff_A_cSCjgSiO6_0),.din(w_dff_A_Ulv1AIIe5_0),.clk(gclk));
	jdff dff_A_cSCjgSiO6_0(.dout(w_dff_A_Rg3GDdbw3_0),.din(w_dff_A_cSCjgSiO6_0),.clk(gclk));
	jdff dff_A_Rg3GDdbw3_0(.dout(w_dff_A_TFxvzmYG6_0),.din(w_dff_A_Rg3GDdbw3_0),.clk(gclk));
	jdff dff_A_TFxvzmYG6_0(.dout(w_dff_A_6TOXXDxv9_0),.din(w_dff_A_TFxvzmYG6_0),.clk(gclk));
	jdff dff_A_6TOXXDxv9_0(.dout(w_dff_A_TYKCbDKs9_0),.din(w_dff_A_6TOXXDxv9_0),.clk(gclk));
	jdff dff_A_TYKCbDKs9_0(.dout(w_dff_A_WQlnJwOw5_0),.din(w_dff_A_TYKCbDKs9_0),.clk(gclk));
	jdff dff_A_WQlnJwOw5_0(.dout(w_dff_A_DktPXKxr7_0),.din(w_dff_A_WQlnJwOw5_0),.clk(gclk));
	jdff dff_A_DktPXKxr7_0(.dout(w_dff_A_oCnjY3oC6_0),.din(w_dff_A_DktPXKxr7_0),.clk(gclk));
	jdff dff_A_oCnjY3oC6_0(.dout(w_dff_A_krxf78v44_0),.din(w_dff_A_oCnjY3oC6_0),.clk(gclk));
	jdff dff_A_krxf78v44_0(.dout(w_dff_A_QpOltkc82_0),.din(w_dff_A_krxf78v44_0),.clk(gclk));
	jdff dff_A_QpOltkc82_0(.dout(w_dff_A_9XmaKbEu5_0),.din(w_dff_A_QpOltkc82_0),.clk(gclk));
	jdff dff_A_9XmaKbEu5_0(.dout(w_dff_A_Bg0I2PMk3_0),.din(w_dff_A_9XmaKbEu5_0),.clk(gclk));
	jdff dff_A_Bg0I2PMk3_0(.dout(w_dff_A_DOtYBabN3_0),.din(w_dff_A_Bg0I2PMk3_0),.clk(gclk));
	jdff dff_A_DOtYBabN3_0(.dout(w_dff_A_S0xPbrrl1_0),.din(w_dff_A_DOtYBabN3_0),.clk(gclk));
	jdff dff_A_S0xPbrrl1_0(.dout(w_dff_A_gr5JutjT0_0),.din(w_dff_A_S0xPbrrl1_0),.clk(gclk));
	jdff dff_A_gr5JutjT0_0(.dout(w_dff_A_FXVMSB5l1_0),.din(w_dff_A_gr5JutjT0_0),.clk(gclk));
	jdff dff_A_FXVMSB5l1_0(.dout(w_dff_A_WWiGWFJq0_0),.din(w_dff_A_FXVMSB5l1_0),.clk(gclk));
	jdff dff_A_WWiGWFJq0_0(.dout(G598),.din(w_dff_A_WWiGWFJq0_0),.clk(gclk));
	jdff dff_A_nrahmVjl6_2(.dout(w_dff_A_gJNmfqdw2_0),.din(w_dff_A_nrahmVjl6_2),.clk(gclk));
	jdff dff_A_gJNmfqdw2_0(.dout(w_dff_A_r4LJK7Qq3_0),.din(w_dff_A_gJNmfqdw2_0),.clk(gclk));
	jdff dff_A_r4LJK7Qq3_0(.dout(w_dff_A_xBT7N27k6_0),.din(w_dff_A_r4LJK7Qq3_0),.clk(gclk));
	jdff dff_A_xBT7N27k6_0(.dout(w_dff_A_77Cebwvq4_0),.din(w_dff_A_xBT7N27k6_0),.clk(gclk));
	jdff dff_A_77Cebwvq4_0(.dout(w_dff_A_DUBoqliQ4_0),.din(w_dff_A_77Cebwvq4_0),.clk(gclk));
	jdff dff_A_DUBoqliQ4_0(.dout(w_dff_A_QpCZgQQK4_0),.din(w_dff_A_DUBoqliQ4_0),.clk(gclk));
	jdff dff_A_QpCZgQQK4_0(.dout(w_dff_A_kexmRSBR3_0),.din(w_dff_A_QpCZgQQK4_0),.clk(gclk));
	jdff dff_A_kexmRSBR3_0(.dout(w_dff_A_FnWcXVaO8_0),.din(w_dff_A_kexmRSBR3_0),.clk(gclk));
	jdff dff_A_FnWcXVaO8_0(.dout(w_dff_A_lTAyseaB6_0),.din(w_dff_A_FnWcXVaO8_0),.clk(gclk));
	jdff dff_A_lTAyseaB6_0(.dout(w_dff_A_nTHi0pZl9_0),.din(w_dff_A_lTAyseaB6_0),.clk(gclk));
	jdff dff_A_nTHi0pZl9_0(.dout(w_dff_A_i0wTYvHg5_0),.din(w_dff_A_nTHi0pZl9_0),.clk(gclk));
	jdff dff_A_i0wTYvHg5_0(.dout(w_dff_A_1MU40sgG8_0),.din(w_dff_A_i0wTYvHg5_0),.clk(gclk));
	jdff dff_A_1MU40sgG8_0(.dout(w_dff_A_RLp9M79N2_0),.din(w_dff_A_1MU40sgG8_0),.clk(gclk));
	jdff dff_A_RLp9M79N2_0(.dout(w_dff_A_i7Iqz03p8_0),.din(w_dff_A_RLp9M79N2_0),.clk(gclk));
	jdff dff_A_i7Iqz03p8_0(.dout(w_dff_A_HJXsng5R6_0),.din(w_dff_A_i7Iqz03p8_0),.clk(gclk));
	jdff dff_A_HJXsng5R6_0(.dout(w_dff_A_nfrFDF2U4_0),.din(w_dff_A_HJXsng5R6_0),.clk(gclk));
	jdff dff_A_nfrFDF2U4_0(.dout(w_dff_A_9oS0Va600_0),.din(w_dff_A_nfrFDF2U4_0),.clk(gclk));
	jdff dff_A_9oS0Va600_0(.dout(w_dff_A_RxNMsRf29_0),.din(w_dff_A_9oS0Va600_0),.clk(gclk));
	jdff dff_A_RxNMsRf29_0(.dout(G610),.din(w_dff_A_RxNMsRf29_0),.clk(gclk));
	jdff dff_A_RHR5feu64_2(.dout(w_dff_A_fF6Xt8aN2_0),.din(w_dff_A_RHR5feu64_2),.clk(gclk));
	jdff dff_A_fF6Xt8aN2_0(.dout(w_dff_A_JqVYQZuN9_0),.din(w_dff_A_fF6Xt8aN2_0),.clk(gclk));
	jdff dff_A_JqVYQZuN9_0(.dout(w_dff_A_H420Pagp6_0),.din(w_dff_A_JqVYQZuN9_0),.clk(gclk));
	jdff dff_A_H420Pagp6_0(.dout(w_dff_A_aXamRz1Q6_0),.din(w_dff_A_H420Pagp6_0),.clk(gclk));
	jdff dff_A_aXamRz1Q6_0(.dout(w_dff_A_lIoPnAyI0_0),.din(w_dff_A_aXamRz1Q6_0),.clk(gclk));
	jdff dff_A_lIoPnAyI0_0(.dout(w_dff_A_kvSIjSbT2_0),.din(w_dff_A_lIoPnAyI0_0),.clk(gclk));
	jdff dff_A_kvSIjSbT2_0(.dout(w_dff_A_up1A3Lm06_0),.din(w_dff_A_kvSIjSbT2_0),.clk(gclk));
	jdff dff_A_up1A3Lm06_0(.dout(w_dff_A_DZlFkdvP0_0),.din(w_dff_A_up1A3Lm06_0),.clk(gclk));
	jdff dff_A_DZlFkdvP0_0(.dout(w_dff_A_C85mTphH5_0),.din(w_dff_A_DZlFkdvP0_0),.clk(gclk));
	jdff dff_A_C85mTphH5_0(.dout(w_dff_A_6ePqGiPn9_0),.din(w_dff_A_C85mTphH5_0),.clk(gclk));
	jdff dff_A_6ePqGiPn9_0(.dout(w_dff_A_4aMRgxII0_0),.din(w_dff_A_6ePqGiPn9_0),.clk(gclk));
	jdff dff_A_4aMRgxII0_0(.dout(w_dff_A_jPfzc2ib4_0),.din(w_dff_A_4aMRgxII0_0),.clk(gclk));
	jdff dff_A_jPfzc2ib4_0(.dout(w_dff_A_ST4ndAa71_0),.din(w_dff_A_jPfzc2ib4_0),.clk(gclk));
	jdff dff_A_ST4ndAa71_0(.dout(w_dff_A_cE1E5OSF7_0),.din(w_dff_A_ST4ndAa71_0),.clk(gclk));
	jdff dff_A_cE1E5OSF7_0(.dout(w_dff_A_E2xsAdWp7_0),.din(w_dff_A_cE1E5OSF7_0),.clk(gclk));
	jdff dff_A_E2xsAdWp7_0(.dout(w_dff_A_zJENpbXn5_0),.din(w_dff_A_E2xsAdWp7_0),.clk(gclk));
	jdff dff_A_zJENpbXn5_0(.dout(G588),.din(w_dff_A_zJENpbXn5_0),.clk(gclk));
	jdff dff_A_QCJjv6qE4_2(.dout(w_dff_A_0noHcg101_0),.din(w_dff_A_QCJjv6qE4_2),.clk(gclk));
	jdff dff_A_0noHcg101_0(.dout(w_dff_A_6wgbPrYP3_0),.din(w_dff_A_0noHcg101_0),.clk(gclk));
	jdff dff_A_6wgbPrYP3_0(.dout(w_dff_A_2Ghlu4Eg8_0),.din(w_dff_A_6wgbPrYP3_0),.clk(gclk));
	jdff dff_A_2Ghlu4Eg8_0(.dout(w_dff_A_cKMaclMw9_0),.din(w_dff_A_2Ghlu4Eg8_0),.clk(gclk));
	jdff dff_A_cKMaclMw9_0(.dout(w_dff_A_7gzxcZtL7_0),.din(w_dff_A_cKMaclMw9_0),.clk(gclk));
	jdff dff_A_7gzxcZtL7_0(.dout(w_dff_A_05TkpdN03_0),.din(w_dff_A_7gzxcZtL7_0),.clk(gclk));
	jdff dff_A_05TkpdN03_0(.dout(w_dff_A_vBGTO0xF7_0),.din(w_dff_A_05TkpdN03_0),.clk(gclk));
	jdff dff_A_vBGTO0xF7_0(.dout(w_dff_A_gFNU69yT3_0),.din(w_dff_A_vBGTO0xF7_0),.clk(gclk));
	jdff dff_A_gFNU69yT3_0(.dout(w_dff_A_lmAvD1OV4_0),.din(w_dff_A_gFNU69yT3_0),.clk(gclk));
	jdff dff_A_lmAvD1OV4_0(.dout(w_dff_A_mDzFsg8Z9_0),.din(w_dff_A_lmAvD1OV4_0),.clk(gclk));
	jdff dff_A_mDzFsg8Z9_0(.dout(w_dff_A_hF25cm8s4_0),.din(w_dff_A_mDzFsg8Z9_0),.clk(gclk));
	jdff dff_A_hF25cm8s4_0(.dout(w_dff_A_uC5iMHRi3_0),.din(w_dff_A_hF25cm8s4_0),.clk(gclk));
	jdff dff_A_uC5iMHRi3_0(.dout(w_dff_A_GI4CL9851_0),.din(w_dff_A_uC5iMHRi3_0),.clk(gclk));
	jdff dff_A_GI4CL9851_0(.dout(w_dff_A_xZFobIqm7_0),.din(w_dff_A_GI4CL9851_0),.clk(gclk));
	jdff dff_A_xZFobIqm7_0(.dout(w_dff_A_09bONyQn2_0),.din(w_dff_A_xZFobIqm7_0),.clk(gclk));
	jdff dff_A_09bONyQn2_0(.dout(w_dff_A_vZUqpITH7_0),.din(w_dff_A_09bONyQn2_0),.clk(gclk));
	jdff dff_A_vZUqpITH7_0(.dout(w_dff_A_Khh3TTeo2_0),.din(w_dff_A_vZUqpITH7_0),.clk(gclk));
	jdff dff_A_Khh3TTeo2_0(.dout(G615),.din(w_dff_A_Khh3TTeo2_0),.clk(gclk));
	jdff dff_A_Dg5KC4an0_2(.dout(w_dff_A_eHVHO0sT1_0),.din(w_dff_A_Dg5KC4an0_2),.clk(gclk));
	jdff dff_A_eHVHO0sT1_0(.dout(w_dff_A_UCT4t5Rf2_0),.din(w_dff_A_eHVHO0sT1_0),.clk(gclk));
	jdff dff_A_UCT4t5Rf2_0(.dout(w_dff_A_jZTUOCdY8_0),.din(w_dff_A_UCT4t5Rf2_0),.clk(gclk));
	jdff dff_A_jZTUOCdY8_0(.dout(w_dff_A_66NDokpo9_0),.din(w_dff_A_jZTUOCdY8_0),.clk(gclk));
	jdff dff_A_66NDokpo9_0(.dout(w_dff_A_u2qcZ0eh1_0),.din(w_dff_A_66NDokpo9_0),.clk(gclk));
	jdff dff_A_u2qcZ0eh1_0(.dout(w_dff_A_miumCsT48_0),.din(w_dff_A_u2qcZ0eh1_0),.clk(gclk));
	jdff dff_A_miumCsT48_0(.dout(w_dff_A_z3shtDXP9_0),.din(w_dff_A_miumCsT48_0),.clk(gclk));
	jdff dff_A_z3shtDXP9_0(.dout(w_dff_A_GgbdXAIj5_0),.din(w_dff_A_z3shtDXP9_0),.clk(gclk));
	jdff dff_A_GgbdXAIj5_0(.dout(w_dff_A_2cWTen6x2_0),.din(w_dff_A_GgbdXAIj5_0),.clk(gclk));
	jdff dff_A_2cWTen6x2_0(.dout(w_dff_A_S48hZHOi3_0),.din(w_dff_A_2cWTen6x2_0),.clk(gclk));
	jdff dff_A_S48hZHOi3_0(.dout(w_dff_A_uIOD6Wp56_0),.din(w_dff_A_S48hZHOi3_0),.clk(gclk));
	jdff dff_A_uIOD6Wp56_0(.dout(w_dff_A_5S5U2Q2c1_0),.din(w_dff_A_uIOD6Wp56_0),.clk(gclk));
	jdff dff_A_5S5U2Q2c1_0(.dout(w_dff_A_A0V4sbjp7_0),.din(w_dff_A_5S5U2Q2c1_0),.clk(gclk));
	jdff dff_A_A0V4sbjp7_0(.dout(w_dff_A_Gb4QojF33_0),.din(w_dff_A_A0V4sbjp7_0),.clk(gclk));
	jdff dff_A_Gb4QojF33_0(.dout(w_dff_A_OOOwFFxb5_0),.din(w_dff_A_Gb4QojF33_0),.clk(gclk));
	jdff dff_A_OOOwFFxb5_0(.dout(w_dff_A_1qyQ6q1M1_0),.din(w_dff_A_OOOwFFxb5_0),.clk(gclk));
	jdff dff_A_1qyQ6q1M1_0(.dout(w_dff_A_e0MEue5I5_0),.din(w_dff_A_1qyQ6q1M1_0),.clk(gclk));
	jdff dff_A_e0MEue5I5_0(.dout(G626),.din(w_dff_A_e0MEue5I5_0),.clk(gclk));
	jdff dff_A_zX1uAcE31_2(.dout(w_dff_A_fw9UzGh89_0),.din(w_dff_A_zX1uAcE31_2),.clk(gclk));
	jdff dff_A_fw9UzGh89_0(.dout(w_dff_A_ZGTPVf9W2_0),.din(w_dff_A_fw9UzGh89_0),.clk(gclk));
	jdff dff_A_ZGTPVf9W2_0(.dout(w_dff_A_DGHH1tyM2_0),.din(w_dff_A_ZGTPVf9W2_0),.clk(gclk));
	jdff dff_A_DGHH1tyM2_0(.dout(w_dff_A_pxCO5q8I4_0),.din(w_dff_A_DGHH1tyM2_0),.clk(gclk));
	jdff dff_A_pxCO5q8I4_0(.dout(w_dff_A_d4sdXjMy7_0),.din(w_dff_A_pxCO5q8I4_0),.clk(gclk));
	jdff dff_A_d4sdXjMy7_0(.dout(w_dff_A_tq84brqH5_0),.din(w_dff_A_d4sdXjMy7_0),.clk(gclk));
	jdff dff_A_tq84brqH5_0(.dout(w_dff_A_QzRkFl9R9_0),.din(w_dff_A_tq84brqH5_0),.clk(gclk));
	jdff dff_A_QzRkFl9R9_0(.dout(w_dff_A_qTlI0DBE0_0),.din(w_dff_A_QzRkFl9R9_0),.clk(gclk));
	jdff dff_A_qTlI0DBE0_0(.dout(w_dff_A_MhIHG7kR8_0),.din(w_dff_A_qTlI0DBE0_0),.clk(gclk));
	jdff dff_A_MhIHG7kR8_0(.dout(w_dff_A_SKHzLK3b9_0),.din(w_dff_A_MhIHG7kR8_0),.clk(gclk));
	jdff dff_A_SKHzLK3b9_0(.dout(w_dff_A_68nPV9O08_0),.din(w_dff_A_SKHzLK3b9_0),.clk(gclk));
	jdff dff_A_68nPV9O08_0(.dout(w_dff_A_c7OrDsHw1_0),.din(w_dff_A_68nPV9O08_0),.clk(gclk));
	jdff dff_A_c7OrDsHw1_0(.dout(w_dff_A_CL1eNI2R0_0),.din(w_dff_A_c7OrDsHw1_0),.clk(gclk));
	jdff dff_A_CL1eNI2R0_0(.dout(w_dff_A_2IPaDmAB2_0),.din(w_dff_A_CL1eNI2R0_0),.clk(gclk));
	jdff dff_A_2IPaDmAB2_0(.dout(w_dff_A_ZPU5Q32r8_0),.din(w_dff_A_2IPaDmAB2_0),.clk(gclk));
	jdff dff_A_ZPU5Q32r8_0(.dout(w_dff_A_J06MSiW32_0),.din(w_dff_A_ZPU5Q32r8_0),.clk(gclk));
	jdff dff_A_J06MSiW32_0(.dout(G632),.din(w_dff_A_J06MSiW32_0),.clk(gclk));
	jdff dff_A_hM9YJ7h17_1(.dout(w_dff_A_1zHWn9Mh3_0),.din(w_dff_A_hM9YJ7h17_1),.clk(gclk));
	jdff dff_A_1zHWn9Mh3_0(.dout(w_dff_A_bncCssNd8_0),.din(w_dff_A_1zHWn9Mh3_0),.clk(gclk));
	jdff dff_A_bncCssNd8_0(.dout(w_dff_A_HJk9iyZJ4_0),.din(w_dff_A_bncCssNd8_0),.clk(gclk));
	jdff dff_A_HJk9iyZJ4_0(.dout(w_dff_A_nBradd275_0),.din(w_dff_A_HJk9iyZJ4_0),.clk(gclk));
	jdff dff_A_nBradd275_0(.dout(w_dff_A_v4H21F0A9_0),.din(w_dff_A_nBradd275_0),.clk(gclk));
	jdff dff_A_v4H21F0A9_0(.dout(w_dff_A_RAFoCmNz3_0),.din(w_dff_A_v4H21F0A9_0),.clk(gclk));
	jdff dff_A_RAFoCmNz3_0(.dout(w_dff_A_ObdjxysS5_0),.din(w_dff_A_RAFoCmNz3_0),.clk(gclk));
	jdff dff_A_ObdjxysS5_0(.dout(w_dff_A_mtTWLdfV8_0),.din(w_dff_A_ObdjxysS5_0),.clk(gclk));
	jdff dff_A_mtTWLdfV8_0(.dout(w_dff_A_PFS7FIlM2_0),.din(w_dff_A_mtTWLdfV8_0),.clk(gclk));
	jdff dff_A_PFS7FIlM2_0(.dout(w_dff_A_iFjQS5Dp9_0),.din(w_dff_A_PFS7FIlM2_0),.clk(gclk));
	jdff dff_A_iFjQS5Dp9_0(.dout(w_dff_A_KoroU8UW1_0),.din(w_dff_A_iFjQS5Dp9_0),.clk(gclk));
	jdff dff_A_KoroU8UW1_0(.dout(w_dff_A_X4pDVrFQ6_0),.din(w_dff_A_KoroU8UW1_0),.clk(gclk));
	jdff dff_A_X4pDVrFQ6_0(.dout(w_dff_A_cgDj8fhF2_0),.din(w_dff_A_X4pDVrFQ6_0),.clk(gclk));
	jdff dff_A_cgDj8fhF2_0(.dout(w_dff_A_FVSw9pZ65_0),.din(w_dff_A_cgDj8fhF2_0),.clk(gclk));
	jdff dff_A_FVSw9pZ65_0(.dout(w_dff_A_covnFvY72_0),.din(w_dff_A_FVSw9pZ65_0),.clk(gclk));
	jdff dff_A_covnFvY72_0(.dout(w_dff_A_LNodNHtu9_0),.din(w_dff_A_covnFvY72_0),.clk(gclk));
	jdff dff_A_LNodNHtu9_0(.dout(w_dff_A_wIdL56Et2_0),.din(w_dff_A_LNodNHtu9_0),.clk(gclk));
	jdff dff_A_wIdL56Et2_0(.dout(w_dff_A_qJbiZyYs6_0),.din(w_dff_A_wIdL56Et2_0),.clk(gclk));
	jdff dff_A_qJbiZyYs6_0(.dout(w_dff_A_vp4rglR89_0),.din(w_dff_A_qJbiZyYs6_0),.clk(gclk));
	jdff dff_A_vp4rglR89_0(.dout(w_dff_A_v8mPjnKV5_0),.din(w_dff_A_vp4rglR89_0),.clk(gclk));
	jdff dff_A_v8mPjnKV5_0(.dout(w_dff_A_sBTcLB2d4_0),.din(w_dff_A_v8mPjnKV5_0),.clk(gclk));
	jdff dff_A_sBTcLB2d4_0(.dout(w_dff_A_E28C4AF21_0),.din(w_dff_A_sBTcLB2d4_0),.clk(gclk));
	jdff dff_A_E28C4AF21_0(.dout(G1002),.din(w_dff_A_E28C4AF21_0),.clk(gclk));
	jdff dff_A_2qWiafb32_1(.dout(w_dff_A_SEkelveQ6_0),.din(w_dff_A_2qWiafb32_1),.clk(gclk));
	jdff dff_A_SEkelveQ6_0(.dout(w_dff_A_syackUCF5_0),.din(w_dff_A_SEkelveQ6_0),.clk(gclk));
	jdff dff_A_syackUCF5_0(.dout(w_dff_A_mZEO4lcH5_0),.din(w_dff_A_syackUCF5_0),.clk(gclk));
	jdff dff_A_mZEO4lcH5_0(.dout(w_dff_A_Qed4fNtD6_0),.din(w_dff_A_mZEO4lcH5_0),.clk(gclk));
	jdff dff_A_Qed4fNtD6_0(.dout(w_dff_A_dnkFVgsd9_0),.din(w_dff_A_Qed4fNtD6_0),.clk(gclk));
	jdff dff_A_dnkFVgsd9_0(.dout(w_dff_A_GzdROERb7_0),.din(w_dff_A_dnkFVgsd9_0),.clk(gclk));
	jdff dff_A_GzdROERb7_0(.dout(w_dff_A_H6pVIzM71_0),.din(w_dff_A_GzdROERb7_0),.clk(gclk));
	jdff dff_A_H6pVIzM71_0(.dout(w_dff_A_fWCT3Tbj0_0),.din(w_dff_A_H6pVIzM71_0),.clk(gclk));
	jdff dff_A_fWCT3Tbj0_0(.dout(w_dff_A_LJittrPQ2_0),.din(w_dff_A_fWCT3Tbj0_0),.clk(gclk));
	jdff dff_A_LJittrPQ2_0(.dout(w_dff_A_O1Ysbbvb8_0),.din(w_dff_A_LJittrPQ2_0),.clk(gclk));
	jdff dff_A_O1Ysbbvb8_0(.dout(w_dff_A_wIAaI4lj1_0),.din(w_dff_A_O1Ysbbvb8_0),.clk(gclk));
	jdff dff_A_wIAaI4lj1_0(.dout(w_dff_A_3AA3RUl77_0),.din(w_dff_A_wIAaI4lj1_0),.clk(gclk));
	jdff dff_A_3AA3RUl77_0(.dout(w_dff_A_epUiVVul2_0),.din(w_dff_A_3AA3RUl77_0),.clk(gclk));
	jdff dff_A_epUiVVul2_0(.dout(w_dff_A_SgiBcpn85_0),.din(w_dff_A_epUiVVul2_0),.clk(gclk));
	jdff dff_A_SgiBcpn85_0(.dout(w_dff_A_lFX3JfSB8_0),.din(w_dff_A_SgiBcpn85_0),.clk(gclk));
	jdff dff_A_lFX3JfSB8_0(.dout(w_dff_A_jsyb64pj3_0),.din(w_dff_A_lFX3JfSB8_0),.clk(gclk));
	jdff dff_A_jsyb64pj3_0(.dout(w_dff_A_jstxn0x46_0),.din(w_dff_A_jsyb64pj3_0),.clk(gclk));
	jdff dff_A_jstxn0x46_0(.dout(w_dff_A_g63k50sU5_0),.din(w_dff_A_jstxn0x46_0),.clk(gclk));
	jdff dff_A_g63k50sU5_0(.dout(w_dff_A_ugv7Mo1N1_0),.din(w_dff_A_g63k50sU5_0),.clk(gclk));
	jdff dff_A_ugv7Mo1N1_0(.dout(w_dff_A_1rfbSUbt9_0),.din(w_dff_A_ugv7Mo1N1_0),.clk(gclk));
	jdff dff_A_1rfbSUbt9_0(.dout(w_dff_A_Kyr4O1qO0_0),.din(w_dff_A_1rfbSUbt9_0),.clk(gclk));
	jdff dff_A_Kyr4O1qO0_0(.dout(w_dff_A_yUdAOVuT6_0),.din(w_dff_A_Kyr4O1qO0_0),.clk(gclk));
	jdff dff_A_yUdAOVuT6_0(.dout(G1004),.din(w_dff_A_yUdAOVuT6_0),.clk(gclk));
	jdff dff_A_wVLt2fwl5_2(.dout(w_dff_A_PZCHGf947_0),.din(w_dff_A_wVLt2fwl5_2),.clk(gclk));
	jdff dff_A_PZCHGf947_0(.dout(w_dff_A_NJ11g6qr5_0),.din(w_dff_A_PZCHGf947_0),.clk(gclk));
	jdff dff_A_NJ11g6qr5_0(.dout(w_dff_A_mWohJyYd5_0),.din(w_dff_A_NJ11g6qr5_0),.clk(gclk));
	jdff dff_A_mWohJyYd5_0(.dout(w_dff_A_EEbexcJG9_0),.din(w_dff_A_mWohJyYd5_0),.clk(gclk));
	jdff dff_A_EEbexcJG9_0(.dout(w_dff_A_7Wvr3adD9_0),.din(w_dff_A_EEbexcJG9_0),.clk(gclk));
	jdff dff_A_7Wvr3adD9_0(.dout(w_dff_A_AnjeX9W55_0),.din(w_dff_A_7Wvr3adD9_0),.clk(gclk));
	jdff dff_A_AnjeX9W55_0(.dout(w_dff_A_JeVX2hpH3_0),.din(w_dff_A_AnjeX9W55_0),.clk(gclk));
	jdff dff_A_JeVX2hpH3_0(.dout(w_dff_A_mQ3pGYN86_0),.din(w_dff_A_JeVX2hpH3_0),.clk(gclk));
	jdff dff_A_mQ3pGYN86_0(.dout(w_dff_A_XYf36Z6f4_0),.din(w_dff_A_mQ3pGYN86_0),.clk(gclk));
	jdff dff_A_XYf36Z6f4_0(.dout(w_dff_A_DzdQewHO0_0),.din(w_dff_A_XYf36Z6f4_0),.clk(gclk));
	jdff dff_A_DzdQewHO0_0(.dout(w_dff_A_RujkW4kl1_0),.din(w_dff_A_DzdQewHO0_0),.clk(gclk));
	jdff dff_A_RujkW4kl1_0(.dout(w_dff_A_6PA3kwT35_0),.din(w_dff_A_RujkW4kl1_0),.clk(gclk));
	jdff dff_A_6PA3kwT35_0(.dout(w_dff_A_zdVWXy3r7_0),.din(w_dff_A_6PA3kwT35_0),.clk(gclk));
	jdff dff_A_zdVWXy3r7_0(.dout(G591),.din(w_dff_A_zdVWXy3r7_0),.clk(gclk));
	jdff dff_A_MzAOxEXW9_2(.dout(w_dff_A_9X3Pn8eE2_0),.din(w_dff_A_MzAOxEXW9_2),.clk(gclk));
	jdff dff_A_9X3Pn8eE2_0(.dout(w_dff_A_qawLeH7P7_0),.din(w_dff_A_9X3Pn8eE2_0),.clk(gclk));
	jdff dff_A_qawLeH7P7_0(.dout(w_dff_A_9Rfmas5U0_0),.din(w_dff_A_qawLeH7P7_0),.clk(gclk));
	jdff dff_A_9Rfmas5U0_0(.dout(w_dff_A_jEfDCNv94_0),.din(w_dff_A_9Rfmas5U0_0),.clk(gclk));
	jdff dff_A_jEfDCNv94_0(.dout(w_dff_A_zk8pjiVS4_0),.din(w_dff_A_jEfDCNv94_0),.clk(gclk));
	jdff dff_A_zk8pjiVS4_0(.dout(w_dff_A_OXsUkfJn6_0),.din(w_dff_A_zk8pjiVS4_0),.clk(gclk));
	jdff dff_A_OXsUkfJn6_0(.dout(w_dff_A_k4j8aSAO1_0),.din(w_dff_A_OXsUkfJn6_0),.clk(gclk));
	jdff dff_A_k4j8aSAO1_0(.dout(w_dff_A_ALiYrbV64_0),.din(w_dff_A_k4j8aSAO1_0),.clk(gclk));
	jdff dff_A_ALiYrbV64_0(.dout(w_dff_A_hAvwYYuR6_0),.din(w_dff_A_ALiYrbV64_0),.clk(gclk));
	jdff dff_A_hAvwYYuR6_0(.dout(w_dff_A_Ma8vgY6H1_0),.din(w_dff_A_hAvwYYuR6_0),.clk(gclk));
	jdff dff_A_Ma8vgY6H1_0(.dout(w_dff_A_hY6M1ezZ6_0),.din(w_dff_A_Ma8vgY6H1_0),.clk(gclk));
	jdff dff_A_hY6M1ezZ6_0(.dout(w_dff_A_B1Joi4kL7_0),.din(w_dff_A_hY6M1ezZ6_0),.clk(gclk));
	jdff dff_A_B1Joi4kL7_0(.dout(w_dff_A_tN8T7bLt9_0),.din(w_dff_A_B1Joi4kL7_0),.clk(gclk));
	jdff dff_A_tN8T7bLt9_0(.dout(w_dff_A_N8vkVn4P5_0),.din(w_dff_A_tN8T7bLt9_0),.clk(gclk));
	jdff dff_A_N8vkVn4P5_0(.dout(G618),.din(w_dff_A_N8vkVn4P5_0),.clk(gclk));
	jdff dff_A_J8PJIiZa7_2(.dout(w_dff_A_UMXLmLoQ3_0),.din(w_dff_A_J8PJIiZa7_2),.clk(gclk));
	jdff dff_A_UMXLmLoQ3_0(.dout(w_dff_A_IwFPbbez8_0),.din(w_dff_A_UMXLmLoQ3_0),.clk(gclk));
	jdff dff_A_IwFPbbez8_0(.dout(w_dff_A_1NNzDRzd3_0),.din(w_dff_A_IwFPbbez8_0),.clk(gclk));
	jdff dff_A_1NNzDRzd3_0(.dout(w_dff_A_LeKReWjO6_0),.din(w_dff_A_1NNzDRzd3_0),.clk(gclk));
	jdff dff_A_LeKReWjO6_0(.dout(w_dff_A_l9rsI4ey3_0),.din(w_dff_A_LeKReWjO6_0),.clk(gclk));
	jdff dff_A_l9rsI4ey3_0(.dout(w_dff_A_cndWKWAL7_0),.din(w_dff_A_l9rsI4ey3_0),.clk(gclk));
	jdff dff_A_cndWKWAL7_0(.dout(w_dff_A_Vmg6RrNA6_0),.din(w_dff_A_cndWKWAL7_0),.clk(gclk));
	jdff dff_A_Vmg6RrNA6_0(.dout(w_dff_A_eLXdqB9e3_0),.din(w_dff_A_Vmg6RrNA6_0),.clk(gclk));
	jdff dff_A_eLXdqB9e3_0(.dout(w_dff_A_3mfnXiYl9_0),.din(w_dff_A_eLXdqB9e3_0),.clk(gclk));
	jdff dff_A_3mfnXiYl9_0(.dout(w_dff_A_LGKsPkIc3_0),.din(w_dff_A_3mfnXiYl9_0),.clk(gclk));
	jdff dff_A_LGKsPkIc3_0(.dout(w_dff_A_DdYiOf791_0),.din(w_dff_A_LGKsPkIc3_0),.clk(gclk));
	jdff dff_A_DdYiOf791_0(.dout(w_dff_A_ZRvPIl9d4_0),.din(w_dff_A_DdYiOf791_0),.clk(gclk));
	jdff dff_A_ZRvPIl9d4_0(.dout(w_dff_A_ApMhF7as7_0),.din(w_dff_A_ZRvPIl9d4_0),.clk(gclk));
	jdff dff_A_ApMhF7as7_0(.dout(G621),.din(w_dff_A_ApMhF7as7_0),.clk(gclk));
	jdff dff_A_hRVgxDpe1_2(.dout(w_dff_A_3BKxgBZc2_0),.din(w_dff_A_hRVgxDpe1_2),.clk(gclk));
	jdff dff_A_3BKxgBZc2_0(.dout(w_dff_A_W9FL22ak9_0),.din(w_dff_A_3BKxgBZc2_0),.clk(gclk));
	jdff dff_A_W9FL22ak9_0(.dout(w_dff_A_5VJjdRjV6_0),.din(w_dff_A_W9FL22ak9_0),.clk(gclk));
	jdff dff_A_5VJjdRjV6_0(.dout(w_dff_A_UwkYKMji2_0),.din(w_dff_A_5VJjdRjV6_0),.clk(gclk));
	jdff dff_A_UwkYKMji2_0(.dout(w_dff_A_ovQ3zXr26_0),.din(w_dff_A_UwkYKMji2_0),.clk(gclk));
	jdff dff_A_ovQ3zXr26_0(.dout(w_dff_A_1T0kapjh0_0),.din(w_dff_A_ovQ3zXr26_0),.clk(gclk));
	jdff dff_A_1T0kapjh0_0(.dout(w_dff_A_ajMJw7G86_0),.din(w_dff_A_1T0kapjh0_0),.clk(gclk));
	jdff dff_A_ajMJw7G86_0(.dout(w_dff_A_NGFkhBio2_0),.din(w_dff_A_ajMJw7G86_0),.clk(gclk));
	jdff dff_A_NGFkhBio2_0(.dout(w_dff_A_ONl7d8SL5_0),.din(w_dff_A_NGFkhBio2_0),.clk(gclk));
	jdff dff_A_ONl7d8SL5_0(.dout(w_dff_A_11F9Sisx4_0),.din(w_dff_A_ONl7d8SL5_0),.clk(gclk));
	jdff dff_A_11F9Sisx4_0(.dout(w_dff_A_dTEu4vA70_0),.din(w_dff_A_11F9Sisx4_0),.clk(gclk));
	jdff dff_A_dTEu4vA70_0(.dout(w_dff_A_54hU4fjU8_0),.din(w_dff_A_dTEu4vA70_0),.clk(gclk));
	jdff dff_A_54hU4fjU8_0(.dout(w_dff_A_1kwP5e1J8_0),.din(w_dff_A_54hU4fjU8_0),.clk(gclk));
	jdff dff_A_1kwP5e1J8_0(.dout(w_dff_A_CGf1GCyk1_0),.din(w_dff_A_1kwP5e1J8_0),.clk(gclk));
	jdff dff_A_CGf1GCyk1_0(.dout(G629),.din(w_dff_A_CGf1GCyk1_0),.clk(gclk));
	jdff dff_A_SdU8Ychv1_1(.dout(w_dff_A_b59BOzON2_0),.din(w_dff_A_SdU8Ychv1_1),.clk(gclk));
	jdff dff_A_b59BOzON2_0(.dout(w_dff_A_5evS7cM61_0),.din(w_dff_A_b59BOzON2_0),.clk(gclk));
	jdff dff_A_5evS7cM61_0(.dout(w_dff_A_VQsZAgLQ5_0),.din(w_dff_A_5evS7cM61_0),.clk(gclk));
	jdff dff_A_VQsZAgLQ5_0(.dout(w_dff_A_fvgTNHTg3_0),.din(w_dff_A_VQsZAgLQ5_0),.clk(gclk));
	jdff dff_A_fvgTNHTg3_0(.dout(w_dff_A_LmxUshWR6_0),.din(w_dff_A_fvgTNHTg3_0),.clk(gclk));
	jdff dff_A_LmxUshWR6_0(.dout(w_dff_A_YLOO6T3Q7_0),.din(w_dff_A_LmxUshWR6_0),.clk(gclk));
	jdff dff_A_YLOO6T3Q7_0(.dout(w_dff_A_FiQgZcED1_0),.din(w_dff_A_YLOO6T3Q7_0),.clk(gclk));
	jdff dff_A_FiQgZcED1_0(.dout(w_dff_A_TPFL85ES4_0),.din(w_dff_A_FiQgZcED1_0),.clk(gclk));
	jdff dff_A_TPFL85ES4_0(.dout(w_dff_A_VOrjK6ku2_0),.din(w_dff_A_TPFL85ES4_0),.clk(gclk));
	jdff dff_A_VOrjK6ku2_0(.dout(w_dff_A_8MPjGdTR8_0),.din(w_dff_A_VOrjK6ku2_0),.clk(gclk));
	jdff dff_A_8MPjGdTR8_0(.dout(w_dff_A_sit0Az727_0),.din(w_dff_A_8MPjGdTR8_0),.clk(gclk));
	jdff dff_A_sit0Az727_0(.dout(w_dff_A_adQgxcG27_0),.din(w_dff_A_sit0Az727_0),.clk(gclk));
	jdff dff_A_adQgxcG27_0(.dout(w_dff_A_LCRA9Brj1_0),.din(w_dff_A_adQgxcG27_0),.clk(gclk));
	jdff dff_A_LCRA9Brj1_0(.dout(w_dff_A_T8BgQUx47_0),.din(w_dff_A_LCRA9Brj1_0),.clk(gclk));
	jdff dff_A_T8BgQUx47_0(.dout(w_dff_A_UBPzdATJ5_0),.din(w_dff_A_T8BgQUx47_0),.clk(gclk));
	jdff dff_A_UBPzdATJ5_0(.dout(w_dff_A_Z0mK3ixY2_0),.din(w_dff_A_UBPzdATJ5_0),.clk(gclk));
	jdff dff_A_Z0mK3ixY2_0(.dout(w_dff_A_5IVW2f2u0_0),.din(w_dff_A_Z0mK3ixY2_0),.clk(gclk));
	jdff dff_A_5IVW2f2u0_0(.dout(w_dff_A_j99qilMN7_0),.din(w_dff_A_5IVW2f2u0_0),.clk(gclk));
	jdff dff_A_j99qilMN7_0(.dout(w_dff_A_DUizNmRJ3_0),.din(w_dff_A_j99qilMN7_0),.clk(gclk));
	jdff dff_A_DUizNmRJ3_0(.dout(G822),.din(w_dff_A_DUizNmRJ3_0),.clk(gclk));
	jdff dff_A_a58wHPnb2_1(.dout(w_dff_A_wYn9j1Et6_0),.din(w_dff_A_a58wHPnb2_1),.clk(gclk));
	jdff dff_A_wYn9j1Et6_0(.dout(w_dff_A_yI9ZSApH4_0),.din(w_dff_A_wYn9j1Et6_0),.clk(gclk));
	jdff dff_A_yI9ZSApH4_0(.dout(w_dff_A_lPSCcV8t7_0),.din(w_dff_A_yI9ZSApH4_0),.clk(gclk));
	jdff dff_A_lPSCcV8t7_0(.dout(w_dff_A_hDKu8tTO6_0),.din(w_dff_A_lPSCcV8t7_0),.clk(gclk));
	jdff dff_A_hDKu8tTO6_0(.dout(w_dff_A_TbUr0Iry2_0),.din(w_dff_A_hDKu8tTO6_0),.clk(gclk));
	jdff dff_A_TbUr0Iry2_0(.dout(w_dff_A_HCRNcGUn5_0),.din(w_dff_A_TbUr0Iry2_0),.clk(gclk));
	jdff dff_A_HCRNcGUn5_0(.dout(w_dff_A_S4LhQc787_0),.din(w_dff_A_HCRNcGUn5_0),.clk(gclk));
	jdff dff_A_S4LhQc787_0(.dout(w_dff_A_NTat5lOP9_0),.din(w_dff_A_S4LhQc787_0),.clk(gclk));
	jdff dff_A_NTat5lOP9_0(.dout(w_dff_A_EaIYQwfe6_0),.din(w_dff_A_NTat5lOP9_0),.clk(gclk));
	jdff dff_A_EaIYQwfe6_0(.dout(w_dff_A_tYebnlEB2_0),.din(w_dff_A_EaIYQwfe6_0),.clk(gclk));
	jdff dff_A_tYebnlEB2_0(.dout(w_dff_A_WGg9h5RS3_0),.din(w_dff_A_tYebnlEB2_0),.clk(gclk));
	jdff dff_A_WGg9h5RS3_0(.dout(w_dff_A_3wl6G3dr5_0),.din(w_dff_A_WGg9h5RS3_0),.clk(gclk));
	jdff dff_A_3wl6G3dr5_0(.dout(w_dff_A_EckDMSF67_0),.din(w_dff_A_3wl6G3dr5_0),.clk(gclk));
	jdff dff_A_EckDMSF67_0(.dout(w_dff_A_MQf5LBrF0_0),.din(w_dff_A_EckDMSF67_0),.clk(gclk));
	jdff dff_A_MQf5LBrF0_0(.dout(G838),.din(w_dff_A_MQf5LBrF0_0),.clk(gclk));
	jdff dff_A_32PGN2ft4_1(.dout(w_dff_A_0NT0t0jJ8_0),.din(w_dff_A_32PGN2ft4_1),.clk(gclk));
	jdff dff_A_0NT0t0jJ8_0(.dout(w_dff_A_WlYMB3uz7_0),.din(w_dff_A_0NT0t0jJ8_0),.clk(gclk));
	jdff dff_A_WlYMB3uz7_0(.dout(w_dff_A_lAlYggaD6_0),.din(w_dff_A_WlYMB3uz7_0),.clk(gclk));
	jdff dff_A_lAlYggaD6_0(.dout(w_dff_A_WclX20pc4_0),.din(w_dff_A_lAlYggaD6_0),.clk(gclk));
	jdff dff_A_WclX20pc4_0(.dout(w_dff_A_6AHVoOgq9_0),.din(w_dff_A_WclX20pc4_0),.clk(gclk));
	jdff dff_A_6AHVoOgq9_0(.dout(w_dff_A_gD65qEXj8_0),.din(w_dff_A_6AHVoOgq9_0),.clk(gclk));
	jdff dff_A_gD65qEXj8_0(.dout(w_dff_A_Te0haAZQ7_0),.din(w_dff_A_gD65qEXj8_0),.clk(gclk));
	jdff dff_A_Te0haAZQ7_0(.dout(w_dff_A_x76ZPAeB7_0),.din(w_dff_A_Te0haAZQ7_0),.clk(gclk));
	jdff dff_A_x76ZPAeB7_0(.dout(w_dff_A_gLnDJxeA3_0),.din(w_dff_A_x76ZPAeB7_0),.clk(gclk));
	jdff dff_A_gLnDJxeA3_0(.dout(w_dff_A_469XsOUb1_0),.din(w_dff_A_gLnDJxeA3_0),.clk(gclk));
	jdff dff_A_469XsOUb1_0(.dout(w_dff_A_XgfTY49g7_0),.din(w_dff_A_469XsOUb1_0),.clk(gclk));
	jdff dff_A_XgfTY49g7_0(.dout(w_dff_A_BWypaNZQ2_0),.din(w_dff_A_XgfTY49g7_0),.clk(gclk));
	jdff dff_A_BWypaNZQ2_0(.dout(w_dff_A_pSruikRH1_0),.din(w_dff_A_BWypaNZQ2_0),.clk(gclk));
	jdff dff_A_pSruikRH1_0(.dout(w_dff_A_nYalfgC52_0),.din(w_dff_A_pSruikRH1_0),.clk(gclk));
	jdff dff_A_nYalfgC52_0(.dout(w_dff_A_hVbPYwVF4_0),.din(w_dff_A_nYalfgC52_0),.clk(gclk));
	jdff dff_A_hVbPYwVF4_0(.dout(w_dff_A_ePx9x8A67_0),.din(w_dff_A_hVbPYwVF4_0),.clk(gclk));
	jdff dff_A_ePx9x8A67_0(.dout(w_dff_A_kyW7fDwR3_0),.din(w_dff_A_ePx9x8A67_0),.clk(gclk));
	jdff dff_A_kyW7fDwR3_0(.dout(G861),.din(w_dff_A_kyW7fDwR3_0),.clk(gclk));
	jdff dff_A_3zZlppPo2_1(.dout(w_dff_A_8weYVMmf7_0),.din(w_dff_A_3zZlppPo2_1),.clk(gclk));
	jdff dff_A_8weYVMmf7_0(.dout(w_dff_A_46xYHbYS7_0),.din(w_dff_A_8weYVMmf7_0),.clk(gclk));
	jdff dff_A_46xYHbYS7_0(.dout(w_dff_A_O8QUlp923_0),.din(w_dff_A_46xYHbYS7_0),.clk(gclk));
	jdff dff_A_O8QUlp923_0(.dout(w_dff_A_qHVTEQ9X1_0),.din(w_dff_A_O8QUlp923_0),.clk(gclk));
	jdff dff_A_qHVTEQ9X1_0(.dout(w_dff_A_LIMCHDzK6_0),.din(w_dff_A_qHVTEQ9X1_0),.clk(gclk));
	jdff dff_A_LIMCHDzK6_0(.dout(w_dff_A_5Tc8NSCd0_0),.din(w_dff_A_LIMCHDzK6_0),.clk(gclk));
	jdff dff_A_5Tc8NSCd0_0(.dout(w_dff_A_fZyzX2971_0),.din(w_dff_A_5Tc8NSCd0_0),.clk(gclk));
	jdff dff_A_fZyzX2971_0(.dout(w_dff_A_BjgDiEph7_0),.din(w_dff_A_fZyzX2971_0),.clk(gclk));
	jdff dff_A_BjgDiEph7_0(.dout(w_dff_A_8ZxZ9coM0_0),.din(w_dff_A_BjgDiEph7_0),.clk(gclk));
	jdff dff_A_8ZxZ9coM0_0(.dout(G623),.din(w_dff_A_8ZxZ9coM0_0),.clk(gclk));
	jdff dff_A_GoqX3tdp4_2(.dout(w_dff_A_I9xItxkS9_0),.din(w_dff_A_GoqX3tdp4_2),.clk(gclk));
	jdff dff_A_I9xItxkS9_0(.dout(w_dff_A_uq9sOmXv4_0),.din(w_dff_A_I9xItxkS9_0),.clk(gclk));
	jdff dff_A_uq9sOmXv4_0(.dout(w_dff_A_tNUsV5H25_0),.din(w_dff_A_uq9sOmXv4_0),.clk(gclk));
	jdff dff_A_tNUsV5H25_0(.dout(w_dff_A_Z3uo7zSo0_0),.din(w_dff_A_tNUsV5H25_0),.clk(gclk));
	jdff dff_A_Z3uo7zSo0_0(.dout(w_dff_A_nrJ2TCgw8_0),.din(w_dff_A_Z3uo7zSo0_0),.clk(gclk));
	jdff dff_A_nrJ2TCgw8_0(.dout(w_dff_A_ct8DkuX10_0),.din(w_dff_A_nrJ2TCgw8_0),.clk(gclk));
	jdff dff_A_ct8DkuX10_0(.dout(w_dff_A_uiLP1dwA9_0),.din(w_dff_A_ct8DkuX10_0),.clk(gclk));
	jdff dff_A_uiLP1dwA9_0(.dout(w_dff_A_ntBSl8Xl6_0),.din(w_dff_A_uiLP1dwA9_0),.clk(gclk));
	jdff dff_A_ntBSl8Xl6_0(.dout(w_dff_A_HabsYJWC9_0),.din(w_dff_A_ntBSl8Xl6_0),.clk(gclk));
	jdff dff_A_HabsYJWC9_0(.dout(w_dff_A_4kUgOLuD8_0),.din(w_dff_A_HabsYJWC9_0),.clk(gclk));
	jdff dff_A_4kUgOLuD8_0(.dout(w_dff_A_QtoxRyzn3_0),.din(w_dff_A_4kUgOLuD8_0),.clk(gclk));
	jdff dff_A_QtoxRyzn3_0(.dout(w_dff_A_2RuDNGB85_0),.din(w_dff_A_QtoxRyzn3_0),.clk(gclk));
	jdff dff_A_2RuDNGB85_0(.dout(w_dff_A_cSpm6UOC1_0),.din(w_dff_A_2RuDNGB85_0),.clk(gclk));
	jdff dff_A_cSpm6UOC1_0(.dout(G722),.din(w_dff_A_cSpm6UOC1_0),.clk(gclk));
	jdff dff_A_J4Jmmsg98_1(.dout(w_dff_A_fu8N7Iyj5_0),.din(w_dff_A_J4Jmmsg98_1),.clk(gclk));
	jdff dff_A_fu8N7Iyj5_0(.dout(w_dff_A_q07gtgke8_0),.din(w_dff_A_fu8N7Iyj5_0),.clk(gclk));
	jdff dff_A_q07gtgke8_0(.dout(w_dff_A_VMTIhTb74_0),.din(w_dff_A_q07gtgke8_0),.clk(gclk));
	jdff dff_A_VMTIhTb74_0(.dout(w_dff_A_yxirF8vl7_0),.din(w_dff_A_VMTIhTb74_0),.clk(gclk));
	jdff dff_A_yxirF8vl7_0(.dout(w_dff_A_7IkhlJY36_0),.din(w_dff_A_yxirF8vl7_0),.clk(gclk));
	jdff dff_A_7IkhlJY36_0(.dout(w_dff_A_i5pzBwBT1_0),.din(w_dff_A_7IkhlJY36_0),.clk(gclk));
	jdff dff_A_i5pzBwBT1_0(.dout(w_dff_A_K4J5kSOj3_0),.din(w_dff_A_i5pzBwBT1_0),.clk(gclk));
	jdff dff_A_K4J5kSOj3_0(.dout(w_dff_A_MEOPsBff9_0),.din(w_dff_A_K4J5kSOj3_0),.clk(gclk));
	jdff dff_A_MEOPsBff9_0(.dout(w_dff_A_eYIqAtBs3_0),.din(w_dff_A_MEOPsBff9_0),.clk(gclk));
	jdff dff_A_eYIqAtBs3_0(.dout(w_dff_A_SpvSlMBR6_0),.din(w_dff_A_eYIqAtBs3_0),.clk(gclk));
	jdff dff_A_SpvSlMBR6_0(.dout(w_dff_A_YM9XQKYJ3_0),.din(w_dff_A_SpvSlMBR6_0),.clk(gclk));
	jdff dff_A_YM9XQKYJ3_0(.dout(w_dff_A_85IV5hjF4_0),.din(w_dff_A_YM9XQKYJ3_0),.clk(gclk));
	jdff dff_A_85IV5hjF4_0(.dout(G832),.din(w_dff_A_85IV5hjF4_0),.clk(gclk));
	jdff dff_A_BZPX3kBd6_1(.dout(w_dff_A_MItrpGh65_0),.din(w_dff_A_BZPX3kBd6_1),.clk(gclk));
	jdff dff_A_MItrpGh65_0(.dout(w_dff_A_IUypSK960_0),.din(w_dff_A_MItrpGh65_0),.clk(gclk));
	jdff dff_A_IUypSK960_0(.dout(w_dff_A_XzVI3ZSR3_0),.din(w_dff_A_IUypSK960_0),.clk(gclk));
	jdff dff_A_XzVI3ZSR3_0(.dout(w_dff_A_f9L7DiAN9_0),.din(w_dff_A_XzVI3ZSR3_0),.clk(gclk));
	jdff dff_A_f9L7DiAN9_0(.dout(w_dff_A_a2K44Dff4_0),.din(w_dff_A_f9L7DiAN9_0),.clk(gclk));
	jdff dff_A_a2K44Dff4_0(.dout(w_dff_A_Y41Fkdox8_0),.din(w_dff_A_a2K44Dff4_0),.clk(gclk));
	jdff dff_A_Y41Fkdox8_0(.dout(w_dff_A_SPgIzt2E7_0),.din(w_dff_A_Y41Fkdox8_0),.clk(gclk));
	jdff dff_A_SPgIzt2E7_0(.dout(w_dff_A_9ssSqLAV8_0),.din(w_dff_A_SPgIzt2E7_0),.clk(gclk));
	jdff dff_A_9ssSqLAV8_0(.dout(w_dff_A_CXWCqIcV7_0),.din(w_dff_A_9ssSqLAV8_0),.clk(gclk));
	jdff dff_A_CXWCqIcV7_0(.dout(w_dff_A_srJsI7k85_0),.din(w_dff_A_CXWCqIcV7_0),.clk(gclk));
	jdff dff_A_srJsI7k85_0(.dout(w_dff_A_ADpst9c51_0),.din(w_dff_A_srJsI7k85_0),.clk(gclk));
	jdff dff_A_ADpst9c51_0(.dout(w_dff_A_rrDLn1se8_0),.din(w_dff_A_ADpst9c51_0),.clk(gclk));
	jdff dff_A_rrDLn1se8_0(.dout(w_dff_A_hLae4ReT4_0),.din(w_dff_A_rrDLn1se8_0),.clk(gclk));
	jdff dff_A_hLae4ReT4_0(.dout(G834),.din(w_dff_A_hLae4ReT4_0),.clk(gclk));
	jdff dff_A_YrJpRzMx9_1(.dout(w_dff_A_vPTUWUZ44_0),.din(w_dff_A_YrJpRzMx9_1),.clk(gclk));
	jdff dff_A_vPTUWUZ44_0(.dout(w_dff_A_4mbCgx3w6_0),.din(w_dff_A_vPTUWUZ44_0),.clk(gclk));
	jdff dff_A_4mbCgx3w6_0(.dout(w_dff_A_k7kLNezn5_0),.din(w_dff_A_4mbCgx3w6_0),.clk(gclk));
	jdff dff_A_k7kLNezn5_0(.dout(w_dff_A_sSAHpwEj7_0),.din(w_dff_A_k7kLNezn5_0),.clk(gclk));
	jdff dff_A_sSAHpwEj7_0(.dout(w_dff_A_JQ7IdnRW4_0),.din(w_dff_A_sSAHpwEj7_0),.clk(gclk));
	jdff dff_A_JQ7IdnRW4_0(.dout(w_dff_A_k9QeNSBi3_0),.din(w_dff_A_JQ7IdnRW4_0),.clk(gclk));
	jdff dff_A_k9QeNSBi3_0(.dout(w_dff_A_V72f7WbK2_0),.din(w_dff_A_k9QeNSBi3_0),.clk(gclk));
	jdff dff_A_V72f7WbK2_0(.dout(w_dff_A_8SZzEg7y1_0),.din(w_dff_A_V72f7WbK2_0),.clk(gclk));
	jdff dff_A_8SZzEg7y1_0(.dout(w_dff_A_ro2KrKeu3_0),.din(w_dff_A_8SZzEg7y1_0),.clk(gclk));
	jdff dff_A_ro2KrKeu3_0(.dout(w_dff_A_oIZkV3059_0),.din(w_dff_A_ro2KrKeu3_0),.clk(gclk));
	jdff dff_A_oIZkV3059_0(.dout(w_dff_A_Rr0bFvnv3_0),.din(w_dff_A_oIZkV3059_0),.clk(gclk));
	jdff dff_A_Rr0bFvnv3_0(.dout(w_dff_A_JwJNc1rY2_0),.din(w_dff_A_Rr0bFvnv3_0),.clk(gclk));
	jdff dff_A_JwJNc1rY2_0(.dout(w_dff_A_oEGW1y4M4_0),.din(w_dff_A_JwJNc1rY2_0),.clk(gclk));
	jdff dff_A_oEGW1y4M4_0(.dout(w_dff_A_jrRy5ZX90_0),.din(w_dff_A_oEGW1y4M4_0),.clk(gclk));
	jdff dff_A_jrRy5ZX90_0(.dout(w_dff_A_KAN7zrM39_0),.din(w_dff_A_jrRy5ZX90_0),.clk(gclk));
	jdff dff_A_KAN7zrM39_0(.dout(G836),.din(w_dff_A_KAN7zrM39_0),.clk(gclk));
	jdff dff_A_P2qeWm9N7_2(.dout(w_dff_A_cqLYJVgY1_0),.din(w_dff_A_P2qeWm9N7_2),.clk(gclk));
	jdff dff_A_cqLYJVgY1_0(.dout(w_dff_A_aNPxrL0N8_0),.din(w_dff_A_cqLYJVgY1_0),.clk(gclk));
	jdff dff_A_aNPxrL0N8_0(.dout(w_dff_A_JheEaVT01_0),.din(w_dff_A_aNPxrL0N8_0),.clk(gclk));
	jdff dff_A_JheEaVT01_0(.dout(w_dff_A_zC9WtCeW4_0),.din(w_dff_A_JheEaVT01_0),.clk(gclk));
	jdff dff_A_zC9WtCeW4_0(.dout(w_dff_A_zr3zYmsV5_0),.din(w_dff_A_zC9WtCeW4_0),.clk(gclk));
	jdff dff_A_zr3zYmsV5_0(.dout(w_dff_A_csHtLnaH5_0),.din(w_dff_A_zr3zYmsV5_0),.clk(gclk));
	jdff dff_A_csHtLnaH5_0(.dout(w_dff_A_GLz5aASv1_0),.din(w_dff_A_csHtLnaH5_0),.clk(gclk));
	jdff dff_A_GLz5aASv1_0(.dout(w_dff_A_wxejWMT14_0),.din(w_dff_A_GLz5aASv1_0),.clk(gclk));
	jdff dff_A_wxejWMT14_0(.dout(w_dff_A_lnS1CrEj9_0),.din(w_dff_A_wxejWMT14_0),.clk(gclk));
	jdff dff_A_lnS1CrEj9_0(.dout(w_dff_A_slRbJA7W9_0),.din(w_dff_A_lnS1CrEj9_0),.clk(gclk));
	jdff dff_A_slRbJA7W9_0(.dout(w_dff_A_71s5LhIN8_0),.din(w_dff_A_slRbJA7W9_0),.clk(gclk));
	jdff dff_A_71s5LhIN8_0(.dout(w_dff_A_HatCxxBI5_0),.din(w_dff_A_71s5LhIN8_0),.clk(gclk));
	jdff dff_A_HatCxxBI5_0(.dout(w_dff_A_AKunThgh7_0),.din(w_dff_A_HatCxxBI5_0),.clk(gclk));
	jdff dff_A_AKunThgh7_0(.dout(G859),.din(w_dff_A_AKunThgh7_0),.clk(gclk));
	jdff dff_A_mblDQHA37_1(.dout(w_dff_A_HJr4ozNT9_0),.din(w_dff_A_mblDQHA37_1),.clk(gclk));
	jdff dff_A_HJr4ozNT9_0(.dout(w_dff_A_t4aSr7M02_0),.din(w_dff_A_HJr4ozNT9_0),.clk(gclk));
	jdff dff_A_t4aSr7M02_0(.dout(w_dff_A_Lzm1nq0E4_0),.din(w_dff_A_t4aSr7M02_0),.clk(gclk));
	jdff dff_A_Lzm1nq0E4_0(.dout(w_dff_A_qo1EGmtQ5_0),.din(w_dff_A_Lzm1nq0E4_0),.clk(gclk));
	jdff dff_A_qo1EGmtQ5_0(.dout(w_dff_A_dBBSXc9N2_0),.din(w_dff_A_qo1EGmtQ5_0),.clk(gclk));
	jdff dff_A_dBBSXc9N2_0(.dout(w_dff_A_Npxmb5Lo1_0),.din(w_dff_A_dBBSXc9N2_0),.clk(gclk));
	jdff dff_A_Npxmb5Lo1_0(.dout(w_dff_A_8xbCYDrK9_0),.din(w_dff_A_Npxmb5Lo1_0),.clk(gclk));
	jdff dff_A_8xbCYDrK9_0(.dout(w_dff_A_V0v7UeVO0_0),.din(w_dff_A_8xbCYDrK9_0),.clk(gclk));
	jdff dff_A_V0v7UeVO0_0(.dout(w_dff_A_sl4C8Jhf8_0),.din(w_dff_A_V0v7UeVO0_0),.clk(gclk));
	jdff dff_A_sl4C8Jhf8_0(.dout(w_dff_A_NMcB3cU60_0),.din(w_dff_A_sl4C8Jhf8_0),.clk(gclk));
	jdff dff_A_NMcB3cU60_0(.dout(w_dff_A_BrjD1oyV2_0),.din(w_dff_A_NMcB3cU60_0),.clk(gclk));
	jdff dff_A_BrjD1oyV2_0(.dout(w_dff_A_woudQSwI3_0),.din(w_dff_A_BrjD1oyV2_0),.clk(gclk));
	jdff dff_A_woudQSwI3_0(.dout(G871),.din(w_dff_A_woudQSwI3_0),.clk(gclk));
	jdff dff_A_xLUN1R8u8_1(.dout(w_dff_A_1pgpu9CU4_0),.din(w_dff_A_xLUN1R8u8_1),.clk(gclk));
	jdff dff_A_1pgpu9CU4_0(.dout(w_dff_A_pHvWiNJH2_0),.din(w_dff_A_1pgpu9CU4_0),.clk(gclk));
	jdff dff_A_pHvWiNJH2_0(.dout(w_dff_A_TxSgeTzU5_0),.din(w_dff_A_pHvWiNJH2_0),.clk(gclk));
	jdff dff_A_TxSgeTzU5_0(.dout(w_dff_A_9IYKVSVY5_0),.din(w_dff_A_TxSgeTzU5_0),.clk(gclk));
	jdff dff_A_9IYKVSVY5_0(.dout(w_dff_A_2ko0mDBe5_0),.din(w_dff_A_9IYKVSVY5_0),.clk(gclk));
	jdff dff_A_2ko0mDBe5_0(.dout(w_dff_A_XQVLFwgm0_0),.din(w_dff_A_2ko0mDBe5_0),.clk(gclk));
	jdff dff_A_XQVLFwgm0_0(.dout(w_dff_A_byuaIsk05_0),.din(w_dff_A_XQVLFwgm0_0),.clk(gclk));
	jdff dff_A_byuaIsk05_0(.dout(w_dff_A_JfdV9wNw2_0),.din(w_dff_A_byuaIsk05_0),.clk(gclk));
	jdff dff_A_JfdV9wNw2_0(.dout(w_dff_A_UqtS7VJR7_0),.din(w_dff_A_JfdV9wNw2_0),.clk(gclk));
	jdff dff_A_UqtS7VJR7_0(.dout(w_dff_A_HLHm30nX3_0),.din(w_dff_A_UqtS7VJR7_0),.clk(gclk));
	jdff dff_A_HLHm30nX3_0(.dout(w_dff_A_VkDpNVKu4_0),.din(w_dff_A_HLHm30nX3_0),.clk(gclk));
	jdff dff_A_VkDpNVKu4_0(.dout(w_dff_A_4qsKLjYg6_0),.din(w_dff_A_VkDpNVKu4_0),.clk(gclk));
	jdff dff_A_4qsKLjYg6_0(.dout(w_dff_A_nXrFq2gP6_0),.din(w_dff_A_4qsKLjYg6_0),.clk(gclk));
	jdff dff_A_nXrFq2gP6_0(.dout(w_dff_A_GLd1uF4g4_0),.din(w_dff_A_nXrFq2gP6_0),.clk(gclk));
	jdff dff_A_GLd1uF4g4_0(.dout(G873),.din(w_dff_A_GLd1uF4g4_0),.clk(gclk));
	jdff dff_A_ze09dhrl2_1(.dout(w_dff_A_GY1YKhKI1_0),.din(w_dff_A_ze09dhrl2_1),.clk(gclk));
	jdff dff_A_GY1YKhKI1_0(.dout(w_dff_A_0bLJJj1N7_0),.din(w_dff_A_GY1YKhKI1_0),.clk(gclk));
	jdff dff_A_0bLJJj1N7_0(.dout(w_dff_A_dpm6sj3J4_0),.din(w_dff_A_0bLJJj1N7_0),.clk(gclk));
	jdff dff_A_dpm6sj3J4_0(.dout(w_dff_A_q7zv4KAr1_0),.din(w_dff_A_dpm6sj3J4_0),.clk(gclk));
	jdff dff_A_q7zv4KAr1_0(.dout(w_dff_A_zNcILBaT1_0),.din(w_dff_A_q7zv4KAr1_0),.clk(gclk));
	jdff dff_A_zNcILBaT1_0(.dout(w_dff_A_um3UCFwv5_0),.din(w_dff_A_zNcILBaT1_0),.clk(gclk));
	jdff dff_A_um3UCFwv5_0(.dout(w_dff_A_Rn2xYR6i9_0),.din(w_dff_A_um3UCFwv5_0),.clk(gclk));
	jdff dff_A_Rn2xYR6i9_0(.dout(w_dff_A_AEgbe3eT1_0),.din(w_dff_A_Rn2xYR6i9_0),.clk(gclk));
	jdff dff_A_AEgbe3eT1_0(.dout(w_dff_A_uyPdBQa33_0),.din(w_dff_A_AEgbe3eT1_0),.clk(gclk));
	jdff dff_A_uyPdBQa33_0(.dout(w_dff_A_HDBvyhYh9_0),.din(w_dff_A_uyPdBQa33_0),.clk(gclk));
	jdff dff_A_HDBvyhYh9_0(.dout(w_dff_A_KnwHuFUu5_0),.din(w_dff_A_HDBvyhYh9_0),.clk(gclk));
	jdff dff_A_KnwHuFUu5_0(.dout(w_dff_A_paBzv8uy5_0),.din(w_dff_A_KnwHuFUu5_0),.clk(gclk));
	jdff dff_A_paBzv8uy5_0(.dout(w_dff_A_NTj0Pi5f6_0),.din(w_dff_A_paBzv8uy5_0),.clk(gclk));
	jdff dff_A_NTj0Pi5f6_0(.dout(w_dff_A_WlVZTu3x2_0),.din(w_dff_A_NTj0Pi5f6_0),.clk(gclk));
	jdff dff_A_WlVZTu3x2_0(.dout(w_dff_A_KkpLYZB45_0),.din(w_dff_A_WlVZTu3x2_0),.clk(gclk));
	jdff dff_A_KkpLYZB45_0(.dout(G875),.din(w_dff_A_KkpLYZB45_0),.clk(gclk));
	jdff dff_A_5ypKyrfN3_1(.dout(w_dff_A_bY06FGMf2_0),.din(w_dff_A_5ypKyrfN3_1),.clk(gclk));
	jdff dff_A_bY06FGMf2_0(.dout(w_dff_A_58dvA11K9_0),.din(w_dff_A_bY06FGMf2_0),.clk(gclk));
	jdff dff_A_58dvA11K9_0(.dout(w_dff_A_gAw9QXNE6_0),.din(w_dff_A_58dvA11K9_0),.clk(gclk));
	jdff dff_A_gAw9QXNE6_0(.dout(w_dff_A_ZYl6oI143_0),.din(w_dff_A_gAw9QXNE6_0),.clk(gclk));
	jdff dff_A_ZYl6oI143_0(.dout(w_dff_A_wYcYkfCu7_0),.din(w_dff_A_ZYl6oI143_0),.clk(gclk));
	jdff dff_A_wYcYkfCu7_0(.dout(w_dff_A_rhYpeoBP0_0),.din(w_dff_A_wYcYkfCu7_0),.clk(gclk));
	jdff dff_A_rhYpeoBP0_0(.dout(w_dff_A_DCkj2Yyc0_0),.din(w_dff_A_rhYpeoBP0_0),.clk(gclk));
	jdff dff_A_DCkj2Yyc0_0(.dout(w_dff_A_aYqoDzMp9_0),.din(w_dff_A_DCkj2Yyc0_0),.clk(gclk));
	jdff dff_A_aYqoDzMp9_0(.dout(w_dff_A_nD7vw8y92_0),.din(w_dff_A_aYqoDzMp9_0),.clk(gclk));
	jdff dff_A_nD7vw8y92_0(.dout(w_dff_A_NVLplX6H2_0),.din(w_dff_A_nD7vw8y92_0),.clk(gclk));
	jdff dff_A_NVLplX6H2_0(.dout(w_dff_A_jwAkuYzq7_0),.din(w_dff_A_NVLplX6H2_0),.clk(gclk));
	jdff dff_A_jwAkuYzq7_0(.dout(w_dff_A_dMmPU1zY1_0),.din(w_dff_A_jwAkuYzq7_0),.clk(gclk));
	jdff dff_A_dMmPU1zY1_0(.dout(w_dff_A_8mjvj9zO9_0),.din(w_dff_A_dMmPU1zY1_0),.clk(gclk));
	jdff dff_A_8mjvj9zO9_0(.dout(w_dff_A_0TjaEGZH2_0),.din(w_dff_A_8mjvj9zO9_0),.clk(gclk));
	jdff dff_A_0TjaEGZH2_0(.dout(w_dff_A_tib2Cl281_0),.din(w_dff_A_0TjaEGZH2_0),.clk(gclk));
	jdff dff_A_tib2Cl281_0(.dout(w_dff_A_nrb8HoE08_0),.din(w_dff_A_tib2Cl281_0),.clk(gclk));
	jdff dff_A_nrb8HoE08_0(.dout(G877),.din(w_dff_A_nrb8HoE08_0),.clk(gclk));
	jdff dff_A_neliHUfR6_1(.dout(w_dff_A_7ttjikvw7_0),.din(w_dff_A_neliHUfR6_1),.clk(gclk));
	jdff dff_A_7ttjikvw7_0(.dout(w_dff_A_0eA05yF12_0),.din(w_dff_A_7ttjikvw7_0),.clk(gclk));
	jdff dff_A_0eA05yF12_0(.dout(w_dff_A_f316JV8P5_0),.din(w_dff_A_0eA05yF12_0),.clk(gclk));
	jdff dff_A_f316JV8P5_0(.dout(w_dff_A_llQ1HV8w3_0),.din(w_dff_A_f316JV8P5_0),.clk(gclk));
	jdff dff_A_llQ1HV8w3_0(.dout(w_dff_A_qzEdIMsg0_0),.din(w_dff_A_llQ1HV8w3_0),.clk(gclk));
	jdff dff_A_qzEdIMsg0_0(.dout(w_dff_A_ooEUXoGn2_0),.din(w_dff_A_qzEdIMsg0_0),.clk(gclk));
	jdff dff_A_ooEUXoGn2_0(.dout(w_dff_A_x543VmWe4_0),.din(w_dff_A_ooEUXoGn2_0),.clk(gclk));
	jdff dff_A_x543VmWe4_0(.dout(w_dff_A_lAbSOpQ00_0),.din(w_dff_A_x543VmWe4_0),.clk(gclk));
	jdff dff_A_lAbSOpQ00_0(.dout(w_dff_A_28wg7lft1_0),.din(w_dff_A_lAbSOpQ00_0),.clk(gclk));
	jdff dff_A_28wg7lft1_0(.dout(w_dff_A_0Hr276hO9_0),.din(w_dff_A_28wg7lft1_0),.clk(gclk));
	jdff dff_A_0Hr276hO9_0(.dout(w_dff_A_mnDWZTTI2_0),.din(w_dff_A_0Hr276hO9_0),.clk(gclk));
	jdff dff_A_mnDWZTTI2_0(.dout(w_dff_A_CeiUXsYt1_0),.din(w_dff_A_mnDWZTTI2_0),.clk(gclk));
	jdff dff_A_CeiUXsYt1_0(.dout(w_dff_A_NlECMc2a2_0),.din(w_dff_A_CeiUXsYt1_0),.clk(gclk));
	jdff dff_A_NlECMc2a2_0(.dout(w_dff_A_mLxXGnTj0_0),.din(w_dff_A_NlECMc2a2_0),.clk(gclk));
	jdff dff_A_mLxXGnTj0_0(.dout(w_dff_A_X1wFQt2W8_0),.din(w_dff_A_mLxXGnTj0_0),.clk(gclk));
	jdff dff_A_X1wFQt2W8_0(.dout(w_dff_A_usXJEJZa3_0),.din(w_dff_A_X1wFQt2W8_0),.clk(gclk));
	jdff dff_A_usXJEJZa3_0(.dout(w_dff_A_wdxWV2EP4_0),.din(w_dff_A_usXJEJZa3_0),.clk(gclk));
	jdff dff_A_wdxWV2EP4_0(.dout(w_dff_A_WudY5Sp28_0),.din(w_dff_A_wdxWV2EP4_0),.clk(gclk));
	jdff dff_A_WudY5Sp28_0(.dout(w_dff_A_pALQTfio4_0),.din(w_dff_A_WudY5Sp28_0),.clk(gclk));
	jdff dff_A_pALQTfio4_0(.dout(G998),.din(w_dff_A_pALQTfio4_0),.clk(gclk));
	jdff dff_A_KTZtqfg71_1(.dout(w_dff_A_JQ0oYLoT5_0),.din(w_dff_A_KTZtqfg71_1),.clk(gclk));
	jdff dff_A_JQ0oYLoT5_0(.dout(w_dff_A_9Aue2sDH9_0),.din(w_dff_A_JQ0oYLoT5_0),.clk(gclk));
	jdff dff_A_9Aue2sDH9_0(.dout(w_dff_A_xXSErffV0_0),.din(w_dff_A_9Aue2sDH9_0),.clk(gclk));
	jdff dff_A_xXSErffV0_0(.dout(w_dff_A_ElVZFpBl4_0),.din(w_dff_A_xXSErffV0_0),.clk(gclk));
	jdff dff_A_ElVZFpBl4_0(.dout(w_dff_A_efKfqH7a0_0),.din(w_dff_A_ElVZFpBl4_0),.clk(gclk));
	jdff dff_A_efKfqH7a0_0(.dout(w_dff_A_v6ULwx0z3_0),.din(w_dff_A_efKfqH7a0_0),.clk(gclk));
	jdff dff_A_v6ULwx0z3_0(.dout(w_dff_A_ZUq3jIUF3_0),.din(w_dff_A_v6ULwx0z3_0),.clk(gclk));
	jdff dff_A_ZUq3jIUF3_0(.dout(w_dff_A_1ujXqndR2_0),.din(w_dff_A_ZUq3jIUF3_0),.clk(gclk));
	jdff dff_A_1ujXqndR2_0(.dout(w_dff_A_UtlVHKJ78_0),.din(w_dff_A_1ujXqndR2_0),.clk(gclk));
	jdff dff_A_UtlVHKJ78_0(.dout(w_dff_A_fde4e3wZ3_0),.din(w_dff_A_UtlVHKJ78_0),.clk(gclk));
	jdff dff_A_fde4e3wZ3_0(.dout(w_dff_A_rt8TLl1A4_0),.din(w_dff_A_fde4e3wZ3_0),.clk(gclk));
	jdff dff_A_rt8TLl1A4_0(.dout(w_dff_A_zwAXs2pp4_0),.din(w_dff_A_rt8TLl1A4_0),.clk(gclk));
	jdff dff_A_zwAXs2pp4_0(.dout(w_dff_A_JqUsGe384_0),.din(w_dff_A_zwAXs2pp4_0),.clk(gclk));
	jdff dff_A_JqUsGe384_0(.dout(w_dff_A_PQrMPFrc2_0),.din(w_dff_A_JqUsGe384_0),.clk(gclk));
	jdff dff_A_PQrMPFrc2_0(.dout(w_dff_A_QsE1JNbt4_0),.din(w_dff_A_PQrMPFrc2_0),.clk(gclk));
	jdff dff_A_QsE1JNbt4_0(.dout(w_dff_A_tKPhJvgs8_0),.din(w_dff_A_QsE1JNbt4_0),.clk(gclk));
	jdff dff_A_tKPhJvgs8_0(.dout(w_dff_A_rPaLxlP80_0),.din(w_dff_A_tKPhJvgs8_0),.clk(gclk));
	jdff dff_A_rPaLxlP80_0(.dout(w_dff_A_qJgPZP9y1_0),.din(w_dff_A_rPaLxlP80_0),.clk(gclk));
	jdff dff_A_qJgPZP9y1_0(.dout(G1000),.din(w_dff_A_qJgPZP9y1_0),.clk(gclk));
	jdff dff_A_oFxVWF266_2(.dout(w_dff_A_9wPjBMDI0_0),.din(w_dff_A_oFxVWF266_2),.clk(gclk));
	jdff dff_A_9wPjBMDI0_0(.dout(w_dff_A_Mjw2P9eH3_0),.din(w_dff_A_9wPjBMDI0_0),.clk(gclk));
	jdff dff_A_Mjw2P9eH3_0(.dout(w_dff_A_ahniAdbA5_0),.din(w_dff_A_Mjw2P9eH3_0),.clk(gclk));
	jdff dff_A_ahniAdbA5_0(.dout(w_dff_A_cJf3CJ8Y8_0),.din(w_dff_A_ahniAdbA5_0),.clk(gclk));
	jdff dff_A_cJf3CJ8Y8_0(.dout(w_dff_A_tw4viNqM8_0),.din(w_dff_A_cJf3CJ8Y8_0),.clk(gclk));
	jdff dff_A_tw4viNqM8_0(.dout(w_dff_A_u2371pY15_0),.din(w_dff_A_tw4viNqM8_0),.clk(gclk));
	jdff dff_A_u2371pY15_0(.dout(w_dff_A_M2Ic8DYe9_0),.din(w_dff_A_u2371pY15_0),.clk(gclk));
	jdff dff_A_M2Ic8DYe9_0(.dout(G575),.din(w_dff_A_M2Ic8DYe9_0),.clk(gclk));
	jdff dff_A_eSkGMLfB8_2(.dout(w_dff_A_Bjhe3bq82_0),.din(w_dff_A_eSkGMLfB8_2),.clk(gclk));
	jdff dff_A_Bjhe3bq82_0(.dout(w_dff_A_OMVhnJ9u7_0),.din(w_dff_A_Bjhe3bq82_0),.clk(gclk));
	jdff dff_A_OMVhnJ9u7_0(.dout(w_dff_A_NftuWoC69_0),.din(w_dff_A_OMVhnJ9u7_0),.clk(gclk));
	jdff dff_A_NftuWoC69_0(.dout(w_dff_A_1GsB7OMm0_0),.din(w_dff_A_NftuWoC69_0),.clk(gclk));
	jdff dff_A_1GsB7OMm0_0(.dout(w_dff_A_kw1x1V6S9_0),.din(w_dff_A_1GsB7OMm0_0),.clk(gclk));
	jdff dff_A_kw1x1V6S9_0(.dout(w_dff_A_9UfzsOYJ1_0),.din(w_dff_A_kw1x1V6S9_0),.clk(gclk));
	jdff dff_A_9UfzsOYJ1_0(.dout(G585),.din(w_dff_A_9UfzsOYJ1_0),.clk(gclk));
	jdff dff_A_IUyZibeU2_2(.dout(w_dff_A_cRRCAO2L6_0),.din(w_dff_A_IUyZibeU2_2),.clk(gclk));
	jdff dff_A_cRRCAO2L6_0(.dout(w_dff_A_svkJMgjO6_0),.din(w_dff_A_cRRCAO2L6_0),.clk(gclk));
	jdff dff_A_svkJMgjO6_0(.dout(w_dff_A_5ugU9kF67_0),.din(w_dff_A_svkJMgjO6_0),.clk(gclk));
	jdff dff_A_5ugU9kF67_0(.dout(w_dff_A_qqoXLBA01_0),.din(w_dff_A_5ugU9kF67_0),.clk(gclk));
	jdff dff_A_qqoXLBA01_0(.dout(w_dff_A_jqb47BX42_0),.din(w_dff_A_qqoXLBA01_0),.clk(gclk));
	jdff dff_A_jqb47BX42_0(.dout(w_dff_A_lA1THRZE0_0),.din(w_dff_A_jqb47BX42_0),.clk(gclk));
	jdff dff_A_lA1THRZE0_0(.dout(w_dff_A_mOyMGvcL5_0),.din(w_dff_A_lA1THRZE0_0),.clk(gclk));
	jdff dff_A_mOyMGvcL5_0(.dout(w_dff_A_51ahXK5G8_0),.din(w_dff_A_mOyMGvcL5_0),.clk(gclk));
	jdff dff_A_51ahXK5G8_0(.dout(w_dff_A_0HRDwkhQ6_0),.din(w_dff_A_51ahXK5G8_0),.clk(gclk));
	jdff dff_A_0HRDwkhQ6_0(.dout(w_dff_A_dIWxw3nm3_0),.din(w_dff_A_0HRDwkhQ6_0),.clk(gclk));
	jdff dff_A_dIWxw3nm3_0(.dout(w_dff_A_PSgSGnz36_0),.din(w_dff_A_dIWxw3nm3_0),.clk(gclk));
	jdff dff_A_PSgSGnz36_0(.dout(G661),.din(w_dff_A_PSgSGnz36_0),.clk(gclk));
	jdff dff_A_cL0EQVCg1_2(.dout(w_dff_A_Dp0FxNQF2_0),.din(w_dff_A_cL0EQVCg1_2),.clk(gclk));
	jdff dff_A_Dp0FxNQF2_0(.dout(w_dff_A_w9Ynxlfk2_0),.din(w_dff_A_Dp0FxNQF2_0),.clk(gclk));
	jdff dff_A_w9Ynxlfk2_0(.dout(w_dff_A_i95OBmFU3_0),.din(w_dff_A_w9Ynxlfk2_0),.clk(gclk));
	jdff dff_A_i95OBmFU3_0(.dout(w_dff_A_AX8U6Buc9_0),.din(w_dff_A_i95OBmFU3_0),.clk(gclk));
	jdff dff_A_AX8U6Buc9_0(.dout(w_dff_A_2EiIwpA04_0),.din(w_dff_A_AX8U6Buc9_0),.clk(gclk));
	jdff dff_A_2EiIwpA04_0(.dout(w_dff_A_W5mBCs2L4_0),.din(w_dff_A_2EiIwpA04_0),.clk(gclk));
	jdff dff_A_W5mBCs2L4_0(.dout(w_dff_A_bLo8VeWw5_0),.din(w_dff_A_W5mBCs2L4_0),.clk(gclk));
	jdff dff_A_bLo8VeWw5_0(.dout(w_dff_A_kS2MxYg51_0),.din(w_dff_A_bLo8VeWw5_0),.clk(gclk));
	jdff dff_A_kS2MxYg51_0(.dout(w_dff_A_6g9mpdPq0_0),.din(w_dff_A_kS2MxYg51_0),.clk(gclk));
	jdff dff_A_6g9mpdPq0_0(.dout(w_dff_A_wlRpliVa4_0),.din(w_dff_A_6g9mpdPq0_0),.clk(gclk));
	jdff dff_A_wlRpliVa4_0(.dout(w_dff_A_k7Y6xbUH1_0),.din(w_dff_A_wlRpliVa4_0),.clk(gclk));
	jdff dff_A_k7Y6xbUH1_0(.dout(G693),.din(w_dff_A_k7Y6xbUH1_0),.clk(gclk));
	jdff dff_A_IGyoSSEu8_2(.dout(w_dff_A_fnYfrLi49_0),.din(w_dff_A_IGyoSSEu8_2),.clk(gclk));
	jdff dff_A_fnYfrLi49_0(.dout(w_dff_A_07csGbv03_0),.din(w_dff_A_fnYfrLi49_0),.clk(gclk));
	jdff dff_A_07csGbv03_0(.dout(w_dff_A_V8THRWGJ7_0),.din(w_dff_A_07csGbv03_0),.clk(gclk));
	jdff dff_A_V8THRWGJ7_0(.dout(w_dff_A_u1LgeGkp8_0),.din(w_dff_A_V8THRWGJ7_0),.clk(gclk));
	jdff dff_A_u1LgeGkp8_0(.dout(w_dff_A_O0C8QJB56_0),.din(w_dff_A_u1LgeGkp8_0),.clk(gclk));
	jdff dff_A_O0C8QJB56_0(.dout(w_dff_A_6Seknxoa1_0),.din(w_dff_A_O0C8QJB56_0),.clk(gclk));
	jdff dff_A_6Seknxoa1_0(.dout(w_dff_A_gXRfmuoD9_0),.din(w_dff_A_6Seknxoa1_0),.clk(gclk));
	jdff dff_A_gXRfmuoD9_0(.dout(G747),.din(w_dff_A_gXRfmuoD9_0),.clk(gclk));
	jdff dff_A_56RrwCqu2_2(.dout(w_dff_A_XSBLuAK12_0),.din(w_dff_A_56RrwCqu2_2),.clk(gclk));
	jdff dff_A_XSBLuAK12_0(.dout(w_dff_A_TkCiHhqg2_0),.din(w_dff_A_XSBLuAK12_0),.clk(gclk));
	jdff dff_A_TkCiHhqg2_0(.dout(w_dff_A_iBUqbdgB6_0),.din(w_dff_A_TkCiHhqg2_0),.clk(gclk));
	jdff dff_A_iBUqbdgB6_0(.dout(w_dff_A_rqyikVq48_0),.din(w_dff_A_iBUqbdgB6_0),.clk(gclk));
	jdff dff_A_rqyikVq48_0(.dout(w_dff_A_rCYhtEKy0_0),.din(w_dff_A_rqyikVq48_0),.clk(gclk));
	jdff dff_A_rCYhtEKy0_0(.dout(w_dff_A_LoCEBRb97_0),.din(w_dff_A_rCYhtEKy0_0),.clk(gclk));
	jdff dff_A_LoCEBRb97_0(.dout(w_dff_A_tQ2JJ1wQ9_0),.din(w_dff_A_LoCEBRb97_0),.clk(gclk));
	jdff dff_A_tQ2JJ1wQ9_0(.dout(w_dff_A_3qtcbthX2_0),.din(w_dff_A_tQ2JJ1wQ9_0),.clk(gclk));
	jdff dff_A_3qtcbthX2_0(.dout(G752),.din(w_dff_A_3qtcbthX2_0),.clk(gclk));
	jdff dff_A_wwQGevd50_2(.dout(w_dff_A_LuCCvnEv7_0),.din(w_dff_A_wwQGevd50_2),.clk(gclk));
	jdff dff_A_LuCCvnEv7_0(.dout(w_dff_A_iOewLQyw8_0),.din(w_dff_A_LuCCvnEv7_0),.clk(gclk));
	jdff dff_A_iOewLQyw8_0(.dout(w_dff_A_J6hqywOG7_0),.din(w_dff_A_iOewLQyw8_0),.clk(gclk));
	jdff dff_A_J6hqywOG7_0(.dout(w_dff_A_i38oytxA1_0),.din(w_dff_A_J6hqywOG7_0),.clk(gclk));
	jdff dff_A_i38oytxA1_0(.dout(w_dff_A_EiYP8uzZ8_0),.din(w_dff_A_i38oytxA1_0),.clk(gclk));
	jdff dff_A_EiYP8uzZ8_0(.dout(w_dff_A_JMo9xqPC4_0),.din(w_dff_A_EiYP8uzZ8_0),.clk(gclk));
	jdff dff_A_JMo9xqPC4_0(.dout(w_dff_A_NHRKJE9o0_0),.din(w_dff_A_JMo9xqPC4_0),.clk(gclk));
	jdff dff_A_NHRKJE9o0_0(.dout(w_dff_A_vck6t0Ls7_0),.din(w_dff_A_NHRKJE9o0_0),.clk(gclk));
	jdff dff_A_vck6t0Ls7_0(.dout(w_dff_A_BCkQIoXj5_0),.din(w_dff_A_vck6t0Ls7_0),.clk(gclk));
	jdff dff_A_BCkQIoXj5_0(.dout(w_dff_A_zCFXhFnS0_0),.din(w_dff_A_BCkQIoXj5_0),.clk(gclk));
	jdff dff_A_zCFXhFnS0_0(.dout(G757),.din(w_dff_A_zCFXhFnS0_0),.clk(gclk));
	jdff dff_A_keQaPtPi2_2(.dout(w_dff_A_GuMAt2f15_0),.din(w_dff_A_keQaPtPi2_2),.clk(gclk));
	jdff dff_A_GuMAt2f15_0(.dout(w_dff_A_awe276pv0_0),.din(w_dff_A_GuMAt2f15_0),.clk(gclk));
	jdff dff_A_awe276pv0_0(.dout(w_dff_A_6vyJ4y485_0),.din(w_dff_A_awe276pv0_0),.clk(gclk));
	jdff dff_A_6vyJ4y485_0(.dout(w_dff_A_L2bcmLza9_0),.din(w_dff_A_6vyJ4y485_0),.clk(gclk));
	jdff dff_A_L2bcmLza9_0(.dout(w_dff_A_fUGivxGM4_0),.din(w_dff_A_L2bcmLza9_0),.clk(gclk));
	jdff dff_A_fUGivxGM4_0(.dout(w_dff_A_o0JrcGDO4_0),.din(w_dff_A_fUGivxGM4_0),.clk(gclk));
	jdff dff_A_o0JrcGDO4_0(.dout(w_dff_A_cYm2RJ1k5_0),.din(w_dff_A_o0JrcGDO4_0),.clk(gclk));
	jdff dff_A_cYm2RJ1k5_0(.dout(w_dff_A_uzM1zUeL4_0),.din(w_dff_A_cYm2RJ1k5_0),.clk(gclk));
	jdff dff_A_uzM1zUeL4_0(.dout(w_dff_A_tIXEG92T5_0),.din(w_dff_A_uzM1zUeL4_0),.clk(gclk));
	jdff dff_A_tIXEG92T5_0(.dout(G762),.din(w_dff_A_tIXEG92T5_0),.clk(gclk));
	jdff dff_A_7oyN7Kg98_2(.dout(w_dff_A_yrqbt1aF4_0),.din(w_dff_A_7oyN7Kg98_2),.clk(gclk));
	jdff dff_A_yrqbt1aF4_0(.dout(w_dff_A_15HlcQp52_0),.din(w_dff_A_yrqbt1aF4_0),.clk(gclk));
	jdff dff_A_15HlcQp52_0(.dout(w_dff_A_1LRZ8Qgk5_0),.din(w_dff_A_15HlcQp52_0),.clk(gclk));
	jdff dff_A_1LRZ8Qgk5_0(.dout(w_dff_A_eh7ZjtDn5_0),.din(w_dff_A_1LRZ8Qgk5_0),.clk(gclk));
	jdff dff_A_eh7ZjtDn5_0(.dout(w_dff_A_jjTVRLTX2_0),.din(w_dff_A_eh7ZjtDn5_0),.clk(gclk));
	jdff dff_A_jjTVRLTX2_0(.dout(w_dff_A_Q9ukMb3J0_0),.din(w_dff_A_jjTVRLTX2_0),.clk(gclk));
	jdff dff_A_Q9ukMb3J0_0(.dout(w_dff_A_GTOmaDn06_0),.din(w_dff_A_Q9ukMb3J0_0),.clk(gclk));
	jdff dff_A_GTOmaDn06_0(.dout(G787),.din(w_dff_A_GTOmaDn06_0),.clk(gclk));
	jdff dff_A_HwrRny5T3_2(.dout(w_dff_A_IZXO5wd74_0),.din(w_dff_A_HwrRny5T3_2),.clk(gclk));
	jdff dff_A_IZXO5wd74_0(.dout(w_dff_A_R1pQn5dn0_0),.din(w_dff_A_IZXO5wd74_0),.clk(gclk));
	jdff dff_A_R1pQn5dn0_0(.dout(w_dff_A_kWHmk5Ik3_0),.din(w_dff_A_R1pQn5dn0_0),.clk(gclk));
	jdff dff_A_kWHmk5Ik3_0(.dout(w_dff_A_E7lF4cOj9_0),.din(w_dff_A_kWHmk5Ik3_0),.clk(gclk));
	jdff dff_A_E7lF4cOj9_0(.dout(w_dff_A_LaEpSJrB2_0),.din(w_dff_A_E7lF4cOj9_0),.clk(gclk));
	jdff dff_A_LaEpSJrB2_0(.dout(w_dff_A_mT5BA4oI3_0),.din(w_dff_A_LaEpSJrB2_0),.clk(gclk));
	jdff dff_A_mT5BA4oI3_0(.dout(w_dff_A_erYO3d858_0),.din(w_dff_A_mT5BA4oI3_0),.clk(gclk));
	jdff dff_A_erYO3d858_0(.dout(w_dff_A_KWCJk61z9_0),.din(w_dff_A_erYO3d858_0),.clk(gclk));
	jdff dff_A_KWCJk61z9_0(.dout(G792),.din(w_dff_A_KWCJk61z9_0),.clk(gclk));
	jdff dff_A_hBJRCEio6_2(.dout(w_dff_A_4lWHOGkr7_0),.din(w_dff_A_hBJRCEio6_2),.clk(gclk));
	jdff dff_A_4lWHOGkr7_0(.dout(w_dff_A_R7L5ePMw5_0),.din(w_dff_A_4lWHOGkr7_0),.clk(gclk));
	jdff dff_A_R7L5ePMw5_0(.dout(w_dff_A_EonOOZV55_0),.din(w_dff_A_R7L5ePMw5_0),.clk(gclk));
	jdff dff_A_EonOOZV55_0(.dout(w_dff_A_z2Y2UXP12_0),.din(w_dff_A_EonOOZV55_0),.clk(gclk));
	jdff dff_A_z2Y2UXP12_0(.dout(w_dff_A_6M29mEZe3_0),.din(w_dff_A_z2Y2UXP12_0),.clk(gclk));
	jdff dff_A_6M29mEZe3_0(.dout(w_dff_A_35N0HQvi8_0),.din(w_dff_A_6M29mEZe3_0),.clk(gclk));
	jdff dff_A_35N0HQvi8_0(.dout(w_dff_A_nxmcxN7M2_0),.din(w_dff_A_35N0HQvi8_0),.clk(gclk));
	jdff dff_A_nxmcxN7M2_0(.dout(w_dff_A_pkA0WnTx7_0),.din(w_dff_A_nxmcxN7M2_0),.clk(gclk));
	jdff dff_A_pkA0WnTx7_0(.dout(w_dff_A_UyNzVoq93_0),.din(w_dff_A_pkA0WnTx7_0),.clk(gclk));
	jdff dff_A_UyNzVoq93_0(.dout(w_dff_A_YPP1kP491_0),.din(w_dff_A_UyNzVoq93_0),.clk(gclk));
	jdff dff_A_YPP1kP491_0(.dout(G797),.din(w_dff_A_YPP1kP491_0),.clk(gclk));
	jdff dff_A_kRGQhKKq4_2(.dout(w_dff_A_WIc5xmtn9_0),.din(w_dff_A_kRGQhKKq4_2),.clk(gclk));
	jdff dff_A_WIc5xmtn9_0(.dout(w_dff_A_BZfoMNOJ8_0),.din(w_dff_A_WIc5xmtn9_0),.clk(gclk));
	jdff dff_A_BZfoMNOJ8_0(.dout(w_dff_A_OKVU27gA8_0),.din(w_dff_A_BZfoMNOJ8_0),.clk(gclk));
	jdff dff_A_OKVU27gA8_0(.dout(w_dff_A_6M90IALQ6_0),.din(w_dff_A_OKVU27gA8_0),.clk(gclk));
	jdff dff_A_6M90IALQ6_0(.dout(w_dff_A_22v3171a1_0),.din(w_dff_A_6M90IALQ6_0),.clk(gclk));
	jdff dff_A_22v3171a1_0(.dout(w_dff_A_pnzLAGUv5_0),.din(w_dff_A_22v3171a1_0),.clk(gclk));
	jdff dff_A_pnzLAGUv5_0(.dout(w_dff_A_MrILsDGm1_0),.din(w_dff_A_pnzLAGUv5_0),.clk(gclk));
	jdff dff_A_MrILsDGm1_0(.dout(w_dff_A_QaFzE0QM7_0),.din(w_dff_A_MrILsDGm1_0),.clk(gclk));
	jdff dff_A_QaFzE0QM7_0(.dout(w_dff_A_OZueif6j5_0),.din(w_dff_A_QaFzE0QM7_0),.clk(gclk));
	jdff dff_A_OZueif6j5_0(.dout(G802),.din(w_dff_A_OZueif6j5_0),.clk(gclk));
	jdff dff_A_wjAAGGZN0_2(.dout(w_dff_A_g6WAay8Z1_0),.din(w_dff_A_wjAAGGZN0_2),.clk(gclk));
	jdff dff_A_g6WAay8Z1_0(.dout(w_dff_A_JHpN8vBq4_0),.din(w_dff_A_g6WAay8Z1_0),.clk(gclk));
	jdff dff_A_JHpN8vBq4_0(.dout(w_dff_A_kPOWcMVs8_0),.din(w_dff_A_JHpN8vBq4_0),.clk(gclk));
	jdff dff_A_kPOWcMVs8_0(.dout(w_dff_A_reObvyOt0_0),.din(w_dff_A_kPOWcMVs8_0),.clk(gclk));
	jdff dff_A_reObvyOt0_0(.dout(w_dff_A_mX0XWHp30_0),.din(w_dff_A_reObvyOt0_0),.clk(gclk));
	jdff dff_A_mX0XWHp30_0(.dout(w_dff_A_kFMhfeua5_0),.din(w_dff_A_mX0XWHp30_0),.clk(gclk));
	jdff dff_A_kFMhfeua5_0(.dout(G642),.din(w_dff_A_kFMhfeua5_0),.clk(gclk));
	jdff dff_A_kbovglEb0_2(.dout(w_dff_A_kYSdAvvG4_0),.din(w_dff_A_kbovglEb0_2),.clk(gclk));
	jdff dff_A_kYSdAvvG4_0(.dout(w_dff_A_aF8eCFso6_0),.din(w_dff_A_kYSdAvvG4_0),.clk(gclk));
	jdff dff_A_aF8eCFso6_0(.dout(w_dff_A_GjRz2egv7_0),.din(w_dff_A_aF8eCFso6_0),.clk(gclk));
	jdff dff_A_GjRz2egv7_0(.dout(w_dff_A_AwlHth9f5_0),.din(w_dff_A_GjRz2egv7_0),.clk(gclk));
	jdff dff_A_AwlHth9f5_0(.dout(w_dff_A_LviuiotL2_0),.din(w_dff_A_AwlHth9f5_0),.clk(gclk));
	jdff dff_A_LviuiotL2_0(.dout(w_dff_A_AINrNPxn4_0),.din(w_dff_A_LviuiotL2_0),.clk(gclk));
	jdff dff_A_AINrNPxn4_0(.dout(w_dff_A_rE8qxiW14_0),.din(w_dff_A_AINrNPxn4_0),.clk(gclk));
	jdff dff_A_rE8qxiW14_0(.dout(w_dff_A_u3zsD5KS2_0),.din(w_dff_A_rE8qxiW14_0),.clk(gclk));
	jdff dff_A_u3zsD5KS2_0(.dout(w_dff_A_fxDlBdr66_0),.din(w_dff_A_u3zsD5KS2_0),.clk(gclk));
	jdff dff_A_fxDlBdr66_0(.dout(G664),.din(w_dff_A_fxDlBdr66_0),.clk(gclk));
	jdff dff_A_ss9SJ2Xo4_2(.dout(w_dff_A_P0Dx8lPm9_0),.din(w_dff_A_ss9SJ2Xo4_2),.clk(gclk));
	jdff dff_A_P0Dx8lPm9_0(.dout(w_dff_A_0Etvfc4Q2_0),.din(w_dff_A_P0Dx8lPm9_0),.clk(gclk));
	jdff dff_A_0Etvfc4Q2_0(.dout(w_dff_A_qFpBRhTS2_0),.din(w_dff_A_0Etvfc4Q2_0),.clk(gclk));
	jdff dff_A_qFpBRhTS2_0(.dout(w_dff_A_zdbF1X6j9_0),.din(w_dff_A_qFpBRhTS2_0),.clk(gclk));
	jdff dff_A_zdbF1X6j9_0(.dout(w_dff_A_4yIGQfuL3_0),.din(w_dff_A_zdbF1X6j9_0),.clk(gclk));
	jdff dff_A_4yIGQfuL3_0(.dout(w_dff_A_pXW0sItH6_0),.din(w_dff_A_4yIGQfuL3_0),.clk(gclk));
	jdff dff_A_pXW0sItH6_0(.dout(w_dff_A_Ox42J1yh8_0),.din(w_dff_A_pXW0sItH6_0),.clk(gclk));
	jdff dff_A_Ox42J1yh8_0(.dout(w_dff_A_pU10xJRe7_0),.din(w_dff_A_Ox42J1yh8_0),.clk(gclk));
	jdff dff_A_pU10xJRe7_0(.dout(w_dff_A_sK2mi3pL2_0),.din(w_dff_A_pU10xJRe7_0),.clk(gclk));
	jdff dff_A_sK2mi3pL2_0(.dout(G667),.din(w_dff_A_sK2mi3pL2_0),.clk(gclk));
	jdff dff_A_tBBw127J7_2(.dout(w_dff_A_oYjsusMY9_0),.din(w_dff_A_tBBw127J7_2),.clk(gclk));
	jdff dff_A_oYjsusMY9_0(.dout(w_dff_A_CytBECid0_0),.din(w_dff_A_oYjsusMY9_0),.clk(gclk));
	jdff dff_A_CytBECid0_0(.dout(w_dff_A_IhNYKsG56_0),.din(w_dff_A_CytBECid0_0),.clk(gclk));
	jdff dff_A_IhNYKsG56_0(.dout(w_dff_A_1ual1f6d6_0),.din(w_dff_A_IhNYKsG56_0),.clk(gclk));
	jdff dff_A_1ual1f6d6_0(.dout(w_dff_A_cdKTJHI05_0),.din(w_dff_A_1ual1f6d6_0),.clk(gclk));
	jdff dff_A_cdKTJHI05_0(.dout(w_dff_A_FkZIukp17_0),.din(w_dff_A_cdKTJHI05_0),.clk(gclk));
	jdff dff_A_FkZIukp17_0(.dout(w_dff_A_qzhJV5k79_0),.din(w_dff_A_FkZIukp17_0),.clk(gclk));
	jdff dff_A_qzhJV5k79_0(.dout(w_dff_A_ogcvh6NP5_0),.din(w_dff_A_qzhJV5k79_0),.clk(gclk));
	jdff dff_A_ogcvh6NP5_0(.dout(G670),.din(w_dff_A_ogcvh6NP5_0),.clk(gclk));
	jdff dff_A_FJ4eLE8y0_2(.dout(w_dff_A_PYdsn7pj3_0),.din(w_dff_A_FJ4eLE8y0_2),.clk(gclk));
	jdff dff_A_PYdsn7pj3_0(.dout(w_dff_A_DHmYaf239_0),.din(w_dff_A_PYdsn7pj3_0),.clk(gclk));
	jdff dff_A_DHmYaf239_0(.dout(w_dff_A_7mmAos5b6_0),.din(w_dff_A_DHmYaf239_0),.clk(gclk));
	jdff dff_A_7mmAos5b6_0(.dout(w_dff_A_9KSwdT595_0),.din(w_dff_A_7mmAos5b6_0),.clk(gclk));
	jdff dff_A_9KSwdT595_0(.dout(w_dff_A_FoxYZBO38_0),.din(w_dff_A_9KSwdT595_0),.clk(gclk));
	jdff dff_A_FoxYZBO38_0(.dout(G676),.din(w_dff_A_FoxYZBO38_0),.clk(gclk));
	jdff dff_A_aPMm9gZk7_2(.dout(w_dff_A_3d66GSyw0_0),.din(w_dff_A_aPMm9gZk7_2),.clk(gclk));
	jdff dff_A_3d66GSyw0_0(.dout(w_dff_A_6f2ZC6wu8_0),.din(w_dff_A_3d66GSyw0_0),.clk(gclk));
	jdff dff_A_6f2ZC6wu8_0(.dout(w_dff_A_G0NcBXiA6_0),.din(w_dff_A_6f2ZC6wu8_0),.clk(gclk));
	jdff dff_A_G0NcBXiA6_0(.dout(w_dff_A_ray4PLmV4_0),.din(w_dff_A_G0NcBXiA6_0),.clk(gclk));
	jdff dff_A_ray4PLmV4_0(.dout(w_dff_A_e1CuurEu2_0),.din(w_dff_A_ray4PLmV4_0),.clk(gclk));
	jdff dff_A_e1CuurEu2_0(.dout(w_dff_A_aZGTDgYD1_0),.din(w_dff_A_e1CuurEu2_0),.clk(gclk));
	jdff dff_A_aZGTDgYD1_0(.dout(w_dff_A_fOOG70532_0),.din(w_dff_A_aZGTDgYD1_0),.clk(gclk));
	jdff dff_A_fOOG70532_0(.dout(w_dff_A_HSBN9R1w9_0),.din(w_dff_A_fOOG70532_0),.clk(gclk));
	jdff dff_A_HSBN9R1w9_0(.dout(w_dff_A_7QjQD5T44_0),.din(w_dff_A_HSBN9R1w9_0),.clk(gclk));
	jdff dff_A_7QjQD5T44_0(.dout(G696),.din(w_dff_A_7QjQD5T44_0),.clk(gclk));
	jdff dff_A_E416vl2P8_2(.dout(w_dff_A_P2jh8dN06_0),.din(w_dff_A_E416vl2P8_2),.clk(gclk));
	jdff dff_A_P2jh8dN06_0(.dout(w_dff_A_crW3mDMJ7_0),.din(w_dff_A_P2jh8dN06_0),.clk(gclk));
	jdff dff_A_crW3mDMJ7_0(.dout(w_dff_A_D00Sfr7D3_0),.din(w_dff_A_crW3mDMJ7_0),.clk(gclk));
	jdff dff_A_D00Sfr7D3_0(.dout(w_dff_A_sVFNQS8M3_0),.din(w_dff_A_D00Sfr7D3_0),.clk(gclk));
	jdff dff_A_sVFNQS8M3_0(.dout(w_dff_A_Q4v9FAB68_0),.din(w_dff_A_sVFNQS8M3_0),.clk(gclk));
	jdff dff_A_Q4v9FAB68_0(.dout(w_dff_A_ZWBjnRSv6_0),.din(w_dff_A_Q4v9FAB68_0),.clk(gclk));
	jdff dff_A_ZWBjnRSv6_0(.dout(w_dff_A_Zk63SCOk5_0),.din(w_dff_A_ZWBjnRSv6_0),.clk(gclk));
	jdff dff_A_Zk63SCOk5_0(.dout(w_dff_A_J6AimyZZ1_0),.din(w_dff_A_Zk63SCOk5_0),.clk(gclk));
	jdff dff_A_J6AimyZZ1_0(.dout(w_dff_A_gIpfvbWy7_0),.din(w_dff_A_J6AimyZZ1_0),.clk(gclk));
	jdff dff_A_gIpfvbWy7_0(.dout(G699),.din(w_dff_A_gIpfvbWy7_0),.clk(gclk));
	jdff dff_A_88KRnGpV7_2(.dout(w_dff_A_cYNTIumU9_0),.din(w_dff_A_88KRnGpV7_2),.clk(gclk));
	jdff dff_A_cYNTIumU9_0(.dout(w_dff_A_qeJVB7y90_0),.din(w_dff_A_cYNTIumU9_0),.clk(gclk));
	jdff dff_A_qeJVB7y90_0(.dout(w_dff_A_iwUG8mUG7_0),.din(w_dff_A_qeJVB7y90_0),.clk(gclk));
	jdff dff_A_iwUG8mUG7_0(.dout(w_dff_A_Jeo8Nlfx1_0),.din(w_dff_A_iwUG8mUG7_0),.clk(gclk));
	jdff dff_A_Jeo8Nlfx1_0(.dout(w_dff_A_LXsOzG986_0),.din(w_dff_A_Jeo8Nlfx1_0),.clk(gclk));
	jdff dff_A_LXsOzG986_0(.dout(w_dff_A_UnA1ZE3e4_0),.din(w_dff_A_LXsOzG986_0),.clk(gclk));
	jdff dff_A_UnA1ZE3e4_0(.dout(w_dff_A_Ur1W488X2_0),.din(w_dff_A_UnA1ZE3e4_0),.clk(gclk));
	jdff dff_A_Ur1W488X2_0(.dout(w_dff_A_DjupPxtm5_0),.din(w_dff_A_Ur1W488X2_0),.clk(gclk));
	jdff dff_A_DjupPxtm5_0(.dout(G702),.din(w_dff_A_DjupPxtm5_0),.clk(gclk));
	jdff dff_A_oxuB7DjA9_2(.dout(w_dff_A_NxfNV3OH9_0),.din(w_dff_A_oxuB7DjA9_2),.clk(gclk));
	jdff dff_A_NxfNV3OH9_0(.dout(w_dff_A_OGGUHDmq4_0),.din(w_dff_A_NxfNV3OH9_0),.clk(gclk));
	jdff dff_A_OGGUHDmq4_0(.dout(w_dff_A_F598HQwd0_0),.din(w_dff_A_OGGUHDmq4_0),.clk(gclk));
	jdff dff_A_F598HQwd0_0(.dout(w_dff_A_rsCdqn5b3_0),.din(w_dff_A_F598HQwd0_0),.clk(gclk));
	jdff dff_A_rsCdqn5b3_0(.dout(w_dff_A_qIdEvIDR4_0),.din(w_dff_A_rsCdqn5b3_0),.clk(gclk));
	jdff dff_A_qIdEvIDR4_0(.dout(w_dff_A_RuC4hOr78_0),.din(w_dff_A_qIdEvIDR4_0),.clk(gclk));
	jdff dff_A_RuC4hOr78_0(.dout(G818),.din(w_dff_A_RuC4hOr78_0),.clk(gclk));
	jdff dff_A_jvwhkrDN8_2(.dout(w_dff_A_Y8d1aVOm5_0),.din(w_dff_A_jvwhkrDN8_2),.clk(gclk));
	jdff dff_A_Y8d1aVOm5_0(.dout(w_dff_A_WaqFKYA54_0),.din(w_dff_A_Y8d1aVOm5_0),.clk(gclk));
	jdff dff_A_WaqFKYA54_0(.dout(w_dff_A_0kpxCFv33_0),.din(w_dff_A_WaqFKYA54_0),.clk(gclk));
	jdff dff_A_0kpxCFv33_0(.dout(w_dff_A_2ii10nXG5_0),.din(w_dff_A_0kpxCFv33_0),.clk(gclk));
	jdff dff_A_2ii10nXG5_0(.dout(w_dff_A_vgKVjSJ16_0),.din(w_dff_A_2ii10nXG5_0),.clk(gclk));
	jdff dff_A_vgKVjSJ16_0(.dout(w_dff_A_2g2eiFvr1_0),.din(w_dff_A_vgKVjSJ16_0),.clk(gclk));
	jdff dff_A_2g2eiFvr1_0(.dout(w_dff_A_0BRhGLFc0_0),.din(w_dff_A_2g2eiFvr1_0),.clk(gclk));
	jdff dff_A_0BRhGLFc0_0(.dout(w_dff_A_j2omylgn7_0),.din(w_dff_A_0BRhGLFc0_0),.clk(gclk));
	jdff dff_A_j2omylgn7_0(.dout(w_dff_A_NIxKrJk80_0),.din(w_dff_A_j2omylgn7_0),.clk(gclk));
	jdff dff_A_NIxKrJk80_0(.dout(G813),.din(w_dff_A_NIxKrJk80_0),.clk(gclk));
	jdff dff_A_UrnIQvBs9_1(.dout(w_dff_A_z4hFqVTR2_0),.din(w_dff_A_UrnIQvBs9_1),.clk(gclk));
	jdff dff_A_z4hFqVTR2_0(.dout(w_dff_A_6GBVhRSQ7_0),.din(w_dff_A_z4hFqVTR2_0),.clk(gclk));
	jdff dff_A_6GBVhRSQ7_0(.dout(w_dff_A_790Qc8Pg4_0),.din(w_dff_A_6GBVhRSQ7_0),.clk(gclk));
	jdff dff_A_790Qc8Pg4_0(.dout(w_dff_A_SmfxvG303_0),.din(w_dff_A_790Qc8Pg4_0),.clk(gclk));
	jdff dff_A_SmfxvG303_0(.dout(w_dff_A_jqG8pdYj3_0),.din(w_dff_A_SmfxvG303_0),.clk(gclk));
	jdff dff_A_jqG8pdYj3_0(.dout(w_dff_A_piCXS0Pd0_0),.din(w_dff_A_jqG8pdYj3_0),.clk(gclk));
	jdff dff_A_piCXS0Pd0_0(.dout(G824),.din(w_dff_A_piCXS0Pd0_0),.clk(gclk));
	jdff dff_A_Fi5KrCYh7_1(.dout(w_dff_A_XU6G4Rnz6_0),.din(w_dff_A_Fi5KrCYh7_1),.clk(gclk));
	jdff dff_A_XU6G4Rnz6_0(.dout(w_dff_A_FOj9cwjG6_0),.din(w_dff_A_XU6G4Rnz6_0),.clk(gclk));
	jdff dff_A_FOj9cwjG6_0(.dout(w_dff_A_7UcrxjYU9_0),.din(w_dff_A_FOj9cwjG6_0),.clk(gclk));
	jdff dff_A_7UcrxjYU9_0(.dout(w_dff_A_W1WjV6JE5_0),.din(w_dff_A_7UcrxjYU9_0),.clk(gclk));
	jdff dff_A_W1WjV6JE5_0(.dout(w_dff_A_4GH99eSJ4_0),.din(w_dff_A_W1WjV6JE5_0),.clk(gclk));
	jdff dff_A_4GH99eSJ4_0(.dout(w_dff_A_Acvk601o3_0),.din(w_dff_A_4GH99eSJ4_0),.clk(gclk));
	jdff dff_A_Acvk601o3_0(.dout(w_dff_A_w03832J53_0),.din(w_dff_A_Acvk601o3_0),.clk(gclk));
	jdff dff_A_w03832J53_0(.dout(G826),.din(w_dff_A_w03832J53_0),.clk(gclk));
	jdff dff_A_5bYRvP0i0_1(.dout(w_dff_A_sfPU4EOk3_0),.din(w_dff_A_5bYRvP0i0_1),.clk(gclk));
	jdff dff_A_sfPU4EOk3_0(.dout(w_dff_A_BlEsbe956_0),.din(w_dff_A_sfPU4EOk3_0),.clk(gclk));
	jdff dff_A_BlEsbe956_0(.dout(w_dff_A_h3Ni1l6T0_0),.din(w_dff_A_BlEsbe956_0),.clk(gclk));
	jdff dff_A_h3Ni1l6T0_0(.dout(w_dff_A_EydOHUhY4_0),.din(w_dff_A_h3Ni1l6T0_0),.clk(gclk));
	jdff dff_A_EydOHUhY4_0(.dout(w_dff_A_7h98kp6x0_0),.din(w_dff_A_EydOHUhY4_0),.clk(gclk));
	jdff dff_A_7h98kp6x0_0(.dout(w_dff_A_whgDnFsH7_0),.din(w_dff_A_7h98kp6x0_0),.clk(gclk));
	jdff dff_A_whgDnFsH7_0(.dout(G828),.din(w_dff_A_whgDnFsH7_0),.clk(gclk));
	jdff dff_A_RKhsEVmw6_1(.dout(w_dff_A_Ps8KofOz1_0),.din(w_dff_A_RKhsEVmw6_1),.clk(gclk));
	jdff dff_A_Ps8KofOz1_0(.dout(w_dff_A_uOYJOAMV8_0),.din(w_dff_A_Ps8KofOz1_0),.clk(gclk));
	jdff dff_A_uOYJOAMV8_0(.dout(w_dff_A_KzkGDMLA5_0),.din(w_dff_A_uOYJOAMV8_0),.clk(gclk));
	jdff dff_A_KzkGDMLA5_0(.dout(w_dff_A_N3n9LPEy2_0),.din(w_dff_A_KzkGDMLA5_0),.clk(gclk));
	jdff dff_A_N3n9LPEy2_0(.dout(w_dff_A_mA14aquq8_0),.din(w_dff_A_N3n9LPEy2_0),.clk(gclk));
	jdff dff_A_mA14aquq8_0(.dout(w_dff_A_GHyijkEL1_0),.din(w_dff_A_mA14aquq8_0),.clk(gclk));
	jdff dff_A_GHyijkEL1_0(.dout(w_dff_A_V6fy43pr2_0),.din(w_dff_A_GHyijkEL1_0),.clk(gclk));
	jdff dff_A_V6fy43pr2_0(.dout(w_dff_A_R4gtxDkT9_0),.din(w_dff_A_V6fy43pr2_0),.clk(gclk));
	jdff dff_A_R4gtxDkT9_0(.dout(w_dff_A_zcwqaNIL1_0),.din(w_dff_A_R4gtxDkT9_0),.clk(gclk));
	jdff dff_A_zcwqaNIL1_0(.dout(w_dff_A_P3klW2aS8_0),.din(w_dff_A_zcwqaNIL1_0),.clk(gclk));
	jdff dff_A_P3klW2aS8_0(.dout(w_dff_A_grsRAp8K6_0),.din(w_dff_A_P3klW2aS8_0),.clk(gclk));
	jdff dff_A_grsRAp8K6_0(.dout(G830),.din(w_dff_A_grsRAp8K6_0),.clk(gclk));
	jdff dff_A_vafD6ff48_2(.dout(w_dff_A_NHbc80Du1_0),.din(w_dff_A_vafD6ff48_2),.clk(gclk));
	jdff dff_A_NHbc80Du1_0(.dout(w_dff_A_GjT1u7DS1_0),.din(w_dff_A_NHbc80Du1_0),.clk(gclk));
	jdff dff_A_GjT1u7DS1_0(.dout(w_dff_A_egeNTtbU8_0),.din(w_dff_A_GjT1u7DS1_0),.clk(gclk));
	jdff dff_A_egeNTtbU8_0(.dout(w_dff_A_lZi2bb4Y7_0),.din(w_dff_A_egeNTtbU8_0),.clk(gclk));
	jdff dff_A_lZi2bb4Y7_0(.dout(w_dff_A_WSu8YH2N6_0),.din(w_dff_A_lZi2bb4Y7_0),.clk(gclk));
	jdff dff_A_WSu8YH2N6_0(.dout(w_dff_A_YgU5vIS79_0),.din(w_dff_A_WSu8YH2N6_0),.clk(gclk));
	jdff dff_A_YgU5vIS79_0(.dout(w_dff_A_yLvlILzf0_0),.din(w_dff_A_YgU5vIS79_0),.clk(gclk));
	jdff dff_A_yLvlILzf0_0(.dout(w_dff_A_6H7heQwo1_0),.din(w_dff_A_yLvlILzf0_0),.clk(gclk));
	jdff dff_A_6H7heQwo1_0(.dout(w_dff_A_WDpuXTtO2_0),.din(w_dff_A_6H7heQwo1_0),.clk(gclk));
	jdff dff_A_WDpuXTtO2_0(.dout(w_dff_A_iYgPbrkt8_0),.din(w_dff_A_WDpuXTtO2_0),.clk(gclk));
	jdff dff_A_iYgPbrkt8_0(.dout(w_dff_A_cJaLg3Re5_0),.din(w_dff_A_iYgPbrkt8_0),.clk(gclk));
	jdff dff_A_cJaLg3Re5_0(.dout(w_dff_A_wJrX1xWD4_0),.din(w_dff_A_cJaLg3Re5_0),.clk(gclk));
	jdff dff_A_wJrX1xWD4_0(.dout(w_dff_A_aeYc1dxD1_0),.din(w_dff_A_wJrX1xWD4_0),.clk(gclk));
	jdff dff_A_aeYc1dxD1_0(.dout(w_dff_A_GlxHJIEL1_0),.din(w_dff_A_aeYc1dxD1_0),.clk(gclk));
	jdff dff_A_GlxHJIEL1_0(.dout(w_dff_A_d4XYNGRD4_0),.din(w_dff_A_GlxHJIEL1_0),.clk(gclk));
	jdff dff_A_d4XYNGRD4_0(.dout(w_dff_A_sEelVtlB0_0),.din(w_dff_A_d4XYNGRD4_0),.clk(gclk));
	jdff dff_A_sEelVtlB0_0(.dout(G854),.din(w_dff_A_sEelVtlB0_0),.clk(gclk));
	jdff dff_A_MInp1sVP2_1(.dout(w_dff_A_spmEkXTn4_0),.din(w_dff_A_MInp1sVP2_1),.clk(gclk));
	jdff dff_A_spmEkXTn4_0(.dout(w_dff_A_jWlY2xyu9_0),.din(w_dff_A_spmEkXTn4_0),.clk(gclk));
	jdff dff_A_jWlY2xyu9_0(.dout(w_dff_A_NOkych6E0_0),.din(w_dff_A_jWlY2xyu9_0),.clk(gclk));
	jdff dff_A_NOkych6E0_0(.dout(w_dff_A_4ojF5srM0_0),.din(w_dff_A_NOkych6E0_0),.clk(gclk));
	jdff dff_A_4ojF5srM0_0(.dout(w_dff_A_Zf2BjFUE2_0),.din(w_dff_A_4ojF5srM0_0),.clk(gclk));
	jdff dff_A_Zf2BjFUE2_0(.dout(G863),.din(w_dff_A_Zf2BjFUE2_0),.clk(gclk));
	jdff dff_A_cJBm3tzC8_1(.dout(w_dff_A_TTTwWwf34_0),.din(w_dff_A_cJBm3tzC8_1),.clk(gclk));
	jdff dff_A_TTTwWwf34_0(.dout(w_dff_A_LhvBKKL64_0),.din(w_dff_A_TTTwWwf34_0),.clk(gclk));
	jdff dff_A_LhvBKKL64_0(.dout(w_dff_A_28qXxs1M3_0),.din(w_dff_A_LhvBKKL64_0),.clk(gclk));
	jdff dff_A_28qXxs1M3_0(.dout(w_dff_A_eFsPG5Va8_0),.din(w_dff_A_28qXxs1M3_0),.clk(gclk));
	jdff dff_A_eFsPG5Va8_0(.dout(w_dff_A_Il93Y7Ju3_0),.din(w_dff_A_eFsPG5Va8_0),.clk(gclk));
	jdff dff_A_Il93Y7Ju3_0(.dout(w_dff_A_so1IeFct6_0),.din(w_dff_A_Il93Y7Ju3_0),.clk(gclk));
	jdff dff_A_so1IeFct6_0(.dout(w_dff_A_JRyMNrnF2_0),.din(w_dff_A_so1IeFct6_0),.clk(gclk));
	jdff dff_A_JRyMNrnF2_0(.dout(w_dff_A_G5tlOvfn8_0),.din(w_dff_A_JRyMNrnF2_0),.clk(gclk));
	jdff dff_A_G5tlOvfn8_0(.dout(G865),.din(w_dff_A_G5tlOvfn8_0),.clk(gclk));
	jdff dff_A_CZVTd2RE5_1(.dout(w_dff_A_wlNhtr8z1_0),.din(w_dff_A_CZVTd2RE5_1),.clk(gclk));
	jdff dff_A_wlNhtr8z1_0(.dout(w_dff_A_4ixODqpk9_0),.din(w_dff_A_wlNhtr8z1_0),.clk(gclk));
	jdff dff_A_4ixODqpk9_0(.dout(w_dff_A_j3eFymXy2_0),.din(w_dff_A_4ixODqpk9_0),.clk(gclk));
	jdff dff_A_j3eFymXy2_0(.dout(w_dff_A_Z2ZM1x5n9_0),.din(w_dff_A_j3eFymXy2_0),.clk(gclk));
	jdff dff_A_Z2ZM1x5n9_0(.dout(w_dff_A_okzo6YL03_0),.din(w_dff_A_Z2ZM1x5n9_0),.clk(gclk));
	jdff dff_A_okzo6YL03_0(.dout(w_dff_A_bM3xybTO2_0),.din(w_dff_A_okzo6YL03_0),.clk(gclk));
	jdff dff_A_bM3xybTO2_0(.dout(G867),.din(w_dff_A_bM3xybTO2_0),.clk(gclk));
	jdff dff_A_j23ZqMUB9_1(.dout(w_dff_A_BripIcQc4_0),.din(w_dff_A_j23ZqMUB9_1),.clk(gclk));
	jdff dff_A_BripIcQc4_0(.dout(w_dff_A_nkxwIEI26_0),.din(w_dff_A_BripIcQc4_0),.clk(gclk));
	jdff dff_A_nkxwIEI26_0(.dout(w_dff_A_7thvBMRw5_0),.din(w_dff_A_nkxwIEI26_0),.clk(gclk));
	jdff dff_A_7thvBMRw5_0(.dout(w_dff_A_W4DvVmCP1_0),.din(w_dff_A_7thvBMRw5_0),.clk(gclk));
	jdff dff_A_W4DvVmCP1_0(.dout(w_dff_A_Eda2cVrQ1_0),.din(w_dff_A_W4DvVmCP1_0),.clk(gclk));
	jdff dff_A_Eda2cVrQ1_0(.dout(w_dff_A_raUYjNWG4_0),.din(w_dff_A_Eda2cVrQ1_0),.clk(gclk));
	jdff dff_A_raUYjNWG4_0(.dout(w_dff_A_NscxkqwB6_0),.din(w_dff_A_raUYjNWG4_0),.clk(gclk));
	jdff dff_A_NscxkqwB6_0(.dout(w_dff_A_Qz1Vf87J9_0),.din(w_dff_A_NscxkqwB6_0),.clk(gclk));
	jdff dff_A_Qz1Vf87J9_0(.dout(w_dff_A_0lvFX9Rn9_0),.din(w_dff_A_Qz1Vf87J9_0),.clk(gclk));
	jdff dff_A_0lvFX9Rn9_0(.dout(G869),.din(w_dff_A_0lvFX9Rn9_0),.clk(gclk));
	jdff dff_A_2XGOUCxJ2_2(.dout(w_dff_A_L4YhNQt45_0),.din(w_dff_A_2XGOUCxJ2_2),.clk(gclk));
	jdff dff_A_L4YhNQt45_0(.dout(w_dff_A_LZr3Dsus0_0),.din(w_dff_A_L4YhNQt45_0),.clk(gclk));
	jdff dff_A_LZr3Dsus0_0(.dout(w_dff_A_23BSm3Fp3_0),.din(w_dff_A_LZr3Dsus0_0),.clk(gclk));
	jdff dff_A_23BSm3Fp3_0(.dout(G712),.din(w_dff_A_23BSm3Fp3_0),.clk(gclk));
	jdff dff_A_fDdSOlMD0_2(.dout(w_dff_A_SN76x4gC2_0),.din(w_dff_A_fDdSOlMD0_2),.clk(gclk));
	jdff dff_A_SN76x4gC2_0(.dout(w_dff_A_iJYymryz2_0),.din(w_dff_A_SN76x4gC2_0),.clk(gclk));
	jdff dff_A_iJYymryz2_0(.dout(G727),.din(w_dff_A_iJYymryz2_0),.clk(gclk));
	jdff dff_A_5eIRg5hX3_2(.dout(w_dff_A_aaW5Ixtd9_0),.din(w_dff_A_5eIRg5hX3_2),.clk(gclk));
	jdff dff_A_aaW5Ixtd9_0(.dout(w_dff_A_jYli0LbD5_0),.din(w_dff_A_aaW5Ixtd9_0),.clk(gclk));
	jdff dff_A_jYli0LbD5_0(.dout(w_dff_A_82A8IQ7J9_0),.din(w_dff_A_jYli0LbD5_0),.clk(gclk));
	jdff dff_A_82A8IQ7J9_0(.dout(G732),.din(w_dff_A_82A8IQ7J9_0),.clk(gclk));
	jdff dff_A_sYyisCNw9_2(.dout(w_dff_A_uwf4jsWY1_0),.din(w_dff_A_sYyisCNw9_2),.clk(gclk));
	jdff dff_A_uwf4jsWY1_0(.dout(w_dff_A_fvUwqR9F9_0),.din(w_dff_A_uwf4jsWY1_0),.clk(gclk));
	jdff dff_A_fvUwqR9F9_0(.dout(w_dff_A_igVS6zOD9_0),.din(w_dff_A_fvUwqR9F9_0),.clk(gclk));
	jdff dff_A_igVS6zOD9_0(.dout(G737),.din(w_dff_A_igVS6zOD9_0),.clk(gclk));
	jdff dff_A_jLaVIWAZ5_2(.dout(w_dff_A_zobrglLG5_0),.din(w_dff_A_jLaVIWAZ5_2),.clk(gclk));
	jdff dff_A_zobrglLG5_0(.dout(w_dff_A_8BKcmYGu9_0),.din(w_dff_A_zobrglLG5_0),.clk(gclk));
	jdff dff_A_8BKcmYGu9_0(.dout(w_dff_A_CRzGPY5k9_0),.din(w_dff_A_8BKcmYGu9_0),.clk(gclk));
	jdff dff_A_CRzGPY5k9_0(.dout(w_dff_A_fMd2qyrI0_0),.din(w_dff_A_CRzGPY5k9_0),.clk(gclk));
	jdff dff_A_fMd2qyrI0_0(.dout(G742),.din(w_dff_A_fMd2qyrI0_0),.clk(gclk));
	jdff dff_A_jHQxUsEJ2_2(.dout(w_dff_A_VJVUz5976_0),.din(w_dff_A_jHQxUsEJ2_2),.clk(gclk));
	jdff dff_A_VJVUz5976_0(.dout(w_dff_A_QSIPoHGe8_0),.din(w_dff_A_VJVUz5976_0),.clk(gclk));
	jdff dff_A_QSIPoHGe8_0(.dout(w_dff_A_W8Hw7NkO9_0),.din(w_dff_A_QSIPoHGe8_0),.clk(gclk));
	jdff dff_A_W8Hw7NkO9_0(.dout(G772),.din(w_dff_A_W8Hw7NkO9_0),.clk(gclk));
	jdff dff_A_nrcvRrKO0_2(.dout(w_dff_A_T2CRHUaN5_0),.din(w_dff_A_nrcvRrKO0_2),.clk(gclk));
	jdff dff_A_T2CRHUaN5_0(.dout(w_dff_A_CRb5XH6s3_0),.din(w_dff_A_T2CRHUaN5_0),.clk(gclk));
	jdff dff_A_CRb5XH6s3_0(.dout(w_dff_A_BeeoD6W52_0),.din(w_dff_A_CRb5XH6s3_0),.clk(gclk));
	jdff dff_A_BeeoD6W52_0(.dout(G777),.din(w_dff_A_BeeoD6W52_0),.clk(gclk));
	jdff dff_A_7DtcfDVl6_2(.dout(w_dff_A_SpizzXDb1_0),.din(w_dff_A_7DtcfDVl6_2),.clk(gclk));
	jdff dff_A_SpizzXDb1_0(.dout(w_dff_A_9Ei9FrSA4_0),.din(w_dff_A_SpizzXDb1_0),.clk(gclk));
	jdff dff_A_9Ei9FrSA4_0(.dout(w_dff_A_uoq4p2iG1_0),.din(w_dff_A_9Ei9FrSA4_0),.clk(gclk));
	jdff dff_A_uoq4p2iG1_0(.dout(w_dff_A_G8XakyhD1_0),.din(w_dff_A_uoq4p2iG1_0),.clk(gclk));
	jdff dff_A_G8XakyhD1_0(.dout(G782),.din(w_dff_A_G8XakyhD1_0),.clk(gclk));
	jdff dff_A_P32bXcZR1_2(.dout(w_dff_A_zJ9g5eMu7_0),.din(w_dff_A_P32bXcZR1_2),.clk(gclk));
	jdff dff_A_zJ9g5eMu7_0(.dout(w_dff_A_49XX6y1L1_0),.din(w_dff_A_zJ9g5eMu7_0),.clk(gclk));
	jdff dff_A_49XX6y1L1_0(.dout(w_dff_A_nB1rVZ1i2_0),.din(w_dff_A_49XX6y1L1_0),.clk(gclk));
	jdff dff_A_nB1rVZ1i2_0(.dout(G645),.din(w_dff_A_nB1rVZ1i2_0),.clk(gclk));
	jdff dff_A_7lXH9BOj8_2(.dout(w_dff_A_O2WopYZH8_0),.din(w_dff_A_7lXH9BOj8_2),.clk(gclk));
	jdff dff_A_O2WopYZH8_0(.dout(w_dff_A_BTztYjhw3_0),.din(w_dff_A_O2WopYZH8_0),.clk(gclk));
	jdff dff_A_BTztYjhw3_0(.dout(G648),.din(w_dff_A_BTztYjhw3_0),.clk(gclk));
	jdff dff_A_6ondWxNN6_2(.dout(w_dff_A_RJ2UJ6Ua3_0),.din(w_dff_A_6ondWxNN6_2),.clk(gclk));
	jdff dff_A_RJ2UJ6Ua3_0(.dout(w_dff_A_SmIMZAQG8_0),.din(w_dff_A_RJ2UJ6Ua3_0),.clk(gclk));
	jdff dff_A_SmIMZAQG8_0(.dout(G651),.din(w_dff_A_SmIMZAQG8_0),.clk(gclk));
	jdff dff_A_EW50mF6G8_2(.dout(w_dff_A_ToC18BX84_0),.din(w_dff_A_EW50mF6G8_2),.clk(gclk));
	jdff dff_A_ToC18BX84_0(.dout(G654),.din(w_dff_A_ToC18BX84_0),.clk(gclk));
	jdff dff_A_qtIVFaz20_2(.dout(w_dff_A_sohk3fe49_0),.din(w_dff_A_qtIVFaz20_2),.clk(gclk));
	jdff dff_A_sohk3fe49_0(.dout(w_dff_A_DL8HlS531_0),.din(w_dff_A_sohk3fe49_0),.clk(gclk));
	jdff dff_A_DL8HlS531_0(.dout(w_dff_A_Y83qaQXm3_0),.din(w_dff_A_DL8HlS531_0),.clk(gclk));
	jdff dff_A_Y83qaQXm3_0(.dout(G679),.din(w_dff_A_Y83qaQXm3_0),.clk(gclk));
	jdff dff_A_SZppPzwU8_2(.dout(w_dff_A_KWQ3KdOQ2_0),.din(w_dff_A_SZppPzwU8_2),.clk(gclk));
	jdff dff_A_KWQ3KdOQ2_0(.dout(w_dff_A_DduDY9mV2_0),.din(w_dff_A_KWQ3KdOQ2_0),.clk(gclk));
	jdff dff_A_DduDY9mV2_0(.dout(G682),.din(w_dff_A_DduDY9mV2_0),.clk(gclk));
	jdff dff_A_EjeCPIAX3_2(.dout(w_dff_A_lSRPRseG4_0),.din(w_dff_A_EjeCPIAX3_2),.clk(gclk));
	jdff dff_A_lSRPRseG4_0(.dout(w_dff_A_wmPkw9R00_0),.din(w_dff_A_lSRPRseG4_0),.clk(gclk));
	jdff dff_A_wmPkw9R00_0(.dout(G685),.din(w_dff_A_wmPkw9R00_0),.clk(gclk));
	jdff dff_A_NyJ1LQKr6_2(.dout(w_dff_A_J5tMnEw31_0),.din(w_dff_A_NyJ1LQKr6_2),.clk(gclk));
	jdff dff_A_J5tMnEw31_0(.dout(w_dff_A_s8pDORCC1_0),.din(w_dff_A_J5tMnEw31_0),.clk(gclk));
	jdff dff_A_s8pDORCC1_0(.dout(G688),.din(w_dff_A_s8pDORCC1_0),.clk(gclk));
	jdff dff_A_VYoWKH9V5_2(.dout(w_dff_A_iQeJaTKS7_0),.din(w_dff_A_VYoWKH9V5_2),.clk(gclk));
	jdff dff_A_iQeJaTKS7_0(.dout(w_dff_A_pjJjMj0F8_0),.din(w_dff_A_iQeJaTKS7_0),.clk(gclk));
	jdff dff_A_pjJjMj0F8_0(.dout(w_dff_A_Sd2CgZtn5_0),.din(w_dff_A_pjJjMj0F8_0),.clk(gclk));
	jdff dff_A_Sd2CgZtn5_0(.dout(w_dff_A_PUbC0Vfa6_0),.din(w_dff_A_Sd2CgZtn5_0),.clk(gclk));
	jdff dff_A_PUbC0Vfa6_0(.dout(w_dff_A_uX9slJXe3_0),.din(w_dff_A_PUbC0Vfa6_0),.clk(gclk));
	jdff dff_A_uX9slJXe3_0(.dout(G843),.din(w_dff_A_uX9slJXe3_0),.clk(gclk));
	jdff dff_A_6B9aVpnN0_2(.dout(w_dff_A_ZMGT75uD3_0),.din(w_dff_A_6B9aVpnN0_2),.clk(gclk));
	jdff dff_A_ZMGT75uD3_0(.dout(w_dff_A_C32bfpmL1_0),.din(w_dff_A_ZMGT75uD3_0),.clk(gclk));
	jdff dff_A_C32bfpmL1_0(.dout(w_dff_A_jHkqsqtz0_0),.din(w_dff_A_C32bfpmL1_0),.clk(gclk));
	jdff dff_A_jHkqsqtz0_0(.dout(w_dff_A_gPiOw7G95_0),.din(w_dff_A_jHkqsqtz0_0),.clk(gclk));
	jdff dff_A_gPiOw7G95_0(.dout(w_dff_A_cscWtQnO0_0),.din(w_dff_A_gPiOw7G95_0),.clk(gclk));
	jdff dff_A_cscWtQnO0_0(.dout(G882),.din(w_dff_A_cscWtQnO0_0),.clk(gclk));
	jdff dff_A_xjst1swX1_2(.dout(G767),.din(w_dff_A_xjst1swX1_2),.clk(gclk));
	jdff dff_A_73jqJqeU4_2(.dout(G807),.din(w_dff_A_73jqJqeU4_2),.clk(gclk));
endmodule

