/*
gf_bar:
	jspl: 655
	jspl3: 1145
	jnot: 7
	jdff: 1244
	jand: 1478
	jor: 1474

Summary:
	jspl: 655
	jspl3: 1145
	jnot: 7
	jdff: 1244
	jand: 1478
	jor: 1474

The maximum logic level gap of any gate:
	gf_bar: 13
*/

module gf_bar(gclk, a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28, a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42, a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56, a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70, a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84, a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98, a99, a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110, a111, a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122, a123, a124, a125, a126, a127, shift0, shift1, shift2, shift3, shift4, shift5, shift6, result0, result1, result2, result3, result4, result5, result6, result7, result8, result9, result10, result11, result12, result13, result14, result15, result16, result17, result18, result19, result20, result21, result22, result23, result24, result25, result26, result27, result28, result29, result30, result31, result32, result33, result34, result35, result36, result37, result38, result39, result40, result41, result42, result43, result44, result45, result46, result47, result48, result49, result50, result51, result52, result53, result54, result55, result56, result57, result58, result59, result60, result61, result62, result63, result64, result65, result66, result67, result68, result69, result70, result71, result72, result73, result74, result75, result76, result77, result78, result79, result80, result81, result82, result83, result84, result85, result86, result87, result88, result89, result90, result91, result92, result93, result94, result95, result96, result97, result98, result99, result100, result101, result102, result103, result104, result105, result106, result107, result108, result109, result110, result111, result112, result113, result114, result115, result116, result117, result118, result119, result120, result121, result122, result123, result124, result125, result126, result127);
	input gclk;
	input a0;
	input a1;
	input a2;
	input a3;
	input a4;
	input a5;
	input a6;
	input a7;
	input a8;
	input a9;
	input a10;
	input a11;
	input a12;
	input a13;
	input a14;
	input a15;
	input a16;
	input a17;
	input a18;
	input a19;
	input a20;
	input a21;
	input a22;
	input a23;
	input a24;
	input a25;
	input a26;
	input a27;
	input a28;
	input a29;
	input a30;
	input a31;
	input a32;
	input a33;
	input a34;
	input a35;
	input a36;
	input a37;
	input a38;
	input a39;
	input a40;
	input a41;
	input a42;
	input a43;
	input a44;
	input a45;
	input a46;
	input a47;
	input a48;
	input a49;
	input a50;
	input a51;
	input a52;
	input a53;
	input a54;
	input a55;
	input a56;
	input a57;
	input a58;
	input a59;
	input a60;
	input a61;
	input a62;
	input a63;
	input a64;
	input a65;
	input a66;
	input a67;
	input a68;
	input a69;
	input a70;
	input a71;
	input a72;
	input a73;
	input a74;
	input a75;
	input a76;
	input a77;
	input a78;
	input a79;
	input a80;
	input a81;
	input a82;
	input a83;
	input a84;
	input a85;
	input a86;
	input a87;
	input a88;
	input a89;
	input a90;
	input a91;
	input a92;
	input a93;
	input a94;
	input a95;
	input a96;
	input a97;
	input a98;
	input a99;
	input a100;
	input a101;
	input a102;
	input a103;
	input a104;
	input a105;
	input a106;
	input a107;
	input a108;
	input a109;
	input a110;
	input a111;
	input a112;
	input a113;
	input a114;
	input a115;
	input a116;
	input a117;
	input a118;
	input a119;
	input a120;
	input a121;
	input a122;
	input a123;
	input a124;
	input a125;
	input a126;
	input a127;
	input shift0;
	input shift1;
	input shift2;
	input shift3;
	input shift4;
	input shift5;
	input shift6;
	output result0;
	output result1;
	output result2;
	output result3;
	output result4;
	output result5;
	output result6;
	output result7;
	output result8;
	output result9;
	output result10;
	output result11;
	output result12;
	output result13;
	output result14;
	output result15;
	output result16;
	output result17;
	output result18;
	output result19;
	output result20;
	output result21;
	output result22;
	output result23;
	output result24;
	output result25;
	output result26;
	output result27;
	output result28;
	output result29;
	output result30;
	output result31;
	output result32;
	output result33;
	output result34;
	output result35;
	output result36;
	output result37;
	output result38;
	output result39;
	output result40;
	output result41;
	output result42;
	output result43;
	output result44;
	output result45;
	output result46;
	output result47;
	output result48;
	output result49;
	output result50;
	output result51;
	output result52;
	output result53;
	output result54;
	output result55;
	output result56;
	output result57;
	output result58;
	output result59;
	output result60;
	output result61;
	output result62;
	output result63;
	output result64;
	output result65;
	output result66;
	output result67;
	output result68;
	output result69;
	output result70;
	output result71;
	output result72;
	output result73;
	output result74;
	output result75;
	output result76;
	output result77;
	output result78;
	output result79;
	output result80;
	output result81;
	output result82;
	output result83;
	output result84;
	output result85;
	output result86;
	output result87;
	output result88;
	output result89;
	output result90;
	output result91;
	output result92;
	output result93;
	output result94;
	output result95;
	output result96;
	output result97;
	output result98;
	output result99;
	output result100;
	output result101;
	output result102;
	output result103;
	output result104;
	output result105;
	output result106;
	output result107;
	output result108;
	output result109;
	output result110;
	output result111;
	output result112;
	output result113;
	output result114;
	output result115;
	output result116;
	output result117;
	output result118;
	output result119;
	output result120;
	output result121;
	output result122;
	output result123;
	output result124;
	output result125;
	output result126;
	output result127;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1837;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1849;
	wire n1850;
	wire n1851;
	wire n1852;
	wire n1853;
	wire n1854;
	wire n1855;
	wire n1856;
	wire n1857;
	wire n1858;
	wire n1859;
	wire n1860;
	wire n1861;
	wire n1862;
	wire n1863;
	wire n1864;
	wire n1865;
	wire n1866;
	wire n1867;
	wire n1868;
	wire n1869;
	wire n1870;
	wire n1871;
	wire n1872;
	wire n1873;
	wire n1874;
	wire n1875;
	wire n1876;
	wire n1877;
	wire n1878;
	wire n1879;
	wire n1880;
	wire n1881;
	wire n1882;
	wire n1883;
	wire n1884;
	wire n1885;
	wire n1886;
	wire n1887;
	wire n1888;
	wire n1889;
	wire n1890;
	wire n1891;
	wire n1892;
	wire n1893;
	wire n1894;
	wire n1895;
	wire n1896;
	wire n1897;
	wire n1898;
	wire n1899;
	wire n1900;
	wire n1901;
	wire n1902;
	wire n1903;
	wire n1904;
	wire n1905;
	wire n1906;
	wire n1907;
	wire n1908;
	wire n1909;
	wire n1910;
	wire n1911;
	wire n1912;
	wire n1913;
	wire n1914;
	wire n1915;
	wire n1916;
	wire n1917;
	wire n1918;
	wire n1919;
	wire n1920;
	wire n1922;
	wire n1923;
	wire n1924;
	wire n1925;
	wire n1926;
	wire n1927;
	wire n1928;
	wire n1929;
	wire n1930;
	wire n1931;
	wire n1932;
	wire n1933;
	wire n1934;
	wire n1935;
	wire n1936;
	wire n1937;
	wire n1938;
	wire n1939;
	wire n1940;
	wire n1941;
	wire n1942;
	wire n1943;
	wire n1944;
	wire n1945;
	wire n1946;
	wire n1947;
	wire n1948;
	wire n1949;
	wire n1950;
	wire n1951;
	wire n1952;
	wire n1953;
	wire n1954;
	wire n1955;
	wire n1956;
	wire n1957;
	wire n1958;
	wire n1959;
	wire n1960;
	wire n1961;
	wire n1962;
	wire n1963;
	wire n1964;
	wire n1965;
	wire n1966;
	wire n1967;
	wire n1968;
	wire n1969;
	wire n1970;
	wire n1971;
	wire n1972;
	wire n1973;
	wire n1974;
	wire n1975;
	wire n1976;
	wire n1977;
	wire n1978;
	wire n1979;
	wire n1980;
	wire n1981;
	wire n1982;
	wire n1983;
	wire n1984;
	wire n1985;
	wire n1986;
	wire n1987;
	wire n1988;
	wire n1989;
	wire n1990;
	wire n1991;
	wire n1992;
	wire n1993;
	wire n1995;
	wire n1996;
	wire n1997;
	wire n1998;
	wire n1999;
	wire n2000;
	wire n2001;
	wire n2002;
	wire n2003;
	wire n2004;
	wire n2005;
	wire n2006;
	wire n2007;
	wire n2008;
	wire n2009;
	wire n2010;
	wire n2011;
	wire n2012;
	wire n2013;
	wire n2014;
	wire n2015;
	wire n2016;
	wire n2017;
	wire n2018;
	wire n2019;
	wire n2020;
	wire n2021;
	wire n2022;
	wire n2023;
	wire n2024;
	wire n2025;
	wire n2026;
	wire n2027;
	wire n2028;
	wire n2029;
	wire n2030;
	wire n2031;
	wire n2032;
	wire n2033;
	wire n2034;
	wire n2035;
	wire n2036;
	wire n2037;
	wire n2038;
	wire n2039;
	wire n2040;
	wire n2041;
	wire n2042;
	wire n2043;
	wire n2044;
	wire n2045;
	wire n2046;
	wire n2047;
	wire n2048;
	wire n2049;
	wire n2050;
	wire n2051;
	wire n2052;
	wire n2053;
	wire n2054;
	wire n2055;
	wire n2056;
	wire n2057;
	wire n2058;
	wire n2059;
	wire n2060;
	wire n2061;
	wire n2062;
	wire n2063;
	wire n2064;
	wire n2065;
	wire n2066;
	wire n2068;
	wire n2069;
	wire n2070;
	wire n2071;
	wire n2072;
	wire n2073;
	wire n2074;
	wire n2075;
	wire n2076;
	wire n2077;
	wire n2078;
	wire n2079;
	wire n2080;
	wire n2081;
	wire n2082;
	wire n2083;
	wire n2084;
	wire n2085;
	wire n2086;
	wire n2087;
	wire n2088;
	wire n2089;
	wire n2090;
	wire n2091;
	wire n2092;
	wire n2093;
	wire n2094;
	wire n2095;
	wire n2096;
	wire n2097;
	wire n2098;
	wire n2099;
	wire n2100;
	wire n2101;
	wire n2102;
	wire n2103;
	wire n2104;
	wire n2105;
	wire n2106;
	wire n2107;
	wire n2108;
	wire n2109;
	wire n2110;
	wire n2111;
	wire n2112;
	wire n2113;
	wire n2114;
	wire n2115;
	wire n2116;
	wire n2117;
	wire n2118;
	wire n2119;
	wire n2120;
	wire n2121;
	wire n2122;
	wire n2123;
	wire n2124;
	wire n2125;
	wire n2126;
	wire n2127;
	wire n2128;
	wire n2129;
	wire n2130;
	wire n2131;
	wire n2132;
	wire n2133;
	wire n2134;
	wire n2135;
	wire n2136;
	wire n2137;
	wire n2138;
	wire n2139;
	wire n2141;
	wire n2142;
	wire n2143;
	wire n2144;
	wire n2145;
	wire n2146;
	wire n2147;
	wire n2148;
	wire n2149;
	wire n2150;
	wire n2151;
	wire n2152;
	wire n2153;
	wire n2154;
	wire n2155;
	wire n2156;
	wire n2157;
	wire n2158;
	wire n2159;
	wire n2160;
	wire n2161;
	wire n2162;
	wire n2163;
	wire n2164;
	wire n2165;
	wire n2166;
	wire n2167;
	wire n2168;
	wire n2169;
	wire n2170;
	wire n2171;
	wire n2172;
	wire n2173;
	wire n2174;
	wire n2175;
	wire n2176;
	wire n2177;
	wire n2178;
	wire n2179;
	wire n2180;
	wire n2181;
	wire n2182;
	wire n2183;
	wire n2184;
	wire n2185;
	wire n2186;
	wire n2187;
	wire n2188;
	wire n2189;
	wire n2190;
	wire n2191;
	wire n2192;
	wire n2193;
	wire n2194;
	wire n2195;
	wire n2196;
	wire n2197;
	wire n2198;
	wire n2199;
	wire n2200;
	wire n2201;
	wire n2202;
	wire n2203;
	wire n2204;
	wire n2205;
	wire n2206;
	wire n2207;
	wire n2208;
	wire n2209;
	wire n2210;
	wire n2211;
	wire n2212;
	wire n2214;
	wire n2215;
	wire n2216;
	wire n2217;
	wire n2218;
	wire n2219;
	wire n2220;
	wire n2221;
	wire n2222;
	wire n2223;
	wire n2224;
	wire n2225;
	wire n2226;
	wire n2227;
	wire n2228;
	wire n2229;
	wire n2231;
	wire n2232;
	wire n2233;
	wire n2234;
	wire n2235;
	wire n2236;
	wire n2237;
	wire n2238;
	wire n2239;
	wire n2240;
	wire n2241;
	wire n2242;
	wire n2243;
	wire n2244;
	wire n2245;
	wire n2246;
	wire n2248;
	wire n2249;
	wire n2250;
	wire n2251;
	wire n2252;
	wire n2253;
	wire n2254;
	wire n2255;
	wire n2256;
	wire n2257;
	wire n2258;
	wire n2259;
	wire n2260;
	wire n2261;
	wire n2262;
	wire n2263;
	wire n2265;
	wire n2266;
	wire n2267;
	wire n2268;
	wire n2269;
	wire n2270;
	wire n2271;
	wire n2272;
	wire n2273;
	wire n2274;
	wire n2275;
	wire n2276;
	wire n2277;
	wire n2278;
	wire n2279;
	wire n2280;
	wire n2282;
	wire n2283;
	wire n2284;
	wire n2285;
	wire n2286;
	wire n2287;
	wire n2288;
	wire n2289;
	wire n2290;
	wire n2291;
	wire n2292;
	wire n2293;
	wire n2294;
	wire n2295;
	wire n2296;
	wire n2297;
	wire n2299;
	wire n2300;
	wire n2301;
	wire n2302;
	wire n2303;
	wire n2304;
	wire n2305;
	wire n2306;
	wire n2307;
	wire n2308;
	wire n2309;
	wire n2310;
	wire n2311;
	wire n2312;
	wire n2313;
	wire n2314;
	wire n2316;
	wire n2317;
	wire n2318;
	wire n2319;
	wire n2320;
	wire n2321;
	wire n2322;
	wire n2323;
	wire n2324;
	wire n2325;
	wire n2326;
	wire n2327;
	wire n2328;
	wire n2329;
	wire n2330;
	wire n2331;
	wire n2333;
	wire n2334;
	wire n2335;
	wire n2336;
	wire n2337;
	wire n2338;
	wire n2339;
	wire n2340;
	wire n2341;
	wire n2342;
	wire n2343;
	wire n2344;
	wire n2345;
	wire n2346;
	wire n2347;
	wire n2348;
	wire n2350;
	wire n2351;
	wire n2352;
	wire n2353;
	wire n2354;
	wire n2355;
	wire n2356;
	wire n2357;
	wire n2358;
	wire n2359;
	wire n2360;
	wire n2361;
	wire n2362;
	wire n2363;
	wire n2364;
	wire n2365;
	wire n2367;
	wire n2368;
	wire n2369;
	wire n2370;
	wire n2371;
	wire n2372;
	wire n2373;
	wire n2374;
	wire n2375;
	wire n2376;
	wire n2377;
	wire n2378;
	wire n2379;
	wire n2380;
	wire n2381;
	wire n2382;
	wire n2384;
	wire n2385;
	wire n2386;
	wire n2387;
	wire n2388;
	wire n2389;
	wire n2390;
	wire n2391;
	wire n2392;
	wire n2393;
	wire n2394;
	wire n2395;
	wire n2396;
	wire n2397;
	wire n2398;
	wire n2399;
	wire n2401;
	wire n2402;
	wire n2403;
	wire n2404;
	wire n2405;
	wire n2406;
	wire n2407;
	wire n2408;
	wire n2409;
	wire n2410;
	wire n2411;
	wire n2412;
	wire n2413;
	wire n2414;
	wire n2415;
	wire n2416;
	wire n2418;
	wire n2419;
	wire n2420;
	wire n2421;
	wire n2422;
	wire n2423;
	wire n2424;
	wire n2425;
	wire n2426;
	wire n2427;
	wire n2428;
	wire n2429;
	wire n2430;
	wire n2431;
	wire n2432;
	wire n2433;
	wire n2435;
	wire n2436;
	wire n2437;
	wire n2438;
	wire n2439;
	wire n2440;
	wire n2441;
	wire n2442;
	wire n2443;
	wire n2444;
	wire n2445;
	wire n2446;
	wire n2447;
	wire n2448;
	wire n2449;
	wire n2450;
	wire n2452;
	wire n2453;
	wire n2454;
	wire n2455;
	wire n2456;
	wire n2457;
	wire n2458;
	wire n2459;
	wire n2460;
	wire n2461;
	wire n2462;
	wire n2463;
	wire n2464;
	wire n2465;
	wire n2466;
	wire n2467;
	wire n2469;
	wire n2470;
	wire n2471;
	wire n2472;
	wire n2473;
	wire n2474;
	wire n2475;
	wire n2476;
	wire n2477;
	wire n2478;
	wire n2479;
	wire n2480;
	wire n2481;
	wire n2482;
	wire n2483;
	wire n2484;
	wire n2486;
	wire n2487;
	wire n2488;
	wire n2489;
	wire n2490;
	wire n2491;
	wire n2492;
	wire n2493;
	wire n2494;
	wire n2495;
	wire n2496;
	wire n2497;
	wire n2498;
	wire n2499;
	wire n2500;
	wire n2501;
	wire n2503;
	wire n2504;
	wire n2505;
	wire n2506;
	wire n2507;
	wire n2508;
	wire n2509;
	wire n2510;
	wire n2511;
	wire n2512;
	wire n2513;
	wire n2514;
	wire n2515;
	wire n2516;
	wire n2517;
	wire n2518;
	wire n2520;
	wire n2521;
	wire n2522;
	wire n2523;
	wire n2524;
	wire n2525;
	wire n2526;
	wire n2527;
	wire n2528;
	wire n2529;
	wire n2530;
	wire n2531;
	wire n2532;
	wire n2533;
	wire n2534;
	wire n2535;
	wire n2537;
	wire n2538;
	wire n2539;
	wire n2540;
	wire n2541;
	wire n2542;
	wire n2543;
	wire n2544;
	wire n2545;
	wire n2546;
	wire n2547;
	wire n2548;
	wire n2549;
	wire n2550;
	wire n2551;
	wire n2552;
	wire n2554;
	wire n2555;
	wire n2556;
	wire n2557;
	wire n2558;
	wire n2559;
	wire n2560;
	wire n2561;
	wire n2562;
	wire n2563;
	wire n2564;
	wire n2565;
	wire n2566;
	wire n2567;
	wire n2568;
	wire n2569;
	wire n2571;
	wire n2572;
	wire n2573;
	wire n2574;
	wire n2575;
	wire n2576;
	wire n2577;
	wire n2578;
	wire n2579;
	wire n2580;
	wire n2581;
	wire n2582;
	wire n2583;
	wire n2584;
	wire n2585;
	wire n2586;
	wire n2588;
	wire n2589;
	wire n2590;
	wire n2591;
	wire n2592;
	wire n2593;
	wire n2594;
	wire n2595;
	wire n2596;
	wire n2597;
	wire n2598;
	wire n2599;
	wire n2600;
	wire n2601;
	wire n2602;
	wire n2603;
	wire n2605;
	wire n2606;
	wire n2607;
	wire n2608;
	wire n2609;
	wire n2610;
	wire n2611;
	wire n2612;
	wire n2613;
	wire n2614;
	wire n2615;
	wire n2616;
	wire n2617;
	wire n2618;
	wire n2619;
	wire n2620;
	wire n2622;
	wire n2623;
	wire n2624;
	wire n2625;
	wire n2626;
	wire n2627;
	wire n2628;
	wire n2629;
	wire n2630;
	wire n2631;
	wire n2632;
	wire n2633;
	wire n2634;
	wire n2635;
	wire n2636;
	wire n2637;
	wire n2639;
	wire n2640;
	wire n2641;
	wire n2642;
	wire n2643;
	wire n2644;
	wire n2645;
	wire n2646;
	wire n2647;
	wire n2648;
	wire n2649;
	wire n2650;
	wire n2651;
	wire n2652;
	wire n2653;
	wire n2654;
	wire n2656;
	wire n2657;
	wire n2658;
	wire n2659;
	wire n2660;
	wire n2661;
	wire n2662;
	wire n2663;
	wire n2664;
	wire n2665;
	wire n2666;
	wire n2667;
	wire n2668;
	wire n2669;
	wire n2670;
	wire n2671;
	wire n2673;
	wire n2674;
	wire n2675;
	wire n2676;
	wire n2677;
	wire n2678;
	wire n2679;
	wire n2680;
	wire n2681;
	wire n2682;
	wire n2683;
	wire n2684;
	wire n2685;
	wire n2686;
	wire n2687;
	wire n2688;
	wire n2690;
	wire n2691;
	wire n2692;
	wire n2693;
	wire n2694;
	wire n2695;
	wire n2696;
	wire n2697;
	wire n2698;
	wire n2699;
	wire n2700;
	wire n2701;
	wire n2702;
	wire n2703;
	wire n2704;
	wire n2705;
	wire n2707;
	wire n2708;
	wire n2709;
	wire n2710;
	wire n2711;
	wire n2712;
	wire n2713;
	wire n2714;
	wire n2715;
	wire n2716;
	wire n2717;
	wire n2718;
	wire n2719;
	wire n2720;
	wire n2721;
	wire n2722;
	wire n2724;
	wire n2725;
	wire n2726;
	wire n2727;
	wire n2728;
	wire n2729;
	wire n2730;
	wire n2731;
	wire n2732;
	wire n2733;
	wire n2734;
	wire n2735;
	wire n2736;
	wire n2737;
	wire n2738;
	wire n2739;
	wire n2741;
	wire n2742;
	wire n2743;
	wire n2744;
	wire n2745;
	wire n2746;
	wire n2747;
	wire n2748;
	wire n2749;
	wire n2750;
	wire n2751;
	wire n2752;
	wire n2753;
	wire n2754;
	wire n2755;
	wire n2756;
	wire n2758;
	wire n2759;
	wire n2760;
	wire n2761;
	wire n2762;
	wire n2763;
	wire n2764;
	wire n2765;
	wire n2766;
	wire n2767;
	wire n2768;
	wire n2769;
	wire n2770;
	wire n2771;
	wire n2772;
	wire n2773;
	wire n2775;
	wire n2776;
	wire n2777;
	wire n2778;
	wire n2779;
	wire n2780;
	wire n2781;
	wire n2782;
	wire n2783;
	wire n2784;
	wire n2785;
	wire n2786;
	wire n2787;
	wire n2788;
	wire n2789;
	wire n2790;
	wire n2792;
	wire n2793;
	wire n2794;
	wire n2795;
	wire n2796;
	wire n2797;
	wire n2798;
	wire n2799;
	wire n2800;
	wire n2801;
	wire n2802;
	wire n2803;
	wire n2804;
	wire n2805;
	wire n2806;
	wire n2807;
	wire n2809;
	wire n2810;
	wire n2811;
	wire n2812;
	wire n2813;
	wire n2814;
	wire n2815;
	wire n2816;
	wire n2817;
	wire n2818;
	wire n2819;
	wire n2820;
	wire n2821;
	wire n2822;
	wire n2823;
	wire n2824;
	wire n2826;
	wire n2827;
	wire n2828;
	wire n2829;
	wire n2830;
	wire n2831;
	wire n2832;
	wire n2833;
	wire n2834;
	wire n2835;
	wire n2836;
	wire n2837;
	wire n2838;
	wire n2839;
	wire n2840;
	wire n2841;
	wire n2843;
	wire n2844;
	wire n2845;
	wire n2846;
	wire n2847;
	wire n2848;
	wire n2849;
	wire n2850;
	wire n2851;
	wire n2852;
	wire n2853;
	wire n2854;
	wire n2855;
	wire n2856;
	wire n2857;
	wire n2858;
	wire n2860;
	wire n2861;
	wire n2862;
	wire n2863;
	wire n2864;
	wire n2865;
	wire n2866;
	wire n2867;
	wire n2868;
	wire n2869;
	wire n2870;
	wire n2871;
	wire n2872;
	wire n2873;
	wire n2874;
	wire n2875;
	wire n2877;
	wire n2878;
	wire n2879;
	wire n2880;
	wire n2881;
	wire n2882;
	wire n2883;
	wire n2884;
	wire n2885;
	wire n2886;
	wire n2887;
	wire n2888;
	wire n2889;
	wire n2890;
	wire n2891;
	wire n2892;
	wire n2894;
	wire n2895;
	wire n2896;
	wire n2897;
	wire n2898;
	wire n2899;
	wire n2900;
	wire n2901;
	wire n2902;
	wire n2903;
	wire n2904;
	wire n2905;
	wire n2906;
	wire n2907;
	wire n2908;
	wire n2909;
	wire n2911;
	wire n2912;
	wire n2913;
	wire n2914;
	wire n2915;
	wire n2916;
	wire n2917;
	wire n2918;
	wire n2919;
	wire n2920;
	wire n2921;
	wire n2922;
	wire n2923;
	wire n2924;
	wire n2925;
	wire n2926;
	wire n2928;
	wire n2929;
	wire n2930;
	wire n2931;
	wire n2932;
	wire n2933;
	wire n2934;
	wire n2935;
	wire n2936;
	wire n2937;
	wire n2938;
	wire n2939;
	wire n2940;
	wire n2941;
	wire n2942;
	wire n2943;
	wire n2945;
	wire n2946;
	wire n2947;
	wire n2948;
	wire n2949;
	wire n2950;
	wire n2951;
	wire n2952;
	wire n2953;
	wire n2954;
	wire n2955;
	wire n2956;
	wire n2957;
	wire n2958;
	wire n2959;
	wire n2960;
	wire n2962;
	wire n2963;
	wire n2964;
	wire n2965;
	wire n2966;
	wire n2967;
	wire n2968;
	wire n2969;
	wire n2970;
	wire n2971;
	wire n2972;
	wire n2973;
	wire n2974;
	wire n2975;
	wire n2976;
	wire n2977;
	wire n2979;
	wire n2980;
	wire n2981;
	wire n2982;
	wire n2983;
	wire n2984;
	wire n2985;
	wire n2986;
	wire n2987;
	wire n2988;
	wire n2989;
	wire n2990;
	wire n2991;
	wire n2992;
	wire n2993;
	wire n2994;
	wire n2996;
	wire n2997;
	wire n2998;
	wire n2999;
	wire n3000;
	wire n3001;
	wire n3002;
	wire n3003;
	wire n3004;
	wire n3005;
	wire n3006;
	wire n3007;
	wire n3008;
	wire n3009;
	wire n3010;
	wire n3011;
	wire n3013;
	wire n3014;
	wire n3015;
	wire n3016;
	wire n3017;
	wire n3018;
	wire n3019;
	wire n3020;
	wire n3021;
	wire n3022;
	wire n3023;
	wire n3024;
	wire n3025;
	wire n3026;
	wire n3027;
	wire n3028;
	wire n3030;
	wire n3031;
	wire n3033;
	wire n3034;
	wire n3036;
	wire n3037;
	wire n3039;
	wire n3040;
	wire n3042;
	wire n3043;
	wire n3045;
	wire n3046;
	wire n3048;
	wire n3049;
	wire n3051;
	wire n3052;
	wire n3054;
	wire n3055;
	wire n3057;
	wire n3058;
	wire n3060;
	wire n3061;
	wire n3063;
	wire n3064;
	wire n3066;
	wire n3067;
	wire n3069;
	wire n3070;
	wire n3072;
	wire n3073;
	wire n3075;
	wire n3076;
	wire n3078;
	wire n3079;
	wire n3081;
	wire n3082;
	wire n3084;
	wire n3085;
	wire n3087;
	wire n3088;
	wire n3090;
	wire n3091;
	wire n3093;
	wire n3094;
	wire n3096;
	wire n3097;
	wire n3099;
	wire n3100;
	wire n3102;
	wire n3103;
	wire n3105;
	wire n3106;
	wire n3108;
	wire n3109;
	wire n3111;
	wire n3112;
	wire n3114;
	wire n3115;
	wire n3117;
	wire n3118;
	wire n3120;
	wire n3121;
	wire n3123;
	wire n3124;
	wire n3126;
	wire n3127;
	wire n3129;
	wire n3130;
	wire n3132;
	wire n3133;
	wire n3135;
	wire n3136;
	wire n3138;
	wire n3139;
	wire n3141;
	wire n3142;
	wire n3144;
	wire n3145;
	wire n3147;
	wire n3148;
	wire n3150;
	wire n3151;
	wire n3153;
	wire n3154;
	wire n3156;
	wire n3157;
	wire n3159;
	wire n3160;
	wire n3162;
	wire n3163;
	wire n3165;
	wire n3166;
	wire n3168;
	wire n3169;
	wire n3171;
	wire n3172;
	wire n3174;
	wire n3175;
	wire n3177;
	wire n3178;
	wire n3180;
	wire n3181;
	wire n3183;
	wire n3184;
	wire n3186;
	wire n3187;
	wire n3189;
	wire n3190;
	wire n3192;
	wire n3193;
	wire n3195;
	wire n3196;
	wire n3198;
	wire n3199;
	wire n3201;
	wire n3202;
	wire n3204;
	wire n3205;
	wire n3207;
	wire n3208;
	wire n3210;
	wire n3211;
	wire n3213;
	wire n3214;
	wire n3216;
	wire n3217;
	wire n3219;
	wire n3220;
	wire [1:0] w_a0_0;
	wire [1:0] w_a1_0;
	wire [1:0] w_a2_0;
	wire [1:0] w_a3_0;
	wire [1:0] w_a4_0;
	wire [1:0] w_a5_0;
	wire [1:0] w_a6_0;
	wire [1:0] w_a7_0;
	wire [1:0] w_a8_0;
	wire [1:0] w_a9_0;
	wire [1:0] w_a10_0;
	wire [1:0] w_a11_0;
	wire [1:0] w_a12_0;
	wire [1:0] w_a13_0;
	wire [1:0] w_a14_0;
	wire [1:0] w_a15_0;
	wire [1:0] w_a16_0;
	wire [1:0] w_a17_0;
	wire [1:0] w_a18_0;
	wire [1:0] w_a19_0;
	wire [1:0] w_a20_0;
	wire [1:0] w_a21_0;
	wire [1:0] w_a22_0;
	wire [1:0] w_a23_0;
	wire [1:0] w_a24_0;
	wire [1:0] w_a25_0;
	wire [1:0] w_a26_0;
	wire [1:0] w_a27_0;
	wire [1:0] w_a28_0;
	wire [1:0] w_a29_0;
	wire [1:0] w_a30_0;
	wire [1:0] w_a31_0;
	wire [1:0] w_a32_0;
	wire [1:0] w_a33_0;
	wire [1:0] w_a34_0;
	wire [1:0] w_a35_0;
	wire [1:0] w_a36_0;
	wire [1:0] w_a37_0;
	wire [1:0] w_a38_0;
	wire [1:0] w_a39_0;
	wire [1:0] w_a40_0;
	wire [1:0] w_a41_0;
	wire [1:0] w_a42_0;
	wire [1:0] w_a43_0;
	wire [1:0] w_a44_0;
	wire [1:0] w_a45_0;
	wire [1:0] w_a46_0;
	wire [1:0] w_a47_0;
	wire [1:0] w_a48_0;
	wire [1:0] w_a49_0;
	wire [1:0] w_a50_0;
	wire [1:0] w_a51_0;
	wire [1:0] w_a52_0;
	wire [1:0] w_a53_0;
	wire [1:0] w_a54_0;
	wire [1:0] w_a55_0;
	wire [1:0] w_a56_0;
	wire [1:0] w_a57_0;
	wire [1:0] w_a58_0;
	wire [1:0] w_a59_0;
	wire [1:0] w_a60_0;
	wire [1:0] w_a61_0;
	wire [1:0] w_a62_0;
	wire [1:0] w_a63_0;
	wire [1:0] w_a64_0;
	wire [1:0] w_a65_0;
	wire [1:0] w_a66_0;
	wire [1:0] w_a67_0;
	wire [1:0] w_a68_0;
	wire [1:0] w_a69_0;
	wire [1:0] w_a70_0;
	wire [1:0] w_a71_0;
	wire [1:0] w_a72_0;
	wire [1:0] w_a73_0;
	wire [1:0] w_a74_0;
	wire [1:0] w_a75_0;
	wire [1:0] w_a76_0;
	wire [1:0] w_a77_0;
	wire [1:0] w_a78_0;
	wire [1:0] w_a79_0;
	wire [1:0] w_a80_0;
	wire [1:0] w_a81_0;
	wire [1:0] w_a82_0;
	wire [1:0] w_a83_0;
	wire [1:0] w_a84_0;
	wire [1:0] w_a85_0;
	wire [1:0] w_a86_0;
	wire [1:0] w_a87_0;
	wire [1:0] w_a88_0;
	wire [1:0] w_a89_0;
	wire [1:0] w_a90_0;
	wire [1:0] w_a91_0;
	wire [1:0] w_a92_0;
	wire [1:0] w_a93_0;
	wire [1:0] w_a94_0;
	wire [1:0] w_a95_0;
	wire [1:0] w_a96_0;
	wire [1:0] w_a97_0;
	wire [1:0] w_a98_0;
	wire [1:0] w_a99_0;
	wire [1:0] w_a100_0;
	wire [1:0] w_a101_0;
	wire [1:0] w_a102_0;
	wire [1:0] w_a103_0;
	wire [1:0] w_a104_0;
	wire [1:0] w_a105_0;
	wire [1:0] w_a106_0;
	wire [1:0] w_a107_0;
	wire [1:0] w_a108_0;
	wire [1:0] w_a109_0;
	wire [1:0] w_a110_0;
	wire [1:0] w_a111_0;
	wire [1:0] w_a112_0;
	wire [1:0] w_a113_0;
	wire [1:0] w_a114_0;
	wire [1:0] w_a115_0;
	wire [1:0] w_a116_0;
	wire [1:0] w_a117_0;
	wire [1:0] w_a118_0;
	wire [1:0] w_a119_0;
	wire [1:0] w_a120_0;
	wire [1:0] w_a121_0;
	wire [1:0] w_a122_0;
	wire [1:0] w_a123_0;
	wire [1:0] w_a124_0;
	wire [1:0] w_a125_0;
	wire [1:0] w_a126_0;
	wire [1:0] w_a127_0;
	wire [2:0] w_shift0_0;
	wire [2:0] w_shift0_1;
	wire [2:0] w_shift0_2;
	wire [2:0] w_shift0_3;
	wire [2:0] w_shift0_4;
	wire [2:0] w_shift0_5;
	wire [2:0] w_shift0_6;
	wire [2:0] w_shift0_7;
	wire [2:0] w_shift0_8;
	wire [2:0] w_shift0_9;
	wire [2:0] w_shift0_10;
	wire [2:0] w_shift0_11;
	wire [2:0] w_shift0_12;
	wire [2:0] w_shift0_13;
	wire [2:0] w_shift0_14;
	wire [2:0] w_shift0_15;
	wire [2:0] w_shift0_16;
	wire [2:0] w_shift0_17;
	wire [2:0] w_shift0_18;
	wire [2:0] w_shift0_19;
	wire [2:0] w_shift0_20;
	wire [2:0] w_shift0_21;
	wire [2:0] w_shift0_22;
	wire [2:0] w_shift0_23;
	wire [2:0] w_shift0_24;
	wire [2:0] w_shift0_25;
	wire [2:0] w_shift0_26;
	wire [2:0] w_shift0_27;
	wire [2:0] w_shift0_28;
	wire [2:0] w_shift0_29;
	wire [2:0] w_shift0_30;
	wire [2:0] w_shift0_31;
	wire [2:0] w_shift0_32;
	wire [2:0] w_shift0_33;
	wire [2:0] w_shift0_34;
	wire [2:0] w_shift0_35;
	wire [2:0] w_shift0_36;
	wire [2:0] w_shift0_37;
	wire [2:0] w_shift0_38;
	wire [2:0] w_shift0_39;
	wire [2:0] w_shift0_40;
	wire [2:0] w_shift0_41;
	wire [2:0] w_shift0_42;
	wire [2:0] w_shift0_43;
	wire [2:0] w_shift0_44;
	wire [2:0] w_shift0_45;
	wire [2:0] w_shift0_46;
	wire [2:0] w_shift0_47;
	wire [2:0] w_shift0_48;
	wire [2:0] w_shift0_49;
	wire [2:0] w_shift0_50;
	wire [2:0] w_shift0_51;
	wire [2:0] w_shift0_52;
	wire [2:0] w_shift0_53;
	wire [2:0] w_shift0_54;
	wire [2:0] w_shift0_55;
	wire [2:0] w_shift0_56;
	wire [2:0] w_shift0_57;
	wire [2:0] w_shift0_58;
	wire [2:0] w_shift0_59;
	wire [2:0] w_shift0_60;
	wire [2:0] w_shift0_61;
	wire [2:0] w_shift0_62;
	wire [2:0] w_shift0_63;
	wire [2:0] w_shift1_0;
	wire [2:0] w_shift1_1;
	wire [2:0] w_shift1_2;
	wire [2:0] w_shift1_3;
	wire [2:0] w_shift1_4;
	wire [2:0] w_shift1_5;
	wire [2:0] w_shift1_6;
	wire [2:0] w_shift1_7;
	wire [2:0] w_shift1_8;
	wire [2:0] w_shift1_9;
	wire [2:0] w_shift1_10;
	wire [2:0] w_shift1_11;
	wire [2:0] w_shift1_12;
	wire [2:0] w_shift1_13;
	wire [2:0] w_shift1_14;
	wire [2:0] w_shift1_15;
	wire [2:0] w_shift1_16;
	wire [2:0] w_shift1_17;
	wire [2:0] w_shift1_18;
	wire [2:0] w_shift1_19;
	wire [2:0] w_shift1_20;
	wire [2:0] w_shift1_21;
	wire [2:0] w_shift1_22;
	wire [2:0] w_shift1_23;
	wire [2:0] w_shift1_24;
	wire [2:0] w_shift1_25;
	wire [2:0] w_shift1_26;
	wire [2:0] w_shift1_27;
	wire [2:0] w_shift1_28;
	wire [2:0] w_shift1_29;
	wire [2:0] w_shift1_30;
	wire [2:0] w_shift1_31;
	wire [2:0] w_shift1_32;
	wire [2:0] w_shift1_33;
	wire [2:0] w_shift1_34;
	wire [2:0] w_shift1_35;
	wire [2:0] w_shift1_36;
	wire [2:0] w_shift1_37;
	wire [2:0] w_shift1_38;
	wire [2:0] w_shift1_39;
	wire [2:0] w_shift1_40;
	wire [2:0] w_shift1_41;
	wire [2:0] w_shift1_42;
	wire [2:0] w_shift1_43;
	wire [2:0] w_shift1_44;
	wire [2:0] w_shift1_45;
	wire [2:0] w_shift1_46;
	wire [2:0] w_shift1_47;
	wire [2:0] w_shift1_48;
	wire [2:0] w_shift1_49;
	wire [2:0] w_shift1_50;
	wire [2:0] w_shift1_51;
	wire [2:0] w_shift1_52;
	wire [2:0] w_shift1_53;
	wire [2:0] w_shift1_54;
	wire [2:0] w_shift1_55;
	wire [2:0] w_shift1_56;
	wire [2:0] w_shift1_57;
	wire [2:0] w_shift1_58;
	wire [2:0] w_shift1_59;
	wire [2:0] w_shift1_60;
	wire [2:0] w_shift1_61;
	wire [2:0] w_shift1_62;
	wire [2:0] w_shift1_63;
	wire [2:0] w_shift2_0;
	wire [2:0] w_shift3_0;
	wire [2:0] w_shift4_0;
	wire [2:0] w_shift5_0;
	wire [2:0] w_shift6_0;
	wire [2:0] w_shift6_1;
	wire [2:0] w_shift6_2;
	wire [2:0] w_shift6_3;
	wire [2:0] w_shift6_4;
	wire [2:0] w_shift6_5;
	wire [2:0] w_shift6_6;
	wire [2:0] w_shift6_7;
	wire [2:0] w_shift6_8;
	wire [2:0] w_shift6_9;
	wire [2:0] w_shift6_10;
	wire [2:0] w_shift6_11;
	wire [2:0] w_shift6_12;
	wire [2:0] w_shift6_13;
	wire [2:0] w_shift6_14;
	wire [2:0] w_shift6_15;
	wire [2:0] w_shift6_16;
	wire [2:0] w_shift6_17;
	wire [2:0] w_shift6_18;
	wire [2:0] w_shift6_19;
	wire [2:0] w_shift6_20;
	wire [2:0] w_shift6_21;
	wire [2:0] w_shift6_22;
	wire [2:0] w_shift6_23;
	wire [2:0] w_shift6_24;
	wire [2:0] w_shift6_25;
	wire [2:0] w_shift6_26;
	wire [2:0] w_shift6_27;
	wire [2:0] w_shift6_28;
	wire [2:0] w_shift6_29;
	wire [2:0] w_shift6_30;
	wire [2:0] w_shift6_31;
	wire [2:0] w_shift6_32;
	wire [2:0] w_shift6_33;
	wire [2:0] w_shift6_34;
	wire [2:0] w_shift6_35;
	wire [2:0] w_shift6_36;
	wire [2:0] w_shift6_37;
	wire [2:0] w_shift6_38;
	wire [2:0] w_shift6_39;
	wire [2:0] w_shift6_40;
	wire [2:0] w_shift6_41;
	wire [2:0] w_shift6_42;
	wire [2:0] w_shift6_43;
	wire [2:0] w_shift6_44;
	wire [2:0] w_shift6_45;
	wire [2:0] w_shift6_46;
	wire [2:0] w_shift6_47;
	wire [2:0] w_shift6_48;
	wire [2:0] w_shift6_49;
	wire [2:0] w_shift6_50;
	wire [2:0] w_shift6_51;
	wire [2:0] w_shift6_52;
	wire [2:0] w_shift6_53;
	wire [2:0] w_shift6_54;
	wire [2:0] w_shift6_55;
	wire [2:0] w_shift6_56;
	wire [2:0] w_shift6_57;
	wire [2:0] w_shift6_58;
	wire [2:0] w_shift6_59;
	wire [2:0] w_shift6_60;
	wire [2:0] w_shift6_61;
	wire [2:0] w_shift6_62;
	wire [2:0] w_shift6_63;
	wire [2:0] w_n263_0;
	wire [2:0] w_n263_1;
	wire [2:0] w_n263_2;
	wire [2:0] w_n263_3;
	wire [2:0] w_n263_4;
	wire [2:0] w_n263_5;
	wire [2:0] w_n263_6;
	wire [2:0] w_n263_7;
	wire [2:0] w_n263_8;
	wire [2:0] w_n263_9;
	wire [2:0] w_n263_10;
	wire [2:0] w_n263_11;
	wire [2:0] w_n263_12;
	wire [2:0] w_n263_13;
	wire [2:0] w_n263_14;
	wire [2:0] w_n263_15;
	wire [2:0] w_n263_16;
	wire [2:0] w_n263_17;
	wire [2:0] w_n263_18;
	wire [2:0] w_n263_19;
	wire [2:0] w_n263_20;
	wire [2:0] w_n263_21;
	wire [2:0] w_n263_22;
	wire [2:0] w_n263_23;
	wire [2:0] w_n263_24;
	wire [2:0] w_n263_25;
	wire [2:0] w_n263_26;
	wire [2:0] w_n263_27;
	wire [2:0] w_n263_28;
	wire [2:0] w_n263_29;
	wire [2:0] w_n263_30;
	wire [2:0] w_n263_31;
	wire [2:0] w_n263_32;
	wire [2:0] w_n263_33;
	wire [2:0] w_n263_34;
	wire [2:0] w_n263_35;
	wire [2:0] w_n263_36;
	wire [2:0] w_n263_37;
	wire [2:0] w_n263_38;
	wire [2:0] w_n263_39;
	wire [2:0] w_n263_40;
	wire [2:0] w_n263_41;
	wire [2:0] w_n263_42;
	wire [2:0] w_n263_43;
	wire [2:0] w_n263_44;
	wire [2:0] w_n263_45;
	wire [2:0] w_n263_46;
	wire [2:0] w_n263_47;
	wire [2:0] w_n263_48;
	wire [2:0] w_n263_49;
	wire [2:0] w_n263_50;
	wire [2:0] w_n263_51;
	wire [2:0] w_n263_52;
	wire [2:0] w_n263_53;
	wire [2:0] w_n263_54;
	wire [2:0] w_n263_55;
	wire [2:0] w_n263_56;
	wire [2:0] w_n263_57;
	wire [2:0] w_n263_58;
	wire [2:0] w_n263_59;
	wire [2:0] w_n263_60;
	wire [2:0] w_n263_61;
	wire [2:0] w_n263_62;
	wire [1:0] w_n263_63;
	wire [1:0] w_n264_0;
	wire [2:0] w_n265_0;
	wire [2:0] w_n265_1;
	wire [2:0] w_n265_2;
	wire [2:0] w_n265_3;
	wire [2:0] w_n265_4;
	wire [2:0] w_n265_5;
	wire [2:0] w_n265_6;
	wire [2:0] w_n265_7;
	wire [2:0] w_n265_8;
	wire [2:0] w_n265_9;
	wire [2:0] w_n265_10;
	wire [2:0] w_n265_11;
	wire [2:0] w_n265_12;
	wire [2:0] w_n265_13;
	wire [2:0] w_n265_14;
	wire [2:0] w_n265_15;
	wire [2:0] w_n265_16;
	wire [2:0] w_n265_17;
	wire [2:0] w_n265_18;
	wire [2:0] w_n265_19;
	wire [2:0] w_n265_20;
	wire [2:0] w_n265_21;
	wire [2:0] w_n265_22;
	wire [2:0] w_n265_23;
	wire [2:0] w_n265_24;
	wire [2:0] w_n265_25;
	wire [2:0] w_n265_26;
	wire [2:0] w_n265_27;
	wire [2:0] w_n265_28;
	wire [2:0] w_n265_29;
	wire [2:0] w_n265_30;
	wire [2:0] w_n265_31;
	wire [2:0] w_n265_32;
	wire [2:0] w_n265_33;
	wire [2:0] w_n265_34;
	wire [2:0] w_n265_35;
	wire [2:0] w_n265_36;
	wire [2:0] w_n265_37;
	wire [2:0] w_n265_38;
	wire [2:0] w_n265_39;
	wire [2:0] w_n265_40;
	wire [2:0] w_n265_41;
	wire [2:0] w_n265_42;
	wire [2:0] w_n265_43;
	wire [2:0] w_n265_44;
	wire [2:0] w_n265_45;
	wire [2:0] w_n265_46;
	wire [2:0] w_n265_47;
	wire [2:0] w_n265_48;
	wire [2:0] w_n265_49;
	wire [2:0] w_n265_50;
	wire [2:0] w_n265_51;
	wire [2:0] w_n265_52;
	wire [2:0] w_n265_53;
	wire [2:0] w_n265_54;
	wire [2:0] w_n265_55;
	wire [2:0] w_n265_56;
	wire [2:0] w_n265_57;
	wire [2:0] w_n265_58;
	wire [2:0] w_n265_59;
	wire [2:0] w_n265_60;
	wire [2:0] w_n265_61;
	wire [2:0] w_n265_62;
	wire [1:0] w_n265_63;
	wire [1:0] w_n266_0;
	wire [2:0] w_n267_0;
	wire [2:0] w_n267_1;
	wire [2:0] w_n267_2;
	wire [2:0] w_n267_3;
	wire [2:0] w_n267_4;
	wire [2:0] w_n267_5;
	wire [2:0] w_n267_6;
	wire [2:0] w_n267_7;
	wire [2:0] w_n267_8;
	wire [2:0] w_n267_9;
	wire [2:0] w_n267_10;
	wire [2:0] w_n267_11;
	wire [2:0] w_n267_12;
	wire [2:0] w_n267_13;
	wire [2:0] w_n267_14;
	wire [2:0] w_n267_15;
	wire [2:0] w_n267_16;
	wire [2:0] w_n267_17;
	wire [2:0] w_n267_18;
	wire [2:0] w_n267_19;
	wire [2:0] w_n267_20;
	wire [2:0] w_n267_21;
	wire [2:0] w_n267_22;
	wire [2:0] w_n267_23;
	wire [2:0] w_n267_24;
	wire [2:0] w_n267_25;
	wire [2:0] w_n267_26;
	wire [2:0] w_n267_27;
	wire [2:0] w_n267_28;
	wire [2:0] w_n267_29;
	wire [2:0] w_n267_30;
	wire [2:0] w_n267_31;
	wire [2:0] w_n267_32;
	wire [2:0] w_n267_33;
	wire [2:0] w_n267_34;
	wire [2:0] w_n267_35;
	wire [2:0] w_n267_36;
	wire [2:0] w_n267_37;
	wire [2:0] w_n267_38;
	wire [2:0] w_n267_39;
	wire [2:0] w_n267_40;
	wire [2:0] w_n267_41;
	wire [2:0] w_n267_42;
	wire [2:0] w_n267_43;
	wire [2:0] w_n267_44;
	wire [2:0] w_n267_45;
	wire [2:0] w_n267_46;
	wire [2:0] w_n267_47;
	wire [2:0] w_n267_48;
	wire [2:0] w_n267_49;
	wire [2:0] w_n267_50;
	wire [2:0] w_n267_51;
	wire [2:0] w_n267_52;
	wire [2:0] w_n267_53;
	wire [2:0] w_n267_54;
	wire [2:0] w_n267_55;
	wire [2:0] w_n267_56;
	wire [2:0] w_n267_57;
	wire [2:0] w_n267_58;
	wire [2:0] w_n267_59;
	wire [2:0] w_n267_60;
	wire [2:0] w_n267_61;
	wire [2:0] w_n267_62;
	wire [1:0] w_n267_63;
	wire [2:0] w_n269_0;
	wire [2:0] w_n269_1;
	wire [2:0] w_n269_2;
	wire [2:0] w_n269_3;
	wire [2:0] w_n269_4;
	wire [2:0] w_n269_5;
	wire [2:0] w_n269_6;
	wire [2:0] w_n269_7;
	wire [2:0] w_n269_8;
	wire [2:0] w_n269_9;
	wire [2:0] w_n269_10;
	wire [2:0] w_n269_11;
	wire [2:0] w_n269_12;
	wire [2:0] w_n269_13;
	wire [2:0] w_n269_14;
	wire [2:0] w_n269_15;
	wire [2:0] w_n269_16;
	wire [2:0] w_n269_17;
	wire [2:0] w_n269_18;
	wire [2:0] w_n269_19;
	wire [2:0] w_n269_20;
	wire [2:0] w_n269_21;
	wire [2:0] w_n269_22;
	wire [2:0] w_n269_23;
	wire [2:0] w_n269_24;
	wire [2:0] w_n269_25;
	wire [2:0] w_n269_26;
	wire [2:0] w_n269_27;
	wire [2:0] w_n269_28;
	wire [2:0] w_n269_29;
	wire [2:0] w_n269_30;
	wire [2:0] w_n269_31;
	wire [2:0] w_n269_32;
	wire [2:0] w_n269_33;
	wire [2:0] w_n269_34;
	wire [2:0] w_n269_35;
	wire [2:0] w_n269_36;
	wire [2:0] w_n269_37;
	wire [2:0] w_n269_38;
	wire [2:0] w_n269_39;
	wire [2:0] w_n269_40;
	wire [2:0] w_n269_41;
	wire [2:0] w_n269_42;
	wire [2:0] w_n269_43;
	wire [2:0] w_n269_44;
	wire [2:0] w_n269_45;
	wire [2:0] w_n269_46;
	wire [2:0] w_n269_47;
	wire [2:0] w_n269_48;
	wire [2:0] w_n269_49;
	wire [2:0] w_n269_50;
	wire [2:0] w_n269_51;
	wire [2:0] w_n269_52;
	wire [2:0] w_n269_53;
	wire [2:0] w_n269_54;
	wire [2:0] w_n269_55;
	wire [2:0] w_n269_56;
	wire [2:0] w_n269_57;
	wire [2:0] w_n269_58;
	wire [2:0] w_n269_59;
	wire [2:0] w_n269_60;
	wire [2:0] w_n269_61;
	wire [2:0] w_n269_62;
	wire [1:0] w_n269_63;
	wire [1:0] w_n271_0;
	wire [2:0] w_n273_0;
	wire [2:0] w_n273_1;
	wire [2:0] w_n273_2;
	wire [2:0] w_n273_3;
	wire [2:0] w_n273_4;
	wire [2:0] w_n273_5;
	wire [2:0] w_n273_6;
	wire [2:0] w_n273_7;
	wire [2:0] w_n273_8;
	wire [2:0] w_n273_9;
	wire [2:0] w_n273_10;
	wire [2:0] w_n273_11;
	wire [2:0] w_n273_12;
	wire [2:0] w_n273_13;
	wire [2:0] w_n273_14;
	wire [2:0] w_n273_15;
	wire [2:0] w_n273_16;
	wire [2:0] w_n273_17;
	wire [2:0] w_n273_18;
	wire [2:0] w_n273_19;
	wire [2:0] w_n273_20;
	wire [2:0] w_n273_21;
	wire [2:0] w_n273_22;
	wire [2:0] w_n273_23;
	wire [2:0] w_n273_24;
	wire [2:0] w_n273_25;
	wire [2:0] w_n273_26;
	wire [2:0] w_n273_27;
	wire [2:0] w_n273_28;
	wire [2:0] w_n273_29;
	wire [2:0] w_n273_30;
	wire [2:0] w_n273_31;
	wire [2:0] w_n273_32;
	wire [2:0] w_n273_33;
	wire [2:0] w_n273_34;
	wire [2:0] w_n273_35;
	wire [2:0] w_n273_36;
	wire [2:0] w_n273_37;
	wire [2:0] w_n273_38;
	wire [2:0] w_n273_39;
	wire [2:0] w_n273_40;
	wire [2:0] w_n273_41;
	wire [2:0] w_n273_42;
	wire [2:0] w_n273_43;
	wire [2:0] w_n273_44;
	wire [2:0] w_n273_45;
	wire [2:0] w_n273_46;
	wire [2:0] w_n273_47;
	wire [2:0] w_n273_48;
	wire [2:0] w_n273_49;
	wire [2:0] w_n273_50;
	wire [2:0] w_n273_51;
	wire [2:0] w_n273_52;
	wire [2:0] w_n273_53;
	wire [2:0] w_n273_54;
	wire [2:0] w_n273_55;
	wire [2:0] w_n273_56;
	wire [2:0] w_n273_57;
	wire [2:0] w_n273_58;
	wire [2:0] w_n273_59;
	wire [2:0] w_n273_60;
	wire [2:0] w_n273_61;
	wire [2:0] w_n273_62;
	wire [1:0] w_n273_63;
	wire [1:0] w_n276_0;
	wire [2:0] w_n278_0;
	wire [1:0] w_n278_1;
	wire [1:0] w_n280_0;
	wire [2:0] w_n281_0;
	wire [2:0] w_n281_1;
	wire [2:0] w_n281_2;
	wire [2:0] w_n281_3;
	wire [2:0] w_n281_4;
	wire [2:0] w_n281_5;
	wire [2:0] w_n281_6;
	wire [2:0] w_n281_7;
	wire [2:0] w_n281_8;
	wire [2:0] w_n281_9;
	wire [2:0] w_n281_10;
	wire [2:0] w_n281_11;
	wire [2:0] w_n281_12;
	wire [2:0] w_n281_13;
	wire [2:0] w_n281_14;
	wire [2:0] w_n281_15;
	wire [2:0] w_n281_16;
	wire [2:0] w_n281_17;
	wire [2:0] w_n281_18;
	wire [2:0] w_n281_19;
	wire [2:0] w_n281_20;
	wire [2:0] w_n281_21;
	wire [2:0] w_n281_22;
	wire [2:0] w_n281_23;
	wire [2:0] w_n281_24;
	wire [2:0] w_n281_25;
	wire [2:0] w_n281_26;
	wire [2:0] w_n281_27;
	wire [2:0] w_n281_28;
	wire [2:0] w_n281_29;
	wire [2:0] w_n281_30;
	wire [2:0] w_n281_31;
	wire [2:0] w_n281_32;
	wire [2:0] w_n281_33;
	wire [2:0] w_n281_34;
	wire [2:0] w_n281_35;
	wire [2:0] w_n281_36;
	wire [2:0] w_n281_37;
	wire [2:0] w_n281_38;
	wire [2:0] w_n281_39;
	wire [2:0] w_n281_40;
	wire [2:0] w_n281_41;
	wire [2:0] w_n281_42;
	wire [2:0] w_n281_43;
	wire [2:0] w_n281_44;
	wire [2:0] w_n281_45;
	wire [2:0] w_n281_46;
	wire [2:0] w_n281_47;
	wire [2:0] w_n281_48;
	wire [2:0] w_n281_49;
	wire [2:0] w_n281_50;
	wire [2:0] w_n281_51;
	wire [2:0] w_n281_52;
	wire [2:0] w_n281_53;
	wire [2:0] w_n281_54;
	wire [2:0] w_n281_55;
	wire [2:0] w_n281_56;
	wire [2:0] w_n281_57;
	wire [2:0] w_n281_58;
	wire [2:0] w_n281_59;
	wire [2:0] w_n281_60;
	wire [2:0] w_n281_61;
	wire [2:0] w_n281_62;
	wire [1:0] w_n281_63;
	wire [1:0] w_n284_0;
	wire [1:0] w_n288_0;
	wire [2:0] w_n290_0;
	wire [1:0] w_n290_1;
	wire [2:0] w_n292_0;
	wire [2:0] w_n292_1;
	wire [2:0] w_n292_2;
	wire [2:0] w_n292_3;
	wire [2:0] w_n292_4;
	wire [2:0] w_n292_5;
	wire [2:0] w_n292_6;
	wire [2:0] w_n292_7;
	wire [2:0] w_n292_8;
	wire [2:0] w_n292_9;
	wire [2:0] w_n292_10;
	wire [2:0] w_n292_11;
	wire [2:0] w_n292_12;
	wire [2:0] w_n292_13;
	wire [2:0] w_n292_14;
	wire [2:0] w_n292_15;
	wire [2:0] w_n292_16;
	wire [2:0] w_n292_17;
	wire [2:0] w_n292_18;
	wire [2:0] w_n292_19;
	wire [2:0] w_n292_20;
	wire [2:0] w_n292_21;
	wire [2:0] w_n292_22;
	wire [2:0] w_n292_23;
	wire [2:0] w_n292_24;
	wire [2:0] w_n292_25;
	wire [2:0] w_n292_26;
	wire [2:0] w_n292_27;
	wire [2:0] w_n292_28;
	wire [2:0] w_n292_29;
	wire [2:0] w_n292_30;
	wire [2:0] w_n292_31;
	wire [2:0] w_n292_32;
	wire [2:0] w_n292_33;
	wire [2:0] w_n292_34;
	wire [2:0] w_n292_35;
	wire [2:0] w_n292_36;
	wire [2:0] w_n292_37;
	wire [2:0] w_n292_38;
	wire [2:0] w_n292_39;
	wire [2:0] w_n292_40;
	wire [2:0] w_n292_41;
	wire [2:0] w_n292_42;
	wire [2:0] w_n292_43;
	wire [2:0] w_n292_44;
	wire [2:0] w_n292_45;
	wire [2:0] w_n292_46;
	wire [2:0] w_n292_47;
	wire [2:0] w_n292_48;
	wire [2:0] w_n292_49;
	wire [2:0] w_n292_50;
	wire [2:0] w_n292_51;
	wire [2:0] w_n292_52;
	wire [2:0] w_n292_53;
	wire [2:0] w_n292_54;
	wire [2:0] w_n292_55;
	wire [2:0] w_n292_56;
	wire [2:0] w_n292_57;
	wire [2:0] w_n292_58;
	wire [2:0] w_n292_59;
	wire [2:0] w_n292_60;
	wire [2:0] w_n292_61;
	wire [2:0] w_n292_62;
	wire [1:0] w_n292_63;
	wire [1:0] w_n295_0;
	wire [1:0] w_n299_0;
	wire [2:0] w_n301_0;
	wire [1:0] w_n301_1;
	wire [2:0] w_n304_0;
	wire [2:0] w_n304_1;
	wire [2:0] w_n304_2;
	wire [2:0] w_n304_3;
	wire [2:0] w_n304_4;
	wire [2:0] w_n304_5;
	wire [2:0] w_n304_6;
	wire [2:0] w_n304_7;
	wire [2:0] w_n304_8;
	wire [2:0] w_n304_9;
	wire [2:0] w_n304_10;
	wire [2:0] w_n304_11;
	wire [2:0] w_n304_12;
	wire [2:0] w_n304_13;
	wire [2:0] w_n304_14;
	wire [2:0] w_n304_15;
	wire [2:0] w_n304_16;
	wire [2:0] w_n304_17;
	wire [2:0] w_n304_18;
	wire [2:0] w_n304_19;
	wire [2:0] w_n304_20;
	wire [2:0] w_n304_21;
	wire [2:0] w_n304_22;
	wire [2:0] w_n304_23;
	wire [2:0] w_n304_24;
	wire [2:0] w_n304_25;
	wire [2:0] w_n304_26;
	wire [2:0] w_n304_27;
	wire [2:0] w_n304_28;
	wire [2:0] w_n304_29;
	wire [2:0] w_n304_30;
	wire [2:0] w_n304_31;
	wire [2:0] w_n304_32;
	wire [2:0] w_n304_33;
	wire [2:0] w_n304_34;
	wire [2:0] w_n304_35;
	wire [2:0] w_n304_36;
	wire [2:0] w_n304_37;
	wire [2:0] w_n304_38;
	wire [2:0] w_n304_39;
	wire [2:0] w_n304_40;
	wire [2:0] w_n304_41;
	wire [2:0] w_n304_42;
	wire [2:0] w_n304_43;
	wire [2:0] w_n304_44;
	wire [2:0] w_n304_45;
	wire [2:0] w_n304_46;
	wire [2:0] w_n304_47;
	wire [2:0] w_n304_48;
	wire [2:0] w_n304_49;
	wire [2:0] w_n304_50;
	wire [2:0] w_n304_51;
	wire [2:0] w_n304_52;
	wire [2:0] w_n304_53;
	wire [2:0] w_n304_54;
	wire [2:0] w_n304_55;
	wire [2:0] w_n304_56;
	wire [2:0] w_n304_57;
	wire [2:0] w_n304_58;
	wire [2:0] w_n304_59;
	wire [2:0] w_n304_60;
	wire [2:0] w_n304_61;
	wire [2:0] w_n304_62;
	wire [1:0] w_n304_63;
	wire [1:0] w_n307_0;
	wire [1:0] w_n311_0;
	wire [2:0] w_n313_0;
	wire [1:0] w_n313_1;
	wire [2:0] w_n316_0;
	wire [1:0] w_n316_1;
	wire [1:0] w_n318_0;
	wire [2:0] w_n319_0;
	wire [2:0] w_n319_1;
	wire [2:0] w_n319_2;
	wire [2:0] w_n319_3;
	wire [2:0] w_n319_4;
	wire [2:0] w_n319_5;
	wire [2:0] w_n319_6;
	wire [2:0] w_n319_7;
	wire [2:0] w_n319_8;
	wire [2:0] w_n319_9;
	wire [2:0] w_n319_10;
	wire [2:0] w_n319_11;
	wire [2:0] w_n319_12;
	wire [2:0] w_n319_13;
	wire [2:0] w_n319_14;
	wire [2:0] w_n319_15;
	wire [2:0] w_n319_16;
	wire [2:0] w_n319_17;
	wire [2:0] w_n319_18;
	wire [2:0] w_n319_19;
	wire [2:0] w_n319_20;
	wire [2:0] w_n319_21;
	wire [2:0] w_n319_22;
	wire [2:0] w_n319_23;
	wire [2:0] w_n319_24;
	wire [2:0] w_n319_25;
	wire [2:0] w_n319_26;
	wire [2:0] w_n319_27;
	wire [2:0] w_n319_28;
	wire [2:0] w_n319_29;
	wire [2:0] w_n319_30;
	wire [2:0] w_n319_31;
	wire [2:0] w_n319_32;
	wire [2:0] w_n319_33;
	wire [2:0] w_n319_34;
	wire [2:0] w_n319_35;
	wire [2:0] w_n319_36;
	wire [2:0] w_n319_37;
	wire [2:0] w_n319_38;
	wire [2:0] w_n319_39;
	wire [2:0] w_n319_40;
	wire [2:0] w_n319_41;
	wire [2:0] w_n319_42;
	wire [2:0] w_n319_43;
	wire [2:0] w_n319_44;
	wire [2:0] w_n319_45;
	wire [2:0] w_n319_46;
	wire [2:0] w_n319_47;
	wire [2:0] w_n319_48;
	wire [2:0] w_n319_49;
	wire [2:0] w_n319_50;
	wire [2:0] w_n319_51;
	wire [2:0] w_n319_52;
	wire [2:0] w_n319_53;
	wire [2:0] w_n319_54;
	wire [2:0] w_n319_55;
	wire [2:0] w_n319_56;
	wire [2:0] w_n319_57;
	wire [2:0] w_n319_58;
	wire [2:0] w_n319_59;
	wire [2:0] w_n319_60;
	wire [2:0] w_n319_61;
	wire [2:0] w_n319_62;
	wire [1:0] w_n319_63;
	wire [1:0] w_n322_0;
	wire [1:0] w_n326_0;
	wire [2:0] w_n328_0;
	wire [1:0] w_n328_1;
	wire [1:0] w_n332_0;
	wire [1:0] w_n336_0;
	wire [2:0] w_n338_0;
	wire [1:0] w_n338_1;
	wire [1:0] w_n342_0;
	wire [1:0] w_n346_0;
	wire [2:0] w_n348_0;
	wire [1:0] w_n348_1;
	wire [1:0] w_n353_0;
	wire [1:0] w_n357_0;
	wire [2:0] w_n359_0;
	wire [1:0] w_n359_1;
	wire [2:0] w_n362_0;
	wire [1:0] w_n362_1;
	wire [2:0] w_n364_0;
	wire [2:0] w_n364_1;
	wire [2:0] w_n364_2;
	wire [2:0] w_n364_3;
	wire [2:0] w_n364_4;
	wire [2:0] w_n364_5;
	wire [2:0] w_n364_6;
	wire [2:0] w_n364_7;
	wire [2:0] w_n364_8;
	wire [2:0] w_n364_9;
	wire [2:0] w_n364_10;
	wire [2:0] w_n364_11;
	wire [2:0] w_n364_12;
	wire [2:0] w_n364_13;
	wire [2:0] w_n364_14;
	wire [2:0] w_n364_15;
	wire [2:0] w_n364_16;
	wire [2:0] w_n364_17;
	wire [2:0] w_n364_18;
	wire [2:0] w_n364_19;
	wire [2:0] w_n364_20;
	wire [2:0] w_n364_21;
	wire [2:0] w_n364_22;
	wire [2:0] w_n364_23;
	wire [2:0] w_n364_24;
	wire [2:0] w_n364_25;
	wire [2:0] w_n364_26;
	wire [2:0] w_n364_27;
	wire [2:0] w_n364_28;
	wire [2:0] w_n364_29;
	wire [2:0] w_n364_30;
	wire [2:0] w_n364_31;
	wire [2:0] w_n364_32;
	wire [2:0] w_n364_33;
	wire [2:0] w_n364_34;
	wire [2:0] w_n364_35;
	wire [2:0] w_n364_36;
	wire [2:0] w_n364_37;
	wire [2:0] w_n364_38;
	wire [2:0] w_n364_39;
	wire [2:0] w_n364_40;
	wire [2:0] w_n364_41;
	wire [2:0] w_n364_42;
	wire [2:0] w_n364_43;
	wire [2:0] w_n364_44;
	wire [2:0] w_n364_45;
	wire [2:0] w_n364_46;
	wire [2:0] w_n364_47;
	wire [2:0] w_n364_48;
	wire [2:0] w_n364_49;
	wire [2:0] w_n364_50;
	wire [2:0] w_n364_51;
	wire [2:0] w_n364_52;
	wire [2:0] w_n364_53;
	wire [2:0] w_n364_54;
	wire [2:0] w_n364_55;
	wire [2:0] w_n364_56;
	wire [2:0] w_n364_57;
	wire [2:0] w_n364_58;
	wire [2:0] w_n364_59;
	wire [2:0] w_n364_60;
	wire [2:0] w_n364_61;
	wire [2:0] w_n364_62;
	wire [1:0] w_n364_63;
	wire [1:0] w_n367_0;
	wire [1:0] w_n371_0;
	wire [2:0] w_n373_0;
	wire [1:0] w_n373_1;
	wire [1:0] w_n377_0;
	wire [1:0] w_n381_0;
	wire [2:0] w_n383_0;
	wire [1:0] w_n383_1;
	wire [1:0] w_n387_0;
	wire [1:0] w_n391_0;
	wire [2:0] w_n393_0;
	wire [1:0] w_n393_1;
	wire [1:0] w_n398_0;
	wire [1:0] w_n402_0;
	wire [2:0] w_n404_0;
	wire [1:0] w_n404_1;
	wire [2:0] w_n407_0;
	wire [1:0] w_n407_1;
	wire [2:0] w_n410_0;
	wire [2:0] w_n410_1;
	wire [2:0] w_n410_2;
	wire [2:0] w_n410_3;
	wire [2:0] w_n410_4;
	wire [2:0] w_n410_5;
	wire [2:0] w_n410_6;
	wire [2:0] w_n410_7;
	wire [2:0] w_n410_8;
	wire [2:0] w_n410_9;
	wire [2:0] w_n410_10;
	wire [2:0] w_n410_11;
	wire [2:0] w_n410_12;
	wire [2:0] w_n410_13;
	wire [2:0] w_n410_14;
	wire [2:0] w_n410_15;
	wire [2:0] w_n410_16;
	wire [2:0] w_n410_17;
	wire [2:0] w_n410_18;
	wire [2:0] w_n410_19;
	wire [2:0] w_n410_20;
	wire [2:0] w_n410_21;
	wire [2:0] w_n410_22;
	wire [2:0] w_n410_23;
	wire [2:0] w_n410_24;
	wire [2:0] w_n410_25;
	wire [2:0] w_n410_26;
	wire [2:0] w_n410_27;
	wire [2:0] w_n410_28;
	wire [2:0] w_n410_29;
	wire [2:0] w_n410_30;
	wire [2:0] w_n410_31;
	wire [2:0] w_n410_32;
	wire [2:0] w_n410_33;
	wire [2:0] w_n410_34;
	wire [2:0] w_n410_35;
	wire [2:0] w_n410_36;
	wire [2:0] w_n410_37;
	wire [2:0] w_n410_38;
	wire [2:0] w_n410_39;
	wire [2:0] w_n410_40;
	wire [2:0] w_n410_41;
	wire [2:0] w_n410_42;
	wire [2:0] w_n410_43;
	wire [2:0] w_n410_44;
	wire [2:0] w_n410_45;
	wire [2:0] w_n410_46;
	wire [2:0] w_n410_47;
	wire [2:0] w_n410_48;
	wire [2:0] w_n410_49;
	wire [2:0] w_n410_50;
	wire [2:0] w_n410_51;
	wire [2:0] w_n410_52;
	wire [2:0] w_n410_53;
	wire [2:0] w_n410_54;
	wire [2:0] w_n410_55;
	wire [2:0] w_n410_56;
	wire [2:0] w_n410_57;
	wire [2:0] w_n410_58;
	wire [2:0] w_n410_59;
	wire [2:0] w_n410_60;
	wire [2:0] w_n410_61;
	wire [2:0] w_n410_62;
	wire [1:0] w_n410_63;
	wire [1:0] w_n413_0;
	wire [1:0] w_n417_0;
	wire [2:0] w_n419_0;
	wire [1:0] w_n419_1;
	wire [1:0] w_n423_0;
	wire [1:0] w_n427_0;
	wire [2:0] w_n429_0;
	wire [1:0] w_n429_1;
	wire [1:0] w_n433_0;
	wire [1:0] w_n437_0;
	wire [2:0] w_n439_0;
	wire [1:0] w_n439_1;
	wire [1:0] w_n444_0;
	wire [1:0] w_n448_0;
	wire [2:0] w_n450_0;
	wire [1:0] w_n450_1;
	wire [2:0] w_n453_0;
	wire [1:0] w_n453_1;
	wire [1:0] w_n456_0;
	wire [1:0] w_n460_0;
	wire [1:0] w_n464_0;
	wire [2:0] w_n466_0;
	wire [1:0] w_n466_1;
	wire [1:0] w_n470_0;
	wire [1:0] w_n474_0;
	wire [2:0] w_n476_0;
	wire [1:0] w_n476_1;
	wire [1:0] w_n480_0;
	wire [1:0] w_n484_0;
	wire [2:0] w_n486_0;
	wire [1:0] w_n486_1;
	wire [1:0] w_n491_0;
	wire [1:0] w_n495_0;
	wire [2:0] w_n497_0;
	wire [1:0] w_n497_1;
	wire [2:0] w_n500_0;
	wire [1:0] w_n500_1;
	wire [1:0] w_n504_0;
	wire [1:0] w_n508_0;
	wire [2:0] w_n510_0;
	wire [1:0] w_n510_1;
	wire [1:0] w_n514_0;
	wire [1:0] w_n518_0;
	wire [2:0] w_n520_0;
	wire [1:0] w_n520_1;
	wire [1:0] w_n524_0;
	wire [1:0] w_n528_0;
	wire [2:0] w_n530_0;
	wire [1:0] w_n530_1;
	wire [1:0] w_n535_0;
	wire [1:0] w_n539_0;
	wire [2:0] w_n541_0;
	wire [1:0] w_n541_1;
	wire [2:0] w_n544_0;
	wire [1:0] w_n544_1;
	wire [1:0] w_n548_0;
	wire [1:0] w_n552_0;
	wire [2:0] w_n554_0;
	wire [1:0] w_n554_1;
	wire [1:0] w_n558_0;
	wire [1:0] w_n562_0;
	wire [2:0] w_n564_0;
	wire [1:0] w_n564_1;
	wire [1:0] w_n568_0;
	wire [1:0] w_n572_0;
	wire [2:0] w_n574_0;
	wire [1:0] w_n574_1;
	wire [1:0] w_n579_0;
	wire [1:0] w_n583_0;
	wire [2:0] w_n585_0;
	wire [1:0] w_n585_1;
	wire [2:0] w_n588_0;
	wire [1:0] w_n588_1;
	wire [1:0] w_n593_0;
	wire [1:0] w_n597_0;
	wire [2:0] w_n599_0;
	wire [1:0] w_n599_1;
	wire [1:0] w_n603_0;
	wire [1:0] w_n607_0;
	wire [2:0] w_n609_0;
	wire [1:0] w_n609_1;
	wire [1:0] w_n613_0;
	wire [1:0] w_n617_0;
	wire [2:0] w_n619_0;
	wire [1:0] w_n619_1;
	wire [1:0] w_n624_0;
	wire [1:0] w_n628_0;
	wire [2:0] w_n630_0;
	wire [1:0] w_n630_1;
	wire [2:0] w_n633_0;
	wire [1:0] w_n633_1;
	wire [1:0] w_n636_0;
	wire [1:0] w_n641_0;
	wire [1:0] w_n645_0;
	wire [2:0] w_n647_0;
	wire [1:0] w_n647_1;
	wire [1:0] w_n651_0;
	wire [1:0] w_n655_0;
	wire [2:0] w_n657_0;
	wire [1:0] w_n657_1;
	wire [1:0] w_n661_0;
	wire [1:0] w_n665_0;
	wire [2:0] w_n667_0;
	wire [1:0] w_n667_1;
	wire [1:0] w_n672_0;
	wire [1:0] w_n676_0;
	wire [2:0] w_n678_0;
	wire [1:0] w_n678_1;
	wire [2:0] w_n681_0;
	wire [1:0] w_n681_1;
	wire [1:0] w_n685_0;
	wire [1:0] w_n689_0;
	wire [2:0] w_n691_0;
	wire [1:0] w_n691_1;
	wire [1:0] w_n695_0;
	wire [1:0] w_n699_0;
	wire [2:0] w_n701_0;
	wire [1:0] w_n701_1;
	wire [1:0] w_n705_0;
	wire [1:0] w_n709_0;
	wire [2:0] w_n711_0;
	wire [1:0] w_n711_1;
	wire [1:0] w_n716_0;
	wire [1:0] w_n720_0;
	wire [2:0] w_n722_0;
	wire [1:0] w_n722_1;
	wire [2:0] w_n725_0;
	wire [1:0] w_n725_1;
	wire [1:0] w_n729_0;
	wire [1:0] w_n733_0;
	wire [2:0] w_n735_0;
	wire [1:0] w_n735_1;
	wire [1:0] w_n739_0;
	wire [1:0] w_n743_0;
	wire [2:0] w_n745_0;
	wire [1:0] w_n745_1;
	wire [1:0] w_n749_0;
	wire [1:0] w_n753_0;
	wire [2:0] w_n755_0;
	wire [1:0] w_n755_1;
	wire [1:0] w_n760_0;
	wire [1:0] w_n764_0;
	wire [2:0] w_n766_0;
	wire [1:0] w_n766_1;
	wire [2:0] w_n769_0;
	wire [1:0] w_n769_1;
	wire [1:0] w_n774_0;
	wire [1:0] w_n778_0;
	wire [2:0] w_n780_0;
	wire [1:0] w_n780_1;
	wire [1:0] w_n784_0;
	wire [1:0] w_n788_0;
	wire [2:0] w_n790_0;
	wire [1:0] w_n790_1;
	wire [1:0] w_n794_0;
	wire [1:0] w_n798_0;
	wire [2:0] w_n800_0;
	wire [1:0] w_n800_1;
	wire [1:0] w_n805_0;
	wire [1:0] w_n809_0;
	wire [2:0] w_n811_0;
	wire [1:0] w_n811_1;
	wire [2:0] w_n814_0;
	wire [1:0] w_n814_1;
	wire [1:0] w_n817_0;
	wire [1:0] w_n821_0;
	wire [1:0] w_n825_0;
	wire [2:0] w_n827_0;
	wire [1:0] w_n827_1;
	wire [1:0] w_n831_0;
	wire [1:0] w_n835_0;
	wire [2:0] w_n837_0;
	wire [1:0] w_n837_1;
	wire [1:0] w_n841_0;
	wire [1:0] w_n845_0;
	wire [2:0] w_n847_0;
	wire [1:0] w_n847_1;
	wire [1:0] w_n852_0;
	wire [1:0] w_n856_0;
	wire [2:0] w_n858_0;
	wire [1:0] w_n858_1;
	wire [2:0] w_n861_0;
	wire [1:0] w_n861_1;
	wire [1:0] w_n865_0;
	wire [1:0] w_n869_0;
	wire [2:0] w_n871_0;
	wire [1:0] w_n871_1;
	wire [1:0] w_n875_0;
	wire [1:0] w_n879_0;
	wire [2:0] w_n881_0;
	wire [1:0] w_n881_1;
	wire [1:0] w_n885_0;
	wire [1:0] w_n889_0;
	wire [2:0] w_n891_0;
	wire [1:0] w_n891_1;
	wire [1:0] w_n896_0;
	wire [1:0] w_n900_0;
	wire [2:0] w_n902_0;
	wire [1:0] w_n902_1;
	wire [2:0] w_n905_0;
	wire [1:0] w_n905_1;
	wire [1:0] w_n909_0;
	wire [1:0] w_n913_0;
	wire [2:0] w_n915_0;
	wire [1:0] w_n915_1;
	wire [1:0] w_n919_0;
	wire [1:0] w_n923_0;
	wire [2:0] w_n925_0;
	wire [1:0] w_n925_1;
	wire [1:0] w_n929_0;
	wire [1:0] w_n933_0;
	wire [2:0] w_n935_0;
	wire [1:0] w_n935_1;
	wire [1:0] w_n940_0;
	wire [1:0] w_n944_0;
	wire [2:0] w_n946_0;
	wire [1:0] w_n946_1;
	wire [2:0] w_n949_0;
	wire [1:0] w_n949_1;
	wire [1:0] w_n954_0;
	wire [1:0] w_n958_0;
	wire [2:0] w_n960_0;
	wire [1:0] w_n960_1;
	wire [1:0] w_n964_0;
	wire [1:0] w_n968_0;
	wire [2:0] w_n970_0;
	wire [1:0] w_n970_1;
	wire [1:0] w_n974_0;
	wire [1:0] w_n978_0;
	wire [2:0] w_n980_0;
	wire [1:0] w_n980_1;
	wire [1:0] w_n985_0;
	wire [1:0] w_n989_0;
	wire [2:0] w_n991_0;
	wire [1:0] w_n991_1;
	wire [2:0] w_n994_0;
	wire [1:0] w_n994_1;
	wire [1:0] w_n997_0;
	wire [2:0] w_n1002_0;
	wire [1:0] w_n1002_1;
	wire [2:0] w_n1006_0;
	wire [1:0] w_n1006_1;
	wire [2:0] w_n1010_0;
	wire [1:0] w_n1010_1;
	wire [2:0] w_n1015_0;
	wire [1:0] w_n1015_1;
	wire [2:0] w_n1018_0;
	wire [1:0] w_n1018_1;
	wire [2:0] w_n1022_0;
	wire [1:0] w_n1022_1;
	wire [2:0] w_n1026_0;
	wire [1:0] w_n1026_1;
	wire [2:0] w_n1030_0;
	wire [1:0] w_n1030_1;
	wire [2:0] w_n1035_0;
	wire [1:0] w_n1035_1;
	wire [2:0] w_n1038_0;
	wire [1:0] w_n1038_1;
	wire [2:0] w_n1042_0;
	wire [1:0] w_n1042_1;
	wire [2:0] w_n1046_0;
	wire [1:0] w_n1046_1;
	wire [2:0] w_n1050_0;
	wire [1:0] w_n1050_1;
	wire [2:0] w_n1055_0;
	wire [1:0] w_n1055_1;
	wire [2:0] w_n1058_0;
	wire [1:0] w_n1058_1;
	wire [2:0] w_n1063_0;
	wire [1:0] w_n1063_1;
	wire [2:0] w_n1067_0;
	wire [1:0] w_n1067_1;
	wire [2:0] w_n1071_0;
	wire [1:0] w_n1071_1;
	wire [2:0] w_n1076_0;
	wire [1:0] w_n1076_1;
	wire [2:0] w_n1079_0;
	wire [1:0] w_n1079_1;
	wire [1:0] w_n1082_0;
	wire [2:0] w_n1086_0;
	wire [1:0] w_n1086_1;
	wire [2:0] w_n1090_0;
	wire [1:0] w_n1090_1;
	wire [2:0] w_n1094_0;
	wire [1:0] w_n1094_1;
	wire [2:0] w_n1099_0;
	wire [1:0] w_n1099_1;
	wire [2:0] w_n1102_0;
	wire [1:0] w_n1102_1;
	wire [2:0] w_n1106_0;
	wire [1:0] w_n1106_1;
	wire [2:0] w_n1110_0;
	wire [1:0] w_n1110_1;
	wire [2:0] w_n1114_0;
	wire [1:0] w_n1114_1;
	wire [2:0] w_n1119_0;
	wire [1:0] w_n1119_1;
	wire [2:0] w_n1122_0;
	wire [1:0] w_n1122_1;
	wire [2:0] w_n1126_0;
	wire [1:0] w_n1126_1;
	wire [2:0] w_n1130_0;
	wire [1:0] w_n1130_1;
	wire [2:0] w_n1134_0;
	wire [1:0] w_n1134_1;
	wire [2:0] w_n1139_0;
	wire [1:0] w_n1139_1;
	wire [2:0] w_n1142_0;
	wire [1:0] w_n1142_1;
	wire [2:0] w_n1147_0;
	wire [1:0] w_n1147_1;
	wire [2:0] w_n1151_0;
	wire [1:0] w_n1151_1;
	wire [2:0] w_n1155_0;
	wire [1:0] w_n1155_1;
	wire [2:0] w_n1160_0;
	wire [1:0] w_n1160_1;
	wire [2:0] w_n1163_0;
	wire [1:0] w_n1163_1;
	wire [1:0] w_n1166_0;
	wire [2:0] w_n1171_0;
	wire [1:0] w_n1171_1;
	wire [2:0] w_n1175_0;
	wire [1:0] w_n1175_1;
	wire [2:0] w_n1179_0;
	wire [1:0] w_n1179_1;
	wire [2:0] w_n1184_0;
	wire [1:0] w_n1184_1;
	wire [2:0] w_n1187_0;
	wire [1:0] w_n1187_1;
	wire [2:0] w_n1191_0;
	wire [1:0] w_n1191_1;
	wire [2:0] w_n1195_0;
	wire [1:0] w_n1195_1;
	wire [2:0] w_n1199_0;
	wire [1:0] w_n1199_1;
	wire [2:0] w_n1204_0;
	wire [1:0] w_n1204_1;
	wire [2:0] w_n1207_0;
	wire [1:0] w_n1207_1;
	wire [2:0] w_n1211_0;
	wire [1:0] w_n1211_1;
	wire [2:0] w_n1215_0;
	wire [1:0] w_n1215_1;
	wire [2:0] w_n1219_0;
	wire [1:0] w_n1219_1;
	wire [2:0] w_n1224_0;
	wire [1:0] w_n1224_1;
	wire [2:0] w_n1227_0;
	wire [1:0] w_n1227_1;
	wire [2:0] w_n1232_0;
	wire [1:0] w_n1232_1;
	wire [2:0] w_n1236_0;
	wire [1:0] w_n1236_1;
	wire [2:0] w_n1240_0;
	wire [1:0] w_n1240_1;
	wire [2:0] w_n1245_0;
	wire [1:0] w_n1245_1;
	wire [2:0] w_n1248_0;
	wire [1:0] w_n1248_1;
	wire [1:0] w_n1251_0;
	wire [2:0] w_n1255_0;
	wire [1:0] w_n1255_1;
	wire [2:0] w_n1259_0;
	wire [1:0] w_n1259_1;
	wire [2:0] w_n1263_0;
	wire [1:0] w_n1263_1;
	wire [2:0] w_n1268_0;
	wire [1:0] w_n1268_1;
	wire [2:0] w_n1271_0;
	wire [1:0] w_n1271_1;
	wire [2:0] w_n1275_0;
	wire [1:0] w_n1275_1;
	wire [2:0] w_n1279_0;
	wire [1:0] w_n1279_1;
	wire [2:0] w_n1283_0;
	wire [1:0] w_n1283_1;
	wire [2:0] w_n1288_0;
	wire [1:0] w_n1288_1;
	wire [2:0] w_n1291_0;
	wire [1:0] w_n1291_1;
	wire [2:0] w_n1295_0;
	wire [1:0] w_n1295_1;
	wire [2:0] w_n1299_0;
	wire [1:0] w_n1299_1;
	wire [2:0] w_n1303_0;
	wire [1:0] w_n1303_1;
	wire [2:0] w_n1308_0;
	wire [1:0] w_n1308_1;
	wire [2:0] w_n1311_0;
	wire [1:0] w_n1311_1;
	wire [2:0] w_n1316_0;
	wire [1:0] w_n1316_1;
	wire [2:0] w_n1320_0;
	wire [1:0] w_n1320_1;
	wire [2:0] w_n1324_0;
	wire [1:0] w_n1324_1;
	wire [2:0] w_n1329_0;
	wire [1:0] w_n1329_1;
	wire [2:0] w_n1332_0;
	wire [1:0] w_n1332_1;
	wire [1:0] w_n1335_0;
	wire [2:0] w_n1344_0;
	wire [1:0] w_n1344_1;
	wire [2:0] w_n1352_0;
	wire [1:0] w_n1352_1;
	wire [2:0] w_n1360_0;
	wire [1:0] w_n1360_1;
	wire [2:0] w_n1369_0;
	wire [1:0] w_n1369_1;
	wire [1:0] w_n1372_0;
	wire [2:0] w_n1380_0;
	wire [1:0] w_n1380_1;
	wire [2:0] w_n1388_0;
	wire [1:0] w_n1388_1;
	wire [2:0] w_n1396_0;
	wire [1:0] w_n1396_1;
	wire [2:0] w_n1405_0;
	wire [1:0] w_n1405_1;
	wire [1:0] w_n1408_0;
	wire [2:0] w_n1417_0;
	wire [1:0] w_n1417_1;
	wire [2:0] w_n1425_0;
	wire [1:0] w_n1425_1;
	wire [2:0] w_n1433_0;
	wire [1:0] w_n1433_1;
	wire [2:0] w_n1442_0;
	wire [1:0] w_n1442_1;
	wire [1:0] w_n1445_0;
	wire [2:0] w_n1453_0;
	wire [1:0] w_n1453_1;
	wire [2:0] w_n1461_0;
	wire [1:0] w_n1461_1;
	wire [2:0] w_n1469_0;
	wire [1:0] w_n1469_1;
	wire [2:0] w_n1478_0;
	wire [1:0] w_n1478_1;
	wire [1:0] w_n1481_0;
	wire [2:0] w_n1490_0;
	wire [1:0] w_n1490_1;
	wire [2:0] w_n1498_0;
	wire [1:0] w_n1498_1;
	wire [2:0] w_n1506_0;
	wire [1:0] w_n1506_1;
	wire [2:0] w_n1515_0;
	wire [1:0] w_n1515_1;
	wire [1:0] w_n1518_0;
	wire [2:0] w_n1526_0;
	wire [1:0] w_n1526_1;
	wire [2:0] w_n1534_0;
	wire [1:0] w_n1534_1;
	wire [2:0] w_n1542_0;
	wire [1:0] w_n1542_1;
	wire [2:0] w_n1551_0;
	wire [1:0] w_n1551_1;
	wire [1:0] w_n1554_0;
	wire [2:0] w_n1563_0;
	wire [1:0] w_n1563_1;
	wire [2:0] w_n1571_0;
	wire [1:0] w_n1571_1;
	wire [2:0] w_n1579_0;
	wire [1:0] w_n1579_1;
	wire [2:0] w_n1588_0;
	wire [1:0] w_n1588_1;
	wire [1:0] w_n1591_0;
	wire [2:0] w_n1599_0;
	wire [1:0] w_n1599_1;
	wire [2:0] w_n1607_0;
	wire [1:0] w_n1607_1;
	wire [2:0] w_n1615_0;
	wire [1:0] w_n1615_1;
	wire [2:0] w_n1624_0;
	wire [1:0] w_n1624_1;
	wire [1:0] w_n1627_0;
	wire [2:0] w_n1636_0;
	wire [1:0] w_n1636_1;
	wire [2:0] w_n1644_0;
	wire [1:0] w_n1644_1;
	wire [2:0] w_n1652_0;
	wire [1:0] w_n1652_1;
	wire [2:0] w_n1661_0;
	wire [1:0] w_n1661_1;
	wire [1:0] w_n1664_0;
	wire [2:0] w_n1672_0;
	wire [1:0] w_n1672_1;
	wire [2:0] w_n1680_0;
	wire [1:0] w_n1680_1;
	wire [2:0] w_n1688_0;
	wire [1:0] w_n1688_1;
	wire [2:0] w_n1697_0;
	wire [1:0] w_n1697_1;
	wire [1:0] w_n1700_0;
	wire [2:0] w_n1709_0;
	wire [1:0] w_n1709_1;
	wire [2:0] w_n1717_0;
	wire [1:0] w_n1717_1;
	wire [2:0] w_n1725_0;
	wire [1:0] w_n1725_1;
	wire [2:0] w_n1734_0;
	wire [1:0] w_n1734_1;
	wire [1:0] w_n1737_0;
	wire [2:0] w_n1745_0;
	wire [1:0] w_n1745_1;
	wire [2:0] w_n1753_0;
	wire [1:0] w_n1753_1;
	wire [2:0] w_n1761_0;
	wire [1:0] w_n1761_1;
	wire [2:0] w_n1770_0;
	wire [1:0] w_n1770_1;
	wire [1:0] w_n1773_0;
	wire [2:0] w_n1782_0;
	wire [1:0] w_n1782_1;
	wire [2:0] w_n1790_0;
	wire [1:0] w_n1790_1;
	wire [2:0] w_n1798_0;
	wire [1:0] w_n1798_1;
	wire [2:0] w_n1807_0;
	wire [1:0] w_n1807_1;
	wire [1:0] w_n1810_0;
	wire [2:0] w_n1818_0;
	wire [1:0] w_n1818_1;
	wire [2:0] w_n1826_0;
	wire [1:0] w_n1826_1;
	wire [2:0] w_n1834_0;
	wire [1:0] w_n1834_1;
	wire [2:0] w_n1843_0;
	wire [1:0] w_n1843_1;
	wire [1:0] w_n1846_0;
	wire [2:0] w_n1855_0;
	wire [1:0] w_n1855_1;
	wire [2:0] w_n1863_0;
	wire [1:0] w_n1863_1;
	wire [2:0] w_n1871_0;
	wire [1:0] w_n1871_1;
	wire [2:0] w_n1880_0;
	wire [1:0] w_n1880_1;
	wire [1:0] w_n1883_0;
	wire [2:0] w_n1891_0;
	wire [1:0] w_n1891_1;
	wire [2:0] w_n1899_0;
	wire [1:0] w_n1899_1;
	wire [2:0] w_n1907_0;
	wire [1:0] w_n1907_1;
	wire [2:0] w_n1916_0;
	wire [1:0] w_n1916_1;
	wire [1:0] w_n1919_0;
	wire [2:0] w_n1928_0;
	wire [1:0] w_n1928_1;
	wire [2:0] w_n1936_0;
	wire [1:0] w_n1936_1;
	wire [2:0] w_n1944_0;
	wire [1:0] w_n1944_1;
	wire [2:0] w_n1953_0;
	wire [1:0] w_n1953_1;
	wire [1:0] w_n1956_0;
	wire [2:0] w_n1964_0;
	wire [1:0] w_n1964_1;
	wire [2:0] w_n1972_0;
	wire [1:0] w_n1972_1;
	wire [2:0] w_n1980_0;
	wire [1:0] w_n1980_1;
	wire [2:0] w_n1989_0;
	wire [1:0] w_n1989_1;
	wire [1:0] w_n1992_0;
	wire [2:0] w_n2001_0;
	wire [1:0] w_n2001_1;
	wire [2:0] w_n2009_0;
	wire [1:0] w_n2009_1;
	wire [2:0] w_n2017_0;
	wire [1:0] w_n2017_1;
	wire [2:0] w_n2026_0;
	wire [1:0] w_n2026_1;
	wire [1:0] w_n2029_0;
	wire [2:0] w_n2037_0;
	wire [1:0] w_n2037_1;
	wire [2:0] w_n2045_0;
	wire [1:0] w_n2045_1;
	wire [2:0] w_n2053_0;
	wire [1:0] w_n2053_1;
	wire [2:0] w_n2062_0;
	wire [1:0] w_n2062_1;
	wire [1:0] w_n2065_0;
	wire [2:0] w_n2074_0;
	wire [1:0] w_n2074_1;
	wire [2:0] w_n2082_0;
	wire [1:0] w_n2082_1;
	wire [2:0] w_n2090_0;
	wire [1:0] w_n2090_1;
	wire [2:0] w_n2099_0;
	wire [1:0] w_n2099_1;
	wire [1:0] w_n2102_0;
	wire [2:0] w_n2110_0;
	wire [1:0] w_n2110_1;
	wire [2:0] w_n2118_0;
	wire [1:0] w_n2118_1;
	wire [2:0] w_n2126_0;
	wire [1:0] w_n2126_1;
	wire [2:0] w_n2135_0;
	wire [1:0] w_n2135_1;
	wire [1:0] w_n2138_0;
	wire [2:0] w_n2147_0;
	wire [1:0] w_n2147_1;
	wire [2:0] w_n2155_0;
	wire [1:0] w_n2155_1;
	wire [2:0] w_n2163_0;
	wire [1:0] w_n2163_1;
	wire [2:0] w_n2172_0;
	wire [1:0] w_n2172_1;
	wire [1:0] w_n2175_0;
	wire [2:0] w_n2183_0;
	wire [1:0] w_n2183_1;
	wire [2:0] w_n2191_0;
	wire [1:0] w_n2191_1;
	wire [2:0] w_n2199_0;
	wire [1:0] w_n2199_1;
	wire [2:0] w_n2208_0;
	wire [1:0] w_n2208_1;
	wire [1:0] w_n2211_0;
	wire [1:0] w_n2220_0;
	wire [1:0] w_n2228_0;
	wire [1:0] w_n2237_0;
	wire [1:0] w_n2245_0;
	wire [1:0] w_n2254_0;
	wire [1:0] w_n2262_0;
	wire [1:0] w_n2271_0;
	wire [1:0] w_n2279_0;
	wire [1:0] w_n2288_0;
	wire [1:0] w_n2296_0;
	wire [1:0] w_n2305_0;
	wire [1:0] w_n2313_0;
	wire [1:0] w_n2322_0;
	wire [1:0] w_n2330_0;
	wire [1:0] w_n2339_0;
	wire [1:0] w_n2347_0;
	wire [1:0] w_n2356_0;
	wire [1:0] w_n2364_0;
	wire [1:0] w_n2373_0;
	wire [1:0] w_n2381_0;
	wire [1:0] w_n2390_0;
	wire [1:0] w_n2398_0;
	wire [1:0] w_n2407_0;
	wire [1:0] w_n2415_0;
	wire [1:0] w_n2424_0;
	wire [1:0] w_n2432_0;
	wire [1:0] w_n2441_0;
	wire [1:0] w_n2449_0;
	wire [1:0] w_n2458_0;
	wire [1:0] w_n2466_0;
	wire [1:0] w_n2475_0;
	wire [1:0] w_n2483_0;
	wire [1:0] w_n2492_0;
	wire [1:0] w_n2500_0;
	wire [1:0] w_n2509_0;
	wire [1:0] w_n2517_0;
	wire [1:0] w_n2526_0;
	wire [1:0] w_n2534_0;
	wire [1:0] w_n2543_0;
	wire [1:0] w_n2551_0;
	wire [1:0] w_n2560_0;
	wire [1:0] w_n2568_0;
	wire [1:0] w_n2577_0;
	wire [1:0] w_n2585_0;
	wire [1:0] w_n2594_0;
	wire [1:0] w_n2602_0;
	wire [1:0] w_n2611_0;
	wire [1:0] w_n2619_0;
	wire [1:0] w_n2628_0;
	wire [1:0] w_n2636_0;
	wire [1:0] w_n2645_0;
	wire [1:0] w_n2653_0;
	wire [1:0] w_n2662_0;
	wire [1:0] w_n2670_0;
	wire [1:0] w_n2679_0;
	wire [1:0] w_n2687_0;
	wire [1:0] w_n2696_0;
	wire [1:0] w_n2704_0;
	wire [1:0] w_n2713_0;
	wire [1:0] w_n2721_0;
	wire [1:0] w_n2730_0;
	wire [1:0] w_n2738_0;
	wire [1:0] w_n2747_0;
	wire [1:0] w_n2755_0;
	wire [1:0] w_n2764_0;
	wire [1:0] w_n2772_0;
	wire [1:0] w_n2781_0;
	wire [1:0] w_n2789_0;
	wire [1:0] w_n2798_0;
	wire [1:0] w_n2806_0;
	wire [1:0] w_n2815_0;
	wire [1:0] w_n2823_0;
	wire [1:0] w_n2832_0;
	wire [1:0] w_n2840_0;
	wire [1:0] w_n2849_0;
	wire [1:0] w_n2857_0;
	wire [1:0] w_n2866_0;
	wire [1:0] w_n2874_0;
	wire [1:0] w_n2883_0;
	wire [1:0] w_n2891_0;
	wire [1:0] w_n2900_0;
	wire [1:0] w_n2908_0;
	wire [1:0] w_n2917_0;
	wire [1:0] w_n2925_0;
	wire [1:0] w_n2934_0;
	wire [1:0] w_n2942_0;
	wire [1:0] w_n2951_0;
	wire [1:0] w_n2959_0;
	wire [1:0] w_n2968_0;
	wire [1:0] w_n2976_0;
	wire [1:0] w_n2985_0;
	wire [1:0] w_n2993_0;
	wire [1:0] w_n3002_0;
	wire [1:0] w_n3010_0;
	wire [1:0] w_n3019_0;
	wire [1:0] w_n3027_0;
	wire w_dff_B_g1C06Xx82_1;
	wire w_dff_B_IqnWAkCL7_1;
	wire w_dff_B_HpkFhe6A1_0;
	wire w_dff_B_JoZ9Tb4V2_1;
	wire w_dff_B_UCm236lc9_1;
	wire w_dff_B_xuHcFHr59_0;
	wire w_dff_B_T8KfLGzT2_1;
	wire w_dff_B_E17iQHOA7_1;
	wire w_dff_B_gRp8Ggs88_0;
	wire w_dff_B_lIe0sgd26_1;
	wire w_dff_B_WfEiqaoK6_1;
	wire w_dff_B_cjYulRxp8_0;
	wire w_dff_B_D8gYIS3H8_1;
	wire w_dff_B_ZbjPw7uh6_1;
	wire w_dff_B_NanY4bA49_0;
	wire w_dff_B_2N8mDzIw8_1;
	wire w_dff_B_wVw0jevq6_1;
	wire w_dff_B_U2b0FtDF4_0;
	wire w_dff_B_wMj82kuC6_1;
	wire w_dff_B_x7FH33QW3_1;
	wire w_dff_B_PVP23snq0_0;
	wire w_dff_B_rYsrBV0W6_1;
	wire w_dff_B_e8li2tLE4_1;
	wire w_dff_B_5urLXsyC3_0;
	wire w_dff_B_G1whR9533_1;
	wire w_dff_B_yt8yq8iV8_1;
	wire w_dff_B_ckbM7ytb5_0;
	wire w_dff_B_35ZYj0rt8_1;
	wire w_dff_B_4hGgm3Et5_1;
	wire w_dff_B_lMbt7F9W4_0;
	wire w_dff_B_XDdD7kux4_1;
	wire w_dff_B_koWa50FX4_1;
	wire w_dff_B_qygv1SxQ7_0;
	wire w_dff_B_HMAOWoZm1_1;
	wire w_dff_B_emjTCb4j0_1;
	wire w_dff_B_i5x16gKI7_0;
	wire w_dff_B_VchOax7E1_1;
	wire w_dff_B_1dMdFzNe2_1;
	wire w_dff_B_F4EsfGDJ5_0;
	wire w_dff_B_uBXblJmV0_1;
	wire w_dff_B_MXNCDc511_1;
	wire w_dff_B_c0oDU8DR9_0;
	wire w_dff_B_CMZG07on5_1;
	wire w_dff_B_oaC8QtX88_1;
	wire w_dff_B_1GbEw4ra1_0;
	wire w_dff_B_J8H21Ve13_1;
	wire w_dff_B_zMcDdjhX8_1;
	wire w_dff_B_nrM5oNz77_0;
	wire w_dff_B_xentm9ut9_1;
	wire w_dff_B_qvsR5x1d9_1;
	wire w_dff_B_9vGQxAeC7_0;
	wire w_dff_B_116dGzVJ3_1;
	wire w_dff_B_NPGtS0aV6_1;
	wire w_dff_B_8IFA9uxn4_0;
	wire w_dff_B_ecb1o3A97_1;
	wire w_dff_B_LLMoJvwo6_1;
	wire w_dff_B_nuqFSaDm4_0;
	wire w_dff_B_9ymwhC0x0_1;
	wire w_dff_B_robiVxRf4_1;
	wire w_dff_B_OGeIt0NV8_0;
	wire w_dff_B_iE2eMepW7_1;
	wire w_dff_B_cP0exCf09_1;
	wire w_dff_B_g96jNHdJ1_0;
	wire w_dff_B_dBor2d8J6_1;
	wire w_dff_B_ETLDoBFx5_1;
	wire w_dff_B_h1n7C7xB6_0;
	wire w_dff_B_bimxITUi8_1;
	wire w_dff_B_55Edj9Zy7_1;
	wire w_dff_B_NmnoyRaM2_0;
	wire w_dff_B_zNZVTUNb4_1;
	wire w_dff_B_2a5xp3cf3_1;
	wire w_dff_B_m1xLLlKS6_0;
	wire w_dff_B_gs2vDvNb3_1;
	wire w_dff_B_Mfbpq3wo7_1;
	wire w_dff_B_BVk4GIky4_0;
	wire w_dff_B_bLoygNGB6_1;
	wire w_dff_B_hOzIDkh54_1;
	wire w_dff_B_fhJ1mx9l9_0;
	wire w_dff_B_zlxKaspI7_1;
	wire w_dff_B_xuIIATgQ1_1;
	wire w_dff_B_SZs8Qcod0_0;
	wire w_dff_B_PYWeaYGl5_1;
	wire w_dff_B_KLVuGhgh7_1;
	wire w_dff_B_enD4tXYE6_0;
	wire w_dff_B_hCq4zkgr3_1;
	wire w_dff_B_UhGdGDuw2_1;
	wire w_dff_B_Sbji6ZfD0_0;
	wire w_dff_B_j9l6F43z2_1;
	wire w_dff_B_PRxlyw9O6_1;
	wire w_dff_B_OcNBDkyx2_0;
	wire w_dff_B_EFRg9bZf6_1;
	wire w_dff_B_qCuGtxRb1_1;
	wire w_dff_B_o8z0a3BH8_0;
	wire w_dff_B_Vvjm6PZZ6_1;
	wire w_dff_B_ipvPNgWN6_1;
	wire w_dff_B_IfHCHb0m5_0;
	wire w_dff_B_m0ZRsxqR5_1;
	wire w_dff_B_1rfsyViv6_1;
	wire w_dff_B_BoPmVl8N6_0;
	wire w_dff_B_Qo4ZEKl62_1;
	wire w_dff_B_ShHJJsvM6_1;
	wire w_dff_B_8LcbiD876_0;
	wire w_dff_B_61TsfZBo0_1;
	wire w_dff_B_H5LQYE1i4_1;
	wire w_dff_B_ZV0RQbIM7_0;
	wire w_dff_B_IN0A43qU2_1;
	wire w_dff_B_DNWcCaNq6_1;
	wire w_dff_B_WKMYwIeP6_0;
	wire w_dff_B_9Yjqugh99_1;
	wire w_dff_B_wMTGnKcB8_1;
	wire w_dff_B_wQeft8uk8_0;
	wire w_dff_B_vsZalWtc9_1;
	wire w_dff_B_reajkNSh8_1;
	wire w_dff_B_nGRQaI5L2_0;
	wire w_dff_B_ZeRdUNCn5_1;
	wire w_dff_B_vqYPtKNk8_1;
	wire w_dff_B_bAkFKoGi1_0;
	wire w_dff_B_mD3g0jyP8_1;
	wire w_dff_B_QbZh5GTu1_1;
	wire w_dff_B_bvqaMLGq4_0;
	wire w_dff_B_dwolWk1u4_1;
	wire w_dff_B_aJJeIIHt4_1;
	wire w_dff_B_CzywkDtF3_0;
	wire w_dff_B_3VkjLdoL6_1;
	wire w_dff_B_VTYfoZ241_1;
	wire w_dff_B_YX9OTQX74_0;
	wire w_dff_B_RKy8dYIb6_1;
	wire w_dff_B_hCssqM0Q9_1;
	wire w_dff_B_rl1ZH6TR5_0;
	wire w_dff_B_dEI03NQy2_1;
	wire w_dff_B_qJOt6bhg1_1;
	wire w_dff_B_dV3x719y6_0;
	wire w_dff_B_4wh24KR08_1;
	wire w_dff_B_G4Ih9Qr33_1;
	wire w_dff_B_Oi4X5sPK9_0;
	wire w_dff_B_pn4CGLHa1_1;
	wire w_dff_B_UQHrQaep4_1;
	wire w_dff_B_bc3S7ENI2_0;
	wire w_dff_B_KP72rsrz6_1;
	wire w_dff_B_7yGKMDYQ1_1;
	wire w_dff_B_wTfreXba5_0;
	wire w_dff_B_euyAe64v7_1;
	wire w_dff_B_xTJkLHWE4_1;
	wire w_dff_B_Xvu7oEBw8_0;
	wire w_dff_B_yYkEEkM38_1;
	wire w_dff_B_WHlDTliR9_1;
	wire w_dff_B_Bh0cWlsK3_0;
	wire w_dff_B_6a8xIgi53_1;
	wire w_dff_B_2kENvoBC8_1;
	wire w_dff_B_0uemW6GM9_0;
	wire w_dff_B_Y5BvixUE0_1;
	wire w_dff_B_8SRP66dE1_1;
	wire w_dff_B_GNedNEEq9_0;
	wire w_dff_B_uYRKYk1g1_1;
	wire w_dff_B_eD6zHKXZ0_1;
	wire w_dff_B_McwzmPqr1_0;
	wire w_dff_B_uoF5tk2m6_1;
	wire w_dff_B_h3eJu9OU0_1;
	wire w_dff_B_u47osZBz0_0;
	wire w_dff_B_Q4JjspNz1_1;
	wire w_dff_B_ywtVITPN8_1;
	wire w_dff_B_oYfAcDzV7_0;
	wire w_dff_B_rHT2H57k2_1;
	wire w_dff_B_otiiGruG4_1;
	wire w_dff_B_rGaC2c9d4_0;
	wire w_dff_B_W01oYgIo0_1;
	wire w_dff_B_6L9GTXRb7_1;
	wire w_dff_B_SqgF1FXp2_0;
	wire w_dff_B_zcrvu5Ei2_1;
	wire w_dff_B_uHPHRthA7_1;
	wire w_dff_B_rkzRbhOh1_0;
	wire w_dff_B_6bzhAcri5_1;
	wire w_dff_B_99mKSXMI6_1;
	wire w_dff_B_dk5lNsOw9_0;
	wire w_dff_B_aJNLwn6g4_1;
	wire w_dff_B_liuz3nrk5_1;
	wire w_dff_B_H5CDb6oE6_0;
	wire w_dff_B_Hb9wmUcB0_1;
	wire w_dff_B_KAogdi844_1;
	wire w_dff_B_SGLp9wMj4_0;
	wire w_dff_B_GHCPb6rq3_1;
	wire w_dff_B_DnS9XDKT8_1;
	wire w_dff_B_M6qUBrYh2_0;
	wire w_dff_B_DQwxqxQg4_1;
	wire w_dff_B_MG0suzb56_1;
	wire w_dff_B_RgGRMQHE6_0;
	wire w_dff_B_kJ3dij4h6_1;
	wire w_dff_B_9qAu6CEv6_1;
	wire w_dff_B_lNX9XknG9_0;
	wire w_dff_B_uOv1uSkF3_1;
	wire w_dff_B_D9FffPJm6_1;
	wire w_dff_B_q2S1c17p8_0;
	wire w_dff_B_rjprWWua0_1;
	wire w_dff_B_yVPVbjPP6_1;
	wire w_dff_B_9iVsnI3Y0_0;
	wire w_dff_B_Ho3L4MC88_1;
	wire w_dff_B_a3CGe7202_1;
	wire w_dff_B_bTy0068r1_0;
	wire w_dff_B_PjliAp9l8_1;
	wire w_dff_B_19lEeWUB7_1;
	wire w_dff_B_7kVOx8kZ8_0;
	wire w_dff_B_qmiGF2fS5_1;
	wire w_dff_B_7HQfPZQp1_1;
	wire w_dff_B_boPyw8vw4_0;
	wire w_dff_B_YHhQGkIh3_1;
	wire w_dff_B_ky9JnIJa0_1;
	wire w_dff_B_YFkbXwkf8_0;
	wire w_dff_B_8PGIHgI10_1;
	wire w_dff_B_FwE6F5NN2_1;
	wire w_dff_B_9obNFDpn5_0;
	wire w_dff_B_muxmvvbB9_1;
	wire w_dff_B_4eITFKR93_1;
	wire w_dff_B_YdezcyHU5_0;
	wire w_dff_B_Fjv5O2Ty2_1;
	wire w_dff_B_f6wrL0AW5_1;
	wire w_dff_B_0hEDWuI26_0;
	wire w_dff_B_jM0CcFoY3_1;
	wire w_dff_B_0Z3CSdIH1_1;
	wire w_dff_B_qB6dFw1e2_0;
	wire w_dff_B_H34hZ62M9_1;
	wire w_dff_B_f4xDkURy7_1;
	wire w_dff_B_u3F8t7vU1_0;
	wire w_dff_B_1MNqUUdQ1_1;
	wire w_dff_B_OQ4nf9FB4_1;
	wire w_dff_B_huflLVnU8_0;
	wire w_dff_B_BrGOasGm4_1;
	wire w_dff_B_N2r3icPs2_1;
	wire w_dff_B_X8hTW4sa2_0;
	wire w_dff_B_QbSsgr8h7_1;
	wire w_dff_B_nr95JRAm8_1;
	wire w_dff_B_aEdf5wZc7_0;
	wire w_dff_B_zI2Kpgg59_1;
	wire w_dff_B_nkiDrsDo7_1;
	wire w_dff_B_C34EYOny8_0;
	wire w_dff_B_z59wLket6_1;
	wire w_dff_B_b7uSIuaZ4_1;
	wire w_dff_B_YWRYZVvo7_0;
	wire w_dff_B_rZQte5bu0_1;
	wire w_dff_B_CrXB06rb5_1;
	wire w_dff_B_496Qayul4_0;
	wire w_dff_B_TbgNN2S95_1;
	wire w_dff_B_V9UeSrPZ8_1;
	wire w_dff_B_gh9Bjk4K5_0;
	wire w_dff_B_3X0mNpgI5_1;
	wire w_dff_B_uj3d5Aa12_1;
	wire w_dff_B_Onbv6u1X0_0;
	wire w_dff_B_sr510KQA8_1;
	wire w_dff_B_edIm3HEo0_1;
	wire w_dff_B_ocQxDi7i4_0;
	wire w_dff_B_CTjIjAr87_1;
	wire w_dff_B_Sy8fXmtO9_1;
	wire w_dff_B_ZqWDHNKl8_0;
	wire w_dff_B_xoKU3Id01_1;
	wire w_dff_B_SBRBhiff0_1;
	wire w_dff_B_rW47TtDh5_0;
	wire w_dff_B_bfjtPOIV7_1;
	wire w_dff_B_4prvR3SB9_1;
	wire w_dff_B_ujybVo5m3_0;
	wire w_dff_B_T8PVOLJC4_1;
	wire w_dff_B_nh3K4oM22_1;
	wire w_dff_B_AJta4V6q0_0;
	wire w_dff_B_sZXkuFTi7_1;
	wire w_dff_B_43izO5SG7_1;
	wire w_dff_B_x80yLBcc3_0;
	wire w_dff_B_KAgkIkQn7_1;
	wire w_dff_B_UO0r7WtK8_1;
	wire w_dff_B_4o1boigc1_0;
	wire w_dff_B_Ys0zWwiN3_1;
	wire w_dff_B_tFBmKSHU9_1;
	wire w_dff_B_A0PnvmfU3_0;
	wire w_dff_B_20SCvLSX5_1;
	wire w_dff_B_8tVKfkLJ8_1;
	wire w_dff_B_YxqWpnGO2_0;
	wire w_dff_B_JeoVcAtz5_1;
	wire w_dff_B_DbMsD6I55_1;
	wire w_dff_B_0BpUHJ8f5_0;
	wire w_dff_B_sIRvNoS55_1;
	wire w_dff_B_wOKdUDwI7_1;
	wire w_dff_B_jFPT1jCW9_0;
	wire w_dff_B_gLUxUchn8_1;
	wire w_dff_B_TEUMczxJ9_1;
	wire w_dff_B_3WWymGYL5_0;
	wire w_dff_B_AgREMfxR4_1;
	wire w_dff_B_kLVUkxdA1_1;
	wire w_dff_B_iXl7YkEZ9_0;
	wire w_dff_B_X3cYN9Mx0_1;
	wire w_dff_B_4gZnAB7L0_1;
	wire w_dff_B_JOnwcef08_0;
	wire w_dff_B_FephHzNx3_1;
	wire w_dff_B_feWNsbf75_1;
	wire w_dff_B_cjjRtxAq5_0;
	wire w_dff_B_uhfGFFCT8_1;
	wire w_dff_B_3JQdqvgr9_1;
	wire w_dff_B_i4pJGpHe3_0;
	wire w_dff_B_focNT7rN2_1;
	wire w_dff_B_9yHQ4G319_1;
	wire w_dff_B_J66uxfix0_0;
	wire w_dff_B_MKxh3gBh9_1;
	wire w_dff_B_wrKJCLHE2_1;
	wire w_dff_B_WaH1Qvu22_0;
	wire w_dff_B_kWkTLlgn2_1;
	wire w_dff_B_zEG94JNY7_1;
	wire w_dff_B_YzMLCC1i0_0;
	wire w_dff_B_UZmCgTSI6_1;
	wire w_dff_B_cZrHVwDG1_1;
	wire w_dff_B_9CCHJG3I8_0;
	wire w_dff_B_VuxjLPID6_1;
	wire w_dff_B_T9dm59OW2_1;
	wire w_dff_B_PoFkE5wX0_0;
	wire w_dff_B_xGeMO9BU0_1;
	wire w_dff_B_faRWqwxy6_1;
	wire w_dff_B_TkhLCRu23_0;
	wire w_dff_B_a0UUqY5s8_1;
	wire w_dff_B_ENIICq2y3_1;
	wire w_dff_B_GF88rIeY2_0;
	wire w_dff_B_IuTIilJs1_1;
	wire w_dff_B_BFVo2AC79_1;
	wire w_dff_B_AsSN8oxv0_0;
	wire w_dff_B_2WZlsVjY4_1;
	wire w_dff_B_T0GGtFnc1_1;
	wire w_dff_B_jeXu3sy45_0;
	wire w_dff_B_kkOZ5FN67_1;
	wire w_dff_B_5U4XzmXQ9_1;
	wire w_dff_B_poR6M3NX3_0;
	wire w_dff_B_FSunM1fL8_1;
	wire w_dff_B_Mx9XTvKw1_1;
	wire w_dff_B_XJJ0p5Hv1_0;
	wire w_dff_B_kRocFKSE5_1;
	wire w_dff_B_pD3SBYZu7_1;
	wire w_dff_B_R3YJSblS2_0;
	wire w_dff_B_UM9TQzFB4_1;
	wire w_dff_B_NPOXfZNT9_1;
	wire w_dff_B_kk7LeyAl5_0;
	wire w_dff_B_egJRPEu89_1;
	wire w_dff_B_pWTH2BSY6_1;
	wire w_dff_B_MoX53rZY3_0;
	wire w_dff_B_dE1wqsEz3_1;
	wire w_dff_B_EhiM211Y3_1;
	wire w_dff_B_rOHLQUyL7_0;
	wire w_dff_B_Dq3Q0i4O2_1;
	wire w_dff_B_HBaastiB7_1;
	wire w_dff_B_RbwjiVQc5_0;
	wire w_dff_B_YfL9hMuc0_1;
	wire w_dff_B_fvmWPNeu8_1;
	wire w_dff_B_56NlZhYE3_0;
	wire w_dff_B_MIhQQiDJ8_1;
	wire w_dff_B_n4s9MQBi8_1;
	wire w_dff_B_Tp0JK1jz6_0;
	wire w_dff_B_0j7GEJgP0_1;
	wire w_dff_B_h6gd19k23_1;
	wire w_dff_B_YOJR5kVR6_0;
	wire w_dff_B_UDDJjihN1_1;
	wire w_dff_B_CJe3LNGD1_1;
	wire w_dff_B_YCE8fMWj4_0;
	wire w_dff_B_cpHbBKmC5_1;
	wire w_dff_B_ZhWqQhPZ3_1;
	wire w_dff_B_ZGWEitvM6_0;
	wire w_dff_B_yRqUJEnE2_1;
	wire w_dff_B_sQ1XAWmU2_1;
	wire w_dff_B_aeg3cgRf4_0;
	wire w_dff_B_iDyOIIGT5_1;
	wire w_dff_B_oMk1KklB2_1;
	wire w_dff_B_hh4D6Ws52_0;
	wire w_dff_B_3iGzd9JX6_1;
	wire w_dff_B_n9pUpmqm8_1;
	wire w_dff_B_qG7CcZVr6_0;
	wire w_dff_B_6A2FPn0t3_1;
	wire w_dff_B_gws8z3LA1_1;
	wire w_dff_B_5ldzfQYi3_0;
	wire w_dff_B_MaGlQa950_1;
	wire w_dff_B_3KDdwdBk3_1;
	wire w_dff_B_xnBRSN2N3_0;
	wire w_dff_B_djcKn61M3_1;
	wire w_dff_B_wnQLWcq32_1;
	wire w_dff_B_BlDVNLBK7_0;
	wire w_dff_B_WOEkBFSe2_1;
	wire w_dff_B_4OEclSdP1_1;
	wire w_dff_B_vGLAXmG71_0;
	wire w_dff_B_9RJGWIrd7_1;
	wire w_dff_B_XrRsKiC06_1;
	wire w_dff_B_B3HjuQuU9_0;
	wire w_dff_B_FZxU42WT4_1;
	wire w_dff_B_y7xezhI94_1;
	wire w_dff_B_hGQAN2Ud3_0;
	wire w_dff_B_mUIeIU2P5_1;
	wire w_dff_B_v6S0pnWU5_1;
	wire w_dff_B_bxZjKYFc1_0;
	wire w_dff_B_hBgbUGtR7_1;
	wire w_dff_B_6KHWH1Jh5_1;
	wire w_dff_B_xB4q2Qjw2_0;
	wire w_dff_B_YUDdw4H56_1;
	wire w_dff_B_L4laJNFt4_1;
	wire w_dff_B_NyFPXIyr2_0;
	wire w_dff_B_T1FtALzk3_1;
	wire w_dff_B_VMQQNRP08_1;
	wire w_dff_B_SOdTOQwU7_0;
	wire w_dff_B_86vXx9XN1_1;
	wire w_dff_B_vvMFgqlf6_1;
	wire w_dff_B_B2NxBOMf3_0;
	wire w_dff_B_GxdybRXV1_1;
	wire w_dff_B_82FVcnT81_1;
	wire w_dff_B_t5k4kQhB6_0;
	wire w_dff_B_cBR00QJg3_1;
	wire w_dff_B_ycfnNlTi5_1;
	wire w_dff_B_hZx5Rp366_0;
	wire w_dff_B_6ZMF23I40_1;
	wire w_dff_B_VGg8A4KJ8_1;
	wire w_dff_B_Qp7R6Ppv0_0;
	wire w_dff_B_rBcQrI584_1;
	wire w_dff_B_GEI0pHLe2_1;
	wire w_dff_B_7IMUWZDl2_0;
	wire w_dff_B_9QCGOelP1_1;
	wire w_dff_B_bz9R4FL06_1;
	wire w_dff_B_1DoTDJze9_0;
	wire w_dff_B_tcxmG4DG5_1;
	wire w_dff_B_StgGyzNM1_1;
	wire w_dff_B_hknLRKEp8_0;
	wire w_dff_B_d95Y6bnw1_1;
	wire w_dff_B_gfiTS28a2_1;
	wire w_dff_B_1OEUfKzK8_0;
	wire w_dff_B_gO2pJsJg3_1;
	wire w_dff_B_EtA1Bwgh7_1;
	wire w_dff_B_Yji0C1js9_0;
	wire w_dff_B_4bWQ8Y4U4_1;
	wire w_dff_B_IEnkpo8q6_1;
	wire w_dff_B_IHsLOWpC2_0;
	wire w_dff_B_Onbogkyx1_1;
	wire w_dff_B_DD4YCshY8_1;
	wire w_dff_B_RWQCZSD81_0;
	wire w_dff_B_kDPvPpoP4_1;
	wire w_dff_B_wO6CPyKc2_1;
	wire w_dff_B_70rd1kZT3_0;
	wire w_dff_B_rzbj5T0z1_1;
	wire w_dff_B_EMAK944C1_1;
	wire w_dff_B_PIEA6oQH3_0;
	wire w_dff_B_IFtLjBZF6_1;
	wire w_dff_B_Y9K3ClDR7_1;
	wire w_dff_B_8BngNbgd0_0;
	wire w_dff_B_I7aht90O4_1;
	wire w_dff_B_3wuBCOe82_1;
	wire w_dff_B_mfvk1noa9_0;
	wire w_dff_B_98IgX14T0_1;
	wire w_dff_B_O9cfa67M4_1;
	wire w_dff_B_LuB7p5DQ9_0;
	wire w_dff_B_Djzz0kY27_1;
	wire w_dff_B_ObVd5VZ58_1;
	wire w_dff_B_z89m836x9_0;
	wire w_dff_B_okhOeJHm0_1;
	wire w_dff_B_KrkdkH7l9_1;
	wire w_dff_B_iymvmlfM2_0;
	wire w_dff_B_QmqB7p2U9_1;
	wire w_dff_B_QwBaURrl5_1;
	wire w_dff_B_D9fLjXBM7_0;
	wire w_dff_B_1ZtuVlls5_1;
	wire w_dff_B_FRrwnx3T2_1;
	wire w_dff_B_7Xuq5K5W5_0;
	wire w_dff_B_3k65QdRj2_1;
	wire w_dff_B_XnPkPJHe3_1;
	wire w_dff_B_RAvhSOHM5_0;
	wire w_dff_B_1pacFc5A9_1;
	wire w_dff_B_yogMl37H5_1;
	wire w_dff_B_DqhQ5BMC9_0;
	wire w_dff_B_uet8h9lm8_1;
	wire w_dff_B_hozR8B1v3_1;
	wire w_dff_B_FQAQqQ3K2_0;
	wire w_dff_B_61j1RiBO5_1;
	wire w_dff_B_V651QdOo9_1;
	wire w_dff_B_4FGpBViq2_0;
	wire w_dff_B_9fZ3rJLb9_1;
	wire w_dff_B_r38PTKb32_1;
	wire w_dff_B_49MrkuEv1_0;
	wire w_dff_B_dswNJH0Q3_1;
	wire w_dff_B_HZGcZQx65_1;
	wire w_dff_B_HuZqe8R86_0;
	wire w_dff_B_5z6ntGRA1_1;
	wire w_dff_B_LnFLsAV69_1;
	wire w_dff_B_XQRJK8hI2_0;
	wire w_dff_B_3YFfs46K3_1;
	wire w_dff_B_FMefJS5z4_1;
	wire w_dff_B_ldonzCFe9_0;
	wire w_dff_B_V5RqNucF7_1;
	wire w_dff_B_Y88xVshG7_1;
	wire w_dff_B_FHH2yJSp7_0;
	wire w_dff_B_HrXKvA0r3_1;
	wire w_dff_B_3p3FQbxZ2_1;
	wire w_dff_B_FDc46lRH6_0;
	wire w_dff_B_QI6jOKro7_1;
	wire w_dff_B_CBcSyyyU8_1;
	wire w_dff_B_JNJO4QOP3_0;
	wire w_dff_B_q2uZc8Gj9_1;
	wire w_dff_B_qYzkE5Ne5_1;
	wire w_dff_B_7JX91FRK1_0;
	wire w_dff_B_pVLlfeWJ1_1;
	wire w_dff_B_JL4G19Qr8_1;
	wire w_dff_B_yYHiuxfW3_0;
	wire w_dff_B_6w4rnDi74_1;
	wire w_dff_B_QeKRpaxT3_1;
	wire w_dff_B_KwAJ2y101_0;
	wire w_dff_B_hWACObTH0_1;
	wire w_dff_B_ZHHldruu7_1;
	wire w_dff_B_hTzDDnzK8_0;
	wire w_dff_B_cnGtcmvV7_1;
	wire w_dff_B_HugGMlsl5_1;
	wire w_dff_B_yoRicxHq6_0;
	wire w_dff_B_Yp5MvGc20_1;
	wire w_dff_B_fkSCvyox5_1;
	wire w_dff_B_LderWme62_0;
	wire w_dff_B_ql79bxwE5_1;
	wire w_dff_B_Dr5Rgvhi0_1;
	wire w_dff_B_4lNWY1Cp4_0;
	wire w_dff_B_ZJ7t2wem9_1;
	wire w_dff_B_qU6FUjGM9_1;
	wire w_dff_B_PjZlxOwU2_0;
	wire w_dff_B_pcpEuBTO7_1;
	wire w_dff_B_ZRpp3rBP5_1;
	wire w_dff_B_D3k26w8o6_0;
	wire w_dff_B_LCRp0Mdl8_1;
	wire w_dff_B_l9iXkasH1_1;
	wire w_dff_B_znXfgxXr4_0;
	wire w_dff_B_vzerBgVm3_1;
	wire w_dff_B_m13q85Av4_1;
	wire w_dff_B_CGPI3dHX3_0;
	wire w_dff_B_4rpiYas84_1;
	wire w_dff_B_ZxgD49R90_1;
	wire w_dff_B_jew2rhCp7_0;
	wire w_dff_B_N8RSnojY1_1;
	wire w_dff_B_qvZOCGkh7_1;
	wire w_dff_B_K6ULNMp38_0;
	wire w_dff_B_A6DxkfPQ0_1;
	wire w_dff_B_ykEXxVEF6_1;
	wire w_dff_B_ZGsJLjTO8_0;
	wire w_dff_B_cryE1Kd60_1;
	wire w_dff_B_9liRMWfx0_1;
	wire w_dff_B_vqKakcLX8_0;
	wire w_dff_B_tl3HbU9G6_1;
	wire w_dff_B_aGDLZ7hj2_1;
	wire w_dff_B_qHBfuMtU9_0;
	wire w_dff_B_EZu2XAm08_1;
	wire w_dff_B_WSOvahUp7_1;
	wire w_dff_B_YOOdvGcg9_0;
	wire w_dff_B_8wkgG7hP0_1;
	wire w_dff_B_f0Wxj4yd8_1;
	wire w_dff_B_yLZkh10I4_0;
	wire w_dff_B_CGqmudAv9_1;
	wire w_dff_B_lhOl7scJ0_1;
	wire w_dff_B_c2phCQGi0_0;
	wire w_dff_B_2YQMWR6R4_1;
	wire w_dff_B_QBBmk80V1_1;
	wire w_dff_B_U4CRJqxg3_0;
	wire w_dff_B_BJhaO4Sm1_1;
	wire w_dff_B_fPXeCm1I9_1;
	wire w_dff_B_GJ9JITL81_0;
	wire w_dff_B_CXBZKziI3_1;
	wire w_dff_B_9A8x5XsH6_1;
	wire w_dff_B_yS8ELcW17_0;
	wire w_dff_B_mfY5h3s66_1;
	wire w_dff_B_m7kHuDJE5_1;
	wire w_dff_B_fPFHHo2p6_0;
	wire w_dff_B_TbHcYDTX8_1;
	wire w_dff_B_OZhIiuq18_1;
	wire w_dff_B_ZgZcwHQk4_0;
	wire w_dff_B_l03Q91CO4_1;
	wire w_dff_B_FiNXkb9Y6_1;
	wire w_dff_B_02mnb2b89_0;
	wire w_dff_B_aui4nqcb5_1;
	wire w_dff_B_RIw4JiM62_1;
	wire w_dff_B_aQl6SJho8_0;
	wire w_dff_B_1ALoBJ3i8_1;
	wire w_dff_B_PPfha8iG0_1;
	wire w_dff_B_t7mqydWt3_0;
	wire w_dff_B_cZyPlB1Q5_1;
	wire w_dff_B_OSsMJ08H1_1;
	wire w_dff_B_L33fN8wm0_0;
	wire w_dff_B_LseYXHtZ6_1;
	wire w_dff_B_Vexy9pSD4_1;
	wire w_dff_B_PEtYO2nZ2_0;
	wire w_dff_B_ojgVuRDt2_1;
	wire w_dff_B_iuUN1MS12_1;
	wire w_dff_B_DXN0HrMN5_0;
	wire w_dff_B_t1LazA034_1;
	wire w_dff_B_Fg5kkHG93_1;
	wire w_dff_B_kjyfZ68B8_0;
	wire w_dff_B_QWQqj8xb4_1;
	wire w_dff_B_XgKuybAs2_1;
	wire w_dff_B_N0xQg3RU2_0;
	wire w_dff_B_DtzcDB6d0_1;
	wire w_dff_B_3w20PdWI5_1;
	wire w_dff_B_0KacSSWA2_0;
	wire w_dff_B_VnJASxDh2_1;
	wire w_dff_B_LOWVhPMa9_1;
	wire w_dff_B_K2r8C8Bi4_0;
	wire w_dff_B_0RpO4pcF0_1;
	wire w_dff_B_vZrVtr4g8_1;
	wire w_dff_B_aP2Vzczj8_0;
	wire w_dff_B_FPwWCjoV9_1;
	wire w_dff_B_buHD2ggE4_1;
	wire w_dff_B_XBiAr6HB6_0;
	wire w_dff_B_PCbR2CMZ5_1;
	wire w_dff_B_vFRPZe0E7_1;
	wire w_dff_B_lFefcJ9l1_0;
	wire w_dff_B_pgKvcWnY5_1;
	wire w_dff_B_Fa5UygcP0_1;
	wire w_dff_B_nUofu0Ki0_0;
	wire w_dff_B_nyJTp72i1_1;
	wire w_dff_B_ZIGeXFC22_1;
	wire w_dff_B_iXUqkg6b0_0;
	wire w_dff_B_ySBpqbGv9_1;
	wire w_dff_B_QmpjNxjn9_1;
	wire w_dff_B_XA3R5mLm5_0;
	wire w_dff_B_szz47Hzv6_1;
	wire w_dff_B_iky6qif53_1;
	wire w_dff_B_1jugmf9a1_0;
	wire w_dff_B_22ihCfHP1_1;
	wire w_dff_B_Z0mTHOxn2_1;
	wire w_dff_B_XXULzUgH7_0;
	wire w_dff_B_iCqvrP4J6_1;
	wire w_dff_B_BBYKbmq80_1;
	wire w_dff_B_bqScnAXr8_0;
	wire w_dff_B_xxdAL6Gg1_1;
	wire w_dff_B_ICBxgeIV7_1;
	wire w_dff_B_YljleBFN9_0;
	wire w_dff_B_V7meLCNO7_1;
	wire w_dff_B_12bjiM417_1;
	wire w_dff_B_WWcxEztL0_0;
	wire w_dff_B_5rVmUIn50_1;
	wire w_dff_B_FCK49IvL3_1;
	wire w_dff_B_a27ha2GA3_0;
	wire w_dff_B_ucTIwyaU5_1;
	wire w_dff_B_z6Mk3N4z7_1;
	wire w_dff_B_CwRb6Zdg9_0;
	wire w_dff_B_M7HzpFLq5_1;
	wire w_dff_B_cC9wJqdw1_1;
	wire w_dff_B_u3s452In8_0;
	wire w_dff_B_GWN1KlHz0_1;
	wire w_dff_B_8sKYsfXN5_1;
	wire w_dff_B_qzNhIp991_0;
	wire w_dff_B_Ur6ue7jr2_1;
	wire w_dff_B_BhqJTvgw6_1;
	wire w_dff_B_6p5HSVjj5_0;
	wire w_dff_B_OyEk1U2B4_1;
	wire w_dff_B_wM0cwS0E2_1;
	wire w_dff_B_eFTihvvF4_0;
	wire w_dff_B_4rqFI4Gy5_1;
	wire w_dff_B_mQYVjC3V5_1;
	wire w_dff_B_W1m7NuUn4_0;
	wire w_dff_B_z3S3oK5g3_1;
	wire w_dff_B_U7tofJv50_1;
	wire w_dff_B_LXLqwXQf5_0;
	wire w_dff_B_NPxcAtcs0_1;
	wire w_dff_B_NGb1Pgpk3_1;
	wire w_dff_B_vaIk44ui8_0;
	wire w_dff_B_SW6s5Ekj1_1;
	wire w_dff_B_HWXL2sOJ4_1;
	wire w_dff_B_IpfWp5MV0_0;
	wire w_dff_B_gSBDtJ4S1_1;
	wire w_dff_B_0KDHoTdV3_1;
	wire w_dff_B_fOzLotLx0_0;
	wire w_dff_B_m2ferJHn8_1;
	wire w_dff_B_HYrPEvnV5_1;
	wire w_dff_B_osWnsPAs4_0;
	wire w_dff_B_zRQsCoKt9_1;
	wire w_dff_B_vVdaNbcH6_1;
	wire w_dff_B_EyWT0czp2_0;
	wire w_dff_B_pTGLz1Ga5_1;
	wire w_dff_B_BUCvsxNO3_1;
	wire w_dff_B_lnxYEnyW2_0;
	wire w_dff_B_WVMYNQRc8_1;
	wire w_dff_B_EQkAxmtM8_1;
	wire w_dff_B_g3hpVPxg1_0;
	wire w_dff_B_L2tsbO6u6_1;
	wire w_dff_B_75VVNHvJ2_1;
	wire w_dff_B_UgfuBzO50_0;
	wire w_dff_B_6uroEMmR5_1;
	wire w_dff_B_Y7YtLhzO6_1;
	wire w_dff_B_D38jD0K72_0;
	wire w_dff_B_AQTDvday7_1;
	wire w_dff_B_lH0Rc6Lf0_1;
	wire w_dff_B_U5D9P6Db9_0;
	wire w_dff_B_mUqQUmBj9_1;
	wire w_dff_B_JqSHsLGG2_1;
	wire w_dff_B_id4K03Wa5_0;
	wire w_dff_B_jMNibkDP1_1;
	wire w_dff_B_6iCFG5SY4_1;
	wire w_dff_B_l2iJDWqD9_0;
	wire w_dff_B_RE1qjwxi1_1;
	wire w_dff_B_174ZvsxD2_1;
	wire w_dff_B_Tg33vzS97_0;
	wire w_dff_B_Sdr4G0ZW3_1;
	wire w_dff_B_h8DUDHPi9_1;
	wire w_dff_B_92yjbt7N5_0;
	wire w_dff_B_gXXxnHFS1_1;
	wire w_dff_B_slVYtXoH6_1;
	wire w_dff_B_zURs38kR5_0;
	wire w_dff_B_0I265xjZ5_1;
	wire w_dff_B_MNkhRkVJ2_1;
	wire w_dff_B_mNvo9h4e6_0;
	wire w_dff_B_HegFkakD8_1;
	wire w_dff_B_tbWgCQ7T5_1;
	wire w_dff_B_0gJiH3OV1_0;
	wire w_dff_B_Bb2LQOX46_1;
	wire w_dff_B_VbO6w6zD2_1;
	wire w_dff_B_3s6AjRKb2_0;
	wire w_dff_B_0f5VWSQ93_1;
	wire w_dff_B_Z7fK2rF58_1;
	wire w_dff_B_M8RJIFvs4_0;
	wire w_dff_B_T1dMgkpZ6_1;
	wire w_dff_B_rD7Jx1Kl7_1;
	wire w_dff_B_Q96lHp3o5_0;
	wire w_dff_B_xoinFbqO8_1;
	wire w_dff_B_yEJJMF8P9_1;
	wire w_dff_B_m0Sng1PW4_0;
	wire w_dff_B_MdIApfCQ7_1;
	wire w_dff_B_46as8xFJ1_1;
	wire w_dff_B_JGDoXU1T7_0;
	wire w_dff_B_8SdLIGhZ4_1;
	wire w_dff_B_sqwDOK3F5_1;
	wire w_dff_B_wXVKtnh13_1;
	wire w_dff_B_jlhhO1862_1;
	wire w_dff_B_xqLjxEhE3_1;
	wire w_dff_B_gnnLsEbL7_1;
	wire w_dff_B_LvNxJLXv2_1;
	wire w_dff_B_1erSQF5v5_1;
	wire w_dff_B_73zz0aOP0_1;
	wire w_dff_B_kx18ekQ99_1;
	wire w_dff_B_PVvmUK9a6_0;
	wire w_dff_B_RDrOvlHB2_1;
	wire w_dff_B_lrsiFJkx2_1;
	wire w_dff_B_3XYmQ7xa1_1;
	wire w_dff_B_kbso0kek4_1;
	wire w_dff_B_a2qEd9k26_1;
	wire w_dff_B_KkZUlkQY5_1;
	wire w_dff_B_gUpOzecm7_1;
	wire w_dff_B_qDiElXBG9_1;
	wire w_dff_B_peT3tE445_1;
	wire w_dff_B_FFv3MKX02_1;
	wire w_dff_B_0oY8yfNB8_0;
	wire w_dff_B_USEsFc4E6_1;
	wire w_dff_B_qxZUuMrc2_1;
	wire w_dff_B_bUuUbKk52_1;
	wire w_dff_B_0JQMoqEd2_1;
	wire w_dff_B_DBajLoEy0_1;
	wire w_dff_B_oANUBuw89_1;
	wire w_dff_B_ZtYCSpfs0_1;
	wire w_dff_B_kMwsZSDe0_1;
	wire w_dff_B_v0bLqLBi4_1;
	wire w_dff_B_pvT9nqua2_1;
	wire w_dff_B_tozgo1T96_0;
	wire w_dff_B_DgWSqdmm5_1;
	wire w_dff_B_eNbCbCNd4_1;
	wire w_dff_B_pBoU1aAC0_1;
	wire w_dff_B_G73nas932_1;
	wire w_dff_B_oX8bH2f69_1;
	wire w_dff_B_Nhlo4skL5_1;
	wire w_dff_B_LxADl0g43_1;
	wire w_dff_B_0RsxGrIy5_1;
	wire w_dff_B_N69ZWpDm5_1;
	wire w_dff_B_kUjye1l65_1;
	wire w_dff_B_hIuzRHwv3_0;
	wire w_dff_B_2dW9nCZU7_1;
	wire w_dff_B_ylFxSofU1_1;
	wire w_dff_B_Jtue7Ywt4_0;
	wire w_dff_B_rGGKJFCI5_1;
	wire w_dff_B_H3GTqRv49_1;
	wire w_dff_B_8ry3nHbt8_1;
	wire w_dff_B_nAuGj7r26_1;
	wire w_dff_B_ZCt0lbDj7_1;
	wire w_dff_B_qGz8nn0O6_1;
	wire w_dff_B_qCna0wrc1_1;
	wire w_dff_B_1MK5rQm16_1;
	wire w_dff_B_N2gd7BK42_1;
	wire w_dff_B_hk70EXhB4_1;
	wire w_dff_B_fnNiVSQg0_0;
	wire w_dff_B_zn2dswtc8_1;
	wire w_dff_B_J9KIgtCx9_1;
	wire w_dff_B_YlyhWCe47_1;
	wire w_dff_B_pbjsvJRU0_1;
	wire w_dff_B_1NL5v4dj1_1;
	wire w_dff_B_cHVmEYYS1_1;
	wire w_dff_B_tmydoCWx9_1;
	wire w_dff_B_dSDMYpiX8_1;
	wire w_dff_B_yWsrWUVz8_1;
	wire w_dff_B_PJjnjmSe8_1;
	wire w_dff_B_b8CiSugl5_0;
	wire w_dff_B_4u4V4i842_1;
	wire w_dff_B_HatNyVWj5_1;
	wire w_dff_B_EftOFYUE7_1;
	wire w_dff_B_OFdIWwF79_1;
	wire w_dff_B_of9B41I48_1;
	wire w_dff_B_ZQDJ7Ux87_1;
	wire w_dff_B_HdRHntcb1_1;
	wire w_dff_B_LlIFSUYG1_1;
	wire w_dff_B_ga74nord4_1;
	wire w_dff_B_vg76XKpv7_1;
	wire w_dff_B_rECqHm9H4_0;
	wire w_dff_B_EdOZ8SLX0_1;
	wire w_dff_B_qelqFzvL8_1;
	wire w_dff_B_Y1FGDnUK0_1;
	wire w_dff_B_OXno1hik8_1;
	wire w_dff_B_r7LsM7Df4_1;
	wire w_dff_B_e7wXA7DB3_1;
	wire w_dff_B_psoYtpqQ6_1;
	wire w_dff_B_hHESg9fo8_1;
	wire w_dff_B_sukwBUro7_1;
	wire w_dff_B_qIVWh7nJ2_1;
	wire w_dff_B_b2g877Zq9_0;
	wire w_dff_B_nVt1r1Pg4_1;
	wire w_dff_B_3n3bcFZF0_1;
	wire w_dff_B_yFXClqjf2_0;
	wire w_dff_B_lGKQzauE6_1;
	wire w_dff_A_4pYXSgZQ4_0;
	wire w_dff_A_eOY9af3E1_1;
	wire w_dff_B_b1xub7d40_1;
	wire w_dff_A_jsqcgtqV5_0;
	wire w_dff_A_Tf7v1fro5_1;
	wire w_dff_B_qUAu1S6Q0_1;
	wire w_dff_A_I7gyfdFq9_0;
	wire w_dff_A_NA9ziZSD5_1;
	wire w_dff_B_BcmFF8576_1;
	wire w_dff_A_3gOkgdes3_0;
	wire w_dff_A_tD9nMY0t2_1;
	wire w_dff_B_Q6hzBaEe4_1;
	wire w_dff_A_bhAqClr40_0;
	wire w_dff_A_qYdmnUej7_1;
	wire w_dff_B_ZwKVErzE1_1;
	wire w_dff_A_SwhSpGG03_0;
	wire w_dff_A_yYiuMmAx6_1;
	wire w_dff_B_i0X0OPVY5_1;
	wire w_dff_A_aYzwVtdH1_0;
	wire w_dff_A_9PjzwdE12_1;
	wire w_dff_B_sqLFKCT85_1;
	wire w_dff_A_ipr72ra02_0;
	wire w_dff_A_APWgC3dM4_1;
	wire w_dff_B_f7q9HcgA4_1;
	wire w_dff_B_rUo3KNte8_1;
	wire w_dff_B_QlNfdnSh4_0;
	wire w_dff_B_WSLDAw9h6_1;
	wire w_dff_A_Xt1EtlJu1_0;
	wire w_dff_A_Pe361rYG6_1;
	wire w_dff_B_yG764QYf5_1;
	wire w_dff_A_8B97r3VV0_0;
	wire w_dff_A_RTG96NZT0_1;
	wire w_dff_B_42tADvHd7_1;
	wire w_dff_A_wSYwKQKp9_0;
	wire w_dff_A_OiMf06K86_1;
	wire w_dff_B_KImY48fm3_1;
	wire w_dff_A_FxenSOIp9_0;
	wire w_dff_A_X1Lfnzwj8_1;
	wire w_dff_B_XT5fswlN8_1;
	wire w_dff_A_5fD5AaYw7_0;
	wire w_dff_A_TrlnadzK5_1;
	wire w_dff_B_uvuIOWOm0_1;
	wire w_dff_A_i8HqUX7H4_0;
	wire w_dff_A_OcSdyoQr6_1;
	wire w_dff_B_8NBshqAL6_1;
	wire w_dff_A_p4g9Yx0Z8_0;
	wire w_dff_A_OxxYjRfR3_1;
	wire w_dff_B_NrGt6CJe2_1;
	wire w_dff_A_nt5Btme91_0;
	wire w_dff_A_uSzz6U2s7_1;
	wire w_dff_B_xgjTbxSc2_1;
	wire w_dff_B_zacrjjWS4_1;
	wire w_dff_B_5qLGuZg58_0;
	wire w_dff_B_py7Eagjp9_1;
	wire w_dff_A_4h0NH7LH3_0;
	wire w_dff_A_amGWYNxX5_1;
	wire w_dff_B_8EZYNZap4_1;
	wire w_dff_A_HbBmurSs9_0;
	wire w_dff_A_3E0UAqQJ7_1;
	wire w_dff_B_1lzHYFyY3_1;
	wire w_dff_A_BB5cJRhF0_0;
	wire w_dff_A_x0WLNzz69_1;
	wire w_dff_B_iPHr0LC45_1;
	wire w_dff_A_KWIu5I4M0_0;
	wire w_dff_A_NhWoqlJE7_1;
	wire w_dff_B_LzHuIvWe7_1;
	wire w_dff_A_x1m5wCkQ3_0;
	wire w_dff_A_fFCBlUt64_1;
	wire w_dff_B_mXMNmnXD2_1;
	wire w_dff_A_tioEWBSH6_0;
	wire w_dff_A_iMM7uM3x0_1;
	wire w_dff_B_Qru46Pym3_1;
	wire w_dff_A_a4SNezFT6_0;
	wire w_dff_A_bbcJxZ647_1;
	wire w_dff_B_LyBW2d6f4_1;
	wire w_dff_A_3R8e6hTN0_0;
	wire w_dff_A_nyGrOAiO3_1;
	wire w_dff_B_vJXNk5uA4_1;
	wire w_dff_B_DlowA4MC0_1;
	wire w_dff_B_bqhhQYEO8_0;
	wire w_dff_B_FIhTqrhf7_1;
	wire w_dff_A_RGJo87rH1_0;
	wire w_dff_A_4GIKWQI35_1;
	wire w_dff_B_745QdKaB0_1;
	wire w_dff_A_aqMYVpgr1_0;
	wire w_dff_A_bKqOvwAI6_1;
	wire w_dff_B_g2UrCknn7_1;
	wire w_dff_A_SKaaili94_0;
	wire w_dff_A_nSHI3wrB2_1;
	wire w_dff_B_K0Y4km6g5_1;
	wire w_dff_A_kGWQUzm74_0;
	wire w_dff_A_q0xtfwdX5_1;
	wire w_dff_B_dyfUBpGV8_1;
	wire w_dff_A_lRhC755p2_0;
	wire w_dff_A_ECSpmsBT6_1;
	wire w_dff_B_sskXJKkD8_1;
	wire w_dff_A_aEQEN3Xf2_0;
	wire w_dff_A_vTXKnj262_1;
	wire w_dff_B_43V9h6ET3_1;
	wire w_dff_A_2Aq7vbmA8_0;
	wire w_dff_A_OqgJmqtR1_1;
	wire w_dff_B_rF98fik62_1;
	wire w_dff_A_qYADieKW4_0;
	wire w_dff_A_p4ahpbAJ4_1;
	wire w_dff_B_spBzN65s6_1;
	wire w_dff_B_o6DVcVCt5_1;
	wire w_dff_B_ClAbqRb96_0;
	wire w_dff_B_aUU9y1mb9_1;
	wire w_dff_B_uSl1DoMb4_1;
	wire w_dff_B_TnrR4rFy8_0;
	wire w_dff_B_Np9QaPFa9_1;
	wire w_dff_A_hUN70b8y2_0;
	wire w_dff_A_dUrA3tEd2_1;
	wire w_dff_B_PH0lI8405_1;
	wire w_dff_A_XF2Yyt4V5_0;
	wire w_dff_A_bTr2Cfs06_1;
	wire w_dff_B_JkVSSvVk5_1;
	wire w_dff_A_4hVRVXx43_0;
	wire w_dff_A_IeX7m3QI0_1;
	wire w_dff_B_tarZfy621_1;
	wire w_dff_A_wkaxuBD72_0;
	wire w_dff_A_7OB6oRqA1_1;
	wire w_dff_B_mYmJWWo27_1;
	wire w_dff_A_we9q0Jad5_0;
	wire w_dff_A_VjN2Qliq0_1;
	wire w_dff_B_sBdhvQYX3_1;
	wire w_dff_A_O8Ze6Upb1_0;
	wire w_dff_A_Z0uMSCcz9_1;
	wire w_dff_B_upysfaBQ0_1;
	wire w_dff_A_VKlsC5cZ2_0;
	wire w_dff_A_Wwy7IlhU6_1;
	wire w_dff_B_1VoqRzDF0_1;
	wire w_dff_A_Dkax2EMe2_0;
	wire w_dff_A_qtRk7Icw0_1;
	wire w_dff_B_DMqPlBFe5_3;
	wire w_dff_B_jUEppjKS7_3;
	wire w_dff_B_NzBHWWlV2_3;
	wire w_dff_B_WUQO6yvK5_3;
	wire w_dff_B_inBTF3Cj2_3;
	wire w_dff_B_1nYZ6e8Z1_3;
	wire w_dff_B_ypPvMaYr6_3;
	wire w_dff_B_rk8XASRI6_1;
	wire w_dff_B_871fhSZh8_1;
	wire w_dff_B_Ewoal9ki5_0;
	wire w_dff_B_DGgUZnJK3_1;
	wire w_dff_A_rcrknBQy7_0;
	wire w_dff_A_PUmUpuIX0_1;
	wire w_dff_B_uICq5SCD7_1;
	wire w_dff_A_JPoE7RgR9_0;
	wire w_dff_A_KS7aaRbG4_1;
	wire w_dff_B_fsEUZG1w2_1;
	wire w_dff_A_JozpVLIs7_0;
	wire w_dff_A_P7ahRfJd1_1;
	wire w_dff_B_Wz80cizW6_1;
	wire w_dff_A_g47baKUj6_0;
	wire w_dff_A_2LdNMFjs0_1;
	wire w_dff_B_6YxyaqYr2_1;
	wire w_dff_A_5wvWWH0g3_0;
	wire w_dff_A_2ewe9RPU2_1;
	wire w_dff_B_aBi3tGKD9_1;
	wire w_dff_A_V7FH9gfr3_0;
	wire w_dff_A_IhAADU2o4_1;
	wire w_dff_B_oi8DblKT5_1;
	wire w_dff_A_aZ8WAfFs3_0;
	wire w_dff_A_jaLZbcNB9_1;
	wire w_dff_B_h6051X5M0_1;
	wire w_dff_A_vcWxBCo84_0;
	wire w_dff_A_n7nis0rM6_1;
	wire w_dff_B_9BosVVVW8_3;
	wire w_dff_B_y1OvB6m63_3;
	wire w_dff_B_pGhbj1re6_3;
	wire w_dff_B_e40Q35VS4_3;
	wire w_dff_B_qGUjWA5Y0_3;
	wire w_dff_B_NOMuLjAk2_3;
	wire w_dff_B_EZWknVjS0_3;
	wire w_dff_B_F1l9p9yf4_3;
	wire w_dff_B_jTlFOYMo5_1;
	wire w_dff_B_5fVocIcW4_1;
	wire w_dff_B_sdDWXqfe3_0;
	wire w_dff_B_Pj71flbm8_1;
	wire w_dff_A_FL8rfjir2_0;
	wire w_dff_A_7GZZbsWq5_1;
	wire w_dff_B_xpd5mGRp3_1;
	wire w_dff_A_JsBVmPGJ3_0;
	wire w_dff_A_LpS4cIVI1_1;
	wire w_dff_B_MFGGkqzk7_1;
	wire w_dff_A_HqaVWGpG4_0;
	wire w_dff_A_EfquT9R57_1;
	wire w_dff_B_gXNcxvia2_1;
	wire w_dff_A_6rr88UQ06_0;
	wire w_dff_A_IjOIf2Vv3_1;
	wire w_dff_B_o7JVhuzP9_1;
	wire w_dff_A_ypOJA4Mn4_0;
	wire w_dff_A_ECU7ndwr9_1;
	wire w_dff_B_a5mabnqU6_1;
	wire w_dff_A_z9RlMpd06_0;
	wire w_dff_A_OrPlTNw66_1;
	wire w_dff_B_DVmtjqsy4_1;
	wire w_dff_A_yNeInT2q0_0;
	wire w_dff_A_yjHZSHH70_1;
	wire w_dff_B_TF8VuoJz5_1;
	wire w_dff_A_ixqoCv1I6_0;
	wire w_dff_A_AvFtfhSE5_1;
	wire w_dff_B_CxYsv1cW2_3;
	wire w_dff_B_qeWyi0A84_3;
	wire w_dff_B_81YZhcyd8_3;
	wire w_dff_B_KLxrtH251_3;
	wire w_dff_B_1oN0NPYh2_3;
	wire w_dff_B_FM0LHf2p9_3;
	wire w_dff_B_eLdE6Tba8_3;
	wire w_dff_B_2BfiXtTV3_1;
	wire w_dff_B_wKhuxg1O7_1;
	wire w_dff_B_sFr9dA5r6_0;
	wire w_dff_B_v2guYC8y6_1;
	wire w_dff_A_HmdqNm8g4_0;
	wire w_dff_A_8mgBZIQg7_1;
	wire w_dff_B_0oLZnUPh4_1;
	wire w_dff_A_ruJEv85L7_0;
	wire w_dff_A_zbNXoOqW6_1;
	wire w_dff_B_T6FhMLOl0_3;
	wire w_dff_B_2lyKqjFZ9_3;
	wire w_dff_B_L3XqwQjn4_3;
	wire w_dff_B_PK6M6bQk2_1;
	wire w_dff_A_qerx9cuT9_0;
	wire w_dff_A_MCBIUaBq2_1;
	wire w_dff_B_YqCEMGkj8_1;
	wire w_dff_A_x9iScKCA1_0;
	wire w_dff_A_mAgVgHU16_1;
	wire w_dff_B_3n7FITo24_3;
	wire w_dff_B_2lzJbilg4_3;
	wire w_dff_B_bi8l2YH76_3;
	wire w_dff_B_H2R9KPX95_3;
	wire w_dff_B_tfJFhTxG8_1;
	wire w_dff_A_xNYvrMCm0_0;
	wire w_dff_A_0nnYYHF55_1;
	wire w_dff_B_SLXi6sqx0_1;
	wire w_dff_A_TEmwG3XJ6_0;
	wire w_dff_A_r5bZU0Yn6_1;
	wire w_dff_B_x2mt324E2_3;
	wire w_dff_B_rnaB24hv3_3;
	wire w_dff_B_FULzpxU81_3;
	wire w_dff_B_HKuzR6c52_1;
	wire w_dff_A_AY4LJMyP2_0;
	wire w_dff_A_td3IjRBo8_1;
	wire w_dff_B_5jw3Llau0_3;
	wire w_dff_B_AMEaIxgs6_3;
	wire w_dff_A_e2KaJXa04_0;
	wire w_dff_A_vpG9IxaZ1_0;
	wire w_dff_A_hDIMdffy1_0;
	wire w_dff_A_1Z7k3zc65_2;
	wire w_dff_A_OmMWeXIQ2_2;
	wire w_dff_A_bMqTrhbp3_2;
	wire w_dff_A_RC8wWg7O0_0;
	wire w_dff_A_hcEVGi5I5_0;
	wire w_dff_A_9kI7kVaC9_0;
	wire w_dff_A_ATtTd43D2_1;
	wire w_dff_A_VgBYN22x4_1;
	wire w_dff_A_rtDyqCOd8_1;
	wire w_dff_A_aJMy0lZt4_0;
	wire w_dff_A_1KxTcwcD2_0;
	wire w_dff_A_imsCNVkT2_0;
	wire w_dff_A_MyYUwFlP4_2;
	wire w_dff_A_dyImM1rh4_2;
	wire w_dff_A_mDIUIck97_2;
	wire w_dff_A_88LexBq42_0;
	wire w_dff_A_NqFXEflt2_0;
	wire w_dff_A_VLfOiBZL1_0;
	wire w_dff_A_zcodIgwo3_1;
	wire w_dff_A_anpED3qE4_1;
	wire w_dff_A_LfupF43K8_1;
	wire w_dff_B_innup2oD0_1;
	wire w_dff_A_Nsc29slm7_0;
	wire w_dff_A_S63Jgp8X2_1;
	wire w_dff_A_FxTfk7bY2_1;
	wire w_dff_A_MOLsVTew2_1;
	wire w_dff_A_2auC8Ory6_1;
	wire w_dff_A_4rP6ARZQ0_2;
	wire w_dff_A_Mwoc0Tgp8_2;
	wire w_dff_A_ewMNBLer3_2;
	wire w_dff_B_3XLTqWEN0_3;
	wire w_dff_B_mkxpvy5v7_3;
	wire w_dff_B_BzJqvu7e0_3;
	wire w_dff_A_6q7NhxpC3_1;
	wire w_dff_A_iZkaQ2vc3_2;
	wire w_dff_B_cWtJz30h3_3;
	wire w_dff_B_JG7qnRyB1_3;
	wire w_dff_B_odhJBSIE1_3;
	wire w_dff_B_7rQcpyIn7_3;
	wire w_dff_B_TNFpLTFg8_3;
	wire w_dff_B_zRdqDAAF6_3;
	wire w_dff_B_cE1lYXHF5_3;
	wire w_dff_A_6JmKMWA78_2;
	wire w_dff_A_kHgVQNIK1_1;
	wire w_dff_B_D1MyPfrQ5_3;
	wire w_dff_B_TlEknDsx1_3;
	wire w_dff_B_7lDjzph70_3;
	wire w_dff_B_rFdjlMZD1_3;
	wire w_dff_B_cpeRMzaJ8_3;
	wire w_dff_B_ZPRNw5ou6_3;
	wire w_dff_B_LUTSYlbD1_3;
	wire w_dff_B_SchMfHZx3_3;
	wire w_dff_B_lPjXFL1b0_3;
	wire w_dff_B_rFFecGf23_3;
	wire w_dff_B_wnnGE9y38_3;
	wire w_dff_B_auwam0s87_3;
	wire w_dff_A_yAJH0Bn31_0;
	wire w_dff_A_UgEDVB5a1_0;
	wire w_dff_A_cXfHOD8n6_0;
	wire w_dff_A_BJ1qMqCb1_0;
	wire w_dff_A_KvzloDZH6_0;
	wire w_dff_A_DlfBdeCe3_0;
	wire w_dff_A_Mw1W6pyL3_0;
	wire w_dff_A_7I6ciW9d6_0;
	wire w_dff_A_k0l05ikN7_0;
	wire w_dff_A_8CG9Zvle8_0;
	wire w_dff_A_O19qIvxa8_0;
	wire w_dff_A_1lSULzdc6_0;
	wire w_dff_A_bqhDMCvs6_0;
	wire w_dff_A_asXnvvCp1_1;
	wire w_dff_A_7MV0wofZ2_1;
	wire w_dff_A_YYodgnKE3_1;
	wire w_dff_A_OAQAKcMT7_1;
	wire w_dff_A_a6OmcwGy4_1;
	wire w_dff_A_7awDuIx24_1;
	wire w_dff_A_zHovBbBN9_1;
	wire w_dff_A_GEHCN80u4_1;
	wire w_dff_A_5v7paUrI6_1;
	wire w_dff_A_gm71wfmI4_1;
	wire w_dff_A_rlnw4zxw4_1;
	wire w_dff_A_ntqqrbQY5_1;
	wire w_dff_A_QEbkLJAp3_1;
	wire w_dff_A_yTLlrHtH8_0;
	wire w_dff_A_6WbT2UZz4_0;
	wire w_dff_A_s0Zks23c4_0;
	wire w_dff_A_KVbybT3z0_0;
	wire w_dff_A_sUerBJWF3_0;
	wire w_dff_A_KwRqLfUv4_0;
	wire w_dff_A_MPQc3Pdx9_0;
	wire w_dff_A_kc3JFFaF5_0;
	wire w_dff_A_kDlzFewf6_0;
	wire w_dff_A_RtiDpvgr1_0;
	wire w_dff_A_Fex9r6ri9_0;
	wire w_dff_A_wIe7t5VD4_0;
	wire w_dff_A_SkPkN92h4_0;
	wire w_dff_A_VI5eUidT5_1;
	wire w_dff_A_NWadLbxG1_1;
	wire w_dff_A_zqTuj6v83_1;
	wire w_dff_A_peXhlYT34_1;
	wire w_dff_A_7giuYgW11_1;
	wire w_dff_A_Sg3rSI1a8_1;
	wire w_dff_A_FWlwrulx5_1;
	wire w_dff_A_kFQVZGOf6_1;
	wire w_dff_A_gMPxVi5q6_1;
	wire w_dff_A_aWYGTbjE2_1;
	wire w_dff_A_xz481dg06_1;
	wire w_dff_A_9TqyH9XI9_1;
	wire w_dff_A_GnocIZ4d7_1;
	wire w_dff_A_CxgjtJf25_0;
	wire w_dff_A_aqwxP7733_0;
	wire w_dff_A_QaxrS6Bk7_0;
	wire w_dff_A_QR95RoFe4_0;
	wire w_dff_A_zc0yCe6x6_0;
	wire w_dff_A_ds5wZAaK9_0;
	wire w_dff_A_JHwHU07f3_0;
	wire w_dff_A_tQvjFbhx2_0;
	wire w_dff_A_7l4ZZ3Oy4_0;
	wire w_dff_A_JJ01ICRq4_0;
	wire w_dff_A_eYY6o3js5_0;
	wire w_dff_A_QMLCc8ja8_0;
	wire w_dff_A_ilrk8ITG9_0;
	wire w_dff_A_9KEoRETL5_2;
	wire w_dff_A_xQz8WY0T2_2;
	wire w_dff_A_VqmGKOO02_2;
	wire w_dff_A_Hgg1ozR90_2;
	wire w_dff_A_wQQikEXv7_2;
	wire w_dff_A_mf1pd0do8_2;
	wire w_dff_A_B4U2IVCW5_2;
	wire w_dff_A_WzNzoCIq5_2;
	wire w_dff_A_50ekwJrz5_2;
	wire w_dff_A_YxGiN22x4_2;
	wire w_dff_A_Ly6xRXqK6_2;
	wire w_dff_A_uudtF6AE7_2;
	wire w_dff_A_NGTUJztT7_2;
	wire w_dff_A_OEfCsjIo7_0;
	wire w_dff_A_moDPj9Iq5_0;
	wire w_dff_A_ltgJltH36_0;
	wire w_dff_A_sb6j7kem3_0;
	wire w_dff_A_iQ2BsceM8_0;
	wire w_dff_A_5sYHyqNT2_0;
	wire w_dff_A_KFLXylHK7_0;
	wire w_dff_A_bLaMM5ge3_0;
	wire w_dff_A_tFBeomrf2_0;
	wire w_dff_A_RfTcGk5e1_0;
	wire w_dff_A_SG4k4aTM0_0;
	wire w_dff_A_7akYvcM92_0;
	wire w_dff_A_LF7uoH3p0_0;
	wire w_dff_A_OYJcZjJL1_1;
	wire w_dff_A_wsTqhXUy8_1;
	wire w_dff_A_OsgiMFyk8_1;
	wire w_dff_A_3UlkHgJ53_1;
	wire w_dff_A_qpXxM72y4_1;
	wire w_dff_A_INOTK3000_1;
	wire w_dff_A_c48fOM751_1;
	wire w_dff_A_yIPwSEAS6_1;
	wire w_dff_A_uZDh0bOA9_1;
	wire w_dff_A_s2JklApE7_1;
	wire w_dff_A_Vg7e5cJ63_1;
	wire w_dff_A_mn4QwLaf2_1;
	wire w_dff_A_yhw6Bu9C1_1;
	wire w_dff_A_d0HlFfEt8_1;
	wire w_dff_A_0KHUZMz38_1;
	wire w_dff_A_WOA0ZQHw3_1;
	wire w_dff_A_nn1kfmOP4_1;
	wire w_dff_A_wlxdjjOG7_1;
	wire w_dff_A_hx4tVmIK8_1;
	wire w_dff_A_UyHOTMnZ3_1;
	wire w_dff_A_ITcnN2XY5_1;
	wire w_dff_A_VbtfVEBv5_1;
	wire w_dff_A_dr5pNRNJ3_1;
	wire w_dff_A_SBbXK7hb5_1;
	wire w_dff_A_GQoVLGyR6_1;
	wire w_dff_A_khYPEM4x6_1;
	wire w_dff_A_2TQqs4AQ5_2;
	wire w_dff_A_6LJGIMCL8_2;
	wire w_dff_A_bI9SQkqI0_2;
	wire w_dff_A_XbM50qoe5_2;
	wire w_dff_A_OlXmRDr23_2;
	wire w_dff_A_tYxLAhIr1_2;
	wire w_dff_A_MxFCGgOe5_2;
	wire w_dff_A_ujp1IjfH8_2;
	wire w_dff_A_chwKj2SQ7_2;
	wire w_dff_A_4gtYzkjf5_2;
	wire w_dff_A_8Of7GbxQ4_2;
	wire w_dff_A_s1NI9TQu9_2;
	wire w_dff_A_eLfj31eX1_2;
	jnot g0000(.din(w_shift6_63[2]),.dout(n263),.clk(gclk));
	jnot g0001(.din(w_shift4_0[2]),.dout(n264),.clk(gclk));
	jand g0002(.dina(w_shift5_0[2]),.dinb(w_n264_0[1]),.dout(n265),.clk(gclk));
	jnot g0003(.din(w_shift3_0[2]),.dout(n266),.clk(gclk));
	jand g0004(.dina(w_n266_0[1]),.dinb(w_shift2_0[2]),.dout(n267),.clk(gclk));
	jor g0005(.dina(w_shift0_63[2]),.dinb(w_a28_0[1]),.dout(n268),.clk(gclk));
	jnot g0006(.din(w_shift0_63[1]),.dout(n269),.clk(gclk));
	jor g0007(.dina(w_n269_63[1]),.dinb(w_a27_0[1]),.dout(n270),.clk(gclk));
	jand g0008(.dina(n270),.dinb(w_dff_B_HatNyVWj5_1),.dout(n271),.clk(gclk));
	jor g0009(.dina(w_n271_0[1]),.dinb(w_shift1_63[2]),.dout(n272),.clk(gclk));
	jnot g0010(.din(w_shift1_63[1]),.dout(n273),.clk(gclk));
	jor g0011(.dina(w_shift0_63[0]),.dinb(w_a26_0[1]),.dout(n274),.clk(gclk));
	jor g0012(.dina(w_n269_63[0]),.dinb(w_a25_0[1]),.dout(n275),.clk(gclk));
	jand g0013(.dina(n275),.dinb(w_dff_B_EftOFYUE7_1),.dout(n276),.clk(gclk));
	jor g0014(.dina(w_n276_0[1]),.dinb(w_n273_63[1]),.dout(n277),.clk(gclk));
	jand g0015(.dina(n277),.dinb(n272),.dout(n278),.clk(gclk));
	jand g0016(.dina(w_n278_1[1]),.dinb(w_n267_63[1]),.dout(n279),.clk(gclk));
	jnot g0017(.din(w_shift2_0[1]),.dout(n280),.clk(gclk));
	jand g0018(.dina(w_shift3_0[1]),.dinb(w_n280_0[1]),.dout(n281),.clk(gclk));
	jor g0019(.dina(w_shift0_62[2]),.dinb(w_a24_0[1]),.dout(n282),.clk(gclk));
	jor g0020(.dina(w_n269_62[2]),.dinb(w_a23_0[1]),.dout(n283),.clk(gclk));
	jand g0021(.dina(n283),.dinb(w_dff_B_OFdIWwF79_1),.dout(n284),.clk(gclk));
	jor g0022(.dina(w_n284_0[1]),.dinb(w_shift1_63[0]),.dout(n285),.clk(gclk));
	jor g0023(.dina(w_shift0_62[1]),.dinb(w_a22_0[1]),.dout(n286),.clk(gclk));
	jor g0024(.dina(w_n269_62[1]),.dinb(w_a21_0[1]),.dout(n287),.clk(gclk));
	jand g0025(.dina(n287),.dinb(w_dff_B_of9B41I48_1),.dout(n288),.clk(gclk));
	jor g0026(.dina(w_n288_0[1]),.dinb(w_n273_63[0]),.dout(n289),.clk(gclk));
	jand g0027(.dina(n289),.dinb(n285),.dout(n290),.clk(gclk));
	jand g0028(.dina(w_n290_1[1]),.dinb(w_n281_63[1]),.dout(n291),.clk(gclk));
	jand g0029(.dina(w_shift3_0[0]),.dinb(w_shift2_0[0]),.dout(n292),.clk(gclk));
	jor g0030(.dina(w_shift0_62[0]),.dinb(w_a20_0[1]),.dout(n293),.clk(gclk));
	jor g0031(.dina(w_n269_62[0]),.dinb(w_a19_0[1]),.dout(n294),.clk(gclk));
	jand g0032(.dina(n294),.dinb(w_dff_B_ZQDJ7Ux87_1),.dout(n295),.clk(gclk));
	jor g0033(.dina(w_n295_0[1]),.dinb(w_shift1_62[2]),.dout(n296),.clk(gclk));
	jor g0034(.dina(w_shift0_61[2]),.dinb(w_a18_0[1]),.dout(n297),.clk(gclk));
	jor g0035(.dina(w_n269_61[2]),.dinb(w_a17_0[1]),.dout(n298),.clk(gclk));
	jand g0036(.dina(n298),.dinb(w_dff_B_HdRHntcb1_1),.dout(n299),.clk(gclk));
	jor g0037(.dina(w_n299_0[1]),.dinb(w_n273_62[2]),.dout(n300),.clk(gclk));
	jand g0038(.dina(n300),.dinb(n296),.dout(n301),.clk(gclk));
	jand g0039(.dina(w_n301_1[1]),.dinb(w_n292_63[1]),.dout(n302),.clk(gclk));
	jor g0040(.dina(n302),.dinb(n291),.dout(n303),.clk(gclk));
	jand g0041(.dina(w_n266_0[0]),.dinb(w_n280_0[0]),.dout(n304),.clk(gclk));
	jor g0042(.dina(w_shift0_61[1]),.dinb(w_a32_0[1]),.dout(n305),.clk(gclk));
	jor g0043(.dina(w_n269_61[1]),.dinb(w_a31_0[1]),.dout(n306),.clk(gclk));
	jand g0044(.dina(n306),.dinb(w_dff_B_pbjsvJRU0_1),.dout(n307),.clk(gclk));
	jor g0045(.dina(w_n307_0[1]),.dinb(w_shift1_62[1]),.dout(n308),.clk(gclk));
	jor g0046(.dina(w_shift0_61[0]),.dinb(w_a30_0[1]),.dout(n309),.clk(gclk));
	jor g0047(.dina(w_n269_61[0]),.dinb(w_a29_0[1]),.dout(n310),.clk(gclk));
	jand g0048(.dina(n310),.dinb(w_dff_B_4u4V4i842_1),.dout(n311),.clk(gclk));
	jor g0049(.dina(w_n311_0[1]),.dinb(w_n273_62[1]),.dout(n312),.clk(gclk));
	jand g0050(.dina(n312),.dinb(n308),.dout(n313),.clk(gclk));
	jand g0051(.dina(w_n313_1[1]),.dinb(w_n304_63[1]),.dout(n314),.clk(gclk));
	jor g0052(.dina(w_dff_B_GF88rIeY2_0),.dinb(n303),.dout(n315),.clk(gclk));
	jor g0053(.dina(n315),.dinb(w_dff_B_ENIICq2y3_1),.dout(n316),.clk(gclk));
	jand g0054(.dina(w_n316_1[1]),.dinb(w_n265_63[1]),.dout(n317),.clk(gclk));
	jnot g0055(.din(w_shift5_0[1]),.dout(n318),.clk(gclk));
	jand g0056(.dina(w_n318_0[1]),.dinb(w_shift4_0[1]),.dout(n319),.clk(gclk));
	jor g0057(.dina(w_shift0_60[2]),.dinb(w_a36_0[1]),.dout(n320),.clk(gclk));
	jor g0058(.dina(w_n269_60[2]),.dinb(w_a35_0[1]),.dout(n321),.clk(gclk));
	jand g0059(.dina(n321),.dinb(w_dff_B_cHVmEYYS1_1),.dout(n322),.clk(gclk));
	jor g0060(.dina(w_n322_0[1]),.dinb(w_shift1_62[0]),.dout(n323),.clk(gclk));
	jor g0061(.dina(w_shift0_60[1]),.dinb(w_a34_0[1]),.dout(n324),.clk(gclk));
	jor g0062(.dina(w_n269_60[1]),.dinb(w_a33_0[1]),.dout(n325),.clk(gclk));
	jand g0063(.dina(n325),.dinb(w_dff_B_YlyhWCe47_1),.dout(n326),.clk(gclk));
	jor g0064(.dina(w_n326_0[1]),.dinb(w_n273_62[0]),.dout(n327),.clk(gclk));
	jand g0065(.dina(n327),.dinb(n323),.dout(n328),.clk(gclk));
	jand g0066(.dina(w_n328_1[1]),.dinb(w_n292_63[0]),.dout(n329),.clk(gclk));
	jor g0067(.dina(w_shift0_60[0]),.dinb(w_a40_0[1]),.dout(n330),.clk(gclk));
	jor g0068(.dina(w_n269_60[0]),.dinb(w_a39_0[1]),.dout(n331),.clk(gclk));
	jand g0069(.dina(n331),.dinb(w_dff_B_dSDMYpiX8_1),.dout(n332),.clk(gclk));
	jand g0070(.dina(w_n332_0[1]),.dinb(w_n273_61[2]),.dout(n333),.clk(gclk));
	jor g0071(.dina(w_shift0_59[2]),.dinb(w_a38_0[1]),.dout(n334),.clk(gclk));
	jor g0072(.dina(w_n269_59[2]),.dinb(w_a37_0[1]),.dout(n335),.clk(gclk));
	jand g0073(.dina(n335),.dinb(w_dff_B_1NL5v4dj1_1),.dout(n336),.clk(gclk));
	jand g0074(.dina(w_n336_0[1]),.dinb(w_shift1_61[2]),.dout(n337),.clk(gclk));
	jor g0075(.dina(n337),.dinb(n333),.dout(n338),.clk(gclk));
	jand g0076(.dina(w_n338_1[1]),.dinb(w_n281_63[0]),.dout(n339),.clk(gclk));
	jor g0077(.dina(w_shift0_59[1]),.dinb(w_a44_0[1]),.dout(n340),.clk(gclk));
	jor g0078(.dina(w_n269_59[1]),.dinb(w_a43_0[1]),.dout(n341),.clk(gclk));
	jand g0079(.dina(n341),.dinb(w_dff_B_zn2dswtc8_1),.dout(n342),.clk(gclk));
	jor g0080(.dina(w_n342_0[1]),.dinb(w_shift1_61[1]),.dout(n343),.clk(gclk));
	jor g0081(.dina(w_shift0_59[0]),.dinb(w_a42_0[1]),.dout(n344),.clk(gclk));
	jor g0082(.dina(w_n269_59[0]),.dinb(w_a41_0[1]),.dout(n345),.clk(gclk));
	jand g0083(.dina(n345),.dinb(w_dff_B_tmydoCWx9_1),.dout(n346),.clk(gclk));
	jor g0084(.dina(w_n346_0[1]),.dinb(w_n273_61[1]),.dout(n347),.clk(gclk));
	jand g0085(.dina(n347),.dinb(n343),.dout(n348),.clk(gclk));
	jand g0086(.dina(w_n348_1[1]),.dinb(w_n267_63[0]),.dout(n349),.clk(gclk));
	jor g0087(.dina(n349),.dinb(n339),.dout(n350),.clk(gclk));
	jor g0088(.dina(w_shift0_58[2]),.dinb(w_a48_0[1]),.dout(n351),.clk(gclk));
	jor g0089(.dina(w_n269_58[2]),.dinb(w_a47_0[1]),.dout(n352),.clk(gclk));
	jand g0090(.dina(n352),.dinb(w_dff_B_H3GTqRv49_1),.dout(n353),.clk(gclk));
	jor g0091(.dina(w_n353_0[1]),.dinb(w_shift1_61[0]),.dout(n354),.clk(gclk));
	jor g0092(.dina(w_shift0_58[1]),.dinb(w_a46_0[1]),.dout(n355),.clk(gclk));
	jor g0093(.dina(w_n269_58[1]),.dinb(w_a45_0[1]),.dout(n356),.clk(gclk));
	jand g0094(.dina(n356),.dinb(w_dff_B_J9KIgtCx9_1),.dout(n357),.clk(gclk));
	jor g0095(.dina(w_n357_0[1]),.dinb(w_n273_61[0]),.dout(n358),.clk(gclk));
	jand g0096(.dina(n358),.dinb(n354),.dout(n359),.clk(gclk));
	jand g0097(.dina(w_n359_1[1]),.dinb(w_n304_63[0]),.dout(n360),.clk(gclk));
	jor g0098(.dina(w_dff_B_TkhLCRu23_0),.dinb(n350),.dout(n361),.clk(gclk));
	jor g0099(.dina(n361),.dinb(w_dff_B_faRWqwxy6_1),.dout(n362),.clk(gclk));
	jand g0100(.dina(w_n362_1[1]),.dinb(w_n319_63[1]),.dout(n363),.clk(gclk));
	jand g0101(.dina(w_n318_0[0]),.dinb(w_n264_0[0]),.dout(n364),.clk(gclk));
	jor g0102(.dina(w_shift0_58[0]),.dinb(w_a64_0[1]),.dout(n365),.clk(gclk));
	jor g0103(.dina(w_n269_58[0]),.dinb(w_a63_0[1]),.dout(n366),.clk(gclk));
	jand g0104(.dina(n366),.dinb(w_dff_B_jlhhO1862_1),.dout(n367),.clk(gclk));
	jor g0105(.dina(w_n367_0[1]),.dinb(w_shift1_60[2]),.dout(n368),.clk(gclk));
	jor g0106(.dina(w_shift0_57[2]),.dinb(w_a62_0[1]),.dout(n369),.clk(gclk));
	jor g0107(.dina(w_n269_57[2]),.dinb(w_a61_0[1]),.dout(n370),.clk(gclk));
	jand g0108(.dina(n370),.dinb(w_dff_B_qCna0wrc1_1),.dout(n371),.clk(gclk));
	jor g0109(.dina(w_n371_0[1]),.dinb(w_n273_60[2]),.dout(n372),.clk(gclk));
	jand g0110(.dina(n372),.dinb(n368),.dout(n373),.clk(gclk));
	jand g0111(.dina(w_n373_1[1]),.dinb(w_n304_62[2]),.dout(n374),.clk(gclk));
	jor g0112(.dina(w_shift0_57[1]),.dinb(w_a56_0[1]),.dout(n375),.clk(gclk));
	jor g0113(.dina(w_n269_57[1]),.dinb(w_a55_0[1]),.dout(n376),.clk(gclk));
	jand g0114(.dina(n376),.dinb(w_dff_B_nAuGj7r26_1),.dout(n377),.clk(gclk));
	jor g0115(.dina(w_n377_0[1]),.dinb(w_shift1_60[1]),.dout(n378),.clk(gclk));
	jor g0116(.dina(w_shift0_57[0]),.dinb(w_a54_0[1]),.dout(n379),.clk(gclk));
	jor g0117(.dina(w_n269_57[0]),.dinb(w_a53_0[1]),.dout(n380),.clk(gclk));
	jand g0118(.dina(n380),.dinb(w_dff_B_ZCt0lbDj7_1),.dout(n381),.clk(gclk));
	jor g0119(.dina(w_n381_0[1]),.dinb(w_n273_60[1]),.dout(n382),.clk(gclk));
	jand g0120(.dina(n382),.dinb(n378),.dout(n383),.clk(gclk));
	jand g0121(.dina(w_n383_1[1]),.dinb(w_n281_62[2]),.dout(n384),.clk(gclk));
	jor g0122(.dina(w_shift0_56[2]),.dinb(w_a60_0[1]),.dout(n385),.clk(gclk));
	jor g0123(.dina(w_n269_56[2]),.dinb(w_a59_0[1]),.dout(n386),.clk(gclk));
	jand g0124(.dina(n386),.dinb(w_dff_B_1MK5rQm16_1),.dout(n387),.clk(gclk));
	jor g0125(.dina(w_n387_0[1]),.dinb(w_shift1_60[0]),.dout(n388),.clk(gclk));
	jor g0126(.dina(w_shift0_56[1]),.dinb(w_a58_0[1]),.dout(n389),.clk(gclk));
	jor g0127(.dina(w_n269_56[1]),.dinb(w_a57_0[1]),.dout(n390),.clk(gclk));
	jand g0128(.dina(n390),.dinb(w_dff_B_8ry3nHbt8_1),.dout(n391),.clk(gclk));
	jor g0129(.dina(w_n391_0[1]),.dinb(w_n273_60[0]),.dout(n392),.clk(gclk));
	jand g0130(.dina(n392),.dinb(n388),.dout(n393),.clk(gclk));
	jand g0131(.dina(w_n393_1[1]),.dinb(w_n267_62[2]),.dout(n394),.clk(gclk));
	jor g0132(.dina(n394),.dinb(n384),.dout(n395),.clk(gclk));
	jor g0133(.dina(w_shift0_56[0]),.dinb(w_a52_0[1]),.dout(n396),.clk(gclk));
	jor g0134(.dina(w_n269_56[0]),.dinb(w_a51_0[1]),.dout(n397),.clk(gclk));
	jand g0135(.dina(n397),.dinb(w_dff_B_qGz8nn0O6_1),.dout(n398),.clk(gclk));
	jor g0136(.dina(w_n398_0[1]),.dinb(w_shift1_59[2]),.dout(n399),.clk(gclk));
	jor g0137(.dina(w_shift0_55[2]),.dinb(w_a50_0[1]),.dout(n400),.clk(gclk));
	jor g0138(.dina(w_n269_55[2]),.dinb(w_a49_0[1]),.dout(n401),.clk(gclk));
	jand g0139(.dina(n401),.dinb(w_dff_B_rGGKJFCI5_1),.dout(n402),.clk(gclk));
	jor g0140(.dina(w_n402_0[1]),.dinb(w_n273_59[2]),.dout(n403),.clk(gclk));
	jand g0141(.dina(n403),.dinb(n399),.dout(n404),.clk(gclk));
	jand g0142(.dina(w_n404_1[1]),.dinb(w_n292_62[2]),.dout(n405),.clk(gclk));
	jor g0143(.dina(w_dff_B_YzMLCC1i0_0),.dinb(n395),.dout(n406),.clk(gclk));
	jor g0144(.dina(n406),.dinb(w_dff_B_zEG94JNY7_1),.dout(n407),.clk(gclk));
	jand g0145(.dina(w_n407_1[1]),.dinb(w_n364_63[1]),.dout(n408),.clk(gclk));
	jor g0146(.dina(n408),.dinb(n363),.dout(n409),.clk(gclk));
	jand g0147(.dina(w_shift5_0[0]),.dinb(w_shift4_0[0]),.dout(n410),.clk(gclk));
	jor g0148(.dina(w_shift0_55[1]),.dinb(w_a12_0[1]),.dout(n411),.clk(gclk));
	jor g0149(.dina(w_n269_55[1]),.dinb(w_a11_0[1]),.dout(n412),.clk(gclk));
	jand g0150(.dina(n412),.dinb(w_dff_B_hHESg9fo8_1),.dout(n413),.clk(gclk));
	jor g0151(.dina(w_n413_0[1]),.dinb(w_shift1_59[1]),.dout(n414),.clk(gclk));
	jor g0152(.dina(w_shift0_55[0]),.dinb(w_a10_0[1]),.dout(n415),.clk(gclk));
	jor g0153(.dina(w_n269_55[0]),.dinb(w_a9_0[1]),.dout(n416),.clk(gclk));
	jand g0154(.dina(n416),.dinb(w_dff_B_EdOZ8SLX0_1),.dout(n417),.clk(gclk));
	jor g0155(.dina(w_n417_0[1]),.dinb(w_n273_59[1]),.dout(n418),.clk(gclk));
	jand g0156(.dina(n418),.dinb(n414),.dout(n419),.clk(gclk));
	jand g0157(.dina(w_n419_1[1]),.dinb(w_n267_62[1]),.dout(n420),.clk(gclk));
	jor g0158(.dina(w_shift0_54[2]),.dinb(w_a8_0[1]),.dout(n421),.clk(gclk));
	jor g0159(.dina(w_n269_54[2]),.dinb(w_a7_0[1]),.dout(n422),.clk(gclk));
	jand g0160(.dina(n422),.dinb(w_dff_B_qelqFzvL8_1),.dout(n423),.clk(gclk));
	jor g0161(.dina(w_n423_0[1]),.dinb(w_shift1_59[0]),.dout(n424),.clk(gclk));
	jor g0162(.dina(w_shift0_54[1]),.dinb(w_a6_0[1]),.dout(n425),.clk(gclk));
	jor g0163(.dina(w_n269_54[1]),.dinb(w_a5_0[1]),.dout(n426),.clk(gclk));
	jand g0164(.dina(n426),.dinb(w_dff_B_r7LsM7Df4_1),.dout(n427),.clk(gclk));
	jor g0165(.dina(w_n427_0[1]),.dinb(w_n273_59[0]),.dout(n428),.clk(gclk));
	jand g0166(.dina(n428),.dinb(n424),.dout(n429),.clk(gclk));
	jand g0167(.dina(w_n429_1[1]),.dinb(w_n281_62[1]),.dout(n430),.clk(gclk));
	jor g0168(.dina(w_shift0_54[0]),.dinb(w_a4_0[1]),.dout(n431),.clk(gclk));
	jor g0169(.dina(w_n269_54[0]),.dinb(w_a3_0[1]),.dout(n432),.clk(gclk));
	jand g0170(.dina(n432),.dinb(w_dff_B_e7wXA7DB3_1),.dout(n433),.clk(gclk));
	jor g0171(.dina(w_n433_0[1]),.dinb(w_shift1_58[2]),.dout(n434),.clk(gclk));
	jor g0172(.dina(w_shift0_53[2]),.dinb(w_a2_0[1]),.dout(n435),.clk(gclk));
	jor g0173(.dina(w_n269_53[2]),.dinb(w_a1_0[1]),.dout(n436),.clk(gclk));
	jand g0174(.dina(n436),.dinb(w_dff_B_Y1FGDnUK0_1),.dout(n437),.clk(gclk));
	jor g0175(.dina(w_n437_0[1]),.dinb(w_n273_58[2]),.dout(n438),.clk(gclk));
	jand g0176(.dina(n438),.dinb(n434),.dout(n439),.clk(gclk));
	jand g0177(.dina(w_n439_1[1]),.dinb(w_n292_62[1]),.dout(n440),.clk(gclk));
	jor g0178(.dina(n440),.dinb(n430),.dout(n441),.clk(gclk));
	jor g0179(.dina(w_shift0_53[1]),.dinb(w_a16_0[1]),.dout(n442),.clk(gclk));
	jor g0180(.dina(w_n269_53[1]),.dinb(w_a15_0[1]),.dout(n443),.clk(gclk));
	jand g0181(.dina(n443),.dinb(w_dff_B_LlIFSUYG1_1),.dout(n444),.clk(gclk));
	jor g0182(.dina(w_n444_0[1]),.dinb(w_shift1_58[1]),.dout(n445),.clk(gclk));
	jor g0183(.dina(w_shift0_53[0]),.dinb(w_a14_0[1]),.dout(n446),.clk(gclk));
	jor g0184(.dina(w_n269_53[0]),.dinb(w_a13_0[1]),.dout(n447),.clk(gclk));
	jand g0185(.dina(n447),.dinb(w_dff_B_psoYtpqQ6_1),.dout(n448),.clk(gclk));
	jor g0186(.dina(w_n448_0[1]),.dinb(w_n273_58[1]),.dout(n449),.clk(gclk));
	jand g0187(.dina(n449),.dinb(n445),.dout(n450),.clk(gclk));
	jand g0188(.dina(w_n450_1[1]),.dinb(w_n304_62[1]),.dout(n451),.clk(gclk));
	jor g0189(.dina(w_dff_B_AsSN8oxv0_0),.dinb(n441),.dout(n452),.clk(gclk));
	jor g0190(.dina(n452),.dinb(w_dff_B_BFVo2AC79_1),.dout(n453),.clk(gclk));
	jand g0191(.dina(w_n453_1[1]),.dinb(w_n410_63[1]),.dout(n454),.clk(gclk));
	jor g0192(.dina(w_dff_B_HpkFhe6A1_0),.dinb(n409),.dout(n455),.clk(gclk));
	jor g0193(.dina(n455),.dinb(w_dff_B_IqnWAkCL7_1),.dout(n456),.clk(gclk));
	jor g0194(.dina(w_n456_0[1]),.dinb(w_n263_63[1]),.dout(n457),.clk(gclk));
	jor g0195(.dina(w_shift0_52[2]),.dinb(w_a68_0[1]),.dout(n458),.clk(gclk));
	jor g0196(.dina(w_n269_52[2]),.dinb(w_a67_0[1]),.dout(n459),.clk(gclk));
	jand g0197(.dina(n459),.dinb(w_dff_B_gnnLsEbL7_1),.dout(n460),.clk(gclk));
	jor g0198(.dina(w_n460_0[1]),.dinb(w_shift1_58[0]),.dout(n461),.clk(gclk));
	jor g0199(.dina(w_shift0_52[1]),.dinb(w_a66_0[1]),.dout(n462),.clk(gclk));
	jor g0200(.dina(w_n269_52[1]),.dinb(w_a65_0[1]),.dout(n463),.clk(gclk));
	jand g0201(.dina(n463),.dinb(w_dff_B_wXVKtnh13_1),.dout(n464),.clk(gclk));
	jor g0202(.dina(w_n464_0[1]),.dinb(w_n273_58[0]),.dout(n465),.clk(gclk));
	jand g0203(.dina(n465),.dinb(n461),.dout(n466),.clk(gclk));
	jand g0204(.dina(w_n466_1[1]),.dinb(w_n292_62[0]),.dout(n467),.clk(gclk));
	jor g0205(.dina(w_shift0_52[0]),.dinb(w_a72_0[1]),.dout(n468),.clk(gclk));
	jor g0206(.dina(w_n269_52[0]),.dinb(w_a71_0[1]),.dout(n469),.clk(gclk));
	jand g0207(.dina(n469),.dinb(w_dff_B_sqwDOK3F5_1),.dout(n470),.clk(gclk));
	jor g0208(.dina(w_n470_0[1]),.dinb(w_shift1_57[2]),.dout(n471),.clk(gclk));
	jor g0209(.dina(w_shift0_51[2]),.dinb(w_a70_0[1]),.dout(n472),.clk(gclk));
	jor g0210(.dina(w_n269_51[2]),.dinb(w_a69_0[1]),.dout(n473),.clk(gclk));
	jand g0211(.dina(n473),.dinb(w_dff_B_xqLjxEhE3_1),.dout(n474),.clk(gclk));
	jor g0212(.dina(w_n474_0[1]),.dinb(w_n273_57[2]),.dout(n475),.clk(gclk));
	jand g0213(.dina(n475),.dinb(n471),.dout(n476),.clk(gclk));
	jand g0214(.dina(w_n476_1[1]),.dinb(w_n281_62[0]),.dout(n477),.clk(gclk));
	jor g0215(.dina(w_shift0_51[1]),.dinb(w_a76_0[1]),.dout(n478),.clk(gclk));
	jor g0216(.dina(w_n269_51[1]),.dinb(w_a75_0[1]),.dout(n479),.clk(gclk));
	jand g0217(.dina(n479),.dinb(w_dff_B_1erSQF5v5_1),.dout(n480),.clk(gclk));
	jor g0218(.dina(w_n480_0[1]),.dinb(w_shift1_57[1]),.dout(n481),.clk(gclk));
	jor g0219(.dina(w_shift0_51[0]),.dinb(w_a74_0[1]),.dout(n482),.clk(gclk));
	jor g0220(.dina(w_n269_51[0]),.dinb(w_a73_0[1]),.dout(n483),.clk(gclk));
	jand g0221(.dina(n483),.dinb(w_dff_B_8SdLIGhZ4_1),.dout(n484),.clk(gclk));
	jor g0222(.dina(w_n484_0[1]),.dinb(w_n273_57[1]),.dout(n485),.clk(gclk));
	jand g0223(.dina(n485),.dinb(n481),.dout(n486),.clk(gclk));
	jand g0224(.dina(w_n486_1[1]),.dinb(w_n267_62[0]),.dout(n487),.clk(gclk));
	jor g0225(.dina(n487),.dinb(n477),.dout(n488),.clk(gclk));
	jor g0226(.dina(w_shift0_50[2]),.dinb(w_a80_0[1]),.dout(n489),.clk(gclk));
	jor g0227(.dina(w_n269_50[2]),.dinb(w_a79_0[1]),.dout(n490),.clk(gclk));
	jand g0228(.dina(n490),.dinb(w_dff_B_qDiElXBG9_1),.dout(n491),.clk(gclk));
	jor g0229(.dina(w_n491_0[1]),.dinb(w_shift1_57[0]),.dout(n492),.clk(gclk));
	jor g0230(.dina(w_shift0_50[1]),.dinb(w_a78_0[1]),.dout(n493),.clk(gclk));
	jor g0231(.dina(w_n269_50[1]),.dinb(w_a77_0[1]),.dout(n494),.clk(gclk));
	jand g0232(.dina(n494),.dinb(w_dff_B_LvNxJLXv2_1),.dout(n495),.clk(gclk));
	jor g0233(.dina(w_n495_0[1]),.dinb(w_n273_57[0]),.dout(n496),.clk(gclk));
	jand g0234(.dina(n496),.dinb(n492),.dout(n497),.clk(gclk));
	jand g0235(.dina(w_n497_1[1]),.dinb(w_n304_62[0]),.dout(n498),.clk(gclk));
	jor g0236(.dina(w_dff_B_i4pJGpHe3_0),.dinb(n488),.dout(n499),.clk(gclk));
	jor g0237(.dina(n499),.dinb(w_dff_B_3JQdqvgr9_1),.dout(n500),.clk(gclk));
	jand g0238(.dina(w_n500_1[1]),.dinb(w_n410_63[0]),.dout(n501),.clk(gclk));
	jor g0239(.dina(w_shift0_50[0]),.dinb(w_a100_0[1]),.dout(n502),.clk(gclk));
	jor g0240(.dina(w_n269_50[0]),.dinb(w_a99_0[1]),.dout(n503),.clk(gclk));
	jand g0241(.dina(n503),.dinb(w_dff_B_oANUBuw89_1),.dout(n504),.clk(gclk));
	jor g0242(.dina(w_n504_0[1]),.dinb(w_shift1_56[2]),.dout(n505),.clk(gclk));
	jor g0243(.dina(w_shift0_49[2]),.dinb(w_a98_0[1]),.dout(n506),.clk(gclk));
	jor g0244(.dina(w_n269_49[2]),.dinb(w_a97_0[1]),.dout(n507),.clk(gclk));
	jand g0245(.dina(n507),.dinb(w_dff_B_ZtYCSpfs0_1),.dout(n508),.clk(gclk));
	jor g0246(.dina(w_n508_0[1]),.dinb(w_n273_56[2]),.dout(n509),.clk(gclk));
	jand g0247(.dina(n509),.dinb(n505),.dout(n510),.clk(gclk));
	jand g0248(.dina(w_n510_1[1]),.dinb(w_n292_61[2]),.dout(n511),.clk(gclk));
	jor g0249(.dina(w_shift0_49[1]),.dinb(w_a104_0[1]),.dout(n512),.clk(gclk));
	jor g0250(.dina(w_n269_49[1]),.dinb(w_a103_0[1]),.dout(n513),.clk(gclk));
	jand g0251(.dina(n513),.dinb(w_dff_B_0JQMoqEd2_1),.dout(n514),.clk(gclk));
	jor g0252(.dina(w_n514_0[1]),.dinb(w_shift1_56[1]),.dout(n515),.clk(gclk));
	jor g0253(.dina(w_shift0_49[0]),.dinb(w_a102_0[1]),.dout(n516),.clk(gclk));
	jor g0254(.dina(w_n269_49[0]),.dinb(w_a101_0[1]),.dout(n517),.clk(gclk));
	jand g0255(.dina(n517),.dinb(w_dff_B_DBajLoEy0_1),.dout(n518),.clk(gclk));
	jor g0256(.dina(w_n518_0[1]),.dinb(w_n273_56[1]),.dout(n519),.clk(gclk));
	jand g0257(.dina(n519),.dinb(n515),.dout(n520),.clk(gclk));
	jand g0258(.dina(w_n520_1[1]),.dinb(w_n281_61[2]),.dout(n521),.clk(gclk));
	jor g0259(.dina(w_shift0_48[2]),.dinb(w_a108_0[1]),.dout(n522),.clk(gclk));
	jor g0260(.dina(w_n269_48[2]),.dinb(w_a107_0[1]),.dout(n523),.clk(gclk));
	jand g0261(.dina(n523),.dinb(w_dff_B_qxZUuMrc2_1),.dout(n524),.clk(gclk));
	jor g0262(.dina(w_n524_0[1]),.dinb(w_shift1_56[0]),.dout(n525),.clk(gclk));
	jor g0263(.dina(w_shift0_48[1]),.dinb(w_a106_0[1]),.dout(n526),.clk(gclk));
	jor g0264(.dina(w_n269_48[1]),.dinb(w_a105_0[1]),.dout(n527),.clk(gclk));
	jand g0265(.dina(n527),.dinb(w_dff_B_bUuUbKk52_1),.dout(n528),.clk(gclk));
	jor g0266(.dina(w_n528_0[1]),.dinb(w_n273_56[0]),.dout(n529),.clk(gclk));
	jand g0267(.dina(n529),.dinb(n525),.dout(n530),.clk(gclk));
	jand g0268(.dina(w_n530_1[1]),.dinb(w_n267_61[2]),.dout(n531),.clk(gclk));
	jor g0269(.dina(n531),.dinb(n521),.dout(n532),.clk(gclk));
	jor g0270(.dina(w_shift0_48[0]),.dinb(w_a112_0[1]),.dout(n533),.clk(gclk));
	jor g0271(.dina(w_n269_48[0]),.dinb(w_a111_0[1]),.dout(n534),.clk(gclk));
	jand g0272(.dina(n534),.dinb(w_dff_B_eNbCbCNd4_1),.dout(n535),.clk(gclk));
	jor g0273(.dina(w_n535_0[1]),.dinb(w_shift1_55[2]),.dout(n536),.clk(gclk));
	jor g0274(.dina(w_shift0_47[2]),.dinb(w_a110_0[1]),.dout(n537),.clk(gclk));
	jor g0275(.dina(w_n269_47[2]),.dinb(w_a109_0[1]),.dout(n538),.clk(gclk));
	jand g0276(.dina(n538),.dinb(w_dff_B_USEsFc4E6_1),.dout(n539),.clk(gclk));
	jor g0277(.dina(w_n539_0[1]),.dinb(w_n273_55[2]),.dout(n540),.clk(gclk));
	jand g0278(.dina(n540),.dinb(n536),.dout(n541),.clk(gclk));
	jand g0279(.dina(w_n541_1[1]),.dinb(w_n304_61[2]),.dout(n542),.clk(gclk));
	jor g0280(.dina(w_dff_B_WaH1Qvu22_0),.dinb(n532),.dout(n543),.clk(gclk));
	jor g0281(.dina(n543),.dinb(w_dff_B_wrKJCLHE2_1),.dout(n544),.clk(gclk));
	jand g0282(.dina(w_n544_1[1]),.dinb(w_n319_63[0]),.dout(n545),.clk(gclk));
	jor g0283(.dina(w_shift0_47[1]),.dinb(w_a92_0[1]),.dout(n546),.clk(gclk));
	jor g0284(.dina(w_n269_47[1]),.dinb(w_a91_0[1]),.dout(n547),.clk(gclk));
	jand g0285(.dina(n547),.dinb(w_dff_B_lrsiFJkx2_1),.dout(n548),.clk(gclk));
	jor g0286(.dina(w_n548_0[1]),.dinb(w_shift1_55[1]),.dout(n549),.clk(gclk));
	jor g0287(.dina(w_shift0_47[0]),.dinb(w_a90_0[1]),.dout(n550),.clk(gclk));
	jor g0288(.dina(w_n269_47[0]),.dinb(w_a89_0[1]),.dout(n551),.clk(gclk));
	jand g0289(.dina(n551),.dinb(w_dff_B_3XYmQ7xa1_1),.dout(n552),.clk(gclk));
	jor g0290(.dina(w_n552_0[1]),.dinb(w_n273_55[1]),.dout(n553),.clk(gclk));
	jand g0291(.dina(n553),.dinb(n549),.dout(n554),.clk(gclk));
	jand g0292(.dina(w_n554_1[1]),.dinb(w_n267_61[1]),.dout(n555),.clk(gclk));
	jor g0293(.dina(w_shift0_46[2]),.dinb(w_a88_0[1]),.dout(n556),.clk(gclk));
	jor g0294(.dina(w_n269_46[2]),.dinb(w_a87_0[1]),.dout(n557),.clk(gclk));
	jand g0295(.dina(n557),.dinb(w_dff_B_kbso0kek4_1),.dout(n558),.clk(gclk));
	jor g0296(.dina(w_n558_0[1]),.dinb(w_shift1_55[0]),.dout(n559),.clk(gclk));
	jor g0297(.dina(w_shift0_46[1]),.dinb(w_a86_0[1]),.dout(n560),.clk(gclk));
	jor g0298(.dina(w_n269_46[1]),.dinb(w_a85_0[1]),.dout(n561),.clk(gclk));
	jand g0299(.dina(n561),.dinb(w_dff_B_a2qEd9k26_1),.dout(n562),.clk(gclk));
	jor g0300(.dina(w_n562_0[1]),.dinb(w_n273_55[0]),.dout(n563),.clk(gclk));
	jand g0301(.dina(n563),.dinb(n559),.dout(n564),.clk(gclk));
	jand g0302(.dina(w_n564_1[1]),.dinb(w_n281_61[1]),.dout(n565),.clk(gclk));
	jor g0303(.dina(w_shift0_46[0]),.dinb(w_a84_0[1]),.dout(n566),.clk(gclk));
	jor g0304(.dina(w_n269_46[0]),.dinb(w_a83_0[1]),.dout(n567),.clk(gclk));
	jand g0305(.dina(n567),.dinb(w_dff_B_KkZUlkQY5_1),.dout(n568),.clk(gclk));
	jor g0306(.dina(w_n568_0[1]),.dinb(w_shift1_54[2]),.dout(n569),.clk(gclk));
	jor g0307(.dina(w_shift0_45[2]),.dinb(w_a82_0[1]),.dout(n570),.clk(gclk));
	jor g0308(.dina(w_n269_45[2]),.dinb(w_a81_0[1]),.dout(n571),.clk(gclk));
	jand g0309(.dina(n571),.dinb(w_dff_B_gUpOzecm7_1),.dout(n572),.clk(gclk));
	jor g0310(.dina(w_n572_0[1]),.dinb(w_n273_54[2]),.dout(n573),.clk(gclk));
	jand g0311(.dina(n573),.dinb(n569),.dout(n574),.clk(gclk));
	jand g0312(.dina(w_n574_1[1]),.dinb(w_n292_61[1]),.dout(n575),.clk(gclk));
	jor g0313(.dina(n575),.dinb(n565),.dout(n576),.clk(gclk));
	jor g0314(.dina(w_shift0_45[1]),.dinb(w_a96_0[1]),.dout(n577),.clk(gclk));
	jor g0315(.dina(w_n269_45[1]),.dinb(w_a95_0[1]),.dout(n578),.clk(gclk));
	jand g0316(.dina(n578),.dinb(w_dff_B_kMwsZSDe0_1),.dout(n579),.clk(gclk));
	jor g0317(.dina(w_n579_0[1]),.dinb(w_shift1_54[1]),.dout(n580),.clk(gclk));
	jor g0318(.dina(w_shift0_45[0]),.dinb(w_a94_0[1]),.dout(n581),.clk(gclk));
	jor g0319(.dina(w_n269_45[0]),.dinb(w_a93_0[1]),.dout(n582),.clk(gclk));
	jand g0320(.dina(n582),.dinb(w_dff_B_RDrOvlHB2_1),.dout(n583),.clk(gclk));
	jor g0321(.dina(w_n583_0[1]),.dinb(w_n273_54[1]),.dout(n584),.clk(gclk));
	jand g0322(.dina(n584),.dinb(n580),.dout(n585),.clk(gclk));
	jand g0323(.dina(w_n585_1[1]),.dinb(w_n304_61[1]),.dout(n586),.clk(gclk));
	jor g0324(.dina(w_dff_B_J66uxfix0_0),.dinb(n576),.dout(n587),.clk(gclk));
	jor g0325(.dina(n587),.dinb(w_dff_B_9yHQ4G319_1),.dout(n588),.clk(gclk));
	jand g0326(.dina(w_n588_1[1]),.dinb(w_n265_63[0]),.dout(n589),.clk(gclk));
	jor g0327(.dina(n589),.dinb(n545),.dout(n590),.clk(gclk));
	jor g0328(.dina(w_shift0_44[2]),.dinb(w_a124_0[1]),.dout(n591),.clk(gclk));
	jor g0329(.dina(w_n269_44[2]),.dinb(w_a123_0[1]),.dout(n592),.clk(gclk));
	jand g0330(.dina(n592),.dinb(w_dff_B_0RsxGrIy5_1),.dout(n593),.clk(gclk));
	jor g0331(.dina(w_n593_0[1]),.dinb(w_shift1_54[0]),.dout(n594),.clk(gclk));
	jor g0332(.dina(w_shift0_44[1]),.dinb(w_a122_0[1]),.dout(n595),.clk(gclk));
	jor g0333(.dina(w_n269_44[1]),.dinb(w_a121_0[1]),.dout(n596),.clk(gclk));
	jand g0334(.dina(n596),.dinb(w_dff_B_pBoU1aAC0_1),.dout(n597),.clk(gclk));
	jor g0335(.dina(w_n597_0[1]),.dinb(w_n273_54[0]),.dout(n598),.clk(gclk));
	jand g0336(.dina(n598),.dinb(n594),.dout(n599),.clk(gclk));
	jand g0337(.dina(w_n599_1[1]),.dinb(w_n267_61[0]),.dout(n600),.clk(gclk));
	jor g0338(.dina(w_shift0_44[0]),.dinb(w_a120_0[1]),.dout(n601),.clk(gclk));
	jor g0339(.dina(w_n269_44[0]),.dinb(w_a119_0[1]),.dout(n602),.clk(gclk));
	jand g0340(.dina(n602),.dinb(w_dff_B_G73nas932_1),.dout(n603),.clk(gclk));
	jor g0341(.dina(w_n603_0[1]),.dinb(w_shift1_53[2]),.dout(n604),.clk(gclk));
	jor g0342(.dina(w_shift0_43[2]),.dinb(w_a118_0[1]),.dout(n605),.clk(gclk));
	jor g0343(.dina(w_n269_43[2]),.dinb(w_a117_0[1]),.dout(n606),.clk(gclk));
	jand g0344(.dina(n606),.dinb(w_dff_B_oX8bH2f69_1),.dout(n607),.clk(gclk));
	jor g0345(.dina(w_n607_0[1]),.dinb(w_n273_53[2]),.dout(n608),.clk(gclk));
	jand g0346(.dina(n608),.dinb(n604),.dout(n609),.clk(gclk));
	jand g0347(.dina(w_n609_1[1]),.dinb(w_n281_61[0]),.dout(n610),.clk(gclk));
	jor g0348(.dina(w_shift0_43[1]),.dinb(w_a116_0[1]),.dout(n611),.clk(gclk));
	jor g0349(.dina(w_n269_43[1]),.dinb(w_a115_0[1]),.dout(n612),.clk(gclk));
	jand g0350(.dina(n612),.dinb(w_dff_B_Nhlo4skL5_1),.dout(n613),.clk(gclk));
	jor g0351(.dina(w_n613_0[1]),.dinb(w_shift1_53[1]),.dout(n614),.clk(gclk));
	jor g0352(.dina(w_shift0_43[0]),.dinb(w_a114_0[1]),.dout(n615),.clk(gclk));
	jor g0353(.dina(w_n269_43[0]),.dinb(w_a113_0[1]),.dout(n616),.clk(gclk));
	jand g0354(.dina(n616),.dinb(w_dff_B_DgWSqdmm5_1),.dout(n617),.clk(gclk));
	jor g0355(.dina(w_n617_0[1]),.dinb(w_n273_53[1]),.dout(n618),.clk(gclk));
	jand g0356(.dina(n618),.dinb(n614),.dout(n619),.clk(gclk));
	jand g0357(.dina(w_n619_1[1]),.dinb(w_n292_61[0]),.dout(n620),.clk(gclk));
	jor g0358(.dina(n620),.dinb(n610),.dout(n621),.clk(gclk));
	jor g0359(.dina(w_shift0_42[2]),.dinb(w_a0_0[1]),.dout(n622),.clk(gclk));
	jor g0360(.dina(w_n269_42[2]),.dinb(w_a127_0[1]),.dout(n623),.clk(gclk));
	jand g0361(.dina(n623),.dinb(w_dff_B_OXno1hik8_1),.dout(n624),.clk(gclk));
	jor g0362(.dina(w_n624_0[1]),.dinb(w_shift1_53[0]),.dout(n625),.clk(gclk));
	jor g0363(.dina(w_shift0_42[1]),.dinb(w_a126_0[1]),.dout(n626),.clk(gclk));
	jor g0364(.dina(w_n269_42[1]),.dinb(w_a125_0[1]),.dout(n627),.clk(gclk));
	jand g0365(.dina(n627),.dinb(w_dff_B_LxADl0g43_1),.dout(n628),.clk(gclk));
	jor g0366(.dina(w_n628_0[1]),.dinb(w_n273_53[0]),.dout(n629),.clk(gclk));
	jand g0367(.dina(n629),.dinb(n625),.dout(n630),.clk(gclk));
	jand g0368(.dina(w_n630_1[1]),.dinb(w_n304_61[0]),.dout(n631),.clk(gclk));
	jor g0369(.dina(w_dff_B_PoFkE5wX0_0),.dinb(n621),.dout(n632),.clk(gclk));
	jor g0370(.dina(n632),.dinb(w_dff_B_T9dm59OW2_1),.dout(n633),.clk(gclk));
	jand g0371(.dina(w_n633_1[1]),.dinb(w_n364_63[0]),.dout(n634),.clk(gclk));
	jor g0372(.dina(w_dff_B_xuHcFHr59_0),.dinb(n590),.dout(n635),.clk(gclk));
	jor g0373(.dina(n635),.dinb(w_dff_B_UCm236lc9_1),.dout(n636),.clk(gclk));
	jor g0374(.dina(w_n636_0[1]),.dinb(w_shift6_63[1]),.dout(n637),.clk(gclk));
	jand g0375(.dina(n637),.dinb(n457),.dout(result0),.clk(gclk));
	jor g0376(.dina(w_shift0_42[0]),.dinb(w_a61_0[0]),.dout(n639),.clk(gclk));
	jor g0377(.dina(w_n269_42[0]),.dinb(w_a60_0[0]),.dout(n640),.clk(gclk));
	jand g0378(.dina(n640),.dinb(w_dff_B_0oLZnUPh4_1),.dout(n641),.clk(gclk));
	jand g0379(.dina(w_n641_0[1]),.dinb(w_n273_52[2]),.dout(n642),.clk(gclk));
	jor g0380(.dina(w_shift0_41[2]),.dinb(w_a59_0[0]),.dout(n643),.clk(gclk));
	jor g0381(.dina(w_n269_41[2]),.dinb(w_a58_0[0]),.dout(n644),.clk(gclk));
	jand g0382(.dina(n644),.dinb(w_dff_B_HKuzR6c52_1),.dout(n645),.clk(gclk));
	jand g0383(.dina(w_n645_0[1]),.dinb(w_shift1_52[2]),.dout(n646),.clk(gclk));
	jor g0384(.dina(n646),.dinb(n642),.dout(n647),.clk(gclk));
	jand g0385(.dina(w_n647_1[1]),.dinb(w_n267_60[2]),.dout(n648),.clk(gclk));
	jor g0386(.dina(w_shift0_41[1]),.dinb(w_a57_0[0]),.dout(n649),.clk(gclk));
	jor g0387(.dina(w_n269_41[1]),.dinb(w_a56_0[0]),.dout(n650),.clk(gclk));
	jand g0388(.dina(n650),.dinb(w_dff_B_innup2oD0_1),.dout(n651),.clk(gclk));
	jand g0389(.dina(w_n651_0[1]),.dinb(w_n273_52[1]),.dout(n652),.clk(gclk));
	jor g0390(.dina(w_shift0_41[0]),.dinb(w_a55_0[0]),.dout(n653),.clk(gclk));
	jor g0391(.dina(w_n269_41[0]),.dinb(w_a54_0[0]),.dout(n654),.clk(gclk));
	jand g0392(.dina(n654),.dinb(w_dff_B_tfJFhTxG8_1),.dout(n655),.clk(gclk));
	jand g0393(.dina(w_n655_0[1]),.dinb(w_shift1_52[1]),.dout(n656),.clk(gclk));
	jor g0394(.dina(n656),.dinb(n652),.dout(n657),.clk(gclk));
	jand g0395(.dina(w_n657_1[1]),.dinb(w_n281_60[2]),.dout(n658),.clk(gclk));
	jor g0396(.dina(w_shift0_40[2]),.dinb(w_a53_0[0]),.dout(n659),.clk(gclk));
	jor g0397(.dina(w_n269_40[2]),.dinb(w_a52_0[0]),.dout(n660),.clk(gclk));
	jand g0398(.dina(n660),.dinb(w_dff_B_SLXi6sqx0_1),.dout(n661),.clk(gclk));
	jand g0399(.dina(w_n661_0[1]),.dinb(w_n273_52[0]),.dout(n662),.clk(gclk));
	jor g0400(.dina(w_shift0_40[1]),.dinb(w_a51_0[0]),.dout(n663),.clk(gclk));
	jor g0401(.dina(w_n269_40[1]),.dinb(w_a50_0[0]),.dout(n664),.clk(gclk));
	jand g0402(.dina(n664),.dinb(w_dff_B_PK6M6bQk2_1),.dout(n665),.clk(gclk));
	jand g0403(.dina(w_n665_0[1]),.dinb(w_shift1_52[0]),.dout(n666),.clk(gclk));
	jor g0404(.dina(n666),.dinb(n662),.dout(n667),.clk(gclk));
	jand g0405(.dina(w_n667_1[1]),.dinb(w_n292_60[2]),.dout(n668),.clk(gclk));
	jor g0406(.dina(n668),.dinb(n658),.dout(n669),.clk(gclk));
	jor g0407(.dina(w_shift0_40[0]),.dinb(w_a65_0[0]),.dout(n670),.clk(gclk));
	jor g0408(.dina(w_n269_40[0]),.dinb(w_a64_0[0]),.dout(n671),.clk(gclk));
	jand g0409(.dina(n671),.dinb(w_dff_B_sqLFKCT85_1),.dout(n672),.clk(gclk));
	jand g0410(.dina(w_n672_0[1]),.dinb(w_n273_51[2]),.dout(n673),.clk(gclk));
	jor g0411(.dina(w_shift0_39[2]),.dinb(w_a63_0[0]),.dout(n674),.clk(gclk));
	jor g0412(.dina(w_n269_39[2]),.dinb(w_a62_0[0]),.dout(n675),.clk(gclk));
	jand g0413(.dina(n675),.dinb(w_dff_B_v2guYC8y6_1),.dout(n676),.clk(gclk));
	jand g0414(.dina(w_n676_0[1]),.dinb(w_shift1_51[2]),.dout(n677),.clk(gclk));
	jor g0415(.dina(n677),.dinb(n673),.dout(n678),.clk(gclk));
	jand g0416(.dina(w_n678_1[1]),.dinb(w_n304_60[2]),.dout(n679),.clk(gclk));
	jor g0417(.dina(w_dff_B_poR6M3NX3_0),.dinb(n669),.dout(n680),.clk(gclk));
	jor g0418(.dina(n680),.dinb(w_dff_B_5U4XzmXQ9_1),.dout(n681),.clk(gclk));
	jand g0419(.dina(w_n681_1[1]),.dinb(w_n364_62[2]),.dout(n682),.clk(gclk));
	jor g0420(.dina(w_shift0_39[1]),.dinb(w_a21_0[0]),.dout(n683),.clk(gclk));
	jor g0421(.dina(w_n269_39[1]),.dinb(w_a20_0[0]),.dout(n684),.clk(gclk));
	jand g0422(.dina(n684),.dinb(w_dff_B_a5mabnqU6_1),.dout(n685),.clk(gclk));
	jand g0423(.dina(w_n685_0[1]),.dinb(w_n273_51[1]),.dout(n686),.clk(gclk));
	jor g0424(.dina(w_shift0_39[0]),.dinb(w_a19_0[0]),.dout(n687),.clk(gclk));
	jor g0425(.dina(w_n269_39[0]),.dinb(w_a18_0[0]),.dout(n688),.clk(gclk));
	jand g0426(.dina(n688),.dinb(w_dff_B_MFGGkqzk7_1),.dout(n689),.clk(gclk));
	jand g0427(.dina(w_n689_0[1]),.dinb(w_shift1_51[1]),.dout(n690),.clk(gclk));
	jor g0428(.dina(n690),.dinb(n686),.dout(n691),.clk(gclk));
	jand g0429(.dina(w_n691_1[1]),.dinb(w_n292_60[1]),.dout(n692),.clk(gclk));
	jor g0430(.dina(w_shift0_38[2]),.dinb(w_a25_0[0]),.dout(n693),.clk(gclk));
	jor g0431(.dina(w_n269_38[2]),.dinb(w_a24_0[0]),.dout(n694),.clk(gclk));
	jand g0432(.dina(n694),.dinb(w_dff_B_xpd5mGRp3_1),.dout(n695),.clk(gclk));
	jand g0433(.dina(w_n695_0[1]),.dinb(w_n273_51[0]),.dout(n696),.clk(gclk));
	jor g0434(.dina(w_shift0_38[1]),.dinb(w_a23_0[0]),.dout(n697),.clk(gclk));
	jor g0435(.dina(w_n269_38[1]),.dinb(w_a22_0[0]),.dout(n698),.clk(gclk));
	jand g0436(.dina(n698),.dinb(w_dff_B_o7JVhuzP9_1),.dout(n699),.clk(gclk));
	jand g0437(.dina(w_n699_0[1]),.dinb(w_shift1_51[0]),.dout(n700),.clk(gclk));
	jor g0438(.dina(n700),.dinb(n696),.dout(n701),.clk(gclk));
	jand g0439(.dina(w_n701_1[1]),.dinb(w_n281_60[1]),.dout(n702),.clk(gclk));
	jor g0440(.dina(w_shift0_38[0]),.dinb(w_a29_0[0]),.dout(n703),.clk(gclk));
	jor g0441(.dina(w_n269_38[0]),.dinb(w_a28_0[0]),.dout(n704),.clk(gclk));
	jand g0442(.dina(n704),.dinb(w_dff_B_TF8VuoJz5_1),.dout(n705),.clk(gclk));
	jand g0443(.dina(w_n705_0[1]),.dinb(w_n273_50[2]),.dout(n706),.clk(gclk));
	jor g0444(.dina(w_shift0_37[2]),.dinb(w_a27_0[0]),.dout(n707),.clk(gclk));
	jor g0445(.dina(w_n269_37[2]),.dinb(w_a26_0[0]),.dout(n708),.clk(gclk));
	jand g0446(.dina(n708),.dinb(w_dff_B_Pj71flbm8_1),.dout(n709),.clk(gclk));
	jand g0447(.dina(w_n709_0[1]),.dinb(w_shift1_50[2]),.dout(n710),.clk(gclk));
	jor g0448(.dina(n710),.dinb(n706),.dout(n711),.clk(gclk));
	jand g0449(.dina(w_n711_1[1]),.dinb(w_n267_60[1]),.dout(n712),.clk(gclk));
	jor g0450(.dina(n712),.dinb(n702),.dout(n713),.clk(gclk));
	jor g0451(.dina(w_shift0_37[1]),.dinb(w_a33_0[0]),.dout(n714),.clk(gclk));
	jor g0452(.dina(w_n269_37[1]),.dinb(w_a32_0[0]),.dout(n715),.clk(gclk));
	jand g0453(.dina(n715),.dinb(w_dff_B_tarZfy621_1),.dout(n716),.clk(gclk));
	jand g0454(.dina(w_n716_0[1]),.dinb(w_n273_50[1]),.dout(n717),.clk(gclk));
	jor g0455(.dina(w_shift0_37[0]),.dinb(w_a31_0[0]),.dout(n718),.clk(gclk));
	jor g0456(.dina(w_n269_37[0]),.dinb(w_a30_0[0]),.dout(n719),.clk(gclk));
	jand g0457(.dina(n719),.dinb(w_dff_B_DVmtjqsy4_1),.dout(n720),.clk(gclk));
	jand g0458(.dina(w_n720_0[1]),.dinb(w_shift1_50[1]),.dout(n721),.clk(gclk));
	jor g0459(.dina(n721),.dinb(n717),.dout(n722),.clk(gclk));
	jand g0460(.dina(w_n722_1[1]),.dinb(w_n304_60[1]),.dout(n723),.clk(gclk));
	jor g0461(.dina(w_dff_B_56NlZhYE3_0),.dinb(n713),.dout(n724),.clk(gclk));
	jor g0462(.dina(n724),.dinb(w_dff_B_fvmWPNeu8_1),.dout(n725),.clk(gclk));
	jand g0463(.dina(w_n725_1[1]),.dinb(w_n265_62[2]),.dout(n726),.clk(gclk));
	jor g0464(.dina(w_shift0_36[2]),.dinb(w_a17_0[0]),.dout(n727),.clk(gclk));
	jor g0465(.dina(w_n269_36[2]),.dinb(w_a16_0[0]),.dout(n728),.clk(gclk));
	jand g0466(.dina(n728),.dinb(w_dff_B_gXNcxvia2_1),.dout(n729),.clk(gclk));
	jand g0467(.dina(w_n729_0[1]),.dinb(w_n273_50[0]),.dout(n730),.clk(gclk));
	jor g0468(.dina(w_shift0_36[1]),.dinb(w_a15_0[0]),.dout(n731),.clk(gclk));
	jor g0469(.dina(w_n269_36[1]),.dinb(w_a14_0[0]),.dout(n732),.clk(gclk));
	jand g0470(.dina(n732),.dinb(w_dff_B_oi8DblKT5_1),.dout(n733),.clk(gclk));
	jand g0471(.dina(w_n733_0[1]),.dinb(w_shift1_50[0]),.dout(n734),.clk(gclk));
	jor g0472(.dina(n734),.dinb(n730),.dout(n735),.clk(gclk));
	jand g0473(.dina(w_n735_1[1]),.dinb(w_n304_60[0]),.dout(n736),.clk(gclk));
	jor g0474(.dina(w_shift0_36[0]),.dinb(w_a9_0[0]),.dout(n737),.clk(gclk));
	jor g0475(.dina(w_n269_36[0]),.dinb(w_a8_0[0]),.dout(n738),.clk(gclk));
	jand g0476(.dina(n738),.dinb(w_dff_B_uICq5SCD7_1),.dout(n739),.clk(gclk));
	jand g0477(.dina(w_n739_0[1]),.dinb(w_n273_49[2]),.dout(n740),.clk(gclk));
	jor g0478(.dina(w_shift0_35[2]),.dinb(w_a7_0[0]),.dout(n741),.clk(gclk));
	jor g0479(.dina(w_n269_35[2]),.dinb(w_a6_0[0]),.dout(n742),.clk(gclk));
	jand g0480(.dina(n742),.dinb(w_dff_B_6YxyaqYr2_1),.dout(n743),.clk(gclk));
	jand g0481(.dina(w_n743_0[1]),.dinb(w_shift1_49[2]),.dout(n744),.clk(gclk));
	jor g0482(.dina(n744),.dinb(n740),.dout(n745),.clk(gclk));
	jand g0483(.dina(w_n745_1[1]),.dinb(w_n281_60[0]),.dout(n746),.clk(gclk));
	jor g0484(.dina(w_shift0_35[1]),.dinb(w_a5_0[0]),.dout(n747),.clk(gclk));
	jor g0485(.dina(w_n269_35[1]),.dinb(w_a4_0[0]),.dout(n748),.clk(gclk));
	jand g0486(.dina(n748),.dinb(w_dff_B_aBi3tGKD9_1),.dout(n749),.clk(gclk));
	jand g0487(.dina(w_n749_0[1]),.dinb(w_n273_49[1]),.dout(n750),.clk(gclk));
	jor g0488(.dina(w_shift0_35[0]),.dinb(w_a3_0[0]),.dout(n751),.clk(gclk));
	jor g0489(.dina(w_n269_35[0]),.dinb(w_a2_0[0]),.dout(n752),.clk(gclk));
	jand g0490(.dina(n752),.dinb(w_dff_B_fsEUZG1w2_1),.dout(n753),.clk(gclk));
	jand g0491(.dina(w_n753_0[1]),.dinb(w_shift1_49[1]),.dout(n754),.clk(gclk));
	jor g0492(.dina(n754),.dinb(n750),.dout(n755),.clk(gclk));
	jand g0493(.dina(w_n755_1[1]),.dinb(w_n292_60[0]),.dout(n756),.clk(gclk));
	jor g0494(.dina(n756),.dinb(n746),.dout(n757),.clk(gclk));
	jor g0495(.dina(w_shift0_34[2]),.dinb(w_a13_0[0]),.dout(n758),.clk(gclk));
	jor g0496(.dina(w_n269_34[2]),.dinb(w_a12_0[0]),.dout(n759),.clk(gclk));
	jand g0497(.dina(n759),.dinb(w_dff_B_h6051X5M0_1),.dout(n760),.clk(gclk));
	jand g0498(.dina(w_n760_0[1]),.dinb(w_n273_49[0]),.dout(n761),.clk(gclk));
	jor g0499(.dina(w_shift0_34[1]),.dinb(w_a11_0[0]),.dout(n762),.clk(gclk));
	jor g0500(.dina(w_n269_34[1]),.dinb(w_a10_0[0]),.dout(n763),.clk(gclk));
	jand g0501(.dina(n763),.dinb(w_dff_B_DGgUZnJK3_1),.dout(n764),.clk(gclk));
	jand g0502(.dina(w_n764_0[1]),.dinb(w_shift1_49[0]),.dout(n765),.clk(gclk));
	jor g0503(.dina(n765),.dinb(n761),.dout(n766),.clk(gclk));
	jand g0504(.dina(w_n766_1[1]),.dinb(w_n267_60[0]),.dout(n767),.clk(gclk));
	jor g0505(.dina(w_dff_B_RbwjiVQc5_0),.dinb(n757),.dout(n768),.clk(gclk));
	jor g0506(.dina(n768),.dinb(w_dff_B_HBaastiB7_1),.dout(n769),.clk(gclk));
	jand g0507(.dina(w_n769_1[1]),.dinb(w_n410_62[2]),.dout(n770),.clk(gclk));
	jor g0508(.dina(n770),.dinb(n726),.dout(n771),.clk(gclk));
	jor g0509(.dina(w_shift0_34[0]),.dinb(w_a37_0[0]),.dout(n772),.clk(gclk));
	jor g0510(.dina(w_n269_34[0]),.dinb(w_a36_0[0]),.dout(n773),.clk(gclk));
	jand g0511(.dina(n773),.dinb(w_dff_B_sBdhvQYX3_1),.dout(n774),.clk(gclk));
	jand g0512(.dina(w_n774_0[1]),.dinb(w_n273_48[2]),.dout(n775),.clk(gclk));
	jor g0513(.dina(w_shift0_33[2]),.dinb(w_a35_0[0]),.dout(n776),.clk(gclk));
	jor g0514(.dina(w_n269_33[2]),.dinb(w_a34_0[0]),.dout(n777),.clk(gclk));
	jand g0515(.dina(n777),.dinb(w_dff_B_JkVSSvVk5_1),.dout(n778),.clk(gclk));
	jand g0516(.dina(w_n778_0[1]),.dinb(w_shift1_48[2]),.dout(n779),.clk(gclk));
	jor g0517(.dina(n779),.dinb(n775),.dout(n780),.clk(gclk));
	jand g0518(.dina(w_n780_1[1]),.dinb(w_n292_59[2]),.dout(n781),.clk(gclk));
	jor g0519(.dina(w_shift0_33[1]),.dinb(w_a39_0[0]),.dout(n782),.clk(gclk));
	jor g0520(.dina(w_n269_33[1]),.dinb(w_a38_0[0]),.dout(n783),.clk(gclk));
	jand g0521(.dina(n783),.dinb(w_dff_B_mYmJWWo27_1),.dout(n784),.clk(gclk));
	jor g0522(.dina(w_n784_0[1]),.dinb(w_n273_48[1]),.dout(n785),.clk(gclk));
	jor g0523(.dina(w_shift0_33[0]),.dinb(w_a41_0[0]),.dout(n786),.clk(gclk));
	jor g0524(.dina(w_n269_33[0]),.dinb(w_a40_0[0]),.dout(n787),.clk(gclk));
	jand g0525(.dina(n787),.dinb(w_dff_B_1VoqRzDF0_1),.dout(n788),.clk(gclk));
	jor g0526(.dina(w_n788_0[1]),.dinb(w_shift1_48[1]),.dout(n789),.clk(gclk));
	jand g0527(.dina(n789),.dinb(n785),.dout(n790),.clk(gclk));
	jand g0528(.dina(w_n790_1[1]),.dinb(w_n281_59[2]),.dout(n791),.clk(gclk));
	jor g0529(.dina(w_shift0_32[2]),.dinb(w_a45_0[0]),.dout(n792),.clk(gclk));
	jor g0530(.dina(w_n269_32[2]),.dinb(w_a44_0[0]),.dout(n793),.clk(gclk));
	jand g0531(.dina(n793),.dinb(w_dff_B_Np9QaPFa9_1),.dout(n794),.clk(gclk));
	jor g0532(.dina(w_n794_0[1]),.dinb(w_shift1_48[0]),.dout(n795),.clk(gclk));
	jor g0533(.dina(w_shift0_32[1]),.dinb(w_a43_0[0]),.dout(n796),.clk(gclk));
	jor g0534(.dina(w_n269_32[1]),.dinb(w_a42_0[0]),.dout(n797),.clk(gclk));
	jand g0535(.dina(n797),.dinb(w_dff_B_upysfaBQ0_1),.dout(n798),.clk(gclk));
	jor g0536(.dina(w_n798_0[1]),.dinb(w_n273_48[0]),.dout(n799),.clk(gclk));
	jand g0537(.dina(n799),.dinb(n795),.dout(n800),.clk(gclk));
	jand g0538(.dina(w_n800_1[1]),.dinb(w_n267_59[2]),.dout(n801),.clk(gclk));
	jor g0539(.dina(n801),.dinb(n791),.dout(n802),.clk(gclk));
	jor g0540(.dina(w_shift0_32[0]),.dinb(w_a49_0[0]),.dout(n803),.clk(gclk));
	jor g0541(.dina(w_n269_32[0]),.dinb(w_a48_0[0]),.dout(n804),.clk(gclk));
	jand g0542(.dina(n804),.dinb(w_dff_B_YqCEMGkj8_1),.dout(n805),.clk(gclk));
	jand g0543(.dina(w_n805_0[1]),.dinb(w_n273_47[2]),.dout(n806),.clk(gclk));
	jor g0544(.dina(w_shift0_31[2]),.dinb(w_a47_0[0]),.dout(n807),.clk(gclk));
	jor g0545(.dina(w_n269_31[2]),.dinb(w_a46_0[0]),.dout(n808),.clk(gclk));
	jand g0546(.dina(n808),.dinb(w_dff_B_PH0lI8405_1),.dout(n809),.clk(gclk));
	jand g0547(.dina(w_n809_0[1]),.dinb(w_shift1_47[2]),.dout(n810),.clk(gclk));
	jor g0548(.dina(n810),.dinb(n806),.dout(n811),.clk(gclk));
	jand g0549(.dina(w_n811_1[1]),.dinb(w_n304_59[2]),.dout(n812),.clk(gclk));
	jor g0550(.dina(w_dff_B_rOHLQUyL7_0),.dinb(n802),.dout(n813),.clk(gclk));
	jor g0551(.dina(n813),.dinb(w_dff_B_EhiM211Y3_1),.dout(n814),.clk(gclk));
	jand g0552(.dina(w_n814_1[1]),.dinb(w_n319_62[2]),.dout(n815),.clk(gclk));
	jor g0553(.dina(w_dff_B_gRp8Ggs88_0),.dinb(n771),.dout(n816),.clk(gclk));
	jor g0554(.dina(n816),.dinb(w_dff_B_E17iQHOA7_1),.dout(n817),.clk(gclk));
	jor g0555(.dina(w_n817_0[1]),.dinb(w_n263_63[0]),.dout(n818),.clk(gclk));
	jor g0556(.dina(w_shift0_31[1]),.dinb(w_a69_0[0]),.dout(n819),.clk(gclk));
	jor g0557(.dina(w_n269_31[1]),.dinb(w_a68_0[0]),.dout(n820),.clk(gclk));
	jand g0558(.dina(n820),.dinb(w_dff_B_ZwKVErzE1_1),.dout(n821),.clk(gclk));
	jand g0559(.dina(w_n821_0[1]),.dinb(w_n273_47[1]),.dout(n822),.clk(gclk));
	jor g0560(.dina(w_shift0_31[0]),.dinb(w_a67_0[0]),.dout(n823),.clk(gclk));
	jor g0561(.dina(w_n269_31[0]),.dinb(w_a66_0[0]),.dout(n824),.clk(gclk));
	jand g0562(.dina(n824),.dinb(w_dff_B_i0X0OPVY5_1),.dout(n825),.clk(gclk));
	jand g0563(.dina(w_n825_0[1]),.dinb(w_shift1_47[1]),.dout(n826),.clk(gclk));
	jor g0564(.dina(n826),.dinb(n822),.dout(n827),.clk(gclk));
	jand g0565(.dina(w_n827_1[1]),.dinb(w_n292_59[1]),.dout(n828),.clk(gclk));
	jor g0566(.dina(w_shift0_30[2]),.dinb(w_a73_0[0]),.dout(n829),.clk(gclk));
	jor g0567(.dina(w_n269_30[2]),.dinb(w_a72_0[0]),.dout(n830),.clk(gclk));
	jand g0568(.dina(n830),.dinb(w_dff_B_BcmFF8576_1),.dout(n831),.clk(gclk));
	jand g0569(.dina(w_n831_0[1]),.dinb(w_n273_47[0]),.dout(n832),.clk(gclk));
	jor g0570(.dina(w_shift0_30[1]),.dinb(w_a71_0[0]),.dout(n833),.clk(gclk));
	jor g0571(.dina(w_n269_30[1]),.dinb(w_a70_0[0]),.dout(n834),.clk(gclk));
	jand g0572(.dina(n834),.dinb(w_dff_B_Q6hzBaEe4_1),.dout(n835),.clk(gclk));
	jand g0573(.dina(w_n835_0[1]),.dinb(w_shift1_47[0]),.dout(n836),.clk(gclk));
	jor g0574(.dina(n836),.dinb(n832),.dout(n837),.clk(gclk));
	jand g0575(.dina(w_n837_1[1]),.dinb(w_n281_59[1]),.dout(n838),.clk(gclk));
	jor g0576(.dina(w_shift0_30[0]),.dinb(w_a77_0[0]),.dout(n839),.clk(gclk));
	jor g0577(.dina(w_n269_30[0]),.dinb(w_a76_0[0]),.dout(n840),.clk(gclk));
	jand g0578(.dina(n840),.dinb(w_dff_B_b1xub7d40_1),.dout(n841),.clk(gclk));
	jand g0579(.dina(w_n841_0[1]),.dinb(w_n273_46[2]),.dout(n842),.clk(gclk));
	jor g0580(.dina(w_shift0_29[2]),.dinb(w_a75_0[0]),.dout(n843),.clk(gclk));
	jor g0581(.dina(w_n269_29[2]),.dinb(w_a74_0[0]),.dout(n844),.clk(gclk));
	jand g0582(.dina(n844),.dinb(w_dff_B_qUAu1S6Q0_1),.dout(n845),.clk(gclk));
	jand g0583(.dina(w_n845_0[1]),.dinb(w_shift1_46[2]),.dout(n846),.clk(gclk));
	jor g0584(.dina(n846),.dinb(n842),.dout(n847),.clk(gclk));
	jand g0585(.dina(w_n847_1[1]),.dinb(w_n267_59[1]),.dout(n848),.clk(gclk));
	jor g0586(.dina(n848),.dinb(n838),.dout(n849),.clk(gclk));
	jor g0587(.dina(w_shift0_29[1]),.dinb(w_a81_0[0]),.dout(n850),.clk(gclk));
	jor g0588(.dina(w_n269_29[1]),.dinb(w_a80_0[0]),.dout(n851),.clk(gclk));
	jand g0589(.dina(n851),.dinb(w_dff_B_KImY48fm3_1),.dout(n852),.clk(gclk));
	jand g0590(.dina(w_n852_0[1]),.dinb(w_n273_46[1]),.dout(n853),.clk(gclk));
	jor g0591(.dina(w_shift0_29[0]),.dinb(w_a79_0[0]),.dout(n854),.clk(gclk));
	jor g0592(.dina(w_n269_29[0]),.dinb(w_a78_0[0]),.dout(n855),.clk(gclk));
	jand g0593(.dina(n855),.dinb(w_dff_B_lGKQzauE6_1),.dout(n856),.clk(gclk));
	jand g0594(.dina(w_n856_0[1]),.dinb(w_shift1_46[1]),.dout(n857),.clk(gclk));
	jor g0595(.dina(n857),.dinb(n853),.dout(n858),.clk(gclk));
	jand g0596(.dina(w_n858_1[1]),.dinb(w_n304_59[1]),.dout(n859),.clk(gclk));
	jor g0597(.dina(w_dff_B_kk7LeyAl5_0),.dinb(n849),.dout(n860),.clk(gclk));
	jor g0598(.dina(n860),.dinb(w_dff_B_NPOXfZNT9_1),.dout(n861),.clk(gclk));
	jand g0599(.dina(w_n861_1[1]),.dinb(w_n410_62[1]),.dout(n862),.clk(gclk));
	jor g0600(.dina(w_shift0_28[2]),.dinb(w_a101_0[0]),.dout(n863),.clk(gclk));
	jor g0601(.dina(w_n269_28[2]),.dinb(w_a100_0[0]),.dout(n864),.clk(gclk));
	jand g0602(.dina(n864),.dinb(w_dff_B_mXMNmnXD2_1),.dout(n865),.clk(gclk));
	jand g0603(.dina(w_n865_0[1]),.dinb(w_n273_46[0]),.dout(n866),.clk(gclk));
	jor g0604(.dina(w_shift0_28[1]),.dinb(w_a99_0[0]),.dout(n867),.clk(gclk));
	jor g0605(.dina(w_n269_28[1]),.dinb(w_a98_0[0]),.dout(n868),.clk(gclk));
	jand g0606(.dina(n868),.dinb(w_dff_B_py7Eagjp9_1),.dout(n869),.clk(gclk));
	jand g0607(.dina(w_n869_0[1]),.dinb(w_shift1_46[0]),.dout(n870),.clk(gclk));
	jor g0608(.dina(n870),.dinb(n866),.dout(n871),.clk(gclk));
	jand g0609(.dina(w_n871_1[1]),.dinb(w_n292_59[0]),.dout(n872),.clk(gclk));
	jor g0610(.dina(w_shift0_28[0]),.dinb(w_a105_0[0]),.dout(n873),.clk(gclk));
	jor g0611(.dina(w_n269_28[0]),.dinb(w_a104_0[0]),.dout(n874),.clk(gclk));
	jand g0612(.dina(n874),.dinb(w_dff_B_iPHr0LC45_1),.dout(n875),.clk(gclk));
	jand g0613(.dina(w_n875_0[1]),.dinb(w_n273_45[2]),.dout(n876),.clk(gclk));
	jor g0614(.dina(w_shift0_27[2]),.dinb(w_a103_0[0]),.dout(n877),.clk(gclk));
	jor g0615(.dina(w_n269_27[2]),.dinb(w_a102_0[0]),.dout(n878),.clk(gclk));
	jand g0616(.dina(n878),.dinb(w_dff_B_LzHuIvWe7_1),.dout(n879),.clk(gclk));
	jand g0617(.dina(w_n879_0[1]),.dinb(w_shift1_45[2]),.dout(n880),.clk(gclk));
	jor g0618(.dina(n880),.dinb(n876),.dout(n881),.clk(gclk));
	jand g0619(.dina(w_n881_1[1]),.dinb(w_n281_59[0]),.dout(n882),.clk(gclk));
	jor g0620(.dina(w_shift0_27[1]),.dinb(w_a109_0[0]),.dout(n883),.clk(gclk));
	jor g0621(.dina(w_n269_27[1]),.dinb(w_a108_0[0]),.dout(n884),.clk(gclk));
	jand g0622(.dina(n884),.dinb(w_dff_B_LyBW2d6f4_1),.dout(n885),.clk(gclk));
	jand g0623(.dina(w_n885_0[1]),.dinb(w_n273_45[1]),.dout(n886),.clk(gclk));
	jor g0624(.dina(w_shift0_27[0]),.dinb(w_a107_0[0]),.dout(n887),.clk(gclk));
	jor g0625(.dina(w_n269_27[0]),.dinb(w_a106_0[0]),.dout(n888),.clk(gclk));
	jand g0626(.dina(n888),.dinb(w_dff_B_1lzHYFyY3_1),.dout(n889),.clk(gclk));
	jand g0627(.dina(w_n889_0[1]),.dinb(w_shift1_45[1]),.dout(n890),.clk(gclk));
	jor g0628(.dina(n890),.dinb(n886),.dout(n891),.clk(gclk));
	jand g0629(.dina(w_n891_1[1]),.dinb(w_n267_59[0]),.dout(n892),.clk(gclk));
	jor g0630(.dina(n892),.dinb(n882),.dout(n893),.clk(gclk));
	jor g0631(.dina(w_shift0_26[2]),.dinb(w_a113_0[0]),.dout(n894),.clk(gclk));
	jor g0632(.dina(w_n269_26[2]),.dinb(w_a112_0[0]),.dout(n895),.clk(gclk));
	jand g0633(.dina(n895),.dinb(w_dff_B_745QdKaB0_1),.dout(n896),.clk(gclk));
	jand g0634(.dina(w_n896_0[1]),.dinb(w_n273_45[0]),.dout(n897),.clk(gclk));
	jor g0635(.dina(w_shift0_26[1]),.dinb(w_a111_0[0]),.dout(n898),.clk(gclk));
	jor g0636(.dina(w_n269_26[1]),.dinb(w_a110_0[0]),.dout(n899),.clk(gclk));
	jand g0637(.dina(n899),.dinb(w_dff_B_Qru46Pym3_1),.dout(n900),.clk(gclk));
	jand g0638(.dina(w_n900_0[1]),.dinb(w_shift1_45[0]),.dout(n901),.clk(gclk));
	jor g0639(.dina(n901),.dinb(n897),.dout(n902),.clk(gclk));
	jand g0640(.dina(w_n902_1[1]),.dinb(w_n304_59[0]),.dout(n903),.clk(gclk));
	jor g0641(.dina(w_dff_B_XJJ0p5Hv1_0),.dinb(n893),.dout(n904),.clk(gclk));
	jor g0642(.dina(n904),.dinb(w_dff_B_Mx9XTvKw1_1),.dout(n905),.clk(gclk));
	jand g0643(.dina(w_n905_1[1]),.dinb(w_n319_62[1]),.dout(n906),.clk(gclk));
	jor g0644(.dina(w_shift0_26[0]),.dinb(w_a85_0[0]),.dout(n907),.clk(gclk));
	jor g0645(.dina(w_n269_26[0]),.dinb(w_a84_0[0]),.dout(n908),.clk(gclk));
	jand g0646(.dina(n908),.dinb(w_dff_B_uvuIOWOm0_1),.dout(n909),.clk(gclk));
	jand g0647(.dina(w_n909_0[1]),.dinb(w_n273_44[2]),.dout(n910),.clk(gclk));
	jor g0648(.dina(w_shift0_25[2]),.dinb(w_a83_0[0]),.dout(n911),.clk(gclk));
	jor g0649(.dina(w_n269_25[2]),.dinb(w_a82_0[0]),.dout(n912),.clk(gclk));
	jand g0650(.dina(n912),.dinb(w_dff_B_42tADvHd7_1),.dout(n913),.clk(gclk));
	jand g0651(.dina(w_n913_0[1]),.dinb(w_shift1_44[2]),.dout(n914),.clk(gclk));
	jor g0652(.dina(n914),.dinb(n910),.dout(n915),.clk(gclk));
	jand g0653(.dina(w_n915_1[1]),.dinb(w_n292_58[2]),.dout(n916),.clk(gclk));
	jor g0654(.dina(w_shift0_25[1]),.dinb(w_a89_0[0]),.dout(n917),.clk(gclk));
	jor g0655(.dina(w_n269_25[1]),.dinb(w_a88_0[0]),.dout(n918),.clk(gclk));
	jand g0656(.dina(n918),.dinb(w_dff_B_NrGt6CJe2_1),.dout(n919),.clk(gclk));
	jand g0657(.dina(w_n919_0[1]),.dinb(w_n273_44[1]),.dout(n920),.clk(gclk));
	jor g0658(.dina(w_shift0_25[0]),.dinb(w_a87_0[0]),.dout(n921),.clk(gclk));
	jor g0659(.dina(w_n269_25[0]),.dinb(w_a86_0[0]),.dout(n922),.clk(gclk));
	jand g0660(.dina(n922),.dinb(w_dff_B_XT5fswlN8_1),.dout(n923),.clk(gclk));
	jand g0661(.dina(w_n923_0[1]),.dinb(w_shift1_44[1]),.dout(n924),.clk(gclk));
	jor g0662(.dina(n924),.dinb(n920),.dout(n925),.clk(gclk));
	jand g0663(.dina(w_n925_1[1]),.dinb(w_n281_58[2]),.dout(n926),.clk(gclk));
	jor g0664(.dina(w_shift0_24[2]),.dinb(w_a93_0[0]),.dout(n927),.clk(gclk));
	jor g0665(.dina(w_n269_24[2]),.dinb(w_a92_0[0]),.dout(n928),.clk(gclk));
	jand g0666(.dina(n928),.dinb(w_dff_B_yG764QYf5_1),.dout(n929),.clk(gclk));
	jand g0667(.dina(w_n929_0[1]),.dinb(w_n273_44[0]),.dout(n930),.clk(gclk));
	jor g0668(.dina(w_shift0_24[1]),.dinb(w_a91_0[0]),.dout(n931),.clk(gclk));
	jor g0669(.dina(w_n269_24[1]),.dinb(w_a90_0[0]),.dout(n932),.clk(gclk));
	jand g0670(.dina(n932),.dinb(w_dff_B_8NBshqAL6_1),.dout(n933),.clk(gclk));
	jand g0671(.dina(w_n933_0[1]),.dinb(w_shift1_44[0]),.dout(n934),.clk(gclk));
	jor g0672(.dina(n934),.dinb(n930),.dout(n935),.clk(gclk));
	jand g0673(.dina(w_n935_1[1]),.dinb(w_n267_58[2]),.dout(n936),.clk(gclk));
	jor g0674(.dina(n936),.dinb(n926),.dout(n937),.clk(gclk));
	jor g0675(.dina(w_shift0_24[0]),.dinb(w_a97_0[0]),.dout(n938),.clk(gclk));
	jor g0676(.dina(w_n269_24[0]),.dinb(w_a96_0[0]),.dout(n939),.clk(gclk));
	jand g0677(.dina(n939),.dinb(w_dff_B_8EZYNZap4_1),.dout(n940),.clk(gclk));
	jand g0678(.dina(w_n940_0[1]),.dinb(w_n273_43[2]),.dout(n941),.clk(gclk));
	jor g0679(.dina(w_shift0_23[2]),.dinb(w_a95_0[0]),.dout(n942),.clk(gclk));
	jor g0680(.dina(w_n269_23[2]),.dinb(w_a94_0[0]),.dout(n943),.clk(gclk));
	jand g0681(.dina(n943),.dinb(w_dff_B_WSLDAw9h6_1),.dout(n944),.clk(gclk));
	jand g0682(.dina(w_n944_0[1]),.dinb(w_shift1_43[2]),.dout(n945),.clk(gclk));
	jor g0683(.dina(n945),.dinb(n941),.dout(n946),.clk(gclk));
	jand g0684(.dina(w_n946_1[1]),.dinb(w_n304_58[2]),.dout(n947),.clk(gclk));
	jor g0685(.dina(w_dff_B_R3YJSblS2_0),.dinb(n937),.dout(n948),.clk(gclk));
	jor g0686(.dina(n948),.dinb(w_dff_B_pD3SBYZu7_1),.dout(n949),.clk(gclk));
	jand g0687(.dina(w_n949_1[1]),.dinb(w_n265_62[1]),.dout(n950),.clk(gclk));
	jor g0688(.dina(n950),.dinb(n906),.dout(n951),.clk(gclk));
	jor g0689(.dina(w_shift0_23[1]),.dinb(w_a125_0[0]),.dout(n952),.clk(gclk));
	jor g0690(.dina(w_n269_23[1]),.dinb(w_a124_0[0]),.dout(n953),.clk(gclk));
	jand g0691(.dina(n953),.dinb(w_dff_B_rF98fik62_1),.dout(n954),.clk(gclk));
	jand g0692(.dina(w_n954_0[1]),.dinb(w_n273_43[1]),.dout(n955),.clk(gclk));
	jor g0693(.dina(w_shift0_23[0]),.dinb(w_a123_0[0]),.dout(n956),.clk(gclk));
	jor g0694(.dina(w_n269_23[0]),.dinb(w_a122_0[0]),.dout(n957),.clk(gclk));
	jand g0695(.dina(n957),.dinb(w_dff_B_g2UrCknn7_1),.dout(n958),.clk(gclk));
	jand g0696(.dina(w_n958_0[1]),.dinb(w_shift1_43[1]),.dout(n959),.clk(gclk));
	jor g0697(.dina(n959),.dinb(n955),.dout(n960),.clk(gclk));
	jand g0698(.dina(w_n960_1[1]),.dinb(w_n267_58[1]),.dout(n961),.clk(gclk));
	jor g0699(.dina(w_shift0_22[2]),.dinb(w_a121_0[0]),.dout(n962),.clk(gclk));
	jor g0700(.dina(w_n269_22[2]),.dinb(w_a120_0[0]),.dout(n963),.clk(gclk));
	jand g0701(.dina(n963),.dinb(w_dff_B_K0Y4km6g5_1),.dout(n964),.clk(gclk));
	jand g0702(.dina(w_n964_0[1]),.dinb(w_n273_43[0]),.dout(n965),.clk(gclk));
	jor g0703(.dina(w_shift0_22[1]),.dinb(w_a119_0[0]),.dout(n966),.clk(gclk));
	jor g0704(.dina(w_n269_22[1]),.dinb(w_a118_0[0]),.dout(n967),.clk(gclk));
	jand g0705(.dina(n967),.dinb(w_dff_B_dyfUBpGV8_1),.dout(n968),.clk(gclk));
	jand g0706(.dina(w_n968_0[1]),.dinb(w_shift1_43[0]),.dout(n969),.clk(gclk));
	jor g0707(.dina(n969),.dinb(n965),.dout(n970),.clk(gclk));
	jand g0708(.dina(w_n970_1[1]),.dinb(w_n281_58[1]),.dout(n971),.clk(gclk));
	jor g0709(.dina(w_shift0_22[0]),.dinb(w_a117_0[0]),.dout(n972),.clk(gclk));
	jor g0710(.dina(w_n269_22[0]),.dinb(w_a116_0[0]),.dout(n973),.clk(gclk));
	jand g0711(.dina(n973),.dinb(w_dff_B_sskXJKkD8_1),.dout(n974),.clk(gclk));
	jand g0712(.dina(w_n974_0[1]),.dinb(w_n273_42[2]),.dout(n975),.clk(gclk));
	jor g0713(.dina(w_shift0_21[2]),.dinb(w_a115_0[0]),.dout(n976),.clk(gclk));
	jor g0714(.dina(w_n269_21[2]),.dinb(w_a114_0[0]),.dout(n977),.clk(gclk));
	jand g0715(.dina(n977),.dinb(w_dff_B_FIhTqrhf7_1),.dout(n978),.clk(gclk));
	jand g0716(.dina(w_n978_0[1]),.dinb(w_shift1_42[2]),.dout(n979),.clk(gclk));
	jor g0717(.dina(n979),.dinb(n975),.dout(n980),.clk(gclk));
	jand g0718(.dina(w_n980_1[1]),.dinb(w_n292_58[1]),.dout(n981),.clk(gclk));
	jor g0719(.dina(n981),.dinb(n971),.dout(n982),.clk(gclk));
	jor g0720(.dina(w_shift0_21[1]),.dinb(w_a1_0[0]),.dout(n983),.clk(gclk));
	jor g0721(.dina(w_n269_21[1]),.dinb(w_a0_0[0]),.dout(n984),.clk(gclk));
	jand g0722(.dina(n984),.dinb(w_dff_B_Wz80cizW6_1),.dout(n985),.clk(gclk));
	jand g0723(.dina(w_n985_0[1]),.dinb(w_n273_42[1]),.dout(n986),.clk(gclk));
	jor g0724(.dina(w_shift0_21[0]),.dinb(w_a127_0[0]),.dout(n987),.clk(gclk));
	jor g0725(.dina(w_n269_21[0]),.dinb(w_a126_0[0]),.dout(n988),.clk(gclk));
	jand g0726(.dina(n988),.dinb(w_dff_B_43V9h6ET3_1),.dout(n989),.clk(gclk));
	jand g0727(.dina(w_n989_0[1]),.dinb(w_shift1_42[1]),.dout(n990),.clk(gclk));
	jor g0728(.dina(n990),.dinb(n986),.dout(n991),.clk(gclk));
	jand g0729(.dina(w_n991_1[1]),.dinb(w_n304_58[1]),.dout(n992),.clk(gclk));
	jor g0730(.dina(w_dff_B_Tp0JK1jz6_0),.dinb(n982),.dout(n993),.clk(gclk));
	jor g0731(.dina(n993),.dinb(w_dff_B_n4s9MQBi8_1),.dout(n994),.clk(gclk));
	jand g0732(.dina(w_n994_1[1]),.dinb(w_n364_62[1]),.dout(n995),.clk(gclk));
	jor g0733(.dina(w_dff_B_cjYulRxp8_0),.dinb(n951),.dout(n996),.clk(gclk));
	jor g0734(.dina(n996),.dinb(w_dff_B_WfEiqaoK6_1),.dout(n997),.clk(gclk));
	jor g0735(.dina(w_n997_0[1]),.dinb(w_shift6_63[0]),.dout(n998),.clk(gclk));
	jand g0736(.dina(n998),.dinb(n818),.dout(result1),.clk(gclk));
	jor g0737(.dina(w_n357_0[0]),.dinb(w_shift1_42[0]),.dout(n1000),.clk(gclk));
	jor g0738(.dina(w_n342_0[0]),.dinb(w_n273_42[0]),.dout(n1001),.clk(gclk));
	jand g0739(.dina(n1001),.dinb(n1000),.dout(n1002),.clk(gclk));
	jand g0740(.dina(w_n1002_1[1]),.dinb(w_n267_58[0]),.dout(n1003),.clk(gclk));
	jor g0741(.dina(w_n332_0[0]),.dinb(w_n273_41[2]),.dout(n1004),.clk(gclk));
	jor g0742(.dina(w_n346_0[0]),.dinb(w_shift1_41[2]),.dout(n1005),.clk(gclk));
	jand g0743(.dina(n1005),.dinb(n1004),.dout(n1006),.clk(gclk));
	jand g0744(.dina(w_n1006_1[1]),.dinb(w_n281_58[0]),.dout(n1007),.clk(gclk));
	jor g0745(.dina(w_n322_0[0]),.dinb(w_n273_41[1]),.dout(n1008),.clk(gclk));
	jor g0746(.dina(w_n336_0[0]),.dinb(w_shift1_41[1]),.dout(n1009),.clk(gclk));
	jand g0747(.dina(n1009),.dinb(n1008),.dout(n1010),.clk(gclk));
	jand g0748(.dina(w_n1010_1[1]),.dinb(w_n292_58[0]),.dout(n1011),.clk(gclk));
	jor g0749(.dina(n1011),.dinb(n1007),.dout(n1012),.clk(gclk));
	jor g0750(.dina(w_n353_0[0]),.dinb(w_n273_41[0]),.dout(n1013),.clk(gclk));
	jor g0751(.dina(w_n402_0[0]),.dinb(w_shift1_41[0]),.dout(n1014),.clk(gclk));
	jand g0752(.dina(n1014),.dinb(n1013),.dout(n1015),.clk(gclk));
	jand g0753(.dina(w_n1015_1[1]),.dinb(w_n304_58[0]),.dout(n1016),.clk(gclk));
	jor g0754(.dina(w_dff_B_vGLAXmG71_0),.dinb(n1012),.dout(n1017),.clk(gclk));
	jor g0755(.dina(n1017),.dinb(w_dff_B_4OEclSdP1_1),.dout(n1018),.clk(gclk));
	jand g0756(.dina(w_n1018_1[1]),.dinb(w_n319_62[0]),.dout(n1019),.clk(gclk));
	jor g0757(.dina(w_n295_0[0]),.dinb(w_n273_40[2]),.dout(n1020),.clk(gclk));
	jor g0758(.dina(w_n288_0[0]),.dinb(w_shift1_40[2]),.dout(n1021),.clk(gclk));
	jand g0759(.dina(n1021),.dinb(n1020),.dout(n1022),.clk(gclk));
	jand g0760(.dina(w_n1022_1[1]),.dinb(w_n292_57[2]),.dout(n1023),.clk(gclk));
	jor g0761(.dina(w_n284_0[0]),.dinb(w_n273_40[1]),.dout(n1024),.clk(gclk));
	jor g0762(.dina(w_n276_0[0]),.dinb(w_shift1_40[1]),.dout(n1025),.clk(gclk));
	jand g0763(.dina(n1025),.dinb(n1024),.dout(n1026),.clk(gclk));
	jand g0764(.dina(w_n1026_1[1]),.dinb(w_n281_57[2]),.dout(n1027),.clk(gclk));
	jor g0765(.dina(w_n271_0[0]),.dinb(w_n273_40[0]),.dout(n1028),.clk(gclk));
	jor g0766(.dina(w_n311_0[0]),.dinb(w_shift1_40[0]),.dout(n1029),.clk(gclk));
	jand g0767(.dina(n1029),.dinb(n1028),.dout(n1030),.clk(gclk));
	jand g0768(.dina(w_n1030_1[1]),.dinb(w_n267_57[2]),.dout(n1031),.clk(gclk));
	jor g0769(.dina(n1031),.dinb(n1027),.dout(n1032),.clk(gclk));
	jor g0770(.dina(w_n307_0[0]),.dinb(w_n273_39[2]),.dout(n1033),.clk(gclk));
	jor g0771(.dina(w_n326_0[0]),.dinb(w_shift1_39[2]),.dout(n1034),.clk(gclk));
	jand g0772(.dina(n1034),.dinb(n1033),.dout(n1035),.clk(gclk));
	jand g0773(.dina(w_n1035_1[1]),.dinb(w_n304_57[2]),.dout(n1036),.clk(gclk));
	jor g0774(.dina(w_dff_B_BlDVNLBK7_0),.dinb(n1032),.dout(n1037),.clk(gclk));
	jor g0775(.dina(n1037),.dinb(w_dff_B_wnQLWcq32_1),.dout(n1038),.clk(gclk));
	jand g0776(.dina(w_n1038_1[1]),.dinb(w_n265_62[0]),.dout(n1039),.clk(gclk));
	jor g0777(.dina(w_n444_0[0]),.dinb(w_n273_39[1]),.dout(n1040),.clk(gclk));
	jor g0778(.dina(w_n299_0[0]),.dinb(w_shift1_39[1]),.dout(n1041),.clk(gclk));
	jand g0779(.dina(n1041),.dinb(n1040),.dout(n1042),.clk(gclk));
	jand g0780(.dina(w_n1042_1[1]),.dinb(w_n304_57[1]),.dout(n1043),.clk(gclk));
	jor g0781(.dina(w_n423_0[0]),.dinb(w_n273_39[0]),.dout(n1044),.clk(gclk));
	jor g0782(.dina(w_n417_0[0]),.dinb(w_shift1_39[0]),.dout(n1045),.clk(gclk));
	jand g0783(.dina(n1045),.dinb(n1044),.dout(n1046),.clk(gclk));
	jand g0784(.dina(w_n1046_1[1]),.dinb(w_n281_57[1]),.dout(n1047),.clk(gclk));
	jor g0785(.dina(w_n413_0[0]),.dinb(w_n273_38[2]),.dout(n1048),.clk(gclk));
	jor g0786(.dina(w_n448_0[0]),.dinb(w_shift1_38[2]),.dout(n1049),.clk(gclk));
	jand g0787(.dina(n1049),.dinb(n1048),.dout(n1050),.clk(gclk));
	jand g0788(.dina(w_n1050_1[1]),.dinb(w_n267_57[1]),.dout(n1051),.clk(gclk));
	jor g0789(.dina(n1051),.dinb(n1047),.dout(n1052),.clk(gclk));
	jor g0790(.dina(w_n433_0[0]),.dinb(w_n273_38[1]),.dout(n1053),.clk(gclk));
	jor g0791(.dina(w_n427_0[0]),.dinb(w_shift1_38[1]),.dout(n1054),.clk(gclk));
	jand g0792(.dina(n1054),.dinb(n1053),.dout(n1055),.clk(gclk));
	jand g0793(.dina(w_n1055_1[1]),.dinb(w_n292_57[1]),.dout(n1056),.clk(gclk));
	jor g0794(.dina(w_dff_B_xnBRSN2N3_0),.dinb(n1052),.dout(n1057),.clk(gclk));
	jor g0795(.dina(n1057),.dinb(w_dff_B_3KDdwdBk3_1),.dout(n1058),.clk(gclk));
	jand g0796(.dina(w_n1058_1[1]),.dinb(w_n410_62[0]),.dout(n1059),.clk(gclk));
	jor g0797(.dina(n1059),.dinb(n1039),.dout(n1060),.clk(gclk));
	jor g0798(.dina(w_n398_0[0]),.dinb(w_n273_38[0]),.dout(n1061),.clk(gclk));
	jor g0799(.dina(w_n381_0[0]),.dinb(w_shift1_38[0]),.dout(n1062),.clk(gclk));
	jand g0800(.dina(n1062),.dinb(n1061),.dout(n1063),.clk(gclk));
	jand g0801(.dina(w_n1063_1[1]),.dinb(w_n292_57[0]),.dout(n1064),.clk(gclk));
	jor g0802(.dina(w_n377_0[0]),.dinb(w_n273_37[2]),.dout(n1065),.clk(gclk));
	jor g0803(.dina(w_n391_0[0]),.dinb(w_shift1_37[2]),.dout(n1066),.clk(gclk));
	jand g0804(.dina(n1066),.dinb(n1065),.dout(n1067),.clk(gclk));
	jand g0805(.dina(w_n1067_1[1]),.dinb(w_n281_57[0]),.dout(n1068),.clk(gclk));
	jor g0806(.dina(w_n387_0[0]),.dinb(w_n273_37[1]),.dout(n1069),.clk(gclk));
	jor g0807(.dina(w_n371_0[0]),.dinb(w_shift1_37[1]),.dout(n1070),.clk(gclk));
	jand g0808(.dina(n1070),.dinb(n1069),.dout(n1071),.clk(gclk));
	jand g0809(.dina(w_n1071_1[1]),.dinb(w_n267_57[0]),.dout(n1072),.clk(gclk));
	jor g0810(.dina(n1072),.dinb(n1068),.dout(n1073),.clk(gclk));
	jor g0811(.dina(w_n367_0[0]),.dinb(w_n273_37[0]),.dout(n1074),.clk(gclk));
	jor g0812(.dina(w_n464_0[0]),.dinb(w_shift1_37[0]),.dout(n1075),.clk(gclk));
	jand g0813(.dina(n1075),.dinb(n1074),.dout(n1076),.clk(gclk));
	jand g0814(.dina(w_n1076_1[1]),.dinb(w_n304_57[0]),.dout(n1077),.clk(gclk));
	jor g0815(.dina(w_dff_B_hh4D6Ws52_0),.dinb(n1073),.dout(n1078),.clk(gclk));
	jor g0816(.dina(n1078),.dinb(w_dff_B_oMk1KklB2_1),.dout(n1079),.clk(gclk));
	jand g0817(.dina(w_n1079_1[1]),.dinb(w_n364_62[0]),.dout(n1080),.clk(gclk));
	jor g0818(.dina(w_dff_B_NanY4bA49_0),.dinb(n1060),.dout(n1081),.clk(gclk));
	jor g0819(.dina(n1081),.dinb(w_dff_B_ZbjPw7uh6_1),.dout(n1082),.clk(gclk));
	jor g0820(.dina(w_n1082_0[1]),.dinb(w_n263_62[2]),.dout(n1083),.clk(gclk));
	jor g0821(.dina(w_n480_0[0]),.dinb(w_n273_36[2]),.dout(n1084),.clk(gclk));
	jor g0822(.dina(w_n495_0[0]),.dinb(w_shift1_36[2]),.dout(n1085),.clk(gclk));
	jand g0823(.dina(n1085),.dinb(n1084),.dout(n1086),.clk(gclk));
	jand g0824(.dina(w_n1086_1[1]),.dinb(w_n267_56[2]),.dout(n1087),.clk(gclk));
	jor g0825(.dina(w_n470_0[0]),.dinb(w_n273_36[1]),.dout(n1088),.clk(gclk));
	jor g0826(.dina(w_n484_0[0]),.dinb(w_shift1_36[1]),.dout(n1089),.clk(gclk));
	jand g0827(.dina(n1089),.dinb(n1088),.dout(n1090),.clk(gclk));
	jand g0828(.dina(w_n1090_1[1]),.dinb(w_n281_56[2]),.dout(n1091),.clk(gclk));
	jor g0829(.dina(w_n460_0[0]),.dinb(w_n273_36[0]),.dout(n1092),.clk(gclk));
	jor g0830(.dina(w_n474_0[0]),.dinb(w_shift1_36[0]),.dout(n1093),.clk(gclk));
	jand g0831(.dina(n1093),.dinb(n1092),.dout(n1094),.clk(gclk));
	jand g0832(.dina(w_n1094_1[1]),.dinb(w_n292_56[2]),.dout(n1095),.clk(gclk));
	jor g0833(.dina(n1095),.dinb(n1091),.dout(n1096),.clk(gclk));
	jor g0834(.dina(w_n491_0[0]),.dinb(w_n273_35[2]),.dout(n1097),.clk(gclk));
	jor g0835(.dina(w_n572_0[0]),.dinb(w_shift1_35[2]),.dout(n1098),.clk(gclk));
	jand g0836(.dina(n1098),.dinb(n1097),.dout(n1099),.clk(gclk));
	jand g0837(.dina(w_n1099_1[1]),.dinb(w_n304_56[2]),.dout(n1100),.clk(gclk));
	jor g0838(.dina(w_dff_B_ZGWEitvM6_0),.dinb(n1096),.dout(n1101),.clk(gclk));
	jor g0839(.dina(n1101),.dinb(w_dff_B_ZhWqQhPZ3_1),.dout(n1102),.clk(gclk));
	jand g0840(.dina(w_n1102_1[1]),.dinb(w_n410_61[2]),.dout(n1103),.clk(gclk));
	jor g0841(.dina(w_n535_0[0]),.dinb(w_n273_35[1]),.dout(n1104),.clk(gclk));
	jor g0842(.dina(w_n617_0[0]),.dinb(w_shift1_35[1]),.dout(n1105),.clk(gclk));
	jand g0843(.dina(n1105),.dinb(n1104),.dout(n1106),.clk(gclk));
	jand g0844(.dina(w_n1106_1[1]),.dinb(w_n304_56[1]),.dout(n1107),.clk(gclk));
	jor g0845(.dina(w_n514_0[0]),.dinb(w_n273_35[0]),.dout(n1108),.clk(gclk));
	jor g0846(.dina(w_n528_0[0]),.dinb(w_shift1_35[0]),.dout(n1109),.clk(gclk));
	jand g0847(.dina(n1109),.dinb(n1108),.dout(n1110),.clk(gclk));
	jand g0848(.dina(w_n1110_1[1]),.dinb(w_n281_56[1]),.dout(n1111),.clk(gclk));
	jor g0849(.dina(w_n504_0[0]),.dinb(w_n273_34[2]),.dout(n1112),.clk(gclk));
	jor g0850(.dina(w_n518_0[0]),.dinb(w_shift1_34[2]),.dout(n1113),.clk(gclk));
	jand g0851(.dina(n1113),.dinb(n1112),.dout(n1114),.clk(gclk));
	jand g0852(.dina(w_n1114_1[1]),.dinb(w_n292_56[1]),.dout(n1115),.clk(gclk));
	jor g0853(.dina(n1115),.dinb(n1111),.dout(n1116),.clk(gclk));
	jor g0854(.dina(w_n524_0[0]),.dinb(w_n273_34[1]),.dout(n1117),.clk(gclk));
	jor g0855(.dina(w_n539_0[0]),.dinb(w_shift1_34[1]),.dout(n1118),.clk(gclk));
	jand g0856(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jand g0857(.dina(w_n1119_1[1]),.dinb(w_n267_56[1]),.dout(n1120),.clk(gclk));
	jor g0858(.dina(w_dff_B_YCE8fMWj4_0),.dinb(n1116),.dout(n1121),.clk(gclk));
	jor g0859(.dina(n1121),.dinb(w_dff_B_CJe3LNGD1_1),.dout(n1122),.clk(gclk));
	jand g0860(.dina(w_n1122_1[1]),.dinb(w_n319_61[2]),.dout(n1123),.clk(gclk));
	jor g0861(.dina(w_n624_0[0]),.dinb(w_n273_34[0]),.dout(n1124),.clk(gclk));
	jor g0862(.dina(w_n437_0[0]),.dinb(w_shift1_34[0]),.dout(n1125),.clk(gclk));
	jand g0863(.dina(n1125),.dinb(n1124),.dout(n1126),.clk(gclk));
	jand g0864(.dina(w_n1126_1[1]),.dinb(w_n304_56[0]),.dout(n1127),.clk(gclk));
	jor g0865(.dina(w_n603_0[0]),.dinb(w_n273_33[2]),.dout(n1128),.clk(gclk));
	jor g0866(.dina(w_n597_0[0]),.dinb(w_shift1_33[2]),.dout(n1129),.clk(gclk));
	jand g0867(.dina(n1129),.dinb(n1128),.dout(n1130),.clk(gclk));
	jand g0868(.dina(w_n1130_1[1]),.dinb(w_n281_56[0]),.dout(n1131),.clk(gclk));
	jor g0869(.dina(w_n593_0[0]),.dinb(w_n273_33[1]),.dout(n1132),.clk(gclk));
	jor g0870(.dina(w_n628_0[0]),.dinb(w_shift1_33[1]),.dout(n1133),.clk(gclk));
	jand g0871(.dina(n1133),.dinb(n1132),.dout(n1134),.clk(gclk));
	jand g0872(.dina(w_n1134_1[1]),.dinb(w_n267_56[0]),.dout(n1135),.clk(gclk));
	jor g0873(.dina(n1135),.dinb(n1131),.dout(n1136),.clk(gclk));
	jor g0874(.dina(w_n613_0[0]),.dinb(w_n273_33[0]),.dout(n1137),.clk(gclk));
	jor g0875(.dina(w_n607_0[0]),.dinb(w_shift1_33[0]),.dout(n1138),.clk(gclk));
	jand g0876(.dina(n1138),.dinb(n1137),.dout(n1139),.clk(gclk));
	jand g0877(.dina(w_n1139_1[1]),.dinb(w_n292_56[0]),.dout(n1140),.clk(gclk));
	jor g0878(.dina(w_dff_B_5ldzfQYi3_0),.dinb(n1136),.dout(n1141),.clk(gclk));
	jor g0879(.dina(n1141),.dinb(w_dff_B_gws8z3LA1_1),.dout(n1142),.clk(gclk));
	jand g0880(.dina(w_n1142_1[1]),.dinb(w_n364_61[2]),.dout(n1143),.clk(gclk));
	jor g0881(.dina(n1143),.dinb(n1123),.dout(n1144),.clk(gclk));
	jor g0882(.dina(w_n568_0[0]),.dinb(w_n273_32[2]),.dout(n1145),.clk(gclk));
	jor g0883(.dina(w_n562_0[0]),.dinb(w_shift1_32[2]),.dout(n1146),.clk(gclk));
	jand g0884(.dina(n1146),.dinb(n1145),.dout(n1147),.clk(gclk));
	jand g0885(.dina(w_n1147_1[1]),.dinb(w_n292_55[2]),.dout(n1148),.clk(gclk));
	jor g0886(.dina(w_n558_0[0]),.dinb(w_n273_32[1]),.dout(n1149),.clk(gclk));
	jor g0887(.dina(w_n552_0[0]),.dinb(w_shift1_32[1]),.dout(n1150),.clk(gclk));
	jand g0888(.dina(n1150),.dinb(n1149),.dout(n1151),.clk(gclk));
	jand g0889(.dina(w_n1151_1[1]),.dinb(w_n281_55[2]),.dout(n1152),.clk(gclk));
	jor g0890(.dina(w_n548_0[0]),.dinb(w_n273_32[0]),.dout(n1153),.clk(gclk));
	jor g0891(.dina(w_n583_0[0]),.dinb(w_shift1_32[0]),.dout(n1154),.clk(gclk));
	jand g0892(.dina(n1154),.dinb(n1153),.dout(n1155),.clk(gclk));
	jand g0893(.dina(w_n1155_1[1]),.dinb(w_n267_55[2]),.dout(n1156),.clk(gclk));
	jor g0894(.dina(n1156),.dinb(n1152),.dout(n1157),.clk(gclk));
	jor g0895(.dina(w_n579_0[0]),.dinb(w_n273_31[2]),.dout(n1158),.clk(gclk));
	jor g0896(.dina(w_n508_0[0]),.dinb(w_shift1_31[2]),.dout(n1159),.clk(gclk));
	jand g0897(.dina(n1159),.dinb(n1158),.dout(n1160),.clk(gclk));
	jand g0898(.dina(w_n1160_1[1]),.dinb(w_n304_55[2]),.dout(n1161),.clk(gclk));
	jor g0899(.dina(w_dff_B_aeg3cgRf4_0),.dinb(n1157),.dout(n1162),.clk(gclk));
	jor g0900(.dina(n1162),.dinb(w_dff_B_sQ1XAWmU2_1),.dout(n1163),.clk(gclk));
	jand g0901(.dina(w_n1163_1[1]),.dinb(w_n265_61[2]),.dout(n1164),.clk(gclk));
	jor g0902(.dina(w_dff_B_U2b0FtDF4_0),.dinb(n1144),.dout(n1165),.clk(gclk));
	jor g0903(.dina(n1165),.dinb(w_dff_B_wVw0jevq6_1),.dout(n1166),.clk(gclk));
	jor g0904(.dina(w_n1166_0[1]),.dinb(w_shift6_62[2]),.dout(n1167),.clk(gclk));
	jand g0905(.dina(n1167),.dinb(n1083),.dout(result2),.clk(gclk));
	jand g0906(.dina(w_n661_0[0]),.dinb(w_shift1_31[1]),.dout(n1169),.clk(gclk));
	jand g0907(.dina(w_n655_0[0]),.dinb(w_n273_31[1]),.dout(n1170),.clk(gclk));
	jor g0908(.dina(n1170),.dinb(n1169),.dout(n1171),.clk(gclk));
	jand g0909(.dina(w_n1171_1[1]),.dinb(w_n292_55[1]),.dout(n1172),.clk(gclk));
	jand g0910(.dina(w_n651_0[0]),.dinb(w_shift1_31[0]),.dout(n1173),.clk(gclk));
	jand g0911(.dina(w_n645_0[0]),.dinb(w_n273_31[0]),.dout(n1174),.clk(gclk));
	jor g0912(.dina(n1174),.dinb(n1173),.dout(n1175),.clk(gclk));
	jand g0913(.dina(w_n1175_1[1]),.dinb(w_n281_55[1]),.dout(n1176),.clk(gclk));
	jand g0914(.dina(w_n641_0[0]),.dinb(w_shift1_30[2]),.dout(n1177),.clk(gclk));
	jand g0915(.dina(w_n676_0[0]),.dinb(w_n273_30[2]),.dout(n1178),.clk(gclk));
	jor g0916(.dina(n1178),.dinb(n1177),.dout(n1179),.clk(gclk));
	jand g0917(.dina(w_n1179_1[1]),.dinb(w_n267_55[1]),.dout(n1180),.clk(gclk));
	jor g0918(.dina(n1180),.dinb(n1176),.dout(n1181),.clk(gclk));
	jand g0919(.dina(w_n672_0[0]),.dinb(w_shift1_30[1]),.dout(n1182),.clk(gclk));
	jand g0920(.dina(w_n825_0[0]),.dinb(w_n273_30[1]),.dout(n1183),.clk(gclk));
	jor g0921(.dina(n1183),.dinb(n1182),.dout(n1184),.clk(gclk));
	jand g0922(.dina(w_n1184_1[1]),.dinb(w_n304_55[1]),.dout(n1185),.clk(gclk));
	jor g0923(.dina(w_dff_B_NyFPXIyr2_0),.dinb(n1181),.dout(n1186),.clk(gclk));
	jor g0924(.dina(n1186),.dinb(w_dff_B_L4laJNFt4_1),.dout(n1187),.clk(gclk));
	jand g0925(.dina(w_n1187_1[1]),.dinb(w_n364_61[1]),.dout(n1188),.clk(gclk));
	jand g0926(.dina(w_n716_0[0]),.dinb(w_shift1_30[0]),.dout(n1189),.clk(gclk));
	jand g0927(.dina(w_n778_0[0]),.dinb(w_n273_30[0]),.dout(n1190),.clk(gclk));
	jor g0928(.dina(n1190),.dinb(n1189),.dout(n1191),.clk(gclk));
	jand g0929(.dina(w_n1191_1[1]),.dinb(w_n304_55[0]),.dout(n1192),.clk(gclk));
	jand g0930(.dina(w_n695_0[0]),.dinb(w_shift1_29[2]),.dout(n1193),.clk(gclk));
	jand g0931(.dina(w_n709_0[0]),.dinb(w_n273_29[2]),.dout(n1194),.clk(gclk));
	jor g0932(.dina(n1194),.dinb(n1193),.dout(n1195),.clk(gclk));
	jand g0933(.dina(w_n1195_1[1]),.dinb(w_n281_55[0]),.dout(n1196),.clk(gclk));
	jand g0934(.dina(w_n685_0[0]),.dinb(w_shift1_29[1]),.dout(n1197),.clk(gclk));
	jand g0935(.dina(w_n699_0[0]),.dinb(w_n273_29[1]),.dout(n1198),.clk(gclk));
	jor g0936(.dina(n1198),.dinb(n1197),.dout(n1199),.clk(gclk));
	jand g0937(.dina(w_n1199_1[1]),.dinb(w_n292_55[0]),.dout(n1200),.clk(gclk));
	jor g0938(.dina(n1200),.dinb(n1196),.dout(n1201),.clk(gclk));
	jand g0939(.dina(w_n705_0[0]),.dinb(w_shift1_29[0]),.dout(n1202),.clk(gclk));
	jand g0940(.dina(w_n720_0[0]),.dinb(w_n273_29[0]),.dout(n1203),.clk(gclk));
	jor g0941(.dina(n1203),.dinb(n1202),.dout(n1204),.clk(gclk));
	jand g0942(.dina(w_n1204_1[1]),.dinb(w_n267_55[0]),.dout(n1205),.clk(gclk));
	jor g0943(.dina(w_dff_B_t5k4kQhB6_0),.dinb(n1201),.dout(n1206),.clk(gclk));
	jor g0944(.dina(n1206),.dinb(w_dff_B_82FVcnT81_1),.dout(n1207),.clk(gclk));
	jand g0945(.dina(w_n1207_1[1]),.dinb(w_n265_61[1]),.dout(n1208),.clk(gclk));
	jand g0946(.dina(w_n729_0[0]),.dinb(w_shift1_28[2]),.dout(n1209),.clk(gclk));
	jand g0947(.dina(w_n689_0[0]),.dinb(w_n273_28[2]),.dout(n1210),.clk(gclk));
	jor g0948(.dina(n1210),.dinb(n1209),.dout(n1211),.clk(gclk));
	jand g0949(.dina(w_n1211_1[1]),.dinb(w_n304_54[2]),.dout(n1212),.clk(gclk));
	jand g0950(.dina(w_n739_0[0]),.dinb(w_shift1_28[1]),.dout(n1213),.clk(gclk));
	jand g0951(.dina(w_n764_0[0]),.dinb(w_n273_28[1]),.dout(n1214),.clk(gclk));
	jor g0952(.dina(n1214),.dinb(n1213),.dout(n1215),.clk(gclk));
	jand g0953(.dina(w_n1215_1[1]),.dinb(w_n281_54[2]),.dout(n1216),.clk(gclk));
	jand g0954(.dina(w_n760_0[0]),.dinb(w_shift1_28[0]),.dout(n1217),.clk(gclk));
	jand g0955(.dina(w_n733_0[0]),.dinb(w_n273_28[0]),.dout(n1218),.clk(gclk));
	jor g0956(.dina(n1218),.dinb(n1217),.dout(n1219),.clk(gclk));
	jand g0957(.dina(w_n1219_1[1]),.dinb(w_n267_54[2]),.dout(n1220),.clk(gclk));
	jor g0958(.dina(n1220),.dinb(n1216),.dout(n1221),.clk(gclk));
	jand g0959(.dina(w_n749_0[0]),.dinb(w_shift1_27[2]),.dout(n1222),.clk(gclk));
	jand g0960(.dina(w_n743_0[0]),.dinb(w_n273_27[2]),.dout(n1223),.clk(gclk));
	jor g0961(.dina(n1223),.dinb(n1222),.dout(n1224),.clk(gclk));
	jand g0962(.dina(w_n1224_1[1]),.dinb(w_n292_54[2]),.dout(n1225),.clk(gclk));
	jor g0963(.dina(w_dff_B_hZx5Rp366_0),.dinb(n1221),.dout(n1226),.clk(gclk));
	jor g0964(.dina(n1226),.dinb(w_dff_B_ycfnNlTi5_1),.dout(n1227),.clk(gclk));
	jand g0965(.dina(w_n1227_1[1]),.dinb(w_n410_61[1]),.dout(n1228),.clk(gclk));
	jor g0966(.dina(n1228),.dinb(n1208),.dout(n1229),.clk(gclk));
	jand g0967(.dina(w_n774_0[0]),.dinb(w_shift1_27[1]),.dout(n1230),.clk(gclk));
	jand g0968(.dina(w_n784_0[0]),.dinb(w_n273_27[1]),.dout(n1231),.clk(gclk));
	jor g0969(.dina(n1231),.dinb(n1230),.dout(n1232),.clk(gclk));
	jand g0970(.dina(w_n1232_1[1]),.dinb(w_n292_54[1]),.dout(n1233),.clk(gclk));
	jand g0971(.dina(w_n788_0[0]),.dinb(w_shift1_27[0]),.dout(n1234),.clk(gclk));
	jand g0972(.dina(w_n798_0[0]),.dinb(w_n273_27[0]),.dout(n1235),.clk(gclk));
	jor g0973(.dina(n1235),.dinb(n1234),.dout(n1236),.clk(gclk));
	jand g0974(.dina(w_n1236_1[1]),.dinb(w_n281_54[1]),.dout(n1237),.clk(gclk));
	jor g0975(.dina(w_n809_0[0]),.dinb(w_shift1_26[2]),.dout(n1238),.clk(gclk));
	jor g0976(.dina(w_n794_0[0]),.dinb(w_n273_26[2]),.dout(n1239),.clk(gclk));
	jand g0977(.dina(n1239),.dinb(n1238),.dout(n1240),.clk(gclk));
	jand g0978(.dina(w_n1240_1[1]),.dinb(w_n267_54[1]),.dout(n1241),.clk(gclk));
	jor g0979(.dina(n1241),.dinb(n1237),.dout(n1242),.clk(gclk));
	jand g0980(.dina(w_n805_0[0]),.dinb(w_shift1_26[1]),.dout(n1243),.clk(gclk));
	jand g0981(.dina(w_n665_0[0]),.dinb(w_n273_26[1]),.dout(n1244),.clk(gclk));
	jor g0982(.dina(n1244),.dinb(n1243),.dout(n1245),.clk(gclk));
	jand g0983(.dina(w_n1245_1[1]),.dinb(w_n304_54[1]),.dout(n1246),.clk(gclk));
	jor g0984(.dina(w_dff_B_Qp7R6Ppv0_0),.dinb(n1242),.dout(n1247),.clk(gclk));
	jor g0985(.dina(n1247),.dinb(w_dff_B_VGg8A4KJ8_1),.dout(n1248),.clk(gclk));
	jand g0986(.dina(w_n1248_1[1]),.dinb(w_n319_61[1]),.dout(n1249),.clk(gclk));
	jor g0987(.dina(w_dff_B_PVP23snq0_0),.dinb(n1229),.dout(n1250),.clk(gclk));
	jor g0988(.dina(n1250),.dinb(w_dff_B_x7FH33QW3_1),.dout(n1251),.clk(gclk));
	jor g0989(.dina(w_n1251_0[1]),.dinb(w_n263_62[1]),.dout(n1252),.clk(gclk));
	jand g0990(.dina(w_n896_0[0]),.dinb(w_shift1_26[0]),.dout(n1253),.clk(gclk));
	jand g0991(.dina(w_n978_0[0]),.dinb(w_n273_26[0]),.dout(n1254),.clk(gclk));
	jor g0992(.dina(n1254),.dinb(n1253),.dout(n1255),.clk(gclk));
	jand g0993(.dina(w_n1255_1[1]),.dinb(w_n304_54[0]),.dout(n1256),.clk(gclk));
	jand g0994(.dina(w_n875_0[0]),.dinb(w_shift1_25[2]),.dout(n1257),.clk(gclk));
	jand g0995(.dina(w_n889_0[0]),.dinb(w_n273_25[2]),.dout(n1258),.clk(gclk));
	jor g0996(.dina(n1258),.dinb(n1257),.dout(n1259),.clk(gclk));
	jand g0997(.dina(w_n1259_1[1]),.dinb(w_n281_54[0]),.dout(n1260),.clk(gclk));
	jand g0998(.dina(w_n885_0[0]),.dinb(w_shift1_25[1]),.dout(n1261),.clk(gclk));
	jand g0999(.dina(w_n900_0[0]),.dinb(w_n273_25[1]),.dout(n1262),.clk(gclk));
	jor g1000(.dina(n1262),.dinb(n1261),.dout(n1263),.clk(gclk));
	jand g1001(.dina(w_n1263_1[1]),.dinb(w_n267_54[0]),.dout(n1264),.clk(gclk));
	jor g1002(.dina(n1264),.dinb(n1260),.dout(n1265),.clk(gclk));
	jand g1003(.dina(w_n865_0[0]),.dinb(w_shift1_25[0]),.dout(n1266),.clk(gclk));
	jand g1004(.dina(w_n879_0[0]),.dinb(w_n273_25[0]),.dout(n1267),.clk(gclk));
	jor g1005(.dina(n1267),.dinb(n1266),.dout(n1268),.clk(gclk));
	jand g1006(.dina(w_n1268_1[1]),.dinb(w_n292_54[0]),.dout(n1269),.clk(gclk));
	jor g1007(.dina(w_dff_B_hGQAN2Ud3_0),.dinb(n1265),.dout(n1270),.clk(gclk));
	jor g1008(.dina(n1270),.dinb(w_dff_B_y7xezhI94_1),.dout(n1271),.clk(gclk));
	jand g1009(.dina(w_n1271_1[1]),.dinb(w_n319_61[0]),.dout(n1272),.clk(gclk));
	jand g1010(.dina(w_n852_0[0]),.dinb(w_shift1_24[2]),.dout(n1273),.clk(gclk));
	jand g1011(.dina(w_n913_0[0]),.dinb(w_n273_24[2]),.dout(n1274),.clk(gclk));
	jor g1012(.dina(n1274),.dinb(n1273),.dout(n1275),.clk(gclk));
	jand g1013(.dina(w_n1275_1[1]),.dinb(w_n304_53[2]),.dout(n1276),.clk(gclk));
	jand g1014(.dina(w_n831_0[0]),.dinb(w_shift1_24[1]),.dout(n1277),.clk(gclk));
	jand g1015(.dina(w_n845_0[0]),.dinb(w_n273_24[1]),.dout(n1278),.clk(gclk));
	jor g1016(.dina(n1278),.dinb(n1277),.dout(n1279),.clk(gclk));
	jand g1017(.dina(w_n1279_1[1]),.dinb(w_n281_53[2]),.dout(n1280),.clk(gclk));
	jand g1018(.dina(w_n841_0[0]),.dinb(w_shift1_24[0]),.dout(n1281),.clk(gclk));
	jand g1019(.dina(w_n856_0[0]),.dinb(w_n273_24[0]),.dout(n1282),.clk(gclk));
	jor g1020(.dina(n1282),.dinb(n1281),.dout(n1283),.clk(gclk));
	jand g1021(.dina(w_n1283_1[1]),.dinb(w_n267_53[2]),.dout(n1284),.clk(gclk));
	jor g1022(.dina(n1284),.dinb(n1280),.dout(n1285),.clk(gclk));
	jand g1023(.dina(w_n821_0[0]),.dinb(w_shift1_23[2]),.dout(n1286),.clk(gclk));
	jand g1024(.dina(w_n835_0[0]),.dinb(w_n273_23[2]),.dout(n1287),.clk(gclk));
	jor g1025(.dina(n1287),.dinb(n1286),.dout(n1288),.clk(gclk));
	jand g1026(.dina(w_n1288_1[1]),.dinb(w_n292_53[2]),.dout(n1289),.clk(gclk));
	jor g1027(.dina(w_dff_B_bxZjKYFc1_0),.dinb(n1285),.dout(n1290),.clk(gclk));
	jor g1028(.dina(n1290),.dinb(w_dff_B_v6S0pnWU5_1),.dout(n1291),.clk(gclk));
	jand g1029(.dina(w_n1291_1[1]),.dinb(w_n410_61[0]),.dout(n1292),.clk(gclk));
	jand g1030(.dina(w_n974_0[0]),.dinb(w_shift1_23[1]),.dout(n1293),.clk(gclk));
	jand g1031(.dina(w_n968_0[0]),.dinb(w_n273_23[1]),.dout(n1294),.clk(gclk));
	jor g1032(.dina(n1294),.dinb(n1293),.dout(n1295),.clk(gclk));
	jand g1033(.dina(w_n1295_1[1]),.dinb(w_n292_53[1]),.dout(n1296),.clk(gclk));
	jand g1034(.dina(w_n964_0[0]),.dinb(w_shift1_23[0]),.dout(n1297),.clk(gclk));
	jand g1035(.dina(w_n958_0[0]),.dinb(w_n273_23[0]),.dout(n1298),.clk(gclk));
	jor g1036(.dina(n1298),.dinb(n1297),.dout(n1299),.clk(gclk));
	jand g1037(.dina(w_n1299_1[1]),.dinb(w_n281_53[1]),.dout(n1300),.clk(gclk));
	jand g1038(.dina(w_n954_0[0]),.dinb(w_shift1_22[2]),.dout(n1301),.clk(gclk));
	jand g1039(.dina(w_n989_0[0]),.dinb(w_n273_22[2]),.dout(n1302),.clk(gclk));
	jor g1040(.dina(n1302),.dinb(n1301),.dout(n1303),.clk(gclk));
	jand g1041(.dina(w_n1303_1[1]),.dinb(w_n267_53[1]),.dout(n1304),.clk(gclk));
	jor g1042(.dina(n1304),.dinb(n1300),.dout(n1305),.clk(gclk));
	jand g1043(.dina(w_n985_0[0]),.dinb(w_shift1_22[1]),.dout(n1306),.clk(gclk));
	jand g1044(.dina(w_n753_0[0]),.dinb(w_n273_22[1]),.dout(n1307),.clk(gclk));
	jor g1045(.dina(n1307),.dinb(n1306),.dout(n1308),.clk(gclk));
	jand g1046(.dina(w_n1308_1[1]),.dinb(w_n304_53[1]),.dout(n1309),.clk(gclk));
	jor g1047(.dina(w_dff_B_B2NxBOMf3_0),.dinb(n1305),.dout(n1310),.clk(gclk));
	jor g1048(.dina(n1310),.dinb(w_dff_B_vvMFgqlf6_1),.dout(n1311),.clk(gclk));
	jand g1049(.dina(w_n1311_1[1]),.dinb(w_n364_61[0]),.dout(n1312),.clk(gclk));
	jor g1050(.dina(n1312),.dinb(n1292),.dout(n1313),.clk(gclk));
	jand g1051(.dina(w_n940_0[0]),.dinb(w_shift1_22[0]),.dout(n1314),.clk(gclk));
	jand g1052(.dina(w_n869_0[0]),.dinb(w_n273_22[0]),.dout(n1315),.clk(gclk));
	jor g1053(.dina(n1315),.dinb(n1314),.dout(n1316),.clk(gclk));
	jand g1054(.dina(w_n1316_1[1]),.dinb(w_n304_53[0]),.dout(n1317),.clk(gclk));
	jand g1055(.dina(w_n919_0[0]),.dinb(w_shift1_21[2]),.dout(n1318),.clk(gclk));
	jand g1056(.dina(w_n933_0[0]),.dinb(w_n273_21[2]),.dout(n1319),.clk(gclk));
	jor g1057(.dina(n1319),.dinb(n1318),.dout(n1320),.clk(gclk));
	jand g1058(.dina(w_n1320_1[1]),.dinb(w_n281_53[0]),.dout(n1321),.clk(gclk));
	jand g1059(.dina(w_n929_0[0]),.dinb(w_shift1_21[1]),.dout(n1322),.clk(gclk));
	jand g1060(.dina(w_n944_0[0]),.dinb(w_n273_21[1]),.dout(n1323),.clk(gclk));
	jor g1061(.dina(n1323),.dinb(n1322),.dout(n1324),.clk(gclk));
	jand g1062(.dina(w_n1324_1[1]),.dinb(w_n267_53[0]),.dout(n1325),.clk(gclk));
	jor g1063(.dina(n1325),.dinb(n1321),.dout(n1326),.clk(gclk));
	jand g1064(.dina(w_n909_0[0]),.dinb(w_shift1_21[0]),.dout(n1327),.clk(gclk));
	jand g1065(.dina(w_n923_0[0]),.dinb(w_n273_21[0]),.dout(n1328),.clk(gclk));
	jor g1066(.dina(n1328),.dinb(n1327),.dout(n1329),.clk(gclk));
	jand g1067(.dina(w_n1329_1[1]),.dinb(w_n292_53[0]),.dout(n1330),.clk(gclk));
	jor g1068(.dina(w_dff_B_xB4q2Qjw2_0),.dinb(n1326),.dout(n1331),.clk(gclk));
	jor g1069(.dina(n1331),.dinb(w_dff_B_6KHWH1Jh5_1),.dout(n1332),.clk(gclk));
	jand g1070(.dina(w_n1332_1[1]),.dinb(w_n265_61[0]),.dout(n1333),.clk(gclk));
	jor g1071(.dina(w_dff_B_5urLXsyC3_0),.dinb(n1313),.dout(n1334),.clk(gclk));
	jor g1072(.dina(n1334),.dinb(w_dff_B_e8li2tLE4_1),.dout(n1335),.clk(gclk));
	jor g1073(.dina(w_n1335_0[1]),.dinb(w_shift6_62[1]),.dout(n1336),.clk(gclk));
	jand g1074(.dina(n1336),.dinb(n1252),.dout(result3),.clk(gclk));
	jand g1075(.dina(w_n383_1[0]),.dinb(w_n292_52[2]),.dout(n1338),.clk(gclk));
	jand g1076(.dina(w_n393_1[0]),.dinb(w_n281_52[2]),.dout(n1339),.clk(gclk));
	jand g1077(.dina(w_n373_1[0]),.dinb(w_n267_52[2]),.dout(n1340),.clk(gclk));
	jor g1078(.dina(n1340),.dinb(n1339),.dout(n1341),.clk(gclk));
	jand g1079(.dina(w_n466_1[0]),.dinb(w_n304_52[2]),.dout(n1342),.clk(gclk));
	jor g1080(.dina(w_dff_B_1OEUfKzK8_0),.dinb(n1341),.dout(n1343),.clk(gclk));
	jor g1081(.dina(n1343),.dinb(w_dff_B_gfiTS28a2_1),.dout(n1344),.clk(gclk));
	jand g1082(.dina(w_n1344_1[1]),.dinb(w_n364_60[2]),.dout(n1345),.clk(gclk));
	jand g1083(.dina(w_n450_1[0]),.dinb(w_n267_52[1]),.dout(n1346),.clk(gclk));
	jand g1084(.dina(w_n419_1[0]),.dinb(w_n281_52[1]),.dout(n1347),.clk(gclk));
	jand g1085(.dina(w_n429_1[0]),.dinb(w_n292_52[1]),.dout(n1348),.clk(gclk));
	jor g1086(.dina(n1348),.dinb(n1347),.dout(n1349),.clk(gclk));
	jand g1087(.dina(w_n304_52[1]),.dinb(w_n301_1[0]),.dout(n1350),.clk(gclk));
	jor g1088(.dina(w_dff_B_PIEA6oQH3_0),.dinb(n1349),.dout(n1351),.clk(gclk));
	jor g1089(.dina(n1351),.dinb(w_dff_B_EMAK944C1_1),.dout(n1352),.clk(gclk));
	jand g1090(.dina(w_n1352_1[1]),.dinb(w_n410_60[2]),.dout(n1353),.clk(gclk));
	jand g1091(.dina(w_n328_1[0]),.dinb(w_n304_52[0]),.dout(n1354),.clk(gclk));
	jand g1092(.dina(w_n281_52[0]),.dinb(w_n278_1[0]),.dout(n1355),.clk(gclk));
	jand g1093(.dina(w_n292_52[0]),.dinb(w_n290_1[0]),.dout(n1356),.clk(gclk));
	jor g1094(.dina(n1356),.dinb(n1355),.dout(n1357),.clk(gclk));
	jand g1095(.dina(w_n313_1[0]),.dinb(w_n267_52[0]),.dout(n1358),.clk(gclk));
	jor g1096(.dina(w_dff_B_8BngNbgd0_0),.dinb(n1357),.dout(n1359),.clk(gclk));
	jor g1097(.dina(n1359),.dinb(w_dff_B_Y9K3ClDR7_1),.dout(n1360),.clk(gclk));
	jand g1098(.dina(w_n1360_1[1]),.dinb(w_n265_60[2]),.dout(n1361),.clk(gclk));
	jor g1099(.dina(n1361),.dinb(n1353),.dout(n1362),.clk(gclk));
	jand g1100(.dina(w_n359_1[0]),.dinb(w_n267_51[2]),.dout(n1363),.clk(gclk));
	jand g1101(.dina(w_n348_1[0]),.dinb(w_n281_51[2]),.dout(n1364),.clk(gclk));
	jand g1102(.dina(w_n338_1[0]),.dinb(w_n292_51[2]),.dout(n1365),.clk(gclk));
	jor g1103(.dina(n1365),.dinb(n1364),.dout(n1366),.clk(gclk));
	jand g1104(.dina(w_n404_1[0]),.dinb(w_n304_51[2]),.dout(n1367),.clk(gclk));
	jor g1105(.dina(w_dff_B_RWQCZSD81_0),.dinb(n1366),.dout(n1368),.clk(gclk));
	jor g1106(.dina(n1368),.dinb(w_dff_B_DD4YCshY8_1),.dout(n1369),.clk(gclk));
	jand g1107(.dina(w_n1369_1[1]),.dinb(w_n319_60[2]),.dout(n1370),.clk(gclk));
	jor g1108(.dina(w_dff_B_ckbM7ytb5_0),.dinb(n1362),.dout(n1371),.clk(gclk));
	jor g1109(.dina(n1371),.dinb(w_dff_B_yt8yq8iV8_1),.dout(n1372),.clk(gclk));
	jor g1110(.dina(w_n1372_0[1]),.dinb(w_n263_62[0]),.dout(n1373),.clk(gclk));
	jand g1111(.dina(w_n585_1[0]),.dinb(w_n267_51[1]),.dout(n1374),.clk(gclk));
	jand g1112(.dina(w_n554_1[0]),.dinb(w_n281_51[1]),.dout(n1375),.clk(gclk));
	jand g1113(.dina(w_n564_1[0]),.dinb(w_n292_51[1]),.dout(n1376),.clk(gclk));
	jor g1114(.dina(n1376),.dinb(n1375),.dout(n1377),.clk(gclk));
	jand g1115(.dina(w_n510_1[0]),.dinb(w_n304_51[1]),.dout(n1378),.clk(gclk));
	jor g1116(.dina(w_dff_B_Yji0C1js9_0),.dinb(n1377),.dout(n1379),.clk(gclk));
	jor g1117(.dina(n1379),.dinb(w_dff_B_EtA1Bwgh7_1),.dout(n1380),.clk(gclk));
	jand g1118(.dina(w_n1380_1[1]),.dinb(w_n265_60[1]),.dout(n1381),.clk(gclk));
	jand g1119(.dina(w_n619_1[0]),.dinb(w_n304_51[0]),.dout(n1382),.clk(gclk));
	jand g1120(.dina(w_n530_1[0]),.dinb(w_n281_51[0]),.dout(n1383),.clk(gclk));
	jand g1121(.dina(w_n541_1[0]),.dinb(w_n267_51[0]),.dout(n1384),.clk(gclk));
	jor g1122(.dina(n1384),.dinb(n1383),.dout(n1385),.clk(gclk));
	jand g1123(.dina(w_n520_1[0]),.dinb(w_n292_51[0]),.dout(n1386),.clk(gclk));
	jor g1124(.dina(w_dff_B_hknLRKEp8_0),.dinb(n1385),.dout(n1387),.clk(gclk));
	jor g1125(.dina(n1387),.dinb(w_dff_B_StgGyzNM1_1),.dout(n1388),.clk(gclk));
	jand g1126(.dina(w_n1388_1[1]),.dinb(w_n319_60[1]),.dout(n1389),.clk(gclk));
	jand g1127(.dina(w_n439_1[0]),.dinb(w_n304_50[2]),.dout(n1390),.clk(gclk));
	jand g1128(.dina(w_n599_1[0]),.dinb(w_n281_50[2]),.dout(n1391),.clk(gclk));
	jand g1129(.dina(w_n609_1[0]),.dinb(w_n292_50[2]),.dout(n1392),.clk(gclk));
	jor g1130(.dina(n1392),.dinb(n1391),.dout(n1393),.clk(gclk));
	jand g1131(.dina(w_n630_1[0]),.dinb(w_n267_50[2]),.dout(n1394),.clk(gclk));
	jor g1132(.dina(w_dff_B_70rd1kZT3_0),.dinb(n1393),.dout(n1395),.clk(gclk));
	jor g1133(.dina(n1395),.dinb(w_dff_B_wO6CPyKc2_1),.dout(n1396),.clk(gclk));
	jand g1134(.dina(w_n1396_1[1]),.dinb(w_n364_60[1]),.dout(n1397),.clk(gclk));
	jor g1135(.dina(n1397),.dinb(n1389),.dout(n1398),.clk(gclk));
	jand g1136(.dina(w_n574_1[0]),.dinb(w_n304_50[1]),.dout(n1399),.clk(gclk));
	jand g1137(.dina(w_n486_1[0]),.dinb(w_n281_50[1]),.dout(n1400),.clk(gclk));
	jand g1138(.dina(w_n497_1[0]),.dinb(w_n267_50[1]),.dout(n1401),.clk(gclk));
	jor g1139(.dina(n1401),.dinb(n1400),.dout(n1402),.clk(gclk));
	jand g1140(.dina(w_n476_1[0]),.dinb(w_n292_50[1]),.dout(n1403),.clk(gclk));
	jor g1141(.dina(w_dff_B_1DoTDJze9_0),.dinb(n1402),.dout(n1404),.clk(gclk));
	jor g1142(.dina(n1404),.dinb(w_dff_B_bz9R4FL06_1),.dout(n1405),.clk(gclk));
	jand g1143(.dina(w_n1405_1[1]),.dinb(w_n410_60[1]),.dout(n1406),.clk(gclk));
	jor g1144(.dina(w_dff_B_lMbt7F9W4_0),.dinb(n1398),.dout(n1407),.clk(gclk));
	jor g1145(.dina(n1407),.dinb(w_dff_B_4hGgm3Et5_1),.dout(n1408),.clk(gclk));
	jor g1146(.dina(w_n1408_0[1]),.dinb(w_shift6_62[0]),.dout(n1409),.clk(gclk));
	jand g1147(.dina(n1409),.dinb(n1373),.dout(result4),.clk(gclk));
	jand g1148(.dina(w_n667_1[0]),.dinb(w_n304_50[0]),.dout(n1411),.clk(gclk));
	jand g1149(.dina(w_n800_1[0]),.dinb(w_n281_50[0]),.dout(n1412),.clk(gclk));
	jand g1150(.dina(w_n790_1[0]),.dinb(w_n292_50[0]),.dout(n1413),.clk(gclk));
	jor g1151(.dina(n1413),.dinb(n1412),.dout(n1414),.clk(gclk));
	jand g1152(.dina(w_n811_1[0]),.dinb(w_n267_50[0]),.dout(n1415),.clk(gclk));
	jor g1153(.dina(w_dff_B_4FGpBViq2_0),.dinb(n1414),.dout(n1416),.clk(gclk));
	jor g1154(.dina(n1416),.dinb(w_dff_B_V651QdOo9_1),.dout(n1417),.clk(gclk));
	jand g1155(.dina(w_n1417_1[1]),.dinb(w_n319_60[0]),.dout(n1418),.clk(gclk));
	jand g1156(.dina(w_n745_1[0]),.dinb(w_n292_49[2]),.dout(n1419),.clk(gclk));
	jand g1157(.dina(w_n766_1[0]),.dinb(w_n281_49[2]),.dout(n1420),.clk(gclk));
	jand g1158(.dina(w_n735_1[0]),.dinb(w_n267_49[2]),.dout(n1421),.clk(gclk));
	jor g1159(.dina(n1421),.dinb(n1420),.dout(n1422),.clk(gclk));
	jand g1160(.dina(w_n691_1[0]),.dinb(w_n304_49[2]),.dout(n1423),.clk(gclk));
	jor g1161(.dina(w_dff_B_FQAQqQ3K2_0),.dinb(n1422),.dout(n1424),.clk(gclk));
	jor g1162(.dina(n1424),.dinb(w_dff_B_hozR8B1v3_1),.dout(n1425),.clk(gclk));
	jand g1163(.dina(w_n1425_1[1]),.dinb(w_n410_60[0]),.dout(n1426),.clk(gclk));
	jand g1164(.dina(w_n701_1[0]),.dinb(w_n292_49[1]),.dout(n1427),.clk(gclk));
	jand g1165(.dina(w_n711_1[0]),.dinb(w_n281_49[1]),.dout(n1428),.clk(gclk));
	jand g1166(.dina(w_n722_1[0]),.dinb(w_n267_49[1]),.dout(n1429),.clk(gclk));
	jor g1167(.dina(n1429),.dinb(n1428),.dout(n1430),.clk(gclk));
	jand g1168(.dina(w_n780_1[0]),.dinb(w_n304_49[1]),.dout(n1431),.clk(gclk));
	jor g1169(.dina(w_dff_B_DqhQ5BMC9_0),.dinb(n1430),.dout(n1432),.clk(gclk));
	jor g1170(.dina(n1432),.dinb(w_dff_B_yogMl37H5_1),.dout(n1433),.clk(gclk));
	jand g1171(.dina(w_n1433_1[1]),.dinb(w_n265_60[0]),.dout(n1434),.clk(gclk));
	jor g1172(.dina(n1434),.dinb(n1426),.dout(n1435),.clk(gclk));
	jand g1173(.dina(w_n827_1[0]),.dinb(w_n304_49[0]),.dout(n1436),.clk(gclk));
	jand g1174(.dina(w_n647_1[0]),.dinb(w_n281_49[0]),.dout(n1437),.clk(gclk));
	jand g1175(.dina(w_n678_1[0]),.dinb(w_n267_49[0]),.dout(n1438),.clk(gclk));
	jor g1176(.dina(n1438),.dinb(n1437),.dout(n1439),.clk(gclk));
	jand g1177(.dina(w_n657_1[0]),.dinb(w_n292_49[0]),.dout(n1440),.clk(gclk));
	jor g1178(.dina(w_dff_B_iymvmlfM2_0),.dinb(n1439),.dout(n1441),.clk(gclk));
	jor g1179(.dina(n1441),.dinb(w_dff_B_KrkdkH7l9_1),.dout(n1442),.clk(gclk));
	jand g1180(.dina(w_n1442_1[1]),.dinb(w_n364_60[0]),.dout(n1443),.clk(gclk));
	jor g1181(.dina(w_dff_B_qygv1SxQ7_0),.dinb(n1435),.dout(n1444),.clk(gclk));
	jor g1182(.dina(n1444),.dinb(w_dff_B_koWa50FX4_1),.dout(n1445),.clk(gclk));
	jor g1183(.dina(w_n1445_0[1]),.dinb(w_n263_61[2]),.dout(n1446),.clk(gclk));
	jand g1184(.dina(w_n837_1[0]),.dinb(w_n292_48[2]),.dout(n1447),.clk(gclk));
	jand g1185(.dina(w_n847_1[0]),.dinb(w_n281_48[2]),.dout(n1448),.clk(gclk));
	jand g1186(.dina(w_n858_1[0]),.dinb(w_n267_48[2]),.dout(n1449),.clk(gclk));
	jor g1187(.dina(n1449),.dinb(n1448),.dout(n1450),.clk(gclk));
	jand g1188(.dina(w_n915_1[0]),.dinb(w_n304_48[2]),.dout(n1451),.clk(gclk));
	jor g1189(.dina(w_dff_B_D9fLjXBM7_0),.dinb(n1450),.dout(n1452),.clk(gclk));
	jor g1190(.dina(n1452),.dinb(w_dff_B_QwBaURrl5_1),.dout(n1453),.clk(gclk));
	jand g1191(.dina(w_n1453_1[1]),.dinb(w_n410_59[2]),.dout(n1454),.clk(gclk));
	jand g1192(.dina(w_n980_1[0]),.dinb(w_n304_48[1]),.dout(n1455),.clk(gclk));
	jand g1193(.dina(w_n891_1[0]),.dinb(w_n281_48[1]),.dout(n1456),.clk(gclk));
	jand g1194(.dina(w_n881_1[0]),.dinb(w_n292_48[1]),.dout(n1457),.clk(gclk));
	jor g1195(.dina(n1457),.dinb(n1456),.dout(n1458),.clk(gclk));
	jand g1196(.dina(w_n902_1[0]),.dinb(w_n267_48[1]),.dout(n1459),.clk(gclk));
	jor g1197(.dina(w_dff_B_LuB7p5DQ9_0),.dinb(n1458),.dout(n1460),.clk(gclk));
	jor g1198(.dina(n1460),.dinb(w_dff_B_O9cfa67M4_1),.dout(n1461),.clk(gclk));
	jand g1199(.dina(w_n1461_1[1]),.dinb(w_n319_59[2]),.dout(n1462),.clk(gclk));
	jand g1200(.dina(w_n871_1[0]),.dinb(w_n304_48[0]),.dout(n1463),.clk(gclk));
	jand g1201(.dina(w_n935_1[0]),.dinb(w_n281_48[0]),.dout(n1464),.clk(gclk));
	jand g1202(.dina(w_n925_1[0]),.dinb(w_n292_48[0]),.dout(n1465),.clk(gclk));
	jor g1203(.dina(n1465),.dinb(n1464),.dout(n1466),.clk(gclk));
	jand g1204(.dina(w_n946_1[0]),.dinb(w_n267_48[0]),.dout(n1467),.clk(gclk));
	jor g1205(.dina(w_dff_B_z89m836x9_0),.dinb(n1466),.dout(n1468),.clk(gclk));
	jor g1206(.dina(n1468),.dinb(w_dff_B_ObVd5VZ58_1),.dout(n1469),.clk(gclk));
	jand g1207(.dina(w_n1469_1[1]),.dinb(w_n265_59[2]),.dout(n1470),.clk(gclk));
	jor g1208(.dina(n1470),.dinb(n1462),.dout(n1471),.clk(gclk));
	jand g1209(.dina(w_n755_1[0]),.dinb(w_n304_47[2]),.dout(n1472),.clk(gclk));
	jand g1210(.dina(w_n960_1[0]),.dinb(w_n281_47[2]),.dout(n1473),.clk(gclk));
	jand g1211(.dina(w_n970_1[0]),.dinb(w_n292_47[2]),.dout(n1474),.clk(gclk));
	jor g1212(.dina(n1474),.dinb(n1473),.dout(n1475),.clk(gclk));
	jand g1213(.dina(w_n991_1[0]),.dinb(w_n267_47[2]),.dout(n1476),.clk(gclk));
	jor g1214(.dina(w_dff_B_RAvhSOHM5_0),.dinb(n1475),.dout(n1477),.clk(gclk));
	jor g1215(.dina(n1477),.dinb(w_dff_B_XnPkPJHe3_1),.dout(n1478),.clk(gclk));
	jand g1216(.dina(w_n1478_1[1]),.dinb(w_n364_59[2]),.dout(n1479),.clk(gclk));
	jor g1217(.dina(w_dff_B_i5x16gKI7_0),.dinb(n1471),.dout(n1480),.clk(gclk));
	jor g1218(.dina(n1480),.dinb(w_dff_B_emjTCb4j0_1),.dout(n1481),.clk(gclk));
	jor g1219(.dina(w_n1481_0[1]),.dinb(w_shift6_61[2]),.dout(n1482),.clk(gclk));
	jand g1220(.dina(n1482),.dinb(n1446),.dout(result5),.clk(gclk));
	jand g1221(.dina(w_n1010_1[0]),.dinb(w_n304_47[1]),.dout(n1484),.clk(gclk));
	jand g1222(.dina(w_n1030_1[0]),.dinb(w_n281_47[1]),.dout(n1485),.clk(gclk));
	jand g1223(.dina(w_n1026_1[0]),.dinb(w_n292_47[1]),.dout(n1486),.clk(gclk));
	jor g1224(.dina(n1486),.dinb(n1485),.dout(n1487),.clk(gclk));
	jand g1225(.dina(w_n1035_1[0]),.dinb(w_n267_47[1]),.dout(n1488),.clk(gclk));
	jor g1226(.dina(w_dff_B_JNJO4QOP3_0),.dinb(n1487),.dout(n1489),.clk(gclk));
	jor g1227(.dina(n1489),.dinb(w_dff_B_CBcSyyyU8_1),.dout(n1490),.clk(gclk));
	jand g1228(.dina(w_n1490_1[1]),.dinb(w_n265_59[1]),.dout(n1491),.clk(gclk));
	jand g1229(.dina(w_n1042_1[0]),.dinb(w_n267_47[0]),.dout(n1492),.clk(gclk));
	jand g1230(.dina(w_n1050_1[0]),.dinb(w_n281_47[0]),.dout(n1493),.clk(gclk));
	jand g1231(.dina(w_n1046_1[0]),.dinb(w_n292_47[0]),.dout(n1494),.clk(gclk));
	jor g1232(.dina(n1494),.dinb(n1493),.dout(n1495),.clk(gclk));
	jand g1233(.dina(w_n1022_1[0]),.dinb(w_n304_47[0]),.dout(n1496),.clk(gclk));
	jor g1234(.dina(w_dff_B_yYHiuxfW3_0),.dinb(n1495),.dout(n1497),.clk(gclk));
	jor g1235(.dina(n1497),.dinb(w_dff_B_JL4G19Qr8_1),.dout(n1498),.clk(gclk));
	jand g1236(.dina(w_n1498_1[1]),.dinb(w_n410_59[1]),.dout(n1499),.clk(gclk));
	jand g1237(.dina(w_n1076_1[0]),.dinb(w_n267_46[2]),.dout(n1500),.clk(gclk));
	jand g1238(.dina(w_n1071_1[0]),.dinb(w_n281_46[2]),.dout(n1501),.clk(gclk));
	jand g1239(.dina(w_n1067_1[0]),.dinb(w_n292_46[2]),.dout(n1502),.clk(gclk));
	jor g1240(.dina(n1502),.dinb(n1501),.dout(n1503),.clk(gclk));
	jand g1241(.dina(w_n1094_1[0]),.dinb(w_n304_46[2]),.dout(n1504),.clk(gclk));
	jor g1242(.dina(w_dff_B_ldonzCFe9_0),.dinb(n1503),.dout(n1505),.clk(gclk));
	jor g1243(.dina(n1505),.dinb(w_dff_B_FMefJS5z4_1),.dout(n1506),.clk(gclk));
	jand g1244(.dina(w_n1506_1[1]),.dinb(w_n364_59[1]),.dout(n1507),.clk(gclk));
	jor g1245(.dina(n1507),.dinb(n1499),.dout(n1508),.clk(gclk));
	jand g1246(.dina(w_n1063_1[0]),.dinb(w_n304_46[1]),.dout(n1509),.clk(gclk));
	jand g1247(.dina(w_n1002_1[0]),.dinb(w_n281_46[1]),.dout(n1510),.clk(gclk));
	jand g1248(.dina(w_n1015_1[0]),.dinb(w_n267_46[1]),.dout(n1511),.clk(gclk));
	jor g1249(.dina(n1511),.dinb(n1510),.dout(n1512),.clk(gclk));
	jand g1250(.dina(w_n1006_1[0]),.dinb(w_n292_46[1]),.dout(n1513),.clk(gclk));
	jor g1251(.dina(w_dff_B_KwAJ2y101_0),.dinb(n1512),.dout(n1514),.clk(gclk));
	jor g1252(.dina(n1514),.dinb(w_dff_B_QeKRpaxT3_1),.dout(n1515),.clk(gclk));
	jand g1253(.dina(w_n1515_1[1]),.dinb(w_n319_59[1]),.dout(n1516),.clk(gclk));
	jor g1254(.dina(w_dff_B_F4EsfGDJ5_0),.dinb(n1508),.dout(n1517),.clk(gclk));
	jor g1255(.dina(n1517),.dinb(w_dff_B_1dMdFzNe2_1),.dout(n1518),.clk(gclk));
	jor g1256(.dina(w_n1518_0[1]),.dinb(w_n263_61[1]),.dout(n1519),.clk(gclk));
	jand g1257(.dina(w_n1147_1[0]),.dinb(w_n304_46[0]),.dout(n1520),.clk(gclk));
	jand g1258(.dina(w_n1086_1[0]),.dinb(w_n281_46[0]),.dout(n1521),.clk(gclk));
	jand g1259(.dina(w_n1099_1[0]),.dinb(w_n267_46[0]),.dout(n1522),.clk(gclk));
	jor g1260(.dina(n1522),.dinb(n1521),.dout(n1523),.clk(gclk));
	jand g1261(.dina(w_n1090_1[0]),.dinb(w_n292_46[0]),.dout(n1524),.clk(gclk));
	jor g1262(.dina(w_dff_B_HuZqe8R86_0),.dinb(n1523),.dout(n1525),.clk(gclk));
	jor g1263(.dina(n1525),.dinb(w_dff_B_HZGcZQx65_1),.dout(n1526),.clk(gclk));
	jand g1264(.dina(w_n1526_1[1]),.dinb(w_n410_59[0]),.dout(n1527),.clk(gclk));
	jand g1265(.dina(w_n1106_1[0]),.dinb(w_n267_45[2]),.dout(n1528),.clk(gclk));
	jand g1266(.dina(w_n1119_1[0]),.dinb(w_n281_45[2]),.dout(n1529),.clk(gclk));
	jand g1267(.dina(w_n1110_1[0]),.dinb(w_n292_45[2]),.dout(n1530),.clk(gclk));
	jor g1268(.dina(n1530),.dinb(n1529),.dout(n1531),.clk(gclk));
	jand g1269(.dina(w_n1139_1[0]),.dinb(w_n304_45[2]),.dout(n1532),.clk(gclk));
	jor g1270(.dina(w_dff_B_FHH2yJSp7_0),.dinb(n1531),.dout(n1533),.clk(gclk));
	jor g1271(.dina(n1533),.dinb(w_dff_B_Y88xVshG7_1),.dout(n1534),.clk(gclk));
	jand g1272(.dina(w_n1534_1[1]),.dinb(w_n319_59[0]),.dout(n1535),.clk(gclk));
	jand g1273(.dina(w_n1055_1[0]),.dinb(w_n304_45[1]),.dout(n1536),.clk(gclk));
	jand g1274(.dina(w_n1134_1[0]),.dinb(w_n281_45[1]),.dout(n1537),.clk(gclk));
	jand g1275(.dina(w_n1126_1[0]),.dinb(w_n267_45[1]),.dout(n1538),.clk(gclk));
	jor g1276(.dina(n1538),.dinb(n1537),.dout(n1539),.clk(gclk));
	jand g1277(.dina(w_n1130_1[0]),.dinb(w_n292_45[1]),.dout(n1540),.clk(gclk));
	jor g1278(.dina(w_dff_B_7JX91FRK1_0),.dinb(n1539),.dout(n1541),.clk(gclk));
	jor g1279(.dina(n1541),.dinb(w_dff_B_qYzkE5Ne5_1),.dout(n1542),.clk(gclk));
	jand g1280(.dina(w_n1542_1[1]),.dinb(w_n364_59[0]),.dout(n1543),.clk(gclk));
	jor g1281(.dina(n1543),.dinb(n1535),.dout(n1544),.clk(gclk));
	jand g1282(.dina(w_n1151_1[0]),.dinb(w_n292_45[0]),.dout(n1545),.clk(gclk));
	jand g1283(.dina(w_n1155_1[0]),.dinb(w_n281_45[0]),.dout(n1546),.clk(gclk));
	jand g1284(.dina(w_n1160_1[0]),.dinb(w_n267_45[0]),.dout(n1547),.clk(gclk));
	jor g1285(.dina(n1547),.dinb(n1546),.dout(n1548),.clk(gclk));
	jand g1286(.dina(w_n1114_1[0]),.dinb(w_n304_45[0]),.dout(n1549),.clk(gclk));
	jor g1287(.dina(w_dff_B_XQRJK8hI2_0),.dinb(n1548),.dout(n1550),.clk(gclk));
	jor g1288(.dina(n1550),.dinb(w_dff_B_LnFLsAV69_1),.dout(n1551),.clk(gclk));
	jand g1289(.dina(w_n1551_1[1]),.dinb(w_n265_59[0]),.dout(n1552),.clk(gclk));
	jor g1290(.dina(w_dff_B_c0oDU8DR9_0),.dinb(n1544),.dout(n1553),.clk(gclk));
	jor g1291(.dina(n1553),.dinb(w_dff_B_MXNCDc511_1),.dout(n1554),.clk(gclk));
	jor g1292(.dina(w_n1554_0[1]),.dinb(w_shift6_61[1]),.dout(n1555),.clk(gclk));
	jand g1293(.dina(n1555),.dinb(n1519),.dout(result6),.clk(gclk));
	jand g1294(.dina(w_n1191_1[0]),.dinb(w_n267_44[2]),.dout(n1557),.clk(gclk));
	jand g1295(.dina(w_n1204_1[0]),.dinb(w_n281_44[2]),.dout(n1558),.clk(gclk));
	jand g1296(.dina(w_n1195_1[0]),.dinb(w_n292_44[2]),.dout(n1559),.clk(gclk));
	jor g1297(.dina(n1559),.dinb(n1558),.dout(n1560),.clk(gclk));
	jand g1298(.dina(w_n1232_1[0]),.dinb(w_n304_44[2]),.dout(n1561),.clk(gclk));
	jor g1299(.dina(w_dff_B_jew2rhCp7_0),.dinb(n1560),.dout(n1562),.clk(gclk));
	jor g1300(.dina(n1562),.dinb(w_dff_B_ZxgD49R90_1),.dout(n1563),.clk(gclk));
	jand g1301(.dina(w_n1563_1[1]),.dinb(w_n265_58[2]),.dout(n1564),.clk(gclk));
	jand g1302(.dina(w_n1199_1[0]),.dinb(w_n304_44[1]),.dout(n1565),.clk(gclk));
	jand g1303(.dina(w_n1219_1[0]),.dinb(w_n281_44[1]),.dout(n1566),.clk(gclk));
	jand g1304(.dina(w_n1211_1[0]),.dinb(w_n267_44[1]),.dout(n1567),.clk(gclk));
	jor g1305(.dina(n1567),.dinb(n1566),.dout(n1568),.clk(gclk));
	jand g1306(.dina(w_n1215_1[0]),.dinb(w_n292_44[1]),.dout(n1569),.clk(gclk));
	jor g1307(.dina(w_dff_B_K6ULNMp38_0),.dinb(n1568),.dout(n1570),.clk(gclk));
	jor g1308(.dina(n1570),.dinb(w_dff_B_qvZOCGkh7_1),.dout(n1571),.clk(gclk));
	jand g1309(.dina(w_n1571_1[1]),.dinb(w_n410_58[2]),.dout(n1572),.clk(gclk));
	jand g1310(.dina(w_n1184_1[0]),.dinb(w_n267_44[0]),.dout(n1573),.clk(gclk));
	jand g1311(.dina(w_n1179_1[0]),.dinb(w_n281_44[0]),.dout(n1574),.clk(gclk));
	jand g1312(.dina(w_n1175_1[0]),.dinb(w_n292_44[0]),.dout(n1575),.clk(gclk));
	jor g1313(.dina(n1575),.dinb(n1574),.dout(n1576),.clk(gclk));
	jand g1314(.dina(w_n1288_1[0]),.dinb(w_n304_44[0]),.dout(n1577),.clk(gclk));
	jor g1315(.dina(w_dff_B_PjZlxOwU2_0),.dinb(n1576),.dout(n1578),.clk(gclk));
	jor g1316(.dina(n1578),.dinb(w_dff_B_qU6FUjGM9_1),.dout(n1579),.clk(gclk));
	jand g1317(.dina(w_n1579_1[1]),.dinb(w_n364_58[2]),.dout(n1580),.clk(gclk));
	jor g1318(.dina(n1580),.dinb(n1572),.dout(n1581),.clk(gclk));
	jand g1319(.dina(w_n1240_1[0]),.dinb(w_n281_43[2]),.dout(n1582),.clk(gclk));
	jand g1320(.dina(w_n1171_1[0]),.dinb(w_n304_43[2]),.dout(n1583),.clk(gclk));
	jand g1321(.dina(w_n1236_1[0]),.dinb(w_n292_43[2]),.dout(n1584),.clk(gclk));
	jor g1322(.dina(n1584),.dinb(n1583),.dout(n1585),.clk(gclk));
	jand g1323(.dina(w_n1245_1[0]),.dinb(w_n267_43[2]),.dout(n1586),.clk(gclk));
	jor g1324(.dina(w_dff_B_znXfgxXr4_0),.dinb(n1585),.dout(n1587),.clk(gclk));
	jor g1325(.dina(n1587),.dinb(w_dff_B_l9iXkasH1_1),.dout(n1588),.clk(gclk));
	jand g1326(.dina(w_n1588_1[1]),.dinb(w_n319_58[2]),.dout(n1589),.clk(gclk));
	jor g1327(.dina(w_dff_B_1GbEw4ra1_0),.dinb(n1581),.dout(n1590),.clk(gclk));
	jor g1328(.dina(n1590),.dinb(w_dff_B_oaC8QtX88_1),.dout(n1591),.clk(gclk));
	jor g1329(.dina(w_n1591_0[1]),.dinb(w_n263_61[0]),.dout(n1592),.clk(gclk));
	jand g1330(.dina(w_n1329_1[0]),.dinb(w_n304_43[1]),.dout(n1593),.clk(gclk));
	jand g1331(.dina(w_n1283_1[0]),.dinb(w_n281_43[1]),.dout(n1594),.clk(gclk));
	jand g1332(.dina(w_n1279_1[0]),.dinb(w_n292_43[1]),.dout(n1595),.clk(gclk));
	jor g1333(.dina(n1595),.dinb(n1594),.dout(n1596),.clk(gclk));
	jand g1334(.dina(w_n1275_1[0]),.dinb(w_n267_43[1]),.dout(n1597),.clk(gclk));
	jor g1335(.dina(w_dff_B_LderWme62_0),.dinb(n1596),.dout(n1598),.clk(gclk));
	jor g1336(.dina(n1598),.dinb(w_dff_B_fkSCvyox5_1),.dout(n1599),.clk(gclk));
	jand g1337(.dina(w_n1599_1[1]),.dinb(w_n410_58[1]),.dout(n1600),.clk(gclk));
	jand g1338(.dina(w_n1255_1[0]),.dinb(w_n267_43[0]),.dout(n1601),.clk(gclk));
	jand g1339(.dina(w_n1263_1[0]),.dinb(w_n281_43[0]),.dout(n1602),.clk(gclk));
	jand g1340(.dina(w_n1259_1[0]),.dinb(w_n292_43[0]),.dout(n1603),.clk(gclk));
	jor g1341(.dina(n1603),.dinb(n1602),.dout(n1604),.clk(gclk));
	jand g1342(.dina(w_n1295_1[0]),.dinb(w_n304_43[0]),.dout(n1605),.clk(gclk));
	jor g1343(.dina(w_dff_B_yoRicxHq6_0),.dinb(n1604),.dout(n1606),.clk(gclk));
	jor g1344(.dina(n1606),.dinb(w_dff_B_HugGMlsl5_1),.dout(n1607),.clk(gclk));
	jand g1345(.dina(w_n1607_1[1]),.dinb(w_n319_58[1]),.dout(n1608),.clk(gclk));
	jand g1346(.dina(w_n1268_1[0]),.dinb(w_n304_42[2]),.dout(n1609),.clk(gclk));
	jand g1347(.dina(w_n1324_1[0]),.dinb(w_n281_42[2]),.dout(n1610),.clk(gclk));
	jand g1348(.dina(w_n1316_1[0]),.dinb(w_n267_42[2]),.dout(n1611),.clk(gclk));
	jor g1349(.dina(n1611),.dinb(n1610),.dout(n1612),.clk(gclk));
	jand g1350(.dina(w_n1320_1[0]),.dinb(w_n292_42[2]),.dout(n1613),.clk(gclk));
	jor g1351(.dina(w_dff_B_4lNWY1Cp4_0),.dinb(n1612),.dout(n1614),.clk(gclk));
	jor g1352(.dina(n1614),.dinb(w_dff_B_Dr5Rgvhi0_1),.dout(n1615),.clk(gclk));
	jand g1353(.dina(w_n1615_1[1]),.dinb(w_n265_58[1]),.dout(n1616),.clk(gclk));
	jor g1354(.dina(n1616),.dinb(n1608),.dout(n1617),.clk(gclk));
	jand g1355(.dina(w_n1308_1[0]),.dinb(w_n267_42[1]),.dout(n1618),.clk(gclk));
	jand g1356(.dina(w_n1303_1[0]),.dinb(w_n281_42[1]),.dout(n1619),.clk(gclk));
	jand g1357(.dina(w_n1299_1[0]),.dinb(w_n292_42[1]),.dout(n1620),.clk(gclk));
	jor g1358(.dina(n1620),.dinb(n1619),.dout(n1621),.clk(gclk));
	jand g1359(.dina(w_n1224_1[0]),.dinb(w_n304_42[1]),.dout(n1622),.clk(gclk));
	jor g1360(.dina(w_dff_B_CGPI3dHX3_0),.dinb(n1621),.dout(n1623),.clk(gclk));
	jor g1361(.dina(n1623),.dinb(w_dff_B_m13q85Av4_1),.dout(n1624),.clk(gclk));
	jand g1362(.dina(w_n1624_1[1]),.dinb(w_n364_58[1]),.dout(n1625),.clk(gclk));
	jor g1363(.dina(w_dff_B_nrM5oNz77_0),.dinb(n1617),.dout(n1626),.clk(gclk));
	jor g1364(.dina(n1626),.dinb(w_dff_B_zMcDdjhX8_1),.dout(n1627),.clk(gclk));
	jor g1365(.dina(w_n1627_0[1]),.dinb(w_shift6_61[0]),.dout(n1628),.clk(gclk));
	jand g1366(.dina(n1628),.dinb(n1592),.dout(result7),.clk(gclk));
	jand g1367(.dina(w_n292_42[0]),.dinb(w_n278_0[2]),.dout(n1630),.clk(gclk));
	jand g1368(.dina(w_n313_0[2]),.dinb(w_n281_42[0]),.dout(n1631),.clk(gclk));
	jand g1369(.dina(w_n328_0[2]),.dinb(w_n267_42[0]),.dout(n1632),.clk(gclk));
	jor g1370(.dina(n1632),.dinb(n1631),.dout(n1633),.clk(gclk));
	jand g1371(.dina(w_n338_0[2]),.dinb(w_n304_42[0]),.dout(n1634),.clk(gclk));
	jor g1372(.dina(w_dff_B_yS8ELcW17_0),.dinb(n1633),.dout(n1635),.clk(gclk));
	jor g1373(.dina(n1635),.dinb(w_dff_B_9A8x5XsH6_1),.dout(n1636),.clk(gclk));
	jand g1374(.dina(w_n1636_1[1]),.dinb(w_n265_58[0]),.dout(n1637),.clk(gclk));
	jand g1375(.dina(w_n304_41[2]),.dinb(w_n290_0[2]),.dout(n1638),.clk(gclk));
	jand g1376(.dina(w_n450_0[2]),.dinb(w_n281_41[2]),.dout(n1639),.clk(gclk));
	jand g1377(.dina(w_n301_0[2]),.dinb(w_n267_41[2]),.dout(n1640),.clk(gclk));
	jor g1378(.dina(n1640),.dinb(n1639),.dout(n1641),.clk(gclk));
	jand g1379(.dina(w_n419_0[2]),.dinb(w_n292_41[2]),.dout(n1642),.clk(gclk));
	jor g1380(.dina(w_dff_B_GJ9JITL81_0),.dinb(n1641),.dout(n1643),.clk(gclk));
	jor g1381(.dina(n1643),.dinb(w_dff_B_fPXeCm1I9_1),.dout(n1644),.clk(gclk));
	jand g1382(.dina(w_n1644_1[1]),.dinb(w_n410_58[0]),.dout(n1645),.clk(gclk));
	jand g1383(.dina(w_n476_0[2]),.dinb(w_n304_41[1]),.dout(n1646),.clk(gclk));
	jand g1384(.dina(w_n373_0[2]),.dinb(w_n281_41[1]),.dout(n1647),.clk(gclk));
	jand g1385(.dina(w_n393_0[2]),.dinb(w_n292_41[1]),.dout(n1648),.clk(gclk));
	jor g1386(.dina(n1648),.dinb(n1647),.dout(n1649),.clk(gclk));
	jand g1387(.dina(w_n466_0[2]),.dinb(w_n267_41[1]),.dout(n1650),.clk(gclk));
	jor g1388(.dina(w_dff_B_vqKakcLX8_0),.dinb(n1649),.dout(n1651),.clk(gclk));
	jor g1389(.dina(n1651),.dinb(w_dff_B_9liRMWfx0_1),.dout(n1652),.clk(gclk));
	jand g1390(.dina(w_n1652_1[1]),.dinb(w_n364_58[0]),.dout(n1653),.clk(gclk));
	jor g1391(.dina(n1653),.dinb(n1645),.dout(n1654),.clk(gclk));
	jand g1392(.dina(w_n348_0[2]),.dinb(w_n292_41[0]),.dout(n1655),.clk(gclk));
	jand g1393(.dina(w_n359_0[2]),.dinb(w_n281_41[0]),.dout(n1656),.clk(gclk));
	jand g1394(.dina(w_n404_0[2]),.dinb(w_n267_41[0]),.dout(n1657),.clk(gclk));
	jor g1395(.dina(n1657),.dinb(n1656),.dout(n1658),.clk(gclk));
	jand g1396(.dina(w_n383_0[2]),.dinb(w_n304_41[0]),.dout(n1659),.clk(gclk));
	jor g1397(.dina(w_dff_B_U4CRJqxg3_0),.dinb(n1658),.dout(n1660),.clk(gclk));
	jor g1398(.dina(n1660),.dinb(w_dff_B_QBBmk80V1_1),.dout(n1661),.clk(gclk));
	jand g1399(.dina(w_n1661_1[1]),.dinb(w_n319_58[0]),.dout(n1662),.clk(gclk));
	jor g1400(.dina(w_dff_B_9vGQxAeC7_0),.dinb(n1654),.dout(n1663),.clk(gclk));
	jor g1401(.dina(n1663),.dinb(w_dff_B_qvsR5x1d9_1),.dout(n1664),.clk(gclk));
	jor g1402(.dina(w_n1664_0[1]),.dinb(w_n263_60[2]),.dout(n1665),.clk(gclk));
	jand g1403(.dina(w_n486_0[2]),.dinb(w_n292_40[2]),.dout(n1666),.clk(gclk));
	jand g1404(.dina(w_n497_0[2]),.dinb(w_n281_40[2]),.dout(n1667),.clk(gclk));
	jand g1405(.dina(w_n574_0[2]),.dinb(w_n267_40[2]),.dout(n1668),.clk(gclk));
	jor g1406(.dina(n1668),.dinb(n1667),.dout(n1669),.clk(gclk));
	jand g1407(.dina(w_n564_0[2]),.dinb(w_n304_40[2]),.dout(n1670),.clk(gclk));
	jor g1408(.dina(w_dff_B_qHBfuMtU9_0),.dinb(n1669),.dout(n1671),.clk(gclk));
	jor g1409(.dina(n1671),.dinb(w_dff_B_aGDLZ7hj2_1),.dout(n1672),.clk(gclk));
	jand g1410(.dina(w_n1672_1[1]),.dinb(w_n410_57[2]),.dout(n1673),.clk(gclk));
	jand g1411(.dina(w_n609_0[2]),.dinb(w_n304_40[1]),.dout(n1674),.clk(gclk));
	jand g1412(.dina(w_n541_0[2]),.dinb(w_n281_40[1]),.dout(n1675),.clk(gclk));
	jand g1413(.dina(w_n530_0[2]),.dinb(w_n292_40[1]),.dout(n1676),.clk(gclk));
	jor g1414(.dina(n1676),.dinb(n1675),.dout(n1677),.clk(gclk));
	jand g1415(.dina(w_n619_0[2]),.dinb(w_n267_40[1]),.dout(n1678),.clk(gclk));
	jor g1416(.dina(w_dff_B_yLZkh10I4_0),.dinb(n1677),.dout(n1679),.clk(gclk));
	jor g1417(.dina(n1679),.dinb(w_dff_B_f0Wxj4yd8_1),.dout(n1680),.clk(gclk));
	jand g1418(.dina(w_n1680_1[1]),.dinb(w_n319_57[2]),.dout(n1681),.clk(gclk));
	jand g1419(.dina(w_n439_0[2]),.dinb(w_n267_40[0]),.dout(n1682),.clk(gclk));
	jand g1420(.dina(w_n630_0[2]),.dinb(w_n281_40[0]),.dout(n1683),.clk(gclk));
	jand g1421(.dina(w_n599_0[2]),.dinb(w_n292_40[0]),.dout(n1684),.clk(gclk));
	jor g1422(.dina(n1684),.dinb(n1683),.dout(n1685),.clk(gclk));
	jand g1423(.dina(w_n429_0[2]),.dinb(w_n304_40[0]),.dout(n1686),.clk(gclk));
	jor g1424(.dina(w_dff_B_fPFHHo2p6_0),.dinb(n1685),.dout(n1687),.clk(gclk));
	jor g1425(.dina(n1687),.dinb(w_dff_B_m7kHuDJE5_1),.dout(n1688),.clk(gclk));
	jand g1426(.dina(w_n1688_1[1]),.dinb(w_n364_57[2]),.dout(n1689),.clk(gclk));
	jor g1427(.dina(n1689),.dinb(n1681),.dout(n1690),.clk(gclk));
	jand g1428(.dina(w_n554_0[2]),.dinb(w_n292_39[2]),.dout(n1691),.clk(gclk));
	jand g1429(.dina(w_n585_0[2]),.dinb(w_n281_39[2]),.dout(n1692),.clk(gclk));
	jand g1430(.dina(w_n510_0[2]),.dinb(w_n267_39[2]),.dout(n1693),.clk(gclk));
	jor g1431(.dina(n1693),.dinb(n1692),.dout(n1694),.clk(gclk));
	jand g1432(.dina(w_n520_0[2]),.dinb(w_n304_39[2]),.dout(n1695),.clk(gclk));
	jor g1433(.dina(w_dff_B_YOOdvGcg9_0),.dinb(n1694),.dout(n1696),.clk(gclk));
	jor g1434(.dina(n1696),.dinb(w_dff_B_WSOvahUp7_1),.dout(n1697),.clk(gclk));
	jand g1435(.dina(w_n1697_1[1]),.dinb(w_n265_57[2]),.dout(n1698),.clk(gclk));
	jor g1436(.dina(w_dff_B_8IFA9uxn4_0),.dinb(n1690),.dout(n1699),.clk(gclk));
	jor g1437(.dina(n1699),.dinb(w_dff_B_NPGtS0aV6_1),.dout(n1700),.clk(gclk));
	jor g1438(.dina(w_n1700_0[1]),.dinb(w_shift6_60[2]),.dout(n1701),.clk(gclk));
	jand g1439(.dina(n1701),.dinb(n1665),.dout(result8),.clk(gclk));
	jand g1440(.dina(w_n647_0[2]),.dinb(w_n292_39[1]),.dout(n1703),.clk(gclk));
	jand g1441(.dina(w_n678_0[2]),.dinb(w_n281_39[1]),.dout(n1704),.clk(gclk));
	jand g1442(.dina(w_n827_0[2]),.dinb(w_n267_39[1]),.dout(n1705),.clk(gclk));
	jor g1443(.dina(n1705),.dinb(n1704),.dout(n1706),.clk(gclk));
	jand g1444(.dina(w_n837_0[2]),.dinb(w_n304_39[1]),.dout(n1707),.clk(gclk));
	jor g1445(.dina(w_dff_B_02mnb2b89_0),.dinb(n1706),.dout(n1708),.clk(gclk));
	jor g1446(.dina(n1708),.dinb(w_dff_B_FiNXkb9Y6_1),.dout(n1709),.clk(gclk));
	jand g1447(.dina(w_n1709_1[1]),.dinb(w_n364_57[1]),.dout(n1710),.clk(gclk));
	jand g1448(.dina(w_n701_0[2]),.dinb(w_n304_39[0]),.dout(n1711),.clk(gclk));
	jand g1449(.dina(w_n735_0[2]),.dinb(w_n281_39[0]),.dout(n1712),.clk(gclk));
	jand g1450(.dina(w_n766_0[2]),.dinb(w_n292_39[0]),.dout(n1713),.clk(gclk));
	jor g1451(.dina(n1713),.dinb(n1712),.dout(n1714),.clk(gclk));
	jand g1452(.dina(w_n691_0[2]),.dinb(w_n267_39[0]),.dout(n1715),.clk(gclk));
	jor g1453(.dina(w_dff_B_0KacSSWA2_0),.dinb(n1714),.dout(n1716),.clk(gclk));
	jor g1454(.dina(n1716),.dinb(w_dff_B_3w20PdWI5_1),.dout(n1717),.clk(gclk));
	jand g1455(.dina(w_n1717_1[1]),.dinb(w_n410_57[1]),.dout(n1718),.clk(gclk));
	jand g1456(.dina(w_n711_0[2]),.dinb(w_n292_38[2]),.dout(n1719),.clk(gclk));
	jand g1457(.dina(w_n722_0[2]),.dinb(w_n281_38[2]),.dout(n1720),.clk(gclk));
	jand g1458(.dina(w_n780_0[2]),.dinb(w_n267_38[2]),.dout(n1721),.clk(gclk));
	jor g1459(.dina(n1721),.dinb(n1720),.dout(n1722),.clk(gclk));
	jand g1460(.dina(w_n790_0[2]),.dinb(w_n304_38[2]),.dout(n1723),.clk(gclk));
	jor g1461(.dina(w_dff_B_N0xQg3RU2_0),.dinb(n1722),.dout(n1724),.clk(gclk));
	jor g1462(.dina(n1724),.dinb(w_dff_B_XgKuybAs2_1),.dout(n1725),.clk(gclk));
	jand g1463(.dina(w_n1725_1[1]),.dinb(w_n265_57[1]),.dout(n1726),.clk(gclk));
	jor g1464(.dina(n1726),.dinb(n1718),.dout(n1727),.clk(gclk));
	jand g1465(.dina(w_n800_0[2]),.dinb(w_n292_38[1]),.dout(n1728),.clk(gclk));
	jand g1466(.dina(w_n811_0[2]),.dinb(w_n281_38[1]),.dout(n1729),.clk(gclk));
	jand g1467(.dina(w_n667_0[2]),.dinb(w_n267_38[1]),.dout(n1730),.clk(gclk));
	jor g1468(.dina(n1730),.dinb(n1729),.dout(n1731),.clk(gclk));
	jand g1469(.dina(w_n657_0[2]),.dinb(w_n304_38[1]),.dout(n1732),.clk(gclk));
	jor g1470(.dina(w_dff_B_DXN0HrMN5_0),.dinb(n1731),.dout(n1733),.clk(gclk));
	jor g1471(.dina(n1733),.dinb(w_dff_B_iuUN1MS12_1),.dout(n1734),.clk(gclk));
	jand g1472(.dina(w_n1734_1[1]),.dinb(w_n319_57[1]),.dout(n1735),.clk(gclk));
	jor g1473(.dina(w_dff_B_nuqFSaDm4_0),.dinb(n1727),.dout(n1736),.clk(gclk));
	jor g1474(.dina(n1736),.dinb(w_dff_B_LLMoJvwo6_1),.dout(n1737),.clk(gclk));
	jor g1475(.dina(w_n1737_0[1]),.dinb(w_n263_60[1]),.dout(n1738),.clk(gclk));
	jand g1476(.dina(w_n881_0[2]),.dinb(w_n304_38[0]),.dout(n1739),.clk(gclk));
	jand g1477(.dina(w_n946_0[2]),.dinb(w_n281_38[0]),.dout(n1740),.clk(gclk));
	jand g1478(.dina(w_n935_0[2]),.dinb(w_n292_38[0]),.dout(n1741),.clk(gclk));
	jor g1479(.dina(n1741),.dinb(n1740),.dout(n1742),.clk(gclk));
	jand g1480(.dina(w_n871_0[2]),.dinb(w_n267_38[0]),.dout(n1743),.clk(gclk));
	jor g1481(.dina(w_dff_B_t7mqydWt3_0),.dinb(n1742),.dout(n1744),.clk(gclk));
	jor g1482(.dina(n1744),.dinb(w_dff_B_PPfha8iG0_1),.dout(n1745),.clk(gclk));
	jand g1483(.dina(w_n1745_1[1]),.dinb(w_n265_57[0]),.dout(n1746),.clk(gclk));
	jand g1484(.dina(w_n891_0[2]),.dinb(w_n292_37[2]),.dout(n1747),.clk(gclk));
	jand g1485(.dina(w_n902_0[2]),.dinb(w_n281_37[2]),.dout(n1748),.clk(gclk));
	jand g1486(.dina(w_n980_0[2]),.dinb(w_n267_37[2]),.dout(n1749),.clk(gclk));
	jor g1487(.dina(n1749),.dinb(n1748),.dout(n1750),.clk(gclk));
	jand g1488(.dina(w_n970_0[2]),.dinb(w_n304_37[2]),.dout(n1751),.clk(gclk));
	jor g1489(.dina(w_dff_B_aQl6SJho8_0),.dinb(n1750),.dout(n1752),.clk(gclk));
	jor g1490(.dina(n1752),.dinb(w_dff_B_RIw4JiM62_1),.dout(n1753),.clk(gclk));
	jand g1491(.dina(w_n1753_1[1]),.dinb(w_n319_57[0]),.dout(n1754),.clk(gclk));
	jand g1492(.dina(w_n960_0[2]),.dinb(w_n292_37[1]),.dout(n1755),.clk(gclk));
	jand g1493(.dina(w_n991_0[2]),.dinb(w_n281_37[1]),.dout(n1756),.clk(gclk));
	jand g1494(.dina(w_n755_0[2]),.dinb(w_n267_37[1]),.dout(n1757),.clk(gclk));
	jor g1495(.dina(n1757),.dinb(n1756),.dout(n1758),.clk(gclk));
	jand g1496(.dina(w_n745_0[2]),.dinb(w_n304_37[1]),.dout(n1759),.clk(gclk));
	jor g1497(.dina(w_dff_B_kjyfZ68B8_0),.dinb(n1758),.dout(n1760),.clk(gclk));
	jor g1498(.dina(n1760),.dinb(w_dff_B_Fg5kkHG93_1),.dout(n1761),.clk(gclk));
	jand g1499(.dina(w_n1761_1[1]),.dinb(w_n364_57[0]),.dout(n1762),.clk(gclk));
	jor g1500(.dina(n1762),.dinb(n1754),.dout(n1763),.clk(gclk));
	jand g1501(.dina(w_n847_0[2]),.dinb(w_n292_37[0]),.dout(n1764),.clk(gclk));
	jand g1502(.dina(w_n858_0[2]),.dinb(w_n281_37[0]),.dout(n1765),.clk(gclk));
	jand g1503(.dina(w_n915_0[2]),.dinb(w_n267_37[0]),.dout(n1766),.clk(gclk));
	jor g1504(.dina(n1766),.dinb(n1765),.dout(n1767),.clk(gclk));
	jand g1505(.dina(w_n925_0[2]),.dinb(w_n304_37[0]),.dout(n1768),.clk(gclk));
	jor g1506(.dina(w_dff_B_L33fN8wm0_0),.dinb(n1767),.dout(n1769),.clk(gclk));
	jor g1507(.dina(n1769),.dinb(w_dff_B_OSsMJ08H1_1),.dout(n1770),.clk(gclk));
	jand g1508(.dina(w_n1770_1[1]),.dinb(w_n410_57[0]),.dout(n1771),.clk(gclk));
	jor g1509(.dina(w_dff_B_OGeIt0NV8_0),.dinb(n1763),.dout(n1772),.clk(gclk));
	jor g1510(.dina(n1772),.dinb(w_dff_B_robiVxRf4_1),.dout(n1773),.clk(gclk));
	jor g1511(.dina(w_n1773_0[1]),.dinb(w_shift6_60[1]),.dout(n1774),.clk(gclk));
	jand g1512(.dina(n1774),.dinb(n1738),.dout(result9),.clk(gclk));
	jand g1513(.dina(w_n1067_0[2]),.dinb(w_n304_36[2]),.dout(n1776),.clk(gclk));
	jand g1514(.dina(w_n1015_0[2]),.dinb(w_n281_36[2]),.dout(n1777),.clk(gclk));
	jand g1515(.dina(w_n1002_0[2]),.dinb(w_n292_36[2]),.dout(n1778),.clk(gclk));
	jor g1516(.dina(n1778),.dinb(n1777),.dout(n1779),.clk(gclk));
	jand g1517(.dina(w_n1063_0[2]),.dinb(w_n267_36[2]),.dout(n1780),.clk(gclk));
	jor g1518(.dina(w_dff_B_XA3R5mLm5_0),.dinb(n1779),.dout(n1781),.clk(gclk));
	jor g1519(.dina(n1781),.dinb(w_dff_B_QmpjNxjn9_1),.dout(n1782),.clk(gclk));
	jand g1520(.dina(w_n1782_1[1]),.dinb(w_n319_56[2]),.dout(n1783),.clk(gclk));
	jand g1521(.dina(w_n1022_0[2]),.dinb(w_n267_36[1]),.dout(n1784),.clk(gclk));
	jand g1522(.dina(w_n1042_0[2]),.dinb(w_n281_36[1]),.dout(n1785),.clk(gclk));
	jand g1523(.dina(w_n1050_0[2]),.dinb(w_n292_36[1]),.dout(n1786),.clk(gclk));
	jor g1524(.dina(n1786),.dinb(n1785),.dout(n1787),.clk(gclk));
	jand g1525(.dina(w_n1026_0[2]),.dinb(w_n304_36[1]),.dout(n1788),.clk(gclk));
	jor g1526(.dina(w_dff_B_XXULzUgH7_0),.dinb(n1787),.dout(n1789),.clk(gclk));
	jor g1527(.dina(n1789),.dinb(w_dff_B_Z0mTHOxn2_1),.dout(n1790),.clk(gclk));
	jand g1528(.dina(w_n1790_1[1]),.dinb(w_n410_56[2]),.dout(n1791),.clk(gclk));
	jand g1529(.dina(w_n1010_0[2]),.dinb(w_n267_36[0]),.dout(n1792),.clk(gclk));
	jand g1530(.dina(w_n1035_0[2]),.dinb(w_n281_36[0]),.dout(n1793),.clk(gclk));
	jand g1531(.dina(w_n1030_0[2]),.dinb(w_n292_36[0]),.dout(n1794),.clk(gclk));
	jor g1532(.dina(n1794),.dinb(n1793),.dout(n1795),.clk(gclk));
	jand g1533(.dina(w_n1006_0[2]),.dinb(w_n304_36[0]),.dout(n1796),.clk(gclk));
	jor g1534(.dina(w_dff_B_1jugmf9a1_0),.dinb(n1795),.dout(n1797),.clk(gclk));
	jor g1535(.dina(n1797),.dinb(w_dff_B_iky6qif53_1),.dout(n1798),.clk(gclk));
	jand g1536(.dina(w_n1798_1[1]),.dinb(w_n265_56[2]),.dout(n1799),.clk(gclk));
	jor g1537(.dina(n1799),.dinb(n1791),.dout(n1800),.clk(gclk));
	jand g1538(.dina(w_n1090_0[2]),.dinb(w_n304_35[2]),.dout(n1801),.clk(gclk));
	jand g1539(.dina(w_n1076_0[2]),.dinb(w_n281_35[2]),.dout(n1802),.clk(gclk));
	jand g1540(.dina(w_n1071_0[2]),.dinb(w_n292_35[2]),.dout(n1803),.clk(gclk));
	jor g1541(.dina(n1803),.dinb(n1802),.dout(n1804),.clk(gclk));
	jand g1542(.dina(w_n1094_0[2]),.dinb(w_n267_35[2]),.dout(n1805),.clk(gclk));
	jor g1543(.dina(w_dff_B_nUofu0Ki0_0),.dinb(n1804),.dout(n1806),.clk(gclk));
	jor g1544(.dina(n1806),.dinb(w_dff_B_Fa5UygcP0_1),.dout(n1807),.clk(gclk));
	jand g1545(.dina(w_n1807_1[1]),.dinb(w_n364_56[2]),.dout(n1808),.clk(gclk));
	jor g1546(.dina(w_dff_B_g96jNHdJ1_0),.dinb(n1800),.dout(n1809),.clk(gclk));
	jor g1547(.dina(n1809),.dinb(w_dff_B_cP0exCf09_1),.dout(n1810),.clk(gclk));
	jor g1548(.dina(w_n1810_0[1]),.dinb(w_n263_60[0]),.dout(n1811),.clk(gclk));
	jand g1549(.dina(w_n1046_0[2]),.dinb(w_n304_35[1]),.dout(n1812),.clk(gclk));
	jand g1550(.dina(w_n1126_0[2]),.dinb(w_n281_35[1]),.dout(n1813),.clk(gclk));
	jand g1551(.dina(w_n1055_0[2]),.dinb(w_n267_35[1]),.dout(n1814),.clk(gclk));
	jor g1552(.dina(n1814),.dinb(n1813),.dout(n1815),.clk(gclk));
	jand g1553(.dina(w_n1134_0[2]),.dinb(w_n292_35[1]),.dout(n1816),.clk(gclk));
	jor g1554(.dina(w_dff_B_bqScnAXr8_0),.dinb(n1815),.dout(n1817),.clk(gclk));
	jor g1555(.dina(n1817),.dinb(w_dff_B_BBYKbmq80_1),.dout(n1818),.clk(gclk));
	jand g1556(.dina(w_n1818_1[1]),.dinb(w_n364_56[1]),.dout(n1819),.clk(gclk));
	jand g1557(.dina(w_n1119_0[2]),.dinb(w_n292_35[0]),.dout(n1820),.clk(gclk));
	jand g1558(.dina(w_n1106_0[2]),.dinb(w_n281_35[0]),.dout(n1821),.clk(gclk));
	jand g1559(.dina(w_n1139_0[2]),.dinb(w_n267_35[0]),.dout(n1822),.clk(gclk));
	jor g1560(.dina(n1822),.dinb(n1821),.dout(n1823),.clk(gclk));
	jand g1561(.dina(w_n1130_0[2]),.dinb(w_n304_35[0]),.dout(n1824),.clk(gclk));
	jor g1562(.dina(w_dff_B_aP2Vzczj8_0),.dinb(n1823),.dout(n1825),.clk(gclk));
	jor g1563(.dina(n1825),.dinb(w_dff_B_vZrVtr4g8_1),.dout(n1826),.clk(gclk));
	jand g1564(.dina(w_n1826_1[1]),.dinb(w_n319_56[1]),.dout(n1827),.clk(gclk));
	jand g1565(.dina(w_n1110_0[2]),.dinb(w_n304_34[2]),.dout(n1828),.clk(gclk));
	jand g1566(.dina(w_n1160_0[2]),.dinb(w_n281_34[2]),.dout(n1829),.clk(gclk));
	jand g1567(.dina(w_n1114_0[2]),.dinb(w_n267_34[2]),.dout(n1830),.clk(gclk));
	jor g1568(.dina(n1830),.dinb(n1829),.dout(n1831),.clk(gclk));
	jand g1569(.dina(w_n1155_0[2]),.dinb(w_n292_34[2]),.dout(n1832),.clk(gclk));
	jor g1570(.dina(w_dff_B_lFefcJ9l1_0),.dinb(n1831),.dout(n1833),.clk(gclk));
	jor g1571(.dina(n1833),.dinb(w_dff_B_vFRPZe0E7_1),.dout(n1834),.clk(gclk));
	jand g1572(.dina(w_n1834_1[1]),.dinb(w_n265_56[1]),.dout(n1835),.clk(gclk));
	jor g1573(.dina(n1835),.dinb(n1827),.dout(n1836),.clk(gclk));
	jand g1574(.dina(w_n1151_0[2]),.dinb(w_n304_34[1]),.dout(n1837),.clk(gclk));
	jand g1575(.dina(w_n1099_0[2]),.dinb(w_n281_34[1]),.dout(n1838),.clk(gclk));
	jand g1576(.dina(w_n1086_0[2]),.dinb(w_n292_34[1]),.dout(n1839),.clk(gclk));
	jor g1577(.dina(n1839),.dinb(n1838),.dout(n1840),.clk(gclk));
	jand g1578(.dina(w_n1147_0[2]),.dinb(w_n267_34[1]),.dout(n1841),.clk(gclk));
	jor g1579(.dina(w_dff_B_XBiAr6HB6_0),.dinb(n1840),.dout(n1842),.clk(gclk));
	jor g1580(.dina(n1842),.dinb(w_dff_B_buHD2ggE4_1),.dout(n1843),.clk(gclk));
	jand g1581(.dina(w_n1843_1[1]),.dinb(w_n410_56[1]),.dout(n1844),.clk(gclk));
	jor g1582(.dina(w_dff_B_h1n7C7xB6_0),.dinb(n1836),.dout(n1845),.clk(gclk));
	jor g1583(.dina(n1845),.dinb(w_dff_B_ETLDoBFx5_1),.dout(n1846),.clk(gclk));
	jor g1584(.dina(w_n1846_0[1]),.dinb(w_shift6_60[0]),.dout(n1847),.clk(gclk));
	jand g1585(.dina(n1847),.dinb(n1811),.dout(result10),.clk(gclk));
	jand g1586(.dina(w_n1245_0[2]),.dinb(w_n281_34[0]),.dout(n1849),.clk(gclk));
	jand g1587(.dina(w_n1171_0[2]),.dinb(w_n267_34[0]),.dout(n1850),.clk(gclk));
	jand g1588(.dina(w_n1240_0[2]),.dinb(w_n292_34[0]),.dout(n1851),.clk(gclk));
	jor g1589(.dina(n1851),.dinb(n1850),.dout(n1852),.clk(gclk));
	jand g1590(.dina(w_n1175_0[2]),.dinb(w_n304_34[0]),.dout(n1853),.clk(gclk));
	jor g1591(.dina(w_dff_B_6p5HSVjj5_0),.dinb(n1852),.dout(n1854),.clk(gclk));
	jor g1592(.dina(n1854),.dinb(w_dff_B_BhqJTvgw6_1),.dout(n1855),.clk(gclk));
	jand g1593(.dina(w_n1855_1[1]),.dinb(w_n319_56[0]),.dout(n1856),.clk(gclk));
	jand g1594(.dina(w_n1195_0[2]),.dinb(w_n304_33[2]),.dout(n1857),.clk(gclk));
	jand g1595(.dina(w_n1211_0[2]),.dinb(w_n281_33[2]),.dout(n1858),.clk(gclk));
	jand g1596(.dina(w_n1219_0[2]),.dinb(w_n292_33[2]),.dout(n1859),.clk(gclk));
	jor g1597(.dina(n1859),.dinb(n1858),.dout(n1860),.clk(gclk));
	jand g1598(.dina(w_n1199_0[2]),.dinb(w_n267_33[2]),.dout(n1861),.clk(gclk));
	jor g1599(.dina(w_dff_B_W1m7NuUn4_0),.dinb(n1860),.dout(n1862),.clk(gclk));
	jor g1600(.dina(n1862),.dinb(w_dff_B_mQYVjC3V5_1),.dout(n1863),.clk(gclk));
	jand g1601(.dina(w_n1863_1[1]),.dinb(w_n410_56[0]),.dout(n1864),.clk(gclk));
	jand g1602(.dina(w_n1236_0[2]),.dinb(w_n304_33[1]),.dout(n1865),.clk(gclk));
	jand g1603(.dina(w_n1191_0[2]),.dinb(w_n281_33[1]),.dout(n1866),.clk(gclk));
	jand g1604(.dina(w_n1204_0[2]),.dinb(w_n292_33[1]),.dout(n1867),.clk(gclk));
	jor g1605(.dina(n1867),.dinb(n1866),.dout(n1868),.clk(gclk));
	jand g1606(.dina(w_n1232_0[2]),.dinb(w_n267_33[1]),.dout(n1869),.clk(gclk));
	jor g1607(.dina(w_dff_B_LXLqwXQf5_0),.dinb(n1868),.dout(n1870),.clk(gclk));
	jor g1608(.dina(n1870),.dinb(w_dff_B_U7tofJv50_1),.dout(n1871),.clk(gclk));
	jand g1609(.dina(w_n1871_1[1]),.dinb(w_n265_56[0]),.dout(n1872),.clk(gclk));
	jor g1610(.dina(n1872),.dinb(n1864),.dout(n1873),.clk(gclk));
	jand g1611(.dina(w_n1279_0[2]),.dinb(w_n304_33[0]),.dout(n1874),.clk(gclk));
	jand g1612(.dina(w_n1184_0[2]),.dinb(w_n281_33[0]),.dout(n1875),.clk(gclk));
	jand g1613(.dina(w_n1288_0[2]),.dinb(w_n267_33[0]),.dout(n1876),.clk(gclk));
	jor g1614(.dina(n1876),.dinb(n1875),.dout(n1877),.clk(gclk));
	jand g1615(.dina(w_n1179_0[2]),.dinb(w_n292_33[0]),.dout(n1878),.clk(gclk));
	jor g1616(.dina(w_dff_B_WWcxEztL0_0),.dinb(n1877),.dout(n1879),.clk(gclk));
	jor g1617(.dina(n1879),.dinb(w_dff_B_12bjiM417_1),.dout(n1880),.clk(gclk));
	jand g1618(.dina(w_n1880_1[1]),.dinb(w_n364_56[0]),.dout(n1881),.clk(gclk));
	jor g1619(.dina(w_dff_B_NmnoyRaM2_0),.dinb(n1873),.dout(n1882),.clk(gclk));
	jor g1620(.dina(n1882),.dinb(w_dff_B_55Edj9Zy7_1),.dout(n1883),.clk(gclk));
	jor g1621(.dina(w_n1883_0[1]),.dinb(w_n263_59[2]),.dout(n1884),.clk(gclk));
	jand g1622(.dina(w_n1320_0[2]),.dinb(w_n304_32[2]),.dout(n1885),.clk(gclk));
	jand g1623(.dina(w_n1275_0[2]),.dinb(w_n281_32[2]),.dout(n1886),.clk(gclk));
	jand g1624(.dina(w_n1283_0[2]),.dinb(w_n292_32[2]),.dout(n1887),.clk(gclk));
	jor g1625(.dina(n1887),.dinb(n1886),.dout(n1888),.clk(gclk));
	jand g1626(.dina(w_n1329_0[2]),.dinb(w_n267_32[2]),.dout(n1889),.clk(gclk));
	jor g1627(.dina(w_dff_B_a27ha2GA3_0),.dinb(n1888),.dout(n1890),.clk(gclk));
	jor g1628(.dina(n1890),.dinb(w_dff_B_FCK49IvL3_1),.dout(n1891),.clk(gclk));
	jand g1629(.dina(w_n1891_1[1]),.dinb(w_n410_55[2]),.dout(n1892),.clk(gclk));
	jand g1630(.dina(w_n1299_0[2]),.dinb(w_n304_32[1]),.dout(n1893),.clk(gclk));
	jand g1631(.dina(w_n1255_0[2]),.dinb(w_n281_32[1]),.dout(n1894),.clk(gclk));
	jand g1632(.dina(w_n1263_0[2]),.dinb(w_n292_32[1]),.dout(n1895),.clk(gclk));
	jor g1633(.dina(n1895),.dinb(n1894),.dout(n1896),.clk(gclk));
	jand g1634(.dina(w_n1295_0[2]),.dinb(w_n267_32[1]),.dout(n1897),.clk(gclk));
	jor g1635(.dina(w_dff_B_u3s452In8_0),.dinb(n1896),.dout(n1898),.clk(gclk));
	jor g1636(.dina(n1898),.dinb(w_dff_B_cC9wJqdw1_1),.dout(n1899),.clk(gclk));
	jand g1637(.dina(w_n1899_1[1]),.dinb(w_n319_55[2]),.dout(n1900),.clk(gclk));
	jand g1638(.dina(w_n1259_0[2]),.dinb(w_n304_32[0]),.dout(n1901),.clk(gclk));
	jand g1639(.dina(w_n1316_0[2]),.dinb(w_n281_32[0]),.dout(n1902),.clk(gclk));
	jand g1640(.dina(w_n1324_0[2]),.dinb(w_n292_32[0]),.dout(n1903),.clk(gclk));
	jor g1641(.dina(n1903),.dinb(n1902),.dout(n1904),.clk(gclk));
	jand g1642(.dina(w_n1268_0[2]),.dinb(w_n267_32[0]),.dout(n1905),.clk(gclk));
	jor g1643(.dina(w_dff_B_CwRb6Zdg9_0),.dinb(n1904),.dout(n1906),.clk(gclk));
	jor g1644(.dina(n1906),.dinb(w_dff_B_z6Mk3N4z7_1),.dout(n1907),.clk(gclk));
	jand g1645(.dina(w_n1907_1[1]),.dinb(w_n265_55[2]),.dout(n1908),.clk(gclk));
	jor g1646(.dina(n1908),.dinb(n1900),.dout(n1909),.clk(gclk));
	jand g1647(.dina(w_n1303_0[2]),.dinb(w_n292_31[2]),.dout(n1910),.clk(gclk));
	jand g1648(.dina(w_n1308_0[2]),.dinb(w_n281_31[2]),.dout(n1911),.clk(gclk));
	jand g1649(.dina(w_n1224_0[2]),.dinb(w_n267_31[2]),.dout(n1912),.clk(gclk));
	jor g1650(.dina(n1912),.dinb(n1911),.dout(n1913),.clk(gclk));
	jand g1651(.dina(w_n1215_0[2]),.dinb(w_n304_31[2]),.dout(n1914),.clk(gclk));
	jor g1652(.dina(w_dff_B_eFTihvvF4_0),.dinb(n1913),.dout(n1915),.clk(gclk));
	jor g1653(.dina(n1915),.dinb(w_dff_B_wM0cwS0E2_1),.dout(n1916),.clk(gclk));
	jand g1654(.dina(w_n1916_1[1]),.dinb(w_n364_55[2]),.dout(n1917),.clk(gclk));
	jor g1655(.dina(w_dff_B_m1xLLlKS6_0),.dinb(n1909),.dout(n1918),.clk(gclk));
	jor g1656(.dina(n1918),.dinb(w_dff_B_2a5xp3cf3_1),.dout(n1919),.clk(gclk));
	jor g1657(.dina(w_n1919_0[1]),.dinb(w_shift6_59[2]),.dout(n1920),.clk(gclk));
	jand g1658(.dina(n1920),.dinb(n1884),.dout(result11),.clk(gclk));
	jand g1659(.dina(w_n348_0[1]),.dinb(w_n304_31[1]),.dout(n1922),.clk(gclk));
	jand g1660(.dina(w_n328_0[1]),.dinb(w_n281_31[1]),.dout(n1923),.clk(gclk));
	jand g1661(.dina(w_n313_0[1]),.dinb(w_n292_31[1]),.dout(n1924),.clk(gclk));
	jor g1662(.dina(n1924),.dinb(n1923),.dout(n1925),.clk(gclk));
	jand g1663(.dina(w_n338_0[1]),.dinb(w_n267_31[1]),.dout(n1926),.clk(gclk));
	jor g1664(.dina(w_dff_B_U5D9P6Db9_0),.dinb(n1925),.dout(n1927),.clk(gclk));
	jor g1665(.dina(n1927),.dinb(w_dff_B_lH0Rc6Lf0_1),.dout(n1928),.clk(gclk));
	jand g1666(.dina(w_n1928_1[1]),.dinb(w_n265_55[1]),.dout(n1929),.clk(gclk));
	jand g1667(.dina(w_n304_31[0]),.dinb(w_n278_0[1]),.dout(n1930),.clk(gclk));
	jand g1668(.dina(w_n301_0[1]),.dinb(w_n281_31[0]),.dout(n1931),.clk(gclk));
	jand g1669(.dina(w_n450_0[1]),.dinb(w_n292_31[0]),.dout(n1932),.clk(gclk));
	jor g1670(.dina(n1932),.dinb(n1931),.dout(n1933),.clk(gclk));
	jand g1671(.dina(w_n290_0[1]),.dinb(w_n267_31[0]),.dout(n1934),.clk(gclk));
	jor g1672(.dina(w_dff_B_D38jD0K72_0),.dinb(n1933),.dout(n1935),.clk(gclk));
	jor g1673(.dina(n1935),.dinb(w_dff_B_Y7YtLhzO6_1),.dout(n1936),.clk(gclk));
	jand g1674(.dina(w_n1936_1[1]),.dinb(w_n410_55[1]),.dout(n1937),.clk(gclk));
	jand g1675(.dina(w_n486_0[1]),.dinb(w_n304_30[2]),.dout(n1938),.clk(gclk));
	jand g1676(.dina(w_n466_0[1]),.dinb(w_n281_30[2]),.dout(n1939),.clk(gclk));
	jand g1677(.dina(w_n476_0[1]),.dinb(w_n267_30[2]),.dout(n1940),.clk(gclk));
	jor g1678(.dina(n1940),.dinb(n1939),.dout(n1941),.clk(gclk));
	jand g1679(.dina(w_n373_0[1]),.dinb(w_n292_30[2]),.dout(n1942),.clk(gclk));
	jor g1680(.dina(w_dff_B_IpfWp5MV0_0),.dinb(n1941),.dout(n1943),.clk(gclk));
	jor g1681(.dina(n1943),.dinb(w_dff_B_HWXL2sOJ4_1),.dout(n1944),.clk(gclk));
	jand g1682(.dina(w_n1944_1[1]),.dinb(w_n364_55[1]),.dout(n1945),.clk(gclk));
	jor g1683(.dina(n1945),.dinb(n1937),.dout(n1946),.clk(gclk));
	jand g1684(.dina(w_n393_0[1]),.dinb(w_n304_30[1]),.dout(n1947),.clk(gclk));
	jand g1685(.dina(w_n404_0[1]),.dinb(w_n281_30[1]),.dout(n1948),.clk(gclk));
	jand g1686(.dina(w_n383_0[1]),.dinb(w_n267_30[1]),.dout(n1949),.clk(gclk));
	jor g1687(.dina(n1949),.dinb(n1948),.dout(n1950),.clk(gclk));
	jand g1688(.dina(w_n359_0[1]),.dinb(w_n292_30[1]),.dout(n1951),.clk(gclk));
	jor g1689(.dina(w_dff_B_g3hpVPxg1_0),.dinb(n1950),.dout(n1952),.clk(gclk));
	jor g1690(.dina(n1952),.dinb(w_dff_B_EQkAxmtM8_1),.dout(n1953),.clk(gclk));
	jand g1691(.dina(w_n1953_1[1]),.dinb(w_n319_55[1]),.dout(n1954),.clk(gclk));
	jor g1692(.dina(w_dff_B_BVk4GIky4_0),.dinb(n1946),.dout(n1955),.clk(gclk));
	jor g1693(.dina(n1955),.dinb(w_dff_B_Mfbpq3wo7_1),.dout(n1956),.clk(gclk));
	jor g1694(.dina(w_n1956_0[1]),.dinb(w_n263_59[1]),.dout(n1957),.clk(gclk));
	jand g1695(.dina(w_n419_0[1]),.dinb(w_n304_30[0]),.dout(n1958),.clk(gclk));
	jand g1696(.dina(w_n439_0[1]),.dinb(w_n281_30[0]),.dout(n1959),.clk(gclk));
	jand g1697(.dina(w_n630_0[1]),.dinb(w_n292_30[0]),.dout(n1960),.clk(gclk));
	jor g1698(.dina(n1960),.dinb(n1959),.dout(n1961),.clk(gclk));
	jand g1699(.dina(w_n429_0[1]),.dinb(w_n267_30[0]),.dout(n1962),.clk(gclk));
	jor g1700(.dina(w_dff_B_UgfuBzO50_0),.dinb(n1961),.dout(n1963),.clk(gclk));
	jor g1701(.dina(n1963),.dinb(w_dff_B_75VVNHvJ2_1),.dout(n1964),.clk(gclk));
	jand g1702(.dina(w_n1964_1[1]),.dinb(w_n364_55[0]),.dout(n1965),.clk(gclk));
	jand g1703(.dina(w_n599_0[1]),.dinb(w_n304_29[2]),.dout(n1966),.clk(gclk));
	jand g1704(.dina(w_n619_0[1]),.dinb(w_n281_29[2]),.dout(n1967),.clk(gclk));
	jand g1705(.dina(w_n609_0[1]),.dinb(w_n267_29[2]),.dout(n1968),.clk(gclk));
	jor g1706(.dina(n1968),.dinb(n1967),.dout(n1969),.clk(gclk));
	jand g1707(.dina(w_n541_0[1]),.dinb(w_n292_29[2]),.dout(n1970),.clk(gclk));
	jor g1708(.dina(w_dff_B_fOzLotLx0_0),.dinb(n1969),.dout(n1971),.clk(gclk));
	jor g1709(.dina(n1971),.dinb(w_dff_B_0KDHoTdV3_1),.dout(n1972),.clk(gclk));
	jand g1710(.dina(w_n1972_1[1]),.dinb(w_n319_55[0]),.dout(n1973),.clk(gclk));
	jand g1711(.dina(w_n530_0[1]),.dinb(w_n304_29[1]),.dout(n1974),.clk(gclk));
	jand g1712(.dina(w_n510_0[1]),.dinb(w_n281_29[1]),.dout(n1975),.clk(gclk));
	jand g1713(.dina(w_n585_0[1]),.dinb(w_n292_29[1]),.dout(n1976),.clk(gclk));
	jor g1714(.dina(n1976),.dinb(n1975),.dout(n1977),.clk(gclk));
	jand g1715(.dina(w_n520_0[1]),.dinb(w_n267_29[1]),.dout(n1978),.clk(gclk));
	jor g1716(.dina(w_dff_B_osWnsPAs4_0),.dinb(n1977),.dout(n1979),.clk(gclk));
	jor g1717(.dina(n1979),.dinb(w_dff_B_HYrPEvnV5_1),.dout(n1980),.clk(gclk));
	jand g1718(.dina(w_n1980_1[1]),.dinb(w_n265_55[0]),.dout(n1981),.clk(gclk));
	jor g1719(.dina(n1981),.dinb(n1973),.dout(n1982),.clk(gclk));
	jand g1720(.dina(w_n554_0[1]),.dinb(w_n304_29[0]),.dout(n1983),.clk(gclk));
	jand g1721(.dina(w_n574_0[1]),.dinb(w_n281_29[0]),.dout(n1984),.clk(gclk));
	jand g1722(.dina(w_n564_0[1]),.dinb(w_n267_29[0]),.dout(n1985),.clk(gclk));
	jor g1723(.dina(n1985),.dinb(n1984),.dout(n1986),.clk(gclk));
	jand g1724(.dina(w_n497_0[1]),.dinb(w_n292_29[0]),.dout(n1987),.clk(gclk));
	jor g1725(.dina(w_dff_B_EyWT0czp2_0),.dinb(n1986),.dout(n1988),.clk(gclk));
	jor g1726(.dina(n1988),.dinb(w_dff_B_vVdaNbcH6_1),.dout(n1989),.clk(gclk));
	jand g1727(.dina(w_n1989_1[1]),.dinb(w_n410_55[0]),.dout(n1990),.clk(gclk));
	jor g1728(.dina(w_dff_B_fhJ1mx9l9_0),.dinb(n1982),.dout(n1991),.clk(gclk));
	jor g1729(.dina(n1991),.dinb(w_dff_B_hOzIDkh54_1),.dout(n1992),.clk(gclk));
	jor g1730(.dina(w_n1992_0[1]),.dinb(w_shift6_59[1]),.dout(n1993),.clk(gclk));
	jand g1731(.dina(n1993),.dinb(n1957),.dout(result12),.clk(gclk));
	jand g1732(.dina(w_n790_0[1]),.dinb(w_n267_28[2]),.dout(n1995),.clk(gclk));
	jand g1733(.dina(w_n780_0[1]),.dinb(w_n281_28[2]),.dout(n1996),.clk(gclk));
	jand g1734(.dina(w_n722_0[1]),.dinb(w_n292_28[2]),.dout(n1997),.clk(gclk));
	jor g1735(.dina(n1997),.dinb(n1996),.dout(n1998),.clk(gclk));
	jand g1736(.dina(w_n800_0[1]),.dinb(w_n304_28[2]),.dout(n1999),.clk(gclk));
	jor g1737(.dina(w_dff_B_0gJiH3OV1_0),.dinb(n1998),.dout(n2000),.clk(gclk));
	jor g1738(.dina(n2000),.dinb(w_dff_B_tbWgCQ7T5_1),.dout(n2001),.clk(gclk));
	jand g1739(.dina(w_n2001_1[1]),.dinb(w_n265_54[2]),.dout(n2002),.clk(gclk));
	jand g1740(.dina(w_n711_0[1]),.dinb(w_n304_28[1]),.dout(n2003),.clk(gclk));
	jand g1741(.dina(w_n691_0[1]),.dinb(w_n281_28[1]),.dout(n2004),.clk(gclk));
	jand g1742(.dina(w_n735_0[1]),.dinb(w_n292_28[1]),.dout(n2005),.clk(gclk));
	jor g1743(.dina(n2005),.dinb(n2004),.dout(n2006),.clk(gclk));
	jand g1744(.dina(w_n701_0[1]),.dinb(w_n267_28[1]),.dout(n2007),.clk(gclk));
	jor g1745(.dina(w_dff_B_M8RJIFvs4_0),.dinb(n2006),.dout(n2008),.clk(gclk));
	jor g1746(.dina(n2008),.dinb(w_dff_B_Z7fK2rF58_1),.dout(n2009),.clk(gclk));
	jand g1747(.dina(w_n2009_1[1]),.dinb(w_n410_54[2]),.dout(n2010),.clk(gclk));
	jand g1748(.dina(w_n847_0[1]),.dinb(w_n304_28[0]),.dout(n2011),.clk(gclk));
	jand g1749(.dina(w_n827_0[1]),.dinb(w_n281_28[0]),.dout(n2012),.clk(gclk));
	jand g1750(.dina(w_n678_0[1]),.dinb(w_n292_28[0]),.dout(n2013),.clk(gclk));
	jor g1751(.dina(n2013),.dinb(n2012),.dout(n2014),.clk(gclk));
	jand g1752(.dina(w_n837_0[1]),.dinb(w_n267_28[0]),.dout(n2015),.clk(gclk));
	jor g1753(.dina(w_dff_B_l2iJDWqD9_0),.dinb(n2014),.dout(n2016),.clk(gclk));
	jor g1754(.dina(n2016),.dinb(w_dff_B_6iCFG5SY4_1),.dout(n2017),.clk(gclk));
	jand g1755(.dina(w_n2017_1[1]),.dinb(w_n364_54[2]),.dout(n2018),.clk(gclk));
	jor g1756(.dina(n2018),.dinb(n2010),.dout(n2019),.clk(gclk));
	jand g1757(.dina(w_n657_0[1]),.dinb(w_n267_27[2]),.dout(n2020),.clk(gclk));
	jand g1758(.dina(w_n667_0[1]),.dinb(w_n281_27[2]),.dout(n2021),.clk(gclk));
	jand g1759(.dina(w_n811_0[1]),.dinb(w_n292_27[2]),.dout(n2022),.clk(gclk));
	jor g1760(.dina(n2022),.dinb(n2021),.dout(n2023),.clk(gclk));
	jand g1761(.dina(w_n647_0[1]),.dinb(w_n304_27[2]),.dout(n2024),.clk(gclk));
	jor g1762(.dina(w_dff_B_Q96lHp3o5_0),.dinb(n2023),.dout(n2025),.clk(gclk));
	jor g1763(.dina(n2025),.dinb(w_dff_B_rD7Jx1Kl7_1),.dout(n2026),.clk(gclk));
	jand g1764(.dina(w_n2026_1[1]),.dinb(w_n319_54[2]),.dout(n2027),.clk(gclk));
	jor g1765(.dina(w_dff_B_SZs8Qcod0_0),.dinb(n2019),.dout(n2028),.clk(gclk));
	jor g1766(.dina(n2028),.dinb(w_dff_B_xuIIATgQ1_1),.dout(n2029),.clk(gclk));
	jor g1767(.dina(w_n2029_0[1]),.dinb(w_n263_59[0]),.dout(n2030),.clk(gclk));
	jand g1768(.dina(w_n935_0[1]),.dinb(w_n304_27[1]),.dout(n2031),.clk(gclk));
	jand g1769(.dina(w_n915_0[1]),.dinb(w_n281_27[1]),.dout(n2032),.clk(gclk));
	jand g1770(.dina(w_n925_0[1]),.dinb(w_n267_27[1]),.dout(n2033),.clk(gclk));
	jor g1771(.dina(n2033),.dinb(n2032),.dout(n2034),.clk(gclk));
	jand g1772(.dina(w_n858_0[1]),.dinb(w_n292_27[1]),.dout(n2035),.clk(gclk));
	jor g1773(.dina(w_dff_B_zURs38kR5_0),.dinb(n2034),.dout(n2036),.clk(gclk));
	jor g1774(.dina(n2036),.dinb(w_dff_B_slVYtXoH6_1),.dout(n2037),.clk(gclk));
	jand g1775(.dina(w_n2037_1[1]),.dinb(w_n410_54[1]),.dout(n2038),.clk(gclk));
	jand g1776(.dina(w_n960_0[1]),.dinb(w_n304_27[0]),.dout(n2039),.clk(gclk));
	jand g1777(.dina(w_n980_0[1]),.dinb(w_n281_27[0]),.dout(n2040),.clk(gclk));
	jand g1778(.dina(w_n902_0[1]),.dinb(w_n292_27[0]),.dout(n2041),.clk(gclk));
	jor g1779(.dina(n2041),.dinb(n2040),.dout(n2042),.clk(gclk));
	jand g1780(.dina(w_n970_0[1]),.dinb(w_n267_27[0]),.dout(n2043),.clk(gclk));
	jor g1781(.dina(w_dff_B_Tg33vzS97_0),.dinb(n2042),.dout(n2044),.clk(gclk));
	jor g1782(.dina(n2044),.dinb(w_dff_B_174ZvsxD2_1),.dout(n2045),.clk(gclk));
	jand g1783(.dina(w_n2045_1[1]),.dinb(w_n319_54[1]),.dout(n2046),.clk(gclk));
	jand g1784(.dina(w_n766_0[1]),.dinb(w_n304_26[2]),.dout(n2047),.clk(gclk));
	jand g1785(.dina(w_n755_0[1]),.dinb(w_n281_26[2]),.dout(n2048),.clk(gclk));
	jand g1786(.dina(w_n991_0[1]),.dinb(w_n292_26[2]),.dout(n2049),.clk(gclk));
	jor g1787(.dina(n2049),.dinb(n2048),.dout(n2050),.clk(gclk));
	jand g1788(.dina(w_n745_0[1]),.dinb(w_n267_26[2]),.dout(n2051),.clk(gclk));
	jor g1789(.dina(w_dff_B_3s6AjRKb2_0),.dinb(n2050),.dout(n2052),.clk(gclk));
	jor g1790(.dina(n2052),.dinb(w_dff_B_VbO6w6zD2_1),.dout(n2053),.clk(gclk));
	jand g1791(.dina(w_n2053_1[1]),.dinb(w_n364_54[1]),.dout(n2054),.clk(gclk));
	jor g1792(.dina(n2054),.dinb(n2046),.dout(n2055),.clk(gclk));
	jand g1793(.dina(w_n881_0[1]),.dinb(w_n267_26[1]),.dout(n2056),.clk(gclk));
	jand g1794(.dina(w_n871_0[1]),.dinb(w_n281_26[1]),.dout(n2057),.clk(gclk));
	jand g1795(.dina(w_n946_0[1]),.dinb(w_n292_26[1]),.dout(n2058),.clk(gclk));
	jor g1796(.dina(n2058),.dinb(n2057),.dout(n2059),.clk(gclk));
	jand g1797(.dina(w_n891_0[1]),.dinb(w_n304_26[1]),.dout(n2060),.clk(gclk));
	jor g1798(.dina(w_dff_B_92yjbt7N5_0),.dinb(n2059),.dout(n2061),.clk(gclk));
	jor g1799(.dina(n2061),.dinb(w_dff_B_h8DUDHPi9_1),.dout(n2062),.clk(gclk));
	jand g1800(.dina(w_n2062_1[1]),.dinb(w_n265_54[1]),.dout(n2063),.clk(gclk));
	jor g1801(.dina(w_dff_B_enD4tXYE6_0),.dinb(n2055),.dout(n2064),.clk(gclk));
	jor g1802(.dina(n2064),.dinb(w_dff_B_KLVuGhgh7_1),.dout(n2065),.clk(gclk));
	jor g1803(.dina(w_n2065_0[1]),.dinb(w_shift6_59[0]),.dout(n2066),.clk(gclk));
	jand g1804(.dina(n2066),.dinb(n2030),.dout(result13),.clk(gclk));
	jand g1805(.dina(w_n1071_0[1]),.dinb(w_n304_26[0]),.dout(n2068),.clk(gclk));
	jand g1806(.dina(w_n1063_0[1]),.dinb(w_n281_26[0]),.dout(n2069),.clk(gclk));
	jand g1807(.dina(w_n1067_0[1]),.dinb(w_n267_26[0]),.dout(n2070),.clk(gclk));
	jor g1808(.dina(n2070),.dinb(n2069),.dout(n2071),.clk(gclk));
	jand g1809(.dina(w_n1015_0[1]),.dinb(w_n292_26[0]),.dout(n2072),.clk(gclk));
	jor g1810(.dina(w_dff_B_Jtue7Ywt4_0),.dinb(n2071),.dout(n2073),.clk(gclk));
	jor g1811(.dina(n2073),.dinb(w_dff_B_ylFxSofU1_1),.dout(n2074),.clk(gclk));
	jand g1812(.dina(w_n2074_1[1]),.dinb(w_n319_54[0]),.dout(n2075),.clk(gclk));
	jand g1813(.dina(w_n1042_0[1]),.dinb(w_n292_25[2]),.dout(n2076),.clk(gclk));
	jand g1814(.dina(w_n1022_0[1]),.dinb(w_n281_25[2]),.dout(n2077),.clk(gclk));
	jand g1815(.dina(w_n1026_0[1]),.dinb(w_n267_25[2]),.dout(n2078),.clk(gclk));
	jor g1816(.dina(n2078),.dinb(n2077),.dout(n2079),.clk(gclk));
	jand g1817(.dina(w_n1030_0[1]),.dinb(w_n304_25[2]),.dout(n2080),.clk(gclk));
	jor g1818(.dina(w_dff_B_b8CiSugl5_0),.dinb(n2079),.dout(n2081),.clk(gclk));
	jor g1819(.dina(n2081),.dinb(w_dff_B_PJjnjmSe8_1),.dout(n2082),.clk(gclk));
	jand g1820(.dina(w_n2082_1[1]),.dinb(w_n410_54[0]),.dout(n2083),.clk(gclk));
	jand g1821(.dina(w_n1086_0[1]),.dinb(w_n304_25[1]),.dout(n2084),.clk(gclk));
	jand g1822(.dina(w_n1094_0[1]),.dinb(w_n281_25[1]),.dout(n2085),.clk(gclk));
	jand g1823(.dina(w_n1076_0[1]),.dinb(w_n292_25[1]),.dout(n2086),.clk(gclk));
	jor g1824(.dina(n2086),.dinb(n2085),.dout(n2087),.clk(gclk));
	jand g1825(.dina(w_n1090_0[1]),.dinb(w_n267_25[1]),.dout(n2088),.clk(gclk));
	jor g1826(.dina(w_dff_B_JGDoXU1T7_0),.dinb(n2087),.dout(n2089),.clk(gclk));
	jor g1827(.dina(n2089),.dinb(w_dff_B_46as8xFJ1_1),.dout(n2090),.clk(gclk));
	jand g1828(.dina(w_n2090_1[1]),.dinb(w_n364_54[0]),.dout(n2091),.clk(gclk));
	jor g1829(.dina(n2091),.dinb(n2083),.dout(n2092),.clk(gclk));
	jand g1830(.dina(w_n1006_0[1]),.dinb(w_n267_25[0]),.dout(n2093),.clk(gclk));
	jand g1831(.dina(w_n1010_0[1]),.dinb(w_n281_25[0]),.dout(n2094),.clk(gclk));
	jand g1832(.dina(w_n1035_0[1]),.dinb(w_n292_25[0]),.dout(n2095),.clk(gclk));
	jor g1833(.dina(n2095),.dinb(n2094),.dout(n2096),.clk(gclk));
	jand g1834(.dina(w_n1002_0[1]),.dinb(w_n304_25[0]),.dout(n2097),.clk(gclk));
	jor g1835(.dina(w_dff_B_fnNiVSQg0_0),.dinb(n2096),.dout(n2098),.clk(gclk));
	jor g1836(.dina(n2098),.dinb(w_dff_B_hk70EXhB4_1),.dout(n2099),.clk(gclk));
	jand g1837(.dina(w_n2099_1[1]),.dinb(w_n265_54[0]),.dout(n2100),.clk(gclk));
	jor g1838(.dina(w_dff_B_Sbji6ZfD0_0),.dinb(n2092),.dout(n2101),.clk(gclk));
	jor g1839(.dina(n2101),.dinb(w_dff_B_UhGdGDuw2_1),.dout(n2102),.clk(gclk));
	jor g1840(.dina(w_n2102_0[1]),.dinb(w_n263_58[2]),.dout(n2103),.clk(gclk));
	jand g1841(.dina(w_n1160_0[1]),.dinb(w_n292_24[2]),.dout(n2104),.clk(gclk));
	jand g1842(.dina(w_n1114_0[1]),.dinb(w_n281_24[2]),.dout(n2105),.clk(gclk));
	jand g1843(.dina(w_n1110_0[1]),.dinb(w_n267_24[2]),.dout(n2106),.clk(gclk));
	jor g1844(.dina(n2106),.dinb(n2105),.dout(n2107),.clk(gclk));
	jand g1845(.dina(w_n1119_0[1]),.dinb(w_n304_24[2]),.dout(n2108),.clk(gclk));
	jor g1846(.dina(w_dff_B_0oY8yfNB8_0),.dinb(n2107),.dout(n2109),.clk(gclk));
	jor g1847(.dina(n2109),.dinb(w_dff_B_FFv3MKX02_1),.dout(n2110),.clk(gclk));
	jand g1848(.dina(w_n2110_1[1]),.dinb(w_n265_53[2]),.dout(n2111),.clk(gclk));
	jand g1849(.dina(w_n1134_0[1]),.dinb(w_n304_24[1]),.dout(n2112),.clk(gclk));
	jand g1850(.dina(w_n1139_0[1]),.dinb(w_n281_24[1]),.dout(n2113),.clk(gclk));
	jand g1851(.dina(w_n1130_0[1]),.dinb(w_n267_24[1]),.dout(n2114),.clk(gclk));
	jor g1852(.dina(n2114),.dinb(n2113),.dout(n2115),.clk(gclk));
	jand g1853(.dina(w_n1106_0[1]),.dinb(w_n292_24[1]),.dout(n2116),.clk(gclk));
	jor g1854(.dina(w_dff_B_tozgo1T96_0),.dinb(n2115),.dout(n2117),.clk(gclk));
	jor g1855(.dina(n2117),.dinb(w_dff_B_pvT9nqua2_1),.dout(n2118),.clk(gclk));
	jand g1856(.dina(w_n2118_1[1]),.dinb(w_n319_53[2]),.dout(n2119),.clk(gclk));
	jand g1857(.dina(w_n1050_0[1]),.dinb(w_n304_24[0]),.dout(n2120),.clk(gclk));
	jand g1858(.dina(w_n1055_0[1]),.dinb(w_n281_24[0]),.dout(n2121),.clk(gclk));
	jand g1859(.dina(w_n1126_0[1]),.dinb(w_n292_24[0]),.dout(n2122),.clk(gclk));
	jor g1860(.dina(n2122),.dinb(n2121),.dout(n2123),.clk(gclk));
	jand g1861(.dina(w_n1046_0[1]),.dinb(w_n267_24[0]),.dout(n2124),.clk(gclk));
	jor g1862(.dina(w_dff_B_rECqHm9H4_0),.dinb(n2123),.dout(n2125),.clk(gclk));
	jor g1863(.dina(n2125),.dinb(w_dff_B_vg76XKpv7_1),.dout(n2126),.clk(gclk));
	jand g1864(.dina(w_n2126_1[1]),.dinb(w_n364_53[2]),.dout(n2127),.clk(gclk));
	jor g1865(.dina(n2127),.dinb(n2119),.dout(n2128),.clk(gclk));
	jand g1866(.dina(w_n1099_0[1]),.dinb(w_n292_23[2]),.dout(n2129),.clk(gclk));
	jand g1867(.dina(w_n1147_0[1]),.dinb(w_n281_23[2]),.dout(n2130),.clk(gclk));
	jand g1868(.dina(w_n1151_0[1]),.dinb(w_n267_23[2]),.dout(n2131),.clk(gclk));
	jor g1869(.dina(n2131),.dinb(n2130),.dout(n2132),.clk(gclk));
	jand g1870(.dina(w_n1155_0[1]),.dinb(w_n304_23[2]),.dout(n2133),.clk(gclk));
	jor g1871(.dina(w_dff_B_PVvmUK9a6_0),.dinb(n2132),.dout(n2134),.clk(gclk));
	jor g1872(.dina(n2134),.dinb(w_dff_B_kx18ekQ99_1),.dout(n2135),.clk(gclk));
	jand g1873(.dina(w_n2135_1[1]),.dinb(w_n410_53[2]),.dout(n2136),.clk(gclk));
	jor g1874(.dina(w_dff_B_OcNBDkyx2_0),.dinb(n2128),.dout(n2137),.clk(gclk));
	jor g1875(.dina(n2137),.dinb(w_dff_B_PRxlyw9O6_1),.dout(n2138),.clk(gclk));
	jor g1876(.dina(w_n2138_0[1]),.dinb(w_shift6_58[2]),.dout(n2139),.clk(gclk));
	jand g1877(.dina(n2139),.dinb(n2103),.dout(result14),.clk(gclk));
	jand g1878(.dina(w_n1175_0[1]),.dinb(w_n267_23[1]),.dout(n2141),.clk(gclk));
	jand g1879(.dina(w_n1171_0[1]),.dinb(w_n281_23[1]),.dout(n2142),.clk(gclk));
	jand g1880(.dina(w_n1245_0[1]),.dinb(w_n292_23[1]),.dout(n2143),.clk(gclk));
	jor g1881(.dina(n2143),.dinb(n2142),.dout(n2144),.clk(gclk));
	jand g1882(.dina(w_n1179_0[1]),.dinb(w_n304_23[1]),.dout(n2145),.clk(gclk));
	jor g1883(.dina(w_dff_B_sFr9dA5r6_0),.dinb(n2144),.dout(n2146),.clk(gclk));
	jor g1884(.dina(n2146),.dinb(w_dff_B_wKhuxg1O7_1),.dout(n2147),.clk(gclk));
	jand g1885(.dina(w_n2147_1[1]),.dinb(w_n319_53[1]),.dout(n2148),.clk(gclk));
	jand g1886(.dina(w_n1204_0[1]),.dinb(w_n304_23[0]),.dout(n2149),.clk(gclk));
	jand g1887(.dina(w_n1199_0[1]),.dinb(w_n281_23[0]),.dout(n2150),.clk(gclk));
	jand g1888(.dina(w_n1211_0[1]),.dinb(w_n292_23[0]),.dout(n2151),.clk(gclk));
	jor g1889(.dina(n2151),.dinb(n2150),.dout(n2152),.clk(gclk));
	jand g1890(.dina(w_n1195_0[1]),.dinb(w_n267_23[0]),.dout(n2153),.clk(gclk));
	jor g1891(.dina(w_dff_B_sdDWXqfe3_0),.dinb(n2152),.dout(n2154),.clk(gclk));
	jor g1892(.dina(n2154),.dinb(w_dff_B_5fVocIcW4_1),.dout(n2155),.clk(gclk));
	jand g1893(.dina(w_n2155_1[1]),.dinb(w_n410_53[1]),.dout(n2156),.clk(gclk));
	jand g1894(.dina(w_n1236_0[1]),.dinb(w_n267_22[2]),.dout(n2157),.clk(gclk));
	jand g1895(.dina(w_n1232_0[1]),.dinb(w_n281_22[2]),.dout(n2158),.clk(gclk));
	jand g1896(.dina(w_n1191_0[1]),.dinb(w_n292_22[2]),.dout(n2159),.clk(gclk));
	jor g1897(.dina(n2159),.dinb(n2158),.dout(n2160),.clk(gclk));
	jand g1898(.dina(w_n1240_0[1]),.dinb(w_n304_22[2]),.dout(n2161),.clk(gclk));
	jor g1899(.dina(w_dff_B_TnrR4rFy8_0),.dinb(n2160),.dout(n2162),.clk(gclk));
	jor g1900(.dina(n2162),.dinb(w_dff_B_uSl1DoMb4_1),.dout(n2163),.clk(gclk));
	jand g1901(.dina(w_n2163_1[1]),.dinb(w_n265_53[1]),.dout(n2164),.clk(gclk));
	jor g1902(.dina(n2164),.dinb(n2156),.dout(n2165),.clk(gclk));
	jand g1903(.dina(w_n1184_0[1]),.dinb(w_n292_22[1]),.dout(n2166),.clk(gclk));
	jand g1904(.dina(w_n1288_0[1]),.dinb(w_n281_22[1]),.dout(n2167),.clk(gclk));
	jand g1905(.dina(w_n1279_0[1]),.dinb(w_n267_22[1]),.dout(n2168),.clk(gclk));
	jor g1906(.dina(n2168),.dinb(n2167),.dout(n2169),.clk(gclk));
	jand g1907(.dina(w_n1283_0[1]),.dinb(w_n304_22[1]),.dout(n2170),.clk(gclk));
	jor g1908(.dina(w_dff_B_yFXClqjf2_0),.dinb(n2169),.dout(n2171),.clk(gclk));
	jor g1909(.dina(n2171),.dinb(w_dff_B_3n3bcFZF0_1),.dout(n2172),.clk(gclk));
	jand g1910(.dina(w_n2172_1[1]),.dinb(w_n364_53[1]),.dout(n2173),.clk(gclk));
	jor g1911(.dina(w_dff_B_o8z0a3BH8_0),.dinb(n2165),.dout(n2174),.clk(gclk));
	jor g1912(.dina(n2174),.dinb(w_dff_B_qCuGtxRb1_1),.dout(n2175),.clk(gclk));
	jor g1913(.dina(w_n2175_0[1]),.dinb(w_n263_58[1]),.dout(n2176),.clk(gclk));
	jand g1914(.dina(w_n1219_0[1]),.dinb(w_n304_22[0]),.dout(n2177),.clk(gclk));
	jand g1915(.dina(w_n1224_0[1]),.dinb(w_n281_22[0]),.dout(n2178),.clk(gclk));
	jand g1916(.dina(w_n1308_0[1]),.dinb(w_n292_22[0]),.dout(n2179),.clk(gclk));
	jor g1917(.dina(n2179),.dinb(n2178),.dout(n2180),.clk(gclk));
	jand g1918(.dina(w_n1215_0[1]),.dinb(w_n267_22[0]),.dout(n2181),.clk(gclk));
	jor g1919(.dina(w_dff_B_Ewoal9ki5_0),.dinb(n2180),.dout(n2182),.clk(gclk));
	jor g1920(.dina(n2182),.dinb(w_dff_B_871fhSZh8_1),.dout(n2183),.clk(gclk));
	jand g1921(.dina(w_n2183_1[1]),.dinb(w_n364_53[0]),.dout(n2184),.clk(gclk));
	jand g1922(.dina(w_n1303_0[1]),.dinb(w_n304_21[2]),.dout(n2185),.clk(gclk));
	jand g1923(.dina(w_n1295_0[1]),.dinb(w_n281_21[2]),.dout(n2186),.clk(gclk));
	jand g1924(.dina(w_n1299_0[1]),.dinb(w_n267_21[2]),.dout(n2187),.clk(gclk));
	jor g1925(.dina(n2187),.dinb(n2186),.dout(n2188),.clk(gclk));
	jand g1926(.dina(w_n1255_0[1]),.dinb(w_n292_21[2]),.dout(n2189),.clk(gclk));
	jor g1927(.dina(w_dff_B_bqhhQYEO8_0),.dinb(n2188),.dout(n2190),.clk(gclk));
	jor g1928(.dina(n2190),.dinb(w_dff_B_DlowA4MC0_1),.dout(n2191),.clk(gclk));
	jand g1929(.dina(w_n2191_1[1]),.dinb(w_n319_53[0]),.dout(n2192),.clk(gclk));
	jand g1930(.dina(w_n1263_0[1]),.dinb(w_n304_21[1]),.dout(n2193),.clk(gclk));
	jand g1931(.dina(w_n1268_0[1]),.dinb(w_n281_21[1]),.dout(n2194),.clk(gclk));
	jand g1932(.dina(w_n1259_0[1]),.dinb(w_n267_21[1]),.dout(n2195),.clk(gclk));
	jor g1933(.dina(n2195),.dinb(n2194),.dout(n2196),.clk(gclk));
	jand g1934(.dina(w_n1316_0[1]),.dinb(w_n292_21[1]),.dout(n2197),.clk(gclk));
	jor g1935(.dina(w_dff_B_5qLGuZg58_0),.dinb(n2196),.dout(n2198),.clk(gclk));
	jor g1936(.dina(n2198),.dinb(w_dff_B_zacrjjWS4_1),.dout(n2199),.clk(gclk));
	jand g1937(.dina(w_n2199_1[1]),.dinb(w_n265_53[0]),.dout(n2200),.clk(gclk));
	jor g1938(.dina(n2200),.dinb(n2192),.dout(n2201),.clk(gclk));
	jand g1939(.dina(w_n1320_0[1]),.dinb(w_n267_21[0]),.dout(n2202),.clk(gclk));
	jand g1940(.dina(w_n1329_0[1]),.dinb(w_n281_21[0]),.dout(n2203),.clk(gclk));
	jand g1941(.dina(w_n1275_0[1]),.dinb(w_n292_21[0]),.dout(n2204),.clk(gclk));
	jor g1942(.dina(n2204),.dinb(n2203),.dout(n2205),.clk(gclk));
	jand g1943(.dina(w_n1324_0[1]),.dinb(w_n304_21[0]),.dout(n2206),.clk(gclk));
	jor g1944(.dina(w_dff_B_QlNfdnSh4_0),.dinb(n2205),.dout(n2207),.clk(gclk));
	jor g1945(.dina(n2207),.dinb(w_dff_B_rUo3KNte8_1),.dout(n2208),.clk(gclk));
	jand g1946(.dina(w_n2208_1[1]),.dinb(w_n410_53[0]),.dout(n2209),.clk(gclk));
	jor g1947(.dina(w_dff_B_IfHCHb0m5_0),.dinb(n2201),.dout(n2210),.clk(gclk));
	jor g1948(.dina(n2210),.dinb(w_dff_B_ipvPNgWN6_1),.dout(n2211),.clk(gclk));
	jor g1949(.dina(w_n2211_0[1]),.dinb(w_shift6_58[1]),.dout(n2212),.clk(gclk));
	jand g1950(.dina(n2212),.dinb(n2176),.dout(result15),.clk(gclk));
	jand g1951(.dina(w_n407_1[0]),.dinb(w_n319_52[2]),.dout(n2214),.clk(gclk));
	jand g1952(.dina(w_n362_1[0]),.dinb(w_n265_52[2]),.dout(n2215),.clk(gclk));
	jand g1953(.dina(w_n410_52[2]),.dinb(w_n316_1[0]),.dout(n2216),.clk(gclk));
	jor g1954(.dina(n2216),.dinb(n2215),.dout(n2217),.clk(gclk));
	jand g1955(.dina(w_n500_1[0]),.dinb(w_n364_52[2]),.dout(n2218),.clk(gclk));
	jor g1956(.dina(w_dff_B_BoPmVl8N6_0),.dinb(n2217),.dout(n2219),.clk(gclk));
	jor g1957(.dina(n2219),.dinb(w_dff_B_1rfsyViv6_1),.dout(n2220),.clk(gclk));
	jor g1958(.dina(w_n2220_0[1]),.dinb(w_n263_58[0]),.dout(n2221),.clk(gclk));
	jand g1959(.dina(w_n588_1[0]),.dinb(w_n410_52[1]),.dout(n2222),.clk(gclk));
	jand g1960(.dina(w_n633_1[0]),.dinb(w_n319_52[1]),.dout(n2223),.clk(gclk));
	jand g1961(.dina(w_n544_1[0]),.dinb(w_n265_52[1]),.dout(n2224),.clk(gclk));
	jor g1962(.dina(n2224),.dinb(n2223),.dout(n2225),.clk(gclk));
	jand g1963(.dina(w_n453_1[0]),.dinb(w_n364_52[1]),.dout(n2226),.clk(gclk));
	jor g1964(.dina(w_dff_B_8LcbiD876_0),.dinb(n2225),.dout(n2227),.clk(gclk));
	jor g1965(.dina(n2227),.dinb(w_dff_B_ShHJJsvM6_1),.dout(n2228),.clk(gclk));
	jor g1966(.dina(w_n2228_0[1]),.dinb(w_shift6_58[0]),.dout(n2229),.clk(gclk));
	jand g1967(.dina(n2229),.dinb(n2221),.dout(result16),.clk(gclk));
	jand g1968(.dina(w_n814_1[0]),.dinb(w_n265_52[0]),.dout(n2231),.clk(gclk));
	jand g1969(.dina(w_n725_1[0]),.dinb(w_n410_52[0]),.dout(n2232),.clk(gclk));
	jand g1970(.dina(w_n861_1[0]),.dinb(w_n364_52[0]),.dout(n2233),.clk(gclk));
	jor g1971(.dina(n2233),.dinb(n2232),.dout(n2234),.clk(gclk));
	jand g1972(.dina(w_n681_1[0]),.dinb(w_n319_52[0]),.dout(n2235),.clk(gclk));
	jor g1973(.dina(w_dff_B_ZV0RQbIM7_0),.dinb(n2234),.dout(n2236),.clk(gclk));
	jor g1974(.dina(n2236),.dinb(w_dff_B_H5LQYE1i4_1),.dout(n2237),.clk(gclk));
	jor g1975(.dina(w_n2237_0[1]),.dinb(w_n263_57[2]),.dout(n2238),.clk(gclk));
	jand g1976(.dina(w_n769_1[0]),.dinb(w_n364_51[2]),.dout(n2239),.clk(gclk));
	jand g1977(.dina(w_n994_1[0]),.dinb(w_n319_51[2]),.dout(n2240),.clk(gclk));
	jand g1978(.dina(w_n905_1[0]),.dinb(w_n265_51[2]),.dout(n2241),.clk(gclk));
	jor g1979(.dina(n2241),.dinb(n2240),.dout(n2242),.clk(gclk));
	jand g1980(.dina(w_n949_1[0]),.dinb(w_n410_51[2]),.dout(n2243),.clk(gclk));
	jor g1981(.dina(w_dff_B_WKMYwIeP6_0),.dinb(n2242),.dout(n2244),.clk(gclk));
	jor g1982(.dina(n2244),.dinb(w_dff_B_DNWcCaNq6_1),.dout(n2245),.clk(gclk));
	jor g1983(.dina(w_n2245_0[1]),.dinb(w_shift6_57[2]),.dout(n2246),.clk(gclk));
	jand g1984(.dina(n2246),.dinb(n2238),.dout(result17),.clk(gclk));
	jand g1985(.dina(w_n1102_1[0]),.dinb(w_n364_51[1]),.dout(n2248),.clk(gclk));
	jand g1986(.dina(w_n1038_1[0]),.dinb(w_n410_51[1]),.dout(n2249),.clk(gclk));
	jand g1987(.dina(w_n1018_1[0]),.dinb(w_n265_51[1]),.dout(n2250),.clk(gclk));
	jor g1988(.dina(n2250),.dinb(n2249),.dout(n2251),.clk(gclk));
	jand g1989(.dina(w_n1079_1[0]),.dinb(w_n319_51[1]),.dout(n2252),.clk(gclk));
	jor g1990(.dina(w_dff_B_wQeft8uk8_0),.dinb(n2251),.dout(n2253),.clk(gclk));
	jor g1991(.dina(n2253),.dinb(w_dff_B_wMTGnKcB8_1),.dout(n2254),.clk(gclk));
	jor g1992(.dina(w_n2254_0[1]),.dinb(w_n263_57[1]),.dout(n2255),.clk(gclk));
	jand g1993(.dina(w_n1058_1[0]),.dinb(w_n364_51[0]),.dout(n2256),.clk(gclk));
	jand g1994(.dina(w_n1142_1[0]),.dinb(w_n319_51[0]),.dout(n2257),.clk(gclk));
	jand g1995(.dina(w_n1122_1[0]),.dinb(w_n265_51[0]),.dout(n2258),.clk(gclk));
	jor g1996(.dina(n2258),.dinb(n2257),.dout(n2259),.clk(gclk));
	jand g1997(.dina(w_n1163_1[0]),.dinb(w_n410_51[0]),.dout(n2260),.clk(gclk));
	jor g1998(.dina(w_dff_B_nGRQaI5L2_0),.dinb(n2259),.dout(n2261),.clk(gclk));
	jor g1999(.dina(n2261),.dinb(w_dff_B_reajkNSh8_1),.dout(n2262),.clk(gclk));
	jor g2000(.dina(w_n2262_0[1]),.dinb(w_shift6_57[1]),.dout(n2263),.clk(gclk));
	jand g2001(.dina(n2263),.dinb(n2255),.dout(result18),.clk(gclk));
	jand g2002(.dina(w_n1187_1[0]),.dinb(w_n319_50[2]),.dout(n2265),.clk(gclk));
	jand g2003(.dina(w_n1248_1[0]),.dinb(w_n265_50[2]),.dout(n2266),.clk(gclk));
	jand g2004(.dina(w_n1207_1[0]),.dinb(w_n410_50[2]),.dout(n2267),.clk(gclk));
	jor g2005(.dina(n2267),.dinb(n2266),.dout(n2268),.clk(gclk));
	jand g2006(.dina(w_n1291_1[0]),.dinb(w_n364_50[2]),.dout(n2269),.clk(gclk));
	jor g2007(.dina(w_dff_B_bAkFKoGi1_0),.dinb(n2268),.dout(n2270),.clk(gclk));
	jor g2008(.dina(n2270),.dinb(w_dff_B_vqYPtKNk8_1),.dout(n2271),.clk(gclk));
	jor g2009(.dina(w_n2271_0[1]),.dinb(w_n263_57[0]),.dout(n2272),.clk(gclk));
	jand g2010(.dina(w_n1271_1[0]),.dinb(w_n265_50[1]),.dout(n2273),.clk(gclk));
	jand g2011(.dina(w_n1227_1[0]),.dinb(w_n364_50[1]),.dout(n2274),.clk(gclk));
	jand g2012(.dina(w_n1311_1[0]),.dinb(w_n319_50[1]),.dout(n2275),.clk(gclk));
	jor g2013(.dina(n2275),.dinb(n2274),.dout(n2276),.clk(gclk));
	jand g2014(.dina(w_n1332_1[0]),.dinb(w_n410_50[1]),.dout(n2277),.clk(gclk));
	jor g2015(.dina(w_dff_B_bvqaMLGq4_0),.dinb(n2276),.dout(n2278),.clk(gclk));
	jor g2016(.dina(n2278),.dinb(w_dff_B_QbZh5GTu1_1),.dout(n2279),.clk(gclk));
	jor g2017(.dina(w_n2279_0[1]),.dinb(w_shift6_57[0]),.dout(n2280),.clk(gclk));
	jand g2018(.dina(n2280),.dinb(n2272),.dout(result19),.clk(gclk));
	jand g2019(.dina(w_n1405_1[0]),.dinb(w_n364_50[0]),.dout(n2282),.clk(gclk));
	jand g2020(.dina(w_n1344_1[0]),.dinb(w_n319_50[0]),.dout(n2283),.clk(gclk));
	jand g2021(.dina(w_n1360_1[0]),.dinb(w_n410_50[0]),.dout(n2284),.clk(gclk));
	jor g2022(.dina(n2284),.dinb(n2283),.dout(n2285),.clk(gclk));
	jand g2023(.dina(w_n1369_1[0]),.dinb(w_n265_50[0]),.dout(n2286),.clk(gclk));
	jor g2024(.dina(w_dff_B_CzywkDtF3_0),.dinb(n2285),.dout(n2287),.clk(gclk));
	jor g2025(.dina(n2287),.dinb(w_dff_B_aJJeIIHt4_1),.dout(n2288),.clk(gclk));
	jor g2026(.dina(w_n2288_0[1]),.dinb(w_n263_56[2]),.dout(n2289),.clk(gclk));
	jand g2027(.dina(w_n1380_1[0]),.dinb(w_n410_49[2]),.dout(n2290),.clk(gclk));
	jand g2028(.dina(w_n1396_1[0]),.dinb(w_n319_49[2]),.dout(n2291),.clk(gclk));
	jand g2029(.dina(w_n1388_1[0]),.dinb(w_n265_49[2]),.dout(n2292),.clk(gclk));
	jor g2030(.dina(n2292),.dinb(n2291),.dout(n2293),.clk(gclk));
	jand g2031(.dina(w_n1352_1[0]),.dinb(w_n364_49[2]),.dout(n2294),.clk(gclk));
	jor g2032(.dina(w_dff_B_YX9OTQX74_0),.dinb(n2293),.dout(n2295),.clk(gclk));
	jor g2033(.dina(n2295),.dinb(w_dff_B_VTYfoZ241_1),.dout(n2296),.clk(gclk));
	jor g2034(.dina(w_n2296_0[1]),.dinb(w_shift6_56[2]),.dout(n2297),.clk(gclk));
	jand g2035(.dina(n2297),.dinb(n2289),.dout(result20),.clk(gclk));
	jand g2036(.dina(w_n1417_1[0]),.dinb(w_n265_49[1]),.dout(n2299),.clk(gclk));
	jand g2037(.dina(w_n1442_1[0]),.dinb(w_n319_49[1]),.dout(n2300),.clk(gclk));
	jand g2038(.dina(w_n1433_1[0]),.dinb(w_n410_49[1]),.dout(n2301),.clk(gclk));
	jor g2039(.dina(n2301),.dinb(n2300),.dout(n2302),.clk(gclk));
	jand g2040(.dina(w_n1453_1[0]),.dinb(w_n364_49[1]),.dout(n2303),.clk(gclk));
	jor g2041(.dina(w_dff_B_rl1ZH6TR5_0),.dinb(n2302),.dout(n2304),.clk(gclk));
	jor g2042(.dina(n2304),.dinb(w_dff_B_hCssqM0Q9_1),.dout(n2305),.clk(gclk));
	jor g2043(.dina(w_n2305_0[1]),.dinb(w_n263_56[1]),.dout(n2306),.clk(gclk));
	jand g2044(.dina(w_n1469_1[0]),.dinb(w_n410_49[0]),.dout(n2307),.clk(gclk));
	jand g2045(.dina(w_n1478_1[0]),.dinb(w_n319_49[0]),.dout(n2308),.clk(gclk));
	jand g2046(.dina(w_n1425_1[0]),.dinb(w_n364_49[0]),.dout(n2309),.clk(gclk));
	jor g2047(.dina(n2309),.dinb(n2308),.dout(n2310),.clk(gclk));
	jand g2048(.dina(w_n1461_1[0]),.dinb(w_n265_49[0]),.dout(n2311),.clk(gclk));
	jor g2049(.dina(w_dff_B_dV3x719y6_0),.dinb(n2310),.dout(n2312),.clk(gclk));
	jor g2050(.dina(n2312),.dinb(w_dff_B_qJOt6bhg1_1),.dout(n2313),.clk(gclk));
	jor g2051(.dina(w_n2313_0[1]),.dinb(w_shift6_56[1]),.dout(n2314),.clk(gclk));
	jand g2052(.dina(n2314),.dinb(n2306),.dout(result21),.clk(gclk));
	jand g2053(.dina(w_n1515_1[0]),.dinb(w_n265_48[2]),.dout(n2316),.clk(gclk));
	jand g2054(.dina(w_n1506_1[0]),.dinb(w_n319_48[2]),.dout(n2317),.clk(gclk));
	jand g2055(.dina(w_n1490_1[0]),.dinb(w_n410_48[2]),.dout(n2318),.clk(gclk));
	jor g2056(.dina(n2318),.dinb(n2317),.dout(n2319),.clk(gclk));
	jand g2057(.dina(w_n1526_1[0]),.dinb(w_n364_48[2]),.dout(n2320),.clk(gclk));
	jor g2058(.dina(w_dff_B_Oi4X5sPK9_0),.dinb(n2319),.dout(n2321),.clk(gclk));
	jor g2059(.dina(n2321),.dinb(w_dff_B_G4Ih9Qr33_1),.dout(n2322),.clk(gclk));
	jor g2060(.dina(w_n2322_0[1]),.dinb(w_n263_56[0]),.dout(n2323),.clk(gclk));
	jand g2061(.dina(w_n1551_1[0]),.dinb(w_n410_48[1]),.dout(n2324),.clk(gclk));
	jand g2062(.dina(w_n1542_1[0]),.dinb(w_n319_48[1]),.dout(n2325),.clk(gclk));
	jand g2063(.dina(w_n1534_1[0]),.dinb(w_n265_48[1]),.dout(n2326),.clk(gclk));
	jor g2064(.dina(n2326),.dinb(n2325),.dout(n2327),.clk(gclk));
	jand g2065(.dina(w_n1498_1[0]),.dinb(w_n364_48[1]),.dout(n2328),.clk(gclk));
	jor g2066(.dina(w_dff_B_bc3S7ENI2_0),.dinb(n2327),.dout(n2329),.clk(gclk));
	jor g2067(.dina(n2329),.dinb(w_dff_B_UQHrQaep4_1),.dout(n2330),.clk(gclk));
	jor g2068(.dina(w_n2330_0[1]),.dinb(w_shift6_56[0]),.dout(n2331),.clk(gclk));
	jand g2069(.dina(n2331),.dinb(n2323),.dout(result22),.clk(gclk));
	jand g2070(.dina(w_n1588_1[0]),.dinb(w_n265_48[0]),.dout(n2333),.clk(gclk));
	jand g2071(.dina(w_n1599_1[0]),.dinb(w_n364_48[0]),.dout(n2334),.clk(gclk));
	jand g2072(.dina(w_n1579_1[0]),.dinb(w_n319_48[0]),.dout(n2335),.clk(gclk));
	jor g2073(.dina(n2335),.dinb(n2334),.dout(n2336),.clk(gclk));
	jand g2074(.dina(w_n1563_1[0]),.dinb(w_n410_48[0]),.dout(n2337),.clk(gclk));
	jor g2075(.dina(w_dff_B_wTfreXba5_0),.dinb(n2336),.dout(n2338),.clk(gclk));
	jor g2076(.dina(n2338),.dinb(w_dff_B_7yGKMDYQ1_1),.dout(n2339),.clk(gclk));
	jor g2077(.dina(w_n2339_0[1]),.dinb(w_n263_55[2]),.dout(n2340),.clk(gclk));
	jand g2078(.dina(w_n1615_1[0]),.dinb(w_n410_47[2]),.dout(n2341),.clk(gclk));
	jand g2079(.dina(w_n1607_1[0]),.dinb(w_n265_47[2]),.dout(n2342),.clk(gclk));
	jand g2080(.dina(w_n1624_1[0]),.dinb(w_n319_47[2]),.dout(n2343),.clk(gclk));
	jor g2081(.dina(n2343),.dinb(n2342),.dout(n2344),.clk(gclk));
	jand g2082(.dina(w_n1571_1[0]),.dinb(w_n364_47[2]),.dout(n2345),.clk(gclk));
	jor g2083(.dina(w_dff_B_Xvu7oEBw8_0),.dinb(n2344),.dout(n2346),.clk(gclk));
	jor g2084(.dina(n2346),.dinb(w_dff_B_xTJkLHWE4_1),.dout(n2347),.clk(gclk));
	jor g2085(.dina(w_n2347_0[1]),.dinb(w_shift6_55[2]),.dout(n2348),.clk(gclk));
	jand g2086(.dina(n2348),.dinb(n2340),.dout(result23),.clk(gclk));
	jand g2087(.dina(w_n1661_1[0]),.dinb(w_n265_47[1]),.dout(n2350),.clk(gclk));
	jand g2088(.dina(w_n1672_1[0]),.dinb(w_n364_47[1]),.dout(n2351),.clk(gclk));
	jand g2089(.dina(w_n1652_1[0]),.dinb(w_n319_47[1]),.dout(n2352),.clk(gclk));
	jor g2090(.dina(n2352),.dinb(n2351),.dout(n2353),.clk(gclk));
	jand g2091(.dina(w_n1636_1[0]),.dinb(w_n410_47[1]),.dout(n2354),.clk(gclk));
	jor g2092(.dina(w_dff_B_Bh0cWlsK3_0),.dinb(n2353),.dout(n2355),.clk(gclk));
	jor g2093(.dina(n2355),.dinb(w_dff_B_WHlDTliR9_1),.dout(n2356),.clk(gclk));
	jor g2094(.dina(w_n2356_0[1]),.dinb(w_n263_55[1]),.dout(n2357),.clk(gclk));
	jand g2095(.dina(w_n1688_1[0]),.dinb(w_n319_47[0]),.dout(n2358),.clk(gclk));
	jand g2096(.dina(w_n1680_1[0]),.dinb(w_n265_47[0]),.dout(n2359),.clk(gclk));
	jand g2097(.dina(w_n1644_1[0]),.dinb(w_n364_47[0]),.dout(n2360),.clk(gclk));
	jor g2098(.dina(n2360),.dinb(n2359),.dout(n2361),.clk(gclk));
	jand g2099(.dina(w_n1697_1[0]),.dinb(w_n410_47[0]),.dout(n2362),.clk(gclk));
	jor g2100(.dina(w_dff_B_0uemW6GM9_0),.dinb(n2361),.dout(n2363),.clk(gclk));
	jor g2101(.dina(n2363),.dinb(w_dff_B_2kENvoBC8_1),.dout(n2364),.clk(gclk));
	jor g2102(.dina(w_n2364_0[1]),.dinb(w_shift6_55[1]),.dout(n2365),.clk(gclk));
	jand g2103(.dina(n2365),.dinb(n2357),.dout(result24),.clk(gclk));
	jand g2104(.dina(w_n1725_1[0]),.dinb(w_n410_46[2]),.dout(n2367),.clk(gclk));
	jand g2105(.dina(w_n1770_1[0]),.dinb(w_n364_46[2]),.dout(n2368),.clk(gclk));
	jand g2106(.dina(w_n1709_1[0]),.dinb(w_n319_46[2]),.dout(n2369),.clk(gclk));
	jor g2107(.dina(n2369),.dinb(n2368),.dout(n2370),.clk(gclk));
	jand g2108(.dina(w_n1734_1[0]),.dinb(w_n265_46[2]),.dout(n2371),.clk(gclk));
	jor g2109(.dina(w_dff_B_GNedNEEq9_0),.dinb(n2370),.dout(n2372),.clk(gclk));
	jor g2110(.dina(n2372),.dinb(w_dff_B_8SRP66dE1_1),.dout(n2373),.clk(gclk));
	jor g2111(.dina(w_n2373_0[1]),.dinb(w_n263_55[0]),.dout(n2374),.clk(gclk));
	jand g2112(.dina(w_n1761_1[0]),.dinb(w_n319_46[1]),.dout(n2375),.clk(gclk));
	jand g2113(.dina(w_n1753_1[0]),.dinb(w_n265_46[1]),.dout(n2376),.clk(gclk));
	jand g2114(.dina(w_n1717_1[0]),.dinb(w_n364_46[1]),.dout(n2377),.clk(gclk));
	jor g2115(.dina(n2377),.dinb(n2376),.dout(n2378),.clk(gclk));
	jand g2116(.dina(w_n1745_1[0]),.dinb(w_n410_46[1]),.dout(n2379),.clk(gclk));
	jor g2117(.dina(w_dff_B_McwzmPqr1_0),.dinb(n2378),.dout(n2380),.clk(gclk));
	jor g2118(.dina(n2380),.dinb(w_dff_B_eD6zHKXZ0_1),.dout(n2381),.clk(gclk));
	jor g2119(.dina(w_n2381_0[1]),.dinb(w_shift6_55[0]),.dout(n2382),.clk(gclk));
	jand g2120(.dina(n2382),.dinb(n2374),.dout(result25),.clk(gclk));
	jand g2121(.dina(w_n1807_1[0]),.dinb(w_n319_46[0]),.dout(n2384),.clk(gclk));
	jand g2122(.dina(w_n1843_1[0]),.dinb(w_n364_46[0]),.dout(n2385),.clk(gclk));
	jand g2123(.dina(w_n1798_1[0]),.dinb(w_n410_46[0]),.dout(n2386),.clk(gclk));
	jor g2124(.dina(n2386),.dinb(n2385),.dout(n2387),.clk(gclk));
	jand g2125(.dina(w_n1782_1[0]),.dinb(w_n265_46[0]),.dout(n2388),.clk(gclk));
	jor g2126(.dina(w_dff_B_u47osZBz0_0),.dinb(n2387),.dout(n2389),.clk(gclk));
	jor g2127(.dina(n2389),.dinb(w_dff_B_h3eJu9OU0_1),.dout(n2390),.clk(gclk));
	jor g2128(.dina(w_n2390_0[1]),.dinb(w_n263_54[2]),.dout(n2391),.clk(gclk));
	jand g2129(.dina(w_n1834_1[0]),.dinb(w_n410_45[2]),.dout(n2392),.clk(gclk));
	jand g2130(.dina(w_n1818_1[0]),.dinb(w_n319_45[2]),.dout(n2393),.clk(gclk));
	jand g2131(.dina(w_n1826_1[0]),.dinb(w_n265_45[2]),.dout(n2394),.clk(gclk));
	jor g2132(.dina(n2394),.dinb(n2393),.dout(n2395),.clk(gclk));
	jand g2133(.dina(w_n1790_1[0]),.dinb(w_n364_45[2]),.dout(n2396),.clk(gclk));
	jor g2134(.dina(w_dff_B_oYfAcDzV7_0),.dinb(n2395),.dout(n2397),.clk(gclk));
	jor g2135(.dina(n2397),.dinb(w_dff_B_ywtVITPN8_1),.dout(n2398),.clk(gclk));
	jor g2136(.dina(w_n2398_0[1]),.dinb(w_shift6_54[2]),.dout(n2399),.clk(gclk));
	jand g2137(.dina(n2399),.dinb(n2391),.dout(result26),.clk(gclk));
	jand g2138(.dina(w_n1855_1[0]),.dinb(w_n265_45[1]),.dout(n2401),.clk(gclk));
	jand g2139(.dina(w_n1891_1[0]),.dinb(w_n364_45[1]),.dout(n2402),.clk(gclk));
	jand g2140(.dina(w_n1871_1[0]),.dinb(w_n410_45[1]),.dout(n2403),.clk(gclk));
	jor g2141(.dina(n2403),.dinb(n2402),.dout(n2404),.clk(gclk));
	jand g2142(.dina(w_n1880_1[0]),.dinb(w_n319_45[1]),.dout(n2405),.clk(gclk));
	jor g2143(.dina(w_dff_B_rGaC2c9d4_0),.dinb(n2404),.dout(n2406),.clk(gclk));
	jor g2144(.dina(n2406),.dinb(w_dff_B_otiiGruG4_1),.dout(n2407),.clk(gclk));
	jor g2145(.dina(w_n2407_0[1]),.dinb(w_n263_54[1]),.dout(n2408),.clk(gclk));
	jand g2146(.dina(w_n1907_1[0]),.dinb(w_n410_45[0]),.dout(n2409),.clk(gclk));
	jand g2147(.dina(w_n1916_1[0]),.dinb(w_n319_45[0]),.dout(n2410),.clk(gclk));
	jand g2148(.dina(w_n1899_1[0]),.dinb(w_n265_45[0]),.dout(n2411),.clk(gclk));
	jor g2149(.dina(n2411),.dinb(n2410),.dout(n2412),.clk(gclk));
	jand g2150(.dina(w_n1863_1[0]),.dinb(w_n364_45[0]),.dout(n2413),.clk(gclk));
	jor g2151(.dina(w_dff_B_SqgF1FXp2_0),.dinb(n2412),.dout(n2414),.clk(gclk));
	jor g2152(.dina(n2414),.dinb(w_dff_B_6L9GTXRb7_1),.dout(n2415),.clk(gclk));
	jor g2153(.dina(w_n2415_0[1]),.dinb(w_shift6_54[1]),.dout(n2416),.clk(gclk));
	jand g2154(.dina(n2416),.dinb(n2408),.dout(result27),.clk(gclk));
	jand g2155(.dina(w_n1953_1[0]),.dinb(w_n265_44[2]),.dout(n2418),.clk(gclk));
	jand g2156(.dina(w_n1989_1[0]),.dinb(w_n364_44[2]),.dout(n2419),.clk(gclk));
	jand g2157(.dina(w_n1944_1[0]),.dinb(w_n319_44[2]),.dout(n2420),.clk(gclk));
	jor g2158(.dina(n2420),.dinb(n2419),.dout(n2421),.clk(gclk));
	jand g2159(.dina(w_n1928_1[0]),.dinb(w_n410_44[2]),.dout(n2422),.clk(gclk));
	jor g2160(.dina(w_dff_B_rkzRbhOh1_0),.dinb(n2421),.dout(n2423),.clk(gclk));
	jor g2161(.dina(n2423),.dinb(w_dff_B_uHPHRthA7_1),.dout(n2424),.clk(gclk));
	jor g2162(.dina(w_n2424_0[1]),.dinb(w_n263_54[0]),.dout(n2425),.clk(gclk));
	jand g2163(.dina(w_n1972_1[0]),.dinb(w_n265_44[1]),.dout(n2426),.clk(gclk));
	jand g2164(.dina(w_n1964_1[0]),.dinb(w_n319_44[1]),.dout(n2427),.clk(gclk));
	jand g2165(.dina(w_n1936_1[0]),.dinb(w_n364_44[1]),.dout(n2428),.clk(gclk));
	jor g2166(.dina(n2428),.dinb(n2427),.dout(n2429),.clk(gclk));
	jand g2167(.dina(w_n1980_1[0]),.dinb(w_n410_44[1]),.dout(n2430),.clk(gclk));
	jor g2168(.dina(w_dff_B_dk5lNsOw9_0),.dinb(n2429),.dout(n2431),.clk(gclk));
	jor g2169(.dina(n2431),.dinb(w_dff_B_99mKSXMI6_1),.dout(n2432),.clk(gclk));
	jor g2170(.dina(w_n2432_0[1]),.dinb(w_shift6_54[0]),.dout(n2433),.clk(gclk));
	jand g2171(.dina(n2433),.dinb(n2425),.dout(result28),.clk(gclk));
	jand g2172(.dina(w_n2017_1[0]),.dinb(w_n319_44[0]),.dout(n2435),.clk(gclk));
	jand g2173(.dina(w_n2037_1[0]),.dinb(w_n364_44[0]),.dout(n2436),.clk(gclk));
	jand g2174(.dina(w_n2001_1[0]),.dinb(w_n410_44[0]),.dout(n2437),.clk(gclk));
	jor g2175(.dina(n2437),.dinb(n2436),.dout(n2438),.clk(gclk));
	jand g2176(.dina(w_n2026_1[0]),.dinb(w_n265_44[0]),.dout(n2439),.clk(gclk));
	jor g2177(.dina(w_dff_B_H5CDb6oE6_0),.dinb(n2438),.dout(n2440),.clk(gclk));
	jor g2178(.dina(n2440),.dinb(w_dff_B_liuz3nrk5_1),.dout(n2441),.clk(gclk));
	jor g2179(.dina(w_n2441_0[1]),.dinb(w_n263_53[2]),.dout(n2442),.clk(gclk));
	jand g2180(.dina(w_n2062_1[0]),.dinb(w_n410_43[2]),.dout(n2443),.clk(gclk));
	jand g2181(.dina(w_n2053_1[0]),.dinb(w_n319_43[2]),.dout(n2444),.clk(gclk));
	jand g2182(.dina(w_n2045_1[0]),.dinb(w_n265_43[2]),.dout(n2445),.clk(gclk));
	jor g2183(.dina(n2445),.dinb(n2444),.dout(n2446),.clk(gclk));
	jand g2184(.dina(w_n2009_1[0]),.dinb(w_n364_43[2]),.dout(n2447),.clk(gclk));
	jor g2185(.dina(w_dff_B_SGLp9wMj4_0),.dinb(n2446),.dout(n2448),.clk(gclk));
	jor g2186(.dina(n2448),.dinb(w_dff_B_KAogdi844_1),.dout(n2449),.clk(gclk));
	jor g2187(.dina(w_n2449_0[1]),.dinb(w_shift6_53[2]),.dout(n2450),.clk(gclk));
	jand g2188(.dina(n2450),.dinb(n2442),.dout(result29),.clk(gclk));
	jand g2189(.dina(w_n2090_1[0]),.dinb(w_n319_43[1]),.dout(n2452),.clk(gclk));
	jand g2190(.dina(w_n2135_1[0]),.dinb(w_n364_43[1]),.dout(n2453),.clk(gclk));
	jand g2191(.dina(w_n2099_1[0]),.dinb(w_n410_43[1]),.dout(n2454),.clk(gclk));
	jor g2192(.dina(n2454),.dinb(n2453),.dout(n2455),.clk(gclk));
	jand g2193(.dina(w_n2074_1[0]),.dinb(w_n265_43[1]),.dout(n2456),.clk(gclk));
	jor g2194(.dina(w_dff_B_M6qUBrYh2_0),.dinb(n2455),.dout(n2457),.clk(gclk));
	jor g2195(.dina(n2457),.dinb(w_dff_B_DnS9XDKT8_1),.dout(n2458),.clk(gclk));
	jor g2196(.dina(w_n2458_0[1]),.dinb(w_n263_53[1]),.dout(n2459),.clk(gclk));
	jand g2197(.dina(w_n2082_1[0]),.dinb(w_n364_43[0]),.dout(n2460),.clk(gclk));
	jand g2198(.dina(w_n2126_1[0]),.dinb(w_n319_43[0]),.dout(n2461),.clk(gclk));
	jand g2199(.dina(w_n2118_1[0]),.dinb(w_n265_43[0]),.dout(n2462),.clk(gclk));
	jor g2200(.dina(n2462),.dinb(n2461),.dout(n2463),.clk(gclk));
	jand g2201(.dina(w_n2110_1[0]),.dinb(w_n410_43[0]),.dout(n2464),.clk(gclk));
	jor g2202(.dina(w_dff_B_RgGRMQHE6_0),.dinb(n2463),.dout(n2465),.clk(gclk));
	jor g2203(.dina(n2465),.dinb(w_dff_B_MG0suzb56_1),.dout(n2466),.clk(gclk));
	jor g2204(.dina(w_n2466_0[1]),.dinb(w_shift6_53[1]),.dout(n2467),.clk(gclk));
	jand g2205(.dina(n2467),.dinb(n2459),.dout(result30),.clk(gclk));
	jand g2206(.dina(w_n2147_1[0]),.dinb(w_n265_42[2]),.dout(n2469),.clk(gclk));
	jand g2207(.dina(w_n2208_1[0]),.dinb(w_n364_42[2]),.dout(n2470),.clk(gclk));
	jand g2208(.dina(w_n2163_1[0]),.dinb(w_n410_42[2]),.dout(n2471),.clk(gclk));
	jor g2209(.dina(n2471),.dinb(n2470),.dout(n2472),.clk(gclk));
	jand g2210(.dina(w_n2172_1[0]),.dinb(w_n319_42[2]),.dout(n2473),.clk(gclk));
	jor g2211(.dina(w_dff_B_lNX9XknG9_0),.dinb(n2472),.dout(n2474),.clk(gclk));
	jor g2212(.dina(n2474),.dinb(w_dff_B_9qAu6CEv6_1),.dout(n2475),.clk(gclk));
	jor g2213(.dina(w_n2475_0[1]),.dinb(w_n263_53[0]),.dout(n2476),.clk(gclk));
	jand g2214(.dina(w_n2191_1[0]),.dinb(w_n265_42[1]),.dout(n2477),.clk(gclk));
	jand g2215(.dina(w_n2183_1[0]),.dinb(w_n319_42[1]),.dout(n2478),.clk(gclk));
	jand g2216(.dina(w_n2155_1[0]),.dinb(w_n364_42[1]),.dout(n2479),.clk(gclk));
	jor g2217(.dina(n2479),.dinb(n2478),.dout(n2480),.clk(gclk));
	jand g2218(.dina(w_n2199_1[0]),.dinb(w_n410_42[1]),.dout(n2481),.clk(gclk));
	jor g2219(.dina(w_dff_B_q2S1c17p8_0),.dinb(n2480),.dout(n2482),.clk(gclk));
	jor g2220(.dina(n2482),.dinb(w_dff_B_D9FffPJm6_1),.dout(n2483),.clk(gclk));
	jor g2221(.dina(w_n2483_0[1]),.dinb(w_shift6_53[0]),.dout(n2484),.clk(gclk));
	jand g2222(.dina(n2484),.dinb(n2476),.dout(result31),.clk(gclk));
	jand g2223(.dina(w_n500_0[2]),.dinb(w_n319_42[0]),.dout(n2486),.clk(gclk));
	jand g2224(.dina(w_n410_42[0]),.dinb(w_n362_0[2]),.dout(n2487),.clk(gclk));
	jand g2225(.dina(w_n588_0[2]),.dinb(w_n364_42[0]),.dout(n2488),.clk(gclk));
	jor g2226(.dina(n2488),.dinb(n2487),.dout(n2489),.clk(gclk));
	jand g2227(.dina(w_n407_0[2]),.dinb(w_n265_42[0]),.dout(n2490),.clk(gclk));
	jor g2228(.dina(w_dff_B_9iVsnI3Y0_0),.dinb(n2489),.dout(n2491),.clk(gclk));
	jor g2229(.dina(n2491),.dinb(w_dff_B_yVPVbjPP6_1),.dout(n2492),.clk(gclk));
	jor g2230(.dina(w_n2492_0[1]),.dinb(w_n263_52[2]),.dout(n2493),.clk(gclk));
	jand g2231(.dina(w_n633_0[2]),.dinb(w_n265_41[2]),.dout(n2494),.clk(gclk));
	jand g2232(.dina(w_n453_0[2]),.dinb(w_n319_41[2]),.dout(n2495),.clk(gclk));
	jand g2233(.dina(w_n364_41[2]),.dinb(w_n316_0[2]),.dout(n2496),.clk(gclk));
	jor g2234(.dina(n2496),.dinb(n2495),.dout(n2497),.clk(gclk));
	jand g2235(.dina(w_n544_0[2]),.dinb(w_n410_41[2]),.dout(n2498),.clk(gclk));
	jor g2236(.dina(w_dff_B_bTy0068r1_0),.dinb(n2497),.dout(n2499),.clk(gclk));
	jor g2237(.dina(n2499),.dinb(w_dff_B_a3CGe7202_1),.dout(n2500),.clk(gclk));
	jor g2238(.dina(w_n2500_0[1]),.dinb(w_shift6_52[2]),.dout(n2501),.clk(gclk));
	jand g2239(.dina(n2501),.dinb(n2493),.dout(result32),.clk(gclk));
	jand g2240(.dina(w_n861_0[2]),.dinb(w_n319_41[1]),.dout(n2503),.clk(gclk));
	jand g2241(.dina(w_n949_0[2]),.dinb(w_n364_41[1]),.dout(n2504),.clk(gclk));
	jand g2242(.dina(w_n814_0[2]),.dinb(w_n410_41[1]),.dout(n2505),.clk(gclk));
	jor g2243(.dina(n2505),.dinb(n2504),.dout(n2506),.clk(gclk));
	jand g2244(.dina(w_n681_0[2]),.dinb(w_n265_41[1]),.dout(n2507),.clk(gclk));
	jor g2245(.dina(w_dff_B_7kVOx8kZ8_0),.dinb(n2506),.dout(n2508),.clk(gclk));
	jor g2246(.dina(n2508),.dinb(w_dff_B_19lEeWUB7_1),.dout(n2509),.clk(gclk));
	jor g2247(.dina(w_n2509_0[1]),.dinb(w_n263_52[1]),.dout(n2510),.clk(gclk));
	jand g2248(.dina(w_n994_0[2]),.dinb(w_n265_41[0]),.dout(n2511),.clk(gclk));
	jand g2249(.dina(w_n769_0[2]),.dinb(w_n319_41[0]),.dout(n2512),.clk(gclk));
	jand g2250(.dina(w_n725_0[2]),.dinb(w_n364_41[0]),.dout(n2513),.clk(gclk));
	jor g2251(.dina(n2513),.dinb(n2512),.dout(n2514),.clk(gclk));
	jand g2252(.dina(w_n905_0[2]),.dinb(w_n410_41[0]),.dout(n2515),.clk(gclk));
	jor g2253(.dina(w_dff_B_boPyw8vw4_0),.dinb(n2514),.dout(n2516),.clk(gclk));
	jor g2254(.dina(n2516),.dinb(w_dff_B_7HQfPZQp1_1),.dout(n2517),.clk(gclk));
	jor g2255(.dina(w_n2517_0[1]),.dinb(w_shift6_52[1]),.dout(n2518),.clk(gclk));
	jand g2256(.dina(n2518),.dinb(n2510),.dout(result33),.clk(gclk));
	jand g2257(.dina(w_n1079_0[2]),.dinb(w_n265_40[2]),.dout(n2520),.clk(gclk));
	jand g2258(.dina(w_n1163_0[2]),.dinb(w_n364_40[2]),.dout(n2521),.clk(gclk));
	jand g2259(.dina(w_n1102_0[2]),.dinb(w_n319_40[2]),.dout(n2522),.clk(gclk));
	jor g2260(.dina(n2522),.dinb(n2521),.dout(n2523),.clk(gclk));
	jand g2261(.dina(w_n1018_0[2]),.dinb(w_n410_40[2]),.dout(n2524),.clk(gclk));
	jor g2262(.dina(w_dff_B_YFkbXwkf8_0),.dinb(n2523),.dout(n2525),.clk(gclk));
	jor g2263(.dina(n2525),.dinb(w_dff_B_ky9JnIJa0_1),.dout(n2526),.clk(gclk));
	jor g2264(.dina(w_n2526_0[1]),.dinb(w_n263_52[0]),.dout(n2527),.clk(gclk));
	jand g2265(.dina(w_n1122_0[2]),.dinb(w_n410_40[1]),.dout(n2528),.clk(gclk));
	jand g2266(.dina(w_n1058_0[2]),.dinb(w_n319_40[1]),.dout(n2529),.clk(gclk));
	jand g2267(.dina(w_n1142_0[2]),.dinb(w_n265_40[1]),.dout(n2530),.clk(gclk));
	jor g2268(.dina(n2530),.dinb(n2529),.dout(n2531),.clk(gclk));
	jand g2269(.dina(w_n1038_0[2]),.dinb(w_n364_40[1]),.dout(n2532),.clk(gclk));
	jor g2270(.dina(w_dff_B_9obNFDpn5_0),.dinb(n2531),.dout(n2533),.clk(gclk));
	jor g2271(.dina(n2533),.dinb(w_dff_B_FwE6F5NN2_1),.dout(n2534),.clk(gclk));
	jor g2272(.dina(w_n2534_0[1]),.dinb(w_shift6_52[0]),.dout(n2535),.clk(gclk));
	jand g2273(.dina(n2535),.dinb(n2527),.dout(result34),.clk(gclk));
	jand g2274(.dina(w_n1187_0[2]),.dinb(w_n265_40[0]),.dout(n2537),.clk(gclk));
	jand g2275(.dina(w_n1291_0[2]),.dinb(w_n319_40[0]),.dout(n2538),.clk(gclk));
	jand g2276(.dina(w_n1332_0[2]),.dinb(w_n364_40[0]),.dout(n2539),.clk(gclk));
	jor g2277(.dina(n2539),.dinb(n2538),.dout(n2540),.clk(gclk));
	jand g2278(.dina(w_n1248_0[2]),.dinb(w_n410_40[0]),.dout(n2541),.clk(gclk));
	jor g2279(.dina(w_dff_B_YdezcyHU5_0),.dinb(n2540),.dout(n2542),.clk(gclk));
	jor g2280(.dina(n2542),.dinb(w_dff_B_4eITFKR93_1),.dout(n2543),.clk(gclk));
	jor g2281(.dina(w_n2543_0[1]),.dinb(w_n263_51[2]),.dout(n2544),.clk(gclk));
	jand g2282(.dina(w_n1271_0[2]),.dinb(w_n410_39[2]),.dout(n2545),.clk(gclk));
	jand g2283(.dina(w_n1227_0[2]),.dinb(w_n319_39[2]),.dout(n2546),.clk(gclk));
	jand g2284(.dina(w_n1311_0[2]),.dinb(w_n265_39[2]),.dout(n2547),.clk(gclk));
	jor g2285(.dina(n2547),.dinb(n2546),.dout(n2548),.clk(gclk));
	jand g2286(.dina(w_n1207_0[2]),.dinb(w_n364_39[2]),.dout(n2549),.clk(gclk));
	jor g2287(.dina(w_dff_B_0hEDWuI26_0),.dinb(n2548),.dout(n2550),.clk(gclk));
	jor g2288(.dina(n2550),.dinb(w_dff_B_f6wrL0AW5_1),.dout(n2551),.clk(gclk));
	jor g2289(.dina(w_n2551_0[1]),.dinb(w_shift6_51[2]),.dout(n2552),.clk(gclk));
	jand g2290(.dina(n2552),.dinb(n2544),.dout(result35),.clk(gclk));
	jand g2291(.dina(w_n1405_0[2]),.dinb(w_n319_39[1]),.dout(n2554),.clk(gclk));
	jand g2292(.dina(w_n1369_0[2]),.dinb(w_n410_39[1]),.dout(n2555),.clk(gclk));
	jand g2293(.dina(w_n1380_0[2]),.dinb(w_n364_39[1]),.dout(n2556),.clk(gclk));
	jor g2294(.dina(n2556),.dinb(n2555),.dout(n2557),.clk(gclk));
	jand g2295(.dina(w_n1344_0[2]),.dinb(w_n265_39[1]),.dout(n2558),.clk(gclk));
	jor g2296(.dina(w_dff_B_qB6dFw1e2_0),.dinb(n2557),.dout(n2559),.clk(gclk));
	jor g2297(.dina(n2559),.dinb(w_dff_B_0Z3CSdIH1_1),.dout(n2560),.clk(gclk));
	jor g2298(.dina(w_n2560_0[1]),.dinb(w_n263_51[1]),.dout(n2561),.clk(gclk));
	jand g2299(.dina(w_n1396_0[2]),.dinb(w_n265_39[0]),.dout(n2562),.clk(gclk));
	jand g2300(.dina(w_n1352_0[2]),.dinb(w_n319_39[0]),.dout(n2563),.clk(gclk));
	jand g2301(.dina(w_n1360_0[2]),.dinb(w_n364_39[0]),.dout(n2564),.clk(gclk));
	jor g2302(.dina(n2564),.dinb(n2563),.dout(n2565),.clk(gclk));
	jand g2303(.dina(w_n1388_0[2]),.dinb(w_n410_39[0]),.dout(n2566),.clk(gclk));
	jor g2304(.dina(w_dff_B_u3F8t7vU1_0),.dinb(n2565),.dout(n2567),.clk(gclk));
	jor g2305(.dina(n2567),.dinb(w_dff_B_f4xDkURy7_1),.dout(n2568),.clk(gclk));
	jor g2306(.dina(w_n2568_0[1]),.dinb(w_shift6_51[1]),.dout(n2569),.clk(gclk));
	jand g2307(.dina(n2569),.dinb(n2561),.dout(result36),.clk(gclk));
	jand g2308(.dina(w_n1453_0[2]),.dinb(w_n319_38[2]),.dout(n2571),.clk(gclk));
	jand g2309(.dina(w_n1417_0[2]),.dinb(w_n410_38[2]),.dout(n2572),.clk(gclk));
	jand g2310(.dina(w_n1469_0[2]),.dinb(w_n364_38[2]),.dout(n2573),.clk(gclk));
	jor g2311(.dina(n2573),.dinb(n2572),.dout(n2574),.clk(gclk));
	jand g2312(.dina(w_n1442_0[2]),.dinb(w_n265_38[2]),.dout(n2575),.clk(gclk));
	jor g2313(.dina(w_dff_B_huflLVnU8_0),.dinb(n2574),.dout(n2576),.clk(gclk));
	jor g2314(.dina(n2576),.dinb(w_dff_B_OQ4nf9FB4_1),.dout(n2577),.clk(gclk));
	jor g2315(.dina(w_n2577_0[1]),.dinb(w_n263_51[0]),.dout(n2578),.clk(gclk));
	jand g2316(.dina(w_n1461_0[2]),.dinb(w_n410_38[1]),.dout(n2579),.clk(gclk));
	jand g2317(.dina(w_n1425_0[2]),.dinb(w_n319_38[1]),.dout(n2580),.clk(gclk));
	jand g2318(.dina(w_n1433_0[2]),.dinb(w_n364_38[1]),.dout(n2581),.clk(gclk));
	jor g2319(.dina(n2581),.dinb(n2580),.dout(n2582),.clk(gclk));
	jand g2320(.dina(w_n1478_0[2]),.dinb(w_n265_38[1]),.dout(n2583),.clk(gclk));
	jor g2321(.dina(w_dff_B_X8hTW4sa2_0),.dinb(n2582),.dout(n2584),.clk(gclk));
	jor g2322(.dina(n2584),.dinb(w_dff_B_N2r3icPs2_1),.dout(n2585),.clk(gclk));
	jor g2323(.dina(w_n2585_0[1]),.dinb(w_shift6_51[0]),.dout(n2586),.clk(gclk));
	jand g2324(.dina(n2586),.dinb(n2578),.dout(result37),.clk(gclk));
	jand g2325(.dina(w_n1506_0[2]),.dinb(w_n265_38[0]),.dout(n2588),.clk(gclk));
	jand g2326(.dina(w_n1515_0[2]),.dinb(w_n410_38[0]),.dout(n2589),.clk(gclk));
	jand g2327(.dina(w_n1551_0[2]),.dinb(w_n364_38[0]),.dout(n2590),.clk(gclk));
	jor g2328(.dina(n2590),.dinb(n2589),.dout(n2591),.clk(gclk));
	jand g2329(.dina(w_n1526_0[2]),.dinb(w_n319_38[0]),.dout(n2592),.clk(gclk));
	jor g2330(.dina(w_dff_B_aEdf5wZc7_0),.dinb(n2591),.dout(n2593),.clk(gclk));
	jor g2331(.dina(n2593),.dinb(w_dff_B_nr95JRAm8_1),.dout(n2594),.clk(gclk));
	jor g2332(.dina(w_n2594_0[1]),.dinb(w_n263_50[2]),.dout(n2595),.clk(gclk));
	jand g2333(.dina(w_n1534_0[2]),.dinb(w_n410_37[2]),.dout(n2596),.clk(gclk));
	jand g2334(.dina(w_n1498_0[2]),.dinb(w_n319_37[2]),.dout(n2597),.clk(gclk));
	jand g2335(.dina(w_n1542_0[2]),.dinb(w_n265_37[2]),.dout(n2598),.clk(gclk));
	jor g2336(.dina(n2598),.dinb(n2597),.dout(n2599),.clk(gclk));
	jand g2337(.dina(w_n1490_0[2]),.dinb(w_n364_37[2]),.dout(n2600),.clk(gclk));
	jor g2338(.dina(w_dff_B_C34EYOny8_0),.dinb(n2599),.dout(n2601),.clk(gclk));
	jor g2339(.dina(n2601),.dinb(w_dff_B_nkiDrsDo7_1),.dout(n2602),.clk(gclk));
	jor g2340(.dina(w_n2602_0[1]),.dinb(w_shift6_50[2]),.dout(n2603),.clk(gclk));
	jand g2341(.dina(n2603),.dinb(n2595),.dout(result38),.clk(gclk));
	jand g2342(.dina(w_n1588_0[2]),.dinb(w_n410_37[1]),.dout(n2605),.clk(gclk));
	jand g2343(.dina(w_n1599_0[2]),.dinb(w_n319_37[1]),.dout(n2606),.clk(gclk));
	jand g2344(.dina(w_n1579_0[2]),.dinb(w_n265_37[1]),.dout(n2607),.clk(gclk));
	jor g2345(.dina(n2607),.dinb(n2606),.dout(n2608),.clk(gclk));
	jand g2346(.dina(w_n1615_0[2]),.dinb(w_n364_37[1]),.dout(n2609),.clk(gclk));
	jor g2347(.dina(w_dff_B_YWRYZVvo7_0),.dinb(n2608),.dout(n2610),.clk(gclk));
	jor g2348(.dina(n2610),.dinb(w_dff_B_b7uSIuaZ4_1),.dout(n2611),.clk(gclk));
	jor g2349(.dina(w_n2611_0[1]),.dinb(w_n263_50[1]),.dout(n2612),.clk(gclk));
	jand g2350(.dina(w_n1571_0[2]),.dinb(w_n319_37[0]),.dout(n2613),.clk(gclk));
	jand g2351(.dina(w_n1607_0[2]),.dinb(w_n410_37[0]),.dout(n2614),.clk(gclk));
	jand g2352(.dina(w_n1563_0[2]),.dinb(w_n364_37[0]),.dout(n2615),.clk(gclk));
	jor g2353(.dina(n2615),.dinb(n2614),.dout(n2616),.clk(gclk));
	jand g2354(.dina(w_n1624_0[2]),.dinb(w_n265_37[0]),.dout(n2617),.clk(gclk));
	jor g2355(.dina(w_dff_B_496Qayul4_0),.dinb(n2616),.dout(n2618),.clk(gclk));
	jor g2356(.dina(n2618),.dinb(w_dff_B_CrXB06rb5_1),.dout(n2619),.clk(gclk));
	jor g2357(.dina(w_n2619_0[1]),.dinb(w_shift6_50[1]),.dout(n2620),.clk(gclk));
	jand g2358(.dina(n2620),.dinb(n2612),.dout(result39),.clk(gclk));
	jand g2359(.dina(w_n1661_0[2]),.dinb(w_n410_36[2]),.dout(n2622),.clk(gclk));
	jand g2360(.dina(w_n1672_0[2]),.dinb(w_n319_36[2]),.dout(n2623),.clk(gclk));
	jand g2361(.dina(w_n1697_0[2]),.dinb(w_n364_36[2]),.dout(n2624),.clk(gclk));
	jor g2362(.dina(n2624),.dinb(n2623),.dout(n2625),.clk(gclk));
	jand g2363(.dina(w_n1652_0[2]),.dinb(w_n265_36[2]),.dout(n2626),.clk(gclk));
	jor g2364(.dina(w_dff_B_gh9Bjk4K5_0),.dinb(n2625),.dout(n2627),.clk(gclk));
	jor g2365(.dina(n2627),.dinb(w_dff_B_V9UeSrPZ8_1),.dout(n2628),.clk(gclk));
	jor g2366(.dina(w_n2628_0[1]),.dinb(w_n263_50[0]),.dout(n2629),.clk(gclk));
	jand g2367(.dina(w_n1688_0[2]),.dinb(w_n265_36[1]),.dout(n2630),.clk(gclk));
	jand g2368(.dina(w_n1680_0[2]),.dinb(w_n410_36[1]),.dout(n2631),.clk(gclk));
	jand g2369(.dina(w_n1636_0[2]),.dinb(w_n364_36[1]),.dout(n2632),.clk(gclk));
	jor g2370(.dina(n2632),.dinb(n2631),.dout(n2633),.clk(gclk));
	jand g2371(.dina(w_n1644_0[2]),.dinb(w_n319_36[1]),.dout(n2634),.clk(gclk));
	jor g2372(.dina(w_dff_B_Onbv6u1X0_0),.dinb(n2633),.dout(n2635),.clk(gclk));
	jor g2373(.dina(n2635),.dinb(w_dff_B_uj3d5Aa12_1),.dout(n2636),.clk(gclk));
	jor g2374(.dina(w_n2636_0[1]),.dinb(w_shift6_50[0]),.dout(n2637),.clk(gclk));
	jand g2375(.dina(n2637),.dinb(n2629),.dout(result40),.clk(gclk));
	jand g2376(.dina(w_n1709_0[2]),.dinb(w_n265_36[0]),.dout(n2639),.clk(gclk));
	jand g2377(.dina(w_n1770_0[2]),.dinb(w_n319_36[0]),.dout(n2640),.clk(gclk));
	jand g2378(.dina(w_n1745_0[2]),.dinb(w_n364_36[0]),.dout(n2641),.clk(gclk));
	jor g2379(.dina(n2641),.dinb(n2640),.dout(n2642),.clk(gclk));
	jand g2380(.dina(w_n1734_0[2]),.dinb(w_n410_36[0]),.dout(n2643),.clk(gclk));
	jor g2381(.dina(w_dff_B_ocQxDi7i4_0),.dinb(n2642),.dout(n2644),.clk(gclk));
	jor g2382(.dina(n2644),.dinb(w_dff_B_edIm3HEo0_1),.dout(n2645),.clk(gclk));
	jor g2383(.dina(w_n2645_0[1]),.dinb(w_n263_49[2]),.dout(n2646),.clk(gclk));
	jand g2384(.dina(w_n1717_0[2]),.dinb(w_n319_35[2]),.dout(n2647),.clk(gclk));
	jand g2385(.dina(w_n1753_0[2]),.dinb(w_n410_35[2]),.dout(n2648),.clk(gclk));
	jand g2386(.dina(w_n1725_0[2]),.dinb(w_n364_35[2]),.dout(n2649),.clk(gclk));
	jor g2387(.dina(n2649),.dinb(n2648),.dout(n2650),.clk(gclk));
	jand g2388(.dina(w_n1761_0[2]),.dinb(w_n265_35[2]),.dout(n2651),.clk(gclk));
	jor g2389(.dina(w_dff_B_ZqWDHNKl8_0),.dinb(n2650),.dout(n2652),.clk(gclk));
	jor g2390(.dina(n2652),.dinb(w_dff_B_Sy8fXmtO9_1),.dout(n2653),.clk(gclk));
	jor g2391(.dina(w_n2653_0[1]),.dinb(w_shift6_49[2]),.dout(n2654),.clk(gclk));
	jand g2392(.dina(n2654),.dinb(n2646),.dout(result41),.clk(gclk));
	jand g2393(.dina(w_n1782_0[2]),.dinb(w_n410_35[1]),.dout(n2656),.clk(gclk));
	jand g2394(.dina(w_n1843_0[2]),.dinb(w_n319_35[1]),.dout(n2657),.clk(gclk));
	jand g2395(.dina(w_n1834_0[2]),.dinb(w_n364_35[1]),.dout(n2658),.clk(gclk));
	jor g2396(.dina(n2658),.dinb(n2657),.dout(n2659),.clk(gclk));
	jand g2397(.dina(w_n1807_0[2]),.dinb(w_n265_35[1]),.dout(n2660),.clk(gclk));
	jor g2398(.dina(w_dff_B_rW47TtDh5_0),.dinb(n2659),.dout(n2661),.clk(gclk));
	jor g2399(.dina(n2661),.dinb(w_dff_B_SBRBhiff0_1),.dout(n2662),.clk(gclk));
	jor g2400(.dina(w_n2662_0[1]),.dinb(w_n263_49[1]),.dout(n2663),.clk(gclk));
	jand g2401(.dina(w_n1818_0[2]),.dinb(w_n265_35[0]),.dout(n2664),.clk(gclk));
	jand g2402(.dina(w_n1790_0[2]),.dinb(w_n319_35[0]),.dout(n2665),.clk(gclk));
	jand g2403(.dina(w_n1798_0[2]),.dinb(w_n364_35[0]),.dout(n2666),.clk(gclk));
	jor g2404(.dina(n2666),.dinb(n2665),.dout(n2667),.clk(gclk));
	jand g2405(.dina(w_n1826_0[2]),.dinb(w_n410_35[0]),.dout(n2668),.clk(gclk));
	jor g2406(.dina(w_dff_B_ujybVo5m3_0),.dinb(n2667),.dout(n2669),.clk(gclk));
	jor g2407(.dina(n2669),.dinb(w_dff_B_4prvR3SB9_1),.dout(n2670),.clk(gclk));
	jor g2408(.dina(w_n2670_0[1]),.dinb(w_shift6_49[1]),.dout(n2671),.clk(gclk));
	jand g2409(.dina(n2671),.dinb(n2663),.dout(result42),.clk(gclk));
	jand g2410(.dina(w_n1907_0[2]),.dinb(w_n364_34[2]),.dout(n2673),.clk(gclk));
	jand g2411(.dina(w_n1891_0[2]),.dinb(w_n319_34[2]),.dout(n2674),.clk(gclk));
	jand g2412(.dina(w_n1880_0[2]),.dinb(w_n265_34[2]),.dout(n2675),.clk(gclk));
	jor g2413(.dina(n2675),.dinb(n2674),.dout(n2676),.clk(gclk));
	jand g2414(.dina(w_n1855_0[2]),.dinb(w_n410_34[2]),.dout(n2677),.clk(gclk));
	jor g2415(.dina(w_dff_B_AJta4V6q0_0),.dinb(n2676),.dout(n2678),.clk(gclk));
	jor g2416(.dina(n2678),.dinb(w_dff_B_nh3K4oM22_1),.dout(n2679),.clk(gclk));
	jor g2417(.dina(w_n2679_0[1]),.dinb(w_n263_49[0]),.dout(n2680),.clk(gclk));
	jand g2418(.dina(w_n1871_0[2]),.dinb(w_n364_34[1]),.dout(n2681),.clk(gclk));
	jand g2419(.dina(w_n1863_0[2]),.dinb(w_n319_34[1]),.dout(n2682),.clk(gclk));
	jand g2420(.dina(w_n1916_0[2]),.dinb(w_n265_34[1]),.dout(n2683),.clk(gclk));
	jor g2421(.dina(n2683),.dinb(n2682),.dout(n2684),.clk(gclk));
	jand g2422(.dina(w_n1899_0[2]),.dinb(w_n410_34[1]),.dout(n2685),.clk(gclk));
	jor g2423(.dina(w_dff_B_x80yLBcc3_0),.dinb(n2684),.dout(n2686),.clk(gclk));
	jor g2424(.dina(n2686),.dinb(w_dff_B_43izO5SG7_1),.dout(n2687),.clk(gclk));
	jor g2425(.dina(w_n2687_0[1]),.dinb(w_shift6_49[0]),.dout(n2688),.clk(gclk));
	jand g2426(.dina(n2688),.dinb(n2680),.dout(result43),.clk(gclk));
	jand g2427(.dina(w_n1953_0[2]),.dinb(w_n410_34[0]),.dout(n2690),.clk(gclk));
	jand g2428(.dina(w_n1989_0[2]),.dinb(w_n319_34[0]),.dout(n2691),.clk(gclk));
	jand g2429(.dina(w_n1980_0[2]),.dinb(w_n364_34[0]),.dout(n2692),.clk(gclk));
	jor g2430(.dina(n2692),.dinb(n2691),.dout(n2693),.clk(gclk));
	jand g2431(.dina(w_n1944_0[2]),.dinb(w_n265_34[0]),.dout(n2694),.clk(gclk));
	jor g2432(.dina(w_dff_B_4o1boigc1_0),.dinb(n2693),.dout(n2695),.clk(gclk));
	jor g2433(.dina(n2695),.dinb(w_dff_B_UO0r7WtK8_1),.dout(n2696),.clk(gclk));
	jor g2434(.dina(w_n2696_0[1]),.dinb(w_n263_48[2]),.dout(n2697),.clk(gclk));
	jand g2435(.dina(w_n1964_0[2]),.dinb(w_n265_33[2]),.dout(n2698),.clk(gclk));
	jand g2436(.dina(w_n1936_0[2]),.dinb(w_n319_33[2]),.dout(n2699),.clk(gclk));
	jand g2437(.dina(w_n1928_0[2]),.dinb(w_n364_33[2]),.dout(n2700),.clk(gclk));
	jor g2438(.dina(n2700),.dinb(n2699),.dout(n2701),.clk(gclk));
	jand g2439(.dina(w_n1972_0[2]),.dinb(w_n410_33[2]),.dout(n2702),.clk(gclk));
	jor g2440(.dina(w_dff_B_A0PnvmfU3_0),.dinb(n2701),.dout(n2703),.clk(gclk));
	jor g2441(.dina(n2703),.dinb(w_dff_B_tFBmKSHU9_1),.dout(n2704),.clk(gclk));
	jor g2442(.dina(w_n2704_0[1]),.dinb(w_shift6_48[2]),.dout(n2705),.clk(gclk));
	jand g2443(.dina(n2705),.dinb(n2697),.dout(result44),.clk(gclk));
	jand g2444(.dina(w_n2017_0[2]),.dinb(w_n265_33[1]),.dout(n2707),.clk(gclk));
	jand g2445(.dina(w_n2037_0[2]),.dinb(w_n319_33[1]),.dout(n2708),.clk(gclk));
	jand g2446(.dina(w_n2062_0[2]),.dinb(w_n364_33[1]),.dout(n2709),.clk(gclk));
	jor g2447(.dina(n2709),.dinb(n2708),.dout(n2710),.clk(gclk));
	jand g2448(.dina(w_n2026_0[2]),.dinb(w_n410_33[1]),.dout(n2711),.clk(gclk));
	jor g2449(.dina(w_dff_B_YxqWpnGO2_0),.dinb(n2710),.dout(n2712),.clk(gclk));
	jor g2450(.dina(n2712),.dinb(w_dff_B_8tVKfkLJ8_1),.dout(n2713),.clk(gclk));
	jor g2451(.dina(w_n2713_0[1]),.dinb(w_n263_48[1]),.dout(n2714),.clk(gclk));
	jand g2452(.dina(w_n2045_0[2]),.dinb(w_n410_33[0]),.dout(n2715),.clk(gclk));
	jand g2453(.dina(w_n2009_0[2]),.dinb(w_n319_33[0]),.dout(n2716),.clk(gclk));
	jand g2454(.dina(w_n2053_0[2]),.dinb(w_n265_33[0]),.dout(n2717),.clk(gclk));
	jor g2455(.dina(n2717),.dinb(n2716),.dout(n2718),.clk(gclk));
	jand g2456(.dina(w_n2001_0[2]),.dinb(w_n364_33[0]),.dout(n2719),.clk(gclk));
	jor g2457(.dina(w_dff_B_0BpUHJ8f5_0),.dinb(n2718),.dout(n2720),.clk(gclk));
	jor g2458(.dina(n2720),.dinb(w_dff_B_DbMsD6I55_1),.dout(n2721),.clk(gclk));
	jor g2459(.dina(w_n2721_0[1]),.dinb(w_shift6_48[1]),.dout(n2722),.clk(gclk));
	jand g2460(.dina(n2722),.dinb(n2714),.dout(result45),.clk(gclk));
	jand g2461(.dina(w_n2110_0[2]),.dinb(w_n364_32[2]),.dout(n2724),.clk(gclk));
	jand g2462(.dina(w_n2135_0[2]),.dinb(w_n319_32[2]),.dout(n2725),.clk(gclk));
	jand g2463(.dina(w_n2090_0[2]),.dinb(w_n265_32[2]),.dout(n2726),.clk(gclk));
	jor g2464(.dina(n2726),.dinb(n2725),.dout(n2727),.clk(gclk));
	jand g2465(.dina(w_n2074_0[2]),.dinb(w_n410_32[2]),.dout(n2728),.clk(gclk));
	jor g2466(.dina(w_dff_B_jFPT1jCW9_0),.dinb(n2727),.dout(n2729),.clk(gclk));
	jor g2467(.dina(n2729),.dinb(w_dff_B_wOKdUDwI7_1),.dout(n2730),.clk(gclk));
	jor g2468(.dina(w_n2730_0[1]),.dinb(w_n263_48[0]),.dout(n2731),.clk(gclk));
	jand g2469(.dina(w_n2118_0[2]),.dinb(w_n410_32[1]),.dout(n2732),.clk(gclk));
	jand g2470(.dina(w_n2082_0[2]),.dinb(w_n319_32[1]),.dout(n2733),.clk(gclk));
	jand g2471(.dina(w_n2099_0[2]),.dinb(w_n364_32[1]),.dout(n2734),.clk(gclk));
	jor g2472(.dina(n2734),.dinb(n2733),.dout(n2735),.clk(gclk));
	jand g2473(.dina(w_n2126_0[2]),.dinb(w_n265_32[1]),.dout(n2736),.clk(gclk));
	jor g2474(.dina(w_dff_B_3WWymGYL5_0),.dinb(n2735),.dout(n2737),.clk(gclk));
	jor g2475(.dina(n2737),.dinb(w_dff_B_TEUMczxJ9_1),.dout(n2738),.clk(gclk));
	jor g2476(.dina(w_n2738_0[1]),.dinb(w_shift6_48[0]),.dout(n2739),.clk(gclk));
	jand g2477(.dina(n2739),.dinb(n2731),.dout(result46),.clk(gclk));
	jand g2478(.dina(w_n2172_0[2]),.dinb(w_n265_32[0]),.dout(n2741),.clk(gclk));
	jand g2479(.dina(w_n2208_0[2]),.dinb(w_n319_32[0]),.dout(n2742),.clk(gclk));
	jand g2480(.dina(w_n2199_0[2]),.dinb(w_n364_32[0]),.dout(n2743),.clk(gclk));
	jor g2481(.dina(n2743),.dinb(n2742),.dout(n2744),.clk(gclk));
	jand g2482(.dina(w_n2147_0[2]),.dinb(w_n410_32[0]),.dout(n2745),.clk(gclk));
	jor g2483(.dina(w_dff_B_iXl7YkEZ9_0),.dinb(n2744),.dout(n2746),.clk(gclk));
	jor g2484(.dina(n2746),.dinb(w_dff_B_kLVUkxdA1_1),.dout(n2747),.clk(gclk));
	jor g2485(.dina(w_n2747_0[1]),.dinb(w_n263_47[2]),.dout(n2748),.clk(gclk));
	jand g2486(.dina(w_n2191_0[2]),.dinb(w_n410_31[2]),.dout(n2749),.clk(gclk));
	jand g2487(.dina(w_n2155_0[2]),.dinb(w_n319_31[2]),.dout(n2750),.clk(gclk));
	jand g2488(.dina(w_n2163_0[2]),.dinb(w_n364_31[2]),.dout(n2751),.clk(gclk));
	jor g2489(.dina(n2751),.dinb(n2750),.dout(n2752),.clk(gclk));
	jand g2490(.dina(w_n2183_0[2]),.dinb(w_n265_31[2]),.dout(n2753),.clk(gclk));
	jor g2491(.dina(w_dff_B_JOnwcef08_0),.dinb(n2752),.dout(n2754),.clk(gclk));
	jor g2492(.dina(n2754),.dinb(w_dff_B_4gZnAB7L0_1),.dout(n2755),.clk(gclk));
	jor g2493(.dina(w_n2755_0[1]),.dinb(w_shift6_47[2]),.dout(n2756),.clk(gclk));
	jand g2494(.dina(n2756),.dinb(n2748),.dout(result47),.clk(gclk));
	jand g2495(.dina(w_n410_31[1]),.dinb(w_n407_0[1]),.dout(n2758),.clk(gclk));
	jand g2496(.dina(w_n544_0[1]),.dinb(w_n364_31[1]),.dout(n2759),.clk(gclk));
	jand g2497(.dina(w_n588_0[1]),.dinb(w_n319_31[1]),.dout(n2760),.clk(gclk));
	jor g2498(.dina(n2760),.dinb(n2759),.dout(n2761),.clk(gclk));
	jand g2499(.dina(w_n500_0[1]),.dinb(w_n265_31[1]),.dout(n2762),.clk(gclk));
	jor g2500(.dina(w_dff_B_cjjRtxAq5_0),.dinb(n2761),.dout(n2763),.clk(gclk));
	jor g2501(.dina(n2763),.dinb(w_dff_B_feWNsbf75_1),.dout(n2764),.clk(gclk));
	jor g2502(.dina(w_n2764_0[1]),.dinb(w_n263_47[1]),.dout(n2765),.clk(gclk));
	jand g2503(.dina(w_n453_0[1]),.dinb(w_n265_31[0]),.dout(n2766),.clk(gclk));
	jand g2504(.dina(w_n319_31[0]),.dinb(w_n316_0[1]),.dout(n2767),.clk(gclk));
	jand g2505(.dina(w_n364_31[0]),.dinb(w_n362_0[1]),.dout(n2768),.clk(gclk));
	jor g2506(.dina(n2768),.dinb(n2767),.dout(n2769),.clk(gclk));
	jand g2507(.dina(w_n633_0[1]),.dinb(w_n410_31[0]),.dout(n2770),.clk(gclk));
	jor g2508(.dina(w_dff_B_9CCHJG3I8_0),.dinb(n2769),.dout(n2771),.clk(gclk));
	jor g2509(.dina(n2771),.dinb(w_dff_B_cZrHVwDG1_1),.dout(n2772),.clk(gclk));
	jor g2510(.dina(w_n2772_0[1]),.dinb(w_shift6_47[1]),.dout(n2773),.clk(gclk));
	jand g2511(.dina(n2773),.dinb(n2765),.dout(result48),.clk(gclk));
	jand g2512(.dina(w_n861_0[1]),.dinb(w_n265_30[2]),.dout(n2775),.clk(gclk));
	jand g2513(.dina(w_n949_0[1]),.dinb(w_n319_30[2]),.dout(n2776),.clk(gclk));
	jand g2514(.dina(w_n905_0[1]),.dinb(w_n364_30[2]),.dout(n2777),.clk(gclk));
	jor g2515(.dina(n2777),.dinb(n2776),.dout(n2778),.clk(gclk));
	jand g2516(.dina(w_n681_0[1]),.dinb(w_n410_30[2]),.dout(n2779),.clk(gclk));
	jor g2517(.dina(w_dff_B_jeXu3sy45_0),.dinb(n2778),.dout(n2780),.clk(gclk));
	jor g2518(.dina(n2780),.dinb(w_dff_B_T0GGtFnc1_1),.dout(n2781),.clk(gclk));
	jor g2519(.dina(w_n2781_0[1]),.dinb(w_n263_47[0]),.dout(n2782),.clk(gclk));
	jand g2520(.dina(w_n994_0[1]),.dinb(w_n410_30[1]),.dout(n2783),.clk(gclk));
	jand g2521(.dina(w_n725_0[1]),.dinb(w_n319_30[1]),.dout(n2784),.clk(gclk));
	jand g2522(.dina(w_n769_0[1]),.dinb(w_n265_30[1]),.dout(n2785),.clk(gclk));
	jor g2523(.dina(n2785),.dinb(n2784),.dout(n2786),.clk(gclk));
	jand g2524(.dina(w_n814_0[1]),.dinb(w_n364_30[1]),.dout(n2787),.clk(gclk));
	jor g2525(.dina(w_dff_B_MoX53rZY3_0),.dinb(n2786),.dout(n2788),.clk(gclk));
	jor g2526(.dina(n2788),.dinb(w_dff_B_pWTH2BSY6_1),.dout(n2789),.clk(gclk));
	jor g2527(.dina(w_n2789_0[1]),.dinb(w_shift6_47[0]),.dout(n2790),.clk(gclk));
	jand g2528(.dina(n2790),.dinb(n2782),.dout(result49),.clk(gclk));
	jand g2529(.dina(w_n1079_0[1]),.dinb(w_n410_30[0]),.dout(n2792),.clk(gclk));
	jand g2530(.dina(w_n1163_0[1]),.dinb(w_n319_30[0]),.dout(n2793),.clk(gclk));
	jand g2531(.dina(w_n1102_0[1]),.dinb(w_n265_30[0]),.dout(n2794),.clk(gclk));
	jor g2532(.dina(n2794),.dinb(n2793),.dout(n2795),.clk(gclk));
	jand g2533(.dina(w_n1122_0[1]),.dinb(w_n364_30[0]),.dout(n2796),.clk(gclk));
	jor g2534(.dina(w_dff_B_YOJR5kVR6_0),.dinb(n2795),.dout(n2797),.clk(gclk));
	jor g2535(.dina(n2797),.dinb(w_dff_B_h6gd19k23_1),.dout(n2798),.clk(gclk));
	jor g2536(.dina(w_n2798_0[1]),.dinb(w_n263_46[2]),.dout(n2799),.clk(gclk));
	jand g2537(.dina(w_n1018_0[1]),.dinb(w_n364_29[2]),.dout(n2800),.clk(gclk));
	jand g2538(.dina(w_n1038_0[1]),.dinb(w_n319_29[2]),.dout(n2801),.clk(gclk));
	jand g2539(.dina(w_n1058_0[1]),.dinb(w_n265_29[2]),.dout(n2802),.clk(gclk));
	jor g2540(.dina(n2802),.dinb(n2801),.dout(n2803),.clk(gclk));
	jand g2541(.dina(w_n1142_0[1]),.dinb(w_n410_29[2]),.dout(n2804),.clk(gclk));
	jor g2542(.dina(w_dff_B_qG7CcZVr6_0),.dinb(n2803),.dout(n2805),.clk(gclk));
	jor g2543(.dina(n2805),.dinb(w_dff_B_n9pUpmqm8_1),.dout(n2806),.clk(gclk));
	jor g2544(.dina(w_n2806_0[1]),.dinb(w_shift6_46[2]),.dout(n2807),.clk(gclk));
	jand g2545(.dina(n2807),.dinb(n2799),.dout(result50),.clk(gclk));
	jand g2546(.dina(w_n1187_0[1]),.dinb(w_n410_29[1]),.dout(n2809),.clk(gclk));
	jand g2547(.dina(w_n1332_0[1]),.dinb(w_n319_29[1]),.dout(n2810),.clk(gclk));
	jand g2548(.dina(w_n1291_0[1]),.dinb(w_n265_29[1]),.dout(n2811),.clk(gclk));
	jor g2549(.dina(n2811),.dinb(n2810),.dout(n2812),.clk(gclk));
	jand g2550(.dina(w_n1271_0[1]),.dinb(w_n364_29[1]),.dout(n2813),.clk(gclk));
	jor g2551(.dina(w_dff_B_B3HjuQuU9_0),.dinb(n2812),.dout(n2814),.clk(gclk));
	jor g2552(.dina(n2814),.dinb(w_dff_B_XrRsKiC06_1),.dout(n2815),.clk(gclk));
	jor g2553(.dina(w_n2815_0[1]),.dinb(w_n263_46[1]),.dout(n2816),.clk(gclk));
	jand g2554(.dina(w_n1248_0[1]),.dinb(w_n364_29[0]),.dout(n2817),.clk(gclk));
	jand g2555(.dina(w_n1227_0[1]),.dinb(w_n265_29[0]),.dout(n2818),.clk(gclk));
	jand g2556(.dina(w_n1207_0[1]),.dinb(w_n319_29[0]),.dout(n2819),.clk(gclk));
	jor g2557(.dina(n2819),.dinb(n2818),.dout(n2820),.clk(gclk));
	jand g2558(.dina(w_n1311_0[1]),.dinb(w_n410_29[0]),.dout(n2821),.clk(gclk));
	jor g2559(.dina(w_dff_B_SOdTOQwU7_0),.dinb(n2820),.dout(n2822),.clk(gclk));
	jor g2560(.dina(n2822),.dinb(w_dff_B_VMQQNRP08_1),.dout(n2823),.clk(gclk));
	jor g2561(.dina(w_n2823_0[1]),.dinb(w_shift6_46[1]),.dout(n2824),.clk(gclk));
	jand g2562(.dina(n2824),.dinb(n2816),.dout(result51),.clk(gclk));
	jand g2563(.dina(w_n1380_0[1]),.dinb(w_n319_28[2]),.dout(n2826),.clk(gclk));
	jand g2564(.dina(w_n1344_0[1]),.dinb(w_n410_28[2]),.dout(n2827),.clk(gclk));
	jand g2565(.dina(w_n1388_0[1]),.dinb(w_n364_28[2]),.dout(n2828),.clk(gclk));
	jor g2566(.dina(n2828),.dinb(n2827),.dout(n2829),.clk(gclk));
	jand g2567(.dina(w_n1405_0[1]),.dinb(w_n265_28[2]),.dout(n2830),.clk(gclk));
	jor g2568(.dina(w_dff_B_7IMUWZDl2_0),.dinb(n2829),.dout(n2831),.clk(gclk));
	jor g2569(.dina(n2831),.dinb(w_dff_B_GEI0pHLe2_1),.dout(n2832),.clk(gclk));
	jor g2570(.dina(w_n2832_0[1]),.dinb(w_n263_46[0]),.dout(n2833),.clk(gclk));
	jand g2571(.dina(w_n1360_0[1]),.dinb(w_n319_28[1]),.dout(n2834),.clk(gclk));
	jand g2572(.dina(w_n1352_0[1]),.dinb(w_n265_28[1]),.dout(n2835),.clk(gclk));
	jand g2573(.dina(w_n1396_0[1]),.dinb(w_n410_28[1]),.dout(n2836),.clk(gclk));
	jor g2574(.dina(n2836),.dinb(n2835),.dout(n2837),.clk(gclk));
	jand g2575(.dina(w_n1369_0[1]),.dinb(w_n364_28[1]),.dout(n2838),.clk(gclk));
	jor g2576(.dina(w_dff_B_IHsLOWpC2_0),.dinb(n2837),.dout(n2839),.clk(gclk));
	jor g2577(.dina(n2839),.dinb(w_dff_B_IEnkpo8q6_1),.dout(n2840),.clk(gclk));
	jor g2578(.dina(w_n2840_0[1]),.dinb(w_shift6_46[0]),.dout(n2841),.clk(gclk));
	jand g2579(.dina(n2841),.dinb(n2833),.dout(result52),.clk(gclk));
	jand g2580(.dina(w_n1453_0[1]),.dinb(w_n265_28[0]),.dout(n2843),.clk(gclk));
	jand g2581(.dina(w_n1442_0[1]),.dinb(w_n410_28[0]),.dout(n2844),.clk(gclk));
	jand g2582(.dina(w_n1469_0[1]),.dinb(w_n319_28[0]),.dout(n2845),.clk(gclk));
	jor g2583(.dina(n2845),.dinb(n2844),.dout(n2846),.clk(gclk));
	jand g2584(.dina(w_n1461_0[1]),.dinb(w_n364_28[0]),.dout(n2847),.clk(gclk));
	jor g2585(.dina(w_dff_B_mfvk1noa9_0),.dinb(n2846),.dout(n2848),.clk(gclk));
	jor g2586(.dina(n2848),.dinb(w_dff_B_3wuBCOe82_1),.dout(n2849),.clk(gclk));
	jor g2587(.dina(w_n2849_0[1]),.dinb(w_n263_45[2]),.dout(n2850),.clk(gclk));
	jand g2588(.dina(w_n1417_0[1]),.dinb(w_n364_27[2]),.dout(n2851),.clk(gclk));
	jand g2589(.dina(w_n1425_0[1]),.dinb(w_n265_27[2]),.dout(n2852),.clk(gclk));
	jand g2590(.dina(w_n1433_0[1]),.dinb(w_n319_27[2]),.dout(n2853),.clk(gclk));
	jor g2591(.dina(n2853),.dinb(n2852),.dout(n2854),.clk(gclk));
	jand g2592(.dina(w_n1478_0[1]),.dinb(w_n410_27[2]),.dout(n2855),.clk(gclk));
	jor g2593(.dina(w_dff_B_7Xuq5K5W5_0),.dinb(n2854),.dout(n2856),.clk(gclk));
	jor g2594(.dina(n2856),.dinb(w_dff_B_FRrwnx3T2_1),.dout(n2857),.clk(gclk));
	jor g2595(.dina(w_n2857_0[1]),.dinb(w_shift6_45[2]),.dout(n2858),.clk(gclk));
	jand g2596(.dina(n2858),.dinb(n2850),.dout(result53),.clk(gclk));
	jand g2597(.dina(w_n1534_0[1]),.dinb(w_n364_27[1]),.dout(n2860),.clk(gclk));
	jand g2598(.dina(w_n1506_0[1]),.dinb(w_n410_27[1]),.dout(n2861),.clk(gclk));
	jand g2599(.dina(w_n1551_0[1]),.dinb(w_n319_27[1]),.dout(n2862),.clk(gclk));
	jor g2600(.dina(n2862),.dinb(n2861),.dout(n2863),.clk(gclk));
	jand g2601(.dina(w_n1526_0[1]),.dinb(w_n265_27[1]),.dout(n2864),.clk(gclk));
	jor g2602(.dina(w_dff_B_49MrkuEv1_0),.dinb(n2863),.dout(n2865),.clk(gclk));
	jor g2603(.dina(n2865),.dinb(w_dff_B_r38PTKb32_1),.dout(n2866),.clk(gclk));
	jor g2604(.dina(w_n2866_0[1]),.dinb(w_n263_45[1]),.dout(n2867),.clk(gclk));
	jand g2605(.dina(w_n1515_0[1]),.dinb(w_n364_27[0]),.dout(n2868),.clk(gclk));
	jand g2606(.dina(w_n1498_0[1]),.dinb(w_n265_27[0]),.dout(n2869),.clk(gclk));
	jand g2607(.dina(w_n1542_0[1]),.dinb(w_n410_27[0]),.dout(n2870),.clk(gclk));
	jor g2608(.dina(n2870),.dinb(n2869),.dout(n2871),.clk(gclk));
	jand g2609(.dina(w_n1490_0[1]),.dinb(w_n319_27[0]),.dout(n2872),.clk(gclk));
	jor g2610(.dina(w_dff_B_FDc46lRH6_0),.dinb(n2871),.dout(n2873),.clk(gclk));
	jor g2611(.dina(n2873),.dinb(w_dff_B_3p3FQbxZ2_1),.dout(n2874),.clk(gclk));
	jor g2612(.dina(w_n2874_0[1]),.dinb(w_shift6_45[1]),.dout(n2875),.clk(gclk));
	jand g2613(.dina(n2875),.dinb(n2867),.dout(result54),.clk(gclk));
	jand g2614(.dina(w_n1579_0[1]),.dinb(w_n410_26[2]),.dout(n2877),.clk(gclk));
	jand g2615(.dina(w_n1615_0[1]),.dinb(w_n319_26[2]),.dout(n2878),.clk(gclk));
	jand g2616(.dina(w_n1599_0[1]),.dinb(w_n265_26[2]),.dout(n2879),.clk(gclk));
	jor g2617(.dina(n2879),.dinb(n2878),.dout(n2880),.clk(gclk));
	jand g2618(.dina(w_n1607_0[1]),.dinb(w_n364_26[2]),.dout(n2881),.clk(gclk));
	jor g2619(.dina(w_dff_B_hTzDDnzK8_0),.dinb(n2880),.dout(n2882),.clk(gclk));
	jor g2620(.dina(n2882),.dinb(w_dff_B_ZHHldruu7_1),.dout(n2883),.clk(gclk));
	jor g2621(.dina(w_n2883_0[1]),.dinb(w_n263_45[0]),.dout(n2884),.clk(gclk));
	jand g2622(.dina(w_n1571_0[1]),.dinb(w_n265_26[1]),.dout(n2885),.clk(gclk));
	jand g2623(.dina(w_n1563_0[1]),.dinb(w_n319_26[1]),.dout(n2886),.clk(gclk));
	jand g2624(.dina(w_n1624_0[1]),.dinb(w_n410_26[1]),.dout(n2887),.clk(gclk));
	jor g2625(.dina(n2887),.dinb(n2886),.dout(n2888),.clk(gclk));
	jand g2626(.dina(w_n1588_0[1]),.dinb(w_n364_26[1]),.dout(n2889),.clk(gclk));
	jor g2627(.dina(w_dff_B_D3k26w8o6_0),.dinb(n2888),.dout(n2890),.clk(gclk));
	jor g2628(.dina(n2890),.dinb(w_dff_B_ZRpp3rBP5_1),.dout(n2891),.clk(gclk));
	jor g2629(.dina(w_n2891_0[1]),.dinb(w_shift6_45[0]),.dout(n2892),.clk(gclk));
	jand g2630(.dina(n2892),.dinb(n2884),.dout(result55),.clk(gclk));
	jand g2631(.dina(w_n1680_0[1]),.dinb(w_n364_26[0]),.dout(n2894),.clk(gclk));
	jand g2632(.dina(w_n1697_0[1]),.dinb(w_n319_26[0]),.dout(n2895),.clk(gclk));
	jand g2633(.dina(w_n1672_0[1]),.dinb(w_n265_26[0]),.dout(n2896),.clk(gclk));
	jor g2634(.dina(n2896),.dinb(n2895),.dout(n2897),.clk(gclk));
	jand g2635(.dina(w_n1652_0[1]),.dinb(w_n410_26[0]),.dout(n2898),.clk(gclk));
	jor g2636(.dina(w_dff_B_ZGsJLjTO8_0),.dinb(n2897),.dout(n2899),.clk(gclk));
	jor g2637(.dina(n2899),.dinb(w_dff_B_ykEXxVEF6_1),.dout(n2900),.clk(gclk));
	jor g2638(.dina(w_n2900_0[1]),.dinb(w_n263_44[2]),.dout(n2901),.clk(gclk));
	jand g2639(.dina(w_n1688_0[1]),.dinb(w_n410_25[2]),.dout(n2902),.clk(gclk));
	jand g2640(.dina(w_n1636_0[1]),.dinb(w_n319_25[2]),.dout(n2903),.clk(gclk));
	jand g2641(.dina(w_n1644_0[1]),.dinb(w_n265_25[2]),.dout(n2904),.clk(gclk));
	jor g2642(.dina(n2904),.dinb(n2903),.dout(n2905),.clk(gclk));
	jand g2643(.dina(w_n1661_0[1]),.dinb(w_n364_25[2]),.dout(n2906),.clk(gclk));
	jor g2644(.dina(w_dff_B_c2phCQGi0_0),.dinb(n2905),.dout(n2907),.clk(gclk));
	jor g2645(.dina(n2907),.dinb(w_dff_B_lhOl7scJ0_1),.dout(n2908),.clk(gclk));
	jor g2646(.dina(w_n2908_0[1]),.dinb(w_shift6_44[2]),.dout(n2909),.clk(gclk));
	jand g2647(.dina(n2909),.dinb(n2901),.dout(result56),.clk(gclk));
	jand g2648(.dina(w_n1770_0[1]),.dinb(w_n265_25[1]),.dout(n2911),.clk(gclk));
	jand g2649(.dina(w_n1745_0[1]),.dinb(w_n319_25[1]),.dout(n2912),.clk(gclk));
	jand g2650(.dina(w_n1753_0[1]),.dinb(w_n364_25[1]),.dout(n2913),.clk(gclk));
	jor g2651(.dina(n2913),.dinb(n2912),.dout(n2914),.clk(gclk));
	jand g2652(.dina(w_n1709_0[1]),.dinb(w_n410_25[1]),.dout(n2915),.clk(gclk));
	jor g2653(.dina(w_dff_B_ZgZcwHQk4_0),.dinb(n2914),.dout(n2916),.clk(gclk));
	jor g2654(.dina(n2916),.dinb(w_dff_B_OZhIiuq18_1),.dout(n2917),.clk(gclk));
	jor g2655(.dina(w_n2917_0[1]),.dinb(w_n263_44[1]),.dout(n2918),.clk(gclk));
	jand g2656(.dina(w_n1717_0[1]),.dinb(w_n265_25[0]),.dout(n2919),.clk(gclk));
	jand g2657(.dina(w_n1725_0[1]),.dinb(w_n319_25[0]),.dout(n2920),.clk(gclk));
	jand g2658(.dina(w_n1761_0[1]),.dinb(w_n410_25[0]),.dout(n2921),.clk(gclk));
	jor g2659(.dina(n2921),.dinb(n2920),.dout(n2922),.clk(gclk));
	jand g2660(.dina(w_n1734_0[1]),.dinb(w_n364_25[0]),.dout(n2923),.clk(gclk));
	jor g2661(.dina(w_dff_B_PEtYO2nZ2_0),.dinb(n2922),.dout(n2924),.clk(gclk));
	jor g2662(.dina(n2924),.dinb(w_dff_B_Vexy9pSD4_1),.dout(n2925),.clk(gclk));
	jor g2663(.dina(w_n2925_0[1]),.dinb(w_shift6_44[1]),.dout(n2926),.clk(gclk));
	jand g2664(.dina(n2926),.dinb(n2918),.dout(result57),.clk(gclk));
	jand g2665(.dina(w_n1807_0[1]),.dinb(w_n410_24[2]),.dout(n2928),.clk(gclk));
	jand g2666(.dina(w_n1834_0[1]),.dinb(w_n319_24[2]),.dout(n2929),.clk(gclk));
	jand g2667(.dina(w_n1843_0[1]),.dinb(w_n265_24[2]),.dout(n2930),.clk(gclk));
	jor g2668(.dina(n2930),.dinb(n2929),.dout(n2931),.clk(gclk));
	jand g2669(.dina(w_n1826_0[1]),.dinb(w_n364_24[2]),.dout(n2932),.clk(gclk));
	jor g2670(.dina(w_dff_B_K2r8C8Bi4_0),.dinb(n2931),.dout(n2933),.clk(gclk));
	jor g2671(.dina(n2933),.dinb(w_dff_B_LOWVhPMa9_1),.dout(n2934),.clk(gclk));
	jor g2672(.dina(w_n2934_0[1]),.dinb(w_n263_44[0]),.dout(n2935),.clk(gclk));
	jand g2673(.dina(w_n1818_0[1]),.dinb(w_n410_24[1]),.dout(n2936),.clk(gclk));
	jand g2674(.dina(w_n1790_0[1]),.dinb(w_n265_24[1]),.dout(n2937),.clk(gclk));
	jand g2675(.dina(w_n1798_0[1]),.dinb(w_n319_24[1]),.dout(n2938),.clk(gclk));
	jor g2676(.dina(n2938),.dinb(n2937),.dout(n2939),.clk(gclk));
	jand g2677(.dina(w_n1782_0[1]),.dinb(w_n364_24[1]),.dout(n2940),.clk(gclk));
	jor g2678(.dina(w_dff_B_iXUqkg6b0_0),.dinb(n2939),.dout(n2941),.clk(gclk));
	jor g2679(.dina(n2941),.dinb(w_dff_B_ZIGeXFC22_1),.dout(n2942),.clk(gclk));
	jor g2680(.dina(w_n2942_0[1]),.dinb(w_shift6_44[0]),.dout(n2943),.clk(gclk));
	jand g2681(.dina(n2943),.dinb(n2935),.dout(result58),.clk(gclk));
	jand g2682(.dina(w_n1899_0[1]),.dinb(w_n364_24[0]),.dout(n2945),.clk(gclk));
	jand g2683(.dina(w_n1907_0[1]),.dinb(w_n319_24[0]),.dout(n2946),.clk(gclk));
	jand g2684(.dina(w_n1891_0[1]),.dinb(w_n265_24[0]),.dout(n2947),.clk(gclk));
	jor g2685(.dina(n2947),.dinb(n2946),.dout(n2948),.clk(gclk));
	jand g2686(.dina(w_n1880_0[1]),.dinb(w_n410_24[0]),.dout(n2949),.clk(gclk));
	jor g2687(.dina(w_dff_B_YljleBFN9_0),.dinb(n2948),.dout(n2950),.clk(gclk));
	jor g2688(.dina(n2950),.dinb(w_dff_B_ICBxgeIV7_1),.dout(n2951),.clk(gclk));
	jor g2689(.dina(w_n2951_0[1]),.dinb(w_n263_43[2]),.dout(n2952),.clk(gclk));
	jand g2690(.dina(w_n1871_0[1]),.dinb(w_n319_23[2]),.dout(n2953),.clk(gclk));
	jand g2691(.dina(w_n1863_0[1]),.dinb(w_n265_23[2]),.dout(n2954),.clk(gclk));
	jand g2692(.dina(w_n1916_0[1]),.dinb(w_n410_23[2]),.dout(n2955),.clk(gclk));
	jor g2693(.dina(n2955),.dinb(n2954),.dout(n2956),.clk(gclk));
	jand g2694(.dina(w_n1855_0[1]),.dinb(w_n364_23[2]),.dout(n2957),.clk(gclk));
	jor g2695(.dina(w_dff_B_qzNhIp991_0),.dinb(n2956),.dout(n2958),.clk(gclk));
	jor g2696(.dina(n2958),.dinb(w_dff_B_8sKYsfXN5_1),.dout(n2959),.clk(gclk));
	jor g2697(.dina(w_n2959_0[1]),.dinb(w_shift6_43[2]),.dout(n2960),.clk(gclk));
	jand g2698(.dina(n2960),.dinb(n2952),.dout(result59),.clk(gclk));
	jand g2699(.dina(w_n1989_0[1]),.dinb(w_n265_23[1]),.dout(n2962),.clk(gclk));
	jand g2700(.dina(w_n1980_0[1]),.dinb(w_n319_23[1]),.dout(n2963),.clk(gclk));
	jand g2701(.dina(w_n1972_0[1]),.dinb(w_n364_23[1]),.dout(n2964),.clk(gclk));
	jor g2702(.dina(n2964),.dinb(n2963),.dout(n2965),.clk(gclk));
	jand g2703(.dina(w_n1944_0[1]),.dinb(w_n410_23[1]),.dout(n2966),.clk(gclk));
	jor g2704(.dina(w_dff_B_vaIk44ui8_0),.dinb(n2965),.dout(n2967),.clk(gclk));
	jor g2705(.dina(n2967),.dinb(w_dff_B_NGb1Pgpk3_1),.dout(n2968),.clk(gclk));
	jor g2706(.dina(w_n2968_0[1]),.dinb(w_n263_43[1]),.dout(n2969),.clk(gclk));
	jand g2707(.dina(w_n1928_0[1]),.dinb(w_n319_23[0]),.dout(n2970),.clk(gclk));
	jand g2708(.dina(w_n1936_0[1]),.dinb(w_n265_23[0]),.dout(n2971),.clk(gclk));
	jand g2709(.dina(w_n1964_0[1]),.dinb(w_n410_23[0]),.dout(n2972),.clk(gclk));
	jor g2710(.dina(n2972),.dinb(n2971),.dout(n2973),.clk(gclk));
	jand g2711(.dina(w_n1953_0[1]),.dinb(w_n364_23[0]),.dout(n2974),.clk(gclk));
	jor g2712(.dina(w_dff_B_lnxYEnyW2_0),.dinb(n2973),.dout(n2975),.clk(gclk));
	jor g2713(.dina(n2975),.dinb(w_dff_B_BUCvsxNO3_1),.dout(n2976),.clk(gclk));
	jor g2714(.dina(w_n2976_0[1]),.dinb(w_shift6_43[1]),.dout(n2977),.clk(gclk));
	jand g2715(.dina(n2977),.dinb(n2969),.dout(result60),.clk(gclk));
	jand g2716(.dina(w_n2037_0[1]),.dinb(w_n265_22[2]),.dout(n2979),.clk(gclk));
	jand g2717(.dina(w_n2062_0[1]),.dinb(w_n319_22[2]),.dout(n2980),.clk(gclk));
	jand g2718(.dina(w_n2045_0[1]),.dinb(w_n364_22[2]),.dout(n2981),.clk(gclk));
	jor g2719(.dina(n2981),.dinb(n2980),.dout(n2982),.clk(gclk));
	jand g2720(.dina(w_n2017_0[1]),.dinb(w_n410_22[2]),.dout(n2983),.clk(gclk));
	jor g2721(.dina(w_dff_B_id4K03Wa5_0),.dinb(n2982),.dout(n2984),.clk(gclk));
	jor g2722(.dina(n2984),.dinb(w_dff_B_JqSHsLGG2_1),.dout(n2985),.clk(gclk));
	jor g2723(.dina(w_n2985_0[1]),.dinb(w_n263_43[0]),.dout(n2986),.clk(gclk));
	jand g2724(.dina(w_n2026_0[1]),.dinb(w_n364_22[1]),.dout(n2987),.clk(gclk));
	jand g2725(.dina(w_n2009_0[1]),.dinb(w_n265_22[1]),.dout(n2988),.clk(gclk));
	jand g2726(.dina(w_n2053_0[1]),.dinb(w_n410_22[1]),.dout(n2989),.clk(gclk));
	jor g2727(.dina(n2989),.dinb(n2988),.dout(n2990),.clk(gclk));
	jand g2728(.dina(w_n2001_0[1]),.dinb(w_n319_22[1]),.dout(n2991),.clk(gclk));
	jor g2729(.dina(w_dff_B_mNvo9h4e6_0),.dinb(n2990),.dout(n2992),.clk(gclk));
	jor g2730(.dina(n2992),.dinb(w_dff_B_MNkhRkVJ2_1),.dout(n2993),.clk(gclk));
	jor g2731(.dina(w_n2993_0[1]),.dinb(w_shift6_43[0]),.dout(n2994),.clk(gclk));
	jand g2732(.dina(n2994),.dinb(n2986),.dout(result61),.clk(gclk));
	jand g2733(.dina(w_n2118_0[1]),.dinb(w_n364_22[0]),.dout(n2996),.clk(gclk));
	jand g2734(.dina(w_n2110_0[1]),.dinb(w_n319_22[0]),.dout(n2997),.clk(gclk));
	jand g2735(.dina(w_n2135_0[1]),.dinb(w_n265_22[0]),.dout(n2998),.clk(gclk));
	jor g2736(.dina(n2998),.dinb(n2997),.dout(n2999),.clk(gclk));
	jand g2737(.dina(w_n2090_0[1]),.dinb(w_n410_22[0]),.dout(n3000),.clk(gclk));
	jor g2738(.dina(w_dff_B_m0Sng1PW4_0),.dinb(n2999),.dout(n3001),.clk(gclk));
	jor g2739(.dina(n3001),.dinb(w_dff_B_yEJJMF8P9_1),.dout(n3002),.clk(gclk));
	jor g2740(.dina(w_n3002_0[1]),.dinb(w_n263_42[2]),.dout(n3003),.clk(gclk));
	jand g2741(.dina(w_n2126_0[1]),.dinb(w_n410_21[2]),.dout(n3004),.clk(gclk));
	jand g2742(.dina(w_n2082_0[1]),.dinb(w_n265_21[2]),.dout(n3005),.clk(gclk));
	jand g2743(.dina(w_n2099_0[1]),.dinb(w_n319_21[2]),.dout(n3006),.clk(gclk));
	jor g2744(.dina(n3006),.dinb(n3005),.dout(n3007),.clk(gclk));
	jand g2745(.dina(w_n2074_0[1]),.dinb(w_n364_21[2]),.dout(n3008),.clk(gclk));
	jor g2746(.dina(w_dff_B_hIuzRHwv3_0),.dinb(n3007),.dout(n3009),.clk(gclk));
	jor g2747(.dina(n3009),.dinb(w_dff_B_kUjye1l65_1),.dout(n3010),.clk(gclk));
	jor g2748(.dina(w_n3010_0[1]),.dinb(w_shift6_42[2]),.dout(n3011),.clk(gclk));
	jand g2749(.dina(n3011),.dinb(n3003),.dout(result62),.clk(gclk));
	jand g2750(.dina(w_n2191_0[1]),.dinb(w_n364_21[1]),.dout(n3013),.clk(gclk));
	jand g2751(.dina(w_n2199_0[1]),.dinb(w_n319_21[1]),.dout(n3014),.clk(gclk));
	jand g2752(.dina(w_n2208_0[1]),.dinb(w_n265_21[1]),.dout(n3015),.clk(gclk));
	jor g2753(.dina(n3015),.dinb(n3014),.dout(n3016),.clk(gclk));
	jand g2754(.dina(w_n2172_0[1]),.dinb(w_n410_21[1]),.dout(n3017),.clk(gclk));
	jor g2755(.dina(w_dff_B_b2g877Zq9_0),.dinb(n3016),.dout(n3018),.clk(gclk));
	jor g2756(.dina(n3018),.dinb(w_dff_B_qIVWh7nJ2_1),.dout(n3019),.clk(gclk));
	jor g2757(.dina(w_n3019_0[1]),.dinb(w_n263_42[1]),.dout(n3020),.clk(gclk));
	jand g2758(.dina(w_n2147_0[1]),.dinb(w_n364_21[0]),.dout(n3021),.clk(gclk));
	jand g2759(.dina(w_n2155_0[1]),.dinb(w_n265_21[0]),.dout(n3022),.clk(gclk));
	jand g2760(.dina(w_n2183_0[1]),.dinb(w_n410_21[0]),.dout(n3023),.clk(gclk));
	jor g2761(.dina(n3023),.dinb(n3022),.dout(n3024),.clk(gclk));
	jand g2762(.dina(w_n2163_0[1]),.dinb(w_n319_21[0]),.dout(n3025),.clk(gclk));
	jor g2763(.dina(w_dff_B_ClAbqRb96_0),.dinb(n3024),.dout(n3026),.clk(gclk));
	jor g2764(.dina(n3026),.dinb(w_dff_B_o6DVcVCt5_1),.dout(n3027),.clk(gclk));
	jor g2765(.dina(w_n3027_0[1]),.dinb(w_shift6_42[1]),.dout(n3028),.clk(gclk));
	jand g2766(.dina(n3028),.dinb(n3020),.dout(result63),.clk(gclk));
	jor g2767(.dina(w_n636_0[0]),.dinb(w_n263_42[0]),.dout(n3030),.clk(gclk));
	jor g2768(.dina(w_n456_0[0]),.dinb(w_shift6_42[0]),.dout(n3031),.clk(gclk));
	jand g2769(.dina(n3031),.dinb(n3030),.dout(result64),.clk(gclk));
	jor g2770(.dina(w_n997_0[0]),.dinb(w_n263_41[2]),.dout(n3033),.clk(gclk));
	jor g2771(.dina(w_n817_0[0]),.dinb(w_shift6_41[2]),.dout(n3034),.clk(gclk));
	jand g2772(.dina(n3034),.dinb(n3033),.dout(result65),.clk(gclk));
	jor g2773(.dina(w_n1166_0[0]),.dinb(w_n263_41[1]),.dout(n3036),.clk(gclk));
	jor g2774(.dina(w_n1082_0[0]),.dinb(w_shift6_41[1]),.dout(n3037),.clk(gclk));
	jand g2775(.dina(n3037),.dinb(n3036),.dout(result66),.clk(gclk));
	jor g2776(.dina(w_n1335_0[0]),.dinb(w_n263_41[0]),.dout(n3039),.clk(gclk));
	jor g2777(.dina(w_n1251_0[0]),.dinb(w_shift6_41[0]),.dout(n3040),.clk(gclk));
	jand g2778(.dina(n3040),.dinb(n3039),.dout(result67),.clk(gclk));
	jor g2779(.dina(w_n1408_0[0]),.dinb(w_n263_40[2]),.dout(n3042),.clk(gclk));
	jor g2780(.dina(w_n1372_0[0]),.dinb(w_shift6_40[2]),.dout(n3043),.clk(gclk));
	jand g2781(.dina(n3043),.dinb(n3042),.dout(result68),.clk(gclk));
	jor g2782(.dina(w_n1481_0[0]),.dinb(w_n263_40[1]),.dout(n3045),.clk(gclk));
	jor g2783(.dina(w_n1445_0[0]),.dinb(w_shift6_40[1]),.dout(n3046),.clk(gclk));
	jand g2784(.dina(n3046),.dinb(n3045),.dout(result69),.clk(gclk));
	jor g2785(.dina(w_n1554_0[0]),.dinb(w_n263_40[0]),.dout(n3048),.clk(gclk));
	jor g2786(.dina(w_n1518_0[0]),.dinb(w_shift6_40[0]),.dout(n3049),.clk(gclk));
	jand g2787(.dina(n3049),.dinb(n3048),.dout(result70),.clk(gclk));
	jor g2788(.dina(w_n1627_0[0]),.dinb(w_n263_39[2]),.dout(n3051),.clk(gclk));
	jor g2789(.dina(w_n1591_0[0]),.dinb(w_shift6_39[2]),.dout(n3052),.clk(gclk));
	jand g2790(.dina(n3052),.dinb(n3051),.dout(result71),.clk(gclk));
	jor g2791(.dina(w_n1700_0[0]),.dinb(w_n263_39[1]),.dout(n3054),.clk(gclk));
	jor g2792(.dina(w_n1664_0[0]),.dinb(w_shift6_39[1]),.dout(n3055),.clk(gclk));
	jand g2793(.dina(n3055),.dinb(n3054),.dout(result72),.clk(gclk));
	jor g2794(.dina(w_n1773_0[0]),.dinb(w_n263_39[0]),.dout(n3057),.clk(gclk));
	jor g2795(.dina(w_n1737_0[0]),.dinb(w_shift6_39[0]),.dout(n3058),.clk(gclk));
	jand g2796(.dina(n3058),.dinb(n3057),.dout(result73),.clk(gclk));
	jor g2797(.dina(w_n1846_0[0]),.dinb(w_n263_38[2]),.dout(n3060),.clk(gclk));
	jor g2798(.dina(w_n1810_0[0]),.dinb(w_shift6_38[2]),.dout(n3061),.clk(gclk));
	jand g2799(.dina(n3061),.dinb(n3060),.dout(result74),.clk(gclk));
	jor g2800(.dina(w_n1919_0[0]),.dinb(w_n263_38[1]),.dout(n3063),.clk(gclk));
	jor g2801(.dina(w_n1883_0[0]),.dinb(w_shift6_38[1]),.dout(n3064),.clk(gclk));
	jand g2802(.dina(n3064),.dinb(n3063),.dout(result75),.clk(gclk));
	jor g2803(.dina(w_n1992_0[0]),.dinb(w_n263_38[0]),.dout(n3066),.clk(gclk));
	jor g2804(.dina(w_n1956_0[0]),.dinb(w_shift6_38[0]),.dout(n3067),.clk(gclk));
	jand g2805(.dina(n3067),.dinb(n3066),.dout(result76),.clk(gclk));
	jor g2806(.dina(w_n2065_0[0]),.dinb(w_n263_37[2]),.dout(n3069),.clk(gclk));
	jor g2807(.dina(w_n2029_0[0]),.dinb(w_shift6_37[2]),.dout(n3070),.clk(gclk));
	jand g2808(.dina(n3070),.dinb(n3069),.dout(result77),.clk(gclk));
	jor g2809(.dina(w_n2138_0[0]),.dinb(w_n263_37[1]),.dout(n3072),.clk(gclk));
	jor g2810(.dina(w_n2102_0[0]),.dinb(w_shift6_37[1]),.dout(n3073),.clk(gclk));
	jand g2811(.dina(n3073),.dinb(n3072),.dout(result78),.clk(gclk));
	jor g2812(.dina(w_n2211_0[0]),.dinb(w_n263_37[0]),.dout(n3075),.clk(gclk));
	jor g2813(.dina(w_n2175_0[0]),.dinb(w_shift6_37[0]),.dout(n3076),.clk(gclk));
	jand g2814(.dina(n3076),.dinb(n3075),.dout(result79),.clk(gclk));
	jor g2815(.dina(w_n2228_0[0]),.dinb(w_n263_36[2]),.dout(n3078),.clk(gclk));
	jor g2816(.dina(w_n2220_0[0]),.dinb(w_shift6_36[2]),.dout(n3079),.clk(gclk));
	jand g2817(.dina(n3079),.dinb(n3078),.dout(result80),.clk(gclk));
	jor g2818(.dina(w_n2245_0[0]),.dinb(w_n263_36[1]),.dout(n3081),.clk(gclk));
	jor g2819(.dina(w_n2237_0[0]),.dinb(w_shift6_36[1]),.dout(n3082),.clk(gclk));
	jand g2820(.dina(n3082),.dinb(n3081),.dout(result81),.clk(gclk));
	jor g2821(.dina(w_n2262_0[0]),.dinb(w_n263_36[0]),.dout(n3084),.clk(gclk));
	jor g2822(.dina(w_n2254_0[0]),.dinb(w_shift6_36[0]),.dout(n3085),.clk(gclk));
	jand g2823(.dina(n3085),.dinb(n3084),.dout(result82),.clk(gclk));
	jor g2824(.dina(w_n2279_0[0]),.dinb(w_n263_35[2]),.dout(n3087),.clk(gclk));
	jor g2825(.dina(w_n2271_0[0]),.dinb(w_shift6_35[2]),.dout(n3088),.clk(gclk));
	jand g2826(.dina(n3088),.dinb(n3087),.dout(result83),.clk(gclk));
	jor g2827(.dina(w_n2296_0[0]),.dinb(w_n263_35[1]),.dout(n3090),.clk(gclk));
	jor g2828(.dina(w_n2288_0[0]),.dinb(w_shift6_35[1]),.dout(n3091),.clk(gclk));
	jand g2829(.dina(n3091),.dinb(n3090),.dout(result84),.clk(gclk));
	jor g2830(.dina(w_n2313_0[0]),.dinb(w_n263_35[0]),.dout(n3093),.clk(gclk));
	jor g2831(.dina(w_n2305_0[0]),.dinb(w_shift6_35[0]),.dout(n3094),.clk(gclk));
	jand g2832(.dina(n3094),.dinb(n3093),.dout(result85),.clk(gclk));
	jor g2833(.dina(w_n2330_0[0]),.dinb(w_n263_34[2]),.dout(n3096),.clk(gclk));
	jor g2834(.dina(w_n2322_0[0]),.dinb(w_shift6_34[2]),.dout(n3097),.clk(gclk));
	jand g2835(.dina(n3097),.dinb(n3096),.dout(result86),.clk(gclk));
	jor g2836(.dina(w_n2347_0[0]),.dinb(w_n263_34[1]),.dout(n3099),.clk(gclk));
	jor g2837(.dina(w_n2339_0[0]),.dinb(w_shift6_34[1]),.dout(n3100),.clk(gclk));
	jand g2838(.dina(n3100),.dinb(n3099),.dout(result87),.clk(gclk));
	jor g2839(.dina(w_n2364_0[0]),.dinb(w_n263_34[0]),.dout(n3102),.clk(gclk));
	jor g2840(.dina(w_n2356_0[0]),.dinb(w_shift6_34[0]),.dout(n3103),.clk(gclk));
	jand g2841(.dina(n3103),.dinb(n3102),.dout(result88),.clk(gclk));
	jor g2842(.dina(w_n2381_0[0]),.dinb(w_n263_33[2]),.dout(n3105),.clk(gclk));
	jor g2843(.dina(w_n2373_0[0]),.dinb(w_shift6_33[2]),.dout(n3106),.clk(gclk));
	jand g2844(.dina(n3106),.dinb(n3105),.dout(result89),.clk(gclk));
	jor g2845(.dina(w_n2398_0[0]),.dinb(w_n263_33[1]),.dout(n3108),.clk(gclk));
	jor g2846(.dina(w_n2390_0[0]),.dinb(w_shift6_33[1]),.dout(n3109),.clk(gclk));
	jand g2847(.dina(n3109),.dinb(n3108),.dout(result90),.clk(gclk));
	jor g2848(.dina(w_n2415_0[0]),.dinb(w_n263_33[0]),.dout(n3111),.clk(gclk));
	jor g2849(.dina(w_n2407_0[0]),.dinb(w_shift6_33[0]),.dout(n3112),.clk(gclk));
	jand g2850(.dina(n3112),.dinb(n3111),.dout(result91),.clk(gclk));
	jor g2851(.dina(w_n2432_0[0]),.dinb(w_n263_32[2]),.dout(n3114),.clk(gclk));
	jor g2852(.dina(w_n2424_0[0]),.dinb(w_shift6_32[2]),.dout(n3115),.clk(gclk));
	jand g2853(.dina(n3115),.dinb(n3114),.dout(result92),.clk(gclk));
	jor g2854(.dina(w_n2449_0[0]),.dinb(w_n263_32[1]),.dout(n3117),.clk(gclk));
	jor g2855(.dina(w_n2441_0[0]),.dinb(w_shift6_32[1]),.dout(n3118),.clk(gclk));
	jand g2856(.dina(n3118),.dinb(n3117),.dout(result93),.clk(gclk));
	jor g2857(.dina(w_n2466_0[0]),.dinb(w_n263_32[0]),.dout(n3120),.clk(gclk));
	jor g2858(.dina(w_n2458_0[0]),.dinb(w_shift6_32[0]),.dout(n3121),.clk(gclk));
	jand g2859(.dina(n3121),.dinb(n3120),.dout(result94),.clk(gclk));
	jor g2860(.dina(w_n2483_0[0]),.dinb(w_n263_31[2]),.dout(n3123),.clk(gclk));
	jor g2861(.dina(w_n2475_0[0]),.dinb(w_shift6_31[2]),.dout(n3124),.clk(gclk));
	jand g2862(.dina(n3124),.dinb(n3123),.dout(result95),.clk(gclk));
	jor g2863(.dina(w_n2500_0[0]),.dinb(w_n263_31[1]),.dout(n3126),.clk(gclk));
	jor g2864(.dina(w_n2492_0[0]),.dinb(w_shift6_31[1]),.dout(n3127),.clk(gclk));
	jand g2865(.dina(n3127),.dinb(n3126),.dout(result96),.clk(gclk));
	jor g2866(.dina(w_n2517_0[0]),.dinb(w_n263_31[0]),.dout(n3129),.clk(gclk));
	jor g2867(.dina(w_n2509_0[0]),.dinb(w_shift6_31[0]),.dout(n3130),.clk(gclk));
	jand g2868(.dina(n3130),.dinb(n3129),.dout(result97),.clk(gclk));
	jor g2869(.dina(w_n2534_0[0]),.dinb(w_n263_30[2]),.dout(n3132),.clk(gclk));
	jor g2870(.dina(w_n2526_0[0]),.dinb(w_shift6_30[2]),.dout(n3133),.clk(gclk));
	jand g2871(.dina(n3133),.dinb(n3132),.dout(result98),.clk(gclk));
	jor g2872(.dina(w_n2551_0[0]),.dinb(w_n263_30[1]),.dout(n3135),.clk(gclk));
	jor g2873(.dina(w_n2543_0[0]),.dinb(w_shift6_30[1]),.dout(n3136),.clk(gclk));
	jand g2874(.dina(n3136),.dinb(n3135),.dout(result99),.clk(gclk));
	jor g2875(.dina(w_n2568_0[0]),.dinb(w_n263_30[0]),.dout(n3138),.clk(gclk));
	jor g2876(.dina(w_n2560_0[0]),.dinb(w_shift6_30[0]),.dout(n3139),.clk(gclk));
	jand g2877(.dina(n3139),.dinb(n3138),.dout(result100),.clk(gclk));
	jor g2878(.dina(w_n2585_0[0]),.dinb(w_n263_29[2]),.dout(n3141),.clk(gclk));
	jor g2879(.dina(w_n2577_0[0]),.dinb(w_shift6_29[2]),.dout(n3142),.clk(gclk));
	jand g2880(.dina(n3142),.dinb(n3141),.dout(result101),.clk(gclk));
	jor g2881(.dina(w_n2602_0[0]),.dinb(w_n263_29[1]),.dout(n3144),.clk(gclk));
	jor g2882(.dina(w_n2594_0[0]),.dinb(w_shift6_29[1]),.dout(n3145),.clk(gclk));
	jand g2883(.dina(n3145),.dinb(n3144),.dout(result102),.clk(gclk));
	jor g2884(.dina(w_n2619_0[0]),.dinb(w_n263_29[0]),.dout(n3147),.clk(gclk));
	jor g2885(.dina(w_n2611_0[0]),.dinb(w_shift6_29[0]),.dout(n3148),.clk(gclk));
	jand g2886(.dina(n3148),.dinb(n3147),.dout(result103),.clk(gclk));
	jor g2887(.dina(w_n2636_0[0]),.dinb(w_n263_28[2]),.dout(n3150),.clk(gclk));
	jor g2888(.dina(w_n2628_0[0]),.dinb(w_shift6_28[2]),.dout(n3151),.clk(gclk));
	jand g2889(.dina(n3151),.dinb(n3150),.dout(result104),.clk(gclk));
	jor g2890(.dina(w_n2653_0[0]),.dinb(w_n263_28[1]),.dout(n3153),.clk(gclk));
	jor g2891(.dina(w_n2645_0[0]),.dinb(w_shift6_28[1]),.dout(n3154),.clk(gclk));
	jand g2892(.dina(n3154),.dinb(n3153),.dout(result105),.clk(gclk));
	jor g2893(.dina(w_n2670_0[0]),.dinb(w_n263_28[0]),.dout(n3156),.clk(gclk));
	jor g2894(.dina(w_n2662_0[0]),.dinb(w_shift6_28[0]),.dout(n3157),.clk(gclk));
	jand g2895(.dina(n3157),.dinb(n3156),.dout(result106),.clk(gclk));
	jor g2896(.dina(w_n2687_0[0]),.dinb(w_n263_27[2]),.dout(n3159),.clk(gclk));
	jor g2897(.dina(w_n2679_0[0]),.dinb(w_shift6_27[2]),.dout(n3160),.clk(gclk));
	jand g2898(.dina(n3160),.dinb(n3159),.dout(result107),.clk(gclk));
	jor g2899(.dina(w_n2704_0[0]),.dinb(w_n263_27[1]),.dout(n3162),.clk(gclk));
	jor g2900(.dina(w_n2696_0[0]),.dinb(w_shift6_27[1]),.dout(n3163),.clk(gclk));
	jand g2901(.dina(n3163),.dinb(n3162),.dout(result108),.clk(gclk));
	jor g2902(.dina(w_n2721_0[0]),.dinb(w_n263_27[0]),.dout(n3165),.clk(gclk));
	jor g2903(.dina(w_n2713_0[0]),.dinb(w_shift6_27[0]),.dout(n3166),.clk(gclk));
	jand g2904(.dina(n3166),.dinb(n3165),.dout(result109),.clk(gclk));
	jor g2905(.dina(w_n2738_0[0]),.dinb(w_n263_26[2]),.dout(n3168),.clk(gclk));
	jor g2906(.dina(w_n2730_0[0]),.dinb(w_shift6_26[2]),.dout(n3169),.clk(gclk));
	jand g2907(.dina(n3169),.dinb(n3168),.dout(result110),.clk(gclk));
	jor g2908(.dina(w_n2755_0[0]),.dinb(w_n263_26[1]),.dout(n3171),.clk(gclk));
	jor g2909(.dina(w_n2747_0[0]),.dinb(w_shift6_26[1]),.dout(n3172),.clk(gclk));
	jand g2910(.dina(n3172),.dinb(n3171),.dout(result111),.clk(gclk));
	jor g2911(.dina(w_n2772_0[0]),.dinb(w_n263_26[0]),.dout(n3174),.clk(gclk));
	jor g2912(.dina(w_n2764_0[0]),.dinb(w_shift6_26[0]),.dout(n3175),.clk(gclk));
	jand g2913(.dina(n3175),.dinb(n3174),.dout(result112),.clk(gclk));
	jor g2914(.dina(w_n2789_0[0]),.dinb(w_n263_25[2]),.dout(n3177),.clk(gclk));
	jor g2915(.dina(w_n2781_0[0]),.dinb(w_shift6_25[2]),.dout(n3178),.clk(gclk));
	jand g2916(.dina(n3178),.dinb(n3177),.dout(result113),.clk(gclk));
	jor g2917(.dina(w_n2806_0[0]),.dinb(w_n263_25[1]),.dout(n3180),.clk(gclk));
	jor g2918(.dina(w_n2798_0[0]),.dinb(w_shift6_25[1]),.dout(n3181),.clk(gclk));
	jand g2919(.dina(n3181),.dinb(n3180),.dout(result114),.clk(gclk));
	jor g2920(.dina(w_n2823_0[0]),.dinb(w_n263_25[0]),.dout(n3183),.clk(gclk));
	jor g2921(.dina(w_n2815_0[0]),.dinb(w_shift6_25[0]),.dout(n3184),.clk(gclk));
	jand g2922(.dina(n3184),.dinb(n3183),.dout(result115),.clk(gclk));
	jor g2923(.dina(w_n2840_0[0]),.dinb(w_n263_24[2]),.dout(n3186),.clk(gclk));
	jor g2924(.dina(w_n2832_0[0]),.dinb(w_shift6_24[2]),.dout(n3187),.clk(gclk));
	jand g2925(.dina(n3187),.dinb(n3186),.dout(result116),.clk(gclk));
	jor g2926(.dina(w_n2857_0[0]),.dinb(w_n263_24[1]),.dout(n3189),.clk(gclk));
	jor g2927(.dina(w_n2849_0[0]),.dinb(w_shift6_24[1]),.dout(n3190),.clk(gclk));
	jand g2928(.dina(n3190),.dinb(n3189),.dout(result117),.clk(gclk));
	jor g2929(.dina(w_n2874_0[0]),.dinb(w_n263_24[0]),.dout(n3192),.clk(gclk));
	jor g2930(.dina(w_n2866_0[0]),.dinb(w_shift6_24[0]),.dout(n3193),.clk(gclk));
	jand g2931(.dina(n3193),.dinb(n3192),.dout(result118),.clk(gclk));
	jor g2932(.dina(w_n2891_0[0]),.dinb(w_n263_23[2]),.dout(n3195),.clk(gclk));
	jor g2933(.dina(w_n2883_0[0]),.dinb(w_shift6_23[2]),.dout(n3196),.clk(gclk));
	jand g2934(.dina(n3196),.dinb(n3195),.dout(result119),.clk(gclk));
	jor g2935(.dina(w_n2908_0[0]),.dinb(w_n263_23[1]),.dout(n3198),.clk(gclk));
	jor g2936(.dina(w_n2900_0[0]),.dinb(w_shift6_23[1]),.dout(n3199),.clk(gclk));
	jand g2937(.dina(n3199),.dinb(n3198),.dout(result120),.clk(gclk));
	jor g2938(.dina(w_n2925_0[0]),.dinb(w_n263_23[0]),.dout(n3201),.clk(gclk));
	jor g2939(.dina(w_n2917_0[0]),.dinb(w_shift6_23[0]),.dout(n3202),.clk(gclk));
	jand g2940(.dina(n3202),.dinb(n3201),.dout(result121),.clk(gclk));
	jor g2941(.dina(w_n2942_0[0]),.dinb(w_n263_22[2]),.dout(n3204),.clk(gclk));
	jor g2942(.dina(w_n2934_0[0]),.dinb(w_shift6_22[2]),.dout(n3205),.clk(gclk));
	jand g2943(.dina(n3205),.dinb(n3204),.dout(result122),.clk(gclk));
	jor g2944(.dina(w_n2959_0[0]),.dinb(w_n263_22[1]),.dout(n3207),.clk(gclk));
	jor g2945(.dina(w_n2951_0[0]),.dinb(w_shift6_22[1]),.dout(n3208),.clk(gclk));
	jand g2946(.dina(n3208),.dinb(n3207),.dout(result123),.clk(gclk));
	jor g2947(.dina(w_n2976_0[0]),.dinb(w_n263_22[0]),.dout(n3210),.clk(gclk));
	jor g2948(.dina(w_n2968_0[0]),.dinb(w_shift6_22[0]),.dout(n3211),.clk(gclk));
	jand g2949(.dina(n3211),.dinb(n3210),.dout(result124),.clk(gclk));
	jor g2950(.dina(w_n2993_0[0]),.dinb(w_n263_21[2]),.dout(n3213),.clk(gclk));
	jor g2951(.dina(w_n2985_0[0]),.dinb(w_shift6_21[2]),.dout(n3214),.clk(gclk));
	jand g2952(.dina(n3214),.dinb(n3213),.dout(result125),.clk(gclk));
	jor g2953(.dina(w_n3010_0[0]),.dinb(w_n263_21[1]),.dout(n3216),.clk(gclk));
	jor g2954(.dina(w_n3002_0[0]),.dinb(w_shift6_21[1]),.dout(n3217),.clk(gclk));
	jand g2955(.dina(n3217),.dinb(n3216),.dout(result126),.clk(gclk));
	jor g2956(.dina(w_n3027_0[0]),.dinb(w_n263_21[0]),.dout(n3219),.clk(gclk));
	jor g2957(.dina(w_n3019_0[0]),.dinb(w_shift6_21[0]),.dout(n3220),.clk(gclk));
	jand g2958(.dina(n3220),.dinb(n3219),.dout(result127),.clk(gclk));
	jspl jspl_w_a0_0(.douta(w_dff_A_g47baKUj6_0),.doutb(w_a0_0[1]),.din(a0));
	jspl jspl_w_a1_0(.douta(w_a1_0[0]),.doutb(w_dff_A_2LdNMFjs0_1),.din(a1));
	jspl jspl_w_a2_0(.douta(w_dff_A_JozpVLIs7_0),.doutb(w_a2_0[1]),.din(a2));
	jspl jspl_w_a3_0(.douta(w_a3_0[0]),.doutb(w_dff_A_P7ahRfJd1_1),.din(a3));
	jspl jspl_w_a4_0(.douta(w_dff_A_V7FH9gfr3_0),.doutb(w_a4_0[1]),.din(a4));
	jspl jspl_w_a5_0(.douta(w_a5_0[0]),.doutb(w_dff_A_IhAADU2o4_1),.din(a5));
	jspl jspl_w_a6_0(.douta(w_dff_A_5wvWWH0g3_0),.doutb(w_a6_0[1]),.din(a6));
	jspl jspl_w_a7_0(.douta(w_a7_0[0]),.doutb(w_dff_A_2ewe9RPU2_1),.din(a7));
	jspl jspl_w_a8_0(.douta(w_dff_A_JPoE7RgR9_0),.doutb(w_a8_0[1]),.din(a8));
	jspl jspl_w_a9_0(.douta(w_a9_0[0]),.doutb(w_dff_A_KS7aaRbG4_1),.din(a9));
	jspl jspl_w_a10_0(.douta(w_dff_A_rcrknBQy7_0),.doutb(w_a10_0[1]),.din(a10));
	jspl jspl_w_a11_0(.douta(w_a11_0[0]),.doutb(w_dff_A_PUmUpuIX0_1),.din(a11));
	jspl jspl_w_a12_0(.douta(w_dff_A_vcWxBCo84_0),.doutb(w_a12_0[1]),.din(a12));
	jspl jspl_w_a13_0(.douta(w_a13_0[0]),.doutb(w_dff_A_n7nis0rM6_1),.din(a13));
	jspl jspl_w_a14_0(.douta(w_dff_A_aZ8WAfFs3_0),.doutb(w_a14_0[1]),.din(a14));
	jspl jspl_w_a15_0(.douta(w_a15_0[0]),.doutb(w_dff_A_jaLZbcNB9_1),.din(a15));
	jspl jspl_w_a16_0(.douta(w_dff_A_6rr88UQ06_0),.doutb(w_a16_0[1]),.din(a16));
	jspl jspl_w_a17_0(.douta(w_a17_0[0]),.doutb(w_dff_A_IjOIf2Vv3_1),.din(a17));
	jspl jspl_w_a18_0(.douta(w_dff_A_HqaVWGpG4_0),.doutb(w_a18_0[1]),.din(a18));
	jspl jspl_w_a19_0(.douta(w_a19_0[0]),.doutb(w_dff_A_EfquT9R57_1),.din(a19));
	jspl jspl_w_a20_0(.douta(w_dff_A_z9RlMpd06_0),.doutb(w_a20_0[1]),.din(a20));
	jspl jspl_w_a21_0(.douta(w_a21_0[0]),.doutb(w_dff_A_OrPlTNw66_1),.din(a21));
	jspl jspl_w_a22_0(.douta(w_dff_A_ypOJA4Mn4_0),.doutb(w_a22_0[1]),.din(a22));
	jspl jspl_w_a23_0(.douta(w_a23_0[0]),.doutb(w_dff_A_ECU7ndwr9_1),.din(a23));
	jspl jspl_w_a24_0(.douta(w_dff_A_JsBVmPGJ3_0),.doutb(w_a24_0[1]),.din(a24));
	jspl jspl_w_a25_0(.douta(w_a25_0[0]),.doutb(w_dff_A_LpS4cIVI1_1),.din(a25));
	jspl jspl_w_a26_0(.douta(w_dff_A_FL8rfjir2_0),.doutb(w_a26_0[1]),.din(a26));
	jspl jspl_w_a27_0(.douta(w_a27_0[0]),.doutb(w_dff_A_7GZZbsWq5_1),.din(a27));
	jspl jspl_w_a28_0(.douta(w_dff_A_ixqoCv1I6_0),.doutb(w_a28_0[1]),.din(a28));
	jspl jspl_w_a29_0(.douta(w_a29_0[0]),.doutb(w_dff_A_AvFtfhSE5_1),.din(a29));
	jspl jspl_w_a30_0(.douta(w_dff_A_yNeInT2q0_0),.doutb(w_a30_0[1]),.din(a30));
	jspl jspl_w_a31_0(.douta(w_a31_0[0]),.doutb(w_dff_A_yjHZSHH70_1),.din(a31));
	jspl jspl_w_a32_0(.douta(w_dff_A_wkaxuBD72_0),.doutb(w_a32_0[1]),.din(a32));
	jspl jspl_w_a33_0(.douta(w_a33_0[0]),.doutb(w_dff_A_7OB6oRqA1_1),.din(a33));
	jspl jspl_w_a34_0(.douta(w_dff_A_4hVRVXx43_0),.doutb(w_a34_0[1]),.din(a34));
	jspl jspl_w_a35_0(.douta(w_a35_0[0]),.doutb(w_dff_A_IeX7m3QI0_1),.din(a35));
	jspl jspl_w_a36_0(.douta(w_dff_A_O8Ze6Upb1_0),.doutb(w_a36_0[1]),.din(a36));
	jspl jspl_w_a37_0(.douta(w_a37_0[0]),.doutb(w_dff_A_Z0uMSCcz9_1),.din(a37));
	jspl jspl_w_a38_0(.douta(w_dff_A_we9q0Jad5_0),.doutb(w_a38_0[1]),.din(a38));
	jspl jspl_w_a39_0(.douta(w_a39_0[0]),.doutb(w_dff_A_VjN2Qliq0_1),.din(a39));
	jspl jspl_w_a40_0(.douta(w_dff_A_Dkax2EMe2_0),.doutb(w_a40_0[1]),.din(a40));
	jspl jspl_w_a41_0(.douta(w_a41_0[0]),.doutb(w_dff_A_qtRk7Icw0_1),.din(a41));
	jspl jspl_w_a42_0(.douta(w_dff_A_VKlsC5cZ2_0),.doutb(w_a42_0[1]),.din(a42));
	jspl jspl_w_a43_0(.douta(w_a43_0[0]),.doutb(w_dff_A_Wwy7IlhU6_1),.din(a43));
	jspl jspl_w_a44_0(.douta(w_dff_A_hUN70b8y2_0),.doutb(w_a44_0[1]),.din(a44));
	jspl jspl_w_a45_0(.douta(w_a45_0[0]),.doutb(w_dff_A_dUrA3tEd2_1),.din(a45));
	jspl jspl_w_a46_0(.douta(w_dff_A_XF2Yyt4V5_0),.doutb(w_a46_0[1]),.din(a46));
	jspl jspl_w_a47_0(.douta(w_a47_0[0]),.doutb(w_dff_A_bTr2Cfs06_1),.din(a47));
	jspl jspl_w_a48_0(.douta(w_dff_A_x9iScKCA1_0),.doutb(w_a48_0[1]),.din(a48));
	jspl jspl_w_a49_0(.douta(w_a49_0[0]),.doutb(w_dff_A_mAgVgHU16_1),.din(a49));
	jspl jspl_w_a50_0(.douta(w_dff_A_qerx9cuT9_0),.doutb(w_a50_0[1]),.din(a50));
	jspl jspl_w_a51_0(.douta(w_a51_0[0]),.doutb(w_dff_A_MCBIUaBq2_1),.din(a51));
	jspl jspl_w_a52_0(.douta(w_dff_A_TEmwG3XJ6_0),.doutb(w_a52_0[1]),.din(a52));
	jspl jspl_w_a53_0(.douta(w_a53_0[0]),.doutb(w_dff_A_r5bZU0Yn6_1),.din(a53));
	jspl jspl_w_a54_0(.douta(w_dff_A_xNYvrMCm0_0),.doutb(w_a54_0[1]),.din(a54));
	jspl jspl_w_a55_0(.douta(w_a55_0[0]),.doutb(w_dff_A_0nnYYHF55_1),.din(a55));
	jspl jspl_w_a56_0(.douta(w_dff_A_Nsc29slm7_0),.doutb(w_a56_0[1]),.din(a56));
	jspl jspl_w_a57_0(.douta(w_a57_0[0]),.doutb(w_dff_A_S63Jgp8X2_1),.din(a57));
	jspl jspl_w_a58_0(.douta(w_dff_A_AY4LJMyP2_0),.doutb(w_a58_0[1]),.din(a58));
	jspl jspl_w_a59_0(.douta(w_a59_0[0]),.doutb(w_dff_A_td3IjRBo8_1),.din(a59));
	jspl jspl_w_a60_0(.douta(w_dff_A_ruJEv85L7_0),.doutb(w_a60_0[1]),.din(a60));
	jspl jspl_w_a61_0(.douta(w_a61_0[0]),.doutb(w_dff_A_zbNXoOqW6_1),.din(a61));
	jspl jspl_w_a62_0(.douta(w_dff_A_HmdqNm8g4_0),.doutb(w_a62_0[1]),.din(a62));
	jspl jspl_w_a63_0(.douta(w_a63_0[0]),.doutb(w_dff_A_8mgBZIQg7_1),.din(a63));
	jspl jspl_w_a64_0(.douta(w_dff_A_ipr72ra02_0),.doutb(w_a64_0[1]),.din(a64));
	jspl jspl_w_a65_0(.douta(w_a65_0[0]),.doutb(w_dff_A_APWgC3dM4_1),.din(a65));
	jspl jspl_w_a66_0(.douta(w_dff_A_aYzwVtdH1_0),.doutb(w_a66_0[1]),.din(a66));
	jspl jspl_w_a67_0(.douta(w_a67_0[0]),.doutb(w_dff_A_9PjzwdE12_1),.din(a67));
	jspl jspl_w_a68_0(.douta(w_dff_A_SwhSpGG03_0),.doutb(w_a68_0[1]),.din(a68));
	jspl jspl_w_a69_0(.douta(w_a69_0[0]),.doutb(w_dff_A_yYiuMmAx6_1),.din(a69));
	jspl jspl_w_a70_0(.douta(w_dff_A_bhAqClr40_0),.doutb(w_a70_0[1]),.din(a70));
	jspl jspl_w_a71_0(.douta(w_a71_0[0]),.doutb(w_dff_A_qYdmnUej7_1),.din(a71));
	jspl jspl_w_a72_0(.douta(w_dff_A_3gOkgdes3_0),.doutb(w_a72_0[1]),.din(a72));
	jspl jspl_w_a73_0(.douta(w_a73_0[0]),.doutb(w_dff_A_tD9nMY0t2_1),.din(a73));
	jspl jspl_w_a74_0(.douta(w_dff_A_I7gyfdFq9_0),.doutb(w_a74_0[1]),.din(a74));
	jspl jspl_w_a75_0(.douta(w_a75_0[0]),.doutb(w_dff_A_NA9ziZSD5_1),.din(a75));
	jspl jspl_w_a76_0(.douta(w_dff_A_jsqcgtqV5_0),.doutb(w_a76_0[1]),.din(a76));
	jspl jspl_w_a77_0(.douta(w_a77_0[0]),.doutb(w_dff_A_Tf7v1fro5_1),.din(a77));
	jspl jspl_w_a78_0(.douta(w_dff_A_4pYXSgZQ4_0),.doutb(w_a78_0[1]),.din(a78));
	jspl jspl_w_a79_0(.douta(w_a79_0[0]),.doutb(w_dff_A_eOY9af3E1_1),.din(a79));
	jspl jspl_w_a80_0(.douta(w_dff_A_FxenSOIp9_0),.doutb(w_a80_0[1]),.din(a80));
	jspl jspl_w_a81_0(.douta(w_a81_0[0]),.doutb(w_dff_A_X1Lfnzwj8_1),.din(a81));
	jspl jspl_w_a82_0(.douta(w_dff_A_wSYwKQKp9_0),.doutb(w_a82_0[1]),.din(a82));
	jspl jspl_w_a83_0(.douta(w_a83_0[0]),.doutb(w_dff_A_OiMf06K86_1),.din(a83));
	jspl jspl_w_a84_0(.douta(w_dff_A_i8HqUX7H4_0),.doutb(w_a84_0[1]),.din(a84));
	jspl jspl_w_a85_0(.douta(w_a85_0[0]),.doutb(w_dff_A_OcSdyoQr6_1),.din(a85));
	jspl jspl_w_a86_0(.douta(w_dff_A_5fD5AaYw7_0),.doutb(w_a86_0[1]),.din(a86));
	jspl jspl_w_a87_0(.douta(w_a87_0[0]),.doutb(w_dff_A_TrlnadzK5_1),.din(a87));
	jspl jspl_w_a88_0(.douta(w_dff_A_nt5Btme91_0),.doutb(w_a88_0[1]),.din(a88));
	jspl jspl_w_a89_0(.douta(w_a89_0[0]),.doutb(w_dff_A_uSzz6U2s7_1),.din(a89));
	jspl jspl_w_a90_0(.douta(w_dff_A_p4g9Yx0Z8_0),.doutb(w_a90_0[1]),.din(a90));
	jspl jspl_w_a91_0(.douta(w_a91_0[0]),.doutb(w_dff_A_OxxYjRfR3_1),.din(a91));
	jspl jspl_w_a92_0(.douta(w_dff_A_8B97r3VV0_0),.doutb(w_a92_0[1]),.din(a92));
	jspl jspl_w_a93_0(.douta(w_a93_0[0]),.doutb(w_dff_A_RTG96NZT0_1),.din(a93));
	jspl jspl_w_a94_0(.douta(w_dff_A_Xt1EtlJu1_0),.doutb(w_a94_0[1]),.din(a94));
	jspl jspl_w_a95_0(.douta(w_a95_0[0]),.doutb(w_dff_A_Pe361rYG6_1),.din(a95));
	jspl jspl_w_a96_0(.douta(w_dff_A_HbBmurSs9_0),.doutb(w_a96_0[1]),.din(a96));
	jspl jspl_w_a97_0(.douta(w_a97_0[0]),.doutb(w_dff_A_3E0UAqQJ7_1),.din(a97));
	jspl jspl_w_a98_0(.douta(w_dff_A_4h0NH7LH3_0),.doutb(w_a98_0[1]),.din(a98));
	jspl jspl_w_a99_0(.douta(w_a99_0[0]),.doutb(w_dff_A_amGWYNxX5_1),.din(a99));
	jspl jspl_w_a100_0(.douta(w_dff_A_tioEWBSH6_0),.doutb(w_a100_0[1]),.din(a100));
	jspl jspl_w_a101_0(.douta(w_a101_0[0]),.doutb(w_dff_A_iMM7uM3x0_1),.din(a101));
	jspl jspl_w_a102_0(.douta(w_dff_A_x1m5wCkQ3_0),.doutb(w_a102_0[1]),.din(a102));
	jspl jspl_w_a103_0(.douta(w_a103_0[0]),.doutb(w_dff_A_fFCBlUt64_1),.din(a103));
	jspl jspl_w_a104_0(.douta(w_dff_A_KWIu5I4M0_0),.doutb(w_a104_0[1]),.din(a104));
	jspl jspl_w_a105_0(.douta(w_a105_0[0]),.doutb(w_dff_A_NhWoqlJE7_1),.din(a105));
	jspl jspl_w_a106_0(.douta(w_dff_A_BB5cJRhF0_0),.doutb(w_a106_0[1]),.din(a106));
	jspl jspl_w_a107_0(.douta(w_a107_0[0]),.doutb(w_dff_A_x0WLNzz69_1),.din(a107));
	jspl jspl_w_a108_0(.douta(w_dff_A_3R8e6hTN0_0),.doutb(w_a108_0[1]),.din(a108));
	jspl jspl_w_a109_0(.douta(w_a109_0[0]),.doutb(w_dff_A_nyGrOAiO3_1),.din(a109));
	jspl jspl_w_a110_0(.douta(w_dff_A_a4SNezFT6_0),.doutb(w_a110_0[1]),.din(a110));
	jspl jspl_w_a111_0(.douta(w_a111_0[0]),.doutb(w_dff_A_bbcJxZ647_1),.din(a111));
	jspl jspl_w_a112_0(.douta(w_dff_A_aqMYVpgr1_0),.doutb(w_a112_0[1]),.din(a112));
	jspl jspl_w_a113_0(.douta(w_a113_0[0]),.doutb(w_dff_A_bKqOvwAI6_1),.din(a113));
	jspl jspl_w_a114_0(.douta(w_dff_A_RGJo87rH1_0),.doutb(w_a114_0[1]),.din(a114));
	jspl jspl_w_a115_0(.douta(w_a115_0[0]),.doutb(w_dff_A_4GIKWQI35_1),.din(a115));
	jspl jspl_w_a116_0(.douta(w_dff_A_aEQEN3Xf2_0),.doutb(w_a116_0[1]),.din(a116));
	jspl jspl_w_a117_0(.douta(w_a117_0[0]),.doutb(w_dff_A_vTXKnj262_1),.din(a117));
	jspl jspl_w_a118_0(.douta(w_dff_A_lRhC755p2_0),.doutb(w_a118_0[1]),.din(a118));
	jspl jspl_w_a119_0(.douta(w_a119_0[0]),.doutb(w_dff_A_ECSpmsBT6_1),.din(a119));
	jspl jspl_w_a120_0(.douta(w_dff_A_kGWQUzm74_0),.doutb(w_a120_0[1]),.din(a120));
	jspl jspl_w_a121_0(.douta(w_a121_0[0]),.doutb(w_dff_A_q0xtfwdX5_1),.din(a121));
	jspl jspl_w_a122_0(.douta(w_dff_A_SKaaili94_0),.doutb(w_a122_0[1]),.din(a122));
	jspl jspl_w_a123_0(.douta(w_a123_0[0]),.doutb(w_dff_A_nSHI3wrB2_1),.din(a123));
	jspl jspl_w_a124_0(.douta(w_dff_A_qYADieKW4_0),.doutb(w_a124_0[1]),.din(a124));
	jspl jspl_w_a125_0(.douta(w_a125_0[0]),.doutb(w_dff_A_p4ahpbAJ4_1),.din(a125));
	jspl jspl_w_a126_0(.douta(w_dff_A_2Aq7vbmA8_0),.doutb(w_a126_0[1]),.din(a126));
	jspl jspl_w_a127_0(.douta(w_a127_0[0]),.doutb(w_dff_A_OqgJmqtR1_1),.din(a127));
	jspl3 jspl3_w_shift0_0(.douta(w_shift0_0[0]),.doutb(w_shift0_0[1]),.doutc(w_shift0_0[2]),.din(shift0));
	jspl3 jspl3_w_shift0_1(.douta(w_shift0_1[0]),.doutb(w_shift0_1[1]),.doutc(w_shift0_1[2]),.din(w_shift0_0[0]));
	jspl3 jspl3_w_shift0_2(.douta(w_shift0_2[0]),.doutb(w_shift0_2[1]),.doutc(w_shift0_2[2]),.din(w_shift0_0[1]));
	jspl3 jspl3_w_shift0_3(.douta(w_shift0_3[0]),.doutb(w_shift0_3[1]),.doutc(w_shift0_3[2]),.din(w_shift0_0[2]));
	jspl3 jspl3_w_shift0_4(.douta(w_shift0_4[0]),.doutb(w_shift0_4[1]),.doutc(w_shift0_4[2]),.din(w_shift0_1[0]));
	jspl3 jspl3_w_shift0_5(.douta(w_shift0_5[0]),.doutb(w_shift0_5[1]),.doutc(w_shift0_5[2]),.din(w_shift0_1[1]));
	jspl3 jspl3_w_shift0_6(.douta(w_shift0_6[0]),.doutb(w_shift0_6[1]),.doutc(w_shift0_6[2]),.din(w_shift0_1[2]));
	jspl3 jspl3_w_shift0_7(.douta(w_shift0_7[0]),.doutb(w_shift0_7[1]),.doutc(w_shift0_7[2]),.din(w_shift0_2[0]));
	jspl3 jspl3_w_shift0_8(.douta(w_shift0_8[0]),.doutb(w_shift0_8[1]),.doutc(w_shift0_8[2]),.din(w_shift0_2[1]));
	jspl3 jspl3_w_shift0_9(.douta(w_shift0_9[0]),.doutb(w_shift0_9[1]),.doutc(w_shift0_9[2]),.din(w_shift0_2[2]));
	jspl3 jspl3_w_shift0_10(.douta(w_shift0_10[0]),.doutb(w_shift0_10[1]),.doutc(w_shift0_10[2]),.din(w_shift0_3[0]));
	jspl3 jspl3_w_shift0_11(.douta(w_shift0_11[0]),.doutb(w_shift0_11[1]),.doutc(w_shift0_11[2]),.din(w_shift0_3[1]));
	jspl3 jspl3_w_shift0_12(.douta(w_shift0_12[0]),.doutb(w_shift0_12[1]),.doutc(w_shift0_12[2]),.din(w_shift0_3[2]));
	jspl3 jspl3_w_shift0_13(.douta(w_shift0_13[0]),.doutb(w_shift0_13[1]),.doutc(w_shift0_13[2]),.din(w_shift0_4[0]));
	jspl3 jspl3_w_shift0_14(.douta(w_shift0_14[0]),.doutb(w_shift0_14[1]),.doutc(w_shift0_14[2]),.din(w_shift0_4[1]));
	jspl3 jspl3_w_shift0_15(.douta(w_shift0_15[0]),.doutb(w_shift0_15[1]),.doutc(w_shift0_15[2]),.din(w_shift0_4[2]));
	jspl3 jspl3_w_shift0_16(.douta(w_shift0_16[0]),.doutb(w_shift0_16[1]),.doutc(w_shift0_16[2]),.din(w_shift0_5[0]));
	jspl3 jspl3_w_shift0_17(.douta(w_shift0_17[0]),.doutb(w_shift0_17[1]),.doutc(w_shift0_17[2]),.din(w_shift0_5[1]));
	jspl3 jspl3_w_shift0_18(.douta(w_shift0_18[0]),.doutb(w_shift0_18[1]),.doutc(w_shift0_18[2]),.din(w_shift0_5[2]));
	jspl3 jspl3_w_shift0_19(.douta(w_shift0_19[0]),.doutb(w_shift0_19[1]),.doutc(w_shift0_19[2]),.din(w_shift0_6[0]));
	jspl3 jspl3_w_shift0_20(.douta(w_shift0_20[0]),.doutb(w_shift0_20[1]),.doutc(w_shift0_20[2]),.din(w_shift0_6[1]));
	jspl3 jspl3_w_shift0_21(.douta(w_shift0_21[0]),.doutb(w_shift0_21[1]),.doutc(w_shift0_21[2]),.din(w_shift0_6[2]));
	jspl3 jspl3_w_shift0_22(.douta(w_shift0_22[0]),.doutb(w_shift0_22[1]),.doutc(w_shift0_22[2]),.din(w_shift0_7[0]));
	jspl3 jspl3_w_shift0_23(.douta(w_shift0_23[0]),.doutb(w_shift0_23[1]),.doutc(w_shift0_23[2]),.din(w_shift0_7[1]));
	jspl3 jspl3_w_shift0_24(.douta(w_shift0_24[0]),.doutb(w_shift0_24[1]),.doutc(w_shift0_24[2]),.din(w_shift0_7[2]));
	jspl3 jspl3_w_shift0_25(.douta(w_shift0_25[0]),.doutb(w_shift0_25[1]),.doutc(w_shift0_25[2]),.din(w_shift0_8[0]));
	jspl3 jspl3_w_shift0_26(.douta(w_shift0_26[0]),.doutb(w_shift0_26[1]),.doutc(w_shift0_26[2]),.din(w_shift0_8[1]));
	jspl3 jspl3_w_shift0_27(.douta(w_shift0_27[0]),.doutb(w_shift0_27[1]),.doutc(w_shift0_27[2]),.din(w_shift0_8[2]));
	jspl3 jspl3_w_shift0_28(.douta(w_shift0_28[0]),.doutb(w_shift0_28[1]),.doutc(w_shift0_28[2]),.din(w_shift0_9[0]));
	jspl3 jspl3_w_shift0_29(.douta(w_shift0_29[0]),.doutb(w_shift0_29[1]),.doutc(w_shift0_29[2]),.din(w_shift0_9[1]));
	jspl3 jspl3_w_shift0_30(.douta(w_shift0_30[0]),.doutb(w_shift0_30[1]),.doutc(w_shift0_30[2]),.din(w_shift0_9[2]));
	jspl3 jspl3_w_shift0_31(.douta(w_shift0_31[0]),.doutb(w_shift0_31[1]),.doutc(w_shift0_31[2]),.din(w_shift0_10[0]));
	jspl3 jspl3_w_shift0_32(.douta(w_shift0_32[0]),.doutb(w_shift0_32[1]),.doutc(w_shift0_32[2]),.din(w_shift0_10[1]));
	jspl3 jspl3_w_shift0_33(.douta(w_shift0_33[0]),.doutb(w_shift0_33[1]),.doutc(w_shift0_33[2]),.din(w_shift0_10[2]));
	jspl3 jspl3_w_shift0_34(.douta(w_shift0_34[0]),.doutb(w_shift0_34[1]),.doutc(w_shift0_34[2]),.din(w_shift0_11[0]));
	jspl3 jspl3_w_shift0_35(.douta(w_shift0_35[0]),.doutb(w_shift0_35[1]),.doutc(w_shift0_35[2]),.din(w_shift0_11[1]));
	jspl3 jspl3_w_shift0_36(.douta(w_shift0_36[0]),.doutb(w_shift0_36[1]),.doutc(w_shift0_36[2]),.din(w_shift0_11[2]));
	jspl3 jspl3_w_shift0_37(.douta(w_shift0_37[0]),.doutb(w_shift0_37[1]),.doutc(w_shift0_37[2]),.din(w_shift0_12[0]));
	jspl3 jspl3_w_shift0_38(.douta(w_shift0_38[0]),.doutb(w_shift0_38[1]),.doutc(w_shift0_38[2]),.din(w_shift0_12[1]));
	jspl3 jspl3_w_shift0_39(.douta(w_shift0_39[0]),.doutb(w_shift0_39[1]),.doutc(w_shift0_39[2]),.din(w_shift0_12[2]));
	jspl3 jspl3_w_shift0_40(.douta(w_shift0_40[0]),.doutb(w_shift0_40[1]),.doutc(w_shift0_40[2]),.din(w_shift0_13[0]));
	jspl3 jspl3_w_shift0_41(.douta(w_shift0_41[0]),.doutb(w_shift0_41[1]),.doutc(w_shift0_41[2]),.din(w_shift0_13[1]));
	jspl3 jspl3_w_shift0_42(.douta(w_shift0_42[0]),.doutb(w_shift0_42[1]),.doutc(w_shift0_42[2]),.din(w_shift0_13[2]));
	jspl3 jspl3_w_shift0_43(.douta(w_shift0_43[0]),.doutb(w_shift0_43[1]),.doutc(w_shift0_43[2]),.din(w_shift0_14[0]));
	jspl3 jspl3_w_shift0_44(.douta(w_shift0_44[0]),.doutb(w_shift0_44[1]),.doutc(w_shift0_44[2]),.din(w_shift0_14[1]));
	jspl3 jspl3_w_shift0_45(.douta(w_shift0_45[0]),.doutb(w_shift0_45[1]),.doutc(w_shift0_45[2]),.din(w_shift0_14[2]));
	jspl3 jspl3_w_shift0_46(.douta(w_shift0_46[0]),.doutb(w_shift0_46[1]),.doutc(w_shift0_46[2]),.din(w_shift0_15[0]));
	jspl3 jspl3_w_shift0_47(.douta(w_shift0_47[0]),.doutb(w_shift0_47[1]),.doutc(w_shift0_47[2]),.din(w_shift0_15[1]));
	jspl3 jspl3_w_shift0_48(.douta(w_shift0_48[0]),.doutb(w_shift0_48[1]),.doutc(w_shift0_48[2]),.din(w_shift0_15[2]));
	jspl3 jspl3_w_shift0_49(.douta(w_shift0_49[0]),.doutb(w_shift0_49[1]),.doutc(w_shift0_49[2]),.din(w_shift0_16[0]));
	jspl3 jspl3_w_shift0_50(.douta(w_shift0_50[0]),.doutb(w_shift0_50[1]),.doutc(w_shift0_50[2]),.din(w_shift0_16[1]));
	jspl3 jspl3_w_shift0_51(.douta(w_shift0_51[0]),.doutb(w_shift0_51[1]),.doutc(w_shift0_51[2]),.din(w_shift0_16[2]));
	jspl3 jspl3_w_shift0_52(.douta(w_shift0_52[0]),.doutb(w_shift0_52[1]),.doutc(w_shift0_52[2]),.din(w_shift0_17[0]));
	jspl3 jspl3_w_shift0_53(.douta(w_shift0_53[0]),.doutb(w_shift0_53[1]),.doutc(w_shift0_53[2]),.din(w_shift0_17[1]));
	jspl3 jspl3_w_shift0_54(.douta(w_shift0_54[0]),.doutb(w_shift0_54[1]),.doutc(w_shift0_54[2]),.din(w_shift0_17[2]));
	jspl3 jspl3_w_shift0_55(.douta(w_shift0_55[0]),.doutb(w_shift0_55[1]),.doutc(w_shift0_55[2]),.din(w_shift0_18[0]));
	jspl3 jspl3_w_shift0_56(.douta(w_shift0_56[0]),.doutb(w_shift0_56[1]),.doutc(w_shift0_56[2]),.din(w_shift0_18[1]));
	jspl3 jspl3_w_shift0_57(.douta(w_shift0_57[0]),.doutb(w_shift0_57[1]),.doutc(w_shift0_57[2]),.din(w_shift0_18[2]));
	jspl3 jspl3_w_shift0_58(.douta(w_shift0_58[0]),.doutb(w_shift0_58[1]),.doutc(w_shift0_58[2]),.din(w_shift0_19[0]));
	jspl3 jspl3_w_shift0_59(.douta(w_shift0_59[0]),.doutb(w_shift0_59[1]),.doutc(w_shift0_59[2]),.din(w_shift0_19[1]));
	jspl3 jspl3_w_shift0_60(.douta(w_shift0_60[0]),.doutb(w_shift0_60[1]),.doutc(w_shift0_60[2]),.din(w_shift0_19[2]));
	jspl3 jspl3_w_shift0_61(.douta(w_shift0_61[0]),.doutb(w_shift0_61[1]),.doutc(w_shift0_61[2]),.din(w_shift0_20[0]));
	jspl3 jspl3_w_shift0_62(.douta(w_shift0_62[0]),.doutb(w_shift0_62[1]),.doutc(w_shift0_62[2]),.din(w_shift0_20[1]));
	jspl3 jspl3_w_shift0_63(.douta(w_shift0_63[0]),.doutb(w_shift0_63[1]),.doutc(w_shift0_63[2]),.din(w_shift0_20[2]));
	jspl3 jspl3_w_shift1_0(.douta(w_shift1_0[0]),.doutb(w_dff_A_2auC8Ory6_1),.doutc(w_dff_A_ewMNBLer3_2),.din(shift1));
	jspl3 jspl3_w_shift1_1(.douta(w_dff_A_VLfOiBZL1_0),.doutb(w_dff_A_LfupF43K8_1),.doutc(w_shift1_1[2]),.din(w_shift1_0[0]));
	jspl3 jspl3_w_shift1_2(.douta(w_shift1_2[0]),.doutb(w_shift1_2[1]),.doutc(w_shift1_2[2]),.din(w_shift1_0[1]));
	jspl3 jspl3_w_shift1_3(.douta(w_shift1_3[0]),.doutb(w_shift1_3[1]),.doutc(w_shift1_3[2]),.din(w_shift1_0[2]));
	jspl3 jspl3_w_shift1_4(.douta(w_shift1_4[0]),.doutb(w_shift1_4[1]),.doutc(w_shift1_4[2]),.din(w_shift1_1[0]));
	jspl3 jspl3_w_shift1_5(.douta(w_shift1_5[0]),.doutb(w_shift1_5[1]),.doutc(w_shift1_5[2]),.din(w_shift1_1[1]));
	jspl3 jspl3_w_shift1_6(.douta(w_dff_A_imsCNVkT2_0),.doutb(w_shift1_6[1]),.doutc(w_dff_A_mDIUIck97_2),.din(w_shift1_1[2]));
	jspl3 jspl3_w_shift1_7(.douta(w_shift1_7[0]),.doutb(w_shift1_7[1]),.doutc(w_shift1_7[2]),.din(w_shift1_2[0]));
	jspl3 jspl3_w_shift1_8(.douta(w_shift1_8[0]),.doutb(w_shift1_8[1]),.doutc(w_shift1_8[2]),.din(w_shift1_2[1]));
	jspl3 jspl3_w_shift1_9(.douta(w_shift1_9[0]),.doutb(w_shift1_9[1]),.doutc(w_shift1_9[2]),.din(w_shift1_2[2]));
	jspl3 jspl3_w_shift1_10(.douta(w_shift1_10[0]),.doutb(w_shift1_10[1]),.doutc(w_shift1_10[2]),.din(w_shift1_3[0]));
	jspl3 jspl3_w_shift1_11(.douta(w_shift1_11[0]),.doutb(w_shift1_11[1]),.doutc(w_shift1_11[2]),.din(w_shift1_3[1]));
	jspl3 jspl3_w_shift1_12(.douta(w_shift1_12[0]),.doutb(w_shift1_12[1]),.doutc(w_shift1_12[2]),.din(w_shift1_3[2]));
	jspl3 jspl3_w_shift1_13(.douta(w_shift1_13[0]),.doutb(w_shift1_13[1]),.doutc(w_shift1_13[2]),.din(w_shift1_4[0]));
	jspl3 jspl3_w_shift1_14(.douta(w_shift1_14[0]),.doutb(w_shift1_14[1]),.doutc(w_shift1_14[2]),.din(w_shift1_4[1]));
	jspl3 jspl3_w_shift1_15(.douta(w_shift1_15[0]),.doutb(w_shift1_15[1]),.doutc(w_shift1_15[2]),.din(w_shift1_4[2]));
	jspl3 jspl3_w_shift1_16(.douta(w_shift1_16[0]),.doutb(w_shift1_16[1]),.doutc(w_shift1_16[2]),.din(w_shift1_5[0]));
	jspl3 jspl3_w_shift1_17(.douta(w_shift1_17[0]),.doutb(w_shift1_17[1]),.doutc(w_shift1_17[2]),.din(w_shift1_5[1]));
	jspl3 jspl3_w_shift1_18(.douta(w_shift1_18[0]),.doutb(w_shift1_18[1]),.doutc(w_shift1_18[2]),.din(w_shift1_5[2]));
	jspl3 jspl3_w_shift1_19(.douta(w_shift1_19[0]),.doutb(w_shift1_19[1]),.doutc(w_shift1_19[2]),.din(w_shift1_6[0]));
	jspl3 jspl3_w_shift1_20(.douta(w_dff_A_9kI7kVaC9_0),.doutb(w_dff_A_rtDyqCOd8_1),.doutc(w_shift1_20[2]),.din(w_shift1_6[1]));
	jspl3 jspl3_w_shift1_21(.douta(w_shift1_21[0]),.doutb(w_shift1_21[1]),.doutc(w_shift1_21[2]),.din(w_shift1_6[2]));
	jspl3 jspl3_w_shift1_22(.douta(w_shift1_22[0]),.doutb(w_shift1_22[1]),.doutc(w_shift1_22[2]),.din(w_shift1_7[0]));
	jspl3 jspl3_w_shift1_23(.douta(w_shift1_23[0]),.doutb(w_shift1_23[1]),.doutc(w_shift1_23[2]),.din(w_shift1_7[1]));
	jspl3 jspl3_w_shift1_24(.douta(w_shift1_24[0]),.doutb(w_shift1_24[1]),.doutc(w_shift1_24[2]),.din(w_shift1_7[2]));
	jspl3 jspl3_w_shift1_25(.douta(w_shift1_25[0]),.doutb(w_shift1_25[1]),.doutc(w_shift1_25[2]),.din(w_shift1_8[0]));
	jspl3 jspl3_w_shift1_26(.douta(w_shift1_26[0]),.doutb(w_shift1_26[1]),.doutc(w_shift1_26[2]),.din(w_shift1_8[1]));
	jspl3 jspl3_w_shift1_27(.douta(w_shift1_27[0]),.doutb(w_shift1_27[1]),.doutc(w_shift1_27[2]),.din(w_shift1_8[2]));
	jspl3 jspl3_w_shift1_28(.douta(w_shift1_28[0]),.doutb(w_shift1_28[1]),.doutc(w_shift1_28[2]),.din(w_shift1_9[0]));
	jspl3 jspl3_w_shift1_29(.douta(w_shift1_29[0]),.doutb(w_shift1_29[1]),.doutc(w_shift1_29[2]),.din(w_shift1_9[1]));
	jspl3 jspl3_w_shift1_30(.douta(w_shift1_30[0]),.doutb(w_shift1_30[1]),.doutc(w_shift1_30[2]),.din(w_shift1_9[2]));
	jspl3 jspl3_w_shift1_31(.douta(w_shift1_31[0]),.doutb(w_shift1_31[1]),.doutc(w_shift1_31[2]),.din(w_shift1_10[0]));
	jspl3 jspl3_w_shift1_32(.douta(w_shift1_32[0]),.doutb(w_shift1_32[1]),.doutc(w_shift1_32[2]),.din(w_shift1_10[1]));
	jspl3 jspl3_w_shift1_33(.douta(w_shift1_33[0]),.doutb(w_shift1_33[1]),.doutc(w_shift1_33[2]),.din(w_shift1_10[2]));
	jspl3 jspl3_w_shift1_34(.douta(w_shift1_34[0]),.doutb(w_shift1_34[1]),.doutc(w_shift1_34[2]),.din(w_shift1_11[0]));
	jspl3 jspl3_w_shift1_35(.douta(w_shift1_35[0]),.doutb(w_shift1_35[1]),.doutc(w_shift1_35[2]),.din(w_shift1_11[1]));
	jspl3 jspl3_w_shift1_36(.douta(w_shift1_36[0]),.doutb(w_shift1_36[1]),.doutc(w_shift1_36[2]),.din(w_shift1_11[2]));
	jspl3 jspl3_w_shift1_37(.douta(w_shift1_37[0]),.doutb(w_shift1_37[1]),.doutc(w_shift1_37[2]),.din(w_shift1_12[0]));
	jspl3 jspl3_w_shift1_38(.douta(w_shift1_38[0]),.doutb(w_shift1_38[1]),.doutc(w_shift1_38[2]),.din(w_shift1_12[1]));
	jspl3 jspl3_w_shift1_39(.douta(w_shift1_39[0]),.doutb(w_shift1_39[1]),.doutc(w_shift1_39[2]),.din(w_shift1_12[2]));
	jspl3 jspl3_w_shift1_40(.douta(w_shift1_40[0]),.doutb(w_shift1_40[1]),.doutc(w_shift1_40[2]),.din(w_shift1_13[0]));
	jspl3 jspl3_w_shift1_41(.douta(w_shift1_41[0]),.doutb(w_shift1_41[1]),.doutc(w_shift1_41[2]),.din(w_shift1_13[1]));
	jspl3 jspl3_w_shift1_42(.douta(w_shift1_42[0]),.doutb(w_shift1_42[1]),.doutc(w_shift1_42[2]),.din(w_shift1_13[2]));
	jspl3 jspl3_w_shift1_43(.douta(w_shift1_43[0]),.doutb(w_shift1_43[1]),.doutc(w_shift1_43[2]),.din(w_shift1_14[0]));
	jspl3 jspl3_w_shift1_44(.douta(w_shift1_44[0]),.doutb(w_shift1_44[1]),.doutc(w_shift1_44[2]),.din(w_shift1_14[1]));
	jspl3 jspl3_w_shift1_45(.douta(w_shift1_45[0]),.doutb(w_shift1_45[1]),.doutc(w_shift1_45[2]),.din(w_shift1_14[2]));
	jspl3 jspl3_w_shift1_46(.douta(w_shift1_46[0]),.doutb(w_shift1_46[1]),.doutc(w_shift1_46[2]),.din(w_shift1_15[0]));
	jspl3 jspl3_w_shift1_47(.douta(w_shift1_47[0]),.doutb(w_shift1_47[1]),.doutc(w_shift1_47[2]),.din(w_shift1_15[1]));
	jspl3 jspl3_w_shift1_48(.douta(w_shift1_48[0]),.doutb(w_shift1_48[1]),.doutc(w_shift1_48[2]),.din(w_shift1_15[2]));
	jspl3 jspl3_w_shift1_49(.douta(w_shift1_49[0]),.doutb(w_shift1_49[1]),.doutc(w_shift1_49[2]),.din(w_shift1_16[0]));
	jspl3 jspl3_w_shift1_50(.douta(w_shift1_50[0]),.doutb(w_shift1_50[1]),.doutc(w_shift1_50[2]),.din(w_shift1_16[1]));
	jspl3 jspl3_w_shift1_51(.douta(w_shift1_51[0]),.doutb(w_shift1_51[1]),.doutc(w_shift1_51[2]),.din(w_shift1_16[2]));
	jspl3 jspl3_w_shift1_52(.douta(w_shift1_52[0]),.doutb(w_shift1_52[1]),.doutc(w_shift1_52[2]),.din(w_shift1_17[0]));
	jspl3 jspl3_w_shift1_53(.douta(w_shift1_53[0]),.doutb(w_shift1_53[1]),.doutc(w_shift1_53[2]),.din(w_shift1_17[1]));
	jspl3 jspl3_w_shift1_54(.douta(w_shift1_54[0]),.doutb(w_shift1_54[1]),.doutc(w_shift1_54[2]),.din(w_shift1_17[2]));
	jspl3 jspl3_w_shift1_55(.douta(w_shift1_55[0]),.doutb(w_shift1_55[1]),.doutc(w_shift1_55[2]),.din(w_shift1_18[0]));
	jspl3 jspl3_w_shift1_56(.douta(w_shift1_56[0]),.doutb(w_shift1_56[1]),.doutc(w_shift1_56[2]),.din(w_shift1_18[1]));
	jspl3 jspl3_w_shift1_57(.douta(w_shift1_57[0]),.doutb(w_shift1_57[1]),.doutc(w_shift1_57[2]),.din(w_shift1_18[2]));
	jspl3 jspl3_w_shift1_58(.douta(w_shift1_58[0]),.doutb(w_shift1_58[1]),.doutc(w_shift1_58[2]),.din(w_shift1_19[0]));
	jspl3 jspl3_w_shift1_59(.douta(w_shift1_59[0]),.doutb(w_shift1_59[1]),.doutc(w_shift1_59[2]),.din(w_shift1_19[1]));
	jspl3 jspl3_w_shift1_60(.douta(w_shift1_60[0]),.doutb(w_shift1_60[1]),.doutc(w_shift1_60[2]),.din(w_shift1_19[2]));
	jspl3 jspl3_w_shift1_61(.douta(w_shift1_61[0]),.doutb(w_shift1_61[1]),.doutc(w_shift1_61[2]),.din(w_shift1_20[0]));
	jspl3 jspl3_w_shift1_62(.douta(w_shift1_62[0]),.doutb(w_shift1_62[1]),.doutc(w_shift1_62[2]),.din(w_shift1_20[1]));
	jspl3 jspl3_w_shift1_63(.douta(w_dff_A_hDIMdffy1_0),.doutb(w_shift1_63[1]),.doutc(w_dff_A_bMqTrhbp3_2),.din(w_shift1_20[2]));
	jspl3 jspl3_w_shift2_0(.douta(w_shift2_0[0]),.doutb(w_shift2_0[1]),.doutc(w_dff_A_iZkaQ2vc3_2),.din(shift2));
	jspl3 jspl3_w_shift3_0(.douta(w_shift3_0[0]),.doutb(w_dff_A_6q7NhxpC3_1),.doutc(w_shift3_0[2]),.din(shift3));
	jspl3 jspl3_w_shift4_0(.douta(w_shift4_0[0]),.doutb(w_dff_A_kHgVQNIK1_1),.doutc(w_shift4_0[2]),.din(shift4));
	jspl3 jspl3_w_shift5_0(.douta(w_shift5_0[0]),.doutb(w_shift5_0[1]),.doutc(w_dff_A_6JmKMWA78_2),.din(shift5));
	jspl3 jspl3_w_shift6_0(.douta(w_shift6_0[0]),.doutb(w_dff_A_khYPEM4x6_1),.doutc(w_dff_A_eLfj31eX1_2),.din(shift6));
	jspl3 jspl3_w_shift6_1(.douta(w_dff_A_LF7uoH3p0_0),.doutb(w_dff_A_yhw6Bu9C1_1),.doutc(w_shift6_1[2]),.din(w_shift6_0[0]));
	jspl3 jspl3_w_shift6_2(.douta(w_shift6_2[0]),.doutb(w_shift6_2[1]),.doutc(w_shift6_2[2]),.din(w_shift6_0[1]));
	jspl3 jspl3_w_shift6_3(.douta(w_shift6_3[0]),.doutb(w_shift6_3[1]),.doutc(w_shift6_3[2]),.din(w_shift6_0[2]));
	jspl3 jspl3_w_shift6_4(.douta(w_shift6_4[0]),.doutb(w_shift6_4[1]),.doutc(w_shift6_4[2]),.din(w_shift6_1[0]));
	jspl3 jspl3_w_shift6_5(.douta(w_shift6_5[0]),.doutb(w_shift6_5[1]),.doutc(w_shift6_5[2]),.din(w_shift6_1[1]));
	jspl3 jspl3_w_shift6_6(.douta(w_dff_A_ilrk8ITG9_0),.doutb(w_shift6_6[1]),.doutc(w_dff_A_NGTUJztT7_2),.din(w_shift6_1[2]));
	jspl3 jspl3_w_shift6_7(.douta(w_shift6_7[0]),.doutb(w_shift6_7[1]),.doutc(w_shift6_7[2]),.din(w_shift6_2[0]));
	jspl3 jspl3_w_shift6_8(.douta(w_shift6_8[0]),.doutb(w_shift6_8[1]),.doutc(w_shift6_8[2]),.din(w_shift6_2[1]));
	jspl3 jspl3_w_shift6_9(.douta(w_shift6_9[0]),.doutb(w_shift6_9[1]),.doutc(w_shift6_9[2]),.din(w_shift6_2[2]));
	jspl3 jspl3_w_shift6_10(.douta(w_shift6_10[0]),.doutb(w_shift6_10[1]),.doutc(w_shift6_10[2]),.din(w_shift6_3[0]));
	jspl3 jspl3_w_shift6_11(.douta(w_shift6_11[0]),.doutb(w_shift6_11[1]),.doutc(w_shift6_11[2]),.din(w_shift6_3[1]));
	jspl3 jspl3_w_shift6_12(.douta(w_shift6_12[0]),.doutb(w_shift6_12[1]),.doutc(w_shift6_12[2]),.din(w_shift6_3[2]));
	jspl3 jspl3_w_shift6_13(.douta(w_shift6_13[0]),.doutb(w_shift6_13[1]),.doutc(w_shift6_13[2]),.din(w_shift6_4[0]));
	jspl3 jspl3_w_shift6_14(.douta(w_shift6_14[0]),.doutb(w_shift6_14[1]),.doutc(w_shift6_14[2]),.din(w_shift6_4[1]));
	jspl3 jspl3_w_shift6_15(.douta(w_shift6_15[0]),.doutb(w_shift6_15[1]),.doutc(w_shift6_15[2]),.din(w_shift6_4[2]));
	jspl3 jspl3_w_shift6_16(.douta(w_shift6_16[0]),.doutb(w_shift6_16[1]),.doutc(w_shift6_16[2]),.din(w_shift6_5[0]));
	jspl3 jspl3_w_shift6_17(.douta(w_shift6_17[0]),.doutb(w_shift6_17[1]),.doutc(w_shift6_17[2]),.din(w_shift6_5[1]));
	jspl3 jspl3_w_shift6_18(.douta(w_shift6_18[0]),.doutb(w_shift6_18[1]),.doutc(w_shift6_18[2]),.din(w_shift6_5[2]));
	jspl3 jspl3_w_shift6_19(.douta(w_shift6_19[0]),.doutb(w_shift6_19[1]),.doutc(w_shift6_19[2]),.din(w_shift6_6[0]));
	jspl3 jspl3_w_shift6_20(.douta(w_dff_A_SkPkN92h4_0),.doutb(w_dff_A_GnocIZ4d7_1),.doutc(w_shift6_20[2]),.din(w_shift6_6[1]));
	jspl3 jspl3_w_shift6_21(.douta(w_shift6_21[0]),.doutb(w_shift6_21[1]),.doutc(w_shift6_21[2]),.din(w_shift6_6[2]));
	jspl3 jspl3_w_shift6_22(.douta(w_shift6_22[0]),.doutb(w_shift6_22[1]),.doutc(w_shift6_22[2]),.din(w_shift6_7[0]));
	jspl3 jspl3_w_shift6_23(.douta(w_shift6_23[0]),.doutb(w_shift6_23[1]),.doutc(w_shift6_23[2]),.din(w_shift6_7[1]));
	jspl3 jspl3_w_shift6_24(.douta(w_shift6_24[0]),.doutb(w_shift6_24[1]),.doutc(w_shift6_24[2]),.din(w_shift6_7[2]));
	jspl3 jspl3_w_shift6_25(.douta(w_shift6_25[0]),.doutb(w_shift6_25[1]),.doutc(w_shift6_25[2]),.din(w_shift6_8[0]));
	jspl3 jspl3_w_shift6_26(.douta(w_shift6_26[0]),.doutb(w_shift6_26[1]),.doutc(w_shift6_26[2]),.din(w_shift6_8[1]));
	jspl3 jspl3_w_shift6_27(.douta(w_shift6_27[0]),.doutb(w_shift6_27[1]),.doutc(w_shift6_27[2]),.din(w_shift6_8[2]));
	jspl3 jspl3_w_shift6_28(.douta(w_shift6_28[0]),.doutb(w_shift6_28[1]),.doutc(w_shift6_28[2]),.din(w_shift6_9[0]));
	jspl3 jspl3_w_shift6_29(.douta(w_shift6_29[0]),.doutb(w_shift6_29[1]),.doutc(w_shift6_29[2]),.din(w_shift6_9[1]));
	jspl3 jspl3_w_shift6_30(.douta(w_shift6_30[0]),.doutb(w_shift6_30[1]),.doutc(w_shift6_30[2]),.din(w_shift6_9[2]));
	jspl3 jspl3_w_shift6_31(.douta(w_shift6_31[0]),.doutb(w_shift6_31[1]),.doutc(w_shift6_31[2]),.din(w_shift6_10[0]));
	jspl3 jspl3_w_shift6_32(.douta(w_shift6_32[0]),.doutb(w_shift6_32[1]),.doutc(w_shift6_32[2]),.din(w_shift6_10[1]));
	jspl3 jspl3_w_shift6_33(.douta(w_shift6_33[0]),.doutb(w_shift6_33[1]),.doutc(w_shift6_33[2]),.din(w_shift6_10[2]));
	jspl3 jspl3_w_shift6_34(.douta(w_shift6_34[0]),.doutb(w_shift6_34[1]),.doutc(w_shift6_34[2]),.din(w_shift6_11[0]));
	jspl3 jspl3_w_shift6_35(.douta(w_shift6_35[0]),.doutb(w_shift6_35[1]),.doutc(w_shift6_35[2]),.din(w_shift6_11[1]));
	jspl3 jspl3_w_shift6_36(.douta(w_shift6_36[0]),.doutb(w_shift6_36[1]),.doutc(w_shift6_36[2]),.din(w_shift6_11[2]));
	jspl3 jspl3_w_shift6_37(.douta(w_shift6_37[0]),.doutb(w_shift6_37[1]),.doutc(w_shift6_37[2]),.din(w_shift6_12[0]));
	jspl3 jspl3_w_shift6_38(.douta(w_shift6_38[0]),.doutb(w_shift6_38[1]),.doutc(w_shift6_38[2]),.din(w_shift6_12[1]));
	jspl3 jspl3_w_shift6_39(.douta(w_shift6_39[0]),.doutb(w_shift6_39[1]),.doutc(w_shift6_39[2]),.din(w_shift6_12[2]));
	jspl3 jspl3_w_shift6_40(.douta(w_shift6_40[0]),.doutb(w_shift6_40[1]),.doutc(w_shift6_40[2]),.din(w_shift6_13[0]));
	jspl3 jspl3_w_shift6_41(.douta(w_shift6_41[0]),.doutb(w_shift6_41[1]),.doutc(w_shift6_41[2]),.din(w_shift6_13[1]));
	jspl3 jspl3_w_shift6_42(.douta(w_shift6_42[0]),.doutb(w_shift6_42[1]),.doutc(w_shift6_42[2]),.din(w_shift6_13[2]));
	jspl3 jspl3_w_shift6_43(.douta(w_shift6_43[0]),.doutb(w_shift6_43[1]),.doutc(w_shift6_43[2]),.din(w_shift6_14[0]));
	jspl3 jspl3_w_shift6_44(.douta(w_shift6_44[0]),.doutb(w_shift6_44[1]),.doutc(w_shift6_44[2]),.din(w_shift6_14[1]));
	jspl3 jspl3_w_shift6_45(.douta(w_shift6_45[0]),.doutb(w_shift6_45[1]),.doutc(w_shift6_45[2]),.din(w_shift6_14[2]));
	jspl3 jspl3_w_shift6_46(.douta(w_shift6_46[0]),.doutb(w_shift6_46[1]),.doutc(w_shift6_46[2]),.din(w_shift6_15[0]));
	jspl3 jspl3_w_shift6_47(.douta(w_shift6_47[0]),.doutb(w_shift6_47[1]),.doutc(w_shift6_47[2]),.din(w_shift6_15[1]));
	jspl3 jspl3_w_shift6_48(.douta(w_shift6_48[0]),.doutb(w_shift6_48[1]),.doutc(w_shift6_48[2]),.din(w_shift6_15[2]));
	jspl3 jspl3_w_shift6_49(.douta(w_shift6_49[0]),.doutb(w_shift6_49[1]),.doutc(w_shift6_49[2]),.din(w_shift6_16[0]));
	jspl3 jspl3_w_shift6_50(.douta(w_shift6_50[0]),.doutb(w_shift6_50[1]),.doutc(w_shift6_50[2]),.din(w_shift6_16[1]));
	jspl3 jspl3_w_shift6_51(.douta(w_shift6_51[0]),.doutb(w_shift6_51[1]),.doutc(w_shift6_51[2]),.din(w_shift6_16[2]));
	jspl3 jspl3_w_shift6_52(.douta(w_shift6_52[0]),.doutb(w_shift6_52[1]),.doutc(w_shift6_52[2]),.din(w_shift6_17[0]));
	jspl3 jspl3_w_shift6_53(.douta(w_shift6_53[0]),.doutb(w_shift6_53[1]),.doutc(w_shift6_53[2]),.din(w_shift6_17[1]));
	jspl3 jspl3_w_shift6_54(.douta(w_shift6_54[0]),.doutb(w_shift6_54[1]),.doutc(w_shift6_54[2]),.din(w_shift6_17[2]));
	jspl3 jspl3_w_shift6_55(.douta(w_shift6_55[0]),.doutb(w_shift6_55[1]),.doutc(w_shift6_55[2]),.din(w_shift6_18[0]));
	jspl3 jspl3_w_shift6_56(.douta(w_shift6_56[0]),.doutb(w_shift6_56[1]),.doutc(w_shift6_56[2]),.din(w_shift6_18[1]));
	jspl3 jspl3_w_shift6_57(.douta(w_shift6_57[0]),.doutb(w_shift6_57[1]),.doutc(w_shift6_57[2]),.din(w_shift6_18[2]));
	jspl3 jspl3_w_shift6_58(.douta(w_shift6_58[0]),.doutb(w_shift6_58[1]),.doutc(w_shift6_58[2]),.din(w_shift6_19[0]));
	jspl3 jspl3_w_shift6_59(.douta(w_shift6_59[0]),.doutb(w_shift6_59[1]),.doutc(w_shift6_59[2]),.din(w_shift6_19[1]));
	jspl3 jspl3_w_shift6_60(.douta(w_shift6_60[0]),.doutb(w_shift6_60[1]),.doutc(w_shift6_60[2]),.din(w_shift6_19[2]));
	jspl3 jspl3_w_shift6_61(.douta(w_shift6_61[0]),.doutb(w_shift6_61[1]),.doutc(w_shift6_61[2]),.din(w_shift6_20[0]));
	jspl3 jspl3_w_shift6_62(.douta(w_shift6_62[0]),.doutb(w_shift6_62[1]),.doutc(w_shift6_62[2]),.din(w_shift6_20[1]));
	jspl3 jspl3_w_shift6_63(.douta(w_dff_A_bqhDMCvs6_0),.doutb(w_dff_A_QEbkLJAp3_1),.doutc(w_shift6_63[2]),.din(w_shift6_20[2]));
	jspl3 jspl3_w_n263_0(.douta(w_n263_0[0]),.doutb(w_n263_0[1]),.doutc(w_n263_0[2]),.din(w_dff_B_auwam0s87_3));
	jspl3 jspl3_w_n263_1(.douta(w_n263_1[0]),.doutb(w_n263_1[1]),.doutc(w_n263_1[2]),.din(w_n263_0[0]));
	jspl3 jspl3_w_n263_2(.douta(w_n263_2[0]),.doutb(w_n263_2[1]),.doutc(w_n263_2[2]),.din(w_n263_0[1]));
	jspl3 jspl3_w_n263_3(.douta(w_n263_3[0]),.doutb(w_n263_3[1]),.doutc(w_n263_3[2]),.din(w_n263_0[2]));
	jspl3 jspl3_w_n263_4(.douta(w_n263_4[0]),.doutb(w_n263_4[1]),.doutc(w_n263_4[2]),.din(w_n263_1[0]));
	jspl3 jspl3_w_n263_5(.douta(w_n263_5[0]),.doutb(w_n263_5[1]),.doutc(w_n263_5[2]),.din(w_n263_1[1]));
	jspl3 jspl3_w_n263_6(.douta(w_n263_6[0]),.doutb(w_n263_6[1]),.doutc(w_n263_6[2]),.din(w_n263_1[2]));
	jspl3 jspl3_w_n263_7(.douta(w_n263_7[0]),.doutb(w_n263_7[1]),.doutc(w_n263_7[2]),.din(w_n263_2[0]));
	jspl3 jspl3_w_n263_8(.douta(w_n263_8[0]),.doutb(w_n263_8[1]),.doutc(w_n263_8[2]),.din(w_n263_2[1]));
	jspl3 jspl3_w_n263_9(.douta(w_n263_9[0]),.doutb(w_n263_9[1]),.doutc(w_n263_9[2]),.din(w_n263_2[2]));
	jspl3 jspl3_w_n263_10(.douta(w_n263_10[0]),.doutb(w_n263_10[1]),.doutc(w_n263_10[2]),.din(w_n263_3[0]));
	jspl3 jspl3_w_n263_11(.douta(w_n263_11[0]),.doutb(w_n263_11[1]),.doutc(w_n263_11[2]),.din(w_n263_3[1]));
	jspl3 jspl3_w_n263_12(.douta(w_n263_12[0]),.doutb(w_n263_12[1]),.doutc(w_n263_12[2]),.din(w_n263_3[2]));
	jspl3 jspl3_w_n263_13(.douta(w_n263_13[0]),.doutb(w_n263_13[1]),.doutc(w_n263_13[2]),.din(w_n263_4[0]));
	jspl3 jspl3_w_n263_14(.douta(w_n263_14[0]),.doutb(w_n263_14[1]),.doutc(w_n263_14[2]),.din(w_n263_4[1]));
	jspl3 jspl3_w_n263_15(.douta(w_n263_15[0]),.doutb(w_n263_15[1]),.doutc(w_n263_15[2]),.din(w_n263_4[2]));
	jspl3 jspl3_w_n263_16(.douta(w_n263_16[0]),.doutb(w_n263_16[1]),.doutc(w_n263_16[2]),.din(w_n263_5[0]));
	jspl3 jspl3_w_n263_17(.douta(w_n263_17[0]),.doutb(w_n263_17[1]),.doutc(w_n263_17[2]),.din(w_n263_5[1]));
	jspl3 jspl3_w_n263_18(.douta(w_n263_18[0]),.doutb(w_n263_18[1]),.doutc(w_n263_18[2]),.din(w_n263_5[2]));
	jspl3 jspl3_w_n263_19(.douta(w_n263_19[0]),.doutb(w_n263_19[1]),.doutc(w_n263_19[2]),.din(w_n263_6[0]));
	jspl3 jspl3_w_n263_20(.douta(w_n263_20[0]),.doutb(w_n263_20[1]),.doutc(w_n263_20[2]),.din(w_n263_6[1]));
	jspl3 jspl3_w_n263_21(.douta(w_n263_21[0]),.doutb(w_n263_21[1]),.doutc(w_n263_21[2]),.din(w_n263_6[2]));
	jspl3 jspl3_w_n263_22(.douta(w_n263_22[0]),.doutb(w_n263_22[1]),.doutc(w_n263_22[2]),.din(w_n263_7[0]));
	jspl3 jspl3_w_n263_23(.douta(w_n263_23[0]),.doutb(w_n263_23[1]),.doutc(w_n263_23[2]),.din(w_n263_7[1]));
	jspl3 jspl3_w_n263_24(.douta(w_n263_24[0]),.doutb(w_n263_24[1]),.doutc(w_n263_24[2]),.din(w_n263_7[2]));
	jspl3 jspl3_w_n263_25(.douta(w_n263_25[0]),.doutb(w_n263_25[1]),.doutc(w_n263_25[2]),.din(w_n263_8[0]));
	jspl3 jspl3_w_n263_26(.douta(w_n263_26[0]),.doutb(w_n263_26[1]),.doutc(w_n263_26[2]),.din(w_n263_8[1]));
	jspl3 jspl3_w_n263_27(.douta(w_n263_27[0]),.doutb(w_n263_27[1]),.doutc(w_n263_27[2]),.din(w_n263_8[2]));
	jspl3 jspl3_w_n263_28(.douta(w_n263_28[0]),.doutb(w_n263_28[1]),.doutc(w_n263_28[2]),.din(w_n263_9[0]));
	jspl3 jspl3_w_n263_29(.douta(w_n263_29[0]),.doutb(w_n263_29[1]),.doutc(w_n263_29[2]),.din(w_n263_9[1]));
	jspl3 jspl3_w_n263_30(.douta(w_n263_30[0]),.doutb(w_n263_30[1]),.doutc(w_n263_30[2]),.din(w_n263_9[2]));
	jspl3 jspl3_w_n263_31(.douta(w_n263_31[0]),.doutb(w_n263_31[1]),.doutc(w_n263_31[2]),.din(w_n263_10[0]));
	jspl3 jspl3_w_n263_32(.douta(w_n263_32[0]),.doutb(w_n263_32[1]),.doutc(w_n263_32[2]),.din(w_n263_10[1]));
	jspl3 jspl3_w_n263_33(.douta(w_n263_33[0]),.doutb(w_n263_33[1]),.doutc(w_n263_33[2]),.din(w_n263_10[2]));
	jspl3 jspl3_w_n263_34(.douta(w_n263_34[0]),.doutb(w_n263_34[1]),.doutc(w_n263_34[2]),.din(w_n263_11[0]));
	jspl3 jspl3_w_n263_35(.douta(w_n263_35[0]),.doutb(w_n263_35[1]),.doutc(w_n263_35[2]),.din(w_n263_11[1]));
	jspl3 jspl3_w_n263_36(.douta(w_n263_36[0]),.doutb(w_n263_36[1]),.doutc(w_n263_36[2]),.din(w_n263_11[2]));
	jspl3 jspl3_w_n263_37(.douta(w_n263_37[0]),.doutb(w_n263_37[1]),.doutc(w_n263_37[2]),.din(w_n263_12[0]));
	jspl3 jspl3_w_n263_38(.douta(w_n263_38[0]),.doutb(w_n263_38[1]),.doutc(w_n263_38[2]),.din(w_n263_12[1]));
	jspl3 jspl3_w_n263_39(.douta(w_n263_39[0]),.doutb(w_n263_39[1]),.doutc(w_n263_39[2]),.din(w_n263_12[2]));
	jspl3 jspl3_w_n263_40(.douta(w_n263_40[0]),.doutb(w_n263_40[1]),.doutc(w_n263_40[2]),.din(w_n263_13[0]));
	jspl3 jspl3_w_n263_41(.douta(w_n263_41[0]),.doutb(w_n263_41[1]),.doutc(w_n263_41[2]),.din(w_n263_13[1]));
	jspl3 jspl3_w_n263_42(.douta(w_n263_42[0]),.doutb(w_n263_42[1]),.doutc(w_n263_42[2]),.din(w_n263_13[2]));
	jspl3 jspl3_w_n263_43(.douta(w_n263_43[0]),.doutb(w_n263_43[1]),.doutc(w_n263_43[2]),.din(w_n263_14[0]));
	jspl3 jspl3_w_n263_44(.douta(w_n263_44[0]),.doutb(w_n263_44[1]),.doutc(w_n263_44[2]),.din(w_n263_14[1]));
	jspl3 jspl3_w_n263_45(.douta(w_n263_45[0]),.doutb(w_n263_45[1]),.doutc(w_n263_45[2]),.din(w_n263_14[2]));
	jspl3 jspl3_w_n263_46(.douta(w_n263_46[0]),.doutb(w_n263_46[1]),.doutc(w_n263_46[2]),.din(w_n263_15[0]));
	jspl3 jspl3_w_n263_47(.douta(w_n263_47[0]),.doutb(w_n263_47[1]),.doutc(w_n263_47[2]),.din(w_n263_15[1]));
	jspl3 jspl3_w_n263_48(.douta(w_n263_48[0]),.doutb(w_n263_48[1]),.doutc(w_n263_48[2]),.din(w_n263_15[2]));
	jspl3 jspl3_w_n263_49(.douta(w_n263_49[0]),.doutb(w_n263_49[1]),.doutc(w_n263_49[2]),.din(w_n263_16[0]));
	jspl3 jspl3_w_n263_50(.douta(w_n263_50[0]),.doutb(w_n263_50[1]),.doutc(w_n263_50[2]),.din(w_n263_16[1]));
	jspl3 jspl3_w_n263_51(.douta(w_n263_51[0]),.doutb(w_n263_51[1]),.doutc(w_n263_51[2]),.din(w_n263_16[2]));
	jspl3 jspl3_w_n263_52(.douta(w_n263_52[0]),.doutb(w_n263_52[1]),.doutc(w_n263_52[2]),.din(w_n263_17[0]));
	jspl3 jspl3_w_n263_53(.douta(w_n263_53[0]),.doutb(w_n263_53[1]),.doutc(w_n263_53[2]),.din(w_n263_17[1]));
	jspl3 jspl3_w_n263_54(.douta(w_n263_54[0]),.doutb(w_n263_54[1]),.doutc(w_n263_54[2]),.din(w_n263_17[2]));
	jspl3 jspl3_w_n263_55(.douta(w_n263_55[0]),.doutb(w_n263_55[1]),.doutc(w_n263_55[2]),.din(w_n263_18[0]));
	jspl3 jspl3_w_n263_56(.douta(w_n263_56[0]),.doutb(w_n263_56[1]),.doutc(w_n263_56[2]),.din(w_n263_18[1]));
	jspl3 jspl3_w_n263_57(.douta(w_n263_57[0]),.doutb(w_n263_57[1]),.doutc(w_n263_57[2]),.din(w_n263_18[2]));
	jspl3 jspl3_w_n263_58(.douta(w_n263_58[0]),.doutb(w_n263_58[1]),.doutc(w_n263_58[2]),.din(w_n263_19[0]));
	jspl3 jspl3_w_n263_59(.douta(w_n263_59[0]),.doutb(w_n263_59[1]),.doutc(w_n263_59[2]),.din(w_n263_19[1]));
	jspl3 jspl3_w_n263_60(.douta(w_n263_60[0]),.doutb(w_n263_60[1]),.doutc(w_n263_60[2]),.din(w_n263_19[2]));
	jspl3 jspl3_w_n263_61(.douta(w_n263_61[0]),.doutb(w_n263_61[1]),.doutc(w_n263_61[2]),.din(w_n263_20[0]));
	jspl3 jspl3_w_n263_62(.douta(w_n263_62[0]),.doutb(w_n263_62[1]),.doutc(w_n263_62[2]),.din(w_n263_20[1]));
	jspl jspl_w_n263_63(.douta(w_n263_63[0]),.doutb(w_n263_63[1]),.din(w_n263_20[2]));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl3 jspl3_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.doutc(w_n265_0[2]),.din(w_dff_B_eLdE6Tba8_3));
	jspl3 jspl3_w_n265_1(.douta(w_n265_1[0]),.doutb(w_n265_1[1]),.doutc(w_n265_1[2]),.din(w_n265_0[0]));
	jspl3 jspl3_w_n265_2(.douta(w_n265_2[0]),.doutb(w_n265_2[1]),.doutc(w_n265_2[2]),.din(w_n265_0[1]));
	jspl3 jspl3_w_n265_3(.douta(w_n265_3[0]),.doutb(w_n265_3[1]),.doutc(w_n265_3[2]),.din(w_n265_0[2]));
	jspl3 jspl3_w_n265_4(.douta(w_n265_4[0]),.doutb(w_n265_4[1]),.doutc(w_n265_4[2]),.din(w_n265_1[0]));
	jspl3 jspl3_w_n265_5(.douta(w_n265_5[0]),.doutb(w_n265_5[1]),.doutc(w_n265_5[2]),.din(w_n265_1[1]));
	jspl3 jspl3_w_n265_6(.douta(w_n265_6[0]),.doutb(w_n265_6[1]),.doutc(w_n265_6[2]),.din(w_n265_1[2]));
	jspl3 jspl3_w_n265_7(.douta(w_n265_7[0]),.doutb(w_n265_7[1]),.doutc(w_n265_7[2]),.din(w_n265_2[0]));
	jspl3 jspl3_w_n265_8(.douta(w_n265_8[0]),.doutb(w_n265_8[1]),.doutc(w_n265_8[2]),.din(w_n265_2[1]));
	jspl3 jspl3_w_n265_9(.douta(w_n265_9[0]),.doutb(w_n265_9[1]),.doutc(w_n265_9[2]),.din(w_n265_2[2]));
	jspl3 jspl3_w_n265_10(.douta(w_n265_10[0]),.doutb(w_n265_10[1]),.doutc(w_n265_10[2]),.din(w_n265_3[0]));
	jspl3 jspl3_w_n265_11(.douta(w_n265_11[0]),.doutb(w_n265_11[1]),.doutc(w_n265_11[2]),.din(w_n265_3[1]));
	jspl3 jspl3_w_n265_12(.douta(w_n265_12[0]),.doutb(w_n265_12[1]),.doutc(w_n265_12[2]),.din(w_n265_3[2]));
	jspl3 jspl3_w_n265_13(.douta(w_n265_13[0]),.doutb(w_n265_13[1]),.doutc(w_n265_13[2]),.din(w_n265_4[0]));
	jspl3 jspl3_w_n265_14(.douta(w_n265_14[0]),.doutb(w_n265_14[1]),.doutc(w_n265_14[2]),.din(w_n265_4[1]));
	jspl3 jspl3_w_n265_15(.douta(w_n265_15[0]),.doutb(w_n265_15[1]),.doutc(w_n265_15[2]),.din(w_n265_4[2]));
	jspl3 jspl3_w_n265_16(.douta(w_n265_16[0]),.doutb(w_n265_16[1]),.doutc(w_n265_16[2]),.din(w_n265_5[0]));
	jspl3 jspl3_w_n265_17(.douta(w_n265_17[0]),.doutb(w_n265_17[1]),.doutc(w_n265_17[2]),.din(w_n265_5[1]));
	jspl3 jspl3_w_n265_18(.douta(w_n265_18[0]),.doutb(w_n265_18[1]),.doutc(w_n265_18[2]),.din(w_n265_5[2]));
	jspl3 jspl3_w_n265_19(.douta(w_n265_19[0]),.doutb(w_n265_19[1]),.doutc(w_n265_19[2]),.din(w_n265_6[0]));
	jspl3 jspl3_w_n265_20(.douta(w_n265_20[0]),.doutb(w_n265_20[1]),.doutc(w_n265_20[2]),.din(w_n265_6[1]));
	jspl3 jspl3_w_n265_21(.douta(w_n265_21[0]),.doutb(w_n265_21[1]),.doutc(w_n265_21[2]),.din(w_n265_6[2]));
	jspl3 jspl3_w_n265_22(.douta(w_n265_22[0]),.doutb(w_n265_22[1]),.doutc(w_n265_22[2]),.din(w_n265_7[0]));
	jspl3 jspl3_w_n265_23(.douta(w_n265_23[0]),.doutb(w_n265_23[1]),.doutc(w_n265_23[2]),.din(w_n265_7[1]));
	jspl3 jspl3_w_n265_24(.douta(w_n265_24[0]),.doutb(w_n265_24[1]),.doutc(w_n265_24[2]),.din(w_n265_7[2]));
	jspl3 jspl3_w_n265_25(.douta(w_n265_25[0]),.doutb(w_n265_25[1]),.doutc(w_n265_25[2]),.din(w_n265_8[0]));
	jspl3 jspl3_w_n265_26(.douta(w_n265_26[0]),.doutb(w_n265_26[1]),.doutc(w_n265_26[2]),.din(w_n265_8[1]));
	jspl3 jspl3_w_n265_27(.douta(w_n265_27[0]),.doutb(w_n265_27[1]),.doutc(w_n265_27[2]),.din(w_n265_8[2]));
	jspl3 jspl3_w_n265_28(.douta(w_n265_28[0]),.doutb(w_n265_28[1]),.doutc(w_n265_28[2]),.din(w_n265_9[0]));
	jspl3 jspl3_w_n265_29(.douta(w_n265_29[0]),.doutb(w_n265_29[1]),.doutc(w_n265_29[2]),.din(w_n265_9[1]));
	jspl3 jspl3_w_n265_30(.douta(w_n265_30[0]),.doutb(w_n265_30[1]),.doutc(w_n265_30[2]),.din(w_n265_9[2]));
	jspl3 jspl3_w_n265_31(.douta(w_n265_31[0]),.doutb(w_n265_31[1]),.doutc(w_n265_31[2]),.din(w_n265_10[0]));
	jspl3 jspl3_w_n265_32(.douta(w_n265_32[0]),.doutb(w_n265_32[1]),.doutc(w_n265_32[2]),.din(w_n265_10[1]));
	jspl3 jspl3_w_n265_33(.douta(w_n265_33[0]),.doutb(w_n265_33[1]),.doutc(w_n265_33[2]),.din(w_n265_10[2]));
	jspl3 jspl3_w_n265_34(.douta(w_n265_34[0]),.doutb(w_n265_34[1]),.doutc(w_n265_34[2]),.din(w_n265_11[0]));
	jspl3 jspl3_w_n265_35(.douta(w_n265_35[0]),.doutb(w_n265_35[1]),.doutc(w_n265_35[2]),.din(w_n265_11[1]));
	jspl3 jspl3_w_n265_36(.douta(w_n265_36[0]),.doutb(w_n265_36[1]),.doutc(w_n265_36[2]),.din(w_n265_11[2]));
	jspl3 jspl3_w_n265_37(.douta(w_n265_37[0]),.doutb(w_n265_37[1]),.doutc(w_n265_37[2]),.din(w_n265_12[0]));
	jspl3 jspl3_w_n265_38(.douta(w_n265_38[0]),.doutb(w_n265_38[1]),.doutc(w_n265_38[2]),.din(w_n265_12[1]));
	jspl3 jspl3_w_n265_39(.douta(w_n265_39[0]),.doutb(w_n265_39[1]),.doutc(w_n265_39[2]),.din(w_n265_12[2]));
	jspl3 jspl3_w_n265_40(.douta(w_n265_40[0]),.doutb(w_n265_40[1]),.doutc(w_n265_40[2]),.din(w_n265_13[0]));
	jspl3 jspl3_w_n265_41(.douta(w_n265_41[0]),.doutb(w_n265_41[1]),.doutc(w_n265_41[2]),.din(w_n265_13[1]));
	jspl3 jspl3_w_n265_42(.douta(w_n265_42[0]),.doutb(w_n265_42[1]),.doutc(w_n265_42[2]),.din(w_n265_13[2]));
	jspl3 jspl3_w_n265_43(.douta(w_n265_43[0]),.doutb(w_n265_43[1]),.doutc(w_n265_43[2]),.din(w_n265_14[0]));
	jspl3 jspl3_w_n265_44(.douta(w_n265_44[0]),.doutb(w_n265_44[1]),.doutc(w_n265_44[2]),.din(w_n265_14[1]));
	jspl3 jspl3_w_n265_45(.douta(w_n265_45[0]),.doutb(w_n265_45[1]),.doutc(w_n265_45[2]),.din(w_n265_14[2]));
	jspl3 jspl3_w_n265_46(.douta(w_n265_46[0]),.doutb(w_n265_46[1]),.doutc(w_n265_46[2]),.din(w_n265_15[0]));
	jspl3 jspl3_w_n265_47(.douta(w_n265_47[0]),.doutb(w_n265_47[1]),.doutc(w_n265_47[2]),.din(w_n265_15[1]));
	jspl3 jspl3_w_n265_48(.douta(w_n265_48[0]),.doutb(w_n265_48[1]),.doutc(w_n265_48[2]),.din(w_n265_15[2]));
	jspl3 jspl3_w_n265_49(.douta(w_n265_49[0]),.doutb(w_n265_49[1]),.doutc(w_n265_49[2]),.din(w_n265_16[0]));
	jspl3 jspl3_w_n265_50(.douta(w_n265_50[0]),.doutb(w_n265_50[1]),.doutc(w_n265_50[2]),.din(w_n265_16[1]));
	jspl3 jspl3_w_n265_51(.douta(w_n265_51[0]),.doutb(w_n265_51[1]),.doutc(w_n265_51[2]),.din(w_n265_16[2]));
	jspl3 jspl3_w_n265_52(.douta(w_n265_52[0]),.doutb(w_n265_52[1]),.doutc(w_n265_52[2]),.din(w_n265_17[0]));
	jspl3 jspl3_w_n265_53(.douta(w_n265_53[0]),.doutb(w_n265_53[1]),.doutc(w_n265_53[2]),.din(w_n265_17[1]));
	jspl3 jspl3_w_n265_54(.douta(w_n265_54[0]),.doutb(w_n265_54[1]),.doutc(w_n265_54[2]),.din(w_n265_17[2]));
	jspl3 jspl3_w_n265_55(.douta(w_n265_55[0]),.doutb(w_n265_55[1]),.doutc(w_n265_55[2]),.din(w_n265_18[0]));
	jspl3 jspl3_w_n265_56(.douta(w_n265_56[0]),.doutb(w_n265_56[1]),.doutc(w_n265_56[2]),.din(w_n265_18[1]));
	jspl3 jspl3_w_n265_57(.douta(w_n265_57[0]),.doutb(w_n265_57[1]),.doutc(w_n265_57[2]),.din(w_n265_18[2]));
	jspl3 jspl3_w_n265_58(.douta(w_n265_58[0]),.doutb(w_n265_58[1]),.doutc(w_n265_58[2]),.din(w_n265_19[0]));
	jspl3 jspl3_w_n265_59(.douta(w_n265_59[0]),.doutb(w_n265_59[1]),.doutc(w_n265_59[2]),.din(w_n265_19[1]));
	jspl3 jspl3_w_n265_60(.douta(w_n265_60[0]),.doutb(w_n265_60[1]),.doutc(w_n265_60[2]),.din(w_n265_19[2]));
	jspl3 jspl3_w_n265_61(.douta(w_n265_61[0]),.doutb(w_n265_61[1]),.doutc(w_n265_61[2]),.din(w_n265_20[0]));
	jspl3 jspl3_w_n265_62(.douta(w_n265_62[0]),.doutb(w_n265_62[1]),.doutc(w_n265_62[2]),.din(w_n265_20[1]));
	jspl jspl_w_n265_63(.douta(w_n265_63[0]),.doutb(w_n265_63[1]),.din(w_n265_20[2]));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.doutc(w_n267_0[2]),.din(w_dff_B_BzJqvu7e0_3));
	jspl3 jspl3_w_n267_1(.douta(w_n267_1[0]),.doutb(w_n267_1[1]),.doutc(w_n267_1[2]),.din(w_n267_0[0]));
	jspl3 jspl3_w_n267_2(.douta(w_n267_2[0]),.doutb(w_n267_2[1]),.doutc(w_n267_2[2]),.din(w_n267_0[1]));
	jspl3 jspl3_w_n267_3(.douta(w_n267_3[0]),.doutb(w_n267_3[1]),.doutc(w_n267_3[2]),.din(w_n267_0[2]));
	jspl3 jspl3_w_n267_4(.douta(w_n267_4[0]),.doutb(w_n267_4[1]),.doutc(w_n267_4[2]),.din(w_n267_1[0]));
	jspl3 jspl3_w_n267_5(.douta(w_n267_5[0]),.doutb(w_n267_5[1]),.doutc(w_n267_5[2]),.din(w_n267_1[1]));
	jspl3 jspl3_w_n267_6(.douta(w_n267_6[0]),.doutb(w_n267_6[1]),.doutc(w_n267_6[2]),.din(w_n267_1[2]));
	jspl3 jspl3_w_n267_7(.douta(w_n267_7[0]),.doutb(w_n267_7[1]),.doutc(w_n267_7[2]),.din(w_n267_2[0]));
	jspl3 jspl3_w_n267_8(.douta(w_n267_8[0]),.doutb(w_n267_8[1]),.doutc(w_n267_8[2]),.din(w_n267_2[1]));
	jspl3 jspl3_w_n267_9(.douta(w_n267_9[0]),.doutb(w_n267_9[1]),.doutc(w_n267_9[2]),.din(w_n267_2[2]));
	jspl3 jspl3_w_n267_10(.douta(w_n267_10[0]),.doutb(w_n267_10[1]),.doutc(w_n267_10[2]),.din(w_n267_3[0]));
	jspl3 jspl3_w_n267_11(.douta(w_n267_11[0]),.doutb(w_n267_11[1]),.doutc(w_n267_11[2]),.din(w_n267_3[1]));
	jspl3 jspl3_w_n267_12(.douta(w_n267_12[0]),.doutb(w_n267_12[1]),.doutc(w_n267_12[2]),.din(w_n267_3[2]));
	jspl3 jspl3_w_n267_13(.douta(w_n267_13[0]),.doutb(w_n267_13[1]),.doutc(w_n267_13[2]),.din(w_n267_4[0]));
	jspl3 jspl3_w_n267_14(.douta(w_n267_14[0]),.doutb(w_n267_14[1]),.doutc(w_n267_14[2]),.din(w_n267_4[1]));
	jspl3 jspl3_w_n267_15(.douta(w_n267_15[0]),.doutb(w_n267_15[1]),.doutc(w_n267_15[2]),.din(w_n267_4[2]));
	jspl3 jspl3_w_n267_16(.douta(w_n267_16[0]),.doutb(w_n267_16[1]),.doutc(w_n267_16[2]),.din(w_n267_5[0]));
	jspl3 jspl3_w_n267_17(.douta(w_n267_17[0]),.doutb(w_n267_17[1]),.doutc(w_n267_17[2]),.din(w_n267_5[1]));
	jspl3 jspl3_w_n267_18(.douta(w_n267_18[0]),.doutb(w_n267_18[1]),.doutc(w_n267_18[2]),.din(w_n267_5[2]));
	jspl3 jspl3_w_n267_19(.douta(w_n267_19[0]),.doutb(w_n267_19[1]),.doutc(w_n267_19[2]),.din(w_n267_6[0]));
	jspl3 jspl3_w_n267_20(.douta(w_n267_20[0]),.doutb(w_n267_20[1]),.doutc(w_n267_20[2]),.din(w_n267_6[1]));
	jspl3 jspl3_w_n267_21(.douta(w_n267_21[0]),.doutb(w_n267_21[1]),.doutc(w_n267_21[2]),.din(w_n267_6[2]));
	jspl3 jspl3_w_n267_22(.douta(w_n267_22[0]),.doutb(w_n267_22[1]),.doutc(w_n267_22[2]),.din(w_n267_7[0]));
	jspl3 jspl3_w_n267_23(.douta(w_n267_23[0]),.doutb(w_n267_23[1]),.doutc(w_n267_23[2]),.din(w_n267_7[1]));
	jspl3 jspl3_w_n267_24(.douta(w_n267_24[0]),.doutb(w_n267_24[1]),.doutc(w_n267_24[2]),.din(w_n267_7[2]));
	jspl3 jspl3_w_n267_25(.douta(w_n267_25[0]),.doutb(w_n267_25[1]),.doutc(w_n267_25[2]),.din(w_n267_8[0]));
	jspl3 jspl3_w_n267_26(.douta(w_n267_26[0]),.doutb(w_n267_26[1]),.doutc(w_n267_26[2]),.din(w_n267_8[1]));
	jspl3 jspl3_w_n267_27(.douta(w_n267_27[0]),.doutb(w_n267_27[1]),.doutc(w_n267_27[2]),.din(w_n267_8[2]));
	jspl3 jspl3_w_n267_28(.douta(w_n267_28[0]),.doutb(w_n267_28[1]),.doutc(w_n267_28[2]),.din(w_n267_9[0]));
	jspl3 jspl3_w_n267_29(.douta(w_n267_29[0]),.doutb(w_n267_29[1]),.doutc(w_n267_29[2]),.din(w_n267_9[1]));
	jspl3 jspl3_w_n267_30(.douta(w_n267_30[0]),.doutb(w_n267_30[1]),.doutc(w_n267_30[2]),.din(w_n267_9[2]));
	jspl3 jspl3_w_n267_31(.douta(w_n267_31[0]),.doutb(w_n267_31[1]),.doutc(w_n267_31[2]),.din(w_n267_10[0]));
	jspl3 jspl3_w_n267_32(.douta(w_n267_32[0]),.doutb(w_n267_32[1]),.doutc(w_n267_32[2]),.din(w_n267_10[1]));
	jspl3 jspl3_w_n267_33(.douta(w_n267_33[0]),.doutb(w_n267_33[1]),.doutc(w_n267_33[2]),.din(w_n267_10[2]));
	jspl3 jspl3_w_n267_34(.douta(w_n267_34[0]),.doutb(w_n267_34[1]),.doutc(w_n267_34[2]),.din(w_n267_11[0]));
	jspl3 jspl3_w_n267_35(.douta(w_n267_35[0]),.doutb(w_n267_35[1]),.doutc(w_n267_35[2]),.din(w_n267_11[1]));
	jspl3 jspl3_w_n267_36(.douta(w_n267_36[0]),.doutb(w_n267_36[1]),.doutc(w_n267_36[2]),.din(w_n267_11[2]));
	jspl3 jspl3_w_n267_37(.douta(w_n267_37[0]),.doutb(w_n267_37[1]),.doutc(w_n267_37[2]),.din(w_n267_12[0]));
	jspl3 jspl3_w_n267_38(.douta(w_n267_38[0]),.doutb(w_n267_38[1]),.doutc(w_n267_38[2]),.din(w_n267_12[1]));
	jspl3 jspl3_w_n267_39(.douta(w_n267_39[0]),.doutb(w_n267_39[1]),.doutc(w_n267_39[2]),.din(w_n267_12[2]));
	jspl3 jspl3_w_n267_40(.douta(w_n267_40[0]),.doutb(w_n267_40[1]),.doutc(w_n267_40[2]),.din(w_n267_13[0]));
	jspl3 jspl3_w_n267_41(.douta(w_n267_41[0]),.doutb(w_n267_41[1]),.doutc(w_n267_41[2]),.din(w_n267_13[1]));
	jspl3 jspl3_w_n267_42(.douta(w_n267_42[0]),.doutb(w_n267_42[1]),.doutc(w_n267_42[2]),.din(w_n267_13[2]));
	jspl3 jspl3_w_n267_43(.douta(w_n267_43[0]),.doutb(w_n267_43[1]),.doutc(w_n267_43[2]),.din(w_n267_14[0]));
	jspl3 jspl3_w_n267_44(.douta(w_n267_44[0]),.doutb(w_n267_44[1]),.doutc(w_n267_44[2]),.din(w_n267_14[1]));
	jspl3 jspl3_w_n267_45(.douta(w_n267_45[0]),.doutb(w_n267_45[1]),.doutc(w_n267_45[2]),.din(w_n267_14[2]));
	jspl3 jspl3_w_n267_46(.douta(w_n267_46[0]),.doutb(w_n267_46[1]),.doutc(w_n267_46[2]),.din(w_n267_15[0]));
	jspl3 jspl3_w_n267_47(.douta(w_n267_47[0]),.doutb(w_n267_47[1]),.doutc(w_n267_47[2]),.din(w_n267_15[1]));
	jspl3 jspl3_w_n267_48(.douta(w_n267_48[0]),.doutb(w_n267_48[1]),.doutc(w_n267_48[2]),.din(w_n267_15[2]));
	jspl3 jspl3_w_n267_49(.douta(w_n267_49[0]),.doutb(w_n267_49[1]),.doutc(w_n267_49[2]),.din(w_n267_16[0]));
	jspl3 jspl3_w_n267_50(.douta(w_n267_50[0]),.doutb(w_n267_50[1]),.doutc(w_n267_50[2]),.din(w_n267_16[1]));
	jspl3 jspl3_w_n267_51(.douta(w_n267_51[0]),.doutb(w_n267_51[1]),.doutc(w_n267_51[2]),.din(w_n267_16[2]));
	jspl3 jspl3_w_n267_52(.douta(w_n267_52[0]),.doutb(w_n267_52[1]),.doutc(w_n267_52[2]),.din(w_n267_17[0]));
	jspl3 jspl3_w_n267_53(.douta(w_n267_53[0]),.doutb(w_n267_53[1]),.doutc(w_n267_53[2]),.din(w_n267_17[1]));
	jspl3 jspl3_w_n267_54(.douta(w_n267_54[0]),.doutb(w_n267_54[1]),.doutc(w_n267_54[2]),.din(w_n267_17[2]));
	jspl3 jspl3_w_n267_55(.douta(w_n267_55[0]),.doutb(w_n267_55[1]),.doutc(w_n267_55[2]),.din(w_n267_18[0]));
	jspl3 jspl3_w_n267_56(.douta(w_n267_56[0]),.doutb(w_n267_56[1]),.doutc(w_n267_56[2]),.din(w_n267_18[1]));
	jspl3 jspl3_w_n267_57(.douta(w_n267_57[0]),.doutb(w_n267_57[1]),.doutc(w_n267_57[2]),.din(w_n267_18[2]));
	jspl3 jspl3_w_n267_58(.douta(w_n267_58[0]),.doutb(w_n267_58[1]),.doutc(w_n267_58[2]),.din(w_n267_19[0]));
	jspl3 jspl3_w_n267_59(.douta(w_n267_59[0]),.doutb(w_n267_59[1]),.doutc(w_n267_59[2]),.din(w_n267_19[1]));
	jspl3 jspl3_w_n267_60(.douta(w_n267_60[0]),.doutb(w_n267_60[1]),.doutc(w_n267_60[2]),.din(w_n267_19[2]));
	jspl3 jspl3_w_n267_61(.douta(w_n267_61[0]),.doutb(w_n267_61[1]),.doutc(w_n267_61[2]),.din(w_n267_20[0]));
	jspl3 jspl3_w_n267_62(.douta(w_n267_62[0]),.doutb(w_n267_62[1]),.doutc(w_n267_62[2]),.din(w_n267_20[1]));
	jspl jspl_w_n267_63(.douta(w_n267_63[0]),.doutb(w_n267_63[1]),.din(w_n267_20[2]));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.doutc(w_n269_1[2]),.din(w_n269_0[0]));
	jspl3 jspl3_w_n269_2(.douta(w_n269_2[0]),.doutb(w_n269_2[1]),.doutc(w_n269_2[2]),.din(w_n269_0[1]));
	jspl3 jspl3_w_n269_3(.douta(w_n269_3[0]),.doutb(w_n269_3[1]),.doutc(w_n269_3[2]),.din(w_n269_0[2]));
	jspl3 jspl3_w_n269_4(.douta(w_n269_4[0]),.doutb(w_n269_4[1]),.doutc(w_n269_4[2]),.din(w_n269_1[0]));
	jspl3 jspl3_w_n269_5(.douta(w_n269_5[0]),.doutb(w_n269_5[1]),.doutc(w_n269_5[2]),.din(w_n269_1[1]));
	jspl3 jspl3_w_n269_6(.douta(w_n269_6[0]),.doutb(w_n269_6[1]),.doutc(w_n269_6[2]),.din(w_n269_1[2]));
	jspl3 jspl3_w_n269_7(.douta(w_n269_7[0]),.doutb(w_n269_7[1]),.doutc(w_n269_7[2]),.din(w_n269_2[0]));
	jspl3 jspl3_w_n269_8(.douta(w_n269_8[0]),.doutb(w_n269_8[1]),.doutc(w_n269_8[2]),.din(w_n269_2[1]));
	jspl3 jspl3_w_n269_9(.douta(w_n269_9[0]),.doutb(w_n269_9[1]),.doutc(w_n269_9[2]),.din(w_n269_2[2]));
	jspl3 jspl3_w_n269_10(.douta(w_n269_10[0]),.doutb(w_n269_10[1]),.doutc(w_n269_10[2]),.din(w_n269_3[0]));
	jspl3 jspl3_w_n269_11(.douta(w_n269_11[0]),.doutb(w_n269_11[1]),.doutc(w_n269_11[2]),.din(w_n269_3[1]));
	jspl3 jspl3_w_n269_12(.douta(w_n269_12[0]),.doutb(w_n269_12[1]),.doutc(w_n269_12[2]),.din(w_n269_3[2]));
	jspl3 jspl3_w_n269_13(.douta(w_n269_13[0]),.doutb(w_n269_13[1]),.doutc(w_n269_13[2]),.din(w_n269_4[0]));
	jspl3 jspl3_w_n269_14(.douta(w_n269_14[0]),.doutb(w_n269_14[1]),.doutc(w_n269_14[2]),.din(w_n269_4[1]));
	jspl3 jspl3_w_n269_15(.douta(w_n269_15[0]),.doutb(w_n269_15[1]),.doutc(w_n269_15[2]),.din(w_n269_4[2]));
	jspl3 jspl3_w_n269_16(.douta(w_n269_16[0]),.doutb(w_n269_16[1]),.doutc(w_n269_16[2]),.din(w_n269_5[0]));
	jspl3 jspl3_w_n269_17(.douta(w_n269_17[0]),.doutb(w_n269_17[1]),.doutc(w_n269_17[2]),.din(w_n269_5[1]));
	jspl3 jspl3_w_n269_18(.douta(w_n269_18[0]),.doutb(w_n269_18[1]),.doutc(w_n269_18[2]),.din(w_n269_5[2]));
	jspl3 jspl3_w_n269_19(.douta(w_n269_19[0]),.doutb(w_n269_19[1]),.doutc(w_n269_19[2]),.din(w_n269_6[0]));
	jspl3 jspl3_w_n269_20(.douta(w_n269_20[0]),.doutb(w_n269_20[1]),.doutc(w_n269_20[2]),.din(w_n269_6[1]));
	jspl3 jspl3_w_n269_21(.douta(w_n269_21[0]),.doutb(w_n269_21[1]),.doutc(w_n269_21[2]),.din(w_n269_6[2]));
	jspl3 jspl3_w_n269_22(.douta(w_n269_22[0]),.doutb(w_n269_22[1]),.doutc(w_n269_22[2]),.din(w_n269_7[0]));
	jspl3 jspl3_w_n269_23(.douta(w_n269_23[0]),.doutb(w_n269_23[1]),.doutc(w_n269_23[2]),.din(w_n269_7[1]));
	jspl3 jspl3_w_n269_24(.douta(w_n269_24[0]),.doutb(w_n269_24[1]),.doutc(w_n269_24[2]),.din(w_n269_7[2]));
	jspl3 jspl3_w_n269_25(.douta(w_n269_25[0]),.doutb(w_n269_25[1]),.doutc(w_n269_25[2]),.din(w_n269_8[0]));
	jspl3 jspl3_w_n269_26(.douta(w_n269_26[0]),.doutb(w_n269_26[1]),.doutc(w_n269_26[2]),.din(w_n269_8[1]));
	jspl3 jspl3_w_n269_27(.douta(w_n269_27[0]),.doutb(w_n269_27[1]),.doutc(w_n269_27[2]),.din(w_n269_8[2]));
	jspl3 jspl3_w_n269_28(.douta(w_n269_28[0]),.doutb(w_n269_28[1]),.doutc(w_n269_28[2]),.din(w_n269_9[0]));
	jspl3 jspl3_w_n269_29(.douta(w_n269_29[0]),.doutb(w_n269_29[1]),.doutc(w_n269_29[2]),.din(w_n269_9[1]));
	jspl3 jspl3_w_n269_30(.douta(w_n269_30[0]),.doutb(w_n269_30[1]),.doutc(w_n269_30[2]),.din(w_n269_9[2]));
	jspl3 jspl3_w_n269_31(.douta(w_n269_31[0]),.doutb(w_n269_31[1]),.doutc(w_n269_31[2]),.din(w_n269_10[0]));
	jspl3 jspl3_w_n269_32(.douta(w_n269_32[0]),.doutb(w_n269_32[1]),.doutc(w_n269_32[2]),.din(w_n269_10[1]));
	jspl3 jspl3_w_n269_33(.douta(w_n269_33[0]),.doutb(w_n269_33[1]),.doutc(w_n269_33[2]),.din(w_n269_10[2]));
	jspl3 jspl3_w_n269_34(.douta(w_n269_34[0]),.doutb(w_n269_34[1]),.doutc(w_n269_34[2]),.din(w_n269_11[0]));
	jspl3 jspl3_w_n269_35(.douta(w_n269_35[0]),.doutb(w_n269_35[1]),.doutc(w_n269_35[2]),.din(w_n269_11[1]));
	jspl3 jspl3_w_n269_36(.douta(w_n269_36[0]),.doutb(w_n269_36[1]),.doutc(w_n269_36[2]),.din(w_n269_11[2]));
	jspl3 jspl3_w_n269_37(.douta(w_n269_37[0]),.doutb(w_n269_37[1]),.doutc(w_n269_37[2]),.din(w_n269_12[0]));
	jspl3 jspl3_w_n269_38(.douta(w_n269_38[0]),.doutb(w_n269_38[1]),.doutc(w_n269_38[2]),.din(w_n269_12[1]));
	jspl3 jspl3_w_n269_39(.douta(w_n269_39[0]),.doutb(w_n269_39[1]),.doutc(w_n269_39[2]),.din(w_n269_12[2]));
	jspl3 jspl3_w_n269_40(.douta(w_n269_40[0]),.doutb(w_n269_40[1]),.doutc(w_n269_40[2]),.din(w_n269_13[0]));
	jspl3 jspl3_w_n269_41(.douta(w_n269_41[0]),.doutb(w_n269_41[1]),.doutc(w_n269_41[2]),.din(w_n269_13[1]));
	jspl3 jspl3_w_n269_42(.douta(w_n269_42[0]),.doutb(w_n269_42[1]),.doutc(w_n269_42[2]),.din(w_n269_13[2]));
	jspl3 jspl3_w_n269_43(.douta(w_n269_43[0]),.doutb(w_n269_43[1]),.doutc(w_n269_43[2]),.din(w_n269_14[0]));
	jspl3 jspl3_w_n269_44(.douta(w_n269_44[0]),.doutb(w_n269_44[1]),.doutc(w_n269_44[2]),.din(w_n269_14[1]));
	jspl3 jspl3_w_n269_45(.douta(w_n269_45[0]),.doutb(w_n269_45[1]),.doutc(w_n269_45[2]),.din(w_n269_14[2]));
	jspl3 jspl3_w_n269_46(.douta(w_n269_46[0]),.doutb(w_n269_46[1]),.doutc(w_n269_46[2]),.din(w_n269_15[0]));
	jspl3 jspl3_w_n269_47(.douta(w_n269_47[0]),.doutb(w_n269_47[1]),.doutc(w_n269_47[2]),.din(w_n269_15[1]));
	jspl3 jspl3_w_n269_48(.douta(w_n269_48[0]),.doutb(w_n269_48[1]),.doutc(w_n269_48[2]),.din(w_n269_15[2]));
	jspl3 jspl3_w_n269_49(.douta(w_n269_49[0]),.doutb(w_n269_49[1]),.doutc(w_n269_49[2]),.din(w_n269_16[0]));
	jspl3 jspl3_w_n269_50(.douta(w_n269_50[0]),.doutb(w_n269_50[1]),.doutc(w_n269_50[2]),.din(w_n269_16[1]));
	jspl3 jspl3_w_n269_51(.douta(w_n269_51[0]),.doutb(w_n269_51[1]),.doutc(w_n269_51[2]),.din(w_n269_16[2]));
	jspl3 jspl3_w_n269_52(.douta(w_n269_52[0]),.doutb(w_n269_52[1]),.doutc(w_n269_52[2]),.din(w_n269_17[0]));
	jspl3 jspl3_w_n269_53(.douta(w_n269_53[0]),.doutb(w_n269_53[1]),.doutc(w_n269_53[2]),.din(w_n269_17[1]));
	jspl3 jspl3_w_n269_54(.douta(w_n269_54[0]),.doutb(w_n269_54[1]),.doutc(w_n269_54[2]),.din(w_n269_17[2]));
	jspl3 jspl3_w_n269_55(.douta(w_n269_55[0]),.doutb(w_n269_55[1]),.doutc(w_n269_55[2]),.din(w_n269_18[0]));
	jspl3 jspl3_w_n269_56(.douta(w_n269_56[0]),.doutb(w_n269_56[1]),.doutc(w_n269_56[2]),.din(w_n269_18[1]));
	jspl3 jspl3_w_n269_57(.douta(w_n269_57[0]),.doutb(w_n269_57[1]),.doutc(w_n269_57[2]),.din(w_n269_18[2]));
	jspl3 jspl3_w_n269_58(.douta(w_n269_58[0]),.doutb(w_n269_58[1]),.doutc(w_n269_58[2]),.din(w_n269_19[0]));
	jspl3 jspl3_w_n269_59(.douta(w_n269_59[0]),.doutb(w_n269_59[1]),.doutc(w_n269_59[2]),.din(w_n269_19[1]));
	jspl3 jspl3_w_n269_60(.douta(w_n269_60[0]),.doutb(w_n269_60[1]),.doutc(w_n269_60[2]),.din(w_n269_19[2]));
	jspl3 jspl3_w_n269_61(.douta(w_n269_61[0]),.doutb(w_n269_61[1]),.doutc(w_n269_61[2]),.din(w_n269_20[0]));
	jspl3 jspl3_w_n269_62(.douta(w_n269_62[0]),.doutb(w_n269_62[1]),.doutc(w_n269_62[2]),.din(w_n269_20[1]));
	jspl jspl_w_n269_63(.douta(w_n269_63[0]),.doutb(w_n269_63[1]),.din(w_n269_20[2]));
	jspl jspl_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.din(n271));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.doutc(w_n273_0[2]),.din(w_dff_B_AMEaIxgs6_3));
	jspl3 jspl3_w_n273_1(.douta(w_n273_1[0]),.doutb(w_n273_1[1]),.doutc(w_n273_1[2]),.din(w_n273_0[0]));
	jspl3 jspl3_w_n273_2(.douta(w_n273_2[0]),.doutb(w_n273_2[1]),.doutc(w_n273_2[2]),.din(w_n273_0[1]));
	jspl3 jspl3_w_n273_3(.douta(w_n273_3[0]),.doutb(w_n273_3[1]),.doutc(w_n273_3[2]),.din(w_n273_0[2]));
	jspl3 jspl3_w_n273_4(.douta(w_n273_4[0]),.doutb(w_n273_4[1]),.doutc(w_n273_4[2]),.din(w_n273_1[0]));
	jspl3 jspl3_w_n273_5(.douta(w_n273_5[0]),.doutb(w_n273_5[1]),.doutc(w_n273_5[2]),.din(w_n273_1[1]));
	jspl3 jspl3_w_n273_6(.douta(w_n273_6[0]),.doutb(w_n273_6[1]),.doutc(w_n273_6[2]),.din(w_n273_1[2]));
	jspl3 jspl3_w_n273_7(.douta(w_n273_7[0]),.doutb(w_n273_7[1]),.doutc(w_n273_7[2]),.din(w_n273_2[0]));
	jspl3 jspl3_w_n273_8(.douta(w_n273_8[0]),.doutb(w_n273_8[1]),.doutc(w_n273_8[2]),.din(w_n273_2[1]));
	jspl3 jspl3_w_n273_9(.douta(w_n273_9[0]),.doutb(w_n273_9[1]),.doutc(w_n273_9[2]),.din(w_n273_2[2]));
	jspl3 jspl3_w_n273_10(.douta(w_n273_10[0]),.doutb(w_n273_10[1]),.doutc(w_n273_10[2]),.din(w_n273_3[0]));
	jspl3 jspl3_w_n273_11(.douta(w_n273_11[0]),.doutb(w_n273_11[1]),.doutc(w_n273_11[2]),.din(w_n273_3[1]));
	jspl3 jspl3_w_n273_12(.douta(w_n273_12[0]),.doutb(w_n273_12[1]),.doutc(w_n273_12[2]),.din(w_n273_3[2]));
	jspl3 jspl3_w_n273_13(.douta(w_n273_13[0]),.doutb(w_n273_13[1]),.doutc(w_n273_13[2]),.din(w_n273_4[0]));
	jspl3 jspl3_w_n273_14(.douta(w_n273_14[0]),.doutb(w_n273_14[1]),.doutc(w_n273_14[2]),.din(w_n273_4[1]));
	jspl3 jspl3_w_n273_15(.douta(w_n273_15[0]),.doutb(w_n273_15[1]),.doutc(w_n273_15[2]),.din(w_n273_4[2]));
	jspl3 jspl3_w_n273_16(.douta(w_n273_16[0]),.doutb(w_n273_16[1]),.doutc(w_n273_16[2]),.din(w_n273_5[0]));
	jspl3 jspl3_w_n273_17(.douta(w_n273_17[0]),.doutb(w_n273_17[1]),.doutc(w_n273_17[2]),.din(w_n273_5[1]));
	jspl3 jspl3_w_n273_18(.douta(w_n273_18[0]),.doutb(w_n273_18[1]),.doutc(w_n273_18[2]),.din(w_n273_5[2]));
	jspl3 jspl3_w_n273_19(.douta(w_n273_19[0]),.doutb(w_n273_19[1]),.doutc(w_n273_19[2]),.din(w_n273_6[0]));
	jspl3 jspl3_w_n273_20(.douta(w_n273_20[0]),.doutb(w_n273_20[1]),.doutc(w_n273_20[2]),.din(w_n273_6[1]));
	jspl3 jspl3_w_n273_21(.douta(w_n273_21[0]),.doutb(w_n273_21[1]),.doutc(w_n273_21[2]),.din(w_n273_6[2]));
	jspl3 jspl3_w_n273_22(.douta(w_n273_22[0]),.doutb(w_n273_22[1]),.doutc(w_n273_22[2]),.din(w_n273_7[0]));
	jspl3 jspl3_w_n273_23(.douta(w_n273_23[0]),.doutb(w_n273_23[1]),.doutc(w_n273_23[2]),.din(w_n273_7[1]));
	jspl3 jspl3_w_n273_24(.douta(w_n273_24[0]),.doutb(w_n273_24[1]),.doutc(w_n273_24[2]),.din(w_n273_7[2]));
	jspl3 jspl3_w_n273_25(.douta(w_n273_25[0]),.doutb(w_n273_25[1]),.doutc(w_n273_25[2]),.din(w_n273_8[0]));
	jspl3 jspl3_w_n273_26(.douta(w_n273_26[0]),.doutb(w_n273_26[1]),.doutc(w_n273_26[2]),.din(w_n273_8[1]));
	jspl3 jspl3_w_n273_27(.douta(w_n273_27[0]),.doutb(w_n273_27[1]),.doutc(w_n273_27[2]),.din(w_n273_8[2]));
	jspl3 jspl3_w_n273_28(.douta(w_n273_28[0]),.doutb(w_n273_28[1]),.doutc(w_n273_28[2]),.din(w_n273_9[0]));
	jspl3 jspl3_w_n273_29(.douta(w_n273_29[0]),.doutb(w_n273_29[1]),.doutc(w_n273_29[2]),.din(w_n273_9[1]));
	jspl3 jspl3_w_n273_30(.douta(w_n273_30[0]),.doutb(w_n273_30[1]),.doutc(w_n273_30[2]),.din(w_n273_9[2]));
	jspl3 jspl3_w_n273_31(.douta(w_n273_31[0]),.doutb(w_n273_31[1]),.doutc(w_n273_31[2]),.din(w_n273_10[0]));
	jspl3 jspl3_w_n273_32(.douta(w_n273_32[0]),.doutb(w_n273_32[1]),.doutc(w_n273_32[2]),.din(w_n273_10[1]));
	jspl3 jspl3_w_n273_33(.douta(w_n273_33[0]),.doutb(w_n273_33[1]),.doutc(w_n273_33[2]),.din(w_n273_10[2]));
	jspl3 jspl3_w_n273_34(.douta(w_n273_34[0]),.doutb(w_n273_34[1]),.doutc(w_n273_34[2]),.din(w_n273_11[0]));
	jspl3 jspl3_w_n273_35(.douta(w_n273_35[0]),.doutb(w_n273_35[1]),.doutc(w_n273_35[2]),.din(w_n273_11[1]));
	jspl3 jspl3_w_n273_36(.douta(w_n273_36[0]),.doutb(w_n273_36[1]),.doutc(w_n273_36[2]),.din(w_n273_11[2]));
	jspl3 jspl3_w_n273_37(.douta(w_n273_37[0]),.doutb(w_n273_37[1]),.doutc(w_n273_37[2]),.din(w_n273_12[0]));
	jspl3 jspl3_w_n273_38(.douta(w_n273_38[0]),.doutb(w_n273_38[1]),.doutc(w_n273_38[2]),.din(w_n273_12[1]));
	jspl3 jspl3_w_n273_39(.douta(w_n273_39[0]),.doutb(w_n273_39[1]),.doutc(w_n273_39[2]),.din(w_n273_12[2]));
	jspl3 jspl3_w_n273_40(.douta(w_n273_40[0]),.doutb(w_n273_40[1]),.doutc(w_n273_40[2]),.din(w_n273_13[0]));
	jspl3 jspl3_w_n273_41(.douta(w_n273_41[0]),.doutb(w_n273_41[1]),.doutc(w_n273_41[2]),.din(w_n273_13[1]));
	jspl3 jspl3_w_n273_42(.douta(w_n273_42[0]),.doutb(w_n273_42[1]),.doutc(w_n273_42[2]),.din(w_n273_13[2]));
	jspl3 jspl3_w_n273_43(.douta(w_n273_43[0]),.doutb(w_n273_43[1]),.doutc(w_n273_43[2]),.din(w_n273_14[0]));
	jspl3 jspl3_w_n273_44(.douta(w_n273_44[0]),.doutb(w_n273_44[1]),.doutc(w_n273_44[2]),.din(w_n273_14[1]));
	jspl3 jspl3_w_n273_45(.douta(w_n273_45[0]),.doutb(w_n273_45[1]),.doutc(w_n273_45[2]),.din(w_n273_14[2]));
	jspl3 jspl3_w_n273_46(.douta(w_n273_46[0]),.doutb(w_n273_46[1]),.doutc(w_n273_46[2]),.din(w_n273_15[0]));
	jspl3 jspl3_w_n273_47(.douta(w_n273_47[0]),.doutb(w_n273_47[1]),.doutc(w_n273_47[2]),.din(w_n273_15[1]));
	jspl3 jspl3_w_n273_48(.douta(w_n273_48[0]),.doutb(w_n273_48[1]),.doutc(w_n273_48[2]),.din(w_n273_15[2]));
	jspl3 jspl3_w_n273_49(.douta(w_n273_49[0]),.doutb(w_n273_49[1]),.doutc(w_n273_49[2]),.din(w_n273_16[0]));
	jspl3 jspl3_w_n273_50(.douta(w_n273_50[0]),.doutb(w_n273_50[1]),.doutc(w_n273_50[2]),.din(w_n273_16[1]));
	jspl3 jspl3_w_n273_51(.douta(w_n273_51[0]),.doutb(w_n273_51[1]),.doutc(w_n273_51[2]),.din(w_n273_16[2]));
	jspl3 jspl3_w_n273_52(.douta(w_n273_52[0]),.doutb(w_n273_52[1]),.doutc(w_n273_52[2]),.din(w_n273_17[0]));
	jspl3 jspl3_w_n273_53(.douta(w_n273_53[0]),.doutb(w_n273_53[1]),.doutc(w_n273_53[2]),.din(w_n273_17[1]));
	jspl3 jspl3_w_n273_54(.douta(w_n273_54[0]),.doutb(w_n273_54[1]),.doutc(w_n273_54[2]),.din(w_n273_17[2]));
	jspl3 jspl3_w_n273_55(.douta(w_n273_55[0]),.doutb(w_n273_55[1]),.doutc(w_n273_55[2]),.din(w_n273_18[0]));
	jspl3 jspl3_w_n273_56(.douta(w_n273_56[0]),.doutb(w_n273_56[1]),.doutc(w_n273_56[2]),.din(w_n273_18[1]));
	jspl3 jspl3_w_n273_57(.douta(w_n273_57[0]),.doutb(w_n273_57[1]),.doutc(w_n273_57[2]),.din(w_n273_18[2]));
	jspl3 jspl3_w_n273_58(.douta(w_n273_58[0]),.doutb(w_n273_58[1]),.doutc(w_n273_58[2]),.din(w_n273_19[0]));
	jspl3 jspl3_w_n273_59(.douta(w_n273_59[0]),.doutb(w_n273_59[1]),.doutc(w_n273_59[2]),.din(w_n273_19[1]));
	jspl3 jspl3_w_n273_60(.douta(w_n273_60[0]),.doutb(w_n273_60[1]),.doutc(w_n273_60[2]),.din(w_n273_19[2]));
	jspl3 jspl3_w_n273_61(.douta(w_n273_61[0]),.doutb(w_n273_61[1]),.doutc(w_n273_61[2]),.din(w_n273_20[0]));
	jspl3 jspl3_w_n273_62(.douta(w_n273_62[0]),.doutb(w_n273_62[1]),.doutc(w_n273_62[2]),.din(w_n273_20[1]));
	jspl jspl_w_n273_63(.douta(w_n273_63[0]),.doutb(w_n273_63[1]),.din(w_n273_20[2]));
	jspl jspl_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.din(n276));
	jspl3 jspl3_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.doutc(w_n278_0[2]),.din(n278));
	jspl jspl_w_n278_1(.douta(w_n278_1[0]),.doutb(w_n278_1[1]),.din(w_n278_0[0]));
	jspl jspl_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.din(n280));
	jspl3 jspl3_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.doutc(w_n281_0[2]),.din(w_dff_B_FULzpxU81_3));
	jspl3 jspl3_w_n281_1(.douta(w_n281_1[0]),.doutb(w_n281_1[1]),.doutc(w_n281_1[2]),.din(w_n281_0[0]));
	jspl3 jspl3_w_n281_2(.douta(w_n281_2[0]),.doutb(w_n281_2[1]),.doutc(w_n281_2[2]),.din(w_n281_0[1]));
	jspl3 jspl3_w_n281_3(.douta(w_n281_3[0]),.doutb(w_n281_3[1]),.doutc(w_n281_3[2]),.din(w_n281_0[2]));
	jspl3 jspl3_w_n281_4(.douta(w_n281_4[0]),.doutb(w_n281_4[1]),.doutc(w_n281_4[2]),.din(w_n281_1[0]));
	jspl3 jspl3_w_n281_5(.douta(w_n281_5[0]),.doutb(w_n281_5[1]),.doutc(w_n281_5[2]),.din(w_n281_1[1]));
	jspl3 jspl3_w_n281_6(.douta(w_n281_6[0]),.doutb(w_n281_6[1]),.doutc(w_n281_6[2]),.din(w_n281_1[2]));
	jspl3 jspl3_w_n281_7(.douta(w_n281_7[0]),.doutb(w_n281_7[1]),.doutc(w_n281_7[2]),.din(w_n281_2[0]));
	jspl3 jspl3_w_n281_8(.douta(w_n281_8[0]),.doutb(w_n281_8[1]),.doutc(w_n281_8[2]),.din(w_n281_2[1]));
	jspl3 jspl3_w_n281_9(.douta(w_n281_9[0]),.doutb(w_n281_9[1]),.doutc(w_n281_9[2]),.din(w_n281_2[2]));
	jspl3 jspl3_w_n281_10(.douta(w_n281_10[0]),.doutb(w_n281_10[1]),.doutc(w_n281_10[2]),.din(w_n281_3[0]));
	jspl3 jspl3_w_n281_11(.douta(w_n281_11[0]),.doutb(w_n281_11[1]),.doutc(w_n281_11[2]),.din(w_n281_3[1]));
	jspl3 jspl3_w_n281_12(.douta(w_n281_12[0]),.doutb(w_n281_12[1]),.doutc(w_n281_12[2]),.din(w_n281_3[2]));
	jspl3 jspl3_w_n281_13(.douta(w_n281_13[0]),.doutb(w_n281_13[1]),.doutc(w_n281_13[2]),.din(w_n281_4[0]));
	jspl3 jspl3_w_n281_14(.douta(w_n281_14[0]),.doutb(w_n281_14[1]),.doutc(w_n281_14[2]),.din(w_n281_4[1]));
	jspl3 jspl3_w_n281_15(.douta(w_n281_15[0]),.doutb(w_n281_15[1]),.doutc(w_n281_15[2]),.din(w_n281_4[2]));
	jspl3 jspl3_w_n281_16(.douta(w_n281_16[0]),.doutb(w_n281_16[1]),.doutc(w_n281_16[2]),.din(w_n281_5[0]));
	jspl3 jspl3_w_n281_17(.douta(w_n281_17[0]),.doutb(w_n281_17[1]),.doutc(w_n281_17[2]),.din(w_n281_5[1]));
	jspl3 jspl3_w_n281_18(.douta(w_n281_18[0]),.doutb(w_n281_18[1]),.doutc(w_n281_18[2]),.din(w_n281_5[2]));
	jspl3 jspl3_w_n281_19(.douta(w_n281_19[0]),.doutb(w_n281_19[1]),.doutc(w_n281_19[2]),.din(w_n281_6[0]));
	jspl3 jspl3_w_n281_20(.douta(w_n281_20[0]),.doutb(w_n281_20[1]),.doutc(w_n281_20[2]),.din(w_n281_6[1]));
	jspl3 jspl3_w_n281_21(.douta(w_n281_21[0]),.doutb(w_n281_21[1]),.doutc(w_n281_21[2]),.din(w_n281_6[2]));
	jspl3 jspl3_w_n281_22(.douta(w_n281_22[0]),.doutb(w_n281_22[1]),.doutc(w_n281_22[2]),.din(w_n281_7[0]));
	jspl3 jspl3_w_n281_23(.douta(w_n281_23[0]),.doutb(w_n281_23[1]),.doutc(w_n281_23[2]),.din(w_n281_7[1]));
	jspl3 jspl3_w_n281_24(.douta(w_n281_24[0]),.doutb(w_n281_24[1]),.doutc(w_n281_24[2]),.din(w_n281_7[2]));
	jspl3 jspl3_w_n281_25(.douta(w_n281_25[0]),.doutb(w_n281_25[1]),.doutc(w_n281_25[2]),.din(w_n281_8[0]));
	jspl3 jspl3_w_n281_26(.douta(w_n281_26[0]),.doutb(w_n281_26[1]),.doutc(w_n281_26[2]),.din(w_n281_8[1]));
	jspl3 jspl3_w_n281_27(.douta(w_n281_27[0]),.doutb(w_n281_27[1]),.doutc(w_n281_27[2]),.din(w_n281_8[2]));
	jspl3 jspl3_w_n281_28(.douta(w_n281_28[0]),.doutb(w_n281_28[1]),.doutc(w_n281_28[2]),.din(w_n281_9[0]));
	jspl3 jspl3_w_n281_29(.douta(w_n281_29[0]),.doutb(w_n281_29[1]),.doutc(w_n281_29[2]),.din(w_n281_9[1]));
	jspl3 jspl3_w_n281_30(.douta(w_n281_30[0]),.doutb(w_n281_30[1]),.doutc(w_n281_30[2]),.din(w_n281_9[2]));
	jspl3 jspl3_w_n281_31(.douta(w_n281_31[0]),.doutb(w_n281_31[1]),.doutc(w_n281_31[2]),.din(w_n281_10[0]));
	jspl3 jspl3_w_n281_32(.douta(w_n281_32[0]),.doutb(w_n281_32[1]),.doutc(w_n281_32[2]),.din(w_n281_10[1]));
	jspl3 jspl3_w_n281_33(.douta(w_n281_33[0]),.doutb(w_n281_33[1]),.doutc(w_n281_33[2]),.din(w_n281_10[2]));
	jspl3 jspl3_w_n281_34(.douta(w_n281_34[0]),.doutb(w_n281_34[1]),.doutc(w_n281_34[2]),.din(w_n281_11[0]));
	jspl3 jspl3_w_n281_35(.douta(w_n281_35[0]),.doutb(w_n281_35[1]),.doutc(w_n281_35[2]),.din(w_n281_11[1]));
	jspl3 jspl3_w_n281_36(.douta(w_n281_36[0]),.doutb(w_n281_36[1]),.doutc(w_n281_36[2]),.din(w_n281_11[2]));
	jspl3 jspl3_w_n281_37(.douta(w_n281_37[0]),.doutb(w_n281_37[1]),.doutc(w_n281_37[2]),.din(w_n281_12[0]));
	jspl3 jspl3_w_n281_38(.douta(w_n281_38[0]),.doutb(w_n281_38[1]),.doutc(w_n281_38[2]),.din(w_n281_12[1]));
	jspl3 jspl3_w_n281_39(.douta(w_n281_39[0]),.doutb(w_n281_39[1]),.doutc(w_n281_39[2]),.din(w_n281_12[2]));
	jspl3 jspl3_w_n281_40(.douta(w_n281_40[0]),.doutb(w_n281_40[1]),.doutc(w_n281_40[2]),.din(w_n281_13[0]));
	jspl3 jspl3_w_n281_41(.douta(w_n281_41[0]),.doutb(w_n281_41[1]),.doutc(w_n281_41[2]),.din(w_n281_13[1]));
	jspl3 jspl3_w_n281_42(.douta(w_n281_42[0]),.doutb(w_n281_42[1]),.doutc(w_n281_42[2]),.din(w_n281_13[2]));
	jspl3 jspl3_w_n281_43(.douta(w_n281_43[0]),.doutb(w_n281_43[1]),.doutc(w_n281_43[2]),.din(w_n281_14[0]));
	jspl3 jspl3_w_n281_44(.douta(w_n281_44[0]),.doutb(w_n281_44[1]),.doutc(w_n281_44[2]),.din(w_n281_14[1]));
	jspl3 jspl3_w_n281_45(.douta(w_n281_45[0]),.doutb(w_n281_45[1]),.doutc(w_n281_45[2]),.din(w_n281_14[2]));
	jspl3 jspl3_w_n281_46(.douta(w_n281_46[0]),.doutb(w_n281_46[1]),.doutc(w_n281_46[2]),.din(w_n281_15[0]));
	jspl3 jspl3_w_n281_47(.douta(w_n281_47[0]),.doutb(w_n281_47[1]),.doutc(w_n281_47[2]),.din(w_n281_15[1]));
	jspl3 jspl3_w_n281_48(.douta(w_n281_48[0]),.doutb(w_n281_48[1]),.doutc(w_n281_48[2]),.din(w_n281_15[2]));
	jspl3 jspl3_w_n281_49(.douta(w_n281_49[0]),.doutb(w_n281_49[1]),.doutc(w_n281_49[2]),.din(w_n281_16[0]));
	jspl3 jspl3_w_n281_50(.douta(w_n281_50[0]),.doutb(w_n281_50[1]),.doutc(w_n281_50[2]),.din(w_n281_16[1]));
	jspl3 jspl3_w_n281_51(.douta(w_n281_51[0]),.doutb(w_n281_51[1]),.doutc(w_n281_51[2]),.din(w_n281_16[2]));
	jspl3 jspl3_w_n281_52(.douta(w_n281_52[0]),.doutb(w_n281_52[1]),.doutc(w_n281_52[2]),.din(w_n281_17[0]));
	jspl3 jspl3_w_n281_53(.douta(w_n281_53[0]),.doutb(w_n281_53[1]),.doutc(w_n281_53[2]),.din(w_n281_17[1]));
	jspl3 jspl3_w_n281_54(.douta(w_n281_54[0]),.doutb(w_n281_54[1]),.doutc(w_n281_54[2]),.din(w_n281_17[2]));
	jspl3 jspl3_w_n281_55(.douta(w_n281_55[0]),.doutb(w_n281_55[1]),.doutc(w_n281_55[2]),.din(w_n281_18[0]));
	jspl3 jspl3_w_n281_56(.douta(w_n281_56[0]),.doutb(w_n281_56[1]),.doutc(w_n281_56[2]),.din(w_n281_18[1]));
	jspl3 jspl3_w_n281_57(.douta(w_n281_57[0]),.doutb(w_n281_57[1]),.doutc(w_n281_57[2]),.din(w_n281_18[2]));
	jspl3 jspl3_w_n281_58(.douta(w_n281_58[0]),.doutb(w_n281_58[1]),.doutc(w_n281_58[2]),.din(w_n281_19[0]));
	jspl3 jspl3_w_n281_59(.douta(w_n281_59[0]),.doutb(w_n281_59[1]),.doutc(w_n281_59[2]),.din(w_n281_19[1]));
	jspl3 jspl3_w_n281_60(.douta(w_n281_60[0]),.doutb(w_n281_60[1]),.doutc(w_n281_60[2]),.din(w_n281_19[2]));
	jspl3 jspl3_w_n281_61(.douta(w_n281_61[0]),.doutb(w_n281_61[1]),.doutc(w_n281_61[2]),.din(w_n281_20[0]));
	jspl3 jspl3_w_n281_62(.douta(w_n281_62[0]),.doutb(w_n281_62[1]),.doutc(w_n281_62[2]),.din(w_n281_20[1]));
	jspl jspl_w_n281_63(.douta(w_n281_63[0]),.doutb(w_n281_63[1]),.din(w_n281_20[2]));
	jspl jspl_w_n284_0(.douta(w_n284_0[0]),.doutb(w_n284_0[1]),.din(n284));
	jspl jspl_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.din(n288));
	jspl3 jspl3_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.doutc(w_n290_0[2]),.din(n290));
	jspl jspl_w_n290_1(.douta(w_n290_1[0]),.doutb(w_n290_1[1]),.din(w_n290_0[0]));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(w_dff_B_H2R9KPX95_3));
	jspl3 jspl3_w_n292_1(.douta(w_n292_1[0]),.doutb(w_n292_1[1]),.doutc(w_n292_1[2]),.din(w_n292_0[0]));
	jspl3 jspl3_w_n292_2(.douta(w_n292_2[0]),.doutb(w_n292_2[1]),.doutc(w_n292_2[2]),.din(w_n292_0[1]));
	jspl3 jspl3_w_n292_3(.douta(w_n292_3[0]),.doutb(w_n292_3[1]),.doutc(w_n292_3[2]),.din(w_n292_0[2]));
	jspl3 jspl3_w_n292_4(.douta(w_n292_4[0]),.doutb(w_n292_4[1]),.doutc(w_n292_4[2]),.din(w_n292_1[0]));
	jspl3 jspl3_w_n292_5(.douta(w_n292_5[0]),.doutb(w_n292_5[1]),.doutc(w_n292_5[2]),.din(w_n292_1[1]));
	jspl3 jspl3_w_n292_6(.douta(w_n292_6[0]),.doutb(w_n292_6[1]),.doutc(w_n292_6[2]),.din(w_n292_1[2]));
	jspl3 jspl3_w_n292_7(.douta(w_n292_7[0]),.doutb(w_n292_7[1]),.doutc(w_n292_7[2]),.din(w_n292_2[0]));
	jspl3 jspl3_w_n292_8(.douta(w_n292_8[0]),.doutb(w_n292_8[1]),.doutc(w_n292_8[2]),.din(w_n292_2[1]));
	jspl3 jspl3_w_n292_9(.douta(w_n292_9[0]),.doutb(w_n292_9[1]),.doutc(w_n292_9[2]),.din(w_n292_2[2]));
	jspl3 jspl3_w_n292_10(.douta(w_n292_10[0]),.doutb(w_n292_10[1]),.doutc(w_n292_10[2]),.din(w_n292_3[0]));
	jspl3 jspl3_w_n292_11(.douta(w_n292_11[0]),.doutb(w_n292_11[1]),.doutc(w_n292_11[2]),.din(w_n292_3[1]));
	jspl3 jspl3_w_n292_12(.douta(w_n292_12[0]),.doutb(w_n292_12[1]),.doutc(w_n292_12[2]),.din(w_n292_3[2]));
	jspl3 jspl3_w_n292_13(.douta(w_n292_13[0]),.doutb(w_n292_13[1]),.doutc(w_n292_13[2]),.din(w_n292_4[0]));
	jspl3 jspl3_w_n292_14(.douta(w_n292_14[0]),.doutb(w_n292_14[1]),.doutc(w_n292_14[2]),.din(w_n292_4[1]));
	jspl3 jspl3_w_n292_15(.douta(w_n292_15[0]),.doutb(w_n292_15[1]),.doutc(w_n292_15[2]),.din(w_n292_4[2]));
	jspl3 jspl3_w_n292_16(.douta(w_n292_16[0]),.doutb(w_n292_16[1]),.doutc(w_n292_16[2]),.din(w_n292_5[0]));
	jspl3 jspl3_w_n292_17(.douta(w_n292_17[0]),.doutb(w_n292_17[1]),.doutc(w_n292_17[2]),.din(w_n292_5[1]));
	jspl3 jspl3_w_n292_18(.douta(w_n292_18[0]),.doutb(w_n292_18[1]),.doutc(w_n292_18[2]),.din(w_n292_5[2]));
	jspl3 jspl3_w_n292_19(.douta(w_n292_19[0]),.doutb(w_n292_19[1]),.doutc(w_n292_19[2]),.din(w_n292_6[0]));
	jspl3 jspl3_w_n292_20(.douta(w_n292_20[0]),.doutb(w_n292_20[1]),.doutc(w_n292_20[2]),.din(w_n292_6[1]));
	jspl3 jspl3_w_n292_21(.douta(w_n292_21[0]),.doutb(w_n292_21[1]),.doutc(w_n292_21[2]),.din(w_n292_6[2]));
	jspl3 jspl3_w_n292_22(.douta(w_n292_22[0]),.doutb(w_n292_22[1]),.doutc(w_n292_22[2]),.din(w_n292_7[0]));
	jspl3 jspl3_w_n292_23(.douta(w_n292_23[0]),.doutb(w_n292_23[1]),.doutc(w_n292_23[2]),.din(w_n292_7[1]));
	jspl3 jspl3_w_n292_24(.douta(w_n292_24[0]),.doutb(w_n292_24[1]),.doutc(w_n292_24[2]),.din(w_n292_7[2]));
	jspl3 jspl3_w_n292_25(.douta(w_n292_25[0]),.doutb(w_n292_25[1]),.doutc(w_n292_25[2]),.din(w_n292_8[0]));
	jspl3 jspl3_w_n292_26(.douta(w_n292_26[0]),.doutb(w_n292_26[1]),.doutc(w_n292_26[2]),.din(w_n292_8[1]));
	jspl3 jspl3_w_n292_27(.douta(w_n292_27[0]),.doutb(w_n292_27[1]),.doutc(w_n292_27[2]),.din(w_n292_8[2]));
	jspl3 jspl3_w_n292_28(.douta(w_n292_28[0]),.doutb(w_n292_28[1]),.doutc(w_n292_28[2]),.din(w_n292_9[0]));
	jspl3 jspl3_w_n292_29(.douta(w_n292_29[0]),.doutb(w_n292_29[1]),.doutc(w_n292_29[2]),.din(w_n292_9[1]));
	jspl3 jspl3_w_n292_30(.douta(w_n292_30[0]),.doutb(w_n292_30[1]),.doutc(w_n292_30[2]),.din(w_n292_9[2]));
	jspl3 jspl3_w_n292_31(.douta(w_n292_31[0]),.doutb(w_n292_31[1]),.doutc(w_n292_31[2]),.din(w_n292_10[0]));
	jspl3 jspl3_w_n292_32(.douta(w_n292_32[0]),.doutb(w_n292_32[1]),.doutc(w_n292_32[2]),.din(w_n292_10[1]));
	jspl3 jspl3_w_n292_33(.douta(w_n292_33[0]),.doutb(w_n292_33[1]),.doutc(w_n292_33[2]),.din(w_n292_10[2]));
	jspl3 jspl3_w_n292_34(.douta(w_n292_34[0]),.doutb(w_n292_34[1]),.doutc(w_n292_34[2]),.din(w_n292_11[0]));
	jspl3 jspl3_w_n292_35(.douta(w_n292_35[0]),.doutb(w_n292_35[1]),.doutc(w_n292_35[2]),.din(w_n292_11[1]));
	jspl3 jspl3_w_n292_36(.douta(w_n292_36[0]),.doutb(w_n292_36[1]),.doutc(w_n292_36[2]),.din(w_n292_11[2]));
	jspl3 jspl3_w_n292_37(.douta(w_n292_37[0]),.doutb(w_n292_37[1]),.doutc(w_n292_37[2]),.din(w_n292_12[0]));
	jspl3 jspl3_w_n292_38(.douta(w_n292_38[0]),.doutb(w_n292_38[1]),.doutc(w_n292_38[2]),.din(w_n292_12[1]));
	jspl3 jspl3_w_n292_39(.douta(w_n292_39[0]),.doutb(w_n292_39[1]),.doutc(w_n292_39[2]),.din(w_n292_12[2]));
	jspl3 jspl3_w_n292_40(.douta(w_n292_40[0]),.doutb(w_n292_40[1]),.doutc(w_n292_40[2]),.din(w_n292_13[0]));
	jspl3 jspl3_w_n292_41(.douta(w_n292_41[0]),.doutb(w_n292_41[1]),.doutc(w_n292_41[2]),.din(w_n292_13[1]));
	jspl3 jspl3_w_n292_42(.douta(w_n292_42[0]),.doutb(w_n292_42[1]),.doutc(w_n292_42[2]),.din(w_n292_13[2]));
	jspl3 jspl3_w_n292_43(.douta(w_n292_43[0]),.doutb(w_n292_43[1]),.doutc(w_n292_43[2]),.din(w_n292_14[0]));
	jspl3 jspl3_w_n292_44(.douta(w_n292_44[0]),.doutb(w_n292_44[1]),.doutc(w_n292_44[2]),.din(w_n292_14[1]));
	jspl3 jspl3_w_n292_45(.douta(w_n292_45[0]),.doutb(w_n292_45[1]),.doutc(w_n292_45[2]),.din(w_n292_14[2]));
	jspl3 jspl3_w_n292_46(.douta(w_n292_46[0]),.doutb(w_n292_46[1]),.doutc(w_n292_46[2]),.din(w_n292_15[0]));
	jspl3 jspl3_w_n292_47(.douta(w_n292_47[0]),.doutb(w_n292_47[1]),.doutc(w_n292_47[2]),.din(w_n292_15[1]));
	jspl3 jspl3_w_n292_48(.douta(w_n292_48[0]),.doutb(w_n292_48[1]),.doutc(w_n292_48[2]),.din(w_n292_15[2]));
	jspl3 jspl3_w_n292_49(.douta(w_n292_49[0]),.doutb(w_n292_49[1]),.doutc(w_n292_49[2]),.din(w_n292_16[0]));
	jspl3 jspl3_w_n292_50(.douta(w_n292_50[0]),.doutb(w_n292_50[1]),.doutc(w_n292_50[2]),.din(w_n292_16[1]));
	jspl3 jspl3_w_n292_51(.douta(w_n292_51[0]),.doutb(w_n292_51[1]),.doutc(w_n292_51[2]),.din(w_n292_16[2]));
	jspl3 jspl3_w_n292_52(.douta(w_n292_52[0]),.doutb(w_n292_52[1]),.doutc(w_n292_52[2]),.din(w_n292_17[0]));
	jspl3 jspl3_w_n292_53(.douta(w_n292_53[0]),.doutb(w_n292_53[1]),.doutc(w_n292_53[2]),.din(w_n292_17[1]));
	jspl3 jspl3_w_n292_54(.douta(w_n292_54[0]),.doutb(w_n292_54[1]),.doutc(w_n292_54[2]),.din(w_n292_17[2]));
	jspl3 jspl3_w_n292_55(.douta(w_n292_55[0]),.doutb(w_n292_55[1]),.doutc(w_n292_55[2]),.din(w_n292_18[0]));
	jspl3 jspl3_w_n292_56(.douta(w_n292_56[0]),.doutb(w_n292_56[1]),.doutc(w_n292_56[2]),.din(w_n292_18[1]));
	jspl3 jspl3_w_n292_57(.douta(w_n292_57[0]),.doutb(w_n292_57[1]),.doutc(w_n292_57[2]),.din(w_n292_18[2]));
	jspl3 jspl3_w_n292_58(.douta(w_n292_58[0]),.doutb(w_n292_58[1]),.doutc(w_n292_58[2]),.din(w_n292_19[0]));
	jspl3 jspl3_w_n292_59(.douta(w_n292_59[0]),.doutb(w_n292_59[1]),.doutc(w_n292_59[2]),.din(w_n292_19[1]));
	jspl3 jspl3_w_n292_60(.douta(w_n292_60[0]),.doutb(w_n292_60[1]),.doutc(w_n292_60[2]),.din(w_n292_19[2]));
	jspl3 jspl3_w_n292_61(.douta(w_n292_61[0]),.doutb(w_n292_61[1]),.doutc(w_n292_61[2]),.din(w_n292_20[0]));
	jspl3 jspl3_w_n292_62(.douta(w_n292_62[0]),.doutb(w_n292_62[1]),.doutc(w_n292_62[2]),.din(w_n292_20[1]));
	jspl jspl_w_n292_63(.douta(w_n292_63[0]),.doutb(w_n292_63[1]),.din(w_n292_20[2]));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(n295));
	jspl jspl_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.din(n299));
	jspl3 jspl3_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.doutc(w_n301_0[2]),.din(n301));
	jspl jspl_w_n301_1(.douta(w_n301_1[0]),.doutb(w_n301_1[1]),.din(w_n301_0[0]));
	jspl3 jspl3_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.doutc(w_n304_0[2]),.din(w_dff_B_L3XqwQjn4_3));
	jspl3 jspl3_w_n304_1(.douta(w_n304_1[0]),.doutb(w_n304_1[1]),.doutc(w_n304_1[2]),.din(w_n304_0[0]));
	jspl3 jspl3_w_n304_2(.douta(w_n304_2[0]),.doutb(w_n304_2[1]),.doutc(w_n304_2[2]),.din(w_n304_0[1]));
	jspl3 jspl3_w_n304_3(.douta(w_n304_3[0]),.doutb(w_n304_3[1]),.doutc(w_n304_3[2]),.din(w_n304_0[2]));
	jspl3 jspl3_w_n304_4(.douta(w_n304_4[0]),.doutb(w_n304_4[1]),.doutc(w_n304_4[2]),.din(w_n304_1[0]));
	jspl3 jspl3_w_n304_5(.douta(w_n304_5[0]),.doutb(w_n304_5[1]),.doutc(w_n304_5[2]),.din(w_n304_1[1]));
	jspl3 jspl3_w_n304_6(.douta(w_n304_6[0]),.doutb(w_n304_6[1]),.doutc(w_n304_6[2]),.din(w_n304_1[2]));
	jspl3 jspl3_w_n304_7(.douta(w_n304_7[0]),.doutb(w_n304_7[1]),.doutc(w_n304_7[2]),.din(w_n304_2[0]));
	jspl3 jspl3_w_n304_8(.douta(w_n304_8[0]),.doutb(w_n304_8[1]),.doutc(w_n304_8[2]),.din(w_n304_2[1]));
	jspl3 jspl3_w_n304_9(.douta(w_n304_9[0]),.doutb(w_n304_9[1]),.doutc(w_n304_9[2]),.din(w_n304_2[2]));
	jspl3 jspl3_w_n304_10(.douta(w_n304_10[0]),.doutb(w_n304_10[1]),.doutc(w_n304_10[2]),.din(w_n304_3[0]));
	jspl3 jspl3_w_n304_11(.douta(w_n304_11[0]),.doutb(w_n304_11[1]),.doutc(w_n304_11[2]),.din(w_n304_3[1]));
	jspl3 jspl3_w_n304_12(.douta(w_n304_12[0]),.doutb(w_n304_12[1]),.doutc(w_n304_12[2]),.din(w_n304_3[2]));
	jspl3 jspl3_w_n304_13(.douta(w_n304_13[0]),.doutb(w_n304_13[1]),.doutc(w_n304_13[2]),.din(w_n304_4[0]));
	jspl3 jspl3_w_n304_14(.douta(w_n304_14[0]),.doutb(w_n304_14[1]),.doutc(w_n304_14[2]),.din(w_n304_4[1]));
	jspl3 jspl3_w_n304_15(.douta(w_n304_15[0]),.doutb(w_n304_15[1]),.doutc(w_n304_15[2]),.din(w_n304_4[2]));
	jspl3 jspl3_w_n304_16(.douta(w_n304_16[0]),.doutb(w_n304_16[1]),.doutc(w_n304_16[2]),.din(w_n304_5[0]));
	jspl3 jspl3_w_n304_17(.douta(w_n304_17[0]),.doutb(w_n304_17[1]),.doutc(w_n304_17[2]),.din(w_n304_5[1]));
	jspl3 jspl3_w_n304_18(.douta(w_n304_18[0]),.doutb(w_n304_18[1]),.doutc(w_n304_18[2]),.din(w_n304_5[2]));
	jspl3 jspl3_w_n304_19(.douta(w_n304_19[0]),.doutb(w_n304_19[1]),.doutc(w_n304_19[2]),.din(w_n304_6[0]));
	jspl3 jspl3_w_n304_20(.douta(w_n304_20[0]),.doutb(w_n304_20[1]),.doutc(w_n304_20[2]),.din(w_n304_6[1]));
	jspl3 jspl3_w_n304_21(.douta(w_n304_21[0]),.doutb(w_n304_21[1]),.doutc(w_n304_21[2]),.din(w_n304_6[2]));
	jspl3 jspl3_w_n304_22(.douta(w_n304_22[0]),.doutb(w_n304_22[1]),.doutc(w_n304_22[2]),.din(w_n304_7[0]));
	jspl3 jspl3_w_n304_23(.douta(w_n304_23[0]),.doutb(w_n304_23[1]),.doutc(w_n304_23[2]),.din(w_n304_7[1]));
	jspl3 jspl3_w_n304_24(.douta(w_n304_24[0]),.doutb(w_n304_24[1]),.doutc(w_n304_24[2]),.din(w_n304_7[2]));
	jspl3 jspl3_w_n304_25(.douta(w_n304_25[0]),.doutb(w_n304_25[1]),.doutc(w_n304_25[2]),.din(w_n304_8[0]));
	jspl3 jspl3_w_n304_26(.douta(w_n304_26[0]),.doutb(w_n304_26[1]),.doutc(w_n304_26[2]),.din(w_n304_8[1]));
	jspl3 jspl3_w_n304_27(.douta(w_n304_27[0]),.doutb(w_n304_27[1]),.doutc(w_n304_27[2]),.din(w_n304_8[2]));
	jspl3 jspl3_w_n304_28(.douta(w_n304_28[0]),.doutb(w_n304_28[1]),.doutc(w_n304_28[2]),.din(w_n304_9[0]));
	jspl3 jspl3_w_n304_29(.douta(w_n304_29[0]),.doutb(w_n304_29[1]),.doutc(w_n304_29[2]),.din(w_n304_9[1]));
	jspl3 jspl3_w_n304_30(.douta(w_n304_30[0]),.doutb(w_n304_30[1]),.doutc(w_n304_30[2]),.din(w_n304_9[2]));
	jspl3 jspl3_w_n304_31(.douta(w_n304_31[0]),.doutb(w_n304_31[1]),.doutc(w_n304_31[2]),.din(w_n304_10[0]));
	jspl3 jspl3_w_n304_32(.douta(w_n304_32[0]),.doutb(w_n304_32[1]),.doutc(w_n304_32[2]),.din(w_n304_10[1]));
	jspl3 jspl3_w_n304_33(.douta(w_n304_33[0]),.doutb(w_n304_33[1]),.doutc(w_n304_33[2]),.din(w_n304_10[2]));
	jspl3 jspl3_w_n304_34(.douta(w_n304_34[0]),.doutb(w_n304_34[1]),.doutc(w_n304_34[2]),.din(w_n304_11[0]));
	jspl3 jspl3_w_n304_35(.douta(w_n304_35[0]),.doutb(w_n304_35[1]),.doutc(w_n304_35[2]),.din(w_n304_11[1]));
	jspl3 jspl3_w_n304_36(.douta(w_n304_36[0]),.doutb(w_n304_36[1]),.doutc(w_n304_36[2]),.din(w_n304_11[2]));
	jspl3 jspl3_w_n304_37(.douta(w_n304_37[0]),.doutb(w_n304_37[1]),.doutc(w_n304_37[2]),.din(w_n304_12[0]));
	jspl3 jspl3_w_n304_38(.douta(w_n304_38[0]),.doutb(w_n304_38[1]),.doutc(w_n304_38[2]),.din(w_n304_12[1]));
	jspl3 jspl3_w_n304_39(.douta(w_n304_39[0]),.doutb(w_n304_39[1]),.doutc(w_n304_39[2]),.din(w_n304_12[2]));
	jspl3 jspl3_w_n304_40(.douta(w_n304_40[0]),.doutb(w_n304_40[1]),.doutc(w_n304_40[2]),.din(w_n304_13[0]));
	jspl3 jspl3_w_n304_41(.douta(w_n304_41[0]),.doutb(w_n304_41[1]),.doutc(w_n304_41[2]),.din(w_n304_13[1]));
	jspl3 jspl3_w_n304_42(.douta(w_n304_42[0]),.doutb(w_n304_42[1]),.doutc(w_n304_42[2]),.din(w_n304_13[2]));
	jspl3 jspl3_w_n304_43(.douta(w_n304_43[0]),.doutb(w_n304_43[1]),.doutc(w_n304_43[2]),.din(w_n304_14[0]));
	jspl3 jspl3_w_n304_44(.douta(w_n304_44[0]),.doutb(w_n304_44[1]),.doutc(w_n304_44[2]),.din(w_n304_14[1]));
	jspl3 jspl3_w_n304_45(.douta(w_n304_45[0]),.doutb(w_n304_45[1]),.doutc(w_n304_45[2]),.din(w_n304_14[2]));
	jspl3 jspl3_w_n304_46(.douta(w_n304_46[0]),.doutb(w_n304_46[1]),.doutc(w_n304_46[2]),.din(w_n304_15[0]));
	jspl3 jspl3_w_n304_47(.douta(w_n304_47[0]),.doutb(w_n304_47[1]),.doutc(w_n304_47[2]),.din(w_n304_15[1]));
	jspl3 jspl3_w_n304_48(.douta(w_n304_48[0]),.doutb(w_n304_48[1]),.doutc(w_n304_48[2]),.din(w_n304_15[2]));
	jspl3 jspl3_w_n304_49(.douta(w_n304_49[0]),.doutb(w_n304_49[1]),.doutc(w_n304_49[2]),.din(w_n304_16[0]));
	jspl3 jspl3_w_n304_50(.douta(w_n304_50[0]),.doutb(w_n304_50[1]),.doutc(w_n304_50[2]),.din(w_n304_16[1]));
	jspl3 jspl3_w_n304_51(.douta(w_n304_51[0]),.doutb(w_n304_51[1]),.doutc(w_n304_51[2]),.din(w_n304_16[2]));
	jspl3 jspl3_w_n304_52(.douta(w_n304_52[0]),.doutb(w_n304_52[1]),.doutc(w_n304_52[2]),.din(w_n304_17[0]));
	jspl3 jspl3_w_n304_53(.douta(w_n304_53[0]),.doutb(w_n304_53[1]),.doutc(w_n304_53[2]),.din(w_n304_17[1]));
	jspl3 jspl3_w_n304_54(.douta(w_n304_54[0]),.doutb(w_n304_54[1]),.doutc(w_n304_54[2]),.din(w_n304_17[2]));
	jspl3 jspl3_w_n304_55(.douta(w_n304_55[0]),.doutb(w_n304_55[1]),.doutc(w_n304_55[2]),.din(w_n304_18[0]));
	jspl3 jspl3_w_n304_56(.douta(w_n304_56[0]),.doutb(w_n304_56[1]),.doutc(w_n304_56[2]),.din(w_n304_18[1]));
	jspl3 jspl3_w_n304_57(.douta(w_n304_57[0]),.doutb(w_n304_57[1]),.doutc(w_n304_57[2]),.din(w_n304_18[2]));
	jspl3 jspl3_w_n304_58(.douta(w_n304_58[0]),.doutb(w_n304_58[1]),.doutc(w_n304_58[2]),.din(w_n304_19[0]));
	jspl3 jspl3_w_n304_59(.douta(w_n304_59[0]),.doutb(w_n304_59[1]),.doutc(w_n304_59[2]),.din(w_n304_19[1]));
	jspl3 jspl3_w_n304_60(.douta(w_n304_60[0]),.doutb(w_n304_60[1]),.doutc(w_n304_60[2]),.din(w_n304_19[2]));
	jspl3 jspl3_w_n304_61(.douta(w_n304_61[0]),.doutb(w_n304_61[1]),.doutc(w_n304_61[2]),.din(w_n304_20[0]));
	jspl3 jspl3_w_n304_62(.douta(w_n304_62[0]),.doutb(w_n304_62[1]),.doutc(w_n304_62[2]),.din(w_n304_20[1]));
	jspl jspl_w_n304_63(.douta(w_n304_63[0]),.doutb(w_n304_63[1]),.din(w_n304_20[2]));
	jspl jspl_w_n307_0(.douta(w_n307_0[0]),.doutb(w_n307_0[1]),.din(n307));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl3 jspl3_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.doutc(w_n313_0[2]),.din(n313));
	jspl jspl_w_n313_1(.douta(w_n313_1[0]),.doutb(w_n313_1[1]),.din(w_n313_0[0]));
	jspl3 jspl3_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.doutc(w_n316_0[2]),.din(n316));
	jspl jspl_w_n316_1(.douta(w_n316_1[0]),.doutb(w_n316_1[1]),.din(w_n316_0[0]));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.doutc(w_n319_0[2]),.din(w_dff_B_ypPvMaYr6_3));
	jspl3 jspl3_w_n319_1(.douta(w_n319_1[0]),.doutb(w_n319_1[1]),.doutc(w_n319_1[2]),.din(w_n319_0[0]));
	jspl3 jspl3_w_n319_2(.douta(w_n319_2[0]),.doutb(w_n319_2[1]),.doutc(w_n319_2[2]),.din(w_n319_0[1]));
	jspl3 jspl3_w_n319_3(.douta(w_n319_3[0]),.doutb(w_n319_3[1]),.doutc(w_n319_3[2]),.din(w_n319_0[2]));
	jspl3 jspl3_w_n319_4(.douta(w_n319_4[0]),.doutb(w_n319_4[1]),.doutc(w_n319_4[2]),.din(w_n319_1[0]));
	jspl3 jspl3_w_n319_5(.douta(w_n319_5[0]),.doutb(w_n319_5[1]),.doutc(w_n319_5[2]),.din(w_n319_1[1]));
	jspl3 jspl3_w_n319_6(.douta(w_n319_6[0]),.doutb(w_n319_6[1]),.doutc(w_n319_6[2]),.din(w_n319_1[2]));
	jspl3 jspl3_w_n319_7(.douta(w_n319_7[0]),.doutb(w_n319_7[1]),.doutc(w_n319_7[2]),.din(w_n319_2[0]));
	jspl3 jspl3_w_n319_8(.douta(w_n319_8[0]),.doutb(w_n319_8[1]),.doutc(w_n319_8[2]),.din(w_n319_2[1]));
	jspl3 jspl3_w_n319_9(.douta(w_n319_9[0]),.doutb(w_n319_9[1]),.doutc(w_n319_9[2]),.din(w_n319_2[2]));
	jspl3 jspl3_w_n319_10(.douta(w_n319_10[0]),.doutb(w_n319_10[1]),.doutc(w_n319_10[2]),.din(w_n319_3[0]));
	jspl3 jspl3_w_n319_11(.douta(w_n319_11[0]),.doutb(w_n319_11[1]),.doutc(w_n319_11[2]),.din(w_n319_3[1]));
	jspl3 jspl3_w_n319_12(.douta(w_n319_12[0]),.doutb(w_n319_12[1]),.doutc(w_n319_12[2]),.din(w_n319_3[2]));
	jspl3 jspl3_w_n319_13(.douta(w_n319_13[0]),.doutb(w_n319_13[1]),.doutc(w_n319_13[2]),.din(w_n319_4[0]));
	jspl3 jspl3_w_n319_14(.douta(w_n319_14[0]),.doutb(w_n319_14[1]),.doutc(w_n319_14[2]),.din(w_n319_4[1]));
	jspl3 jspl3_w_n319_15(.douta(w_n319_15[0]),.doutb(w_n319_15[1]),.doutc(w_n319_15[2]),.din(w_n319_4[2]));
	jspl3 jspl3_w_n319_16(.douta(w_n319_16[0]),.doutb(w_n319_16[1]),.doutc(w_n319_16[2]),.din(w_n319_5[0]));
	jspl3 jspl3_w_n319_17(.douta(w_n319_17[0]),.doutb(w_n319_17[1]),.doutc(w_n319_17[2]),.din(w_n319_5[1]));
	jspl3 jspl3_w_n319_18(.douta(w_n319_18[0]),.doutb(w_n319_18[1]),.doutc(w_n319_18[2]),.din(w_n319_5[2]));
	jspl3 jspl3_w_n319_19(.douta(w_n319_19[0]),.doutb(w_n319_19[1]),.doutc(w_n319_19[2]),.din(w_n319_6[0]));
	jspl3 jspl3_w_n319_20(.douta(w_n319_20[0]),.doutb(w_n319_20[1]),.doutc(w_n319_20[2]),.din(w_n319_6[1]));
	jspl3 jspl3_w_n319_21(.douta(w_n319_21[0]),.doutb(w_n319_21[1]),.doutc(w_n319_21[2]),.din(w_n319_6[2]));
	jspl3 jspl3_w_n319_22(.douta(w_n319_22[0]),.doutb(w_n319_22[1]),.doutc(w_n319_22[2]),.din(w_n319_7[0]));
	jspl3 jspl3_w_n319_23(.douta(w_n319_23[0]),.doutb(w_n319_23[1]),.doutc(w_n319_23[2]),.din(w_n319_7[1]));
	jspl3 jspl3_w_n319_24(.douta(w_n319_24[0]),.doutb(w_n319_24[1]),.doutc(w_n319_24[2]),.din(w_n319_7[2]));
	jspl3 jspl3_w_n319_25(.douta(w_n319_25[0]),.doutb(w_n319_25[1]),.doutc(w_n319_25[2]),.din(w_n319_8[0]));
	jspl3 jspl3_w_n319_26(.douta(w_n319_26[0]),.doutb(w_n319_26[1]),.doutc(w_n319_26[2]),.din(w_n319_8[1]));
	jspl3 jspl3_w_n319_27(.douta(w_n319_27[0]),.doutb(w_n319_27[1]),.doutc(w_n319_27[2]),.din(w_n319_8[2]));
	jspl3 jspl3_w_n319_28(.douta(w_n319_28[0]),.doutb(w_n319_28[1]),.doutc(w_n319_28[2]),.din(w_n319_9[0]));
	jspl3 jspl3_w_n319_29(.douta(w_n319_29[0]),.doutb(w_n319_29[1]),.doutc(w_n319_29[2]),.din(w_n319_9[1]));
	jspl3 jspl3_w_n319_30(.douta(w_n319_30[0]),.doutb(w_n319_30[1]),.doutc(w_n319_30[2]),.din(w_n319_9[2]));
	jspl3 jspl3_w_n319_31(.douta(w_n319_31[0]),.doutb(w_n319_31[1]),.doutc(w_n319_31[2]),.din(w_n319_10[0]));
	jspl3 jspl3_w_n319_32(.douta(w_n319_32[0]),.doutb(w_n319_32[1]),.doutc(w_n319_32[2]),.din(w_n319_10[1]));
	jspl3 jspl3_w_n319_33(.douta(w_n319_33[0]),.doutb(w_n319_33[1]),.doutc(w_n319_33[2]),.din(w_n319_10[2]));
	jspl3 jspl3_w_n319_34(.douta(w_n319_34[0]),.doutb(w_n319_34[1]),.doutc(w_n319_34[2]),.din(w_n319_11[0]));
	jspl3 jspl3_w_n319_35(.douta(w_n319_35[0]),.doutb(w_n319_35[1]),.doutc(w_n319_35[2]),.din(w_n319_11[1]));
	jspl3 jspl3_w_n319_36(.douta(w_n319_36[0]),.doutb(w_n319_36[1]),.doutc(w_n319_36[2]),.din(w_n319_11[2]));
	jspl3 jspl3_w_n319_37(.douta(w_n319_37[0]),.doutb(w_n319_37[1]),.doutc(w_n319_37[2]),.din(w_n319_12[0]));
	jspl3 jspl3_w_n319_38(.douta(w_n319_38[0]),.doutb(w_n319_38[1]),.doutc(w_n319_38[2]),.din(w_n319_12[1]));
	jspl3 jspl3_w_n319_39(.douta(w_n319_39[0]),.doutb(w_n319_39[1]),.doutc(w_n319_39[2]),.din(w_n319_12[2]));
	jspl3 jspl3_w_n319_40(.douta(w_n319_40[0]),.doutb(w_n319_40[1]),.doutc(w_n319_40[2]),.din(w_n319_13[0]));
	jspl3 jspl3_w_n319_41(.douta(w_n319_41[0]),.doutb(w_n319_41[1]),.doutc(w_n319_41[2]),.din(w_n319_13[1]));
	jspl3 jspl3_w_n319_42(.douta(w_n319_42[0]),.doutb(w_n319_42[1]),.doutc(w_n319_42[2]),.din(w_n319_13[2]));
	jspl3 jspl3_w_n319_43(.douta(w_n319_43[0]),.doutb(w_n319_43[1]),.doutc(w_n319_43[2]),.din(w_n319_14[0]));
	jspl3 jspl3_w_n319_44(.douta(w_n319_44[0]),.doutb(w_n319_44[1]),.doutc(w_n319_44[2]),.din(w_n319_14[1]));
	jspl3 jspl3_w_n319_45(.douta(w_n319_45[0]),.doutb(w_n319_45[1]),.doutc(w_n319_45[2]),.din(w_n319_14[2]));
	jspl3 jspl3_w_n319_46(.douta(w_n319_46[0]),.doutb(w_n319_46[1]),.doutc(w_n319_46[2]),.din(w_n319_15[0]));
	jspl3 jspl3_w_n319_47(.douta(w_n319_47[0]),.doutb(w_n319_47[1]),.doutc(w_n319_47[2]),.din(w_n319_15[1]));
	jspl3 jspl3_w_n319_48(.douta(w_n319_48[0]),.doutb(w_n319_48[1]),.doutc(w_n319_48[2]),.din(w_n319_15[2]));
	jspl3 jspl3_w_n319_49(.douta(w_n319_49[0]),.doutb(w_n319_49[1]),.doutc(w_n319_49[2]),.din(w_n319_16[0]));
	jspl3 jspl3_w_n319_50(.douta(w_n319_50[0]),.doutb(w_n319_50[1]),.doutc(w_n319_50[2]),.din(w_n319_16[1]));
	jspl3 jspl3_w_n319_51(.douta(w_n319_51[0]),.doutb(w_n319_51[1]),.doutc(w_n319_51[2]),.din(w_n319_16[2]));
	jspl3 jspl3_w_n319_52(.douta(w_n319_52[0]),.doutb(w_n319_52[1]),.doutc(w_n319_52[2]),.din(w_n319_17[0]));
	jspl3 jspl3_w_n319_53(.douta(w_n319_53[0]),.doutb(w_n319_53[1]),.doutc(w_n319_53[2]),.din(w_n319_17[1]));
	jspl3 jspl3_w_n319_54(.douta(w_n319_54[0]),.doutb(w_n319_54[1]),.doutc(w_n319_54[2]),.din(w_n319_17[2]));
	jspl3 jspl3_w_n319_55(.douta(w_n319_55[0]),.doutb(w_n319_55[1]),.doutc(w_n319_55[2]),.din(w_n319_18[0]));
	jspl3 jspl3_w_n319_56(.douta(w_n319_56[0]),.doutb(w_n319_56[1]),.doutc(w_n319_56[2]),.din(w_n319_18[1]));
	jspl3 jspl3_w_n319_57(.douta(w_n319_57[0]),.doutb(w_n319_57[1]),.doutc(w_n319_57[2]),.din(w_n319_18[2]));
	jspl3 jspl3_w_n319_58(.douta(w_n319_58[0]),.doutb(w_n319_58[1]),.doutc(w_n319_58[2]),.din(w_n319_19[0]));
	jspl3 jspl3_w_n319_59(.douta(w_n319_59[0]),.doutb(w_n319_59[1]),.doutc(w_n319_59[2]),.din(w_n319_19[1]));
	jspl3 jspl3_w_n319_60(.douta(w_n319_60[0]),.doutb(w_n319_60[1]),.doutc(w_n319_60[2]),.din(w_n319_19[2]));
	jspl3 jspl3_w_n319_61(.douta(w_n319_61[0]),.doutb(w_n319_61[1]),.doutc(w_n319_61[2]),.din(w_n319_20[0]));
	jspl3 jspl3_w_n319_62(.douta(w_n319_62[0]),.doutb(w_n319_62[1]),.doutc(w_n319_62[2]),.din(w_n319_20[1]));
	jspl jspl_w_n319_63(.douta(w_n319_63[0]),.doutb(w_n319_63[1]),.din(w_n319_20[2]));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.din(n326));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n328_1(.douta(w_n328_1[0]),.doutb(w_n328_1[1]),.din(w_n328_0[0]));
	jspl jspl_w_n332_0(.douta(w_n332_0[0]),.doutb(w_n332_0[1]),.din(n332));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl3 jspl3_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.doutc(w_n338_0[2]),.din(n338));
	jspl jspl_w_n338_1(.douta(w_n338_1[0]),.doutb(w_n338_1[1]),.din(w_n338_0[0]));
	jspl jspl_w_n342_0(.douta(w_n342_0[0]),.doutb(w_n342_0[1]),.din(n342));
	jspl jspl_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.din(n346));
	jspl3 jspl3_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.doutc(w_n348_0[2]),.din(n348));
	jspl jspl_w_n348_1(.douta(w_n348_1[0]),.doutb(w_n348_1[1]),.din(w_n348_0[0]));
	jspl jspl_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.din(n353));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl3 jspl3_w_n359_0(.douta(w_n359_0[0]),.doutb(w_n359_0[1]),.doutc(w_n359_0[2]),.din(n359));
	jspl jspl_w_n359_1(.douta(w_n359_1[0]),.doutb(w_n359_1[1]),.din(w_n359_0[0]));
	jspl3 jspl3_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.doutc(w_n362_0[2]),.din(n362));
	jspl jspl_w_n362_1(.douta(w_n362_1[0]),.doutb(w_n362_1[1]),.din(w_n362_0[0]));
	jspl3 jspl3_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.doutc(w_n364_0[2]),.din(w_dff_B_cE1lYXHF5_3));
	jspl3 jspl3_w_n364_1(.douta(w_n364_1[0]),.doutb(w_n364_1[1]),.doutc(w_n364_1[2]),.din(w_n364_0[0]));
	jspl3 jspl3_w_n364_2(.douta(w_n364_2[0]),.doutb(w_n364_2[1]),.doutc(w_n364_2[2]),.din(w_n364_0[1]));
	jspl3 jspl3_w_n364_3(.douta(w_n364_3[0]),.doutb(w_n364_3[1]),.doutc(w_n364_3[2]),.din(w_n364_0[2]));
	jspl3 jspl3_w_n364_4(.douta(w_n364_4[0]),.doutb(w_n364_4[1]),.doutc(w_n364_4[2]),.din(w_n364_1[0]));
	jspl3 jspl3_w_n364_5(.douta(w_n364_5[0]),.doutb(w_n364_5[1]),.doutc(w_n364_5[2]),.din(w_n364_1[1]));
	jspl3 jspl3_w_n364_6(.douta(w_n364_6[0]),.doutb(w_n364_6[1]),.doutc(w_n364_6[2]),.din(w_n364_1[2]));
	jspl3 jspl3_w_n364_7(.douta(w_n364_7[0]),.doutb(w_n364_7[1]),.doutc(w_n364_7[2]),.din(w_n364_2[0]));
	jspl3 jspl3_w_n364_8(.douta(w_n364_8[0]),.doutb(w_n364_8[1]),.doutc(w_n364_8[2]),.din(w_n364_2[1]));
	jspl3 jspl3_w_n364_9(.douta(w_n364_9[0]),.doutb(w_n364_9[1]),.doutc(w_n364_9[2]),.din(w_n364_2[2]));
	jspl3 jspl3_w_n364_10(.douta(w_n364_10[0]),.doutb(w_n364_10[1]),.doutc(w_n364_10[2]),.din(w_n364_3[0]));
	jspl3 jspl3_w_n364_11(.douta(w_n364_11[0]),.doutb(w_n364_11[1]),.doutc(w_n364_11[2]),.din(w_n364_3[1]));
	jspl3 jspl3_w_n364_12(.douta(w_n364_12[0]),.doutb(w_n364_12[1]),.doutc(w_n364_12[2]),.din(w_n364_3[2]));
	jspl3 jspl3_w_n364_13(.douta(w_n364_13[0]),.doutb(w_n364_13[1]),.doutc(w_n364_13[2]),.din(w_n364_4[0]));
	jspl3 jspl3_w_n364_14(.douta(w_n364_14[0]),.doutb(w_n364_14[1]),.doutc(w_n364_14[2]),.din(w_n364_4[1]));
	jspl3 jspl3_w_n364_15(.douta(w_n364_15[0]),.doutb(w_n364_15[1]),.doutc(w_n364_15[2]),.din(w_n364_4[2]));
	jspl3 jspl3_w_n364_16(.douta(w_n364_16[0]),.doutb(w_n364_16[1]),.doutc(w_n364_16[2]),.din(w_n364_5[0]));
	jspl3 jspl3_w_n364_17(.douta(w_n364_17[0]),.doutb(w_n364_17[1]),.doutc(w_n364_17[2]),.din(w_n364_5[1]));
	jspl3 jspl3_w_n364_18(.douta(w_n364_18[0]),.doutb(w_n364_18[1]),.doutc(w_n364_18[2]),.din(w_n364_5[2]));
	jspl3 jspl3_w_n364_19(.douta(w_n364_19[0]),.doutb(w_n364_19[1]),.doutc(w_n364_19[2]),.din(w_n364_6[0]));
	jspl3 jspl3_w_n364_20(.douta(w_n364_20[0]),.doutb(w_n364_20[1]),.doutc(w_n364_20[2]),.din(w_n364_6[1]));
	jspl3 jspl3_w_n364_21(.douta(w_n364_21[0]),.doutb(w_n364_21[1]),.doutc(w_n364_21[2]),.din(w_n364_6[2]));
	jspl3 jspl3_w_n364_22(.douta(w_n364_22[0]),.doutb(w_n364_22[1]),.doutc(w_n364_22[2]),.din(w_n364_7[0]));
	jspl3 jspl3_w_n364_23(.douta(w_n364_23[0]),.doutb(w_n364_23[1]),.doutc(w_n364_23[2]),.din(w_n364_7[1]));
	jspl3 jspl3_w_n364_24(.douta(w_n364_24[0]),.doutb(w_n364_24[1]),.doutc(w_n364_24[2]),.din(w_n364_7[2]));
	jspl3 jspl3_w_n364_25(.douta(w_n364_25[0]),.doutb(w_n364_25[1]),.doutc(w_n364_25[2]),.din(w_n364_8[0]));
	jspl3 jspl3_w_n364_26(.douta(w_n364_26[0]),.doutb(w_n364_26[1]),.doutc(w_n364_26[2]),.din(w_n364_8[1]));
	jspl3 jspl3_w_n364_27(.douta(w_n364_27[0]),.doutb(w_n364_27[1]),.doutc(w_n364_27[2]),.din(w_n364_8[2]));
	jspl3 jspl3_w_n364_28(.douta(w_n364_28[0]),.doutb(w_n364_28[1]),.doutc(w_n364_28[2]),.din(w_n364_9[0]));
	jspl3 jspl3_w_n364_29(.douta(w_n364_29[0]),.doutb(w_n364_29[1]),.doutc(w_n364_29[2]),.din(w_n364_9[1]));
	jspl3 jspl3_w_n364_30(.douta(w_n364_30[0]),.doutb(w_n364_30[1]),.doutc(w_n364_30[2]),.din(w_n364_9[2]));
	jspl3 jspl3_w_n364_31(.douta(w_n364_31[0]),.doutb(w_n364_31[1]),.doutc(w_n364_31[2]),.din(w_n364_10[0]));
	jspl3 jspl3_w_n364_32(.douta(w_n364_32[0]),.doutb(w_n364_32[1]),.doutc(w_n364_32[2]),.din(w_n364_10[1]));
	jspl3 jspl3_w_n364_33(.douta(w_n364_33[0]),.doutb(w_n364_33[1]),.doutc(w_n364_33[2]),.din(w_n364_10[2]));
	jspl3 jspl3_w_n364_34(.douta(w_n364_34[0]),.doutb(w_n364_34[1]),.doutc(w_n364_34[2]),.din(w_n364_11[0]));
	jspl3 jspl3_w_n364_35(.douta(w_n364_35[0]),.doutb(w_n364_35[1]),.doutc(w_n364_35[2]),.din(w_n364_11[1]));
	jspl3 jspl3_w_n364_36(.douta(w_n364_36[0]),.doutb(w_n364_36[1]),.doutc(w_n364_36[2]),.din(w_n364_11[2]));
	jspl3 jspl3_w_n364_37(.douta(w_n364_37[0]),.doutb(w_n364_37[1]),.doutc(w_n364_37[2]),.din(w_n364_12[0]));
	jspl3 jspl3_w_n364_38(.douta(w_n364_38[0]),.doutb(w_n364_38[1]),.doutc(w_n364_38[2]),.din(w_n364_12[1]));
	jspl3 jspl3_w_n364_39(.douta(w_n364_39[0]),.doutb(w_n364_39[1]),.doutc(w_n364_39[2]),.din(w_n364_12[2]));
	jspl3 jspl3_w_n364_40(.douta(w_n364_40[0]),.doutb(w_n364_40[1]),.doutc(w_n364_40[2]),.din(w_n364_13[0]));
	jspl3 jspl3_w_n364_41(.douta(w_n364_41[0]),.doutb(w_n364_41[1]),.doutc(w_n364_41[2]),.din(w_n364_13[1]));
	jspl3 jspl3_w_n364_42(.douta(w_n364_42[0]),.doutb(w_n364_42[1]),.doutc(w_n364_42[2]),.din(w_n364_13[2]));
	jspl3 jspl3_w_n364_43(.douta(w_n364_43[0]),.doutb(w_n364_43[1]),.doutc(w_n364_43[2]),.din(w_n364_14[0]));
	jspl3 jspl3_w_n364_44(.douta(w_n364_44[0]),.doutb(w_n364_44[1]),.doutc(w_n364_44[2]),.din(w_n364_14[1]));
	jspl3 jspl3_w_n364_45(.douta(w_n364_45[0]),.doutb(w_n364_45[1]),.doutc(w_n364_45[2]),.din(w_n364_14[2]));
	jspl3 jspl3_w_n364_46(.douta(w_n364_46[0]),.doutb(w_n364_46[1]),.doutc(w_n364_46[2]),.din(w_n364_15[0]));
	jspl3 jspl3_w_n364_47(.douta(w_n364_47[0]),.doutb(w_n364_47[1]),.doutc(w_n364_47[2]),.din(w_n364_15[1]));
	jspl3 jspl3_w_n364_48(.douta(w_n364_48[0]),.doutb(w_n364_48[1]),.doutc(w_n364_48[2]),.din(w_n364_15[2]));
	jspl3 jspl3_w_n364_49(.douta(w_n364_49[0]),.doutb(w_n364_49[1]),.doutc(w_n364_49[2]),.din(w_n364_16[0]));
	jspl3 jspl3_w_n364_50(.douta(w_n364_50[0]),.doutb(w_n364_50[1]),.doutc(w_n364_50[2]),.din(w_n364_16[1]));
	jspl3 jspl3_w_n364_51(.douta(w_n364_51[0]),.doutb(w_n364_51[1]),.doutc(w_n364_51[2]),.din(w_n364_16[2]));
	jspl3 jspl3_w_n364_52(.douta(w_n364_52[0]),.doutb(w_n364_52[1]),.doutc(w_n364_52[2]),.din(w_n364_17[0]));
	jspl3 jspl3_w_n364_53(.douta(w_n364_53[0]),.doutb(w_n364_53[1]),.doutc(w_n364_53[2]),.din(w_n364_17[1]));
	jspl3 jspl3_w_n364_54(.douta(w_n364_54[0]),.doutb(w_n364_54[1]),.doutc(w_n364_54[2]),.din(w_n364_17[2]));
	jspl3 jspl3_w_n364_55(.douta(w_n364_55[0]),.doutb(w_n364_55[1]),.doutc(w_n364_55[2]),.din(w_n364_18[0]));
	jspl3 jspl3_w_n364_56(.douta(w_n364_56[0]),.doutb(w_n364_56[1]),.doutc(w_n364_56[2]),.din(w_n364_18[1]));
	jspl3 jspl3_w_n364_57(.douta(w_n364_57[0]),.doutb(w_n364_57[1]),.doutc(w_n364_57[2]),.din(w_n364_18[2]));
	jspl3 jspl3_w_n364_58(.douta(w_n364_58[0]),.doutb(w_n364_58[1]),.doutc(w_n364_58[2]),.din(w_n364_19[0]));
	jspl3 jspl3_w_n364_59(.douta(w_n364_59[0]),.doutb(w_n364_59[1]),.doutc(w_n364_59[2]),.din(w_n364_19[1]));
	jspl3 jspl3_w_n364_60(.douta(w_n364_60[0]),.doutb(w_n364_60[1]),.doutc(w_n364_60[2]),.din(w_n364_19[2]));
	jspl3 jspl3_w_n364_61(.douta(w_n364_61[0]),.doutb(w_n364_61[1]),.doutc(w_n364_61[2]),.din(w_n364_20[0]));
	jspl3 jspl3_w_n364_62(.douta(w_n364_62[0]),.doutb(w_n364_62[1]),.doutc(w_n364_62[2]),.din(w_n364_20[1]));
	jspl jspl_w_n364_63(.douta(w_n364_63[0]),.doutb(w_n364_63[1]),.din(w_n364_20[2]));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl3 jspl3_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.doutc(w_n373_0[2]),.din(n373));
	jspl jspl_w_n373_1(.douta(w_n373_1[0]),.doutb(w_n373_1[1]),.din(w_n373_0[0]));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.din(n377));
	jspl jspl_w_n381_0(.douta(w_n381_0[0]),.doutb(w_n381_0[1]),.din(n381));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl jspl_w_n383_1(.douta(w_n383_1[0]),.doutb(w_n383_1[1]),.din(w_n383_0[0]));
	jspl jspl_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.din(n387));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(n391));
	jspl3 jspl3_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.doutc(w_n393_0[2]),.din(n393));
	jspl jspl_w_n393_1(.douta(w_n393_1[0]),.doutb(w_n393_1[1]),.din(w_n393_0[0]));
	jspl jspl_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.din(n398));
	jspl jspl_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.din(n402));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl jspl_w_n404_1(.douta(w_n404_1[0]),.doutb(w_n404_1[1]),.din(w_n404_0[0]));
	jspl3 jspl3_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.doutc(w_n407_0[2]),.din(n407));
	jspl jspl_w_n407_1(.douta(w_n407_1[0]),.doutb(w_n407_1[1]),.din(w_n407_0[0]));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_n410_0[2]),.din(w_dff_B_F1l9p9yf4_3));
	jspl3 jspl3_w_n410_1(.douta(w_n410_1[0]),.doutb(w_n410_1[1]),.doutc(w_n410_1[2]),.din(w_n410_0[0]));
	jspl3 jspl3_w_n410_2(.douta(w_n410_2[0]),.doutb(w_n410_2[1]),.doutc(w_n410_2[2]),.din(w_n410_0[1]));
	jspl3 jspl3_w_n410_3(.douta(w_n410_3[0]),.doutb(w_n410_3[1]),.doutc(w_n410_3[2]),.din(w_n410_0[2]));
	jspl3 jspl3_w_n410_4(.douta(w_n410_4[0]),.doutb(w_n410_4[1]),.doutc(w_n410_4[2]),.din(w_n410_1[0]));
	jspl3 jspl3_w_n410_5(.douta(w_n410_5[0]),.doutb(w_n410_5[1]),.doutc(w_n410_5[2]),.din(w_n410_1[1]));
	jspl3 jspl3_w_n410_6(.douta(w_n410_6[0]),.doutb(w_n410_6[1]),.doutc(w_n410_6[2]),.din(w_n410_1[2]));
	jspl3 jspl3_w_n410_7(.douta(w_n410_7[0]),.doutb(w_n410_7[1]),.doutc(w_n410_7[2]),.din(w_n410_2[0]));
	jspl3 jspl3_w_n410_8(.douta(w_n410_8[0]),.doutb(w_n410_8[1]),.doutc(w_n410_8[2]),.din(w_n410_2[1]));
	jspl3 jspl3_w_n410_9(.douta(w_n410_9[0]),.doutb(w_n410_9[1]),.doutc(w_n410_9[2]),.din(w_n410_2[2]));
	jspl3 jspl3_w_n410_10(.douta(w_n410_10[0]),.doutb(w_n410_10[1]),.doutc(w_n410_10[2]),.din(w_n410_3[0]));
	jspl3 jspl3_w_n410_11(.douta(w_n410_11[0]),.doutb(w_n410_11[1]),.doutc(w_n410_11[2]),.din(w_n410_3[1]));
	jspl3 jspl3_w_n410_12(.douta(w_n410_12[0]),.doutb(w_n410_12[1]),.doutc(w_n410_12[2]),.din(w_n410_3[2]));
	jspl3 jspl3_w_n410_13(.douta(w_n410_13[0]),.doutb(w_n410_13[1]),.doutc(w_n410_13[2]),.din(w_n410_4[0]));
	jspl3 jspl3_w_n410_14(.douta(w_n410_14[0]),.doutb(w_n410_14[1]),.doutc(w_n410_14[2]),.din(w_n410_4[1]));
	jspl3 jspl3_w_n410_15(.douta(w_n410_15[0]),.doutb(w_n410_15[1]),.doutc(w_n410_15[2]),.din(w_n410_4[2]));
	jspl3 jspl3_w_n410_16(.douta(w_n410_16[0]),.doutb(w_n410_16[1]),.doutc(w_n410_16[2]),.din(w_n410_5[0]));
	jspl3 jspl3_w_n410_17(.douta(w_n410_17[0]),.doutb(w_n410_17[1]),.doutc(w_n410_17[2]),.din(w_n410_5[1]));
	jspl3 jspl3_w_n410_18(.douta(w_n410_18[0]),.doutb(w_n410_18[1]),.doutc(w_n410_18[2]),.din(w_n410_5[2]));
	jspl3 jspl3_w_n410_19(.douta(w_n410_19[0]),.doutb(w_n410_19[1]),.doutc(w_n410_19[2]),.din(w_n410_6[0]));
	jspl3 jspl3_w_n410_20(.douta(w_n410_20[0]),.doutb(w_n410_20[1]),.doutc(w_n410_20[2]),.din(w_n410_6[1]));
	jspl3 jspl3_w_n410_21(.douta(w_n410_21[0]),.doutb(w_n410_21[1]),.doutc(w_n410_21[2]),.din(w_n410_6[2]));
	jspl3 jspl3_w_n410_22(.douta(w_n410_22[0]),.doutb(w_n410_22[1]),.doutc(w_n410_22[2]),.din(w_n410_7[0]));
	jspl3 jspl3_w_n410_23(.douta(w_n410_23[0]),.doutb(w_n410_23[1]),.doutc(w_n410_23[2]),.din(w_n410_7[1]));
	jspl3 jspl3_w_n410_24(.douta(w_n410_24[0]),.doutb(w_n410_24[1]),.doutc(w_n410_24[2]),.din(w_n410_7[2]));
	jspl3 jspl3_w_n410_25(.douta(w_n410_25[0]),.doutb(w_n410_25[1]),.doutc(w_n410_25[2]),.din(w_n410_8[0]));
	jspl3 jspl3_w_n410_26(.douta(w_n410_26[0]),.doutb(w_n410_26[1]),.doutc(w_n410_26[2]),.din(w_n410_8[1]));
	jspl3 jspl3_w_n410_27(.douta(w_n410_27[0]),.doutb(w_n410_27[1]),.doutc(w_n410_27[2]),.din(w_n410_8[2]));
	jspl3 jspl3_w_n410_28(.douta(w_n410_28[0]),.doutb(w_n410_28[1]),.doutc(w_n410_28[2]),.din(w_n410_9[0]));
	jspl3 jspl3_w_n410_29(.douta(w_n410_29[0]),.doutb(w_n410_29[1]),.doutc(w_n410_29[2]),.din(w_n410_9[1]));
	jspl3 jspl3_w_n410_30(.douta(w_n410_30[0]),.doutb(w_n410_30[1]),.doutc(w_n410_30[2]),.din(w_n410_9[2]));
	jspl3 jspl3_w_n410_31(.douta(w_n410_31[0]),.doutb(w_n410_31[1]),.doutc(w_n410_31[2]),.din(w_n410_10[0]));
	jspl3 jspl3_w_n410_32(.douta(w_n410_32[0]),.doutb(w_n410_32[1]),.doutc(w_n410_32[2]),.din(w_n410_10[1]));
	jspl3 jspl3_w_n410_33(.douta(w_n410_33[0]),.doutb(w_n410_33[1]),.doutc(w_n410_33[2]),.din(w_n410_10[2]));
	jspl3 jspl3_w_n410_34(.douta(w_n410_34[0]),.doutb(w_n410_34[1]),.doutc(w_n410_34[2]),.din(w_n410_11[0]));
	jspl3 jspl3_w_n410_35(.douta(w_n410_35[0]),.doutb(w_n410_35[1]),.doutc(w_n410_35[2]),.din(w_n410_11[1]));
	jspl3 jspl3_w_n410_36(.douta(w_n410_36[0]),.doutb(w_n410_36[1]),.doutc(w_n410_36[2]),.din(w_n410_11[2]));
	jspl3 jspl3_w_n410_37(.douta(w_n410_37[0]),.doutb(w_n410_37[1]),.doutc(w_n410_37[2]),.din(w_n410_12[0]));
	jspl3 jspl3_w_n410_38(.douta(w_n410_38[0]),.doutb(w_n410_38[1]),.doutc(w_n410_38[2]),.din(w_n410_12[1]));
	jspl3 jspl3_w_n410_39(.douta(w_n410_39[0]),.doutb(w_n410_39[1]),.doutc(w_n410_39[2]),.din(w_n410_12[2]));
	jspl3 jspl3_w_n410_40(.douta(w_n410_40[0]),.doutb(w_n410_40[1]),.doutc(w_n410_40[2]),.din(w_n410_13[0]));
	jspl3 jspl3_w_n410_41(.douta(w_n410_41[0]),.doutb(w_n410_41[1]),.doutc(w_n410_41[2]),.din(w_n410_13[1]));
	jspl3 jspl3_w_n410_42(.douta(w_n410_42[0]),.doutb(w_n410_42[1]),.doutc(w_n410_42[2]),.din(w_n410_13[2]));
	jspl3 jspl3_w_n410_43(.douta(w_n410_43[0]),.doutb(w_n410_43[1]),.doutc(w_n410_43[2]),.din(w_n410_14[0]));
	jspl3 jspl3_w_n410_44(.douta(w_n410_44[0]),.doutb(w_n410_44[1]),.doutc(w_n410_44[2]),.din(w_n410_14[1]));
	jspl3 jspl3_w_n410_45(.douta(w_n410_45[0]),.doutb(w_n410_45[1]),.doutc(w_n410_45[2]),.din(w_n410_14[2]));
	jspl3 jspl3_w_n410_46(.douta(w_n410_46[0]),.doutb(w_n410_46[1]),.doutc(w_n410_46[2]),.din(w_n410_15[0]));
	jspl3 jspl3_w_n410_47(.douta(w_n410_47[0]),.doutb(w_n410_47[1]),.doutc(w_n410_47[2]),.din(w_n410_15[1]));
	jspl3 jspl3_w_n410_48(.douta(w_n410_48[0]),.doutb(w_n410_48[1]),.doutc(w_n410_48[2]),.din(w_n410_15[2]));
	jspl3 jspl3_w_n410_49(.douta(w_n410_49[0]),.doutb(w_n410_49[1]),.doutc(w_n410_49[2]),.din(w_n410_16[0]));
	jspl3 jspl3_w_n410_50(.douta(w_n410_50[0]),.doutb(w_n410_50[1]),.doutc(w_n410_50[2]),.din(w_n410_16[1]));
	jspl3 jspl3_w_n410_51(.douta(w_n410_51[0]),.doutb(w_n410_51[1]),.doutc(w_n410_51[2]),.din(w_n410_16[2]));
	jspl3 jspl3_w_n410_52(.douta(w_n410_52[0]),.doutb(w_n410_52[1]),.doutc(w_n410_52[2]),.din(w_n410_17[0]));
	jspl3 jspl3_w_n410_53(.douta(w_n410_53[0]),.doutb(w_n410_53[1]),.doutc(w_n410_53[2]),.din(w_n410_17[1]));
	jspl3 jspl3_w_n410_54(.douta(w_n410_54[0]),.doutb(w_n410_54[1]),.doutc(w_n410_54[2]),.din(w_n410_17[2]));
	jspl3 jspl3_w_n410_55(.douta(w_n410_55[0]),.doutb(w_n410_55[1]),.doutc(w_n410_55[2]),.din(w_n410_18[0]));
	jspl3 jspl3_w_n410_56(.douta(w_n410_56[0]),.doutb(w_n410_56[1]),.doutc(w_n410_56[2]),.din(w_n410_18[1]));
	jspl3 jspl3_w_n410_57(.douta(w_n410_57[0]),.doutb(w_n410_57[1]),.doutc(w_n410_57[2]),.din(w_n410_18[2]));
	jspl3 jspl3_w_n410_58(.douta(w_n410_58[0]),.doutb(w_n410_58[1]),.doutc(w_n410_58[2]),.din(w_n410_19[0]));
	jspl3 jspl3_w_n410_59(.douta(w_n410_59[0]),.doutb(w_n410_59[1]),.doutc(w_n410_59[2]),.din(w_n410_19[1]));
	jspl3 jspl3_w_n410_60(.douta(w_n410_60[0]),.doutb(w_n410_60[1]),.doutc(w_n410_60[2]),.din(w_n410_19[2]));
	jspl3 jspl3_w_n410_61(.douta(w_n410_61[0]),.doutb(w_n410_61[1]),.doutc(w_n410_61[2]),.din(w_n410_20[0]));
	jspl3 jspl3_w_n410_62(.douta(w_n410_62[0]),.doutb(w_n410_62[1]),.doutc(w_n410_62[2]),.din(w_n410_20[1]));
	jspl jspl_w_n410_63(.douta(w_n410_63[0]),.doutb(w_n410_63[1]),.din(w_n410_20[2]));
	jspl jspl_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.din(n413));
	jspl jspl_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.din(n417));
	jspl3 jspl3_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.doutc(w_n419_0[2]),.din(n419));
	jspl jspl_w_n419_1(.douta(w_n419_1[0]),.doutb(w_n419_1[1]),.din(w_n419_0[0]));
	jspl jspl_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.din(n423));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(n427));
	jspl3 jspl3_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.doutc(w_n429_0[2]),.din(n429));
	jspl jspl_w_n429_1(.douta(w_n429_1[0]),.doutb(w_n429_1[1]),.din(w_n429_0[0]));
	jspl jspl_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.din(n433));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.doutc(w_n439_0[2]),.din(n439));
	jspl jspl_w_n439_1(.douta(w_n439_1[0]),.doutb(w_n439_1[1]),.din(w_n439_0[0]));
	jspl jspl_w_n444_0(.douta(w_n444_0[0]),.doutb(w_n444_0[1]),.din(n444));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.din(n448));
	jspl3 jspl3_w_n450_0(.douta(w_n450_0[0]),.doutb(w_n450_0[1]),.doutc(w_n450_0[2]),.din(n450));
	jspl jspl_w_n450_1(.douta(w_n450_1[0]),.doutb(w_n450_1[1]),.din(w_n450_0[0]));
	jspl3 jspl3_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.doutc(w_n453_0[2]),.din(n453));
	jspl jspl_w_n453_1(.douta(w_n453_1[0]),.doutb(w_n453_1[1]),.din(w_n453_0[0]));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.din(n460));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(n464));
	jspl3 jspl3_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.doutc(w_n466_0[2]),.din(n466));
	jspl jspl_w_n466_1(.douta(w_n466_1[0]),.doutb(w_n466_1[1]),.din(w_n466_0[0]));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(n474));
	jspl3 jspl3_w_n476_0(.douta(w_n476_0[0]),.doutb(w_n476_0[1]),.doutc(w_n476_0[2]),.din(n476));
	jspl jspl_w_n476_1(.douta(w_n476_1[0]),.doutb(w_n476_1[1]),.din(w_n476_0[0]));
	jspl jspl_w_n480_0(.douta(w_n480_0[0]),.doutb(w_n480_0[1]),.din(n480));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl3 jspl3_w_n486_0(.douta(w_n486_0[0]),.doutb(w_n486_0[1]),.doutc(w_n486_0[2]),.din(n486));
	jspl jspl_w_n486_1(.douta(w_n486_1[0]),.doutb(w_n486_1[1]),.din(w_n486_0[0]));
	jspl jspl_w_n491_0(.douta(w_n491_0[0]),.doutb(w_n491_0[1]),.din(n491));
	jspl jspl_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.din(n495));
	jspl3 jspl3_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.doutc(w_n497_0[2]),.din(n497));
	jspl jspl_w_n497_1(.douta(w_n497_1[0]),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl3 jspl3_w_n500_0(.douta(w_n500_0[0]),.doutb(w_n500_0[1]),.doutc(w_n500_0[2]),.din(n500));
	jspl jspl_w_n500_1(.douta(w_n500_1[0]),.doutb(w_n500_1[1]),.din(w_n500_0[0]));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl3 jspl3_w_n510_0(.douta(w_n510_0[0]),.doutb(w_n510_0[1]),.doutc(w_n510_0[2]),.din(n510));
	jspl jspl_w_n510_1(.douta(w_n510_1[0]),.doutb(w_n510_1[1]),.din(w_n510_0[0]));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl3 jspl3_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.doutc(w_n520_0[2]),.din(n520));
	jspl jspl_w_n520_1(.douta(w_n520_1[0]),.doutb(w_n520_1[1]),.din(w_n520_0[0]));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl jspl_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.din(w_n530_0[0]));
	jspl jspl_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.din(n535));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl3 jspl3_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.doutc(w_n541_0[2]),.din(n541));
	jspl jspl_w_n541_1(.douta(w_n541_1[0]),.doutb(w_n541_1[1]),.din(w_n541_0[0]));
	jspl3 jspl3_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.doutc(w_n544_0[2]),.din(n544));
	jspl jspl_w_n544_1(.douta(w_n544_1[0]),.doutb(w_n544_1[1]),.din(w_n544_0[0]));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(n552));
	jspl3 jspl3_w_n554_0(.douta(w_n554_0[0]),.doutb(w_n554_0[1]),.doutc(w_n554_0[2]),.din(n554));
	jspl jspl_w_n554_1(.douta(w_n554_1[0]),.doutb(w_n554_1[1]),.din(w_n554_0[0]));
	jspl jspl_w_n558_0(.douta(w_n558_0[0]),.doutb(w_n558_0[1]),.din(n558));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n564_0(.douta(w_n564_0[0]),.doutb(w_n564_0[1]),.doutc(w_n564_0[2]),.din(n564));
	jspl jspl_w_n564_1(.douta(w_n564_1[0]),.doutb(w_n564_1[1]),.din(w_n564_0[0]));
	jspl jspl_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.din(n568));
	jspl jspl_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.din(n572));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl jspl_w_n574_1(.douta(w_n574_1[0]),.doutb(w_n574_1[1]),.din(w_n574_0[0]));
	jspl jspl_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.din(n579));
	jspl jspl_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.din(n583));
	jspl3 jspl3_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.doutc(w_n585_0[2]),.din(n585));
	jspl jspl_w_n585_1(.douta(w_n585_1[0]),.doutb(w_n585_1[1]),.din(w_n585_0[0]));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl3 jspl3_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.doutc(w_n599_0[2]),.din(n599));
	jspl jspl_w_n599_1(.douta(w_n599_1[0]),.doutb(w_n599_1[1]),.din(w_n599_0[0]));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.doutc(w_n609_0[2]),.din(n609));
	jspl jspl_w_n609_1(.douta(w_n609_1[0]),.doutb(w_n609_1[1]),.din(w_n609_0[0]));
	jspl jspl_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.din(n613));
	jspl jspl_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.din(n617));
	jspl3 jspl3_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.doutc(w_n619_0[2]),.din(n619));
	jspl jspl_w_n619_1(.douta(w_n619_1[0]),.doutb(w_n619_1[1]),.din(w_n619_0[0]));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(n628));
	jspl3 jspl3_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.doutc(w_n630_0[2]),.din(n630));
	jspl jspl_w_n630_1(.douta(w_n630_1[0]),.doutb(w_n630_1[1]),.din(w_n630_0[0]));
	jspl3 jspl3_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.doutc(w_n633_0[2]),.din(n633));
	jspl jspl_w_n633_1(.douta(w_n633_1[0]),.doutb(w_n633_1[1]),.din(w_n633_0[0]));
	jspl jspl_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.din(n636));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl3 jspl3_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.doutc(w_n647_0[2]),.din(n647));
	jspl jspl_w_n647_1(.douta(w_n647_1[0]),.doutb(w_n647_1[1]),.din(w_n647_0[0]));
	jspl jspl_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.din(n651));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl3 jspl3_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.doutc(w_n657_0[2]),.din(n657));
	jspl jspl_w_n657_1(.douta(w_n657_1[0]),.doutb(w_n657_1[1]),.din(w_n657_0[0]));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl jspl_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.din(n665));
	jspl3 jspl3_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.doutc(w_n667_0[2]),.din(n667));
	jspl jspl_w_n667_1(.douta(w_n667_1[0]),.doutb(w_n667_1[1]),.din(w_n667_0[0]));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl3 jspl3_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.doutc(w_n678_0[2]),.din(n678));
	jspl jspl_w_n678_1(.douta(w_n678_1[0]),.doutb(w_n678_1[1]),.din(w_n678_0[0]));
	jspl3 jspl3_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.doutc(w_n681_0[2]),.din(n681));
	jspl jspl_w_n681_1(.douta(w_n681_1[0]),.doutb(w_n681_1[1]),.din(w_n681_0[0]));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl3 jspl3_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.doutc(w_n691_0[2]),.din(n691));
	jspl jspl_w_n691_1(.douta(w_n691_1[0]),.doutb(w_n691_1[1]),.din(w_n691_0[0]));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl3 jspl3_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.doutc(w_n701_0[2]),.din(n701));
	jspl jspl_w_n701_1(.douta(w_n701_1[0]),.doutb(w_n701_1[1]),.din(w_n701_0[0]));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(n709));
	jspl3 jspl3_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.doutc(w_n711_0[2]),.din(n711));
	jspl jspl_w_n711_1(.douta(w_n711_1[0]),.doutb(w_n711_1[1]),.din(w_n711_0[0]));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl3 jspl3_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.doutc(w_n722_0[2]),.din(n722));
	jspl jspl_w_n722_1(.douta(w_n722_1[0]),.doutb(w_n722_1[1]),.din(w_n722_0[0]));
	jspl3 jspl3_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.doutc(w_n725_0[2]),.din(n725));
	jspl jspl_w_n725_1(.douta(w_n725_1[0]),.doutb(w_n725_1[1]),.din(w_n725_0[0]));
	jspl jspl_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.din(n729));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl3 jspl3_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.doutc(w_n735_0[2]),.din(n735));
	jspl jspl_w_n735_1(.douta(w_n735_1[0]),.doutb(w_n735_1[1]),.din(w_n735_0[0]));
	jspl jspl_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.din(n739));
	jspl jspl_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.din(n743));
	jspl3 jspl3_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.doutc(w_n745_0[2]),.din(n745));
	jspl jspl_w_n745_1(.douta(w_n745_1[0]),.doutb(w_n745_1[1]),.din(w_n745_0[0]));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(n749));
	jspl jspl_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.din(n753));
	jspl3 jspl3_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.doutc(w_n755_0[2]),.din(n755));
	jspl jspl_w_n755_1(.douta(w_n755_1[0]),.doutb(w_n755_1[1]),.din(w_n755_0[0]));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(n764));
	jspl3 jspl3_w_n766_0(.douta(w_n766_0[0]),.doutb(w_n766_0[1]),.doutc(w_n766_0[2]),.din(n766));
	jspl jspl_w_n766_1(.douta(w_n766_1[0]),.doutb(w_n766_1[1]),.din(w_n766_0[0]));
	jspl3 jspl3_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.doutc(w_n769_0[2]),.din(n769));
	jspl jspl_w_n769_1(.douta(w_n769_1[0]),.doutb(w_n769_1[1]),.din(w_n769_0[0]));
	jspl jspl_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.din(n774));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl3 jspl3_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.doutc(w_n780_0[2]),.din(n780));
	jspl jspl_w_n780_1(.douta(w_n780_1[0]),.doutb(w_n780_1[1]),.din(w_n780_0[0]));
	jspl jspl_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.din(n784));
	jspl jspl_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.din(n788));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.doutc(w_n790_0[2]),.din(n790));
	jspl jspl_w_n790_1(.douta(w_n790_1[0]),.doutb(w_n790_1[1]),.din(w_n790_0[0]));
	jspl jspl_w_n794_0(.douta(w_n794_0[0]),.doutb(w_n794_0[1]),.din(n794));
	jspl jspl_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.din(n798));
	jspl3 jspl3_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.doutc(w_n800_0[2]),.din(n800));
	jspl jspl_w_n800_1(.douta(w_n800_1[0]),.doutb(w_n800_1[1]),.din(w_n800_0[0]));
	jspl jspl_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl3 jspl3_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.doutc(w_n811_0[2]),.din(n811));
	jspl jspl_w_n811_1(.douta(w_n811_1[0]),.doutb(w_n811_1[1]),.din(w_n811_0[0]));
	jspl3 jspl3_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.doutc(w_n814_0[2]),.din(n814));
	jspl jspl_w_n814_1(.douta(w_n814_1[0]),.doutb(w_n814_1[1]),.din(w_n814_0[0]));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(n817));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(n821));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl3 jspl3_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.doutc(w_n827_0[2]),.din(n827));
	jspl jspl_w_n827_1(.douta(w_n827_1[0]),.doutb(w_n827_1[1]),.din(w_n827_0[0]));
	jspl jspl_w_n831_0(.douta(w_n831_0[0]),.doutb(w_n831_0[1]),.din(n831));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl3 jspl3_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.doutc(w_n837_0[2]),.din(n837));
	jspl jspl_w_n837_1(.douta(w_n837_1[0]),.doutb(w_n837_1[1]),.din(w_n837_0[0]));
	jspl jspl_w_n841_0(.douta(w_n841_0[0]),.doutb(w_n841_0[1]),.din(n841));
	jspl jspl_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.din(n845));
	jspl3 jspl3_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.doutc(w_n847_0[2]),.din(n847));
	jspl jspl_w_n847_1(.douta(w_n847_1[0]),.doutb(w_n847_1[1]),.din(w_n847_0[0]));
	jspl jspl_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.din(n852));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl3 jspl3_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.doutc(w_n858_0[2]),.din(n858));
	jspl jspl_w_n858_1(.douta(w_n858_1[0]),.doutb(w_n858_1[1]),.din(w_n858_0[0]));
	jspl3 jspl3_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.doutc(w_n861_0[2]),.din(n861));
	jspl jspl_w_n861_1(.douta(w_n861_1[0]),.doutb(w_n861_1[1]),.din(w_n861_0[0]));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.din(n865));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl3 jspl3_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.doutc(w_n871_0[2]),.din(n871));
	jspl jspl_w_n871_1(.douta(w_n871_1[0]),.doutb(w_n871_1[1]),.din(w_n871_0[0]));
	jspl jspl_w_n875_0(.douta(w_n875_0[0]),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl3 jspl3_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.doutc(w_n881_0[2]),.din(n881));
	jspl jspl_w_n881_1(.douta(w_n881_1[0]),.doutb(w_n881_1[1]),.din(w_n881_0[0]));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl3 jspl3_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.doutc(w_n891_0[2]),.din(n891));
	jspl jspl_w_n891_1(.douta(w_n891_1[0]),.doutb(w_n891_1[1]),.din(w_n891_0[0]));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(n896));
	jspl jspl_w_n900_0(.douta(w_n900_0[0]),.doutb(w_n900_0[1]),.din(n900));
	jspl3 jspl3_w_n902_0(.douta(w_n902_0[0]),.doutb(w_n902_0[1]),.doutc(w_n902_0[2]),.din(n902));
	jspl jspl_w_n902_1(.douta(w_n902_1[0]),.doutb(w_n902_1[1]),.din(w_n902_0[0]));
	jspl3 jspl3_w_n905_0(.douta(w_n905_0[0]),.doutb(w_n905_0[1]),.doutc(w_n905_0[2]),.din(n905));
	jspl jspl_w_n905_1(.douta(w_n905_1[0]),.doutb(w_n905_1[1]),.din(w_n905_0[0]));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(n913));
	jspl3 jspl3_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.doutc(w_n915_0[2]),.din(n915));
	jspl jspl_w_n915_1(.douta(w_n915_1[0]),.doutb(w_n915_1[1]),.din(w_n915_0[0]));
	jspl jspl_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.din(n919));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(n923));
	jspl3 jspl3_w_n925_0(.douta(w_n925_0[0]),.doutb(w_n925_0[1]),.doutc(w_n925_0[2]),.din(n925));
	jspl jspl_w_n925_1(.douta(w_n925_1[0]),.doutb(w_n925_1[1]),.din(w_n925_0[0]));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(n929));
	jspl jspl_w_n933_0(.douta(w_n933_0[0]),.doutb(w_n933_0[1]),.din(n933));
	jspl3 jspl3_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.doutc(w_n935_0[2]),.din(n935));
	jspl jspl_w_n935_1(.douta(w_n935_1[0]),.doutb(w_n935_1[1]),.din(w_n935_0[0]));
	jspl jspl_w_n940_0(.douta(w_n940_0[0]),.doutb(w_n940_0[1]),.din(n940));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(n944));
	jspl3 jspl3_w_n946_0(.douta(w_n946_0[0]),.doutb(w_n946_0[1]),.doutc(w_n946_0[2]),.din(n946));
	jspl jspl_w_n946_1(.douta(w_n946_1[0]),.doutb(w_n946_1[1]),.din(w_n946_0[0]));
	jspl3 jspl3_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.doutc(w_n949_0[2]),.din(n949));
	jspl jspl_w_n949_1(.douta(w_n949_1[0]),.doutb(w_n949_1[1]),.din(w_n949_0[0]));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n958_0(.douta(w_n958_0[0]),.doutb(w_n958_0[1]),.din(n958));
	jspl3 jspl3_w_n960_0(.douta(w_n960_0[0]),.doutb(w_n960_0[1]),.doutc(w_n960_0[2]),.din(n960));
	jspl jspl_w_n960_1(.douta(w_n960_1[0]),.doutb(w_n960_1[1]),.din(w_n960_0[0]));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n968_0(.douta(w_n968_0[0]),.doutb(w_n968_0[1]),.din(n968));
	jspl3 jspl3_w_n970_0(.douta(w_n970_0[0]),.doutb(w_n970_0[1]),.doutc(w_n970_0[2]),.din(n970));
	jspl jspl_w_n970_1(.douta(w_n970_1[0]),.doutb(w_n970_1[1]),.din(w_n970_0[0]));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n978_0(.douta(w_n978_0[0]),.doutb(w_n978_0[1]),.din(n978));
	jspl3 jspl3_w_n980_0(.douta(w_n980_0[0]),.doutb(w_n980_0[1]),.doutc(w_n980_0[2]),.din(n980));
	jspl jspl_w_n980_1(.douta(w_n980_1[0]),.doutb(w_n980_1[1]),.din(w_n980_0[0]));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl3 jspl3_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.doutc(w_n991_0[2]),.din(n991));
	jspl jspl_w_n991_1(.douta(w_n991_1[0]),.doutb(w_n991_1[1]),.din(w_n991_0[0]));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl jspl_w_n994_1(.douta(w_n994_1[0]),.doutb(w_n994_1[1]),.din(w_n994_0[0]));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.doutc(w_n1002_0[2]),.din(n1002));
	jspl jspl_w_n1002_1(.douta(w_n1002_1[0]),.doutb(w_n1002_1[1]),.din(w_n1002_0[0]));
	jspl3 jspl3_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.doutc(w_n1006_0[2]),.din(n1006));
	jspl jspl_w_n1006_1(.douta(w_n1006_1[0]),.doutb(w_n1006_1[1]),.din(w_n1006_0[0]));
	jspl3 jspl3_w_n1010_0(.douta(w_n1010_0[0]),.doutb(w_n1010_0[1]),.doutc(w_n1010_0[2]),.din(n1010));
	jspl jspl_w_n1010_1(.douta(w_n1010_1[0]),.doutb(w_n1010_1[1]),.din(w_n1010_0[0]));
	jspl3 jspl3_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.doutc(w_n1015_0[2]),.din(n1015));
	jspl jspl_w_n1015_1(.douta(w_n1015_1[0]),.doutb(w_n1015_1[1]),.din(w_n1015_0[0]));
	jspl3 jspl3_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.doutc(w_n1018_0[2]),.din(n1018));
	jspl jspl_w_n1018_1(.douta(w_n1018_1[0]),.doutb(w_n1018_1[1]),.din(w_n1018_0[0]));
	jspl3 jspl3_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.doutc(w_n1022_0[2]),.din(n1022));
	jspl jspl_w_n1022_1(.douta(w_n1022_1[0]),.doutb(w_n1022_1[1]),.din(w_n1022_0[0]));
	jspl3 jspl3_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.doutc(w_n1026_0[2]),.din(n1026));
	jspl jspl_w_n1026_1(.douta(w_n1026_1[0]),.doutb(w_n1026_1[1]),.din(w_n1026_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.doutc(w_n1035_0[2]),.din(n1035));
	jspl jspl_w_n1035_1(.douta(w_n1035_1[0]),.doutb(w_n1035_1[1]),.din(w_n1035_0[0]));
	jspl3 jspl3_w_n1038_0(.douta(w_n1038_0[0]),.doutb(w_n1038_0[1]),.doutc(w_n1038_0[2]),.din(n1038));
	jspl jspl_w_n1038_1(.douta(w_n1038_1[0]),.doutb(w_n1038_1[1]),.din(w_n1038_0[0]));
	jspl3 jspl3_w_n1042_0(.douta(w_n1042_0[0]),.doutb(w_n1042_0[1]),.doutc(w_n1042_0[2]),.din(n1042));
	jspl jspl_w_n1042_1(.douta(w_n1042_1[0]),.doutb(w_n1042_1[1]),.din(w_n1042_0[0]));
	jspl3 jspl3_w_n1046_0(.douta(w_n1046_0[0]),.doutb(w_n1046_0[1]),.doutc(w_n1046_0[2]),.din(n1046));
	jspl jspl_w_n1046_1(.douta(w_n1046_1[0]),.doutb(w_n1046_1[1]),.din(w_n1046_0[0]));
	jspl3 jspl3_w_n1050_0(.douta(w_n1050_0[0]),.doutb(w_n1050_0[1]),.doutc(w_n1050_0[2]),.din(n1050));
	jspl jspl_w_n1050_1(.douta(w_n1050_1[0]),.doutb(w_n1050_1[1]),.din(w_n1050_0[0]));
	jspl3 jspl3_w_n1055_0(.douta(w_n1055_0[0]),.doutb(w_n1055_0[1]),.doutc(w_n1055_0[2]),.din(n1055));
	jspl jspl_w_n1055_1(.douta(w_n1055_1[0]),.doutb(w_n1055_1[1]),.din(w_n1055_0[0]));
	jspl3 jspl3_w_n1058_0(.douta(w_n1058_0[0]),.doutb(w_n1058_0[1]),.doutc(w_n1058_0[2]),.din(n1058));
	jspl jspl_w_n1058_1(.douta(w_n1058_1[0]),.doutb(w_n1058_1[1]),.din(w_n1058_0[0]));
	jspl3 jspl3_w_n1063_0(.douta(w_n1063_0[0]),.doutb(w_n1063_0[1]),.doutc(w_n1063_0[2]),.din(n1063));
	jspl jspl_w_n1063_1(.douta(w_n1063_1[0]),.doutb(w_n1063_1[1]),.din(w_n1063_0[0]));
	jspl3 jspl3_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.doutc(w_n1067_0[2]),.din(n1067));
	jspl jspl_w_n1067_1(.douta(w_n1067_1[0]),.doutb(w_n1067_1[1]),.din(w_n1067_0[0]));
	jspl3 jspl3_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.doutc(w_n1071_0[2]),.din(n1071));
	jspl jspl_w_n1071_1(.douta(w_n1071_1[0]),.doutb(w_n1071_1[1]),.din(w_n1071_0[0]));
	jspl3 jspl3_w_n1076_0(.douta(w_n1076_0[0]),.doutb(w_n1076_0[1]),.doutc(w_n1076_0[2]),.din(n1076));
	jspl jspl_w_n1076_1(.douta(w_n1076_1[0]),.doutb(w_n1076_1[1]),.din(w_n1076_0[0]));
	jspl3 jspl3_w_n1079_0(.douta(w_n1079_0[0]),.doutb(w_n1079_0[1]),.doutc(w_n1079_0[2]),.din(n1079));
	jspl jspl_w_n1079_1(.douta(w_n1079_1[0]),.doutb(w_n1079_1[1]),.din(w_n1079_0[0]));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl3 jspl3_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.doutc(w_n1086_0[2]),.din(n1086));
	jspl jspl_w_n1086_1(.douta(w_n1086_1[0]),.doutb(w_n1086_1[1]),.din(w_n1086_0[0]));
	jspl3 jspl3_w_n1090_0(.douta(w_n1090_0[0]),.doutb(w_n1090_0[1]),.doutc(w_n1090_0[2]),.din(n1090));
	jspl jspl_w_n1090_1(.douta(w_n1090_1[0]),.doutb(w_n1090_1[1]),.din(w_n1090_0[0]));
	jspl3 jspl3_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.doutc(w_n1094_0[2]),.din(n1094));
	jspl jspl_w_n1094_1(.douta(w_n1094_1[0]),.doutb(w_n1094_1[1]),.din(w_n1094_0[0]));
	jspl3 jspl3_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.doutc(w_n1099_0[2]),.din(n1099));
	jspl jspl_w_n1099_1(.douta(w_n1099_1[0]),.doutb(w_n1099_1[1]),.din(w_n1099_0[0]));
	jspl3 jspl3_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.doutc(w_n1102_0[2]),.din(n1102));
	jspl jspl_w_n1102_1(.douta(w_n1102_1[0]),.doutb(w_n1102_1[1]),.din(w_n1102_0[0]));
	jspl3 jspl3_w_n1106_0(.douta(w_n1106_0[0]),.doutb(w_n1106_0[1]),.doutc(w_n1106_0[2]),.din(n1106));
	jspl jspl_w_n1106_1(.douta(w_n1106_1[0]),.doutb(w_n1106_1[1]),.din(w_n1106_0[0]));
	jspl3 jspl3_w_n1110_0(.douta(w_n1110_0[0]),.doutb(w_n1110_0[1]),.doutc(w_n1110_0[2]),.din(n1110));
	jspl jspl_w_n1110_1(.douta(w_n1110_1[0]),.doutb(w_n1110_1[1]),.din(w_n1110_0[0]));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl jspl_w_n1114_1(.douta(w_n1114_1[0]),.doutb(w_n1114_1[1]),.din(w_n1114_0[0]));
	jspl3 jspl3_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.doutc(w_n1119_0[2]),.din(n1119));
	jspl jspl_w_n1119_1(.douta(w_n1119_1[0]),.doutb(w_n1119_1[1]),.din(w_n1119_0[0]));
	jspl3 jspl3_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.doutc(w_n1122_0[2]),.din(n1122));
	jspl jspl_w_n1122_1(.douta(w_n1122_1[0]),.doutb(w_n1122_1[1]),.din(w_n1122_0[0]));
	jspl3 jspl3_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.doutc(w_n1126_0[2]),.din(n1126));
	jspl jspl_w_n1126_1(.douta(w_n1126_1[0]),.doutb(w_n1126_1[1]),.din(w_n1126_0[0]));
	jspl3 jspl3_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.doutc(w_n1130_0[2]),.din(n1130));
	jspl jspl_w_n1130_1(.douta(w_n1130_1[0]),.doutb(w_n1130_1[1]),.din(w_n1130_0[0]));
	jspl3 jspl3_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.doutc(w_n1134_0[2]),.din(n1134));
	jspl jspl_w_n1134_1(.douta(w_n1134_1[0]),.doutb(w_n1134_1[1]),.din(w_n1134_0[0]));
	jspl3 jspl3_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.doutc(w_n1139_0[2]),.din(n1139));
	jspl jspl_w_n1139_1(.douta(w_n1139_1[0]),.doutb(w_n1139_1[1]),.din(w_n1139_0[0]));
	jspl3 jspl3_w_n1142_0(.douta(w_n1142_0[0]),.doutb(w_n1142_0[1]),.doutc(w_n1142_0[2]),.din(n1142));
	jspl jspl_w_n1142_1(.douta(w_n1142_1[0]),.doutb(w_n1142_1[1]),.din(w_n1142_0[0]));
	jspl3 jspl3_w_n1147_0(.douta(w_n1147_0[0]),.doutb(w_n1147_0[1]),.doutc(w_n1147_0[2]),.din(n1147));
	jspl jspl_w_n1147_1(.douta(w_n1147_1[0]),.doutb(w_n1147_1[1]),.din(w_n1147_0[0]));
	jspl3 jspl3_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.doutc(w_n1151_0[2]),.din(n1151));
	jspl jspl_w_n1151_1(.douta(w_n1151_1[0]),.doutb(w_n1151_1[1]),.din(w_n1151_0[0]));
	jspl3 jspl3_w_n1155_0(.douta(w_n1155_0[0]),.doutb(w_n1155_0[1]),.doutc(w_n1155_0[2]),.din(n1155));
	jspl jspl_w_n1155_1(.douta(w_n1155_1[0]),.doutb(w_n1155_1[1]),.din(w_n1155_0[0]));
	jspl3 jspl3_w_n1160_0(.douta(w_n1160_0[0]),.doutb(w_n1160_0[1]),.doutc(w_n1160_0[2]),.din(n1160));
	jspl jspl_w_n1160_1(.douta(w_n1160_1[0]),.doutb(w_n1160_1[1]),.din(w_n1160_0[0]));
	jspl3 jspl3_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.doutc(w_n1163_0[2]),.din(n1163));
	jspl jspl_w_n1163_1(.douta(w_n1163_1[0]),.doutb(w_n1163_1[1]),.din(w_n1163_0[0]));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl3 jspl3_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.doutc(w_n1171_0[2]),.din(n1171));
	jspl jspl_w_n1171_1(.douta(w_n1171_1[0]),.doutb(w_n1171_1[1]),.din(w_n1171_0[0]));
	jspl3 jspl3_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_n1175_0[1]),.doutc(w_n1175_0[2]),.din(n1175));
	jspl jspl_w_n1175_1(.douta(w_n1175_1[0]),.doutb(w_n1175_1[1]),.din(w_n1175_0[0]));
	jspl3 jspl3_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.doutc(w_n1179_0[2]),.din(n1179));
	jspl jspl_w_n1179_1(.douta(w_n1179_1[0]),.doutb(w_n1179_1[1]),.din(w_n1179_0[0]));
	jspl3 jspl3_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.doutc(w_n1184_0[2]),.din(n1184));
	jspl jspl_w_n1184_1(.douta(w_n1184_1[0]),.doutb(w_n1184_1[1]),.din(w_n1184_0[0]));
	jspl3 jspl3_w_n1187_0(.douta(w_n1187_0[0]),.doutb(w_n1187_0[1]),.doutc(w_n1187_0[2]),.din(n1187));
	jspl jspl_w_n1187_1(.douta(w_n1187_1[0]),.doutb(w_n1187_1[1]),.din(w_n1187_0[0]));
	jspl3 jspl3_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.doutc(w_n1191_0[2]),.din(n1191));
	jspl jspl_w_n1191_1(.douta(w_n1191_1[0]),.doutb(w_n1191_1[1]),.din(w_n1191_0[0]));
	jspl3 jspl3_w_n1195_0(.douta(w_n1195_0[0]),.doutb(w_n1195_0[1]),.doutc(w_n1195_0[2]),.din(n1195));
	jspl jspl_w_n1195_1(.douta(w_n1195_1[0]),.doutb(w_n1195_1[1]),.din(w_n1195_0[0]));
	jspl3 jspl3_w_n1199_0(.douta(w_n1199_0[0]),.doutb(w_n1199_0[1]),.doutc(w_n1199_0[2]),.din(n1199));
	jspl jspl_w_n1199_1(.douta(w_n1199_1[0]),.doutb(w_n1199_1[1]),.din(w_n1199_0[0]));
	jspl3 jspl3_w_n1204_0(.douta(w_n1204_0[0]),.doutb(w_n1204_0[1]),.doutc(w_n1204_0[2]),.din(n1204));
	jspl jspl_w_n1204_1(.douta(w_n1204_1[0]),.doutb(w_n1204_1[1]),.din(w_n1204_0[0]));
	jspl3 jspl3_w_n1207_0(.douta(w_n1207_0[0]),.doutb(w_n1207_0[1]),.doutc(w_n1207_0[2]),.din(n1207));
	jspl jspl_w_n1207_1(.douta(w_n1207_1[0]),.doutb(w_n1207_1[1]),.din(w_n1207_0[0]));
	jspl3 jspl3_w_n1211_0(.douta(w_n1211_0[0]),.doutb(w_n1211_0[1]),.doutc(w_n1211_0[2]),.din(n1211));
	jspl jspl_w_n1211_1(.douta(w_n1211_1[0]),.doutb(w_n1211_1[1]),.din(w_n1211_0[0]));
	jspl3 jspl3_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.doutc(w_n1215_0[2]),.din(n1215));
	jspl jspl_w_n1215_1(.douta(w_n1215_1[0]),.doutb(w_n1215_1[1]),.din(w_n1215_0[0]));
	jspl3 jspl3_w_n1219_0(.douta(w_n1219_0[0]),.doutb(w_n1219_0[1]),.doutc(w_n1219_0[2]),.din(n1219));
	jspl jspl_w_n1219_1(.douta(w_n1219_1[0]),.doutb(w_n1219_1[1]),.din(w_n1219_0[0]));
	jspl3 jspl3_w_n1224_0(.douta(w_n1224_0[0]),.doutb(w_n1224_0[1]),.doutc(w_n1224_0[2]),.din(n1224));
	jspl jspl_w_n1224_1(.douta(w_n1224_1[0]),.doutb(w_n1224_1[1]),.din(w_n1224_0[0]));
	jspl3 jspl3_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.doutc(w_n1227_0[2]),.din(n1227));
	jspl jspl_w_n1227_1(.douta(w_n1227_1[0]),.doutb(w_n1227_1[1]),.din(w_n1227_0[0]));
	jspl3 jspl3_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.doutc(w_n1232_0[2]),.din(n1232));
	jspl jspl_w_n1232_1(.douta(w_n1232_1[0]),.doutb(w_n1232_1[1]),.din(w_n1232_0[0]));
	jspl3 jspl3_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.doutc(w_n1236_0[2]),.din(n1236));
	jspl jspl_w_n1236_1(.douta(w_n1236_1[0]),.doutb(w_n1236_1[1]),.din(w_n1236_0[0]));
	jspl3 jspl3_w_n1240_0(.douta(w_n1240_0[0]),.doutb(w_n1240_0[1]),.doutc(w_n1240_0[2]),.din(n1240));
	jspl jspl_w_n1240_1(.douta(w_n1240_1[0]),.doutb(w_n1240_1[1]),.din(w_n1240_0[0]));
	jspl3 jspl3_w_n1245_0(.douta(w_n1245_0[0]),.doutb(w_n1245_0[1]),.doutc(w_n1245_0[2]),.din(n1245));
	jspl jspl_w_n1245_1(.douta(w_n1245_1[0]),.doutb(w_n1245_1[1]),.din(w_n1245_0[0]));
	jspl3 jspl3_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.doutc(w_n1248_0[2]),.din(n1248));
	jspl jspl_w_n1248_1(.douta(w_n1248_1[0]),.doutb(w_n1248_1[1]),.din(w_n1248_0[0]));
	jspl jspl_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.din(n1251));
	jspl3 jspl3_w_n1255_0(.douta(w_n1255_0[0]),.doutb(w_n1255_0[1]),.doutc(w_n1255_0[2]),.din(n1255));
	jspl jspl_w_n1255_1(.douta(w_n1255_1[0]),.doutb(w_n1255_1[1]),.din(w_n1255_0[0]));
	jspl3 jspl3_w_n1259_0(.douta(w_n1259_0[0]),.doutb(w_n1259_0[1]),.doutc(w_n1259_0[2]),.din(n1259));
	jspl jspl_w_n1259_1(.douta(w_n1259_1[0]),.doutb(w_n1259_1[1]),.din(w_n1259_0[0]));
	jspl3 jspl3_w_n1263_0(.douta(w_n1263_0[0]),.doutb(w_n1263_0[1]),.doutc(w_n1263_0[2]),.din(n1263));
	jspl jspl_w_n1263_1(.douta(w_n1263_1[0]),.doutb(w_n1263_1[1]),.din(w_n1263_0[0]));
	jspl3 jspl3_w_n1268_0(.douta(w_n1268_0[0]),.doutb(w_n1268_0[1]),.doutc(w_n1268_0[2]),.din(n1268));
	jspl jspl_w_n1268_1(.douta(w_n1268_1[0]),.doutb(w_n1268_1[1]),.din(w_n1268_0[0]));
	jspl3 jspl3_w_n1271_0(.douta(w_n1271_0[0]),.doutb(w_n1271_0[1]),.doutc(w_n1271_0[2]),.din(n1271));
	jspl jspl_w_n1271_1(.douta(w_n1271_1[0]),.doutb(w_n1271_1[1]),.din(w_n1271_0[0]));
	jspl3 jspl3_w_n1275_0(.douta(w_n1275_0[0]),.doutb(w_n1275_0[1]),.doutc(w_n1275_0[2]),.din(n1275));
	jspl jspl_w_n1275_1(.douta(w_n1275_1[0]),.doutb(w_n1275_1[1]),.din(w_n1275_0[0]));
	jspl3 jspl3_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.doutc(w_n1279_0[2]),.din(n1279));
	jspl jspl_w_n1279_1(.douta(w_n1279_1[0]),.doutb(w_n1279_1[1]),.din(w_n1279_0[0]));
	jspl3 jspl3_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.doutc(w_n1283_0[2]),.din(n1283));
	jspl jspl_w_n1283_1(.douta(w_n1283_1[0]),.doutb(w_n1283_1[1]),.din(w_n1283_0[0]));
	jspl3 jspl3_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.doutc(w_n1288_0[2]),.din(n1288));
	jspl jspl_w_n1288_1(.douta(w_n1288_1[0]),.doutb(w_n1288_1[1]),.din(w_n1288_0[0]));
	jspl3 jspl3_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_n1291_0[1]),.doutc(w_n1291_0[2]),.din(n1291));
	jspl jspl_w_n1291_1(.douta(w_n1291_1[0]),.doutb(w_n1291_1[1]),.din(w_n1291_0[0]));
	jspl3 jspl3_w_n1295_0(.douta(w_n1295_0[0]),.doutb(w_n1295_0[1]),.doutc(w_n1295_0[2]),.din(n1295));
	jspl jspl_w_n1295_1(.douta(w_n1295_1[0]),.doutb(w_n1295_1[1]),.din(w_n1295_0[0]));
	jspl3 jspl3_w_n1299_0(.douta(w_n1299_0[0]),.doutb(w_n1299_0[1]),.doutc(w_n1299_0[2]),.din(n1299));
	jspl jspl_w_n1299_1(.douta(w_n1299_1[0]),.doutb(w_n1299_1[1]),.din(w_n1299_0[0]));
	jspl3 jspl3_w_n1303_0(.douta(w_n1303_0[0]),.doutb(w_n1303_0[1]),.doutc(w_n1303_0[2]),.din(n1303));
	jspl jspl_w_n1303_1(.douta(w_n1303_1[0]),.doutb(w_n1303_1[1]),.din(w_n1303_0[0]));
	jspl3 jspl3_w_n1308_0(.douta(w_n1308_0[0]),.doutb(w_n1308_0[1]),.doutc(w_n1308_0[2]),.din(n1308));
	jspl jspl_w_n1308_1(.douta(w_n1308_1[0]),.doutb(w_n1308_1[1]),.din(w_n1308_0[0]));
	jspl3 jspl3_w_n1311_0(.douta(w_n1311_0[0]),.doutb(w_n1311_0[1]),.doutc(w_n1311_0[2]),.din(n1311));
	jspl jspl_w_n1311_1(.douta(w_n1311_1[0]),.doutb(w_n1311_1[1]),.din(w_n1311_0[0]));
	jspl3 jspl3_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.doutc(w_n1316_0[2]),.din(n1316));
	jspl jspl_w_n1316_1(.douta(w_n1316_1[0]),.doutb(w_n1316_1[1]),.din(w_n1316_0[0]));
	jspl3 jspl3_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.doutc(w_n1320_0[2]),.din(n1320));
	jspl jspl_w_n1320_1(.douta(w_n1320_1[0]),.doutb(w_n1320_1[1]),.din(w_n1320_0[0]));
	jspl3 jspl3_w_n1324_0(.douta(w_n1324_0[0]),.doutb(w_n1324_0[1]),.doutc(w_n1324_0[2]),.din(n1324));
	jspl jspl_w_n1324_1(.douta(w_n1324_1[0]),.doutb(w_n1324_1[1]),.din(w_n1324_0[0]));
	jspl3 jspl3_w_n1329_0(.douta(w_n1329_0[0]),.doutb(w_n1329_0[1]),.doutc(w_n1329_0[2]),.din(n1329));
	jspl jspl_w_n1329_1(.douta(w_n1329_1[0]),.doutb(w_n1329_1[1]),.din(w_n1329_0[0]));
	jspl3 jspl3_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.doutc(w_n1332_0[2]),.din(n1332));
	jspl jspl_w_n1332_1(.douta(w_n1332_1[0]),.doutb(w_n1332_1[1]),.din(w_n1332_0[0]));
	jspl jspl_w_n1335_0(.douta(w_n1335_0[0]),.doutb(w_n1335_0[1]),.din(n1335));
	jspl3 jspl3_w_n1344_0(.douta(w_n1344_0[0]),.doutb(w_n1344_0[1]),.doutc(w_n1344_0[2]),.din(n1344));
	jspl jspl_w_n1344_1(.douta(w_n1344_1[0]),.doutb(w_n1344_1[1]),.din(w_n1344_0[0]));
	jspl3 jspl3_w_n1352_0(.douta(w_n1352_0[0]),.doutb(w_n1352_0[1]),.doutc(w_n1352_0[2]),.din(n1352));
	jspl jspl_w_n1352_1(.douta(w_n1352_1[0]),.doutb(w_n1352_1[1]),.din(w_n1352_0[0]));
	jspl3 jspl3_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.doutc(w_n1360_0[2]),.din(n1360));
	jspl jspl_w_n1360_1(.douta(w_n1360_1[0]),.doutb(w_n1360_1[1]),.din(w_n1360_0[0]));
	jspl3 jspl3_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.doutc(w_n1369_0[2]),.din(n1369));
	jspl jspl_w_n1369_1(.douta(w_n1369_1[0]),.doutb(w_n1369_1[1]),.din(w_n1369_0[0]));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl3 jspl3_w_n1380_0(.douta(w_n1380_0[0]),.doutb(w_n1380_0[1]),.doutc(w_n1380_0[2]),.din(n1380));
	jspl jspl_w_n1380_1(.douta(w_n1380_1[0]),.doutb(w_n1380_1[1]),.din(w_n1380_0[0]));
	jspl3 jspl3_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_n1388_0[1]),.doutc(w_n1388_0[2]),.din(n1388));
	jspl jspl_w_n1388_1(.douta(w_n1388_1[0]),.doutb(w_n1388_1[1]),.din(w_n1388_0[0]));
	jspl3 jspl3_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.doutc(w_n1396_0[2]),.din(n1396));
	jspl jspl_w_n1396_1(.douta(w_n1396_1[0]),.doutb(w_n1396_1[1]),.din(w_n1396_0[0]));
	jspl3 jspl3_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.doutc(w_n1405_0[2]),.din(n1405));
	jspl jspl_w_n1405_1(.douta(w_n1405_1[0]),.doutb(w_n1405_1[1]),.din(w_n1405_0[0]));
	jspl jspl_w_n1408_0(.douta(w_n1408_0[0]),.doutb(w_n1408_0[1]),.din(n1408));
	jspl3 jspl3_w_n1417_0(.douta(w_n1417_0[0]),.doutb(w_n1417_0[1]),.doutc(w_n1417_0[2]),.din(n1417));
	jspl jspl_w_n1417_1(.douta(w_n1417_1[0]),.doutb(w_n1417_1[1]),.din(w_n1417_0[0]));
	jspl3 jspl3_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.doutc(w_n1425_0[2]),.din(n1425));
	jspl jspl_w_n1425_1(.douta(w_n1425_1[0]),.doutb(w_n1425_1[1]),.din(w_n1425_0[0]));
	jspl3 jspl3_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.doutc(w_n1433_0[2]),.din(n1433));
	jspl jspl_w_n1433_1(.douta(w_n1433_1[0]),.doutb(w_n1433_1[1]),.din(w_n1433_0[0]));
	jspl3 jspl3_w_n1442_0(.douta(w_n1442_0[0]),.doutb(w_n1442_0[1]),.doutc(w_n1442_0[2]),.din(n1442));
	jspl jspl_w_n1442_1(.douta(w_n1442_1[0]),.doutb(w_n1442_1[1]),.din(w_n1442_0[0]));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl3 jspl3_w_n1453_0(.douta(w_n1453_0[0]),.doutb(w_n1453_0[1]),.doutc(w_n1453_0[2]),.din(n1453));
	jspl jspl_w_n1453_1(.douta(w_n1453_1[0]),.doutb(w_n1453_1[1]),.din(w_n1453_0[0]));
	jspl3 jspl3_w_n1461_0(.douta(w_n1461_0[0]),.doutb(w_n1461_0[1]),.doutc(w_n1461_0[2]),.din(n1461));
	jspl jspl_w_n1461_1(.douta(w_n1461_1[0]),.doutb(w_n1461_1[1]),.din(w_n1461_0[0]));
	jspl3 jspl3_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.doutc(w_n1469_0[2]),.din(n1469));
	jspl jspl_w_n1469_1(.douta(w_n1469_1[0]),.doutb(w_n1469_1[1]),.din(w_n1469_0[0]));
	jspl3 jspl3_w_n1478_0(.douta(w_n1478_0[0]),.doutb(w_n1478_0[1]),.doutc(w_n1478_0[2]),.din(n1478));
	jspl jspl_w_n1478_1(.douta(w_n1478_1[0]),.doutb(w_n1478_1[1]),.din(w_n1478_0[0]));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(n1481));
	jspl3 jspl3_w_n1490_0(.douta(w_n1490_0[0]),.doutb(w_n1490_0[1]),.doutc(w_n1490_0[2]),.din(n1490));
	jspl jspl_w_n1490_1(.douta(w_n1490_1[0]),.doutb(w_n1490_1[1]),.din(w_n1490_0[0]));
	jspl3 jspl3_w_n1498_0(.douta(w_n1498_0[0]),.doutb(w_n1498_0[1]),.doutc(w_n1498_0[2]),.din(n1498));
	jspl jspl_w_n1498_1(.douta(w_n1498_1[0]),.doutb(w_n1498_1[1]),.din(w_n1498_0[0]));
	jspl3 jspl3_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.doutc(w_n1506_0[2]),.din(n1506));
	jspl jspl_w_n1506_1(.douta(w_n1506_1[0]),.doutb(w_n1506_1[1]),.din(w_n1506_0[0]));
	jspl3 jspl3_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.doutc(w_n1515_0[2]),.din(n1515));
	jspl jspl_w_n1515_1(.douta(w_n1515_1[0]),.doutb(w_n1515_1[1]),.din(w_n1515_0[0]));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl3 jspl3_w_n1526_0(.douta(w_n1526_0[0]),.doutb(w_n1526_0[1]),.doutc(w_n1526_0[2]),.din(n1526));
	jspl jspl_w_n1526_1(.douta(w_n1526_1[0]),.doutb(w_n1526_1[1]),.din(w_n1526_0[0]));
	jspl3 jspl3_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.doutc(w_n1534_0[2]),.din(n1534));
	jspl jspl_w_n1534_1(.douta(w_n1534_1[0]),.doutb(w_n1534_1[1]),.din(w_n1534_0[0]));
	jspl3 jspl3_w_n1542_0(.douta(w_n1542_0[0]),.doutb(w_n1542_0[1]),.doutc(w_n1542_0[2]),.din(n1542));
	jspl jspl_w_n1542_1(.douta(w_n1542_1[0]),.doutb(w_n1542_1[1]),.din(w_n1542_0[0]));
	jspl3 jspl3_w_n1551_0(.douta(w_n1551_0[0]),.doutb(w_n1551_0[1]),.doutc(w_n1551_0[2]),.din(n1551));
	jspl jspl_w_n1551_1(.douta(w_n1551_1[0]),.doutb(w_n1551_1[1]),.din(w_n1551_0[0]));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl3 jspl3_w_n1563_0(.douta(w_n1563_0[0]),.doutb(w_n1563_0[1]),.doutc(w_n1563_0[2]),.din(n1563));
	jspl jspl_w_n1563_1(.douta(w_n1563_1[0]),.doutb(w_n1563_1[1]),.din(w_n1563_0[0]));
	jspl3 jspl3_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.doutc(w_n1571_0[2]),.din(n1571));
	jspl jspl_w_n1571_1(.douta(w_n1571_1[0]),.doutb(w_n1571_1[1]),.din(w_n1571_0[0]));
	jspl3 jspl3_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.doutc(w_n1579_0[2]),.din(n1579));
	jspl jspl_w_n1579_1(.douta(w_n1579_1[0]),.doutb(w_n1579_1[1]),.din(w_n1579_0[0]));
	jspl3 jspl3_w_n1588_0(.douta(w_n1588_0[0]),.doutb(w_n1588_0[1]),.doutc(w_n1588_0[2]),.din(n1588));
	jspl jspl_w_n1588_1(.douta(w_n1588_1[0]),.doutb(w_n1588_1[1]),.din(w_n1588_0[0]));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl3 jspl3_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.doutc(w_n1599_0[2]),.din(n1599));
	jspl jspl_w_n1599_1(.douta(w_n1599_1[0]),.doutb(w_n1599_1[1]),.din(w_n1599_0[0]));
	jspl3 jspl3_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.doutc(w_n1607_0[2]),.din(n1607));
	jspl jspl_w_n1607_1(.douta(w_n1607_1[0]),.doutb(w_n1607_1[1]),.din(w_n1607_0[0]));
	jspl3 jspl3_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.doutc(w_n1615_0[2]),.din(n1615));
	jspl jspl_w_n1615_1(.douta(w_n1615_1[0]),.doutb(w_n1615_1[1]),.din(w_n1615_0[0]));
	jspl3 jspl3_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.doutc(w_n1624_0[2]),.din(n1624));
	jspl jspl_w_n1624_1(.douta(w_n1624_1[0]),.doutb(w_n1624_1[1]),.din(w_n1624_0[0]));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl3 jspl3_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.doutc(w_n1636_0[2]),.din(n1636));
	jspl jspl_w_n1636_1(.douta(w_n1636_1[0]),.doutb(w_n1636_1[1]),.din(w_n1636_0[0]));
	jspl3 jspl3_w_n1644_0(.douta(w_n1644_0[0]),.doutb(w_n1644_0[1]),.doutc(w_n1644_0[2]),.din(n1644));
	jspl jspl_w_n1644_1(.douta(w_n1644_1[0]),.doutb(w_n1644_1[1]),.din(w_n1644_0[0]));
	jspl3 jspl3_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_n1652_0[1]),.doutc(w_n1652_0[2]),.din(n1652));
	jspl jspl_w_n1652_1(.douta(w_n1652_1[0]),.doutb(w_n1652_1[1]),.din(w_n1652_0[0]));
	jspl3 jspl3_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.doutc(w_n1661_0[2]),.din(n1661));
	jspl jspl_w_n1661_1(.douta(w_n1661_1[0]),.doutb(w_n1661_1[1]),.din(w_n1661_0[0]));
	jspl jspl_w_n1664_0(.douta(w_n1664_0[0]),.doutb(w_n1664_0[1]),.din(n1664));
	jspl3 jspl3_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.doutc(w_n1672_0[2]),.din(n1672));
	jspl jspl_w_n1672_1(.douta(w_n1672_1[0]),.doutb(w_n1672_1[1]),.din(w_n1672_0[0]));
	jspl3 jspl3_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.doutc(w_n1680_0[2]),.din(n1680));
	jspl jspl_w_n1680_1(.douta(w_n1680_1[0]),.doutb(w_n1680_1[1]),.din(w_n1680_0[0]));
	jspl3 jspl3_w_n1688_0(.douta(w_n1688_0[0]),.doutb(w_n1688_0[1]),.doutc(w_n1688_0[2]),.din(n1688));
	jspl jspl_w_n1688_1(.douta(w_n1688_1[0]),.doutb(w_n1688_1[1]),.din(w_n1688_0[0]));
	jspl3 jspl3_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_n1697_0[1]),.doutc(w_n1697_0[2]),.din(n1697));
	jspl jspl_w_n1697_1(.douta(w_n1697_1[0]),.doutb(w_n1697_1[1]),.din(w_n1697_0[0]));
	jspl jspl_w_n1700_0(.douta(w_n1700_0[0]),.doutb(w_n1700_0[1]),.din(n1700));
	jspl3 jspl3_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.doutc(w_n1709_0[2]),.din(n1709));
	jspl jspl_w_n1709_1(.douta(w_n1709_1[0]),.doutb(w_n1709_1[1]),.din(w_n1709_0[0]));
	jspl3 jspl3_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.doutc(w_n1717_0[2]),.din(n1717));
	jspl jspl_w_n1717_1(.douta(w_n1717_1[0]),.doutb(w_n1717_1[1]),.din(w_n1717_0[0]));
	jspl3 jspl3_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.doutc(w_n1725_0[2]),.din(n1725));
	jspl jspl_w_n1725_1(.douta(w_n1725_1[0]),.doutb(w_n1725_1[1]),.din(w_n1725_0[0]));
	jspl3 jspl3_w_n1734_0(.douta(w_n1734_0[0]),.doutb(w_n1734_0[1]),.doutc(w_n1734_0[2]),.din(n1734));
	jspl jspl_w_n1734_1(.douta(w_n1734_1[0]),.doutb(w_n1734_1[1]),.din(w_n1734_0[0]));
	jspl jspl_w_n1737_0(.douta(w_n1737_0[0]),.doutb(w_n1737_0[1]),.din(n1737));
	jspl3 jspl3_w_n1745_0(.douta(w_n1745_0[0]),.doutb(w_n1745_0[1]),.doutc(w_n1745_0[2]),.din(n1745));
	jspl jspl_w_n1745_1(.douta(w_n1745_1[0]),.doutb(w_n1745_1[1]),.din(w_n1745_0[0]));
	jspl3 jspl3_w_n1753_0(.douta(w_n1753_0[0]),.doutb(w_n1753_0[1]),.doutc(w_n1753_0[2]),.din(n1753));
	jspl jspl_w_n1753_1(.douta(w_n1753_1[0]),.doutb(w_n1753_1[1]),.din(w_n1753_0[0]));
	jspl3 jspl3_w_n1761_0(.douta(w_n1761_0[0]),.doutb(w_n1761_0[1]),.doutc(w_n1761_0[2]),.din(n1761));
	jspl jspl_w_n1761_1(.douta(w_n1761_1[0]),.doutb(w_n1761_1[1]),.din(w_n1761_0[0]));
	jspl3 jspl3_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.doutc(w_n1770_0[2]),.din(n1770));
	jspl jspl_w_n1770_1(.douta(w_n1770_1[0]),.doutb(w_n1770_1[1]),.din(w_n1770_0[0]));
	jspl jspl_w_n1773_0(.douta(w_n1773_0[0]),.doutb(w_n1773_0[1]),.din(n1773));
	jspl3 jspl3_w_n1782_0(.douta(w_n1782_0[0]),.doutb(w_n1782_0[1]),.doutc(w_n1782_0[2]),.din(n1782));
	jspl jspl_w_n1782_1(.douta(w_n1782_1[0]),.doutb(w_n1782_1[1]),.din(w_n1782_0[0]));
	jspl3 jspl3_w_n1790_0(.douta(w_n1790_0[0]),.doutb(w_n1790_0[1]),.doutc(w_n1790_0[2]),.din(n1790));
	jspl jspl_w_n1790_1(.douta(w_n1790_1[0]),.doutb(w_n1790_1[1]),.din(w_n1790_0[0]));
	jspl3 jspl3_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.doutc(w_n1798_0[2]),.din(n1798));
	jspl jspl_w_n1798_1(.douta(w_n1798_1[0]),.doutb(w_n1798_1[1]),.din(w_n1798_0[0]));
	jspl3 jspl3_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.doutc(w_n1807_0[2]),.din(n1807));
	jspl jspl_w_n1807_1(.douta(w_n1807_1[0]),.doutb(w_n1807_1[1]),.din(w_n1807_0[0]));
	jspl jspl_w_n1810_0(.douta(w_n1810_0[0]),.doutb(w_n1810_0[1]),.din(n1810));
	jspl3 jspl3_w_n1818_0(.douta(w_n1818_0[0]),.doutb(w_n1818_0[1]),.doutc(w_n1818_0[2]),.din(n1818));
	jspl jspl_w_n1818_1(.douta(w_n1818_1[0]),.doutb(w_n1818_1[1]),.din(w_n1818_0[0]));
	jspl3 jspl3_w_n1826_0(.douta(w_n1826_0[0]),.doutb(w_n1826_0[1]),.doutc(w_n1826_0[2]),.din(n1826));
	jspl jspl_w_n1826_1(.douta(w_n1826_1[0]),.doutb(w_n1826_1[1]),.din(w_n1826_0[0]));
	jspl3 jspl3_w_n1834_0(.douta(w_n1834_0[0]),.doutb(w_n1834_0[1]),.doutc(w_n1834_0[2]),.din(n1834));
	jspl jspl_w_n1834_1(.douta(w_n1834_1[0]),.doutb(w_n1834_1[1]),.din(w_n1834_0[0]));
	jspl3 jspl3_w_n1843_0(.douta(w_n1843_0[0]),.doutb(w_n1843_0[1]),.doutc(w_n1843_0[2]),.din(n1843));
	jspl jspl_w_n1843_1(.douta(w_n1843_1[0]),.doutb(w_n1843_1[1]),.din(w_n1843_0[0]));
	jspl jspl_w_n1846_0(.douta(w_n1846_0[0]),.doutb(w_n1846_0[1]),.din(n1846));
	jspl3 jspl3_w_n1855_0(.douta(w_n1855_0[0]),.doutb(w_n1855_0[1]),.doutc(w_n1855_0[2]),.din(n1855));
	jspl jspl_w_n1855_1(.douta(w_n1855_1[0]),.doutb(w_n1855_1[1]),.din(w_n1855_0[0]));
	jspl3 jspl3_w_n1863_0(.douta(w_n1863_0[0]),.doutb(w_n1863_0[1]),.doutc(w_n1863_0[2]),.din(n1863));
	jspl jspl_w_n1863_1(.douta(w_n1863_1[0]),.doutb(w_n1863_1[1]),.din(w_n1863_0[0]));
	jspl3 jspl3_w_n1871_0(.douta(w_n1871_0[0]),.doutb(w_n1871_0[1]),.doutc(w_n1871_0[2]),.din(n1871));
	jspl jspl_w_n1871_1(.douta(w_n1871_1[0]),.doutb(w_n1871_1[1]),.din(w_n1871_0[0]));
	jspl3 jspl3_w_n1880_0(.douta(w_n1880_0[0]),.doutb(w_n1880_0[1]),.doutc(w_n1880_0[2]),.din(n1880));
	jspl jspl_w_n1880_1(.douta(w_n1880_1[0]),.doutb(w_n1880_1[1]),.din(w_n1880_0[0]));
	jspl jspl_w_n1883_0(.douta(w_n1883_0[0]),.doutb(w_n1883_0[1]),.din(n1883));
	jspl3 jspl3_w_n1891_0(.douta(w_n1891_0[0]),.doutb(w_n1891_0[1]),.doutc(w_n1891_0[2]),.din(n1891));
	jspl jspl_w_n1891_1(.douta(w_n1891_1[0]),.doutb(w_n1891_1[1]),.din(w_n1891_0[0]));
	jspl3 jspl3_w_n1899_0(.douta(w_n1899_0[0]),.doutb(w_n1899_0[1]),.doutc(w_n1899_0[2]),.din(n1899));
	jspl jspl_w_n1899_1(.douta(w_n1899_1[0]),.doutb(w_n1899_1[1]),.din(w_n1899_0[0]));
	jspl3 jspl3_w_n1907_0(.douta(w_n1907_0[0]),.doutb(w_n1907_0[1]),.doutc(w_n1907_0[2]),.din(n1907));
	jspl jspl_w_n1907_1(.douta(w_n1907_1[0]),.doutb(w_n1907_1[1]),.din(w_n1907_0[0]));
	jspl3 jspl3_w_n1916_0(.douta(w_n1916_0[0]),.doutb(w_n1916_0[1]),.doutc(w_n1916_0[2]),.din(n1916));
	jspl jspl_w_n1916_1(.douta(w_n1916_1[0]),.doutb(w_n1916_1[1]),.din(w_n1916_0[0]));
	jspl jspl_w_n1919_0(.douta(w_n1919_0[0]),.doutb(w_n1919_0[1]),.din(n1919));
	jspl3 jspl3_w_n1928_0(.douta(w_n1928_0[0]),.doutb(w_n1928_0[1]),.doutc(w_n1928_0[2]),.din(n1928));
	jspl jspl_w_n1928_1(.douta(w_n1928_1[0]),.doutb(w_n1928_1[1]),.din(w_n1928_0[0]));
	jspl3 jspl3_w_n1936_0(.douta(w_n1936_0[0]),.doutb(w_n1936_0[1]),.doutc(w_n1936_0[2]),.din(n1936));
	jspl jspl_w_n1936_1(.douta(w_n1936_1[0]),.doutb(w_n1936_1[1]),.din(w_n1936_0[0]));
	jspl3 jspl3_w_n1944_0(.douta(w_n1944_0[0]),.doutb(w_n1944_0[1]),.doutc(w_n1944_0[2]),.din(n1944));
	jspl jspl_w_n1944_1(.douta(w_n1944_1[0]),.doutb(w_n1944_1[1]),.din(w_n1944_0[0]));
	jspl3 jspl3_w_n1953_0(.douta(w_n1953_0[0]),.doutb(w_n1953_0[1]),.doutc(w_n1953_0[2]),.din(n1953));
	jspl jspl_w_n1953_1(.douta(w_n1953_1[0]),.doutb(w_n1953_1[1]),.din(w_n1953_0[0]));
	jspl jspl_w_n1956_0(.douta(w_n1956_0[0]),.doutb(w_n1956_0[1]),.din(n1956));
	jspl3 jspl3_w_n1964_0(.douta(w_n1964_0[0]),.doutb(w_n1964_0[1]),.doutc(w_n1964_0[2]),.din(n1964));
	jspl jspl_w_n1964_1(.douta(w_n1964_1[0]),.doutb(w_n1964_1[1]),.din(w_n1964_0[0]));
	jspl3 jspl3_w_n1972_0(.douta(w_n1972_0[0]),.doutb(w_n1972_0[1]),.doutc(w_n1972_0[2]),.din(n1972));
	jspl jspl_w_n1972_1(.douta(w_n1972_1[0]),.doutb(w_n1972_1[1]),.din(w_n1972_0[0]));
	jspl3 jspl3_w_n1980_0(.douta(w_n1980_0[0]),.doutb(w_n1980_0[1]),.doutc(w_n1980_0[2]),.din(n1980));
	jspl jspl_w_n1980_1(.douta(w_n1980_1[0]),.doutb(w_n1980_1[1]),.din(w_n1980_0[0]));
	jspl3 jspl3_w_n1989_0(.douta(w_n1989_0[0]),.doutb(w_n1989_0[1]),.doutc(w_n1989_0[2]),.din(n1989));
	jspl jspl_w_n1989_1(.douta(w_n1989_1[0]),.doutb(w_n1989_1[1]),.din(w_n1989_0[0]));
	jspl jspl_w_n1992_0(.douta(w_n1992_0[0]),.doutb(w_n1992_0[1]),.din(n1992));
	jspl3 jspl3_w_n2001_0(.douta(w_n2001_0[0]),.doutb(w_n2001_0[1]),.doutc(w_n2001_0[2]),.din(n2001));
	jspl jspl_w_n2001_1(.douta(w_n2001_1[0]),.doutb(w_n2001_1[1]),.din(w_n2001_0[0]));
	jspl3 jspl3_w_n2009_0(.douta(w_n2009_0[0]),.doutb(w_n2009_0[1]),.doutc(w_n2009_0[2]),.din(n2009));
	jspl jspl_w_n2009_1(.douta(w_n2009_1[0]),.doutb(w_n2009_1[1]),.din(w_n2009_0[0]));
	jspl3 jspl3_w_n2017_0(.douta(w_n2017_0[0]),.doutb(w_n2017_0[1]),.doutc(w_n2017_0[2]),.din(n2017));
	jspl jspl_w_n2017_1(.douta(w_n2017_1[0]),.doutb(w_n2017_1[1]),.din(w_n2017_0[0]));
	jspl3 jspl3_w_n2026_0(.douta(w_n2026_0[0]),.doutb(w_n2026_0[1]),.doutc(w_n2026_0[2]),.din(n2026));
	jspl jspl_w_n2026_1(.douta(w_n2026_1[0]),.doutb(w_n2026_1[1]),.din(w_n2026_0[0]));
	jspl jspl_w_n2029_0(.douta(w_n2029_0[0]),.doutb(w_n2029_0[1]),.din(n2029));
	jspl3 jspl3_w_n2037_0(.douta(w_n2037_0[0]),.doutb(w_n2037_0[1]),.doutc(w_n2037_0[2]),.din(n2037));
	jspl jspl_w_n2037_1(.douta(w_n2037_1[0]),.doutb(w_n2037_1[1]),.din(w_n2037_0[0]));
	jspl3 jspl3_w_n2045_0(.douta(w_n2045_0[0]),.doutb(w_n2045_0[1]),.doutc(w_n2045_0[2]),.din(n2045));
	jspl jspl_w_n2045_1(.douta(w_n2045_1[0]),.doutb(w_n2045_1[1]),.din(w_n2045_0[0]));
	jspl3 jspl3_w_n2053_0(.douta(w_n2053_0[0]),.doutb(w_n2053_0[1]),.doutc(w_n2053_0[2]),.din(n2053));
	jspl jspl_w_n2053_1(.douta(w_n2053_1[0]),.doutb(w_n2053_1[1]),.din(w_n2053_0[0]));
	jspl3 jspl3_w_n2062_0(.douta(w_n2062_0[0]),.doutb(w_n2062_0[1]),.doutc(w_n2062_0[2]),.din(n2062));
	jspl jspl_w_n2062_1(.douta(w_n2062_1[0]),.doutb(w_n2062_1[1]),.din(w_n2062_0[0]));
	jspl jspl_w_n2065_0(.douta(w_n2065_0[0]),.doutb(w_n2065_0[1]),.din(n2065));
	jspl3 jspl3_w_n2074_0(.douta(w_n2074_0[0]),.doutb(w_n2074_0[1]),.doutc(w_n2074_0[2]),.din(n2074));
	jspl jspl_w_n2074_1(.douta(w_n2074_1[0]),.doutb(w_n2074_1[1]),.din(w_n2074_0[0]));
	jspl3 jspl3_w_n2082_0(.douta(w_n2082_0[0]),.doutb(w_n2082_0[1]),.doutc(w_n2082_0[2]),.din(n2082));
	jspl jspl_w_n2082_1(.douta(w_n2082_1[0]),.doutb(w_n2082_1[1]),.din(w_n2082_0[0]));
	jspl3 jspl3_w_n2090_0(.douta(w_n2090_0[0]),.doutb(w_n2090_0[1]),.doutc(w_n2090_0[2]),.din(n2090));
	jspl jspl_w_n2090_1(.douta(w_n2090_1[0]),.doutb(w_n2090_1[1]),.din(w_n2090_0[0]));
	jspl3 jspl3_w_n2099_0(.douta(w_n2099_0[0]),.doutb(w_n2099_0[1]),.doutc(w_n2099_0[2]),.din(n2099));
	jspl jspl_w_n2099_1(.douta(w_n2099_1[0]),.doutb(w_n2099_1[1]),.din(w_n2099_0[0]));
	jspl jspl_w_n2102_0(.douta(w_n2102_0[0]),.doutb(w_n2102_0[1]),.din(n2102));
	jspl3 jspl3_w_n2110_0(.douta(w_n2110_0[0]),.doutb(w_n2110_0[1]),.doutc(w_n2110_0[2]),.din(n2110));
	jspl jspl_w_n2110_1(.douta(w_n2110_1[0]),.doutb(w_n2110_1[1]),.din(w_n2110_0[0]));
	jspl3 jspl3_w_n2118_0(.douta(w_n2118_0[0]),.doutb(w_n2118_0[1]),.doutc(w_n2118_0[2]),.din(n2118));
	jspl jspl_w_n2118_1(.douta(w_n2118_1[0]),.doutb(w_n2118_1[1]),.din(w_n2118_0[0]));
	jspl3 jspl3_w_n2126_0(.douta(w_n2126_0[0]),.doutb(w_n2126_0[1]),.doutc(w_n2126_0[2]),.din(n2126));
	jspl jspl_w_n2126_1(.douta(w_n2126_1[0]),.doutb(w_n2126_1[1]),.din(w_n2126_0[0]));
	jspl3 jspl3_w_n2135_0(.douta(w_n2135_0[0]),.doutb(w_n2135_0[1]),.doutc(w_n2135_0[2]),.din(n2135));
	jspl jspl_w_n2135_1(.douta(w_n2135_1[0]),.doutb(w_n2135_1[1]),.din(w_n2135_0[0]));
	jspl jspl_w_n2138_0(.douta(w_n2138_0[0]),.doutb(w_n2138_0[1]),.din(n2138));
	jspl3 jspl3_w_n2147_0(.douta(w_n2147_0[0]),.doutb(w_n2147_0[1]),.doutc(w_n2147_0[2]),.din(n2147));
	jspl jspl_w_n2147_1(.douta(w_n2147_1[0]),.doutb(w_n2147_1[1]),.din(w_n2147_0[0]));
	jspl3 jspl3_w_n2155_0(.douta(w_n2155_0[0]),.doutb(w_n2155_0[1]),.doutc(w_n2155_0[2]),.din(n2155));
	jspl jspl_w_n2155_1(.douta(w_n2155_1[0]),.doutb(w_n2155_1[1]),.din(w_n2155_0[0]));
	jspl3 jspl3_w_n2163_0(.douta(w_n2163_0[0]),.doutb(w_n2163_0[1]),.doutc(w_n2163_0[2]),.din(n2163));
	jspl jspl_w_n2163_1(.douta(w_n2163_1[0]),.doutb(w_n2163_1[1]),.din(w_n2163_0[0]));
	jspl3 jspl3_w_n2172_0(.douta(w_n2172_0[0]),.doutb(w_n2172_0[1]),.doutc(w_n2172_0[2]),.din(n2172));
	jspl jspl_w_n2172_1(.douta(w_n2172_1[0]),.doutb(w_n2172_1[1]),.din(w_n2172_0[0]));
	jspl jspl_w_n2175_0(.douta(w_n2175_0[0]),.doutb(w_n2175_0[1]),.din(n2175));
	jspl3 jspl3_w_n2183_0(.douta(w_n2183_0[0]),.doutb(w_n2183_0[1]),.doutc(w_n2183_0[2]),.din(n2183));
	jspl jspl_w_n2183_1(.douta(w_n2183_1[0]),.doutb(w_n2183_1[1]),.din(w_n2183_0[0]));
	jspl3 jspl3_w_n2191_0(.douta(w_n2191_0[0]),.doutb(w_n2191_0[1]),.doutc(w_n2191_0[2]),.din(n2191));
	jspl jspl_w_n2191_1(.douta(w_n2191_1[0]),.doutb(w_n2191_1[1]),.din(w_n2191_0[0]));
	jspl3 jspl3_w_n2199_0(.douta(w_n2199_0[0]),.doutb(w_n2199_0[1]),.doutc(w_n2199_0[2]),.din(n2199));
	jspl jspl_w_n2199_1(.douta(w_n2199_1[0]),.doutb(w_n2199_1[1]),.din(w_n2199_0[0]));
	jspl3 jspl3_w_n2208_0(.douta(w_n2208_0[0]),.doutb(w_n2208_0[1]),.doutc(w_n2208_0[2]),.din(n2208));
	jspl jspl_w_n2208_1(.douta(w_n2208_1[0]),.doutb(w_n2208_1[1]),.din(w_n2208_0[0]));
	jspl jspl_w_n2211_0(.douta(w_n2211_0[0]),.doutb(w_n2211_0[1]),.din(n2211));
	jspl jspl_w_n2220_0(.douta(w_n2220_0[0]),.doutb(w_n2220_0[1]),.din(n2220));
	jspl jspl_w_n2228_0(.douta(w_n2228_0[0]),.doutb(w_n2228_0[1]),.din(n2228));
	jspl jspl_w_n2237_0(.douta(w_n2237_0[0]),.doutb(w_n2237_0[1]),.din(n2237));
	jspl jspl_w_n2245_0(.douta(w_n2245_0[0]),.doutb(w_n2245_0[1]),.din(n2245));
	jspl jspl_w_n2254_0(.douta(w_n2254_0[0]),.doutb(w_n2254_0[1]),.din(n2254));
	jspl jspl_w_n2262_0(.douta(w_n2262_0[0]),.doutb(w_n2262_0[1]),.din(n2262));
	jspl jspl_w_n2271_0(.douta(w_n2271_0[0]),.doutb(w_n2271_0[1]),.din(n2271));
	jspl jspl_w_n2279_0(.douta(w_n2279_0[0]),.doutb(w_n2279_0[1]),.din(n2279));
	jspl jspl_w_n2288_0(.douta(w_n2288_0[0]),.doutb(w_n2288_0[1]),.din(n2288));
	jspl jspl_w_n2296_0(.douta(w_n2296_0[0]),.doutb(w_n2296_0[1]),.din(n2296));
	jspl jspl_w_n2305_0(.douta(w_n2305_0[0]),.doutb(w_n2305_0[1]),.din(n2305));
	jspl jspl_w_n2313_0(.douta(w_n2313_0[0]),.doutb(w_n2313_0[1]),.din(n2313));
	jspl jspl_w_n2322_0(.douta(w_n2322_0[0]),.doutb(w_n2322_0[1]),.din(n2322));
	jspl jspl_w_n2330_0(.douta(w_n2330_0[0]),.doutb(w_n2330_0[1]),.din(n2330));
	jspl jspl_w_n2339_0(.douta(w_n2339_0[0]),.doutb(w_n2339_0[1]),.din(n2339));
	jspl jspl_w_n2347_0(.douta(w_n2347_0[0]),.doutb(w_n2347_0[1]),.din(n2347));
	jspl jspl_w_n2356_0(.douta(w_n2356_0[0]),.doutb(w_n2356_0[1]),.din(n2356));
	jspl jspl_w_n2364_0(.douta(w_n2364_0[0]),.doutb(w_n2364_0[1]),.din(n2364));
	jspl jspl_w_n2373_0(.douta(w_n2373_0[0]),.doutb(w_n2373_0[1]),.din(n2373));
	jspl jspl_w_n2381_0(.douta(w_n2381_0[0]),.doutb(w_n2381_0[1]),.din(n2381));
	jspl jspl_w_n2390_0(.douta(w_n2390_0[0]),.doutb(w_n2390_0[1]),.din(n2390));
	jspl jspl_w_n2398_0(.douta(w_n2398_0[0]),.doutb(w_n2398_0[1]),.din(n2398));
	jspl jspl_w_n2407_0(.douta(w_n2407_0[0]),.doutb(w_n2407_0[1]),.din(n2407));
	jspl jspl_w_n2415_0(.douta(w_n2415_0[0]),.doutb(w_n2415_0[1]),.din(n2415));
	jspl jspl_w_n2424_0(.douta(w_n2424_0[0]),.doutb(w_n2424_0[1]),.din(n2424));
	jspl jspl_w_n2432_0(.douta(w_n2432_0[0]),.doutb(w_n2432_0[1]),.din(n2432));
	jspl jspl_w_n2441_0(.douta(w_n2441_0[0]),.doutb(w_n2441_0[1]),.din(n2441));
	jspl jspl_w_n2449_0(.douta(w_n2449_0[0]),.doutb(w_n2449_0[1]),.din(n2449));
	jspl jspl_w_n2458_0(.douta(w_n2458_0[0]),.doutb(w_n2458_0[1]),.din(n2458));
	jspl jspl_w_n2466_0(.douta(w_n2466_0[0]),.doutb(w_n2466_0[1]),.din(n2466));
	jspl jspl_w_n2475_0(.douta(w_n2475_0[0]),.doutb(w_n2475_0[1]),.din(n2475));
	jspl jspl_w_n2483_0(.douta(w_n2483_0[0]),.doutb(w_n2483_0[1]),.din(n2483));
	jspl jspl_w_n2492_0(.douta(w_n2492_0[0]),.doutb(w_n2492_0[1]),.din(n2492));
	jspl jspl_w_n2500_0(.douta(w_n2500_0[0]),.doutb(w_n2500_0[1]),.din(n2500));
	jspl jspl_w_n2509_0(.douta(w_n2509_0[0]),.doutb(w_n2509_0[1]),.din(n2509));
	jspl jspl_w_n2517_0(.douta(w_n2517_0[0]),.doutb(w_n2517_0[1]),.din(n2517));
	jspl jspl_w_n2526_0(.douta(w_n2526_0[0]),.doutb(w_n2526_0[1]),.din(n2526));
	jspl jspl_w_n2534_0(.douta(w_n2534_0[0]),.doutb(w_n2534_0[1]),.din(n2534));
	jspl jspl_w_n2543_0(.douta(w_n2543_0[0]),.doutb(w_n2543_0[1]),.din(n2543));
	jspl jspl_w_n2551_0(.douta(w_n2551_0[0]),.doutb(w_n2551_0[1]),.din(n2551));
	jspl jspl_w_n2560_0(.douta(w_n2560_0[0]),.doutb(w_n2560_0[1]),.din(n2560));
	jspl jspl_w_n2568_0(.douta(w_n2568_0[0]),.doutb(w_n2568_0[1]),.din(n2568));
	jspl jspl_w_n2577_0(.douta(w_n2577_0[0]),.doutb(w_n2577_0[1]),.din(n2577));
	jspl jspl_w_n2585_0(.douta(w_n2585_0[0]),.doutb(w_n2585_0[1]),.din(n2585));
	jspl jspl_w_n2594_0(.douta(w_n2594_0[0]),.doutb(w_n2594_0[1]),.din(n2594));
	jspl jspl_w_n2602_0(.douta(w_n2602_0[0]),.doutb(w_n2602_0[1]),.din(n2602));
	jspl jspl_w_n2611_0(.douta(w_n2611_0[0]),.doutb(w_n2611_0[1]),.din(n2611));
	jspl jspl_w_n2619_0(.douta(w_n2619_0[0]),.doutb(w_n2619_0[1]),.din(n2619));
	jspl jspl_w_n2628_0(.douta(w_n2628_0[0]),.doutb(w_n2628_0[1]),.din(n2628));
	jspl jspl_w_n2636_0(.douta(w_n2636_0[0]),.doutb(w_n2636_0[1]),.din(n2636));
	jspl jspl_w_n2645_0(.douta(w_n2645_0[0]),.doutb(w_n2645_0[1]),.din(n2645));
	jspl jspl_w_n2653_0(.douta(w_n2653_0[0]),.doutb(w_n2653_0[1]),.din(n2653));
	jspl jspl_w_n2662_0(.douta(w_n2662_0[0]),.doutb(w_n2662_0[1]),.din(n2662));
	jspl jspl_w_n2670_0(.douta(w_n2670_0[0]),.doutb(w_n2670_0[1]),.din(n2670));
	jspl jspl_w_n2679_0(.douta(w_n2679_0[0]),.doutb(w_n2679_0[1]),.din(n2679));
	jspl jspl_w_n2687_0(.douta(w_n2687_0[0]),.doutb(w_n2687_0[1]),.din(n2687));
	jspl jspl_w_n2696_0(.douta(w_n2696_0[0]),.doutb(w_n2696_0[1]),.din(n2696));
	jspl jspl_w_n2704_0(.douta(w_n2704_0[0]),.doutb(w_n2704_0[1]),.din(n2704));
	jspl jspl_w_n2713_0(.douta(w_n2713_0[0]),.doutb(w_n2713_0[1]),.din(n2713));
	jspl jspl_w_n2721_0(.douta(w_n2721_0[0]),.doutb(w_n2721_0[1]),.din(n2721));
	jspl jspl_w_n2730_0(.douta(w_n2730_0[0]),.doutb(w_n2730_0[1]),.din(n2730));
	jspl jspl_w_n2738_0(.douta(w_n2738_0[0]),.doutb(w_n2738_0[1]),.din(n2738));
	jspl jspl_w_n2747_0(.douta(w_n2747_0[0]),.doutb(w_n2747_0[1]),.din(n2747));
	jspl jspl_w_n2755_0(.douta(w_n2755_0[0]),.doutb(w_n2755_0[1]),.din(n2755));
	jspl jspl_w_n2764_0(.douta(w_n2764_0[0]),.doutb(w_n2764_0[1]),.din(n2764));
	jspl jspl_w_n2772_0(.douta(w_n2772_0[0]),.doutb(w_n2772_0[1]),.din(n2772));
	jspl jspl_w_n2781_0(.douta(w_n2781_0[0]),.doutb(w_n2781_0[1]),.din(n2781));
	jspl jspl_w_n2789_0(.douta(w_n2789_0[0]),.doutb(w_n2789_0[1]),.din(n2789));
	jspl jspl_w_n2798_0(.douta(w_n2798_0[0]),.doutb(w_n2798_0[1]),.din(n2798));
	jspl jspl_w_n2806_0(.douta(w_n2806_0[0]),.doutb(w_n2806_0[1]),.din(n2806));
	jspl jspl_w_n2815_0(.douta(w_n2815_0[0]),.doutb(w_n2815_0[1]),.din(n2815));
	jspl jspl_w_n2823_0(.douta(w_n2823_0[0]),.doutb(w_n2823_0[1]),.din(n2823));
	jspl jspl_w_n2832_0(.douta(w_n2832_0[0]),.doutb(w_n2832_0[1]),.din(n2832));
	jspl jspl_w_n2840_0(.douta(w_n2840_0[0]),.doutb(w_n2840_0[1]),.din(n2840));
	jspl jspl_w_n2849_0(.douta(w_n2849_0[0]),.doutb(w_n2849_0[1]),.din(n2849));
	jspl jspl_w_n2857_0(.douta(w_n2857_0[0]),.doutb(w_n2857_0[1]),.din(n2857));
	jspl jspl_w_n2866_0(.douta(w_n2866_0[0]),.doutb(w_n2866_0[1]),.din(n2866));
	jspl jspl_w_n2874_0(.douta(w_n2874_0[0]),.doutb(w_n2874_0[1]),.din(n2874));
	jspl jspl_w_n2883_0(.douta(w_n2883_0[0]),.doutb(w_n2883_0[1]),.din(n2883));
	jspl jspl_w_n2891_0(.douta(w_n2891_0[0]),.doutb(w_n2891_0[1]),.din(n2891));
	jspl jspl_w_n2900_0(.douta(w_n2900_0[0]),.doutb(w_n2900_0[1]),.din(n2900));
	jspl jspl_w_n2908_0(.douta(w_n2908_0[0]),.doutb(w_n2908_0[1]),.din(n2908));
	jspl jspl_w_n2917_0(.douta(w_n2917_0[0]),.doutb(w_n2917_0[1]),.din(n2917));
	jspl jspl_w_n2925_0(.douta(w_n2925_0[0]),.doutb(w_n2925_0[1]),.din(n2925));
	jspl jspl_w_n2934_0(.douta(w_n2934_0[0]),.doutb(w_n2934_0[1]),.din(n2934));
	jspl jspl_w_n2942_0(.douta(w_n2942_0[0]),.doutb(w_n2942_0[1]),.din(n2942));
	jspl jspl_w_n2951_0(.douta(w_n2951_0[0]),.doutb(w_n2951_0[1]),.din(n2951));
	jspl jspl_w_n2959_0(.douta(w_n2959_0[0]),.doutb(w_n2959_0[1]),.din(n2959));
	jspl jspl_w_n2968_0(.douta(w_n2968_0[0]),.doutb(w_n2968_0[1]),.din(n2968));
	jspl jspl_w_n2976_0(.douta(w_n2976_0[0]),.doutb(w_n2976_0[1]),.din(n2976));
	jspl jspl_w_n2985_0(.douta(w_n2985_0[0]),.doutb(w_n2985_0[1]),.din(n2985));
	jspl jspl_w_n2993_0(.douta(w_n2993_0[0]),.doutb(w_n2993_0[1]),.din(n2993));
	jspl jspl_w_n3002_0(.douta(w_n3002_0[0]),.doutb(w_n3002_0[1]),.din(n3002));
	jspl jspl_w_n3010_0(.douta(w_n3010_0[0]),.doutb(w_n3010_0[1]),.din(n3010));
	jspl jspl_w_n3019_0(.douta(w_n3019_0[0]),.doutb(w_n3019_0[1]),.din(n3019));
	jspl jspl_w_n3027_0(.douta(w_n3027_0[0]),.doutb(w_n3027_0[1]),.din(n3027));
	jdff dff_B_g1C06Xx82_1(.din(n317),.dout(w_dff_B_g1C06Xx82_1),.clk(gclk));
	jdff dff_B_IqnWAkCL7_1(.din(w_dff_B_g1C06Xx82_1),.dout(w_dff_B_IqnWAkCL7_1),.clk(gclk));
	jdff dff_B_HpkFhe6A1_0(.din(n454),.dout(w_dff_B_HpkFhe6A1_0),.clk(gclk));
	jdff dff_B_JoZ9Tb4V2_1(.din(n501),.dout(w_dff_B_JoZ9Tb4V2_1),.clk(gclk));
	jdff dff_B_UCm236lc9_1(.din(w_dff_B_JoZ9Tb4V2_1),.dout(w_dff_B_UCm236lc9_1),.clk(gclk));
	jdff dff_B_xuHcFHr59_0(.din(n634),.dout(w_dff_B_xuHcFHr59_0),.clk(gclk));
	jdff dff_B_T8KfLGzT2_1(.din(n682),.dout(w_dff_B_T8KfLGzT2_1),.clk(gclk));
	jdff dff_B_E17iQHOA7_1(.din(w_dff_B_T8KfLGzT2_1),.dout(w_dff_B_E17iQHOA7_1),.clk(gclk));
	jdff dff_B_gRp8Ggs88_0(.din(n815),.dout(w_dff_B_gRp8Ggs88_0),.clk(gclk));
	jdff dff_B_lIe0sgd26_1(.din(n862),.dout(w_dff_B_lIe0sgd26_1),.clk(gclk));
	jdff dff_B_WfEiqaoK6_1(.din(w_dff_B_lIe0sgd26_1),.dout(w_dff_B_WfEiqaoK6_1),.clk(gclk));
	jdff dff_B_cjYulRxp8_0(.din(n995),.dout(w_dff_B_cjYulRxp8_0),.clk(gclk));
	jdff dff_B_D8gYIS3H8_1(.din(n1019),.dout(w_dff_B_D8gYIS3H8_1),.clk(gclk));
	jdff dff_B_ZbjPw7uh6_1(.din(w_dff_B_D8gYIS3H8_1),.dout(w_dff_B_ZbjPw7uh6_1),.clk(gclk));
	jdff dff_B_NanY4bA49_0(.din(n1080),.dout(w_dff_B_NanY4bA49_0),.clk(gclk));
	jdff dff_B_2N8mDzIw8_1(.din(n1103),.dout(w_dff_B_2N8mDzIw8_1),.clk(gclk));
	jdff dff_B_wVw0jevq6_1(.din(w_dff_B_2N8mDzIw8_1),.dout(w_dff_B_wVw0jevq6_1),.clk(gclk));
	jdff dff_B_U2b0FtDF4_0(.din(n1164),.dout(w_dff_B_U2b0FtDF4_0),.clk(gclk));
	jdff dff_B_wMj82kuC6_1(.din(n1188),.dout(w_dff_B_wMj82kuC6_1),.clk(gclk));
	jdff dff_B_x7FH33QW3_1(.din(w_dff_B_wMj82kuC6_1),.dout(w_dff_B_x7FH33QW3_1),.clk(gclk));
	jdff dff_B_PVP23snq0_0(.din(n1249),.dout(w_dff_B_PVP23snq0_0),.clk(gclk));
	jdff dff_B_rYsrBV0W6_1(.din(n1272),.dout(w_dff_B_rYsrBV0W6_1),.clk(gclk));
	jdff dff_B_e8li2tLE4_1(.din(w_dff_B_rYsrBV0W6_1),.dout(w_dff_B_e8li2tLE4_1),.clk(gclk));
	jdff dff_B_5urLXsyC3_0(.din(n1333),.dout(w_dff_B_5urLXsyC3_0),.clk(gclk));
	jdff dff_B_G1whR9533_1(.din(n1345),.dout(w_dff_B_G1whR9533_1),.clk(gclk));
	jdff dff_B_yt8yq8iV8_1(.din(w_dff_B_G1whR9533_1),.dout(w_dff_B_yt8yq8iV8_1),.clk(gclk));
	jdff dff_B_ckbM7ytb5_0(.din(n1370),.dout(w_dff_B_ckbM7ytb5_0),.clk(gclk));
	jdff dff_B_35ZYj0rt8_1(.din(n1381),.dout(w_dff_B_35ZYj0rt8_1),.clk(gclk));
	jdff dff_B_4hGgm3Et5_1(.din(w_dff_B_35ZYj0rt8_1),.dout(w_dff_B_4hGgm3Et5_1),.clk(gclk));
	jdff dff_B_lMbt7F9W4_0(.din(n1406),.dout(w_dff_B_lMbt7F9W4_0),.clk(gclk));
	jdff dff_B_XDdD7kux4_1(.din(n1418),.dout(w_dff_B_XDdD7kux4_1),.clk(gclk));
	jdff dff_B_koWa50FX4_1(.din(w_dff_B_XDdD7kux4_1),.dout(w_dff_B_koWa50FX4_1),.clk(gclk));
	jdff dff_B_qygv1SxQ7_0(.din(n1443),.dout(w_dff_B_qygv1SxQ7_0),.clk(gclk));
	jdff dff_B_HMAOWoZm1_1(.din(n1454),.dout(w_dff_B_HMAOWoZm1_1),.clk(gclk));
	jdff dff_B_emjTCb4j0_1(.din(w_dff_B_HMAOWoZm1_1),.dout(w_dff_B_emjTCb4j0_1),.clk(gclk));
	jdff dff_B_i5x16gKI7_0(.din(n1479),.dout(w_dff_B_i5x16gKI7_0),.clk(gclk));
	jdff dff_B_VchOax7E1_1(.din(n1491),.dout(w_dff_B_VchOax7E1_1),.clk(gclk));
	jdff dff_B_1dMdFzNe2_1(.din(w_dff_B_VchOax7E1_1),.dout(w_dff_B_1dMdFzNe2_1),.clk(gclk));
	jdff dff_B_F4EsfGDJ5_0(.din(n1516),.dout(w_dff_B_F4EsfGDJ5_0),.clk(gclk));
	jdff dff_B_uBXblJmV0_1(.din(n1527),.dout(w_dff_B_uBXblJmV0_1),.clk(gclk));
	jdff dff_B_MXNCDc511_1(.din(w_dff_B_uBXblJmV0_1),.dout(w_dff_B_MXNCDc511_1),.clk(gclk));
	jdff dff_B_c0oDU8DR9_0(.din(n1552),.dout(w_dff_B_c0oDU8DR9_0),.clk(gclk));
	jdff dff_B_CMZG07on5_1(.din(n1564),.dout(w_dff_B_CMZG07on5_1),.clk(gclk));
	jdff dff_B_oaC8QtX88_1(.din(w_dff_B_CMZG07on5_1),.dout(w_dff_B_oaC8QtX88_1),.clk(gclk));
	jdff dff_B_1GbEw4ra1_0(.din(n1589),.dout(w_dff_B_1GbEw4ra1_0),.clk(gclk));
	jdff dff_B_J8H21Ve13_1(.din(n1600),.dout(w_dff_B_J8H21Ve13_1),.clk(gclk));
	jdff dff_B_zMcDdjhX8_1(.din(w_dff_B_J8H21Ve13_1),.dout(w_dff_B_zMcDdjhX8_1),.clk(gclk));
	jdff dff_B_nrM5oNz77_0(.din(n1625),.dout(w_dff_B_nrM5oNz77_0),.clk(gclk));
	jdff dff_B_xentm9ut9_1(.din(n1637),.dout(w_dff_B_xentm9ut9_1),.clk(gclk));
	jdff dff_B_qvsR5x1d9_1(.din(w_dff_B_xentm9ut9_1),.dout(w_dff_B_qvsR5x1d9_1),.clk(gclk));
	jdff dff_B_9vGQxAeC7_0(.din(n1662),.dout(w_dff_B_9vGQxAeC7_0),.clk(gclk));
	jdff dff_B_116dGzVJ3_1(.din(n1673),.dout(w_dff_B_116dGzVJ3_1),.clk(gclk));
	jdff dff_B_NPGtS0aV6_1(.din(w_dff_B_116dGzVJ3_1),.dout(w_dff_B_NPGtS0aV6_1),.clk(gclk));
	jdff dff_B_8IFA9uxn4_0(.din(n1698),.dout(w_dff_B_8IFA9uxn4_0),.clk(gclk));
	jdff dff_B_ecb1o3A97_1(.din(n1710),.dout(w_dff_B_ecb1o3A97_1),.clk(gclk));
	jdff dff_B_LLMoJvwo6_1(.din(w_dff_B_ecb1o3A97_1),.dout(w_dff_B_LLMoJvwo6_1),.clk(gclk));
	jdff dff_B_nuqFSaDm4_0(.din(n1735),.dout(w_dff_B_nuqFSaDm4_0),.clk(gclk));
	jdff dff_B_9ymwhC0x0_1(.din(n1746),.dout(w_dff_B_9ymwhC0x0_1),.clk(gclk));
	jdff dff_B_robiVxRf4_1(.din(w_dff_B_9ymwhC0x0_1),.dout(w_dff_B_robiVxRf4_1),.clk(gclk));
	jdff dff_B_OGeIt0NV8_0(.din(n1771),.dout(w_dff_B_OGeIt0NV8_0),.clk(gclk));
	jdff dff_B_iE2eMepW7_1(.din(n1783),.dout(w_dff_B_iE2eMepW7_1),.clk(gclk));
	jdff dff_B_cP0exCf09_1(.din(w_dff_B_iE2eMepW7_1),.dout(w_dff_B_cP0exCf09_1),.clk(gclk));
	jdff dff_B_g96jNHdJ1_0(.din(n1808),.dout(w_dff_B_g96jNHdJ1_0),.clk(gclk));
	jdff dff_B_dBor2d8J6_1(.din(n1819),.dout(w_dff_B_dBor2d8J6_1),.clk(gclk));
	jdff dff_B_ETLDoBFx5_1(.din(w_dff_B_dBor2d8J6_1),.dout(w_dff_B_ETLDoBFx5_1),.clk(gclk));
	jdff dff_B_h1n7C7xB6_0(.din(n1844),.dout(w_dff_B_h1n7C7xB6_0),.clk(gclk));
	jdff dff_B_bimxITUi8_1(.din(n1856),.dout(w_dff_B_bimxITUi8_1),.clk(gclk));
	jdff dff_B_55Edj9Zy7_1(.din(w_dff_B_bimxITUi8_1),.dout(w_dff_B_55Edj9Zy7_1),.clk(gclk));
	jdff dff_B_NmnoyRaM2_0(.din(n1881),.dout(w_dff_B_NmnoyRaM2_0),.clk(gclk));
	jdff dff_B_zNZVTUNb4_1(.din(n1892),.dout(w_dff_B_zNZVTUNb4_1),.clk(gclk));
	jdff dff_B_2a5xp3cf3_1(.din(w_dff_B_zNZVTUNb4_1),.dout(w_dff_B_2a5xp3cf3_1),.clk(gclk));
	jdff dff_B_m1xLLlKS6_0(.din(n1917),.dout(w_dff_B_m1xLLlKS6_0),.clk(gclk));
	jdff dff_B_gs2vDvNb3_1(.din(n1929),.dout(w_dff_B_gs2vDvNb3_1),.clk(gclk));
	jdff dff_B_Mfbpq3wo7_1(.din(w_dff_B_gs2vDvNb3_1),.dout(w_dff_B_Mfbpq3wo7_1),.clk(gclk));
	jdff dff_B_BVk4GIky4_0(.din(n1954),.dout(w_dff_B_BVk4GIky4_0),.clk(gclk));
	jdff dff_B_bLoygNGB6_1(.din(n1965),.dout(w_dff_B_bLoygNGB6_1),.clk(gclk));
	jdff dff_B_hOzIDkh54_1(.din(w_dff_B_bLoygNGB6_1),.dout(w_dff_B_hOzIDkh54_1),.clk(gclk));
	jdff dff_B_fhJ1mx9l9_0(.din(n1990),.dout(w_dff_B_fhJ1mx9l9_0),.clk(gclk));
	jdff dff_B_zlxKaspI7_1(.din(n2002),.dout(w_dff_B_zlxKaspI7_1),.clk(gclk));
	jdff dff_B_xuIIATgQ1_1(.din(w_dff_B_zlxKaspI7_1),.dout(w_dff_B_xuIIATgQ1_1),.clk(gclk));
	jdff dff_B_SZs8Qcod0_0(.din(n2027),.dout(w_dff_B_SZs8Qcod0_0),.clk(gclk));
	jdff dff_B_PYWeaYGl5_1(.din(n2038),.dout(w_dff_B_PYWeaYGl5_1),.clk(gclk));
	jdff dff_B_KLVuGhgh7_1(.din(w_dff_B_PYWeaYGl5_1),.dout(w_dff_B_KLVuGhgh7_1),.clk(gclk));
	jdff dff_B_enD4tXYE6_0(.din(n2063),.dout(w_dff_B_enD4tXYE6_0),.clk(gclk));
	jdff dff_B_hCq4zkgr3_1(.din(n2075),.dout(w_dff_B_hCq4zkgr3_1),.clk(gclk));
	jdff dff_B_UhGdGDuw2_1(.din(w_dff_B_hCq4zkgr3_1),.dout(w_dff_B_UhGdGDuw2_1),.clk(gclk));
	jdff dff_B_Sbji6ZfD0_0(.din(n2100),.dout(w_dff_B_Sbji6ZfD0_0),.clk(gclk));
	jdff dff_B_j9l6F43z2_1(.din(n2111),.dout(w_dff_B_j9l6F43z2_1),.clk(gclk));
	jdff dff_B_PRxlyw9O6_1(.din(w_dff_B_j9l6F43z2_1),.dout(w_dff_B_PRxlyw9O6_1),.clk(gclk));
	jdff dff_B_OcNBDkyx2_0(.din(n2136),.dout(w_dff_B_OcNBDkyx2_0),.clk(gclk));
	jdff dff_B_EFRg9bZf6_1(.din(n2148),.dout(w_dff_B_EFRg9bZf6_1),.clk(gclk));
	jdff dff_B_qCuGtxRb1_1(.din(w_dff_B_EFRg9bZf6_1),.dout(w_dff_B_qCuGtxRb1_1),.clk(gclk));
	jdff dff_B_o8z0a3BH8_0(.din(n2173),.dout(w_dff_B_o8z0a3BH8_0),.clk(gclk));
	jdff dff_B_Vvjm6PZZ6_1(.din(n2184),.dout(w_dff_B_Vvjm6PZZ6_1),.clk(gclk));
	jdff dff_B_ipvPNgWN6_1(.din(w_dff_B_Vvjm6PZZ6_1),.dout(w_dff_B_ipvPNgWN6_1),.clk(gclk));
	jdff dff_B_IfHCHb0m5_0(.din(n2209),.dout(w_dff_B_IfHCHb0m5_0),.clk(gclk));
	jdff dff_B_m0ZRsxqR5_1(.din(n2214),.dout(w_dff_B_m0ZRsxqR5_1),.clk(gclk));
	jdff dff_B_1rfsyViv6_1(.din(w_dff_B_m0ZRsxqR5_1),.dout(w_dff_B_1rfsyViv6_1),.clk(gclk));
	jdff dff_B_BoPmVl8N6_0(.din(n2218),.dout(w_dff_B_BoPmVl8N6_0),.clk(gclk));
	jdff dff_B_Qo4ZEKl62_1(.din(n2222),.dout(w_dff_B_Qo4ZEKl62_1),.clk(gclk));
	jdff dff_B_ShHJJsvM6_1(.din(w_dff_B_Qo4ZEKl62_1),.dout(w_dff_B_ShHJJsvM6_1),.clk(gclk));
	jdff dff_B_8LcbiD876_0(.din(n2226),.dout(w_dff_B_8LcbiD876_0),.clk(gclk));
	jdff dff_B_61TsfZBo0_1(.din(n2231),.dout(w_dff_B_61TsfZBo0_1),.clk(gclk));
	jdff dff_B_H5LQYE1i4_1(.din(w_dff_B_61TsfZBo0_1),.dout(w_dff_B_H5LQYE1i4_1),.clk(gclk));
	jdff dff_B_ZV0RQbIM7_0(.din(n2235),.dout(w_dff_B_ZV0RQbIM7_0),.clk(gclk));
	jdff dff_B_IN0A43qU2_1(.din(n2239),.dout(w_dff_B_IN0A43qU2_1),.clk(gclk));
	jdff dff_B_DNWcCaNq6_1(.din(w_dff_B_IN0A43qU2_1),.dout(w_dff_B_DNWcCaNq6_1),.clk(gclk));
	jdff dff_B_WKMYwIeP6_0(.din(n2243),.dout(w_dff_B_WKMYwIeP6_0),.clk(gclk));
	jdff dff_B_9Yjqugh99_1(.din(n2248),.dout(w_dff_B_9Yjqugh99_1),.clk(gclk));
	jdff dff_B_wMTGnKcB8_1(.din(w_dff_B_9Yjqugh99_1),.dout(w_dff_B_wMTGnKcB8_1),.clk(gclk));
	jdff dff_B_wQeft8uk8_0(.din(n2252),.dout(w_dff_B_wQeft8uk8_0),.clk(gclk));
	jdff dff_B_vsZalWtc9_1(.din(n2256),.dout(w_dff_B_vsZalWtc9_1),.clk(gclk));
	jdff dff_B_reajkNSh8_1(.din(w_dff_B_vsZalWtc9_1),.dout(w_dff_B_reajkNSh8_1),.clk(gclk));
	jdff dff_B_nGRQaI5L2_0(.din(n2260),.dout(w_dff_B_nGRQaI5L2_0),.clk(gclk));
	jdff dff_B_ZeRdUNCn5_1(.din(n2265),.dout(w_dff_B_ZeRdUNCn5_1),.clk(gclk));
	jdff dff_B_vqYPtKNk8_1(.din(w_dff_B_ZeRdUNCn5_1),.dout(w_dff_B_vqYPtKNk8_1),.clk(gclk));
	jdff dff_B_bAkFKoGi1_0(.din(n2269),.dout(w_dff_B_bAkFKoGi1_0),.clk(gclk));
	jdff dff_B_mD3g0jyP8_1(.din(n2273),.dout(w_dff_B_mD3g0jyP8_1),.clk(gclk));
	jdff dff_B_QbZh5GTu1_1(.din(w_dff_B_mD3g0jyP8_1),.dout(w_dff_B_QbZh5GTu1_1),.clk(gclk));
	jdff dff_B_bvqaMLGq4_0(.din(n2277),.dout(w_dff_B_bvqaMLGq4_0),.clk(gclk));
	jdff dff_B_dwolWk1u4_1(.din(n2282),.dout(w_dff_B_dwolWk1u4_1),.clk(gclk));
	jdff dff_B_aJJeIIHt4_1(.din(w_dff_B_dwolWk1u4_1),.dout(w_dff_B_aJJeIIHt4_1),.clk(gclk));
	jdff dff_B_CzywkDtF3_0(.din(n2286),.dout(w_dff_B_CzywkDtF3_0),.clk(gclk));
	jdff dff_B_3VkjLdoL6_1(.din(n2290),.dout(w_dff_B_3VkjLdoL6_1),.clk(gclk));
	jdff dff_B_VTYfoZ241_1(.din(w_dff_B_3VkjLdoL6_1),.dout(w_dff_B_VTYfoZ241_1),.clk(gclk));
	jdff dff_B_YX9OTQX74_0(.din(n2294),.dout(w_dff_B_YX9OTQX74_0),.clk(gclk));
	jdff dff_B_RKy8dYIb6_1(.din(n2299),.dout(w_dff_B_RKy8dYIb6_1),.clk(gclk));
	jdff dff_B_hCssqM0Q9_1(.din(w_dff_B_RKy8dYIb6_1),.dout(w_dff_B_hCssqM0Q9_1),.clk(gclk));
	jdff dff_B_rl1ZH6TR5_0(.din(n2303),.dout(w_dff_B_rl1ZH6TR5_0),.clk(gclk));
	jdff dff_B_dEI03NQy2_1(.din(n2307),.dout(w_dff_B_dEI03NQy2_1),.clk(gclk));
	jdff dff_B_qJOt6bhg1_1(.din(w_dff_B_dEI03NQy2_1),.dout(w_dff_B_qJOt6bhg1_1),.clk(gclk));
	jdff dff_B_dV3x719y6_0(.din(n2311),.dout(w_dff_B_dV3x719y6_0),.clk(gclk));
	jdff dff_B_4wh24KR08_1(.din(n2316),.dout(w_dff_B_4wh24KR08_1),.clk(gclk));
	jdff dff_B_G4Ih9Qr33_1(.din(w_dff_B_4wh24KR08_1),.dout(w_dff_B_G4Ih9Qr33_1),.clk(gclk));
	jdff dff_B_Oi4X5sPK9_0(.din(n2320),.dout(w_dff_B_Oi4X5sPK9_0),.clk(gclk));
	jdff dff_B_pn4CGLHa1_1(.din(n2324),.dout(w_dff_B_pn4CGLHa1_1),.clk(gclk));
	jdff dff_B_UQHrQaep4_1(.din(w_dff_B_pn4CGLHa1_1),.dout(w_dff_B_UQHrQaep4_1),.clk(gclk));
	jdff dff_B_bc3S7ENI2_0(.din(n2328),.dout(w_dff_B_bc3S7ENI2_0),.clk(gclk));
	jdff dff_B_KP72rsrz6_1(.din(n2333),.dout(w_dff_B_KP72rsrz6_1),.clk(gclk));
	jdff dff_B_7yGKMDYQ1_1(.din(w_dff_B_KP72rsrz6_1),.dout(w_dff_B_7yGKMDYQ1_1),.clk(gclk));
	jdff dff_B_wTfreXba5_0(.din(n2337),.dout(w_dff_B_wTfreXba5_0),.clk(gclk));
	jdff dff_B_euyAe64v7_1(.din(n2341),.dout(w_dff_B_euyAe64v7_1),.clk(gclk));
	jdff dff_B_xTJkLHWE4_1(.din(w_dff_B_euyAe64v7_1),.dout(w_dff_B_xTJkLHWE4_1),.clk(gclk));
	jdff dff_B_Xvu7oEBw8_0(.din(n2345),.dout(w_dff_B_Xvu7oEBw8_0),.clk(gclk));
	jdff dff_B_yYkEEkM38_1(.din(n2350),.dout(w_dff_B_yYkEEkM38_1),.clk(gclk));
	jdff dff_B_WHlDTliR9_1(.din(w_dff_B_yYkEEkM38_1),.dout(w_dff_B_WHlDTliR9_1),.clk(gclk));
	jdff dff_B_Bh0cWlsK3_0(.din(n2354),.dout(w_dff_B_Bh0cWlsK3_0),.clk(gclk));
	jdff dff_B_6a8xIgi53_1(.din(n2358),.dout(w_dff_B_6a8xIgi53_1),.clk(gclk));
	jdff dff_B_2kENvoBC8_1(.din(w_dff_B_6a8xIgi53_1),.dout(w_dff_B_2kENvoBC8_1),.clk(gclk));
	jdff dff_B_0uemW6GM9_0(.din(n2362),.dout(w_dff_B_0uemW6GM9_0),.clk(gclk));
	jdff dff_B_Y5BvixUE0_1(.din(n2367),.dout(w_dff_B_Y5BvixUE0_1),.clk(gclk));
	jdff dff_B_8SRP66dE1_1(.din(w_dff_B_Y5BvixUE0_1),.dout(w_dff_B_8SRP66dE1_1),.clk(gclk));
	jdff dff_B_GNedNEEq9_0(.din(n2371),.dout(w_dff_B_GNedNEEq9_0),.clk(gclk));
	jdff dff_B_uYRKYk1g1_1(.din(n2375),.dout(w_dff_B_uYRKYk1g1_1),.clk(gclk));
	jdff dff_B_eD6zHKXZ0_1(.din(w_dff_B_uYRKYk1g1_1),.dout(w_dff_B_eD6zHKXZ0_1),.clk(gclk));
	jdff dff_B_McwzmPqr1_0(.din(n2379),.dout(w_dff_B_McwzmPqr1_0),.clk(gclk));
	jdff dff_B_uoF5tk2m6_1(.din(n2384),.dout(w_dff_B_uoF5tk2m6_1),.clk(gclk));
	jdff dff_B_h3eJu9OU0_1(.din(w_dff_B_uoF5tk2m6_1),.dout(w_dff_B_h3eJu9OU0_1),.clk(gclk));
	jdff dff_B_u47osZBz0_0(.din(n2388),.dout(w_dff_B_u47osZBz0_0),.clk(gclk));
	jdff dff_B_Q4JjspNz1_1(.din(n2392),.dout(w_dff_B_Q4JjspNz1_1),.clk(gclk));
	jdff dff_B_ywtVITPN8_1(.din(w_dff_B_Q4JjspNz1_1),.dout(w_dff_B_ywtVITPN8_1),.clk(gclk));
	jdff dff_B_oYfAcDzV7_0(.din(n2396),.dout(w_dff_B_oYfAcDzV7_0),.clk(gclk));
	jdff dff_B_rHT2H57k2_1(.din(n2401),.dout(w_dff_B_rHT2H57k2_1),.clk(gclk));
	jdff dff_B_otiiGruG4_1(.din(w_dff_B_rHT2H57k2_1),.dout(w_dff_B_otiiGruG4_1),.clk(gclk));
	jdff dff_B_rGaC2c9d4_0(.din(n2405),.dout(w_dff_B_rGaC2c9d4_0),.clk(gclk));
	jdff dff_B_W01oYgIo0_1(.din(n2409),.dout(w_dff_B_W01oYgIo0_1),.clk(gclk));
	jdff dff_B_6L9GTXRb7_1(.din(w_dff_B_W01oYgIo0_1),.dout(w_dff_B_6L9GTXRb7_1),.clk(gclk));
	jdff dff_B_SqgF1FXp2_0(.din(n2413),.dout(w_dff_B_SqgF1FXp2_0),.clk(gclk));
	jdff dff_B_zcrvu5Ei2_1(.din(n2418),.dout(w_dff_B_zcrvu5Ei2_1),.clk(gclk));
	jdff dff_B_uHPHRthA7_1(.din(w_dff_B_zcrvu5Ei2_1),.dout(w_dff_B_uHPHRthA7_1),.clk(gclk));
	jdff dff_B_rkzRbhOh1_0(.din(n2422),.dout(w_dff_B_rkzRbhOh1_0),.clk(gclk));
	jdff dff_B_6bzhAcri5_1(.din(n2426),.dout(w_dff_B_6bzhAcri5_1),.clk(gclk));
	jdff dff_B_99mKSXMI6_1(.din(w_dff_B_6bzhAcri5_1),.dout(w_dff_B_99mKSXMI6_1),.clk(gclk));
	jdff dff_B_dk5lNsOw9_0(.din(n2430),.dout(w_dff_B_dk5lNsOw9_0),.clk(gclk));
	jdff dff_B_aJNLwn6g4_1(.din(n2435),.dout(w_dff_B_aJNLwn6g4_1),.clk(gclk));
	jdff dff_B_liuz3nrk5_1(.din(w_dff_B_aJNLwn6g4_1),.dout(w_dff_B_liuz3nrk5_1),.clk(gclk));
	jdff dff_B_H5CDb6oE6_0(.din(n2439),.dout(w_dff_B_H5CDb6oE6_0),.clk(gclk));
	jdff dff_B_Hb9wmUcB0_1(.din(n2443),.dout(w_dff_B_Hb9wmUcB0_1),.clk(gclk));
	jdff dff_B_KAogdi844_1(.din(w_dff_B_Hb9wmUcB0_1),.dout(w_dff_B_KAogdi844_1),.clk(gclk));
	jdff dff_B_SGLp9wMj4_0(.din(n2447),.dout(w_dff_B_SGLp9wMj4_0),.clk(gclk));
	jdff dff_B_GHCPb6rq3_1(.din(n2452),.dout(w_dff_B_GHCPb6rq3_1),.clk(gclk));
	jdff dff_B_DnS9XDKT8_1(.din(w_dff_B_GHCPb6rq3_1),.dout(w_dff_B_DnS9XDKT8_1),.clk(gclk));
	jdff dff_B_M6qUBrYh2_0(.din(n2456),.dout(w_dff_B_M6qUBrYh2_0),.clk(gclk));
	jdff dff_B_DQwxqxQg4_1(.din(n2460),.dout(w_dff_B_DQwxqxQg4_1),.clk(gclk));
	jdff dff_B_MG0suzb56_1(.din(w_dff_B_DQwxqxQg4_1),.dout(w_dff_B_MG0suzb56_1),.clk(gclk));
	jdff dff_B_RgGRMQHE6_0(.din(n2464),.dout(w_dff_B_RgGRMQHE6_0),.clk(gclk));
	jdff dff_B_kJ3dij4h6_1(.din(n2469),.dout(w_dff_B_kJ3dij4h6_1),.clk(gclk));
	jdff dff_B_9qAu6CEv6_1(.din(w_dff_B_kJ3dij4h6_1),.dout(w_dff_B_9qAu6CEv6_1),.clk(gclk));
	jdff dff_B_lNX9XknG9_0(.din(n2473),.dout(w_dff_B_lNX9XknG9_0),.clk(gclk));
	jdff dff_B_uOv1uSkF3_1(.din(n2477),.dout(w_dff_B_uOv1uSkF3_1),.clk(gclk));
	jdff dff_B_D9FffPJm6_1(.din(w_dff_B_uOv1uSkF3_1),.dout(w_dff_B_D9FffPJm6_1),.clk(gclk));
	jdff dff_B_q2S1c17p8_0(.din(n2481),.dout(w_dff_B_q2S1c17p8_0),.clk(gclk));
	jdff dff_B_rjprWWua0_1(.din(n2486),.dout(w_dff_B_rjprWWua0_1),.clk(gclk));
	jdff dff_B_yVPVbjPP6_1(.din(w_dff_B_rjprWWua0_1),.dout(w_dff_B_yVPVbjPP6_1),.clk(gclk));
	jdff dff_B_9iVsnI3Y0_0(.din(n2490),.dout(w_dff_B_9iVsnI3Y0_0),.clk(gclk));
	jdff dff_B_Ho3L4MC88_1(.din(n2494),.dout(w_dff_B_Ho3L4MC88_1),.clk(gclk));
	jdff dff_B_a3CGe7202_1(.din(w_dff_B_Ho3L4MC88_1),.dout(w_dff_B_a3CGe7202_1),.clk(gclk));
	jdff dff_B_bTy0068r1_0(.din(n2498),.dout(w_dff_B_bTy0068r1_0),.clk(gclk));
	jdff dff_B_PjliAp9l8_1(.din(n2503),.dout(w_dff_B_PjliAp9l8_1),.clk(gclk));
	jdff dff_B_19lEeWUB7_1(.din(w_dff_B_PjliAp9l8_1),.dout(w_dff_B_19lEeWUB7_1),.clk(gclk));
	jdff dff_B_7kVOx8kZ8_0(.din(n2507),.dout(w_dff_B_7kVOx8kZ8_0),.clk(gclk));
	jdff dff_B_qmiGF2fS5_1(.din(n2511),.dout(w_dff_B_qmiGF2fS5_1),.clk(gclk));
	jdff dff_B_7HQfPZQp1_1(.din(w_dff_B_qmiGF2fS5_1),.dout(w_dff_B_7HQfPZQp1_1),.clk(gclk));
	jdff dff_B_boPyw8vw4_0(.din(n2515),.dout(w_dff_B_boPyw8vw4_0),.clk(gclk));
	jdff dff_B_YHhQGkIh3_1(.din(n2520),.dout(w_dff_B_YHhQGkIh3_1),.clk(gclk));
	jdff dff_B_ky9JnIJa0_1(.din(w_dff_B_YHhQGkIh3_1),.dout(w_dff_B_ky9JnIJa0_1),.clk(gclk));
	jdff dff_B_YFkbXwkf8_0(.din(n2524),.dout(w_dff_B_YFkbXwkf8_0),.clk(gclk));
	jdff dff_B_8PGIHgI10_1(.din(n2528),.dout(w_dff_B_8PGIHgI10_1),.clk(gclk));
	jdff dff_B_FwE6F5NN2_1(.din(w_dff_B_8PGIHgI10_1),.dout(w_dff_B_FwE6F5NN2_1),.clk(gclk));
	jdff dff_B_9obNFDpn5_0(.din(n2532),.dout(w_dff_B_9obNFDpn5_0),.clk(gclk));
	jdff dff_B_muxmvvbB9_1(.din(n2537),.dout(w_dff_B_muxmvvbB9_1),.clk(gclk));
	jdff dff_B_4eITFKR93_1(.din(w_dff_B_muxmvvbB9_1),.dout(w_dff_B_4eITFKR93_1),.clk(gclk));
	jdff dff_B_YdezcyHU5_0(.din(n2541),.dout(w_dff_B_YdezcyHU5_0),.clk(gclk));
	jdff dff_B_Fjv5O2Ty2_1(.din(n2545),.dout(w_dff_B_Fjv5O2Ty2_1),.clk(gclk));
	jdff dff_B_f6wrL0AW5_1(.din(w_dff_B_Fjv5O2Ty2_1),.dout(w_dff_B_f6wrL0AW5_1),.clk(gclk));
	jdff dff_B_0hEDWuI26_0(.din(n2549),.dout(w_dff_B_0hEDWuI26_0),.clk(gclk));
	jdff dff_B_jM0CcFoY3_1(.din(n2554),.dout(w_dff_B_jM0CcFoY3_1),.clk(gclk));
	jdff dff_B_0Z3CSdIH1_1(.din(w_dff_B_jM0CcFoY3_1),.dout(w_dff_B_0Z3CSdIH1_1),.clk(gclk));
	jdff dff_B_qB6dFw1e2_0(.din(n2558),.dout(w_dff_B_qB6dFw1e2_0),.clk(gclk));
	jdff dff_B_H34hZ62M9_1(.din(n2562),.dout(w_dff_B_H34hZ62M9_1),.clk(gclk));
	jdff dff_B_f4xDkURy7_1(.din(w_dff_B_H34hZ62M9_1),.dout(w_dff_B_f4xDkURy7_1),.clk(gclk));
	jdff dff_B_u3F8t7vU1_0(.din(n2566),.dout(w_dff_B_u3F8t7vU1_0),.clk(gclk));
	jdff dff_B_1MNqUUdQ1_1(.din(n2571),.dout(w_dff_B_1MNqUUdQ1_1),.clk(gclk));
	jdff dff_B_OQ4nf9FB4_1(.din(w_dff_B_1MNqUUdQ1_1),.dout(w_dff_B_OQ4nf9FB4_1),.clk(gclk));
	jdff dff_B_huflLVnU8_0(.din(n2575),.dout(w_dff_B_huflLVnU8_0),.clk(gclk));
	jdff dff_B_BrGOasGm4_1(.din(n2579),.dout(w_dff_B_BrGOasGm4_1),.clk(gclk));
	jdff dff_B_N2r3icPs2_1(.din(w_dff_B_BrGOasGm4_1),.dout(w_dff_B_N2r3icPs2_1),.clk(gclk));
	jdff dff_B_X8hTW4sa2_0(.din(n2583),.dout(w_dff_B_X8hTW4sa2_0),.clk(gclk));
	jdff dff_B_QbSsgr8h7_1(.din(n2588),.dout(w_dff_B_QbSsgr8h7_1),.clk(gclk));
	jdff dff_B_nr95JRAm8_1(.din(w_dff_B_QbSsgr8h7_1),.dout(w_dff_B_nr95JRAm8_1),.clk(gclk));
	jdff dff_B_aEdf5wZc7_0(.din(n2592),.dout(w_dff_B_aEdf5wZc7_0),.clk(gclk));
	jdff dff_B_zI2Kpgg59_1(.din(n2596),.dout(w_dff_B_zI2Kpgg59_1),.clk(gclk));
	jdff dff_B_nkiDrsDo7_1(.din(w_dff_B_zI2Kpgg59_1),.dout(w_dff_B_nkiDrsDo7_1),.clk(gclk));
	jdff dff_B_C34EYOny8_0(.din(n2600),.dout(w_dff_B_C34EYOny8_0),.clk(gclk));
	jdff dff_B_z59wLket6_1(.din(n2605),.dout(w_dff_B_z59wLket6_1),.clk(gclk));
	jdff dff_B_b7uSIuaZ4_1(.din(w_dff_B_z59wLket6_1),.dout(w_dff_B_b7uSIuaZ4_1),.clk(gclk));
	jdff dff_B_YWRYZVvo7_0(.din(n2609),.dout(w_dff_B_YWRYZVvo7_0),.clk(gclk));
	jdff dff_B_rZQte5bu0_1(.din(n2613),.dout(w_dff_B_rZQte5bu0_1),.clk(gclk));
	jdff dff_B_CrXB06rb5_1(.din(w_dff_B_rZQte5bu0_1),.dout(w_dff_B_CrXB06rb5_1),.clk(gclk));
	jdff dff_B_496Qayul4_0(.din(n2617),.dout(w_dff_B_496Qayul4_0),.clk(gclk));
	jdff dff_B_TbgNN2S95_1(.din(n2622),.dout(w_dff_B_TbgNN2S95_1),.clk(gclk));
	jdff dff_B_V9UeSrPZ8_1(.din(w_dff_B_TbgNN2S95_1),.dout(w_dff_B_V9UeSrPZ8_1),.clk(gclk));
	jdff dff_B_gh9Bjk4K5_0(.din(n2626),.dout(w_dff_B_gh9Bjk4K5_0),.clk(gclk));
	jdff dff_B_3X0mNpgI5_1(.din(n2630),.dout(w_dff_B_3X0mNpgI5_1),.clk(gclk));
	jdff dff_B_uj3d5Aa12_1(.din(w_dff_B_3X0mNpgI5_1),.dout(w_dff_B_uj3d5Aa12_1),.clk(gclk));
	jdff dff_B_Onbv6u1X0_0(.din(n2634),.dout(w_dff_B_Onbv6u1X0_0),.clk(gclk));
	jdff dff_B_sr510KQA8_1(.din(n2639),.dout(w_dff_B_sr510KQA8_1),.clk(gclk));
	jdff dff_B_edIm3HEo0_1(.din(w_dff_B_sr510KQA8_1),.dout(w_dff_B_edIm3HEo0_1),.clk(gclk));
	jdff dff_B_ocQxDi7i4_0(.din(n2643),.dout(w_dff_B_ocQxDi7i4_0),.clk(gclk));
	jdff dff_B_CTjIjAr87_1(.din(n2647),.dout(w_dff_B_CTjIjAr87_1),.clk(gclk));
	jdff dff_B_Sy8fXmtO9_1(.din(w_dff_B_CTjIjAr87_1),.dout(w_dff_B_Sy8fXmtO9_1),.clk(gclk));
	jdff dff_B_ZqWDHNKl8_0(.din(n2651),.dout(w_dff_B_ZqWDHNKl8_0),.clk(gclk));
	jdff dff_B_xoKU3Id01_1(.din(n2656),.dout(w_dff_B_xoKU3Id01_1),.clk(gclk));
	jdff dff_B_SBRBhiff0_1(.din(w_dff_B_xoKU3Id01_1),.dout(w_dff_B_SBRBhiff0_1),.clk(gclk));
	jdff dff_B_rW47TtDh5_0(.din(n2660),.dout(w_dff_B_rW47TtDh5_0),.clk(gclk));
	jdff dff_B_bfjtPOIV7_1(.din(n2664),.dout(w_dff_B_bfjtPOIV7_1),.clk(gclk));
	jdff dff_B_4prvR3SB9_1(.din(w_dff_B_bfjtPOIV7_1),.dout(w_dff_B_4prvR3SB9_1),.clk(gclk));
	jdff dff_B_ujybVo5m3_0(.din(n2668),.dout(w_dff_B_ujybVo5m3_0),.clk(gclk));
	jdff dff_B_T8PVOLJC4_1(.din(n2673),.dout(w_dff_B_T8PVOLJC4_1),.clk(gclk));
	jdff dff_B_nh3K4oM22_1(.din(w_dff_B_T8PVOLJC4_1),.dout(w_dff_B_nh3K4oM22_1),.clk(gclk));
	jdff dff_B_AJta4V6q0_0(.din(n2677),.dout(w_dff_B_AJta4V6q0_0),.clk(gclk));
	jdff dff_B_sZXkuFTi7_1(.din(n2681),.dout(w_dff_B_sZXkuFTi7_1),.clk(gclk));
	jdff dff_B_43izO5SG7_1(.din(w_dff_B_sZXkuFTi7_1),.dout(w_dff_B_43izO5SG7_1),.clk(gclk));
	jdff dff_B_x80yLBcc3_0(.din(n2685),.dout(w_dff_B_x80yLBcc3_0),.clk(gclk));
	jdff dff_B_KAgkIkQn7_1(.din(n2690),.dout(w_dff_B_KAgkIkQn7_1),.clk(gclk));
	jdff dff_B_UO0r7WtK8_1(.din(w_dff_B_KAgkIkQn7_1),.dout(w_dff_B_UO0r7WtK8_1),.clk(gclk));
	jdff dff_B_4o1boigc1_0(.din(n2694),.dout(w_dff_B_4o1boigc1_0),.clk(gclk));
	jdff dff_B_Ys0zWwiN3_1(.din(n2698),.dout(w_dff_B_Ys0zWwiN3_1),.clk(gclk));
	jdff dff_B_tFBmKSHU9_1(.din(w_dff_B_Ys0zWwiN3_1),.dout(w_dff_B_tFBmKSHU9_1),.clk(gclk));
	jdff dff_B_A0PnvmfU3_0(.din(n2702),.dout(w_dff_B_A0PnvmfU3_0),.clk(gclk));
	jdff dff_B_20SCvLSX5_1(.din(n2707),.dout(w_dff_B_20SCvLSX5_1),.clk(gclk));
	jdff dff_B_8tVKfkLJ8_1(.din(w_dff_B_20SCvLSX5_1),.dout(w_dff_B_8tVKfkLJ8_1),.clk(gclk));
	jdff dff_B_YxqWpnGO2_0(.din(n2711),.dout(w_dff_B_YxqWpnGO2_0),.clk(gclk));
	jdff dff_B_JeoVcAtz5_1(.din(n2715),.dout(w_dff_B_JeoVcAtz5_1),.clk(gclk));
	jdff dff_B_DbMsD6I55_1(.din(w_dff_B_JeoVcAtz5_1),.dout(w_dff_B_DbMsD6I55_1),.clk(gclk));
	jdff dff_B_0BpUHJ8f5_0(.din(n2719),.dout(w_dff_B_0BpUHJ8f5_0),.clk(gclk));
	jdff dff_B_sIRvNoS55_1(.din(n2724),.dout(w_dff_B_sIRvNoS55_1),.clk(gclk));
	jdff dff_B_wOKdUDwI7_1(.din(w_dff_B_sIRvNoS55_1),.dout(w_dff_B_wOKdUDwI7_1),.clk(gclk));
	jdff dff_B_jFPT1jCW9_0(.din(n2728),.dout(w_dff_B_jFPT1jCW9_0),.clk(gclk));
	jdff dff_B_gLUxUchn8_1(.din(n2732),.dout(w_dff_B_gLUxUchn8_1),.clk(gclk));
	jdff dff_B_TEUMczxJ9_1(.din(w_dff_B_gLUxUchn8_1),.dout(w_dff_B_TEUMczxJ9_1),.clk(gclk));
	jdff dff_B_3WWymGYL5_0(.din(n2736),.dout(w_dff_B_3WWymGYL5_0),.clk(gclk));
	jdff dff_B_AgREMfxR4_1(.din(n2741),.dout(w_dff_B_AgREMfxR4_1),.clk(gclk));
	jdff dff_B_kLVUkxdA1_1(.din(w_dff_B_AgREMfxR4_1),.dout(w_dff_B_kLVUkxdA1_1),.clk(gclk));
	jdff dff_B_iXl7YkEZ9_0(.din(n2745),.dout(w_dff_B_iXl7YkEZ9_0),.clk(gclk));
	jdff dff_B_X3cYN9Mx0_1(.din(n2749),.dout(w_dff_B_X3cYN9Mx0_1),.clk(gclk));
	jdff dff_B_4gZnAB7L0_1(.din(w_dff_B_X3cYN9Mx0_1),.dout(w_dff_B_4gZnAB7L0_1),.clk(gclk));
	jdff dff_B_JOnwcef08_0(.din(n2753),.dout(w_dff_B_JOnwcef08_0),.clk(gclk));
	jdff dff_B_FephHzNx3_1(.din(n2758),.dout(w_dff_B_FephHzNx3_1),.clk(gclk));
	jdff dff_B_feWNsbf75_1(.din(w_dff_B_FephHzNx3_1),.dout(w_dff_B_feWNsbf75_1),.clk(gclk));
	jdff dff_B_cjjRtxAq5_0(.din(n2762),.dout(w_dff_B_cjjRtxAq5_0),.clk(gclk));
	jdff dff_B_uhfGFFCT8_1(.din(n467),.dout(w_dff_B_uhfGFFCT8_1),.clk(gclk));
	jdff dff_B_3JQdqvgr9_1(.din(w_dff_B_uhfGFFCT8_1),.dout(w_dff_B_3JQdqvgr9_1),.clk(gclk));
	jdff dff_B_i4pJGpHe3_0(.din(n498),.dout(w_dff_B_i4pJGpHe3_0),.clk(gclk));
	jdff dff_B_focNT7rN2_1(.din(n555),.dout(w_dff_B_focNT7rN2_1),.clk(gclk));
	jdff dff_B_9yHQ4G319_1(.din(w_dff_B_focNT7rN2_1),.dout(w_dff_B_9yHQ4G319_1),.clk(gclk));
	jdff dff_B_J66uxfix0_0(.din(n586),.dout(w_dff_B_J66uxfix0_0),.clk(gclk));
	jdff dff_B_MKxh3gBh9_1(.din(n511),.dout(w_dff_B_MKxh3gBh9_1),.clk(gclk));
	jdff dff_B_wrKJCLHE2_1(.din(w_dff_B_MKxh3gBh9_1),.dout(w_dff_B_wrKJCLHE2_1),.clk(gclk));
	jdff dff_B_WaH1Qvu22_0(.din(n542),.dout(w_dff_B_WaH1Qvu22_0),.clk(gclk));
	jdff dff_B_kWkTLlgn2_1(.din(n374),.dout(w_dff_B_kWkTLlgn2_1),.clk(gclk));
	jdff dff_B_zEG94JNY7_1(.din(w_dff_B_kWkTLlgn2_1),.dout(w_dff_B_zEG94JNY7_1),.clk(gclk));
	jdff dff_B_YzMLCC1i0_0(.din(n405),.dout(w_dff_B_YzMLCC1i0_0),.clk(gclk));
	jdff dff_B_UZmCgTSI6_1(.din(n2766),.dout(w_dff_B_UZmCgTSI6_1),.clk(gclk));
	jdff dff_B_cZrHVwDG1_1(.din(w_dff_B_UZmCgTSI6_1),.dout(w_dff_B_cZrHVwDG1_1),.clk(gclk));
	jdff dff_B_9CCHJG3I8_0(.din(n2770),.dout(w_dff_B_9CCHJG3I8_0),.clk(gclk));
	jdff dff_B_VuxjLPID6_1(.din(n600),.dout(w_dff_B_VuxjLPID6_1),.clk(gclk));
	jdff dff_B_T9dm59OW2_1(.din(w_dff_B_VuxjLPID6_1),.dout(w_dff_B_T9dm59OW2_1),.clk(gclk));
	jdff dff_B_PoFkE5wX0_0(.din(n631),.dout(w_dff_B_PoFkE5wX0_0),.clk(gclk));
	jdff dff_B_xGeMO9BU0_1(.din(n329),.dout(w_dff_B_xGeMO9BU0_1),.clk(gclk));
	jdff dff_B_faRWqwxy6_1(.din(w_dff_B_xGeMO9BU0_1),.dout(w_dff_B_faRWqwxy6_1),.clk(gclk));
	jdff dff_B_TkhLCRu23_0(.din(n360),.dout(w_dff_B_TkhLCRu23_0),.clk(gclk));
	jdff dff_B_a0UUqY5s8_1(.din(n279),.dout(w_dff_B_a0UUqY5s8_1),.clk(gclk));
	jdff dff_B_ENIICq2y3_1(.din(w_dff_B_a0UUqY5s8_1),.dout(w_dff_B_ENIICq2y3_1),.clk(gclk));
	jdff dff_B_GF88rIeY2_0(.din(n314),.dout(w_dff_B_GF88rIeY2_0),.clk(gclk));
	jdff dff_B_IuTIilJs1_1(.din(n420),.dout(w_dff_B_IuTIilJs1_1),.clk(gclk));
	jdff dff_B_BFVo2AC79_1(.din(w_dff_B_IuTIilJs1_1),.dout(w_dff_B_BFVo2AC79_1),.clk(gclk));
	jdff dff_B_AsSN8oxv0_0(.din(n451),.dout(w_dff_B_AsSN8oxv0_0),.clk(gclk));
	jdff dff_B_2WZlsVjY4_1(.din(n2775),.dout(w_dff_B_2WZlsVjY4_1),.clk(gclk));
	jdff dff_B_T0GGtFnc1_1(.din(w_dff_B_2WZlsVjY4_1),.dout(w_dff_B_T0GGtFnc1_1),.clk(gclk));
	jdff dff_B_jeXu3sy45_0(.din(n2779),.dout(w_dff_B_jeXu3sy45_0),.clk(gclk));
	jdff dff_B_kkOZ5FN67_1(.din(n648),.dout(w_dff_B_kkOZ5FN67_1),.clk(gclk));
	jdff dff_B_5U4XzmXQ9_1(.din(w_dff_B_kkOZ5FN67_1),.dout(w_dff_B_5U4XzmXQ9_1),.clk(gclk));
	jdff dff_B_poR6M3NX3_0(.din(n679),.dout(w_dff_B_poR6M3NX3_0),.clk(gclk));
	jdff dff_B_FSunM1fL8_1(.din(n872),.dout(w_dff_B_FSunM1fL8_1),.clk(gclk));
	jdff dff_B_Mx9XTvKw1_1(.din(w_dff_B_FSunM1fL8_1),.dout(w_dff_B_Mx9XTvKw1_1),.clk(gclk));
	jdff dff_B_XJJ0p5Hv1_0(.din(n903),.dout(w_dff_B_XJJ0p5Hv1_0),.clk(gclk));
	jdff dff_B_kRocFKSE5_1(.din(n916),.dout(w_dff_B_kRocFKSE5_1),.clk(gclk));
	jdff dff_B_pD3SBYZu7_1(.din(w_dff_B_kRocFKSE5_1),.dout(w_dff_B_pD3SBYZu7_1),.clk(gclk));
	jdff dff_B_R3YJSblS2_0(.din(n947),.dout(w_dff_B_R3YJSblS2_0),.clk(gclk));
	jdff dff_B_UM9TQzFB4_1(.din(n828),.dout(w_dff_B_UM9TQzFB4_1),.clk(gclk));
	jdff dff_B_NPOXfZNT9_1(.din(w_dff_B_UM9TQzFB4_1),.dout(w_dff_B_NPOXfZNT9_1),.clk(gclk));
	jdff dff_B_kk7LeyAl5_0(.din(n859),.dout(w_dff_B_kk7LeyAl5_0),.clk(gclk));
	jdff dff_B_egJRPEu89_1(.din(n2783),.dout(w_dff_B_egJRPEu89_1),.clk(gclk));
	jdff dff_B_pWTH2BSY6_1(.din(w_dff_B_egJRPEu89_1),.dout(w_dff_B_pWTH2BSY6_1),.clk(gclk));
	jdff dff_B_MoX53rZY3_0(.din(n2787),.dout(w_dff_B_MoX53rZY3_0),.clk(gclk));
	jdff dff_B_dE1wqsEz3_1(.din(n781),.dout(w_dff_B_dE1wqsEz3_1),.clk(gclk));
	jdff dff_B_EhiM211Y3_1(.din(w_dff_B_dE1wqsEz3_1),.dout(w_dff_B_EhiM211Y3_1),.clk(gclk));
	jdff dff_B_rOHLQUyL7_0(.din(n812),.dout(w_dff_B_rOHLQUyL7_0),.clk(gclk));
	jdff dff_B_Dq3Q0i4O2_1(.din(n736),.dout(w_dff_B_Dq3Q0i4O2_1),.clk(gclk));
	jdff dff_B_HBaastiB7_1(.din(w_dff_B_Dq3Q0i4O2_1),.dout(w_dff_B_HBaastiB7_1),.clk(gclk));
	jdff dff_B_RbwjiVQc5_0(.din(n767),.dout(w_dff_B_RbwjiVQc5_0),.clk(gclk));
	jdff dff_B_YfL9hMuc0_1(.din(n692),.dout(w_dff_B_YfL9hMuc0_1),.clk(gclk));
	jdff dff_B_fvmWPNeu8_1(.din(w_dff_B_YfL9hMuc0_1),.dout(w_dff_B_fvmWPNeu8_1),.clk(gclk));
	jdff dff_B_56NlZhYE3_0(.din(n723),.dout(w_dff_B_56NlZhYE3_0),.clk(gclk));
	jdff dff_B_MIhQQiDJ8_1(.din(n961),.dout(w_dff_B_MIhQQiDJ8_1),.clk(gclk));
	jdff dff_B_n4s9MQBi8_1(.din(w_dff_B_MIhQQiDJ8_1),.dout(w_dff_B_n4s9MQBi8_1),.clk(gclk));
	jdff dff_B_Tp0JK1jz6_0(.din(n992),.dout(w_dff_B_Tp0JK1jz6_0),.clk(gclk));
	jdff dff_B_0j7GEJgP0_1(.din(n2792),.dout(w_dff_B_0j7GEJgP0_1),.clk(gclk));
	jdff dff_B_h6gd19k23_1(.din(w_dff_B_0j7GEJgP0_1),.dout(w_dff_B_h6gd19k23_1),.clk(gclk));
	jdff dff_B_YOJR5kVR6_0(.din(n2796),.dout(w_dff_B_YOJR5kVR6_0),.clk(gclk));
	jdff dff_B_UDDJjihN1_1(.din(n1107),.dout(w_dff_B_UDDJjihN1_1),.clk(gclk));
	jdff dff_B_CJe3LNGD1_1(.din(w_dff_B_UDDJjihN1_1),.dout(w_dff_B_CJe3LNGD1_1),.clk(gclk));
	jdff dff_B_YCE8fMWj4_0(.din(n1120),.dout(w_dff_B_YCE8fMWj4_0),.clk(gclk));
	jdff dff_B_cpHbBKmC5_1(.din(n1087),.dout(w_dff_B_cpHbBKmC5_1),.clk(gclk));
	jdff dff_B_ZhWqQhPZ3_1(.din(w_dff_B_cpHbBKmC5_1),.dout(w_dff_B_ZhWqQhPZ3_1),.clk(gclk));
	jdff dff_B_ZGWEitvM6_0(.din(n1100),.dout(w_dff_B_ZGWEitvM6_0),.clk(gclk));
	jdff dff_B_yRqUJEnE2_1(.din(n1148),.dout(w_dff_B_yRqUJEnE2_1),.clk(gclk));
	jdff dff_B_sQ1XAWmU2_1(.din(w_dff_B_yRqUJEnE2_1),.dout(w_dff_B_sQ1XAWmU2_1),.clk(gclk));
	jdff dff_B_aeg3cgRf4_0(.din(n1161),.dout(w_dff_B_aeg3cgRf4_0),.clk(gclk));
	jdff dff_B_iDyOIIGT5_1(.din(n1064),.dout(w_dff_B_iDyOIIGT5_1),.clk(gclk));
	jdff dff_B_oMk1KklB2_1(.din(w_dff_B_iDyOIIGT5_1),.dout(w_dff_B_oMk1KklB2_1),.clk(gclk));
	jdff dff_B_hh4D6Ws52_0(.din(n1077),.dout(w_dff_B_hh4D6Ws52_0),.clk(gclk));
	jdff dff_B_3iGzd9JX6_1(.din(n2800),.dout(w_dff_B_3iGzd9JX6_1),.clk(gclk));
	jdff dff_B_n9pUpmqm8_1(.din(w_dff_B_3iGzd9JX6_1),.dout(w_dff_B_n9pUpmqm8_1),.clk(gclk));
	jdff dff_B_qG7CcZVr6_0(.din(n2804),.dout(w_dff_B_qG7CcZVr6_0),.clk(gclk));
	jdff dff_B_6A2FPn0t3_1(.din(n1127),.dout(w_dff_B_6A2FPn0t3_1),.clk(gclk));
	jdff dff_B_gws8z3LA1_1(.din(w_dff_B_6A2FPn0t3_1),.dout(w_dff_B_gws8z3LA1_1),.clk(gclk));
	jdff dff_B_5ldzfQYi3_0(.din(n1140),.dout(w_dff_B_5ldzfQYi3_0),.clk(gclk));
	jdff dff_B_MaGlQa950_1(.din(n1043),.dout(w_dff_B_MaGlQa950_1),.clk(gclk));
	jdff dff_B_3KDdwdBk3_1(.din(w_dff_B_MaGlQa950_1),.dout(w_dff_B_3KDdwdBk3_1),.clk(gclk));
	jdff dff_B_xnBRSN2N3_0(.din(n1056),.dout(w_dff_B_xnBRSN2N3_0),.clk(gclk));
	jdff dff_B_djcKn61M3_1(.din(n1023),.dout(w_dff_B_djcKn61M3_1),.clk(gclk));
	jdff dff_B_wnQLWcq32_1(.din(w_dff_B_djcKn61M3_1),.dout(w_dff_B_wnQLWcq32_1),.clk(gclk));
	jdff dff_B_BlDVNLBK7_0(.din(n1036),.dout(w_dff_B_BlDVNLBK7_0),.clk(gclk));
	jdff dff_B_WOEkBFSe2_1(.din(n1003),.dout(w_dff_B_WOEkBFSe2_1),.clk(gclk));
	jdff dff_B_4OEclSdP1_1(.din(w_dff_B_WOEkBFSe2_1),.dout(w_dff_B_4OEclSdP1_1),.clk(gclk));
	jdff dff_B_vGLAXmG71_0(.din(n1016),.dout(w_dff_B_vGLAXmG71_0),.clk(gclk));
	jdff dff_B_9RJGWIrd7_1(.din(n2809),.dout(w_dff_B_9RJGWIrd7_1),.clk(gclk));
	jdff dff_B_XrRsKiC06_1(.din(w_dff_B_9RJGWIrd7_1),.dout(w_dff_B_XrRsKiC06_1),.clk(gclk));
	jdff dff_B_B3HjuQuU9_0(.din(n2813),.dout(w_dff_B_B3HjuQuU9_0),.clk(gclk));
	jdff dff_B_FZxU42WT4_1(.din(n1256),.dout(w_dff_B_FZxU42WT4_1),.clk(gclk));
	jdff dff_B_y7xezhI94_1(.din(w_dff_B_FZxU42WT4_1),.dout(w_dff_B_y7xezhI94_1),.clk(gclk));
	jdff dff_B_hGQAN2Ud3_0(.din(n1269),.dout(w_dff_B_hGQAN2Ud3_0),.clk(gclk));
	jdff dff_B_mUIeIU2P5_1(.din(n1276),.dout(w_dff_B_mUIeIU2P5_1),.clk(gclk));
	jdff dff_B_v6S0pnWU5_1(.din(w_dff_B_mUIeIU2P5_1),.dout(w_dff_B_v6S0pnWU5_1),.clk(gclk));
	jdff dff_B_bxZjKYFc1_0(.din(n1289),.dout(w_dff_B_bxZjKYFc1_0),.clk(gclk));
	jdff dff_B_hBgbUGtR7_1(.din(n1317),.dout(w_dff_B_hBgbUGtR7_1),.clk(gclk));
	jdff dff_B_6KHWH1Jh5_1(.din(w_dff_B_hBgbUGtR7_1),.dout(w_dff_B_6KHWH1Jh5_1),.clk(gclk));
	jdff dff_B_xB4q2Qjw2_0(.din(n1330),.dout(w_dff_B_xB4q2Qjw2_0),.clk(gclk));
	jdff dff_B_YUDdw4H56_1(.din(n1172),.dout(w_dff_B_YUDdw4H56_1),.clk(gclk));
	jdff dff_B_L4laJNFt4_1(.din(w_dff_B_YUDdw4H56_1),.dout(w_dff_B_L4laJNFt4_1),.clk(gclk));
	jdff dff_B_NyFPXIyr2_0(.din(n1185),.dout(w_dff_B_NyFPXIyr2_0),.clk(gclk));
	jdff dff_B_T1FtALzk3_1(.din(n2817),.dout(w_dff_B_T1FtALzk3_1),.clk(gclk));
	jdff dff_B_VMQQNRP08_1(.din(w_dff_B_T1FtALzk3_1),.dout(w_dff_B_VMQQNRP08_1),.clk(gclk));
	jdff dff_B_SOdTOQwU7_0(.din(n2821),.dout(w_dff_B_SOdTOQwU7_0),.clk(gclk));
	jdff dff_B_86vXx9XN1_1(.din(n1296),.dout(w_dff_B_86vXx9XN1_1),.clk(gclk));
	jdff dff_B_vvMFgqlf6_1(.din(w_dff_B_86vXx9XN1_1),.dout(w_dff_B_vvMFgqlf6_1),.clk(gclk));
	jdff dff_B_B2NxBOMf3_0(.din(n1309),.dout(w_dff_B_B2NxBOMf3_0),.clk(gclk));
	jdff dff_B_GxdybRXV1_1(.din(n1192),.dout(w_dff_B_GxdybRXV1_1),.clk(gclk));
	jdff dff_B_82FVcnT81_1(.din(w_dff_B_GxdybRXV1_1),.dout(w_dff_B_82FVcnT81_1),.clk(gclk));
	jdff dff_B_t5k4kQhB6_0(.din(n1205),.dout(w_dff_B_t5k4kQhB6_0),.clk(gclk));
	jdff dff_B_cBR00QJg3_1(.din(n1212),.dout(w_dff_B_cBR00QJg3_1),.clk(gclk));
	jdff dff_B_ycfnNlTi5_1(.din(w_dff_B_cBR00QJg3_1),.dout(w_dff_B_ycfnNlTi5_1),.clk(gclk));
	jdff dff_B_hZx5Rp366_0(.din(n1225),.dout(w_dff_B_hZx5Rp366_0),.clk(gclk));
	jdff dff_B_6ZMF23I40_1(.din(n1233),.dout(w_dff_B_6ZMF23I40_1),.clk(gclk));
	jdff dff_B_VGg8A4KJ8_1(.din(w_dff_B_6ZMF23I40_1),.dout(w_dff_B_VGg8A4KJ8_1),.clk(gclk));
	jdff dff_B_Qp7R6Ppv0_0(.din(n1246),.dout(w_dff_B_Qp7R6Ppv0_0),.clk(gclk));
	jdff dff_B_rBcQrI584_1(.din(n2826),.dout(w_dff_B_rBcQrI584_1),.clk(gclk));
	jdff dff_B_GEI0pHLe2_1(.din(w_dff_B_rBcQrI584_1),.dout(w_dff_B_GEI0pHLe2_1),.clk(gclk));
	jdff dff_B_7IMUWZDl2_0(.din(n2830),.dout(w_dff_B_7IMUWZDl2_0),.clk(gclk));
	jdff dff_B_9QCGOelP1_1(.din(n1399),.dout(w_dff_B_9QCGOelP1_1),.clk(gclk));
	jdff dff_B_bz9R4FL06_1(.din(w_dff_B_9QCGOelP1_1),.dout(w_dff_B_bz9R4FL06_1),.clk(gclk));
	jdff dff_B_1DoTDJze9_0(.din(n1403),.dout(w_dff_B_1DoTDJze9_0),.clk(gclk));
	jdff dff_B_tcxmG4DG5_1(.din(n1382),.dout(w_dff_B_tcxmG4DG5_1),.clk(gclk));
	jdff dff_B_StgGyzNM1_1(.din(w_dff_B_tcxmG4DG5_1),.dout(w_dff_B_StgGyzNM1_1),.clk(gclk));
	jdff dff_B_hknLRKEp8_0(.din(n1386),.dout(w_dff_B_hknLRKEp8_0),.clk(gclk));
	jdff dff_B_d95Y6bnw1_1(.din(n1338),.dout(w_dff_B_d95Y6bnw1_1),.clk(gclk));
	jdff dff_B_gfiTS28a2_1(.din(w_dff_B_d95Y6bnw1_1),.dout(w_dff_B_gfiTS28a2_1),.clk(gclk));
	jdff dff_B_1OEUfKzK8_0(.din(n1342),.dout(w_dff_B_1OEUfKzK8_0),.clk(gclk));
	jdff dff_B_gO2pJsJg3_1(.din(n1374),.dout(w_dff_B_gO2pJsJg3_1),.clk(gclk));
	jdff dff_B_EtA1Bwgh7_1(.din(w_dff_B_gO2pJsJg3_1),.dout(w_dff_B_EtA1Bwgh7_1),.clk(gclk));
	jdff dff_B_Yji0C1js9_0(.din(n1378),.dout(w_dff_B_Yji0C1js9_0),.clk(gclk));
	jdff dff_B_4bWQ8Y4U4_1(.din(n2834),.dout(w_dff_B_4bWQ8Y4U4_1),.clk(gclk));
	jdff dff_B_IEnkpo8q6_1(.din(w_dff_B_4bWQ8Y4U4_1),.dout(w_dff_B_IEnkpo8q6_1),.clk(gclk));
	jdff dff_B_IHsLOWpC2_0(.din(n2838),.dout(w_dff_B_IHsLOWpC2_0),.clk(gclk));
	jdff dff_B_Onbogkyx1_1(.din(n1363),.dout(w_dff_B_Onbogkyx1_1),.clk(gclk));
	jdff dff_B_DD4YCshY8_1(.din(w_dff_B_Onbogkyx1_1),.dout(w_dff_B_DD4YCshY8_1),.clk(gclk));
	jdff dff_B_RWQCZSD81_0(.din(n1367),.dout(w_dff_B_RWQCZSD81_0),.clk(gclk));
	jdff dff_B_kDPvPpoP4_1(.din(n1390),.dout(w_dff_B_kDPvPpoP4_1),.clk(gclk));
	jdff dff_B_wO6CPyKc2_1(.din(w_dff_B_kDPvPpoP4_1),.dout(w_dff_B_wO6CPyKc2_1),.clk(gclk));
	jdff dff_B_70rd1kZT3_0(.din(n1394),.dout(w_dff_B_70rd1kZT3_0),.clk(gclk));
	jdff dff_B_rzbj5T0z1_1(.din(n1346),.dout(w_dff_B_rzbj5T0z1_1),.clk(gclk));
	jdff dff_B_EMAK944C1_1(.din(w_dff_B_rzbj5T0z1_1),.dout(w_dff_B_EMAK944C1_1),.clk(gclk));
	jdff dff_B_PIEA6oQH3_0(.din(n1350),.dout(w_dff_B_PIEA6oQH3_0),.clk(gclk));
	jdff dff_B_IFtLjBZF6_1(.din(n1354),.dout(w_dff_B_IFtLjBZF6_1),.clk(gclk));
	jdff dff_B_Y9K3ClDR7_1(.din(w_dff_B_IFtLjBZF6_1),.dout(w_dff_B_Y9K3ClDR7_1),.clk(gclk));
	jdff dff_B_8BngNbgd0_0(.din(n1358),.dout(w_dff_B_8BngNbgd0_0),.clk(gclk));
	jdff dff_B_I7aht90O4_1(.din(n2843),.dout(w_dff_B_I7aht90O4_1),.clk(gclk));
	jdff dff_B_3wuBCOe82_1(.din(w_dff_B_I7aht90O4_1),.dout(w_dff_B_3wuBCOe82_1),.clk(gclk));
	jdff dff_B_mfvk1noa9_0(.din(n2847),.dout(w_dff_B_mfvk1noa9_0),.clk(gclk));
	jdff dff_B_98IgX14T0_1(.din(n1455),.dout(w_dff_B_98IgX14T0_1),.clk(gclk));
	jdff dff_B_O9cfa67M4_1(.din(w_dff_B_98IgX14T0_1),.dout(w_dff_B_O9cfa67M4_1),.clk(gclk));
	jdff dff_B_LuB7p5DQ9_0(.din(n1459),.dout(w_dff_B_LuB7p5DQ9_0),.clk(gclk));
	jdff dff_B_Djzz0kY27_1(.din(n1463),.dout(w_dff_B_Djzz0kY27_1),.clk(gclk));
	jdff dff_B_ObVd5VZ58_1(.din(w_dff_B_Djzz0kY27_1),.dout(w_dff_B_ObVd5VZ58_1),.clk(gclk));
	jdff dff_B_z89m836x9_0(.din(n1467),.dout(w_dff_B_z89m836x9_0),.clk(gclk));
	jdff dff_B_okhOeJHm0_1(.din(n1436),.dout(w_dff_B_okhOeJHm0_1),.clk(gclk));
	jdff dff_B_KrkdkH7l9_1(.din(w_dff_B_okhOeJHm0_1),.dout(w_dff_B_KrkdkH7l9_1),.clk(gclk));
	jdff dff_B_iymvmlfM2_0(.din(n1440),.dout(w_dff_B_iymvmlfM2_0),.clk(gclk));
	jdff dff_B_QmqB7p2U9_1(.din(n1447),.dout(w_dff_B_QmqB7p2U9_1),.clk(gclk));
	jdff dff_B_QwBaURrl5_1(.din(w_dff_B_QmqB7p2U9_1),.dout(w_dff_B_QwBaURrl5_1),.clk(gclk));
	jdff dff_B_D9fLjXBM7_0(.din(n1451),.dout(w_dff_B_D9fLjXBM7_0),.clk(gclk));
	jdff dff_B_1ZtuVlls5_1(.din(n2851),.dout(w_dff_B_1ZtuVlls5_1),.clk(gclk));
	jdff dff_B_FRrwnx3T2_1(.din(w_dff_B_1ZtuVlls5_1),.dout(w_dff_B_FRrwnx3T2_1),.clk(gclk));
	jdff dff_B_7Xuq5K5W5_0(.din(n2855),.dout(w_dff_B_7Xuq5K5W5_0),.clk(gclk));
	jdff dff_B_3k65QdRj2_1(.din(n1472),.dout(w_dff_B_3k65QdRj2_1),.clk(gclk));
	jdff dff_B_XnPkPJHe3_1(.din(w_dff_B_3k65QdRj2_1),.dout(w_dff_B_XnPkPJHe3_1),.clk(gclk));
	jdff dff_B_RAvhSOHM5_0(.din(n1476),.dout(w_dff_B_RAvhSOHM5_0),.clk(gclk));
	jdff dff_B_1pacFc5A9_1(.din(n1427),.dout(w_dff_B_1pacFc5A9_1),.clk(gclk));
	jdff dff_B_yogMl37H5_1(.din(w_dff_B_1pacFc5A9_1),.dout(w_dff_B_yogMl37H5_1),.clk(gclk));
	jdff dff_B_DqhQ5BMC9_0(.din(n1431),.dout(w_dff_B_DqhQ5BMC9_0),.clk(gclk));
	jdff dff_B_uet8h9lm8_1(.din(n1419),.dout(w_dff_B_uet8h9lm8_1),.clk(gclk));
	jdff dff_B_hozR8B1v3_1(.din(w_dff_B_uet8h9lm8_1),.dout(w_dff_B_hozR8B1v3_1),.clk(gclk));
	jdff dff_B_FQAQqQ3K2_0(.din(n1423),.dout(w_dff_B_FQAQqQ3K2_0),.clk(gclk));
	jdff dff_B_61j1RiBO5_1(.din(n1411),.dout(w_dff_B_61j1RiBO5_1),.clk(gclk));
	jdff dff_B_V651QdOo9_1(.din(w_dff_B_61j1RiBO5_1),.dout(w_dff_B_V651QdOo9_1),.clk(gclk));
	jdff dff_B_4FGpBViq2_0(.din(n1415),.dout(w_dff_B_4FGpBViq2_0),.clk(gclk));
	jdff dff_B_9fZ3rJLb9_1(.din(n2860),.dout(w_dff_B_9fZ3rJLb9_1),.clk(gclk));
	jdff dff_B_r38PTKb32_1(.din(w_dff_B_9fZ3rJLb9_1),.dout(w_dff_B_r38PTKb32_1),.clk(gclk));
	jdff dff_B_49MrkuEv1_0(.din(n2864),.dout(w_dff_B_49MrkuEv1_0),.clk(gclk));
	jdff dff_B_dswNJH0Q3_1(.din(n1520),.dout(w_dff_B_dswNJH0Q3_1),.clk(gclk));
	jdff dff_B_HZGcZQx65_1(.din(w_dff_B_dswNJH0Q3_1),.dout(w_dff_B_HZGcZQx65_1),.clk(gclk));
	jdff dff_B_HuZqe8R86_0(.din(n1524),.dout(w_dff_B_HuZqe8R86_0),.clk(gclk));
	jdff dff_B_5z6ntGRA1_1(.din(n1545),.dout(w_dff_B_5z6ntGRA1_1),.clk(gclk));
	jdff dff_B_LnFLsAV69_1(.din(w_dff_B_5z6ntGRA1_1),.dout(w_dff_B_LnFLsAV69_1),.clk(gclk));
	jdff dff_B_XQRJK8hI2_0(.din(n1549),.dout(w_dff_B_XQRJK8hI2_0),.clk(gclk));
	jdff dff_B_3YFfs46K3_1(.din(n1500),.dout(w_dff_B_3YFfs46K3_1),.clk(gclk));
	jdff dff_B_FMefJS5z4_1(.din(w_dff_B_3YFfs46K3_1),.dout(w_dff_B_FMefJS5z4_1),.clk(gclk));
	jdff dff_B_ldonzCFe9_0(.din(n1504),.dout(w_dff_B_ldonzCFe9_0),.clk(gclk));
	jdff dff_B_V5RqNucF7_1(.din(n1528),.dout(w_dff_B_V5RqNucF7_1),.clk(gclk));
	jdff dff_B_Y88xVshG7_1(.din(w_dff_B_V5RqNucF7_1),.dout(w_dff_B_Y88xVshG7_1),.clk(gclk));
	jdff dff_B_FHH2yJSp7_0(.din(n1532),.dout(w_dff_B_FHH2yJSp7_0),.clk(gclk));
	jdff dff_B_HrXKvA0r3_1(.din(n2868),.dout(w_dff_B_HrXKvA0r3_1),.clk(gclk));
	jdff dff_B_3p3FQbxZ2_1(.din(w_dff_B_HrXKvA0r3_1),.dout(w_dff_B_3p3FQbxZ2_1),.clk(gclk));
	jdff dff_B_FDc46lRH6_0(.din(n2872),.dout(w_dff_B_FDc46lRH6_0),.clk(gclk));
	jdff dff_B_QI6jOKro7_1(.din(n1484),.dout(w_dff_B_QI6jOKro7_1),.clk(gclk));
	jdff dff_B_CBcSyyyU8_1(.din(w_dff_B_QI6jOKro7_1),.dout(w_dff_B_CBcSyyyU8_1),.clk(gclk));
	jdff dff_B_JNJO4QOP3_0(.din(n1488),.dout(w_dff_B_JNJO4QOP3_0),.clk(gclk));
	jdff dff_B_q2uZc8Gj9_1(.din(n1536),.dout(w_dff_B_q2uZc8Gj9_1),.clk(gclk));
	jdff dff_B_qYzkE5Ne5_1(.din(w_dff_B_q2uZc8Gj9_1),.dout(w_dff_B_qYzkE5Ne5_1),.clk(gclk));
	jdff dff_B_7JX91FRK1_0(.din(n1540),.dout(w_dff_B_7JX91FRK1_0),.clk(gclk));
	jdff dff_B_pVLlfeWJ1_1(.din(n1492),.dout(w_dff_B_pVLlfeWJ1_1),.clk(gclk));
	jdff dff_B_JL4G19Qr8_1(.din(w_dff_B_pVLlfeWJ1_1),.dout(w_dff_B_JL4G19Qr8_1),.clk(gclk));
	jdff dff_B_yYHiuxfW3_0(.din(n1496),.dout(w_dff_B_yYHiuxfW3_0),.clk(gclk));
	jdff dff_B_6w4rnDi74_1(.din(n1509),.dout(w_dff_B_6w4rnDi74_1),.clk(gclk));
	jdff dff_B_QeKRpaxT3_1(.din(w_dff_B_6w4rnDi74_1),.dout(w_dff_B_QeKRpaxT3_1),.clk(gclk));
	jdff dff_B_KwAJ2y101_0(.din(n1513),.dout(w_dff_B_KwAJ2y101_0),.clk(gclk));
	jdff dff_B_hWACObTH0_1(.din(n2877),.dout(w_dff_B_hWACObTH0_1),.clk(gclk));
	jdff dff_B_ZHHldruu7_1(.din(w_dff_B_hWACObTH0_1),.dout(w_dff_B_ZHHldruu7_1),.clk(gclk));
	jdff dff_B_hTzDDnzK8_0(.din(n2881),.dout(w_dff_B_hTzDDnzK8_0),.clk(gclk));
	jdff dff_B_cnGtcmvV7_1(.din(n1601),.dout(w_dff_B_cnGtcmvV7_1),.clk(gclk));
	jdff dff_B_HugGMlsl5_1(.din(w_dff_B_cnGtcmvV7_1),.dout(w_dff_B_HugGMlsl5_1),.clk(gclk));
	jdff dff_B_yoRicxHq6_0(.din(n1605),.dout(w_dff_B_yoRicxHq6_0),.clk(gclk));
	jdff dff_B_Yp5MvGc20_1(.din(n1593),.dout(w_dff_B_Yp5MvGc20_1),.clk(gclk));
	jdff dff_B_fkSCvyox5_1(.din(w_dff_B_Yp5MvGc20_1),.dout(w_dff_B_fkSCvyox5_1),.clk(gclk));
	jdff dff_B_LderWme62_0(.din(n1597),.dout(w_dff_B_LderWme62_0),.clk(gclk));
	jdff dff_B_ql79bxwE5_1(.din(n1609),.dout(w_dff_B_ql79bxwE5_1),.clk(gclk));
	jdff dff_B_Dr5Rgvhi0_1(.din(w_dff_B_ql79bxwE5_1),.dout(w_dff_B_Dr5Rgvhi0_1),.clk(gclk));
	jdff dff_B_4lNWY1Cp4_0(.din(n1613),.dout(w_dff_B_4lNWY1Cp4_0),.clk(gclk));
	jdff dff_B_ZJ7t2wem9_1(.din(n1573),.dout(w_dff_B_ZJ7t2wem9_1),.clk(gclk));
	jdff dff_B_qU6FUjGM9_1(.din(w_dff_B_ZJ7t2wem9_1),.dout(w_dff_B_qU6FUjGM9_1),.clk(gclk));
	jdff dff_B_PjZlxOwU2_0(.din(n1577),.dout(w_dff_B_PjZlxOwU2_0),.clk(gclk));
	jdff dff_B_pcpEuBTO7_1(.din(n2885),.dout(w_dff_B_pcpEuBTO7_1),.clk(gclk));
	jdff dff_B_ZRpp3rBP5_1(.din(w_dff_B_pcpEuBTO7_1),.dout(w_dff_B_ZRpp3rBP5_1),.clk(gclk));
	jdff dff_B_D3k26w8o6_0(.din(n2889),.dout(w_dff_B_D3k26w8o6_0),.clk(gclk));
	jdff dff_B_LCRp0Mdl8_1(.din(n1582),.dout(w_dff_B_LCRp0Mdl8_1),.clk(gclk));
	jdff dff_B_l9iXkasH1_1(.din(w_dff_B_LCRp0Mdl8_1),.dout(w_dff_B_l9iXkasH1_1),.clk(gclk));
	jdff dff_B_znXfgxXr4_0(.din(n1586),.dout(w_dff_B_znXfgxXr4_0),.clk(gclk));
	jdff dff_B_vzerBgVm3_1(.din(n1618),.dout(w_dff_B_vzerBgVm3_1),.clk(gclk));
	jdff dff_B_m13q85Av4_1(.din(w_dff_B_vzerBgVm3_1),.dout(w_dff_B_m13q85Av4_1),.clk(gclk));
	jdff dff_B_CGPI3dHX3_0(.din(n1622),.dout(w_dff_B_CGPI3dHX3_0),.clk(gclk));
	jdff dff_B_4rpiYas84_1(.din(n1557),.dout(w_dff_B_4rpiYas84_1),.clk(gclk));
	jdff dff_B_ZxgD49R90_1(.din(w_dff_B_4rpiYas84_1),.dout(w_dff_B_ZxgD49R90_1),.clk(gclk));
	jdff dff_B_jew2rhCp7_0(.din(n1561),.dout(w_dff_B_jew2rhCp7_0),.clk(gclk));
	jdff dff_B_N8RSnojY1_1(.din(n1565),.dout(w_dff_B_N8RSnojY1_1),.clk(gclk));
	jdff dff_B_qvZOCGkh7_1(.din(w_dff_B_N8RSnojY1_1),.dout(w_dff_B_qvZOCGkh7_1),.clk(gclk));
	jdff dff_B_K6ULNMp38_0(.din(n1569),.dout(w_dff_B_K6ULNMp38_0),.clk(gclk));
	jdff dff_B_A6DxkfPQ0_1(.din(n2894),.dout(w_dff_B_A6DxkfPQ0_1),.clk(gclk));
	jdff dff_B_ykEXxVEF6_1(.din(w_dff_B_A6DxkfPQ0_1),.dout(w_dff_B_ykEXxVEF6_1),.clk(gclk));
	jdff dff_B_ZGsJLjTO8_0(.din(n2898),.dout(w_dff_B_ZGsJLjTO8_0),.clk(gclk));
	jdff dff_B_cryE1Kd60_1(.din(n1646),.dout(w_dff_B_cryE1Kd60_1),.clk(gclk));
	jdff dff_B_9liRMWfx0_1(.din(w_dff_B_cryE1Kd60_1),.dout(w_dff_B_9liRMWfx0_1),.clk(gclk));
	jdff dff_B_vqKakcLX8_0(.din(n1650),.dout(w_dff_B_vqKakcLX8_0),.clk(gclk));
	jdff dff_B_tl3HbU9G6_1(.din(n1666),.dout(w_dff_B_tl3HbU9G6_1),.clk(gclk));
	jdff dff_B_aGDLZ7hj2_1(.din(w_dff_B_tl3HbU9G6_1),.dout(w_dff_B_aGDLZ7hj2_1),.clk(gclk));
	jdff dff_B_qHBfuMtU9_0(.din(n1670),.dout(w_dff_B_qHBfuMtU9_0),.clk(gclk));
	jdff dff_B_EZu2XAm08_1(.din(n1691),.dout(w_dff_B_EZu2XAm08_1),.clk(gclk));
	jdff dff_B_WSOvahUp7_1(.din(w_dff_B_EZu2XAm08_1),.dout(w_dff_B_WSOvahUp7_1),.clk(gclk));
	jdff dff_B_YOOdvGcg9_0(.din(n1695),.dout(w_dff_B_YOOdvGcg9_0),.clk(gclk));
	jdff dff_B_8wkgG7hP0_1(.din(n1674),.dout(w_dff_B_8wkgG7hP0_1),.clk(gclk));
	jdff dff_B_f0Wxj4yd8_1(.din(w_dff_B_8wkgG7hP0_1),.dout(w_dff_B_f0Wxj4yd8_1),.clk(gclk));
	jdff dff_B_yLZkh10I4_0(.din(n1678),.dout(w_dff_B_yLZkh10I4_0),.clk(gclk));
	jdff dff_B_CGqmudAv9_1(.din(n2902),.dout(w_dff_B_CGqmudAv9_1),.clk(gclk));
	jdff dff_B_lhOl7scJ0_1(.din(w_dff_B_CGqmudAv9_1),.dout(w_dff_B_lhOl7scJ0_1),.clk(gclk));
	jdff dff_B_c2phCQGi0_0(.din(n2906),.dout(w_dff_B_c2phCQGi0_0),.clk(gclk));
	jdff dff_B_2YQMWR6R4_1(.din(n1655),.dout(w_dff_B_2YQMWR6R4_1),.clk(gclk));
	jdff dff_B_QBBmk80V1_1(.din(w_dff_B_2YQMWR6R4_1),.dout(w_dff_B_QBBmk80V1_1),.clk(gclk));
	jdff dff_B_U4CRJqxg3_0(.din(n1659),.dout(w_dff_B_U4CRJqxg3_0),.clk(gclk));
	jdff dff_B_BJhaO4Sm1_1(.din(n1638),.dout(w_dff_B_BJhaO4Sm1_1),.clk(gclk));
	jdff dff_B_fPXeCm1I9_1(.din(w_dff_B_BJhaO4Sm1_1),.dout(w_dff_B_fPXeCm1I9_1),.clk(gclk));
	jdff dff_B_GJ9JITL81_0(.din(n1642),.dout(w_dff_B_GJ9JITL81_0),.clk(gclk));
	jdff dff_B_CXBZKziI3_1(.din(n1630),.dout(w_dff_B_CXBZKziI3_1),.clk(gclk));
	jdff dff_B_9A8x5XsH6_1(.din(w_dff_B_CXBZKziI3_1),.dout(w_dff_B_9A8x5XsH6_1),.clk(gclk));
	jdff dff_B_yS8ELcW17_0(.din(n1634),.dout(w_dff_B_yS8ELcW17_0),.clk(gclk));
	jdff dff_B_mfY5h3s66_1(.din(n1682),.dout(w_dff_B_mfY5h3s66_1),.clk(gclk));
	jdff dff_B_m7kHuDJE5_1(.din(w_dff_B_mfY5h3s66_1),.dout(w_dff_B_m7kHuDJE5_1),.clk(gclk));
	jdff dff_B_fPFHHo2p6_0(.din(n1686),.dout(w_dff_B_fPFHHo2p6_0),.clk(gclk));
	jdff dff_B_TbHcYDTX8_1(.din(n2911),.dout(w_dff_B_TbHcYDTX8_1),.clk(gclk));
	jdff dff_B_OZhIiuq18_1(.din(w_dff_B_TbHcYDTX8_1),.dout(w_dff_B_OZhIiuq18_1),.clk(gclk));
	jdff dff_B_ZgZcwHQk4_0(.din(n2915),.dout(w_dff_B_ZgZcwHQk4_0),.clk(gclk));
	jdff dff_B_l03Q91CO4_1(.din(n1703),.dout(w_dff_B_l03Q91CO4_1),.clk(gclk));
	jdff dff_B_FiNXkb9Y6_1(.din(w_dff_B_l03Q91CO4_1),.dout(w_dff_B_FiNXkb9Y6_1),.clk(gclk));
	jdff dff_B_02mnb2b89_0(.din(n1707),.dout(w_dff_B_02mnb2b89_0),.clk(gclk));
	jdff dff_B_aui4nqcb5_1(.din(n1747),.dout(w_dff_B_aui4nqcb5_1),.clk(gclk));
	jdff dff_B_RIw4JiM62_1(.din(w_dff_B_aui4nqcb5_1),.dout(w_dff_B_RIw4JiM62_1),.clk(gclk));
	jdff dff_B_aQl6SJho8_0(.din(n1751),.dout(w_dff_B_aQl6SJho8_0),.clk(gclk));
	jdff dff_B_1ALoBJ3i8_1(.din(n1739),.dout(w_dff_B_1ALoBJ3i8_1),.clk(gclk));
	jdff dff_B_PPfha8iG0_1(.din(w_dff_B_1ALoBJ3i8_1),.dout(w_dff_B_PPfha8iG0_1),.clk(gclk));
	jdff dff_B_t7mqydWt3_0(.din(n1743),.dout(w_dff_B_t7mqydWt3_0),.clk(gclk));
	jdff dff_B_cZyPlB1Q5_1(.din(n1764),.dout(w_dff_B_cZyPlB1Q5_1),.clk(gclk));
	jdff dff_B_OSsMJ08H1_1(.din(w_dff_B_cZyPlB1Q5_1),.dout(w_dff_B_OSsMJ08H1_1),.clk(gclk));
	jdff dff_B_L33fN8wm0_0(.din(n1768),.dout(w_dff_B_L33fN8wm0_0),.clk(gclk));
	jdff dff_B_LseYXHtZ6_1(.din(n2919),.dout(w_dff_B_LseYXHtZ6_1),.clk(gclk));
	jdff dff_B_Vexy9pSD4_1(.din(w_dff_B_LseYXHtZ6_1),.dout(w_dff_B_Vexy9pSD4_1),.clk(gclk));
	jdff dff_B_PEtYO2nZ2_0(.din(n2923),.dout(w_dff_B_PEtYO2nZ2_0),.clk(gclk));
	jdff dff_B_ojgVuRDt2_1(.din(n1728),.dout(w_dff_B_ojgVuRDt2_1),.clk(gclk));
	jdff dff_B_iuUN1MS12_1(.din(w_dff_B_ojgVuRDt2_1),.dout(w_dff_B_iuUN1MS12_1),.clk(gclk));
	jdff dff_B_DXN0HrMN5_0(.din(n1732),.dout(w_dff_B_DXN0HrMN5_0),.clk(gclk));
	jdff dff_B_t1LazA034_1(.din(n1755),.dout(w_dff_B_t1LazA034_1),.clk(gclk));
	jdff dff_B_Fg5kkHG93_1(.din(w_dff_B_t1LazA034_1),.dout(w_dff_B_Fg5kkHG93_1),.clk(gclk));
	jdff dff_B_kjyfZ68B8_0(.din(n1759),.dout(w_dff_B_kjyfZ68B8_0),.clk(gclk));
	jdff dff_B_QWQqj8xb4_1(.din(n1719),.dout(w_dff_B_QWQqj8xb4_1),.clk(gclk));
	jdff dff_B_XgKuybAs2_1(.din(w_dff_B_QWQqj8xb4_1),.dout(w_dff_B_XgKuybAs2_1),.clk(gclk));
	jdff dff_B_N0xQg3RU2_0(.din(n1723),.dout(w_dff_B_N0xQg3RU2_0),.clk(gclk));
	jdff dff_B_DtzcDB6d0_1(.din(n1711),.dout(w_dff_B_DtzcDB6d0_1),.clk(gclk));
	jdff dff_B_3w20PdWI5_1(.din(w_dff_B_DtzcDB6d0_1),.dout(w_dff_B_3w20PdWI5_1),.clk(gclk));
	jdff dff_B_0KacSSWA2_0(.din(n1715),.dout(w_dff_B_0KacSSWA2_0),.clk(gclk));
	jdff dff_B_VnJASxDh2_1(.din(n2928),.dout(w_dff_B_VnJASxDh2_1),.clk(gclk));
	jdff dff_B_LOWVhPMa9_1(.din(w_dff_B_VnJASxDh2_1),.dout(w_dff_B_LOWVhPMa9_1),.clk(gclk));
	jdff dff_B_K2r8C8Bi4_0(.din(n2932),.dout(w_dff_B_K2r8C8Bi4_0),.clk(gclk));
	jdff dff_B_0RpO4pcF0_1(.din(n1820),.dout(w_dff_B_0RpO4pcF0_1),.clk(gclk));
	jdff dff_B_vZrVtr4g8_1(.din(w_dff_B_0RpO4pcF0_1),.dout(w_dff_B_vZrVtr4g8_1),.clk(gclk));
	jdff dff_B_aP2Vzczj8_0(.din(n1824),.dout(w_dff_B_aP2Vzczj8_0),.clk(gclk));
	jdff dff_B_FPwWCjoV9_1(.din(n1837),.dout(w_dff_B_FPwWCjoV9_1),.clk(gclk));
	jdff dff_B_buHD2ggE4_1(.din(w_dff_B_FPwWCjoV9_1),.dout(w_dff_B_buHD2ggE4_1),.clk(gclk));
	jdff dff_B_XBiAr6HB6_0(.din(n1841),.dout(w_dff_B_XBiAr6HB6_0),.clk(gclk));
	jdff dff_B_PCbR2CMZ5_1(.din(n1828),.dout(w_dff_B_PCbR2CMZ5_1),.clk(gclk));
	jdff dff_B_vFRPZe0E7_1(.din(w_dff_B_PCbR2CMZ5_1),.dout(w_dff_B_vFRPZe0E7_1),.clk(gclk));
	jdff dff_B_lFefcJ9l1_0(.din(n1832),.dout(w_dff_B_lFefcJ9l1_0),.clk(gclk));
	jdff dff_B_pgKvcWnY5_1(.din(n1801),.dout(w_dff_B_pgKvcWnY5_1),.clk(gclk));
	jdff dff_B_Fa5UygcP0_1(.din(w_dff_B_pgKvcWnY5_1),.dout(w_dff_B_Fa5UygcP0_1),.clk(gclk));
	jdff dff_B_nUofu0Ki0_0(.din(n1805),.dout(w_dff_B_nUofu0Ki0_0),.clk(gclk));
	jdff dff_B_nyJTp72i1_1(.din(n2936),.dout(w_dff_B_nyJTp72i1_1),.clk(gclk));
	jdff dff_B_ZIGeXFC22_1(.din(w_dff_B_nyJTp72i1_1),.dout(w_dff_B_ZIGeXFC22_1),.clk(gclk));
	jdff dff_B_iXUqkg6b0_0(.din(n2940),.dout(w_dff_B_iXUqkg6b0_0),.clk(gclk));
	jdff dff_B_ySBpqbGv9_1(.din(n1776),.dout(w_dff_B_ySBpqbGv9_1),.clk(gclk));
	jdff dff_B_QmpjNxjn9_1(.din(w_dff_B_ySBpqbGv9_1),.dout(w_dff_B_QmpjNxjn9_1),.clk(gclk));
	jdff dff_B_XA3R5mLm5_0(.din(n1780),.dout(w_dff_B_XA3R5mLm5_0),.clk(gclk));
	jdff dff_B_szz47Hzv6_1(.din(n1792),.dout(w_dff_B_szz47Hzv6_1),.clk(gclk));
	jdff dff_B_iky6qif53_1(.din(w_dff_B_szz47Hzv6_1),.dout(w_dff_B_iky6qif53_1),.clk(gclk));
	jdff dff_B_1jugmf9a1_0(.din(n1796),.dout(w_dff_B_1jugmf9a1_0),.clk(gclk));
	jdff dff_B_22ihCfHP1_1(.din(n1784),.dout(w_dff_B_22ihCfHP1_1),.clk(gclk));
	jdff dff_B_Z0mTHOxn2_1(.din(w_dff_B_22ihCfHP1_1),.dout(w_dff_B_Z0mTHOxn2_1),.clk(gclk));
	jdff dff_B_XXULzUgH7_0(.din(n1788),.dout(w_dff_B_XXULzUgH7_0),.clk(gclk));
	jdff dff_B_iCqvrP4J6_1(.din(n1812),.dout(w_dff_B_iCqvrP4J6_1),.clk(gclk));
	jdff dff_B_BBYKbmq80_1(.din(w_dff_B_iCqvrP4J6_1),.dout(w_dff_B_BBYKbmq80_1),.clk(gclk));
	jdff dff_B_bqScnAXr8_0(.din(n1816),.dout(w_dff_B_bqScnAXr8_0),.clk(gclk));
	jdff dff_B_xxdAL6Gg1_1(.din(n2945),.dout(w_dff_B_xxdAL6Gg1_1),.clk(gclk));
	jdff dff_B_ICBxgeIV7_1(.din(w_dff_B_xxdAL6Gg1_1),.dout(w_dff_B_ICBxgeIV7_1),.clk(gclk));
	jdff dff_B_YljleBFN9_0(.din(n2949),.dout(w_dff_B_YljleBFN9_0),.clk(gclk));
	jdff dff_B_V7meLCNO7_1(.din(n1874),.dout(w_dff_B_V7meLCNO7_1),.clk(gclk));
	jdff dff_B_12bjiM417_1(.din(w_dff_B_V7meLCNO7_1),.dout(w_dff_B_12bjiM417_1),.clk(gclk));
	jdff dff_B_WWcxEztL0_0(.din(n1878),.dout(w_dff_B_WWcxEztL0_0),.clk(gclk));
	jdff dff_B_5rVmUIn50_1(.din(n1885),.dout(w_dff_B_5rVmUIn50_1),.clk(gclk));
	jdff dff_B_FCK49IvL3_1(.din(w_dff_B_5rVmUIn50_1),.dout(w_dff_B_FCK49IvL3_1),.clk(gclk));
	jdff dff_B_a27ha2GA3_0(.din(n1889),.dout(w_dff_B_a27ha2GA3_0),.clk(gclk));
	jdff dff_B_ucTIwyaU5_1(.din(n1901),.dout(w_dff_B_ucTIwyaU5_1),.clk(gclk));
	jdff dff_B_z6Mk3N4z7_1(.din(w_dff_B_ucTIwyaU5_1),.dout(w_dff_B_z6Mk3N4z7_1),.clk(gclk));
	jdff dff_B_CwRb6Zdg9_0(.din(n1905),.dout(w_dff_B_CwRb6Zdg9_0),.clk(gclk));
	jdff dff_B_M7HzpFLq5_1(.din(n1893),.dout(w_dff_B_M7HzpFLq5_1),.clk(gclk));
	jdff dff_B_cC9wJqdw1_1(.din(w_dff_B_M7HzpFLq5_1),.dout(w_dff_B_cC9wJqdw1_1),.clk(gclk));
	jdff dff_B_u3s452In8_0(.din(n1897),.dout(w_dff_B_u3s452In8_0),.clk(gclk));
	jdff dff_B_GWN1KlHz0_1(.din(n2953),.dout(w_dff_B_GWN1KlHz0_1),.clk(gclk));
	jdff dff_B_8sKYsfXN5_1(.din(w_dff_B_GWN1KlHz0_1),.dout(w_dff_B_8sKYsfXN5_1),.clk(gclk));
	jdff dff_B_qzNhIp991_0(.din(n2957),.dout(w_dff_B_qzNhIp991_0),.clk(gclk));
	jdff dff_B_Ur6ue7jr2_1(.din(n1849),.dout(w_dff_B_Ur6ue7jr2_1),.clk(gclk));
	jdff dff_B_BhqJTvgw6_1(.din(w_dff_B_Ur6ue7jr2_1),.dout(w_dff_B_BhqJTvgw6_1),.clk(gclk));
	jdff dff_B_6p5HSVjj5_0(.din(n1853),.dout(w_dff_B_6p5HSVjj5_0),.clk(gclk));
	jdff dff_B_OyEk1U2B4_1(.din(n1910),.dout(w_dff_B_OyEk1U2B4_1),.clk(gclk));
	jdff dff_B_wM0cwS0E2_1(.din(w_dff_B_OyEk1U2B4_1),.dout(w_dff_B_wM0cwS0E2_1),.clk(gclk));
	jdff dff_B_eFTihvvF4_0(.din(n1914),.dout(w_dff_B_eFTihvvF4_0),.clk(gclk));
	jdff dff_B_4rqFI4Gy5_1(.din(n1857),.dout(w_dff_B_4rqFI4Gy5_1),.clk(gclk));
	jdff dff_B_mQYVjC3V5_1(.din(w_dff_B_4rqFI4Gy5_1),.dout(w_dff_B_mQYVjC3V5_1),.clk(gclk));
	jdff dff_B_W1m7NuUn4_0(.din(n1861),.dout(w_dff_B_W1m7NuUn4_0),.clk(gclk));
	jdff dff_B_z3S3oK5g3_1(.din(n1865),.dout(w_dff_B_z3S3oK5g3_1),.clk(gclk));
	jdff dff_B_U7tofJv50_1(.din(w_dff_B_z3S3oK5g3_1),.dout(w_dff_B_U7tofJv50_1),.clk(gclk));
	jdff dff_B_LXLqwXQf5_0(.din(n1869),.dout(w_dff_B_LXLqwXQf5_0),.clk(gclk));
	jdff dff_B_NPxcAtcs0_1(.din(n2962),.dout(w_dff_B_NPxcAtcs0_1),.clk(gclk));
	jdff dff_B_NGb1Pgpk3_1(.din(w_dff_B_NPxcAtcs0_1),.dout(w_dff_B_NGb1Pgpk3_1),.clk(gclk));
	jdff dff_B_vaIk44ui8_0(.din(n2966),.dout(w_dff_B_vaIk44ui8_0),.clk(gclk));
	jdff dff_B_SW6s5Ekj1_1(.din(n1938),.dout(w_dff_B_SW6s5Ekj1_1),.clk(gclk));
	jdff dff_B_HWXL2sOJ4_1(.din(w_dff_B_SW6s5Ekj1_1),.dout(w_dff_B_HWXL2sOJ4_1),.clk(gclk));
	jdff dff_B_IpfWp5MV0_0(.din(n1942),.dout(w_dff_B_IpfWp5MV0_0),.clk(gclk));
	jdff dff_B_gSBDtJ4S1_1(.din(n1966),.dout(w_dff_B_gSBDtJ4S1_1),.clk(gclk));
	jdff dff_B_0KDHoTdV3_1(.din(w_dff_B_gSBDtJ4S1_1),.dout(w_dff_B_0KDHoTdV3_1),.clk(gclk));
	jdff dff_B_fOzLotLx0_0(.din(n1970),.dout(w_dff_B_fOzLotLx0_0),.clk(gclk));
	jdff dff_B_m2ferJHn8_1(.din(n1974),.dout(w_dff_B_m2ferJHn8_1),.clk(gclk));
	jdff dff_B_HYrPEvnV5_1(.din(w_dff_B_m2ferJHn8_1),.dout(w_dff_B_HYrPEvnV5_1),.clk(gclk));
	jdff dff_B_osWnsPAs4_0(.din(n1978),.dout(w_dff_B_osWnsPAs4_0),.clk(gclk));
	jdff dff_B_zRQsCoKt9_1(.din(n1983),.dout(w_dff_B_zRQsCoKt9_1),.clk(gclk));
	jdff dff_B_vVdaNbcH6_1(.din(w_dff_B_zRQsCoKt9_1),.dout(w_dff_B_vVdaNbcH6_1),.clk(gclk));
	jdff dff_B_EyWT0czp2_0(.din(n1987),.dout(w_dff_B_EyWT0czp2_0),.clk(gclk));
	jdff dff_B_pTGLz1Ga5_1(.din(n2970),.dout(w_dff_B_pTGLz1Ga5_1),.clk(gclk));
	jdff dff_B_BUCvsxNO3_1(.din(w_dff_B_pTGLz1Ga5_1),.dout(w_dff_B_BUCvsxNO3_1),.clk(gclk));
	jdff dff_B_lnxYEnyW2_0(.din(n2974),.dout(w_dff_B_lnxYEnyW2_0),.clk(gclk));
	jdff dff_B_WVMYNQRc8_1(.din(n1947),.dout(w_dff_B_WVMYNQRc8_1),.clk(gclk));
	jdff dff_B_EQkAxmtM8_1(.din(w_dff_B_WVMYNQRc8_1),.dout(w_dff_B_EQkAxmtM8_1),.clk(gclk));
	jdff dff_B_g3hpVPxg1_0(.din(n1951),.dout(w_dff_B_g3hpVPxg1_0),.clk(gclk));
	jdff dff_B_L2tsbO6u6_1(.din(n1958),.dout(w_dff_B_L2tsbO6u6_1),.clk(gclk));
	jdff dff_B_75VVNHvJ2_1(.din(w_dff_B_L2tsbO6u6_1),.dout(w_dff_B_75VVNHvJ2_1),.clk(gclk));
	jdff dff_B_UgfuBzO50_0(.din(n1962),.dout(w_dff_B_UgfuBzO50_0),.clk(gclk));
	jdff dff_B_6uroEMmR5_1(.din(n1930),.dout(w_dff_B_6uroEMmR5_1),.clk(gclk));
	jdff dff_B_Y7YtLhzO6_1(.din(w_dff_B_6uroEMmR5_1),.dout(w_dff_B_Y7YtLhzO6_1),.clk(gclk));
	jdff dff_B_D38jD0K72_0(.din(n1934),.dout(w_dff_B_D38jD0K72_0),.clk(gclk));
	jdff dff_B_AQTDvday7_1(.din(n1922),.dout(w_dff_B_AQTDvday7_1),.clk(gclk));
	jdff dff_B_lH0Rc6Lf0_1(.din(w_dff_B_AQTDvday7_1),.dout(w_dff_B_lH0Rc6Lf0_1),.clk(gclk));
	jdff dff_B_U5D9P6Db9_0(.din(n1926),.dout(w_dff_B_U5D9P6Db9_0),.clk(gclk));
	jdff dff_B_mUqQUmBj9_1(.din(n2979),.dout(w_dff_B_mUqQUmBj9_1),.clk(gclk));
	jdff dff_B_JqSHsLGG2_1(.din(w_dff_B_mUqQUmBj9_1),.dout(w_dff_B_JqSHsLGG2_1),.clk(gclk));
	jdff dff_B_id4K03Wa5_0(.din(n2983),.dout(w_dff_B_id4K03Wa5_0),.clk(gclk));
	jdff dff_B_jMNibkDP1_1(.din(n2011),.dout(w_dff_B_jMNibkDP1_1),.clk(gclk));
	jdff dff_B_6iCFG5SY4_1(.din(w_dff_B_jMNibkDP1_1),.dout(w_dff_B_6iCFG5SY4_1),.clk(gclk));
	jdff dff_B_l2iJDWqD9_0(.din(n2015),.dout(w_dff_B_l2iJDWqD9_0),.clk(gclk));
	jdff dff_B_RE1qjwxi1_1(.din(n2039),.dout(w_dff_B_RE1qjwxi1_1),.clk(gclk));
	jdff dff_B_174ZvsxD2_1(.din(w_dff_B_RE1qjwxi1_1),.dout(w_dff_B_174ZvsxD2_1),.clk(gclk));
	jdff dff_B_Tg33vzS97_0(.din(n2043),.dout(w_dff_B_Tg33vzS97_0),.clk(gclk));
	jdff dff_B_Sdr4G0ZW3_1(.din(n2056),.dout(w_dff_B_Sdr4G0ZW3_1),.clk(gclk));
	jdff dff_B_h8DUDHPi9_1(.din(w_dff_B_Sdr4G0ZW3_1),.dout(w_dff_B_h8DUDHPi9_1),.clk(gclk));
	jdff dff_B_92yjbt7N5_0(.din(n2060),.dout(w_dff_B_92yjbt7N5_0),.clk(gclk));
	jdff dff_B_gXXxnHFS1_1(.din(n2031),.dout(w_dff_B_gXXxnHFS1_1),.clk(gclk));
	jdff dff_B_slVYtXoH6_1(.din(w_dff_B_gXXxnHFS1_1),.dout(w_dff_B_slVYtXoH6_1),.clk(gclk));
	jdff dff_B_zURs38kR5_0(.din(n2035),.dout(w_dff_B_zURs38kR5_0),.clk(gclk));
	jdff dff_B_0I265xjZ5_1(.din(n2987),.dout(w_dff_B_0I265xjZ5_1),.clk(gclk));
	jdff dff_B_MNkhRkVJ2_1(.din(w_dff_B_0I265xjZ5_1),.dout(w_dff_B_MNkhRkVJ2_1),.clk(gclk));
	jdff dff_B_mNvo9h4e6_0(.din(n2991),.dout(w_dff_B_mNvo9h4e6_0),.clk(gclk));
	jdff dff_B_HegFkakD8_1(.din(n1995),.dout(w_dff_B_HegFkakD8_1),.clk(gclk));
	jdff dff_B_tbWgCQ7T5_1(.din(w_dff_B_HegFkakD8_1),.dout(w_dff_B_tbWgCQ7T5_1),.clk(gclk));
	jdff dff_B_0gJiH3OV1_0(.din(n1999),.dout(w_dff_B_0gJiH3OV1_0),.clk(gclk));
	jdff dff_B_Bb2LQOX46_1(.din(n2047),.dout(w_dff_B_Bb2LQOX46_1),.clk(gclk));
	jdff dff_B_VbO6w6zD2_1(.din(w_dff_B_Bb2LQOX46_1),.dout(w_dff_B_VbO6w6zD2_1),.clk(gclk));
	jdff dff_B_3s6AjRKb2_0(.din(n2051),.dout(w_dff_B_3s6AjRKb2_0),.clk(gclk));
	jdff dff_B_0f5VWSQ93_1(.din(n2003),.dout(w_dff_B_0f5VWSQ93_1),.clk(gclk));
	jdff dff_B_Z7fK2rF58_1(.din(w_dff_B_0f5VWSQ93_1),.dout(w_dff_B_Z7fK2rF58_1),.clk(gclk));
	jdff dff_B_M8RJIFvs4_0(.din(n2007),.dout(w_dff_B_M8RJIFvs4_0),.clk(gclk));
	jdff dff_B_T1dMgkpZ6_1(.din(n2020),.dout(w_dff_B_T1dMgkpZ6_1),.clk(gclk));
	jdff dff_B_rD7Jx1Kl7_1(.din(w_dff_B_T1dMgkpZ6_1),.dout(w_dff_B_rD7Jx1Kl7_1),.clk(gclk));
	jdff dff_B_Q96lHp3o5_0(.din(n2024),.dout(w_dff_B_Q96lHp3o5_0),.clk(gclk));
	jdff dff_B_xoinFbqO8_1(.din(n2996),.dout(w_dff_B_xoinFbqO8_1),.clk(gclk));
	jdff dff_B_yEJJMF8P9_1(.din(w_dff_B_xoinFbqO8_1),.dout(w_dff_B_yEJJMF8P9_1),.clk(gclk));
	jdff dff_B_m0Sng1PW4_0(.din(n3000),.dout(w_dff_B_m0Sng1PW4_0),.clk(gclk));
	jdff dff_B_MdIApfCQ7_1(.din(n2084),.dout(w_dff_B_MdIApfCQ7_1),.clk(gclk));
	jdff dff_B_46as8xFJ1_1(.din(w_dff_B_MdIApfCQ7_1),.dout(w_dff_B_46as8xFJ1_1),.clk(gclk));
	jdff dff_B_JGDoXU1T7_0(.din(n2088),.dout(w_dff_B_JGDoXU1T7_0),.clk(gclk));
	jdff dff_B_8SdLIGhZ4_1(.din(n482),.dout(w_dff_B_8SdLIGhZ4_1),.clk(gclk));
	jdff dff_B_sqwDOK3F5_1(.din(n468),.dout(w_dff_B_sqwDOK3F5_1),.clk(gclk));
	jdff dff_B_wXVKtnh13_1(.din(n462),.dout(w_dff_B_wXVKtnh13_1),.clk(gclk));
	jdff dff_B_jlhhO1862_1(.din(n365),.dout(w_dff_B_jlhhO1862_1),.clk(gclk));
	jdff dff_B_xqLjxEhE3_1(.din(n472),.dout(w_dff_B_xqLjxEhE3_1),.clk(gclk));
	jdff dff_B_gnnLsEbL7_1(.din(n458),.dout(w_dff_B_gnnLsEbL7_1),.clk(gclk));
	jdff dff_B_LvNxJLXv2_1(.din(n493),.dout(w_dff_B_LvNxJLXv2_1),.clk(gclk));
	jdff dff_B_1erSQF5v5_1(.din(n478),.dout(w_dff_B_1erSQF5v5_1),.clk(gclk));
	jdff dff_B_73zz0aOP0_1(.din(n2129),.dout(w_dff_B_73zz0aOP0_1),.clk(gclk));
	jdff dff_B_kx18ekQ99_1(.din(w_dff_B_73zz0aOP0_1),.dout(w_dff_B_kx18ekQ99_1),.clk(gclk));
	jdff dff_B_PVvmUK9a6_0(.din(n2133),.dout(w_dff_B_PVvmUK9a6_0),.clk(gclk));
	jdff dff_B_RDrOvlHB2_1(.din(n581),.dout(w_dff_B_RDrOvlHB2_1),.clk(gclk));
	jdff dff_B_lrsiFJkx2_1(.din(n546),.dout(w_dff_B_lrsiFJkx2_1),.clk(gclk));
	jdff dff_B_3XYmQ7xa1_1(.din(n550),.dout(w_dff_B_3XYmQ7xa1_1),.clk(gclk));
	jdff dff_B_kbso0kek4_1(.din(n556),.dout(w_dff_B_kbso0kek4_1),.clk(gclk));
	jdff dff_B_a2qEd9k26_1(.din(n560),.dout(w_dff_B_a2qEd9k26_1),.clk(gclk));
	jdff dff_B_KkZUlkQY5_1(.din(n566),.dout(w_dff_B_KkZUlkQY5_1),.clk(gclk));
	jdff dff_B_gUpOzecm7_1(.din(n570),.dout(w_dff_B_gUpOzecm7_1),.clk(gclk));
	jdff dff_B_qDiElXBG9_1(.din(n489),.dout(w_dff_B_qDiElXBG9_1),.clk(gclk));
	jdff dff_B_peT3tE445_1(.din(n2104),.dout(w_dff_B_peT3tE445_1),.clk(gclk));
	jdff dff_B_FFv3MKX02_1(.din(w_dff_B_peT3tE445_1),.dout(w_dff_B_FFv3MKX02_1),.clk(gclk));
	jdff dff_B_0oY8yfNB8_0(.din(n2108),.dout(w_dff_B_0oY8yfNB8_0),.clk(gclk));
	jdff dff_B_USEsFc4E6_1(.din(n537),.dout(w_dff_B_USEsFc4E6_1),.clk(gclk));
	jdff dff_B_qxZUuMrc2_1(.din(n522),.dout(w_dff_B_qxZUuMrc2_1),.clk(gclk));
	jdff dff_B_bUuUbKk52_1(.din(n526),.dout(w_dff_B_bUuUbKk52_1),.clk(gclk));
	jdff dff_B_0JQMoqEd2_1(.din(n512),.dout(w_dff_B_0JQMoqEd2_1),.clk(gclk));
	jdff dff_B_DBajLoEy0_1(.din(n516),.dout(w_dff_B_DBajLoEy0_1),.clk(gclk));
	jdff dff_B_oANUBuw89_1(.din(n502),.dout(w_dff_B_oANUBuw89_1),.clk(gclk));
	jdff dff_B_ZtYCSpfs0_1(.din(n506),.dout(w_dff_B_ZtYCSpfs0_1),.clk(gclk));
	jdff dff_B_kMwsZSDe0_1(.din(n577),.dout(w_dff_B_kMwsZSDe0_1),.clk(gclk));
	jdff dff_B_v0bLqLBi4_1(.din(n2112),.dout(w_dff_B_v0bLqLBi4_1),.clk(gclk));
	jdff dff_B_pvT9nqua2_1(.din(w_dff_B_v0bLqLBi4_1),.dout(w_dff_B_pvT9nqua2_1),.clk(gclk));
	jdff dff_B_tozgo1T96_0(.din(n2116),.dout(w_dff_B_tozgo1T96_0),.clk(gclk));
	jdff dff_B_DgWSqdmm5_1(.din(n615),.dout(w_dff_B_DgWSqdmm5_1),.clk(gclk));
	jdff dff_B_eNbCbCNd4_1(.din(n533),.dout(w_dff_B_eNbCbCNd4_1),.clk(gclk));
	jdff dff_B_pBoU1aAC0_1(.din(n595),.dout(w_dff_B_pBoU1aAC0_1),.clk(gclk));
	jdff dff_B_G73nas932_1(.din(n601),.dout(w_dff_B_G73nas932_1),.clk(gclk));
	jdff dff_B_oX8bH2f69_1(.din(n605),.dout(w_dff_B_oX8bH2f69_1),.clk(gclk));
	jdff dff_B_Nhlo4skL5_1(.din(n611),.dout(w_dff_B_Nhlo4skL5_1),.clk(gclk));
	jdff dff_B_LxADl0g43_1(.din(n626),.dout(w_dff_B_LxADl0g43_1),.clk(gclk));
	jdff dff_B_0RsxGrIy5_1(.din(n591),.dout(w_dff_B_0RsxGrIy5_1),.clk(gclk));
	jdff dff_B_N69ZWpDm5_1(.din(n3004),.dout(w_dff_B_N69ZWpDm5_1),.clk(gclk));
	jdff dff_B_kUjye1l65_1(.din(w_dff_B_N69ZWpDm5_1),.dout(w_dff_B_kUjye1l65_1),.clk(gclk));
	jdff dff_B_hIuzRHwv3_0(.din(n3008),.dout(w_dff_B_hIuzRHwv3_0),.clk(gclk));
	jdff dff_B_2dW9nCZU7_1(.din(n2068),.dout(w_dff_B_2dW9nCZU7_1),.clk(gclk));
	jdff dff_B_ylFxSofU1_1(.din(w_dff_B_2dW9nCZU7_1),.dout(w_dff_B_ylFxSofU1_1),.clk(gclk));
	jdff dff_B_Jtue7Ywt4_0(.din(n2072),.dout(w_dff_B_Jtue7Ywt4_0),.clk(gclk));
	jdff dff_B_rGGKJFCI5_1(.din(n400),.dout(w_dff_B_rGGKJFCI5_1),.clk(gclk));
	jdff dff_B_H3GTqRv49_1(.din(n351),.dout(w_dff_B_H3GTqRv49_1),.clk(gclk));
	jdff dff_B_8ry3nHbt8_1(.din(n389),.dout(w_dff_B_8ry3nHbt8_1),.clk(gclk));
	jdff dff_B_nAuGj7r26_1(.din(n375),.dout(w_dff_B_nAuGj7r26_1),.clk(gclk));
	jdff dff_B_ZCt0lbDj7_1(.din(n379),.dout(w_dff_B_ZCt0lbDj7_1),.clk(gclk));
	jdff dff_B_qGz8nn0O6_1(.din(n396),.dout(w_dff_B_qGz8nn0O6_1),.clk(gclk));
	jdff dff_B_qCna0wrc1_1(.din(n369),.dout(w_dff_B_qCna0wrc1_1),.clk(gclk));
	jdff dff_B_1MK5rQm16_1(.din(n385),.dout(w_dff_B_1MK5rQm16_1),.clk(gclk));
	jdff dff_B_N2gd7BK42_1(.din(n2093),.dout(w_dff_B_N2gd7BK42_1),.clk(gclk));
	jdff dff_B_hk70EXhB4_1(.din(w_dff_B_N2gd7BK42_1),.dout(w_dff_B_hk70EXhB4_1),.clk(gclk));
	jdff dff_B_fnNiVSQg0_0(.din(n2097),.dout(w_dff_B_fnNiVSQg0_0),.clk(gclk));
	jdff dff_B_zn2dswtc8_1(.din(n340),.dout(w_dff_B_zn2dswtc8_1),.clk(gclk));
	jdff dff_B_J9KIgtCx9_1(.din(n355),.dout(w_dff_B_J9KIgtCx9_1),.clk(gclk));
	jdff dff_B_YlyhWCe47_1(.din(n324),.dout(w_dff_B_YlyhWCe47_1),.clk(gclk));
	jdff dff_B_pbjsvJRU0_1(.din(n305),.dout(w_dff_B_pbjsvJRU0_1),.clk(gclk));
	jdff dff_B_1NL5v4dj1_1(.din(n334),.dout(w_dff_B_1NL5v4dj1_1),.clk(gclk));
	jdff dff_B_cHVmEYYS1_1(.din(n320),.dout(w_dff_B_cHVmEYYS1_1),.clk(gclk));
	jdff dff_B_tmydoCWx9_1(.din(n344),.dout(w_dff_B_tmydoCWx9_1),.clk(gclk));
	jdff dff_B_dSDMYpiX8_1(.din(n330),.dout(w_dff_B_dSDMYpiX8_1),.clk(gclk));
	jdff dff_B_yWsrWUVz8_1(.din(n2076),.dout(w_dff_B_yWsrWUVz8_1),.clk(gclk));
	jdff dff_B_PJjnjmSe8_1(.din(w_dff_B_yWsrWUVz8_1),.dout(w_dff_B_PJjnjmSe8_1),.clk(gclk));
	jdff dff_B_b8CiSugl5_0(.din(n2080),.dout(w_dff_B_b8CiSugl5_0),.clk(gclk));
	jdff dff_B_4u4V4i842_1(.din(n309),.dout(w_dff_B_4u4V4i842_1),.clk(gclk));
	jdff dff_B_HatNyVWj5_1(.din(n268),.dout(w_dff_B_HatNyVWj5_1),.clk(gclk));
	jdff dff_B_EftOFYUE7_1(.din(n274),.dout(w_dff_B_EftOFYUE7_1),.clk(gclk));
	jdff dff_B_OFdIWwF79_1(.din(n282),.dout(w_dff_B_OFdIWwF79_1),.clk(gclk));
	jdff dff_B_of9B41I48_1(.din(n286),.dout(w_dff_B_of9B41I48_1),.clk(gclk));
	jdff dff_B_ZQDJ7Ux87_1(.din(n293),.dout(w_dff_B_ZQDJ7Ux87_1),.clk(gclk));
	jdff dff_B_HdRHntcb1_1(.din(n297),.dout(w_dff_B_HdRHntcb1_1),.clk(gclk));
	jdff dff_B_LlIFSUYG1_1(.din(n442),.dout(w_dff_B_LlIFSUYG1_1),.clk(gclk));
	jdff dff_B_ga74nord4_1(.din(n2120),.dout(w_dff_B_ga74nord4_1),.clk(gclk));
	jdff dff_B_vg76XKpv7_1(.din(w_dff_B_ga74nord4_1),.dout(w_dff_B_vg76XKpv7_1),.clk(gclk));
	jdff dff_B_rECqHm9H4_0(.din(n2124),.dout(w_dff_B_rECqHm9H4_0),.clk(gclk));
	jdff dff_B_EdOZ8SLX0_1(.din(n415),.dout(w_dff_B_EdOZ8SLX0_1),.clk(gclk));
	jdff dff_B_qelqFzvL8_1(.din(n421),.dout(w_dff_B_qelqFzvL8_1),.clk(gclk));
	jdff dff_B_Y1FGDnUK0_1(.din(n435),.dout(w_dff_B_Y1FGDnUK0_1),.clk(gclk));
	jdff dff_B_OXno1hik8_1(.din(n622),.dout(w_dff_B_OXno1hik8_1),.clk(gclk));
	jdff dff_B_r7LsM7Df4_1(.din(n425),.dout(w_dff_B_r7LsM7Df4_1),.clk(gclk));
	jdff dff_B_e7wXA7DB3_1(.din(n431),.dout(w_dff_B_e7wXA7DB3_1),.clk(gclk));
	jdff dff_B_psoYtpqQ6_1(.din(n446),.dout(w_dff_B_psoYtpqQ6_1),.clk(gclk));
	jdff dff_B_hHESg9fo8_1(.din(n411),.dout(w_dff_B_hHESg9fo8_1),.clk(gclk));
	jdff dff_B_sukwBUro7_1(.din(n3013),.dout(w_dff_B_sukwBUro7_1),.clk(gclk));
	jdff dff_B_qIVWh7nJ2_1(.din(w_dff_B_sukwBUro7_1),.dout(w_dff_B_qIVWh7nJ2_1),.clk(gclk));
	jdff dff_B_b2g877Zq9_0(.din(n3017),.dout(w_dff_B_b2g877Zq9_0),.clk(gclk));
	jdff dff_B_nVt1r1Pg4_1(.din(n2166),.dout(w_dff_B_nVt1r1Pg4_1),.clk(gclk));
	jdff dff_B_3n3bcFZF0_1(.din(w_dff_B_nVt1r1Pg4_1),.dout(w_dff_B_3n3bcFZF0_1),.clk(gclk));
	jdff dff_B_yFXClqjf2_0(.din(n2170),.dout(w_dff_B_yFXClqjf2_0),.clk(gclk));
	jdff dff_B_lGKQzauE6_1(.din(n854),.dout(w_dff_B_lGKQzauE6_1),.clk(gclk));
	jdff dff_A_4pYXSgZQ4_0(.dout(w_a78_0[0]),.din(w_dff_A_4pYXSgZQ4_0),.clk(gclk));
	jdff dff_A_eOY9af3E1_1(.dout(w_a79_0[1]),.din(w_dff_A_eOY9af3E1_1),.clk(gclk));
	jdff dff_B_b1xub7d40_1(.din(n839),.dout(w_dff_B_b1xub7d40_1),.clk(gclk));
	jdff dff_A_jsqcgtqV5_0(.dout(w_a76_0[0]),.din(w_dff_A_jsqcgtqV5_0),.clk(gclk));
	jdff dff_A_Tf7v1fro5_1(.dout(w_a77_0[1]),.din(w_dff_A_Tf7v1fro5_1),.clk(gclk));
	jdff dff_B_qUAu1S6Q0_1(.din(n843),.dout(w_dff_B_qUAu1S6Q0_1),.clk(gclk));
	jdff dff_A_I7gyfdFq9_0(.dout(w_a74_0[0]),.din(w_dff_A_I7gyfdFq9_0),.clk(gclk));
	jdff dff_A_NA9ziZSD5_1(.dout(w_a75_0[1]),.din(w_dff_A_NA9ziZSD5_1),.clk(gclk));
	jdff dff_B_BcmFF8576_1(.din(n829),.dout(w_dff_B_BcmFF8576_1),.clk(gclk));
	jdff dff_A_3gOkgdes3_0(.dout(w_a72_0[0]),.din(w_dff_A_3gOkgdes3_0),.clk(gclk));
	jdff dff_A_tD9nMY0t2_1(.dout(w_a73_0[1]),.din(w_dff_A_tD9nMY0t2_1),.clk(gclk));
	jdff dff_B_Q6hzBaEe4_1(.din(n833),.dout(w_dff_B_Q6hzBaEe4_1),.clk(gclk));
	jdff dff_A_bhAqClr40_0(.dout(w_a70_0[0]),.din(w_dff_A_bhAqClr40_0),.clk(gclk));
	jdff dff_A_qYdmnUej7_1(.dout(w_a71_0[1]),.din(w_dff_A_qYdmnUej7_1),.clk(gclk));
	jdff dff_B_ZwKVErzE1_1(.din(n819),.dout(w_dff_B_ZwKVErzE1_1),.clk(gclk));
	jdff dff_A_SwhSpGG03_0(.dout(w_a68_0[0]),.din(w_dff_A_SwhSpGG03_0),.clk(gclk));
	jdff dff_A_yYiuMmAx6_1(.dout(w_a69_0[1]),.din(w_dff_A_yYiuMmAx6_1),.clk(gclk));
	jdff dff_B_i0X0OPVY5_1(.din(n823),.dout(w_dff_B_i0X0OPVY5_1),.clk(gclk));
	jdff dff_A_aYzwVtdH1_0(.dout(w_a66_0[0]),.din(w_dff_A_aYzwVtdH1_0),.clk(gclk));
	jdff dff_A_9PjzwdE12_1(.dout(w_a67_0[1]),.din(w_dff_A_9PjzwdE12_1),.clk(gclk));
	jdff dff_B_sqLFKCT85_1(.din(n670),.dout(w_dff_B_sqLFKCT85_1),.clk(gclk));
	jdff dff_A_ipr72ra02_0(.dout(w_a64_0[0]),.din(w_dff_A_ipr72ra02_0),.clk(gclk));
	jdff dff_A_APWgC3dM4_1(.dout(w_a65_0[1]),.din(w_dff_A_APWgC3dM4_1),.clk(gclk));
	jdff dff_B_f7q9HcgA4_1(.din(n2202),.dout(w_dff_B_f7q9HcgA4_1),.clk(gclk));
	jdff dff_B_rUo3KNte8_1(.din(w_dff_B_f7q9HcgA4_1),.dout(w_dff_B_rUo3KNte8_1),.clk(gclk));
	jdff dff_B_QlNfdnSh4_0(.din(n2206),.dout(w_dff_B_QlNfdnSh4_0),.clk(gclk));
	jdff dff_B_WSLDAw9h6_1(.din(n942),.dout(w_dff_B_WSLDAw9h6_1),.clk(gclk));
	jdff dff_A_Xt1EtlJu1_0(.dout(w_a94_0[0]),.din(w_dff_A_Xt1EtlJu1_0),.clk(gclk));
	jdff dff_A_Pe361rYG6_1(.dout(w_a95_0[1]),.din(w_dff_A_Pe361rYG6_1),.clk(gclk));
	jdff dff_B_yG764QYf5_1(.din(n927),.dout(w_dff_B_yG764QYf5_1),.clk(gclk));
	jdff dff_A_8B97r3VV0_0(.dout(w_a92_0[0]),.din(w_dff_A_8B97r3VV0_0),.clk(gclk));
	jdff dff_A_RTG96NZT0_1(.dout(w_a93_0[1]),.din(w_dff_A_RTG96NZT0_1),.clk(gclk));
	jdff dff_B_42tADvHd7_1(.din(n911),.dout(w_dff_B_42tADvHd7_1),.clk(gclk));
	jdff dff_A_wSYwKQKp9_0(.dout(w_a82_0[0]),.din(w_dff_A_wSYwKQKp9_0),.clk(gclk));
	jdff dff_A_OiMf06K86_1(.dout(w_a83_0[1]),.din(w_dff_A_OiMf06K86_1),.clk(gclk));
	jdff dff_B_KImY48fm3_1(.din(n850),.dout(w_dff_B_KImY48fm3_1),.clk(gclk));
	jdff dff_A_FxenSOIp9_0(.dout(w_a80_0[0]),.din(w_dff_A_FxenSOIp9_0),.clk(gclk));
	jdff dff_A_X1Lfnzwj8_1(.dout(w_a81_0[1]),.din(w_dff_A_X1Lfnzwj8_1),.clk(gclk));
	jdff dff_B_XT5fswlN8_1(.din(n921),.dout(w_dff_B_XT5fswlN8_1),.clk(gclk));
	jdff dff_A_5fD5AaYw7_0(.dout(w_a86_0[0]),.din(w_dff_A_5fD5AaYw7_0),.clk(gclk));
	jdff dff_A_TrlnadzK5_1(.dout(w_a87_0[1]),.din(w_dff_A_TrlnadzK5_1),.clk(gclk));
	jdff dff_B_uvuIOWOm0_1(.din(n907),.dout(w_dff_B_uvuIOWOm0_1),.clk(gclk));
	jdff dff_A_i8HqUX7H4_0(.dout(w_a84_0[0]),.din(w_dff_A_i8HqUX7H4_0),.clk(gclk));
	jdff dff_A_OcSdyoQr6_1(.dout(w_a85_0[1]),.din(w_dff_A_OcSdyoQr6_1),.clk(gclk));
	jdff dff_B_8NBshqAL6_1(.din(n931),.dout(w_dff_B_8NBshqAL6_1),.clk(gclk));
	jdff dff_A_p4g9Yx0Z8_0(.dout(w_a90_0[0]),.din(w_dff_A_p4g9Yx0Z8_0),.clk(gclk));
	jdff dff_A_OxxYjRfR3_1(.dout(w_a91_0[1]),.din(w_dff_A_OxxYjRfR3_1),.clk(gclk));
	jdff dff_B_NrGt6CJe2_1(.din(n917),.dout(w_dff_B_NrGt6CJe2_1),.clk(gclk));
	jdff dff_A_nt5Btme91_0(.dout(w_a88_0[0]),.din(w_dff_A_nt5Btme91_0),.clk(gclk));
	jdff dff_A_uSzz6U2s7_1(.dout(w_a89_0[1]),.din(w_dff_A_uSzz6U2s7_1),.clk(gclk));
	jdff dff_B_xgjTbxSc2_1(.din(n2193),.dout(w_dff_B_xgjTbxSc2_1),.clk(gclk));
	jdff dff_B_zacrjjWS4_1(.din(w_dff_B_xgjTbxSc2_1),.dout(w_dff_B_zacrjjWS4_1),.clk(gclk));
	jdff dff_B_5qLGuZg58_0(.din(n2197),.dout(w_dff_B_5qLGuZg58_0),.clk(gclk));
	jdff dff_B_py7Eagjp9_1(.din(n867),.dout(w_dff_B_py7Eagjp9_1),.clk(gclk));
	jdff dff_A_4h0NH7LH3_0(.dout(w_a98_0[0]),.din(w_dff_A_4h0NH7LH3_0),.clk(gclk));
	jdff dff_A_amGWYNxX5_1(.dout(w_a99_0[1]),.din(w_dff_A_amGWYNxX5_1),.clk(gclk));
	jdff dff_B_8EZYNZap4_1(.din(n938),.dout(w_dff_B_8EZYNZap4_1),.clk(gclk));
	jdff dff_A_HbBmurSs9_0(.dout(w_a96_0[0]),.din(w_dff_A_HbBmurSs9_0),.clk(gclk));
	jdff dff_A_3E0UAqQJ7_1(.dout(w_a97_0[1]),.din(w_dff_A_3E0UAqQJ7_1),.clk(gclk));
	jdff dff_B_1lzHYFyY3_1(.din(n887),.dout(w_dff_B_1lzHYFyY3_1),.clk(gclk));
	jdff dff_A_BB5cJRhF0_0(.dout(w_a106_0[0]),.din(w_dff_A_BB5cJRhF0_0),.clk(gclk));
	jdff dff_A_x0WLNzz69_1(.dout(w_a107_0[1]),.din(w_dff_A_x0WLNzz69_1),.clk(gclk));
	jdff dff_B_iPHr0LC45_1(.din(n873),.dout(w_dff_B_iPHr0LC45_1),.clk(gclk));
	jdff dff_A_KWIu5I4M0_0(.dout(w_a104_0[0]),.din(w_dff_A_KWIu5I4M0_0),.clk(gclk));
	jdff dff_A_NhWoqlJE7_1(.dout(w_a105_0[1]),.din(w_dff_A_NhWoqlJE7_1),.clk(gclk));
	jdff dff_B_LzHuIvWe7_1(.din(n877),.dout(w_dff_B_LzHuIvWe7_1),.clk(gclk));
	jdff dff_A_x1m5wCkQ3_0(.dout(w_a102_0[0]),.din(w_dff_A_x1m5wCkQ3_0),.clk(gclk));
	jdff dff_A_fFCBlUt64_1(.dout(w_a103_0[1]),.din(w_dff_A_fFCBlUt64_1),.clk(gclk));
	jdff dff_B_mXMNmnXD2_1(.din(n863),.dout(w_dff_B_mXMNmnXD2_1),.clk(gclk));
	jdff dff_A_tioEWBSH6_0(.dout(w_a100_0[0]),.din(w_dff_A_tioEWBSH6_0),.clk(gclk));
	jdff dff_A_iMM7uM3x0_1(.dout(w_a101_0[1]),.din(w_dff_A_iMM7uM3x0_1),.clk(gclk));
	jdff dff_B_Qru46Pym3_1(.din(n898),.dout(w_dff_B_Qru46Pym3_1),.clk(gclk));
	jdff dff_A_a4SNezFT6_0(.dout(w_a110_0[0]),.din(w_dff_A_a4SNezFT6_0),.clk(gclk));
	jdff dff_A_bbcJxZ647_1(.dout(w_a111_0[1]),.din(w_dff_A_bbcJxZ647_1),.clk(gclk));
	jdff dff_B_LyBW2d6f4_1(.din(n883),.dout(w_dff_B_LyBW2d6f4_1),.clk(gclk));
	jdff dff_A_3R8e6hTN0_0(.dout(w_a108_0[0]),.din(w_dff_A_3R8e6hTN0_0),.clk(gclk));
	jdff dff_A_nyGrOAiO3_1(.dout(w_a109_0[1]),.din(w_dff_A_nyGrOAiO3_1),.clk(gclk));
	jdff dff_B_vJXNk5uA4_1(.din(n2185),.dout(w_dff_B_vJXNk5uA4_1),.clk(gclk));
	jdff dff_B_DlowA4MC0_1(.din(w_dff_B_vJXNk5uA4_1),.dout(w_dff_B_DlowA4MC0_1),.clk(gclk));
	jdff dff_B_bqhhQYEO8_0(.din(n2189),.dout(w_dff_B_bqhhQYEO8_0),.clk(gclk));
	jdff dff_B_FIhTqrhf7_1(.din(n976),.dout(w_dff_B_FIhTqrhf7_1),.clk(gclk));
	jdff dff_A_RGJo87rH1_0(.dout(w_a114_0[0]),.din(w_dff_A_RGJo87rH1_0),.clk(gclk));
	jdff dff_A_4GIKWQI35_1(.dout(w_a115_0[1]),.din(w_dff_A_4GIKWQI35_1),.clk(gclk));
	jdff dff_B_745QdKaB0_1(.din(n894),.dout(w_dff_B_745QdKaB0_1),.clk(gclk));
	jdff dff_A_aqMYVpgr1_0(.dout(w_a112_0[0]),.din(w_dff_A_aqMYVpgr1_0),.clk(gclk));
	jdff dff_A_bKqOvwAI6_1(.dout(w_a113_0[1]),.din(w_dff_A_bKqOvwAI6_1),.clk(gclk));
	jdff dff_B_g2UrCknn7_1(.din(n956),.dout(w_dff_B_g2UrCknn7_1),.clk(gclk));
	jdff dff_A_SKaaili94_0(.dout(w_a122_0[0]),.din(w_dff_A_SKaaili94_0),.clk(gclk));
	jdff dff_A_nSHI3wrB2_1(.dout(w_a123_0[1]),.din(w_dff_A_nSHI3wrB2_1),.clk(gclk));
	jdff dff_B_K0Y4km6g5_1(.din(n962),.dout(w_dff_B_K0Y4km6g5_1),.clk(gclk));
	jdff dff_A_kGWQUzm74_0(.dout(w_a120_0[0]),.din(w_dff_A_kGWQUzm74_0),.clk(gclk));
	jdff dff_A_q0xtfwdX5_1(.dout(w_a121_0[1]),.din(w_dff_A_q0xtfwdX5_1),.clk(gclk));
	jdff dff_B_dyfUBpGV8_1(.din(n966),.dout(w_dff_B_dyfUBpGV8_1),.clk(gclk));
	jdff dff_A_lRhC755p2_0(.dout(w_a118_0[0]),.din(w_dff_A_lRhC755p2_0),.clk(gclk));
	jdff dff_A_ECSpmsBT6_1(.dout(w_a119_0[1]),.din(w_dff_A_ECSpmsBT6_1),.clk(gclk));
	jdff dff_B_sskXJKkD8_1(.din(n972),.dout(w_dff_B_sskXJKkD8_1),.clk(gclk));
	jdff dff_A_aEQEN3Xf2_0(.dout(w_a116_0[0]),.din(w_dff_A_aEQEN3Xf2_0),.clk(gclk));
	jdff dff_A_vTXKnj262_1(.dout(w_a117_0[1]),.din(w_dff_A_vTXKnj262_1),.clk(gclk));
	jdff dff_B_43V9h6ET3_1(.din(n987),.dout(w_dff_B_43V9h6ET3_1),.clk(gclk));
	jdff dff_A_2Aq7vbmA8_0(.dout(w_a126_0[0]),.din(w_dff_A_2Aq7vbmA8_0),.clk(gclk));
	jdff dff_A_OqgJmqtR1_1(.dout(w_a127_0[1]),.din(w_dff_A_OqgJmqtR1_1),.clk(gclk));
	jdff dff_B_rF98fik62_1(.din(n952),.dout(w_dff_B_rF98fik62_1),.clk(gclk));
	jdff dff_A_qYADieKW4_0(.dout(w_a124_0[0]),.din(w_dff_A_qYADieKW4_0),.clk(gclk));
	jdff dff_A_p4ahpbAJ4_1(.dout(w_a125_0[1]),.din(w_dff_A_p4ahpbAJ4_1),.clk(gclk));
	jdff dff_B_spBzN65s6_1(.din(n3021),.dout(w_dff_B_spBzN65s6_1),.clk(gclk));
	jdff dff_B_o6DVcVCt5_1(.din(w_dff_B_spBzN65s6_1),.dout(w_dff_B_o6DVcVCt5_1),.clk(gclk));
	jdff dff_B_ClAbqRb96_0(.din(n3025),.dout(w_dff_B_ClAbqRb96_0),.clk(gclk));
	jdff dff_B_aUU9y1mb9_1(.din(n2157),.dout(w_dff_B_aUU9y1mb9_1),.clk(gclk));
	jdff dff_B_uSl1DoMb4_1(.din(w_dff_B_aUU9y1mb9_1),.dout(w_dff_B_uSl1DoMb4_1),.clk(gclk));
	jdff dff_B_TnrR4rFy8_0(.din(n2161),.dout(w_dff_B_TnrR4rFy8_0),.clk(gclk));
	jdff dff_B_Np9QaPFa9_1(.din(n792),.dout(w_dff_B_Np9QaPFa9_1),.clk(gclk));
	jdff dff_A_hUN70b8y2_0(.dout(w_a44_0[0]),.din(w_dff_A_hUN70b8y2_0),.clk(gclk));
	jdff dff_A_dUrA3tEd2_1(.dout(w_a45_0[1]),.din(w_dff_A_dUrA3tEd2_1),.clk(gclk));
	jdff dff_B_PH0lI8405_1(.din(n807),.dout(w_dff_B_PH0lI8405_1),.clk(gclk));
	jdff dff_A_XF2Yyt4V5_0(.dout(w_a46_0[0]),.din(w_dff_A_XF2Yyt4V5_0),.clk(gclk));
	jdff dff_A_bTr2Cfs06_1(.dout(w_a47_0[1]),.din(w_dff_A_bTr2Cfs06_1),.clk(gclk));
	jdff dff_B_JkVSSvVk5_1(.din(n776),.dout(w_dff_B_JkVSSvVk5_1),.clk(gclk));
	jdff dff_A_4hVRVXx43_0(.dout(w_a34_0[0]),.din(w_dff_A_4hVRVXx43_0),.clk(gclk));
	jdff dff_A_IeX7m3QI0_1(.dout(w_a35_0[1]),.din(w_dff_A_IeX7m3QI0_1),.clk(gclk));
	jdff dff_B_tarZfy621_1(.din(n714),.dout(w_dff_B_tarZfy621_1),.clk(gclk));
	jdff dff_A_wkaxuBD72_0(.dout(w_a32_0[0]),.din(w_dff_A_wkaxuBD72_0),.clk(gclk));
	jdff dff_A_7OB6oRqA1_1(.dout(w_a33_0[1]),.din(w_dff_A_7OB6oRqA1_1),.clk(gclk));
	jdff dff_B_mYmJWWo27_1(.din(n782),.dout(w_dff_B_mYmJWWo27_1),.clk(gclk));
	jdff dff_A_we9q0Jad5_0(.dout(w_a38_0[0]),.din(w_dff_A_we9q0Jad5_0),.clk(gclk));
	jdff dff_A_VjN2Qliq0_1(.dout(w_a39_0[1]),.din(w_dff_A_VjN2Qliq0_1),.clk(gclk));
	jdff dff_B_sBdhvQYX3_1(.din(n772),.dout(w_dff_B_sBdhvQYX3_1),.clk(gclk));
	jdff dff_A_O8Ze6Upb1_0(.dout(w_a36_0[0]),.din(w_dff_A_O8Ze6Upb1_0),.clk(gclk));
	jdff dff_A_Z0uMSCcz9_1(.dout(w_a37_0[1]),.din(w_dff_A_Z0uMSCcz9_1),.clk(gclk));
	jdff dff_B_upysfaBQ0_1(.din(n796),.dout(w_dff_B_upysfaBQ0_1),.clk(gclk));
	jdff dff_A_VKlsC5cZ2_0(.dout(w_a42_0[0]),.din(w_dff_A_VKlsC5cZ2_0),.clk(gclk));
	jdff dff_A_Wwy7IlhU6_1(.dout(w_a43_0[1]),.din(w_dff_A_Wwy7IlhU6_1),.clk(gclk));
	jdff dff_B_1VoqRzDF0_1(.din(n786),.dout(w_dff_B_1VoqRzDF0_1),.clk(gclk));
	jdff dff_A_Dkax2EMe2_0(.dout(w_a40_0[0]),.din(w_dff_A_Dkax2EMe2_0),.clk(gclk));
	jdff dff_A_qtRk7Icw0_1(.dout(w_a41_0[1]),.din(w_dff_A_qtRk7Icw0_1),.clk(gclk));
	jdff dff_B_DMqPlBFe5_3(.din(n319),.dout(w_dff_B_DMqPlBFe5_3),.clk(gclk));
	jdff dff_B_jUEppjKS7_3(.din(w_dff_B_DMqPlBFe5_3),.dout(w_dff_B_jUEppjKS7_3),.clk(gclk));
	jdff dff_B_NzBHWWlV2_3(.din(w_dff_B_jUEppjKS7_3),.dout(w_dff_B_NzBHWWlV2_3),.clk(gclk));
	jdff dff_B_WUQO6yvK5_3(.din(w_dff_B_NzBHWWlV2_3),.dout(w_dff_B_WUQO6yvK5_3),.clk(gclk));
	jdff dff_B_inBTF3Cj2_3(.din(w_dff_B_WUQO6yvK5_3),.dout(w_dff_B_inBTF3Cj2_3),.clk(gclk));
	jdff dff_B_1nYZ6e8Z1_3(.din(w_dff_B_inBTF3Cj2_3),.dout(w_dff_B_1nYZ6e8Z1_3),.clk(gclk));
	jdff dff_B_ypPvMaYr6_3(.din(w_dff_B_1nYZ6e8Z1_3),.dout(w_dff_B_ypPvMaYr6_3),.clk(gclk));
	jdff dff_B_rk8XASRI6_1(.din(n2177),.dout(w_dff_B_rk8XASRI6_1),.clk(gclk));
	jdff dff_B_871fhSZh8_1(.din(w_dff_B_rk8XASRI6_1),.dout(w_dff_B_871fhSZh8_1),.clk(gclk));
	jdff dff_B_Ewoal9ki5_0(.din(n2181),.dout(w_dff_B_Ewoal9ki5_0),.clk(gclk));
	jdff dff_B_DGgUZnJK3_1(.din(n762),.dout(w_dff_B_DGgUZnJK3_1),.clk(gclk));
	jdff dff_A_rcrknBQy7_0(.dout(w_a10_0[0]),.din(w_dff_A_rcrknBQy7_0),.clk(gclk));
	jdff dff_A_PUmUpuIX0_1(.dout(w_a11_0[1]),.din(w_dff_A_PUmUpuIX0_1),.clk(gclk));
	jdff dff_B_uICq5SCD7_1(.din(n737),.dout(w_dff_B_uICq5SCD7_1),.clk(gclk));
	jdff dff_A_JPoE7RgR9_0(.dout(w_a8_0[0]),.din(w_dff_A_JPoE7RgR9_0),.clk(gclk));
	jdff dff_A_KS7aaRbG4_1(.dout(w_a9_0[1]),.din(w_dff_A_KS7aaRbG4_1),.clk(gclk));
	jdff dff_B_fsEUZG1w2_1(.din(n751),.dout(w_dff_B_fsEUZG1w2_1),.clk(gclk));
	jdff dff_A_JozpVLIs7_0(.dout(w_a2_0[0]),.din(w_dff_A_JozpVLIs7_0),.clk(gclk));
	jdff dff_A_P7ahRfJd1_1(.dout(w_a3_0[1]),.din(w_dff_A_P7ahRfJd1_1),.clk(gclk));
	jdff dff_B_Wz80cizW6_1(.din(n983),.dout(w_dff_B_Wz80cizW6_1),.clk(gclk));
	jdff dff_A_g47baKUj6_0(.dout(w_a0_0[0]),.din(w_dff_A_g47baKUj6_0),.clk(gclk));
	jdff dff_A_2LdNMFjs0_1(.dout(w_a1_0[1]),.din(w_dff_A_2LdNMFjs0_1),.clk(gclk));
	jdff dff_B_6YxyaqYr2_1(.din(n741),.dout(w_dff_B_6YxyaqYr2_1),.clk(gclk));
	jdff dff_A_5wvWWH0g3_0(.dout(w_a6_0[0]),.din(w_dff_A_5wvWWH0g3_0),.clk(gclk));
	jdff dff_A_2ewe9RPU2_1(.dout(w_a7_0[1]),.din(w_dff_A_2ewe9RPU2_1),.clk(gclk));
	jdff dff_B_aBi3tGKD9_1(.din(n747),.dout(w_dff_B_aBi3tGKD9_1),.clk(gclk));
	jdff dff_A_V7FH9gfr3_0(.dout(w_a4_0[0]),.din(w_dff_A_V7FH9gfr3_0),.clk(gclk));
	jdff dff_A_IhAADU2o4_1(.dout(w_a5_0[1]),.din(w_dff_A_IhAADU2o4_1),.clk(gclk));
	jdff dff_B_oi8DblKT5_1(.din(n731),.dout(w_dff_B_oi8DblKT5_1),.clk(gclk));
	jdff dff_A_aZ8WAfFs3_0(.dout(w_a14_0[0]),.din(w_dff_A_aZ8WAfFs3_0),.clk(gclk));
	jdff dff_A_jaLZbcNB9_1(.dout(w_a15_0[1]),.din(w_dff_A_jaLZbcNB9_1),.clk(gclk));
	jdff dff_B_h6051X5M0_1(.din(n758),.dout(w_dff_B_h6051X5M0_1),.clk(gclk));
	jdff dff_A_vcWxBCo84_0(.dout(w_a12_0[0]),.din(w_dff_A_vcWxBCo84_0),.clk(gclk));
	jdff dff_A_n7nis0rM6_1(.dout(w_a13_0[1]),.din(w_dff_A_n7nis0rM6_1),.clk(gclk));
	jdff dff_B_9BosVVVW8_3(.din(n410),.dout(w_dff_B_9BosVVVW8_3),.clk(gclk));
	jdff dff_B_y1OvB6m63_3(.din(w_dff_B_9BosVVVW8_3),.dout(w_dff_B_y1OvB6m63_3),.clk(gclk));
	jdff dff_B_pGhbj1re6_3(.din(w_dff_B_y1OvB6m63_3),.dout(w_dff_B_pGhbj1re6_3),.clk(gclk));
	jdff dff_B_e40Q35VS4_3(.din(w_dff_B_pGhbj1re6_3),.dout(w_dff_B_e40Q35VS4_3),.clk(gclk));
	jdff dff_B_qGUjWA5Y0_3(.din(w_dff_B_e40Q35VS4_3),.dout(w_dff_B_qGUjWA5Y0_3),.clk(gclk));
	jdff dff_B_NOMuLjAk2_3(.din(w_dff_B_qGUjWA5Y0_3),.dout(w_dff_B_NOMuLjAk2_3),.clk(gclk));
	jdff dff_B_EZWknVjS0_3(.din(w_dff_B_NOMuLjAk2_3),.dout(w_dff_B_EZWknVjS0_3),.clk(gclk));
	jdff dff_B_F1l9p9yf4_3(.din(w_dff_B_EZWknVjS0_3),.dout(w_dff_B_F1l9p9yf4_3),.clk(gclk));
	jdff dff_B_jTlFOYMo5_1(.din(n2149),.dout(w_dff_B_jTlFOYMo5_1),.clk(gclk));
	jdff dff_B_5fVocIcW4_1(.din(w_dff_B_jTlFOYMo5_1),.dout(w_dff_B_5fVocIcW4_1),.clk(gclk));
	jdff dff_B_sdDWXqfe3_0(.din(n2153),.dout(w_dff_B_sdDWXqfe3_0),.clk(gclk));
	jdff dff_B_Pj71flbm8_1(.din(n707),.dout(w_dff_B_Pj71flbm8_1),.clk(gclk));
	jdff dff_A_FL8rfjir2_0(.dout(w_a26_0[0]),.din(w_dff_A_FL8rfjir2_0),.clk(gclk));
	jdff dff_A_7GZZbsWq5_1(.dout(w_a27_0[1]),.din(w_dff_A_7GZZbsWq5_1),.clk(gclk));
	jdff dff_B_xpd5mGRp3_1(.din(n693),.dout(w_dff_B_xpd5mGRp3_1),.clk(gclk));
	jdff dff_A_JsBVmPGJ3_0(.dout(w_a24_0[0]),.din(w_dff_A_JsBVmPGJ3_0),.clk(gclk));
	jdff dff_A_LpS4cIVI1_1(.dout(w_a25_0[1]),.din(w_dff_A_LpS4cIVI1_1),.clk(gclk));
	jdff dff_B_MFGGkqzk7_1(.din(n687),.dout(w_dff_B_MFGGkqzk7_1),.clk(gclk));
	jdff dff_A_HqaVWGpG4_0(.dout(w_a18_0[0]),.din(w_dff_A_HqaVWGpG4_0),.clk(gclk));
	jdff dff_A_EfquT9R57_1(.dout(w_a19_0[1]),.din(w_dff_A_EfquT9R57_1),.clk(gclk));
	jdff dff_B_gXNcxvia2_1(.din(n727),.dout(w_dff_B_gXNcxvia2_1),.clk(gclk));
	jdff dff_A_6rr88UQ06_0(.dout(w_a16_0[0]),.din(w_dff_A_6rr88UQ06_0),.clk(gclk));
	jdff dff_A_IjOIf2Vv3_1(.dout(w_a17_0[1]),.din(w_dff_A_IjOIf2Vv3_1),.clk(gclk));
	jdff dff_B_o7JVhuzP9_1(.din(n697),.dout(w_dff_B_o7JVhuzP9_1),.clk(gclk));
	jdff dff_A_ypOJA4Mn4_0(.dout(w_a22_0[0]),.din(w_dff_A_ypOJA4Mn4_0),.clk(gclk));
	jdff dff_A_ECU7ndwr9_1(.dout(w_a23_0[1]),.din(w_dff_A_ECU7ndwr9_1),.clk(gclk));
	jdff dff_B_a5mabnqU6_1(.din(n683),.dout(w_dff_B_a5mabnqU6_1),.clk(gclk));
	jdff dff_A_z9RlMpd06_0(.dout(w_a20_0[0]),.din(w_dff_A_z9RlMpd06_0),.clk(gclk));
	jdff dff_A_OrPlTNw66_1(.dout(w_a21_0[1]),.din(w_dff_A_OrPlTNw66_1),.clk(gclk));
	jdff dff_B_DVmtjqsy4_1(.din(n718),.dout(w_dff_B_DVmtjqsy4_1),.clk(gclk));
	jdff dff_A_yNeInT2q0_0(.dout(w_a30_0[0]),.din(w_dff_A_yNeInT2q0_0),.clk(gclk));
	jdff dff_A_yjHZSHH70_1(.dout(w_a31_0[1]),.din(w_dff_A_yjHZSHH70_1),.clk(gclk));
	jdff dff_B_TF8VuoJz5_1(.din(n703),.dout(w_dff_B_TF8VuoJz5_1),.clk(gclk));
	jdff dff_A_ixqoCv1I6_0(.dout(w_a28_0[0]),.din(w_dff_A_ixqoCv1I6_0),.clk(gclk));
	jdff dff_A_AvFtfhSE5_1(.dout(w_a29_0[1]),.din(w_dff_A_AvFtfhSE5_1),.clk(gclk));
	jdff dff_B_CxYsv1cW2_3(.din(n265),.dout(w_dff_B_CxYsv1cW2_3),.clk(gclk));
	jdff dff_B_qeWyi0A84_3(.din(w_dff_B_CxYsv1cW2_3),.dout(w_dff_B_qeWyi0A84_3),.clk(gclk));
	jdff dff_B_81YZhcyd8_3(.din(w_dff_B_qeWyi0A84_3),.dout(w_dff_B_81YZhcyd8_3),.clk(gclk));
	jdff dff_B_KLxrtH251_3(.din(w_dff_B_81YZhcyd8_3),.dout(w_dff_B_KLxrtH251_3),.clk(gclk));
	jdff dff_B_1oN0NPYh2_3(.din(w_dff_B_KLxrtH251_3),.dout(w_dff_B_1oN0NPYh2_3),.clk(gclk));
	jdff dff_B_FM0LHf2p9_3(.din(w_dff_B_1oN0NPYh2_3),.dout(w_dff_B_FM0LHf2p9_3),.clk(gclk));
	jdff dff_B_eLdE6Tba8_3(.din(w_dff_B_FM0LHf2p9_3),.dout(w_dff_B_eLdE6Tba8_3),.clk(gclk));
	jdff dff_B_2BfiXtTV3_1(.din(n2141),.dout(w_dff_B_2BfiXtTV3_1),.clk(gclk));
	jdff dff_B_wKhuxg1O7_1(.din(w_dff_B_2BfiXtTV3_1),.dout(w_dff_B_wKhuxg1O7_1),.clk(gclk));
	jdff dff_B_sFr9dA5r6_0(.din(n2145),.dout(w_dff_B_sFr9dA5r6_0),.clk(gclk));
	jdff dff_B_v2guYC8y6_1(.din(n674),.dout(w_dff_B_v2guYC8y6_1),.clk(gclk));
	jdff dff_A_HmdqNm8g4_0(.dout(w_a62_0[0]),.din(w_dff_A_HmdqNm8g4_0),.clk(gclk));
	jdff dff_A_8mgBZIQg7_1(.dout(w_a63_0[1]),.din(w_dff_A_8mgBZIQg7_1),.clk(gclk));
	jdff dff_B_0oLZnUPh4_1(.din(n639),.dout(w_dff_B_0oLZnUPh4_1),.clk(gclk));
	jdff dff_A_ruJEv85L7_0(.dout(w_a60_0[0]),.din(w_dff_A_ruJEv85L7_0),.clk(gclk));
	jdff dff_A_zbNXoOqW6_1(.dout(w_a61_0[1]),.din(w_dff_A_zbNXoOqW6_1),.clk(gclk));
	jdff dff_B_T6FhMLOl0_3(.din(n304),.dout(w_dff_B_T6FhMLOl0_3),.clk(gclk));
	jdff dff_B_2lyKqjFZ9_3(.din(w_dff_B_T6FhMLOl0_3),.dout(w_dff_B_2lyKqjFZ9_3),.clk(gclk));
	jdff dff_B_L3XqwQjn4_3(.din(w_dff_B_2lyKqjFZ9_3),.dout(w_dff_B_L3XqwQjn4_3),.clk(gclk));
	jdff dff_B_PK6M6bQk2_1(.din(n663),.dout(w_dff_B_PK6M6bQk2_1),.clk(gclk));
	jdff dff_A_qerx9cuT9_0(.dout(w_a50_0[0]),.din(w_dff_A_qerx9cuT9_0),.clk(gclk));
	jdff dff_A_MCBIUaBq2_1(.dout(w_a51_0[1]),.din(w_dff_A_MCBIUaBq2_1),.clk(gclk));
	jdff dff_B_YqCEMGkj8_1(.din(n803),.dout(w_dff_B_YqCEMGkj8_1),.clk(gclk));
	jdff dff_A_x9iScKCA1_0(.dout(w_a48_0[0]),.din(w_dff_A_x9iScKCA1_0),.clk(gclk));
	jdff dff_A_mAgVgHU16_1(.dout(w_a49_0[1]),.din(w_dff_A_mAgVgHU16_1),.clk(gclk));
	jdff dff_B_3n7FITo24_3(.din(n292),.dout(w_dff_B_3n7FITo24_3),.clk(gclk));
	jdff dff_B_2lzJbilg4_3(.din(w_dff_B_3n7FITo24_3),.dout(w_dff_B_2lzJbilg4_3),.clk(gclk));
	jdff dff_B_bi8l2YH76_3(.din(w_dff_B_2lzJbilg4_3),.dout(w_dff_B_bi8l2YH76_3),.clk(gclk));
	jdff dff_B_H2R9KPX95_3(.din(w_dff_B_bi8l2YH76_3),.dout(w_dff_B_H2R9KPX95_3),.clk(gclk));
	jdff dff_B_tfJFhTxG8_1(.din(n653),.dout(w_dff_B_tfJFhTxG8_1),.clk(gclk));
	jdff dff_A_xNYvrMCm0_0(.dout(w_a54_0[0]),.din(w_dff_A_xNYvrMCm0_0),.clk(gclk));
	jdff dff_A_0nnYYHF55_1(.dout(w_a55_0[1]),.din(w_dff_A_0nnYYHF55_1),.clk(gclk));
	jdff dff_B_SLXi6sqx0_1(.din(n659),.dout(w_dff_B_SLXi6sqx0_1),.clk(gclk));
	jdff dff_A_TEmwG3XJ6_0(.dout(w_a52_0[0]),.din(w_dff_A_TEmwG3XJ6_0),.clk(gclk));
	jdff dff_A_r5bZU0Yn6_1(.dout(w_a53_0[1]),.din(w_dff_A_r5bZU0Yn6_1),.clk(gclk));
	jdff dff_B_x2mt324E2_3(.din(n281),.dout(w_dff_B_x2mt324E2_3),.clk(gclk));
	jdff dff_B_rnaB24hv3_3(.din(w_dff_B_x2mt324E2_3),.dout(w_dff_B_rnaB24hv3_3),.clk(gclk));
	jdff dff_B_FULzpxU81_3(.din(w_dff_B_rnaB24hv3_3),.dout(w_dff_B_FULzpxU81_3),.clk(gclk));
	jdff dff_B_HKuzR6c52_1(.din(n643),.dout(w_dff_B_HKuzR6c52_1),.clk(gclk));
	jdff dff_A_AY4LJMyP2_0(.dout(w_a58_0[0]),.din(w_dff_A_AY4LJMyP2_0),.clk(gclk));
	jdff dff_A_td3IjRBo8_1(.dout(w_a59_0[1]),.din(w_dff_A_td3IjRBo8_1),.clk(gclk));
	jdff dff_B_5jw3Llau0_3(.din(n273),.dout(w_dff_B_5jw3Llau0_3),.clk(gclk));
	jdff dff_B_AMEaIxgs6_3(.din(w_dff_B_5jw3Llau0_3),.dout(w_dff_B_AMEaIxgs6_3),.clk(gclk));
	jdff dff_A_e2KaJXa04_0(.dout(w_shift1_63[0]),.din(w_dff_A_e2KaJXa04_0),.clk(gclk));
	jdff dff_A_vpG9IxaZ1_0(.dout(w_dff_A_e2KaJXa04_0),.din(w_dff_A_vpG9IxaZ1_0),.clk(gclk));
	jdff dff_A_hDIMdffy1_0(.dout(w_dff_A_vpG9IxaZ1_0),.din(w_dff_A_hDIMdffy1_0),.clk(gclk));
	jdff dff_A_1Z7k3zc65_2(.dout(w_shift1_63[2]),.din(w_dff_A_1Z7k3zc65_2),.clk(gclk));
	jdff dff_A_OmMWeXIQ2_2(.dout(w_dff_A_1Z7k3zc65_2),.din(w_dff_A_OmMWeXIQ2_2),.clk(gclk));
	jdff dff_A_bMqTrhbp3_2(.dout(w_dff_A_OmMWeXIQ2_2),.din(w_dff_A_bMqTrhbp3_2),.clk(gclk));
	jdff dff_A_RC8wWg7O0_0(.dout(w_shift1_20[0]),.din(w_dff_A_RC8wWg7O0_0),.clk(gclk));
	jdff dff_A_hcEVGi5I5_0(.dout(w_dff_A_RC8wWg7O0_0),.din(w_dff_A_hcEVGi5I5_0),.clk(gclk));
	jdff dff_A_9kI7kVaC9_0(.dout(w_dff_A_hcEVGi5I5_0),.din(w_dff_A_9kI7kVaC9_0),.clk(gclk));
	jdff dff_A_ATtTd43D2_1(.dout(w_shift1_20[1]),.din(w_dff_A_ATtTd43D2_1),.clk(gclk));
	jdff dff_A_VgBYN22x4_1(.dout(w_dff_A_ATtTd43D2_1),.din(w_dff_A_VgBYN22x4_1),.clk(gclk));
	jdff dff_A_rtDyqCOd8_1(.dout(w_dff_A_VgBYN22x4_1),.din(w_dff_A_rtDyqCOd8_1),.clk(gclk));
	jdff dff_A_aJMy0lZt4_0(.dout(w_shift1_6[0]),.din(w_dff_A_aJMy0lZt4_0),.clk(gclk));
	jdff dff_A_1KxTcwcD2_0(.dout(w_dff_A_aJMy0lZt4_0),.din(w_dff_A_1KxTcwcD2_0),.clk(gclk));
	jdff dff_A_imsCNVkT2_0(.dout(w_dff_A_1KxTcwcD2_0),.din(w_dff_A_imsCNVkT2_0),.clk(gclk));
	jdff dff_A_MyYUwFlP4_2(.dout(w_shift1_6[2]),.din(w_dff_A_MyYUwFlP4_2),.clk(gclk));
	jdff dff_A_dyImM1rh4_2(.dout(w_dff_A_MyYUwFlP4_2),.din(w_dff_A_dyImM1rh4_2),.clk(gclk));
	jdff dff_A_mDIUIck97_2(.dout(w_dff_A_dyImM1rh4_2),.din(w_dff_A_mDIUIck97_2),.clk(gclk));
	jdff dff_A_88LexBq42_0(.dout(w_shift1_1[0]),.din(w_dff_A_88LexBq42_0),.clk(gclk));
	jdff dff_A_NqFXEflt2_0(.dout(w_dff_A_88LexBq42_0),.din(w_dff_A_NqFXEflt2_0),.clk(gclk));
	jdff dff_A_VLfOiBZL1_0(.dout(w_dff_A_NqFXEflt2_0),.din(w_dff_A_VLfOiBZL1_0),.clk(gclk));
	jdff dff_A_zcodIgwo3_1(.dout(w_shift1_1[1]),.din(w_dff_A_zcodIgwo3_1),.clk(gclk));
	jdff dff_A_anpED3qE4_1(.dout(w_dff_A_zcodIgwo3_1),.din(w_dff_A_anpED3qE4_1),.clk(gclk));
	jdff dff_A_LfupF43K8_1(.dout(w_dff_A_anpED3qE4_1),.din(w_dff_A_LfupF43K8_1),.clk(gclk));
	jdff dff_B_innup2oD0_1(.din(n649),.dout(w_dff_B_innup2oD0_1),.clk(gclk));
	jdff dff_A_Nsc29slm7_0(.dout(w_a56_0[0]),.din(w_dff_A_Nsc29slm7_0),.clk(gclk));
	jdff dff_A_S63Jgp8X2_1(.dout(w_a57_0[1]),.din(w_dff_A_S63Jgp8X2_1),.clk(gclk));
	jdff dff_A_FxTfk7bY2_1(.dout(w_shift1_0[1]),.din(w_dff_A_FxTfk7bY2_1),.clk(gclk));
	jdff dff_A_MOLsVTew2_1(.dout(w_dff_A_FxTfk7bY2_1),.din(w_dff_A_MOLsVTew2_1),.clk(gclk));
	jdff dff_A_2auC8Ory6_1(.dout(w_dff_A_MOLsVTew2_1),.din(w_dff_A_2auC8Ory6_1),.clk(gclk));
	jdff dff_A_4rP6ARZQ0_2(.dout(w_shift1_0[2]),.din(w_dff_A_4rP6ARZQ0_2),.clk(gclk));
	jdff dff_A_Mwoc0Tgp8_2(.dout(w_dff_A_4rP6ARZQ0_2),.din(w_dff_A_Mwoc0Tgp8_2),.clk(gclk));
	jdff dff_A_ewMNBLer3_2(.dout(w_dff_A_Mwoc0Tgp8_2),.din(w_dff_A_ewMNBLer3_2),.clk(gclk));
	jdff dff_B_3XLTqWEN0_3(.din(n267),.dout(w_dff_B_3XLTqWEN0_3),.clk(gclk));
	jdff dff_B_mkxpvy5v7_3(.din(w_dff_B_3XLTqWEN0_3),.dout(w_dff_B_mkxpvy5v7_3),.clk(gclk));
	jdff dff_B_BzJqvu7e0_3(.din(w_dff_B_mkxpvy5v7_3),.dout(w_dff_B_BzJqvu7e0_3),.clk(gclk));
	jdff dff_A_6q7NhxpC3_1(.dout(w_shift3_0[1]),.din(w_dff_A_6q7NhxpC3_1),.clk(gclk));
	jdff dff_A_iZkaQ2vc3_2(.dout(w_shift2_0[2]),.din(w_dff_A_iZkaQ2vc3_2),.clk(gclk));
	jdff dff_B_cWtJz30h3_3(.din(n364),.dout(w_dff_B_cWtJz30h3_3),.clk(gclk));
	jdff dff_B_JG7qnRyB1_3(.din(w_dff_B_cWtJz30h3_3),.dout(w_dff_B_JG7qnRyB1_3),.clk(gclk));
	jdff dff_B_odhJBSIE1_3(.din(w_dff_B_JG7qnRyB1_3),.dout(w_dff_B_odhJBSIE1_3),.clk(gclk));
	jdff dff_B_7rQcpyIn7_3(.din(w_dff_B_odhJBSIE1_3),.dout(w_dff_B_7rQcpyIn7_3),.clk(gclk));
	jdff dff_B_TNFpLTFg8_3(.din(w_dff_B_7rQcpyIn7_3),.dout(w_dff_B_TNFpLTFg8_3),.clk(gclk));
	jdff dff_B_zRdqDAAF6_3(.din(w_dff_B_TNFpLTFg8_3),.dout(w_dff_B_zRdqDAAF6_3),.clk(gclk));
	jdff dff_B_cE1lYXHF5_3(.din(w_dff_B_zRdqDAAF6_3),.dout(w_dff_B_cE1lYXHF5_3),.clk(gclk));
	jdff dff_A_6JmKMWA78_2(.dout(w_shift5_0[2]),.din(w_dff_A_6JmKMWA78_2),.clk(gclk));
	jdff dff_A_kHgVQNIK1_1(.dout(w_shift4_0[1]),.din(w_dff_A_kHgVQNIK1_1),.clk(gclk));
	jdff dff_B_D1MyPfrQ5_3(.din(n263),.dout(w_dff_B_D1MyPfrQ5_3),.clk(gclk));
	jdff dff_B_TlEknDsx1_3(.din(w_dff_B_D1MyPfrQ5_3),.dout(w_dff_B_TlEknDsx1_3),.clk(gclk));
	jdff dff_B_7lDjzph70_3(.din(w_dff_B_TlEknDsx1_3),.dout(w_dff_B_7lDjzph70_3),.clk(gclk));
	jdff dff_B_rFdjlMZD1_3(.din(w_dff_B_7lDjzph70_3),.dout(w_dff_B_rFdjlMZD1_3),.clk(gclk));
	jdff dff_B_cpeRMzaJ8_3(.din(w_dff_B_rFdjlMZD1_3),.dout(w_dff_B_cpeRMzaJ8_3),.clk(gclk));
	jdff dff_B_ZPRNw5ou6_3(.din(w_dff_B_cpeRMzaJ8_3),.dout(w_dff_B_ZPRNw5ou6_3),.clk(gclk));
	jdff dff_B_LUTSYlbD1_3(.din(w_dff_B_ZPRNw5ou6_3),.dout(w_dff_B_LUTSYlbD1_3),.clk(gclk));
	jdff dff_B_SchMfHZx3_3(.din(w_dff_B_LUTSYlbD1_3),.dout(w_dff_B_SchMfHZx3_3),.clk(gclk));
	jdff dff_B_lPjXFL1b0_3(.din(w_dff_B_SchMfHZx3_3),.dout(w_dff_B_lPjXFL1b0_3),.clk(gclk));
	jdff dff_B_rFFecGf23_3(.din(w_dff_B_lPjXFL1b0_3),.dout(w_dff_B_rFFecGf23_3),.clk(gclk));
	jdff dff_B_wnnGE9y38_3(.din(w_dff_B_rFFecGf23_3),.dout(w_dff_B_wnnGE9y38_3),.clk(gclk));
	jdff dff_B_auwam0s87_3(.din(w_dff_B_wnnGE9y38_3),.dout(w_dff_B_auwam0s87_3),.clk(gclk));
	jdff dff_A_yAJH0Bn31_0(.dout(w_shift6_63[0]),.din(w_dff_A_yAJH0Bn31_0),.clk(gclk));
	jdff dff_A_UgEDVB5a1_0(.dout(w_dff_A_yAJH0Bn31_0),.din(w_dff_A_UgEDVB5a1_0),.clk(gclk));
	jdff dff_A_cXfHOD8n6_0(.dout(w_dff_A_UgEDVB5a1_0),.din(w_dff_A_cXfHOD8n6_0),.clk(gclk));
	jdff dff_A_BJ1qMqCb1_0(.dout(w_dff_A_cXfHOD8n6_0),.din(w_dff_A_BJ1qMqCb1_0),.clk(gclk));
	jdff dff_A_KvzloDZH6_0(.dout(w_dff_A_BJ1qMqCb1_0),.din(w_dff_A_KvzloDZH6_0),.clk(gclk));
	jdff dff_A_DlfBdeCe3_0(.dout(w_dff_A_KvzloDZH6_0),.din(w_dff_A_DlfBdeCe3_0),.clk(gclk));
	jdff dff_A_Mw1W6pyL3_0(.dout(w_dff_A_DlfBdeCe3_0),.din(w_dff_A_Mw1W6pyL3_0),.clk(gclk));
	jdff dff_A_7I6ciW9d6_0(.dout(w_dff_A_Mw1W6pyL3_0),.din(w_dff_A_7I6ciW9d6_0),.clk(gclk));
	jdff dff_A_k0l05ikN7_0(.dout(w_dff_A_7I6ciW9d6_0),.din(w_dff_A_k0l05ikN7_0),.clk(gclk));
	jdff dff_A_8CG9Zvle8_0(.dout(w_dff_A_k0l05ikN7_0),.din(w_dff_A_8CG9Zvle8_0),.clk(gclk));
	jdff dff_A_O19qIvxa8_0(.dout(w_dff_A_8CG9Zvle8_0),.din(w_dff_A_O19qIvxa8_0),.clk(gclk));
	jdff dff_A_1lSULzdc6_0(.dout(w_dff_A_O19qIvxa8_0),.din(w_dff_A_1lSULzdc6_0),.clk(gclk));
	jdff dff_A_bqhDMCvs6_0(.dout(w_dff_A_1lSULzdc6_0),.din(w_dff_A_bqhDMCvs6_0),.clk(gclk));
	jdff dff_A_asXnvvCp1_1(.dout(w_shift6_63[1]),.din(w_dff_A_asXnvvCp1_1),.clk(gclk));
	jdff dff_A_7MV0wofZ2_1(.dout(w_dff_A_asXnvvCp1_1),.din(w_dff_A_7MV0wofZ2_1),.clk(gclk));
	jdff dff_A_YYodgnKE3_1(.dout(w_dff_A_7MV0wofZ2_1),.din(w_dff_A_YYodgnKE3_1),.clk(gclk));
	jdff dff_A_OAQAKcMT7_1(.dout(w_dff_A_YYodgnKE3_1),.din(w_dff_A_OAQAKcMT7_1),.clk(gclk));
	jdff dff_A_a6OmcwGy4_1(.dout(w_dff_A_OAQAKcMT7_1),.din(w_dff_A_a6OmcwGy4_1),.clk(gclk));
	jdff dff_A_7awDuIx24_1(.dout(w_dff_A_a6OmcwGy4_1),.din(w_dff_A_7awDuIx24_1),.clk(gclk));
	jdff dff_A_zHovBbBN9_1(.dout(w_dff_A_7awDuIx24_1),.din(w_dff_A_zHovBbBN9_1),.clk(gclk));
	jdff dff_A_GEHCN80u4_1(.dout(w_dff_A_zHovBbBN9_1),.din(w_dff_A_GEHCN80u4_1),.clk(gclk));
	jdff dff_A_5v7paUrI6_1(.dout(w_dff_A_GEHCN80u4_1),.din(w_dff_A_5v7paUrI6_1),.clk(gclk));
	jdff dff_A_gm71wfmI4_1(.dout(w_dff_A_5v7paUrI6_1),.din(w_dff_A_gm71wfmI4_1),.clk(gclk));
	jdff dff_A_rlnw4zxw4_1(.dout(w_dff_A_gm71wfmI4_1),.din(w_dff_A_rlnw4zxw4_1),.clk(gclk));
	jdff dff_A_ntqqrbQY5_1(.dout(w_dff_A_rlnw4zxw4_1),.din(w_dff_A_ntqqrbQY5_1),.clk(gclk));
	jdff dff_A_QEbkLJAp3_1(.dout(w_dff_A_ntqqrbQY5_1),.din(w_dff_A_QEbkLJAp3_1),.clk(gclk));
	jdff dff_A_yTLlrHtH8_0(.dout(w_shift6_20[0]),.din(w_dff_A_yTLlrHtH8_0),.clk(gclk));
	jdff dff_A_6WbT2UZz4_0(.dout(w_dff_A_yTLlrHtH8_0),.din(w_dff_A_6WbT2UZz4_0),.clk(gclk));
	jdff dff_A_s0Zks23c4_0(.dout(w_dff_A_6WbT2UZz4_0),.din(w_dff_A_s0Zks23c4_0),.clk(gclk));
	jdff dff_A_KVbybT3z0_0(.dout(w_dff_A_s0Zks23c4_0),.din(w_dff_A_KVbybT3z0_0),.clk(gclk));
	jdff dff_A_sUerBJWF3_0(.dout(w_dff_A_KVbybT3z0_0),.din(w_dff_A_sUerBJWF3_0),.clk(gclk));
	jdff dff_A_KwRqLfUv4_0(.dout(w_dff_A_sUerBJWF3_0),.din(w_dff_A_KwRqLfUv4_0),.clk(gclk));
	jdff dff_A_MPQc3Pdx9_0(.dout(w_dff_A_KwRqLfUv4_0),.din(w_dff_A_MPQc3Pdx9_0),.clk(gclk));
	jdff dff_A_kc3JFFaF5_0(.dout(w_dff_A_MPQc3Pdx9_0),.din(w_dff_A_kc3JFFaF5_0),.clk(gclk));
	jdff dff_A_kDlzFewf6_0(.dout(w_dff_A_kc3JFFaF5_0),.din(w_dff_A_kDlzFewf6_0),.clk(gclk));
	jdff dff_A_RtiDpvgr1_0(.dout(w_dff_A_kDlzFewf6_0),.din(w_dff_A_RtiDpvgr1_0),.clk(gclk));
	jdff dff_A_Fex9r6ri9_0(.dout(w_dff_A_RtiDpvgr1_0),.din(w_dff_A_Fex9r6ri9_0),.clk(gclk));
	jdff dff_A_wIe7t5VD4_0(.dout(w_dff_A_Fex9r6ri9_0),.din(w_dff_A_wIe7t5VD4_0),.clk(gclk));
	jdff dff_A_SkPkN92h4_0(.dout(w_dff_A_wIe7t5VD4_0),.din(w_dff_A_SkPkN92h4_0),.clk(gclk));
	jdff dff_A_VI5eUidT5_1(.dout(w_shift6_20[1]),.din(w_dff_A_VI5eUidT5_1),.clk(gclk));
	jdff dff_A_NWadLbxG1_1(.dout(w_dff_A_VI5eUidT5_1),.din(w_dff_A_NWadLbxG1_1),.clk(gclk));
	jdff dff_A_zqTuj6v83_1(.dout(w_dff_A_NWadLbxG1_1),.din(w_dff_A_zqTuj6v83_1),.clk(gclk));
	jdff dff_A_peXhlYT34_1(.dout(w_dff_A_zqTuj6v83_1),.din(w_dff_A_peXhlYT34_1),.clk(gclk));
	jdff dff_A_7giuYgW11_1(.dout(w_dff_A_peXhlYT34_1),.din(w_dff_A_7giuYgW11_1),.clk(gclk));
	jdff dff_A_Sg3rSI1a8_1(.dout(w_dff_A_7giuYgW11_1),.din(w_dff_A_Sg3rSI1a8_1),.clk(gclk));
	jdff dff_A_FWlwrulx5_1(.dout(w_dff_A_Sg3rSI1a8_1),.din(w_dff_A_FWlwrulx5_1),.clk(gclk));
	jdff dff_A_kFQVZGOf6_1(.dout(w_dff_A_FWlwrulx5_1),.din(w_dff_A_kFQVZGOf6_1),.clk(gclk));
	jdff dff_A_gMPxVi5q6_1(.dout(w_dff_A_kFQVZGOf6_1),.din(w_dff_A_gMPxVi5q6_1),.clk(gclk));
	jdff dff_A_aWYGTbjE2_1(.dout(w_dff_A_gMPxVi5q6_1),.din(w_dff_A_aWYGTbjE2_1),.clk(gclk));
	jdff dff_A_xz481dg06_1(.dout(w_dff_A_aWYGTbjE2_1),.din(w_dff_A_xz481dg06_1),.clk(gclk));
	jdff dff_A_9TqyH9XI9_1(.dout(w_dff_A_xz481dg06_1),.din(w_dff_A_9TqyH9XI9_1),.clk(gclk));
	jdff dff_A_GnocIZ4d7_1(.dout(w_dff_A_9TqyH9XI9_1),.din(w_dff_A_GnocIZ4d7_1),.clk(gclk));
	jdff dff_A_CxgjtJf25_0(.dout(w_shift6_6[0]),.din(w_dff_A_CxgjtJf25_0),.clk(gclk));
	jdff dff_A_aqwxP7733_0(.dout(w_dff_A_CxgjtJf25_0),.din(w_dff_A_aqwxP7733_0),.clk(gclk));
	jdff dff_A_QaxrS6Bk7_0(.dout(w_dff_A_aqwxP7733_0),.din(w_dff_A_QaxrS6Bk7_0),.clk(gclk));
	jdff dff_A_QR95RoFe4_0(.dout(w_dff_A_QaxrS6Bk7_0),.din(w_dff_A_QR95RoFe4_0),.clk(gclk));
	jdff dff_A_zc0yCe6x6_0(.dout(w_dff_A_QR95RoFe4_0),.din(w_dff_A_zc0yCe6x6_0),.clk(gclk));
	jdff dff_A_ds5wZAaK9_0(.dout(w_dff_A_zc0yCe6x6_0),.din(w_dff_A_ds5wZAaK9_0),.clk(gclk));
	jdff dff_A_JHwHU07f3_0(.dout(w_dff_A_ds5wZAaK9_0),.din(w_dff_A_JHwHU07f3_0),.clk(gclk));
	jdff dff_A_tQvjFbhx2_0(.dout(w_dff_A_JHwHU07f3_0),.din(w_dff_A_tQvjFbhx2_0),.clk(gclk));
	jdff dff_A_7l4ZZ3Oy4_0(.dout(w_dff_A_tQvjFbhx2_0),.din(w_dff_A_7l4ZZ3Oy4_0),.clk(gclk));
	jdff dff_A_JJ01ICRq4_0(.dout(w_dff_A_7l4ZZ3Oy4_0),.din(w_dff_A_JJ01ICRq4_0),.clk(gclk));
	jdff dff_A_eYY6o3js5_0(.dout(w_dff_A_JJ01ICRq4_0),.din(w_dff_A_eYY6o3js5_0),.clk(gclk));
	jdff dff_A_QMLCc8ja8_0(.dout(w_dff_A_eYY6o3js5_0),.din(w_dff_A_QMLCc8ja8_0),.clk(gclk));
	jdff dff_A_ilrk8ITG9_0(.dout(w_dff_A_QMLCc8ja8_0),.din(w_dff_A_ilrk8ITG9_0),.clk(gclk));
	jdff dff_A_9KEoRETL5_2(.dout(w_shift6_6[2]),.din(w_dff_A_9KEoRETL5_2),.clk(gclk));
	jdff dff_A_xQz8WY0T2_2(.dout(w_dff_A_9KEoRETL5_2),.din(w_dff_A_xQz8WY0T2_2),.clk(gclk));
	jdff dff_A_VqmGKOO02_2(.dout(w_dff_A_xQz8WY0T2_2),.din(w_dff_A_VqmGKOO02_2),.clk(gclk));
	jdff dff_A_Hgg1ozR90_2(.dout(w_dff_A_VqmGKOO02_2),.din(w_dff_A_Hgg1ozR90_2),.clk(gclk));
	jdff dff_A_wQQikEXv7_2(.dout(w_dff_A_Hgg1ozR90_2),.din(w_dff_A_wQQikEXv7_2),.clk(gclk));
	jdff dff_A_mf1pd0do8_2(.dout(w_dff_A_wQQikEXv7_2),.din(w_dff_A_mf1pd0do8_2),.clk(gclk));
	jdff dff_A_B4U2IVCW5_2(.dout(w_dff_A_mf1pd0do8_2),.din(w_dff_A_B4U2IVCW5_2),.clk(gclk));
	jdff dff_A_WzNzoCIq5_2(.dout(w_dff_A_B4U2IVCW5_2),.din(w_dff_A_WzNzoCIq5_2),.clk(gclk));
	jdff dff_A_50ekwJrz5_2(.dout(w_dff_A_WzNzoCIq5_2),.din(w_dff_A_50ekwJrz5_2),.clk(gclk));
	jdff dff_A_YxGiN22x4_2(.dout(w_dff_A_50ekwJrz5_2),.din(w_dff_A_YxGiN22x4_2),.clk(gclk));
	jdff dff_A_Ly6xRXqK6_2(.dout(w_dff_A_YxGiN22x4_2),.din(w_dff_A_Ly6xRXqK6_2),.clk(gclk));
	jdff dff_A_uudtF6AE7_2(.dout(w_dff_A_Ly6xRXqK6_2),.din(w_dff_A_uudtF6AE7_2),.clk(gclk));
	jdff dff_A_NGTUJztT7_2(.dout(w_dff_A_uudtF6AE7_2),.din(w_dff_A_NGTUJztT7_2),.clk(gclk));
	jdff dff_A_OEfCsjIo7_0(.dout(w_shift6_1[0]),.din(w_dff_A_OEfCsjIo7_0),.clk(gclk));
	jdff dff_A_moDPj9Iq5_0(.dout(w_dff_A_OEfCsjIo7_0),.din(w_dff_A_moDPj9Iq5_0),.clk(gclk));
	jdff dff_A_ltgJltH36_0(.dout(w_dff_A_moDPj9Iq5_0),.din(w_dff_A_ltgJltH36_0),.clk(gclk));
	jdff dff_A_sb6j7kem3_0(.dout(w_dff_A_ltgJltH36_0),.din(w_dff_A_sb6j7kem3_0),.clk(gclk));
	jdff dff_A_iQ2BsceM8_0(.dout(w_dff_A_sb6j7kem3_0),.din(w_dff_A_iQ2BsceM8_0),.clk(gclk));
	jdff dff_A_5sYHyqNT2_0(.dout(w_dff_A_iQ2BsceM8_0),.din(w_dff_A_5sYHyqNT2_0),.clk(gclk));
	jdff dff_A_KFLXylHK7_0(.dout(w_dff_A_5sYHyqNT2_0),.din(w_dff_A_KFLXylHK7_0),.clk(gclk));
	jdff dff_A_bLaMM5ge3_0(.dout(w_dff_A_KFLXylHK7_0),.din(w_dff_A_bLaMM5ge3_0),.clk(gclk));
	jdff dff_A_tFBeomrf2_0(.dout(w_dff_A_bLaMM5ge3_0),.din(w_dff_A_tFBeomrf2_0),.clk(gclk));
	jdff dff_A_RfTcGk5e1_0(.dout(w_dff_A_tFBeomrf2_0),.din(w_dff_A_RfTcGk5e1_0),.clk(gclk));
	jdff dff_A_SG4k4aTM0_0(.dout(w_dff_A_RfTcGk5e1_0),.din(w_dff_A_SG4k4aTM0_0),.clk(gclk));
	jdff dff_A_7akYvcM92_0(.dout(w_dff_A_SG4k4aTM0_0),.din(w_dff_A_7akYvcM92_0),.clk(gclk));
	jdff dff_A_LF7uoH3p0_0(.dout(w_dff_A_7akYvcM92_0),.din(w_dff_A_LF7uoH3p0_0),.clk(gclk));
	jdff dff_A_OYJcZjJL1_1(.dout(w_shift6_1[1]),.din(w_dff_A_OYJcZjJL1_1),.clk(gclk));
	jdff dff_A_wsTqhXUy8_1(.dout(w_dff_A_OYJcZjJL1_1),.din(w_dff_A_wsTqhXUy8_1),.clk(gclk));
	jdff dff_A_OsgiMFyk8_1(.dout(w_dff_A_wsTqhXUy8_1),.din(w_dff_A_OsgiMFyk8_1),.clk(gclk));
	jdff dff_A_3UlkHgJ53_1(.dout(w_dff_A_OsgiMFyk8_1),.din(w_dff_A_3UlkHgJ53_1),.clk(gclk));
	jdff dff_A_qpXxM72y4_1(.dout(w_dff_A_3UlkHgJ53_1),.din(w_dff_A_qpXxM72y4_1),.clk(gclk));
	jdff dff_A_INOTK3000_1(.dout(w_dff_A_qpXxM72y4_1),.din(w_dff_A_INOTK3000_1),.clk(gclk));
	jdff dff_A_c48fOM751_1(.dout(w_dff_A_INOTK3000_1),.din(w_dff_A_c48fOM751_1),.clk(gclk));
	jdff dff_A_yIPwSEAS6_1(.dout(w_dff_A_c48fOM751_1),.din(w_dff_A_yIPwSEAS6_1),.clk(gclk));
	jdff dff_A_uZDh0bOA9_1(.dout(w_dff_A_yIPwSEAS6_1),.din(w_dff_A_uZDh0bOA9_1),.clk(gclk));
	jdff dff_A_s2JklApE7_1(.dout(w_dff_A_uZDh0bOA9_1),.din(w_dff_A_s2JklApE7_1),.clk(gclk));
	jdff dff_A_Vg7e5cJ63_1(.dout(w_dff_A_s2JklApE7_1),.din(w_dff_A_Vg7e5cJ63_1),.clk(gclk));
	jdff dff_A_mn4QwLaf2_1(.dout(w_dff_A_Vg7e5cJ63_1),.din(w_dff_A_mn4QwLaf2_1),.clk(gclk));
	jdff dff_A_yhw6Bu9C1_1(.dout(w_dff_A_mn4QwLaf2_1),.din(w_dff_A_yhw6Bu9C1_1),.clk(gclk));
	jdff dff_A_d0HlFfEt8_1(.dout(w_shift6_0[1]),.din(w_dff_A_d0HlFfEt8_1),.clk(gclk));
	jdff dff_A_0KHUZMz38_1(.dout(w_dff_A_d0HlFfEt8_1),.din(w_dff_A_0KHUZMz38_1),.clk(gclk));
	jdff dff_A_WOA0ZQHw3_1(.dout(w_dff_A_0KHUZMz38_1),.din(w_dff_A_WOA0ZQHw3_1),.clk(gclk));
	jdff dff_A_nn1kfmOP4_1(.dout(w_dff_A_WOA0ZQHw3_1),.din(w_dff_A_nn1kfmOP4_1),.clk(gclk));
	jdff dff_A_wlxdjjOG7_1(.dout(w_dff_A_nn1kfmOP4_1),.din(w_dff_A_wlxdjjOG7_1),.clk(gclk));
	jdff dff_A_hx4tVmIK8_1(.dout(w_dff_A_wlxdjjOG7_1),.din(w_dff_A_hx4tVmIK8_1),.clk(gclk));
	jdff dff_A_UyHOTMnZ3_1(.dout(w_dff_A_hx4tVmIK8_1),.din(w_dff_A_UyHOTMnZ3_1),.clk(gclk));
	jdff dff_A_ITcnN2XY5_1(.dout(w_dff_A_UyHOTMnZ3_1),.din(w_dff_A_ITcnN2XY5_1),.clk(gclk));
	jdff dff_A_VbtfVEBv5_1(.dout(w_dff_A_ITcnN2XY5_1),.din(w_dff_A_VbtfVEBv5_1),.clk(gclk));
	jdff dff_A_dr5pNRNJ3_1(.dout(w_dff_A_VbtfVEBv5_1),.din(w_dff_A_dr5pNRNJ3_1),.clk(gclk));
	jdff dff_A_SBbXK7hb5_1(.dout(w_dff_A_dr5pNRNJ3_1),.din(w_dff_A_SBbXK7hb5_1),.clk(gclk));
	jdff dff_A_GQoVLGyR6_1(.dout(w_dff_A_SBbXK7hb5_1),.din(w_dff_A_GQoVLGyR6_1),.clk(gclk));
	jdff dff_A_khYPEM4x6_1(.dout(w_dff_A_GQoVLGyR6_1),.din(w_dff_A_khYPEM4x6_1),.clk(gclk));
	jdff dff_A_2TQqs4AQ5_2(.dout(w_shift6_0[2]),.din(w_dff_A_2TQqs4AQ5_2),.clk(gclk));
	jdff dff_A_6LJGIMCL8_2(.dout(w_dff_A_2TQqs4AQ5_2),.din(w_dff_A_6LJGIMCL8_2),.clk(gclk));
	jdff dff_A_bI9SQkqI0_2(.dout(w_dff_A_6LJGIMCL8_2),.din(w_dff_A_bI9SQkqI0_2),.clk(gclk));
	jdff dff_A_XbM50qoe5_2(.dout(w_dff_A_bI9SQkqI0_2),.din(w_dff_A_XbM50qoe5_2),.clk(gclk));
	jdff dff_A_OlXmRDr23_2(.dout(w_dff_A_XbM50qoe5_2),.din(w_dff_A_OlXmRDr23_2),.clk(gclk));
	jdff dff_A_tYxLAhIr1_2(.dout(w_dff_A_OlXmRDr23_2),.din(w_dff_A_tYxLAhIr1_2),.clk(gclk));
	jdff dff_A_MxFCGgOe5_2(.dout(w_dff_A_tYxLAhIr1_2),.din(w_dff_A_MxFCGgOe5_2),.clk(gclk));
	jdff dff_A_ujp1IjfH8_2(.dout(w_dff_A_MxFCGgOe5_2),.din(w_dff_A_ujp1IjfH8_2),.clk(gclk));
	jdff dff_A_chwKj2SQ7_2(.dout(w_dff_A_ujp1IjfH8_2),.din(w_dff_A_chwKj2SQ7_2),.clk(gclk));
	jdff dff_A_4gtYzkjf5_2(.dout(w_dff_A_chwKj2SQ7_2),.din(w_dff_A_4gtYzkjf5_2),.clk(gclk));
	jdff dff_A_8Of7GbxQ4_2(.dout(w_dff_A_4gtYzkjf5_2),.din(w_dff_A_8Of7GbxQ4_2),.clk(gclk));
	jdff dff_A_s1NI9TQu9_2(.dout(w_dff_A_8Of7GbxQ4_2),.din(w_dff_A_s1NI9TQu9_2),.clk(gclk));
	jdff dff_A_eLfj31eX1_2(.dout(w_dff_A_s1NI9TQu9_2),.din(w_dff_A_eLfj31eX1_2),.clk(gclk));
endmodule

